// ...
module top(RIb4bfa38_65_b1 ,RIb4bfa38_65_b0 ,RIb4c69c8_39_b1 ,RIb4c69c8_39_b0 ,RIa167a08_1_b1 ,RIa167a08_1_b0 ,RIb4ca3e8_33_b1 ,RIb4ca3e8_33_b0 ,RIa167990_2_b1 ,
		RIa167990_2_b0 ,RIb4c6c20_34_b1 ,RIb4c6c20_34_b0 ,RIa167918_3_b1 ,RIa167918_3_b0 ,RIb4c6ba8_35_b1 ,RIb4c6ba8_35_b0 ,RIa1678a0_4_b1 ,RIa1678a0_4_b0 ,
		RIb4c6b30_36_b1 ,RIb4c6b30_36_b0 ,RIa167828_5_b1 ,RIa167828_5_b0 ,RIb4c6ab8_37_b1 ,RIb4c6ab8_37_b0 ,RIa1677b0_6_b1 ,RIa1677b0_6_b0 ,RIb4c6a40_38_b1 ,
		RIb4c6a40_38_b0 ,RIa167738_7_b1 ,RIa167738_7_b0 ,RIa1676c0_8_b1 ,RIa1676c0_8_b0 ,RIb4c6950_40_b1 ,RIb4c6950_40_b0 ,RIa167648_9_b1 ,RIa167648_9_b0 ,
		RIb4c68d8_41_b1 ,RIb4c68d8_41_b0 ,RIa1675d0_10_b1 ,RIa1675d0_10_b0 ,RIb4c6860_42_b1 ,RIb4c6860_42_b0 ,RIa167558_11_b1 ,RIa167558_11_b0 ,RIb4c67e8_43_b1 ,
		RIb4c67e8_43_b0 ,RIa1674e0_12_b1 ,RIa1674e0_12_b0 ,RIb4c6770_44_b1 ,RIb4c6770_44_b0 ,RIa167468_13_b1 ,RIa167468_13_b0 ,RIb4c3368_45_b1 ,RIb4c3368_45_b0 ,
		RIa1673f0_14_b1 ,RIa1673f0_14_b0 ,RIb4c32f0_46_b1 ,RIb4c32f0_46_b0 ,RIa167378_15_b1 ,RIa167378_15_b0 ,RIb4c3278_47_b1 ,RIb4c3278_47_b0 ,RIa167300_16_b1 ,
		RIa167300_16_b0 ,RIb4c3200_48_b1 ,RIb4c3200_48_b0 ,RIa167288_17_b1 ,RIa167288_17_b0 ,RIb4c3188_49_b1 ,RIb4c3188_49_b0 ,RIa167210_18_b1 ,RIa167210_18_b0 ,
		RIb4c3110_50_b1 ,RIb4c3110_50_b0 ,RIa167198_19_b1 ,RIa167198_19_b0 ,RIb4c3098_51_b1 ,RIb4c3098_51_b0 ,RIa167120_20_b1 ,RIa167120_20_b0 ,RIb4c3020_52_b1 ,
		RIb4c3020_52_b0 ,RIa1670a8_21_b1 ,RIa1670a8_21_b0 ,RIb4c2fa8_53_b1 ,RIb4c2fa8_53_b0 ,RIa167030_22_b1 ,RIa167030_22_b0 ,RIb4c2f30_54_b1 ,RIb4c2f30_54_b0 ,
		RIa166fb8_23_b1 ,RIa166fb8_23_b0 ,RIb4c2eb8_55_b1 ,RIb4c2eb8_55_b0 ,RIa166f40_24_b1 ,RIa166f40_24_b0 ,RIb4c2e40_56_b1 ,RIb4c2e40_56_b0 ,RIa166ec8_25_b1 ,
		RIa166ec8_25_b0 ,RIb4c2dc8_57_b1 ,RIb4c2dc8_57_b0 ,RIa166e50_26_b1 ,RIa166e50_26_b0 ,RIb4c2d50_58_b1 ,RIb4c2d50_58_b0 ,RIa166dd8_27_b1 ,RIa166dd8_27_b0 ,
		RIb4c2cd8_59_b1 ,RIb4c2cd8_59_b0 ,RIa166d60_28_b1 ,RIa166d60_28_b0 ,RIb4c2c60_60_b1 ,RIb4c2c60_60_b0 ,RIa166ce8_29_b1 ,RIa166ce8_29_b0 ,RIb4c2be8_61_b1 ,
		RIb4c2be8_61_b0 ,RIa166c70_30_b1 ,RIa166c70_30_b0 ,RIb4c2b70_62_b1 ,RIb4c2b70_62_b0 ,RIb4ca4d8_31_b1 ,RIb4ca4d8_31_b0 ,RIb4c2af8_63_b1 ,RIb4c2af8_63_b0 ,
		RIb4ca460_32_b1 ,RIb4ca460_32_b0 ,RIb4bfab0_64_b1 ,RIb4bfab0_64_b0 ,RIb4bf948_67_b1 ,RIb4bf948_67_b0 ,RIb4bf9c0_66_b1 ,RIb4bf9c0_66_b0 ,RIb4bf858_69_b1 ,
		RIb4bf858_69_b0 ,RIb4bf8d0_68_b1 ,RIb4bf8d0_68_b0 ,RIb4bf768_71_b1 ,RIb4bf768_71_b0 ,RIb4bf7e0_70_b1 ,RIb4bf7e0_70_b0 ,RIb4bf6f0_72_b1 ,RIb4bf6f0_72_b0 ,
		RIb4bf678_73_b1 ,RIb4bf678_73_b0 ,RIb4bf600_74_b1 ,RIb4bf600_74_b0 ,RIb4bf588_75_b1 ,RIb4bf588_75_b0 ,RIb4bf510_76_b1 ,RIb4bf510_76_b0 ,RIb4bf498_77_b1 ,
		RIb4bf498_77_b0 ,RIb4bf420_78_b1 ,RIb4bf420_78_b0 ,RIb4bf3a8_79_b1 ,RIb4bf3a8_79_b0 ,RIb4bf330_80_b1 ,RIb4bf330_80_b0 ,RIb4bf2b8_81_b1 ,RIb4bf2b8_81_b0 ,
		RIb4bf240_82_b1 ,RIb4bf240_82_b0 ,RIb4bf1c8_83_b1 ,RIb4bf1c8_83_b0 ,RIb4bf150_84_b1 ,RIb4bf150_84_b0 ,RIb4bf0d8_85_b1 ,RIb4bf0d8_85_b0 ,RIb4bf060_86_b1 ,
		RIb4bf060_86_b0 ,RIb4befe8_87_b1 ,RIb4befe8_87_b0 ,RIb4bef70_88_b1 ,RIb4bef70_88_b0 ,RIb4beef8_89_b1 ,RIb4beef8_89_b0 ,RIb4bee80_90_b1 ,RIb4bee80_90_b0 ,
		RIb4bc1f8_91_b1 ,RIb4bc1f8_91_b0 ,RIb4bc180_92_b1 ,RIb4bc180_92_b0 ,RIb4bc108_93_b1 ,RIb4bc108_93_b0 ,RIb4bc090_94_b1 ,RIb4bc090_94_b0 ,RIb4bc018_95_b1 ,
		RIb4bc018_95_b0 ,RIb4bbfa0_96_b1 ,RIb4bbfa0_96_b0 ,R_61_85b54e8_b1 ,R_61_85b54e8_b0 ,R_62_85b5590_b1 ,R_62_85b5590_b0 ,R_63_85b5638_b1 ,R_63_85b5638_b0 ,
		R_64_85b56e0_b1 ,R_64_85b56e0_b0 ,R_65_85b5788_b1 ,R_65_85b5788_b0 ,R_66_85b5830_b1 ,R_66_85b5830_b0 ,R_67_85b58d8_b1 ,R_67_85b58d8_b0 ,R_68_85b5980_b1 ,
		R_68_85b5980_b0 ,R_69_85b5a28_b1 ,R_69_85b5a28_b0 ,R_6a_85b5ad0_b1 ,R_6a_85b5ad0_b0 ,R_6b_85b5b78_b1 ,R_6b_85b5b78_b0 ,R_6c_85b5c20_b1 ,R_6c_85b5c20_b0 ,
		R_6d_85b5cc8_b1 ,R_6d_85b5cc8_b0 ,R_6e_85b5d70_b1 ,R_6e_85b5d70_b0 ,R_6f_85b5e18_b1 ,R_6f_85b5e18_b0 ,R_70_85b5ec0_b1 ,R_70_85b5ec0_b0 ,R_71_85b5f68_b1 ,
		R_71_85b5f68_b0 ,R_72_85b6010_b1 ,R_72_85b6010_b0 ,R_73_85b60b8_b1 ,R_73_85b60b8_b0 ,R_74_85b6160_b1 ,R_74_85b6160_b0 ,R_75_85b6208_b1 ,R_75_85b6208_b0 ,
		R_76_85b62b0_b1 ,R_76_85b62b0_b0 ,R_77_85b6358_b1 ,R_77_85b6358_b0 ,R_78_85b6400_b1 ,R_78_85b6400_b0 ,R_79_85b64a8_b1 ,R_79_85b64a8_b0 ,R_7a_85b6550_b1 ,
		R_7a_85b6550_b0 ,R_7b_85b65f8_b1 ,R_7b_85b65f8_b0 ,R_7c_85b66a0_b1 ,R_7c_85b66a0_b0 ,R_7d_85b6748_b1 ,R_7d_85b6748_b0 ,R_7e_85b67f0_b1 ,R_7e_85b67f0_b0 ,
		R_7f_85b6898_b1 ,R_7f_85b6898_b0 ,R_80_85b6940_b1 ,R_80_85b6940_b0 ,R_81_85b69e8_b1 ,R_81_85b69e8_b0 ,R_82_85b6a90_b1 ,R_82_85b6a90_b0 ,R_83_85b6b38_b1 ,
		R_83_85b6b38_b0 ,R_84_85b6be0_b1 ,R_84_85b6be0_b0 ,R_85_85b6c88_b1 ,R_85_85b6c88_b0 ,R_86_85b6d30_b1 ,R_86_85b6d30_b0 ,R_87_85b6dd8_b1 ,R_87_85b6dd8_b0 ,
		R_88_85b6e80_b1 ,R_88_85b6e80_b0 ,R_89_85b6f28_b1 ,R_89_85b6f28_b0 ,R_8a_85b6fd0_b1 ,R_8a_85b6fd0_b0 ,R_8b_85b7078_b1 ,R_8b_85b7078_b0 ,R_8c_85b7120_b1 ,
		R_8c_85b7120_b0 ,R_8d_85b71c8_b1 ,R_8d_85b71c8_b0 ,R_8e_85b7270_b1 ,R_8e_85b7270_b0 ,R_8f_85b7318_b1 ,R_8f_85b7318_b0 ,R_90_85b73c0_b1 ,R_90_85b73c0_b0 ,
		R_91_85b7468_b1 ,R_91_85b7468_b0 ,R_92_85b7510_b1 ,R_92_85b7510_b0 ,R_93_85b75b8_b1 ,R_93_85b75b8_b0 ,R_94_85b7660_b1 ,R_94_85b7660_b0 ,R_95_85b7708_b1 ,
		R_95_85b7708_b0 ,R_96_85b77b0_b1 ,R_96_85b77b0_b0 ,R_97_85b7858_b1 ,R_97_85b7858_b0 ,R_98_85b7900_b1 ,R_98_85b7900_b0 ,R_99_85b79a8_b1 ,R_99_85b79a8_b0 ,
		R_9a_85b7a50_b1 ,R_9a_85b7a50_b0 );
input RIb4bfa38_65_b1 ,RIb4bfa38_65_b0 ,RIb4c69c8_39_b1 ,RIb4c69c8_39_b0 ,RIa167a08_1_b1 ,RIa167a08_1_b0 ,RIb4ca3e8_33_b1 ,RIb4ca3e8_33_b0 ,RIa167990_2_b1 ,
		RIa167990_2_b0 ,RIb4c6c20_34_b1 ,RIb4c6c20_34_b0 ,RIa167918_3_b1 ,RIa167918_3_b0 ,RIb4c6ba8_35_b1 ,RIb4c6ba8_35_b0 ,RIa1678a0_4_b1 ,RIa1678a0_4_b0 ,
		RIb4c6b30_36_b1 ,RIb4c6b30_36_b0 ,RIa167828_5_b1 ,RIa167828_5_b0 ,RIb4c6ab8_37_b1 ,RIb4c6ab8_37_b0 ,RIa1677b0_6_b1 ,RIa1677b0_6_b0 ,RIb4c6a40_38_b1 ,
		RIb4c6a40_38_b0 ,RIa167738_7_b1 ,RIa167738_7_b0 ,RIa1676c0_8_b1 ,RIa1676c0_8_b0 ,RIb4c6950_40_b1 ,RIb4c6950_40_b0 ,RIa167648_9_b1 ,RIa167648_9_b0 ,
		RIb4c68d8_41_b1 ,RIb4c68d8_41_b0 ,RIa1675d0_10_b1 ,RIa1675d0_10_b0 ,RIb4c6860_42_b1 ,RIb4c6860_42_b0 ,RIa167558_11_b1 ,RIa167558_11_b0 ,RIb4c67e8_43_b1 ,
		RIb4c67e8_43_b0 ,RIa1674e0_12_b1 ,RIa1674e0_12_b0 ,RIb4c6770_44_b1 ,RIb4c6770_44_b0 ,RIa167468_13_b1 ,RIa167468_13_b0 ,RIb4c3368_45_b1 ,RIb4c3368_45_b0 ,
		RIa1673f0_14_b1 ,RIa1673f0_14_b0 ,RIb4c32f0_46_b1 ,RIb4c32f0_46_b0 ,RIa167378_15_b1 ,RIa167378_15_b0 ,RIb4c3278_47_b1 ,RIb4c3278_47_b0 ,RIa167300_16_b1 ,
		RIa167300_16_b0 ,RIb4c3200_48_b1 ,RIb4c3200_48_b0 ,RIa167288_17_b1 ,RIa167288_17_b0 ,RIb4c3188_49_b1 ,RIb4c3188_49_b0 ,RIa167210_18_b1 ,RIa167210_18_b0 ,
		RIb4c3110_50_b1 ,RIb4c3110_50_b0 ,RIa167198_19_b1 ,RIa167198_19_b0 ,RIb4c3098_51_b1 ,RIb4c3098_51_b0 ,RIa167120_20_b1 ,RIa167120_20_b0 ,RIb4c3020_52_b1 ,
		RIb4c3020_52_b0 ,RIa1670a8_21_b1 ,RIa1670a8_21_b0 ,RIb4c2fa8_53_b1 ,RIb4c2fa8_53_b0 ,RIa167030_22_b1 ,RIa167030_22_b0 ,RIb4c2f30_54_b1 ,RIb4c2f30_54_b0 ,
		RIa166fb8_23_b1 ,RIa166fb8_23_b0 ,RIb4c2eb8_55_b1 ,RIb4c2eb8_55_b0 ,RIa166f40_24_b1 ,RIa166f40_24_b0 ,RIb4c2e40_56_b1 ,RIb4c2e40_56_b0 ,RIa166ec8_25_b1 ,
		RIa166ec8_25_b0 ,RIb4c2dc8_57_b1 ,RIb4c2dc8_57_b0 ,RIa166e50_26_b1 ,RIa166e50_26_b0 ,RIb4c2d50_58_b1 ,RIb4c2d50_58_b0 ,RIa166dd8_27_b1 ,RIa166dd8_27_b0 ,
		RIb4c2cd8_59_b1 ,RIb4c2cd8_59_b0 ,RIa166d60_28_b1 ,RIa166d60_28_b0 ,RIb4c2c60_60_b1 ,RIb4c2c60_60_b0 ,RIa166ce8_29_b1 ,RIa166ce8_29_b0 ,RIb4c2be8_61_b1 ,
		RIb4c2be8_61_b0 ,RIa166c70_30_b1 ,RIa166c70_30_b0 ,RIb4c2b70_62_b1 ,RIb4c2b70_62_b0 ,RIb4ca4d8_31_b1 ,RIb4ca4d8_31_b0 ,RIb4c2af8_63_b1 ,RIb4c2af8_63_b0 ,
		RIb4ca460_32_b1 ,RIb4ca460_32_b0 ,RIb4bfab0_64_b1 ,RIb4bfab0_64_b0 ,RIb4bf948_67_b1 ,RIb4bf948_67_b0 ,RIb4bf9c0_66_b1 ,RIb4bf9c0_66_b0 ,RIb4bf858_69_b1 ,
		RIb4bf858_69_b0 ,RIb4bf8d0_68_b1 ,RIb4bf8d0_68_b0 ,RIb4bf768_71_b1 ,RIb4bf768_71_b0 ,RIb4bf7e0_70_b1 ,RIb4bf7e0_70_b0 ,RIb4bf6f0_72_b1 ,RIb4bf6f0_72_b0 ,
		RIb4bf678_73_b1 ,RIb4bf678_73_b0 ,RIb4bf600_74_b1 ,RIb4bf600_74_b0 ,RIb4bf588_75_b1 ,RIb4bf588_75_b0 ,RIb4bf510_76_b1 ,RIb4bf510_76_b0 ,RIb4bf498_77_b1 ,
		RIb4bf498_77_b0 ,RIb4bf420_78_b1 ,RIb4bf420_78_b0 ,RIb4bf3a8_79_b1 ,RIb4bf3a8_79_b0 ,RIb4bf330_80_b1 ,RIb4bf330_80_b0 ,RIb4bf2b8_81_b1 ,RIb4bf2b8_81_b0 ,
		RIb4bf240_82_b1 ,RIb4bf240_82_b0 ,RIb4bf1c8_83_b1 ,RIb4bf1c8_83_b0 ,RIb4bf150_84_b1 ,RIb4bf150_84_b0 ,RIb4bf0d8_85_b1 ,RIb4bf0d8_85_b0 ,RIb4bf060_86_b1 ,
		RIb4bf060_86_b0 ,RIb4befe8_87_b1 ,RIb4befe8_87_b0 ,RIb4bef70_88_b1 ,RIb4bef70_88_b0 ,RIb4beef8_89_b1 ,RIb4beef8_89_b0 ,RIb4bee80_90_b1 ,RIb4bee80_90_b0 ,
		RIb4bc1f8_91_b1 ,RIb4bc1f8_91_b0 ,RIb4bc180_92_b1 ,RIb4bc180_92_b0 ,RIb4bc108_93_b1 ,RIb4bc108_93_b0 ,RIb4bc090_94_b1 ,RIb4bc090_94_b0 ,RIb4bc018_95_b1 ,
		RIb4bc018_95_b0 ,RIb4bbfa0_96_b1 ,RIb4bbfa0_96_b0 ;
output R_61_85b54e8_b1 ,R_61_85b54e8_b0 ,R_62_85b5590_b1 ,R_62_85b5590_b0 ,R_63_85b5638_b1 ,R_63_85b5638_b0 ,R_64_85b56e0_b1 ,R_64_85b56e0_b0 ,R_65_85b5788_b1 ,
		R_65_85b5788_b0 ,R_66_85b5830_b1 ,R_66_85b5830_b0 ,R_67_85b58d8_b1 ,R_67_85b58d8_b0 ,R_68_85b5980_b1 ,R_68_85b5980_b0 ,R_69_85b5a28_b1 ,R_69_85b5a28_b0 ,
		R_6a_85b5ad0_b1 ,R_6a_85b5ad0_b0 ,R_6b_85b5b78_b1 ,R_6b_85b5b78_b0 ,R_6c_85b5c20_b1 ,R_6c_85b5c20_b0 ,R_6d_85b5cc8_b1 ,R_6d_85b5cc8_b0 ,R_6e_85b5d70_b1 ,
		R_6e_85b5d70_b0 ,R_6f_85b5e18_b1 ,R_6f_85b5e18_b0 ,R_70_85b5ec0_b1 ,R_70_85b5ec0_b0 ,R_71_85b5f68_b1 ,R_71_85b5f68_b0 ,R_72_85b6010_b1 ,R_72_85b6010_b0 ,
		R_73_85b60b8_b1 ,R_73_85b60b8_b0 ,R_74_85b6160_b1 ,R_74_85b6160_b0 ,R_75_85b6208_b1 ,R_75_85b6208_b0 ,R_76_85b62b0_b1 ,R_76_85b62b0_b0 ,R_77_85b6358_b1 ,
		R_77_85b6358_b0 ,R_78_85b6400_b1 ,R_78_85b6400_b0 ,R_79_85b64a8_b1 ,R_79_85b64a8_b0 ,R_7a_85b6550_b1 ,R_7a_85b6550_b0 ,R_7b_85b65f8_b1 ,R_7b_85b65f8_b0 ,
		R_7c_85b66a0_b1 ,R_7c_85b66a0_b0 ,R_7d_85b6748_b1 ,R_7d_85b6748_b0 ,R_7e_85b67f0_b1 ,R_7e_85b67f0_b0 ,R_7f_85b6898_b1 ,R_7f_85b6898_b0 ,R_80_85b6940_b1 ,
		R_80_85b6940_b0 ,R_81_85b69e8_b1 ,R_81_85b69e8_b0 ,R_82_85b6a90_b1 ,R_82_85b6a90_b0 ,R_83_85b6b38_b1 ,R_83_85b6b38_b0 ,R_84_85b6be0_b1 ,R_84_85b6be0_b0 ,
		R_85_85b6c88_b1 ,R_85_85b6c88_b0 ,R_86_85b6d30_b1 ,R_86_85b6d30_b0 ,R_87_85b6dd8_b1 ,R_87_85b6dd8_b0 ,R_88_85b6e80_b1 ,R_88_85b6e80_b0 ,R_89_85b6f28_b1 ,
		R_89_85b6f28_b0 ,R_8a_85b6fd0_b1 ,R_8a_85b6fd0_b0 ,R_8b_85b7078_b1 ,R_8b_85b7078_b0 ,R_8c_85b7120_b1 ,R_8c_85b7120_b0 ,R_8d_85b71c8_b1 ,R_8d_85b71c8_b0 ,
		R_8e_85b7270_b1 ,R_8e_85b7270_b0 ,R_8f_85b7318_b1 ,R_8f_85b7318_b0 ,R_90_85b73c0_b1 ,R_90_85b73c0_b0 ,R_91_85b7468_b1 ,R_91_85b7468_b0 ,R_92_85b7510_b1 ,
		R_92_85b7510_b0 ,R_93_85b75b8_b1 ,R_93_85b75b8_b0 ,R_94_85b7660_b1 ,R_94_85b7660_b0 ,R_95_85b7708_b1 ,R_95_85b7708_b0 ,R_96_85b77b0_b1 ,R_96_85b77b0_b0 ,
		R_97_85b7858_b1 ,R_97_85b7858_b0 ,R_98_85b7900_b1 ,R_98_85b7900_b0 ,R_99_85b79a8_b1 ,R_99_85b79a8_b0 ,R_9a_85b7a50_b1 ,R_9a_85b7a50_b0 ;

wire \155_b1 , \155_b0 , \156_N$1_b1 , \156_N$1_b0 , \157_ZERO_b1 , \157_ZERO_b0 , \158_ONE_b1 , \158_ONE_b0 , \159_b1 , \159_b0 , 
		\160_b1 , \160_b0 , \161_b1 , \161_b0 , \162_b1 , \162_b0 , \163_b1 , \163_b0 , \164_b1 , \164_b0 , 
		\165_b1 , \165_b0 , \166_b1 , \166_b0 , \167_b1 , \167_b0 , \168_b1 , \168_b0 , \169_b1 , \169_b0 , 
		\170_b1 , \170_b0 , \171_b1 , \171_b0 , \172_b1 , \172_b0 , \173_b1 , \173_b0 , \174_b1 , \174_b0 , 
		\175_b1 , \175_b0 , \176_b1 , \176_b0 , \177_b1 , \177_b0 , \178_b1 , \178_b0 , \179_b1 , \179_b0 , 
		\180_b1 , \180_b0 , \181_b1 , \181_b0 , \182_b1 , \182_b0 , \183_b1 , \183_b0 , \184_b1 , \184_b0 , 
		\185_b1 , \185_b0 , \186_b1 , \186_b0 , \187_b1 , \187_b0 , \188_b1 , \188_b0 , \189_b1 , \189_b0 , 
		\190_b1 , \190_b0 , \191_b1 , \191_b0 , \192_b1 , \192_b0 , \193_b1 , \193_b0 , \194_b1 , \194_b0 , 
		\195_b1 , \195_b0 , \196_b1 , \196_b0 , \197_b1 , \197_b0 , \198_b1 , \198_b0 , \199_b1 , \199_b0 , 
		\200_b1 , \200_b0 , \201_b1 , \201_b0 , \202_b1 , \202_b0 , \203_b1 , \203_b0 , \204_b1 , \204_b0 , 
		\205_b1 , \205_b0 , \206_b1 , \206_b0 , \207_b1 , \207_b0 , \208_b1 , \208_b0 , \209_b1 , \209_b0 , 
		\210_b1 , \210_b0 , \211_b1 , \211_b0 , \212_b1 , \212_b0 , \213_b1 , \213_b0 , \214_b1 , \214_b0 , 
		\215_b1 , \215_b0 , \216_b1 , \216_b0 , \217_b1 , \217_b0 , \218_b1 , \218_b0 , \219_b1 , \219_b0 , 
		\220_b1 , \220_b0 , \221_b1 , \221_b0 , \222_b1 , \222_b0 , \223_b1 , \223_b0 , \224_b1 , \224_b0 , 
		\225_b1 , \225_b0 , \226_b1 , \226_b0 , \227_b1 , \227_b0 , \228_b1 , \228_b0 , \229_b1 , \229_b0 , 
		\230_b1 , \230_b0 , \231_b1 , \231_b0 , \232_b1 , \232_b0 , \233_b1 , \233_b0 , \234_b1 , \234_b0 , 
		\235_b1 , \235_b0 , \236_b1 , \236_b0 , \237_b1 , \237_b0 , \238_b1 , \238_b0 , \239_b1 , \239_b0 , 
		\240_b1 , \240_b0 , \241_b1 , \241_b0 , \242_b1 , \242_b0 , \243_b1 , \243_b0 , \244_b1 , \244_b0 , 
		\245_b1 , \245_b0 , \246_b1 , \246_b0 , \247_b1 , \247_b0 , \248_b1 , \248_b0 , \249_b1 , \249_b0 , 
		\250_b1 , \250_b0 , \251_b1 , \251_b0 , \252_b1 , \252_b0 , \253_b1 , \253_b0 , \254_b1 , \254_b0 , 
		\255_b1 , \255_b0 , \256_b1 , \256_b0 , \257_b1 , \257_b0 , \258_b1 , \258_b0 , \259_b1 , \259_b0 , 
		\260_b1 , \260_b0 , \261_b1 , \261_b0 , \262_b1 , \262_b0 , \263_b1 , \263_b0 , \264_b1 , \264_b0 , 
		\265_b1 , \265_b0 , \266_b1 , \266_b0 , \267_b1 , \267_b0 , \268_b1 , \268_b0 , \269_b1 , \269_b0 , 
		\270_b1 , \270_b0 , \271_b1 , \271_b0 , \272_b1 , \272_b0 , \273_b1 , \273_b0 , \274_b1 , \274_b0 , 
		\275_b1 , \275_b0 , \276_b1 , \276_b0 , \277_b1 , \277_b0 , \278_b1 , \278_b0 , \279_b1 , \279_b0 , 
		\280_b1 , \280_b0 , \281_b1 , \281_b0 , \282_b1 , \282_b0 , \283_b1 , \283_b0 , \284_b1 , \284_b0 , 
		\285_b1 , \285_b0 , \286_b1 , \286_b0 , \287_b1 , \287_b0 , \288_b1 , \288_b0 , \289_nR13d_b1 , \289_nR13d_b0 , 
		\290_b1 , \290_b0 , \291_nR13c_b1 , \291_nR13c_b0 , \292_b1 , \292_b0 , \293_b1 , \293_b0 , \294_nR13b_b1 , \294_nR13b_b0 , 
		\295_b1 , \295_b0 , \296_b1 , \296_b0 , \297_b1 , \297_b0 , \298_b1 , \298_b0 , \299_b1 , \299_b0 , 
		\300_b1 , \300_b0 , \301_b1 , \301_b0 , \302_b1 , \302_b0 , \303_b1 , \303_b0 , \304_b1 , \304_b0 , 
		\305_b1 , \305_b0 , \306_nR13f_b1 , \306_nR13f_b0 , \307_b1 , \307_b0 , \308_nR13e_b1 , \308_nR13e_b0 , \309_b1 , \309_b0 , 
		\310_b1 , \310_b0 , \311_b1 , \311_b0 , \312_b1 , \312_b0 , \313_b1 , \313_b0 , \314_b1 , \314_b0 , 
		\315_b1 , \315_b0 , \316_b1 , \316_b0 , \317_b1 , \317_b0 , \318_b1 , \318_b0 , \319_b1 , \319_b0 , 
		\320_b1 , \320_b0 , \321_b1 , \321_b0 , \322_b1 , \322_b0 , \323_b1 , \323_b0 , \324_nR141_b1 , \324_nR141_b0 , 
		\325_b1 , \325_b0 , \326_nR140_b1 , \326_nR140_b0 , \327_b1 , \327_b0 , \328_b1 , \328_b0 , \329_b1 , \329_b0 , 
		\330_b1 , \330_b0 , \331_b1 , \331_b0 , \332_b1 , \332_b0 , \333_b1 , \333_b0 , \334_b1 , \334_b0 , 
		\335_b1 , \335_b0 , \336_b1 , \336_b0 , \337_b1 , \337_b0 , \338_b1 , \338_b0 , \339_b1 , \339_b0 , 
		\340_b1 , \340_b0 , \341_b1 , \341_b0 , \342_b1 , \342_b0 , \343_b1 , \343_b0 , \344_nR143_b1 , \344_nR143_b0 , 
		\345_b1 , \345_b0 , \346_nR142_b1 , \346_nR142_b0 , \347_b1 , \347_b0 , \348_b1 , \348_b0 , \349_b1 , \349_b0 , 
		\350_b1 , \350_b0 , \351_b1 , \351_b0 , \352_b1 , \352_b0 , \353_b1 , \353_b0 , \354_b1 , \354_b0 , 
		\355_b1 , \355_b0 , \356_b1 , \356_b0 , \357_b1 , \357_b0 , \358_b1 , \358_b0 , \359_b1 , \359_b0 , 
		\360_b1 , \360_b0 , \361_b1 , \361_b0 , \362_b1 , \362_b0 , \363_b1 , \363_b0 , \364_b1 , \364_b0 , 
		\365_b1 , \365_b0 , \366_b1 , \366_b0 , \367_b1 , \367_b0 , \368_b1 , \368_b0 , \369_b1 , \369_b0 , 
		\370_b1 , \370_b0 , \371_b1 , \371_b0 , \372_b1 , \372_b0 , \373_b1 , \373_b0 , \374_b1 , \374_b0 , 
		\375_b1 , \375_b0 , \376_b1 , \376_b0 , \377_b1 , \377_b0 , \378_b1 , \378_b0 , \379_b1 , \379_b0 , 
		\380_b1 , \380_b0 , \381_b1 , \381_b0 , \382_b1 , \382_b0 , \383_b1 , \383_b0 , \384_b1 , \384_b0 , 
		\385_b1 , \385_b0 , \386_b1 , \386_b0 , \387_b1 , \387_b0 , \388_b1 , \388_b0 , \389_b1 , \389_b0 , 
		\390_b1 , \390_b0 , \391_b1 , \391_b0 , \392_b1 , \392_b0 , \393_b1 , \393_b0 , \394_b1 , \394_b0 , 
		\395_b1 , \395_b0 , \396_b1 , \396_b0 , \397_b1 , \397_b0 , \398_b1 , \398_b0 , \399_b1 , \399_b0 , 
		\400_b1 , \400_b0 , \401_b1 , \401_b0 , \402_b1 , \402_b0 , \403_b1 , \403_b0 , \404_b1 , \404_b0 , 
		\405_b1 , \405_b0 , \406_b1 , \406_b0 , \407_b1 , \407_b0 , \408_b1 , \408_b0 , \409_b1 , \409_b0 , 
		\410_b1 , \410_b0 , \411_b1 , \411_b0 , \412_b1 , \412_b0 , \413_b1 , \413_b0 , \414_b1 , \414_b0 , 
		\415_b1 , \415_b0 , \416_b1 , \416_b0 , \417_b1 , \417_b0 , \418_b1 , \418_b0 , \419_b1 , \419_b0 , 
		\420_b1 , \420_b0 , \421_b1 , \421_b0 , \422_b1 , \422_b0 , \423_b1 , \423_b0 , \424_b1 , \424_b0 , 
		\425_b1 , \425_b0 , \426_b1 , \426_b0 , \427_b1 , \427_b0 , \428_b1 , \428_b0 , \429_b1 , \429_b0 , 
		\430_b1 , \430_b0 , \431_b1 , \431_b0 , \432_b1 , \432_b0 , \433_b1 , \433_b0 , \434_b1 , \434_b0 , 
		\435_b1 , \435_b0 , \436_b1 , \436_b0 , \437_b1 , \437_b0 , \438_b1 , \438_b0 , \439_b1 , \439_b0 , 
		\440_b1 , \440_b0 , \441_b1 , \441_b0 , \442_b1 , \442_b0 , \443_b1 , \443_b0 , \444_b1 , \444_b0 , 
		\445_b1 , \445_b0 , \446_b1 , \446_b0 , \447_b1 , \447_b0 , \448_b1 , \448_b0 , \449_nR13a_b1 , \449_nR13a_b0 , 
		\450_b1 , \450_b0 , \451_nR139_b1 , \451_nR139_b0 , \452_b1 , \452_b0 , \453_b1 , \453_b0 , \454_b1 , \454_b0 , 
		\455_b1 , \455_b0 , \456_b1 , \456_b0 , \457_b1 , \457_b0 , \458_b1 , \458_b0 , \459_b1 , \459_b0 , 
		\460_b1 , \460_b0 , \461_b1 , \461_b0 , \462_b1 , \462_b0 , \463_b1 , \463_b0 , \464_b1 , \464_b0 , 
		\465_b1 , \465_b0 , \466_b1 , \466_b0 , \467_b1 , \467_b0 , \468_b1 , \468_b0 , \469_b1 , \469_b0 , 
		\470_b1 , \470_b0 , \471_b1 , \471_b0 , \472_b1 , \472_b0 , \473_b1 , \473_b0 , \474_b1 , \474_b0 , 
		\475_b1 , \475_b0 , \476_b1 , \476_b0 , \477_b1 , \477_b0 , \478_b1 , \478_b0 , \479_b1 , \479_b0 , 
		\480_b1 , \480_b0 , \481_b1 , \481_b0 , \482_b1 , \482_b0 , \483_b1 , \483_b0 , \484_b1 , \484_b0 , 
		\485_b1 , \485_b0 , \486_b1 , \486_b0 , \487_b1 , \487_b0 , \488_b1 , \488_b0 , \489_b1 , \489_b0 , 
		\490_b1 , \490_b0 , \491_b1 , \491_b0 , \492_b1 , \492_b0 , \493_b1 , \493_b0 , \494_b1 , \494_b0 , 
		\495_b1 , \495_b0 , \496_b1 , \496_b0 , \497_b1 , \497_b0 , \498_b1 , \498_b0 , \499_b1 , \499_b0 , 
		\500_b1 , \500_b0 , \501_b1 , \501_b0 , \502_b1 , \502_b0 , \503_b1 , \503_b0 , \504_b1 , \504_b0 , 
		\505_b1 , \505_b0 , \506_b1 , \506_b0 , \507_b1 , \507_b0 , \508_b1 , \508_b0 , \509_b1 , \509_b0 , 
		\510_b1 , \510_b0 , \511_b1 , \511_b0 , \512_b1 , \512_b0 , \513_b1 , \513_b0 , \514_b1 , \514_b0 , 
		\515_b1 , \515_b0 , \516_b1 , \516_b0 , \517_b1 , \517_b0 , \518_b1 , \518_b0 , \519_b1 , \519_b0 , 
		\520_b1 , \520_b0 , \521_b1 , \521_b0 , \522_b1 , \522_b0 , \523_b1 , \523_b0 , \524_b1 , \524_b0 , 
		\525_b1 , \525_b0 , \526_b1 , \526_b0 , \527_b1 , \527_b0 , \528_b1 , \528_b0 , \529_b1 , \529_b0 , 
		\530_b1 , \530_b0 , \531_b1 , \531_b0 , \532_b1 , \532_b0 , \533_b1 , \533_b0 , \534_b1 , \534_b0 , 
		\535_b1 , \535_b0 , \536_b1 , \536_b0 , \537_b1 , \537_b0 , \538_b1 , \538_b0 , \539_b1 , \539_b0 , 
		\540_b1 , \540_b0 , \541_b1 , \541_b0 , \542_b1 , \542_b0 , \543_b1 , \543_b0 , \544_b1 , \544_b0 , 
		\545_b1 , \545_b0 , \546_b1 , \546_b0 , \547_b1 , \547_b0 , \548_b1 , \548_b0 , \549_b1 , \549_b0 , 
		\550_b1 , \550_b0 , \551_b1 , \551_b0 , \552_b1 , \552_b0 , \553_b1 , \553_b0 , \554_b1 , \554_b0 , 
		\555_nR138_b1 , \555_nR138_b0 , \556_b1 , \556_b0 , \557_nR137_b1 , \557_nR137_b0 , \558_b1 , \558_b0 , \559_b1 , \559_b0 , 
		\560_b1 , \560_b0 , \561_b1 , \561_b0 , \562_b1 , \562_b0 , \563_b1 , \563_b0 , \564_b1 , \564_b0 , 
		\565_b1 , \565_b0 , \566_b1 , \566_b0 , \567_b1 , \567_b0 , \568_b1 , \568_b0 , \569_b1 , \569_b0 , 
		\570_b1 , \570_b0 , \571_b1 , \571_b0 , \572_b1 , \572_b0 , \573_b1 , \573_b0 , \574_b1 , \574_b0 , 
		\575_b1 , \575_b0 , \576_b1 , \576_b0 , \577_b1 , \577_b0 , \578_b1 , \578_b0 , \579_b1 , \579_b0 , 
		\580_b1 , \580_b0 , \581_b1 , \581_b0 , \582_b1 , \582_b0 , \583_b1 , \583_b0 , \584_b1 , \584_b0 , 
		\585_b1 , \585_b0 , \586_b1 , \586_b0 , \587_b1 , \587_b0 , \588_b1 , \588_b0 , \589_b1 , \589_b0 , 
		\590_b1 , \590_b0 , \591_b1 , \591_b0 , \592_b1 , \592_b0 , \593_b1 , \593_b0 , \594_b1 , \594_b0 , 
		\595_b1 , \595_b0 , \596_b1 , \596_b0 , \597_b1 , \597_b0 , \598_b1 , \598_b0 , \599_b1 , \599_b0 , 
		\600_b1 , \600_b0 , \601_b1 , \601_b0 , \602_b1 , \602_b0 , \603_b1 , \603_b0 , \604_b1 , \604_b0 , 
		\605_b1 , \605_b0 , \606_b1 , \606_b0 , \607_b1 , \607_b0 , \608_b1 , \608_b0 , \609_b1 , \609_b0 , 
		\610_b1 , \610_b0 , \611_b1 , \611_b0 , \612_b1 , \612_b0 , \613_b1 , \613_b0 , \614_b1 , \614_b0 , 
		\615_b1 , \615_b0 , \616_b1 , \616_b0 , \617_b1 , \617_b0 , \618_b1 , \618_b0 , \619_b1 , \619_b0 , 
		\620_b1 , \620_b0 , \621_b1 , \621_b0 , \622_b1 , \622_b0 , \623_b1 , \623_b0 , \624_b1 , \624_b0 , 
		\625_b1 , \625_b0 , \626_b1 , \626_b0 , \627_b1 , \627_b0 , \628_b1 , \628_b0 , \629_b1 , \629_b0 , 
		\630_b1 , \630_b0 , \631_b1 , \631_b0 , \632_b1 , \632_b0 , \633_b1 , \633_b0 , \634_b1 , \634_b0 , 
		\635_b1 , \635_b0 , \636_b1 , \636_b0 , \637_b1 , \637_b0 , \638_b1 , \638_b0 , \639_b1 , \639_b0 , 
		\640_b1 , \640_b0 , \641_b1 , \641_b0 , \642_b1 , \642_b0 , \643_b1 , \643_b0 , \644_b1 , \644_b0 , 
		\645_b1 , \645_b0 , \646_b1 , \646_b0 , \647_b1 , \647_b0 , \648_b1 , \648_b0 , \649_b1 , \649_b0 , 
		\650_b1 , \650_b0 , \651_b1 , \651_b0 , \652_b1 , \652_b0 , \653_b1 , \653_b0 , \654_b1 , \654_b0 , 
		\655_b1 , \655_b0 , \656_b1 , \656_b0 , \657_b1 , \657_b0 , \658_b1 , \658_b0 , \659_b1 , \659_b0 , 
		\660_b1 , \660_b0 , \661_b1 , \661_b0 , \662_nR136_b1 , \662_nR136_b0 , \663_b1 , \663_b0 , \664_nR135_b1 , \664_nR135_b0 , 
		\665_b1 , \665_b0 , \666_b1 , \666_b0 , \667_b1 , \667_b0 , \668_b1 , \668_b0 , \669_b1 , \669_b0 , 
		\670_b1 , \670_b0 , \671_b1 , \671_b0 , \672_b1 , \672_b0 , \673_b1 , \673_b0 , \674_b1 , \674_b0 , 
		\675_b1 , \675_b0 , \676_b1 , \676_b0 , \677_b1 , \677_b0 , \678_b1 , \678_b0 , \679_b1 , \679_b0 , 
		\680_b1 , \680_b0 , \681_b1 , \681_b0 , \682_b1 , \682_b0 , \683_b1 , \683_b0 , \684_b1 , \684_b0 , 
		\685_b1 , \685_b0 , \686_b1 , \686_b0 , \687_b1 , \687_b0 , \688_b1 , \688_b0 , \689_b1 , \689_b0 , 
		\690_b1 , \690_b0 , \691_b1 , \691_b0 , \692_b1 , \692_b0 , \693_b1 , \693_b0 , \694_b1 , \694_b0 , 
		\695_b1 , \695_b0 , \696_b1 , \696_b0 , \697_b1 , \697_b0 , \698_b1 , \698_b0 , \699_b1 , \699_b0 , 
		\700_b1 , \700_b0 , \701_b1 , \701_b0 , \702_b1 , \702_b0 , \703_b1 , \703_b0 , \704_b1 , \704_b0 , 
		\705_b1 , \705_b0 , \706_b1 , \706_b0 , \707_b1 , \707_b0 , \708_b1 , \708_b0 , \709_b1 , \709_b0 , 
		\710_b1 , \710_b0 , \711_b1 , \711_b0 , \712_b1 , \712_b0 , \713_b1 , \713_b0 , \714_b1 , \714_b0 , 
		\715_b1 , \715_b0 , \716_b1 , \716_b0 , \717_b1 , \717_b0 , \718_b1 , \718_b0 , \719_b1 , \719_b0 , 
		\720_b1 , \720_b0 , \721_b1 , \721_b0 , \722_b1 , \722_b0 , \723_b1 , \723_b0 , \724_b1 , \724_b0 , 
		\725_b1 , \725_b0 , \726_b1 , \726_b0 , \727_b1 , \727_b0 , \728_b1 , \728_b0 , \729_b1 , \729_b0 , 
		\730_b1 , \730_b0 , \731_b1 , \731_b0 , \732_b1 , \732_b0 , \733_b1 , \733_b0 , \734_b1 , \734_b0 , 
		\735_b1 , \735_b0 , \736_b1 , \736_b0 , \737_b1 , \737_b0 , \738_b1 , \738_b0 , \739_b1 , \739_b0 , 
		\740_b1 , \740_b0 , \741_b1 , \741_b0 , \742_b1 , \742_b0 , \743_b1 , \743_b0 , \744_b1 , \744_b0 , 
		\745_b1 , \745_b0 , \746_b1 , \746_b0 , \747_b1 , \747_b0 , \748_b1 , \748_b0 , \749_b1 , \749_b0 , 
		\750_b1 , \750_b0 , \751_b1 , \751_b0 , \752_b1 , \752_b0 , \753_b1 , \753_b0 , \754_b1 , \754_b0 , 
		\755_b1 , \755_b0 , \756_b1 , \756_b0 , \757_b1 , \757_b0 , \758_b1 , \758_b0 , \759_b1 , \759_b0 , 
		\760_b1 , \760_b0 , \761_b1 , \761_b0 , \762_b1 , \762_b0 , \763_b1 , \763_b0 , \764_b1 , \764_b0 , 
		\765_b1 , \765_b0 , \766_b1 , \766_b0 , \767_b1 , \767_b0 , \768_b1 , \768_b0 , \769_b1 , \769_b0 , 
		\770_b1 , \770_b0 , \771_b1 , \771_b0 , \772_b1 , \772_b0 , \773_b1 , \773_b0 , \774_b1 , \774_b0 , 
		\775_b1 , \775_b0 , \776_b1 , \776_b0 , \777_b1 , \777_b0 , \778_b1 , \778_b0 , \779_b1 , \779_b0 , 
		\780_b1 , \780_b0 , \781_b1 , \781_b0 , \782_b1 , \782_b0 , \783_b1 , \783_b0 , \784_b1 , \784_b0 , 
		\785_b1 , \785_b0 , \786_b1 , \786_b0 , \787_b1 , \787_b0 , \788_b1 , \788_b0 , \789_b1 , \789_b0 , 
		\790_b1 , \790_b0 , \791_b1 , \791_b0 , \792_b1 , \792_b0 , \793_b1 , \793_b0 , \794_b1 , \794_b0 , 
		\795_b1 , \795_b0 , \796_b1 , \796_b0 , \797_b1 , \797_b0 , \798_b1 , \798_b0 , \799_b1 , \799_b0 , 
		\800_b1 , \800_b0 , \801_b1 , \801_b0 , \802_b1 , \802_b0 , \803_b1 , \803_b0 , \804_b1 , \804_b0 , 
		\805_b1 , \805_b0 , \806_b1 , \806_b0 , \807_b1 , \807_b0 , \808_b1 , \808_b0 , \809_b1 , \809_b0 , 
		\810_b1 , \810_b0 , \811_b1 , \811_b0 , \812_nR134_b1 , \812_nR134_b0 , \813_b1 , \813_b0 , \814_nR133_b1 , \814_nR133_b0 , 
		\815_b1 , \815_b0 , \816_b1 , \816_b0 , \817_b1 , \817_b0 , \818_b1 , \818_b0 , \819_b1 , \819_b0 , 
		\820_b1 , \820_b0 , \821_b1 , \821_b0 , \822_b1 , \822_b0 , \823_b1 , \823_b0 , \824_b1 , \824_b0 , 
		\825_b1 , \825_b0 , \826_b1 , \826_b0 , \827_b1 , \827_b0 , \828_b1 , \828_b0 , \829_b1 , \829_b0 , 
		\830_b1 , \830_b0 , \831_b1 , \831_b0 , \832_b1 , \832_b0 , \833_b1 , \833_b0 , \834_b1 , \834_b0 , 
		\835_b1 , \835_b0 , \836_b1 , \836_b0 , \837_b1 , \837_b0 , \838_b1 , \838_b0 , \839_b1 , \839_b0 , 
		\840_b1 , \840_b0 , \841_b1 , \841_b0 , \842_b1 , \842_b0 , \843_b1 , \843_b0 , \844_b1 , \844_b0 , 
		\845_b1 , \845_b0 , \846_b1 , \846_b0 , \847_b1 , \847_b0 , \848_b1 , \848_b0 , \849_b1 , \849_b0 , 
		\850_b1 , \850_b0 , \851_b1 , \851_b0 , \852_b1 , \852_b0 , \853_b1 , \853_b0 , \854_b1 , \854_b0 , 
		\855_b1 , \855_b0 , \856_b1 , \856_b0 , \857_b1 , \857_b0 , \858_b1 , \858_b0 , \859_b1 , \859_b0 , 
		\860_b1 , \860_b0 , \861_b1 , \861_b0 , \862_b1 , \862_b0 , \863_b1 , \863_b0 , \864_b1 , \864_b0 , 
		\865_b1 , \865_b0 , \866_b1 , \866_b0 , \867_b1 , \867_b0 , \868_b1 , \868_b0 , \869_b1 , \869_b0 , 
		\870_b1 , \870_b0 , \871_b1 , \871_b0 , \872_b1 , \872_b0 , \873_b1 , \873_b0 , \874_b1 , \874_b0 , 
		\875_b1 , \875_b0 , \876_b1 , \876_b0 , \877_b1 , \877_b0 , \878_b1 , \878_b0 , \879_b1 , \879_b0 , 
		\880_b1 , \880_b0 , \881_b1 , \881_b0 , \882_b1 , \882_b0 , \883_b1 , \883_b0 , \884_b1 , \884_b0 , 
		\885_b1 , \885_b0 , \886_b1 , \886_b0 , \887_b1 , \887_b0 , \888_b1 , \888_b0 , \889_b1 , \889_b0 , 
		\890_b1 , \890_b0 , \891_b1 , \891_b0 , \892_b1 , \892_b0 , \893_b1 , \893_b0 , \894_b1 , \894_b0 , 
		\895_b1 , \895_b0 , \896_b1 , \896_b0 , \897_b1 , \897_b0 , \898_b1 , \898_b0 , \899_b1 , \899_b0 , 
		\900_b1 , \900_b0 , \901_b1 , \901_b0 , \902_b1 , \902_b0 , \903_b1 , \903_b0 , \904_b1 , \904_b0 , 
		\905_b1 , \905_b0 , \906_b1 , \906_b0 , \907_b1 , \907_b0 , \908_b1 , \908_b0 , \909_b1 , \909_b0 , 
		\910_b1 , \910_b0 , \911_b1 , \911_b0 , \912_b1 , \912_b0 , \913_b1 , \913_b0 , \914_b1 , \914_b0 , 
		\915_b1 , \915_b0 , \916_b1 , \916_b0 , \917_b1 , \917_b0 , \918_b1 , \918_b0 , \919_b1 , \919_b0 , 
		\920_b1 , \920_b0 , \921_b1 , \921_b0 , \922_b1 , \922_b0 , \923_b1 , \923_b0 , \924_b1 , \924_b0 , 
		\925_b1 , \925_b0 , \926_b1 , \926_b0 , \927_b1 , \927_b0 , \928_b1 , \928_b0 , \929_b1 , \929_b0 , 
		\930_b1 , \930_b0 , \931_b1 , \931_b0 , \932_b1 , \932_b0 , \933_b1 , \933_b0 , \934_b1 , \934_b0 , 
		\935_b1 , \935_b0 , \936_b1 , \936_b0 , \937_b1 , \937_b0 , \938_b1 , \938_b0 , \939_b1 , \939_b0 , 
		\940_b1 , \940_b0 , \941_b1 , \941_b0 , \942_b1 , \942_b0 , \943_b1 , \943_b0 , \944_b1 , \944_b0 , 
		\945_b1 , \945_b0 , \946_b1 , \946_b0 , \947_b1 , \947_b0 , \948_b1 , \948_b0 , \949_b1 , \949_b0 , 
		\950_b1 , \950_b0 , \951_b1 , \951_b0 , \952_b1 , \952_b0 , \953_b1 , \953_b0 , \954_b1 , \954_b0 , 
		\955_b1 , \955_b0 , \956_b1 , \956_b0 , \957_b1 , \957_b0 , \958_b1 , \958_b0 , \959_b1 , \959_b0 , 
		\960_b1 , \960_b0 , \961_b1 , \961_b0 , \962_b1 , \962_b0 , \963_b1 , \963_b0 , \964_b1 , \964_b0 , 
		\965_b1 , \965_b0 , \966_b1 , \966_b0 , \967_b1 , \967_b0 , \968_b1 , \968_b0 , \969_b1 , \969_b0 , 
		\970_b1 , \970_b0 , \971_b1 , \971_b0 , \972_b1 , \972_b0 , \973_b1 , \973_b0 , \974_b1 , \974_b0 , 
		\975_b1 , \975_b0 , \976_b1 , \976_b0 , \977_b1 , \977_b0 , \978_nR132_b1 , \978_nR132_b0 , \979_b1 , \979_b0 , 
		\980_nR131_b1 , \980_nR131_b0 , \981_b1 , \981_b0 , \982_b1 , \982_b0 , \983_b1 , \983_b0 , \984_b1 , \984_b0 , 
		\985_b1 , \985_b0 , \986_b1 , \986_b0 , \987_b1 , \987_b0 , \988_b1 , \988_b0 , \989_b1 , \989_b0 , 
		\990_b1 , \990_b0 , \991_b1 , \991_b0 , \992_b1 , \992_b0 , \993_b1 , \993_b0 , \994_b1 , \994_b0 , 
		\995_b1 , \995_b0 , \996_b1 , \996_b0 , \997_b1 , \997_b0 , \998_b1 , \998_b0 , \999_b1 , \999_b0 , 
		\1000_b1 , \1000_b0 , \1001_b1 , \1001_b0 , \1002_b1 , \1002_b0 , \1003_b1 , \1003_b0 , \1004_b1 , \1004_b0 , 
		\1005_b1 , \1005_b0 , \1006_b1 , \1006_b0 , \1007_b1 , \1007_b0 , \1008_b1 , \1008_b0 , \1009_b1 , \1009_b0 , 
		\1010_b1 , \1010_b0 , \1011_b1 , \1011_b0 , \1012_b1 , \1012_b0 , \1013_b1 , \1013_b0 , \1014_b1 , \1014_b0 , 
		\1015_b1 , \1015_b0 , \1016_b1 , \1016_b0 , \1017_b1 , \1017_b0 , \1018_b1 , \1018_b0 , \1019_b1 , \1019_b0 , 
		\1020_b1 , \1020_b0 , \1021_b1 , \1021_b0 , \1022_b1 , \1022_b0 , \1023_b1 , \1023_b0 , \1024_b1 , \1024_b0 , 
		\1025_b1 , \1025_b0 , \1026_b1 , \1026_b0 , \1027_b1 , \1027_b0 , \1028_b1 , \1028_b0 , \1029_b1 , \1029_b0 , 
		\1030_b1 , \1030_b0 , \1031_b1 , \1031_b0 , \1032_b1 , \1032_b0 , \1033_b1 , \1033_b0 , \1034_b1 , \1034_b0 , 
		\1035_b1 , \1035_b0 , \1036_b1 , \1036_b0 , \1037_b1 , \1037_b0 , \1038_b1 , \1038_b0 , \1039_b1 , \1039_b0 , 
		\1040_b1 , \1040_b0 , \1041_b1 , \1041_b0 , \1042_b1 , \1042_b0 , \1043_b1 , \1043_b0 , \1044_b1 , \1044_b0 , 
		\1045_b1 , \1045_b0 , \1046_b1 , \1046_b0 , \1047_b1 , \1047_b0 , \1048_b1 , \1048_b0 , \1049_b1 , \1049_b0 , 
		\1050_b1 , \1050_b0 , \1051_b1 , \1051_b0 , \1052_b1 , \1052_b0 , \1053_b1 , \1053_b0 , \1054_b1 , \1054_b0 , 
		\1055_b1 , \1055_b0 , \1056_b1 , \1056_b0 , \1057_b1 , \1057_b0 , \1058_b1 , \1058_b0 , \1059_b1 , \1059_b0 , 
		\1060_b1 , \1060_b0 , \1061_b1 , \1061_b0 , \1062_b1 , \1062_b0 , \1063_b1 , \1063_b0 , \1064_b1 , \1064_b0 , 
		\1065_b1 , \1065_b0 , \1066_b1 , \1066_b0 , \1067_b1 , \1067_b0 , \1068_b1 , \1068_b0 , \1069_b1 , \1069_b0 , 
		\1070_b1 , \1070_b0 , \1071_b1 , \1071_b0 , \1072_b1 , \1072_b0 , \1073_b1 , \1073_b0 , \1074_b1 , \1074_b0 , 
		\1075_b1 , \1075_b0 , \1076_b1 , \1076_b0 , \1077_b1 , \1077_b0 , \1078_b1 , \1078_b0 , \1079_b1 , \1079_b0 , 
		\1080_b1 , \1080_b0 , \1081_b1 , \1081_b0 , \1082_b1 , \1082_b0 , \1083_b1 , \1083_b0 , \1084_b1 , \1084_b0 , 
		\1085_b1 , \1085_b0 , \1086_b1 , \1086_b0 , \1087_b1 , \1087_b0 , \1088_b1 , \1088_b0 , \1089_b1 , \1089_b0 , 
		\1090_b1 , \1090_b0 , \1091_b1 , \1091_b0 , \1092_b1 , \1092_b0 , \1093_b1 , \1093_b0 , \1094_b1 , \1094_b0 , 
		\1095_b1 , \1095_b0 , \1096_b1 , \1096_b0 , \1097_b1 , \1097_b0 , \1098_b1 , \1098_b0 , \1099_b1 , \1099_b0 , 
		\1100_b1 , \1100_b0 , \1101_b1 , \1101_b0 , \1102_b1 , \1102_b0 , \1103_b1 , \1103_b0 , \1104_b1 , \1104_b0 , 
		\1105_b1 , \1105_b0 , \1106_b1 , \1106_b0 , \1107_b1 , \1107_b0 , \1108_b1 , \1108_b0 , \1109_b1 , \1109_b0 , 
		\1110_b1 , \1110_b0 , \1111_b1 , \1111_b0 , \1112_b1 , \1112_b0 , \1113_b1 , \1113_b0 , \1114_b1 , \1114_b0 , 
		\1115_b1 , \1115_b0 , \1116_b1 , \1116_b0 , \1117_b1 , \1117_b0 , \1118_b1 , \1118_b0 , \1119_b1 , \1119_b0 , 
		\1120_b1 , \1120_b0 , \1121_b1 , \1121_b0 , \1122_b1 , \1122_b0 , \1123_b1 , \1123_b0 , \1124_b1 , \1124_b0 , 
		\1125_b1 , \1125_b0 , \1126_b1 , \1126_b0 , \1127_b1 , \1127_b0 , \1128_b1 , \1128_b0 , \1129_b1 , \1129_b0 , 
		\1130_b1 , \1130_b0 , \1131_b1 , \1131_b0 , \1132_b1 , \1132_b0 , \1133_b1 , \1133_b0 , \1134_b1 , \1134_b0 , 
		\1135_b1 , \1135_b0 , \1136_b1 , \1136_b0 , \1137_b1 , \1137_b0 , \1138_b1 , \1138_b0 , \1139_b1 , \1139_b0 , 
		\1140_b1 , \1140_b0 , \1141_b1 , \1141_b0 , \1142_b1 , \1142_b0 , \1143_b1 , \1143_b0 , \1144_b1 , \1144_b0 , 
		\1145_b1 , \1145_b0 , \1146_b1 , \1146_b0 , \1147_b1 , \1147_b0 , \1148_b1 , \1148_b0 , \1149_b1 , \1149_b0 , 
		\1150_b1 , \1150_b0 , \1151_b1 , \1151_b0 , \1152_b1 , \1152_b0 , \1153_b1 , \1153_b0 , \1154_b1 , \1154_b0 , 
		\1155_b1 , \1155_b0 , \1156_b1 , \1156_b0 , \1157_b1 , \1157_b0 , \1158_b1 , \1158_b0 , \1159_b1 , \1159_b0 , 
		\1160_b1 , \1160_b0 , \1161_b1 , \1161_b0 , \1162_b1 , \1162_b0 , \1163_b1 , \1163_b0 , \1164_b1 , \1164_b0 , 
		\1165_b1 , \1165_b0 , \1166_b1 , \1166_b0 , \1167_b1 , \1167_b0 , \1168_b1 , \1168_b0 , \1169_b1 , \1169_b0 , 
		\1170_b1 , \1170_b0 , \1171_nR130_b1 , \1171_nR130_b0 , \1172_b1 , \1172_b0 , \1173_nR12f_b1 , \1173_nR12f_b0 , \1174_b1 , \1174_b0 , 
		\1175_b1 , \1175_b0 , \1176_b1 , \1176_b0 , \1177_b1 , \1177_b0 , \1178_b1 , \1178_b0 , \1179_b1 , \1179_b0 , 
		\1180_b1 , \1180_b0 , \1181_b1 , \1181_b0 , \1182_b1 , \1182_b0 , \1183_b1 , \1183_b0 , \1184_b1 , \1184_b0 , 
		\1185_b1 , \1185_b0 , \1186_b1 , \1186_b0 , \1187_b1 , \1187_b0 , \1188_b1 , \1188_b0 , \1189_b1 , \1189_b0 , 
		\1190_b1 , \1190_b0 , \1191_b1 , \1191_b0 , \1192_b1 , \1192_b0 , \1193_b1 , \1193_b0 , \1194_b1 , \1194_b0 , 
		\1195_b1 , \1195_b0 , \1196_b1 , \1196_b0 , \1197_b1 , \1197_b0 , \1198_b1 , \1198_b0 , \1199_b1 , \1199_b0 , 
		\1200_b1 , \1200_b0 , \1201_b1 , \1201_b0 , \1202_b1 , \1202_b0 , \1203_b1 , \1203_b0 , \1204_b1 , \1204_b0 , 
		\1205_b1 , \1205_b0 , \1206_b1 , \1206_b0 , \1207_b1 , \1207_b0 , \1208_b1 , \1208_b0 , \1209_b1 , \1209_b0 , 
		\1210_b1 , \1210_b0 , \1211_b1 , \1211_b0 , \1212_b1 , \1212_b0 , \1213_b1 , \1213_b0 , \1214_b1 , \1214_b0 , 
		\1215_b1 , \1215_b0 , \1216_b1 , \1216_b0 , \1217_b1 , \1217_b0 , \1218_b1 , \1218_b0 , \1219_b1 , \1219_b0 , 
		\1220_b1 , \1220_b0 , \1221_b1 , \1221_b0 , \1222_b1 , \1222_b0 , \1223_b1 , \1223_b0 , \1224_b1 , \1224_b0 , 
		\1225_b1 , \1225_b0 , \1226_b1 , \1226_b0 , \1227_b1 , \1227_b0 , \1228_b1 , \1228_b0 , \1229_b1 , \1229_b0 , 
		\1230_b1 , \1230_b0 , \1231_b1 , \1231_b0 , \1232_b1 , \1232_b0 , \1233_b1 , \1233_b0 , \1234_b1 , \1234_b0 , 
		\1235_b1 , \1235_b0 , \1236_b1 , \1236_b0 , \1237_b1 , \1237_b0 , \1238_b1 , \1238_b0 , \1239_b1 , \1239_b0 , 
		\1240_b1 , \1240_b0 , \1241_b1 , \1241_b0 , \1242_b1 , \1242_b0 , \1243_b1 , \1243_b0 , \1244_b1 , \1244_b0 , 
		\1245_b1 , \1245_b0 , \1246_b1 , \1246_b0 , \1247_b1 , \1247_b0 , \1248_b1 , \1248_b0 , \1249_b1 , \1249_b0 , 
		\1250_b1 , \1250_b0 , \1251_b1 , \1251_b0 , \1252_b1 , \1252_b0 , \1253_b1 , \1253_b0 , \1254_b1 , \1254_b0 , 
		\1255_b1 , \1255_b0 , \1256_b1 , \1256_b0 , \1257_b1 , \1257_b0 , \1258_b1 , \1258_b0 , \1259_b1 , \1259_b0 , 
		\1260_b1 , \1260_b0 , \1261_b1 , \1261_b0 , \1262_b1 , \1262_b0 , \1263_b1 , \1263_b0 , \1264_b1 , \1264_b0 , 
		\1265_b1 , \1265_b0 , \1266_b1 , \1266_b0 , \1267_b1 , \1267_b0 , \1268_b1 , \1268_b0 , \1269_b1 , \1269_b0 , 
		\1270_b1 , \1270_b0 , \1271_b1 , \1271_b0 , \1272_b1 , \1272_b0 , \1273_b1 , \1273_b0 , \1274_b1 , \1274_b0 , 
		\1275_b1 , \1275_b0 , \1276_b1 , \1276_b0 , \1277_b1 , \1277_b0 , \1278_b1 , \1278_b0 , \1279_b1 , \1279_b0 , 
		\1280_b1 , \1280_b0 , \1281_b1 , \1281_b0 , \1282_b1 , \1282_b0 , \1283_b1 , \1283_b0 , \1284_b1 , \1284_b0 , 
		\1285_b1 , \1285_b0 , \1286_b1 , \1286_b0 , \1287_b1 , \1287_b0 , \1288_b1 , \1288_b0 , \1289_b1 , \1289_b0 , 
		\1290_b1 , \1290_b0 , \1291_b1 , \1291_b0 , \1292_b1 , \1292_b0 , \1293_b1 , \1293_b0 , \1294_b1 , \1294_b0 , 
		\1295_b1 , \1295_b0 , \1296_b1 , \1296_b0 , \1297_b1 , \1297_b0 , \1298_b1 , \1298_b0 , \1299_b1 , \1299_b0 , 
		\1300_b1 , \1300_b0 , \1301_b1 , \1301_b0 , \1302_b1 , \1302_b0 , \1303_b1 , \1303_b0 , \1304_b1 , \1304_b0 , 
		\1305_b1 , \1305_b0 , \1306_b1 , \1306_b0 , \1307_b1 , \1307_b0 , \1308_b1 , \1308_b0 , \1309_b1 , \1309_b0 , 
		\1310_b1 , \1310_b0 , \1311_b1 , \1311_b0 , \1312_b1 , \1312_b0 , \1313_b1 , \1313_b0 , \1314_b1 , \1314_b0 , 
		\1315_b1 , \1315_b0 , \1316_b1 , \1316_b0 , \1317_b1 , \1317_b0 , \1318_b1 , \1318_b0 , \1319_b1 , \1319_b0 , 
		\1320_b1 , \1320_b0 , \1321_b1 , \1321_b0 , \1322_b1 , \1322_b0 , \1323_b1 , \1323_b0 , \1324_b1 , \1324_b0 , 
		\1325_b1 , \1325_b0 , \1326_b1 , \1326_b0 , \1327_b1 , \1327_b0 , \1328_b1 , \1328_b0 , \1329_b1 , \1329_b0 , 
		\1330_b1 , \1330_b0 , \1331_b1 , \1331_b0 , \1332_b1 , \1332_b0 , \1333_b1 , \1333_b0 , \1334_b1 , \1334_b0 , 
		\1335_b1 , \1335_b0 , \1336_b1 , \1336_b0 , \1337_b1 , \1337_b0 , \1338_b1 , \1338_b0 , \1339_b1 , \1339_b0 , 
		\1340_b1 , \1340_b0 , \1341_b1 , \1341_b0 , \1342_b1 , \1342_b0 , \1343_b1 , \1343_b0 , \1344_b1 , \1344_b0 , 
		\1345_b1 , \1345_b0 , \1346_b1 , \1346_b0 , \1347_b1 , \1347_b0 , \1348_b1 , \1348_b0 , \1349_b1 , \1349_b0 , 
		\1350_b1 , \1350_b0 , \1351_b1 , \1351_b0 , \1352_b1 , \1352_b0 , \1353_b1 , \1353_b0 , \1354_b1 , \1354_b0 , 
		\1355_b1 , \1355_b0 , \1356_b1 , \1356_b0 , \1357_nR12e_b1 , \1357_nR12e_b0 , \1358_b1 , \1358_b0 , \1359_nR12d_b1 , \1359_nR12d_b0 , 
		\1360_b1 , \1360_b0 , \1361_b1 , \1361_b0 , \1362_b1 , \1362_b0 , \1363_b1 , \1363_b0 , \1364_b1 , \1364_b0 , 
		\1365_b1 , \1365_b0 , \1366_b1 , \1366_b0 , \1367_b1 , \1367_b0 , \1368_b1 , \1368_b0 , \1369_b1 , \1369_b0 , 
		\1370_b1 , \1370_b0 , \1371_b1 , \1371_b0 , \1372_b1 , \1372_b0 , \1373_b1 , \1373_b0 , \1374_b1 , \1374_b0 , 
		\1375_b1 , \1375_b0 , \1376_b1 , \1376_b0 , \1377_b1 , \1377_b0 , \1378_b1 , \1378_b0 , \1379_b1 , \1379_b0 , 
		\1380_b1 , \1380_b0 , \1381_b1 , \1381_b0 , \1382_b1 , \1382_b0 , \1383_b1 , \1383_b0 , \1384_b1 , \1384_b0 , 
		\1385_b1 , \1385_b0 , \1386_b1 , \1386_b0 , \1387_b1 , \1387_b0 , \1388_b1 , \1388_b0 , \1389_b1 , \1389_b0 , 
		\1390_b1 , \1390_b0 , \1391_b1 , \1391_b0 , \1392_b1 , \1392_b0 , \1393_b1 , \1393_b0 , \1394_b1 , \1394_b0 , 
		\1395_b1 , \1395_b0 , \1396_b1 , \1396_b0 , \1397_b1 , \1397_b0 , \1398_b1 , \1398_b0 , \1399_b1 , \1399_b0 , 
		\1400_b1 , \1400_b0 , \1401_b1 , \1401_b0 , \1402_b1 , \1402_b0 , \1403_b1 , \1403_b0 , \1404_b1 , \1404_b0 , 
		\1405_b1 , \1405_b0 , \1406_b1 , \1406_b0 , \1407_b1 , \1407_b0 , \1408_b1 , \1408_b0 , \1409_b1 , \1409_b0 , 
		\1410_b1 , \1410_b0 , \1411_b1 , \1411_b0 , \1412_b1 , \1412_b0 , \1413_b1 , \1413_b0 , \1414_b1 , \1414_b0 , 
		\1415_b1 , \1415_b0 , \1416_b1 , \1416_b0 , \1417_b1 , \1417_b0 , \1418_b1 , \1418_b0 , \1419_b1 , \1419_b0 , 
		\1420_b1 , \1420_b0 , \1421_b1 , \1421_b0 , \1422_b1 , \1422_b0 , \1423_b1 , \1423_b0 , \1424_b1 , \1424_b0 , 
		\1425_b1 , \1425_b0 , \1426_b1 , \1426_b0 , \1427_b1 , \1427_b0 , \1428_b1 , \1428_b0 , \1429_b1 , \1429_b0 , 
		\1430_b1 , \1430_b0 , \1431_b1 , \1431_b0 , \1432_b1 , \1432_b0 , \1433_b1 , \1433_b0 , \1434_b1 , \1434_b0 , 
		\1435_b1 , \1435_b0 , \1436_b1 , \1436_b0 , \1437_b1 , \1437_b0 , \1438_b1 , \1438_b0 , \1439_b1 , \1439_b0 , 
		\1440_b1 , \1440_b0 , \1441_b1 , \1441_b0 , \1442_b1 , \1442_b0 , \1443_b1 , \1443_b0 , \1444_b1 , \1444_b0 , 
		\1445_b1 , \1445_b0 , \1446_b1 , \1446_b0 , \1447_b1 , \1447_b0 , \1448_b1 , \1448_b0 , \1449_b1 , \1449_b0 , 
		\1450_b1 , \1450_b0 , \1451_b1 , \1451_b0 , \1452_b1 , \1452_b0 , \1453_b1 , \1453_b0 , \1454_b1 , \1454_b0 , 
		\1455_b1 , \1455_b0 , \1456_b1 , \1456_b0 , \1457_b1 , \1457_b0 , \1458_b1 , \1458_b0 , \1459_b1 , \1459_b0 , 
		\1460_b1 , \1460_b0 , \1461_b1 , \1461_b0 , \1462_b1 , \1462_b0 , \1463_b1 , \1463_b0 , \1464_b1 , \1464_b0 , 
		\1465_b1 , \1465_b0 , \1466_b1 , \1466_b0 , \1467_b1 , \1467_b0 , \1468_b1 , \1468_b0 , \1469_b1 , \1469_b0 , 
		\1470_b1 , \1470_b0 , \1471_b1 , \1471_b0 , \1472_b1 , \1472_b0 , \1473_b1 , \1473_b0 , \1474_b1 , \1474_b0 , 
		\1475_b1 , \1475_b0 , \1476_b1 , \1476_b0 , \1477_b1 , \1477_b0 , \1478_b1 , \1478_b0 , \1479_b1 , \1479_b0 , 
		\1480_b1 , \1480_b0 , \1481_b1 , \1481_b0 , \1482_b1 , \1482_b0 , \1483_b1 , \1483_b0 , \1484_b1 , \1484_b0 , 
		\1485_b1 , \1485_b0 , \1486_b1 , \1486_b0 , \1487_b1 , \1487_b0 , \1488_b1 , \1488_b0 , \1489_b1 , \1489_b0 , 
		\1490_b1 , \1490_b0 , \1491_b1 , \1491_b0 , \1492_b1 , \1492_b0 , \1493_b1 , \1493_b0 , \1494_b1 , \1494_b0 , 
		\1495_b1 , \1495_b0 , \1496_b1 , \1496_b0 , \1497_b1 , \1497_b0 , \1498_b1 , \1498_b0 , \1499_b1 , \1499_b0 , 
		\1500_b1 , \1500_b0 , \1501_b1 , \1501_b0 , \1502_b1 , \1502_b0 , \1503_b1 , \1503_b0 , \1504_b1 , \1504_b0 , 
		\1505_b1 , \1505_b0 , \1506_b1 , \1506_b0 , \1507_b1 , \1507_b0 , \1508_b1 , \1508_b0 , \1509_b1 , \1509_b0 , 
		\1510_b1 , \1510_b0 , \1511_b1 , \1511_b0 , \1512_b1 , \1512_b0 , \1513_b1 , \1513_b0 , \1514_b1 , \1514_b0 , 
		\1515_b1 , \1515_b0 , \1516_b1 , \1516_b0 , \1517_b1 , \1517_b0 , \1518_b1 , \1518_b0 , \1519_b1 , \1519_b0 , 
		\1520_b1 , \1520_b0 , \1521_b1 , \1521_b0 , \1522_b1 , \1522_b0 , \1523_b1 , \1523_b0 , \1524_b1 , \1524_b0 , 
		\1525_b1 , \1525_b0 , \1526_b1 , \1526_b0 , \1527_b1 , \1527_b0 , \1528_b1 , \1528_b0 , \1529_b1 , \1529_b0 , 
		\1530_b1 , \1530_b0 , \1531_b1 , \1531_b0 , \1532_b1 , \1532_b0 , \1533_b1 , \1533_b0 , \1534_b1 , \1534_b0 , 
		\1535_b1 , \1535_b0 , \1536_b1 , \1536_b0 , \1537_b1 , \1537_b0 , \1538_b1 , \1538_b0 , \1539_b1 , \1539_b0 , 
		\1540_b1 , \1540_b0 , \1541_b1 , \1541_b0 , \1542_b1 , \1542_b0 , \1543_b1 , \1543_b0 , \1544_b1 , \1544_b0 , 
		\1545_b1 , \1545_b0 , \1546_b1 , \1546_b0 , \1547_b1 , \1547_b0 , \1548_b1 , \1548_b0 , \1549_b1 , \1549_b0 , 
		\1550_b1 , \1550_b0 , \1551_b1 , \1551_b0 , \1552_b1 , \1552_b0 , \1553_b1 , \1553_b0 , \1554_b1 , \1554_b0 , 
		\1555_b1 , \1555_b0 , \1556_b1 , \1556_b0 , \1557_b1 , \1557_b0 , \1558_b1 , \1558_b0 , \1559_b1 , \1559_b0 , 
		\1560_b1 , \1560_b0 , \1561_b1 , \1561_b0 , \1562_b1 , \1562_b0 , \1563_b1 , \1563_b0 , \1564_b1 , \1564_b0 , 
		\1565_b1 , \1565_b0 , \1566_b1 , \1566_b0 , \1567_b1 , \1567_b0 , \1568_b1 , \1568_b0 , \1569_b1 , \1569_b0 , 
		\1570_b1 , \1570_b0 , \1571_b1 , \1571_b0 , \1572_b1 , \1572_b0 , \1573_b1 , \1573_b0 , \1574_b1 , \1574_b0 , 
		\1575_b1 , \1575_b0 , \1576_b1 , \1576_b0 , \1577_b1 , \1577_b0 , \1578_b1 , \1578_b0 , \1579_b1 , \1579_b0 , 
		\1580_b1 , \1580_b0 , \1581_b1 , \1581_b0 , \1582_b1 , \1582_b0 , \1583_b1 , \1583_b0 , \1584_b1 , \1584_b0 , 
		\1585_b1 , \1585_b0 , \1586_b1 , \1586_b0 , \1587_b1 , \1587_b0 , \1588_b1 , \1588_b0 , \1589_b1 , \1589_b0 , 
		\1590_b1 , \1590_b0 , \1591_b1 , \1591_b0 , \1592_b1 , \1592_b0 , \1593_b1 , \1593_b0 , \1594_b1 , \1594_b0 , 
		\1595_b1 , \1595_b0 , \1596_b1 , \1596_b0 , \1597_b1 , \1597_b0 , \1598_b1 , \1598_b0 , \1599_b1 , \1599_b0 , 
		\1600_b1 , \1600_b0 , \1601_b1 , \1601_b0 , \1602_b1 , \1602_b0 , \1603_b1 , \1603_b0 , \1604_nR12c_b1 , \1604_nR12c_b0 , 
		\1605_b1 , \1605_b0 , \1606_nR12b_b1 , \1606_nR12b_b0 , \1607_b1 , \1607_b0 , \1608_b1 , \1608_b0 , \1609_b1 , \1609_b0 , 
		\1610_b1 , \1610_b0 , \1611_b1 , \1611_b0 , \1612_b1 , \1612_b0 , \1613_b1 , \1613_b0 , \1614_b1 , \1614_b0 , 
		\1615_b1 , \1615_b0 , \1616_b1 , \1616_b0 , \1617_b1 , \1617_b0 , \1618_b1 , \1618_b0 , \1619_b1 , \1619_b0 , 
		\1620_b1 , \1620_b0 , \1621_b1 , \1621_b0 , \1622_b1 , \1622_b0 , \1623_b1 , \1623_b0 , \1624_b1 , \1624_b0 , 
		\1625_b1 , \1625_b0 , \1626_b1 , \1626_b0 , \1627_b1 , \1627_b0 , \1628_b1 , \1628_b0 , \1629_b1 , \1629_b0 , 
		\1630_b1 , \1630_b0 , \1631_b1 , \1631_b0 , \1632_b1 , \1632_b0 , \1633_b1 , \1633_b0 , \1634_b1 , \1634_b0 , 
		\1635_b1 , \1635_b0 , \1636_b1 , \1636_b0 , \1637_b1 , \1637_b0 , \1638_b1 , \1638_b0 , \1639_b1 , \1639_b0 , 
		\1640_b1 , \1640_b0 , \1641_b1 , \1641_b0 , \1642_b1 , \1642_b0 , \1643_b1 , \1643_b0 , \1644_b1 , \1644_b0 , 
		\1645_b1 , \1645_b0 , \1646_b1 , \1646_b0 , \1647_b1 , \1647_b0 , \1648_b1 , \1648_b0 , \1649_b1 , \1649_b0 , 
		\1650_b1 , \1650_b0 , \1651_b1 , \1651_b0 , \1652_b1 , \1652_b0 , \1653_b1 , \1653_b0 , \1654_b1 , \1654_b0 , 
		\1655_b1 , \1655_b0 , \1656_b1 , \1656_b0 , \1657_b1 , \1657_b0 , \1658_b1 , \1658_b0 , \1659_b1 , \1659_b0 , 
		\1660_b1 , \1660_b0 , \1661_b1 , \1661_b0 , \1662_b1 , \1662_b0 , \1663_b1 , \1663_b0 , \1664_b1 , \1664_b0 , 
		\1665_b1 , \1665_b0 , \1666_b1 , \1666_b0 , \1667_b1 , \1667_b0 , \1668_b1 , \1668_b0 , \1669_b1 , \1669_b0 , 
		\1670_b1 , \1670_b0 , \1671_b1 , \1671_b0 , \1672_b1 , \1672_b0 , \1673_b1 , \1673_b0 , \1674_b1 , \1674_b0 , 
		\1675_b1 , \1675_b0 , \1676_b1 , \1676_b0 , \1677_b1 , \1677_b0 , \1678_b1 , \1678_b0 , \1679_b1 , \1679_b0 , 
		\1680_b1 , \1680_b0 , \1681_b1 , \1681_b0 , \1682_b1 , \1682_b0 , \1683_b1 , \1683_b0 , \1684_b1 , \1684_b0 , 
		\1685_b1 , \1685_b0 , \1686_b1 , \1686_b0 , \1687_b1 , \1687_b0 , \1688_b1 , \1688_b0 , \1689_b1 , \1689_b0 , 
		\1690_b1 , \1690_b0 , \1691_b1 , \1691_b0 , \1692_b1 , \1692_b0 , \1693_b1 , \1693_b0 , \1694_b1 , \1694_b0 , 
		\1695_b1 , \1695_b0 , \1696_b1 , \1696_b0 , \1697_b1 , \1697_b0 , \1698_b1 , \1698_b0 , \1699_b1 , \1699_b0 , 
		\1700_b1 , \1700_b0 , \1701_b1 , \1701_b0 , \1702_b1 , \1702_b0 , \1703_b1 , \1703_b0 , \1704_b1 , \1704_b0 , 
		\1705_b1 , \1705_b0 , \1706_b1 , \1706_b0 , \1707_b1 , \1707_b0 , \1708_b1 , \1708_b0 , \1709_b1 , \1709_b0 , 
		\1710_b1 , \1710_b0 , \1711_b1 , \1711_b0 , \1712_b1 , \1712_b0 , \1713_b1 , \1713_b0 , \1714_b1 , \1714_b0 , 
		\1715_b1 , \1715_b0 , \1716_b1 , \1716_b0 , \1717_b1 , \1717_b0 , \1718_b1 , \1718_b0 , \1719_b1 , \1719_b0 , 
		\1720_b1 , \1720_b0 , \1721_b1 , \1721_b0 , \1722_b1 , \1722_b0 , \1723_b1 , \1723_b0 , \1724_b1 , \1724_b0 , 
		\1725_b1 , \1725_b0 , \1726_b1 , \1726_b0 , \1727_b1 , \1727_b0 , \1728_b1 , \1728_b0 , \1729_b1 , \1729_b0 , 
		\1730_b1 , \1730_b0 , \1731_b1 , \1731_b0 , \1732_b1 , \1732_b0 , \1733_b1 , \1733_b0 , \1734_b1 , \1734_b0 , 
		\1735_b1 , \1735_b0 , \1736_b1 , \1736_b0 , \1737_b1 , \1737_b0 , \1738_b1 , \1738_b0 , \1739_b1 , \1739_b0 , 
		\1740_b1 , \1740_b0 , \1741_b1 , \1741_b0 , \1742_b1 , \1742_b0 , \1743_b1 , \1743_b0 , \1744_b1 , \1744_b0 , 
		\1745_b1 , \1745_b0 , \1746_b1 , \1746_b0 , \1747_b1 , \1747_b0 , \1748_b1 , \1748_b0 , \1749_b1 , \1749_b0 , 
		\1750_b1 , \1750_b0 , \1751_b1 , \1751_b0 , \1752_b1 , \1752_b0 , \1753_b1 , \1753_b0 , \1754_b1 , \1754_b0 , 
		\1755_b1 , \1755_b0 , \1756_b1 , \1756_b0 , \1757_b1 , \1757_b0 , \1758_b1 , \1758_b0 , \1759_b1 , \1759_b0 , 
		\1760_b1 , \1760_b0 , \1761_b1 , \1761_b0 , \1762_b1 , \1762_b0 , \1763_b1 , \1763_b0 , \1764_b1 , \1764_b0 , 
		\1765_b1 , \1765_b0 , \1766_b1 , \1766_b0 , \1767_b1 , \1767_b0 , \1768_b1 , \1768_b0 , \1769_b1 , \1769_b0 , 
		\1770_b1 , \1770_b0 , \1771_b1 , \1771_b0 , \1772_b1 , \1772_b0 , \1773_b1 , \1773_b0 , \1774_b1 , \1774_b0 , 
		\1775_b1 , \1775_b0 , \1776_b1 , \1776_b0 , \1777_b1 , \1777_b0 , \1778_b1 , \1778_b0 , \1779_b1 , \1779_b0 , 
		\1780_b1 , \1780_b0 , \1781_b1 , \1781_b0 , \1782_b1 , \1782_b0 , \1783_b1 , \1783_b0 , \1784_b1 , \1784_b0 , 
		\1785_b1 , \1785_b0 , \1786_b1 , \1786_b0 , \1787_b1 , \1787_b0 , \1788_b1 , \1788_b0 , \1789_b1 , \1789_b0 , 
		\1790_b1 , \1790_b0 , \1791_b1 , \1791_b0 , \1792_b1 , \1792_b0 , \1793_b1 , \1793_b0 , \1794_b1 , \1794_b0 , 
		\1795_b1 , \1795_b0 , \1796_b1 , \1796_b0 , \1797_b1 , \1797_b0 , \1798_b1 , \1798_b0 , \1799_b1 , \1799_b0 , 
		\1800_b1 , \1800_b0 , \1801_b1 , \1801_b0 , \1802_b1 , \1802_b0 , \1803_b1 , \1803_b0 , \1804_b1 , \1804_b0 , 
		\1805_b1 , \1805_b0 , \1806_b1 , \1806_b0 , \1807_b1 , \1807_b0 , \1808_b1 , \1808_b0 , \1809_b1 , \1809_b0 , 
		\1810_b1 , \1810_b0 , \1811_b1 , \1811_b0 , \1812_b1 , \1812_b0 , \1813_b1 , \1813_b0 , \1814_b1 , \1814_b0 , 
		\1815_b1 , \1815_b0 , \1816_b1 , \1816_b0 , \1817_b1 , \1817_b0 , \1818_b1 , \1818_b0 , \1819_b1 , \1819_b0 , 
		\1820_b1 , \1820_b0 , \1821_b1 , \1821_b0 , \1822_b1 , \1822_b0 , \1823_b1 , \1823_b0 , \1824_b1 , \1824_b0 , 
		\1825_b1 , \1825_b0 , \1826_b1 , \1826_b0 , \1827_b1 , \1827_b0 , \1828_b1 , \1828_b0 , \1829_nR12a_b1 , \1829_nR12a_b0 , 
		\1830_b1 , \1830_b0 , \1831_nR129_b1 , \1831_nR129_b0 , \1832_b1 , \1832_b0 , \1833_b1 , \1833_b0 , \1834_b1 , \1834_b0 , 
		\1835_b1 , \1835_b0 , \1836_b1 , \1836_b0 , \1837_b1 , \1837_b0 , \1838_b1 , \1838_b0 , \1839_b1 , \1839_b0 , 
		\1840_b1 , \1840_b0 , \1841_b1 , \1841_b0 , \1842_b1 , \1842_b0 , \1843_b1 , \1843_b0 , \1844_b1 , \1844_b0 , 
		\1845_b1 , \1845_b0 , \1846_b1 , \1846_b0 , \1847_b1 , \1847_b0 , \1848_b1 , \1848_b0 , \1849_b1 , \1849_b0 , 
		\1850_b1 , \1850_b0 , \1851_b1 , \1851_b0 , \1852_b1 , \1852_b0 , \1853_b1 , \1853_b0 , \1854_b1 , \1854_b0 , 
		\1855_b1 , \1855_b0 , \1856_b1 , \1856_b0 , \1857_b1 , \1857_b0 , \1858_b1 , \1858_b0 , \1859_b1 , \1859_b0 , 
		\1860_b1 , \1860_b0 , \1861_b1 , \1861_b0 , \1862_b1 , \1862_b0 , \1863_b1 , \1863_b0 , \1864_b1 , \1864_b0 , 
		\1865_b1 , \1865_b0 , \1866_b1 , \1866_b0 , \1867_b1 , \1867_b0 , \1868_b1 , \1868_b0 , \1869_b1 , \1869_b0 , 
		\1870_b1 , \1870_b0 , \1871_b1 , \1871_b0 , \1872_b1 , \1872_b0 , \1873_b1 , \1873_b0 , \1874_b1 , \1874_b0 , 
		\1875_b1 , \1875_b0 , \1876_b1 , \1876_b0 , \1877_b1 , \1877_b0 , \1878_b1 , \1878_b0 , \1879_b1 , \1879_b0 , 
		\1880_b1 , \1880_b0 , \1881_b1 , \1881_b0 , \1882_b1 , \1882_b0 , \1883_b1 , \1883_b0 , \1884_b1 , \1884_b0 , 
		\1885_b1 , \1885_b0 , \1886_b1 , \1886_b0 , \1887_b1 , \1887_b0 , \1888_b1 , \1888_b0 , \1889_b1 , \1889_b0 , 
		\1890_b1 , \1890_b0 , \1891_b1 , \1891_b0 , \1892_b1 , \1892_b0 , \1893_b1 , \1893_b0 , \1894_b1 , \1894_b0 , 
		\1895_b1 , \1895_b0 , \1896_b1 , \1896_b0 , \1897_b1 , \1897_b0 , \1898_b1 , \1898_b0 , \1899_b1 , \1899_b0 , 
		\1900_b1 , \1900_b0 , \1901_b1 , \1901_b0 , \1902_b1 , \1902_b0 , \1903_b1 , \1903_b0 , \1904_b1 , \1904_b0 , 
		\1905_b1 , \1905_b0 , \1906_b1 , \1906_b0 , \1907_b1 , \1907_b0 , \1908_b1 , \1908_b0 , \1909_b1 , \1909_b0 , 
		\1910_b1 , \1910_b0 , \1911_b1 , \1911_b0 , \1912_b1 , \1912_b0 , \1913_b1 , \1913_b0 , \1914_b1 , \1914_b0 , 
		\1915_b1 , \1915_b0 , \1916_b1 , \1916_b0 , \1917_b1 , \1917_b0 , \1918_b1 , \1918_b0 , \1919_b1 , \1919_b0 , 
		\1920_b1 , \1920_b0 , \1921_b1 , \1921_b0 , \1922_b1 , \1922_b0 , \1923_b1 , \1923_b0 , \1924_b1 , \1924_b0 , 
		\1925_b1 , \1925_b0 , \1926_b1 , \1926_b0 , \1927_b1 , \1927_b0 , \1928_b1 , \1928_b0 , \1929_b1 , \1929_b0 , 
		\1930_b1 , \1930_b0 , \1931_b1 , \1931_b0 , \1932_b1 , \1932_b0 , \1933_b1 , \1933_b0 , \1934_b1 , \1934_b0 , 
		\1935_b1 , \1935_b0 , \1936_b1 , \1936_b0 , \1937_b1 , \1937_b0 , \1938_b1 , \1938_b0 , \1939_b1 , \1939_b0 , 
		\1940_b1 , \1940_b0 , \1941_b1 , \1941_b0 , \1942_b1 , \1942_b0 , \1943_b1 , \1943_b0 , \1944_b1 , \1944_b0 , 
		\1945_b1 , \1945_b0 , \1946_b1 , \1946_b0 , \1947_b1 , \1947_b0 , \1948_b1 , \1948_b0 , \1949_b1 , \1949_b0 , 
		\1950_b1 , \1950_b0 , \1951_b1 , \1951_b0 , \1952_b1 , \1952_b0 , \1953_b1 , \1953_b0 , \1954_b1 , \1954_b0 , 
		\1955_b1 , \1955_b0 , \1956_b1 , \1956_b0 , \1957_b1 , \1957_b0 , \1958_b1 , \1958_b0 , \1959_b1 , \1959_b0 , 
		\1960_b1 , \1960_b0 , \1961_b1 , \1961_b0 , \1962_b1 , \1962_b0 , \1963_b1 , \1963_b0 , \1964_b1 , \1964_b0 , 
		\1965_b1 , \1965_b0 , \1966_b1 , \1966_b0 , \1967_b1 , \1967_b0 , \1968_b1 , \1968_b0 , \1969_b1 , \1969_b0 , 
		\1970_b1 , \1970_b0 , \1971_b1 , \1971_b0 , \1972_b1 , \1972_b0 , \1973_b1 , \1973_b0 , \1974_b1 , \1974_b0 , 
		\1975_b1 , \1975_b0 , \1976_b1 , \1976_b0 , \1977_b1 , \1977_b0 , \1978_b1 , \1978_b0 , \1979_b1 , \1979_b0 , 
		\1980_b1 , \1980_b0 , \1981_b1 , \1981_b0 , \1982_b1 , \1982_b0 , \1983_b1 , \1983_b0 , \1984_b1 , \1984_b0 , 
		\1985_b1 , \1985_b0 , \1986_b1 , \1986_b0 , \1987_b1 , \1987_b0 , \1988_b1 , \1988_b0 , \1989_b1 , \1989_b0 , 
		\1990_b1 , \1990_b0 , \1991_b1 , \1991_b0 , \1992_b1 , \1992_b0 , \1993_b1 , \1993_b0 , \1994_b1 , \1994_b0 , 
		\1995_b1 , \1995_b0 , \1996_b1 , \1996_b0 , \1997_b1 , \1997_b0 , \1998_b1 , \1998_b0 , \1999_b1 , \1999_b0 , 
		\2000_b1 , \2000_b0 , \2001_b1 , \2001_b0 , \2002_b1 , \2002_b0 , \2003_b1 , \2003_b0 , \2004_b1 , \2004_b0 , 
		\2005_b1 , \2005_b0 , \2006_b1 , \2006_b0 , \2007_b1 , \2007_b0 , \2008_b1 , \2008_b0 , \2009_b1 , \2009_b0 , 
		\2010_b1 , \2010_b0 , \2011_b1 , \2011_b0 , \2012_b1 , \2012_b0 , \2013_b1 , \2013_b0 , \2014_b1 , \2014_b0 , 
		\2015_b1 , \2015_b0 , \2016_b1 , \2016_b0 , \2017_b1 , \2017_b0 , \2018_b1 , \2018_b0 , \2019_b1 , \2019_b0 , 
		\2020_b1 , \2020_b0 , \2021_b1 , \2021_b0 , \2022_b1 , \2022_b0 , \2023_b1 , \2023_b0 , \2024_b1 , \2024_b0 , 
		\2025_b1 , \2025_b0 , \2026_b1 , \2026_b0 , \2027_b1 , \2027_b0 , \2028_b1 , \2028_b0 , \2029_b1 , \2029_b0 , 
		\2030_b1 , \2030_b0 , \2031_b1 , \2031_b0 , \2032_b1 , \2032_b0 , \2033_b1 , \2033_b0 , \2034_b1 , \2034_b0 , 
		\2035_b1 , \2035_b0 , \2036_b1 , \2036_b0 , \2037_b1 , \2037_b0 , \2038_b1 , \2038_b0 , \2039_b1 , \2039_b0 , 
		\2040_b1 , \2040_b0 , \2041_b1 , \2041_b0 , \2042_b1 , \2042_b0 , \2043_b1 , \2043_b0 , \2044_b1 , \2044_b0 , 
		\2045_b1 , \2045_b0 , \2046_b1 , \2046_b0 , \2047_b1 , \2047_b0 , \2048_b1 , \2048_b0 , \2049_b1 , \2049_b0 , 
		\2050_b1 , \2050_b0 , \2051_b1 , \2051_b0 , \2052_b1 , \2052_b0 , \2053_b1 , \2053_b0 , \2054_b1 , \2054_b0 , 
		\2055_b1 , \2055_b0 , \2056_b1 , \2056_b0 , \2057_b1 , \2057_b0 , \2058_b1 , \2058_b0 , \2059_b1 , \2059_b0 , 
		\2060_b1 , \2060_b0 , \2061_b1 , \2061_b0 , \2062_b1 , \2062_b0 , \2063_b1 , \2063_b0 , \2064_b1 , \2064_b0 , 
		\2065_b1 , \2065_b0 , \2066_b1 , \2066_b0 , \2067_b1 , \2067_b0 , \2068_b1 , \2068_b0 , \2069_b1 , \2069_b0 , 
		\2070_b1 , \2070_b0 , \2071_b1 , \2071_b0 , \2072_b1 , \2072_b0 , \2073_b1 , \2073_b0 , \2074_b1 , \2074_b0 , 
		\2075_b1 , \2075_b0 , \2076_b1 , \2076_b0 , \2077_b1 , \2077_b0 , \2078_b1 , \2078_b0 , \2079_b1 , \2079_b0 , 
		\2080_b1 , \2080_b0 , \2081_b1 , \2081_b0 , \2082_b1 , \2082_b0 , \2083_b1 , \2083_b0 , \2084_b1 , \2084_b0 , 
		\2085_b1 , \2085_b0 , \2086_b1 , \2086_b0 , \2087_b1 , \2087_b0 , \2088_b1 , \2088_b0 , \2089_b1 , \2089_b0 , 
		\2090_b1 , \2090_b0 , \2091_b1 , \2091_b0 , \2092_b1 , \2092_b0 , \2093_b1 , \2093_b0 , \2094_b1 , \2094_b0 , 
		\2095_b1 , \2095_b0 , \2096_b1 , \2096_b0 , \2097_b1 , \2097_b0 , \2098_b1 , \2098_b0 , \2099_b1 , \2099_b0 , 
		\2100_b1 , \2100_b0 , \2101_b1 , \2101_b0 , \2102_b1 , \2102_b0 , \2103_b1 , \2103_b0 , \2104_b1 , \2104_b0 , 
		\2105_b1 , \2105_b0 , \2106_b1 , \2106_b0 , \2107_b1 , \2107_b0 , \2108_b1 , \2108_b0 , \2109_b1 , \2109_b0 , 
		\2110_b1 , \2110_b0 , \2111_b1 , \2111_b0 , \2112_b1 , \2112_b0 , \2113_b1 , \2113_b0 , \2114_b1 , \2114_b0 , 
		\2115_b1 , \2115_b0 , \2116_b1 , \2116_b0 , \2117_b1 , \2117_b0 , \2118_nR128_b1 , \2118_nR128_b0 , \2119_b1 , \2119_b0 , 
		\2120_nR127_b1 , \2120_nR127_b0 , \2121_b1 , \2121_b0 , \2122_b1 , \2122_b0 , \2123_b1 , \2123_b0 , \2124_b1 , \2124_b0 , 
		\2125_b1 , \2125_b0 , \2126_b1 , \2126_b0 , \2127_b1 , \2127_b0 , \2128_b1 , \2128_b0 , \2129_b1 , \2129_b0 , 
		\2130_b1 , \2130_b0 , \2131_b1 , \2131_b0 , \2132_b1 , \2132_b0 , \2133_b1 , \2133_b0 , \2134_b1 , \2134_b0 , 
		\2135_b1 , \2135_b0 , \2136_b1 , \2136_b0 , \2137_b1 , \2137_b0 , \2138_b1 , \2138_b0 , \2139_b1 , \2139_b0 , 
		\2140_b1 , \2140_b0 , \2141_b1 , \2141_b0 , \2142_b1 , \2142_b0 , \2143_b1 , \2143_b0 , \2144_b1 , \2144_b0 , 
		\2145_b1 , \2145_b0 , \2146_b1 , \2146_b0 , \2147_b1 , \2147_b0 , \2148_b1 , \2148_b0 , \2149_b1 , \2149_b0 , 
		\2150_b1 , \2150_b0 , \2151_b1 , \2151_b0 , \2152_b1 , \2152_b0 , \2153_b1 , \2153_b0 , \2154_b1 , \2154_b0 , 
		\2155_b1 , \2155_b0 , \2156_b1 , \2156_b0 , \2157_b1 , \2157_b0 , \2158_b1 , \2158_b0 , \2159_b1 , \2159_b0 , 
		\2160_b1 , \2160_b0 , \2161_b1 , \2161_b0 , \2162_b1 , \2162_b0 , \2163_b1 , \2163_b0 , \2164_b1 , \2164_b0 , 
		\2165_b1 , \2165_b0 , \2166_b1 , \2166_b0 , \2167_b1 , \2167_b0 , \2168_b1 , \2168_b0 , \2169_b1 , \2169_b0 , 
		\2170_b1 , \2170_b0 , \2171_b1 , \2171_b0 , \2172_b1 , \2172_b0 , \2173_b1 , \2173_b0 , \2174_b1 , \2174_b0 , 
		\2175_b1 , \2175_b0 , \2176_b1 , \2176_b0 , \2177_b1 , \2177_b0 , \2178_b1 , \2178_b0 , \2179_b1 , \2179_b0 , 
		\2180_b1 , \2180_b0 , \2181_b1 , \2181_b0 , \2182_b1 , \2182_b0 , \2183_b1 , \2183_b0 , \2184_b1 , \2184_b0 , 
		\2185_b1 , \2185_b0 , \2186_b1 , \2186_b0 , \2187_b1 , \2187_b0 , \2188_b1 , \2188_b0 , \2189_b1 , \2189_b0 , 
		\2190_b1 , \2190_b0 , \2191_b1 , \2191_b0 , \2192_b1 , \2192_b0 , \2193_b1 , \2193_b0 , \2194_b1 , \2194_b0 , 
		\2195_b1 , \2195_b0 , \2196_b1 , \2196_b0 , \2197_b1 , \2197_b0 , \2198_b1 , \2198_b0 , \2199_b1 , \2199_b0 , 
		\2200_b1 , \2200_b0 , \2201_b1 , \2201_b0 , \2202_b1 , \2202_b0 , \2203_b1 , \2203_b0 , \2204_b1 , \2204_b0 , 
		\2205_b1 , \2205_b0 , \2206_b1 , \2206_b0 , \2207_b1 , \2207_b0 , \2208_b1 , \2208_b0 , \2209_b1 , \2209_b0 , 
		\2210_b1 , \2210_b0 , \2211_b1 , \2211_b0 , \2212_b1 , \2212_b0 , \2213_b1 , \2213_b0 , \2214_b1 , \2214_b0 , 
		\2215_b1 , \2215_b0 , \2216_b1 , \2216_b0 , \2217_b1 , \2217_b0 , \2218_b1 , \2218_b0 , \2219_b1 , \2219_b0 , 
		\2220_b1 , \2220_b0 , \2221_b1 , \2221_b0 , \2222_b1 , \2222_b0 , \2223_b1 , \2223_b0 , \2224_b1 , \2224_b0 , 
		\2225_b1 , \2225_b0 , \2226_b1 , \2226_b0 , \2227_b1 , \2227_b0 , \2228_b1 , \2228_b0 , \2229_b1 , \2229_b0 , 
		\2230_b1 , \2230_b0 , \2231_b1 , \2231_b0 , \2232_b1 , \2232_b0 , \2233_b1 , \2233_b0 , \2234_b1 , \2234_b0 , 
		\2235_b1 , \2235_b0 , \2236_b1 , \2236_b0 , \2237_b1 , \2237_b0 , \2238_b1 , \2238_b0 , \2239_b1 , \2239_b0 , 
		\2240_b1 , \2240_b0 , \2241_b1 , \2241_b0 , \2242_b1 , \2242_b0 , \2243_b1 , \2243_b0 , \2244_b1 , \2244_b0 , 
		\2245_b1 , \2245_b0 , \2246_b1 , \2246_b0 , \2247_b1 , \2247_b0 , \2248_b1 , \2248_b0 , \2249_b1 , \2249_b0 , 
		\2250_b1 , \2250_b0 , \2251_b1 , \2251_b0 , \2252_b1 , \2252_b0 , \2253_b1 , \2253_b0 , \2254_b1 , \2254_b0 , 
		\2255_b1 , \2255_b0 , \2256_b1 , \2256_b0 , \2257_b1 , \2257_b0 , \2258_b1 , \2258_b0 , \2259_b1 , \2259_b0 , 
		\2260_b1 , \2260_b0 , \2261_b1 , \2261_b0 , \2262_b1 , \2262_b0 , \2263_b1 , \2263_b0 , \2264_b1 , \2264_b0 , 
		\2265_b1 , \2265_b0 , \2266_b1 , \2266_b0 , \2267_b1 , \2267_b0 , \2268_b1 , \2268_b0 , \2269_b1 , \2269_b0 , 
		\2270_b1 , \2270_b0 , \2271_b1 , \2271_b0 , \2272_b1 , \2272_b0 , \2273_b1 , \2273_b0 , \2274_b1 , \2274_b0 , 
		\2275_b1 , \2275_b0 , \2276_b1 , \2276_b0 , \2277_b1 , \2277_b0 , \2278_b1 , \2278_b0 , \2279_b1 , \2279_b0 , 
		\2280_b1 , \2280_b0 , \2281_b1 , \2281_b0 , \2282_b1 , \2282_b0 , \2283_b1 , \2283_b0 , \2284_b1 , \2284_b0 , 
		\2285_b1 , \2285_b0 , \2286_b1 , \2286_b0 , \2287_b1 , \2287_b0 , \2288_b1 , \2288_b0 , \2289_b1 , \2289_b0 , 
		\2290_b1 , \2290_b0 , \2291_b1 , \2291_b0 , \2292_b1 , \2292_b0 , \2293_b1 , \2293_b0 , \2294_b1 , \2294_b0 , 
		\2295_b1 , \2295_b0 , \2296_b1 , \2296_b0 , \2297_b1 , \2297_b0 , \2298_b1 , \2298_b0 , \2299_b1 , \2299_b0 , 
		\2300_b1 , \2300_b0 , \2301_b1 , \2301_b0 , \2302_b1 , \2302_b0 , \2303_b1 , \2303_b0 , \2304_b1 , \2304_b0 , 
		\2305_b1 , \2305_b0 , \2306_b1 , \2306_b0 , \2307_b1 , \2307_b0 , \2308_b1 , \2308_b0 , \2309_b1 , \2309_b0 , 
		\2310_b1 , \2310_b0 , \2311_b1 , \2311_b0 , \2312_b1 , \2312_b0 , \2313_b1 , \2313_b0 , \2314_b1 , \2314_b0 , 
		\2315_b1 , \2315_b0 , \2316_b1 , \2316_b0 , \2317_b1 , \2317_b0 , \2318_b1 , \2318_b0 , \2319_b1 , \2319_b0 , 
		\2320_b1 , \2320_b0 , \2321_b1 , \2321_b0 , \2322_b1 , \2322_b0 , \2323_b1 , \2323_b0 , \2324_b1 , \2324_b0 , 
		\2325_b1 , \2325_b0 , \2326_b1 , \2326_b0 , \2327_b1 , \2327_b0 , \2328_b1 , \2328_b0 , \2329_b1 , \2329_b0 , 
		\2330_b1 , \2330_b0 , \2331_b1 , \2331_b0 , \2332_b1 , \2332_b0 , \2333_b1 , \2333_b0 , \2334_b1 , \2334_b0 , 
		\2335_b1 , \2335_b0 , \2336_b1 , \2336_b0 , \2337_b1 , \2337_b0 , \2338_b1 , \2338_b0 , \2339_b1 , \2339_b0 , 
		\2340_b1 , \2340_b0 , \2341_b1 , \2341_b0 , \2342_b1 , \2342_b0 , \2343_b1 , \2343_b0 , \2344_b1 , \2344_b0 , 
		\2345_b1 , \2345_b0 , \2346_b1 , \2346_b0 , \2347_b1 , \2347_b0 , \2348_b1 , \2348_b0 , \2349_b1 , \2349_b0 , 
		\2350_b1 , \2350_b0 , \2351_b1 , \2351_b0 , \2352_b1 , \2352_b0 , \2353_b1 , \2353_b0 , \2354_b1 , \2354_b0 , 
		\2355_b1 , \2355_b0 , \2356_b1 , \2356_b0 , \2357_b1 , \2357_b0 , \2358_b1 , \2358_b0 , \2359_b1 , \2359_b0 , 
		\2360_b1 , \2360_b0 , \2361_b1 , \2361_b0 , \2362_b1 , \2362_b0 , \2363_b1 , \2363_b0 , \2364_b1 , \2364_b0 , 
		\2365_b1 , \2365_b0 , \2366_b1 , \2366_b0 , \2367_b1 , \2367_b0 , \2368_nR126_b1 , \2368_nR126_b0 , \2369_b1 , \2369_b0 , 
		\2370_nR125_b1 , \2370_nR125_b0 , \2371_b1 , \2371_b0 , \2372_b1 , \2372_b0 , \2373_b1 , \2373_b0 , \2374_b1 , \2374_b0 , 
		\2375_b1 , \2375_b0 , \2376_b1 , \2376_b0 , \2377_b1 , \2377_b0 , \2378_b1 , \2378_b0 , \2379_b1 , \2379_b0 , 
		\2380_b1 , \2380_b0 , \2381_b1 , \2381_b0 , \2382_b1 , \2382_b0 , \2383_b1 , \2383_b0 , \2384_b1 , \2384_b0 , 
		\2385_b1 , \2385_b0 , \2386_b1 , \2386_b0 , \2387_b1 , \2387_b0 , \2388_b1 , \2388_b0 , \2389_b1 , \2389_b0 , 
		\2390_b1 , \2390_b0 , \2391_b1 , \2391_b0 , \2392_b1 , \2392_b0 , \2393_b1 , \2393_b0 , \2394_b1 , \2394_b0 , 
		\2395_b1 , \2395_b0 , \2396_b1 , \2396_b0 , \2397_b1 , \2397_b0 , \2398_b1 , \2398_b0 , \2399_b1 , \2399_b0 , 
		\2400_b1 , \2400_b0 , \2401_b1 , \2401_b0 , \2402_b1 , \2402_b0 , \2403_b1 , \2403_b0 , \2404_b1 , \2404_b0 , 
		\2405_b1 , \2405_b0 , \2406_b1 , \2406_b0 , \2407_b1 , \2407_b0 , \2408_b1 , \2408_b0 , \2409_b1 , \2409_b0 , 
		\2410_b1 , \2410_b0 , \2411_b1 , \2411_b0 , \2412_b1 , \2412_b0 , \2413_b1 , \2413_b0 , \2414_b1 , \2414_b0 , 
		\2415_b1 , \2415_b0 , \2416_b1 , \2416_b0 , \2417_b1 , \2417_b0 , \2418_b1 , \2418_b0 , \2419_b1 , \2419_b0 , 
		\2420_b1 , \2420_b0 , \2421_b1 , \2421_b0 , \2422_b1 , \2422_b0 , \2423_b1 , \2423_b0 , \2424_b1 , \2424_b0 , 
		\2425_b1 , \2425_b0 , \2426_b1 , \2426_b0 , \2427_b1 , \2427_b0 , \2428_b1 , \2428_b0 , \2429_b1 , \2429_b0 , 
		\2430_b1 , \2430_b0 , \2431_b1 , \2431_b0 , \2432_b1 , \2432_b0 , \2433_b1 , \2433_b0 , \2434_b1 , \2434_b0 , 
		\2435_b1 , \2435_b0 , \2436_b1 , \2436_b0 , \2437_b1 , \2437_b0 , \2438_b1 , \2438_b0 , \2439_b1 , \2439_b0 , 
		\2440_b1 , \2440_b0 , \2441_b1 , \2441_b0 , \2442_b1 , \2442_b0 , \2443_b1 , \2443_b0 , \2444_b1 , \2444_b0 , 
		\2445_b1 , \2445_b0 , \2446_b1 , \2446_b0 , \2447_b1 , \2447_b0 , \2448_b1 , \2448_b0 , \2449_b1 , \2449_b0 , 
		\2450_b1 , \2450_b0 , \2451_b1 , \2451_b0 , \2452_b1 , \2452_b0 , \2453_b1 , \2453_b0 , \2454_b1 , \2454_b0 , 
		\2455_b1 , \2455_b0 , \2456_b1 , \2456_b0 , \2457_b1 , \2457_b0 , \2458_b1 , \2458_b0 , \2459_b1 , \2459_b0 , 
		\2460_b1 , \2460_b0 , \2461_b1 , \2461_b0 , \2462_b1 , \2462_b0 , \2463_b1 , \2463_b0 , \2464_b1 , \2464_b0 , 
		\2465_b1 , \2465_b0 , \2466_b1 , \2466_b0 , \2467_b1 , \2467_b0 , \2468_b1 , \2468_b0 , \2469_b1 , \2469_b0 , 
		\2470_b1 , \2470_b0 , \2471_b1 , \2471_b0 , \2472_b1 , \2472_b0 , \2473_b1 , \2473_b0 , \2474_b1 , \2474_b0 , 
		\2475_b1 , \2475_b0 , \2476_b1 , \2476_b0 , \2477_b1 , \2477_b0 , \2478_b1 , \2478_b0 , \2479_b1 , \2479_b0 , 
		\2480_b1 , \2480_b0 , \2481_b1 , \2481_b0 , \2482_b1 , \2482_b0 , \2483_b1 , \2483_b0 , \2484_b1 , \2484_b0 , 
		\2485_b1 , \2485_b0 , \2486_b1 , \2486_b0 , \2487_b1 , \2487_b0 , \2488_b1 , \2488_b0 , \2489_b1 , \2489_b0 , 
		\2490_b1 , \2490_b0 , \2491_b1 , \2491_b0 , \2492_b1 , \2492_b0 , \2493_b1 , \2493_b0 , \2494_b1 , \2494_b0 , 
		\2495_b1 , \2495_b0 , \2496_b1 , \2496_b0 , \2497_b1 , \2497_b0 , \2498_b1 , \2498_b0 , \2499_b1 , \2499_b0 , 
		\2500_b1 , \2500_b0 , \2501_b1 , \2501_b0 , \2502_b1 , \2502_b0 , \2503_b1 , \2503_b0 , \2504_b1 , \2504_b0 , 
		\2505_b1 , \2505_b0 , \2506_b1 , \2506_b0 , \2507_b1 , \2507_b0 , \2508_b1 , \2508_b0 , \2509_b1 , \2509_b0 , 
		\2510_b1 , \2510_b0 , \2511_b1 , \2511_b0 , \2512_b1 , \2512_b0 , \2513_b1 , \2513_b0 , \2514_b1 , \2514_b0 , 
		\2515_b1 , \2515_b0 , \2516_b1 , \2516_b0 , \2517_b1 , \2517_b0 , \2518_b1 , \2518_b0 , \2519_b1 , \2519_b0 , 
		\2520_b1 , \2520_b0 , \2521_b1 , \2521_b0 , \2522_b1 , \2522_b0 , \2523_b1 , \2523_b0 , \2524_b1 , \2524_b0 , 
		\2525_b1 , \2525_b0 , \2526_b1 , \2526_b0 , \2527_b1 , \2527_b0 , \2528_b1 , \2528_b0 , \2529_b1 , \2529_b0 , 
		\2530_b1 , \2530_b0 , \2531_b1 , \2531_b0 , \2532_b1 , \2532_b0 , \2533_b1 , \2533_b0 , \2534_b1 , \2534_b0 , 
		\2535_b1 , \2535_b0 , \2536_b1 , \2536_b0 , \2537_b1 , \2537_b0 , \2538_b1 , \2538_b0 , \2539_b1 , \2539_b0 , 
		\2540_b1 , \2540_b0 , \2541_b1 , \2541_b0 , \2542_b1 , \2542_b0 , \2543_b1 , \2543_b0 , \2544_b1 , \2544_b0 , 
		\2545_b1 , \2545_b0 , \2546_b1 , \2546_b0 , \2547_b1 , \2547_b0 , \2548_b1 , \2548_b0 , \2549_b1 , \2549_b0 , 
		\2550_b1 , \2550_b0 , \2551_b1 , \2551_b0 , \2552_b1 , \2552_b0 , \2553_b1 , \2553_b0 , \2554_b1 , \2554_b0 , 
		\2555_b1 , \2555_b0 , \2556_b1 , \2556_b0 , \2557_b1 , \2557_b0 , \2558_b1 , \2558_b0 , \2559_b1 , \2559_b0 , 
		\2560_b1 , \2560_b0 , \2561_b1 , \2561_b0 , \2562_b1 , \2562_b0 , \2563_b1 , \2563_b0 , \2564_b1 , \2564_b0 , 
		\2565_b1 , \2565_b0 , \2566_b1 , \2566_b0 , \2567_b1 , \2567_b0 , \2568_b1 , \2568_b0 , \2569_b1 , \2569_b0 , 
		\2570_b1 , \2570_b0 , \2571_b1 , \2571_b0 , \2572_b1 , \2572_b0 , \2573_b1 , \2573_b0 , \2574_b1 , \2574_b0 , 
		\2575_b1 , \2575_b0 , \2576_b1 , \2576_b0 , \2577_b1 , \2577_b0 , \2578_b1 , \2578_b0 , \2579_b1 , \2579_b0 , 
		\2580_b1 , \2580_b0 , \2581_b1 , \2581_b0 , \2582_b1 , \2582_b0 , \2583_b1 , \2583_b0 , \2584_b1 , \2584_b0 , 
		\2585_b1 , \2585_b0 , \2586_b1 , \2586_b0 , \2587_b1 , \2587_b0 , \2588_b1 , \2588_b0 , \2589_b1 , \2589_b0 , 
		\2590_b1 , \2590_b0 , \2591_b1 , \2591_b0 , \2592_b1 , \2592_b0 , \2593_b1 , \2593_b0 , \2594_b1 , \2594_b0 , 
		\2595_b1 , \2595_b0 , \2596_b1 , \2596_b0 , \2597_b1 , \2597_b0 , \2598_b1 , \2598_b0 , \2599_b1 , \2599_b0 , 
		\2600_b1 , \2600_b0 , \2601_b1 , \2601_b0 , \2602_b1 , \2602_b0 , \2603_b1 , \2603_b0 , \2604_b1 , \2604_b0 , 
		\2605_b1 , \2605_b0 , \2606_b1 , \2606_b0 , \2607_b1 , \2607_b0 , \2608_b1 , \2608_b0 , \2609_b1 , \2609_b0 , 
		\2610_b1 , \2610_b0 , \2611_b1 , \2611_b0 , \2612_b1 , \2612_b0 , \2613_b1 , \2613_b0 , \2614_b1 , \2614_b0 , 
		\2615_b1 , \2615_b0 , \2616_b1 , \2616_b0 , \2617_b1 , \2617_b0 , \2618_b1 , \2618_b0 , \2619_b1 , \2619_b0 , 
		\2620_b1 , \2620_b0 , \2621_b1 , \2621_b0 , \2622_b1 , \2622_b0 , \2623_b1 , \2623_b0 , \2624_b1 , \2624_b0 , 
		\2625_b1 , \2625_b0 , \2626_b1 , \2626_b0 , \2627_b1 , \2627_b0 , \2628_b1 , \2628_b0 , \2629_b1 , \2629_b0 , 
		\2630_b1 , \2630_b0 , \2631_b1 , \2631_b0 , \2632_b1 , \2632_b0 , \2633_b1 , \2633_b0 , \2634_b1 , \2634_b0 , 
		\2635_b1 , \2635_b0 , \2636_b1 , \2636_b0 , \2637_b1 , \2637_b0 , \2638_b1 , \2638_b0 , \2639_b1 , \2639_b0 , 
		\2640_b1 , \2640_b0 , \2641_b1 , \2641_b0 , \2642_b1 , \2642_b0 , \2643_b1 , \2643_b0 , \2644_b1 , \2644_b0 , 
		\2645_b1 , \2645_b0 , \2646_b1 , \2646_b0 , \2647_b1 , \2647_b0 , \2648_b1 , \2648_b0 , \2649_b1 , \2649_b0 , 
		\2650_b1 , \2650_b0 , \2651_b1 , \2651_b0 , \2652_b1 , \2652_b0 , \2653_b1 , \2653_b0 , \2654_b1 , \2654_b0 , 
		\2655_b1 , \2655_b0 , \2656_b1 , \2656_b0 , \2657_b1 , \2657_b0 , \2658_b1 , \2658_b0 , \2659_b1 , \2659_b0 , 
		\2660_b1 , \2660_b0 , \2661_b1 , \2661_b0 , \2662_b1 , \2662_b0 , \2663_b1 , \2663_b0 , \2664_b1 , \2664_b0 , 
		\2665_b1 , \2665_b0 , \2666_b1 , \2666_b0 , \2667_b1 , \2667_b0 , \2668_b1 , \2668_b0 , \2669_b1 , \2669_b0 , 
		\2670_b1 , \2670_b0 , \2671_b1 , \2671_b0 , \2672_b1 , \2672_b0 , \2673_b1 , \2673_b0 , \2674_b1 , \2674_b0 , 
		\2675_b1 , \2675_b0 , \2676_b1 , \2676_b0 , \2677_b1 , \2677_b0 , \2678_b1 , \2678_b0 , \2679_b1 , \2679_b0 , 
		\2680_b1 , \2680_b0 , \2681_b1 , \2681_b0 , \2682_b1 , \2682_b0 , \2683_b1 , \2683_b0 , \2684_b1 , \2684_b0 , 
		\2685_b1 , \2685_b0 , \2686_b1 , \2686_b0 , \2687_b1 , \2687_b0 , \2688_b1 , \2688_b0 , \2689_b1 , \2689_b0 , 
		\2690_b1 , \2690_b0 , \2691_b1 , \2691_b0 , \2692_b1 , \2692_b0 , \2693_b1 , \2693_b0 , \2694_b1 , \2694_b0 , 
		\2695_b1 , \2695_b0 , \2696_b1 , \2696_b0 , \2697_b1 , \2697_b0 , \2698_b1 , \2698_b0 , \2699_b1 , \2699_b0 , 
		\2700_b1 , \2700_b0 , \2701_b1 , \2701_b0 , \2702_b1 , \2702_b0 , \2703_b1 , \2703_b0 , \2704_b1 , \2704_b0 , 
		\2705_b1 , \2705_b0 , \2706_b1 , \2706_b0 , \2707_b1 , \2707_b0 , \2708_b1 , \2708_b0 , \2709_b1 , \2709_b0 , 
		\2710_b1 , \2710_b0 , \2711_b1 , \2711_b0 , \2712_b1 , \2712_b0 , \2713_b1 , \2713_b0 , \2714_b1 , \2714_b0 , 
		\2715_b1 , \2715_b0 , \2716_b1 , \2716_b0 , \2717_b1 , \2717_b0 , \2718_b1 , \2718_b0 , \2719_b1 , \2719_b0 , 
		\2720_b1 , \2720_b0 , \2721_b1 , \2721_b0 , \2722_b1 , \2722_b0 , \2723_b1 , \2723_b0 , \2724_b1 , \2724_b0 , 
		\2725_b1 , \2725_b0 , \2726_b1 , \2726_b0 , \2727_b1 , \2727_b0 , \2728_b1 , \2728_b0 , \2729_b1 , \2729_b0 , 
		\2730_b1 , \2730_b0 , \2731_b1 , \2731_b0 , \2732_b1 , \2732_b0 , \2733_b1 , \2733_b0 , \2734_b1 , \2734_b0 , 
		\2735_b1 , \2735_b0 , \2736_b1 , \2736_b0 , \2737_b1 , \2737_b0 , \2738_b1 , \2738_b0 , \2739_b1 , \2739_b0 , 
		\2740_b1 , \2740_b0 , \2741_b1 , \2741_b0 , \2742_b1 , \2742_b0 , \2743_b1 , \2743_b0 , \2744_b1 , \2744_b0 , 
		\2745_b1 , \2745_b0 , \2746_b1 , \2746_b0 , \2747_b1 , \2747_b0 , \2748_b1 , \2748_b0 , \2749_b1 , \2749_b0 , 
		\2750_b1 , \2750_b0 , \2751_b1 , \2751_b0 , \2752_b1 , \2752_b0 , \2753_b1 , \2753_b0 , \2754_b1 , \2754_b0 , 
		\2755_b1 , \2755_b0 , \2756_b1 , \2756_b0 , \2757_b1 , \2757_b0 , \2758_b1 , \2758_b0 , \2759_b1 , \2759_b0 , 
		\2760_b1 , \2760_b0 , \2761_b1 , \2761_b0 , \2762_b1 , \2762_b0 , \2763_b1 , \2763_b0 , \2764_b1 , \2764_b0 , 
		\2765_b1 , \2765_b0 , \2766_b1 , \2766_b0 , \2767_b1 , \2767_b0 , \2768_b1 , \2768_b0 , \2769_b1 , \2769_b0 , 
		\2770_b1 , \2770_b0 , \2771_b1 , \2771_b0 , \2772_b1 , \2772_b0 , \2773_b1 , \2773_b0 , \2774_b1 , \2774_b0 , 
		\2775_b1 , \2775_b0 , \2776_b1 , \2776_b0 , \2777_b1 , \2777_b0 , \2778_b1 , \2778_b0 , \2779_b1 , \2779_b0 , 
		\2780_b1 , \2780_b0 , \2781_b1 , \2781_b0 , \2782_b1 , \2782_b0 , \2783_b1 , \2783_b0 , \2784_b1 , \2784_b0 , 
		\2785_b1 , \2785_b0 , \2786_b1 , \2786_b0 , \2787_b1 , \2787_b0 , \2788_b1 , \2788_b0 , \2789_b1 , \2789_b0 , 
		\2790_b1 , \2790_b0 , \2791_b1 , \2791_b0 , \2792_b1 , \2792_b0 , \2793_b1 , \2793_b0 , \2794_b1 , \2794_b0 , 
		\2795_b1 , \2795_b0 , \2796_b1 , \2796_b0 , \2797_b1 , \2797_b0 , \2798_b1 , \2798_b0 , \2799_b1 , \2799_b0 , 
		\2800_b1 , \2800_b0 , \2801_b1 , \2801_b0 , \2802_b1 , \2802_b0 , \2803_b1 , \2803_b0 , \2804_b1 , \2804_b0 , 
		\2805_b1 , \2805_b0 , \2806_b1 , \2806_b0 , \2807_b1 , \2807_b0 , \2808_b1 , \2808_b0 , \2809_b1 , \2809_b0 , 
		\2810_b1 , \2810_b0 , \2811_b1 , \2811_b0 , \2812_b1 , \2812_b0 , \2813_b1 , \2813_b0 , \2814_b1 , \2814_b0 , 
		\2815_b1 , \2815_b0 , \2816_b1 , \2816_b0 , \2817_b1 , \2817_b0 , \2818_b1 , \2818_b0 , \2819_b1 , \2819_b0 , 
		\2820_b1 , \2820_b0 , \2821_b1 , \2821_b0 , \2822_b1 , \2822_b0 , \2823_b1 , \2823_b0 , \2824_b1 , \2824_b0 , 
		\2825_b1 , \2825_b0 , \2826_b1 , \2826_b0 , \2827_b1 , \2827_b0 , \2828_b1 , \2828_b0 , \2829_b1 , \2829_b0 , 
		\2830_b1 , \2830_b0 , \2831_b1 , \2831_b0 , \2832_b1 , \2832_b0 , \2833_b1 , \2833_b0 , \2834_b1 , \2834_b0 , 
		\2835_b1 , \2835_b0 , \2836_b1 , \2836_b0 , \2837_b1 , \2837_b0 , \2838_b1 , \2838_b0 , \2839_b1 , \2839_b0 , 
		\2840_b1 , \2840_b0 , \2841_b1 , \2841_b0 , \2842_b1 , \2842_b0 , \2843_b1 , \2843_b0 , \2844_b1 , \2844_b0 , 
		\2845_b1 , \2845_b0 , \2846_b1 , \2846_b0 , \2847_b1 , \2847_b0 , \2848_b1 , \2848_b0 , \2849_b1 , \2849_b0 , 
		\2850_b1 , \2850_b0 , \2851_b1 , \2851_b0 , \2852_b1 , \2852_b0 , \2853_b1 , \2853_b0 , \2854_b1 , \2854_b0 , 
		\2855_b1 , \2855_b0 , \2856_b1 , \2856_b0 , \2857_b1 , \2857_b0 , \2858_b1 , \2858_b0 , \2859_b1 , \2859_b0 , 
		\2860_b1 , \2860_b0 , \2861_b1 , \2861_b0 , \2862_b1 , \2862_b0 , \2863_b1 , \2863_b0 , \2864_b1 , \2864_b0 , 
		\2865_b1 , \2865_b0 , \2866_b1 , \2866_b0 , \2867_b1 , \2867_b0 , \2868_b1 , \2868_b0 , \2869_b1 , \2869_b0 , 
		\2870_b1 , \2870_b0 , \2871_b1 , \2871_b0 , \2872_b1 , \2872_b0 , \2873_b1 , \2873_b0 , \2874_b1 , \2874_b0 , 
		\2875_b1 , \2875_b0 , \2876_b1 , \2876_b0 , \2877_b1 , \2877_b0 , \2878_b1 , \2878_b0 , \2879_b1 , \2879_b0 , 
		\2880_b1 , \2880_b0 , \2881_b1 , \2881_b0 , \2882_b1 , \2882_b0 , \2883_b1 , \2883_b0 , \2884_b1 , \2884_b0 , 
		\2885_b1 , \2885_b0 , \2886_b1 , \2886_b0 , \2887_b1 , \2887_b0 , \2888_b1 , \2888_b0 , \2889_b1 , \2889_b0 , 
		\2890_b1 , \2890_b0 , \2891_b1 , \2891_b0 , \2892_b1 , \2892_b0 , \2893_b1 , \2893_b0 , \2894_b1 , \2894_b0 , 
		\2895_b1 , \2895_b0 , \2896_b1 , \2896_b0 , \2897_b1 , \2897_b0 , \2898_b1 , \2898_b0 , \2899_b1 , \2899_b0 , 
		\2900_b1 , \2900_b0 , \2901_b1 , \2901_b0 , \2902_b1 , \2902_b0 , \2903_b1 , \2903_b0 , \2904_b1 , \2904_b0 , 
		\2905_b1 , \2905_b0 , \2906_b1 , \2906_b0 , \2907_b1 , \2907_b0 , \2908_b1 , \2908_b0 , \2909_nR123_b1 , \2909_nR123_b0 , 
		\2910_b1 , \2910_b0 , \2911_b1 , \2911_b0 , \2912_b1 , \2912_b0 , \2913_b1 , \2913_b0 , \2914_b1 , \2914_b0 , 
		\2915_b1 , \2915_b0 , \2916_b1 , \2916_b0 , \2917_b1 , \2917_b0 , \2918_b1 , \2918_b0 , \2919_b1 , \2919_b0 , 
		\2920_b1 , \2920_b0 , \2921_b1 , \2921_b0 , \2922_b1 , \2922_b0 , \2923_b1 , \2923_b0 , \2924_b1 , \2924_b0 , 
		\2925_b1 , \2925_b0 , \2926_b1 , \2926_b0 , \2927_b1 , \2927_b0 , \2928_b1 , \2928_b0 , \2929_b1 , \2929_b0 , 
		\2930_b1 , \2930_b0 , \2931_b1 , \2931_b0 , \2932_b1 , \2932_b0 , \2933_b1 , \2933_b0 , \2934_b1 , \2934_b0 , 
		\2935_b1 , \2935_b0 , \2936_b1 , \2936_b0 , \2937_b1 , \2937_b0 , \2938_b1 , \2938_b0 , \2939_b1 , \2939_b0 , 
		\2940_b1 , \2940_b0 , \2941_b1 , \2941_b0 , \2942_b1 , \2942_b0 , \2943_b1 , \2943_b0 , \2944_b1 , \2944_b0 , 
		\2945_b1 , \2945_b0 , \2946_b1 , \2946_b0 , \2947_b1 , \2947_b0 , \2948_b1 , \2948_b0 , \2949_b1 , \2949_b0 , 
		\2950_b1 , \2950_b0 , \2951_b1 , \2951_b0 , \2952_b1 , \2952_b0 , \2953_b1 , \2953_b0 , \2954_b1 , \2954_b0 , 
		\2955_b1 , \2955_b0 , \2956_b1 , \2956_b0 , \2957_b1 , \2957_b0 , \2958_b1 , \2958_b0 , \2959_b1 , \2959_b0 , 
		\2960_b1 , \2960_b0 , \2961_b1 , \2961_b0 , \2962_b1 , \2962_b0 , \2963_b1 , \2963_b0 , \2964_b1 , \2964_b0 , 
		\2965_b1 , \2965_b0 , \2966_b1 , \2966_b0 , \2967_b1 , \2967_b0 , \2968_b1 , \2968_b0 , \2969_b1 , \2969_b0 , 
		\2970_b1 , \2970_b0 , \2971_b1 , \2971_b0 , \2972_b1 , \2972_b0 , \2973_b1 , \2973_b0 , \2974_b1 , \2974_b0 , 
		\2975_b1 , \2975_b0 , \2976_b1 , \2976_b0 , \2977_b1 , \2977_b0 , \2978_b1 , \2978_b0 , \2979_b1 , \2979_b0 , 
		\2980_b1 , \2980_b0 , \2981_b1 , \2981_b0 , \2982_b1 , \2982_b0 , \2983_b1 , \2983_b0 , \2984_b1 , \2984_b0 , 
		\2985_b1 , \2985_b0 , \2986_b1 , \2986_b0 , \2987_b1 , \2987_b0 , \2988_b1 , \2988_b0 , \2989_b1 , \2989_b0 , 
		\2990_b1 , \2990_b0 , \2991_b1 , \2991_b0 , \2992_b1 , \2992_b0 , \2993_b1 , \2993_b0 , \2994_b1 , \2994_b0 , 
		\2995_b1 , \2995_b0 , \2996_b1 , \2996_b0 , \2997_b1 , \2997_b0 , \2998_b1 , \2998_b0 , \2999_b1 , \2999_b0 , 
		\3000_b1 , \3000_b0 , \3001_b1 , \3001_b0 , \3002_b1 , \3002_b0 , \3003_b1 , \3003_b0 , \3004_b1 , \3004_b0 , 
		\3005_b1 , \3005_b0 , \3006_b1 , \3006_b0 , \3007_b1 , \3007_b0 , \3008_b1 , \3008_b0 , \3009_b1 , \3009_b0 , 
		\3010_b1 , \3010_b0 , \3011_b1 , \3011_b0 , \3012_b1 , \3012_b0 , \3013_b1 , \3013_b0 , \3014_b1 , \3014_b0 , 
		\3015_b1 , \3015_b0 , \3016_b1 , \3016_b0 , \3017_b1 , \3017_b0 , \3018_b1 , \3018_b0 , \3019_b1 , \3019_b0 , 
		\3020_b1 , \3020_b0 , \3021_b1 , \3021_b0 , \3022_b1 , \3022_b0 , \3023_b1 , \3023_b0 , \3024_b1 , \3024_b0 , 
		\3025_b1 , \3025_b0 , \3026_b1 , \3026_b0 , \3027_b1 , \3027_b0 , \3028_b1 , \3028_b0 , \3029_b1 , \3029_b0 , 
		\3030_b1 , \3030_b0 , \3031_b1 , \3031_b0 , \3032_b1 , \3032_b0 , \3033_b1 , \3033_b0 , \3034_b1 , \3034_b0 , 
		\3035_b1 , \3035_b0 , \3036_b1 , \3036_b0 , \3037_b1 , \3037_b0 , \3038_b1 , \3038_b0 , \3039_b1 , \3039_b0 , 
		\3040_b1 , \3040_b0 , \3041_b1 , \3041_b0 , \3042_b1 , \3042_b0 , \3043_b1 , \3043_b0 , \3044_b1 , \3044_b0 , 
		\3045_b1 , \3045_b0 , \3046_b1 , \3046_b0 , \3047_b1 , \3047_b0 , \3048_b1 , \3048_b0 , \3049_b1 , \3049_b0 , 
		\3050_b1 , \3050_b0 , \3051_b1 , \3051_b0 , \3052_b1 , \3052_b0 , \3053_b1 , \3053_b0 , \3054_b1 , \3054_b0 , 
		\3055_b1 , \3055_b0 , \3056_b1 , \3056_b0 , \3057_b1 , \3057_b0 , \3058_b1 , \3058_b0 , \3059_b1 , \3059_b0 , 
		\3060_b1 , \3060_b0 , \3061_b1 , \3061_b0 , \3062_b1 , \3062_b0 , \3063_b1 , \3063_b0 , \3064_b1 , \3064_b0 , 
		\3065_b1 , \3065_b0 , \3066_b1 , \3066_b0 , \3067_b1 , \3067_b0 , \3068_b1 , \3068_b0 , \3069_b1 , \3069_b0 , 
		\3070_b1 , \3070_b0 , \3071_b1 , \3071_b0 , \3072_b1 , \3072_b0 , \3073_b1 , \3073_b0 , \3074_b1 , \3074_b0 , 
		\3075_b1 , \3075_b0 , \3076_b1 , \3076_b0 , \3077_b1 , \3077_b0 , \3078_b1 , \3078_b0 , \3079_b1 , \3079_b0 , 
		\3080_b1 , \3080_b0 , \3081_b1 , \3081_b0 , \3082_b1 , \3082_b0 , \3083_b1 , \3083_b0 , \3084_b1 , \3084_b0 , 
		\3085_b1 , \3085_b0 , \3086_b1 , \3086_b0 , \3087_b1 , \3087_b0 , \3088_b1 , \3088_b0 , \3089_b1 , \3089_b0 , 
		\3090_b1 , \3090_b0 , \3091_b1 , \3091_b0 , \3092_b1 , \3092_b0 , \3093_b1 , \3093_b0 , \3094_b1 , \3094_b0 , 
		\3095_b1 , \3095_b0 , \3096_b1 , \3096_b0 , \3097_b1 , \3097_b0 , \3098_b1 , \3098_b0 , \3099_b1 , \3099_b0 , 
		\3100_b1 , \3100_b0 , \3101_b1 , \3101_b0 , \3102_b1 , \3102_b0 , \3103_b1 , \3103_b0 , \3104_b1 , \3104_b0 , 
		\3105_b1 , \3105_b0 , \3106_b1 , \3106_b0 , \3107_b1 , \3107_b0 , \3108_b1 , \3108_b0 , \3109_b1 , \3109_b0 , 
		\3110_b1 , \3110_b0 , \3111_b1 , \3111_b0 , \3112_b1 , \3112_b0 , \3113_b1 , \3113_b0 , \3114_b1 , \3114_b0 , 
		\3115_b1 , \3115_b0 , \3116_b1 , \3116_b0 , \3117_b1 , \3117_b0 , \3118_b1 , \3118_b0 , \3119_b1 , \3119_b0 , 
		\3120_b1 , \3120_b0 , \3121_b1 , \3121_b0 , \3122_b1 , \3122_b0 , \3123_b1 , \3123_b0 , \3124_b1 , \3124_b0 , 
		\3125_b1 , \3125_b0 , \3126_b1 , \3126_b0 , \3127_b1 , \3127_b0 , \3128_b1 , \3128_b0 , \3129_b1 , \3129_b0 , 
		\3130_b1 , \3130_b0 , \3131_b1 , \3131_b0 , \3132_b1 , \3132_b0 , \3133_b1 , \3133_b0 , \3134_b1 , \3134_b0 , 
		\3135_b1 , \3135_b0 , \3136_b1 , \3136_b0 , \3137_b1 , \3137_b0 , \3138_b1 , \3138_b0 , \3139_b1 , \3139_b0 , 
		\3140_b1 , \3140_b0 , \3141_b1 , \3141_b0 , \3142_b1 , \3142_b0 , \3143_b1 , \3143_b0 , \3144_b1 , \3144_b0 , 
		\3145_b1 , \3145_b0 , \3146_b1 , \3146_b0 , \3147_b1 , \3147_b0 , \3148_b1 , \3148_b0 , \3149_b1 , \3149_b0 , 
		\3150_b1 , \3150_b0 , \3151_b1 , \3151_b0 , \3152_b1 , \3152_b0 , \3153_b1 , \3153_b0 , \3154_b1 , \3154_b0 , 
		\3155_b1 , \3155_b0 , \3156_b1 , \3156_b0 , \3157_b1 , \3157_b0 , \3158_b1 , \3158_b0 , \3159_b1 , \3159_b0 , 
		\3160_b1 , \3160_b0 , \3161_b1 , \3161_b0 , \3162_b1 , \3162_b0 , \3163_b1 , \3163_b0 , \3164_b1 , \3164_b0 , 
		\3165_b1 , \3165_b0 , \3166_b1 , \3166_b0 , \3167_b1 , \3167_b0 , \3168_b1 , \3168_b0 , \3169_b1 , \3169_b0 , 
		\3170_b1 , \3170_b0 , \3171_b1 , \3171_b0 , \3172_b1 , \3172_b0 , \3173_b1 , \3173_b0 , \3174_b1 , \3174_b0 , 
		\3175_b1 , \3175_b0 , \3176_b1 , \3176_b0 , \3177_b1 , \3177_b0 , \3178_b1 , \3178_b0 , \3179_b1 , \3179_b0 , 
		\3180_b1 , \3180_b0 , \3181_b1 , \3181_b0 , \3182_b1 , \3182_b0 , \3183_b1 , \3183_b0 , \3184_b1 , \3184_b0 , 
		\3185_b1 , \3185_b0 , \3186_b1 , \3186_b0 , \3187_b1 , \3187_b0 , \3188_b1 , \3188_b0 , \3189_b1 , \3189_b0 , 
		\3190_b1 , \3190_b0 , \3191_b1 , \3191_b0 , \3192_b1 , \3192_b0 , \3193_b1 , \3193_b0 , \3194_b1 , \3194_b0 , 
		\3195_b1 , \3195_b0 , \3196_b1 , \3196_b0 , \3197_b1 , \3197_b0 , \3198_b1 , \3198_b0 , \3199_b1 , \3199_b0 , 
		\3200_b1 , \3200_b0 , \3201_b1 , \3201_b0 , \3202_b1 , \3202_b0 , \3203_b1 , \3203_b0 , \3204_b1 , \3204_b0 , 
		\3205_b1 , \3205_b0 , \3206_b1 , \3206_b0 , \3207_b1 , \3207_b0 , \3208_b1 , \3208_b0 , \3209_b1 , \3209_b0 , 
		\3210_b1 , \3210_b0 , \3211_b1 , \3211_b0 , \3212_b1 , \3212_b0 , \3213_b1 , \3213_b0 , \3214_b1 , \3214_b0 , 
		\3215_b1 , \3215_b0 , \3216_b1 , \3216_b0 , \3217_b1 , \3217_b0 , \3218_b1 , \3218_b0 , \3219_b1 , \3219_b0 , 
		\3220_b1 , \3220_b0 , \3221_b1 , \3221_b0 , \3222_b1 , \3222_b0 , \3223_b1 , \3223_b0 , \3224_b1 , \3224_b0 , 
		\3225_b1 , \3225_b0 , \3226_b1 , \3226_b0 , \3227_b1 , \3227_b0 , \3228_b1 , \3228_b0 , \3229_b1 , \3229_b0 , 
		\3230_b1 , \3230_b0 , \3231_b1 , \3231_b0 , \3232_b1 , \3232_b0 , \3233_b1 , \3233_b0 , \3234_b1 , \3234_b0 , 
		\3235_b1 , \3235_b0 , \3236_b1 , \3236_b0 , \3237_b1 , \3237_b0 , \3238_b1 , \3238_b0 , \3239_b1 , \3239_b0 , 
		\3240_b1 , \3240_b0 , \3241_b1 , \3241_b0 , \3242_b1 , \3242_b0 , \3243_b1 , \3243_b0 , \3244_b1 , \3244_b0 , 
		\3245_b1 , \3245_b0 , \3246_b1 , \3246_b0 , \3247_b1 , \3247_b0 , \3248_b1 , \3248_b0 , \3249_b1 , \3249_b0 , 
		\3250_b1 , \3250_b0 , \3251_b1 , \3251_b0 , \3252_b1 , \3252_b0 , \3253_b1 , \3253_b0 , \3254_b1 , \3254_b0 , 
		\3255_b1 , \3255_b0 , \3256_b1 , \3256_b0 , \3257_b1 , \3257_b0 , \3258_b1 , \3258_b0 , \3259_b1 , \3259_b0 , 
		\3260_b1 , \3260_b0 , \3261_b1 , \3261_b0 , \3262_b1 , \3262_b0 , \3263_b1 , \3263_b0 , \3264_b1 , \3264_b0 , 
		\3265_b1 , \3265_b0 , \3266_b1 , \3266_b0 , \3267_b1 , \3267_b0 , \3268_b1 , \3268_b0 , \3269_b1 , \3269_b0 , 
		\3270_b1 , \3270_b0 , \3271_b1 , \3271_b0 , \3272_b1 , \3272_b0 , \3273_b1 , \3273_b0 , \3274_b1 , \3274_b0 , 
		\3275_b1 , \3275_b0 , \3276_b1 , \3276_b0 , \3277_b1 , \3277_b0 , \3278_b1 , \3278_b0 , \3279_b1 , \3279_b0 , 
		\3280_b1 , \3280_b0 , \3281_b1 , \3281_b0 , \3282_b1 , \3282_b0 , \3283_b1 , \3283_b0 , \3284_b1 , \3284_b0 , 
		\3285_b1 , \3285_b0 , \3286_b1 , \3286_b0 , \3287_b1 , \3287_b0 , \3288_b1 , \3288_b0 , \3289_b1 , \3289_b0 , 
		\3290_b1 , \3290_b0 , \3291_b1 , \3291_b0 , \3292_b1 , \3292_b0 , \3293_b1 , \3293_b0 , \3294_b1 , \3294_b0 , 
		\3295_b1 , \3295_b0 , \3296_b1 , \3296_b0 , \3297_b1 , \3297_b0 , \3298_b1 , \3298_b0 , \3299_b1 , \3299_b0 , 
		\3300_b1 , \3300_b0 , \3301_b1 , \3301_b0 , \3302_b1 , \3302_b0 , \3303_b1 , \3303_b0 , \3304_b1 , \3304_b0 , 
		\3305_b1 , \3305_b0 , \3306_b1 , \3306_b0 , \3307_b1 , \3307_b0 , \3308_b1 , \3308_b0 , \3309_b1 , \3309_b0 , 
		\3310_b1 , \3310_b0 , \3311_b1 , \3311_b0 , \3312_b1 , \3312_b0 , \3313_b1 , \3313_b0 , \3314_b1 , \3314_b0 , 
		\3315_b1 , \3315_b0 , \3316_b1 , \3316_b0 , \3317_b1 , \3317_b0 , \3318_b1 , \3318_b0 , \3319_b1 , \3319_b0 , 
		\3320_b1 , \3320_b0 , \3321_b1 , \3321_b0 , \3322_b1 , \3322_b0 , \3323_b1 , \3323_b0 , \3324_b1 , \3324_b0 , 
		\3325_b1 , \3325_b0 , \3326_b1 , \3326_b0 , \3327_b1 , \3327_b0 , \3328_b1 , \3328_b0 , \3329_b1 , \3329_b0 , 
		\3330_b1 , \3330_b0 , \3331_b1 , \3331_b0 , \3332_b1 , \3332_b0 , \3333_b1 , \3333_b0 , \3334_b1 , \3334_b0 , 
		\3335_b1 , \3335_b0 , \3336_b1 , \3336_b0 , \3337_b1 , \3337_b0 , \3338_b1 , \3338_b0 , \3339_b1 , \3339_b0 , 
		\3340_b1 , \3340_b0 , \3341_b1 , \3341_b0 , \3342_b1 , \3342_b0 , \3343_b1 , \3343_b0 , \3344_b1 , \3344_b0 , 
		\3345_b1 , \3345_b0 , \3346_b1 , \3346_b0 , \3347_b1 , \3347_b0 , \3348_b1 , \3348_b0 , \3349_b1 , \3349_b0 , 
		\3350_b1 , \3350_b0 , \3351_b1 , \3351_b0 , \3352_b1 , \3352_b0 , \3353_b1 , \3353_b0 , \3354_b1 , \3354_b0 , 
		\3355_b1 , \3355_b0 , \3356_b1 , \3356_b0 , \3357_b1 , \3357_b0 , \3358_b1 , \3358_b0 , \3359_b1 , \3359_b0 , 
		\3360_b1 , \3360_b0 , \3361_b1 , \3361_b0 , \3362_b1 , \3362_b0 , \3363_b1 , \3363_b0 , \3364_b1 , \3364_b0 , 
		\3365_b1 , \3365_b0 , \3366_b1 , \3366_b0 , \3367_b1 , \3367_b0 , \3368_b1 , \3368_b0 , \3369_b1 , \3369_b0 , 
		\3370_b1 , \3370_b0 , \3371_b1 , \3371_b0 , \3372_b1 , \3372_b0 , \3373_b1 , \3373_b0 , \3374_b1 , \3374_b0 , 
		\3375_b1 , \3375_b0 , \3376_b1 , \3376_b0 , \3377_b1 , \3377_b0 , \3378_b1 , \3378_b0 , \3379_b1 , \3379_b0 , 
		\3380_b1 , \3380_b0 , \3381_b1 , \3381_b0 , \3382_b1 , \3382_b0 , \3383_b1 , \3383_b0 , \3384_b1 , \3384_b0 , 
		\3385_b1 , \3385_b0 , \3386_b1 , \3386_b0 , \3387_b1 , \3387_b0 , \3388_b1 , \3388_b0 , \3389_b1 , \3389_b0 , 
		\3390_b1 , \3390_b0 , \3391_b1 , \3391_b0 , \3392_b1 , \3392_b0 , \3393_b1 , \3393_b0 , \3394_b1 , \3394_b0 , 
		\3395_b1 , \3395_b0 , \3396_b1 , \3396_b0 , \3397_b1 , \3397_b0 , \3398_b1 , \3398_b0 , \3399_b1 , \3399_b0 , 
		\3400_b1 , \3400_b0 , \3401_b1 , \3401_b0 , \3402_b1 , \3402_b0 , \3403_b1 , \3403_b0 , \3404_b1 , \3404_b0 , 
		\3405_b1 , \3405_b0 , \3406_b1 , \3406_b0 , \3407_b1 , \3407_b0 , \3408_b1 , \3408_b0 , \3409_b1 , \3409_b0 , 
		\3410_b1 , \3410_b0 , \3411_b1 , \3411_b0 , \3412_b1 , \3412_b0 , \3413_b1 , \3413_b0 , \3414_b1 , \3414_b0 , 
		\3415_b1 , \3415_b0 , \3416_b1 , \3416_b0 , \3417_b1 , \3417_b0 , \3418_b1 , \3418_b0 , \3419_b1 , \3419_b0 , 
		\3420_b1 , \3420_b0 , \3421_b1 , \3421_b0 , \3422_b1 , \3422_b0 , \3423_b1 , \3423_b0 , \3424_b1 , \3424_b0 , 
		\3425_b1 , \3425_b0 , \3426_b1 , \3426_b0 , \3427_b1 , \3427_b0 , \3428_b1 , \3428_b0 , \3429_b1 , \3429_b0 , 
		\3430_b1 , \3430_b0 , \3431_b1 , \3431_b0 , \3432_b1 , \3432_b0 , \3433_b1 , \3433_b0 , \3434_b1 , \3434_b0 , 
		\3435_b1 , \3435_b0 , \3436_b1 , \3436_b0 , \3437_b1 , \3437_b0 , \3438_b1 , \3438_b0 , \3439_b1 , \3439_b0 , 
		\3440_b1 , \3440_b0 , \3441_b1 , \3441_b0 , \3442_b1 , \3442_b0 , \3443_b1 , \3443_b0 , \3444_b1 , \3444_b0 , 
		\3445_b1 , \3445_b0 , \3446_b1 , \3446_b0 , \3447_b1 , \3447_b0 , \3448_b1 , \3448_b0 , \3449_b1 , \3449_b0 , 
		\3450_b1 , \3450_b0 , \3451_b1 , \3451_b0 , \3452_b1 , \3452_b0 , \3453_b1 , \3453_b0 , \3454_b1 , \3454_b0 , 
		\3455_b1 , \3455_b0 , \3456_b1 , \3456_b0 , \3457_b1 , \3457_b0 , \3458_b1 , \3458_b0 , \3459_b1 , \3459_b0 , 
		\3460_b1 , \3460_b0 , \3461_b1 , \3461_b0 , \3462_b1 , \3462_b0 , \3463_b1 , \3463_b0 , \3464_b1 , \3464_b0 , 
		\3465_b1 , \3465_b0 , \3466_b1 , \3466_b0 , \3467_b1 , \3467_b0 , \3468_b1 , \3468_b0 , \3469_b1 , \3469_b0 , 
		\3470_b1 , \3470_b0 , \3471_b1 , \3471_b0 , \3472_b1 , \3472_b0 , \3473_b1 , \3473_b0 , \3474_b1 , \3474_b0 , 
		\3475_b1 , \3475_b0 , \3476_b1 , \3476_b0 , \3477_b1 , \3477_b0 , \3478_b1 , \3478_b0 , \3479_b1 , \3479_b0 , 
		\3480_b1 , \3480_b0 , \3481_b1 , \3481_b0 , \3482_b1 , \3482_b0 , \3483_b1 , \3483_b0 , \3484_b1 , \3484_b0 , 
		\3485_b1 , \3485_b0 , \3486_b1 , \3486_b0 , \3487_b1 , \3487_b0 , \3488_b1 , \3488_b0 , \3489_b1 , \3489_b0 , 
		\3490_b1 , \3490_b0 , \3491_b1 , \3491_b0 , \3492_b1 , \3492_b0 , \3493_b1 , \3493_b0 , \3494_b1 , \3494_b0 , 
		\3495_b1 , \3495_b0 , \3496_b1 , \3496_b0 , \3497_b1 , \3497_b0 , \3498_b1 , \3498_b0 , \3499_b1 , \3499_b0 , 
		\3500_b1 , \3500_b0 , \3501_b1 , \3501_b0 , \3502_b1 , \3502_b0 , \3503_b1 , \3503_b0 , \3504_b1 , \3504_b0 , 
		\3505_b1 , \3505_b0 , \3506_b1 , \3506_b0 , \3507_b1 , \3507_b0 , \3508_b1 , \3508_b0 , \3509_b1 , \3509_b0 , 
		\3510_b1 , \3510_b0 , \3511_b1 , \3511_b0 , \3512_b1 , \3512_b0 , \3513_b1 , \3513_b0 , \3514_b1 , \3514_b0 , 
		\3515_b1 , \3515_b0 , \3516_b1 , \3516_b0 , \3517_b1 , \3517_b0 , \3518_b1 , \3518_b0 , \3519_b1 , \3519_b0 , 
		\3520_b1 , \3520_b0 , \3521_b1 , \3521_b0 , \3522_b1 , \3522_b0 , \3523_b1 , \3523_b0 , \3524_b1 , \3524_b0 , 
		\3525_b1 , \3525_b0 , \3526_b1 , \3526_b0 , \3527_b1 , \3527_b0 , \3528_b1 , \3528_b0 , \3529_b1 , \3529_b0 , 
		\3530_b1 , \3530_b0 , \3531_b1 , \3531_b0 , \3532_b1 , \3532_b0 , \3533_b1 , \3533_b0 , \3534_b1 , \3534_b0 , 
		\3535_b1 , \3535_b0 , \3536_b1 , \3536_b0 , \3537_b1 , \3537_b0 , \3538_b1 , \3538_b0 , \3539_b1 , \3539_b0 , 
		\3540_b1 , \3540_b0 , \3541_b1 , \3541_b0 , \3542_b1 , \3542_b0 , \3543_b1 , \3543_b0 , \3544_b1 , \3544_b0 , 
		\3545_b1 , \3545_b0 , \3546_b1 , \3546_b0 , \3547_b1 , \3547_b0 , \3548_b1 , \3548_b0 , \3549_b1 , \3549_b0 , 
		\3550_b1 , \3550_b0 , \3551_b1 , \3551_b0 , \3552_b1 , \3552_b0 , \3553_b1 , \3553_b0 , \3554_b1 , \3554_b0 , 
		\3555_b1 , \3555_b0 , \3556_b1 , \3556_b0 , \3557_b1 , \3557_b0 , \3558_b1 , \3558_b0 , \3559_b1 , \3559_b0 , 
		\3560_b1 , \3560_b0 , \3561_b1 , \3561_b0 , \3562_b1 , \3562_b0 , \3563_b1 , \3563_b0 , \3564_b1 , \3564_b0 , 
		\3565_b1 , \3565_b0 , \3566_b1 , \3566_b0 , \3567_b1 , \3567_b0 , \3568_b1 , \3568_b0 , \3569_b1 , \3569_b0 , 
		\3570_b1 , \3570_b0 , \3571_b1 , \3571_b0 , \3572_b1 , \3572_b0 , \3573_b1 , \3573_b0 , \3574_b1 , \3574_b0 , 
		\3575_b1 , \3575_b0 , \3576_b1 , \3576_b0 , \3577_b1 , \3577_b0 , \3578_b1 , \3578_b0 , \3579_b1 , \3579_b0 , 
		\3580_b1 , \3580_b0 , \3581_b1 , \3581_b0 , \3582_b1 , \3582_b0 , \3583_b1 , \3583_b0 , \3584_b1 , \3584_b0 , 
		\3585_b1 , \3585_b0 , \3586_b1 , \3586_b0 , \3587_b1 , \3587_b0 , \3588_b1 , \3588_b0 , \3589_b1 , \3589_b0 , 
		\3590_b1 , \3590_b0 , \3591_b1 , \3591_b0 , \3592_b1 , \3592_b0 , \3593_b1 , \3593_b0 , \3594_b1 , \3594_b0 , 
		\3595_b1 , \3595_b0 , \3596_b1 , \3596_b0 , \3597_b1 , \3597_b0 , \3598_b1 , \3598_b0 , \3599_b1 , \3599_b0 , 
		\3600_b1 , \3600_b0 , \3601_b1 , \3601_b0 , \3602_b1 , \3602_b0 , \3603_b1 , \3603_b0 , \3604_b1 , \3604_b0 , 
		\3605_b1 , \3605_b0 , \3606_b1 , \3606_b0 , \3607_b1 , \3607_b0 , \3608_b1 , \3608_b0 , \3609_b1 , \3609_b0 , 
		\3610_b1 , \3610_b0 , \3611_b1 , \3611_b0 , \3612_b1 , \3612_b0 , \3613_b1 , \3613_b0 , \3614_b1 , \3614_b0 , 
		\3615_b1 , \3615_b0 , \3616_b1 , \3616_b0 , \3617_b1 , \3617_b0 , \3618_b1 , \3618_b0 , \3619_b1 , \3619_b0 , 
		\3620_b1 , \3620_b0 , \3621_b1 , \3621_b0 , \3622_b1 , \3622_b0 , \3623_b1 , \3623_b0 , \3624_b1 , \3624_b0 , 
		\3625_b1 , \3625_b0 , \3626_b1 , \3626_b0 , \3627_b1 , \3627_b0 , \3628_b1 , \3628_b0 , \3629_b1 , \3629_b0 , 
		\3630_b1 , \3630_b0 , \3631_b1 , \3631_b0 , \3632_b1 , \3632_b0 , \3633_b1 , \3633_b0 , \3634_b1 , \3634_b0 , 
		\3635_b1 , \3635_b0 , \3636_b1 , \3636_b0 , \3637_b1 , \3637_b0 , \3638_b1 , \3638_b0 , \3639_b1 , \3639_b0 , 
		\3640_b1 , \3640_b0 , \3641_b1 , \3641_b0 , \3642_b1 , \3642_b0 , \3643_b1 , \3643_b0 , \3644_b1 , \3644_b0 , 
		\3645_b1 , \3645_b0 , \3646_b1 , \3646_b0 , \3647_b1 , \3647_b0 , \3648_b1 , \3648_b0 , \3649_b1 , \3649_b0 , 
		\3650_b1 , \3650_b0 , \3651_b1 , \3651_b0 , \3652_b1 , \3652_b0 , \3653_b1 , \3653_b0 , \3654_b1 , \3654_b0 , 
		\3655_b1 , \3655_b0 , \3656_b1 , \3656_b0 , \3657_b1 , \3657_b0 , \3658_b1 , \3658_b0 , \3659_b1 , \3659_b0 , 
		\3660_b1 , \3660_b0 , \3661_b1 , \3661_b0 , \3662_b1 , \3662_b0 , \3663_b1 , \3663_b0 , \3664_b1 , \3664_b0 , 
		\3665_b1 , \3665_b0 , \3666_b1 , \3666_b0 , \3667_b1 , \3667_b0 , \3668_b1 , \3668_b0 , \3669_b1 , \3669_b0 , 
		\3670_b1 , \3670_b0 , \3671_b1 , \3671_b0 , \3672_b1 , \3672_b0 , \3673_b1 , \3673_b0 , \3674_b1 , \3674_b0 , 
		\3675_b1 , \3675_b0 , \3676_b1 , \3676_b0 , \3677_b1 , \3677_b0 , \3678_b1 , \3678_b0 , \3679_b1 , \3679_b0 , 
		\3680_b1 , \3680_b0 , \3681_b1 , \3681_b0 , \3682_b1 , \3682_b0 , \3683_b1 , \3683_b0 , \3684_b1 , \3684_b0 , 
		\3685_b1 , \3685_b0 , \3686_b1 , \3686_b0 , \3687_b1 , \3687_b0 , \3688_b1 , \3688_b0 , \3689_b1 , \3689_b0 , 
		\3690_b1 , \3690_b0 , \3691_b1 , \3691_b0 , \3692_b1 , \3692_b0 , \3693_b1 , \3693_b0 , \3694_b1 , \3694_b0 , 
		\3695_b1 , \3695_b0 , \3696_b1 , \3696_b0 , \3697_b1 , \3697_b0 , \3698_b1 , \3698_b0 , \3699_b1 , \3699_b0 , 
		\3700_b1 , \3700_b0 , \3701_b1 , \3701_b0 , \3702_b1 , \3702_b0 , \3703_b1 , \3703_b0 , \3704_b1 , \3704_b0 , 
		\3705_b1 , \3705_b0 , \3706_b1 , \3706_b0 , \3707_b1 , \3707_b0 , \3708_b1 , \3708_b0 , \3709_b1 , \3709_b0 , 
		\3710_b1 , \3710_b0 , \3711_b1 , \3711_b0 , \3712_b1 , \3712_b0 , \3713_b1 , \3713_b0 , \3714_b1 , \3714_b0 , 
		\3715_b1 , \3715_b0 , \3716_b1 , \3716_b0 , \3717_b1 , \3717_b0 , \3718_b1 , \3718_b0 , \3719_b1 , \3719_b0 , 
		\3720_b1 , \3720_b0 , \3721_b1 , \3721_b0 , \3722_b1 , \3722_b0 , \3723_b1 , \3723_b0 , \3724_b1 , \3724_b0 , 
		\3725_b1 , \3725_b0 , \3726_b1 , \3726_b0 , \3727_b1 , \3727_b0 , \3728_b1 , \3728_b0 , \3729_b1 , \3729_b0 , 
		\3730_b1 , \3730_b0 , \3731_b1 , \3731_b0 , \3732_b1 , \3732_b0 , \3733_b1 , \3733_b0 , \3734_b1 , \3734_b0 , 
		\3735_b1 , \3735_b0 , \3736_b1 , \3736_b0 , \3737_b1 , \3737_b0 , \3738_b1 , \3738_b0 , \3739_b1 , \3739_b0 , 
		\3740_b1 , \3740_b0 , \3741_b1 , \3741_b0 , \3742_b1 , \3742_b0 , \3743_b1 , \3743_b0 , \3744_b1 , \3744_b0 , 
		\3745_b1 , \3745_b0 , \3746_b1 , \3746_b0 , \3747_b1 , \3747_b0 , \3748_b1 , \3748_b0 , \3749_b1 , \3749_b0 , 
		\3750_b1 , \3750_b0 , \3751_b1 , \3751_b0 , \3752_b1 , \3752_b0 , \3753_b1 , \3753_b0 , \3754_b1 , \3754_b0 , 
		\3755_b1 , \3755_b0 , \3756_b1 , \3756_b0 , \3757_b1 , \3757_b0 , \3758_b1 , \3758_b0 , \3759_b1 , \3759_b0 , 
		\3760_b1 , \3760_b0 , \3761_b1 , \3761_b0 , \3762_b1 , \3762_b0 , \3763_b1 , \3763_b0 , \3764_b1 , \3764_b0 , 
		\3765_b1 , \3765_b0 , \3766_b1 , \3766_b0 , \3767_b1 , \3767_b0 , \3768_b1 , \3768_b0 , \3769_b1 , \3769_b0 , 
		\3770_b1 , \3770_b0 , \3771_b1 , \3771_b0 , \3772_b1 , \3772_b0 , \3773_b1 , \3773_b0 , \3774_b1 , \3774_b0 , 
		\3775_b1 , \3775_b0 , \3776_b1 , \3776_b0 , \3777_b1 , \3777_b0 , \3778_b1 , \3778_b0 , \3779_b1 , \3779_b0 , 
		\3780_b1 , \3780_b0 , \3781_b1 , \3781_b0 , \3782_b1 , \3782_b0 , \3783_b1 , \3783_b0 , \3784_b1 , \3784_b0 , 
		\3785_b1 , \3785_b0 , \3786_b1 , \3786_b0 , \3787_b1 , \3787_b0 , \3788_b1 , \3788_b0 , \3789_b1 , \3789_b0 , 
		\3790_b1 , \3790_b0 , \3791_b1 , \3791_b0 , \3792_b1 , \3792_b0 , \3793_b1 , \3793_b0 , \3794_b1 , \3794_b0 , 
		\3795_b1 , \3795_b0 , \3796_b1 , \3796_b0 , \3797_b1 , \3797_b0 , \3798_b1 , \3798_b0 , \3799_b1 , \3799_b0 , 
		\3800_b1 , \3800_b0 , \3801_b1 , \3801_b0 , \3802_b1 , \3802_b0 , \3803_b1 , \3803_b0 , \3804_b1 , \3804_b0 , 
		\3805_b1 , \3805_b0 , \3806_b1 , \3806_b0 , \3807_b1 , \3807_b0 , \3808_b1 , \3808_b0 , \3809_b1 , \3809_b0 , 
		\3810_b1 , \3810_b0 , \3811_b1 , \3811_b0 , \3812_b1 , \3812_b0 , \3813_b1 , \3813_b0 , \3814_b1 , \3814_b0 , 
		\3815_b1 , \3815_b0 , \3816_b1 , \3816_b0 , \3817_b1 , \3817_b0 , \3818_b1 , \3818_b0 , \3819_b1 , \3819_b0 , 
		\3820_b1 , \3820_b0 , \3821_b1 , \3821_b0 , \3822_b1 , \3822_b0 , \3823_b1 , \3823_b0 , \3824_b1 , \3824_b0 , 
		\3825_b1 , \3825_b0 , \3826_b1 , \3826_b0 , \3827_b1 , \3827_b0 , \3828_b1 , \3828_b0 , \3829_b1 , \3829_b0 , 
		\3830_b1 , \3830_b0 , \3831_b1 , \3831_b0 , \3832_b1 , \3832_b0 , \3833_b1 , \3833_b0 , \3834_b1 , \3834_b0 , 
		\3835_b1 , \3835_b0 , \3836_b1 , \3836_b0 , \3837_b1 , \3837_b0 , \3838_b1 , \3838_b0 , \3839_b1 , \3839_b0 , 
		\3840_b1 , \3840_b0 , \3841_b1 , \3841_b0 , \3842_b1 , \3842_b0 , \3843_b1 , \3843_b0 , \3844_b1 , \3844_b0 , 
		\3845_b1 , \3845_b0 , \3846_b1 , \3846_b0 , \3847_b1 , \3847_b0 , \3848_b1 , \3848_b0 , \3849_b1 , \3849_b0 , 
		\3850_b1 , \3850_b0 , \3851_b1 , \3851_b0 , \3852_b1 , \3852_b0 , \3853_b1 , \3853_b0 , \3854_b1 , \3854_b0 , 
		\3855_b1 , \3855_b0 , \3856_b1 , \3856_b0 , \3857_b1 , \3857_b0 , \3858_b1 , \3858_b0 , \3859_b1 , \3859_b0 , 
		\3860_b1 , \3860_b0 , \3861_b1 , \3861_b0 , \3862_b1 , \3862_b0 , \3863_b1 , \3863_b0 , \3864_b1 , \3864_b0 , 
		\3865_b1 , \3865_b0 , \3866_b1 , \3866_b0 , \3867_b1 , \3867_b0 , \3868_b1 , \3868_b0 , \3869_b1 , \3869_b0 , 
		\3870_b1 , \3870_b0 , \3871_b1 , \3871_b0 , \3872_b1 , \3872_b0 , \3873_b1 , \3873_b0 , \3874_b1 , \3874_b0 , 
		\3875_b1 , \3875_b0 , \3876_b1 , \3876_b0 , \3877_b1 , \3877_b0 , \3878_b1 , \3878_b0 , \3879_b1 , \3879_b0 , 
		\3880_b1 , \3880_b0 , \3881_b1 , \3881_b0 , \3882_b1 , \3882_b0 , \3883_b1 , \3883_b0 , \3884_b1 , \3884_b0 , 
		\3885_b1 , \3885_b0 , \3886_b1 , \3886_b0 , \3887_b1 , \3887_b0 , \3888_b1 , \3888_b0 , \3889_b1 , \3889_b0 , 
		\3890_b1 , \3890_b0 , \3891_b1 , \3891_b0 , \3892_b1 , \3892_b0 , \3893_b1 , \3893_b0 , \3894_b1 , \3894_b0 , 
		\3895_b1 , \3895_b0 , \3896_b1 , \3896_b0 , \3897_b1 , \3897_b0 , \3898_b1 , \3898_b0 , \3899_b1 , \3899_b0 , 
		\3900_b1 , \3900_b0 , \3901_b1 , \3901_b0 , \3902_b1 , \3902_b0 , \3903_b1 , \3903_b0 , \3904_b1 , \3904_b0 , 
		\3905_b1 , \3905_b0 , \3906_b1 , \3906_b0 , \3907_b1 , \3907_b0 , \3908_b1 , \3908_b0 , \3909_b1 , \3909_b0 , 
		\3910_b1 , \3910_b0 , \3911_b1 , \3911_b0 , \3912_b1 , \3912_b0 , \3913_b1 , \3913_b0 , \3914_b1 , \3914_b0 , 
		\3915_b1 , \3915_b0 , \3916_b1 , \3916_b0 , \3917_b1 , \3917_b0 , \3918_b1 , \3918_b0 , \3919_b1 , \3919_b0 , 
		\3920_b1 , \3920_b0 , \3921_b1 , \3921_b0 , \3922_b1 , \3922_b0 , \3923_b1 , \3923_b0 , \3924_b1 , \3924_b0 , 
		\3925_b1 , \3925_b0 , \3926_b1 , \3926_b0 , \3927_b1 , \3927_b0 , \3928_b1 , \3928_b0 , \3929_b1 , \3929_b0 , 
		\3930_b1 , \3930_b0 , \3931_b1 , \3931_b0 , \3932_b1 , \3932_b0 , \3933_b1 , \3933_b0 , \3934_b1 , \3934_b0 , 
		\3935_b1 , \3935_b0 , \3936_b1 , \3936_b0 , \3937_b1 , \3937_b0 , \3938_b1 , \3938_b0 , \3939_b1 , \3939_b0 , 
		\3940_b1 , \3940_b0 , \3941_b1 , \3941_b0 , \3942_b1 , \3942_b0 , \3943_b1 , \3943_b0 , \3944_b1 , \3944_b0 , 
		\3945_b1 , \3945_b0 , \3946_b1 , \3946_b0 , \3947_b1 , \3947_b0 , \3948_b1 , \3948_b0 , \3949_b1 , \3949_b0 , 
		\3950_b1 , \3950_b0 , \3951_b1 , \3951_b0 , \3952_b1 , \3952_b0 , \3953_b1 , \3953_b0 , \3954_b1 , \3954_b0 , 
		\3955_b1 , \3955_b0 , \3956_b1 , \3956_b0 , \3957_b1 , \3957_b0 , \3958_b1 , \3958_b0 , \3959_b1 , \3959_b0 , 
		\3960_b1 , \3960_b0 , \3961_b1 , \3961_b0 , \3962_b1 , \3962_b0 , \3963_b1 , \3963_b0 , \3964_b1 , \3964_b0 , 
		\3965_b1 , \3965_b0 , \3966_b1 , \3966_b0 , \3967_b1 , \3967_b0 , \3968_b1 , \3968_b0 , \3969_b1 , \3969_b0 , 
		\3970_b1 , \3970_b0 , \3971_b1 , \3971_b0 , \3972_b1 , \3972_b0 , \3973_b1 , \3973_b0 , \3974_b1 , \3974_b0 , 
		\3975_b1 , \3975_b0 , \3976_b1 , \3976_b0 , \3977_b1 , \3977_b0 , \3978_b1 , \3978_b0 , \3979_b1 , \3979_b0 , 
		\3980_b1 , \3980_b0 , \3981_b1 , \3981_b0 , \3982_b1 , \3982_b0 , \3983_b1 , \3983_b0 , \3984_b1 , \3984_b0 , 
		\3985_b1 , \3985_b0 , \3986_b1 , \3986_b0 , \3987_b1 , \3987_b0 , \3988_b1 , \3988_b0 , \3989_b1 , \3989_b0 , 
		\3990_b1 , \3990_b0 , \3991_b1 , \3991_b0 , \3992_b1 , \3992_b0 , \3993_b1 , \3993_b0 , \3994_b1 , \3994_b0 , 
		\3995_b1 , \3995_b0 , \3996_b1 , \3996_b0 , \3997_b1 , \3997_b0 , \3998_b1 , \3998_b0 , \3999_b1 , \3999_b0 , 
		\4000_b1 , \4000_b0 , \4001_b1 , \4001_b0 , \4002_b1 , \4002_b0 , \4003_b1 , \4003_b0 , \4004_b1 , \4004_b0 , 
		\4005_b1 , \4005_b0 , \4006_b1 , \4006_b0 , \4007_b1 , \4007_b0 , \4008_b1 , \4008_b0 , \4009_b1 , \4009_b0 , 
		\4010_b1 , \4010_b0 , \4011_b1 , \4011_b0 , \4012_b1 , \4012_b0 , \4013_b1 , \4013_b0 , \4014_b1 , \4014_b0 , 
		\4015_b1 , \4015_b0 , \4016_b1 , \4016_b0 , \4017_b1 , \4017_b0 , \4018_b1 , \4018_b0 , \4019_b1 , \4019_b0 , 
		\4020_b1 , \4020_b0 , \4021_b1 , \4021_b0 , \4022_b1 , \4022_b0 , \4023_b1 , \4023_b0 , \4024_b1 , \4024_b0 , 
		\4025_b1 , \4025_b0 , \4026_b1 , \4026_b0 , \4027_b1 , \4027_b0 , \4028_b1 , \4028_b0 , \4029_b1 , \4029_b0 , 
		\4030_b1 , \4030_b0 , \4031_b1 , \4031_b0 , \4032_b1 , \4032_b0 , \4033_b1 , \4033_b0 , \4034_b1 , \4034_b0 , 
		\4035_b1 , \4035_b0 , \4036_b1 , \4036_b0 , \4037_b1 , \4037_b0 , \4038_b1 , \4038_b0 , \4039_b1 , \4039_b0 , 
		\4040_b1 , \4040_b0 , \4041_b1 , \4041_b0 , \4042_b1 , \4042_b0 , \4043_b1 , \4043_b0 , \4044_b1 , \4044_b0 , 
		\4045_b1 , \4045_b0 , \4046_b1 , \4046_b0 , \4047_b1 , \4047_b0 , \4048_b1 , \4048_b0 , \4049_b1 , \4049_b0 , 
		\4050_b1 , \4050_b0 , \4051_b1 , \4051_b0 , \4052_b1 , \4052_b0 , \4053_b1 , \4053_b0 , \4054_b1 , \4054_b0 , 
		\4055_b1 , \4055_b0 , \4056_b1 , \4056_b0 , \4057_b1 , \4057_b0 , \4058_b1 , \4058_b0 , \4059_b1 , \4059_b0 , 
		\4060_b1 , \4060_b0 , \4061_b1 , \4061_b0 , \4062_b1 , \4062_b0 , \4063_b1 , \4063_b0 , \4064_b1 , \4064_b0 , 
		\4065_b1 , \4065_b0 , \4066_b1 , \4066_b0 , \4067_b1 , \4067_b0 , \4068_b1 , \4068_b0 , \4069_b1 , \4069_b0 , 
		\4070_b1 , \4070_b0 , \4071_b1 , \4071_b0 , \4072_b1 , \4072_b0 , \4073_b1 , \4073_b0 , \4074_b1 , \4074_b0 , 
		\4075_b1 , \4075_b0 , \4076_b1 , \4076_b0 , \4077_b1 , \4077_b0 , \4078_b1 , \4078_b0 , \4079_b1 , \4079_b0 , 
		\4080_b1 , \4080_b0 , \4081_b1 , \4081_b0 , \4082_b1 , \4082_b0 , \4083_b1 , \4083_b0 , \4084_b1 , \4084_b0 , 
		\4085_b1 , \4085_b0 , \4086_b1 , \4086_b0 , \4087_b1 , \4087_b0 , \4088_b1 , \4088_b0 , \4089_b1 , \4089_b0 , 
		\4090_b1 , \4090_b0 , \4091_b1 , \4091_b0 , \4092_b1 , \4092_b0 , \4093_b1 , \4093_b0 , \4094_b1 , \4094_b0 , 
		\4095_b1 , \4095_b0 , \4096_b1 , \4096_b0 , \4097_b1 , \4097_b0 , \4098_b1 , \4098_b0 , \4099_b1 , \4099_b0 , 
		\4100_b1 , \4100_b0 , \4101_b1 , \4101_b0 , \4102_b1 , \4102_b0 , \4103_b1 , \4103_b0 , \4104_b1 , \4104_b0 , 
		\4105_b1 , \4105_b0 , \4106_b1 , \4106_b0 , \4107_b1 , \4107_b0 , \4108_b1 , \4108_b0 , \4109_b1 , \4109_b0 , 
		\4110_b1 , \4110_b0 , \4111_b1 , \4111_b0 , \4112_b1 , \4112_b0 , \4113_b1 , \4113_b0 , \4114_b1 , \4114_b0 , 
		\4115_b1 , \4115_b0 , \4116_b1 , \4116_b0 , \4117_b1 , \4117_b0 , \4118_b1 , \4118_b0 , \4119_b1 , \4119_b0 , 
		\4120_b1 , \4120_b0 , \4121_b1 , \4121_b0 , \4122_b1 , \4122_b0 , \4123_b1 , \4123_b0 , \4124_b1 , \4124_b0 , 
		\4125_b1 , \4125_b0 , \4126_b1 , \4126_b0 , \4127_b1 , \4127_b0 , \4128_b1 , \4128_b0 , \4129_b1 , \4129_b0 , 
		\4130_b1 , \4130_b0 , \4131_b1 , \4131_b0 , \4132_b1 , \4132_b0 , \4133_b1 , \4133_b0 , \4134_b1 , \4134_b0 , 
		\4135_b1 , \4135_b0 , \4136_b1 , \4136_b0 , \4137_b1 , \4137_b0 , \4138_b1 , \4138_b0 , \4139_b1 , \4139_b0 , 
		\4140_b1 , \4140_b0 , \4141_b1 , \4141_b0 , \4142_b1 , \4142_b0 , \4143_b1 , \4143_b0 , \4144_b1 , \4144_b0 , 
		\4145_b1 , \4145_b0 , \4146_b1 , \4146_b0 , \4147_b1 , \4147_b0 , \4148_b1 , \4148_b0 , \4149_b1 , \4149_b0 , 
		\4150_b1 , \4150_b0 , \4151_b1 , \4151_b0 , \4152_b1 , \4152_b0 , \4153_b1 , \4153_b0 , \4154_b1 , \4154_b0 , 
		\4155_b1 , \4155_b0 , \4156_b1 , \4156_b0 , \4157_b1 , \4157_b0 , \4158_b1 , \4158_b0 , \4159_b1 , \4159_b0 , 
		\4160_b1 , \4160_b0 , \4161_b1 , \4161_b0 , \4162_b1 , \4162_b0 , \4163_b1 , \4163_b0 , \4164_b1 , \4164_b0 , 
		\4165_b1 , \4165_b0 , \4166_b1 , \4166_b0 , \4167_b1 , \4167_b0 , \4168_b1 , \4168_b0 , \4169_b1 , \4169_b0 , 
		\4170_b1 , \4170_b0 , \4171_b1 , \4171_b0 , \4172_b1 , \4172_b0 , \4173_b1 , \4173_b0 , \4174_b1 , \4174_b0 , 
		\4175_b1 , \4175_b0 , \4176_b1 , \4176_b0 , \4177_b1 , \4177_b0 , \4178_b1 , \4178_b0 , \4179_b1 , \4179_b0 , 
		\4180_b1 , \4180_b0 , \4181_b1 , \4181_b0 , \4182_b1 , \4182_b0 , \4183_b1 , \4183_b0 , \4184_b1 , \4184_b0 , 
		\4185_b1 , \4185_b0 , \4186_b1 , \4186_b0 , \4187_b1 , \4187_b0 , \4188_b1 , \4188_b0 , \4189_b1 , \4189_b0 , 
		\4190_b1 , \4190_b0 , \4191_b1 , \4191_b0 , \4192_b1 , \4192_b0 , \4193_b1 , \4193_b0 , \4194_b1 , \4194_b0 , 
		\4195_b1 , \4195_b0 , \4196_b1 , \4196_b0 , \4197_b1 , \4197_b0 , \4198_b1 , \4198_b0 , \4199_b1 , \4199_b0 , 
		\4200_b1 , \4200_b0 , \4201_b1 , \4201_b0 , \4202_b1 , \4202_b0 , \4203_b1 , \4203_b0 , \4204_b1 , \4204_b0 , 
		\4205_b1 , \4205_b0 , \4206_b1 , \4206_b0 , \4207_b1 , \4207_b0 , \4208_b1 , \4208_b0 , \4209_b1 , \4209_b0 , 
		\4210_b1 , \4210_b0 , \4211_b1 , \4211_b0 , \4212_b1 , \4212_b0 , \4213_b1 , \4213_b0 , \4214_b1 , \4214_b0 , 
		\4215_b1 , \4215_b0 , \4216_b1 , \4216_b0 , \4217_b1 , \4217_b0 , \4218_b1 , \4218_b0 , \4219_b1 , \4219_b0 , 
		\4220_b1 , \4220_b0 , \4221_b1 , \4221_b0 , \4222_b1 , \4222_b0 , \4223_b1 , \4223_b0 , \4224_b1 , \4224_b0 , 
		\4225_b1 , \4225_b0 , \4226_b1 , \4226_b0 , \4227_b1 , \4227_b0 , \4228_b1 , \4228_b0 , \4229_b1 , \4229_b0 , 
		\4230_b1 , \4230_b0 , \4231_b1 , \4231_b0 , \4232_b1 , \4232_b0 , \4233_b1 , \4233_b0 , \4234_b1 , \4234_b0 , 
		\4235_b1 , \4235_b0 , \4236_b1 , \4236_b0 , \4237_b1 , \4237_b0 , \4238_b1 , \4238_b0 , \4239_b1 , \4239_b0 , 
		\4240_b1 , \4240_b0 , \4241_b1 , \4241_b0 , \4242_b1 , \4242_b0 , \4243_b1 , \4243_b0 , \4244_b1 , \4244_b0 , 
		\4245_b1 , \4245_b0 , \4246_b1 , \4246_b0 , \4247_b1 , \4247_b0 , \4248_b1 , \4248_b0 , \4249_b1 , \4249_b0 , 
		\4250_b1 , \4250_b0 , \4251_b1 , \4251_b0 , \4252_b1 , \4252_b0 , \4253_b1 , \4253_b0 , \4254_b1 , \4254_b0 , 
		\4255_b1 , \4255_b0 , \4256_b1 , \4256_b0 , \4257_b1 , \4257_b0 , \4258_b1 , \4258_b0 , \4259_b1 , \4259_b0 , 
		\4260_b1 , \4260_b0 , \4261_b1 , \4261_b0 , \4262_b1 , \4262_b0 , \4263_b1 , \4263_b0 , \4264_b1 , \4264_b0 , 
		\4265_b1 , \4265_b0 , \4266_b1 , \4266_b0 , \4267_b1 , \4267_b0 , \4268_b1 , \4268_b0 , \4269_b1 , \4269_b0 , 
		\4270_b1 , \4270_b0 , \4271_b1 , \4271_b0 , \4272_b1 , \4272_b0 , \4273_b1 , \4273_b0 , \4274_b1 , \4274_b0 , 
		\4275_b1 , \4275_b0 , \4276_b1 , \4276_b0 , \4277_b1 , \4277_b0 , \4278_b1 , \4278_b0 , \4279_b1 , \4279_b0 , 
		\4280_b1 , \4280_b0 , \4281_b1 , \4281_b0 , \4282_b1 , \4282_b0 , \4283_b1 , \4283_b0 , \4284_b1 , \4284_b0 , 
		\4285_b1 , \4285_b0 , \4286_b1 , \4286_b0 , \4287_b1 , \4287_b0 , \4288_b1 , \4288_b0 , \4289_b1 , \4289_b0 , 
		\4290_b1 , \4290_b0 , \4291_b1 , \4291_b0 , \4292_b1 , \4292_b0 , \4293_b1 , \4293_b0 , \4294_b1 , \4294_b0 , 
		\4295_b1 , \4295_b0 , \4296_b1 , \4296_b0 , \4297_b1 , \4297_b0 , \4298_b1 , \4298_b0 , \4299_b1 , \4299_b0 , 
		\4300_b1 , \4300_b0 , \4301_b1 , \4301_b0 , \4302_b1 , \4302_b0 , \4303_b1 , \4303_b0 , \4304_b1 , \4304_b0 , 
		\4305_b1 , \4305_b0 , \4306_b1 , \4306_b0 , \4307_b1 , \4307_b0 , \4308_b1 , \4308_b0 , \4309_b1 , \4309_b0 , 
		\4310_b1 , \4310_b0 , \4311_b1 , \4311_b0 , \4312_b1 , \4312_b0 , \4313_b1 , \4313_b0 , \4314_b1 , \4314_b0 , 
		\4315_b1 , \4315_b0 , \4316_b1 , \4316_b0 , \4317_b1 , \4317_b0 , \4318_b1 , \4318_b0 , \4319_b1 , \4319_b0 , 
		\4320_b1 , \4320_b0 , \4321_b1 , \4321_b0 , \4322_b1 , \4322_b0 , \4323_b1 , \4323_b0 , \4324_b1 , \4324_b0 , 
		\4325_b1 , \4325_b0 , \4326_b1 , \4326_b0 , \4327_b1 , \4327_b0 , \4328_b1 , \4328_b0 , \4329_b1 , \4329_b0 , 
		\4330_b1 , \4330_b0 , \4331_b1 , \4331_b0 , \4332_b1 , \4332_b0 , \4333_b1 , \4333_b0 , \4334_b1 , \4334_b0 , 
		\4335_b1 , \4335_b0 , \4336_b1 , \4336_b0 , \4337_b1 , \4337_b0 , \4338_b1 , \4338_b0 , \4339_b1 , \4339_b0 , 
		\4340_b1 , \4340_b0 , \4341_b1 , \4341_b0 , \4342_b1 , \4342_b0 , \4343_b1 , \4343_b0 , \4344_b1 , \4344_b0 , 
		\4345_b1 , \4345_b0 , \4346_b1 , \4346_b0 , \4347_b1 , \4347_b0 , \4348_b1 , \4348_b0 , \4349_b1 , \4349_b0 , 
		\4350_b1 , \4350_b0 , \4351_b1 , \4351_b0 , \4352_b1 , \4352_b0 , \4353_b1 , \4353_b0 , \4354_b1 , \4354_b0 , 
		\4355_b1 , \4355_b0 , \4356_b1 , \4356_b0 , \4357_b1 , \4357_b0 , \4358_b1 , \4358_b0 , \4359_b1 , \4359_b0 , 
		\4360_b1 , \4360_b0 , \4361_b1 , \4361_b0 , \4362_b1 , \4362_b0 , \4363_b1 , \4363_b0 , \4364_b1 , \4364_b0 , 
		\4365_b1 , \4365_b0 , \4366_b1 , \4366_b0 , \4367_b1 , \4367_b0 , \4368_b1 , \4368_b0 , \4369_b1 , \4369_b0 , 
		\4370_b1 , \4370_b0 , \4371_b1 , \4371_b0 , \4372_b1 , \4372_b0 , \4373_b1 , \4373_b0 , \4374_b1 , \4374_b0 , 
		\4375_b1 , \4375_b0 , \4376_b1 , \4376_b0 , \4377_b1 , \4377_b0 , \4378_b1 , \4378_b0 , \4379_b1 , \4379_b0 , 
		\4380_b1 , \4380_b0 , \4381_b1 , \4381_b0 , \4382_b1 , \4382_b0 , \4383_b1 , \4383_b0 , \4384_b1 , \4384_b0 , 
		\4385_b1 , \4385_b0 , \4386_b1 , \4386_b0 , \4387_b1 , \4387_b0 , \4388_b1 , \4388_b0 , \4389_b1 , \4389_b0 , 
		\4390_b1 , \4390_b0 , \4391_b1 , \4391_b0 , \4392_b1 , \4392_b0 , \4393_b1 , \4393_b0 , \4394_b1 , \4394_b0 , 
		\4395_b1 , \4395_b0 , \4396_b1 , \4396_b0 , \4397_b1 , \4397_b0 , \4398_b1 , \4398_b0 , \4399_b1 , \4399_b0 , 
		\4400_b1 , \4400_b0 , \4401_b1 , \4401_b0 , \4402_b1 , \4402_b0 , \4403_b1 , \4403_b0 , \4404_b1 , \4404_b0 , 
		\4405_b1 , \4405_b0 , \4406_b1 , \4406_b0 , \4407_b1 , \4407_b0 , \4408_b1 , \4408_b0 , \4409_b1 , \4409_b0 , 
		\4410_b1 , \4410_b0 , \4411_b1 , \4411_b0 , \4412_b1 , \4412_b0 , \4413_b1 , \4413_b0 , \4414_b1 , \4414_b0 , 
		\4415_b1 , \4415_b0 , \4416_b1 , \4416_b0 , \4417_b1 , \4417_b0 , \4418_b1 , \4418_b0 , \4419_b1 , \4419_b0 , 
		\4420_b1 , \4420_b0 , \4421_b1 , \4421_b0 , \4422_b1 , \4422_b0 , \4423_b1 , \4423_b0 , \4424_b1 , \4424_b0 , 
		\4425_b1 , \4425_b0 , \4426_b1 , \4426_b0 , \4427_b1 , \4427_b0 , \4428_b1 , \4428_b0 , \4429_b1 , \4429_b0 , 
		\4430_b1 , \4430_b0 , \4431_b1 , \4431_b0 , \4432_b1 , \4432_b0 , \4433_b1 , \4433_b0 , \4434_b1 , \4434_b0 , 
		\4435_b1 , \4435_b0 , \4436_b1 , \4436_b0 , \4437_b1 , \4437_b0 , \4438_b1 , \4438_b0 , \4439_b1 , \4439_b0 , 
		\4440_b1 , \4440_b0 , \4441_b1 , \4441_b0 , \4442_b1 , \4442_b0 , \4443_b1 , \4443_b0 , \4444_b1 , \4444_b0 , 
		\4445_b1 , \4445_b0 , \4446_b1 , \4446_b0 , \4447_b1 , \4447_b0 , \4448_b1 , \4448_b0 , \4449_b1 , \4449_b0 , 
		\4450_b1 , \4450_b0 , \4451_b1 , \4451_b0 , \4452_b1 , \4452_b0 , \4453_b1 , \4453_b0 , \4454_b1 , \4454_b0 , 
		\4455_b1 , \4455_b0 , \4456_b1 , \4456_b0 , \4457_b1 , \4457_b0 , \4458_b1 , \4458_b0 , \4459_b1 , \4459_b0 , 
		\4460_b1 , \4460_b0 , \4461_b1 , \4461_b0 , \4462_b1 , \4462_b0 , \4463_b1 , \4463_b0 , \4464_b1 , \4464_b0 , 
		\4465_b1 , \4465_b0 , \4466_b1 , \4466_b0 , \4467_b1 , \4467_b0 , \4468_b1 , \4468_b0 , \4469_b1 , \4469_b0 , 
		\4470_b1 , \4470_b0 , \4471_b1 , \4471_b0 , \4472_b1 , \4472_b0 , \4473_b1 , \4473_b0 , \4474_b1 , \4474_b0 , 
		\4475_b1 , \4475_b0 , \4476_b1 , \4476_b0 , \4477_b1 , \4477_b0 , \4478_b1 , \4478_b0 , \4479_b1 , \4479_b0 , 
		\4480_b1 , \4480_b0 , \4481_b1 , \4481_b0 , \4482_b1 , \4482_b0 , \4483_b1 , \4483_b0 , \4484_b1 , \4484_b0 , 
		\4485_b1 , \4485_b0 , \4486_b1 , \4486_b0 , \4487_b1 , \4487_b0 , \4488_b1 , \4488_b0 , \4489_b1 , \4489_b0 , 
		\4490_b1 , \4490_b0 , \4491_b1 , \4491_b0 , \4492_b1 , \4492_b0 , \4493_b1 , \4493_b0 , \4494_b1 , \4494_b0 , 
		\4495_b1 , \4495_b0 , \4496_b1 , \4496_b0 , \4497_b1 , \4497_b0 , \4498_b1 , \4498_b0 , \4499_b1 , \4499_b0 , 
		\4500_b1 , \4500_b0 , \4501_b1 , \4501_b0 , \4502_b1 , \4502_b0 , \4503_b1 , \4503_b0 , \4504_b1 , \4504_b0 , 
		\4505_b1 , \4505_b0 , \4506_b1 , \4506_b0 , \4507_b1 , \4507_b0 , \4508_b1 , \4508_b0 , \4509_b1 , \4509_b0 , 
		\4510_b1 , \4510_b0 , \4511_b1 , \4511_b0 , \4512_b1 , \4512_b0 , \4513_b1 , \4513_b0 , \4514_b1 , \4514_b0 , 
		\4515_b1 , \4515_b0 , \4516_b1 , \4516_b0 , \4517_b1 , \4517_b0 , \4518_b1 , \4518_b0 , \4519_b1 , \4519_b0 , 
		\4520_b1 , \4520_b0 , \4521_b1 , \4521_b0 , \4522_b1 , \4522_b0 , \4523_b1 , \4523_b0 , \4524_b1 , \4524_b0 , 
		\4525_b1 , \4525_b0 , \4526_b1 , \4526_b0 , \4527_b1 , \4527_b0 , \4528_b1 , \4528_b0 , \4529_b1 , \4529_b0 , 
		\4530_b1 , \4530_b0 , \4531_b1 , \4531_b0 , \4532_b1 , \4532_b0 , \4533_b1 , \4533_b0 , \4534_b1 , \4534_b0 , 
		\4535_b1 , \4535_b0 , \4536_b1 , \4536_b0 , \4537_b1 , \4537_b0 , \4538_b1 , \4538_b0 , \4539_b1 , \4539_b0 , 
		\4540_b1 , \4540_b0 , \4541_b1 , \4541_b0 , \4542_b1 , \4542_b0 , \4543_b1 , \4543_b0 , \4544_b1 , \4544_b0 , 
		\4545_b1 , \4545_b0 , \4546_b1 , \4546_b0 , \4547_b1 , \4547_b0 , \4548_b1 , \4548_b0 , \4549_b1 , \4549_b0 , 
		\4550_b1 , \4550_b0 , \4551_b1 , \4551_b0 , \4552_b1 , \4552_b0 , \4553_b1 , \4553_b0 , \4554_b1 , \4554_b0 , 
		\4555_b1 , \4555_b0 , \4556_b1 , \4556_b0 , \4557_b1 , \4557_b0 , \4558_b1 , \4558_b0 , \4559_b1 , \4559_b0 , 
		\4560_b1 , \4560_b0 , \4561_b1 , \4561_b0 , \4562_b1 , \4562_b0 , \4563_b1 , \4563_b0 , \4564_b1 , \4564_b0 , 
		\4565_b1 , \4565_b0 , \4566_b1 , \4566_b0 , \4567_b1 , \4567_b0 , \4568_b1 , \4568_b0 , \4569_b1 , \4569_b0 , 
		\4570_b1 , \4570_b0 , \4571_b1 , \4571_b0 , \4572_b1 , \4572_b0 , \4573_b1 , \4573_b0 , \4574_b1 , \4574_b0 , 
		\4575_b1 , \4575_b0 , \4576_b1 , \4576_b0 , \4577_b1 , \4577_b0 , \4578_b1 , \4578_b0 , \4579_b1 , \4579_b0 , 
		\4580_b1 , \4580_b0 , \4581_b1 , \4581_b0 , \4582_b1 , \4582_b0 , \4583_b1 , \4583_b0 , \4584_b1 , \4584_b0 , 
		\4585_b1 , \4585_b0 , \4586_b1 , \4586_b0 , \4587_b1 , \4587_b0 , \4588_b1 , \4588_b0 , \4589_b1 , \4589_b0 , 
		\4590_b1 , \4590_b0 , \4591_b1 , \4591_b0 , \4592_b1 , \4592_b0 , \4593_b1 , \4593_b0 , \4594_b1 , \4594_b0 , 
		\4595_b1 , \4595_b0 , \4596_b1 , \4596_b0 , \4597_b1 , \4597_b0 , \4598_b1 , \4598_b0 , \4599_b1 , \4599_b0 , 
		\4600_b1 , \4600_b0 , \4601_b1 , \4601_b0 , \4602_b1 , \4602_b0 , \4603_b1 , \4603_b0 , \4604_b1 , \4604_b0 , 
		\4605_b1 , \4605_b0 , \4606_b1 , \4606_b0 , \4607_b1 , \4607_b0 , \4608_b1 , \4608_b0 , \4609_b1 , \4609_b0 , 
		\4610_b1 , \4610_b0 , \4611_b1 , \4611_b0 , \4612_b1 , \4612_b0 , \4613_b1 , \4613_b0 , \4614_b1 , \4614_b0 , 
		\4615_b1 , \4615_b0 , \4616_b1 , \4616_b0 , \4617_b1 , \4617_b0 , \4618_b1 , \4618_b0 , \4619_b1 , \4619_b0 , 
		\4620_b1 , \4620_b0 , \4621_b1 , \4621_b0 , \4622_b1 , \4622_b0 , \4623_b1 , \4623_b0 , \4624_b1 , \4624_b0 , 
		\4625_b1 , \4625_b0 , \4626_b1 , \4626_b0 , \4627_b1 , \4627_b0 , \4628_b1 , \4628_b0 , \4629_b1 , \4629_b0 , 
		\4630_b1 , \4630_b0 , \4631_b1 , \4631_b0 , \4632_b1 , \4632_b0 , \4633_b1 , \4633_b0 , \4634_b1 , \4634_b0 , 
		\4635_b1 , \4635_b0 , \4636_b1 , \4636_b0 , \4637_b1 , \4637_b0 , \4638_b1 , \4638_b0 , \4639_b1 , \4639_b0 , 
		\4640_b1 , \4640_b0 , \4641_b1 , \4641_b0 , \4642_b1 , \4642_b0 , \4643_b1 , \4643_b0 , \4644_b1 , \4644_b0 , 
		\4645_b1 , \4645_b0 , \4646_b1 , \4646_b0 , \4647_b1 , \4647_b0 , \4648_b1 , \4648_b0 , \4649_b1 , \4649_b0 , 
		\4650_b1 , \4650_b0 , \4651_b1 , \4651_b0 , \4652_b1 , \4652_b0 , \4653_b1 , \4653_b0 , \4654_b1 , \4654_b0 , 
		\4655_b1 , \4655_b0 , \4656_b1 , \4656_b0 , \4657_b1 , \4657_b0 , \4658_b1 , \4658_b0 , \4659_b1 , \4659_b0 , 
		\4660_b1 , \4660_b0 , \4661_b1 , \4661_b0 , \4662_b1 , \4662_b0 , \4663_b1 , \4663_b0 , \4664_b1 , \4664_b0 , 
		\4665_b1 , \4665_b0 , \4666_b1 , \4666_b0 , \4667_b1 , \4667_b0 , \4668_b1 , \4668_b0 , \4669_b1 , \4669_b0 , 
		\4670_b1 , \4670_b0 , \4671_b1 , \4671_b0 , \4672_b1 , \4672_b0 , \4673_b1 , \4673_b0 , \4674_b1 , \4674_b0 , 
		\4675_b1 , \4675_b0 , \4676_b1 , \4676_b0 , \4677_b1 , \4677_b0 , \4678_b1 , \4678_b0 , \4679_b1 , \4679_b0 , 
		\4680_b1 , \4680_b0 , \4681_b1 , \4681_b0 , \4682_b1 , \4682_b0 , \4683_b1 , \4683_b0 , \4684_b1 , \4684_b0 , 
		\4685_b1 , \4685_b0 , \4686_b1 , \4686_b0 , \4687_b1 , \4687_b0 , \4688_b1 , \4688_b0 , \4689_b1 , \4689_b0 , 
		\4690_b1 , \4690_b0 , \4691_b1 , \4691_b0 , \4692_b1 , \4692_b0 , \4693_b1 , \4693_b0 , \4694_b1 , \4694_b0 , 
		\4695_b1 , \4695_b0 , \4696_b1 , \4696_b0 , \4697_b1 , \4697_b0 , \4698_b1 , \4698_b0 , \4699_b1 , \4699_b0 , 
		\4700_b1 , \4700_b0 , \4701_b1 , \4701_b0 , \4702_b1 , \4702_b0 , \4703_b1 , \4703_b0 , \4704_b1 , \4704_b0 , 
		\4705_b1 , \4705_b0 , \4706_b1 , \4706_b0 , \4707_b1 , \4707_b0 , \4708_b1 , \4708_b0 , \4709_b1 , \4709_b0 , 
		\4710_b1 , \4710_b0 , \4711_b1 , \4711_b0 , \4712_b1 , \4712_b0 , \4713_b1 , \4713_b0 , \4714_b1 , \4714_b0 , 
		\4715_b1 , \4715_b0 , \4716_b1 , \4716_b0 , \4717_b1 , \4717_b0 , \4718_b1 , \4718_b0 , \4719_b1 , \4719_b0 , 
		\4720_b1 , \4720_b0 , \4721_b1 , \4721_b0 , \4722_b1 , \4722_b0 , \4723_b1 , \4723_b0 , \4724_b1 , \4724_b0 , 
		\4725_b1 , \4725_b0 , \4726_b1 , \4726_b0 , \4727_b1 , \4727_b0 , \4728_b1 , \4728_b0 , \4729_b1 , \4729_b0 , 
		\4730_b1 , \4730_b0 , \4731_b1 , \4731_b0 , \4732_b1 , \4732_b0 , \4733_b1 , \4733_b0 , \4734_b1 , \4734_b0 , 
		\4735_b1 , \4735_b0 , \4736_b1 , \4736_b0 , \4737_b1 , \4737_b0 , \4738_b1 , \4738_b0 , \4739_b1 , \4739_b0 , 
		\4740_b1 , \4740_b0 , \4741_b1 , \4741_b0 , \4742_b1 , \4742_b0 , \4743_b1 , \4743_b0 , \4744_b1 , \4744_b0 , 
		\4745_b1 , \4745_b0 , \4746_b1 , \4746_b0 , \4747_b1 , \4747_b0 , \4748_b1 , \4748_b0 , \4749_b1 , \4749_b0 , 
		\4750_b1 , \4750_b0 , \4751_b1 , \4751_b0 , \4752_b1 , \4752_b0 , \4753_b1 , \4753_b0 , \4754_b1 , \4754_b0 , 
		\4755_b1 , \4755_b0 , \4756_b1 , \4756_b0 , \4757_b1 , \4757_b0 , \4758_b1 , \4758_b0 , \4759_b1 , \4759_b0 , 
		\4760_b1 , \4760_b0 , \4761_b1 , \4761_b0 , \4762_b1 , \4762_b0 , \4763_b1 , \4763_b0 , \4764_b1 , \4764_b0 , 
		\4765_b1 , \4765_b0 , \4766_b1 , \4766_b0 , \4767_b1 , \4767_b0 , \4768_b1 , \4768_b0 , \4769_b1 , \4769_b0 , 
		\4770_b1 , \4770_b0 , \4771_b1 , \4771_b0 , \4772_b1 , \4772_b0 , \4773_b1 , \4773_b0 , \4774_b1 , \4774_b0 , 
		\4775_b1 , \4775_b0 , \4776_b1 , \4776_b0 , \4777_b1 , \4777_b0 , \4778_b1 , \4778_b0 , \4779_b1 , \4779_b0 , 
		\4780_b1 , \4780_b0 , \4781_b1 , \4781_b0 , \4782_b1 , \4782_b0 , \4783_b1 , \4783_b0 , \4784_b1 , \4784_b0 , 
		\4785_b1 , \4785_b0 , \4786_b1 , \4786_b0 , \4787_b1 , \4787_b0 , \4788_b1 , \4788_b0 , \4789_b1 , \4789_b0 , 
		\4790_b1 , \4790_b0 , \4791_b1 , \4791_b0 , \4792_b1 , \4792_b0 , \4793_b1 , \4793_b0 , \4794_b1 , \4794_b0 , 
		\4795_b1 , \4795_b0 , \4796_b1 , \4796_b0 , \4797_b1 , \4797_b0 , \4798_b1 , \4798_b0 , \4799_b1 , \4799_b0 , 
		\4800_b1 , \4800_b0 , \4801_b1 , \4801_b0 , \4802_b1 , \4802_b0 , \4803_b1 , \4803_b0 , \4804_b1 , \4804_b0 , 
		\4805_b1 , \4805_b0 , \4806_b1 , \4806_b0 , \4807_b1 , \4807_b0 , \4808_b1 , \4808_b0 , \4809_b1 , \4809_b0 , 
		\4810_b1 , \4810_b0 , \4811_b1 , \4811_b0 , \4812_b1 , \4812_b0 , \4813_b1 , \4813_b0 , \4814_b1 , \4814_b0 , 
		\4815_b1 , \4815_b0 , \4816_b1 , \4816_b0 , \4817_b1 , \4817_b0 , \4818_b1 , \4818_b0 , \4819_b1 , \4819_b0 , 
		\4820_b1 , \4820_b0 , \4821_b1 , \4821_b0 , \4822_b1 , \4822_b0 , \4823_b1 , \4823_b0 , \4824_b1 , \4824_b0 , 
		\4825_b1 , \4825_b0 , \4826_b1 , \4826_b0 , \4827_b1 , \4827_b0 , \4828_b1 , \4828_b0 , \4829_b1 , \4829_b0 , 
		\4830_b1 , \4830_b0 , \4831_b1 , \4831_b0 , \4832_b1 , \4832_b0 , \4833_b1 , \4833_b0 , \4834_b1 , \4834_b0 , 
		\4835_b1 , \4835_b0 , \4836_b1 , \4836_b0 , \4837_b1 , \4837_b0 , \4838_b1 , \4838_b0 , \4839_b1 , \4839_b0 , 
		\4840_b1 , \4840_b0 , \4841_b1 , \4841_b0 , \4842_b1 , \4842_b0 , \4843_b1 , \4843_b0 , \4844_b1 , \4844_b0 , 
		\4845_b1 , \4845_b0 , \4846_b1 , \4846_b0 , \4847_b1 , \4847_b0 , \4848_b1 , \4848_b0 , \4849_b1 , \4849_b0 , 
		\4850_b1 , \4850_b0 , \4851_b1 , \4851_b0 , \4852_b1 , \4852_b0 , \4853_b1 , \4853_b0 , \4854_b1 , \4854_b0 , 
		\4855_b1 , \4855_b0 , \4856_b1 , \4856_b0 , \4857_b1 , \4857_b0 , \4858_b1 , \4858_b0 , \4859_b1 , \4859_b0 , 
		\4860_b1 , \4860_b0 , \4861_b1 , \4861_b0 , \4862_b1 , \4862_b0 , \4863_b1 , \4863_b0 , \4864_b1 , \4864_b0 , 
		\4865_b1 , \4865_b0 , \4866_b1 , \4866_b0 , \4867_b1 , \4867_b0 , \4868_b1 , \4868_b0 , \4869_b1 , \4869_b0 , 
		\4870_b1 , \4870_b0 , \4871_b1 , \4871_b0 , \4872_b1 , \4872_b0 , \4873_b1 , \4873_b0 , \4874_b1 , \4874_b0 , 
		\4875_b1 , \4875_b0 , \4876_b1 , \4876_b0 , \4877_b1 , \4877_b0 , \4878_b1 , \4878_b0 , \4879_b1 , \4879_b0 , 
		\4880_b1 , \4880_b0 , \4881_b1 , \4881_b0 , \4882_b1 , \4882_b0 , \4883_b1 , \4883_b0 , \4884_b1 , \4884_b0 , 
		\4885_b1 , \4885_b0 , \4886_b1 , \4886_b0 , \4887_b1 , \4887_b0 , \4888_b1 , \4888_b0 , \4889_b1 , \4889_b0 , 
		\4890_b1 , \4890_b0 , \4891_b1 , \4891_b0 , \4892_b1 , \4892_b0 , \4893_b1 , \4893_b0 , \4894_b1 , \4894_b0 , 
		\4895_b1 , \4895_b0 , \4896_b1 , \4896_b0 , \4897_b1 , \4897_b0 , \4898_b1 , \4898_b0 , \4899_b1 , \4899_b0 , 
		\4900_b1 , \4900_b0 , \4901_b1 , \4901_b0 , \4902_b1 , \4902_b0 , \4903_b1 , \4903_b0 , \4904_b1 , \4904_b0 , 
		\4905_b1 , \4905_b0 , \4906_b1 , \4906_b0 , \4907_b1 , \4907_b0 , \4908_b1 , \4908_b0 , \4909_b1 , \4909_b0 , 
		\4910_b1 , \4910_b0 , \4911_b1 , \4911_b0 , \4912_b1 , \4912_b0 , \4913_b1 , \4913_b0 , \4914_b1 , \4914_b0 , 
		\4915_b1 , \4915_b0 , \4916_b1 , \4916_b0 , \4917_b1 , \4917_b0 , \4918_b1 , \4918_b0 , \4919_b1 , \4919_b0 , 
		\4920_b1 , \4920_b0 , \4921_b1 , \4921_b0 , \4922_b1 , \4922_b0 , \4923_b1 , \4923_b0 , \4924_b1 , \4924_b0 , 
		\4925_b1 , \4925_b0 , \4926_b1 , \4926_b0 , \4927_b1 , \4927_b0 , \4928_b1 , \4928_b0 , \4929_b1 , \4929_b0 , 
		\4930_b1 , \4930_b0 , \4931_b1 , \4931_b0 , \4932_b1 , \4932_b0 , \4933_b1 , \4933_b0 , \4934_b1 , \4934_b0 , 
		\4935_b1 , \4935_b0 , \4936_b1 , \4936_b0 , \4937_b1 , \4937_b0 , \4938_b1 , \4938_b0 , \4939_b1 , \4939_b0 , 
		\4940_b1 , \4940_b0 , \4941_b1 , \4941_b0 , \4942_b1 , \4942_b0 , \4943_b1 , \4943_b0 , \4944_b1 , \4944_b0 , 
		\4945_b1 , \4945_b0 , \4946_b1 , \4946_b0 , \4947_b1 , \4947_b0 , \4948_b1 , \4948_b0 , \4949_b1 , \4949_b0 , 
		\4950_b1 , \4950_b0 , \4951_b1 , \4951_b0 , \4952_b1 , \4952_b0 , \4953_b1 , \4953_b0 , \4954_b1 , \4954_b0 , 
		\4955_b1 , \4955_b0 , \4956_b1 , \4956_b0 , \4957_b1 , \4957_b0 , \4958_b1 , \4958_b0 , \4959_b1 , \4959_b0 , 
		\4960_b1 , \4960_b0 , \4961_b1 , \4961_b0 , \4962_b1 , \4962_b0 , \4963_b1 , \4963_b0 , \4964_b1 , \4964_b0 , 
		\4965_b1 , \4965_b0 , \4966_b1 , \4966_b0 , \4967_b1 , \4967_b0 , \4968_b1 , \4968_b0 , \4969_b1 , \4969_b0 , 
		\4970_b1 , \4970_b0 , \4971_b1 , \4971_b0 , \4972_b1 , \4972_b0 , \4973_b1 , \4973_b0 , \4974_b1 , \4974_b0 , 
		\4975_b1 , \4975_b0 , \4976_b1 , \4976_b0 , \4977_b1 , \4977_b0 , \4978_b1 , \4978_b0 , \4979_b1 , \4979_b0 , 
		\4980_b1 , \4980_b0 , \4981_b1 , \4981_b0 , \4982_b1 , \4982_b0 , \4983_b1 , \4983_b0 , \4984_b1 , \4984_b0 , 
		\4985_b1 , \4985_b0 , \4986_b1 , \4986_b0 , \4987_b1 , \4987_b0 , \4988_b1 , \4988_b0 , \4989_b1 , \4989_b0 , 
		\4990_b1 , \4990_b0 , \4991_b1 , \4991_b0 , \4992_b1 , \4992_b0 , \4993_b1 , \4993_b0 , \4994_b1 , \4994_b0 , 
		\4995_b1 , \4995_b0 , \4996_b1 , \4996_b0 , \4997_b1 , \4997_b0 , \4998_b1 , \4998_b0 , \4999_b1 , \4999_b0 , 
		\5000_b1 , \5000_b0 , \5001_b1 , \5001_b0 , \5002_b1 , \5002_b0 , \5003_b1 , \5003_b0 , \5004_b1 , \5004_b0 , 
		\5005_b1 , \5005_b0 , \5006_b1 , \5006_b0 , \5007_b1 , \5007_b0 , \5008_b1 , \5008_b0 , \5009_b1 , \5009_b0 , 
		\5010_b1 , \5010_b0 , \5011_b1 , \5011_b0 , \5012_b1 , \5012_b0 , \5013_b1 , \5013_b0 , \5014_b1 , \5014_b0 , 
		\5015_b1 , \5015_b0 , \5016_b1 , \5016_b0 , \5017_b1 , \5017_b0 , \5018_b1 , \5018_b0 , \5019_b1 , \5019_b0 , 
		\5020_b1 , \5020_b0 , \5021_b1 , \5021_b0 , \5022_b1 , \5022_b0 , \5023_b1 , \5023_b0 , \5024_b1 , \5024_b0 , 
		\5025_b1 , \5025_b0 , \5026_b1 , \5026_b0 , \5027_b1 , \5027_b0 , \5028_b1 , \5028_b0 , \5029_b1 , \5029_b0 , 
		\5030_b1 , \5030_b0 , \5031_b1 , \5031_b0 , \5032_b1 , \5032_b0 , \5033_b1 , \5033_b0 , \5034_b1 , \5034_b0 , 
		\5035_b1 , \5035_b0 , \5036_b1 , \5036_b0 , \5037_b1 , \5037_b0 , \5038_b1 , \5038_b0 , \5039_b1 , \5039_b0 , 
		\5040_b1 , \5040_b0 , \5041_b1 , \5041_b0 , \5042_b1 , \5042_b0 , \5043_b1 , \5043_b0 , \5044_b1 , \5044_b0 , 
		\5045_b1 , \5045_b0 , \5046_b1 , \5046_b0 , \5047_b1 , \5047_b0 , \5048_b1 , \5048_b0 , \5049_b1 , \5049_b0 , 
		\5050_b1 , \5050_b0 , \5051_b1 , \5051_b0 , \5052_b1 , \5052_b0 , \5053_b1 , \5053_b0 , \5054_b1 , \5054_b0 , 
		\5055_b1 , \5055_b0 , \5056_b1 , \5056_b0 , \5057_b1 , \5057_b0 , \5058_b1 , \5058_b0 , \5059_b1 , \5059_b0 , 
		\5060_b1 , \5060_b0 , \5061_b1 , \5061_b0 , \5062_b1 , \5062_b0 , \5063_b1 , \5063_b0 , \5064_b1 , \5064_b0 , 
		\5065_b1 , \5065_b0 , \5066_b1 , \5066_b0 , \5067_b1 , \5067_b0 , \5068_b1 , \5068_b0 , \5069_b1 , \5069_b0 , 
		\5070_b1 , \5070_b0 , \5071_b1 , \5071_b0 , \5072_b1 , \5072_b0 , \5073_b1 , \5073_b0 , \5074_b1 , \5074_b0 , 
		\5075_b1 , \5075_b0 , \5076_b1 , \5076_b0 , \5077_b1 , \5077_b0 , \5078_b1 , \5078_b0 , \5079_b1 , \5079_b0 , 
		\5080_b1 , \5080_b0 , \5081_b1 , \5081_b0 , \5082_b1 , \5082_b0 , \5083_b1 , \5083_b0 , \5084_b1 , \5084_b0 , 
		\5085_b1 , \5085_b0 , \5086_b1 , \5086_b0 , \5087_b1 , \5087_b0 , \5088_b1 , \5088_b0 , \5089_b1 , \5089_b0 , 
		\5090_b1 , \5090_b0 , \5091_b1 , \5091_b0 , \5092_b1 , \5092_b0 , \5093_b1 , \5093_b0 , \5094_b1 , \5094_b0 , 
		\5095_b1 , \5095_b0 , \5096_b1 , \5096_b0 , \5097_b1 , \5097_b0 , \5098_b1 , \5098_b0 , \5099_b1 , \5099_b0 , 
		\5100_b1 , \5100_b0 , \5101_b1 , \5101_b0 , \5102_b1 , \5102_b0 , \5103_b1 , \5103_b0 , \5104_b1 , \5104_b0 , 
		\5105_b1 , \5105_b0 , \5106_b1 , \5106_b0 , \5107_b1 , \5107_b0 , \5108_b1 , \5108_b0 , \5109_b1 , \5109_b0 , 
		\5110_b1 , \5110_b0 , \5111_b1 , \5111_b0 , \5112_b1 , \5112_b0 , \5113_b1 , \5113_b0 , \5114_b1 , \5114_b0 , 
		\5115_b1 , \5115_b0 , \5116_b1 , \5116_b0 , \5117_b1 , \5117_b0 , \5118_b1 , \5118_b0 , \5119_b1 , \5119_b0 , 
		\5120_b1 , \5120_b0 , \5121_b1 , \5121_b0 , \5122_b1 , \5122_b0 , \5123_b1 , \5123_b0 , \5124_b1 , \5124_b0 , 
		\5125_b1 , \5125_b0 , \5126_b1 , \5126_b0 , \5127_b1 , \5127_b0 , \5128_b1 , \5128_b0 , \5129_b1 , \5129_b0 , 
		\5130_b1 , \5130_b0 , \5131_b1 , \5131_b0 , \5132_b1 , \5132_b0 , \5133_b1 , \5133_b0 , \5134_b1 , \5134_b0 , 
		\5135_b1 , \5135_b0 , \5136_b1 , \5136_b0 , \5137_b1 , \5137_b0 , \5138_b1 , \5138_b0 , \5139_b1 , \5139_b0 , 
		\5140_b1 , \5140_b0 , \5141_b1 , \5141_b0 , \5142_b1 , \5142_b0 , \5143_b1 , \5143_b0 , \5144_b1 , \5144_b0 , 
		\5145_b1 , \5145_b0 , \5146_b1 , \5146_b0 , \5147_b1 , \5147_b0 , \5148_b1 , \5148_b0 , \5149_b1 , \5149_b0 , 
		\5150_b1 , \5150_b0 , \5151_b1 , \5151_b0 , \5152_b1 , \5152_b0 , \5153_b1 , \5153_b0 , \5154_b1 , \5154_b0 , 
		\5155_b1 , \5155_b0 , \5156_b1 , \5156_b0 , \5157_b1 , \5157_b0 , \5158_b1 , \5158_b0 , \5159_b1 , \5159_b0 , 
		\5160_b1 , \5160_b0 , \5161_b1 , \5161_b0 , \5162_b1 , \5162_b0 , \5163_b1 , \5163_b0 , \5164_b1 , \5164_b0 , 
		\5165_b1 , \5165_b0 , \5166_b1 , \5166_b0 , \5167_b1 , \5167_b0 , \5168_b1 , \5168_b0 , \5169_b1 , \5169_b0 , 
		\5170_b1 , \5170_b0 , \5171_b1 , \5171_b0 , \5172_b1 , \5172_b0 , \5173_b1 , \5173_b0 , \5174_b1 , \5174_b0 , 
		\5175_b1 , \5175_b0 , \5176_b1 , \5176_b0 , \5177_b1 , \5177_b0 , \5178_b1 , \5178_b0 , \5179_b1 , \5179_b0 , 
		\5180_b1 , \5180_b0 , \5181_b1 , \5181_b0 , \5182_b1 , \5182_b0 , \5183_b1 , \5183_b0 , \5184_b1 , \5184_b0 , 
		\5185_b1 , \5185_b0 , \5186_b1 , \5186_b0 , \5187_b1 , \5187_b0 , \5188_b1 , \5188_b0 , \5189_b1 , \5189_b0 , 
		\5190_b1 , \5190_b0 , \5191_b1 , \5191_b0 , \5192_b1 , \5192_b0 , \5193_b1 , \5193_b0 , \5194_b1 , \5194_b0 , 
		\5195_b1 , \5195_b0 , \5196_b1 , \5196_b0 , \5197_b1 , \5197_b0 , \5198_b1 , \5198_b0 , \5199_b1 , \5199_b0 , 
		\5200_b1 , \5200_b0 , \5201_b1 , \5201_b0 , \5202_b1 , \5202_b0 , \5203_b1 , \5203_b0 , \5204_b1 , \5204_b0 , 
		\5205_b1 , \5205_b0 , \5206_b1 , \5206_b0 , \5207_b1 , \5207_b0 , \5208_b1 , \5208_b0 , \5209_b1 , \5209_b0 , 
		\5210_b1 , \5210_b0 , \5211_b1 , \5211_b0 , \5212_b1 , \5212_b0 , \5213_b1 , \5213_b0 , \5214_b1 , \5214_b0 , 
		\5215_b1 , \5215_b0 , \5216_b1 , \5216_b0 , \5217_b1 , \5217_b0 , \5218_b1 , \5218_b0 , \5219_b1 , \5219_b0 , 
		\5220_b1 , \5220_b0 , \5221_b1 , \5221_b0 , \5222_b1 , \5222_b0 , \5223_b1 , \5223_b0 , \5224_b1 , \5224_b0 , 
		\5225_b1 , \5225_b0 , \5226_b1 , \5226_b0 , \5227_b1 , \5227_b0 , \5228_b1 , \5228_b0 , \5229_b1 , \5229_b0 , 
		\5230_b1 , \5230_b0 , \5231_b1 , \5231_b0 , \5232_b1 , \5232_b0 , \5233_b1 , \5233_b0 , \5234_b1 , \5234_b0 , 
		\5235_b1 , \5235_b0 , \5236_b1 , \5236_b0 , \5237_b1 , \5237_b0 , \5238_b1 , \5238_b0 , \5239_b1 , \5239_b0 , 
		\5240_b1 , \5240_b0 , \5241_b1 , \5241_b0 , \5242_b1 , \5242_b0 , \5243_b1 , \5243_b0 , \5244_b1 , \5244_b0 , 
		\5245_b1 , \5245_b0 , \5246_b1 , \5246_b0 , \5247_b1 , \5247_b0 , \5248_b1 , \5248_b0 , \5249_b1 , \5249_b0 , 
		\5250_b1 , \5250_b0 , \5251_b1 , \5251_b0 , \5252_b1 , \5252_b0 , \5253_b1 , \5253_b0 , \5254_b1 , \5254_b0 , 
		\5255_b1 , \5255_b0 , \5256_b1 , \5256_b0 , \5257_b1 , \5257_b0 , \5258_b1 , \5258_b0 , \5259_b1 , \5259_b0 , 
		\5260_b1 , \5260_b0 , \5261_b1 , \5261_b0 , \5262_b1 , \5262_b0 , \5263_b1 , \5263_b0 , \5264_b1 , \5264_b0 , 
		\5265_b1 , \5265_b0 , \5266_b1 , \5266_b0 , \5267_b1 , \5267_b0 , \5268_b1 , \5268_b0 , \5269_b1 , \5269_b0 , 
		\5270_b1 , \5270_b0 , \5271_b1 , \5271_b0 , \5272_b1 , \5272_b0 , \5273_b1 , \5273_b0 , \5274_b1 , \5274_b0 , 
		\5275_b1 , \5275_b0 , \5276_b1 , \5276_b0 , \5277_b1 , \5277_b0 , \5278_b1 , \5278_b0 , \5279_b1 , \5279_b0 , 
		\5280_b1 , \5280_b0 , \5281_b1 , \5281_b0 , \5282_b1 , \5282_b0 , \5283_b1 , \5283_b0 , \5284_b1 , \5284_b0 , 
		\5285_b1 , \5285_b0 , \5286_b1 , \5286_b0 , \5287_b1 , \5287_b0 , \5288_b1 , \5288_b0 , \5289_b1 , \5289_b0 , 
		\5290_b1 , \5290_b0 , \5291_b1 , \5291_b0 , \5292_b1 , \5292_b0 , \5293_b1 , \5293_b0 , \5294_b1 , \5294_b0 , 
		\5295_b1 , \5295_b0 , \5296_b1 , \5296_b0 , \5297_b1 , \5297_b0 , \5298_b1 , \5298_b0 , \5299_b1 , \5299_b0 , 
		\5300_b1 , \5300_b0 , \5301_b1 , \5301_b0 , \5302_b1 , \5302_b0 , \5303_b1 , \5303_b0 , \5304_b1 , \5304_b0 , 
		\5305_b1 , \5305_b0 , \5306_b1 , \5306_b0 , \5307_b1 , \5307_b0 , \5308_b1 , \5308_b0 , \5309_b1 , \5309_b0 , 
		\5310_b1 , \5310_b0 , \5311_b1 , \5311_b0 , \5312_b1 , \5312_b0 , \5313_b1 , \5313_b0 , \5314_b1 , \5314_b0 , 
		\5315_b1 , \5315_b0 , \5316_b1 , \5316_b0 , \5317_b1 , \5317_b0 , \5318_b1 , \5318_b0 , \5319_b1 , \5319_b0 , 
		\5320_b1 , \5320_b0 , \5321_b1 , \5321_b0 , \5322_b1 , \5322_b0 , \5323_b1 , \5323_b0 , \5324_b1 , \5324_b0 , 
		\5325_b1 , \5325_b0 , \5326_b1 , \5326_b0 , \5327_b1 , \5327_b0 , \5328_b1 , \5328_b0 , \5329_b1 , \5329_b0 , 
		\5330_b1 , \5330_b0 , \5331_b1 , \5331_b0 , \5332_b1 , \5332_b0 , \5333_b1 , \5333_b0 , \5334_b1 , \5334_b0 , 
		\5335_b1 , \5335_b0 , \5336_b1 , \5336_b0 , \5337_b1 , \5337_b0 , \5338_b1 , \5338_b0 , \5339_b1 , \5339_b0 , 
		\5340_b1 , \5340_b0 , \5341_b1 , \5341_b0 , \5342_b1 , \5342_b0 , \5343_b1 , \5343_b0 , \5344_b1 , \5344_b0 , 
		\5345_b1 , \5345_b0 , \5346_b1 , \5346_b0 , \5347_b1 , \5347_b0 , \5348_b1 , \5348_b0 , \5349_b1 , \5349_b0 , 
		\5350_b1 , \5350_b0 , \5351_b1 , \5351_b0 , \5352_b1 , \5352_b0 , \5353_b1 , \5353_b0 , \5354_b1 , \5354_b0 , 
		\5355_b1 , \5355_b0 , \5356_b1 , \5356_b0 , \5357_b1 , \5357_b0 , \5358_b1 , \5358_b0 , \5359_b1 , \5359_b0 , 
		\5360_b1 , \5360_b0 , \5361_b1 , \5361_b0 , \5362_b1 , \5362_b0 , \5363_b1 , \5363_b0 , \5364_b1 , \5364_b0 , 
		\5365_b1 , \5365_b0 , \5366_b1 , \5366_b0 , \5367_b1 , \5367_b0 , \5368_b1 , \5368_b0 , \5369_b1 , \5369_b0 , 
		\5370_b1 , \5370_b0 , \5371_b1 , \5371_b0 , \5372_b1 , \5372_b0 , \5373_b1 , \5373_b0 , \5374_b1 , \5374_b0 , 
		\5375_b1 , \5375_b0 , \5376_b1 , \5376_b0 , \5377_b1 , \5377_b0 , \5378_b1 , \5378_b0 , \5379_b1 , \5379_b0 , 
		\5380_b1 , \5380_b0 , \5381_b1 , \5381_b0 , \5382_b1 , \5382_b0 , \5383_b1 , \5383_b0 , \5384_b1 , \5384_b0 , 
		\5385_b1 , \5385_b0 , \5386_b1 , \5386_b0 , \5387_b1 , \5387_b0 , \5388_b1 , \5388_b0 , \5389_b1 , \5389_b0 , 
		\5390_b1 , \5390_b0 , \5391_b1 , \5391_b0 , \5392_b1 , \5392_b0 , \5393_b1 , \5393_b0 , \5394_b1 , \5394_b0 , 
		\5395_b1 , \5395_b0 , \5396_b1 , \5396_b0 , \5397_b1 , \5397_b0 , \5398_b1 , \5398_b0 , \5399_b1 , \5399_b0 , 
		\5400_b1 , \5400_b0 , \5401_b1 , \5401_b0 , \5402_b1 , \5402_b0 , \5403_b1 , \5403_b0 , \5404_b1 , \5404_b0 , 
		\5405_b1 , \5405_b0 , \5406_b1 , \5406_b0 , \5407_b1 , \5407_b0 , \5408_b1 , \5408_b0 , \5409_b1 , \5409_b0 , 
		\5410_b1 , \5410_b0 , \5411_b1 , \5411_b0 , \5412_b1 , \5412_b0 , \5413_b1 , \5413_b0 , \5414_b1 , \5414_b0 , 
		\5415_b1 , \5415_b0 , \5416_b1 , \5416_b0 , \5417_b1 , \5417_b0 , \5418_b1 , \5418_b0 , \5419_b1 , \5419_b0 , 
		\5420_b1 , \5420_b0 , \5421_b1 , \5421_b0 , \5422_b1 , \5422_b0 , \5423_b1 , \5423_b0 , \5424_b1 , \5424_b0 , 
		\5425_b1 , \5425_b0 , \5426_b1 , \5426_b0 , \5427_b1 , \5427_b0 , \5428_b1 , \5428_b0 , \5429_b1 , \5429_b0 , 
		\5430_b1 , \5430_b0 , \5431_b1 , \5431_b0 , \5432_b1 , \5432_b0 , \5433_b1 , \5433_b0 , \5434_b1 , \5434_b0 , 
		\5435_b1 , \5435_b0 , \5436_b1 , \5436_b0 , \5437_b1 , \5437_b0 , \5438_b1 , \5438_b0 , \5439_b1 , \5439_b0 , 
		\5440_b1 , \5440_b0 , \5441_b1 , \5441_b0 , \5442_b1 , \5442_b0 , \5443_b1 , \5443_b0 , \5444_b1 , \5444_b0 , 
		\5445_b1 , \5445_b0 , \5446_b1 , \5446_b0 , \5447_b1 , \5447_b0 , \5448_b1 , \5448_b0 , \5449_b1 , \5449_b0 , 
		\5450_b1 , \5450_b0 , \5451_b1 , \5451_b0 , \5452_b1 , \5452_b0 , \5453_b1 , \5453_b0 , \5454_b1 , \5454_b0 , 
		\5455_b1 , \5455_b0 , \5456_b1 , \5456_b0 , \5457_b1 , \5457_b0 , \5458_b1 , \5458_b0 , \5459_b1 , \5459_b0 , 
		\5460_b1 , \5460_b0 , \5461_b1 , \5461_b0 , \5462_b1 , \5462_b0 , \5463_b1 , \5463_b0 , \5464_b1 , \5464_b0 , 
		\5465_b1 , \5465_b0 , \5466_b1 , \5466_b0 , \5467_b1 , \5467_b0 , \5468_b1 , \5468_b0 , \5469_b1 , \5469_b0 , 
		\5470_b1 , \5470_b0 , \5471_b1 , \5471_b0 , \5472_b1 , \5472_b0 , \5473_b1 , \5473_b0 , \5474_b1 , \5474_b0 , 
		\5475_b1 , \5475_b0 , \5476_b1 , \5476_b0 , \5477_b1 , \5477_b0 , \5478_b1 , \5478_b0 , \5479_b1 , \5479_b0 , 
		\5480_b1 , \5480_b0 , \5481_b1 , \5481_b0 , \5482_b1 , \5482_b0 , \5483_b1 , \5483_b0 , \5484_b1 , \5484_b0 , 
		\5485_b1 , \5485_b0 , \5486_b1 , \5486_b0 , \5487_b1 , \5487_b0 , \5488_b1 , \5488_b0 , \5489_b1 , \5489_b0 , 
		\5490_b1 , \5490_b0 , \5491_b1 , \5491_b0 , \5492_b1 , \5492_b0 , \5493_b1 , \5493_b0 , \5494_b1 , \5494_b0 , 
		\5495_b1 , \5495_b0 , \5496_b1 , \5496_b0 , \5497_b1 , \5497_b0 , \5498_b1 , \5498_b0 , \5499_b1 , \5499_b0 , 
		\5500_b1 , \5500_b0 , \5501_b1 , \5501_b0 , \5502_b1 , \5502_b0 , \5503_b1 , \5503_b0 , \5504_b1 , \5504_b0 , 
		\5505_b1 , \5505_b0 , \5506_b1 , \5506_b0 , \5507_b1 , \5507_b0 , \5508_b1 , \5508_b0 , \5509_b1 , \5509_b0 , 
		\5510_b1 , \5510_b0 , \5511_b1 , \5511_b0 , \5512_b1 , \5512_b0 , \5513_b1 , \5513_b0 , \5514_b1 , \5514_b0 , 
		\5515_b1 , \5515_b0 , \5516_b1 , \5516_b0 , \5517_b1 , \5517_b0 , \5518_b1 , \5518_b0 , \5519_b1 , \5519_b0 , 
		\5520_b1 , \5520_b0 , \5521_b1 , \5521_b0 , \5522_b1 , \5522_b0 , \5523_b1 , \5523_b0 , \5524_b1 , \5524_b0 , 
		\5525_b1 , \5525_b0 , \5526_b1 , \5526_b0 , \5527_b1 , \5527_b0 , \5528_b1 , \5528_b0 , \5529_b1 , \5529_b0 , 
		\5530_b1 , \5530_b0 , \5531_b1 , \5531_b0 , \5532_b1 , \5532_b0 , \5533_b1 , \5533_b0 , \5534_b1 , \5534_b0 , 
		\5535_b1 , \5535_b0 , \5536_b1 , \5536_b0 , \5537_b1 , \5537_b0 , \5538_b1 , \5538_b0 , \5539_b1 , \5539_b0 , 
		\5540_b1 , \5540_b0 , \5541_b1 , \5541_b0 , \5542_b1 , \5542_b0 , \5543_b1 , \5543_b0 , \5544_b1 , \5544_b0 , 
		\5545_b1 , \5545_b0 , \5546_b1 , \5546_b0 , \5547_b1 , \5547_b0 , \5548_b1 , \5548_b0 , \5549_b1 , \5549_b0 , 
		\5550_b1 , \5550_b0 , \5551_b1 , \5551_b0 , \5552_b1 , \5552_b0 , \5553_b1 , \5553_b0 , \5554_b1 , \5554_b0 , 
		\5555_b1 , \5555_b0 , \5556_b1 , \5556_b0 , \5557_b1 , \5557_b0 , \5558_b1 , \5558_b0 , \5559_b1 , \5559_b0 , 
		\5560_b1 , \5560_b0 , \5561_b1 , \5561_b0 , \5562_b1 , \5562_b0 , \5563_b1 , \5563_b0 , \5564_b1 , \5564_b0 , 
		\5565_b1 , \5565_b0 , \5566_b1 , \5566_b0 , \5567_b1 , \5567_b0 , \5568_b1 , \5568_b0 , \5569_b1 , \5569_b0 , 
		\5570_b1 , \5570_b0 , \5571_b1 , \5571_b0 , \5572_b1 , \5572_b0 , \5573_b1 , \5573_b0 , \5574_b1 , \5574_b0 , 
		\5575_b1 , \5575_b0 , \5576_b1 , \5576_b0 , \5577_b1 , \5577_b0 , \5578_b1 , \5578_b0 , \5579_b1 , \5579_b0 , 
		\5580_b1 , \5580_b0 , \5581_b1 , \5581_b0 , \5582_b1 , \5582_b0 , \5583_b1 , \5583_b0 , \5584_b1 , \5584_b0 , 
		\5585_b1 , \5585_b0 , \5586_b1 , \5586_b0 , \5587_b1 , \5587_b0 , \5588_b1 , \5588_b0 , \5589_b1 , \5589_b0 , 
		\5590_b1 , \5590_b0 , \5591_b1 , \5591_b0 , \5592_b1 , \5592_b0 , \5593_b1 , \5593_b0 , \5594_b1 , \5594_b0 , 
		\5595_b1 , \5595_b0 , \5596_b1 , \5596_b0 , \5597_b1 , \5597_b0 , \5598_b1 , \5598_b0 , \5599_b1 , \5599_b0 , 
		\5600_b1 , \5600_b0 , \5601_b1 , \5601_b0 , \5602_b1 , \5602_b0 , \5603_b1 , \5603_b0 , \5604_b1 , \5604_b0 , 
		\5605_b1 , \5605_b0 , \5606_b1 , \5606_b0 , \5607_b1 , \5607_b0 , \5608_b1 , \5608_b0 , \5609_b1 , \5609_b0 , 
		\5610_b1 , \5610_b0 , \5611_b1 , \5611_b0 , \5612_b1 , \5612_b0 , \5613_b1 , \5613_b0 , \5614_b1 , \5614_b0 , 
		\5615_b1 , \5615_b0 , \5616_b1 , \5616_b0 , \5617_b1 , \5617_b0 , \5618_b1 , \5618_b0 , \5619_b1 , \5619_b0 , 
		\5620_b1 , \5620_b0 , \5621_b1 , \5621_b0 , \5622_b1 , \5622_b0 , \5623_b1 , \5623_b0 , \5624_b1 , \5624_b0 , 
		\5625_b1 , \5625_b0 , \5626_b1 , \5626_b0 , \5627_b1 , \5627_b0 , \5628_b1 , \5628_b0 , \5629_b1 , \5629_b0 , 
		\5630_b1 , \5630_b0 , \5631_b1 , \5631_b0 , \5632_b1 , \5632_b0 , \5633_b1 , \5633_b0 , \5634_b1 , \5634_b0 , 
		\5635_b1 , \5635_b0 , \5636_b1 , \5636_b0 , \5637_b1 , \5637_b0 , \5638_b1 , \5638_b0 , \5639_b1 , \5639_b0 , 
		\5640_b1 , \5640_b0 , \5641_b1 , \5641_b0 , \5642_b1 , \5642_b0 , \5643_b1 , \5643_b0 , \5644_b1 , \5644_b0 , 
		\5645_b1 , \5645_b0 , \5646_b1 , \5646_b0 , \5647_b1 , \5647_b0 , \5648_b1 , \5648_b0 , \5649_b1 , \5649_b0 , 
		\5650_b1 , \5650_b0 , \5651_b1 , \5651_b0 , \5652_b1 , \5652_b0 , \5653_b1 , \5653_b0 , \5654_b1 , \5654_b0 , 
		\5655_b1 , \5655_b0 , \5656_b1 , \5656_b0 , \5657_b1 , \5657_b0 , \5658_b1 , \5658_b0 , \5659_b1 , \5659_b0 , 
		\5660_b1 , \5660_b0 , \5661_b1 , \5661_b0 , \5662_b1 , \5662_b0 , \5663_b1 , \5663_b0 , \5664_b1 , \5664_b0 , 
		\5665_b1 , \5665_b0 , \5666_b1 , \5666_b0 , \5667_b1 , \5667_b0 , \5668_b1 , \5668_b0 , \5669_b1 , \5669_b0 , 
		\5670_b1 , \5670_b0 , \5671_b1 , \5671_b0 , \5672_b1 , \5672_b0 , \5673_b1 , \5673_b0 , \5674_b1 , \5674_b0 , 
		\5675_b1 , \5675_b0 , \5676_b1 , \5676_b0 , \5677_b1 , \5677_b0 , \5678_b1 , \5678_b0 , \5679_b1 , \5679_b0 , 
		\5680_b1 , \5680_b0 , \5681_b1 , \5681_b0 , \5682_b1 , \5682_b0 , \5683_b1 , \5683_b0 , \5684_b1 , \5684_b0 , 
		\5685_b1 , \5685_b0 , \5686_b1 , \5686_b0 , \5687_b1 , \5687_b0 , \5688_b1 , \5688_b0 , \5689_b1 , \5689_b0 , 
		\5690_b1 , \5690_b0 , \5691_b1 , \5691_b0 , \5692_b1 , \5692_b0 , \5693_b1 , \5693_b0 , \5694_b1 , \5694_b0 , 
		\5695_b1 , \5695_b0 , \5696_b1 , \5696_b0 , \5697_b1 , \5697_b0 , \5698_b1 , \5698_b0 , \5699_b1 , \5699_b0 , 
		\5700_b1 , \5700_b0 , \5701_b1 , \5701_b0 , \5702_b1 , \5702_b0 , \5703_b1 , \5703_b0 , \5704_b1 , \5704_b0 , 
		\5705_b1 , \5705_b0 , \5706_b1 , \5706_b0 , \5707_b1 , \5707_b0 , \5708_b1 , \5708_b0 , \5709_b1 , \5709_b0 , 
		\5710_b1 , \5710_b0 , \5711_b1 , \5711_b0 , \5712_b1 , \5712_b0 , \5713_b1 , \5713_b0 , \5714_b1 , \5714_b0 , 
		\5715_b1 , \5715_b0 , \5716_b1 , \5716_b0 , \5717_b1 , \5717_b0 , \5718_b1 , \5718_b0 , \5719_b1 , \5719_b0 , 
		\5720_b1 , \5720_b0 , \5721_b1 , \5721_b0 , \5722_b1 , \5722_b0 , \5723_b1 , \5723_b0 , \5724_b1 , \5724_b0 , 
		\5725_b1 , \5725_b0 , \5726_b1 , \5726_b0 , \5727_b1 , \5727_b0 , \5728_b1 , \5728_b0 , \5729_b1 , \5729_b0 , 
		\5730_b1 , \5730_b0 , \5731_b1 , \5731_b0 , \5732_b1 , \5732_b0 , \5733_b1 , \5733_b0 , \5734_b1 , \5734_b0 , 
		\5735_b1 , \5735_b0 , \5736_b1 , \5736_b0 , \5737_b1 , \5737_b0 , \5738_b1 , \5738_b0 , \5739_b1 , \5739_b0 , 
		\5740_b1 , \5740_b0 , \5741_b1 , \5741_b0 , \5742_b1 , \5742_b0 , \5743_b1 , \5743_b0 , \5744_b1 , \5744_b0 , 
		\5745_b1 , \5745_b0 , \5746_b1 , \5746_b0 , \5747_b1 , \5747_b0 , \5748_b1 , \5748_b0 , \5749_b1 , \5749_b0 , 
		\5750_b1 , \5750_b0 , \5751_b1 , \5751_b0 , \5752_b1 , \5752_b0 , \5753_b1 , \5753_b0 , \5754_b1 , \5754_b0 , 
		\5755_b1 , \5755_b0 , \5756_b1 , \5756_b0 , \5757_b1 , \5757_b0 , \5758_b1 , \5758_b0 , \5759_b1 , \5759_b0 , 
		\5760_b1 , \5760_b0 , \5761_b1 , \5761_b0 , \5762_b1 , \5762_b0 , \5763_b1 , \5763_b0 , \5764_b1 , \5764_b0 , 
		\5765_b1 , \5765_b0 , \5766_b1 , \5766_b0 , \5767_b1 , \5767_b0 , \5768_b1 , \5768_b0 , \5769_b1 , \5769_b0 , 
		\5770_b1 , \5770_b0 , \5771_b1 , \5771_b0 , \5772_b1 , \5772_b0 , \5773_b1 , \5773_b0 , \5774_b1 , \5774_b0 , 
		\5775_b1 , \5775_b0 , \5776_b1 , \5776_b0 , \5777_b1 , \5777_b0 , \5778_b1 , \5778_b0 , \5779_b1 , \5779_b0 , 
		\5780_b1 , \5780_b0 , \5781_b1 , \5781_b0 , \5782_b1 , \5782_b0 , \5783_b1 , \5783_b0 , \5784_b1 , \5784_b0 , 
		\5785_b1 , \5785_b0 , \5786_b1 , \5786_b0 , \5787_b1 , \5787_b0 , \5788_b1 , \5788_b0 , \5789_b1 , \5789_b0 , 
		\5790_b1 , \5790_b0 , \5791_b1 , \5791_b0 , \5792_b1 , \5792_b0 , \5793_b1 , \5793_b0 , \5794_b1 , \5794_b0 , 
		\5795_b1 , \5795_b0 , \5796_b1 , \5796_b0 , \5797_b1 , \5797_b0 , \5798_b1 , \5798_b0 , \5799_b1 , \5799_b0 , 
		\5800_b1 , \5800_b0 , \5801_b1 , \5801_b0 , \5802_b1 , \5802_b0 , \5803_b1 , \5803_b0 , \5804_b1 , \5804_b0 , 
		\5805_b1 , \5805_b0 , \5806_b1 , \5806_b0 , \5807_b1 , \5807_b0 , \5808_b1 , \5808_b0 , \5809_b1 , \5809_b0 , 
		\5810_b1 , \5810_b0 , \5811_b1 , \5811_b0 , \5812_b1 , \5812_b0 , \5813_b1 , \5813_b0 , \5814_b1 , \5814_b0 , 
		\5815_b1 , \5815_b0 , \5816_b1 , \5816_b0 , \5817_b1 , \5817_b0 , \5818_b1 , \5818_b0 , \5819_b1 , \5819_b0 , 
		\5820_b1 , \5820_b0 , \5821_b1 , \5821_b0 , \5822_b1 , \5822_b0 , \5823_b1 , \5823_b0 , \5824_b1 , \5824_b0 , 
		\5825_b1 , \5825_b0 , \5826_b1 , \5826_b0 , \5827_b1 , \5827_b0 , \5828_b1 , \5828_b0 , \5829_b1 , \5829_b0 , 
		\5830_b1 , \5830_b0 , \5831_b1 , \5831_b0 , \5832_b1 , \5832_b0 , \5833_b1 , \5833_b0 , \5834_b1 , \5834_b0 , 
		\5835_b1 , \5835_b0 , \5836_b1 , \5836_b0 , \5837_b1 , \5837_b0 , \5838_b1 , \5838_b0 , \5839_b1 , \5839_b0 , 
		\5840_b1 , \5840_b0 , \5841_b1 , \5841_b0 , \5842_b1 , \5842_b0 , \5843_b1 , \5843_b0 , \5844_b1 , \5844_b0 , 
		\5845_b1 , \5845_b0 , \5846_b1 , \5846_b0 , \5847_b1 , \5847_b0 , \5848_b1 , \5848_b0 , \5849_b1 , \5849_b0 , 
		\5850_b1 , \5850_b0 , \5851_b1 , \5851_b0 , \5852_b1 , \5852_b0 , \5853_b1 , \5853_b0 , \5854_b1 , \5854_b0 , 
		\5855_b1 , \5855_b0 , \5856_b1 , \5856_b0 , \5857_b1 , \5857_b0 , \5858_b1 , \5858_b0 , \5859_b1 , \5859_b0 , 
		\5860_b1 , \5860_b0 , \5861_b1 , \5861_b0 , \5862_b1 , \5862_b0 , \5863_b1 , \5863_b0 , \5864_b1 , \5864_b0 , 
		\5865_b1 , \5865_b0 , \5866_b1 , \5866_b0 , \5867_b1 , \5867_b0 , \5868_b1 , \5868_b0 , \5869_b1 , \5869_b0 , 
		\5870_b1 , \5870_b0 , \5871_b1 , \5871_b0 , \5872_b1 , \5872_b0 , \5873_b1 , \5873_b0 , \5874_b1 , \5874_b0 , 
		\5875_b1 , \5875_b0 , \5876_b1 , \5876_b0 , \5877_b1 , \5877_b0 , \5878_b1 , \5878_b0 , \5879_b1 , \5879_b0 , 
		\5880_b1 , \5880_b0 , \5881_b1 , \5881_b0 , \5882_b1 , \5882_b0 , \5883_b1 , \5883_b0 , \5884_b1 , \5884_b0 , 
		\5885_b1 , \5885_b0 , \5886_b1 , \5886_b0 , \5887_b1 , \5887_b0 , \5888_b1 , \5888_b0 , \5889_b1 , \5889_b0 , 
		\5890_b1 , \5890_b0 , \5891_b1 , \5891_b0 , \5892_b1 , \5892_b0 , \5893_b1 , \5893_b0 , \5894_b1 , \5894_b0 , 
		\5895_b1 , \5895_b0 , \5896_b1 , \5896_b0 , \5897_b1 , \5897_b0 , \5898_b1 , \5898_b0 , \5899_b1 , \5899_b0 , 
		\5900_b1 , \5900_b0 , \5901_b1 , \5901_b0 , \5902_b1 , \5902_b0 , \5903_b1 , \5903_b0 , \5904_b1 , \5904_b0 , 
		\5905_b1 , \5905_b0 , \5906_b1 , \5906_b0 , \5907_b1 , \5907_b0 , \5908_b1 , \5908_b0 , \5909_b1 , \5909_b0 , 
		\5910_b1 , \5910_b0 , \5911_b1 , \5911_b0 , \5912_b1 , \5912_b0 , \5913_b1 , \5913_b0 , \5914_b1 , \5914_b0 , 
		\5915_b1 , \5915_b0 , \5916_b1 , \5916_b0 , \5917_b1 , \5917_b0 , \5918_b1 , \5918_b0 , \5919_b1 , \5919_b0 , 
		\5920_b1 , \5920_b0 , \5921_b1 , \5921_b0 , \5922_b1 , \5922_b0 , \5923_b1 , \5923_b0 , \5924_b1 , \5924_b0 , 
		\5925_b1 , \5925_b0 , \5926_b1 , \5926_b0 , \5927_b1 , \5927_b0 , \5928_b1 , \5928_b0 , \5929_b1 , \5929_b0 , 
		\5930_b1 , \5930_b0 , \5931_b1 , \5931_b0 , \5932_b1 , \5932_b0 , \5933_b1 , \5933_b0 , \5934_b1 , \5934_b0 , 
		\5935_b1 , \5935_b0 , \5936_b1 , \5936_b0 , \5937_b1 , \5937_b0 , \5938_b1 , \5938_b0 , \5939_b1 , \5939_b0 , 
		\5940_b1 , \5940_b0 , \5941_b1 , \5941_b0 , \5942_b1 , \5942_b0 , \5943_b1 , \5943_b0 , \5944_b1 , \5944_b0 , 
		\5945_b1 , \5945_b0 , \5946_b1 , \5946_b0 , \5947_b1 , \5947_b0 , \5948_b1 , \5948_b0 , \5949_b1 , \5949_b0 , 
		\5950_b1 , \5950_b0 , \5951_b1 , \5951_b0 , \5952_b1 , \5952_b0 , \5953_b1 , \5953_b0 , \5954_b1 , \5954_b0 , 
		\5955_b1 , \5955_b0 , \5956_b1 , \5956_b0 , \5957_b1 , \5957_b0 , \5958_b1 , \5958_b0 , \5959_b1 , \5959_b0 , 
		\5960_b1 , \5960_b0 , \5961_b1 , \5961_b0 , \5962_b1 , \5962_b0 , \5963_b1 , \5963_b0 , \5964_b1 , \5964_b0 , 
		\5965_b1 , \5965_b0 , \5966_b1 , \5966_b0 , \5967_b1 , \5967_b0 , \5968_b1 , \5968_b0 , \5969_b1 , \5969_b0 , 
		\5970_b1 , \5970_b0 , \5971_b1 , \5971_b0 , \5972_b1 , \5972_b0 , \5973_b1 , \5973_b0 , \5974_b1 , \5974_b0 , 
		\5975_b1 , \5975_b0 , \5976_b1 , \5976_b0 , \5977_b1 , \5977_b0 , \5978_b1 , \5978_b0 , \5979_b1 , \5979_b0 , 
		\5980_b1 , \5980_b0 , \5981_b1 , \5981_b0 , \5982_b1 , \5982_b0 , \5983_b1 , \5983_b0 , \5984_b1 , \5984_b0 , 
		\5985_b1 , \5985_b0 , \5986_b1 , \5986_b0 , \5987_b1 , \5987_b0 , \5988_b1 , \5988_b0 , \5989_b1 , \5989_b0 , 
		\5990_b1 , \5990_b0 , \5991_b1 , \5991_b0 , \5992_b1 , \5992_b0 , \5993_b1 , \5993_b0 , \5994_b1 , \5994_b0 , 
		\5995_b1 , \5995_b0 , \5996_b1 , \5996_b0 , \5997_b1 , \5997_b0 , \5998_b1 , \5998_b0 , \5999_b1 , \5999_b0 , 
		\6000_b1 , \6000_b0 , \6001_b1 , \6001_b0 , \6002_b1 , \6002_b0 , \6003_b1 , \6003_b0 , \6004_b1 , \6004_b0 , 
		\6005_b1 , \6005_b0 , \6006_b1 , \6006_b0 , \6007_b1 , \6007_b0 , \6008_b1 , \6008_b0 , \6009_b1 , \6009_b0 , 
		\6010_b1 , \6010_b0 , \6011_b1 , \6011_b0 , \6012_b1 , \6012_b0 , \6013_b1 , \6013_b0 , \6014_b1 , \6014_b0 , 
		\6015_b1 , \6015_b0 , \6016_b1 , \6016_b0 , \6017_b1 , \6017_b0 , \6018_b1 , \6018_b0 , \6019_b1 , \6019_b0 , 
		\6020_b1 , \6020_b0 , \6021_b1 , \6021_b0 , \6022_b1 , \6022_b0 , \6023_b1 , \6023_b0 , \6024_b1 , \6024_b0 , 
		\6025_b1 , \6025_b0 , \6026_b1 , \6026_b0 , \6027_b1 , \6027_b0 , \6028_b1 , \6028_b0 , \6029_b1 , \6029_b0 , 
		\6030_b1 , \6030_b0 , \6031_b1 , \6031_b0 , \6032_b1 , \6032_b0 , \6033_b1 , \6033_b0 , \6034_b1 , \6034_b0 , 
		\6035_b1 , \6035_b0 , \6036_b1 , \6036_b0 , \6037_b1 , \6037_b0 , \6038_b1 , \6038_b0 , \6039_b1 , \6039_b0 , 
		\6040_b1 , \6040_b0 , \6041_b1 , \6041_b0 , \6042_b1 , \6042_b0 , \6043_b1 , \6043_b0 , \6044_b1 , \6044_b0 , 
		\6045_b1 , \6045_b0 , \6046_b1 , \6046_b0 , \6047_b1 , \6047_b0 , \6048_b1 , \6048_b0 , \6049_b1 , \6049_b0 , 
		\6050_b1 , \6050_b0 , \6051_b1 , \6051_b0 , \6052_b1 , \6052_b0 , \6053_b1 , \6053_b0 , \6054_b1 , \6054_b0 , 
		\6055_b1 , \6055_b0 , \6056_b1 , \6056_b0 , \6057_b1 , \6057_b0 , \6058_b1 , \6058_b0 , \6059_b1 , \6059_b0 , 
		\6060_b1 , \6060_b0 , \6061_b1 , \6061_b0 , \6062_b1 , \6062_b0 , \6063_b1 , \6063_b0 , \6064_b1 , \6064_b0 , 
		\6065_b1 , \6065_b0 , \6066_b1 , \6066_b0 , \6067_b1 , \6067_b0 , \6068_b1 , \6068_b0 , \6069_b1 , \6069_b0 , 
		\6070_b1 , \6070_b0 , \6071_b1 , \6071_b0 , \6072_b1 , \6072_b0 , \6073_b1 , \6073_b0 , \6074_b1 , \6074_b0 , 
		\6075_b1 , \6075_b0 , \6076_b1 , \6076_b0 , \6077_b1 , \6077_b0 , \6078_b1 , \6078_b0 , \6079_b1 , \6079_b0 , 
		\6080_b1 , \6080_b0 , \6081_b1 , \6081_b0 , \6082_b1 , \6082_b0 , \6083_b1 , \6083_b0 , \6084_b1 , \6084_b0 , 
		\6085_b1 , \6085_b0 , \6086_b1 , \6086_b0 , \6087_b1 , \6087_b0 , \6088_b1 , \6088_b0 , \6089_b1 , \6089_b0 , 
		\6090_b1 , \6090_b0 , \6091_b1 , \6091_b0 , \6092_b1 , \6092_b0 , \6093_b1 , \6093_b0 , \6094_b1 , \6094_b0 , 
		\6095_b1 , \6095_b0 , \6096_b1 , \6096_b0 , \6097_b1 , \6097_b0 , \6098_b1 , \6098_b0 , \6099_b1 , \6099_b0 , 
		\6100_b1 , \6100_b0 , \6101_b1 , \6101_b0 , \6102_b1 , \6102_b0 , \6103_b1 , \6103_b0 , \6104_b1 , \6104_b0 , 
		\6105_b1 , \6105_b0 , \6106_b1 , \6106_b0 , \6107_b1 , \6107_b0 , \6108_b1 , \6108_b0 , \6109_b1 , \6109_b0 , 
		\6110_b1 , \6110_b0 , \6111_b1 , \6111_b0 , \6112_b1 , \6112_b0 , \6113_b1 , \6113_b0 , \6114_b1 , \6114_b0 , 
		\6115_b1 , \6115_b0 , \6116_b1 , \6116_b0 , \6117_b1 , \6117_b0 , \6118_b1 , \6118_b0 , \6119_b1 , \6119_b0 , 
		\6120_b1 , \6120_b0 , \6121_b1 , \6121_b0 , \6122_b1 , \6122_b0 , \6123_b1 , \6123_b0 , \6124_b1 , \6124_b0 , 
		\6125_b1 , \6125_b0 , \6126_b1 , \6126_b0 , \6127_b1 , \6127_b0 , \6128_b1 , \6128_b0 , \6129_b1 , \6129_b0 , 
		\6130_b1 , \6130_b0 , \6131_b1 , \6131_b0 , \6132_b1 , \6132_b0 , \6133_b1 , \6133_b0 , \6134_b1 , \6134_b0 , 
		\6135_b1 , \6135_b0 , \6136_b1 , \6136_b0 , \6137_b1 , \6137_b0 , \6138_b1 , \6138_b0 , \6139_b1 , \6139_b0 , 
		\6140_b1 , \6140_b0 , \6141_b1 , \6141_b0 , \6142_b1 , \6142_b0 , \6143_b1 , \6143_b0 , \6144_b1 , \6144_b0 , 
		\6145_b1 , \6145_b0 , \6146_b1 , \6146_b0 , \6147_b1 , \6147_b0 , \6148_b1 , \6148_b0 , \6149_b1 , \6149_b0 , 
		\6150_b1 , \6150_b0 , \6151_b1 , \6151_b0 , \6152_b1 , \6152_b0 , \6153_b1 , \6153_b0 , \6154_b1 , \6154_b0 , 
		\6155_b1 , \6155_b0 , \6156_b1 , \6156_b0 , \6157_b1 , \6157_b0 , \6158_b1 , \6158_b0 , \6159_b1 , \6159_b0 , 
		\6160_b1 , \6160_b0 , \6161_b1 , \6161_b0 , \6162_b1 , \6162_b0 , \6163_b1 , \6163_b0 , \6164_b1 , \6164_b0 , 
		\6165_b1 , \6165_b0 , \6166_b1 , \6166_b0 , \6167_b1 , \6167_b0 , \6168_b1 , \6168_b0 , \6169_b1 , \6169_b0 , 
		\6170_b1 , \6170_b0 , \6171_b1 , \6171_b0 , \6172_b1 , \6172_b0 , \6173_b1 , \6173_b0 , \6174_b1 , \6174_b0 , 
		\6175_b1 , \6175_b0 , \6176_b1 , \6176_b0 , \6177_b1 , \6177_b0 , \6178_b1 , \6178_b0 , \6179_b1 , \6179_b0 , 
		\6180_b1 , \6180_b0 , \6181_b1 , \6181_b0 , \6182_b1 , \6182_b0 , \6183_b1 , \6183_b0 , \6184_b1 , \6184_b0 , 
		\6185_b1 , \6185_b0 , \6186_b1 , \6186_b0 , \6187_b1 , \6187_b0 , \6188_b1 , \6188_b0 , \6189_b1 , \6189_b0 , 
		\6190_b1 , \6190_b0 , \6191_b1 , \6191_b0 , \6192_b1 , \6192_b0 , \6193_b1 , \6193_b0 , \6194_b1 , \6194_b0 , 
		\6195_b1 , \6195_b0 , \6196_b1 , \6196_b0 , \6197_b1 , \6197_b0 , \6198_b1 , \6198_b0 , \6199_b1 , \6199_b0 , 
		\6200_b1 , \6200_b0 , \6201_b1 , \6201_b0 , \6202_b1 , \6202_b0 , \6203_b1 , \6203_b0 , \6204_b1 , \6204_b0 , 
		\6205_b1 , \6205_b0 , \6206_b1 , \6206_b0 , \6207_b1 , \6207_b0 , \6208_b1 , \6208_b0 , \6209_b1 , \6209_b0 , 
		\6210_b1 , \6210_b0 , \6211_b1 , \6211_b0 , \6212_b1 , \6212_b0 , \6213_b1 , \6213_b0 , \6214_b1 , \6214_b0 , 
		\6215_b1 , \6215_b0 , \6216_b1 , \6216_b0 , \6217_b1 , \6217_b0 , \6218_b1 , \6218_b0 , \6219_b1 , \6219_b0 , 
		\6220_b1 , \6220_b0 , \6221_b1 , \6221_b0 , \6222_b1 , \6222_b0 , \6223_b1 , \6223_b0 , \6224_b1 , \6224_b0 , 
		\6225_b1 , \6225_b0 , \6226_b1 , \6226_b0 , \6227_b1 , \6227_b0 , \6228_b1 , \6228_b0 , \6229_b1 , \6229_b0 , 
		\6230_b1 , \6230_b0 , \6231_b1 , \6231_b0 , \6232_b1 , \6232_b0 , \6233_b1 , \6233_b0 , \6234_b1 , \6234_b0 , 
		\6235_b1 , \6235_b0 , \6236_b1 , \6236_b0 , \6237_b1 , \6237_b0 , \6238_b1 , \6238_b0 , \6239_b1 , \6239_b0 , 
		\6240_b1 , \6240_b0 , \6241_b1 , \6241_b0 , \6242_b1 , \6242_b0 , \6243_b1 , \6243_b0 , \6244_b1 , \6244_b0 , 
		\6245_b1 , \6245_b0 , \6246_b1 , \6246_b0 , \6247_b1 , \6247_b0 , \6248_b1 , \6248_b0 , \6249_b1 , \6249_b0 , 
		\6250_b1 , \6250_b0 , \6251_b1 , \6251_b0 , \6252_b1 , \6252_b0 , \6253_b1 , \6253_b0 , \6254_b1 , \6254_b0 , 
		\6255_b1 , \6255_b0 , \6256_b1 , \6256_b0 , \6257_b1 , \6257_b0 , \6258_b1 , \6258_b0 , \6259_b1 , \6259_b0 , 
		\6260_b1 , \6260_b0 , \6261_b1 , \6261_b0 , \6262_b1 , \6262_b0 , \6263_b1 , \6263_b0 , \6264_b1 , \6264_b0 , 
		\6265_b1 , \6265_b0 , \6266_b1 , \6266_b0 , \6267_b1 , \6267_b0 , \6268_b1 , \6268_b0 , \6269_b1 , \6269_b0 , 
		\6270_b1 , \6270_b0 , \6271_b1 , \6271_b0 , \6272_b1 , \6272_b0 , \6273_b1 , \6273_b0 , \6274_b1 , \6274_b0 , 
		\6275_b1 , \6275_b0 , \6276_b1 , \6276_b0 , \6277_b1 , \6277_b0 , \6278_b1 , \6278_b0 , \6279_b1 , \6279_b0 , 
		\6280_b1 , \6280_b0 , \6281_b1 , \6281_b0 , \6282_b1 , \6282_b0 , \6283_b1 , \6283_b0 , \6284_b1 , \6284_b0 , 
		\6285_b1 , \6285_b0 , \6286_b1 , \6286_b0 , \6287_b1 , \6287_b0 , \6288_b1 , \6288_b0 , \6289_b1 , \6289_b0 , 
		\6290_b1 , \6290_b0 , \6291_b1 , \6291_b0 , \6292_b1 , \6292_b0 , \6293_b1 , \6293_b0 , \6294_b1 , \6294_b0 , 
		\6295_b1 , \6295_b0 , \6296_b1 , \6296_b0 , \6297_b1 , \6297_b0 , \6298_b1 , \6298_b0 , \6299_b1 , \6299_b0 , 
		\6300_b1 , \6300_b0 , \6301_b1 , \6301_b0 , \6302_b1 , \6302_b0 , \6303_b1 , \6303_b0 , \6304_b1 , \6304_b0 , 
		\6305_b1 , \6305_b0 , \6306_b1 , \6306_b0 , \6307_b1 , \6307_b0 , \6308_b1 , \6308_b0 , \6309_b1 , \6309_b0 , 
		\6310_b1 , \6310_b0 , \6311_b1 , \6311_b0 , \6312_b1 , \6312_b0 , \6313_b1 , \6313_b0 , \6314_b1 , \6314_b0 , 
		\6315_b1 , \6315_b0 , \6316_b1 , \6316_b0 , \6317_b1 , \6317_b0 , \6318_b1 , \6318_b0 , \6319_b1 , \6319_b0 , 
		\6320_b1 , \6320_b0 , \6321_b1 , \6321_b0 , \6322_b1 , \6322_b0 , \6323_b1 , \6323_b0 , \6324_b1 , \6324_b0 , 
		\6325_b1 , \6325_b0 , \6326_b1 , \6326_b0 , \6327_b1 , \6327_b0 , \6328_b1 , \6328_b0 , \6329_b1 , \6329_b0 , 
		\6330_b1 , \6330_b0 , \6331_b1 , \6331_b0 , \6332_b1 , \6332_b0 , \6333_b1 , \6333_b0 , \6334_b1 , \6334_b0 , 
		\6335_b1 , \6335_b0 , \6336_b1 , \6336_b0 , \6337_b1 , \6337_b0 , \6338_b1 , \6338_b0 , \6339_b1 , \6339_b0 , 
		\6340_b1 , \6340_b0 , \6341_b1 , \6341_b0 , \6342_b1 , \6342_b0 , \6343_b1 , \6343_b0 , \6344_b1 , \6344_b0 , 
		\6345_b1 , \6345_b0 , \6346_b1 , \6346_b0 , \6347_b1 , \6347_b0 , \6348_b1 , \6348_b0 , \6349_b1 , \6349_b0 , 
		\6350_b1 , \6350_b0 , \6351_b1 , \6351_b0 , \6352_b1 , \6352_b0 , \6353_b1 , \6353_b0 , \6354_b1 , \6354_b0 , 
		\6355_b1 , \6355_b0 , \6356_b1 , \6356_b0 , \6357_b1 , \6357_b0 , \6358_b1 , \6358_b0 , \6359_b1 , \6359_b0 , 
		\6360_b1 , \6360_b0 , \6361_b1 , \6361_b0 , \6362_b1 , \6362_b0 , \6363_b1 , \6363_b0 , \6364_b1 , \6364_b0 , 
		\6365_b1 , \6365_b0 , \6366_b1 , \6366_b0 , \6367_b1 , \6367_b0 , \6368_b1 , \6368_b0 , \6369_b1 , \6369_b0 , 
		\6370_b1 , \6370_b0 , \6371_b1 , \6371_b0 , \6372_b1 , \6372_b0 , \6373_b1 , \6373_b0 , \6374_b1 , \6374_b0 , 
		\6375_b1 , \6375_b0 , \6376_b1 , \6376_b0 , \6377_b1 , \6377_b0 , \6378_b1 , \6378_b0 , \6379_b1 , \6379_b0 , 
		\6380_b1 , \6380_b0 , \6381_b1 , \6381_b0 , \6382_b1 , \6382_b0 , \6383_b1 , \6383_b0 , \6384_b1 , \6384_b0 , 
		\6385_b1 , \6385_b0 , \6386_b1 , \6386_b0 , \6387_b1 , \6387_b0 , \6388_b1 , \6388_b0 , \6389_b1 , \6389_b0 , 
		\6390_b1 , \6390_b0 , \6391_b1 , \6391_b0 , \6392_b1 , \6392_b0 , \6393_b1 , \6393_b0 , \6394_b1 , \6394_b0 , 
		\6395_b1 , \6395_b0 , \6396_b1 , \6396_b0 , \6397_b1 , \6397_b0 , \6398_b1 , \6398_b0 , \6399_b1 , \6399_b0 , 
		\6400_b1 , \6400_b0 , \6401_b1 , \6401_b0 , \6402_b1 , \6402_b0 , \6403_b1 , \6403_b0 , \6404_b1 , \6404_b0 , 
		\6405_b1 , \6405_b0 , \6406_b1 , \6406_b0 , \6407_b1 , \6407_b0 , \6408_b1 , \6408_b0 , \6409_b1 , \6409_b0 , 
		\6410_b1 , \6410_b0 , \6411_b1 , \6411_b0 , \6412_b1 , \6412_b0 , \6413_b1 , \6413_b0 , \6414_b1 , \6414_b0 , 
		\6415_b1 , \6415_b0 , \6416_b1 , \6416_b0 , \6417_b1 , \6417_b0 , \6418_b1 , \6418_b0 , \6419_b1 , \6419_b0 , 
		\6420_b1 , \6420_b0 , \6421_b1 , \6421_b0 , \6422_b1 , \6422_b0 , \6423_b1 , \6423_b0 , \6424_b1 , \6424_b0 , 
		\6425_b1 , \6425_b0 , \6426_b1 , \6426_b0 , \6427_b1 , \6427_b0 , \6428_b1 , \6428_b0 , \6429_b1 , \6429_b0 , 
		\6430_b1 , \6430_b0 , \6431_b1 , \6431_b0 , \6432_b1 , \6432_b0 , \6433_b1 , \6433_b0 , \6434_b1 , \6434_b0 , 
		\6435_b1 , \6435_b0 , \6436_b1 , \6436_b0 , \6437_b1 , \6437_b0 , \6438_b1 , \6438_b0 , \6439_b1 , \6439_b0 , 
		\6440_b1 , \6440_b0 , \6441_b1 , \6441_b0 , \6442_b1 , \6442_b0 , \6443_b1 , \6443_b0 , \6444_b1 , \6444_b0 , 
		\6445_b1 , \6445_b0 , \6446_b1 , \6446_b0 , \6447_b1 , \6447_b0 , \6448_b1 , \6448_b0 , \6449_b1 , \6449_b0 , 
		\6450_b1 , \6450_b0 , \6451_b1 , \6451_b0 , \6452_b1 , \6452_b0 , \6453_b1 , \6453_b0 , \6454_b1 , \6454_b0 , 
		\6455_b1 , \6455_b0 , \6456_b1 , \6456_b0 , \6457_b1 , \6457_b0 , \6458_b1 , \6458_b0 , \6459_b1 , \6459_b0 , 
		\6460_b1 , \6460_b0 , \6461_b1 , \6461_b0 , \6462_b1 , \6462_b0 , \6463_b1 , \6463_b0 , \6464_b1 , \6464_b0 , 
		\6465_b1 , \6465_b0 , \6466_b1 , \6466_b0 , \6467_b1 , \6467_b0 , \6468_b1 , \6468_b0 , \6469_b1 , \6469_b0 , 
		\6470_b1 , \6470_b0 , \6471_b1 , \6471_b0 , \6472_b1 , \6472_b0 , \6473_b1 , \6473_b0 , \6474_b1 , \6474_b0 , 
		\6475_b1 , \6475_b0 , \6476_b1 , \6476_b0 , \6477_b1 , \6477_b0 , \6478_b1 , \6478_b0 , \6479_b1 , \6479_b0 , 
		\6480_b1 , \6480_b0 , \6481_b1 , \6481_b0 , \6482_b1 , \6482_b0 , \6483_b1 , \6483_b0 , \6484_b1 , \6484_b0 , 
		\6485_b1 , \6485_b0 , \6486_b1 , \6486_b0 , \6487_b1 , \6487_b0 , \6488_b1 , \6488_b0 , \6489_b1 , \6489_b0 , 
		\6490_b1 , \6490_b0 , \6491_b1 , \6491_b0 , \6492_b1 , \6492_b0 , \6493_b1 , \6493_b0 , \6494_b1 , \6494_b0 , 
		\6495_b1 , \6495_b0 , \6496_b1 , \6496_b0 , \6497_b1 , \6497_b0 , \6498_b1 , \6498_b0 , \6499_b1 , \6499_b0 , 
		\6500_b1 , \6500_b0 , \6501_b1 , \6501_b0 , \6502_b1 , \6502_b0 , \6503_b1 , \6503_b0 , \6504_b1 , \6504_b0 , 
		\6505_b1 , \6505_b0 , \6506_b1 , \6506_b0 , \6507_b1 , \6507_b0 , \6508_b1 , \6508_b0 , \6509_b1 , \6509_b0 , 
		\6510_b1 , \6510_b0 , \6511_b1 , \6511_b0 , \6512_b1 , \6512_b0 , \6513_b1 , \6513_b0 , \6514_b1 , \6514_b0 , 
		\6515_b1 , \6515_b0 , \6516_b1 , \6516_b0 , \6517_b1 , \6517_b0 , \6518_b1 , \6518_b0 , \6519_b1 , \6519_b0 , 
		\6520_b1 , \6520_b0 , \6521_b1 , \6521_b0 , \6522_b1 , \6522_b0 , \6523_b1 , \6523_b0 , \6524_b1 , \6524_b0 , 
		\6525_b1 , \6525_b0 , \6526_b1 , \6526_b0 , \6527_b1 , \6527_b0 , \6528_b1 , \6528_b0 , \6529_b1 , \6529_b0 , 
		\6530_b1 , \6530_b0 , \6531_b1 , \6531_b0 , \6532_b1 , \6532_b0 , \6533_b1 , \6533_b0 , \6534_b1 , \6534_b0 , 
		\6535_b1 , \6535_b0 , \6536_b1 , \6536_b0 , \6537_b1 , \6537_b0 , \6538_b1 , \6538_b0 , \6539_b1 , \6539_b0 , 
		\6540_b1 , \6540_b0 , \6541_b1 , \6541_b0 , \6542_b1 , \6542_b0 , \6543_b1 , \6543_b0 , \6544_b1 , \6544_b0 , 
		\6545_b1 , \6545_b0 , \6546_b1 , \6546_b0 , \6547_b1 , \6547_b0 , \6548_b1 , \6548_b0 , \6549_b1 , \6549_b0 , 
		\6550_b1 , \6550_b0 , \6551_b1 , \6551_b0 , \6552_b1 , \6552_b0 , \6553_b1 , \6553_b0 , \6554_b1 , \6554_b0 , 
		\6555_b1 , \6555_b0 , \6556_b1 , \6556_b0 , \6557_b1 , \6557_b0 , \6558_b1 , \6558_b0 , \6559_b1 , \6559_b0 , 
		\6560_b1 , \6560_b0 , \6561_b1 , \6561_b0 , \6562_b1 , \6562_b0 , \6563_b1 , \6563_b0 , \6564_b1 , \6564_b0 , 
		\6565_b1 , \6565_b0 , \6566_b1 , \6566_b0 , \6567_b1 , \6567_b0 , \6568_b1 , \6568_b0 , \6569_b1 , \6569_b0 , 
		\6570_b1 , \6570_b0 , \6571_b1 , \6571_b0 , \6572_b1 , \6572_b0 , \6573_b1 , \6573_b0 , \6574_b1 , \6574_b0 , 
		\6575_b1 , \6575_b0 , \6576_b1 , \6576_b0 , \6577_b1 , \6577_b0 , \6578_b1 , \6578_b0 , \6579_b1 , \6579_b0 , 
		\6580_b1 , \6580_b0 , \6581_b1 , \6581_b0 , \6582_b1 , \6582_b0 , \6583_b1 , \6583_b0 , \6584_b1 , \6584_b0 , 
		\6585_b1 , \6585_b0 , \6586_b1 , \6586_b0 , \6587_b1 , \6587_b0 , \6588_b1 , \6588_b0 , \6589_b1 , \6589_b0 , 
		\6590_b1 , \6590_b0 , \6591_b1 , \6591_b0 , \6592_b1 , \6592_b0 , \6593_b1 , \6593_b0 , \6594_b1 , \6594_b0 , 
		\6595_b1 , \6595_b0 , \6596_b1 , \6596_b0 , \6597_b1 , \6597_b0 , \6598_b1 , \6598_b0 , \6599_b1 , \6599_b0 , 
		\6600_b1 , \6600_b0 , \6601_b1 , \6601_b0 , \6602_b1 , \6602_b0 , \6603_b1 , \6603_b0 , \6604_b1 , \6604_b0 , 
		\6605_b1 , \6605_b0 , \6606_b1 , \6606_b0 , \6607_b1 , \6607_b0 , \6608_b1 , \6608_b0 , \6609_b1 , \6609_b0 , 
		\6610_b1 , \6610_b0 , \6611_b1 , \6611_b0 , \6612_b1 , \6612_b0 , \6613_b1 , \6613_b0 , \6614_b1 , \6614_b0 , 
		\6615_b1 , \6615_b0 , \6616_b1 , \6616_b0 , \6617_b1 , \6617_b0 , \6618_b1 , \6618_b0 , \6619_b1 , \6619_b0 , 
		\6620_b1 , \6620_b0 , \6621_b1 , \6621_b0 , \6622_b1 , \6622_b0 , \6623_b1 , \6623_b0 , \6624_b1 , \6624_b0 , 
		\6625_b1 , \6625_b0 , \6626_b1 , \6626_b0 , \6627_b1 , \6627_b0 , \6628_b1 , \6628_b0 , \6629_b1 , \6629_b0 , 
		\6630_b1 , \6630_b0 , \6631_b1 , \6631_b0 , \6632_b1 , \6632_b0 , \6633_b1 , \6633_b0 , \6634_b1 , \6634_b0 , 
		\6635_b1 , \6635_b0 , \6636_b1 , \6636_b0 , \6637_b1 , \6637_b0 , \6638_b1 , \6638_b0 , \6639_b1 , \6639_b0 , 
		\6640_b1 , \6640_b0 , \6641_b1 , \6641_b0 , \6642_b1 , \6642_b0 , \6643_b1 , \6643_b0 , \6644_b1 , \6644_b0 , 
		\6645_b1 , \6645_b0 , \6646_b1 , \6646_b0 , \6647_b1 , \6647_b0 , \6648_b1 , \6648_b0 , \6649_b1 , \6649_b0 , 
		\6650_b1 , \6650_b0 , \6651_b1 , \6651_b0 , \6652_b1 , \6652_b0 , \6653_b1 , \6653_b0 , \6654_b1 , \6654_b0 , 
		\6655_b1 , \6655_b0 , \6656_b1 , \6656_b0 , \6657_b1 , \6657_b0 , \6658_b1 , \6658_b0 , \6659_b1 , \6659_b0 , 
		\6660_b1 , \6660_b0 , \6661_b1 , \6661_b0 , \6662_b1 , \6662_b0 , \6663_b1 , \6663_b0 , \6664_b1 , \6664_b0 , 
		\6665_b1 , \6665_b0 , \6666_b1 , \6666_b0 , \6667_b1 , \6667_b0 , \6668_b1 , \6668_b0 , \6669_b1 , \6669_b0 , 
		\6670_b1 , \6670_b0 , \6671_b1 , \6671_b0 , \6672_b1 , \6672_b0 , \6673_b1 , \6673_b0 , \6674_b1 , \6674_b0 , 
		\6675_b1 , \6675_b0 , \6676_b1 , \6676_b0 , \6677_b1 , \6677_b0 , \6678_b1 , \6678_b0 , \6679_b1 , \6679_b0 , 
		\6680_b1 , \6680_b0 , \6681_b1 , \6681_b0 , \6682_b1 , \6682_b0 , \6683_b1 , \6683_b0 , \6684_b1 , \6684_b0 , 
		\6685_b1 , \6685_b0 , \6686_b1 , \6686_b0 , \6687_b1 , \6687_b0 , \6688_b1 , \6688_b0 , \6689_b1 , \6689_b0 , 
		\6690_b1 , \6690_b0 , \6691_b1 , \6691_b0 , \6692_b1 , \6692_b0 , \6693_b1 , \6693_b0 , \6694_b1 , \6694_b0 , 
		\6695_b1 , \6695_b0 , \6696_b1 , \6696_b0 , \6697_b1 , \6697_b0 , \6698_b1 , \6698_b0 , \6699_b1 , \6699_b0 , 
		\6700_b1 , \6700_b0 , \6701_b1 , \6701_b0 , \6702_b1 , \6702_b0 , \6703_b1 , \6703_b0 , \6704_b1 , \6704_b0 , 
		\6705_b1 , \6705_b0 , \6706_b1 , \6706_b0 , \6707_b1 , \6707_b0 , \6708_b1 , \6708_b0 , \6709_b1 , \6709_b0 , 
		\6710_b1 , \6710_b0 , \6711_b1 , \6711_b0 , \6712_b1 , \6712_b0 , \6713_b1 , \6713_b0 , \6714_b1 , \6714_b0 , 
		\6715_b1 , \6715_b0 , \6716_b1 , \6716_b0 , \6717_b1 , \6717_b0 , \6718_b1 , \6718_b0 , \6719_b1 , \6719_b0 , 
		\6720_b1 , \6720_b0 , \6721_b1 , \6721_b0 , \6722_b1 , \6722_b0 , \6723_b1 , \6723_b0 , \6724_b1 , \6724_b0 , 
		\6725_b1 , \6725_b0 , \6726_b1 , \6726_b0 , \6727_b1 , \6727_b0 , \6728_b1 , \6728_b0 , \6729_b1 , \6729_b0 , 
		\6730_b1 , \6730_b0 , \6731_b1 , \6731_b0 , \6732_b1 , \6732_b0 , \6733_b1 , \6733_b0 , \6734_b1 , \6734_b0 , 
		\6735_b1 , \6735_b0 , \6736_b1 , \6736_b0 , \6737_b1 , \6737_b0 , \6738_b1 , \6738_b0 , \6739_b1 , \6739_b0 , 
		\6740_b1 , \6740_b0 , \6741_b1 , \6741_b0 , \6742_b1 , \6742_b0 , \6743_b1 , \6743_b0 , \6744_b1 , \6744_b0 , 
		\6745_b1 , \6745_b0 , \6746_b1 , \6746_b0 , \6747_b1 , \6747_b0 , \6748_b1 , \6748_b0 , \6749_b1 , \6749_b0 , 
		\6750_b1 , \6750_b0 , \6751_b1 , \6751_b0 , \6752_b1 , \6752_b0 , \6753_b1 , \6753_b0 , \6754_b1 , \6754_b0 , 
		\6755_b1 , \6755_b0 , \6756_b1 , \6756_b0 , \6757_b1 , \6757_b0 , \6758_b1 , \6758_b0 , \6759_b1 , \6759_b0 , 
		\6760_b1 , \6760_b0 , \6761_b1 , \6761_b0 , \6762_b1 , \6762_b0 , \6763_b1 , \6763_b0 , \6764_b1 , \6764_b0 , 
		\6765_b1 , \6765_b0 , \6766_b1 , \6766_b0 , \6767_b1 , \6767_b0 , \6768_b1 , \6768_b0 , \6769_b1 , \6769_b0 , 
		\6770_b1 , \6770_b0 , \6771_b1 , \6771_b0 , \6772_b1 , \6772_b0 , \6773_b1 , \6773_b0 , \6774_b1 , \6774_b0 , 
		\6775_b1 , \6775_b0 , \6776_b1 , \6776_b0 , \6777_b1 , \6777_b0 , \6778_b1 , \6778_b0 , \6779_b1 , \6779_b0 , 
		\6780_b1 , \6780_b0 , \6781_b1 , \6781_b0 , \6782_b1 , \6782_b0 , \6783_b1 , \6783_b0 , \6784_b1 , \6784_b0 , 
		\6785_b1 , \6785_b0 , \6786_b1 , \6786_b0 , \6787_b1 , \6787_b0 , \6788_b1 , \6788_b0 , \6789_b1 , \6789_b0 , 
		\6790_b1 , \6790_b0 , \6791_b1 , \6791_b0 , \6792_b1 , \6792_b0 , \6793_b1 , \6793_b0 , \6794_b1 , \6794_b0 , 
		\6795_b1 , \6795_b0 , \6796_b1 , \6796_b0 , \6797_b1 , \6797_b0 , \6798_b1 , \6798_b0 , \6799_b1 , \6799_b0 , 
		\6800_b1 , \6800_b0 , \6801_b1 , \6801_b0 , \6802_b1 , \6802_b0 , \6803_b1 , \6803_b0 , \6804_b1 , \6804_b0 , 
		\6805_b1 , \6805_b0 , \6806_b1 , \6806_b0 , \6807_b1 , \6807_b0 , \6808_b1 , \6808_b0 , \6809_b1 , \6809_b0 , 
		\6810_b1 , \6810_b0 , \6811_b1 , \6811_b0 , \6812_b1 , \6812_b0 , \6813_b1 , \6813_b0 , \6814_b1 , \6814_b0 , 
		\6815_b1 , \6815_b0 , \6816_b1 , \6816_b0 , \6817_b1 , \6817_b0 , \6818_b1 , \6818_b0 , \6819_b1 , \6819_b0 , 
		\6820_b1 , \6820_b0 , \6821_b1 , \6821_b0 , \6822_b1 , \6822_b0 , \6823_b1 , \6823_b0 , \6824_b1 , \6824_b0 , 
		\6825_b1 , \6825_b0 , \6826_b1 , \6826_b0 , \6827_b1 , \6827_b0 , \6828_b1 , \6828_b0 , \6829_b1 , \6829_b0 , 
		\6830_b1 , \6830_b0 , \6831_b1 , \6831_b0 , \6832_b1 , \6832_b0 , \6833_b1 , \6833_b0 , \6834_b1 , \6834_b0 , 
		\6835_b1 , \6835_b0 , \6836_b1 , \6836_b0 , \6837_b1 , \6837_b0 , \6838_b1 , \6838_b0 , \6839_b1 , \6839_b0 , 
		\6840_b1 , \6840_b0 , \6841_b1 , \6841_b0 , \6842_b1 , \6842_b0 , \6843_b1 , \6843_b0 , \6844_b1 , \6844_b0 , 
		\6845_b1 , \6845_b0 , \6846_b1 , \6846_b0 , \6847_b1 , \6847_b0 , \6848_b1 , \6848_b0 , \6849_b1 , \6849_b0 , 
		\6850_b1 , \6850_b0 , \6851_b1 , \6851_b0 , \6852_b1 , \6852_b0 , \6853_b1 , \6853_b0 , \6854_b1 , \6854_b0 , 
		\6855_b1 , \6855_b0 , \6856_b1 , \6856_b0 , \6857_b1 , \6857_b0 , \6858_b1 , \6858_b0 , \6859_b1 , \6859_b0 , 
		\6860_b1 , \6860_b0 , \6861_b1 , \6861_b0 , \6862_b1 , \6862_b0 , \6863_b1 , \6863_b0 , \6864_b1 , \6864_b0 , 
		\6865_b1 , \6865_b0 , \6866_b1 , \6866_b0 , \6867_b1 , \6867_b0 , \6868_b1 , \6868_b0 , \6869_b1 , \6869_b0 , 
		\6870_b1 , \6870_b0 , \6871_b1 , \6871_b0 , \6872_b1 , \6872_b0 , \6873_b1 , \6873_b0 , \6874_b1 , \6874_b0 , 
		\6875_b1 , \6875_b0 , \6876_b1 , \6876_b0 , \6877_b1 , \6877_b0 , \6878_b1 , \6878_b0 , \6879_b1 , \6879_b0 , 
		\6880_b1 , \6880_b0 , \6881_b1 , \6881_b0 , \6882_b1 , \6882_b0 , \6883_b1 , \6883_b0 , \6884_b1 , \6884_b0 , 
		\6885_b1 , \6885_b0 , \6886_b1 , \6886_b0 , \6887_b1 , \6887_b0 , \6888_b1 , \6888_b0 , \6889_b1 , \6889_b0 , 
		\6890_b1 , \6890_b0 , \6891_b1 , \6891_b0 , \6892_b1 , \6892_b0 , \6893_b1 , \6893_b0 , \6894_b1 , \6894_b0 , 
		\6895_b1 , \6895_b0 , \6896_b1 , \6896_b0 , \6897_b1 , \6897_b0 , \6898_b1 , \6898_b0 , \6899_b1 , \6899_b0 , 
		\6900_b1 , \6900_b0 , \6901_b1 , \6901_b0 , \6902_b1 , \6902_b0 , \6903_b1 , \6903_b0 , \6904_b1 , \6904_b0 , 
		\6905_b1 , \6905_b0 , \6906_b1 , \6906_b0 , \6907_b1 , \6907_b0 , \6908_b1 , \6908_b0 , \6909_b1 , \6909_b0 , 
		\6910_b1 , \6910_b0 , \6911_b1 , \6911_b0 , \6912_b1 , \6912_b0 , \6913_b1 , \6913_b0 , \6914_b1 , \6914_b0 , 
		\6915_b1 , \6915_b0 , \6916_b1 , \6916_b0 , \6917_b1 , \6917_b0 , \6918_b1 , \6918_b0 , \6919_b1 , \6919_b0 , 
		\6920_b1 , \6920_b0 , \6921_b1 , \6921_b0 , \6922_b1 , \6922_b0 , \6923_b1 , \6923_b0 , \6924_b1 , \6924_b0 , 
		\6925_b1 , \6925_b0 , \6926_b1 , \6926_b0 , \6927_b1 , \6927_b0 , \6928_b1 , \6928_b0 , \6929_b1 , \6929_b0 , 
		\6930_b1 , \6930_b0 , \6931_b1 , \6931_b0 , \6932_b1 , \6932_b0 , \6933_b1 , \6933_b0 , \6934_b1 , \6934_b0 , 
		\6935_b1 , \6935_b0 , \6936_b1 , \6936_b0 , \6937_b1 , \6937_b0 , \6938_b1 , \6938_b0 , \6939_b1 , \6939_b0 , 
		\6940_b1 , \6940_b0 , \6941_b1 , \6941_b0 , \6942_b1 , \6942_b0 , \6943_b1 , \6943_b0 , \6944_b1 , \6944_b0 , 
		\6945_b1 , \6945_b0 , \6946_b1 , \6946_b0 , \6947_b1 , \6947_b0 , \6948_b1 , \6948_b0 , \6949_b1 , \6949_b0 , 
		\6950_b1 , \6950_b0 , \6951_b1 , \6951_b0 , \6952_b1 , \6952_b0 , \6953_b1 , \6953_b0 , \6954_b1 , \6954_b0 , 
		\6955_b1 , \6955_b0 , \6956_b1 , \6956_b0 , \6957_b1 , \6957_b0 , \6958_b1 , \6958_b0 , \6959_b1 , \6959_b0 , 
		\6960_b1 , \6960_b0 , \6961_b1 , \6961_b0 , \6962_b1 , \6962_b0 , \6963_b1 , \6963_b0 , \6964_b1 , \6964_b0 , 
		\6965_b1 , \6965_b0 , \6966_b1 , \6966_b0 , \6967_b1 , \6967_b0 , \6968_b1 , \6968_b0 , \6969_b1 , \6969_b0 , 
		\6970_b1 , \6970_b0 , \6971_b1 , \6971_b0 , \6972_b1 , \6972_b0 , \6973_b1 , \6973_b0 , \6974_b1 , \6974_b0 , 
		\6975_b1 , \6975_b0 , \6976_b1 , \6976_b0 , \6977_b1 , \6977_b0 , \6978_b1 , \6978_b0 , \6979_b1 , \6979_b0 , 
		\6980_b1 , \6980_b0 , \6981_b1 , \6981_b0 , \6982_b1 , \6982_b0 , \6983_b1 , \6983_b0 , \6984_b1 , \6984_b0 , 
		\6985_b1 , \6985_b0 , \6986_b1 , \6986_b0 , \6987_b1 , \6987_b0 , \6988_b1 , \6988_b0 , \6989_b1 , \6989_b0 , 
		\6990_b1 , \6990_b0 , \6991_b1 , \6991_b0 , \6992_b1 , \6992_b0 , \6993_b1 , \6993_b0 , \6994_b1 , \6994_b0 , 
		\6995_b1 , \6995_b0 , \6996_b1 , \6996_b0 , \6997_b1 , \6997_b0 , \6998_b1 , \6998_b0 , \6999_b1 , \6999_b0 , 
		\7000_b1 , \7000_b0 , \7001_b1 , \7001_b0 , \7002_b1 , \7002_b0 , \7003_b1 , \7003_b0 , \7004_b1 , \7004_b0 , 
		\7005_b1 , \7005_b0 , \7006_b1 , \7006_b0 , \7007_b1 , \7007_b0 , \7008_b1 , \7008_b0 , \7009_b1 , \7009_b0 , 
		\7010_b1 , \7010_b0 , \7011_b1 , \7011_b0 , \7012_b1 , \7012_b0 , \7013_b1 , \7013_b0 , \7014_b1 , \7014_b0 , 
		\7015_b1 , \7015_b0 , \7016_b1 , \7016_b0 , \7017_b1 , \7017_b0 , \7018_b1 , \7018_b0 , \7019_b1 , \7019_b0 , 
		\7020_b1 , \7020_b0 , \7021_b1 , \7021_b0 , \7022_b1 , \7022_b0 , \7023_b1 , \7023_b0 , \7024_b1 , \7024_b0 , 
		\7025_b1 , \7025_b0 , \7026_b1 , \7026_b0 , \7027_b1 , \7027_b0 , \7028_b1 , \7028_b0 , \7029_b1 , \7029_b0 , 
		\7030_b1 , \7030_b0 , \7031_b1 , \7031_b0 , \7032_b1 , \7032_b0 , \7033_b1 , \7033_b0 , \7034_b1 , \7034_b0 , 
		\7035_b1 , \7035_b0 , \7036_b1 , \7036_b0 , \7037_b1 , \7037_b0 , \7038_b1 , \7038_b0 , \7039_b1 , \7039_b0 , 
		\7040_b1 , \7040_b0 , \7041_b1 , \7041_b0 , \7042_b1 , \7042_b0 , \7043_b1 , \7043_b0 , \7044_b1 , \7044_b0 , 
		\7045_b1 , \7045_b0 , \7046_b1 , \7046_b0 , \7047_b1 , \7047_b0 , \7048_b1 , \7048_b0 , \7049_b1 , \7049_b0 , 
		\7050_b1 , \7050_b0 , \7051_b1 , \7051_b0 , \7052_b1 , \7052_b0 , \7053_b1 , \7053_b0 , \7054_b1 , \7054_b0 , 
		\7055_b1 , \7055_b0 , \7056_b1 , \7056_b0 , \7057_b1 , \7057_b0 , \7058_b1 , \7058_b0 , \7059_b1 , \7059_b0 , 
		\7060_b1 , \7060_b0 , \7061_b1 , \7061_b0 , \7062_b1 , \7062_b0 , \7063_b1 , \7063_b0 , \7064_b1 , \7064_b0 , 
		\7065_b1 , \7065_b0 , \7066_b1 , \7066_b0 , \7067_b1 , \7067_b0 , \7068_b1 , \7068_b0 , \7069_b1 , \7069_b0 , 
		\7070_b1 , \7070_b0 , \7071_b1 , \7071_b0 , \7072_b1 , \7072_b0 , \7073_b1 , \7073_b0 , \7074_b1 , \7074_b0 , 
		\7075_b1 , \7075_b0 , \7076_b1 , \7076_b0 , \7077_b1 , \7077_b0 , \7078_b1 , \7078_b0 , \7079_b1 , \7079_b0 , 
		\7080_b1 , \7080_b0 , \7081_b1 , \7081_b0 , \7082_b1 , \7082_b0 , \7083_b1 , \7083_b0 , \7084_b1 , \7084_b0 , 
		\7085_b1 , \7085_b0 , \7086_b1 , \7086_b0 , \7087_b1 , \7087_b0 , \7088_b1 , \7088_b0 , \7089_b1 , \7089_b0 , 
		\7090_b1 , \7090_b0 , \7091_b1 , \7091_b0 , \7092_b1 , \7092_b0 , \7093_b1 , \7093_b0 , \7094_b1 , \7094_b0 , 
		\7095_b1 , \7095_b0 , \7096_b1 , \7096_b0 , \7097_b1 , \7097_b0 , \7098_b1 , \7098_b0 , \7099_b1 , \7099_b0 , 
		\7100_b1 , \7100_b0 , \7101_b1 , \7101_b0 , \7102_b1 , \7102_b0 , \7103_b1 , \7103_b0 , \7104_b1 , \7104_b0 , 
		\7105_b1 , \7105_b0 , \7106_b1 , \7106_b0 , \7107_b1 , \7107_b0 , \7108_b1 , \7108_b0 , \7109_b1 , \7109_b0 , 
		\7110_b1 , \7110_b0 , \7111_b1 , \7111_b0 , \7112_b1 , \7112_b0 , \7113_b1 , \7113_b0 , \7114_b1 , \7114_b0 , 
		\7115_b1 , \7115_b0 , \7116_b1 , \7116_b0 , \7117_b1 , \7117_b0 , \7118_b1 , \7118_b0 , \7119_b1 , \7119_b0 , 
		\7120_b1 , \7120_b0 , \7121_b1 , \7121_b0 , \7122_b1 , \7122_b0 , \7123_b1 , \7123_b0 , \7124_b1 , \7124_b0 , 
		\7125_b1 , \7125_b0 , \7126_b1 , \7126_b0 , \7127_b1 , \7127_b0 , \7128_b1 , \7128_b0 , \7129_b1 , \7129_b0 , 
		\7130_b1 , \7130_b0 , \7131_b1 , \7131_b0 , \7132_b1 , \7132_b0 , \7133_b1 , \7133_b0 , \7134_b1 , \7134_b0 , 
		\7135_b1 , \7135_b0 , \7136_b1 , \7136_b0 , \7137_b1 , \7137_b0 , \7138_b1 , \7138_b0 , \7139_b1 , \7139_b0 , 
		\7140_b1 , \7140_b0 , \7141_b1 , \7141_b0 , \7142_b1 , \7142_b0 , \7143_b1 , \7143_b0 , \7144_b1 , \7144_b0 , 
		\7145_b1 , \7145_b0 , \7146_b1 , \7146_b0 , \7147_b1 , \7147_b0 , \7148_b1 , \7148_b0 , \7149_b1 , \7149_b0 , 
		\7150_b1 , \7150_b0 , \7151_b1 , \7151_b0 , \7152_b1 , \7152_b0 , \7153_b1 , \7153_b0 , \7154_b1 , \7154_b0 , 
		\7155_b1 , \7155_b0 , \7156_b1 , \7156_b0 , \7157_b1 , \7157_b0 , \7158_b1 , \7158_b0 , \7159_b1 , \7159_b0 , 
		\7160_b1 , \7160_b0 , \7161_b1 , \7161_b0 , \7162_b1 , \7162_b0 , \7163_b1 , \7163_b0 , \7164_b1 , \7164_b0 , 
		\7165_b1 , \7165_b0 , \7166_b1 , \7166_b0 , \7167_b1 , \7167_b0 , \7168_b1 , \7168_b0 , \7169_b1 , \7169_b0 , 
		\7170_b1 , \7170_b0 , \7171_b1 , \7171_b0 , \7172_b1 , \7172_b0 , \7173_b1 , \7173_b0 , \7174_b1 , \7174_b0 , 
		\7175_b1 , \7175_b0 , \7176_b1 , \7176_b0 , \7177_b1 , \7177_b0 , \7178_b1 , \7178_b0 , \7179_b1 , \7179_b0 , 
		\7180_b1 , \7180_b0 , \7181_b1 , \7181_b0 , \7182_b1 , \7182_b0 , \7183_b1 , \7183_b0 , \7184_b1 , \7184_b0 , 
		\7185_b1 , \7185_b0 , \7186_b1 , \7186_b0 , \7187_b1 , \7187_b0 , \7188_b1 , \7188_b0 , \7189_b1 , \7189_b0 , 
		\7190_b1 , \7190_b0 , \7191_b1 , \7191_b0 , \7192_b1 , \7192_b0 , \7193_b1 , \7193_b0 , \7194_b1 , \7194_b0 , 
		\7195_b1 , \7195_b0 , \7196_b1 , \7196_b0 , \7197_b1 , \7197_b0 , \7198_b1 , \7198_b0 , \7199_b1 , \7199_b0 , 
		\7200_b1 , \7200_b0 , \7201_b1 , \7201_b0 , \7202_b1 , \7202_b0 , \7203_b1 , \7203_b0 , \7204_b1 , \7204_b0 , 
		\7205_b1 , \7205_b0 , \7206_b1 , \7206_b0 , \7207_b1 , \7207_b0 , \7208_b1 , \7208_b0 , \7209_b1 , \7209_b0 , 
		\7210_b1 , \7210_b0 , \7211_b1 , \7211_b0 , \7212_b1 , \7212_b0 , \7213_b1 , \7213_b0 , \7214_b1 , \7214_b0 , 
		\7215_b1 , \7215_b0 , \7216_b1 , \7216_b0 , \7217_b1 , \7217_b0 , \7218_b1 , \7218_b0 , \7219_b1 , \7219_b0 , 
		\7220_b1 , \7220_b0 , \7221_b1 , \7221_b0 , \7222_b1 , \7222_b0 , \7223_b1 , \7223_b0 , \7224_b1 , \7224_b0 , 
		\7225_b1 , \7225_b0 , \7226_b1 , \7226_b0 , \7227_b1 , \7227_b0 , \7228_b1 , \7228_b0 , \7229_b1 , \7229_b0 , 
		\7230_b1 , \7230_b0 , \7231_b1 , \7231_b0 , \7232_b1 , \7232_b0 , \7233_b1 , \7233_b0 , \7234_b1 , \7234_b0 , 
		\7235_b1 , \7235_b0 , \7236_b1 , \7236_b0 , \7237_b1 , \7237_b0 , \7238_b1 , \7238_b0 , \7239_b1 , \7239_b0 , 
		\7240_b1 , \7240_b0 , \7241_b1 , \7241_b0 , \7242_b1 , \7242_b0 , \7243_b1 , \7243_b0 , \7244_b1 , \7244_b0 , 
		\7245_b1 , \7245_b0 , \7246_b1 , \7246_b0 , \7247_b1 , \7247_b0 , \7248_b1 , \7248_b0 , \7249_b1 , \7249_b0 , 
		\7250_b1 , \7250_b0 , \7251_b1 , \7251_b0 , \7252_b1 , \7252_b0 , \7253_b1 , \7253_b0 , \7254_b1 , \7254_b0 , 
		\7255_b1 , \7255_b0 , \7256_b1 , \7256_b0 , \7257_b1 , \7257_b0 , \7258_b1 , \7258_b0 , \7259_b1 , \7259_b0 , 
		\7260_b1 , \7260_b0 , \7261_b1 , \7261_b0 , \7262_b1 , \7262_b0 , \7263_b1 , \7263_b0 , \7264_b1 , \7264_b0 , 
		\7265_b1 , \7265_b0 , \7266_b1 , \7266_b0 , \7267_b1 , \7267_b0 , \7268_b1 , \7268_b0 , \7269_b1 , \7269_b0 , 
		\7270_b1 , \7270_b0 , \7271_b1 , \7271_b0 , \7272_b1 , \7272_b0 , \7273_b1 , \7273_b0 , \7274_b1 , \7274_b0 , 
		\7275_b1 , \7275_b0 , \7276_b1 , \7276_b0 , \7277_b1 , \7277_b0 , \7278_b1 , \7278_b0 , \7279_b1 , \7279_b0 , 
		\7280_b1 , \7280_b0 , \7281_b1 , \7281_b0 , \7282_b1 , \7282_b0 , \7283_b1 , \7283_b0 , \7284_b1 , \7284_b0 , 
		\7285_b1 , \7285_b0 , \7286_b1 , \7286_b0 , \7287_b1 , \7287_b0 , \7288_b1 , \7288_b0 , \7289_b1 , \7289_b0 , 
		\7290_b1 , \7290_b0 , \7291_b1 , \7291_b0 , \7292_b1 , \7292_b0 , \7293_b1 , \7293_b0 , \7294_b1 , \7294_b0 , 
		\7295_b1 , \7295_b0 , \7296_b1 , \7296_b0 , \7297_b1 , \7297_b0 , \7298_b1 , \7298_b0 , \7299_b1 , \7299_b0 , 
		\7300_b1 , \7300_b0 , \7301_b1 , \7301_b0 , \7302_b1 , \7302_b0 , \7303_b1 , \7303_b0 , \7304_b1 , \7304_b0 , 
		\7305_b1 , \7305_b0 , \7306_b1 , \7306_b0 , \7307_b1 , \7307_b0 , \7308_b1 , \7308_b0 , \7309_b1 , \7309_b0 , 
		\7310_b1 , \7310_b0 , \7311_b1 , \7311_b0 , \7312_b1 , \7312_b0 , \7313_b1 , \7313_b0 , \7314_b1 , \7314_b0 , 
		\7315_b1 , \7315_b0 , \7316_b1 , \7316_b0 , \7317_b1 , \7317_b0 , \7318_b1 , \7318_b0 , \7319_b1 , \7319_b0 , 
		\7320_b1 , \7320_b0 , \7321_b1 , \7321_b0 , \7322_b1 , \7322_b0 , \7323_b1 , \7323_b0 , \7324_b1 , \7324_b0 , 
		\7325_b1 , \7325_b0 , \7326_b1 , \7326_b0 , \7327_b1 , \7327_b0 , \7328_b1 , \7328_b0 , \7329_b1 , \7329_b0 , 
		\7330_b1 , \7330_b0 , \7331_b1 , \7331_b0 , \7332_b1 , \7332_b0 , \7333_b1 , \7333_b0 , \7334_b1 , \7334_b0 , 
		\7335_b1 , \7335_b0 , \7336_b1 , \7336_b0 , \7337_b1 , \7337_b0 , \7338_b1 , \7338_b0 , \7339_b1 , \7339_b0 , 
		\7340_b1 , \7340_b0 , \7341_b1 , \7341_b0 , \7342_b1 , \7342_b0 , \7343_b1 , \7343_b0 , \7344_b1 , \7344_b0 , 
		\7345_b1 , \7345_b0 , \7346_b1 , \7346_b0 , \7347_b1 , \7347_b0 , \7348_b1 , \7348_b0 , \7349_b1 , \7349_b0 , 
		\7350_b1 , \7350_b0 , \7351_b1 , \7351_b0 , \7352_b1 , \7352_b0 , \7353_b1 , \7353_b0 , \7354_b1 , \7354_b0 , 
		\7355_b1 , \7355_b0 , \7356_b1 , \7356_b0 , \7357_b1 , \7357_b0 , \7358_b1 , \7358_b0 , \7359_b1 , \7359_b0 , 
		\7360_b1 , \7360_b0 , \7361_b1 , \7361_b0 , \7362_b1 , \7362_b0 , \7363_b1 , \7363_b0 , \7364_b1 , \7364_b0 , 
		\7365_b1 , \7365_b0 , \7366_b1 , \7366_b0 , \7367_b1 , \7367_b0 , \7368_b1 , \7368_b0 , \7369_b1 , \7369_b0 , 
		\7370_b1 , \7370_b0 , \7371_b1 , \7371_b0 , \7372_b1 , \7372_b0 , \7373_b1 , \7373_b0 , \7374_b1 , \7374_b0 , 
		\7375_b1 , \7375_b0 , \7376_b1 , \7376_b0 , \7377_b1 , \7377_b0 , \7378_b1 , \7378_b0 , \7379_b1 , \7379_b0 , 
		\7380_b1 , \7380_b0 , \7381_b1 , \7381_b0 , \7382_b1 , \7382_b0 , \7383_b1 , \7383_b0 , \7384_b1 , \7384_b0 , 
		\7385_b1 , \7385_b0 , \7386_b1 , \7386_b0 , \7387_b1 , \7387_b0 , \7388_b1 , \7388_b0 , \7389_b1 , \7389_b0 , 
		\7390_b1 , \7390_b0 , \7391_b1 , \7391_b0 , \7392_b1 , \7392_b0 , \7393_b1 , \7393_b0 , \7394_b1 , \7394_b0 , 
		\7395_b1 , \7395_b0 , \7396_b1 , \7396_b0 , \7397_b1 , \7397_b0 , \7398_b1 , \7398_b0 , \7399_b1 , \7399_b0 , 
		\7400_b1 , \7400_b0 , \7401_b1 , \7401_b0 , \7402_b1 , \7402_b0 , \7403_b1 , \7403_b0 , \7404_b1 , \7404_b0 , 
		\7405_b1 , \7405_b0 , \7406_b1 , \7406_b0 , \7407_b1 , \7407_b0 , \7408_b1 , \7408_b0 , \7409_b1 , \7409_b0 , 
		\7410_b1 , \7410_b0 , \7411_b1 , \7411_b0 , \7412_b1 , \7412_b0 , \7413_b1 , \7413_b0 , \7414_b1 , \7414_b0 , 
		\7415_b1 , \7415_b0 , \7416_b1 , \7416_b0 , \7417_b1 , \7417_b0 , \7418_b1 , \7418_b0 , \7419_b1 , \7419_b0 , 
		\7420_b1 , \7420_b0 , \7421_b1 , \7421_b0 , \7422_b1 , \7422_b0 , \7423_b1 , \7423_b0 , \7424_b1 , \7424_b0 , 
		\7425_b1 , \7425_b0 , \7426_b1 , \7426_b0 , \7427_b1 , \7427_b0 , \7428_b1 , \7428_b0 , \7429_b1 , \7429_b0 , 
		\7430_b1 , \7430_b0 , \7431_b1 , \7431_b0 , \7432_b1 , \7432_b0 , \7433_b1 , \7433_b0 , \7434_b1 , \7434_b0 , 
		\7435_b1 , \7435_b0 , \7436_b1 , \7436_b0 , \7437_b1 , \7437_b0 , \7438_b1 , \7438_b0 , \7439_b1 , \7439_b0 , 
		\7440_b1 , \7440_b0 , \7441_b1 , \7441_b0 , \7442_b1 , \7442_b0 , \7443_b1 , \7443_b0 , \7444_b1 , \7444_b0 , 
		\7445_b1 , \7445_b0 , \7446_b1 , \7446_b0 , \7447_b1 , \7447_b0 , \7448_b1 , \7448_b0 , \7449_b1 , \7449_b0 , 
		\7450_b1 , \7450_b0 , \7451_b1 , \7451_b0 , \7452_b1 , \7452_b0 , \7453_b1 , \7453_b0 , \7454_b1 , \7454_b0 , 
		\7455_b1 , \7455_b0 , \7456_b1 , \7456_b0 , \7457_b1 , \7457_b0 , \7458_b1 , \7458_b0 , \7459_b1 , \7459_b0 , 
		\7460_b1 , \7460_b0 , \7461_b1 , \7461_b0 , \7462_b1 , \7462_b0 , \7463_b1 , \7463_b0 , \7464_b1 , \7464_b0 , 
		\7465_b1 , \7465_b0 , \7466_b1 , \7466_b0 , \7467_b1 , \7467_b0 , \7468_b1 , \7468_b0 , \7469_b1 , \7469_b0 , 
		\7470_b1 , \7470_b0 , \7471_b1 , \7471_b0 , \7472_b1 , \7472_b0 , \7473_b1 , \7473_b0 , \7474_b1 , \7474_b0 , 
		\7475_b1 , \7475_b0 , \7476_b1 , \7476_b0 , \7477_b1 , \7477_b0 , \7478_b1 , \7478_b0 , \7479_b1 , \7479_b0 , 
		\7480_b1 , \7480_b0 , \7481_b1 , \7481_b0 , \7482_b1 , \7482_b0 , \7483_b1 , \7483_b0 , \7484_b1 , \7484_b0 , 
		\7485_b1 , \7485_b0 , \7486_b1 , \7486_b0 , \7487_b1 , \7487_b0 , \7488_b1 , \7488_b0 , \7489_b1 , \7489_b0 , 
		\7490_b1 , \7490_b0 , \7491_b1 , \7491_b0 , \7492_b1 , \7492_b0 , \7493_b1 , \7493_b0 , \7494_b1 , \7494_b0 , 
		\7495_b1 , \7495_b0 , \7496_b1 , \7496_b0 , \7497_b1 , \7497_b0 , \7498_b1 , \7498_b0 , \7499_b1 , \7499_b0 , 
		\7500_b1 , \7500_b0 , \7501_b1 , \7501_b0 , \7502_b1 , \7502_b0 , \7503_b1 , \7503_b0 , \7504_b1 , \7504_b0 , 
		\7505_b1 , \7505_b0 , \7506_b1 , \7506_b0 , \7507_b1 , \7507_b0 , \7508_b1 , \7508_b0 , \7509_b1 , \7509_b0 , 
		\7510_b1 , \7510_b0 , \7511_b1 , \7511_b0 , \7512_b1 , \7512_b0 , \7513_b1 , \7513_b0 , \7514_b1 , \7514_b0 , 
		\7515_b1 , \7515_b0 , \7516_b1 , \7516_b0 , \7517_b1 , \7517_b0 , \7518_b1 , \7518_b0 , \7519_b1 , \7519_b0 , 
		\7520_b1 , \7520_b0 , \7521_b1 , \7521_b0 , \7522_b1 , \7522_b0 , \7523_b1 , \7523_b0 , \7524_b1 , \7524_b0 , 
		\7525_b1 , \7525_b0 , \7526_b1 , \7526_b0 , \7527_b1 , \7527_b0 , \7528_b1 , \7528_b0 , \7529_b1 , \7529_b0 , 
		\7530_b1 , \7530_b0 , \7531_b1 , \7531_b0 , \7532_b1 , \7532_b0 , \7533_b1 , \7533_b0 , \7534_b1 , \7534_b0 , 
		\7535_b1 , \7535_b0 , \7536_b1 , \7536_b0 , \7537_b1 , \7537_b0 , \7538_b1 , \7538_b0 , \7539_b1 , \7539_b0 , 
		\7540_b1 , \7540_b0 , \7541_b1 , \7541_b0 , \7542_b1 , \7542_b0 , \7543_b1 , \7543_b0 , \7544_b1 , \7544_b0 , 
		\7545_b1 , \7545_b0 , \7546_b1 , \7546_b0 , \7547_b1 , \7547_b0 , \7548_b1 , \7548_b0 , \7549_b1 , \7549_b0 , 
		\7550_b1 , \7550_b0 , \7551_b1 , \7551_b0 , \7552_b1 , \7552_b0 , \7553_b1 , \7553_b0 , \7554_b1 , \7554_b0 , 
		\7555_b1 , \7555_b0 , \7556_b1 , \7556_b0 , \7557_b1 , \7557_b0 , \7558_b1 , \7558_b0 , \7559_b1 , \7559_b0 , 
		\7560_b1 , \7560_b0 , \7561_b1 , \7561_b0 , \7562_b1 , \7562_b0 , \7563_b1 , \7563_b0 , \7564_b1 , \7564_b0 , 
		\7565_b1 , \7565_b0 , \7566_b1 , \7566_b0 , \7567_b1 , \7567_b0 , \7568_b1 , \7568_b0 , \7569_b1 , \7569_b0 , 
		\7570_b1 , \7570_b0 , \7571_b1 , \7571_b0 , \7572_b1 , \7572_b0 , \7573_b1 , \7573_b0 , \7574_b1 , \7574_b0 , 
		\7575_b1 , \7575_b0 , \7576_b1 , \7576_b0 , \7577_b1 , \7577_b0 , \7578_b1 , \7578_b0 , \7579_b1 , \7579_b0 , 
		\7580_b1 , \7580_b0 , \7581_b1 , \7581_b0 , \7582_b1 , \7582_b0 , \7583_b1 , \7583_b0 , \7584_b1 , \7584_b0 , 
		\7585_b1 , \7585_b0 , \7586_b1 , \7586_b0 , \7587_b1 , \7587_b0 , \7588_b1 , \7588_b0 , \7589_b1 , \7589_b0 , 
		\7590_b1 , \7590_b0 , \7591_b1 , \7591_b0 , \7592_b1 , \7592_b0 , \7593_b1 , \7593_b0 , \7594_b1 , \7594_b0 , 
		\7595_b1 , \7595_b0 , \7596_b1 , \7596_b0 , \7597_b1 , \7597_b0 , \7598_b1 , \7598_b0 , \7599_b1 , \7599_b0 , 
		\7600_b1 , \7600_b0 , \7601_b1 , \7601_b0 , \7602_b1 , \7602_b0 , \7603_b1 , \7603_b0 , \7604_b1 , \7604_b0 , 
		\7605_b1 , \7605_b0 , \7606_b1 , \7606_b0 , \7607_b1 , \7607_b0 , \7608_b1 , \7608_b0 , \7609_b1 , \7609_b0 , 
		\7610_b1 , \7610_b0 , \7611_b1 , \7611_b0 , \7612_b1 , \7612_b0 , \7613_b1 , \7613_b0 , \7614_b1 , \7614_b0 , 
		\7615_b1 , \7615_b0 , \7616_b1 , \7616_b0 , \7617_b1 , \7617_b0 , \7618_b1 , \7618_b0 , \7619_b1 , \7619_b0 , 
		\7620_b1 , \7620_b0 , \7621_b1 , \7621_b0 , \7622_b1 , \7622_b0 , \7623_b1 , \7623_b0 , \7624_b1 , \7624_b0 , 
		\7625_b1 , \7625_b0 , \7626_b1 , \7626_b0 , \7627_b1 , \7627_b0 , \7628_b1 , \7628_b0 , \7629_b1 , \7629_b0 , 
		\7630_b1 , \7630_b0 , \7631_b1 , \7631_b0 , \7632_b1 , \7632_b0 , \7633_b1 , \7633_b0 , \7634_b1 , \7634_b0 , 
		\7635_b1 , \7635_b0 , \7636_b1 , \7636_b0 , \7637_b1 , \7637_b0 , \7638_b1 , \7638_b0 , \7639_b1 , \7639_b0 , 
		\7640_b1 , \7640_b0 , \7641_b1 , \7641_b0 , \7642_b1 , \7642_b0 , \7643_b1 , \7643_b0 , \7644_b1 , \7644_b0 , 
		\7645_b1 , \7645_b0 , \7646_b1 , \7646_b0 , \7647_b1 , \7647_b0 , \7648_b1 , \7648_b0 , \7649_b1 , \7649_b0 , 
		\7650_b1 , \7650_b0 , \7651_b1 , \7651_b0 , \7652_b1 , \7652_b0 , \7653_b1 , \7653_b0 , \7654_b1 , \7654_b0 , 
		\7655_b1 , \7655_b0 , \7656_b1 , \7656_b0 , \7657_b1 , \7657_b0 , \7658_b1 , \7658_b0 , \7659_b1 , \7659_b0 , 
		\7660_b1 , \7660_b0 , \7661_b1 , \7661_b0 , \7662_b1 , \7662_b0 , \7663_b1 , \7663_b0 , \7664_b1 , \7664_b0 , 
		\7665_b1 , \7665_b0 , \7666_b1 , \7666_b0 , \7667_b1 , \7667_b0 , \7668_b1 , \7668_b0 , \7669_b1 , \7669_b0 , 
		\7670_b1 , \7670_b0 , \7671_b1 , \7671_b0 , \7672_b1 , \7672_b0 , \7673_b1 , \7673_b0 , \7674_b1 , \7674_b0 , 
		\7675_b1 , \7675_b0 , \7676_b1 , \7676_b0 , \7677_b1 , \7677_b0 , \7678_b1 , \7678_b0 , \7679_b1 , \7679_b0 , 
		\7680_b1 , \7680_b0 , \7681_b1 , \7681_b0 , \7682_b1 , \7682_b0 , \7683_b1 , \7683_b0 , \7684_b1 , \7684_b0 , 
		\7685_b1 , \7685_b0 , \7686_b1 , \7686_b0 , \7687_b1 , \7687_b0 , \7688_b1 , \7688_b0 , \7689_b1 , \7689_b0 , 
		\7690_b1 , \7690_b0 , \7691_b1 , \7691_b0 , \7692_b1 , \7692_b0 , \7693_b1 , \7693_b0 , \7694_b1 , \7694_b0 , 
		\7695_b1 , \7695_b0 , \7696_b1 , \7696_b0 , \7697_b1 , \7697_b0 , \7698_b1 , \7698_b0 , \7699_b1 , \7699_b0 , 
		\7700_b1 , \7700_b0 , \7701_b1 , \7701_b0 , \7702_b1 , \7702_b0 , \7703_b1 , \7703_b0 , \7704_b1 , \7704_b0 , 
		\7705_b1 , \7705_b0 , \7706_b1 , \7706_b0 , \7707_b1 , \7707_b0 , \7708_b1 , \7708_b0 , \7709_b1 , \7709_b0 , 
		\7710_b1 , \7710_b0 , \7711_b1 , \7711_b0 , \7712_b1 , \7712_b0 , \7713_b1 , \7713_b0 , \7714_b1 , \7714_b0 , 
		\7715_b1 , \7715_b0 , \7716_b1 , \7716_b0 , \7717_b1 , \7717_b0 , \7718_b1 , \7718_b0 , \7719_b1 , \7719_b0 , 
		\7720_b1 , \7720_b0 , \7721_b1 , \7721_b0 , \7722_b1 , \7722_b0 , \7723_b1 , \7723_b0 , \7724_b1 , \7724_b0 , 
		\7725_b1 , \7725_b0 , \7726_b1 , \7726_b0 , \7727_b1 , \7727_b0 , \7728_b1 , \7728_b0 , \7729_b1 , \7729_b0 , 
		\7730_b1 , \7730_b0 , \7731_b1 , \7731_b0 , \7732_b1 , \7732_b0 , \7733_b1 , \7733_b0 , \7734_b1 , \7734_b0 , 
		\7735_b1 , \7735_b0 , \7736_b1 , \7736_b0 , \7737_b1 , \7737_b0 , \7738_b1 , \7738_b0 , \7739_b1 , \7739_b0 , 
		\7740_b1 , \7740_b0 , \7741_b1 , \7741_b0 , \7742_b1 , \7742_b0 , \7743_b1 , \7743_b0 , \7744_b1 , \7744_b0 , 
		\7745_b1 , \7745_b0 , \7746_b1 , \7746_b0 , \7747_b1 , \7747_b0 , \7748_b1 , \7748_b0 , \7749_b1 , \7749_b0 , 
		\7750_b1 , \7750_b0 , \7751_b1 , \7751_b0 , \7752_b1 , \7752_b0 , \7753_b1 , \7753_b0 , \7754_b1 , \7754_b0 , 
		\7755_b1 , \7755_b0 , \7756_b1 , \7756_b0 , \7757_b1 , \7757_b0 , \7758_b1 , \7758_b0 , \7759_b1 , \7759_b0 , 
		\7760_b1 , \7760_b0 , \7761_b1 , \7761_b0 , \7762_b1 , \7762_b0 , \7763_b1 , \7763_b0 , \7764_b1 , \7764_b0 , 
		\7765_b1 , \7765_b0 , \7766_b1 , \7766_b0 , \7767_b1 , \7767_b0 , \7768_b1 , \7768_b0 , \7769_b1 , \7769_b0 , 
		\7770_b1 , \7770_b0 , \7771_b1 , \7771_b0 , \7772_b1 , \7772_b0 , \7773_b1 , \7773_b0 , \7774_b1 , \7774_b0 , 
		\7775_b1 , \7775_b0 , \7776_b1 , \7776_b0 , \7777_b1 , \7777_b0 , \7778_b1 , \7778_b0 , \7779_b1 , \7779_b0 , 
		\7780_b1 , \7780_b0 , \7781_b1 , \7781_b0 , \7782_b1 , \7782_b0 , \7783_b1 , \7783_b0 , \7784_b1 , \7784_b0 , 
		\7785_b1 , \7785_b0 , \7786_b1 , \7786_b0 , \7787_b1 , \7787_b0 , \7788_b1 , \7788_b0 , \7789_b1 , \7789_b0 , 
		\7790_b1 , \7790_b0 , \7791_b1 , \7791_b0 , \7792_b1 , \7792_b0 , \7793_b1 , \7793_b0 , \7794_b1 , \7794_b0 , 
		\7795_b1 , \7795_b0 , \7796_b1 , \7796_b0 , \7797_b1 , \7797_b0 , \7798_b1 , \7798_b0 , \7799_b1 , \7799_b0 , 
		\7800_b1 , \7800_b0 , \7801_b1 , \7801_b0 , \7802_b1 , \7802_b0 , \7803_b1 , \7803_b0 , \7804_b1 , \7804_b0 , 
		\7805_b1 , \7805_b0 , \7806_b1 , \7806_b0 , \7807_b1 , \7807_b0 , \7808_b1 , \7808_b0 , \7809_b1 , \7809_b0 , 
		\7810_b1 , \7810_b0 , \7811_b1 , \7811_b0 , \7812_b1 , \7812_b0 , \7813_b1 , \7813_b0 , \7814_b1 , \7814_b0 , 
		\7815_b1 , \7815_b0 , \7816_b1 , \7816_b0 , \7817_b1 , \7817_b0 , \7818_b1 , \7818_b0 , \7819_b1 , \7819_b0 , 
		\7820_b1 , \7820_b0 , \7821_b1 , \7821_b0 , \7822_b1 , \7822_b0 , \7823_b1 , \7823_b0 , \7824_b1 , \7824_b0 , 
		\7825_b1 , \7825_b0 , \7826_b1 , \7826_b0 , \7827_b1 , \7827_b0 , \7828_b1 , \7828_b0 , \7829_b1 , \7829_b0 , 
		\7830_b1 , \7830_b0 , \7831_b1 , \7831_b0 , \7832_b1 , \7832_b0 , \7833_b1 , \7833_b0 , \7834_b1 , \7834_b0 , 
		\7835_b1 , \7835_b0 , \7836_b1 , \7836_b0 , \7837_b1 , \7837_b0 , \7838_b1 , \7838_b0 , \7839_b1 , \7839_b0 , 
		\7840_b1 , \7840_b0 , \7841_b1 , \7841_b0 , \7842_b1 , \7842_b0 , \7843_b1 , \7843_b0 , \7844_b1 , \7844_b0 , 
		\7845_b1 , \7845_b0 , \7846_b1 , \7846_b0 , \7847_b1 , \7847_b0 , \7848_b1 , \7848_b0 , \7849_b1 , \7849_b0 , 
		\7850_b1 , \7850_b0 , \7851_b1 , \7851_b0 , \7852_b1 , \7852_b0 , \7853_b1 , \7853_b0 , \7854_b1 , \7854_b0 , 
		\7855_b1 , \7855_b0 , \7856_b1 , \7856_b0 , \7857_b1 , \7857_b0 , \7858_b1 , \7858_b0 , \7859_b1 , \7859_b0 , 
		\7860_b1 , \7860_b0 , \7861_b1 , \7861_b0 , \7862_b1 , \7862_b0 , \7863_b1 , \7863_b0 , \7864_b1 , \7864_b0 , 
		\7865_b1 , \7865_b0 , \7866_b1 , \7866_b0 , \7867_b1 , \7867_b0 , \7868_b1 , \7868_b0 , \7869_b1 , \7869_b0 , 
		\7870_b1 , \7870_b0 , \7871_b1 , \7871_b0 , \7872_b1 , \7872_b0 , \7873_b1 , \7873_b0 , \7874_b1 , \7874_b0 , 
		\7875_b1 , \7875_b0 , \7876_b1 , \7876_b0 , \7877_b1 , \7877_b0 , \7878_b1 , \7878_b0 , \7879_b1 , \7879_b0 , 
		\7880_b1 , \7880_b0 , \7881_b1 , \7881_b0 , \7882_b1 , \7882_b0 , \7883_b1 , \7883_b0 , \7884_b1 , \7884_b0 , 
		\7885_b1 , \7885_b0 , \7886_b1 , \7886_b0 , \7887_b1 , \7887_b0 , \7888_b1 , \7888_b0 , \7889_b1 , \7889_b0 , 
		\7890_b1 , \7890_b0 , \7891_b1 , \7891_b0 , \7892_b1 , \7892_b0 , \7893_b1 , \7893_b0 , \7894_b1 , \7894_b0 , 
		\7895_b1 , \7895_b0 , \7896_b1 , \7896_b0 , \7897_b1 , \7897_b0 , \7898_b1 , \7898_b0 , \7899_b1 , \7899_b0 , 
		\7900_b1 , \7900_b0 , \7901_b1 , \7901_b0 , \7902_b1 , \7902_b0 , \7903_b1 , \7903_b0 , \7904_b1 , \7904_b0 , 
		\7905_b1 , \7905_b0 , \7906_b1 , \7906_b0 , \7907_b1 , \7907_b0 , \7908_b1 , \7908_b0 , \7909_b1 , \7909_b0 , 
		\7910_b1 , \7910_b0 , \7911_b1 , \7911_b0 , \7912_b1 , \7912_b0 , \7913_b1 , \7913_b0 , \7914_b1 , \7914_b0 , 
		\7915_b1 , \7915_b0 , \7916_b1 , \7916_b0 , \7917_b1 , \7917_b0 , \7918_b1 , \7918_b0 , \7919_b1 , \7919_b0 , 
		\7920_b1 , \7920_b0 , \7921_b1 , \7921_b0 , \7922_b1 , \7922_b0 , \7923_b1 , \7923_b0 , \7924_b1 , \7924_b0 , 
		\7925_b1 , \7925_b0 , \7926_b1 , \7926_b0 , \7927_b1 , \7927_b0 , \7928_b1 , \7928_b0 , \7929_b1 , \7929_b0 , 
		\7930_b1 , \7930_b0 , \7931_b1 , \7931_b0 , \7932_b1 , \7932_b0 , \7933_b1 , \7933_b0 , \7934_b1 , \7934_b0 , 
		\7935_b1 , \7935_b0 , \7936_b1 , \7936_b0 , \7937_b1 , \7937_b0 , \7938_b1 , \7938_b0 , \7939_b1 , \7939_b0 , 
		\7940_b1 , \7940_b0 , \7941_b1 , \7941_b0 , \7942_b1 , \7942_b0 , \7943_b1 , \7943_b0 , \7944_b1 , \7944_b0 , 
		\7945_b1 , \7945_b0 , \7946_b1 , \7946_b0 , \7947_b1 , \7947_b0 , \7948_b1 , \7948_b0 , \7949_b1 , \7949_b0 , 
		\7950_b1 , \7950_b0 , \7951_b1 , \7951_b0 , \7952_b1 , \7952_b0 , \7953_b1 , \7953_b0 , \7954_b1 , \7954_b0 , 
		\7955_b1 , \7955_b0 , \7956_b1 , \7956_b0 , \7957_b1 , \7957_b0 , \7958_b1 , \7958_b0 , \7959_b1 , \7959_b0 , 
		\7960_b1 , \7960_b0 , \7961_b1 , \7961_b0 , \7962_b1 , \7962_b0 , \7963_b1 , \7963_b0 , \7964_b1 , \7964_b0 , 
		\7965_b1 , \7965_b0 , \7966_b1 , \7966_b0 , \7967_b1 , \7967_b0 , \7968_b1 , \7968_b0 , \7969_b1 , \7969_b0 , 
		\7970_b1 , \7970_b0 , \7971_b1 , \7971_b0 , \7972_b1 , \7972_b0 , \7973_b1 , \7973_b0 , \7974_b1 , \7974_b0 , 
		\7975_b1 , \7975_b0 , \7976_b1 , \7976_b0 , \7977_b1 , \7977_b0 , \7978_b1 , \7978_b0 , \7979_b1 , \7979_b0 , 
		\7980_b1 , \7980_b0 , \7981_b1 , \7981_b0 , \7982_b1 , \7982_b0 , \7983_b1 , \7983_b0 , \7984_b1 , \7984_b0 , 
		\7985_b1 , \7985_b0 , \7986_b1 , \7986_b0 , \7987_b1 , \7987_b0 , \7988_b1 , \7988_b0 , \7989_b1 , \7989_b0 , 
		\7990_b1 , \7990_b0 , \7991_b1 , \7991_b0 , \7992_b1 , \7992_b0 , \7993_b1 , \7993_b0 , \7994_b1 , \7994_b0 , 
		\7995_b1 , \7995_b0 , \7996_b1 , \7996_b0 , \7997_b1 , \7997_b0 , \7998_b1 , \7998_b0 , \7999_b1 , \7999_b0 , 
		\8000_b1 , \8000_b0 , \8001_b1 , \8001_b0 , \8002_b1 , \8002_b0 , \8003_b1 , \8003_b0 , \8004_b1 , \8004_b0 , 
		\8005_b1 , \8005_b0 , \8006_b1 , \8006_b0 , \8007_b1 , \8007_b0 , \8008_b1 , \8008_b0 , \8009_b1 , \8009_b0 , 
		\8010_b1 , \8010_b0 , \8011_b1 , \8011_b0 , \8012_b1 , \8012_b0 , \8013_b1 , \8013_b0 , \8014_b1 , \8014_b0 , 
		\8015_b1 , \8015_b0 , \8016_b1 , \8016_b0 , \8017_b1 , \8017_b0 , \8018_b1 , \8018_b0 , \8019_b1 , \8019_b0 , 
		\8020_b1 , \8020_b0 , \8021_b1 , \8021_b0 , \8022_b1 , \8022_b0 , \8023_b1 , \8023_b0 , \8024_b1 , \8024_b0 , 
		\8025_b1 , \8025_b0 , \8026_b1 , \8026_b0 , \8027_b1 , \8027_b0 , \8028_b1 , \8028_b0 , \8029_b1 , \8029_b0 , 
		\8030_b1 , \8030_b0 , \8031_b1 , \8031_b0 , \8032_b1 , \8032_b0 , \8033_b1 , \8033_b0 , \8034_b1 , \8034_b0 , 
		\8035_b1 , \8035_b0 , \8036_b1 , \8036_b0 , \8037_b1 , \8037_b0 , \8038_b1 , \8038_b0 , \8039_b1 , \8039_b0 , 
		\8040_b1 , \8040_b0 , \8041_b1 , \8041_b0 , \8042_b1 , \8042_b0 , \8043_b1 , \8043_b0 , \8044_b1 , \8044_b0 , 
		\8045_b1 , \8045_b0 , \8046_b1 , \8046_b0 , \8047_b1 , \8047_b0 , \8048_b1 , \8048_b0 , \8049_b1 , \8049_b0 , 
		\8050_b1 , \8050_b0 , \8051_b1 , \8051_b0 , \8052_b1 , \8052_b0 , \8053_b1 , \8053_b0 , \8054_b1 , \8054_b0 , 
		\8055_b1 , \8055_b0 , \8056_b1 , \8056_b0 , \8057_b1 , \8057_b0 , \8058_b1 , \8058_b0 , \8059_b1 , \8059_b0 , 
		\8060_b1 , \8060_b0 , \8061_b1 , \8061_b0 , \8062_b1 , \8062_b0 , \8063_b1 , \8063_b0 , \8064_b1 , \8064_b0 , 
		\8065_b1 , \8065_b0 , \8066_b1 , \8066_b0 , \8067_b1 , \8067_b0 , \8068_b1 , \8068_b0 , \8069_b1 , \8069_b0 , 
		\8070_b1 , \8070_b0 , \8071_b1 , \8071_b0 , \8072_b1 , \8072_b0 , \8073_b1 , \8073_b0 , \8074_b1 , \8074_b0 , 
		\8075_b1 , \8075_b0 , \8076_b1 , \8076_b0 , \8077_b1 , \8077_b0 , \8078_b1 , \8078_b0 , \8079_b1 , \8079_b0 , 
		\8080_b1 , \8080_b0 , \8081_b1 , \8081_b0 , \8082_b1 , \8082_b0 , \8083_b1 , \8083_b0 , \8084_b1 , \8084_b0 , 
		\8085_b1 , \8085_b0 , \8086_b1 , \8086_b0 , \8087_b1 , \8087_b0 , \8088_b1 , \8088_b0 , \8089_b1 , \8089_b0 , 
		\8090_b1 , \8090_b0 , \8091_b1 , \8091_b0 , \8092_b1 , \8092_b0 , \8093_b1 , \8093_b0 , \8094_b1 , \8094_b0 , 
		\8095_b1 , \8095_b0 , \8096_b1 , \8096_b0 , \8097_b1 , \8097_b0 , \8098_b1 , \8098_b0 , \8099_b1 , \8099_b0 , 
		\8100_b1 , \8100_b0 , \8101_b1 , \8101_b0 , \8102_b1 , \8102_b0 , \8103_b1 , \8103_b0 , \8104_b1 , \8104_b0 , 
		\8105_b1 , \8105_b0 , \8106_b1 , \8106_b0 , \8107_b1 , \8107_b0 , \8108_b1 , \8108_b0 , \8109_b1 , \8109_b0 , 
		\8110_b1 , \8110_b0 , \8111_b1 , \8111_b0 , \8112_b1 , \8112_b0 , \8113_b1 , \8113_b0 , \8114_b1 , \8114_b0 , 
		\8115_b1 , \8115_b0 , \8116_b1 , \8116_b0 , \8117_b1 , \8117_b0 , \8118_b1 , \8118_b0 , \8119_b1 , \8119_b0 , 
		\8120_b1 , \8120_b0 , \8121_b1 , \8121_b0 , \8122_b1 , \8122_b0 , \8123_b1 , \8123_b0 , \8124_b1 , \8124_b0 , 
		\8125_b1 , \8125_b0 , \8126_b1 , \8126_b0 , \8127_b1 , \8127_b0 , \8128_b1 , \8128_b0 , \8129_b1 , \8129_b0 , 
		\8130_b1 , \8130_b0 , \8131_b1 , \8131_b0 , \8132_b1 , \8132_b0 , \8133_b1 , \8133_b0 , \8134_b1 , \8134_b0 , 
		\8135_b1 , \8135_b0 , \8136_b1 , \8136_b0 , \8137_b1 , \8137_b0 , \8138_b1 , \8138_b0 , \8139_b1 , \8139_b0 , 
		\8140_b1 , \8140_b0 , \8141_b1 , \8141_b0 , \8142_b1 , \8142_b0 , \8143_b1 , \8143_b0 , \8144_b1 , \8144_b0 , 
		\8145_b1 , \8145_b0 , \8146_b1 , \8146_b0 , \8147_b1 , \8147_b0 , \8148_b1 , \8148_b0 , \8149_b1 , \8149_b0 , 
		\8150_b1 , \8150_b0 , \8151_b1 , \8151_b0 , \8152_b1 , \8152_b0 , \8153_b1 , \8153_b0 , \8154_b1 , \8154_b0 , 
		\8155_b1 , \8155_b0 , \8156_b1 , \8156_b0 , \8157_b1 , \8157_b0 , \8158_b1 , \8158_b0 , \8159_b1 , \8159_b0 , 
		\8160_b1 , \8160_b0 , \8161_b1 , \8161_b0 , \8162_b1 , \8162_b0 , \8163_b1 , \8163_b0 , \8164_b1 , \8164_b0 , 
		\8165_b1 , \8165_b0 , \8166_b1 , \8166_b0 , \8167_b1 , \8167_b0 , \8168_b1 , \8168_b0 , \8169_b1 , \8169_b0 , 
		\8170_b1 , \8170_b0 , \8171_b1 , \8171_b0 , \8172_b1 , \8172_b0 , \8173_b1 , \8173_b0 , \8174_b1 , \8174_b0 , 
		\8175_b1 , \8175_b0 , \8176_b1 , \8176_b0 , \8177_b1 , \8177_b0 , \8178_b1 , \8178_b0 , \8179_b1 , \8179_b0 , 
		\8180_b1 , \8180_b0 , \8181_b1 , \8181_b0 , \8182_b1 , \8182_b0 , \8183_b1 , \8183_b0 , \8184_b1 , \8184_b0 , 
		\8185_b1 , \8185_b0 , \8186_b1 , \8186_b0 , \8187_b1 , \8187_b0 , \8188_b1 , \8188_b0 , \8189_b1 , \8189_b0 , 
		\8190_b1 , \8190_b0 , \8191_b1 , \8191_b0 , \8192_b1 , \8192_b0 , \8193_b1 , \8193_b0 , \8194_b1 , \8194_b0 , 
		\8195_b1 , \8195_b0 , \8196_b1 , \8196_b0 , \8197_b1 , \8197_b0 , \8198_b1 , \8198_b0 , \8199_b1 , \8199_b0 , 
		\8200_b1 , \8200_b0 , \8201_b1 , \8201_b0 , \8202_b1 , \8202_b0 , \8203_b1 , \8203_b0 , \8204_b1 , \8204_b0 , 
		\8205_b1 , \8205_b0 , \8206_b1 , \8206_b0 , \8207_b1 , \8207_b0 , \8208_b1 , \8208_b0 , \8209_b1 , \8209_b0 , 
		\8210_b1 , \8210_b0 , \8211_b1 , \8211_b0 , \8212_b1 , \8212_b0 , \8213_b1 , \8213_b0 , \8214_b1 , \8214_b0 , 
		\8215_b1 , \8215_b0 , \8216_b1 , \8216_b0 , \8217_b1 , \8217_b0 , \8218_b1 , \8218_b0 , \8219_b1 , \8219_b0 , 
		\8220_b1 , \8220_b0 , \8221_b1 , \8221_b0 , \8222_b1 , \8222_b0 , \8223_b1 , \8223_b0 , \8224_b1 , \8224_b0 , 
		\8225_b1 , \8225_b0 , \8226_b1 , \8226_b0 , \8227_b1 , \8227_b0 , \8228_b1 , \8228_b0 , \8229_b1 , \8229_b0 , 
		\8230_b1 , \8230_b0 , \8231_b1 , \8231_b0 , \8232_b1 , \8232_b0 , \8233_b1 , \8233_b0 , \8234_b1 , \8234_b0 , 
		\8235_b1 , \8235_b0 , \8236_b1 , \8236_b0 , \8237_b1 , \8237_b0 , \8238_b1 , \8238_b0 , \8239_b1 , \8239_b0 , 
		\8240_b1 , \8240_b0 , \8241_b1 , \8241_b0 , \8242_b1 , \8242_b0 , \8243_b1 , \8243_b0 , \8244_b1 , \8244_b0 , 
		\8245_b1 , \8245_b0 , \8246_b1 , \8246_b0 , \8247_b1 , \8247_b0 , \8248_b1 , \8248_b0 , \8249_b1 , \8249_b0 , 
		\8250_b1 , \8250_b0 , \8251_b1 , \8251_b0 , \8252_b1 , \8252_b0 , \8253_b1 , \8253_b0 , \8254_b1 , \8254_b0 , 
		\8255_b1 , \8255_b0 , \8256_b1 , \8256_b0 , \8257_b1 , \8257_b0 , \8258_b1 , \8258_b0 , \8259_b1 , \8259_b0 , 
		\8260_b1 , \8260_b0 , \8261_b1 , \8261_b0 , \8262_b1 , \8262_b0 , \8263_b1 , \8263_b0 , \8264_b1 , \8264_b0 , 
		\8265_b1 , \8265_b0 , \8266_b1 , \8266_b0 , \8267_b1 , \8267_b0 , \8268_b1 , \8268_b0 , \8269_b1 , \8269_b0 , 
		\8270_b1 , \8270_b0 , \8271_b1 , \8271_b0 , \8272_b1 , \8272_b0 , \8273_b1 , \8273_b0 , \8274_b1 , \8274_b0 , 
		\8275_b1 , \8275_b0 , \8276_b1 , \8276_b0 , \8277_b1 , \8277_b0 , \8278_b1 , \8278_b0 , \8279_b1 , \8279_b0 , 
		\8280_b1 , \8280_b0 , \8281_b1 , \8281_b0 , \8282_b1 , \8282_b0 , \8283_b1 , \8283_b0 , \8284_b1 , \8284_b0 , 
		\8285_b1 , \8285_b0 , \8286_b1 , \8286_b0 , \8287_b1 , \8287_b0 , \8288_b1 , \8288_b0 , \8289_b1 , \8289_b0 , 
		\8290_b1 , \8290_b0 , \8291_b1 , \8291_b0 , \8292_b1 , \8292_b0 , \8293_b1 , \8293_b0 , \8294_b1 , \8294_b0 , 
		\8295_b1 , \8295_b0 , \8296_b1 , \8296_b0 , \8297_b1 , \8297_b0 , \8298_b1 , \8298_b0 , \8299_b1 , \8299_b0 , 
		\8300_b1 , \8300_b0 , \8301_b1 , \8301_b0 , \8302_b1 , \8302_b0 , \8303_b1 , \8303_b0 , \8304_b1 , \8304_b0 , 
		\8305_b1 , \8305_b0 , \8306_b1 , \8306_b0 , \8307_b1 , \8307_b0 , \8308_b1 , \8308_b0 , \8309_b1 , \8309_b0 , 
		\8310_b1 , \8310_b0 , \8311_b1 , \8311_b0 , \8312_b1 , \8312_b0 , \8313_b1 , \8313_b0 , \8314_b1 , \8314_b0 , 
		\8315_b1 , \8315_b0 , \8316_b1 , \8316_b0 , \8317_b1 , \8317_b0 , \8318_b1 , \8318_b0 , \8319_b1 , \8319_b0 , 
		\8320_b1 , \8320_b0 , \8321_b1 , \8321_b0 , \8322_b1 , \8322_b0 , \8323_b1 , \8323_b0 , \8324_b1 , \8324_b0 , 
		\8325_b1 , \8325_b0 , \8326_b1 , \8326_b0 , \8327_b1 , \8327_b0 , \8328_b1 , \8328_b0 , \8329_b1 , \8329_b0 , 
		\8330_b1 , \8330_b0 , \8331_b1 , \8331_b0 , \8332_b1 , \8332_b0 , \8333_b1 , \8333_b0 , \8334_b1 , \8334_b0 , 
		\8335_b1 , \8335_b0 , \8336_b1 , \8336_b0 , \8337_b1 , \8337_b0 , \8338_b1 , \8338_b0 , \8339_b1 , \8339_b0 , 
		\8340_b1 , \8340_b0 , \8341_b1 , \8341_b0 , \8342_b1 , \8342_b0 , \8343_b1 , \8343_b0 , \8344_b1 , \8344_b0 , 
		\8345_b1 , \8345_b0 , \8346_b1 , \8346_b0 , \8347_b1 , \8347_b0 , \8348_b1 , \8348_b0 , \8349_b1 , \8349_b0 , 
		\8350_b1 , \8350_b0 , \8351_b1 , \8351_b0 , \8352_b1 , \8352_b0 , \8353_b1 , \8353_b0 , \8354_b1 , \8354_b0 , 
		\8355_b1 , \8355_b0 , \8356_b1 , \8356_b0 , \8357_b1 , \8357_b0 , \8358_b1 , \8358_b0 , \8359_b1 , \8359_b0 , 
		\8360_b1 , \8360_b0 , \8361_b1 , \8361_b0 , \8362_b1 , \8362_b0 , \8363_b1 , \8363_b0 , \8364_b1 , \8364_b0 , 
		\8365_b1 , \8365_b0 , \8366_b1 , \8366_b0 , \8367_b1 , \8367_b0 , \8368_b1 , \8368_b0 , \8369_b1 , \8369_b0 , 
		\8370_b1 , \8370_b0 , \8371_b1 , \8371_b0 , \8372_b1 , \8372_b0 , \8373_b1 , \8373_b0 , \8374_b1 , \8374_b0 , 
		\8375_b1 , \8375_b0 , \8376_b1 , \8376_b0 , \8377_b1 , \8377_b0 , \8378_b1 , \8378_b0 , \8379_b1 , \8379_b0 , 
		\8380_b1 , \8380_b0 , \8381_b1 , \8381_b0 , \8382_b1 , \8382_b0 , \8383_b1 , \8383_b0 , \8384_b1 , \8384_b0 , 
		\8385_b1 , \8385_b0 , \8386_b1 , \8386_b0 , \8387_b1 , \8387_b0 , \8388_b1 , \8388_b0 , \8389_b1 , \8389_b0 , 
		\8390_b1 , \8390_b0 , \8391_b1 , \8391_b0 , \8392_b1 , \8392_b0 , \8393_b1 , \8393_b0 , \8394_b1 , \8394_b0 , 
		\8395_b1 , \8395_b0 , \8396_b1 , \8396_b0 , \8397_b1 , \8397_b0 , \8398_b1 , \8398_b0 , \8399_b1 , \8399_b0 , 
		\8400_b1 , \8400_b0 , \8401_b1 , \8401_b0 , \8402_b1 , \8402_b0 , \8403_b1 , \8403_b0 , \8404_b1 , \8404_b0 , 
		\8405_b1 , \8405_b0 , \8406_b1 , \8406_b0 , \8407_b1 , \8407_b0 , \8408_b1 , \8408_b0 , \8409_b1 , \8409_b0 , 
		\8410_b1 , \8410_b0 , \8411_b1 , \8411_b0 , \8412_b1 , \8412_b0 , \8413_b1 , \8413_b0 , \8414_b1 , \8414_b0 , 
		\8415_b1 , \8415_b0 , \8416_b1 , \8416_b0 , \8417_b1 , \8417_b0 , \8418_b1 , \8418_b0 , \8419_b1 , \8419_b0 , 
		\8420_b1 , \8420_b0 , \8421_b1 , \8421_b0 , \8422_b1 , \8422_b0 , \8423_b1 , \8423_b0 , \8424_b1 , \8424_b0 , 
		\8425_b1 , \8425_b0 , \8426_b1 , \8426_b0 , \8427_b1 , \8427_b0 , \8428_b1 , \8428_b0 , \8429_b1 , \8429_b0 , 
		\8430_b1 , \8430_b0 , \8431_b1 , \8431_b0 , \8432_b1 , \8432_b0 , \8433_b1 , \8433_b0 , \8434_b1 , \8434_b0 , 
		\8435_b1 , \8435_b0 , \8436_b1 , \8436_b0 , \8437_b1 , \8437_b0 , \8438_b1 , \8438_b0 , \8439_b1 , \8439_b0 , 
		\8440_b1 , \8440_b0 , \8441_b1 , \8441_b0 , \8442_b1 , \8442_b0 , \8443_b1 , \8443_b0 , \8444_b1 , \8444_b0 , 
		\8445_b1 , \8445_b0 , \8446_b1 , \8446_b0 , \8447_b1 , \8447_b0 , \8448_b1 , \8448_b0 , \8449_b1 , \8449_b0 , 
		\8450_b1 , \8450_b0 , \8451_b1 , \8451_b0 , \8452_b1 , \8452_b0 , \8453_b1 , \8453_b0 , \8454_b1 , \8454_b0 , 
		\8455_b1 , \8455_b0 , \8456_b1 , \8456_b0 , \8457_b1 , \8457_b0 , \8458_b1 , \8458_b0 , \8459_b1 , \8459_b0 , 
		\8460_b1 , \8460_b0 , \8461_b1 , \8461_b0 , \8462_b1 , \8462_b0 , \8463_b1 , \8463_b0 , \8464_b1 , \8464_b0 , 
		\8465_b1 , \8465_b0 , \8466_b1 , \8466_b0 , \8467_b1 , \8467_b0 , \8468_b1 , \8468_b0 , \8469_b1 , \8469_b0 , 
		\8470_b1 , \8470_b0 , \8471_b1 , \8471_b0 , \8472_b1 , \8472_b0 , \8473_b1 , \8473_b0 , \8474_b1 , \8474_b0 , 
		\8475_b1 , \8475_b0 , \8476_b1 , \8476_b0 , \8477_b1 , \8477_b0 , \8478_b1 , \8478_b0 , \8479_b1 , \8479_b0 , 
		\8480_b1 , \8480_b0 , \8481_b1 , \8481_b0 , \8482_b1 , \8482_b0 , \8483_b1 , \8483_b0 , \8484_b1 , \8484_b0 , 
		\8485_b1 , \8485_b0 , \8486_b1 , \8486_b0 , \8487_b1 , \8487_b0 , \8488_b1 , \8488_b0 , \8489_b1 , \8489_b0 , 
		\8490_b1 , \8490_b0 , \8491_b1 , \8491_b0 , \8492_b1 , \8492_b0 , \8493_b1 , \8493_b0 , \8494_b1 , \8494_b0 , 
		\8495_b1 , \8495_b0 , \8496_b1 , \8496_b0 , \8497_b1 , \8497_b0 , \8498_b1 , \8498_b0 , \8499_b1 , \8499_b0 , 
		\8500_b1 , \8500_b0 , \8501_b1 , \8501_b0 , \8502_b1 , \8502_b0 , \8503_b1 , \8503_b0 , \8504_b1 , \8504_b0 , 
		\8505_b1 , \8505_b0 , \8506_b1 , \8506_b0 , \8507_b1 , \8507_b0 , \8508_b1 , \8508_b0 , \8509_b1 , \8509_b0 , 
		\8510_b1 , \8510_b0 , \8511_b1 , \8511_b0 , \8512_b1 , \8512_b0 , \8513_b1 , \8513_b0 , \8514_b1 , \8514_b0 , 
		\8515_b1 , \8515_b0 , \8516_b1 , \8516_b0 , \8517_b1 , \8517_b0 , \8518_b1 , \8518_b0 , \8519_b1 , \8519_b0 , 
		\8520_b1 , \8520_b0 , \8521_b1 , \8521_b0 , \8522_b1 , \8522_b0 , \8523_b1 , \8523_b0 , \8524_b1 , \8524_b0 , 
		\8525_b1 , \8525_b0 , \8526_b1 , \8526_b0 , \8527_b1 , \8527_b0 , \8528_b1 , \8528_b0 , \8529_b1 , \8529_b0 , 
		\8530_b1 , \8530_b0 , \8531_b1 , \8531_b0 , \8532_b1 , \8532_b0 , \8533_b1 , \8533_b0 , \8534_b1 , \8534_b0 , 
		\8535_b1 , \8535_b0 , \8536_b1 , \8536_b0 , \8537_b1 , \8537_b0 , \8538_b1 , \8538_b0 , \8539_b1 , \8539_b0 , 
		\8540_b1 , \8540_b0 , \8541_b1 , \8541_b0 , \8542_b1 , \8542_b0 , \8543_b1 , \8543_b0 , \8544_b1 , \8544_b0 , 
		\8545_b1 , \8545_b0 , \8546_b1 , \8546_b0 , \8547_b1 , \8547_b0 , \8548_b1 , \8548_b0 , \8549_b1 , \8549_b0 , 
		\8550_b1 , \8550_b0 , \8551_b1 , \8551_b0 , \8552_b1 , \8552_b0 , \8553_b1 , \8553_b0 , \8554_b1 , \8554_b0 , 
		\8555_b1 , \8555_b0 , \8556_b1 , \8556_b0 , \8557_b1 , \8557_b0 , \8558_b1 , \8558_b0 , \8559_b1 , \8559_b0 , 
		\8560_b1 , \8560_b0 , \8561_b1 , \8561_b0 , \8562_b1 , \8562_b0 , \8563_b1 , \8563_b0 , \8564_b1 , \8564_b0 , 
		\8565_b1 , \8565_b0 , \8566_b1 , \8566_b0 , \8567_b1 , \8567_b0 , \8568_b1 , \8568_b0 , \8569_b1 , \8569_b0 , 
		\8570_b1 , \8570_b0 , \8571_b1 , \8571_b0 , \8572_b1 , \8572_b0 , \8573_b1 , \8573_b0 , \8574_b1 , \8574_b0 , 
		\8575_b1 , \8575_b0 , \8576_b1 , \8576_b0 , \8577_b1 , \8577_b0 , \8578_b1 , \8578_b0 , \8579_b1 , \8579_b0 , 
		\8580_b1 , \8580_b0 , \8581_b1 , \8581_b0 , \8582_b1 , \8582_b0 , \8583_b1 , \8583_b0 , \8584_b1 , \8584_b0 , 
		\8585_b1 , \8585_b0 , \8586_b1 , \8586_b0 , \8587_b1 , \8587_b0 , \8588_b1 , \8588_b0 , \8589_b1 , \8589_b0 , 
		\8590_b1 , \8590_b0 , \8591_b1 , \8591_b0 , \8592_b1 , \8592_b0 , \8593_b1 , \8593_b0 , \8594_b1 , \8594_b0 , 
		\8595_b1 , \8595_b0 , \8596_b1 , \8596_b0 , \8597_b1 , \8597_b0 , \8598_b1 , \8598_b0 , \8599_b1 , \8599_b0 , 
		\8600_b1 , \8600_b0 , \8601_b1 , \8601_b0 , \8602_b1 , \8602_b0 , \8603_b1 , \8603_b0 , \8604_b1 , \8604_b0 , 
		\8605_b1 , \8605_b0 , \8606_b1 , \8606_b0 , \8607_b1 , \8607_b0 , \8608_b1 , \8608_b0 , \8609_b1 , \8609_b0 , 
		\8610_b1 , \8610_b0 , \8611_b1 , \8611_b0 , \8612_b1 , \8612_b0 , \8613_b1 , \8613_b0 , \8614_b1 , \8614_b0 , 
		\8615_b1 , \8615_b0 , \8616_b1 , \8616_b0 , \8617_b1 , \8617_b0 , \8618_b1 , \8618_b0 , \8619_b1 , \8619_b0 , 
		\8620_b1 , \8620_b0 , \8621_b1 , \8621_b0 , \8622_b1 , \8622_b0 , \8623_b1 , \8623_b0 , \8624_b1 , \8624_b0 , 
		\8625_b1 , \8625_b0 , \8626_b1 , \8626_b0 , \8627_b1 , \8627_b0 , \8628_b1 , \8628_b0 , \8629_b1 , \8629_b0 , 
		\8630_b1 , \8630_b0 , \8631_b1 , \8631_b0 , \8632_b1 , \8632_b0 , \8633_b1 , \8633_b0 , \8634_b1 , \8634_b0 , 
		\8635_b1 , \8635_b0 , \8636_b1 , \8636_b0 , \8637_b1 , \8637_b0 , \8638_b1 , \8638_b0 , \8639_b1 , \8639_b0 , 
		\8640_b1 , \8640_b0 , \8641_b1 , \8641_b0 , \8642_b1 , \8642_b0 , \8643_b1 , \8643_b0 , \8644_b1 , \8644_b0 , 
		\8645_b1 , \8645_b0 , \8646_b1 , \8646_b0 , \8647_b1 , \8647_b0 , \8648_b1 , \8648_b0 , \8649_b1 , \8649_b0 , 
		\8650_b1 , \8650_b0 , \8651_b1 , \8651_b0 , \8652_b1 , \8652_b0 , \8653_b1 , \8653_b0 , \8654_b1 , \8654_b0 , 
		\8655_b1 , \8655_b0 , \8656_b1 , \8656_b0 , \8657_b1 , \8657_b0 , \8658_b1 , \8658_b0 , \8659_b1 , \8659_b0 , 
		\8660_b1 , \8660_b0 , \8661_b1 , \8661_b0 , \8662_b1 , \8662_b0 , \8663_b1 , \8663_b0 , \8664_b1 , \8664_b0 , 
		\8665_b1 , \8665_b0 , \8666_b1 , \8666_b0 , \8667_b1 , \8667_b0 , \8668_b1 , \8668_b0 , \8669_b1 , \8669_b0 , 
		\8670_b1 , \8670_b0 , \8671_b1 , \8671_b0 , \8672_b1 , \8672_b0 , \8673_b1 , \8673_b0 , \8674_b1 , \8674_b0 , 
		\8675_b1 , \8675_b0 , \8676_b1 , \8676_b0 , \8677_b1 , \8677_b0 , \8678_b1 , \8678_b0 , \8679_b1 , \8679_b0 , 
		\8680_b1 , \8680_b0 , \8681_b1 , \8681_b0 , \8682_b1 , \8682_b0 , \8683_b1 , \8683_b0 , \8684_b1 , \8684_b0 , 
		\8685_b1 , \8685_b0 , \8686_b1 , \8686_b0 , \8687_b1 , \8687_b0 , \8688_b1 , \8688_b0 , \8689_b1 , \8689_b0 , 
		\8690_b1 , \8690_b0 , \8691_b1 , \8691_b0 , \8692_b1 , \8692_b0 , \8693_b1 , \8693_b0 , \8694_b1 , \8694_b0 , 
		\8695_b1 , \8695_b0 , \8696_b1 , \8696_b0 , \8697_b1 , \8697_b0 , \8698_b1 , \8698_b0 , \8699_b1 , \8699_b0 , 
		\8700_b1 , \8700_b0 , \8701_b1 , \8701_b0 , \8702_b1 , \8702_b0 , \8703_b1 , \8703_b0 , \8704_b1 , \8704_b0 , 
		\8705_b1 , \8705_b0 , \8706_b1 , \8706_b0 , \8707_b1 , \8707_b0 , \8708_b1 , \8708_b0 , \8709_b1 , \8709_b0 , 
		\8710_b1 , \8710_b0 , \8711_b1 , \8711_b0 , \8712_b1 , \8712_b0 , \8713_b1 , \8713_b0 , \8714_b1 , \8714_b0 , 
		\8715_b1 , \8715_b0 , \8716_b1 , \8716_b0 , \8717_b1 , \8717_b0 , \8718_b1 , \8718_b0 , \8719_b1 , \8719_b0 , 
		\8720_b1 , \8720_b0 , \8721_b1 , \8721_b0 , \8722_b1 , \8722_b0 , \8723_b1 , \8723_b0 , \8724_b1 , \8724_b0 , 
		\8725_b1 , \8725_b0 , \8726_b1 , \8726_b0 , \8727_b1 , \8727_b0 , \8728_b1 , \8728_b0 , \8729_b1 , \8729_b0 , 
		\8730_b1 , \8730_b0 , \8731_b1 , \8731_b0 , \8732_b1 , \8732_b0 , \8733_b1 , \8733_b0 , \8734_b1 , \8734_b0 , 
		\8735_b1 , \8735_b0 , \8736_b1 , \8736_b0 , \8737_b1 , \8737_b0 , \8738_b1 , \8738_b0 , \8739_b1 , \8739_b0 , 
		\8740_b1 , \8740_b0 , \8741_b1 , \8741_b0 , \8742_b1 , \8742_b0 , \8743_b1 , \8743_b0 , \8744_b1 , \8744_b0 , 
		\8745_b1 , \8745_b0 , \8746_b1 , \8746_b0 , \8747_b1 , \8747_b0 , \8748_b1 , \8748_b0 , \8749_b1 , \8749_b0 , 
		\8750_b1 , \8750_b0 , \8751_b1 , \8751_b0 , \8752_b1 , \8752_b0 , \8753_b1 , \8753_b0 , \8754_b1 , \8754_b0 , 
		\8755_b1 , \8755_b0 , \8756_b1 , \8756_b0 , \8757_b1 , \8757_b0 , \8758_b1 , \8758_b0 , \8759_b1 , \8759_b0 , 
		\8760_b1 , \8760_b0 , \8761_b1 , \8761_b0 , \8762_b1 , \8762_b0 , \8763_b1 , \8763_b0 , \8764_b1 , \8764_b0 , 
		\8765_b1 , \8765_b0 , \8766_b1 , \8766_b0 , \8767_b1 , \8767_b0 , \8768_b1 , \8768_b0 , \8769_b1 , \8769_b0 , 
		\8770_b1 , \8770_b0 , \8771_b1 , \8771_b0 , \8772_b1 , \8772_b0 , \8773_b1 , \8773_b0 , \8774_b1 , \8774_b0 , 
		\8775_b1 , \8775_b0 , \8776_b1 , \8776_b0 , \8777_b1 , \8777_b0 , \8778_b1 , \8778_b0 , \8779_b1 , \8779_b0 , 
		\8780_b1 , \8780_b0 , \8781_b1 , \8781_b0 , \8782_b1 , \8782_b0 , \8783_b1 , \8783_b0 , \8784_b1 , \8784_b0 , 
		\8785_b1 , \8785_b0 , \8786_b1 , \8786_b0 , \8787_b1 , \8787_b0 , \8788_b1 , \8788_b0 , \8789_b1 , \8789_b0 , 
		\8790_b1 , \8790_b0 , \8791_b1 , \8791_b0 , \8792_b1 , \8792_b0 , \8793_b1 , \8793_b0 , \8794_b1 , \8794_b0 , 
		\8795_b1 , \8795_b0 , \8796_b1 , \8796_b0 , \8797_b1 , \8797_b0 , \8798_b1 , \8798_b0 , \8799_b1 , \8799_b0 , 
		\8800_b1 , \8800_b0 , \8801_b1 , \8801_b0 , \8802_b1 , \8802_b0 , \8803_b1 , \8803_b0 , \8804_b1 , \8804_b0 , 
		\8805_b1 , \8805_b0 , \8806_b1 , \8806_b0 , \8807_b1 , \8807_b0 , \8808_b1 , \8808_b0 , \8809_b1 , \8809_b0 , 
		\8810_b1 , \8810_b0 , \8811_b1 , \8811_b0 , \8812_b1 , \8812_b0 , \8813_b1 , \8813_b0 , \8814_b1 , \8814_b0 , 
		\8815_b1 , \8815_b0 , \8816_b1 , \8816_b0 , \8817_b1 , \8817_b0 , \8818_b1 , \8818_b0 , \8819_b1 , \8819_b0 , 
		\8820_b1 , \8820_b0 , \8821_b1 , \8821_b0 , \8822_b1 , \8822_b0 , \8823_b1 , \8823_b0 , \8824_b1 , \8824_b0 , 
		\8825_b1 , \8825_b0 , \8826_b1 , \8826_b0 , \8827_b1 , \8827_b0 , \8828_b1 , \8828_b0 , \8829_b1 , \8829_b0 , 
		\8830_b1 , \8830_b0 , \8831_b1 , \8831_b0 , \8832_b1 , \8832_b0 , \8833_b1 , \8833_b0 , \8834_b1 , \8834_b0 , 
		\8835_b1 , \8835_b0 , \8836_b1 , \8836_b0 , \8837_b1 , \8837_b0 , \8838_b1 , \8838_b0 , \8839_b1 , \8839_b0 , 
		\8840_b1 , \8840_b0 , \8841_b1 , \8841_b0 , \8842_b1 , \8842_b0 , \8843_b1 , \8843_b0 , \8844_b1 , \8844_b0 , 
		\8845_b1 , \8845_b0 , \8846_b1 , \8846_b0 , \8847_b1 , \8847_b0 , \8848_b1 , \8848_b0 , \8849_b1 , \8849_b0 , 
		\8850_b1 , \8850_b0 , \8851_b1 , \8851_b0 , \8852_b1 , \8852_b0 , \8853_b1 , \8853_b0 , \8854_b1 , \8854_b0 , 
		\8855_b1 , \8855_b0 , \8856_b1 , \8856_b0 , \8857_b1 , \8857_b0 , \8858_b1 , \8858_b0 , \8859_b1 , \8859_b0 , 
		\8860_b1 , \8860_b0 , \8861_b1 , \8861_b0 , \8862_b1 , \8862_b0 , \8863_b1 , \8863_b0 , \8864_b1 , \8864_b0 , 
		\8865_b1 , \8865_b0 , \8866_b1 , \8866_b0 , \8867_b1 , \8867_b0 , \8868_b1 , \8868_b0 , \8869_b1 , \8869_b0 , 
		\8870_b1 , \8870_b0 , \8871_b1 , \8871_b0 , \8872_b1 , \8872_b0 , \8873_b1 , \8873_b0 , \8874_b1 , \8874_b0 , 
		\8875_b1 , \8875_b0 , \8876_b1 , \8876_b0 , \8877_b1 , \8877_b0 , \8878_b1 , \8878_b0 , \8879_b1 , \8879_b0 , 
		\8880_b1 , \8880_b0 , \8881_b1 , \8881_b0 , \8882_b1 , \8882_b0 , \8883_b1 , \8883_b0 , \8884_b1 , \8884_b0 , 
		\8885_b1 , \8885_b0 , \8886_b1 , \8886_b0 , \8887_b1 , \8887_b0 , \8888_b1 , \8888_b0 , \8889_b1 , \8889_b0 , 
		\8890_b1 , \8890_b0 , \8891_b1 , \8891_b0 , \8892_b1 , \8892_b0 , \8893_b1 , \8893_b0 , \8894_b1 , \8894_b0 , 
		\8895_b1 , \8895_b0 , \8896_b1 , \8896_b0 , \8897_b1 , \8897_b0 , \8898_b1 , \8898_b0 , \8899_b1 , \8899_b0 , 
		\8900_b1 , \8900_b0 , \8901_b1 , \8901_b0 , \8902_b1 , \8902_b0 , \8903_b1 , \8903_b0 , \8904_b1 , \8904_b0 , 
		\8905_b1 , \8905_b0 , \8906_b1 , \8906_b0 , \8907_b1 , \8907_b0 , \8908_b1 , \8908_b0 , \8909_b1 , \8909_b0 , 
		\8910_b1 , \8910_b0 , \8911_b1 , \8911_b0 , \8912_b1 , \8912_b0 , \8913_b1 , \8913_b0 , \8914_b1 , \8914_b0 , 
		\8915_b1 , \8915_b0 , \8916_b1 , \8916_b0 , \8917_b1 , \8917_b0 , \8918_b1 , \8918_b0 , \8919_b1 , \8919_b0 , 
		\8920_b1 , \8920_b0 , \8921_b1 , \8921_b0 , \8922_b1 , \8922_b0 , \8923_b1 , \8923_b0 , \8924_b1 , \8924_b0 , 
		\8925_b1 , \8925_b0 , \8926_b1 , \8926_b0 , \8927_b1 , \8927_b0 , \8928_b1 , \8928_b0 , \8929_b1 , \8929_b0 , 
		\8930_b1 , \8930_b0 , \8931_b1 , \8931_b0 , \8932_b1 , \8932_b0 , \8933_b1 , \8933_b0 , \8934_b1 , \8934_b0 , 
		\8935_b1 , \8935_b0 , \8936_b1 , \8936_b0 , \8937_b1 , \8937_b0 , \8938_b1 , \8938_b0 , \8939_b1 , \8939_b0 , 
		\8940_b1 , \8940_b0 , \8941_b1 , \8941_b0 , \8942_b1 , \8942_b0 , \8943_b1 , \8943_b0 , \8944_b1 , \8944_b0 , 
		\8945_b1 , \8945_b0 , \8946_b1 , \8946_b0 , \8947_b1 , \8947_b0 , \8948_b1 , \8948_b0 , \8949_b1 , \8949_b0 , 
		\8950_b1 , \8950_b0 , \8951_b1 , \8951_b0 , \8952_b1 , \8952_b0 , \8953_b1 , \8953_b0 , \8954_b1 , \8954_b0 , 
		\8955_b1 , \8955_b0 , \8956_b1 , \8956_b0 , \8957_b1 , \8957_b0 , \8958_b1 , \8958_b0 , \8959_b1 , \8959_b0 , 
		\8960_b1 , \8960_b0 , \8961_b1 , \8961_b0 , \8962_b1 , \8962_b0 , \8963_b1 , \8963_b0 , \8964_b1 , \8964_b0 , 
		\8965_b1 , \8965_b0 , \8966_b1 , \8966_b0 , \8967_b1 , \8967_b0 , \8968_b1 , \8968_b0 , \8969_b1 , \8969_b0 , 
		\8970_b1 , \8970_b0 , \8971_b1 , \8971_b0 , \8972_b1 , \8972_b0 , \8973_b1 , \8973_b0 , \8974_b1 , \8974_b0 , 
		\8975_b1 , \8975_b0 , \8976_b1 , \8976_b0 , \8977_b1 , \8977_b0 , \8978_b1 , \8978_b0 , \8979_b1 , \8979_b0 , 
		\8980_b1 , \8980_b0 , \8981_b1 , \8981_b0 , \8982_b1 , \8982_b0 , \8983_b1 , \8983_b0 , \8984_b1 , \8984_b0 , 
		\8985_b1 , \8985_b0 , \8986_b1 , \8986_b0 , \8987_b1 , \8987_b0 , \8988_b1 , \8988_b0 , \8989_b1 , \8989_b0 , 
		\8990_b1 , \8990_b0 , \8991_b1 , \8991_b0 , \8992_b1 , \8992_b0 , \8993_b1 , \8993_b0 , \8994_b1 , \8994_b0 , 
		\8995_b1 , \8995_b0 , \8996_b1 , \8996_b0 , \8997_b1 , \8997_b0 , \8998_b1 , \8998_b0 , \8999_b1 , \8999_b0 , 
		\9000_b1 , \9000_b0 , \9001_b1 , \9001_b0 , \9002_b1 , \9002_b0 , \9003_b1 , \9003_b0 , \9004_b1 , \9004_b0 , 
		\9005_b1 , \9005_b0 , \9006_b1 , \9006_b0 , \9007_b1 , \9007_b0 , \9008_b1 , \9008_b0 , \9009_b1 , \9009_b0 , 
		\9010_b1 , \9010_b0 , \9011_b1 , \9011_b0 , \9012_b1 , \9012_b0 , \9013_b1 , \9013_b0 , \9014_b1 , \9014_b0 , 
		\9015_b1 , \9015_b0 , \9016_b1 , \9016_b0 , \9017_b1 , \9017_b0 , \9018_b1 , \9018_b0 , \9019_b1 , \9019_b0 , 
		\9020_b1 , \9020_b0 , \9021_b1 , \9021_b0 , \9022_b1 , \9022_b0 , \9023_b1 , \9023_b0 , \9024_b1 , \9024_b0 , 
		\9025_b1 , \9025_b0 , \9026_b1 , \9026_b0 , \9027_b1 , \9027_b0 , \9028_b1 , \9028_b0 , \9029_b1 , \9029_b0 , 
		\9030_b1 , \9030_b0 , \9031_b1 , \9031_b0 , \9032_b1 , \9032_b0 , \9033_b1 , \9033_b0 , \9034_b1 , \9034_b0 , 
		\9035_b1 , \9035_b0 , \9036_b1 , \9036_b0 , \9037_b1 , \9037_b0 , \9038_b1 , \9038_b0 , \9039_b1 , \9039_b0 , 
		\9040_b1 , \9040_b0 , \9041_b1 , \9041_b0 , \9042_b1 , \9042_b0 , \9043_b1 , \9043_b0 , \9044_b1 , \9044_b0 , 
		\9045_b1 , \9045_b0 , \9046_b1 , \9046_b0 , \9047_b1 , \9047_b0 , \9048_b1 , \9048_b0 , \9049_b1 , \9049_b0 , 
		\9050_b1 , \9050_b0 , \9051_b1 , \9051_b0 , \9052_b1 , \9052_b0 , \9053_b1 , \9053_b0 , \9054_b1 , \9054_b0 , 
		\9055_b1 , \9055_b0 , \9056_b1 , \9056_b0 , \9057_b1 , \9057_b0 , \9058_b1 , \9058_b0 , \9059_b1 , \9059_b0 , 
		\9060_b1 , \9060_b0 , \9061_b1 , \9061_b0 , \9062_b1 , \9062_b0 , \9063_b1 , \9063_b0 , \9064_b1 , \9064_b0 , 
		\9065_b1 , \9065_b0 , \9066_b1 , \9066_b0 , \9067_b1 , \9067_b0 , \9068_b1 , \9068_b0 , \9069_b1 , \9069_b0 , 
		\9070_b1 , \9070_b0 , \9071_b1 , \9071_b0 , \9072_b1 , \9072_b0 , \9073_b1 , \9073_b0 , \9074_b1 , \9074_b0 , 
		\9075_b1 , \9075_b0 , \9076_b1 , \9076_b0 , \9077_b1 , \9077_b0 , \9078_b1 , \9078_b0 , \9079_b1 , \9079_b0 , 
		\9080_b1 , \9080_b0 , \9081_b1 , \9081_b0 , \9082_b1 , \9082_b0 , \9083_b1 , \9083_b0 , \9084_b1 , \9084_b0 , 
		\9085_b1 , \9085_b0 , \9086_b1 , \9086_b0 , \9087_b1 , \9087_b0 , \9088_b1 , \9088_b0 , \9089_b1 , \9089_b0 , 
		\9090_b1 , \9090_b0 , \9091_b1 , \9091_b0 , \9092_b1 , \9092_b0 , \9093_b1 , \9093_b0 , \9094_b1 , \9094_b0 , 
		\9095_b1 , \9095_b0 , \9096_b1 , \9096_b0 , \9097_b1 , \9097_b0 , \9098_b1 , \9098_b0 , \9099_b1 , \9099_b0 , 
		\9100_b1 , \9100_b0 , \9101_b1 , \9101_b0 , \9102_b1 , \9102_b0 , \9103_b1 , \9103_b0 , \9104_b1 , \9104_b0 , 
		\9105_b1 , \9105_b0 , \9106_b1 , \9106_b0 , \9107_b1 , \9107_b0 , \9108_b1 , \9108_b0 , \9109_b1 , \9109_b0 , 
		\9110_b1 , \9110_b0 , \9111_b1 , \9111_b0 , \9112_b1 , \9112_b0 , \9113_b1 , \9113_b0 , \9114_b1 , \9114_b0 , 
		\9115_b1 , \9115_b0 , \9116_b1 , \9116_b0 , \9117_b1 , \9117_b0 , \9118_b1 , \9118_b0 , \9119_b1 , \9119_b0 , 
		\9120_b1 , \9120_b0 , \9121_b1 , \9121_b0 , \9122_b1 , \9122_b0 , \9123_b1 , \9123_b0 , \9124_b1 , \9124_b0 , 
		\9125_b1 , \9125_b0 , \9126_b1 , \9126_b0 , \9127_b1 , \9127_b0 , \9128_b1 , \9128_b0 , \9129_b1 , \9129_b0 , 
		\9130_b1 , \9130_b0 , \9131_b1 , \9131_b0 , \9132_b1 , \9132_b0 , \9133_b1 , \9133_b0 , \9134_b1 , \9134_b0 , 
		\9135_b1 , \9135_b0 , \9136_b1 , \9136_b0 , \9137_b1 , \9137_b0 , \9138_b1 , \9138_b0 , \9139_b1 , \9139_b0 , 
		\9140_b1 , \9140_b0 , \9141_b1 , \9141_b0 , \9142_b1 , \9142_b0 , \9143_b1 , \9143_b0 , \9144_b1 , \9144_b0 , 
		\9145_b1 , \9145_b0 , \9146_b1 , \9146_b0 , \9147_b1 , \9147_b0 , \9148_b1 , \9148_b0 , \9149_b1 , \9149_b0 , 
		\9150_b1 , \9150_b0 , \9151_b1 , \9151_b0 , \9152_b1 , \9152_b0 , \9153_b1 , \9153_b0 , \9154_b1 , \9154_b0 , 
		\9155_b1 , \9155_b0 , \9156_b1 , \9156_b0 , \9157_b1 , \9157_b0 , \9158_b1 , \9158_b0 , \9159_b1 , \9159_b0 , 
		\9160_b1 , \9160_b0 , \9161_b1 , \9161_b0 , \9162_b1 , \9162_b0 , \9163_b1 , \9163_b0 , \9164_b1 , \9164_b0 , 
		\9165_b1 , \9165_b0 , \9166_b1 , \9166_b0 , \9167_b1 , \9167_b0 , \9168_b1 , \9168_b0 , \9169_b1 , \9169_b0 , 
		\9170_b1 , \9170_b0 , \9171_b1 , \9171_b0 , \9172_b1 , \9172_b0 , \9173_b1 , \9173_b0 , \9174_b1 , \9174_b0 , 
		\9175_b1 , \9175_b0 , \9176_b1 , \9176_b0 , \9177_b1 , \9177_b0 , \9178_b1 , \9178_b0 , \9179_b1 , \9179_b0 , 
		\9180_b1 , \9180_b0 , \9181_b1 , \9181_b0 , \9182_b1 , \9182_b0 , \9183_b1 , \9183_b0 , \9184_b1 , \9184_b0 , 
		\9185_b1 , \9185_b0 , \9186_b1 , \9186_b0 , \9187_b1 , \9187_b0 , \9188_b1 , \9188_b0 , \9189_b1 , \9189_b0 , 
		\9190_b1 , \9190_b0 , \9191_b1 , \9191_b0 , \9192_b1 , \9192_b0 , \9193_b1 , \9193_b0 , \9194_b1 , \9194_b0 , 
		\9195_b1 , \9195_b0 , \9196_b1 , \9196_b0 , \9197_b1 , \9197_b0 , \9198_b1 , \9198_b0 , \9199_b1 , \9199_b0 , 
		\9200_b1 , \9200_b0 , \9201_b1 , \9201_b0 , \9202_b1 , \9202_b0 , \9203_b1 , \9203_b0 , \9204_b1 , \9204_b0 , 
		\9205_b1 , \9205_b0 , \9206_b1 , \9206_b0 , \9207_b1 , \9207_b0 , \9208_b1 , \9208_b0 , \9209_b1 , \9209_b0 , 
		\9210_b1 , \9210_b0 , \9211_b1 , \9211_b0 , \9212_b1 , \9212_b0 , \9213_b1 , \9213_b0 , \9214_b1 , \9214_b0 , 
		\9215_b1 , \9215_b0 , \9216_b1 , \9216_b0 , \9217_b1 , \9217_b0 , \9218_b1 , \9218_b0 , \9219_b1 , \9219_b0 , 
		\9220_b1 , \9220_b0 , \9221_b1 , \9221_b0 , \9222_b1 , \9222_b0 , \9223_b1 , \9223_b0 , \9224_b1 , \9224_b0 , 
		\9225_b1 , \9225_b0 , \9226_b1 , \9226_b0 , \9227_b1 , \9227_b0 , \9228_b1 , \9228_b0 , \9229_b1 , \9229_b0 , 
		\9230_b1 , \9230_b0 , \9231_b1 , \9231_b0 , \9232_b1 , \9232_b0 , \9233_b1 , \9233_b0 , \9234_b1 , \9234_b0 , 
		\9235_b1 , \9235_b0 , \9236_b1 , \9236_b0 , \9237_b1 , \9237_b0 , \9238_b1 , \9238_b0 , \9239_b1 , \9239_b0 , 
		\9240_b1 , \9240_b0 , \9241_b1 , \9241_b0 , \9242_b1 , \9242_b0 , \9243_b1 , \9243_b0 , \9244_b1 , \9244_b0 , 
		\9245_b1 , \9245_b0 , \9246_b1 , \9246_b0 , \9247_b1 , \9247_b0 , \9248_b1 , \9248_b0 , \9249_b1 , \9249_b0 , 
		\9250_b1 , \9250_b0 , \9251_b1 , \9251_b0 , \9252_b1 , \9252_b0 , \9253_b1 , \9253_b0 , \9254_b1 , \9254_b0 , 
		\9255_b1 , \9255_b0 , \9256_b1 , \9256_b0 , \9257_b1 , \9257_b0 , \9258_b1 , \9258_b0 , \9259_b1 , \9259_b0 , 
		\9260_b1 , \9260_b0 , \9261_b1 , \9261_b0 , \9262_b1 , \9262_b0 , \9263_b1 , \9263_b0 , \9264_b1 , \9264_b0 , 
		\9265_b1 , \9265_b0 , \9266_b1 , \9266_b0 , \9267_b1 , \9267_b0 , \9268_b1 , \9268_b0 , \9269_b1 , \9269_b0 , 
		\9270_b1 , \9270_b0 , \9271_b1 , \9271_b0 , \9272_b1 , \9272_b0 , \9273_b1 , \9273_b0 , \9274_b1 , \9274_b0 , 
		\9275_b1 , \9275_b0 , \9276_b1 , \9276_b0 , \9277_b1 , \9277_b0 , \9278_b1 , \9278_b0 , \9279_b1 , \9279_b0 , 
		\9280_b1 , \9280_b0 , \9281_b1 , \9281_b0 , \9282_b1 , \9282_b0 , \9283_b1 , \9283_b0 , \9284_b1 , \9284_b0 , 
		\9285_b1 , \9285_b0 , \9286_b1 , \9286_b0 , \9287_b1 , \9287_b0 , \9288_b1 , \9288_b0 , \9289_b1 , \9289_b0 , 
		\9290_b1 , \9290_b0 , \9291_b1 , \9291_b0 , \9292_b1 , \9292_b0 , \9293_b1 , \9293_b0 , \9294_b1 , \9294_b0 , 
		\9295_b1 , \9295_b0 , \9296_b1 , \9296_b0 , \9297_b1 , \9297_b0 , \9298_b1 , \9298_b0 , \9299_b1 , \9299_b0 , 
		\9300_b1 , \9300_b0 , \9301_b1 , \9301_b0 , \9302_b1 , \9302_b0 , \9303_b1 , \9303_b0 , \9304_b1 , \9304_b0 , 
		\9305_b1 , \9305_b0 , \9306_b1 , \9306_b0 , \9307_b1 , \9307_b0 , \9308_b1 , \9308_b0 , \9309_b1 , \9309_b0 , 
		\9310_b1 , \9310_b0 , \9311_b1 , \9311_b0 , \9312_b1 , \9312_b0 , \9313_b1 , \9313_b0 , \9314_b1 , \9314_b0 , 
		\9315_b1 , \9315_b0 , \9316_b1 , \9316_b0 , \9317_b1 , \9317_b0 , \9318_b1 , \9318_b0 , \9319_b1 , \9319_b0 , 
		\9320_b1 , \9320_b0 , \9321_b1 , \9321_b0 , \9322_b1 , \9322_b0 , \9323_b1 , \9323_b0 , \9324_b1 , \9324_b0 , 
		\9325_b1 , \9325_b0 , \9326_b1 , \9326_b0 , \9327_b1 , \9327_b0 , \9328_b1 , \9328_b0 , \9329_b1 , \9329_b0 , 
		\9330_b1 , \9330_b0 , \9331_b1 , \9331_b0 , \9332_b1 , \9332_b0 , \9333_b1 , \9333_b0 , \9334_b1 , \9334_b0 , 
		\9335_b1 , \9335_b0 , \9336_b1 , \9336_b0 , \9337_b1 , \9337_b0 , \9338_b1 , \9338_b0 , \9339_b1 , \9339_b0 , 
		\9340_b1 , \9340_b0 , \9341_b1 , \9341_b0 , \9342_b1 , \9342_b0 , \9343_b1 , \9343_b0 , \9344_b1 , \9344_b0 , 
		\9345_b1 , \9345_b0 , \9346_b1 , \9346_b0 , \9347_b1 , \9347_b0 , \9348_b1 , \9348_b0 , \9349_b1 , \9349_b0 , 
		\9350_b1 , \9350_b0 , \9351_b1 , \9351_b0 , \9352_b1 , \9352_b0 , \9353_b1 , \9353_b0 , \9354_b1 , \9354_b0 , 
		\9355_b1 , \9355_b0 , \9356_b1 , \9356_b0 , \9357_b1 , \9357_b0 , \9358_b1 , \9358_b0 , \9359_b1 , \9359_b0 , 
		\9360_b1 , \9360_b0 , \9361_b1 , \9361_b0 , \9362_b1 , \9362_b0 , \9363_b1 , \9363_b0 , \9364_b1 , \9364_b0 , 
		\9365_b1 , \9365_b0 , \9366_b1 , \9366_b0 , \9367_b1 , \9367_b0 , \9368_b1 , \9368_b0 , \9369_b1 , \9369_b0 , 
		\9370_b1 , \9370_b0 , \9371_b1 , \9371_b0 , \9372_b1 , \9372_b0 , \9373_b1 , \9373_b0 , \9374_b1 , \9374_b0 , 
		\9375_b1 , \9375_b0 , \9376_b1 , \9376_b0 , \9377_b1 , \9377_b0 , \9378_b1 , \9378_b0 , \9379_b1 , \9379_b0 , 
		\9380_b1 , \9380_b0 , \9381_b1 , \9381_b0 , \9382_b1 , \9382_b0 , \9383_b1 , \9383_b0 , \9384_b1 , \9384_b0 , 
		\9385_b1 , \9385_b0 , \9386_b1 , \9386_b0 , \9387_b1 , \9387_b0 , \9388_b1 , \9388_b0 , \9389_b1 , \9389_b0 , 
		\9390_b1 , \9390_b0 , \9391_b1 , \9391_b0 , \9392_b1 , \9392_b0 , \9393_b1 , \9393_b0 , \9394_b1 , \9394_b0 , 
		\9395_b1 , \9395_b0 , \9396_b1 , \9396_b0 , \9397_b1 , \9397_b0 , \9398_b1 , \9398_b0 , \9399_b1 , \9399_b0 , 
		\9400_b1 , \9400_b0 , \9401_b1 , \9401_b0 , \9402_b1 , \9402_b0 , \9403_b1 , \9403_b0 , \9404_b1 , \9404_b0 , 
		\9405_b1 , \9405_b0 , \9406_b1 , \9406_b0 , \9407_b1 , \9407_b0 , \9408_b1 , \9408_b0 , \9409_b1 , \9409_b0 , 
		\9410_b1 , \9410_b0 , \9411_b1 , \9411_b0 , \9412_b1 , \9412_b0 , \9413_b1 , \9413_b0 , \9414_b1 , \9414_b0 , 
		\9415_b1 , \9415_b0 , \9416_b1 , \9416_b0 , \9417_b1 , \9417_b0 , \9418_b1 , \9418_b0 , \9419_b1 , \9419_b0 , 
		\9420_b1 , \9420_b0 , \9421_b1 , \9421_b0 , \9422_b1 , \9422_b0 , \9423_b1 , \9423_b0 , \9424_b1 , \9424_b0 , 
		\9425_b1 , \9425_b0 , \9426_b1 , \9426_b0 , \9427_b1 , \9427_b0 , \9428_b1 , \9428_b0 , \9429_b1 , \9429_b0 , 
		\9430_b1 , \9430_b0 , \9431_b1 , \9431_b0 , \9432_b1 , \9432_b0 , \9433_b1 , \9433_b0 , \9434_b1 , \9434_b0 , 
		\9435_b1 , \9435_b0 , \9436_b1 , \9436_b0 , \9437_b1 , \9437_b0 , \9438_b1 , \9438_b0 , \9439_b1 , \9439_b0 , 
		\9440_b1 , \9440_b0 , \9441_b1 , \9441_b0 , \9442_b1 , \9442_b0 , \9443_b1 , \9443_b0 , \9444_b1 , \9444_b0 , 
		\9445_b1 , \9445_b0 , \9446_b1 , \9446_b0 , \9447_b1 , \9447_b0 , \9448_b1 , \9448_b0 , \9449_b1 , \9449_b0 , 
		\9450_b1 , \9450_b0 , \9451_b1 , \9451_b0 , \9452_b1 , \9452_b0 , \9453_b1 , \9453_b0 , \9454_b1 , \9454_b0 , 
		\9455_b1 , \9455_b0 , \9456_b1 , \9456_b0 , \9457_b1 , \9457_b0 , \9458_b1 , \9458_b0 , \9459_b1 , \9459_b0 , 
		\9460_b1 , \9460_b0 , \9461_b1 , \9461_b0 , \9462_b1 , \9462_b0 , \9463_b1 , \9463_b0 , \9464_b1 , \9464_b0 , 
		\9465_b1 , \9465_b0 , \9466_b1 , \9466_b0 , \9467_b1 , \9467_b0 , \9468_b1 , \9468_b0 , \9469_b1 , \9469_b0 , 
		\9470_b1 , \9470_b0 , \9471_b1 , \9471_b0 , \9472_b1 , \9472_b0 , \9473_b1 , \9473_b0 , \9474_b1 , \9474_b0 , 
		\9475_b1 , \9475_b0 , \9476_b1 , \9476_b0 , \9477_b1 , \9477_b0 , \9478_b1 , \9478_b0 , \9479_b1 , \9479_b0 , 
		\9480_b1 , \9480_b0 , \9481_b1 , \9481_b0 , \9482_b1 , \9482_b0 , \9483_b1 , \9483_b0 , \9484_b1 , \9484_b0 , 
		\9485_b1 , \9485_b0 , \9486_b1 , \9486_b0 , \9487_b1 , \9487_b0 , \9488_b1 , \9488_b0 , \9489_b1 , \9489_b0 , 
		\9490_b1 , \9490_b0 , \9491_b1 , \9491_b0 , \9492_b1 , \9492_b0 , \9493_b1 , \9493_b0 , \9494_b1 , \9494_b0 , 
		\9495_b1 , \9495_b0 , \9496_b1 , \9496_b0 , \9497_b1 , \9497_b0 , \9498_b1 , \9498_b0 , \9499_b1 , \9499_b0 , 
		\9500_b1 , \9500_b0 , \9501_b1 , \9501_b0 , \9502_b1 , \9502_b0 , \9503_b1 , \9503_b0 , \9504_b1 , \9504_b0 , 
		\9505_b1 , \9505_b0 , \9506_b1 , \9506_b0 , \9507_b1 , \9507_b0 , \9508_b1 , \9508_b0 , \9509_b1 , \9509_b0 , 
		\9510_b1 , \9510_b0 , \9511_b1 , \9511_b0 , \9512_b1 , \9512_b0 , \9513_b1 , \9513_b0 , \9514_b1 , \9514_b0 , 
		\9515_b1 , \9515_b0 , \9516_b1 , \9516_b0 , \9517_b1 , \9517_b0 , \9518_b1 , \9518_b0 , \9519_b1 , \9519_b0 , 
		\9520_b1 , \9520_b0 , \9521_b1 , \9521_b0 , \9522_b1 , \9522_b0 , \9523_b1 , \9523_b0 , \9524_b1 , \9524_b0 , 
		\9525_b1 , \9525_b0 , \9526_b1 , \9526_b0 , \9527_b1 , \9527_b0 , \9528_b1 , \9528_b0 , \9529_b1 , \9529_b0 , 
		\9530_b1 , \9530_b0 , \9531_b1 , \9531_b0 , \9532_b1 , \9532_b0 , \9533_b1 , \9533_b0 , \9534_b1 , \9534_b0 , 
		\9535_b1 , \9535_b0 , \9536_b1 , \9536_b0 , \9537_b1 , \9537_b0 , \9538_b1 , \9538_b0 , \9539_b1 , \9539_b0 , 
		\9540_b1 , \9540_b0 , \9541_b1 , \9541_b0 , \9542_b1 , \9542_b0 , \9543_b1 , \9543_b0 , \9544_b1 , \9544_b0 , 
		\9545_b1 , \9545_b0 , \9546_b1 , \9546_b0 , \9547_b1 , \9547_b0 , \9548_b1 , \9548_b0 , \9549_b1 , \9549_b0 , 
		\9550_b1 , \9550_b0 , \9551_b1 , \9551_b0 , \9552_b1 , \9552_b0 , \9553_b1 , \9553_b0 , \9554_b1 , \9554_b0 , 
		\9555_b1 , \9555_b0 , \9556_b1 , \9556_b0 , \9557_b1 , \9557_b0 , \9558_b1 , \9558_b0 , \9559_b1 , \9559_b0 , 
		\9560_b1 , \9560_b0 , \9561_b1 , \9561_b0 , \9562_b1 , \9562_b0 , \9563_b1 , \9563_b0 , \9564_b1 , \9564_b0 , 
		\9565_b1 , \9565_b0 , \9566_b1 , \9566_b0 , \9567_b1 , \9567_b0 , \9568_b1 , \9568_b0 , \9569_b1 , \9569_b0 , 
		\9570_b1 , \9570_b0 , \9571_b1 , \9571_b0 , \9572_b1 , \9572_b0 , \9573_b1 , \9573_b0 , \9574_b1 , \9574_b0 , 
		\9575_b1 , \9575_b0 , \9576_b1 , \9576_b0 , \9577_b1 , \9577_b0 , \9578_b1 , \9578_b0 , \9579_b1 , \9579_b0 , 
		\9580_b1 , \9580_b0 , \9581_b1 , \9581_b0 , \9582_b1 , \9582_b0 , \9583_b1 , \9583_b0 , \9584_b1 , \9584_b0 , 
		\9585_b1 , \9585_b0 , \9586_b1 , \9586_b0 , \9587_b1 , \9587_b0 , \9588_b1 , \9588_b0 , \9589_b1 , \9589_b0 , 
		\9590_b1 , \9590_b0 , \9591_b1 , \9591_b0 , \9592_b1 , \9592_b0 , \9593_b1 , \9593_b0 , \9594_b1 , \9594_b0 , 
		\9595_b1 , \9595_b0 , \9596_b1 , \9596_b0 , \9597_b1 , \9597_b0 , \9598_b1 , \9598_b0 , \9599_b1 , \9599_b0 , 
		\9600_b1 , \9600_b0 , \9601_b1 , \9601_b0 , \9602_b1 , \9602_b0 , \9603_b1 , \9603_b0 , \9604_b1 , \9604_b0 , 
		\9605_b1 , \9605_b0 , \9606_b1 , \9606_b0 , \9607_b1 , \9607_b0 , \9608_b1 , \9608_b0 , \9609_b1 , \9609_b0 , 
		\9610_b1 , \9610_b0 , \9611_b1 , \9611_b0 , \9612_b1 , \9612_b0 , \9613_b1 , \9613_b0 , \9614_b1 , \9614_b0 , 
		\9615_b1 , \9615_b0 , \9616_b1 , \9616_b0 , \9617_b1 , \9617_b0 , \9618_b1 , \9618_b0 , \9619_b1 , \9619_b0 , 
		\9620_b1 , \9620_b0 , \9621_b1 , \9621_b0 , \9622_b1 , \9622_b0 , \9623_b1 , \9623_b0 , \9624_b1 , \9624_b0 , 
		\9625_b1 , \9625_b0 , \9626_b1 , \9626_b0 , \9627_b1 , \9627_b0 , \9628_b1 , \9628_b0 , \9629_b1 , \9629_b0 , 
		\9630_b1 , \9630_b0 , \9631_b1 , \9631_b0 , \9632_b1 , \9632_b0 , \9633_b1 , \9633_b0 , \9634_b1 , \9634_b0 , 
		\9635_b1 , \9635_b0 , \9636_b1 , \9636_b0 , \9637_b1 , \9637_b0 , \9638_b1 , \9638_b0 , \9639_b1 , \9639_b0 , 
		\9640_b1 , \9640_b0 , \9641_b1 , \9641_b0 , \9642_b1 , \9642_b0 , \9643_b1 , \9643_b0 , \9644_b1 , \9644_b0 , 
		\9645_b1 , \9645_b0 , \9646_b1 , \9646_b0 , \9647_b1 , \9647_b0 , \9648_b1 , \9648_b0 , \9649_b1 , \9649_b0 , 
		\9650_b1 , \9650_b0 , \9651_b1 , \9651_b0 , \9652_b1 , \9652_b0 , \9653_b1 , \9653_b0 , \9654_b1 , \9654_b0 , 
		\9655_b1 , \9655_b0 , \9656_b1 , \9656_b0 , \9657_b1 , \9657_b0 , \9658_b1 , \9658_b0 , \9659_b1 , \9659_b0 , 
		\9660_b1 , \9660_b0 , \9661_b1 , \9661_b0 , \9662_b1 , \9662_b0 , \9663_b1 , \9663_b0 , \9664_b1 , \9664_b0 , 
		\9665_b1 , \9665_b0 , \9666_b1 , \9666_b0 , \9667_b1 , \9667_b0 , \9668_b1 , \9668_b0 , \9669_b1 , \9669_b0 , 
		\9670_b1 , \9670_b0 , \9671_b1 , \9671_b0 , \9672_b1 , \9672_b0 , \9673_b1 , \9673_b0 , \9674_b1 , \9674_b0 , 
		\9675_b1 , \9675_b0 , \9676_b1 , \9676_b0 , \9677_b1 , \9677_b0 , \9678_b1 , \9678_b0 , \9679_b1 , \9679_b0 , 
		\9680_b1 , \9680_b0 , \9681_b1 , \9681_b0 , \9682_b1 , \9682_b0 , \9683_b1 , \9683_b0 , \9684_b1 , \9684_b0 , 
		\9685_b1 , \9685_b0 , \9686_b1 , \9686_b0 , \9687_b1 , \9687_b0 , \9688_b1 , \9688_b0 , \9689_b1 , \9689_b0 , 
		\9690_b1 , \9690_b0 , \9691_b1 , \9691_b0 , \9692_b1 , \9692_b0 , \9693_b1 , \9693_b0 , \9694_b1 , \9694_b0 , 
		\9695_b1 , \9695_b0 , \9696_b1 , \9696_b0 , \9697_b1 , \9697_b0 , \9698_b1 , \9698_b0 , \9699_b1 , \9699_b0 , 
		\9700_b1 , \9700_b0 , \9701_b1 , \9701_b0 , \9702_b1 , \9702_b0 , \9703_b1 , \9703_b0 , \9704_b1 , \9704_b0 , 
		\9705_b1 , \9705_b0 , \9706_b1 , \9706_b0 , \9707_b1 , \9707_b0 , \9708_b1 , \9708_b0 , \9709_b1 , \9709_b0 , 
		\9710_b1 , \9710_b0 , \9711_b1 , \9711_b0 , \9712_b1 , \9712_b0 , \9713_b1 , \9713_b0 , \9714_b1 , \9714_b0 , 
		\9715_b1 , \9715_b0 , \9716_b1 , \9716_b0 , \9717_b1 , \9717_b0 , \9718_b1 , \9718_b0 , \9719_b1 , \9719_b0 , 
		\9720_b1 , \9720_b0 , \9721_b1 , \9721_b0 , \9722_b1 , \9722_b0 , \9723_b1 , \9723_b0 , \9724_b1 , \9724_b0 , 
		\9725_b1 , \9725_b0 , \9726_b1 , \9726_b0 , \9727_b1 , \9727_b0 , \9728_b1 , \9728_b0 , \9729_b1 , \9729_b0 , 
		\9730_b1 , \9730_b0 , \9731_b1 , \9731_b0 , \9732_b1 , \9732_b0 , \9733_b1 , \9733_b0 , \9734_b1 , \9734_b0 , 
		\9735_b1 , \9735_b0 , \9736_b1 , \9736_b0 , \9737_b1 , \9737_b0 , \9738_b1 , \9738_b0 , \9739_b1 , \9739_b0 , 
		\9740_b1 , \9740_b0 , \9741_b1 , \9741_b0 , \9742_b1 , \9742_b0 , \9743_b1 , \9743_b0 , \9744_b1 , \9744_b0 , 
		\9745_b1 , \9745_b0 , \9746_b1 , \9746_b0 , \9747_b1 , \9747_b0 , \9748_b1 , \9748_b0 , \9749_b1 , \9749_b0 , 
		\9750_b1 , \9750_b0 , \9751_b1 , \9751_b0 , \9752_b1 , \9752_b0 , \9753_b1 , \9753_b0 , \9754_b1 , \9754_b0 , 
		\9755_b1 , \9755_b0 , \9756_b1 , \9756_b0 , \9757_b1 , \9757_b0 , \9758_b1 , \9758_b0 , \9759_b1 , \9759_b0 , 
		\9760_b1 , \9760_b0 , \9761_b1 , \9761_b0 , \9762_b1 , \9762_b0 , \9763_b1 , \9763_b0 , \9764_b1 , \9764_b0 , 
		\9765_b1 , \9765_b0 , \9766_b1 , \9766_b0 , \9767_b1 , \9767_b0 , \9768_b1 , \9768_b0 , \9769_b1 , \9769_b0 , 
		\9770_b1 , \9770_b0 , \9771_b1 , \9771_b0 , \9772_b1 , \9772_b0 , \9773_b1 , \9773_b0 , \9774_b1 , \9774_b0 , 
		\9775_b1 , \9775_b0 , \9776_b1 , \9776_b0 , \9777_b1 , \9777_b0 , \9778_b1 , \9778_b0 , \9779_b1 , \9779_b0 , 
		\9780_b1 , \9780_b0 , \9781_b1 , \9781_b0 , \9782_b1 , \9782_b0 , \9783_b1 , \9783_b0 , \9784_b1 , \9784_b0 , 
		\9785_b1 , \9785_b0 , \9786_b1 , \9786_b0 , \9787_b1 , \9787_b0 , \9788_b1 , \9788_b0 , \9789_b1 , \9789_b0 , 
		\9790_b1 , \9790_b0 , \9791_b1 , \9791_b0 , \9792_b1 , \9792_b0 , \9793_b1 , \9793_b0 , \9794_b1 , \9794_b0 , 
		\9795_b1 , \9795_b0 , \9796_b1 , \9796_b0 , \9797_b1 , \9797_b0 , \9798_b1 , \9798_b0 , \9799_b1 , \9799_b0 , 
		\9800_b1 , \9800_b0 , \9801_b1 , \9801_b0 , \9802_b1 , \9802_b0 , \9803_b1 , \9803_b0 , \9804_b1 , \9804_b0 , 
		\9805_b1 , \9805_b0 , \9806_b1 , \9806_b0 , \9807_b1 , \9807_b0 , \9808_b1 , \9808_b0 , \9809_b1 , \9809_b0 , 
		\9810_b1 , \9810_b0 , \9811_b1 , \9811_b0 , \9812_b1 , \9812_b0 , \9813_b1 , \9813_b0 , \9814_b1 , \9814_b0 , 
		\9815_b1 , \9815_b0 , \9816_b1 , \9816_b0 , \9817_b1 , \9817_b0 , \9818_b1 , \9818_b0 , \9819_b1 , \9819_b0 , 
		\9820_b1 , \9820_b0 , \9821_b1 , \9821_b0 , \9822_b1 , \9822_b0 , \9823_b1 , \9823_b0 , \9824_b1 , \9824_b0 , 
		\9825_b1 , \9825_b0 , \9826_b1 , \9826_b0 , \9827_b1 , \9827_b0 , \9828_b1 , \9828_b0 , \9829_b1 , \9829_b0 , 
		\9830_b1 , \9830_b0 , \9831_b1 , \9831_b0 , \9832_b1 , \9832_b0 , \9833_b1 , \9833_b0 , \9834_b1 , \9834_b0 , 
		\9835_b1 , \9835_b0 , \9836_b1 , \9836_b0 , \9837_b1 , \9837_b0 , \9838_b1 , \9838_b0 , \9839_b1 , \9839_b0 , 
		\9840_b1 , \9840_b0 , \9841_b1 , \9841_b0 , \9842_b1 , \9842_b0 , \9843_b1 , \9843_b0 , \9844_b1 , \9844_b0 , 
		\9845_b1 , \9845_b0 , \9846_b1 , \9846_b0 , \9847_b1 , \9847_b0 , \9848_b1 , \9848_b0 , \9849_b1 , \9849_b0 , 
		\9850_b1 , \9850_b0 , \9851_b1 , \9851_b0 , \9852_b1 , \9852_b0 , \9853_b1 , \9853_b0 , \9854_b1 , \9854_b0 , 
		\9855_b1 , \9855_b0 , \9856_b1 , \9856_b0 , \9857_b1 , \9857_b0 , \9858_b1 , \9858_b0 , \9859_b1 , \9859_b0 , 
		\9860_b1 , \9860_b0 , \9861_b1 , \9861_b0 , \9862_b1 , \9862_b0 , \9863_b1 , \9863_b0 , \9864_b1 , \9864_b0 , 
		\9865_b1 , \9865_b0 , \9866_b1 , \9866_b0 , \9867_b1 , \9867_b0 , \9868_b1 , \9868_b0 , \9869_b1 , \9869_b0 , 
		\9870_b1 , \9870_b0 , \9871_b1 , \9871_b0 , \9872_b1 , \9872_b0 , \9873_b1 , \9873_b0 , \9874_b1 , \9874_b0 , 
		\9875_b1 , \9875_b0 , \9876_b1 , \9876_b0 , \9877_b1 , \9877_b0 , \9878_b1 , \9878_b0 , \9879_b1 , \9879_b0 , 
		\9880_b1 , \9880_b0 , \9881_b1 , \9881_b0 , \9882_b1 , \9882_b0 , \9883_b1 , \9883_b0 , \9884_b1 , \9884_b0 , 
		\9885_b1 , \9885_b0 , \9886_b1 , \9886_b0 , \9887_b1 , \9887_b0 , \9888_b1 , \9888_b0 , \9889_b1 , \9889_b0 , 
		\9890_b1 , \9890_b0 , \9891_b1 , \9891_b0 , \9892_b1 , \9892_b0 , \9893_b1 , \9893_b0 , \9894_b1 , \9894_b0 , 
		\9895_b1 , \9895_b0 , \9896_b1 , \9896_b0 , \9897_b1 , \9897_b0 , \9898_b1 , \9898_b0 , \9899_b1 , \9899_b0 , 
		\9900_b1 , \9900_b0 , \9901_b1 , \9901_b0 , \9902_b1 , \9902_b0 , \9903_b1 , \9903_b0 , \9904_b1 , \9904_b0 , 
		\9905_b1 , \9905_b0 , \9906_b1 , \9906_b0 , \9907_b1 , \9907_b0 , \9908_b1 , \9908_b0 , \9909_b1 , \9909_b0 , 
		\9910_b1 , \9910_b0 , \9911_b1 , \9911_b0 , \9912_b1 , \9912_b0 , \9913_b1 , \9913_b0 , \9914_b1 , \9914_b0 , 
		\9915_b1 , \9915_b0 , \9916_b1 , \9916_b0 , \9917_b1 , \9917_b0 , \9918_b1 , \9918_b0 , \9919_b1 , \9919_b0 , 
		\9920_b1 , \9920_b0 , \9921_b1 , \9921_b0 , \9922_b1 , \9922_b0 , \9923_b1 , \9923_b0 , \9924_b1 , \9924_b0 , 
		\9925_b1 , \9925_b0 , \9926_b1 , \9926_b0 , \9927_b1 , \9927_b0 , \9928_b1 , \9928_b0 , \9929_b1 , \9929_b0 , 
		\9930_b1 , \9930_b0 , \9931_b1 , \9931_b0 , \9932_b1 , \9932_b0 , \9933_b1 , \9933_b0 , \9934_b1 , \9934_b0 , 
		\9935_b1 , \9935_b0 , \9936_b1 , \9936_b0 , \9937_b1 , \9937_b0 , \9938_b1 , \9938_b0 , \9939_b1 , \9939_b0 , 
		\9940_b1 , \9940_b0 , \9941_b1 , \9941_b0 , \9942_b1 , \9942_b0 , \9943_b1 , \9943_b0 , \9944_b1 , \9944_b0 , 
		\9945_b1 , \9945_b0 , \9946_b1 , \9946_b0 , \9947_b1 , \9947_b0 , \9948_b1 , \9948_b0 , \9949_b1 , \9949_b0 , 
		\9950_b1 , \9950_b0 , \9951_b1 , \9951_b0 , \9952_b1 , \9952_b0 , \9953_b1 , \9953_b0 , \9954_b1 , \9954_b0 , 
		\9955_b1 , \9955_b0 , \9956_b1 , \9956_b0 , \9957_b1 , \9957_b0 , \9958_b1 , \9958_b0 , \9959_b1 , \9959_b0 , 
		\9960_b1 , \9960_b0 , \9961_b1 , \9961_b0 , \9962_b1 , \9962_b0 , \9963_b1 , \9963_b0 , \9964_b1 , \9964_b0 , 
		\9965_b1 , \9965_b0 , \9966_b1 , \9966_b0 , \9967_b1 , \9967_b0 , \9968_b1 , \9968_b0 , \9969_b1 , \9969_b0 , 
		\9970_b1 , \9970_b0 , \9971_b1 , \9971_b0 , \9972_b1 , \9972_b0 , \9973_b1 , \9973_b0 , \9974_b1 , \9974_b0 , 
		\9975_b1 , \9975_b0 , \9976_b1 , \9976_b0 , \9977_b1 , \9977_b0 , \9978_b1 , \9978_b0 , \9979_b1 , \9979_b0 , 
		\9980_b1 , \9980_b0 , \9981_b1 , \9981_b0 , \9982_b1 , \9982_b0 , \9983_b1 , \9983_b0 , \9984_b1 , \9984_b0 , 
		\9985_b1 , \9985_b0 , \9986_b1 , \9986_b0 , \9987_b1 , \9987_b0 , \9988_b1 , \9988_b0 , \9989_b1 , \9989_b0 , 
		\9990_b1 , \9990_b0 , \9991_b1 , \9991_b0 , \9992_b1 , \9992_b0 , \9993_b1 , \9993_b0 , \9994_b1 , \9994_b0 , 
		\9995_b1 , \9995_b0 , \9996_b1 , \9996_b0 , \9997_b1 , \9997_b0 , \9998_b1 , \9998_b0 , \9999_b1 , \9999_b0 , 
		\10000_b1 , \10000_b0 , \10001_b1 , \10001_b0 , \10002_b1 , \10002_b0 , \10003_b1 , \10003_b0 , \10004_b1 , \10004_b0 , 
		\10005_b1 , \10005_b0 , \10006_b1 , \10006_b0 , \10007_b1 , \10007_b0 , \10008_b1 , \10008_b0 , \10009_b1 , \10009_b0 , 
		\10010_b1 , \10010_b0 , \10011_b1 , \10011_b0 , \10012_b1 , \10012_b0 , \10013_b1 , \10013_b0 , \10014_b1 , \10014_b0 , 
		\10015_b1 , \10015_b0 , \10016_b1 , \10016_b0 , \10017_b1 , \10017_b0 , \10018_b1 , \10018_b0 , \10019_b1 , \10019_b0 , 
		\10020_b1 , \10020_b0 , \10021_b1 , \10021_b0 , \10022_b1 , \10022_b0 , \10023_b1 , \10023_b0 , \10024_b1 , \10024_b0 , 
		\10025_b1 , \10025_b0 , \10026_b1 , \10026_b0 , \10027_b1 , \10027_b0 , \10028_b1 , \10028_b0 , \10029_b1 , \10029_b0 , 
		\10030_b1 , \10030_b0 , \10031_b1 , \10031_b0 , \10032_b1 , \10032_b0 , \10033_b1 , \10033_b0 , \10034_b1 , \10034_b0 , 
		\10035_b1 , \10035_b0 , \10036_b1 , \10036_b0 , \10037_b1 , \10037_b0 , \10038_b1 , \10038_b0 , \10039_b1 , \10039_b0 , 
		\10040_b1 , \10040_b0 , \10041_b1 , \10041_b0 , \10042_b1 , \10042_b0 , \10043_b1 , \10043_b0 , \10044_b1 , \10044_b0 , 
		\10045_b1 , \10045_b0 , \10046_b1 , \10046_b0 , \10047_b1 , \10047_b0 , \10048_b1 , \10048_b0 , \10049_b1 , \10049_b0 , 
		\10050_b1 , \10050_b0 , \10051_b1 , \10051_b0 , \10052_b1 , \10052_b0 , \10053_b1 , \10053_b0 , \10054_b1 , \10054_b0 , 
		\10055_b1 , \10055_b0 , \10056_b1 , \10056_b0 , \10057_b1 , \10057_b0 , \10058_b1 , \10058_b0 , \10059_b1 , \10059_b0 , 
		\10060_b1 , \10060_b0 , \10061_b1 , \10061_b0 , \10062_b1 , \10062_b0 , \10063_b1 , \10063_b0 , \10064_b1 , \10064_b0 , 
		\10065_b1 , \10065_b0 , \10066_b1 , \10066_b0 , \10067_b1 , \10067_b0 , \10068_b1 , \10068_b0 , \10069_b1 , \10069_b0 , 
		\10070_b1 , \10070_b0 , \10071_b1 , \10071_b0 , \10072_b1 , \10072_b0 , \10073_b1 , \10073_b0 , \10074_b1 , \10074_b0 , 
		\10075_b1 , \10075_b0 , \10076_b1 , \10076_b0 , \10077_b1 , \10077_b0 , \10078_b1 , \10078_b0 , \10079_b1 , \10079_b0 , 
		\10080_b1 , \10080_b0 , \10081_b1 , \10081_b0 , \10082_b1 , \10082_b0 , \10083_b1 , \10083_b0 , \10084_b1 , \10084_b0 , 
		\10085_b1 , \10085_b0 , \10086_b1 , \10086_b0 , \10087_b1 , \10087_b0 , \10088_b1 , \10088_b0 , \10089_b1 , \10089_b0 , 
		\10090_b1 , \10090_b0 , \10091_b1 , \10091_b0 , \10092_b1 , \10092_b0 , \10093_b1 , \10093_b0 , \10094_b1 , \10094_b0 , 
		\10095_b1 , \10095_b0 , \10096_b1 , \10096_b0 , \10097_b1 , \10097_b0 , \10098_b1 , \10098_b0 , \10099_b1 , \10099_b0 , 
		\10100_b1 , \10100_b0 , \10101_b1 , \10101_b0 , \10102_b1 , \10102_b0 , \10103_b1 , \10103_b0 , \10104_b1 , \10104_b0 , 
		\10105_b1 , \10105_b0 , \10106_b1 , \10106_b0 , \10107_b1 , \10107_b0 , \10108_b1 , \10108_b0 , \10109_b1 , \10109_b0 , 
		\10110_b1 , \10110_b0 , \10111_b1 , \10111_b0 , \10112_b1 , \10112_b0 , \10113_b1 , \10113_b0 , \10114_b1 , \10114_b0 , 
		\10115_b1 , \10115_b0 , \10116_b1 , \10116_b0 , \10117_b1 , \10117_b0 , \10118_b1 , \10118_b0 , \10119_b1 , \10119_b0 , 
		\10120_b1 , \10120_b0 , \10121_b1 , \10121_b0 , \10122_b1 , \10122_b0 , \10123_b1 , \10123_b0 , \10124_b1 , \10124_b0 , 
		\10125_b1 , \10125_b0 , \10126_b1 , \10126_b0 , \10127_b1 , \10127_b0 , \10128_b1 , \10128_b0 , \10129_b1 , \10129_b0 , 
		\10130_b1 , \10130_b0 , \10131_b1 , \10131_b0 , \10132_b1 , \10132_b0 , \10133_b1 , \10133_b0 , \10134_b1 , \10134_b0 , 
		\10135_b1 , \10135_b0 , \10136_b1 , \10136_b0 , \10137_b1 , \10137_b0 , \10138_b1 , \10138_b0 , \10139_b1 , \10139_b0 , 
		\10140_b1 , \10140_b0 , \10141_b1 , \10141_b0 , \10142_b1 , \10142_b0 , \10143_b1 , \10143_b0 , \10144_b1 , \10144_b0 , 
		\10145_b1 , \10145_b0 , \10146_b1 , \10146_b0 , \10147_b1 , \10147_b0 , \10148_b1 , \10148_b0 , \10149_b1 , \10149_b0 , 
		\10150_b1 , \10150_b0 , \10151_b1 , \10151_b0 , \10152_b1 , \10152_b0 , \10153_b1 , \10153_b0 , \10154_b1 , \10154_b0 , 
		\10155_b1 , \10155_b0 , \10156_b1 , \10156_b0 , \10157_b1 , \10157_b0 , \10158_b1 , \10158_b0 , \10159_b1 , \10159_b0 , 
		\10160_b1 , \10160_b0 , \10161_b1 , \10161_b0 , \10162_b1 , \10162_b0 , \10163_b1 , \10163_b0 , \10164_b1 , \10164_b0 , 
		\10165_b1 , \10165_b0 , \10166_b1 , \10166_b0 , \10167_b1 , \10167_b0 , \10168_b1 , \10168_b0 , \10169_b1 , \10169_b0 , 
		\10170_b1 , \10170_b0 , \10171_b1 , \10171_b0 , \10172_b1 , \10172_b0 , \10173_b1 , \10173_b0 , \10174_b1 , \10174_b0 , 
		\10175_b1 , \10175_b0 , \10176_b1 , \10176_b0 , \10177_b1 , \10177_b0 , \10178_b1 , \10178_b0 , \10179_b1 , \10179_b0 , 
		\10180_b1 , \10180_b0 , \10181_b1 , \10181_b0 , \10182_b1 , \10182_b0 , \10183_b1 , \10183_b0 , \10184_b1 , \10184_b0 , 
		\10185_b1 , \10185_b0 , \10186_b1 , \10186_b0 , \10187_b1 , \10187_b0 , \10188_b1 , \10188_b0 , \10189_b1 , \10189_b0 , 
		\10190_b1 , \10190_b0 , \10191_b1 , \10191_b0 , \10192_b1 , \10192_b0 , \10193_b1 , \10193_b0 , \10194_b1 , \10194_b0 , 
		\10195_b1 , \10195_b0 , \10196_b1 , \10196_b0 , \10197_b1 , \10197_b0 , \10198_b1 , \10198_b0 , \10199_b1 , \10199_b0 , 
		\10200_b1 , \10200_b0 , \10201_b1 , \10201_b0 , \10202_b1 , \10202_b0 , \10203_b1 , \10203_b0 , \10204_b1 , \10204_b0 , 
		\10205_b1 , \10205_b0 , \10206_b1 , \10206_b0 , \10207_b1 , \10207_b0 , \10208_b1 , \10208_b0 , \10209_b1 , \10209_b0 , 
		\10210_b1 , \10210_b0 , \10211_b1 , \10211_b0 , \10212_b1 , \10212_b0 , \10213_b1 , \10213_b0 , \10214_b1 , \10214_b0 , 
		\10215_b1 , \10215_b0 , \10216_b1 , \10216_b0 , \10217_b1 , \10217_b0 , \10218_b1 , \10218_b0 , \10219_b1 , \10219_b0 , 
		\10220_b1 , \10220_b0 , \10221_b1 , \10221_b0 , \10222_b1 , \10222_b0 , \10223_b1 , \10223_b0 , \10224_b1 , \10224_b0 , 
		\10225_b1 , \10225_b0 , \10226_b1 , \10226_b0 , \10227_b1 , \10227_b0 , \10228_b1 , \10228_b0 , \10229_b1 , \10229_b0 , 
		\10230_b1 , \10230_b0 , \10231_b1 , \10231_b0 , \10232_b1 , \10232_b0 , \10233_b1 , \10233_b0 , \10234_b1 , \10234_b0 , 
		\10235_b1 , \10235_b0 , \10236_b1 , \10236_b0 , \10237_b1 , \10237_b0 , \10238_b1 , \10238_b0 , \10239_b1 , \10239_b0 , 
		\10240_b1 , \10240_b0 , \10241_b1 , \10241_b0 , \10242_b1 , \10242_b0 , \10243_b1 , \10243_b0 , \10244_b1 , \10244_b0 , 
		\10245_b1 , \10245_b0 , \10246_b1 , \10246_b0 , \10247_b1 , \10247_b0 , \10248_b1 , \10248_b0 , \10249_b1 , \10249_b0 , 
		\10250_b1 , \10250_b0 , \10251_b1 , \10251_b0 , \10252_b1 , \10252_b0 , \10253_b1 , \10253_b0 , \10254_b1 , \10254_b0 , 
		\10255_b1 , \10255_b0 , \10256_b1 , \10256_b0 , \10257_b1 , \10257_b0 , \10258_b1 , \10258_b0 , \10259_b1 , \10259_b0 , 
		\10260_b1 , \10260_b0 , \10261_b1 , \10261_b0 , \10262_b1 , \10262_b0 , \10263_b1 , \10263_b0 , \10264_b1 , \10264_b0 , 
		\10265_b1 , \10265_b0 , \10266_b1 , \10266_b0 , \10267_b1 , \10267_b0 , \10268_b1 , \10268_b0 , \10269_b1 , \10269_b0 , 
		\10270_b1 , \10270_b0 , \10271_b1 , \10271_b0 , \10272_b1 , \10272_b0 , \10273_b1 , \10273_b0 , \10274_b1 , \10274_b0 , 
		\10275_b1 , \10275_b0 , \10276_b1 , \10276_b0 , \10277_b1 , \10277_b0 , \10278_b1 , \10278_b0 , \10279_b1 , \10279_b0 , 
		\10280_b1 , \10280_b0 , \10281_b1 , \10281_b0 , \10282_b1 , \10282_b0 , \10283_b1 , \10283_b0 , \10284_b1 , \10284_b0 , 
		\10285_b1 , \10285_b0 , \10286_b1 , \10286_b0 , \10287_b1 , \10287_b0 , \10288_b1 , \10288_b0 , \10289_b1 , \10289_b0 , 
		\10290_b1 , \10290_b0 , \10291_b1 , \10291_b0 , \10292_b1 , \10292_b0 , \10293_b1 , \10293_b0 , \10294_b1 , \10294_b0 , 
		\10295_b1 , \10295_b0 , \10296_b1 , \10296_b0 , \10297_b1 , \10297_b0 , \10298_b1 , \10298_b0 , \10299_b1 , \10299_b0 , 
		\10300_b1 , \10300_b0 , \10301_b1 , \10301_b0 , \10302_b1 , \10302_b0 , \10303_b1 , \10303_b0 , \10304_b1 , \10304_b0 , 
		\10305_b1 , \10305_b0 , \10306_b1 , \10306_b0 , \10307_b1 , \10307_b0 , \10308_b1 , \10308_b0 , \10309_b1 , \10309_b0 , 
		\10310_b1 , \10310_b0 , \10311_b1 , \10311_b0 , \10312_b1 , \10312_b0 , \10313_b1 , \10313_b0 , \10314_b1 , \10314_b0 , 
		\10315_b1 , \10315_b0 , \10316_b1 , \10316_b0 , \10317_b1 , \10317_b0 , \10318_b1 , \10318_b0 , \10319_b1 , \10319_b0 , 
		\10320_b1 , \10320_b0 , \10321_b1 , \10321_b0 , \10322_b1 , \10322_b0 , \10323_b1 , \10323_b0 , \10324_b1 , \10324_b0 , 
		\10325_b1 , \10325_b0 , \10326_b1 , \10326_b0 , \10327_b1 , \10327_b0 , \10328_b1 , \10328_b0 , \10329_b1 , \10329_b0 , 
		\10330_b1 , \10330_b0 , \10331_b1 , \10331_b0 , \10332_b1 , \10332_b0 , \10333_b1 , \10333_b0 , \10334_b1 , \10334_b0 , 
		\10335_b1 , \10335_b0 , \10336_b1 , \10336_b0 , \10337_b1 , \10337_b0 , \10338_b1 , \10338_b0 , \10339_b1 , \10339_b0 , 
		\10340_b1 , \10340_b0 , \10341_b1 , \10341_b0 , \10342_b1 , \10342_b0 , \10343_b1 , \10343_b0 , \10344_b1 , \10344_b0 , 
		\10345_b1 , \10345_b0 , \10346_b1 , \10346_b0 , \10347_b1 , \10347_b0 , \10348_b1 , \10348_b0 , \10349_b1 , \10349_b0 , 
		\10350_b1 , \10350_b0 , \10351_b1 , \10351_b0 , \10352_b1 , \10352_b0 , \10353_b1 , \10353_b0 , \10354_b1 , \10354_b0 , 
		\10355_b1 , \10355_b0 , \10356_b1 , \10356_b0 , \10357_b1 , \10357_b0 , \10358_b1 , \10358_b0 , \10359_b1 , \10359_b0 , 
		\10360_b1 , \10360_b0 , \10361_b1 , \10361_b0 , \10362_b1 , \10362_b0 , \10363_b1 , \10363_b0 , \10364_b1 , \10364_b0 , 
		\10365_b1 , \10365_b0 , \10366_b1 , \10366_b0 , \10367_b1 , \10367_b0 , \10368_b1 , \10368_b0 , \10369_b1 , \10369_b0 , 
		\10370_b1 , \10370_b0 , \10371_b1 , \10371_b0 , \10372_b1 , \10372_b0 , \10373_b1 , \10373_b0 , \10374_b1 , \10374_b0 , 
		\10375_b1 , \10375_b0 , \10376_b1 , \10376_b0 , \10377_b1 , \10377_b0 , \10378_b1 , \10378_b0 , \10379_b1 , \10379_b0 , 
		\10380_b1 , \10380_b0 , \10381_b1 , \10381_b0 , \10382_b1 , \10382_b0 , \10383_b1 , \10383_b0 , \10384_b1 , \10384_b0 , 
		\10385_b1 , \10385_b0 , \10386_b1 , \10386_b0 , \10387_b1 , \10387_b0 , \10388_b1 , \10388_b0 , \10389_b1 , \10389_b0 , 
		\10390_b1 , \10390_b0 , \10391_b1 , \10391_b0 , \10392_b1 , \10392_b0 , \10393_b1 , \10393_b0 , \10394_b1 , \10394_b0 , 
		\10395_b1 , \10395_b0 , \10396_b1 , \10396_b0 , \10397_b1 , \10397_b0 , \10398_b1 , \10398_b0 , \10399_b1 , \10399_b0 , 
		\10400_b1 , \10400_b0 , \10401_b1 , \10401_b0 , \10402_b1 , \10402_b0 , \10403_b1 , \10403_b0 , \10404_b1 , \10404_b0 , 
		\10405_b1 , \10405_b0 , \10406_b1 , \10406_b0 , \10407_b1 , \10407_b0 , \10408_b1 , \10408_b0 , \10409_b1 , \10409_b0 , 
		\10410_b1 , \10410_b0 , \10411_b1 , \10411_b0 , \10412_b1 , \10412_b0 , \10413_b1 , \10413_b0 , \10414_b1 , \10414_b0 , 
		\10415_b1 , \10415_b0 , \10416_b1 , \10416_b0 , \10417_b1 , \10417_b0 , \10418_b1 , \10418_b0 , \10419_b1 , \10419_b0 , 
		\10420_b1 , \10420_b0 , \10421_b1 , \10421_b0 , \10422_b1 , \10422_b0 , \10423_b1 , \10423_b0 , \10424_b1 , \10424_b0 , 
		\10425_b1 , \10425_b0 , \10426_b1 , \10426_b0 , \10427_b1 , \10427_b0 , \10428_b1 , \10428_b0 , \10429_b1 , \10429_b0 , 
		\10430_b1 , \10430_b0 , \10431_b1 , \10431_b0 , \10432_b1 , \10432_b0 , \10433_b1 , \10433_b0 , \10434_b1 , \10434_b0 , 
		\10435_b1 , \10435_b0 , \10436_b1 , \10436_b0 , \10437_b1 , \10437_b0 , \10438_b1 , \10438_b0 , \10439_b1 , \10439_b0 , 
		\10440_b1 , \10440_b0 , \10441_b1 , \10441_b0 , \10442_b1 , \10442_b0 , \10443_b1 , \10443_b0 , \10444_b1 , \10444_b0 , 
		\10445_b1 , \10445_b0 , \10446_b1 , \10446_b0 , \10447_b1 , \10447_b0 , \10448_b1 , \10448_b0 , \10449_b1 , \10449_b0 , 
		\10450_b1 , \10450_b0 , \10451_b1 , \10451_b0 , \10452_b1 , \10452_b0 , \10453_b1 , \10453_b0 , \10454_b1 , \10454_b0 , 
		\10455_b1 , \10455_b0 , \10456_b1 , \10456_b0 , \10457_b1 , \10457_b0 , \10458_b1 , \10458_b0 , \10459_b1 , \10459_b0 , 
		\10460_b1 , \10460_b0 , \10461_b1 , \10461_b0 , \10462_b1 , \10462_b0 , \10463_b1 , \10463_b0 , \10464_b1 , \10464_b0 , 
		\10465_b1 , \10465_b0 , \10466_b1 , \10466_b0 , \10467_b1 , \10467_b0 , \10468_b1 , \10468_b0 , \10469_b1 , \10469_b0 , 
		\10470_b1 , \10470_b0 , \10471_b1 , \10471_b0 , \10472_b1 , \10472_b0 , \10473_b1 , \10473_b0 , \10474_b1 , \10474_b0 , 
		\10475_b1 , \10475_b0 , \10476_b1 , \10476_b0 , \10477_b1 , \10477_b0 , \10478_b1 , \10478_b0 , \10479_b1 , \10479_b0 , 
		\10480_b1 , \10480_b0 , \10481_b1 , \10481_b0 , \10482_b1 , \10482_b0 , \10483_b1 , \10483_b0 , \10484_b1 , \10484_b0 , 
		\10485_b1 , \10485_b0 , \10486_b1 , \10486_b0 , \10487_b1 , \10487_b0 , \10488_b1 , \10488_b0 , \10489_b1 , \10489_b0 , 
		\10490_b1 , \10490_b0 , \10491_b1 , \10491_b0 , \10492_b1 , \10492_b0 , \10493_b1 , \10493_b0 , \10494_b1 , \10494_b0 , 
		\10495_b1 , \10495_b0 , \10496_b1 , \10496_b0 , \10497_b1 , \10497_b0 , \10498_b1 , \10498_b0 , \10499_b1 , \10499_b0 , 
		\10500_b1 , \10500_b0 , \10501_b1 , \10501_b0 , \10502_b1 , \10502_b0 , \10503_b1 , \10503_b0 , \10504_b1 , \10504_b0 , 
		\10505_b1 , \10505_b0 , \10506_b1 , \10506_b0 , \10507_b1 , \10507_b0 , \10508_b1 , \10508_b0 , \10509_b1 , \10509_b0 , 
		\10510_b1 , \10510_b0 , \10511_b1 , \10511_b0 , \10512_b1 , \10512_b0 , \10513_b1 , \10513_b0 , \10514_b1 , \10514_b0 , 
		\10515_b1 , \10515_b0 , \10516_b1 , \10516_b0 , \10517_b1 , \10517_b0 , \10518_b1 , \10518_b0 , \10519_b1 , \10519_b0 , 
		\10520_b1 , \10520_b0 , \10521_b1 , \10521_b0 , \10522_b1 , \10522_b0 , \10523_b1 , \10523_b0 , \10524_b1 , \10524_b0 , 
		\10525_b1 , \10525_b0 , \10526_b1 , \10526_b0 , \10527_b1 , \10527_b0 , \10528_b1 , \10528_b0 , \10529_b1 , \10529_b0 , 
		\10530_b1 , \10530_b0 , \10531_b1 , \10531_b0 , \10532_b1 , \10532_b0 , \10533_b1 , \10533_b0 , \10534_b1 , \10534_b0 , 
		\10535_b1 , \10535_b0 , \10536_b1 , \10536_b0 , \10537_b1 , \10537_b0 , \10538_b1 , \10538_b0 , \10539_b1 , \10539_b0 , 
		\10540_b1 , \10540_b0 , \10541_b1 , \10541_b0 , \10542_b1 , \10542_b0 , \10543_b1 , \10543_b0 , \10544_b1 , \10544_b0 , 
		\10545_b1 , \10545_b0 , \10546_b1 , \10546_b0 , \10547_b1 , \10547_b0 , \10548_b1 , \10548_b0 , \10549_b1 , \10549_b0 , 
		\10550_b1 , \10550_b0 , \10551_b1 , \10551_b0 , \10552_b1 , \10552_b0 , \10553_b1 , \10553_b0 , \10554_b1 , \10554_b0 , 
		\10555_b1 , \10555_b0 , \10556_b1 , \10556_b0 , \10557_b1 , \10557_b0 , \10558_b1 , \10558_b0 , \10559_b1 , \10559_b0 , 
		\10560_b1 , \10560_b0 , \10561_b1 , \10561_b0 , \10562_b1 , \10562_b0 , \10563_b1 , \10563_b0 , \10564_b1 , \10564_b0 , 
		\10565_b1 , \10565_b0 , \10566_b1 , \10566_b0 , \10567_b1 , \10567_b0 , \10568_b1 , \10568_b0 , \10569_b1 , \10569_b0 , 
		\10570_b1 , \10570_b0 , \10571_b1 , \10571_b0 , \10572_b1 , \10572_b0 , \10573_b1 , \10573_b0 , \10574_b1 , \10574_b0 , 
		\10575_b1 , \10575_b0 , \10576_b1 , \10576_b0 , \10577_b1 , \10577_b0 , \10578_b1 , \10578_b0 , \10579_b1 , \10579_b0 , 
		\10580_b1 , \10580_b0 , \10581_b1 , \10581_b0 , \10582_b1 , \10582_b0 , \10583_b1 , \10583_b0 , \10584_b1 , \10584_b0 , 
		\10585_b1 , \10585_b0 , \10586_b1 , \10586_b0 , \10587_b1 , \10587_b0 , \10588_b1 , \10588_b0 , \10589_b1 , \10589_b0 , 
		\10590_b1 , \10590_b0 , \10591_b1 , \10591_b0 , \10592_b1 , \10592_b0 , \10593_b1 , \10593_b0 , \10594_b1 , \10594_b0 , 
		\10595_b1 , \10595_b0 , \10596_b1 , \10596_b0 , \10597_b1 , \10597_b0 , \10598_b1 , \10598_b0 , \10599_b1 , \10599_b0 , 
		\10600_b1 , \10600_b0 , \10601_b1 , \10601_b0 , \10602_b1 , \10602_b0 , \10603_b1 , \10603_b0 , \10604_b1 , \10604_b0 , 
		\10605_b1 , \10605_b0 , \10606_b1 , \10606_b0 , \10607_b1 , \10607_b0 , \10608_b1 , \10608_b0 , \10609_b1 , \10609_b0 , 
		\10610_b1 , \10610_b0 , \10611_b1 , \10611_b0 , \10612_b1 , \10612_b0 , \10613_b1 , \10613_b0 , \10614_b1 , \10614_b0 , 
		\10615_b1 , \10615_b0 , \10616_b1 , \10616_b0 , \10617_b1 , \10617_b0 , \10618_b1 , \10618_b0 , \10619_b1 , \10619_b0 , 
		\10620_b1 , \10620_b0 , \10621_b1 , \10621_b0 , \10622_b1 , \10622_b0 , \10623_b1 , \10623_b0 , \10624_b1 , \10624_b0 , 
		\10625_b1 , \10625_b0 , \10626_b1 , \10626_b0 , \10627_b1 , \10627_b0 , \10628_b1 , \10628_b0 , \10629_b1 , \10629_b0 , 
		\10630_b1 , \10630_b0 , \10631_b1 , \10631_b0 , \10632_b1 , \10632_b0 , \10633_b1 , \10633_b0 , \10634_b1 , \10634_b0 , 
		\10635_b1 , \10635_b0 , \10636_b1 , \10636_b0 , \10637_b1 , \10637_b0 , \10638_b1 , \10638_b0 , \10639_b1 , \10639_b0 , 
		\10640_b1 , \10640_b0 , \10641_b1 , \10641_b0 , \10642_b1 , \10642_b0 , \10643_b1 , \10643_b0 , \10644_b1 , \10644_b0 , 
		\10645_b1 , \10645_b0 , \10646_b1 , \10646_b0 , \10647_b1 , \10647_b0 , \10648_b1 , \10648_b0 , \10649_b1 , \10649_b0 , 
		\10650_b1 , \10650_b0 , \10651_b1 , \10651_b0 , \10652_b1 , \10652_b0 , \10653_b1 , \10653_b0 , \10654_b1 , \10654_b0 , 
		\10655_b1 , \10655_b0 , \10656_b1 , \10656_b0 , \10657_b1 , \10657_b0 , \10658_b1 , \10658_b0 , \10659_b1 , \10659_b0 , 
		\10660_b1 , \10660_b0 , \10661_b1 , \10661_b0 , \10662_b1 , \10662_b0 , \10663_b1 , \10663_b0 , \10664_b1 , \10664_b0 , 
		\10665_b1 , \10665_b0 , \10666_b1 , \10666_b0 , \10667_b1 , \10667_b0 , \10668_b1 , \10668_b0 , \10669_b1 , \10669_b0 , 
		\10670_b1 , \10670_b0 , \10671_b1 , \10671_b0 , \10672_b1 , \10672_b0 , \10673_b1 , \10673_b0 , \10674_b1 , \10674_b0 , 
		\10675_b1 , \10675_b0 , \10676_b1 , \10676_b0 , \10677_b1 , \10677_b0 , \10678_b1 , \10678_b0 , \10679_b1 , \10679_b0 , 
		\10680_b1 , \10680_b0 , \10681_b1 , \10681_b0 , \10682_b1 , \10682_b0 , \10683_b1 , \10683_b0 , \10684_b1 , \10684_b0 , 
		\10685_b1 , \10685_b0 , \10686_b1 , \10686_b0 , \10687_b1 , \10687_b0 , \10688_b1 , \10688_b0 , \10689_b1 , \10689_b0 , 
		\10690_b1 , \10690_b0 , \10691_b1 , \10691_b0 , \10692_b1 , \10692_b0 , \10693_b1 , \10693_b0 , \10694_b1 , \10694_b0 , 
		\10695_b1 , \10695_b0 , \10696_b1 , \10696_b0 , \10697_b1 , \10697_b0 , \10698_b1 , \10698_b0 , \10699_b1 , \10699_b0 , 
		\10700_b1 , \10700_b0 , \10701_b1 , \10701_b0 , \10702_b1 , \10702_b0 , \10703_b1 , \10703_b0 , \10704_b1 , \10704_b0 , 
		\10705_b1 , \10705_b0 , \10706_b1 , \10706_b0 , \10707_b1 , \10707_b0 , \10708_b1 , \10708_b0 , \10709_b1 , \10709_b0 , 
		\10710_b1 , \10710_b0 , \10711_b1 , \10711_b0 , \10712_b1 , \10712_b0 , \10713_b1 , \10713_b0 , \10714_b1 , \10714_b0 , 
		\10715_b1 , \10715_b0 , \10716_b1 , \10716_b0 , \10717_b1 , \10717_b0 , \10718_b1 , \10718_b0 , \10719_b1 , \10719_b0 , 
		\10720_b1 , \10720_b0 , \10721_b1 , \10721_b0 , \10722_b1 , \10722_b0 , \10723_b1 , \10723_b0 , \10724_b1 , \10724_b0 , 
		\10725_b1 , \10725_b0 , \10726_b1 , \10726_b0 , \10727_b1 , \10727_b0 , \10728_b1 , \10728_b0 , \10729_b1 , \10729_b0 , 
		\10730_b1 , \10730_b0 , \10731_b1 , \10731_b0 , \10732_b1 , \10732_b0 , \10733_b1 , \10733_b0 , \10734_b1 , \10734_b0 , 
		\10735_b1 , \10735_b0 , \10736_b1 , \10736_b0 , \10737_b1 , \10737_b0 , \10738_b1 , \10738_b0 , \10739_b1 , \10739_b0 , 
		\10740_b1 , \10740_b0 , \10741_b1 , \10741_b0 , \10742_b1 , \10742_b0 , \10743_b1 , \10743_b0 , \10744_b1 , \10744_b0 , 
		\10745_b1 , \10745_b0 , \10746_b1 , \10746_b0 , \10747_b1 , \10747_b0 , \10748_b1 , \10748_b0 , \10749_b1 , \10749_b0 , 
		\10750_b1 , \10750_b0 , \10751_b1 , \10751_b0 , \10752_b1 , \10752_b0 , \10753_b1 , \10753_b0 , \10754_b1 , \10754_b0 , 
		\10755_b1 , \10755_b0 , \10756_b1 , \10756_b0 , \10757_b1 , \10757_b0 , \10758_b1 , \10758_b0 , \10759_b1 , \10759_b0 , 
		\10760_b1 , \10760_b0 , \10761_b1 , \10761_b0 , \10762_b1 , \10762_b0 , \10763_b1 , \10763_b0 , \10764_b1 , \10764_b0 , 
		\10765_b1 , \10765_b0 , \10766_b1 , \10766_b0 , \10767_b1 , \10767_b0 , \10768_b1 , \10768_b0 , \10769_b1 , \10769_b0 , 
		\10770_b1 , \10770_b0 , \10771_b1 , \10771_b0 , \10772_b1 , \10772_b0 , \10773_b1 , \10773_b0 , \10774_b1 , \10774_b0 , 
		\10775_b1 , \10775_b0 , \10776_b1 , \10776_b0 , \10777_b1 , \10777_b0 , \10778_b1 , \10778_b0 , \10779_b1 , \10779_b0 , 
		\10780_b1 , \10780_b0 , \10781_b1 , \10781_b0 , \10782_b1 , \10782_b0 , \10783_b1 , \10783_b0 , \10784_b1 , \10784_b0 , 
		\10785_b1 , \10785_b0 , \10786_b1 , \10786_b0 , \10787_b1 , \10787_b0 , \10788_b1 , \10788_b0 , \10789_b1 , \10789_b0 , 
		\10790_b1 , \10790_b0 , \10791_b1 , \10791_b0 , \10792_b1 , \10792_b0 , \10793_b1 , \10793_b0 , \10794_b1 , \10794_b0 , 
		\10795_b1 , \10795_b0 , \10796_b1 , \10796_b0 , \10797_b1 , \10797_b0 , \10798_b1 , \10798_b0 , \10799_b1 , \10799_b0 , 
		\10800_b1 , \10800_b0 , \10801_b1 , \10801_b0 , \10802_b1 , \10802_b0 , \10803_b1 , \10803_b0 , \10804_b1 , \10804_b0 , 
		\10805_b1 , \10805_b0 , \10806_b1 , \10806_b0 , \10807_b1 , \10807_b0 , \10808_b1 , \10808_b0 , \10809_b1 , \10809_b0 , 
		\10810_b1 , \10810_b0 , \10811_b1 , \10811_b0 , \10812_b1 , \10812_b0 , \10813_b1 , \10813_b0 , \10814_b1 , \10814_b0 , 
		\10815_b1 , \10815_b0 , \10816_b1 , \10816_b0 , \10817_b1 , \10817_b0 , \10818_b1 , \10818_b0 , \10819_b1 , \10819_b0 , 
		\10820_b1 , \10820_b0 , \10821_b1 , \10821_b0 , \10822_b1 , \10822_b0 , \10823_b1 , \10823_b0 , \10824_b1 , \10824_b0 , 
		\10825_b1 , \10825_b0 , \10826_b1 , \10826_b0 , \10827_b1 , \10827_b0 , \10828_b1 , \10828_b0 , \10829_b1 , \10829_b0 , 
		\10830_b1 , \10830_b0 , \10831_b1 , \10831_b0 , \10832_b1 , \10832_b0 , \10833_b1 , \10833_b0 , \10834_b1 , \10834_b0 , 
		\10835_b1 , \10835_b0 , \10836_b1 , \10836_b0 , \10837_b1 , \10837_b0 , \10838_b1 , \10838_b0 , \10839_b1 , \10839_b0 , 
		\10840_b1 , \10840_b0 , \10841_b1 , \10841_b0 , \10842_b1 , \10842_b0 , \10843_b1 , \10843_b0 , \10844_b1 , \10844_b0 , 
		\10845_b1 , \10845_b0 , \10846_b1 , \10846_b0 , \10847_b1 , \10847_b0 , \10848_b1 , \10848_b0 , \10849_b1 , \10849_b0 , 
		\10850_b1 , \10850_b0 , \10851_b1 , \10851_b0 , \10852_b1 , \10852_b0 , \10853_b1 , \10853_b0 , \10854_b1 , \10854_b0 , 
		\10855_b1 , \10855_b0 , \10856_b1 , \10856_b0 , \10857_b1 , \10857_b0 , \10858_b1 , \10858_b0 , \10859_b1 , \10859_b0 , 
		\10860_b1 , \10860_b0 , \10861_b1 , \10861_b0 , \10862_b1 , \10862_b0 , \10863_b1 , \10863_b0 , \10864_b1 , \10864_b0 , 
		\10865_b1 , \10865_b0 , \10866_b1 , \10866_b0 , \10867_b1 , \10867_b0 , \10868_b1 , \10868_b0 , \10869_b1 , \10869_b0 , 
		\10870_b1 , \10870_b0 , \10871_b1 , \10871_b0 , \10872_b1 , \10872_b0 , \10873_b1 , \10873_b0 , \10874_b1 , \10874_b0 , 
		\10875_b1 , \10875_b0 , \10876_b1 , \10876_b0 , \10877_b1 , \10877_b0 , \10878_b1 , \10878_b0 , \10879_b1 , \10879_b0 , 
		\10880_b1 , \10880_b0 , \10881_b1 , \10881_b0 , \10882_b1 , \10882_b0 , \10883_b1 , \10883_b0 , \10884_b1 , \10884_b0 , 
		\10885_b1 , \10885_b0 , \10886_b1 , \10886_b0 , \10887_b1 , \10887_b0 , \10888_b1 , \10888_b0 , \10889_b1 , \10889_b0 , 
		\10890_b1 , \10890_b0 , \10891_b1 , \10891_b0 , \10892_b1 , \10892_b0 , \10893_b1 , \10893_b0 , \10894_b1 , \10894_b0 , 
		\10895_b1 , \10895_b0 , \10896_b1 , \10896_b0 , \10897_b1 , \10897_b0 , \10898_b1 , \10898_b0 , \10899_b1 , \10899_b0 , 
		\10900_b1 , \10900_b0 , \10901_b1 , \10901_b0 , \10902_b1 , \10902_b0 , \10903_b1 , \10903_b0 , \10904_b1 , \10904_b0 , 
		\10905_b1 , \10905_b0 , \10906_b1 , \10906_b0 , \10907_b1 , \10907_b0 , \10908_b1 , \10908_b0 , \10909_b1 , \10909_b0 , 
		\10910_b1 , \10910_b0 , \10911_b1 , \10911_b0 , \10912_b1 , \10912_b0 , \10913_b1 , \10913_b0 , \10914_b1 , \10914_b0 , 
		\10915_b1 , \10915_b0 , \10916_b1 , \10916_b0 , \10917_b1 , \10917_b0 , \10918_b1 , \10918_b0 , \10919_b1 , \10919_b0 , 
		\10920_b1 , \10920_b0 , \10921_b1 , \10921_b0 , \10922_b1 , \10922_b0 , \10923_b1 , \10923_b0 , \10924_b1 , \10924_b0 , 
		\10925_b1 , \10925_b0 , \10926_b1 , \10926_b0 , \10927_b1 , \10927_b0 , \10928_b1 , \10928_b0 , \10929_b1 , \10929_b0 , 
		\10930_b1 , \10930_b0 , \10931_b1 , \10931_b0 , \10932_b1 , \10932_b0 , \10933_b1 , \10933_b0 , \10934_b1 , \10934_b0 , 
		\10935_b1 , \10935_b0 , \10936_b1 , \10936_b0 , \10937_b1 , \10937_b0 , \10938_b1 , \10938_b0 , \10939_b1 , \10939_b0 , 
		\10940_b1 , \10940_b0 , \10941_b1 , \10941_b0 , \10942_b1 , \10942_b0 , \10943_b1 , \10943_b0 , \10944_b1 , \10944_b0 , 
		\10945_b1 , \10945_b0 , \10946_b1 , \10946_b0 , \10947_b1 , \10947_b0 , \10948_b1 , \10948_b0 , \10949_b1 , \10949_b0 , 
		\10950_b1 , \10950_b0 , \10951_b1 , \10951_b0 , \10952_b1 , \10952_b0 , \10953_b1 , \10953_b0 , \10954_b1 , \10954_b0 , 
		\10955_b1 , \10955_b0 , \10956_b1 , \10956_b0 , \10957_b1 , \10957_b0 , \10958_b1 , \10958_b0 , \10959_b1 , \10959_b0 , 
		\10960_b1 , \10960_b0 , \10961_b1 , \10961_b0 , \10962_b1 , \10962_b0 , \10963_b1 , \10963_b0 , \10964_b1 , \10964_b0 , 
		\10965_b1 , \10965_b0 , \10966_b1 , \10966_b0 , \10967_b1 , \10967_b0 , \10968_b1 , \10968_b0 , \10969_b1 , \10969_b0 , 
		\10970_b1 , \10970_b0 , \10971_b1 , \10971_b0 , \10972_b1 , \10972_b0 , \10973_b1 , \10973_b0 , \10974_b1 , \10974_b0 , 
		\10975_b1 , \10975_b0 , \10976_b1 , \10976_b0 , \10977_b1 , \10977_b0 , \10978_b1 , \10978_b0 , \10979_b1 , \10979_b0 , 
		\10980_b1 , \10980_b0 , \10981_b1 , \10981_b0 , \10982_b1 , \10982_b0 , \10983_b1 , \10983_b0 , \10984_b1 , \10984_b0 , 
		\10985_b1 , \10985_b0 , \10986_b1 , \10986_b0 , \10987_b1 , \10987_b0 , \10988_b1 , \10988_b0 , \10989_b1 , \10989_b0 , 
		\10990_b1 , \10990_b0 , \10991_b1 , \10991_b0 , \10992_b1 , \10992_b0 , \10993_b1 , \10993_b0 , \10994_b1 , \10994_b0 , 
		\10995_b1 , \10995_b0 , \10996_b1 , \10996_b0 , \10997_b1 , \10997_b0 , \10998_b1 , \10998_b0 , \10999_b1 , \10999_b0 , 
		\11000_b1 , \11000_b0 , \11001_b1 , \11001_b0 , \11002_b1 , \11002_b0 , \11003_b1 , \11003_b0 , \11004_b1 , \11004_b0 , 
		\11005_b1 , \11005_b0 , \11006_b1 , \11006_b0 , \11007_b1 , \11007_b0 , \11008_b1 , \11008_b0 , \11009_b1 , \11009_b0 , 
		\11010_b1 , \11010_b0 , \11011_b1 , \11011_b0 , \11012_b1 , \11012_b0 , \11013_b1 , \11013_b0 , \11014_b1 , \11014_b0 , 
		\11015_b1 , \11015_b0 , \11016_b1 , \11016_b0 , \11017_b1 , \11017_b0 , \11018_b1 , \11018_b0 , \11019_b1 , \11019_b0 , 
		\11020_b1 , \11020_b0 , \11021_b1 , \11021_b0 , \11022_b1 , \11022_b0 , \11023_b1 , \11023_b0 , \11024_b1 , \11024_b0 , 
		\11025_b1 , \11025_b0 , \11026_b1 , \11026_b0 , \11027_b1 , \11027_b0 , \11028_b1 , \11028_b0 , \11029_b1 , \11029_b0 , 
		\11030_b1 , \11030_b0 , \11031_b1 , \11031_b0 , \11032_b1 , \11032_b0 , \11033_b1 , \11033_b0 , \11034_b1 , \11034_b0 , 
		\11035_b1 , \11035_b0 , \11036_b1 , \11036_b0 , \11037_b1 , \11037_b0 , \11038_b1 , \11038_b0 , \11039_b1 , \11039_b0 , 
		\11040_b1 , \11040_b0 , \11041_b1 , \11041_b0 , \11042_b1 , \11042_b0 , \11043_b1 , \11043_b0 , \11044_b1 , \11044_b0 , 
		\11045_b1 , \11045_b0 , \11046_b1 , \11046_b0 , \11047_b1 , \11047_b0 , \11048_b1 , \11048_b0 , \11049_b1 , \11049_b0 , 
		\11050_b1 , \11050_b0 , \11051_b1 , \11051_b0 , \11052_b1 , \11052_b0 , \11053_b1 , \11053_b0 , \11054_b1 , \11054_b0 , 
		\11055_b1 , \11055_b0 , \11056_b1 , \11056_b0 , \11057_b1 , \11057_b0 , \11058_b1 , \11058_b0 , \11059_b1 , \11059_b0 , 
		\11060_b1 , \11060_b0 , \11061_b1 , \11061_b0 , \11062_b1 , \11062_b0 , \11063_b1 , \11063_b0 , \11064_b1 , \11064_b0 , 
		\11065_b1 , \11065_b0 , \11066_b1 , \11066_b0 , \11067_b1 , \11067_b0 , \11068_b1 , \11068_b0 , \11069_b1 , \11069_b0 , 
		\11070_b1 , \11070_b0 , \11071_b1 , \11071_b0 , \11072_b1 , \11072_b0 , \11073_b1 , \11073_b0 , \11074_b1 , \11074_b0 , 
		\11075_b1 , \11075_b0 , \11076_b1 , \11076_b0 , \11077_b1 , \11077_b0 , \11078_b1 , \11078_b0 , \11079_b1 , \11079_b0 , 
		\11080_b1 , \11080_b0 , \11081_b1 , \11081_b0 , \11082_b1 , \11082_b0 , \11083_b1 , \11083_b0 , \11084_b1 , \11084_b0 , 
		\11085_b1 , \11085_b0 , \11086_b1 , \11086_b0 , \11087_b1 , \11087_b0 , \11088_b1 , \11088_b0 , \11089_b1 , \11089_b0 , 
		\11090_b1 , \11090_b0 , \11091_b1 , \11091_b0 , \11092_b1 , \11092_b0 , \11093_b1 , \11093_b0 , \11094_b1 , \11094_b0 , 
		\11095_b1 , \11095_b0 , \11096_b1 , \11096_b0 , \11097_b1 , \11097_b0 , \11098_b1 , \11098_b0 , \11099_b1 , \11099_b0 , 
		\11100_b1 , \11100_b0 , \11101_b1 , \11101_b0 , \11102_b1 , \11102_b0 , \11103_b1 , \11103_b0 , \11104_b1 , \11104_b0 , 
		\11105_b1 , \11105_b0 , \11106_b1 , \11106_b0 , \11107_b1 , \11107_b0 , \11108_b1 , \11108_b0 , \11109_b1 , \11109_b0 , 
		\11110_b1 , \11110_b0 , \11111_b1 , \11111_b0 , \11112_b1 , \11112_b0 , \11113_b1 , \11113_b0 , \11114_b1 , \11114_b0 , 
		\11115_b1 , \11115_b0 , \11116_b1 , \11116_b0 , \11117_b1 , \11117_b0 , \11118_b1 , \11118_b0 , \11119_b1 , \11119_b0 , 
		\11120_b1 , \11120_b0 , \11121_b1 , \11121_b0 , \11122_b1 , \11122_b0 , \11123_b1 , \11123_b0 , \11124_b1 , \11124_b0 , 
		\11125_b1 , \11125_b0 , \11126_b1 , \11126_b0 , \11127_b1 , \11127_b0 , \11128_b1 , \11128_b0 , \11129_b1 , \11129_b0 , 
		\11130_b1 , \11130_b0 , \11131_b1 , \11131_b0 , \11132_b1 , \11132_b0 , \11133_b1 , \11133_b0 , \11134_b1 , \11134_b0 , 
		\11135_b1 , \11135_b0 , \11136_b1 , \11136_b0 , \11137_b1 , \11137_b0 , \11138_b1 , \11138_b0 , \11139_b1 , \11139_b0 , 
		\11140_b1 , \11140_b0 , \11141_b1 , \11141_b0 , \11142_b1 , \11142_b0 , \11143_b1 , \11143_b0 , \11144_b1 , \11144_b0 , 
		\11145_b1 , \11145_b0 , \11146_b1 , \11146_b0 , \11147_b1 , \11147_b0 , \11148_b1 , \11148_b0 , \11149_b1 , \11149_b0 , 
		\11150_b1 , \11150_b0 , \11151_b1 , \11151_b0 , \11152_b1 , \11152_b0 , \11153_b1 , \11153_b0 , \11154_b1 , \11154_b0 , 
		\11155_b1 , \11155_b0 , \11156_b1 , \11156_b0 , \11157_b1 , \11157_b0 , \11158_b1 , \11158_b0 , \11159_b1 , \11159_b0 , 
		\11160_b1 , \11160_b0 , \11161_b1 , \11161_b0 , \11162_b1 , \11162_b0 , \11163_b1 , \11163_b0 , \11164_b1 , \11164_b0 , 
		\11165_b1 , \11165_b0 , \11166_b1 , \11166_b0 , \11167_b1 , \11167_b0 , \11168_b1 , \11168_b0 , \11169_b1 , \11169_b0 , 
		\11170_b1 , \11170_b0 , \11171_b1 , \11171_b0 , \11172_b1 , \11172_b0 , \11173_b1 , \11173_b0 , \11174_b1 , \11174_b0 , 
		\11175_b1 , \11175_b0 , \11176_b1 , \11176_b0 , \11177_b1 , \11177_b0 , \11178_b1 , \11178_b0 , \11179_b1 , \11179_b0 , 
		\11180_b1 , \11180_b0 , \11181_b1 , \11181_b0 , \11182_b1 , \11182_b0 , \11183_b1 , \11183_b0 , \11184_b1 , \11184_b0 , 
		\11185_b1 , \11185_b0 , \11186_b1 , \11186_b0 , \11187_b1 , \11187_b0 , \11188_b1 , \11188_b0 , \11189_b1 , \11189_b0 , 
		\11190_b1 , \11190_b0 , \11191_b1 , \11191_b0 , \11192_b1 , \11192_b0 , \11193_b1 , \11193_b0 , \11194_b1 , \11194_b0 , 
		\11195_b1 , \11195_b0 , \11196_b1 , \11196_b0 , \11197_b1 , \11197_b0 , \11198_b1 , \11198_b0 , \11199_b1 , \11199_b0 , 
		\11200_b1 , \11200_b0 , \11201_b1 , \11201_b0 , \11202_b1 , \11202_b0 , \11203_b1 , \11203_b0 , \11204_b1 , \11204_b0 , 
		\11205_b1 , \11205_b0 , \11206_b1 , \11206_b0 , \11207_b1 , \11207_b0 , \11208_b1 , \11208_b0 , \11209_b1 , \11209_b0 , 
		\11210_b1 , \11210_b0 , \11211_b1 , \11211_b0 , \11212_b1 , \11212_b0 , \11213_b1 , \11213_b0 , \11214_b1 , \11214_b0 , 
		\11215_b1 , \11215_b0 , \11216_b1 , \11216_b0 , \11217_b1 , \11217_b0 , \11218_b1 , \11218_b0 , \11219_b1 , \11219_b0 , 
		\11220_b1 , \11220_b0 , \11221_b1 , \11221_b0 , \11222_b1 , \11222_b0 , \11223_b1 , \11223_b0 , \11224_b1 , \11224_b0 , 
		\11225_b1 , \11225_b0 , \11226_b1 , \11226_b0 , \11227_b1 , \11227_b0 , \11228_b1 , \11228_b0 , \11229_b1 , \11229_b0 , 
		\11230_b1 , \11230_b0 , \11231_b1 , \11231_b0 , \11232_b1 , \11232_b0 , \11233_b1 , \11233_b0 , \11234_b1 , \11234_b0 , 
		\11235_b1 , \11235_b0 , \11236_b1 , \11236_b0 , \11237_b1 , \11237_b0 , \11238_b1 , \11238_b0 , \11239_b1 , \11239_b0 , 
		\11240_b1 , \11240_b0 , \11241_b1 , \11241_b0 , \11242_b1 , \11242_b0 , \11243_b1 , \11243_b0 , \11244_b1 , \11244_b0 , 
		\11245_b1 , \11245_b0 , \11246_b1 , \11246_b0 , \11247_b1 , \11247_b0 , \11248_b1 , \11248_b0 , \11249_b1 , \11249_b0 , 
		\11250_b1 , \11250_b0 , \11251_b1 , \11251_b0 , \11252_b1 , \11252_b0 , \11253_b1 , \11253_b0 , \11254_b1 , \11254_b0 , 
		\11255_b1 , \11255_b0 , \11256_b1 , \11256_b0 , \11257_b1 , \11257_b0 , \11258_b1 , \11258_b0 , \11259_b1 , \11259_b0 , 
		\11260_b1 , \11260_b0 , \11261_b1 , \11261_b0 , \11262_b1 , \11262_b0 , \11263_b1 , \11263_b0 , \11264_b1 , \11264_b0 , 
		\11265_b1 , \11265_b0 , \11266_b1 , \11266_b0 , \11267_b1 , \11267_b0 , \11268_b1 , \11268_b0 , \11269_b1 , \11269_b0 , 
		\11270_b1 , \11270_b0 , \11271_b1 , \11271_b0 , \11272_b1 , \11272_b0 , \11273_b1 , \11273_b0 , \11274_b1 , \11274_b0 , 
		\11275_b1 , \11275_b0 , \11276_b1 , \11276_b0 , \11277_b1 , \11277_b0 , \11278_b1 , \11278_b0 , \11279_b1 , \11279_b0 , 
		\11280_b1 , \11280_b0 , \11281_b1 , \11281_b0 , \11282_b1 , \11282_b0 , \11283_b1 , \11283_b0 , \11284_b1 , \11284_b0 , 
		\11285_b1 , \11285_b0 , \11286_b1 , \11286_b0 , \11287_b1 , \11287_b0 , \11288_b1 , \11288_b0 , \11289_b1 , \11289_b0 , 
		\11290_b1 , \11290_b0 , \11291_b1 , \11291_b0 , \11292_b1 , \11292_b0 , \11293_b1 , \11293_b0 , \11294_b1 , \11294_b0 , 
		\11295_b1 , \11295_b0 , \11296_b1 , \11296_b0 , \11297_b1 , \11297_b0 , \11298_b1 , \11298_b0 , \11299_b1 , \11299_b0 , 
		\11300_b1 , \11300_b0 , \11301_b1 , \11301_b0 , \11302_b1 , \11302_b0 , \11303_b1 , \11303_b0 , \11304_b1 , \11304_b0 , 
		\11305_b1 , \11305_b0 , \11306_b1 , \11306_b0 , \11307_b1 , \11307_b0 , \11308_b1 , \11308_b0 , \11309_b1 , \11309_b0 , 
		\11310_b1 , \11310_b0 , \11311_b1 , \11311_b0 , \11312_b1 , \11312_b0 , \11313_b1 , \11313_b0 , \11314_b1 , \11314_b0 , 
		\11315_b1 , \11315_b0 , \11316_b1 , \11316_b0 , \11317_b1 , \11317_b0 , \11318_b1 , \11318_b0 , \11319_b1 , \11319_b0 , 
		\11320_b1 , \11320_b0 , \11321_b1 , \11321_b0 , \11322_b1 , \11322_b0 , \11323_b1 , \11323_b0 , \11324_b1 , \11324_b0 , 
		\11325_b1 , \11325_b0 , \11326_b1 , \11326_b0 , \11327_b1 , \11327_b0 , \11328_b1 , \11328_b0 , \11329_b1 , \11329_b0 , 
		\11330_b1 , \11330_b0 , \11331_b1 , \11331_b0 , \11332_b1 , \11332_b0 , \11333_b1 , \11333_b0 , \11334_b1 , \11334_b0 , 
		\11335_b1 , \11335_b0 , \11336_b1 , \11336_b0 , \11337_b1 , \11337_b0 , \11338_b1 , \11338_b0 , \11339_b1 , \11339_b0 , 
		\11340_b1 , \11340_b0 , \11341_b1 , \11341_b0 , \11342_b1 , \11342_b0 , \11343_b1 , \11343_b0 , \11344_b1 , \11344_b0 , 
		\11345_b1 , \11345_b0 , \11346_b1 , \11346_b0 , \11347_b1 , \11347_b0 , \11348_b1 , \11348_b0 , \11349_b1 , \11349_b0 , 
		\11350_b1 , \11350_b0 , \11351_b1 , \11351_b0 , \11352_b1 , \11352_b0 , \11353_b1 , \11353_b0 , \11354_b1 , \11354_b0 , 
		\11355_b1 , \11355_b0 , \11356_b1 , \11356_b0 , \11357_b1 , \11357_b0 , \11358_b1 , \11358_b0 , \11359_b1 , \11359_b0 , 
		\11360_b1 , \11360_b0 , \11361_b1 , \11361_b0 , \11362_b1 , \11362_b0 , \11363_b1 , \11363_b0 , \11364_b1 , \11364_b0 , 
		\11365_b1 , \11365_b0 , \11366_b1 , \11366_b0 , \11367_b1 , \11367_b0 , \11368_b1 , \11368_b0 , \11369_b1 , \11369_b0 , 
		\11370_b1 , \11370_b0 , \11371_b1 , \11371_b0 , \11372_b1 , \11372_b0 , \11373_b1 , \11373_b0 , \11374_b1 , \11374_b0 , 
		\11375_b1 , \11375_b0 , \11376_b1 , \11376_b0 , \11377_b1 , \11377_b0 , \11378_b1 , \11378_b0 , \11379_b1 , \11379_b0 , 
		\11380_b1 , \11380_b0 , \11381_b1 , \11381_b0 , \11382_b1 , \11382_b0 , \11383_b1 , \11383_b0 , \11384_b1 , \11384_b0 , 
		\11385_b1 , \11385_b0 , \11386_b1 , \11386_b0 , \11387_b1 , \11387_b0 , \11388_b1 , \11388_b0 , \11389_b1 , \11389_b0 , 
		\11390_b1 , \11390_b0 , \11391_b1 , \11391_b0 , \11392_b1 , \11392_b0 , \11393_b1 , \11393_b0 , \11394_b1 , \11394_b0 , 
		\11395_b1 , \11395_b0 , \11396_b1 , \11396_b0 , \11397_b1 , \11397_b0 , \11398_b1 , \11398_b0 , \11399_b1 , \11399_b0 , 
		\11400_b1 , \11400_b0 , \11401_b1 , \11401_b0 , \11402_b1 , \11402_b0 , \11403_b1 , \11403_b0 , \11404_b1 , \11404_b0 , 
		\11405_b1 , \11405_b0 , \11406_b1 , \11406_b0 , \11407_b1 , \11407_b0 , \11408_b1 , \11408_b0 , \11409_b1 , \11409_b0 , 
		\11410_b1 , \11410_b0 , \11411_b1 , \11411_b0 , \11412_b1 , \11412_b0 , \11413_b1 , \11413_b0 , \11414_b1 , \11414_b0 , 
		\11415_b1 , \11415_b0 , \11416_b1 , \11416_b0 , \11417_b1 , \11417_b0 , \11418_b1 , \11418_b0 , \11419_b1 , \11419_b0 , 
		\11420_b1 , \11420_b0 , \11421_b1 , \11421_b0 , \11422_b1 , \11422_b0 , \11423_b1 , \11423_b0 , \11424_b1 , \11424_b0 , 
		\11425_b1 , \11425_b0 , \11426_b1 , \11426_b0 , \11427_b1 , \11427_b0 , \11428_b1 , \11428_b0 , \11429_b1 , \11429_b0 , 
		\11430_b1 , \11430_b0 , \11431_b1 , \11431_b0 , \11432_b1 , \11432_b0 , \11433_b1 , \11433_b0 , \11434_b1 , \11434_b0 , 
		\11435_b1 , \11435_b0 , \11436_b1 , \11436_b0 , \11437_b1 , \11437_b0 , \11438_b1 , \11438_b0 , \11439_b1 , \11439_b0 , 
		\11440_b1 , \11440_b0 , \11441_b1 , \11441_b0 , \11442_b1 , \11442_b0 , \11443_b1 , \11443_b0 , \11444_b1 , \11444_b0 , 
		\11445_b1 , \11445_b0 , \11446_b1 , \11446_b0 , \11447_b1 , \11447_b0 , \11448_b1 , \11448_b0 , \11449_b1 , \11449_b0 , 
		\11450_b1 , \11450_b0 , \11451_b1 , \11451_b0 , \11452_b1 , \11452_b0 , \11453_b1 , \11453_b0 , \11454_b1 , \11454_b0 , 
		\11455_b1 , \11455_b0 , \11456_b1 , \11456_b0 , \11457_b1 , \11457_b0 , \11458_b1 , \11458_b0 , \11459_b1 , \11459_b0 , 
		\11460_b1 , \11460_b0 , \11461_b1 , \11461_b0 , \11462_b1 , \11462_b0 , \11463_b1 , \11463_b0 , \11464_b1 , \11464_b0 , 
		\11465_b1 , \11465_b0 , \11466_b1 , \11466_b0 , \11467_b1 , \11467_b0 , \11468_b1 , \11468_b0 , \11469_b1 , \11469_b0 , 
		\11470_b1 , \11470_b0 , \11471_b1 , \11471_b0 , \11472_b1 , \11472_b0 , \11473_b1 , \11473_b0 , \11474_b1 , \11474_b0 , 
		\11475_b1 , \11475_b0 , \11476_b1 , \11476_b0 , \11477_b1 , \11477_b0 , \11478_b1 , \11478_b0 , \11479_b1 , \11479_b0 , 
		\11480_b1 , \11480_b0 , \11481_b1 , \11481_b0 , \11482_b1 , \11482_b0 , \11483_b1 , \11483_b0 , \11484_b1 , \11484_b0 , 
		\11485_b1 , \11485_b0 , \11486_b1 , \11486_b0 , \11487_b1 , \11487_b0 , \11488_b1 , \11488_b0 , \11489_b1 , \11489_b0 , 
		\11490_b1 , \11490_b0 , \11491_b1 , \11491_b0 , \11492_b1 , \11492_b0 , \11493_b1 , \11493_b0 , \11494_b1 , \11494_b0 , 
		\11495_b1 , \11495_b0 , \11496_b1 , \11496_b0 , \11497_b1 , \11497_b0 , \11498_b1 , \11498_b0 , \11499_b1 , \11499_b0 , 
		\11500_b1 , \11500_b0 , \11501_b1 , \11501_b0 , \11502_b1 , \11502_b0 , \11503_b1 , \11503_b0 , \11504_b1 , \11504_b0 , 
		\11505_b1 , \11505_b0 , \11506_b1 , \11506_b0 , \11507_b1 , \11507_b0 , \11508_b1 , \11508_b0 , \11509_b1 , \11509_b0 , 
		\11510_b1 , \11510_b0 , \11511_b1 , \11511_b0 , \11512_b1 , \11512_b0 , \11513_b1 , \11513_b0 , \11514_b1 , \11514_b0 , 
		\11515_b1 , \11515_b0 , \11516_b1 , \11516_b0 , \11517_b1 , \11517_b0 , \11518_b1 , \11518_b0 , \11519_b1 , \11519_b0 , 
		\11520_b1 , \11520_b0 , \11521_b1 , \11521_b0 , \11522_b1 , \11522_b0 , \11523_b1 , \11523_b0 , \11524_b1 , \11524_b0 , 
		\11525_b1 , \11525_b0 , \11526_b1 , \11526_b0 , \11527_b1 , \11527_b0 , \11528_b1 , \11528_b0 , \11529_b1 , \11529_b0 , 
		\11530_b1 , \11530_b0 , \11531_b1 , \11531_b0 , \11532_b1 , \11532_b0 , \11533_b1 , \11533_b0 , \11534_b1 , \11534_b0 , 
		\11535_b1 , \11535_b0 , \11536_b1 , \11536_b0 , \11537_b1 , \11537_b0 , \11538_b1 , \11538_b0 , \11539_b1 , \11539_b0 , 
		\11540_b1 , \11540_b0 , \11541_b1 , \11541_b0 , \11542_b1 , \11542_b0 , \11543_b1 , \11543_b0 , \11544_b1 , \11544_b0 , 
		\11545_b1 , \11545_b0 , \11546_b1 , \11546_b0 , \11547_b1 , \11547_b0 , \11548_b1 , \11548_b0 , \11549_b1 , \11549_b0 , 
		\11550_b1 , \11550_b0 , \11551_b1 , \11551_b0 , \11552_b1 , \11552_b0 , \11553_b1 , \11553_b0 , \11554_b1 , \11554_b0 , 
		\11555_b1 , \11555_b0 , \11556_b1 , \11556_b0 , \11557_b1 , \11557_b0 , \11558_b1 , \11558_b0 , \11559_b1 , \11559_b0 , 
		\11560_b1 , \11560_b0 , \11561_b1 , \11561_b0 , \11562_b1 , \11562_b0 , \11563_b1 , \11563_b0 , \11564_b1 , \11564_b0 , 
		\11565_b1 , \11565_b0 , \11566_b1 , \11566_b0 , \11567_b1 , \11567_b0 , \11568_b1 , \11568_b0 , \11569_b1 , \11569_b0 , 
		\11570_b1 , \11570_b0 , \11571_b1 , \11571_b0 , \11572_b1 , \11572_b0 , \11573_b1 , \11573_b0 , \11574_b1 , \11574_b0 , 
		\11575_b1 , \11575_b0 , \11576_b1 , \11576_b0 , \11577_b1 , \11577_b0 , \11578_b1 , \11578_b0 , \11579_b1 , \11579_b0 , 
		\11580_b1 , \11580_b0 , \11581_b1 , \11581_b0 , \11582_b1 , \11582_b0 , \11583_b1 , \11583_b0 , \11584_b1 , \11584_b0 , 
		\11585_b1 , \11585_b0 , \11586_b1 , \11586_b0 , \11587_b1 , \11587_b0 , \11588_b1 , \11588_b0 , \11589_b1 , \11589_b0 , 
		\11590_b1 , \11590_b0 , \11591_b1 , \11591_b0 , \11592_b1 , \11592_b0 , \11593_b1 , \11593_b0 , \11594_b1 , \11594_b0 , 
		\11595_b1 , \11595_b0 , \11596_b1 , \11596_b0 , \11597_b1 , \11597_b0 , \11598_b1 , \11598_b0 , \11599_b1 , \11599_b0 , 
		\11600_b1 , \11600_b0 , \11601_b1 , \11601_b0 , \11602_b1 , \11602_b0 , \11603_b1 , \11603_b0 , \11604_b1 , \11604_b0 , 
		\11605_b1 , \11605_b0 , \11606_b1 , \11606_b0 , \11607_b1 , \11607_b0 , \11608_b1 , \11608_b0 , \11609_b1 , \11609_b0 , 
		\11610_b1 , \11610_b0 , \11611_b1 , \11611_b0 , \11612_b1 , \11612_b0 , \11613_b1 , \11613_b0 , \11614_b1 , \11614_b0 , 
		\11615_b1 , \11615_b0 , \11616_b1 , \11616_b0 , \11617_b1 , \11617_b0 , \11618_b1 , \11618_b0 , \11619_b1 , \11619_b0 , 
		\11620_b1 , \11620_b0 , \11621_b1 , \11621_b0 , \11622_b1 , \11622_b0 , \11623_b1 , \11623_b0 , \11624_b1 , \11624_b0 , 
		\11625_b1 , \11625_b0 , \11626_b1 , \11626_b0 , \11627_b1 , \11627_b0 , \11628_b1 , \11628_b0 , \11629_b1 , \11629_b0 , 
		\11630_b1 , \11630_b0 , \11631_b1 , \11631_b0 , \11632_b1 , \11632_b0 , \11633_b1 , \11633_b0 , \11634_b1 , \11634_b0 , 
		\11635_b1 , \11635_b0 , \11636_b1 , \11636_b0 , \11637_b1 , \11637_b0 , \11638_b1 , \11638_b0 , \11639_b1 , \11639_b0 , 
		\11640_b1 , \11640_b0 , \11641_b1 , \11641_b0 , \11642_b1 , \11642_b0 , \11643_b1 , \11643_b0 , \11644_b1 , \11644_b0 , 
		\11645_b1 , \11645_b0 , \11646_b1 , \11646_b0 , \11647_b1 , \11647_b0 , \11648_b1 , \11648_b0 , \11649_b1 , \11649_b0 , 
		\11650_b1 , \11650_b0 , \11651_b1 , \11651_b0 , \11652_b1 , \11652_b0 , \11653_b1 , \11653_b0 , \11654_b1 , \11654_b0 , 
		\11655_b1 , \11655_b0 , \11656_b1 , \11656_b0 , \11657_b1 , \11657_b0 , \11658_b1 , \11658_b0 , \11659_b1 , \11659_b0 , 
		\11660_b1 , \11660_b0 , \11661_b1 , \11661_b0 , \11662_b1 , \11662_b0 , \11663_b1 , \11663_b0 , \11664_b1 , \11664_b0 , 
		\11665_b1 , \11665_b0 , \11666_b1 , \11666_b0 , \11667_b1 , \11667_b0 , \11668_b1 , \11668_b0 , \11669_b1 , \11669_b0 , 
		\11670_b1 , \11670_b0 , \11671_b1 , \11671_b0 , \11672_b1 , \11672_b0 , \11673_b1 , \11673_b0 , \11674_b1 , \11674_b0 , 
		\11675_b1 , \11675_b0 , \11676_b1 , \11676_b0 , \11677_b1 , \11677_b0 , \11678_b1 , \11678_b0 , \11679_b1 , \11679_b0 , 
		\11680_b1 , \11680_b0 , \11681_b1 , \11681_b0 , \11682_b1 , \11682_b0 , \11683_b1 , \11683_b0 , \11684_b1 , \11684_b0 , 
		\11685_b1 , \11685_b0 , \11686_b1 , \11686_b0 , \11687_b1 , \11687_b0 , \11688_b1 , \11688_b0 , \11689_b1 , \11689_b0 , 
		\11690_b1 , \11690_b0 , \11691_b1 , \11691_b0 , \11692_b1 , \11692_b0 , \11693_b1 , \11693_b0 , \11694_b1 , \11694_b0 , 
		\11695_b1 , \11695_b0 , \11696_b1 , \11696_b0 , \11697_b1 , \11697_b0 , \11698_b1 , \11698_b0 , \11699_b1 , \11699_b0 , 
		\11700_b1 , \11700_b0 , \11701_b1 , \11701_b0 , \11702_b1 , \11702_b0 , \11703_b1 , \11703_b0 , \11704_b1 , \11704_b0 , 
		\11705_b1 , \11705_b0 , \11706_b1 , \11706_b0 , \11707_b1 , \11707_b0 , \11708_b1 , \11708_b0 , \11709_b1 , \11709_b0 , 
		\11710_b1 , \11710_b0 , \11711_b1 , \11711_b0 , \11712_b1 , \11712_b0 , \11713_b1 , \11713_b0 , \11714_b1 , \11714_b0 , 
		\11715_b1 , \11715_b0 , \11716_b1 , \11716_b0 , \11717_b1 , \11717_b0 , \11718_b1 , \11718_b0 , \11719_b1 , \11719_b0 , 
		\11720_b1 , \11720_b0 , \11721_b1 , \11721_b0 , \11722_b1 , \11722_b0 , \11723_b1 , \11723_b0 , \11724_b1 , \11724_b0 , 
		\11725_b1 , \11725_b0 , \11726_b1 , \11726_b0 , \11727_b1 , \11727_b0 , \11728_b1 , \11728_b0 , \11729_b1 , \11729_b0 , 
		\11730_b1 , \11730_b0 , \11731_b1 , \11731_b0 , \11732_b1 , \11732_b0 , \11733_b1 , \11733_b0 , \11734_b1 , \11734_b0 , 
		\11735_b1 , \11735_b0 , \11736_b1 , \11736_b0 , \11737_b1 , \11737_b0 , \11738_b1 , \11738_b0 , \11739_b1 , \11739_b0 , 
		\11740_b1 , \11740_b0 , \11741_b1 , \11741_b0 , \11742_b1 , \11742_b0 , \11743_b1 , \11743_b0 , \11744_b1 , \11744_b0 , 
		\11745_b1 , \11745_b0 , \11746_b1 , \11746_b0 , \11747_b1 , \11747_b0 , \11748_b1 , \11748_b0 , \11749_b1 , \11749_b0 , 
		\11750_b1 , \11750_b0 , \11751_b1 , \11751_b0 , \11752_b1 , \11752_b0 , \11753_b1 , \11753_b0 , \11754_b1 , \11754_b0 , 
		\11755_b1 , \11755_b0 , \11756_b1 , \11756_b0 , \11757_b1 , \11757_b0 , \11758_b1 , \11758_b0 , \11759_b1 , \11759_b0 , 
		\11760_b1 , \11760_b0 , \11761_b1 , \11761_b0 , \11762_b1 , \11762_b0 , \11763_b1 , \11763_b0 , \11764_b1 , \11764_b0 , 
		\11765_b1 , \11765_b0 , \11766_b1 , \11766_b0 , \11767_b1 , \11767_b0 , \11768_b1 , \11768_b0 , \11769_b1 , \11769_b0 , 
		\11770_b1 , \11770_b0 , \11771_b1 , \11771_b0 , \11772_b1 , \11772_b0 , \11773_b1 , \11773_b0 , \11774_b1 , \11774_b0 , 
		\11775_b1 , \11775_b0 , \11776_b1 , \11776_b0 , \11777_b1 , \11777_b0 , \11778_b1 , \11778_b0 , \11779_b1 , \11779_b0 , 
		\11780_b1 , \11780_b0 , \11781_b1 , \11781_b0 , \11782_b1 , \11782_b0 , \11783_b1 , \11783_b0 , \11784_b1 , \11784_b0 , 
		\11785_b1 , \11785_b0 , \11786_b1 , \11786_b0 , \11787_b1 , \11787_b0 , \11788_b1 , \11788_b0 , \11789_b1 , \11789_b0 , 
		\11790_b1 , \11790_b0 , \11791_b1 , \11791_b0 , \11792_b1 , \11792_b0 , \11793_b1 , \11793_b0 , \11794_b1 , \11794_b0 , 
		\11795_b1 , \11795_b0 , \11796_b1 , \11796_b0 , \11797_b1 , \11797_b0 , \11798_b1 , \11798_b0 , \11799_b1 , \11799_b0 , 
		\11800_b1 , \11800_b0 , \11801_b1 , \11801_b0 , \11802_b1 , \11802_b0 , \11803_b1 , \11803_b0 , \11804_b1 , \11804_b0 , 
		\11805_b1 , \11805_b0 , \11806_b1 , \11806_b0 , \11807_b1 , \11807_b0 , \11808_b1 , \11808_b0 , \11809_b1 , \11809_b0 , 
		\11810_b1 , \11810_b0 , \11811_b1 , \11811_b0 , \11812_b1 , \11812_b0 , \11813_b1 , \11813_b0 , \11814_b1 , \11814_b0 , 
		\11815_b1 , \11815_b0 , \11816_b1 , \11816_b0 , \11817_b1 , \11817_b0 , \11818_b1 , \11818_b0 , \11819_b1 , \11819_b0 , 
		\11820_b1 , \11820_b0 , \11821_b1 , \11821_b0 , \11822_b1 , \11822_b0 , \11823_b1 , \11823_b0 , \11824_b1 , \11824_b0 , 
		\11825_b1 , \11825_b0 , \11826_b1 , \11826_b0 , \11827_b1 , \11827_b0 , \11828_b1 , \11828_b0 , \11829_b1 , \11829_b0 , 
		\11830_b1 , \11830_b0 , \11831_b1 , \11831_b0 , \11832_b1 , \11832_b0 , \11833_b1 , \11833_b0 , \11834_b1 , \11834_b0 , 
		\11835_b1 , \11835_b0 , \11836_b1 , \11836_b0 , \11837_b1 , \11837_b0 , \11838_b1 , \11838_b0 , \11839_b1 , \11839_b0 , 
		\11840_b1 , \11840_b0 , \11841_b1 , \11841_b0 , \11842_b1 , \11842_b0 , \11843_b1 , \11843_b0 , \11844_b1 , \11844_b0 , 
		\11845_b1 , \11845_b0 , \11846_b1 , \11846_b0 , \11847_b1 , \11847_b0 , \11848_b1 , \11848_b0 , \11849_b1 , \11849_b0 , 
		\11850_b1 , \11850_b0 , \11851_b1 , \11851_b0 , \11852_b1 , \11852_b0 , \11853_b1 , \11853_b0 , \11854_b1 , \11854_b0 , 
		\11855_b1 , \11855_b0 , \11856_b1 , \11856_b0 , \11857_b1 , \11857_b0 , \11858_b1 , \11858_b0 , \11859_b1 , \11859_b0 , 
		\11860_b1 , \11860_b0 , \11861_b1 , \11861_b0 , \11862_b1 , \11862_b0 , \11863_b1 , \11863_b0 , \11864_b1 , \11864_b0 , 
		\11865_b1 , \11865_b0 , \11866_b1 , \11866_b0 , \11867_b1 , \11867_b0 , \11868_b1 , \11868_b0 , \11869_b1 , \11869_b0 , 
		\11870_b1 , \11870_b0 , \11871_b1 , \11871_b0 , \11872_b1 , \11872_b0 , \11873_b1 , \11873_b0 , \11874_b1 , \11874_b0 , 
		\11875_b1 , \11875_b0 , \11876_b1 , \11876_b0 , \11877_b1 , \11877_b0 , \11878_b1 , \11878_b0 , \11879_b1 , \11879_b0 , 
		\11880_b1 , \11880_b0 , \11881_b1 , \11881_b0 , \11882_b1 , \11882_b0 , \11883_b1 , \11883_b0 , \11884_b1 , \11884_b0 , 
		\11885_b1 , \11885_b0 , \11886_b1 , \11886_b0 , \11887_b1 , \11887_b0 , \11888_b1 , \11888_b0 , \11889_b1 , \11889_b0 , 
		\11890_b1 , \11890_b0 , \11891_b1 , \11891_b0 , \11892_b1 , \11892_b0 , \11893_b1 , \11893_b0 , \11894_b1 , \11894_b0 , 
		\11895_b1 , \11895_b0 , \11896_b1 , \11896_b0 , \11897_b1 , \11897_b0 , \11898_b1 , \11898_b0 , \11899_b1 , \11899_b0 , 
		\11900_b1 , \11900_b0 , \11901_b1 , \11901_b0 , \11902_b1 , \11902_b0 , \11903_b1 , \11903_b0 , \11904_b1 , \11904_b0 , 
		\11905_b1 , \11905_b0 , \11906_b1 , \11906_b0 , \11907_b1 , \11907_b0 , \11908_b1 , \11908_b0 , \11909_b1 , \11909_b0 , 
		\11910_b1 , \11910_b0 , \11911_b1 , \11911_b0 , \11912_b1 , \11912_b0 , \11913_b1 , \11913_b0 , \11914_b1 , \11914_b0 , 
		\11915_b1 , \11915_b0 , \11916_b1 , \11916_b0 , \11917_b1 , \11917_b0 , \11918_b1 , \11918_b0 , \11919_b1 , \11919_b0 , 
		\11920_b1 , \11920_b0 , \11921_b1 , \11921_b0 , \11922_b1 , \11922_b0 , \11923_b1 , \11923_b0 , \11924_b1 , \11924_b0 , 
		\11925_b1 , \11925_b0 , \11926_b1 , \11926_b0 , \11927_b1 , \11927_b0 , \11928_b1 , \11928_b0 , \11929_b1 , \11929_b0 , 
		\11930_b1 , \11930_b0 , \11931_b1 , \11931_b0 , \11932_b1 , \11932_b0 , \11933_b1 , \11933_b0 , \11934_b1 , \11934_b0 , 
		\11935_b1 , \11935_b0 , \11936_b1 , \11936_b0 , \11937_b1 , \11937_b0 , \11938_b1 , \11938_b0 , \11939_b1 , \11939_b0 , 
		\11940_b1 , \11940_b0 , \11941_b1 , \11941_b0 , \11942_b1 , \11942_b0 , \11943_b1 , \11943_b0 , \11944_b1 , \11944_b0 , 
		\11945_b1 , \11945_b0 , \11946_b1 , \11946_b0 , \11947_b1 , \11947_b0 , \11948_b1 , \11948_b0 , \11949_b1 , \11949_b0 , 
		\11950_b1 , \11950_b0 , \11951_b1 , \11951_b0 , \11952_b1 , \11952_b0 , \11953_b1 , \11953_b0 , \11954_b1 , \11954_b0 , 
		\11955_b1 , \11955_b0 , \11956_b1 , \11956_b0 , \11957_b1 , \11957_b0 , \11958_b1 , \11958_b0 , \11959_b1 , \11959_b0 , 
		\11960_b1 , \11960_b0 , \11961_b1 , \11961_b0 , \11962_b1 , \11962_b0 , \11963_b1 , \11963_b0 , \11964_b1 , \11964_b0 , 
		\11965_b1 , \11965_b0 , \11966_b1 , \11966_b0 , \11967_b1 , \11967_b0 , \11968_b1 , \11968_b0 , \11969_b1 , \11969_b0 , 
		\11970_b1 , \11970_b0 , \11971_b1 , \11971_b0 , \11972_b1 , \11972_b0 , \11973_b1 , \11973_b0 , \11974_b1 , \11974_b0 , 
		\11975_b1 , \11975_b0 , \11976_b1 , \11976_b0 , \11977_b1 , \11977_b0 , \11978_b1 , \11978_b0 , \11979_b1 , \11979_b0 , 
		\11980_b1 , \11980_b0 , \11981_b1 , \11981_b0 , \11982_b1 , \11982_b0 , \11983_b1 , \11983_b0 , \11984_b1 , \11984_b0 , 
		\11985_b1 , \11985_b0 , \11986_b1 , \11986_b0 , \11987_b1 , \11987_b0 , \11988_b1 , \11988_b0 , \11989_b1 , \11989_b0 , 
		\11990_b1 , \11990_b0 , \11991_b1 , \11991_b0 , \11992_b1 , \11992_b0 , \11993_b1 , \11993_b0 , \11994_b1 , \11994_b0 , 
		\11995_b1 , \11995_b0 , \11996_b1 , \11996_b0 , \11997_b1 , \11997_b0 , \11998_b1 , \11998_b0 , \11999_b1 , \11999_b0 , 
		\12000_b1 , \12000_b0 , \12001_b1 , \12001_b0 , \12002_b1 , \12002_b0 , \12003_b1 , \12003_b0 , \12004_b1 , \12004_b0 , 
		\12005_b1 , \12005_b0 , \12006_b1 , \12006_b0 , \12007_b1 , \12007_b0 , \12008_b1 , \12008_b0 , \12009_b1 , \12009_b0 , 
		\12010_b1 , \12010_b0 , \12011_b1 , \12011_b0 , \12012_b1 , \12012_b0 , \12013_b1 , \12013_b0 , \12014_b1 , \12014_b0 , 
		\12015_b1 , \12015_b0 , \12016_b1 , \12016_b0 , \12017_b1 , \12017_b0 , \12018_b1 , \12018_b0 , \12019_b1 , \12019_b0 , 
		\12020_b1 , \12020_b0 , \12021_b1 , \12021_b0 , \12022_b1 , \12022_b0 , \12023_b1 , \12023_b0 , \12024_b1 , \12024_b0 , 
		\12025_b1 , \12025_b0 , \12026_b1 , \12026_b0 , \12027_b1 , \12027_b0 , \12028_b1 , \12028_b0 , \12029_b1 , \12029_b0 , 
		\12030_b1 , \12030_b0 , \12031_b1 , \12031_b0 , \12032_b1 , \12032_b0 , \12033_b1 , \12033_b0 , \12034_b1 , \12034_b0 , 
		\12035_b1 , \12035_b0 , \12036_b1 , \12036_b0 , \12037_b1 , \12037_b0 , \12038_b1 , \12038_b0 , \12039_b1 , \12039_b0 , 
		\12040_b1 , \12040_b0 , \12041_b1 , \12041_b0 , \12042_b1 , \12042_b0 , \12043_b1 , \12043_b0 , \12044_b1 , \12044_b0 , 
		\12045_b1 , \12045_b0 , \12046_b1 , \12046_b0 , \12047_b1 , \12047_b0 , \12048_b1 , \12048_b0 , \12049_b1 , \12049_b0 , 
		\12050_b1 , \12050_b0 , \12051_b1 , \12051_b0 , \12052_b1 , \12052_b0 , \12053_b1 , \12053_b0 , \12054_b1 , \12054_b0 , 
		\12055_b1 , \12055_b0 , \12056_b1 , \12056_b0 , \12057_b1 , \12057_b0 , \12058_b1 , \12058_b0 , \12059_b1 , \12059_b0 , 
		\12060_b1 , \12060_b0 , \12061_b1 , \12061_b0 , \12062_b1 , \12062_b0 , \12063_b1 , \12063_b0 , \12064_b1 , \12064_b0 , 
		\12065_b1 , \12065_b0 , \12066_b1 , \12066_b0 , \12067_b1 , \12067_b0 , \12068_b1 , \12068_b0 , \12069_b1 , \12069_b0 , 
		\12070_b1 , \12070_b0 , \12071_b1 , \12071_b0 , \12072_b1 , \12072_b0 , \12073_b1 , \12073_b0 , \12074_b1 , \12074_b0 , 
		\12075_b1 , \12075_b0 , \12076_b1 , \12076_b0 , \12077_b1 , \12077_b0 , \12078_b1 , \12078_b0 , \12079_b1 , \12079_b0 , 
		\12080_b1 , \12080_b0 , \12081_b1 , \12081_b0 , \12082_b1 , \12082_b0 , \12083_b1 , \12083_b0 , \12084_b1 , \12084_b0 , 
		\12085_b1 , \12085_b0 , \12086_b1 , \12086_b0 , \12087_b1 , \12087_b0 , \12088_b1 , \12088_b0 , \12089_b1 , \12089_b0 , 
		\12090_b1 , \12090_b0 , \12091_b1 , \12091_b0 , \12092_b1 , \12092_b0 , \12093_b1 , \12093_b0 , \12094_b1 , \12094_b0 , 
		\12095_b1 , \12095_b0 , \12096_b1 , \12096_b0 , \12097_b1 , \12097_b0 , \12098_b1 , \12098_b0 , \12099_b1 , \12099_b0 , 
		\12100_b1 , \12100_b0 , \12101_b1 , \12101_b0 , \12102_b1 , \12102_b0 , \12103_b1 , \12103_b0 , \12104_b1 , \12104_b0 , 
		\12105_b1 , \12105_b0 , \12106_b1 , \12106_b0 , \12107_b1 , \12107_b0 , \12108_b1 , \12108_b0 , \12109_b1 , \12109_b0 , 
		\12110_b1 , \12110_b0 , \12111_b1 , \12111_b0 , \12112_b1 , \12112_b0 , \12113_b1 , \12113_b0 , \12114_b1 , \12114_b0 , 
		\12115_b1 , \12115_b0 , \12116_b1 , \12116_b0 , \12117_b1 , \12117_b0 , \12118_b1 , \12118_b0 , \12119_b1 , \12119_b0 , 
		\12120_b1 , \12120_b0 , \12121_b1 , \12121_b0 , \12122_b1 , \12122_b0 , \12123_b1 , \12123_b0 , \12124_b1 , \12124_b0 , 
		\12125_b1 , \12125_b0 , \12126_b1 , \12126_b0 , \12127_b1 , \12127_b0 , \12128_b1 , \12128_b0 , \12129_b1 , \12129_b0 , 
		\12130_b1 , \12130_b0 , \12131_b1 , \12131_b0 , \12132_b1 , \12132_b0 , \12133_b1 , \12133_b0 , \12134_b1 , \12134_b0 , 
		\12135_b1 , \12135_b0 , \12136_b1 , \12136_b0 , \12137_b1 , \12137_b0 , \12138_b1 , \12138_b0 , \12139_b1 , \12139_b0 , 
		\12140_b1 , \12140_b0 , \12141_b1 , \12141_b0 , \12142_b1 , \12142_b0 , \12143_b1 , \12143_b0 , \12144_b1 , \12144_b0 , 
		\12145_b1 , \12145_b0 , \12146_b1 , \12146_b0 , \12147_b1 , \12147_b0 , \12148_b1 , \12148_b0 , \12149_b1 , \12149_b0 , 
		\12150_b1 , \12150_b0 , \12151_b1 , \12151_b0 , \12152_b1 , \12152_b0 , \12153_b1 , \12153_b0 , \12154_b1 , \12154_b0 , 
		\12155_b1 , \12155_b0 , \12156_b1 , \12156_b0 , \12157_b1 , \12157_b0 , \12158_b1 , \12158_b0 , \12159_b1 , \12159_b0 , 
		\12160_b1 , \12160_b0 , \12161_b1 , \12161_b0 , \12162_b1 , \12162_b0 , \12163_b1 , \12163_b0 , \12164_b1 , \12164_b0 , 
		\12165_b1 , \12165_b0 , \12166_b1 , \12166_b0 , \12167_b1 , \12167_b0 , \12168_b1 , \12168_b0 , \12169_b1 , \12169_b0 , 
		\12170_b1 , \12170_b0 , \12171_b1 , \12171_b0 , \12172_b1 , \12172_b0 , \12173_b1 , \12173_b0 , \12174_b1 , \12174_b0 , 
		\12175_b1 , \12175_b0 , \12176_b1 , \12176_b0 , \12177_b1 , \12177_b0 , \12178_b1 , \12178_b0 , \12179_b1 , \12179_b0 , 
		\12180_b1 , \12180_b0 , \12181_b1 , \12181_b0 , \12182_b1 , \12182_b0 , \12183_b1 , \12183_b0 , \12184_b1 , \12184_b0 , 
		\12185_b1 , \12185_b0 , \12186_b1 , \12186_b0 , \12187_b1 , \12187_b0 , \12188_b1 , \12188_b0 , \12189_b1 , \12189_b0 , 
		\12190_b1 , \12190_b0 , \12191_b1 , \12191_b0 , \12192_b1 , \12192_b0 , \12193_b1 , \12193_b0 , \12194_b1 , \12194_b0 , 
		\12195_b1 , \12195_b0 , \12196_b1 , \12196_b0 , \12197_b1 , \12197_b0 , \12198_b1 , \12198_b0 , \12199_b1 , \12199_b0 , 
		\12200_b1 , \12200_b0 , \12201_b1 , \12201_b0 , \12202_b1 , \12202_b0 , \12203_b1 , \12203_b0 , \12204_b1 , \12204_b0 , 
		\12205_b1 , \12205_b0 , \12206_b1 , \12206_b0 , \12207_b1 , \12207_b0 , \12208_b1 , \12208_b0 , \12209_b1 , \12209_b0 , 
		\12210_b1 , \12210_b0 , \12211_b1 , \12211_b0 , \12212_b1 , \12212_b0 , \12213_b1 , \12213_b0 , \12214_b1 , \12214_b0 , 
		\12215_b1 , \12215_b0 , \12216_b1 , \12216_b0 , \12217_b1 , \12217_b0 , \12218_b1 , \12218_b0 , \12219_b1 , \12219_b0 , 
		\12220_b1 , \12220_b0 , \12221_b1 , \12221_b0 , \12222_b1 , \12222_b0 , \12223_b1 , \12223_b0 , \12224_b1 , \12224_b0 , 
		\12225_b1 , \12225_b0 , \12226_b1 , \12226_b0 , \12227_b1 , \12227_b0 , \12228_b1 , \12228_b0 , \12229_b1 , \12229_b0 , 
		\12230_b1 , \12230_b0 , \12231_b1 , \12231_b0 , \12232_b1 , \12232_b0 , \12233_b1 , \12233_b0 , \12234_b1 , \12234_b0 , 
		\12235_b1 , \12235_b0 , \12236_b1 , \12236_b0 , \12237_b1 , \12237_b0 , \12238_b1 , \12238_b0 , \12239_b1 , \12239_b0 , 
		\12240_b1 , \12240_b0 , \12241_b1 , \12241_b0 , \12242_b1 , \12242_b0 , \12243_b1 , \12243_b0 , \12244_b1 , \12244_b0 , 
		\12245_b1 , \12245_b0 , \12246_b1 , \12246_b0 , \12247_b1 , \12247_b0 , \12248_b1 , \12248_b0 , \12249_b1 , \12249_b0 , 
		\12250_b1 , \12250_b0 , \12251_b1 , \12251_b0 , \12252_b1 , \12252_b0 , \12253_b1 , \12253_b0 , \12254_b1 , \12254_b0 , 
		\12255_b1 , \12255_b0 , \12256_b1 , \12256_b0 , \12257_b1 , \12257_b0 , \12258_b1 , \12258_b0 , \12259_b1 , \12259_b0 , 
		\12260_b1 , \12260_b0 , \12261_b1 , \12261_b0 , \12262_b1 , \12262_b0 , \12263_b1 , \12263_b0 , \12264_b1 , \12264_b0 , 
		\12265_b1 , \12265_b0 , \12266_b1 , \12266_b0 , \12267_b1 , \12267_b0 , \12268_b1 , \12268_b0 , \12269_b1 , \12269_b0 , 
		\12270_b1 , \12270_b0 , \12271_b1 , \12271_b0 , \12272_b1 , \12272_b0 , \12273_b1 , \12273_b0 , \12274_b1 , \12274_b0 , 
		\12275_b1 , \12275_b0 , \12276_b1 , \12276_b0 , \12277_b1 , \12277_b0 , \12278_b1 , \12278_b0 , \12279_b1 , \12279_b0 , 
		\12280_b1 , \12280_b0 , \12281_b1 , \12281_b0 , \12282_b1 , \12282_b0 , \12283_b1 , \12283_b0 , \12284_b1 , \12284_b0 , 
		\12285_b1 , \12285_b0 , \12286_b1 , \12286_b0 , \12287_b1 , \12287_b0 , \12288_b1 , \12288_b0 , \12289_b1 , \12289_b0 , 
		\12290_b1 , \12290_b0 , \12291_b1 , \12291_b0 , \12292_b1 , \12292_b0 , \12293_b1 , \12293_b0 , \12294_b1 , \12294_b0 , 
		\12295_b1 , \12295_b0 , \12296_b1 , \12296_b0 , \12297_b1 , \12297_b0 , \12298_b1 , \12298_b0 , \12299_b1 , \12299_b0 , 
		\12300_b1 , \12300_b0 , \12301_b1 , \12301_b0 , \12302_b1 , \12302_b0 , \12303_b1 , \12303_b0 , \12304_b1 , \12304_b0 , 
		\12305_b1 , \12305_b0 , \12306_b1 , \12306_b0 , \12307_b1 , \12307_b0 , \12308_b1 , \12308_b0 , \12309_b1 , \12309_b0 , 
		\12310_b1 , \12310_b0 , \12311_b1 , \12311_b0 , \12312_b1 , \12312_b0 , \12313_b1 , \12313_b0 , \12314_b1 , \12314_b0 , 
		\12315_b1 , \12315_b0 , \12316_b1 , \12316_b0 , \12317_b1 , \12317_b0 , \12318_b1 , \12318_b0 , \12319_b1 , \12319_b0 , 
		\12320_b1 , \12320_b0 , \12321_b1 , \12321_b0 , \12322_b1 , \12322_b0 , \12323_b1 , \12323_b0 , \12324_b1 , \12324_b0 , 
		\12325_b1 , \12325_b0 , \12326_b1 , \12326_b0 , \12327_b1 , \12327_b0 , \12328_b1 , \12328_b0 , \12329_b1 , \12329_b0 , 
		\12330_b1 , \12330_b0 , \12331_b1 , \12331_b0 , \12332_b1 , \12332_b0 , \12333_b1 , \12333_b0 , \12334_b1 , \12334_b0 , 
		\12335_b1 , \12335_b0 , \12336_b1 , \12336_b0 , \12337_b1 , \12337_b0 , \12338_b1 , \12338_b0 , \12339_b1 , \12339_b0 , 
		\12340_b1 , \12340_b0 , \12341_b1 , \12341_b0 , \12342_b1 , \12342_b0 , \12343_b1 , \12343_b0 , \12344_b1 , \12344_b0 , 
		\12345_b1 , \12345_b0 , \12346_b1 , \12346_b0 , \12347_b1 , \12347_b0 , \12348_b1 , \12348_b0 , \12349_b1 , \12349_b0 , 
		\12350_b1 , \12350_b0 , \12351_b1 , \12351_b0 , \12352_b1 , \12352_b0 , \12353_b1 , \12353_b0 , \12354_b1 , \12354_b0 , 
		\12355_b1 , \12355_b0 , \12356_b1 , \12356_b0 , \12357_b1 , \12357_b0 , \12358_b1 , \12358_b0 , \12359_b1 , \12359_b0 , 
		\12360_b1 , \12360_b0 , \12361_b1 , \12361_b0 , \12362_b1 , \12362_b0 , \12363_b1 , \12363_b0 , \12364_b1 , \12364_b0 , 
		\12365_b1 , \12365_b0 , \12366_b1 , \12366_b0 , \12367_b1 , \12367_b0 , \12368_b1 , \12368_b0 , \12369_b1 , \12369_b0 , 
		\12370_b1 , \12370_b0 , \12371_b1 , \12371_b0 , \12372_b1 , \12372_b0 , \12373_b1 , \12373_b0 , \12374_b1 , \12374_b0 , 
		\12375_b1 , \12375_b0 , \12376_b1 , \12376_b0 , \12377_b1 , \12377_b0 , \12378_b1 , \12378_b0 , \12379_b1 , \12379_b0 , 
		\12380_b1 , \12380_b0 , \12381_b1 , \12381_b0 , \12382_b1 , \12382_b0 , \12383_b1 , \12383_b0 , \12384_b1 , \12384_b0 , 
		\12385_b1 , \12385_b0 , \12386_b1 , \12386_b0 , \12387_b1 , \12387_b0 , \12388_b1 , \12388_b0 , \12389_b1 , \12389_b0 , 
		\12390_b1 , \12390_b0 , \12391_b1 , \12391_b0 , \12392_b1 , \12392_b0 , \12393_b1 , \12393_b0 , \12394_b1 , \12394_b0 , 
		\12395_b1 , \12395_b0 , \12396_b1 , \12396_b0 , \12397_b1 , \12397_b0 , \12398_b1 , \12398_b0 , \12399_b1 , \12399_b0 , 
		\12400_b1 , \12400_b0 , \12401_b1 , \12401_b0 , \12402_b1 , \12402_b0 , \12403_b1 , \12403_b0 , \12404_b1 , \12404_b0 , 
		\12405_b1 , \12405_b0 , \12406_b1 , \12406_b0 , \12407_b1 , \12407_b0 , \12408_b1 , \12408_b0 , \12409_b1 , \12409_b0 , 
		\12410_b1 , \12410_b0 , \12411_b1 , \12411_b0 , \12412_b1 , \12412_b0 , \12413_b1 , \12413_b0 , \12414_b1 , \12414_b0 , 
		\12415_b1 , \12415_b0 , \12416_b1 , \12416_b0 , \12417_b1 , \12417_b0 , \12418_b1 , \12418_b0 , \12419_b1 , \12419_b0 , 
		\12420_b1 , \12420_b0 , \12421_b1 , \12421_b0 , \12422_b1 , \12422_b0 , \12423_b1 , \12423_b0 , \12424_b1 , \12424_b0 , 
		\12425_b1 , \12425_b0 , \12426_b1 , \12426_b0 , \12427_b1 , \12427_b0 , \12428_b1 , \12428_b0 , \12429_b1 , \12429_b0 , 
		\12430_b1 , \12430_b0 , \12431_b1 , \12431_b0 , \12432_b1 , \12432_b0 , \12433_b1 , \12433_b0 , \12434_b1 , \12434_b0 , 
		\12435_b1 , \12435_b0 , \12436_b1 , \12436_b0 , \12437_b1 , \12437_b0 , \12438_b1 , \12438_b0 , \12439_b1 , \12439_b0 , 
		\12440_b1 , \12440_b0 , \12441_b1 , \12441_b0 , \12442_b1 , \12442_b0 , \12443_b1 , \12443_b0 , \12444_b1 , \12444_b0 , 
		\12445_b1 , \12445_b0 , \12446_b1 , \12446_b0 , \12447_b1 , \12447_b0 , \12448_b1 , \12448_b0 , \12449_b1 , \12449_b0 , 
		\12450_b1 , \12450_b0 , \12451_b1 , \12451_b0 , \12452_b1 , \12452_b0 , \12453_b1 , \12453_b0 , \12454_b1 , \12454_b0 , 
		\12455_b1 , \12455_b0 , \12456_b1 , \12456_b0 , \12457_b1 , \12457_b0 , \12458_b1 , \12458_b0 , \12459_b1 , \12459_b0 , 
		\12460_b1 , \12460_b0 , \12461_b1 , \12461_b0 , \12462_b1 , \12462_b0 , \12463_b1 , \12463_b0 , \12464_b1 , \12464_b0 , 
		\12465_b1 , \12465_b0 , \12466_b1 , \12466_b0 , \12467_b1 , \12467_b0 , \12468_b1 , \12468_b0 , \12469_b1 , \12469_b0 , 
		\12470_b1 , \12470_b0 , \12471_b1 , \12471_b0 , \12472_b1 , \12472_b0 , \12473_b1 , \12473_b0 , \12474_b1 , \12474_b0 , 
		\12475_b1 , \12475_b0 , \12476_b1 , \12476_b0 , \12477_b1 , \12477_b0 , \12478_b1 , \12478_b0 , \12479_b1 , \12479_b0 , 
		\12480_b1 , \12480_b0 , \12481_b1 , \12481_b0 , \12482_b1 , \12482_b0 , \12483_b1 , \12483_b0 , \12484_b1 , \12484_b0 , 
		\12485_b1 , \12485_b0 , \12486_b1 , \12486_b0 , \12487_b1 , \12487_b0 , \12488_b1 , \12488_b0 , \12489_b1 , \12489_b0 , 
		\12490_b1 , \12490_b0 , \12491_b1 , \12491_b0 , \12492_b1 , \12492_b0 , \12493_b1 , \12493_b0 , \12494_b1 , \12494_b0 , 
		\12495_b1 , \12495_b0 , \12496_b1 , \12496_b0 , \12497_b1 , \12497_b0 , \12498_b1 , \12498_b0 , \12499_b1 , \12499_b0 , 
		\12500_b1 , \12500_b0 , \12501_b1 , \12501_b0 , \12502_b1 , \12502_b0 , \12503_b1 , \12503_b0 , \12504_b1 , \12504_b0 , 
		\12505_b1 , \12505_b0 , \12506_b1 , \12506_b0 , \12507_b1 , \12507_b0 , \12508_b1 , \12508_b0 , \12509_b1 , \12509_b0 , 
		\12510_b1 , \12510_b0 , \12511_b1 , \12511_b0 , \12512_b1 , \12512_b0 , \12513_b1 , \12513_b0 , \12514_b1 , \12514_b0 , 
		\12515_b1 , \12515_b0 , \12516_b1 , \12516_b0 , \12517_b1 , \12517_b0 , \12518_b1 , \12518_b0 , \12519_b1 , \12519_b0 , 
		\12520_b1 , \12520_b0 , \12521_b1 , \12521_b0 , \12522_b1 , \12522_b0 , \12523_b1 , \12523_b0 , \12524_b1 , \12524_b0 , 
		\12525_b1 , \12525_b0 , \12526_b1 , \12526_b0 , \12527_b1 , \12527_b0 , \12528_b1 , \12528_b0 , \12529_b1 , \12529_b0 , 
		\12530_b1 , \12530_b0 , \12531_b1 , \12531_b0 , \12532_b1 , \12532_b0 , \12533_b1 , \12533_b0 , \12534_b1 , \12534_b0 , 
		\12535_b1 , \12535_b0 , \12536_b1 , \12536_b0 , \12537_b1 , \12537_b0 , \12538_b1 , \12538_b0 , \12539_b1 , \12539_b0 , 
		\12540_b1 , \12540_b0 , \12541_b1 , \12541_b0 , \12542_b1 , \12542_b0 , \12543_b1 , \12543_b0 , \12544_b1 , \12544_b0 , 
		\12545_b1 , \12545_b0 , \12546_b1 , \12546_b0 , \12547_b1 , \12547_b0 , \12548_b1 , \12548_b0 , \12549_b1 , \12549_b0 , 
		\12550_b1 , \12550_b0 , \12551_b1 , \12551_b0 , \12552_b1 , \12552_b0 , \12553_b1 , \12553_b0 , \12554_b1 , \12554_b0 , 
		\12555_b1 , \12555_b0 , \12556_b1 , \12556_b0 , \12557_b1 , \12557_b0 , \12558_b1 , \12558_b0 , \12559_b1 , \12559_b0 , 
		\12560_b1 , \12560_b0 , \12561_b1 , \12561_b0 , \12562_b1 , \12562_b0 , \12563_b1 , \12563_b0 , \12564_b1 , \12564_b0 , 
		\12565_b1 , \12565_b0 , \12566_b1 , \12566_b0 , \12567_b1 , \12567_b0 , \12568_b1 , \12568_b0 , \12569_b1 , \12569_b0 , 
		\12570_b1 , \12570_b0 , \12571_b1 , \12571_b0 , \12572_b1 , \12572_b0 , \12573_b1 , \12573_b0 , \12574_b1 , \12574_b0 , 
		\12575_b1 , \12575_b0 , \12576_b1 , \12576_b0 , \12577_b1 , \12577_b0 , \12578_b1 , \12578_b0 , \12579_b1 , \12579_b0 , 
		\12580_b1 , \12580_b0 , \12581_b1 , \12581_b0 , \12582_b1 , \12582_b0 , \12583_b1 , \12583_b0 , \12584_b1 , \12584_b0 , 
		\12585_b1 , \12585_b0 , \12586_b1 , \12586_b0 , \12587_b1 , \12587_b0 , \12588_b1 , \12588_b0 , \12589_b1 , \12589_b0 , 
		\12590_b1 , \12590_b0 , \12591_b1 , \12591_b0 , \12592_b1 , \12592_b0 , \12593_b1 , \12593_b0 , \12594_b1 , \12594_b0 , 
		\12595_b1 , \12595_b0 , \12596_b1 , \12596_b0 , \12597_b1 , \12597_b0 , \12598_b1 , \12598_b0 , \12599_b1 , \12599_b0 , 
		\12600_b1 , \12600_b0 , \12601_b1 , \12601_b0 , \12602_b1 , \12602_b0 , \12603_b1 , \12603_b0 , \12604_b1 , \12604_b0 , 
		\12605_b1 , \12605_b0 , \12606_b1 , \12606_b0 , \12607_b1 , \12607_b0 , \12608_b1 , \12608_b0 , \12609_b1 , \12609_b0 , 
		\12610_b1 , \12610_b0 , \12611_b1 , \12611_b0 , \12612_b1 , \12612_b0 , \12613_b1 , \12613_b0 , \12614_b1 , \12614_b0 , 
		\12615_b1 , \12615_b0 , \12616_b1 , \12616_b0 , \12617_b1 , \12617_b0 , \12618_b1 , \12618_b0 , \12619_b1 , \12619_b0 , 
		\12620_b1 , \12620_b0 , \12621_b1 , \12621_b0 , \12622_b1 , \12622_b0 , \12623_b1 , \12623_b0 , \12624_b1 , \12624_b0 , 
		\12625_b1 , \12625_b0 , \12626_b1 , \12626_b0 , \12627_b1 , \12627_b0 , \12628_b1 , \12628_b0 , \12629_b1 , \12629_b0 , 
		\12630_b1 , \12630_b0 , \12631_b1 , \12631_b0 , \12632_b1 , \12632_b0 , \12633_b1 , \12633_b0 , \12634_b1 , \12634_b0 , 
		\12635_b1 , \12635_b0 , \12636_b1 , \12636_b0 , \12637_b1 , \12637_b0 , \12638_b1 , \12638_b0 , \12639_b1 , \12639_b0 , 
		\12640_b1 , \12640_b0 , \12641_b1 , \12641_b0 , \12642_b1 , \12642_b0 , \12643_b1 , \12643_b0 , \12644_b1 , \12644_b0 , 
		\12645_b1 , \12645_b0 , \12646_b1 , \12646_b0 , \12647_b1 , \12647_b0 , \12648_b1 , \12648_b0 , \12649_b1 , \12649_b0 , 
		\12650_b1 , \12650_b0 , \12651_b1 , \12651_b0 , \12652_b1 , \12652_b0 , \12653_b1 , \12653_b0 , \12654_b1 , \12654_b0 , 
		\12655_b1 , \12655_b0 , \12656_b1 , \12656_b0 , \12657_b1 , \12657_b0 , \12658_b1 , \12658_b0 , \12659_b1 , \12659_b0 , 
		\12660_b1 , \12660_b0 , \12661_b1 , \12661_b0 , \12662_b1 , \12662_b0 , \12663_b1 , \12663_b0 , \12664_b1 , \12664_b0 , 
		\12665_b1 , \12665_b0 , \12666_b1 , \12666_b0 , \12667_b1 , \12667_b0 , \12668_b1 , \12668_b0 , \12669_b1 , \12669_b0 , 
		\12670_b1 , \12670_b0 , \12671_b1 , \12671_b0 , \12672_b1 , \12672_b0 , \12673_b1 , \12673_b0 , \12674_b1 , \12674_b0 , 
		\12675_b1 , \12675_b0 , \12676_b1 , \12676_b0 , \12677_b1 , \12677_b0 , \12678_b1 , \12678_b0 , \12679_b1 , \12679_b0 , 
		\12680_b1 , \12680_b0 , \12681_b1 , \12681_b0 , \12682_b1 , \12682_b0 , \12683_b1 , \12683_b0 , \12684_b1 , \12684_b0 , 
		\12685_b1 , \12685_b0 , \12686_b1 , \12686_b0 , \12687_b1 , \12687_b0 , \12688_b1 , \12688_b0 , \12689_b1 , \12689_b0 , 
		\12690_b1 , \12690_b0 , \12691_b1 , \12691_b0 , \12692_b1 , \12692_b0 , \12693_b1 , \12693_b0 , \12694_b1 , \12694_b0 , 
		\12695_b1 , \12695_b0 , \12696_b1 , \12696_b0 , \12697_b1 , \12697_b0 , \12698_b1 , \12698_b0 , \12699_b1 , \12699_b0 , 
		\12700_b1 , \12700_b0 , \12701_b1 , \12701_b0 , \12702_b1 , \12702_b0 , \12703_b1 , \12703_b0 , \12704_b1 , \12704_b0 , 
		\12705_b1 , \12705_b0 , \12706_b1 , \12706_b0 , \12707_b1 , \12707_b0 , \12708_b1 , \12708_b0 , \12709_b1 , \12709_b0 , 
		\12710_b1 , \12710_b0 , \12711_b1 , \12711_b0 , \12712_b1 , \12712_b0 , \12713_b1 , \12713_b0 , \12714_b1 , \12714_b0 , 
		\12715_b1 , \12715_b0 , \12716_b1 , \12716_b0 , \12717_b1 , \12717_b0 , \12718_b1 , \12718_b0 , \12719_b1 , \12719_b0 , 
		\12720_b1 , \12720_b0 , \12721_b1 , \12721_b0 , \12722_b1 , \12722_b0 , \12723_b1 , \12723_b0 , \12724_b1 , \12724_b0 , 
		\12725_b1 , \12725_b0 , \12726_b1 , \12726_b0 , \12727_b1 , \12727_b0 , \12728_b1 , \12728_b0 , \12729_b1 , \12729_b0 , 
		\12730_b1 , \12730_b0 , \12731_b1 , \12731_b0 , \12732_b1 , \12732_b0 , \12733_b1 , \12733_b0 , \12734_b1 , \12734_b0 , 
		\12735_b1 , \12735_b0 , \12736_b1 , \12736_b0 , \12737_b1 , \12737_b0 , \12738_b1 , \12738_b0 , \12739_b1 , \12739_b0 , 
		\12740_b1 , \12740_b0 , \12741_b1 , \12741_b0 , \12742_b1 , \12742_b0 , \12743_b1 , \12743_b0 , \12744_b1 , \12744_b0 , 
		\12745_b1 , \12745_b0 , \12746_b1 , \12746_b0 , \12747_b1 , \12747_b0 , \12748_b1 , \12748_b0 , \12749_b1 , \12749_b0 , 
		\12750_b1 , \12750_b0 , \12751_b1 , \12751_b0 , \12752_b1 , \12752_b0 , \12753_b1 , \12753_b0 , \12754_b1 , \12754_b0 , 
		\12755_b1 , \12755_b0 , \12756_b1 , \12756_b0 , \12757_b1 , \12757_b0 , \12758_b1 , \12758_b0 , \12759_b1 , \12759_b0 , 
		\12760_b1 , \12760_b0 , \12761_b1 , \12761_b0 , \12762_b1 , \12762_b0 , \12763_b1 , \12763_b0 , \12764_b1 , \12764_b0 , 
		\12765_b1 , \12765_b0 , \12766_b1 , \12766_b0 , \12767_b1 , \12767_b0 , \12768_b1 , \12768_b0 , \12769_b1 , \12769_b0 , 
		\12770_b1 , \12770_b0 , \12771_b1 , \12771_b0 , \12772_b1 , \12772_b0 , \12773_b1 , \12773_b0 , \12774_b1 , \12774_b0 , 
		\12775_b1 , \12775_b0 , \12776_b1 , \12776_b0 , \12777_b1 , \12777_b0 , \12778_b1 , \12778_b0 , \12779_b1 , \12779_b0 , 
		\12780_b1 , \12780_b0 , \12781_b1 , \12781_b0 , \12782_b1 , \12782_b0 , \12783_b1 , \12783_b0 , \12784_b1 , \12784_b0 , 
		\12785_b1 , \12785_b0 , \12786_b1 , \12786_b0 , \12787_b1 , \12787_b0 , \12788_b1 , \12788_b0 , \12789_b1 , \12789_b0 , 
		\12790_b1 , \12790_b0 , \12791_b1 , \12791_b0 , \12792_b1 , \12792_b0 , \12793_b1 , \12793_b0 , \12794_b1 , \12794_b0 , 
		\12795_b1 , \12795_b0 , \12796_b1 , \12796_b0 , \12797_b1 , \12797_b0 , \12798_b1 , \12798_b0 , \12799_b1 , \12799_b0 , 
		\12800_b1 , \12800_b0 , \12801_b1 , \12801_b0 , \12802_b1 , \12802_b0 , \12803_b1 , \12803_b0 , \12804_b1 , \12804_b0 , 
		\12805_b1 , \12805_b0 , \12806_b1 , \12806_b0 , \12807_b1 , \12807_b0 , \12808_b1 , \12808_b0 , \12809_b1 , \12809_b0 , 
		\12810_b1 , \12810_b0 , \12811_b1 , \12811_b0 , \12812_b1 , \12812_b0 , \12813_b1 , \12813_b0 , \12814_b1 , \12814_b0 , 
		\12815_b1 , \12815_b0 , \12816_b1 , \12816_b0 , \12817_b1 , \12817_b0 , \12818_b1 , \12818_b0 , \12819_b1 , \12819_b0 , 
		\12820_b1 , \12820_b0 , \12821_b1 , \12821_b0 , \12822_b1 , \12822_b0 , \12823_b1 , \12823_b0 , \12824_b1 , \12824_b0 , 
		\12825_b1 , \12825_b0 , \12826_b1 , \12826_b0 , \12827_b1 , \12827_b0 , \12828_b1 , \12828_b0 , \12829_b1 , \12829_b0 , 
		\12830_b1 , \12830_b0 , \12831_b1 , \12831_b0 , \12832_b1 , \12832_b0 , \12833_b1 , \12833_b0 , \12834_b1 , \12834_b0 , 
		\12835_b1 , \12835_b0 , \12836_b1 , \12836_b0 , \12837_b1 , \12837_b0 , \12838_b1 , \12838_b0 , \12839_b1 , \12839_b0 , 
		\12840_b1 , \12840_b0 , \12841_b1 , \12841_b0 , \12842_b1 , \12842_b0 , \12843_b1 , \12843_b0 , \12844_b1 , \12844_b0 , 
		\12845_b1 , \12845_b0 , \12846_b1 , \12846_b0 , \12847_b1 , \12847_b0 , \12848_b1 , \12848_b0 , \12849_b1 , \12849_b0 , 
		\12850_b1 , \12850_b0 , \12851_b1 , \12851_b0 , \12852_b1 , \12852_b0 , \12853_b1 , \12853_b0 , \12854_b1 , \12854_b0 , 
		\12855_b1 , \12855_b0 , \12856_b1 , \12856_b0 , \12857_b1 , \12857_b0 , \12858_b1 , \12858_b0 , \12859_b1 , \12859_b0 , 
		\12860_b1 , \12860_b0 , \12861_b1 , \12861_b0 , \12862_b1 , \12862_b0 , \12863_b1 , \12863_b0 , \12864_b1 , \12864_b0 , 
		\12865_b1 , \12865_b0 , \12866_b1 , \12866_b0 , \12867_b1 , \12867_b0 , \12868_b1 , \12868_b0 , \12869_b1 , \12869_b0 , 
		\12870_b1 , \12870_b0 , \12871_b1 , \12871_b0 , \12872_b1 , \12872_b0 , \12873_b1 , \12873_b0 , \12874_b1 , \12874_b0 , 
		\12875_b1 , \12875_b0 , \12876_b1 , \12876_b0 , \12877_b1 , \12877_b0 , \12878_b1 , \12878_b0 , \12879_b1 , \12879_b0 , 
		\12880_b1 , \12880_b0 , \12881_b1 , \12881_b0 , \12882_b1 , \12882_b0 , \12883_b1 , \12883_b0 , \12884_b1 , \12884_b0 , 
		\12885_b1 , \12885_b0 , \12886_b1 , \12886_b0 , \12887_b1 , \12887_b0 , \12888_b1 , \12888_b0 , \12889_b1 , \12889_b0 , 
		\12890_b1 , \12890_b0 , \12891_b1 , \12891_b0 , \12892_b1 , \12892_b0 , \12893_b1 , \12893_b0 , \12894_b1 , \12894_b0 , 
		\12895_b1 , \12895_b0 , \12896_b1 , \12896_b0 , \12897_b1 , \12897_b0 , \12898_b1 , \12898_b0 , \12899_b1 , \12899_b0 , 
		\12900_b1 , \12900_b0 , \12901_b1 , \12901_b0 , \12902_b1 , \12902_b0 , \12903_b1 , \12903_b0 , \12904_b1 , \12904_b0 , 
		\12905_b1 , \12905_b0 , \12906_b1 , \12906_b0 , \12907_b1 , \12907_b0 , \12908_b1 , \12908_b0 , \12909_b1 , \12909_b0 , 
		\12910_b1 , \12910_b0 , \12911_b1 , \12911_b0 , \12912_b1 , \12912_b0 , \12913_b1 , \12913_b0 , \12914_b1 , \12914_b0 , 
		\12915_b1 , \12915_b0 , \12916_b1 , \12916_b0 , \12917_b1 , \12917_b0 , \12918_b1 , \12918_b0 , \12919_b1 , \12919_b0 , 
		\12920_b1 , \12920_b0 , \12921_b1 , \12921_b0 , \12922_b1 , \12922_b0 , \12923_b1 , \12923_b0 , \12924_b1 , \12924_b0 , 
		\12925_b1 , \12925_b0 , \12926_b1 , \12926_b0 , \12927_b1 , \12927_b0 , \12928_b1 , \12928_b0 , \12929_b1 , \12929_b0 , 
		\12930_b1 , \12930_b0 , \12931_b1 , \12931_b0 , \12932_b1 , \12932_b0 , \12933_b1 , \12933_b0 , \12934_b1 , \12934_b0 , 
		\12935_b1 , \12935_b0 , \12936_b1 , \12936_b0 , \12937_b1 , \12937_b0 , \12938_b1 , \12938_b0 , \12939_b1 , \12939_b0 , 
		\12940_b1 , \12940_b0 , \12941_b1 , \12941_b0 , \12942_b1 , \12942_b0 , \12943_b1 , \12943_b0 , \12944_b1 , \12944_b0 , 
		\12945_b1 , \12945_b0 , \12946_b1 , \12946_b0 , \12947_b1 , \12947_b0 , \12948_b1 , \12948_b0 , \12949_b1 , \12949_b0 , 
		\12950_b1 , \12950_b0 , \12951_b1 , \12951_b0 , \12952_b1 , \12952_b0 , \12953_b1 , \12953_b0 , \12954_b1 , \12954_b0 , 
		\12955_b1 , \12955_b0 , \12956_b1 , \12956_b0 , \12957_b1 , \12957_b0 , \12958_b1 , \12958_b0 , \12959_b1 , \12959_b0 , 
		\12960_b1 , \12960_b0 , \12961_b1 , \12961_b0 , \12962_b1 , \12962_b0 , \12963_b1 , \12963_b0 , \12964_b1 , \12964_b0 , 
		\12965_b1 , \12965_b0 , \12966_b1 , \12966_b0 , \12967_b1 , \12967_b0 , \12968_b1 , \12968_b0 , \12969_b1 , \12969_b0 , 
		\12970_b1 , \12970_b0 , \12971_b1 , \12971_b0 , \12972_b1 , \12972_b0 , \12973_b1 , \12973_b0 , \12974_b1 , \12974_b0 , 
		\12975_b1 , \12975_b0 , \12976_b1 , \12976_b0 , \12977_b1 , \12977_b0 , \12978_b1 , \12978_b0 , \12979_b1 , \12979_b0 , 
		\12980_b1 , \12980_b0 , \12981_b1 , \12981_b0 , \12982_b1 , \12982_b0 , \12983_b1 , \12983_b0 , \12984_b1 , \12984_b0 , 
		\12985_b1 , \12985_b0 , \12986_b1 , \12986_b0 , \12987_b1 , \12987_b0 , \12988_b1 , \12988_b0 , \12989_b1 , \12989_b0 , 
		\12990_b1 , \12990_b0 , \12991_b1 , \12991_b0 , \12992_b1 , \12992_b0 , \12993_b1 , \12993_b0 , \12994_b1 , \12994_b0 , 
		\12995_b1 , \12995_b0 , \12996_b1 , \12996_b0 , \12997_b1 , \12997_b0 , \12998_b1 , \12998_b0 , \12999_b1 , \12999_b0 , 
		\13000_b1 , \13000_b0 , \13001_b1 , \13001_b0 , \13002_b1 , \13002_b0 , \13003_b1 , \13003_b0 , \13004_b1 , \13004_b0 , 
		\13005_b1 , \13005_b0 , \13006_b1 , \13006_b0 , \13007_b1 , \13007_b0 , \13008_b1 , \13008_b0 , \13009_b1 , \13009_b0 , 
		\13010_b1 , \13010_b0 , \13011_b1 , \13011_b0 , \13012_b1 , \13012_b0 , \13013_b1 , \13013_b0 , \13014_b1 , \13014_b0 , 
		\13015_b1 , \13015_b0 , \13016_b1 , \13016_b0 , \13017_b1 , \13017_b0 , \13018_b1 , \13018_b0 , \13019_b1 , \13019_b0 , 
		\13020_b1 , \13020_b0 , \13021_b1 , \13021_b0 , \13022_b1 , \13022_b0 , \13023_b1 , \13023_b0 , \13024_b1 , \13024_b0 , 
		\13025_b1 , \13025_b0 , \13026_b1 , \13026_b0 , \13027_b1 , \13027_b0 , \13028_b1 , \13028_b0 , \13029_b1 , \13029_b0 , 
		\13030_b1 , \13030_b0 , \13031_b1 , \13031_b0 , \13032_b1 , \13032_b0 , \13033_b1 , \13033_b0 , \13034_b1 , \13034_b0 , 
		\13035_b1 , \13035_b0 , \13036_b1 , \13036_b0 , \13037_b1 , \13037_b0 , \13038_b1 , \13038_b0 , \13039_b1 , \13039_b0 , 
		\13040_b1 , \13040_b0 , \13041_b1 , \13041_b0 , \13042_b1 , \13042_b0 , \13043_b1 , \13043_b0 , \13044_b1 , \13044_b0 , 
		\13045_b1 , \13045_b0 , \13046_b1 , \13046_b0 , \13047_b1 , \13047_b0 , \13048_b1 , \13048_b0 , \13049_b1 , \13049_b0 , 
		\13050_b1 , \13050_b0 , \13051_b1 , \13051_b0 , \13052_b1 , \13052_b0 , \13053_b1 , \13053_b0 , \13054_b1 , \13054_b0 , 
		\13055_b1 , \13055_b0 , \13056_b1 , \13056_b0 , \13057_b1 , \13057_b0 , \13058_b1 , \13058_b0 , \13059_b1 , \13059_b0 , 
		\13060_b1 , \13060_b0 , \13061_b1 , \13061_b0 , \13062_b1 , \13062_b0 , \13063_b1 , \13063_b0 , \13064_b1 , \13064_b0 , 
		\13065_b1 , \13065_b0 , \13066_b1 , \13066_b0 , \13067_b1 , \13067_b0 , \13068_b1 , \13068_b0 , \13069_b1 , \13069_b0 , 
		\13070_b1 , \13070_b0 , \13071_b1 , \13071_b0 , \13072_b1 , \13072_b0 , \13073_b1 , \13073_b0 , \13074_b1 , \13074_b0 , 
		\13075_b1 , \13075_b0 , \13076_b1 , \13076_b0 , \13077_b1 , \13077_b0 , \13078_b1 , \13078_b0 , \13079_b1 , \13079_b0 , 
		\13080_b1 , \13080_b0 , \13081_b1 , \13081_b0 , \13082_b1 , \13082_b0 , \13083_b1 , \13083_b0 , \13084_b1 , \13084_b0 , 
		\13085_b1 , \13085_b0 , \13086_b1 , \13086_b0 , \13087_b1 , \13087_b0 , \13088_b1 , \13088_b0 , \13089_b1 , \13089_b0 , 
		\13090_b1 , \13090_b0 , \13091_b1 , \13091_b0 , \13092_b1 , \13092_b0 , \13093_b1 , \13093_b0 , \13094_b1 , \13094_b0 , 
		\13095_b1 , \13095_b0 , \13096_b1 , \13096_b0 , \13097_b1 , \13097_b0 , \13098_b1 , \13098_b0 , \13099_b1 , \13099_b0 , 
		\13100_b1 , \13100_b0 , \13101_b1 , \13101_b0 , \13102_b1 , \13102_b0 , \13103_b1 , \13103_b0 , \13104_b1 , \13104_b0 , 
		\13105_b1 , \13105_b0 , \13106_b1 , \13106_b0 , \13107_b1 , \13107_b0 , \13108_b1 , \13108_b0 , \13109_b1 , \13109_b0 , 
		\13110_b1 , \13110_b0 , \13111_b1 , \13111_b0 , \13112_b1 , \13112_b0 , \13113_b1 , \13113_b0 , \13114_b1 , \13114_b0 , 
		\13115_b1 , \13115_b0 , \13116_b1 , \13116_b0 , \13117_b1 , \13117_b0 , \13118_b1 , \13118_b0 , \13119_b1 , \13119_b0 , 
		\13120_b1 , \13120_b0 , \13121_b1 , \13121_b0 , \13122_b1 , \13122_b0 , \13123_b1 , \13123_b0 , \13124_b1 , \13124_b0 , 
		\13125_b1 , \13125_b0 , \13126_b1 , \13126_b0 , \13127_b1 , \13127_b0 , \13128_b1 , \13128_b0 , \13129_b1 , \13129_b0 , 
		\13130_b1 , \13130_b0 , \13131_b1 , \13131_b0 , \13132_b1 , \13132_b0 , \13133_b1 , \13133_b0 , \13134_b1 , \13134_b0 , 
		\13135_b1 , \13135_b0 , \13136_b1 , \13136_b0 , \13137_b1 , \13137_b0 , \13138_b1 , \13138_b0 , \13139_b1 , \13139_b0 , 
		\13140_b1 , \13140_b0 , \13141_b1 , \13141_b0 , \13142_b1 , \13142_b0 , \13143_b1 , \13143_b0 , \13144_b1 , \13144_b0 , 
		\13145_b1 , \13145_b0 , \13146_b1 , \13146_b0 , \13147_b1 , \13147_b0 , \13148_b1 , \13148_b0 , \13149_b1 , \13149_b0 , 
		\13150_b1 , \13150_b0 , \13151_b1 , \13151_b0 , \13152_b1 , \13152_b0 , \13153_b1 , \13153_b0 , \13154_b1 , \13154_b0 , 
		\13155_b1 , \13155_b0 , \13156_b1 , \13156_b0 , \13157_b1 , \13157_b0 , \13158_b1 , \13158_b0 , \13159_b1 , \13159_b0 , 
		\13160_b1 , \13160_b0 , \13161_b1 , \13161_b0 , \13162_b1 , \13162_b0 , \13163_b1 , \13163_b0 , \13164_b1 , \13164_b0 , 
		\13165_b1 , \13165_b0 , \13166_b1 , \13166_b0 , \13167_b1 , \13167_b0 , \13168_b1 , \13168_b0 , \13169_b1 , \13169_b0 , 
		\13170_b1 , \13170_b0 , \13171_b1 , \13171_b0 , \13172_b1 , \13172_b0 , \13173_b1 , \13173_b0 , \13174_b1 , \13174_b0 , 
		\13175_b1 , \13175_b0 , \13176_b1 , \13176_b0 , \13177_b1 , \13177_b0 , \13178_b1 , \13178_b0 , \13179_b1 , \13179_b0 , 
		\13180_b1 , \13180_b0 , \13181_b1 , \13181_b0 , \13182_b1 , \13182_b0 , \13183_b1 , \13183_b0 , \13184_b1 , \13184_b0 , 
		\13185_b1 , \13185_b0 , \13186_b1 , \13186_b0 , \13187_b1 , \13187_b0 , \13188_b1 , \13188_b0 , \13189_b1 , \13189_b0 , 
		\13190_b1 , \13190_b0 , \13191_b1 , \13191_b0 , \13192_b1 , \13192_b0 , \13193_b1 , \13193_b0 , \13194_b1 , \13194_b0 , 
		\13195_b1 , \13195_b0 , \13196_b1 , \13196_b0 , \13197_b1 , \13197_b0 , \13198_b1 , \13198_b0 , \13199_b1 , \13199_b0 , 
		\13200_b1 , \13200_b0 , \13201_b1 , \13201_b0 , \13202_b1 , \13202_b0 , \13203_b1 , \13203_b0 , \13204_b1 , \13204_b0 , 
		\13205_b1 , \13205_b0 , \13206_b1 , \13206_b0 , \13207_b1 , \13207_b0 , \13208_b1 , \13208_b0 , \13209_b1 , \13209_b0 , 
		\13210_b1 , \13210_b0 , \13211_b1 , \13211_b0 , \13212_b1 , \13212_b0 , \13213_b1 , \13213_b0 , \13214_b1 , \13214_b0 , 
		\13215_b1 , \13215_b0 , \13216_b1 , \13216_b0 , \13217_b1 , \13217_b0 , \13218_b1 , \13218_b0 , \13219_b1 , \13219_b0 , 
		\13220_b1 , \13220_b0 , \13221_b1 , \13221_b0 , \13222_b1 , \13222_b0 , \13223_b1 , \13223_b0 , \13224_b1 , \13224_b0 , 
		\13225_b1 , \13225_b0 , \13226_b1 , \13226_b0 , \13227_b1 , \13227_b0 , \13228_b1 , \13228_b0 , \13229_b1 , \13229_b0 , 
		\13230_b1 , \13230_b0 , \13231_b1 , \13231_b0 , \13232_b1 , \13232_b0 , \13233_b1 , \13233_b0 , \13234_b1 , \13234_b0 , 
		\13235_b1 , \13235_b0 , \13236_b1 , \13236_b0 , \13237_b1 , \13237_b0 , \13238_b1 , \13238_b0 , \13239_b1 , \13239_b0 , 
		\13240_b1 , \13240_b0 , \13241_b1 , \13241_b0 , \13242_b1 , \13242_b0 , \13243_b1 , \13243_b0 , \13244_b1 , \13244_b0 , 
		\13245_b1 , \13245_b0 , \13246_b1 , \13246_b0 , \13247_b1 , \13247_b0 , \13248_b1 , \13248_b0 , \13249_b1 , \13249_b0 , 
		\13250_b1 , \13250_b0 , \13251_b1 , \13251_b0 , \13252_b1 , \13252_b0 , \13253_b1 , \13253_b0 , \13254_b1 , \13254_b0 , 
		\13255_b1 , \13255_b0 , \13256_b1 , \13256_b0 , \13257_b1 , \13257_b0 , \13258_b1 , \13258_b0 , \13259_b1 , \13259_b0 , 
		\13260_b1 , \13260_b0 , \13261_b1 , \13261_b0 , \13262_b1 , \13262_b0 , \13263_b1 , \13263_b0 , \13264_b1 , \13264_b0 , 
		\13265_b1 , \13265_b0 , \13266_b1 , \13266_b0 , \13267_b1 , \13267_b0 , \13268_b1 , \13268_b0 , \13269_b1 , \13269_b0 , 
		\13270_b1 , \13270_b0 , \13271_b1 , \13271_b0 , \13272_b1 , \13272_b0 , \13273_b1 , \13273_b0 , \13274_b1 , \13274_b0 , 
		\13275_b1 , \13275_b0 , \13276_b1 , \13276_b0 , \13277_b1 , \13277_b0 , \13278_b1 , \13278_b0 , \13279_b1 , \13279_b0 , 
		\13280_b1 , \13280_b0 , \13281_b1 , \13281_b0 , \13282_b1 , \13282_b0 , \13283_b1 , \13283_b0 , \13284_b1 , \13284_b0 , 
		\13285_b1 , \13285_b0 , \13286_b1 , \13286_b0 , \13287_b1 , \13287_b0 , \13288_b1 , \13288_b0 , \13289_b1 , \13289_b0 , 
		\13290_b1 , \13290_b0 , \13291_b1 , \13291_b0 , \13292_b1 , \13292_b0 , \13293_b1 , \13293_b0 , \13294_b1 , \13294_b0 , 
		\13295_b1 , \13295_b0 , \13296_b1 , \13296_b0 , \13297_b1 , \13297_b0 , \13298_b1 , \13298_b0 , \13299_b1 , \13299_b0 , 
		\13300_b1 , \13300_b0 , \13301_b1 , \13301_b0 , \13302_b1 , \13302_b0 , \13303_b1 , \13303_b0 , \13304_b1 , \13304_b0 , 
		\13305_b1 , \13305_b0 , \13306_b1 , \13306_b0 , \13307_b1 , \13307_b0 , \13308_b1 , \13308_b0 , \13309_b1 , \13309_b0 , 
		\13310_b1 , \13310_b0 , \13311_b1 , \13311_b0 , \13312_b1 , \13312_b0 , \13313_b1 , \13313_b0 , \13314_b1 , \13314_b0 , 
		\13315_b1 , \13315_b0 , \13316_b1 , \13316_b0 , \13317_b1 , \13317_b0 , \13318_b1 , \13318_b0 , \13319_b1 , \13319_b0 , 
		\13320_b1 , \13320_b0 , \13321_b1 , \13321_b0 , \13322_b1 , \13322_b0 , \13323_b1 , \13323_b0 , \13324_b1 , \13324_b0 , 
		\13325_b1 , \13325_b0 , \13326_b1 , \13326_b0 , \13327_b1 , \13327_b0 , \13328_b1 , \13328_b0 , \13329_b1 , \13329_b0 , 
		\13330_b1 , \13330_b0 , \13331_b1 , \13331_b0 , \13332_b1 , \13332_b0 , \13333_b1 , \13333_b0 , \13334_b1 , \13334_b0 , 
		\13335_b1 , \13335_b0 , \13336_b1 , \13336_b0 , \13337_b1 , \13337_b0 , \13338_b1 , \13338_b0 , \13339_b1 , \13339_b0 , 
		\13340_b1 , \13340_b0 , \13341_b1 , \13341_b0 , \13342_b1 , \13342_b0 , \13343_b1 , \13343_b0 , \13344_b1 , \13344_b0 , 
		\13345_b1 , \13345_b0 , \13346_b1 , \13346_b0 , \13347_b1 , \13347_b0 , \13348_b1 , \13348_b0 , \13349_b1 , \13349_b0 , 
		\13350_b1 , \13350_b0 , \13351_b1 , \13351_b0 , \13352_b1 , \13352_b0 , \13353_b1 , \13353_b0 , \13354_b1 , \13354_b0 , 
		\13355_b1 , \13355_b0 , \13356_b1 , \13356_b0 , \13357_b1 , \13357_b0 , \13358_b1 , \13358_b0 , \13359_b1 , \13359_b0 , 
		\13360_b1 , \13360_b0 , \13361_b1 , \13361_b0 , \13362_b1 , \13362_b0 , \13363_b1 , \13363_b0 , \13364_b1 , \13364_b0 , 
		\13365_b1 , \13365_b0 , \13366_b1 , \13366_b0 , \13367_b1 , \13367_b0 , \13368_b1 , \13368_b0 , \13369_b1 , \13369_b0 , 
		\13370_b1 , \13370_b0 , \13371_b1 , \13371_b0 , \13372_b1 , \13372_b0 , \13373_b1 , \13373_b0 , \13374_b1 , \13374_b0 , 
		\13375_b1 , \13375_b0 , \13376_b1 , \13376_b0 , \13377_b1 , \13377_b0 , \13378_b1 , \13378_b0 , \13379_b1 , \13379_b0 , 
		\13380_b1 , \13380_b0 , \13381_b1 , \13381_b0 , \13382_b1 , \13382_b0 , \13383_b1 , \13383_b0 , \13384_b1 , \13384_b0 , 
		\13385_b1 , \13385_b0 , \13386_b1 , \13386_b0 , \13387_b1 , \13387_b0 , \13388_b1 , \13388_b0 , \13389_b1 , \13389_b0 , 
		\13390_b1 , \13390_b0 , \13391_b1 , \13391_b0 , \13392_b1 , \13392_b0 , \13393_b1 , \13393_b0 , \13394_b1 , \13394_b0 , 
		\13395_b1 , \13395_b0 , \13396_b1 , \13396_b0 , \13397_b1 , \13397_b0 , \13398_b1 , \13398_b0 , \13399_b1 , \13399_b0 , 
		\13400_b1 , \13400_b0 , \13401_b1 , \13401_b0 , \13402_b1 , \13402_b0 , \13403_b1 , \13403_b0 , \13404_b1 , \13404_b0 , 
		\13405_b1 , \13405_b0 , \13406_b1 , \13406_b0 , \13407_b1 , \13407_b0 , \13408_b1 , \13408_b0 , \13409_b1 , \13409_b0 , 
		\13410_b1 , \13410_b0 , \13411_b1 , \13411_b0 , \13412_b1 , \13412_b0 , \13413_b1 , \13413_b0 , \13414_b1 , \13414_b0 , 
		\13415_b1 , \13415_b0 , \13416_b1 , \13416_b0 , \13417_b1 , \13417_b0 , \13418_b1 , \13418_b0 , \13419_b1 , \13419_b0 , 
		\13420_b1 , \13420_b0 , \13421_b1 , \13421_b0 , \13422_b1 , \13422_b0 , \13423_b1 , \13423_b0 , \13424_b1 , \13424_b0 , 
		\13425_b1 , \13425_b0 , \13426_b1 , \13426_b0 , \13427_b1 , \13427_b0 , \13428_b1 , \13428_b0 , \13429_b1 , \13429_b0 , 
		\13430_b1 , \13430_b0 , \13431_b1 , \13431_b0 , \13432_b1 , \13432_b0 , \13433_b1 , \13433_b0 , \13434_b1 , \13434_b0 , 
		\13435_b1 , \13435_b0 , \13436_b1 , \13436_b0 , \13437_b1 , \13437_b0 , \13438_b1 , \13438_b0 , \13439_b1 , \13439_b0 , 
		\13440_b1 , \13440_b0 , \13441_b1 , \13441_b0 , \13442_b1 , \13442_b0 , \13443_b1 , \13443_b0 , \13444_b1 , \13444_b0 , 
		\13445_b1 , \13445_b0 , \13446_b1 , \13446_b0 , \13447_b1 , \13447_b0 , \13448_b1 , \13448_b0 , \13449_b1 , \13449_b0 , 
		\13450_b1 , \13450_b0 , \13451_b1 , \13451_b0 , \13452_b1 , \13452_b0 , \13453_b1 , \13453_b0 , \13454_b1 , \13454_b0 , 
		\13455_b1 , \13455_b0 , \13456_b1 , \13456_b0 , \13457_b1 , \13457_b0 , \13458_b1 , \13458_b0 , \13459_b1 , \13459_b0 , 
		\13460_b1 , \13460_b0 , \13461_b1 , \13461_b0 , \13462_b1 , \13462_b0 , \13463_b1 , \13463_b0 , \13464_b1 , \13464_b0 , 
		\13465_b1 , \13465_b0 , \13466_b1 , \13466_b0 , \13467_b1 , \13467_b0 , \13468_b1 , \13468_b0 , \13469_b1 , \13469_b0 , 
		\13470_b1 , \13470_b0 , \13471_b1 , \13471_b0 , \13472_b1 , \13472_b0 , \13473_b1 , \13473_b0 , \13474_b1 , \13474_b0 , 
		\13475_b1 , \13475_b0 , \13476_b1 , \13476_b0 , \13477_b1 , \13477_b0 , \13478_b1 , \13478_b0 , \13479_b1 , \13479_b0 , 
		\13480_b1 , \13480_b0 , \13481_b1 , \13481_b0 , \13482_b1 , \13482_b0 , \13483_b1 , \13483_b0 , \13484_b1 , \13484_b0 , 
		\13485_b1 , \13485_b0 , \13486_b1 , \13486_b0 , \13487_b1 , \13487_b0 , \13488_b1 , \13488_b0 , \13489_b1 , \13489_b0 , 
		\13490_b1 , \13490_b0 , \13491_b1 , \13491_b0 , \13492_b1 , \13492_b0 , \13493_b1 , \13493_b0 , \13494_b1 , \13494_b0 , 
		\13495_b1 , \13495_b0 , \13496_b1 , \13496_b0 , \13497_b1 , \13497_b0 , \13498_b1 , \13498_b0 , \13499_b1 , \13499_b0 , 
		\13500_b1 , \13500_b0 , \13501_b1 , \13501_b0 , \13502_b1 , \13502_b0 , \13503_b1 , \13503_b0 , \13504_b1 , \13504_b0 , 
		\13505_b1 , \13505_b0 , \13506_b1 , \13506_b0 , \13507_b1 , \13507_b0 , \13508_b1 , \13508_b0 , \13509_b1 , \13509_b0 , 
		\13510_b1 , \13510_b0 , \13511_b1 , \13511_b0 , \13512_b1 , \13512_b0 , \13513_b1 , \13513_b0 , \13514_b1 , \13514_b0 , 
		\13515_b1 , \13515_b0 , \13516_b1 , \13516_b0 , \13517_b1 , \13517_b0 , \13518_b1 , \13518_b0 , \13519_b1 , \13519_b0 , 
		\13520_b1 , \13520_b0 , \13521_b1 , \13521_b0 , \13522_b1 , \13522_b0 , \13523_b1 , \13523_b0 , \13524_b1 , \13524_b0 , 
		\13525_b1 , \13525_b0 , \13526_b1 , \13526_b0 , \13527_b1 , \13527_b0 , \13528_b1 , \13528_b0 , \13529_b1 , \13529_b0 , 
		\13530_b1 , \13530_b0 , \13531_b1 , \13531_b0 , \13532_b1 , \13532_b0 , \13533_b1 , \13533_b0 , \13534_b1 , \13534_b0 , 
		\13535_b1 , \13535_b0 , \13536_b1 , \13536_b0 , \13537_b1 , \13537_b0 , \13538_b1 , \13538_b0 , \13539_b1 , \13539_b0 , 
		\13540_b1 , \13540_b0 , \13541_b1 , \13541_b0 , \13542_b1 , \13542_b0 , \13543_b1 , \13543_b0 , \13544_b1 , \13544_b0 , 
		\13545_b1 , \13545_b0 , \13546_b1 , \13546_b0 , \13547_b1 , \13547_b0 , \13548_b1 , \13548_b0 , \13549_b1 , \13549_b0 , 
		\13550_b1 , \13550_b0 , \13551_b1 , \13551_b0 , \13552_b1 , \13552_b0 , \13553_b1 , \13553_b0 , \13554_b1 , \13554_b0 , 
		\13555_b1 , \13555_b0 , \13556_b1 , \13556_b0 , \13557_b1 , \13557_b0 , \13558_b1 , \13558_b0 , \13559_b1 , \13559_b0 , 
		\13560_b1 , \13560_b0 , \13561_b1 , \13561_b0 , \13562_b1 , \13562_b0 , \13563_b1 , \13563_b0 , \13564_b1 , \13564_b0 , 
		\13565_b1 , \13565_b0 , \13566_b1 , \13566_b0 , \13567_b1 , \13567_b0 , \13568_b1 , \13568_b0 , \13569_b1 , \13569_b0 , 
		\13570_b1 , \13570_b0 , \13571_b1 , \13571_b0 , \13572_b1 , \13572_b0 , \13573_b1 , \13573_b0 , \13574_b1 , \13574_b0 , 
		\13575_b1 , \13575_b0 , \13576_b1 , \13576_b0 , \13577_b1 , \13577_b0 , \13578_b1 , \13578_b0 , \13579_b1 , \13579_b0 , 
		\13580_b1 , \13580_b0 , \13581_b1 , \13581_b0 , \13582_b1 , \13582_b0 , \13583_b1 , \13583_b0 , \13584_b1 , \13584_b0 , 
		\13585_b1 , \13585_b0 , \13586_b1 , \13586_b0 , \13587_b1 , \13587_b0 , \13588_b1 , \13588_b0 , \13589_b1 , \13589_b0 , 
		\13590_b1 , \13590_b0 , \13591_b1 , \13591_b0 , \13592_b1 , \13592_b0 , \13593_b1 , \13593_b0 , \13594_b1 , \13594_b0 , 
		\13595_b1 , \13595_b0 , \13596_b1 , \13596_b0 , \13597_b1 , \13597_b0 , \13598_b1 , \13598_b0 , \13599_b1 , \13599_b0 , 
		\13600_b1 , \13600_b0 , \13601_b1 , \13601_b0 , \13602_b1 , \13602_b0 , \13603_b1 , \13603_b0 , \13604_b1 , \13604_b0 , 
		\13605_b1 , \13605_b0 , \13606_b1 , \13606_b0 , \13607_b1 , \13607_b0 , \13608_b1 , \13608_b0 , \13609_b1 , \13609_b0 , 
		\13610_b1 , \13610_b0 , \13611_b1 , \13611_b0 , \13612_b1 , \13612_b0 , \13613_b1 , \13613_b0 , \13614_b1 , \13614_b0 , 
		\13615_b1 , \13615_b0 , \13616_b1 , \13616_b0 , \13617_b1 , \13617_b0 , \13618_b1 , \13618_b0 , \13619_b1 , \13619_b0 , 
		\13620_b1 , \13620_b0 , \13621_b1 , \13621_b0 , \13622_b1 , \13622_b0 , \13623_b1 , \13623_b0 , \13624_b1 , \13624_b0 , 
		\13625_b1 , \13625_b0 , \13626_b1 , \13626_b0 , \13627_b1 , \13627_b0 , \13628_b1 , \13628_b0 , \13629_b1 , \13629_b0 , 
		\13630_b1 , \13630_b0 , \13631_b1 , \13631_b0 , \13632_b1 , \13632_b0 , \13633_b1 , \13633_b0 , \13634_b1 , \13634_b0 , 
		\13635_b1 , \13635_b0 , \13636_b1 , \13636_b0 , \13637_b1 , \13637_b0 , \13638_b1 , \13638_b0 , \13639_b1 , \13639_b0 , 
		\13640_b1 , \13640_b0 , \13641_b1 , \13641_b0 , \13642_b1 , \13642_b0 , \13643_b1 , \13643_b0 , \13644_b1 , \13644_b0 , 
		\13645_b1 , \13645_b0 , \13646_b1 , \13646_b0 , \13647_b1 , \13647_b0 , \13648_b1 , \13648_b0 , \13649_b1 , \13649_b0 , 
		\13650_b1 , \13650_b0 , \13651_b1 , \13651_b0 , \13652_b1 , \13652_b0 , \13653_b1 , \13653_b0 , \13654_b1 , \13654_b0 , 
		\13655_b1 , \13655_b0 , \13656_b1 , \13656_b0 , \13657_b1 , \13657_b0 , \13658_b1 , \13658_b0 , \13659_b1 , \13659_b0 , 
		\13660_b1 , \13660_b0 , \13661_b1 , \13661_b0 , \13662_b1 , \13662_b0 , \13663_b1 , \13663_b0 , \13664_b1 , \13664_b0 , 
		\13665_b1 , \13665_b0 , \13666_b1 , \13666_b0 , \13667_b1 , \13667_b0 , \13668_b1 , \13668_b0 , \13669_b1 , \13669_b0 , 
		\13670_b1 , \13670_b0 , \13671_b1 , \13671_b0 , \13672_b1 , \13672_b0 , \13673_b1 , \13673_b0 , \13674_b1 , \13674_b0 , 
		\13675_b1 , \13675_b0 , \13676_b1 , \13676_b0 , \13677_b1 , \13677_b0 , \13678_b1 , \13678_b0 , \13679_b1 , \13679_b0 , 
		\13680_b1 , \13680_b0 , \13681_b1 , \13681_b0 , \13682_b1 , \13682_b0 , \13683_b1 , \13683_b0 , \13684_b1 , \13684_b0 , 
		\13685_b1 , \13685_b0 , \13686_b1 , \13686_b0 , \13687_b1 , \13687_b0 , \13688_b1 , \13688_b0 , \13689_b1 , \13689_b0 , 
		\13690_b1 , \13690_b0 , \13691_b1 , \13691_b0 , \13692_b1 , \13692_b0 , \13693_b1 , \13693_b0 , \13694_b1 , \13694_b0 , 
		\13695_b1 , \13695_b0 , \13696_b1 , \13696_b0 , \13697_b1 , \13697_b0 , \13698_b1 , \13698_b0 , \13699_b1 , \13699_b0 , 
		\13700_b1 , \13700_b0 , \13701_b1 , \13701_b0 , \13702_b1 , \13702_b0 , \13703_b1 , \13703_b0 , \13704_b1 , \13704_b0 , 
		\13705_b1 , \13705_b0 , \13706_b1 , \13706_b0 , \13707_b1 , \13707_b0 , \13708_b1 , \13708_b0 , \13709_b1 , \13709_b0 , 
		\13710_b1 , \13710_b0 , \13711_b1 , \13711_b0 , \13712_b1 , \13712_b0 , \13713_b1 , \13713_b0 , \13714_b1 , \13714_b0 , 
		\13715_b1 , \13715_b0 , \13716_b1 , \13716_b0 , \13717_b1 , \13717_b0 , \13718_b1 , \13718_b0 , \13719_b1 , \13719_b0 , 
		\13720_b1 , \13720_b0 , \13721_b1 , \13721_b0 , \13722_b1 , \13722_b0 , \13723_b1 , \13723_b0 , \13724_b1 , \13724_b0 , 
		\13725_b1 , \13725_b0 , \13726_b1 , \13726_b0 , \13727_b1 , \13727_b0 , \13728_b1 , \13728_b0 , \13729_b1 , \13729_b0 , 
		\13730_b1 , \13730_b0 , \13731_b1 , \13731_b0 , \13732_b1 , \13732_b0 , \13733_b1 , \13733_b0 , \13734_b1 , \13734_b0 , 
		\13735_b1 , \13735_b0 , \13736_b1 , \13736_b0 , \13737_b1 , \13737_b0 , \13738_b1 , \13738_b0 , \13739_b1 , \13739_b0 , 
		\13740_b1 , \13740_b0 , \13741_b1 , \13741_b0 , \13742_b1 , \13742_b0 , \13743_b1 , \13743_b0 , \13744_b1 , \13744_b0 , 
		\13745_b1 , \13745_b0 , \13746_b1 , \13746_b0 , \13747_b1 , \13747_b0 , \13748_b1 , \13748_b0 , \13749_b1 , \13749_b0 , 
		\13750_b1 , \13750_b0 , \13751_b1 , \13751_b0 , \13752_b1 , \13752_b0 , \13753_b1 , \13753_b0 , \13754_b1 , \13754_b0 , 
		\13755_b1 , \13755_b0 , \13756_b1 , \13756_b0 , \13757_b1 , \13757_b0 , \13758_b1 , \13758_b0 , \13759_b1 , \13759_b0 , 
		\13760_b1 , \13760_b0 , \13761_b1 , \13761_b0 , \13762_b1 , \13762_b0 , \13763_b1 , \13763_b0 , \13764_b1 , \13764_b0 , 
		\13765_b1 , \13765_b0 , \13766_b1 , \13766_b0 , \13767_b1 , \13767_b0 , \13768_b1 , \13768_b0 , \13769_b1 , \13769_b0 , 
		\13770_b1 , \13770_b0 , \13771_b1 , \13771_b0 , \13772_b1 , \13772_b0 , \13773_b1 , \13773_b0 , \13774_b1 , \13774_b0 , 
		\13775_b1 , \13775_b0 , \13776_b1 , \13776_b0 , \13777_b1 , \13777_b0 , \13778_b1 , \13778_b0 , \13779_b1 , \13779_b0 , 
		\13780_b1 , \13780_b0 , \13781_b1 , \13781_b0 , \13782_b1 , \13782_b0 , \13783_b1 , \13783_b0 , \13784_b1 , \13784_b0 , 
		\13785_b1 , \13785_b0 , \13786_b1 , \13786_b0 , \13787_b1 , \13787_b0 , \13788_b1 , \13788_b0 , \13789_b1 , \13789_b0 , 
		\13790_b1 , \13790_b0 , \13791_b1 , \13791_b0 , \13792_b1 , \13792_b0 , \13793_b1 , \13793_b0 , \13794_b1 , \13794_b0 , 
		\13795_b1 , \13795_b0 , \13796_b1 , \13796_b0 , \13797_b1 , \13797_b0 , \13798_b1 , \13798_b0 , \13799_b1 , \13799_b0 , 
		\13800_b1 , \13800_b0 , \13801_b1 , \13801_b0 , \13802_b1 , \13802_b0 , \13803_b1 , \13803_b0 , \13804_b1 , \13804_b0 , 
		\13805_b1 , \13805_b0 , \13806_b1 , \13806_b0 , \13807_b1 , \13807_b0 , \13808_b1 , \13808_b0 , \13809_b1 , \13809_b0 , 
		\13810_b1 , \13810_b0 , \13811_b1 , \13811_b0 , \13812_b1 , \13812_b0 , \13813_b1 , \13813_b0 , \13814_b1 , \13814_b0 , 
		\13815_b1 , \13815_b0 , \13816_b1 , \13816_b0 , \13817_b1 , \13817_b0 , \13818_b1 , \13818_b0 , \13819_b1 , \13819_b0 , 
		\13820_b1 , \13820_b0 , \13821_b1 , \13821_b0 , \13822_b1 , \13822_b0 , \13823_b1 , \13823_b0 , \13824_b1 , \13824_b0 , 
		\13825_b1 , \13825_b0 , \13826_b1 , \13826_b0 , \13827_b1 , \13827_b0 , \13828_b1 , \13828_b0 , \13829_b1 , \13829_b0 , 
		\13830_b1 , \13830_b0 , \13831_b1 , \13831_b0 , \13832_b1 , \13832_b0 , \13833_b1 , \13833_b0 , \13834_b1 , \13834_b0 , 
		\13835_b1 , \13835_b0 , \13836_b1 , \13836_b0 , \13837_b1 , \13837_b0 , \13838_b1 , \13838_b0 , \13839_b1 , \13839_b0 , 
		\13840_b1 , \13840_b0 , \13841_b1 , \13841_b0 , \13842_b1 , \13842_b0 , \13843_b1 , \13843_b0 , \13844_b1 , \13844_b0 , 
		\13845_b1 , \13845_b0 , \13846_b1 , \13846_b0 , \13847_b1 , \13847_b0 , \13848_b1 , \13848_b0 , \13849_b1 , \13849_b0 , 
		\13850_b1 , \13850_b0 , \13851_b1 , \13851_b0 , \13852_b1 , \13852_b0 , \13853_b1 , \13853_b0 , \13854_b1 , \13854_b0 , 
		\13855_b1 , \13855_b0 , \13856_b1 , \13856_b0 , \13857_b1 , \13857_b0 , \13858_b1 , \13858_b0 , \13859_b1 , \13859_b0 , 
		\13860_b1 , \13860_b0 , \13861_b1 , \13861_b0 , \13862_b1 , \13862_b0 , \13863_b1 , \13863_b0 , \13864_b1 , \13864_b0 , 
		\13865_b1 , \13865_b0 , \13866_b1 , \13866_b0 , \13867_b1 , \13867_b0 , \13868_b1 , \13868_b0 , \13869_b1 , \13869_b0 , 
		\13870_b1 , \13870_b0 , \13871_b1 , \13871_b0 , \13872_b1 , \13872_b0 , \13873_b1 , \13873_b0 , \13874_b1 , \13874_b0 , 
		\13875_b1 , \13875_b0 , \13876_b1 , \13876_b0 , \13877_b1 , \13877_b0 , \13878_b1 , \13878_b0 , \13879_b1 , \13879_b0 , 
		\13880_b1 , \13880_b0 , \13881_b1 , \13881_b0 , \13882_b1 , \13882_b0 , \13883_b1 , \13883_b0 , \13884_b1 , \13884_b0 , 
		\13885_b1 , \13885_b0 , \13886_b1 , \13886_b0 , \13887_b1 , \13887_b0 , \13888_b1 , \13888_b0 , \13889_b1 , \13889_b0 , 
		\13890_b1 , \13890_b0 , \13891_b1 , \13891_b0 , \13892_b1 , \13892_b0 , \13893_b1 , \13893_b0 , \13894_b1 , \13894_b0 , 
		\13895_b1 , \13895_b0 , \13896_b1 , \13896_b0 , \13897_b1 , \13897_b0 , \13898_b1 , \13898_b0 , \13899_b1 , \13899_b0 , 
		\13900_b1 , \13900_b0 , \13901_b1 , \13901_b0 , \13902_b1 , \13902_b0 , \13903_b1 , \13903_b0 , \13904_b1 , \13904_b0 , 
		\13905_b1 , \13905_b0 , \13906_b1 , \13906_b0 , \13907_b1 , \13907_b0 , \13908_b1 , \13908_b0 , \13909_b1 , \13909_b0 , 
		\13910_b1 , \13910_b0 , \13911_b1 , \13911_b0 , \13912_b1 , \13912_b0 , \13913_b1 , \13913_b0 , \13914_b1 , \13914_b0 , 
		\13915_b1 , \13915_b0 , \13916_b1 , \13916_b0 , \13917_b1 , \13917_b0 , \13918_b1 , \13918_b0 , \13919_b1 , \13919_b0 , 
		\13920_b1 , \13920_b0 , \13921_b1 , \13921_b0 , \13922_b1 , \13922_b0 , \13923_b1 , \13923_b0 , \13924_b1 , \13924_b0 , 
		\13925_b1 , \13925_b0 , \13926_b1 , \13926_b0 , \13927_b1 , \13927_b0 , \13928_b1 , \13928_b0 , \13929_b1 , \13929_b0 , 
		\13930_b1 , \13930_b0 , \13931_b1 , \13931_b0 , \13932_b1 , \13932_b0 , \13933_b1 , \13933_b0 , \13934_b1 , \13934_b0 , 
		\13935_b1 , \13935_b0 , \13936_b1 , \13936_b0 , \13937_b1 , \13937_b0 , \13938_b1 , \13938_b0 , \13939_b1 , \13939_b0 , 
		\13940_b1 , \13940_b0 , \13941_b1 , \13941_b0 , \13942_b1 , \13942_b0 , \13943_b1 , \13943_b0 , \13944_b1 , \13944_b0 , 
		\13945_b1 , \13945_b0 , \13946_b1 , \13946_b0 , \13947_b1 , \13947_b0 , \13948_b1 , \13948_b0 , \13949_b1 , \13949_b0 , 
		\13950_b1 , \13950_b0 , \13951_b1 , \13951_b0 , \13952_b1 , \13952_b0 , \13953_b1 , \13953_b0 , \13954_b1 , \13954_b0 , 
		\13955_b1 , \13955_b0 , \13956_b1 , \13956_b0 , \13957_b1 , \13957_b0 , \13958_b1 , \13958_b0 , \13959_b1 , \13959_b0 , 
		\13960_b1 , \13960_b0 , \13961_b1 , \13961_b0 , \13962_b1 , \13962_b0 , \13963_b1 , \13963_b0 , \13964_b1 , \13964_b0 , 
		\13965_b1 , \13965_b0 , \13966_b1 , \13966_b0 , \13967_b1 , \13967_b0 , \13968_b1 , \13968_b0 , \13969_b1 , \13969_b0 , 
		\13970_b1 , \13970_b0 , \13971_b1 , \13971_b0 , \13972_b1 , \13972_b0 , \13973_b1 , \13973_b0 , \13974_b1 , \13974_b0 , 
		\13975_b1 , \13975_b0 , \13976_b1 , \13976_b0 , \13977_b1 , \13977_b0 , \13978_b1 , \13978_b0 , \13979_b1 , \13979_b0 , 
		\13980_b1 , \13980_b0 , \13981_b1 , \13981_b0 , \13982_b1 , \13982_b0 , \13983_b1 , \13983_b0 , \13984_b1 , \13984_b0 , 
		\13985_b1 , \13985_b0 , \13986_b1 , \13986_b0 , \13987_b1 , \13987_b0 , \13988_b1 , \13988_b0 , \13989_b1 , \13989_b0 , 
		\13990_b1 , \13990_b0 , \13991_b1 , \13991_b0 , \13992_b1 , \13992_b0 , \13993_b1 , \13993_b0 , \13994_b1 , \13994_b0 , 
		\13995_b1 , \13995_b0 , \13996_b1 , \13996_b0 , \13997_b1 , \13997_b0 , \13998_b1 , \13998_b0 , \13999_b1 , \13999_b0 , 
		\14000_b1 , \14000_b0 , \14001_b1 , \14001_b0 , \14002_b1 , \14002_b0 , \14003_b1 , \14003_b0 , \14004_b1 , \14004_b0 , 
		\14005_b1 , \14005_b0 , \14006_b1 , \14006_b0 , \14007_b1 , \14007_b0 , \14008_b1 , \14008_b0 , \14009_b1 , \14009_b0 , 
		\14010_b1 , \14010_b0 , \14011_b1 , \14011_b0 , \14012_b1 , \14012_b0 , \14013_b1 , \14013_b0 , \14014_b1 , \14014_b0 , 
		\14015_b1 , \14015_b0 , \14016_b1 , \14016_b0 , \14017_b1 , \14017_b0 , \14018_b1 , \14018_b0 , \14019_b1 , \14019_b0 , 
		\14020_b1 , \14020_b0 , \14021_b1 , \14021_b0 , \14022_b1 , \14022_b0 , \14023_b1 , \14023_b0 , \14024_b1 , \14024_b0 , 
		\14025_b1 , \14025_b0 , \14026_b1 , \14026_b0 , \14027_b1 , \14027_b0 , \14028_b1 , \14028_b0 , \14029_b1 , \14029_b0 , 
		\14030_b1 , \14030_b0 , \14031_b1 , \14031_b0 , \14032_b1 , \14032_b0 , \14033_b1 , \14033_b0 , \14034_b1 , \14034_b0 , 
		\14035_b1 , \14035_b0 , \14036_b1 , \14036_b0 , \14037_b1 , \14037_b0 , \14038_b1 , \14038_b0 , \14039_b1 , \14039_b0 , 
		\14040_b1 , \14040_b0 , \14041_b1 , \14041_b0 , \14042_b1 , \14042_b0 , \14043_b1 , \14043_b0 , \14044_b1 , \14044_b0 , 
		\14045_b1 , \14045_b0 , \14046_b1 , \14046_b0 , \14047_b1 , \14047_b0 , \14048_b1 , \14048_b0 , \14049_b1 , \14049_b0 , 
		\14050_b1 , \14050_b0 , \14051_b1 , \14051_b0 , \14052_b1 , \14052_b0 , \14053_b1 , \14053_b0 , \14054_b1 , \14054_b0 , 
		\14055_b1 , \14055_b0 , \14056_b1 , \14056_b0 , \14057_b1 , \14057_b0 , \14058_b1 , \14058_b0 , \14059_b1 , \14059_b0 , 
		\14060_b1 , \14060_b0 , \14061_b1 , \14061_b0 , \14062_b1 , \14062_b0 , \14063_b1 , \14063_b0 , \14064_b1 , \14064_b0 , 
		\14065_b1 , \14065_b0 , \14066_b1 , \14066_b0 , \14067_b1 , \14067_b0 , \14068_b1 , \14068_b0 , \14069_b1 , \14069_b0 , 
		\14070_b1 , \14070_b0 , \14071_b1 , \14071_b0 , \14072_b1 , \14072_b0 , \14073_b1 , \14073_b0 , \14074_b1 , \14074_b0 , 
		\14075_b1 , \14075_b0 , \14076_b1 , \14076_b0 , \14077_b1 , \14077_b0 , \14078_b1 , \14078_b0 , \14079_b1 , \14079_b0 , 
		\14080_b1 , \14080_b0 , \14081_b1 , \14081_b0 , \14082_b1 , \14082_b0 , \14083_b1 , \14083_b0 , \14084_b1 , \14084_b0 , 
		\14085_b1 , \14085_b0 , \14086_b1 , \14086_b0 , \14087_b1 , \14087_b0 , \14088_b1 , \14088_b0 , \14089_b1 , \14089_b0 , 
		\14090_b1 , \14090_b0 , \14091_b1 , \14091_b0 , \14092_b1 , \14092_b0 , \14093_b1 , \14093_b0 , \14094_b1 , \14094_b0 , 
		\14095_b1 , \14095_b0 , \14096_b1 , \14096_b0 , \14097_b1 , \14097_b0 , \14098_b1 , \14098_b0 , \14099_b1 , \14099_b0 , 
		\14100_b1 , \14100_b0 , \14101_b1 , \14101_b0 , \14102_b1 , \14102_b0 , \14103_b1 , \14103_b0 , \14104_b1 , \14104_b0 , 
		\14105_b1 , \14105_b0 , \14106_b1 , \14106_b0 , \14107_b1 , \14107_b0 , \14108_b1 , \14108_b0 , \14109_b1 , \14109_b0 , 
		\14110_b1 , \14110_b0 , \14111_b1 , \14111_b0 , \14112_b1 , \14112_b0 , \14113_b1 , \14113_b0 , \14114_b1 , \14114_b0 , 
		\14115_b1 , \14115_b0 , \14116_b1 , \14116_b0 , \14117_b1 , \14117_b0 , \14118_b1 , \14118_b0 , \14119_b1 , \14119_b0 , 
		\14120_b1 , \14120_b0 , \14121_b1 , \14121_b0 , \14122_b1 , \14122_b0 , \14123_b1 , \14123_b0 , \14124_b1 , \14124_b0 , 
		\14125_b1 , \14125_b0 , \14126_b1 , \14126_b0 , \14127_b1 , \14127_b0 , \14128_b1 , \14128_b0 , \14129_b1 , \14129_b0 , 
		\14130_b1 , \14130_b0 , \14131_b1 , \14131_b0 , \14132_b1 , \14132_b0 , \14133_b1 , \14133_b0 , \14134_b1 , \14134_b0 , 
		\14135_b1 , \14135_b0 , \14136_b1 , \14136_b0 , \14137_b1 , \14137_b0 , \14138_b1 , \14138_b0 , \14139_b1 , \14139_b0 , 
		\14140_b1 , \14140_b0 , \14141_b1 , \14141_b0 , \14142_b1 , \14142_b0 , \14143_b1 , \14143_b0 , \14144_b1 , \14144_b0 , 
		\14145_b1 , \14145_b0 , \14146_b1 , \14146_b0 , \14147_b1 , \14147_b0 , \14148_b1 , \14148_b0 , \14149_b1 , \14149_b0 , 
		\14150_b1 , \14150_b0 , \14151_b1 , \14151_b0 , \14152_b1 , \14152_b0 , \14153_b1 , \14153_b0 , \14154_b1 , \14154_b0 , 
		\14155_b1 , \14155_b0 , \14156_b1 , \14156_b0 , \14157_b1 , \14157_b0 , \14158_b1 , \14158_b0 , \14159_b1 , \14159_b0 , 
		\14160_b1 , \14160_b0 , \14161_b1 , \14161_b0 , \14162_b1 , \14162_b0 , \14163_b1 , \14163_b0 , \14164_b1 , \14164_b0 , 
		\14165_b1 , \14165_b0 , \14166_b1 , \14166_b0 , \14167_b1 , \14167_b0 , \14168_b1 , \14168_b0 , \14169_b1 , \14169_b0 , 
		\14170_b1 , \14170_b0 , \14171_b1 , \14171_b0 , \14172_b1 , \14172_b0 , \14173_b1 , \14173_b0 , \14174_b1 , \14174_b0 , 
		\14175_b1 , \14175_b0 , \14176_b1 , \14176_b0 , \14177_b1 , \14177_b0 , \14178_b1 , \14178_b0 , \14179_b1 , \14179_b0 , 
		\14180_b1 , \14180_b0 , \14181_b1 , \14181_b0 , \14182_b1 , \14182_b0 , \14183_b1 , \14183_b0 , \14184_b1 , \14184_b0 , 
		\14185_b1 , \14185_b0 , \14186_b1 , \14186_b0 , \14187_b1 , \14187_b0 , \14188_b1 , \14188_b0 , \14189_b1 , \14189_b0 , 
		\14190_b1 , \14190_b0 , \14191_b1 , \14191_b0 , \14192_b1 , \14192_b0 , \14193_b1 , \14193_b0 , \14194_b1 , \14194_b0 , 
		\14195_b1 , \14195_b0 , \14196_b1 , \14196_b0 , \14197_b1 , \14197_b0 , \14198_b1 , \14198_b0 , \14199_b1 , \14199_b0 , 
		\14200_b1 , \14200_b0 , \14201_b1 , \14201_b0 , \14202_b1 , \14202_b0 , \14203_b1 , \14203_b0 , \14204_b1 , \14204_b0 , 
		\14205_b1 , \14205_b0 , \14206_b1 , \14206_b0 , \14207_b1 , \14207_b0 , \14208_b1 , \14208_b0 , \14209_b1 , \14209_b0 , 
		\14210_b1 , \14210_b0 , \14211_b1 , \14211_b0 , \14212_b1 , \14212_b0 , \14213_b1 , \14213_b0 , \14214_b1 , \14214_b0 , 
		\14215_b1 , \14215_b0 , \14216_b1 , \14216_b0 , \14217_b1 , \14217_b0 , \14218_b1 , \14218_b0 , \14219_b1 , \14219_b0 , 
		\14220_b1 , \14220_b0 , \14221_b1 , \14221_b0 , \14222_b1 , \14222_b0 , \14223_b1 , \14223_b0 , \14224_b1 , \14224_b0 , 
		\14225_b1 , \14225_b0 , \14226_b1 , \14226_b0 , \14227_b1 , \14227_b0 , \14228_b1 , \14228_b0 , \14229_b1 , \14229_b0 , 
		\14230_b1 , \14230_b0 , \14231_b1 , \14231_b0 , \14232_b1 , \14232_b0 , \14233_b1 , \14233_b0 , \14234_b1 , \14234_b0 , 
		\14235_b1 , \14235_b0 , \14236_b1 , \14236_b0 , \14237_b1 , \14237_b0 , \14238_b1 , \14238_b0 , \14239_b1 , \14239_b0 , 
		\14240_b1 , \14240_b0 , \14241_b1 , \14241_b0 , \14242_b1 , \14242_b0 , \14243_b1 , \14243_b0 , \14244_b1 , \14244_b0 , 
		\14245_b1 , \14245_b0 , \14246_b1 , \14246_b0 , \14247_b1 , \14247_b0 , \14248_b1 , \14248_b0 , \14249_b1 , \14249_b0 , 
		\14250_b1 , \14250_b0 , \14251_b1 , \14251_b0 , \14252_b1 , \14252_b0 , \14253_b1 , \14253_b0 , \14254_b1 , \14254_b0 , 
		\14255_b1 , \14255_b0 , \14256_b1 , \14256_b0 , \14257_b1 , \14257_b0 , \14258_b1 , \14258_b0 , \14259_b1 , \14259_b0 , 
		\14260_b1 , \14260_b0 , \14261_b1 , \14261_b0 , \14262_b1 , \14262_b0 , \14263_b1 , \14263_b0 , \14264_b1 , \14264_b0 , 
		\14265_b1 , \14265_b0 , \14266_b1 , \14266_b0 , \14267_b1 , \14267_b0 , \14268_b1 , \14268_b0 , \14269_b1 , \14269_b0 , 
		\14270_b1 , \14270_b0 , \14271_b1 , \14271_b0 , \14272_b1 , \14272_b0 , \14273_b1 , \14273_b0 , \14274_b1 , \14274_b0 , 
		\14275_b1 , \14275_b0 , \14276_b1 , \14276_b0 , \14277_b1 , \14277_b0 , \14278_b1 , \14278_b0 , \14279_b1 , \14279_b0 , 
		\14280_b1 , \14280_b0 , \14281_b1 , \14281_b0 , \14282_b1 , \14282_b0 , \14283_b1 , \14283_b0 , \14284_b1 , \14284_b0 , 
		\14285_b1 , \14285_b0 , \14286_b1 , \14286_b0 , \14287_b1 , \14287_b0 , \14288_b1 , \14288_b0 , \14289_b1 , \14289_b0 , 
		\14290_b1 , \14290_b0 , \14291_b1 , \14291_b0 , \14292_b1 , \14292_b0 , \14293_b1 , \14293_b0 , \14294_b1 , \14294_b0 , 
		\14295_b1 , \14295_b0 , \14296_b1 , \14296_b0 , \14297_b1 , \14297_b0 , \14298_b1 , \14298_b0 , \14299_b1 , \14299_b0 , 
		\14300_b1 , \14300_b0 , \14301_b1 , \14301_b0 , \14302_b1 , \14302_b0 , \14303_b1 , \14303_b0 , \14304_b1 , \14304_b0 , 
		\14305_b1 , \14305_b0 , \14306_b1 , \14306_b0 , \14307_b1 , \14307_b0 , \14308_b1 , \14308_b0 , \14309_b1 , \14309_b0 , 
		\14310_b1 , \14310_b0 , \14311_b1 , \14311_b0 , \14312_b1 , \14312_b0 , \14313_b1 , \14313_b0 , \14314_b1 , \14314_b0 , 
		\14315_b1 , \14315_b0 , \14316_b1 , \14316_b0 , \14317_b1 , \14317_b0 , \14318_b1 , \14318_b0 , \14319_b1 , \14319_b0 , 
		\14320_b1 , \14320_b0 , \14321_b1 , \14321_b0 , \14322_b1 , \14322_b0 , \14323_b1 , \14323_b0 , \14324_b1 , \14324_b0 , 
		\14325_b1 , \14325_b0 , \14326_b1 , \14326_b0 , \14327_b1 , \14327_b0 , \14328_b1 , \14328_b0 , \14329_b1 , \14329_b0 , 
		\14330_b1 , \14330_b0 , \14331_b1 , \14331_b0 , \14332_b1 , \14332_b0 , \14333_b1 , \14333_b0 , \14334_b1 , \14334_b0 , 
		\14335_b1 , \14335_b0 , \14336_b1 , \14336_b0 , \14337_b1 , \14337_b0 , \14338_b1 , \14338_b0 , \14339_b1 , \14339_b0 , 
		\14340_b1 , \14340_b0 , \14341_b1 , \14341_b0 , \14342_b1 , \14342_b0 , \14343_b1 , \14343_b0 , \14344_b1 , \14344_b0 , 
		\14345_b1 , \14345_b0 , \14346_b1 , \14346_b0 , \14347_b1 , \14347_b0 , \14348_b1 , \14348_b0 , \14349_b1 , \14349_b0 , 
		\14350_b1 , \14350_b0 , \14351_b1 , \14351_b0 , \14352_b1 , \14352_b0 , \14353_b1 , \14353_b0 , \14354_b1 , \14354_b0 , 
		\14355_b1 , \14355_b0 , \14356_b1 , \14356_b0 , \14357_b1 , \14357_b0 , \14358_b1 , \14358_b0 , \14359_b1 , \14359_b0 , 
		\14360_b1 , \14360_b0 , \14361_b1 , \14361_b0 , \14362_b1 , \14362_b0 , \14363_b1 , \14363_b0 , \14364_b1 , \14364_b0 , 
		\14365_b1 , \14365_b0 , \14366_b1 , \14366_b0 , \14367_b1 , \14367_b0 , \14368_b1 , \14368_b0 , \14369_b1 , \14369_b0 , 
		\14370_b1 , \14370_b0 , \14371_b1 , \14371_b0 , \14372_b1 , \14372_b0 , \14373_b1 , \14373_b0 , \14374_b1 , \14374_b0 , 
		\14375_b1 , \14375_b0 , \14376_b1 , \14376_b0 , \14377_b1 , \14377_b0 , \14378_b1 , \14378_b0 , \14379_b1 , \14379_b0 , 
		\14380_b1 , \14380_b0 , \14381_b1 , \14381_b0 , \14382_b1 , \14382_b0 , \14383_b1 , \14383_b0 , \14384_b1 , \14384_b0 , 
		\14385_b1 , \14385_b0 , \14386_b1 , \14386_b0 , \14387_b1 , \14387_b0 , \14388_b1 , \14388_b0 , \14389_b1 , \14389_b0 , 
		\14390_b1 , \14390_b0 , \14391_b1 , \14391_b0 , \14392_b1 , \14392_b0 , \14393_b1 , \14393_b0 , \14394_b1 , \14394_b0 , 
		\14395_b1 , \14395_b0 , \14396_b1 , \14396_b0 , \14397_b1 , \14397_b0 , \14398_b1 , \14398_b0 , \14399_b1 , \14399_b0 , 
		\14400_b1 , \14400_b0 , \14401_b1 , \14401_b0 , \14402_b1 , \14402_b0 , \14403_b1 , \14403_b0 , \14404_b1 , \14404_b0 , 
		\14405_b1 , \14405_b0 , \14406_b1 , \14406_b0 , \14407_b1 , \14407_b0 , \14408_b1 , \14408_b0 , \14409_b1 , \14409_b0 , 
		\14410_b1 , \14410_b0 , \14411_b1 , \14411_b0 , \14412_b1 , \14412_b0 , \14413_b1 , \14413_b0 , \14414_b1 , \14414_b0 , 
		\14415_b1 , \14415_b0 , \14416_b1 , \14416_b0 , \14417_b1 , \14417_b0 , \14418_b1 , \14418_b0 , \14419_b1 , \14419_b0 , 
		\14420_b1 , \14420_b0 , \14421_b1 , \14421_b0 , \14422_b1 , \14422_b0 , \14423_b1 , \14423_b0 , \14424_b1 , \14424_b0 , 
		\14425_b1 , \14425_b0 , \14426_b1 , \14426_b0 , \14427_b1 , \14427_b0 , \14428_b1 , \14428_b0 , \14429_b1 , \14429_b0 , 
		\14430_b1 , \14430_b0 , \14431_b1 , \14431_b0 , \14432_b1 , \14432_b0 , \14433_b1 , \14433_b0 , \14434_b1 , \14434_b0 , 
		\14435_b1 , \14435_b0 , \14436_b1 , \14436_b0 , \14437_b1 , \14437_b0 , \14438_b1 , \14438_b0 , \14439_b1 , \14439_b0 , 
		\14440_b1 , \14440_b0 , \14441_b1 , \14441_b0 , \14442_b1 , \14442_b0 , \14443_b1 , \14443_b0 , \14444_b1 , \14444_b0 , 
		\14445_b1 , \14445_b0 , \14446_b1 , \14446_b0 , \14447_b1 , \14447_b0 , \14448_b1 , \14448_b0 , \14449_b1 , \14449_b0 , 
		\14450_b1 , \14450_b0 , \14451_b1 , \14451_b0 , \14452_b1 , \14452_b0 , \14453_b1 , \14453_b0 , \14454_b1 , \14454_b0 , 
		\14455_b1 , \14455_b0 , \14456_b1 , \14456_b0 , \14457_b1 , \14457_b0 , \14458_b1 , \14458_b0 , \14459_b1 , \14459_b0 , 
		\14460_b1 , \14460_b0 , \14461_b1 , \14461_b0 , \14462_b1 , \14462_b0 , \14463_b1 , \14463_b0 , \14464_b1 , \14464_b0 , 
		\14465_b1 , \14465_b0 , \14466_b1 , \14466_b0 , \14467_b1 , \14467_b0 , \14468_b1 , \14468_b0 , \14469_b1 , \14469_b0 , 
		\14470_b1 , \14470_b0 , \14471_b1 , \14471_b0 , \14472_b1 , \14472_b0 , \14473_b1 , \14473_b0 , \14474_b1 , \14474_b0 , 
		\14475_b1 , \14475_b0 , \14476_b1 , \14476_b0 , \14477_b1 , \14477_b0 , \14478_b1 , \14478_b0 , \14479_b1 , \14479_b0 , 
		\14480_b1 , \14480_b0 , \14481_b1 , \14481_b0 , \14482_b1 , \14482_b0 , \14483_b1 , \14483_b0 , \14484_b1 , \14484_b0 , 
		\14485_b1 , \14485_b0 , \14486_b1 , \14486_b0 , \14487_b1 , \14487_b0 , \14488_b1 , \14488_b0 , \14489_b1 , \14489_b0 , 
		\14490_b1 , \14490_b0 , \14491_b1 , \14491_b0 , \14492_b1 , \14492_b0 , \14493_b1 , \14493_b0 , \14494_b1 , \14494_b0 , 
		\14495_b1 , \14495_b0 , \14496_b1 , \14496_b0 , \14497_b1 , \14497_b0 , \14498_b1 , \14498_b0 , \14499_b1 , \14499_b0 , 
		\14500_b1 , \14500_b0 , \14501_b1 , \14501_b0 , \14502_b1 , \14502_b0 , \14503_b1 , \14503_b0 , \14504_b1 , \14504_b0 , 
		\14505_b1 , \14505_b0 , \14506_b1 , \14506_b0 , \14507_b1 , \14507_b0 , \14508_b1 , \14508_b0 , \14509_b1 , \14509_b0 , 
		\14510_b1 , \14510_b0 , \14511_b1 , \14511_b0 , \14512_b1 , \14512_b0 , \14513_b1 , \14513_b0 , \14514_b1 , \14514_b0 , 
		\14515_b1 , \14515_b0 , \14516_b1 , \14516_b0 , \14517_b1 , \14517_b0 , \14518_b1 , \14518_b0 , \14519_b1 , \14519_b0 , 
		\14520_b1 , \14520_b0 , \14521_b1 , \14521_b0 , \14522_b1 , \14522_b0 , \14523_b1 , \14523_b0 , \14524_b1 , \14524_b0 , 
		\14525_b1 , \14525_b0 , \14526_b1 , \14526_b0 , \14527_b1 , \14527_b0 , \14528_b1 , \14528_b0 , \14529_b1 , \14529_b0 , 
		\14530_b1 , \14530_b0 , \14531_b1 , \14531_b0 , \14532_b1 , \14532_b0 , \14533_b1 , \14533_b0 , \14534_b1 , \14534_b0 , 
		\14535_b1 , \14535_b0 , \14536_b1 , \14536_b0 , \14537_b1 , \14537_b0 , \14538_b1 , \14538_b0 , \14539_b1 , \14539_b0 , 
		\14540_b1 , \14540_b0 , \14541_b1 , \14541_b0 , \14542_b1 , \14542_b0 , \14543_b1 , \14543_b0 , \14544_b1 , \14544_b0 , 
		\14545_b1 , \14545_b0 , \14546_b1 , \14546_b0 , \14547_b1 , \14547_b0 , \14548_b1 , \14548_b0 , \14549_b1 , \14549_b0 , 
		\14550_b1 , \14550_b0 , \14551_b1 , \14551_b0 , \14552_b1 , \14552_b0 , \14553_b1 , \14553_b0 , \14554_b1 , \14554_b0 , 
		\14555_b1 , \14555_b0 , \14556_b1 , \14556_b0 , \14557_b1 , \14557_b0 , \14558_b1 , \14558_b0 , \14559_b1 , \14559_b0 , 
		\14560_b1 , \14560_b0 , \14561_b1 , \14561_b0 , \14562_b1 , \14562_b0 , \14563_b1 , \14563_b0 , \14564_b1 , \14564_b0 , 
		\14565_b1 , \14565_b0 , \14566_b1 , \14566_b0 , \14567_b1 , \14567_b0 , \14568_b1 , \14568_b0 , \14569_b1 , \14569_b0 , 
		\14570_b1 , \14570_b0 , \14571_b1 , \14571_b0 , \14572_b1 , \14572_b0 , \14573_b1 , \14573_b0 , \14574_b1 , \14574_b0 , 
		\14575_b1 , \14575_b0 , \14576_b1 , \14576_b0 , \14577_b1 , \14577_b0 , \14578_b1 , \14578_b0 , \14579_b1 , \14579_b0 , 
		\14580_b1 , \14580_b0 , \14581_b1 , \14581_b0 , \14582_b1 , \14582_b0 , \14583_b1 , \14583_b0 , \14584_b1 , \14584_b0 , 
		\14585_b1 , \14585_b0 , \14586_b1 , \14586_b0 , \14587_b1 , \14587_b0 , \14588_b1 , \14588_b0 , \14589_b1 , \14589_b0 , 
		\14590_b1 , \14590_b0 , \14591_b1 , \14591_b0 , \14592_b1 , \14592_b0 , \14593_b1 , \14593_b0 , \14594_b1 , \14594_b0 , 
		\14595_b1 , \14595_b0 , \14596_b1 , \14596_b0 , \14597_b1 , \14597_b0 , \14598_b1 , \14598_b0 , \14599_b1 , \14599_b0 , 
		\14600_b1 , \14600_b0 , \14601_b1 , \14601_b0 , \14602_b1 , \14602_b0 , \14603_b1 , \14603_b0 , \14604_b1 , \14604_b0 , 
		\14605_b1 , \14605_b0 , \14606_b1 , \14606_b0 , \14607_b1 , \14607_b0 , \14608_b1 , \14608_b0 , \14609_b1 , \14609_b0 , 
		\14610_b1 , \14610_b0 , \14611_b1 , \14611_b0 , \14612_b1 , \14612_b0 , \14613_b1 , \14613_b0 , \14614_b1 , \14614_b0 , 
		\14615_b1 , \14615_b0 , \14616_b1 , \14616_b0 , \14617_b1 , \14617_b0 , \14618_b1 , \14618_b0 , \14619_b1 , \14619_b0 , 
		\14620_b1 , \14620_b0 , \14621_b1 , \14621_b0 , \14622_b1 , \14622_b0 , \14623_b1 , \14623_b0 , \14624_b1 , \14624_b0 , 
		\14625_b1 , \14625_b0 , \14626_b1 , \14626_b0 , \14627_b1 , \14627_b0 , \14628_b1 , \14628_b0 , \14629_b1 , \14629_b0 , 
		\14630_b1 , \14630_b0 , \14631_b1 , \14631_b0 , \14632_b1 , \14632_b0 , \14633_b1 , \14633_b0 , \14634_b1 , \14634_b0 , 
		\14635_b1 , \14635_b0 , \14636_b1 , \14636_b0 , \14637_b1 , \14637_b0 , \14638_b1 , \14638_b0 , \14639_b1 , \14639_b0 , 
		\14640_b1 , \14640_b0 , \14641_b1 , \14641_b0 , \14642_b1 , \14642_b0 , \14643_b1 , \14643_b0 , \14644_b1 , \14644_b0 , 
		\14645_b1 , \14645_b0 , \14646_b1 , \14646_b0 , \14647_b1 , \14647_b0 , \14648_b1 , \14648_b0 , \14649_b1 , \14649_b0 , 
		\14650_b1 , \14650_b0 , \14651_b1 , \14651_b0 , \14652_b1 , \14652_b0 , \14653_b1 , \14653_b0 , \14654_b1 , \14654_b0 , 
		\14655_b1 , \14655_b0 , \14656_b1 , \14656_b0 , \14657_b1 , \14657_b0 , \14658_b1 , \14658_b0 , \14659_b1 , \14659_b0 , 
		\14660_b1 , \14660_b0 , \14661_b1 , \14661_b0 , \14662_b1 , \14662_b0 , \14663_b1 , \14663_b0 , \14664_b1 , \14664_b0 , 
		\14665_b1 , \14665_b0 , \14666_b1 , \14666_b0 , \14667_b1 , \14667_b0 , \14668_b1 , \14668_b0 , \14669_b1 , \14669_b0 , 
		\14670_b1 , \14670_b0 , \14671_b1 , \14671_b0 , \14672_b1 , \14672_b0 , \14673_b1 , \14673_b0 , \14674_b1 , \14674_b0 , 
		\14675_b1 , \14675_b0 , \14676_b1 , \14676_b0 , \14677_b1 , \14677_b0 , \14678_b1 , \14678_b0 , \14679_b1 , \14679_b0 , 
		\14680_b1 , \14680_b0 , \14681_b1 , \14681_b0 , \14682_b1 , \14682_b0 , \14683_b1 , \14683_b0 , \14684_b1 , \14684_b0 , 
		\14685_b1 , \14685_b0 , \14686_b1 , \14686_b0 , \14687_b1 , \14687_b0 , \14688_b1 , \14688_b0 , \14689_b1 , \14689_b0 , 
		\14690_b1 , \14690_b0 , \14691_b1 , \14691_b0 , \14692_b1 , \14692_b0 , \14693_b1 , \14693_b0 , \14694_b1 , \14694_b0 , 
		\14695_b1 , \14695_b0 , \14696_b1 , \14696_b0 , \14697_b1 , \14697_b0 , \14698_b1 , \14698_b0 , \14699_b1 , \14699_b0 , 
		\14700_b1 , \14700_b0 , \14701_b1 , \14701_b0 , \14702_b1 , \14702_b0 , \14703_b1 , \14703_b0 , \14704_b1 , \14704_b0 , 
		\14705_b1 , \14705_b0 , \14706_b1 , \14706_b0 , \14707_b1 , \14707_b0 , \14708_b1 , \14708_b0 , \14709_b1 , \14709_b0 , 
		\14710_b1 , \14710_b0 , \14711_b1 , \14711_b0 , \14712_b1 , \14712_b0 , \14713_b1 , \14713_b0 , \14714_b1 , \14714_b0 , 
		\14715_b1 , \14715_b0 , \14716_b1 , \14716_b0 , \14717_b1 , \14717_b0 , \14718_b1 , \14718_b0 , \14719_b1 , \14719_b0 , 
		\14720_b1 , \14720_b0 , \14721_b1 , \14721_b0 , \14722_b1 , \14722_b0 , \14723_b1 , \14723_b0 , \14724_b1 , \14724_b0 , 
		\14725_b1 , \14725_b0 , \14726_b1 , \14726_b0 , \14727_b1 , \14727_b0 , \14728_b1 , \14728_b0 , \14729_b1 , \14729_b0 , 
		\14730_b1 , \14730_b0 , \14731_b1 , \14731_b0 , \14732_b1 , \14732_b0 , \14733_b1 , \14733_b0 , \14734_b1 , \14734_b0 , 
		\14735_b1 , \14735_b0 , \14736_b1 , \14736_b0 , \14737_b1 , \14737_b0 , \14738_b1 , \14738_b0 , \14739_b1 , \14739_b0 , 
		\14740_b1 , \14740_b0 , \14741_b1 , \14741_b0 , \14742_b1 , \14742_b0 , \14743_b1 , \14743_b0 , \14744_b1 , \14744_b0 , 
		\14745_b1 , \14745_b0 , \14746_b1 , \14746_b0 , \14747_b1 , \14747_b0 , \14748_b1 , \14748_b0 , \14749_b1 , \14749_b0 , 
		\14750_b1 , \14750_b0 , \14751_b1 , \14751_b0 , \14752_b1 , \14752_b0 , \14753_b1 , \14753_b0 , \14754_b1 , \14754_b0 , 
		\14755_b1 , \14755_b0 , \14756_b1 , \14756_b0 , \14757_b1 , \14757_b0 , \14758_b1 , \14758_b0 , \14759_b1 , \14759_b0 , 
		\14760_b1 , \14760_b0 , \14761_b1 , \14761_b0 , \14762_b1 , \14762_b0 , \14763_b1 , \14763_b0 , \14764_b1 , \14764_b0 , 
		\14765_b1 , \14765_b0 , \14766_b1 , \14766_b0 , \14767_b1 , \14767_b0 , \14768_b1 , \14768_b0 , \14769_b1 , \14769_b0 , 
		\14770_b1 , \14770_b0 , \14771_b1 , \14771_b0 , \14772_b1 , \14772_b0 , \14773_b1 , \14773_b0 , \14774_b1 , \14774_b0 , 
		\14775_b1 , \14775_b0 , \14776_b1 , \14776_b0 , \14777_b1 , \14777_b0 , \14778_b1 , \14778_b0 , \14779_b1 , \14779_b0 , 
		\14780_b1 , \14780_b0 , \14781_b1 , \14781_b0 , \14782_b1 , \14782_b0 , \14783_b1 , \14783_b0 , \14784_b1 , \14784_b0 , 
		\14785_b1 , \14785_b0 , \14786_b1 , \14786_b0 , \14787_b1 , \14787_b0 , \14788_b1 , \14788_b0 , \14789_b1 , \14789_b0 , 
		\14790_b1 , \14790_b0 , \14791_b1 , \14791_b0 , \14792_b1 , \14792_b0 , \14793_b1 , \14793_b0 , \14794_b1 , \14794_b0 , 
		\14795_b1 , \14795_b0 , \14796_b1 , \14796_b0 , \14797_b1 , \14797_b0 , \14798_b1 , \14798_b0 , \14799_b1 , \14799_b0 , 
		\14800_b1 , \14800_b0 , \14801_b1 , \14801_b0 , \14802_b1 , \14802_b0 , \14803_b1 , \14803_b0 , \14804_b1 , \14804_b0 , 
		\14805_b1 , \14805_b0 , \14806_b1 , \14806_b0 , \14807_b1 , \14807_b0 , \14808_b1 , \14808_b0 , \14809_b1 , \14809_b0 , 
		\14810_b1 , \14810_b0 , \14811_b1 , \14811_b0 , \14812_b1 , \14812_b0 , \14813_b1 , \14813_b0 , \14814_b1 , \14814_b0 , 
		\14815_b1 , \14815_b0 , \14816_b1 , \14816_b0 , \14817_b1 , \14817_b0 , \14818_b1 , \14818_b0 , \14819_b1 , \14819_b0 , 
		\14820_b1 , \14820_b0 , \14821_b1 , \14821_b0 , \14822_b1 , \14822_b0 , \14823_b1 , \14823_b0 , \14824_b1 , \14824_b0 , 
		\14825_b1 , \14825_b0 , \14826_b1 , \14826_b0 , \14827_b1 , \14827_b0 , \14828_b1 , \14828_b0 , \14829_b1 , \14829_b0 , 
		\14830_b1 , \14830_b0 , \14831_b1 , \14831_b0 , \14832_b1 , \14832_b0 , \14833_b1 , \14833_b0 , \14834_b1 , \14834_b0 , 
		\14835_b1 , \14835_b0 , \14836_b1 , \14836_b0 , \14837_b1 , \14837_b0 , \14838_b1 , \14838_b0 , \14839_b1 , \14839_b0 , 
		\14840_b1 , \14840_b0 , \14841_b1 , \14841_b0 , \14842_b1 , \14842_b0 , \14843_b1 , \14843_b0 , \14844_b1 , \14844_b0 , 
		\14845_b1 , \14845_b0 , \14846_b1 , \14846_b0 , \14847_b1 , \14847_b0 , \14848_b1 , \14848_b0 , \14849_b1 , \14849_b0 , 
		\14850_b1 , \14850_b0 , \14851_b1 , \14851_b0 , \14852_b1 , \14852_b0 , \14853_b1 , \14853_b0 , \14854_b1 , \14854_b0 , 
		\14855_b1 , \14855_b0 , \14856_b1 , \14856_b0 , \14857_b1 , \14857_b0 , \14858_b1 , \14858_b0 , \14859_b1 , \14859_b0 , 
		\14860_b1 , \14860_b0 , \14861_b1 , \14861_b0 , \14862_b1 , \14862_b0 , \14863_b1 , \14863_b0 , \14864_b1 , \14864_b0 , 
		\14865_b1 , \14865_b0 , \14866_b1 , \14866_b0 , \14867_b1 , \14867_b0 , \14868_b1 , \14868_b0 , \14869_b1 , \14869_b0 , 
		\14870_b1 , \14870_b0 , \14871_b1 , \14871_b0 , \14872_b1 , \14872_b0 , \14873_b1 , \14873_b0 , \14874_b1 , \14874_b0 , 
		\14875_b1 , \14875_b0 , \14876_b1 , \14876_b0 , \14877_b1 , \14877_b0 , \14878_b1 , \14878_b0 , \14879_b1 , \14879_b0 , 
		\14880_b1 , \14880_b0 , \14881_b1 , \14881_b0 , \14882_b1 , \14882_b0 , \14883_b1 , \14883_b0 , \14884_b1 , \14884_b0 , 
		\14885_b1 , \14885_b0 , \14886_b1 , \14886_b0 , \14887_b1 , \14887_b0 , \14888_b1 , \14888_b0 , \14889_b1 , \14889_b0 , 
		\14890_b1 , \14890_b0 , \14891_b1 , \14891_b0 , \14892_b1 , \14892_b0 , \14893_b1 , \14893_b0 , \14894_b1 , \14894_b0 , 
		\14895_b1 , \14895_b0 , \14896_b1 , \14896_b0 , \14897_b1 , \14897_b0 , \14898_b1 , \14898_b0 , \14899_b1 , \14899_b0 , 
		\14900_b1 , \14900_b0 , \14901_b1 , \14901_b0 , \14902_b1 , \14902_b0 , \14903_b1 , \14903_b0 , \14904_b1 , \14904_b0 , 
		\14905_b1 , \14905_b0 , \14906_b1 , \14906_b0 , \14907_b1 , \14907_b0 , \14908_b1 , \14908_b0 , \14909_b1 , \14909_b0 , 
		\14910_b1 , \14910_b0 , \14911_b1 , \14911_b0 , \14912_b1 , \14912_b0 , \14913_b1 , \14913_b0 , \14914_b1 , \14914_b0 , 
		\14915_b1 , \14915_b0 , \14916_b1 , \14916_b0 , \14917_b1 , \14917_b0 , \14918_b1 , \14918_b0 , \14919_b1 , \14919_b0 , 
		\14920_b1 , \14920_b0 , \14921_b1 , \14921_b0 , \14922_b1 , \14922_b0 , \14923_b1 , \14923_b0 , \14924_b1 , \14924_b0 , 
		\14925_b1 , \14925_b0 , \14926_b1 , \14926_b0 , \14927_b1 , \14927_b0 , \14928_b1 , \14928_b0 , \14929_b1 , \14929_b0 , 
		\14930_b1 , \14930_b0 , \14931_b1 , \14931_b0 , \14932_b1 , \14932_b0 , \14933_b1 , \14933_b0 , \14934_b1 , \14934_b0 , 
		\14935_b1 , \14935_b0 , \14936_b1 , \14936_b0 , \14937_b1 , \14937_b0 , \14938_b1 , \14938_b0 , \14939_b1 , \14939_b0 , 
		\14940_b1 , \14940_b0 , \14941_b1 , \14941_b0 , \14942_b1 , \14942_b0 , \14943_b1 , \14943_b0 , \14944_b1 , \14944_b0 , 
		\14945_b1 , \14945_b0 , \14946_b1 , \14946_b0 , \14947_b1 , \14947_b0 , \14948_b1 , \14948_b0 , \14949_b1 , \14949_b0 , 
		\14950_b1 , \14950_b0 , \14951_b1 , \14951_b0 , \14952_b1 , \14952_b0 , \14953_b1 , \14953_b0 , \14954_b1 , \14954_b0 , 
		\14955_b1 , \14955_b0 , \14956_b1 , \14956_b0 , \14957_b1 , \14957_b0 , \14958_b1 , \14958_b0 , \14959_b1 , \14959_b0 , 
		\14960_b1 , \14960_b0 , \14961_b1 , \14961_b0 , \14962_b1 , \14962_b0 , \14963_b1 , \14963_b0 , \14964_b1 , \14964_b0 , 
		\14965_b1 , \14965_b0 , \14966_b1 , \14966_b0 , \14967_b1 , \14967_b0 , \14968_b1 , \14968_b0 , \14969_b1 , \14969_b0 , 
		\14970_b1 , \14970_b0 , \14971_b1 , \14971_b0 , \14972_b1 , \14972_b0 , \14973_b1 , \14973_b0 , \14974_b1 , \14974_b0 , 
		\14975_b1 , \14975_b0 , \14976_b1 , \14976_b0 , \14977_b1 , \14977_b0 , \14978_b1 , \14978_b0 , \14979_b1 , \14979_b0 , 
		\14980_b1 , \14980_b0 , \14981_b1 , \14981_b0 , \14982_b1 , \14982_b0 , \14983_b1 , \14983_b0 , \14984_b1 , \14984_b0 , 
		\14985_b1 , \14985_b0 , \14986_b1 , \14986_b0 , \14987_b1 , \14987_b0 , \14988_b1 , \14988_b0 , \14989_b1 , \14989_b0 , 
		\14990_b1 , \14990_b0 , \14991_b1 , \14991_b0 , \14992_b1 , \14992_b0 , \14993_b1 , \14993_b0 , \14994_b1 , \14994_b0 , 
		\14995_b1 , \14995_b0 , \14996_b1 , \14996_b0 , \14997_b1 , \14997_b0 , \14998_b1 , \14998_b0 , \14999_b1 , \14999_b0 , 
		\15000_b1 , \15000_b0 , \15001_b1 , \15001_b0 , \15002_b1 , \15002_b0 , \15003_b1 , \15003_b0 , \15004_b1 , \15004_b0 , 
		\15005_b1 , \15005_b0 , \15006_b1 , \15006_b0 , \15007_b1 , \15007_b0 , \15008_b1 , \15008_b0 , \15009_b1 , \15009_b0 , 
		\15010_b1 , \15010_b0 , \15011_b1 , \15011_b0 , \15012_b1 , \15012_b0 , \15013_b1 , \15013_b0 , \15014_b1 , \15014_b0 , 
		\15015_b1 , \15015_b0 , \15016_b1 , \15016_b0 , \15017_b1 , \15017_b0 , \15018_b1 , \15018_b0 , \15019_b1 , \15019_b0 , 
		\15020_b1 , \15020_b0 , \15021_b1 , \15021_b0 , \15022_b1 , \15022_b0 , \15023_b1 , \15023_b0 , \15024_b1 , \15024_b0 , 
		\15025_b1 , \15025_b0 , \15026_b1 , \15026_b0 , \15027_b1 , \15027_b0 , \15028_b1 , \15028_b0 , \15029_b1 , \15029_b0 , 
		\15030_b1 , \15030_b0 , \15031_b1 , \15031_b0 , w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , 
		w_6 , w_7 , w_8 , w_9 , w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , 
		w_16 , w_17 , w_18 , w_19 , w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , 
		w_26 , w_27 , w_28 , w_29 , w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , 
		w_36 , w_37 , w_38 , w_39 , w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , 
		w_46 , w_47 , w_48 , w_49 , w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , 
		w_56 , w_57 , w_58 , w_59 , w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , 
		w_66 , w_67 , w_68 , w_69 , w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , 
		w_76 , w_77 , w_78 , w_79 , w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , 
		w_86 , w_87 , w_88 , w_89 , w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , 
		w_96 , w_97 , w_98 , w_99 , w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , 
		w_106 , w_107 , w_108 , w_109 , w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , 
		w_116 , w_117 , w_118 , w_119 , w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , 
		w_126 , w_127 , w_128 , w_129 , w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , 
		w_136 , w_137 , w_138 , w_139 , w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , 
		w_146 , w_147 , w_148 , w_149 , w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , 
		w_156 , w_157 , w_158 , w_159 , w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , 
		w_166 , w_167 , w_168 , w_169 , w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , 
		w_176 , w_177 , w_178 , w_179 , w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , 
		w_186 , w_187 , w_188 , w_189 , w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , 
		w_196 , w_197 , w_198 , w_199 , w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , 
		w_206 , w_207 , w_208 , w_209 , w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , 
		w_216 , w_217 , w_218 , w_219 , w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , 
		w_226 , w_227 , w_228 , w_229 , w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , 
		w_236 , w_237 , w_238 , w_239 , w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , 
		w_246 , w_247 , w_248 , w_249 , w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , 
		w_256 , w_257 , w_258 , w_259 , w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , 
		w_266 , w_267 , w_268 , w_269 , w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , 
		w_276 , w_277 , w_278 , w_279 , w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , 
		w_286 , w_287 , w_288 , w_289 , w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , 
		w_296 , w_297 , w_298 , w_299 , w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , 
		w_306 , w_307 , w_308 , w_309 , w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , 
		w_316 , w_317 , w_318 , w_319 , w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , 
		w_326 , w_327 , w_328 , w_329 , w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , 
		w_336 , w_337 , w_338 , w_339 , w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , 
		w_346 , w_347 , w_348 , w_349 , w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , 
		w_356 , w_357 , w_358 , w_359 , w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , 
		w_366 , w_367 , w_368 , w_369 , w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , 
		w_376 , w_377 , w_378 , w_379 , w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , 
		w_386 , w_387 , w_388 , w_389 , w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , 
		w_396 , w_397 , w_398 , w_399 , w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , 
		w_406 , w_407 , w_408 , w_409 , w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , 
		w_416 , w_417 , w_418 , w_419 , w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , 
		w_426 , w_427 , w_428 , w_429 , w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , 
		w_436 , w_437 , w_438 , w_439 , w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , 
		w_446 , w_447 , w_448 , w_449 , w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , 
		w_456 , w_457 , w_458 , w_459 , w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , 
		w_466 , w_467 , w_468 , w_469 , w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , 
		w_476 , w_477 , w_478 , w_479 , w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , 
		w_486 , w_487 , w_488 , w_489 , w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , 
		w_496 , w_497 , w_498 , w_499 , w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , 
		w_506 , w_507 , w_508 , w_509 , w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , 
		w_516 , w_517 , w_518 , w_519 , w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , 
		w_526 , w_527 , w_528 , w_529 , w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , 
		w_536 , w_537 , w_538 , w_539 , w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , 
		w_546 , w_547 , w_548 , w_549 , w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , 
		w_556 , w_557 , w_558 , w_559 , w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , 
		w_566 , w_567 , w_568 , w_569 , w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , 
		w_576 , w_577 , w_578 , w_579 , w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , 
		w_586 , w_587 , w_588 , w_589 , w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , 
		w_596 , w_597 , w_598 , w_599 , w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , 
		w_606 , w_607 , w_608 , w_609 , w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , 
		w_616 , w_617 , w_618 , w_619 , w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , 
		w_626 , w_627 , w_628 , w_629 , w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , 
		w_636 , w_637 , w_638 , w_639 , w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , 
		w_646 , w_647 , w_648 , w_649 , w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , 
		w_656 , w_657 , w_658 , w_659 , w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , 
		w_666 , w_667 , w_668 , w_669 , w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , 
		w_676 , w_677 , w_678 , w_679 , w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , 
		w_686 , w_687 , w_688 , w_689 , w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , 
		w_696 , w_697 , w_698 , w_699 , w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , 
		w_706 , w_707 , w_708 , w_709 , w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , 
		w_716 , w_717 , w_718 , w_719 , w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , 
		w_726 , w_727 , w_728 , w_729 , w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , 
		w_736 , w_737 , w_738 , w_739 , w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , 
		w_746 , w_747 , w_748 , w_749 , w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , 
		w_756 , w_757 , w_758 , w_759 , w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , 
		w_766 , w_767 , w_768 , w_769 , w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , 
		w_776 , w_777 , w_778 , w_779 , w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , 
		w_786 , w_787 , w_788 , w_789 , w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , 
		w_796 , w_797 , w_798 , w_799 , w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , 
		w_806 , w_807 , w_808 , w_809 , w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , 
		w_816 , w_817 , w_818 , w_819 , w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , 
		w_826 , w_827 , w_828 , w_829 , w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , 
		w_836 , w_837 , w_838 , w_839 , w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , 
		w_846 , w_847 , w_848 , w_849 , w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , 
		w_856 , w_857 , w_858 , w_859 , w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , 
		w_866 , w_867 , w_868 , w_869 , w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , 
		w_876 , w_877 , w_878 , w_879 , w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , 
		w_886 , w_887 , w_888 , w_889 , w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , 
		w_896 , w_897 , w_898 , w_899 , w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , 
		w_906 , w_907 , w_908 , w_909 , w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , 
		w_916 , w_917 , w_918 , w_919 , w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , 
		w_926 , w_927 , w_928 , w_929 , w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , 
		w_936 , w_937 , w_938 , w_939 , w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , 
		w_946 , w_947 , w_948 , w_949 , w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , 
		w_956 , w_957 , w_958 , w_959 , w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , 
		w_966 , w_967 , w_968 , w_969 , w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , 
		w_976 , w_977 , w_978 , w_979 , w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , 
		w_986 , w_987 , w_988 , w_989 , w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , 
		w_996 , w_997 , w_998 , w_999 , w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , 
		w_1006 , w_1007 , w_1008 , w_1009 , w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , 
		w_1016 , w_1017 , w_1018 , w_1019 , w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , 
		w_1026 , w_1027 , w_1028 , w_1029 , w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , 
		w_1036 , w_1037 , w_1038 , w_1039 , w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , 
		w_1046 , w_1047 , w_1048 , w_1049 , w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , 
		w_1056 , w_1057 , w_1058 , w_1059 , w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , 
		w_1066 , w_1067 , w_1068 , w_1069 , w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , 
		w_1076 , w_1077 , w_1078 , w_1079 , w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , 
		w_1086 , w_1087 , w_1088 , w_1089 , w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , 
		w_1096 , w_1097 , w_1098 , w_1099 , w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , 
		w_1106 , w_1107 , w_1108 , w_1109 , w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , 
		w_1116 , w_1117 , w_1118 , w_1119 , w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , 
		w_1126 , w_1127 , w_1128 , w_1129 , w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , 
		w_1136 , w_1137 , w_1138 , w_1139 , w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , 
		w_1146 , w_1147 , w_1148 , w_1149 , w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , 
		w_1156 , w_1157 , w_1158 , w_1159 , w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , 
		w_1166 , w_1167 , w_1168 , w_1169 , w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , 
		w_1176 , w_1177 , w_1178 , w_1179 , w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , 
		w_1186 , w_1187 , w_1188 , w_1189 , w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , 
		w_1196 , w_1197 , w_1198 , w_1199 , w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , 
		w_1206 , w_1207 , w_1208 , w_1209 , w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , 
		w_1216 , w_1217 , w_1218 , w_1219 , w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , 
		w_1226 , w_1227 , w_1228 , w_1229 , w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , 
		w_1236 , w_1237 , w_1238 , w_1239 , w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , 
		w_1246 , w_1247 , w_1248 , w_1249 , w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , 
		w_1256 , w_1257 , w_1258 , w_1259 , w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , 
		w_1266 , w_1267 , w_1268 , w_1269 , w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , 
		w_1276 , w_1277 , w_1278 , w_1279 , w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , 
		w_1286 , w_1287 , w_1288 , w_1289 , w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , 
		w_1296 , w_1297 , w_1298 , w_1299 , w_1300 , w_1301 , w_1302 , w_1303 , w_1304 , w_1305 , 
		w_1306 , w_1307 , w_1308 , w_1309 , w_1310 , w_1311 , w_1312 , w_1313 , w_1314 , w_1315 , 
		w_1316 , w_1317 , w_1318 , w_1319 , w_1320 , w_1321 , w_1322 , w_1323 , w_1324 , w_1325 , 
		w_1326 , w_1327 , w_1328 , w_1329 , w_1330 , w_1331 , w_1332 , w_1333 , w_1334 , w_1335 , 
		w_1336 , w_1337 , w_1338 , w_1339 , w_1340 , w_1341 , w_1342 , w_1343 , w_1344 , w_1345 , 
		w_1346 , w_1347 , w_1348 , w_1349 , w_1350 , w_1351 , w_1352 , w_1353 , w_1354 , w_1355 , 
		w_1356 , w_1357 , w_1358 , w_1359 , w_1360 , w_1361 , w_1362 , w_1363 , w_1364 , w_1365 , 
		w_1366 , w_1367 , w_1368 , w_1369 , w_1370 , w_1371 , w_1372 , w_1373 , w_1374 , w_1375 , 
		w_1376 , w_1377 , w_1378 , w_1379 , w_1380 , w_1381 , w_1382 , w_1383 , w_1384 , w_1385 , 
		w_1386 , w_1387 , w_1388 , w_1389 , w_1390 , w_1391 , w_1392 , w_1393 , w_1394 , w_1395 , 
		w_1396 , w_1397 , w_1398 , w_1399 , w_1400 , w_1401 , w_1402 , w_1403 , w_1404 , w_1405 , 
		w_1406 , w_1407 , w_1408 , w_1409 , w_1410 , w_1411 , w_1412 , w_1413 , w_1414 , w_1415 , 
		w_1416 , w_1417 , w_1418 , w_1419 , w_1420 , w_1421 , w_1422 , w_1423 , w_1424 , w_1425 , 
		w_1426 , w_1427 , w_1428 , w_1429 , w_1430 , w_1431 , w_1432 , w_1433 , w_1434 , w_1435 , 
		w_1436 , w_1437 , w_1438 , w_1439 , w_1440 , w_1441 , w_1442 , w_1443 , w_1444 , w_1445 , 
		w_1446 , w_1447 , w_1448 , w_1449 , w_1450 , w_1451 , w_1452 , w_1453 , w_1454 , w_1455 , 
		w_1456 , w_1457 , w_1458 , w_1459 , w_1460 , w_1461 , w_1462 , w_1463 , w_1464 , w_1465 , 
		w_1466 , w_1467 , w_1468 , w_1469 , w_1470 , w_1471 , w_1472 , w_1473 , w_1474 , w_1475 , 
		w_1476 , w_1477 , w_1478 , w_1479 , w_1480 , w_1481 , w_1482 , w_1483 , w_1484 , w_1485 , 
		w_1486 , w_1487 , w_1488 , w_1489 , w_1490 , w_1491 , w_1492 , w_1493 , w_1494 , w_1495 , 
		w_1496 , w_1497 , w_1498 , w_1499 , w_1500 , w_1501 , w_1502 , w_1503 , w_1504 , w_1505 , 
		w_1506 , w_1507 , w_1508 , w_1509 , w_1510 , w_1511 , w_1512 , w_1513 , w_1514 , w_1515 , 
		w_1516 , w_1517 , w_1518 , w_1519 , w_1520 , w_1521 , w_1522 , w_1523 , w_1524 , w_1525 , 
		w_1526 , w_1527 , w_1528 , w_1529 , w_1530 , w_1531 , w_1532 , w_1533 , w_1534 , w_1535 , 
		w_1536 , w_1537 , w_1538 , w_1539 , w_1540 , w_1541 , w_1542 , w_1543 , w_1544 , w_1545 , 
		w_1546 , w_1547 , w_1548 , w_1549 , w_1550 , w_1551 , w_1552 , w_1553 , w_1554 , w_1555 , 
		w_1556 , w_1557 , w_1558 , w_1559 , w_1560 , w_1561 , w_1562 , w_1563 , w_1564 , w_1565 , 
		w_1566 , w_1567 , w_1568 , w_1569 , w_1570 , w_1571 , w_1572 , w_1573 , w_1574 , w_1575 , 
		w_1576 , w_1577 , w_1578 , w_1579 , w_1580 , w_1581 , w_1582 , w_1583 , w_1584 , w_1585 , 
		w_1586 , w_1587 , w_1588 , w_1589 , w_1590 , w_1591 , w_1592 , w_1593 , w_1594 , w_1595 , 
		w_1596 , w_1597 , w_1598 , w_1599 , w_1600 , w_1601 , w_1602 , w_1603 , w_1604 , w_1605 , 
		w_1606 , w_1607 , w_1608 , w_1609 , w_1610 , w_1611 , w_1612 , w_1613 , w_1614 , w_1615 , 
		w_1616 , w_1617 , w_1618 , w_1619 , w_1620 , w_1621 , w_1622 , w_1623 , w_1624 , w_1625 , 
		w_1626 , w_1627 , w_1628 , w_1629 , w_1630 , w_1631 , w_1632 , w_1633 , w_1634 , w_1635 , 
		w_1636 , w_1637 , w_1638 , w_1639 , w_1640 , w_1641 , w_1642 , w_1643 , w_1644 , w_1645 , 
		w_1646 , w_1647 , w_1648 , w_1649 , w_1650 , w_1651 , w_1652 , w_1653 , w_1654 , w_1655 , 
		w_1656 , w_1657 , w_1658 , w_1659 , w_1660 , w_1661 , w_1662 , w_1663 , w_1664 , w_1665 , 
		w_1666 , w_1667 , w_1668 , w_1669 , w_1670 , w_1671 , w_1672 , w_1673 , w_1674 , w_1675 , 
		w_1676 , w_1677 , w_1678 , w_1679 , w_1680 , w_1681 , w_1682 , w_1683 , w_1684 , w_1685 , 
		w_1686 , w_1687 , w_1688 , w_1689 , w_1690 , w_1691 , w_1692 , w_1693 , w_1694 , w_1695 , 
		w_1696 , w_1697 , w_1698 , w_1699 , w_1700 , w_1701 , w_1702 , w_1703 , w_1704 , w_1705 , 
		w_1706 , w_1707 , w_1708 , w_1709 , w_1710 , w_1711 , w_1712 , w_1713 , w_1714 , w_1715 , 
		w_1716 , w_1717 , w_1718 , w_1719 , w_1720 , w_1721 , w_1722 , w_1723 , w_1724 , w_1725 , 
		w_1726 , w_1727 , w_1728 , w_1729 , w_1730 , w_1731 , w_1732 , w_1733 , w_1734 , w_1735 , 
		w_1736 , w_1737 , w_1738 , w_1739 , w_1740 , w_1741 , w_1742 , w_1743 , w_1744 , w_1745 , 
		w_1746 , w_1747 , w_1748 , w_1749 , w_1750 , w_1751 , w_1752 , w_1753 , w_1754 , w_1755 , 
		w_1756 , w_1757 , w_1758 , w_1759 , w_1760 , w_1761 , w_1762 , w_1763 , w_1764 , w_1765 , 
		w_1766 , w_1767 , w_1768 , w_1769 , w_1770 , w_1771 , w_1772 , w_1773 , w_1774 , w_1775 , 
		w_1776 , w_1777 , w_1778 , w_1779 , w_1780 , w_1781 , w_1782 , w_1783 , w_1784 , w_1785 , 
		w_1786 , w_1787 , w_1788 , w_1789 , w_1790 , w_1791 , w_1792 , w_1793 , w_1794 , w_1795 , 
		w_1796 , w_1797 , w_1798 , w_1799 , w_1800 , w_1801 , w_1802 , w_1803 , w_1804 , w_1805 , 
		w_1806 , w_1807 , w_1808 , w_1809 , w_1810 , w_1811 , w_1812 , w_1813 , w_1814 , w_1815 , 
		w_1816 , w_1817 , w_1818 , w_1819 , w_1820 , w_1821 , w_1822 , w_1823 , w_1824 , w_1825 , 
		w_1826 , w_1827 , w_1828 , w_1829 , w_1830 , w_1831 , w_1832 , w_1833 , w_1834 , w_1835 , 
		w_1836 , w_1837 , w_1838 , w_1839 , w_1840 , w_1841 , w_1842 , w_1843 , w_1844 , w_1845 , 
		w_1846 , w_1847 , w_1848 , w_1849 , w_1850 , w_1851 , w_1852 , w_1853 , w_1854 , w_1855 , 
		w_1856 , w_1857 , w_1858 , w_1859 , w_1860 , w_1861 , w_1862 , w_1863 , w_1864 , w_1865 , 
		w_1866 , w_1867 , w_1868 , w_1869 , w_1870 , w_1871 , w_1872 , w_1873 , w_1874 , w_1875 , 
		w_1876 , w_1877 , w_1878 , w_1879 , w_1880 , w_1881 , w_1882 , w_1883 , w_1884 , w_1885 , 
		w_1886 , w_1887 , w_1888 , w_1889 , w_1890 , w_1891 , w_1892 , w_1893 , w_1894 , w_1895 , 
		w_1896 , w_1897 , w_1898 , w_1899 , w_1900 , w_1901 , w_1902 , w_1903 , w_1904 , w_1905 , 
		w_1906 , w_1907 , w_1908 , w_1909 , w_1910 , w_1911 , w_1912 , w_1913 , w_1914 , w_1915 , 
		w_1916 , w_1917 , w_1918 , w_1919 , w_1920 , w_1921 , w_1922 , w_1923 , w_1924 , w_1925 , 
		w_1926 , w_1927 , w_1928 , w_1929 , w_1930 , w_1931 , w_1932 , w_1933 , w_1934 , w_1935 , 
		w_1936 , w_1937 , w_1938 , w_1939 , w_1940 , w_1941 , w_1942 , w_1943 , w_1944 , w_1945 , 
		w_1946 , w_1947 , w_1948 , w_1949 , w_1950 , w_1951 , w_1952 , w_1953 , w_1954 , w_1955 , 
		w_1956 , w_1957 , w_1958 , w_1959 , w_1960 , w_1961 , w_1962 , w_1963 , w_1964 , w_1965 , 
		w_1966 , w_1967 , w_1968 , w_1969 , w_1970 , w_1971 , w_1972 , w_1973 , w_1974 , w_1975 , 
		w_1976 , w_1977 , w_1978 , w_1979 , w_1980 , w_1981 , w_1982 , w_1983 , w_1984 , w_1985 , 
		w_1986 , w_1987 , w_1988 , w_1989 , w_1990 , w_1991 , w_1992 , w_1993 , w_1994 , w_1995 , 
		w_1996 , w_1997 , w_1998 , w_1999 , w_2000 , w_2001 , w_2002 , w_2003 , w_2004 , w_2005 , 
		w_2006 , w_2007 , w_2008 , w_2009 , w_2010 , w_2011 , w_2012 , w_2013 , w_2014 , w_2015 , 
		w_2016 , w_2017 , w_2018 , w_2019 , w_2020 , w_2021 , w_2022 , w_2023 , w_2024 , w_2025 , 
		w_2026 , w_2027 , w_2028 , w_2029 , w_2030 , w_2031 , w_2032 , w_2033 , w_2034 , w_2035 , 
		w_2036 , w_2037 , w_2038 , w_2039 , w_2040 , w_2041 , w_2042 , w_2043 , w_2044 , w_2045 , 
		w_2046 , w_2047 , w_2048 , w_2049 , w_2050 , w_2051 , w_2052 , w_2053 , w_2054 , w_2055 , 
		w_2056 , w_2057 , w_2058 , w_2059 , w_2060 , w_2061 , w_2062 , w_2063 , w_2064 , w_2065 , 
		w_2066 , w_2067 , w_2068 , w_2069 , w_2070 , w_2071 , w_2072 , w_2073 , w_2074 , w_2075 , 
		w_2076 , w_2077 , w_2078 , w_2079 , w_2080 , w_2081 , w_2082 , w_2083 , w_2084 , w_2085 , 
		w_2086 , w_2087 , w_2088 , w_2089 , w_2090 , w_2091 , w_2092 , w_2093 , w_2094 , w_2095 , 
		w_2096 , w_2097 , w_2098 , w_2099 , w_2100 , w_2101 , w_2102 , w_2103 , w_2104 , w_2105 , 
		w_2106 , w_2107 , w_2108 , w_2109 , w_2110 , w_2111 , w_2112 , w_2113 , w_2114 , w_2115 , 
		w_2116 , w_2117 , w_2118 , w_2119 , w_2120 , w_2121 , w_2122 , w_2123 , w_2124 , w_2125 , 
		w_2126 , w_2127 , w_2128 , w_2129 , w_2130 , w_2131 , w_2132 , w_2133 , w_2134 , w_2135 , 
		w_2136 , w_2137 , w_2138 , w_2139 , w_2140 , w_2141 , w_2142 , w_2143 , w_2144 , w_2145 , 
		w_2146 , w_2147 , w_2148 , w_2149 , w_2150 , w_2151 , w_2152 , w_2153 , w_2154 , w_2155 , 
		w_2156 , w_2157 , w_2158 , w_2159 , w_2160 , w_2161 , w_2162 , w_2163 , w_2164 , w_2165 , 
		w_2166 , w_2167 , w_2168 , w_2169 , w_2170 , w_2171 , w_2172 , w_2173 , w_2174 , w_2175 , 
		w_2176 , w_2177 , w_2178 , w_2179 , w_2180 , w_2181 , w_2182 , w_2183 , w_2184 , w_2185 , 
		w_2186 , w_2187 , w_2188 , w_2189 , w_2190 , w_2191 , w_2192 , w_2193 , w_2194 , w_2195 , 
		w_2196 , w_2197 , w_2198 , w_2199 , w_2200 , w_2201 , w_2202 , w_2203 , w_2204 , w_2205 , 
		w_2206 , w_2207 , w_2208 , w_2209 , w_2210 , w_2211 , w_2212 , w_2213 , w_2214 , w_2215 , 
		w_2216 , w_2217 , w_2218 , w_2219 , w_2220 , w_2221 , w_2222 , w_2223 , w_2224 , w_2225 , 
		w_2226 , w_2227 , w_2228 , w_2229 , w_2230 , w_2231 , w_2232 , w_2233 , w_2234 , w_2235 , 
		w_2236 , w_2237 , w_2238 , w_2239 , w_2240 , w_2241 , w_2242 , w_2243 , w_2244 , w_2245 , 
		w_2246 , w_2247 , w_2248 , w_2249 , w_2250 , w_2251 , w_2252 , w_2253 , w_2254 , w_2255 , 
		w_2256 , w_2257 , w_2258 , w_2259 , w_2260 , w_2261 , w_2262 , w_2263 , w_2264 , w_2265 , 
		w_2266 , w_2267 , w_2268 , w_2269 , w_2270 , w_2271 , w_2272 , w_2273 , w_2274 , w_2275 , 
		w_2276 , w_2277 , w_2278 , w_2279 , w_2280 , w_2281 , w_2282 , w_2283 , w_2284 , w_2285 , 
		w_2286 , w_2287 , w_2288 , w_2289 , w_2290 , w_2291 , w_2292 , w_2293 , w_2294 , w_2295 , 
		w_2296 , w_2297 , w_2298 , w_2299 , w_2300 , w_2301 , w_2302 , w_2303 , w_2304 , w_2305 , 
		w_2306 , w_2307 , w_2308 , w_2309 , w_2310 , w_2311 , w_2312 , w_2313 , w_2314 , w_2315 , 
		w_2316 , w_2317 , w_2318 , w_2319 , w_2320 , w_2321 , w_2322 , w_2323 , w_2324 , w_2325 , 
		w_2326 , w_2327 , w_2328 , w_2329 , w_2330 , w_2331 , w_2332 , w_2333 , w_2334 , w_2335 , 
		w_2336 , w_2337 , w_2338 , w_2339 , w_2340 , w_2341 , w_2342 , w_2343 , w_2344 , w_2345 , 
		w_2346 , w_2347 , w_2348 , w_2349 , w_2350 , w_2351 , w_2352 , w_2353 , w_2354 , w_2355 , 
		w_2356 , w_2357 , w_2358 , w_2359 , w_2360 , w_2361 , w_2362 , w_2363 , w_2364 , w_2365 , 
		w_2366 , w_2367 , w_2368 , w_2369 , w_2370 , w_2371 , w_2372 , w_2373 , w_2374 , w_2375 , 
		w_2376 , w_2377 , w_2378 , w_2379 , w_2380 , w_2381 , w_2382 , w_2383 , w_2384 , w_2385 , 
		w_2386 , w_2387 , w_2388 , w_2389 , w_2390 , w_2391 , w_2392 , w_2393 , w_2394 , w_2395 , 
		w_2396 , w_2397 , w_2398 , w_2399 , w_2400 , w_2401 , w_2402 , w_2403 , w_2404 , w_2405 , 
		w_2406 , w_2407 , w_2408 , w_2409 , w_2410 , w_2411 , w_2412 , w_2413 , w_2414 , w_2415 , 
		w_2416 , w_2417 , w_2418 , w_2419 , w_2420 , w_2421 , w_2422 , w_2423 , w_2424 , w_2425 , 
		w_2426 , w_2427 , w_2428 , w_2429 , w_2430 , w_2431 , w_2432 , w_2433 , w_2434 , w_2435 , 
		w_2436 , w_2437 , w_2438 , w_2439 , w_2440 , w_2441 , w_2442 , w_2443 , w_2444 , w_2445 , 
		w_2446 , w_2447 , w_2448 , w_2449 , w_2450 , w_2451 , w_2452 , w_2453 , w_2454 , w_2455 , 
		w_2456 , w_2457 , w_2458 , w_2459 , w_2460 , w_2461 , w_2462 , w_2463 , w_2464 , w_2465 , 
		w_2466 , w_2467 , w_2468 , w_2469 , w_2470 , w_2471 , w_2472 , w_2473 , w_2474 , w_2475 , 
		w_2476 , w_2477 , w_2478 , w_2479 , w_2480 , w_2481 , w_2482 , w_2483 , w_2484 , w_2485 , 
		w_2486 , w_2487 , w_2488 , w_2489 , w_2490 , w_2491 , w_2492 , w_2493 , w_2494 , w_2495 , 
		w_2496 , w_2497 , w_2498 , w_2499 , w_2500 , w_2501 , w_2502 , w_2503 , w_2504 , w_2505 , 
		w_2506 , w_2507 , w_2508 , w_2509 , w_2510 , w_2511 , w_2512 , w_2513 , w_2514 , w_2515 , 
		w_2516 , w_2517 , w_2518 , w_2519 , w_2520 , w_2521 , w_2522 , w_2523 , w_2524 , w_2525 , 
		w_2526 , w_2527 , w_2528 , w_2529 , w_2530 , w_2531 , w_2532 , w_2533 , w_2534 , w_2535 , 
		w_2536 , w_2537 , w_2538 , w_2539 , w_2540 , w_2541 , w_2542 , w_2543 , w_2544 , w_2545 , 
		w_2546 , w_2547 , w_2548 , w_2549 , w_2550 , w_2551 , w_2552 , w_2553 , w_2554 , w_2555 , 
		w_2556 , w_2557 , w_2558 , w_2559 , w_2560 , w_2561 , w_2562 , w_2563 , w_2564 , w_2565 , 
		w_2566 , w_2567 , w_2568 , w_2569 , w_2570 , w_2571 , w_2572 , w_2573 , w_2574 , w_2575 , 
		w_2576 , w_2577 , w_2578 , w_2579 , w_2580 , w_2581 , w_2582 , w_2583 , w_2584 , w_2585 , 
		w_2586 , w_2587 , w_2588 , w_2589 , w_2590 , w_2591 , w_2592 , w_2593 , w_2594 , w_2595 , 
		w_2596 , w_2597 , w_2598 , w_2599 , w_2600 , w_2601 , w_2602 , w_2603 , w_2604 , w_2605 , 
		w_2606 , w_2607 , w_2608 , w_2609 , w_2610 , w_2611 , w_2612 , w_2613 , w_2614 , w_2615 , 
		w_2616 , w_2617 , w_2618 , w_2619 , w_2620 , w_2621 , w_2622 , w_2623 , w_2624 , w_2625 , 
		w_2626 , w_2627 , w_2628 , w_2629 , w_2630 , w_2631 , w_2632 , w_2633 , w_2634 , w_2635 , 
		w_2636 , w_2637 , w_2638 , w_2639 , w_2640 , w_2641 , w_2642 , w_2643 , w_2644 , w_2645 , 
		w_2646 , w_2647 , w_2648 , w_2649 , w_2650 , w_2651 , w_2652 , w_2653 , w_2654 , w_2655 , 
		w_2656 , w_2657 , w_2658 , w_2659 , w_2660 , w_2661 , w_2662 , w_2663 , w_2664 , w_2665 , 
		w_2666 , w_2667 , w_2668 , w_2669 , w_2670 , w_2671 , w_2672 , w_2673 , w_2674 , w_2675 , 
		w_2676 , w_2677 , w_2678 , w_2679 , w_2680 , w_2681 , w_2682 , w_2683 , w_2684 , w_2685 , 
		w_2686 , w_2687 , w_2688 , w_2689 , w_2690 , w_2691 , w_2692 , w_2693 , w_2694 , w_2695 , 
		w_2696 , w_2697 , w_2698 , w_2699 , w_2700 , w_2701 , w_2702 , w_2703 , w_2704 , w_2705 , 
		w_2706 , w_2707 , w_2708 , w_2709 , w_2710 , w_2711 , w_2712 , w_2713 , w_2714 , w_2715 , 
		w_2716 , w_2717 , w_2718 , w_2719 , w_2720 , w_2721 , w_2722 , w_2723 , w_2724 , w_2725 , 
		w_2726 , w_2727 , w_2728 , w_2729 , w_2730 , w_2731 , w_2732 , w_2733 , w_2734 , w_2735 , 
		w_2736 , w_2737 , w_2738 , w_2739 , w_2740 , w_2741 , w_2742 , w_2743 , w_2744 , w_2745 , 
		w_2746 , w_2747 , w_2748 , w_2749 , w_2750 , w_2751 , w_2752 , w_2753 , w_2754 , w_2755 , 
		w_2756 , w_2757 , w_2758 , w_2759 , w_2760 , w_2761 , w_2762 , w_2763 , w_2764 , w_2765 , 
		w_2766 , w_2767 , w_2768 , w_2769 , w_2770 , w_2771 , w_2772 , w_2773 , w_2774 , w_2775 , 
		w_2776 , w_2777 , w_2778 , w_2779 , w_2780 , w_2781 , w_2782 , w_2783 , w_2784 , w_2785 , 
		w_2786 , w_2787 , w_2788 , w_2789 , w_2790 , w_2791 , w_2792 , w_2793 , w_2794 , w_2795 , 
		w_2796 , w_2797 , w_2798 , w_2799 , w_2800 , w_2801 , w_2802 , w_2803 , w_2804 , w_2805 , 
		w_2806 , w_2807 , w_2808 , w_2809 , w_2810 , w_2811 , w_2812 , w_2813 , w_2814 , w_2815 , 
		w_2816 , w_2817 , w_2818 , w_2819 , w_2820 , w_2821 , w_2822 , w_2823 , w_2824 , w_2825 , 
		w_2826 , w_2827 , w_2828 , w_2829 , w_2830 , w_2831 , w_2832 , w_2833 , w_2834 , w_2835 , 
		w_2836 , w_2837 , w_2838 , w_2839 , w_2840 , w_2841 , w_2842 , w_2843 , w_2844 , w_2845 , 
		w_2846 , w_2847 , w_2848 , w_2849 , w_2850 , w_2851 , w_2852 , w_2853 , w_2854 , w_2855 , 
		w_2856 , w_2857 , w_2858 , w_2859 , w_2860 , w_2861 , w_2862 , w_2863 , w_2864 , w_2865 , 
		w_2866 , w_2867 , w_2868 , w_2869 , w_2870 , w_2871 , w_2872 , w_2873 , w_2874 , w_2875 , 
		w_2876 , w_2877 , w_2878 , w_2879 , w_2880 , w_2881 , w_2882 , w_2883 , w_2884 , w_2885 , 
		w_2886 , w_2887 , w_2888 , w_2889 , w_2890 , w_2891 , w_2892 , w_2893 , w_2894 , w_2895 , 
		w_2896 , w_2897 , w_2898 , w_2899 , w_2900 , w_2901 , w_2902 , w_2903 , w_2904 , w_2905 , 
		w_2906 , w_2907 , w_2908 , w_2909 , w_2910 , w_2911 , w_2912 , w_2913 , w_2914 , w_2915 , 
		w_2916 , w_2917 , w_2918 , w_2919 , w_2920 , w_2921 , w_2922 , w_2923 , w_2924 , w_2925 , 
		w_2926 , w_2927 , w_2928 , w_2929 , w_2930 , w_2931 , w_2932 , w_2933 , w_2934 , w_2935 , 
		w_2936 , w_2937 , w_2938 , w_2939 , w_2940 , w_2941 , w_2942 , w_2943 , w_2944 , w_2945 , 
		w_2946 , w_2947 , w_2948 , w_2949 , w_2950 , w_2951 , w_2952 , w_2953 , w_2954 , w_2955 , 
		w_2956 , w_2957 , w_2958 , w_2959 , w_2960 , w_2961 , w_2962 , w_2963 , w_2964 , w_2965 , 
		w_2966 , w_2967 , w_2968 , w_2969 , w_2970 , w_2971 , w_2972 , w_2973 , w_2974 , w_2975 , 
		w_2976 , w_2977 , w_2978 , w_2979 , w_2980 , w_2981 , w_2982 , w_2983 , w_2984 , w_2985 , 
		w_2986 , w_2987 , w_2988 , w_2989 , w_2990 , w_2991 , w_2992 , w_2993 , w_2994 , w_2995 , 
		w_2996 , w_2997 , w_2998 , w_2999 , w_3000 , w_3001 , w_3002 , w_3003 , w_3004 , w_3005 , 
		w_3006 , w_3007 , w_3008 , w_3009 , w_3010 , w_3011 , w_3012 , w_3013 , w_3014 , w_3015 , 
		w_3016 , w_3017 , w_3018 , w_3019 , w_3020 , w_3021 , w_3022 , w_3023 , w_3024 , w_3025 , 
		w_3026 , w_3027 , w_3028 , w_3029 , w_3030 , w_3031 , w_3032 , w_3033 , w_3034 , w_3035 , 
		w_3036 , w_3037 , w_3038 , w_3039 , w_3040 , w_3041 , w_3042 , w_3043 , w_3044 , w_3045 , 
		w_3046 , w_3047 , w_3048 , w_3049 , w_3050 , w_3051 , w_3052 , w_3053 , w_3054 , w_3055 , 
		w_3056 , w_3057 , w_3058 , w_3059 , w_3060 , w_3061 , w_3062 , w_3063 , w_3064 , w_3065 , 
		w_3066 , w_3067 , w_3068 , w_3069 , w_3070 , w_3071 , w_3072 , w_3073 , w_3074 , w_3075 , 
		w_3076 , w_3077 , w_3078 , w_3079 , w_3080 , w_3081 , w_3082 , w_3083 , w_3084 , w_3085 , 
		w_3086 , w_3087 , w_3088 , w_3089 , w_3090 , w_3091 , w_3092 , w_3093 , w_3094 , w_3095 , 
		w_3096 , w_3097 , w_3098 , w_3099 , w_3100 , w_3101 , w_3102 , w_3103 , w_3104 , w_3105 , 
		w_3106 , w_3107 , w_3108 , w_3109 , w_3110 , w_3111 , w_3112 , w_3113 , w_3114 , w_3115 , 
		w_3116 , w_3117 , w_3118 , w_3119 , w_3120 , w_3121 , w_3122 , w_3123 , w_3124 , w_3125 , 
		w_3126 , w_3127 , w_3128 , w_3129 , w_3130 , w_3131 , w_3132 , w_3133 , w_3134 , w_3135 , 
		w_3136 , w_3137 , w_3138 , w_3139 , w_3140 , w_3141 , w_3142 , w_3143 , w_3144 , w_3145 , 
		w_3146 , w_3147 , w_3148 , w_3149 , w_3150 , w_3151 , w_3152 , w_3153 , w_3154 , w_3155 , 
		w_3156 , w_3157 , w_3158 , w_3159 , w_3160 , w_3161 , w_3162 , w_3163 , w_3164 , w_3165 , 
		w_3166 , w_3167 , w_3168 , w_3169 , w_3170 , w_3171 , w_3172 , w_3173 , w_3174 , w_3175 , 
		w_3176 , w_3177 , w_3178 , w_3179 , w_3180 , w_3181 , w_3182 , w_3183 , w_3184 , w_3185 , 
		w_3186 , w_3187 , w_3188 , w_3189 , w_3190 , w_3191 , w_3192 , w_3193 , w_3194 , w_3195 , 
		w_3196 , w_3197 , w_3198 , w_3199 , w_3200 , w_3201 , w_3202 , w_3203 , w_3204 , w_3205 , 
		w_3206 , w_3207 , w_3208 , w_3209 , w_3210 , w_3211 , w_3212 , w_3213 , w_3214 , w_3215 , 
		w_3216 , w_3217 , w_3218 , w_3219 , w_3220 , w_3221 , w_3222 , w_3223 , w_3224 , w_3225 , 
		w_3226 , w_3227 , w_3228 , w_3229 , w_3230 , w_3231 , w_3232 , w_3233 , w_3234 , w_3235 , 
		w_3236 , w_3237 , w_3238 , w_3239 , w_3240 , w_3241 , w_3242 , w_3243 , w_3244 , w_3245 , 
		w_3246 , w_3247 , w_3248 , w_3249 , w_3250 , w_3251 , w_3252 , w_3253 , w_3254 , w_3255 , 
		w_3256 , w_3257 , w_3258 , w_3259 , w_3260 , w_3261 , w_3262 , w_3263 , w_3264 , w_3265 , 
		w_3266 , w_3267 , w_3268 , w_3269 , w_3270 , w_3271 , w_3272 , w_3273 , w_3274 , w_3275 , 
		w_3276 , w_3277 , w_3278 , w_3279 , w_3280 , w_3281 , w_3282 , w_3283 , w_3284 , w_3285 , 
		w_3286 , w_3287 , w_3288 , w_3289 , w_3290 , w_3291 , w_3292 , w_3293 , w_3294 , w_3295 , 
		w_3296 , w_3297 , w_3298 , w_3299 , w_3300 , w_3301 , w_3302 , w_3303 , w_3304 , w_3305 , 
		w_3306 , w_3307 , w_3308 , w_3309 , w_3310 , w_3311 , w_3312 , w_3313 , w_3314 , w_3315 , 
		w_3316 , w_3317 , w_3318 , w_3319 , w_3320 , w_3321 , w_3322 , w_3323 , w_3324 , w_3325 , 
		w_3326 , w_3327 , w_3328 , w_3329 , w_3330 , w_3331 , w_3332 , w_3333 , w_3334 , w_3335 , 
		w_3336 , w_3337 , w_3338 , w_3339 , w_3340 , w_3341 , w_3342 , w_3343 , w_3344 , w_3345 , 
		w_3346 , w_3347 , w_3348 , w_3349 , w_3350 , w_3351 , w_3352 , w_3353 , w_3354 , w_3355 , 
		w_3356 , w_3357 , w_3358 , w_3359 , w_3360 , w_3361 , w_3362 , w_3363 , w_3364 , w_3365 , 
		w_3366 , w_3367 , w_3368 , w_3369 , w_3370 , w_3371 , w_3372 , w_3373 , w_3374 , w_3375 , 
		w_3376 , w_3377 , w_3378 , w_3379 , w_3380 , w_3381 , w_3382 , w_3383 , w_3384 , w_3385 , 
		w_3386 , w_3387 , w_3388 , w_3389 , w_3390 , w_3391 , w_3392 , w_3393 , w_3394 , w_3395 , 
		w_3396 , w_3397 , w_3398 , w_3399 , w_3400 , w_3401 , w_3402 , w_3403 , w_3404 , w_3405 , 
		w_3406 , w_3407 , w_3408 , w_3409 , w_3410 , w_3411 , w_3412 , w_3413 , w_3414 , w_3415 , 
		w_3416 , w_3417 , w_3418 , w_3419 , w_3420 , w_3421 , w_3422 , w_3423 , w_3424 , w_3425 , 
		w_3426 , w_3427 , w_3428 , w_3429 , w_3430 , w_3431 , w_3432 , w_3433 , w_3434 , w_3435 , 
		w_3436 , w_3437 , w_3438 , w_3439 , w_3440 , w_3441 , w_3442 , w_3443 , w_3444 , w_3445 , 
		w_3446 , w_3447 , w_3448 , w_3449 , w_3450 , w_3451 , w_3452 , w_3453 , w_3454 , w_3455 , 
		w_3456 , w_3457 , w_3458 , w_3459 , w_3460 , w_3461 , w_3462 , w_3463 , w_3464 , w_3465 , 
		w_3466 , w_3467 , w_3468 , w_3469 , w_3470 , w_3471 , w_3472 , w_3473 , w_3474 , w_3475 , 
		w_3476 , w_3477 , w_3478 , w_3479 , w_3480 , w_3481 , w_3482 , w_3483 , w_3484 , w_3485 , 
		w_3486 , w_3487 , w_3488 , w_3489 , w_3490 , w_3491 , w_3492 , w_3493 , w_3494 , w_3495 , 
		w_3496 , w_3497 , w_3498 , w_3499 , w_3500 , w_3501 , w_3502 , w_3503 , w_3504 , w_3505 , 
		w_3506 , w_3507 , w_3508 , w_3509 , w_3510 , w_3511 , w_3512 , w_3513 , w_3514 , w_3515 , 
		w_3516 , w_3517 , w_3518 , w_3519 , w_3520 , w_3521 , w_3522 , w_3523 , w_3524 , w_3525 , 
		w_3526 , w_3527 , w_3528 , w_3529 , w_3530 , w_3531 , w_3532 , w_3533 , w_3534 , w_3535 , 
		w_3536 , w_3537 , w_3538 , w_3539 , w_3540 , w_3541 , w_3542 , w_3543 , w_3544 , w_3545 , 
		w_3546 , w_3547 , w_3548 , w_3549 , w_3550 , w_3551 , w_3552 , w_3553 , w_3554 , w_3555 , 
		w_3556 , w_3557 , w_3558 , w_3559 , w_3560 , w_3561 , w_3562 , w_3563 , w_3564 , w_3565 , 
		w_3566 , w_3567 , w_3568 , w_3569 , w_3570 , w_3571 , w_3572 , w_3573 , w_3574 , w_3575 , 
		w_3576 , w_3577 , w_3578 , w_3579 , w_3580 , w_3581 , w_3582 , w_3583 , w_3584 , w_3585 , 
		w_3586 , w_3587 , w_3588 , w_3589 , w_3590 , w_3591 , w_3592 , w_3593 , w_3594 , w_3595 , 
		w_3596 , w_3597 , w_3598 , w_3599 , w_3600 , w_3601 , w_3602 , w_3603 , w_3604 , w_3605 , 
		w_3606 , w_3607 , w_3608 , w_3609 , w_3610 , w_3611 , w_3612 , w_3613 , w_3614 , w_3615 , 
		w_3616 , w_3617 , w_3618 , w_3619 , w_3620 , w_3621 , w_3622 , w_3623 , w_3624 , w_3625 , 
		w_3626 , w_3627 , w_3628 , w_3629 , w_3630 , w_3631 , w_3632 , w_3633 , w_3634 , w_3635 , 
		w_3636 , w_3637 , w_3638 , w_3639 , w_3640 , w_3641 , w_3642 , w_3643 , w_3644 , w_3645 , 
		w_3646 , w_3647 , w_3648 , w_3649 , w_3650 , w_3651 , w_3652 , w_3653 , w_3654 , w_3655 , 
		w_3656 , w_3657 , w_3658 , w_3659 , w_3660 , w_3661 , w_3662 , w_3663 , w_3664 , w_3665 , 
		w_3666 , w_3667 , w_3668 , w_3669 , w_3670 , w_3671 , w_3672 , w_3673 , w_3674 , w_3675 , 
		w_3676 , w_3677 , w_3678 , w_3679 , w_3680 , w_3681 , w_3682 , w_3683 , w_3684 , w_3685 , 
		w_3686 , w_3687 , w_3688 , w_3689 , w_3690 , w_3691 , w_3692 , w_3693 , w_3694 , w_3695 , 
		w_3696 , w_3697 , w_3698 , w_3699 , w_3700 , w_3701 , w_3702 , w_3703 , w_3704 , w_3705 , 
		w_3706 , w_3707 , w_3708 , w_3709 , w_3710 , w_3711 , w_3712 , w_3713 , w_3714 , w_3715 , 
		w_3716 , w_3717 , w_3718 , w_3719 , w_3720 , w_3721 , w_3722 , w_3723 , w_3724 , w_3725 , 
		w_3726 , w_3727 , w_3728 , w_3729 , w_3730 , w_3731 , w_3732 , w_3733 , w_3734 , w_3735 , 
		w_3736 , w_3737 , w_3738 , w_3739 , w_3740 , w_3741 , w_3742 , w_3743 , w_3744 , w_3745 , 
		w_3746 , w_3747 , w_3748 , w_3749 , w_3750 , w_3751 , w_3752 , w_3753 , w_3754 , w_3755 , 
		w_3756 , w_3757 , w_3758 , w_3759 , w_3760 , w_3761 , w_3762 , w_3763 , w_3764 , w_3765 , 
		w_3766 , w_3767 , w_3768 , w_3769 , w_3770 , w_3771 , w_3772 , w_3773 , w_3774 , w_3775 , 
		w_3776 , w_3777 , w_3778 , w_3779 , w_3780 , w_3781 , w_3782 , w_3783 , w_3784 , w_3785 , 
		w_3786 , w_3787 , w_3788 , w_3789 , w_3790 , w_3791 , w_3792 , w_3793 , w_3794 , w_3795 , 
		w_3796 , w_3797 , w_3798 , w_3799 , w_3800 , w_3801 , w_3802 , w_3803 , w_3804 , w_3805 , 
		w_3806 , w_3807 , w_3808 , w_3809 , w_3810 , w_3811 , w_3812 , w_3813 , w_3814 , w_3815 , 
		w_3816 , w_3817 , w_3818 , w_3819 , w_3820 , w_3821 , w_3822 , w_3823 , w_3824 , w_3825 , 
		w_3826 , w_3827 , w_3828 , w_3829 , w_3830 , w_3831 , w_3832 , w_3833 , w_3834 , w_3835 , 
		w_3836 , w_3837 , w_3838 , w_3839 , w_3840 , w_3841 , w_3842 , w_3843 , w_3844 , w_3845 , 
		w_3846 , w_3847 , w_3848 , w_3849 , w_3850 , w_3851 , w_3852 , w_3853 , w_3854 , w_3855 , 
		w_3856 , w_3857 , w_3858 , w_3859 , w_3860 , w_3861 , w_3862 , w_3863 , w_3864 , w_3865 , 
		w_3866 , w_3867 , w_3868 , w_3869 , w_3870 , w_3871 , w_3872 , w_3873 , w_3874 , w_3875 , 
		w_3876 , w_3877 , w_3878 , w_3879 , w_3880 , w_3881 , w_3882 , w_3883 , w_3884 , w_3885 , 
		w_3886 , w_3887 , w_3888 , w_3889 , w_3890 , w_3891 , w_3892 , w_3893 , w_3894 , w_3895 , 
		w_3896 , w_3897 , w_3898 , w_3899 , w_3900 , w_3901 , w_3902 , w_3903 , w_3904 , w_3905 , 
		w_3906 , w_3907 , w_3908 , w_3909 , w_3910 , w_3911 , w_3912 , w_3913 , w_3914 , w_3915 , 
		w_3916 , w_3917 , w_3918 , w_3919 , w_3920 , w_3921 , w_3922 , w_3923 , w_3924 , w_3925 , 
		w_3926 , w_3927 , w_3928 , w_3929 , w_3930 , w_3931 , w_3932 , w_3933 , w_3934 , w_3935 , 
		w_3936 , w_3937 , w_3938 , w_3939 , w_3940 , w_3941 , w_3942 , w_3943 , w_3944 , w_3945 , 
		w_3946 , w_3947 , w_3948 , w_3949 , w_3950 , w_3951 , w_3952 , w_3953 , w_3954 , w_3955 , 
		w_3956 , w_3957 , w_3958 , w_3959 , w_3960 , w_3961 , w_3962 , w_3963 , w_3964 , w_3965 , 
		w_3966 , w_3967 , w_3968 , w_3969 , w_3970 , w_3971 , w_3972 , w_3973 , w_3974 , w_3975 , 
		w_3976 , w_3977 , w_3978 , w_3979 , w_3980 , w_3981 , w_3982 , w_3983 , w_3984 , w_3985 , 
		w_3986 , w_3987 , w_3988 , w_3989 , w_3990 , w_3991 , w_3992 , w_3993 , w_3994 , w_3995 , 
		w_3996 , w_3997 , w_3998 , w_3999 , w_4000 , w_4001 , w_4002 , w_4003 , w_4004 , w_4005 , 
		w_4006 , w_4007 , w_4008 , w_4009 , w_4010 , w_4011 , w_4012 , w_4013 , w_4014 , w_4015 , 
		w_4016 , w_4017 , w_4018 , w_4019 , w_4020 , w_4021 , w_4022 , w_4023 , w_4024 , w_4025 , 
		w_4026 , w_4027 , w_4028 , w_4029 , w_4030 , w_4031 , w_4032 , w_4033 , w_4034 , w_4035 , 
		w_4036 , w_4037 , w_4038 , w_4039 , w_4040 , w_4041 , w_4042 , w_4043 , w_4044 , w_4045 , 
		w_4046 , w_4047 , w_4048 , w_4049 , w_4050 , w_4051 , w_4052 , w_4053 , w_4054 , w_4055 , 
		w_4056 , w_4057 , w_4058 , w_4059 , w_4060 , w_4061 , w_4062 , w_4063 , w_4064 , w_4065 , 
		w_4066 , w_4067 , w_4068 , w_4069 , w_4070 , w_4071 , w_4072 , w_4073 , w_4074 , w_4075 , 
		w_4076 , w_4077 , w_4078 , w_4079 , w_4080 , w_4081 , w_4082 , w_4083 , w_4084 , w_4085 , 
		w_4086 , w_4087 , w_4088 , w_4089 , w_4090 , w_4091 , w_4092 , w_4093 , w_4094 , w_4095 , 
		w_4096 , w_4097 , w_4098 , w_4099 , w_4100 , w_4101 , w_4102 , w_4103 , w_4104 , w_4105 , 
		w_4106 , w_4107 , w_4108 , w_4109 , w_4110 , w_4111 , w_4112 , w_4113 , w_4114 , w_4115 , 
		w_4116 , w_4117 , w_4118 , w_4119 , w_4120 , w_4121 , w_4122 , w_4123 , w_4124 , w_4125 , 
		w_4126 , w_4127 , w_4128 , w_4129 , w_4130 , w_4131 , w_4132 , w_4133 , w_4134 , w_4135 , 
		w_4136 , w_4137 , w_4138 , w_4139 , w_4140 , w_4141 , w_4142 , w_4143 , w_4144 , w_4145 , 
		w_4146 , w_4147 , w_4148 , w_4149 , w_4150 , w_4151 , w_4152 , w_4153 , w_4154 , w_4155 , 
		w_4156 , w_4157 , w_4158 , w_4159 , w_4160 , w_4161 , w_4162 , w_4163 , w_4164 , w_4165 , 
		w_4166 , w_4167 , w_4168 , w_4169 , w_4170 , w_4171 , w_4172 , w_4173 , w_4174 , w_4175 , 
		w_4176 , w_4177 , w_4178 , w_4179 , w_4180 , w_4181 , w_4182 , w_4183 , w_4184 , w_4185 , 
		w_4186 , w_4187 , w_4188 , w_4189 , w_4190 , w_4191 , w_4192 , w_4193 , w_4194 , w_4195 , 
		w_4196 , w_4197 , w_4198 , w_4199 , w_4200 , w_4201 , w_4202 , w_4203 , w_4204 , w_4205 , 
		w_4206 , w_4207 , w_4208 , w_4209 , w_4210 , w_4211 , w_4212 , w_4213 , w_4214 , w_4215 , 
		w_4216 , w_4217 , w_4218 , w_4219 , w_4220 , w_4221 , w_4222 , w_4223 , w_4224 , w_4225 , 
		w_4226 , w_4227 , w_4228 , w_4229 , w_4230 , w_4231 , w_4232 , w_4233 , w_4234 , w_4235 , 
		w_4236 , w_4237 , w_4238 , w_4239 , w_4240 , w_4241 , w_4242 , w_4243 , w_4244 , w_4245 , 
		w_4246 , w_4247 , w_4248 , w_4249 , w_4250 , w_4251 , w_4252 , w_4253 , w_4254 , w_4255 , 
		w_4256 , w_4257 , w_4258 , w_4259 , w_4260 , w_4261 , w_4262 , w_4263 , w_4264 , w_4265 , 
		w_4266 , w_4267 , w_4268 , w_4269 , w_4270 , w_4271 , w_4272 , w_4273 , w_4274 , w_4275 , 
		w_4276 , w_4277 , w_4278 , w_4279 , w_4280 , w_4281 , w_4282 , w_4283 , w_4284 , w_4285 , 
		w_4286 , w_4287 , w_4288 , w_4289 , w_4290 , w_4291 , w_4292 , w_4293 , w_4294 , w_4295 , 
		w_4296 , w_4297 , w_4298 , w_4299 , w_4300 , w_4301 , w_4302 , w_4303 , w_4304 , w_4305 , 
		w_4306 , w_4307 , w_4308 , w_4309 , w_4310 , w_4311 , w_4312 , w_4313 , w_4314 , w_4315 , 
		w_4316 , w_4317 , w_4318 , w_4319 , w_4320 , w_4321 , w_4322 , w_4323 , w_4324 , w_4325 , 
		w_4326 , w_4327 , w_4328 , w_4329 , w_4330 , w_4331 , w_4332 , w_4333 , w_4334 , w_4335 , 
		w_4336 , w_4337 , w_4338 , w_4339 , w_4340 , w_4341 , w_4342 , w_4343 , w_4344 , w_4345 , 
		w_4346 , w_4347 , w_4348 , w_4349 , w_4350 , w_4351 , w_4352 , w_4353 , w_4354 , w_4355 , 
		w_4356 , w_4357 , w_4358 , w_4359 , w_4360 , w_4361 , w_4362 , w_4363 , w_4364 , w_4365 , 
		w_4366 , w_4367 , w_4368 , w_4369 , w_4370 , w_4371 , w_4372 , w_4373 , w_4374 , w_4375 , 
		w_4376 , w_4377 , w_4378 , w_4379 , w_4380 , w_4381 , w_4382 , w_4383 , w_4384 , w_4385 , 
		w_4386 , w_4387 , w_4388 , w_4389 , w_4390 , w_4391 , w_4392 , w_4393 , w_4394 , w_4395 , 
		w_4396 , w_4397 , w_4398 , w_4399 , w_4400 , w_4401 , w_4402 , w_4403 , w_4404 , w_4405 , 
		w_4406 , w_4407 , w_4408 , w_4409 , w_4410 , w_4411 , w_4412 , w_4413 , w_4414 , w_4415 , 
		w_4416 , w_4417 , w_4418 , w_4419 , w_4420 , w_4421 , w_4422 , w_4423 , w_4424 , w_4425 , 
		w_4426 , w_4427 , w_4428 , w_4429 , w_4430 , w_4431 , w_4432 , w_4433 , w_4434 , w_4435 , 
		w_4436 , w_4437 , w_4438 , w_4439 , w_4440 , w_4441 , w_4442 , w_4443 , w_4444 , w_4445 , 
		w_4446 , w_4447 , w_4448 , w_4449 , w_4450 , w_4451 , w_4452 , w_4453 , w_4454 , w_4455 , 
		w_4456 , w_4457 , w_4458 , w_4459 , w_4460 , w_4461 , w_4462 , w_4463 , w_4464 , w_4465 , 
		w_4466 , w_4467 , w_4468 , w_4469 , w_4470 , w_4471 , w_4472 , w_4473 , w_4474 , w_4475 , 
		w_4476 , w_4477 , w_4478 , w_4479 , w_4480 , w_4481 , w_4482 , w_4483 , w_4484 , w_4485 , 
		w_4486 , w_4487 , w_4488 , w_4489 , w_4490 , w_4491 , w_4492 , w_4493 , w_4494 , w_4495 , 
		w_4496 , w_4497 , w_4498 , w_4499 , w_4500 , w_4501 , w_4502 , w_4503 , w_4504 , w_4505 , 
		w_4506 , w_4507 , w_4508 , w_4509 , w_4510 , w_4511 , w_4512 , w_4513 , w_4514 , w_4515 , 
		w_4516 , w_4517 , w_4518 , w_4519 , w_4520 , w_4521 , w_4522 , w_4523 , w_4524 , w_4525 , 
		w_4526 , w_4527 , w_4528 , w_4529 , w_4530 , w_4531 , w_4532 , w_4533 , w_4534 , w_4535 , 
		w_4536 , w_4537 , w_4538 , w_4539 , w_4540 , w_4541 , w_4542 , w_4543 , w_4544 , w_4545 , 
		w_4546 , w_4547 , w_4548 , w_4549 , w_4550 , w_4551 , w_4552 , w_4553 , w_4554 , w_4555 , 
		w_4556 , w_4557 , w_4558 , w_4559 , w_4560 , w_4561 , w_4562 , w_4563 , w_4564 , w_4565 , 
		w_4566 , w_4567 , w_4568 , w_4569 , w_4570 , w_4571 , w_4572 , w_4573 , w_4574 , w_4575 , 
		w_4576 , w_4577 , w_4578 , w_4579 , w_4580 , w_4581 , w_4582 , w_4583 , w_4584 , w_4585 , 
		w_4586 , w_4587 , w_4588 , w_4589 , w_4590 , w_4591 , w_4592 , w_4593 , w_4594 , w_4595 , 
		w_4596 , w_4597 , w_4598 , w_4599 , w_4600 , w_4601 , w_4602 , w_4603 , w_4604 , w_4605 , 
		w_4606 , w_4607 , w_4608 , w_4609 , w_4610 , w_4611 , w_4612 , w_4613 , w_4614 , w_4615 , 
		w_4616 , w_4617 , w_4618 , w_4619 , w_4620 , w_4621 , w_4622 , w_4623 , w_4624 , w_4625 , 
		w_4626 , w_4627 , w_4628 , w_4629 , w_4630 , w_4631 , w_4632 , w_4633 , w_4634 , w_4635 , 
		w_4636 , w_4637 , w_4638 , w_4639 , w_4640 , w_4641 , w_4642 , w_4643 , w_4644 , w_4645 , 
		w_4646 , w_4647 , w_4648 , w_4649 , w_4650 , w_4651 , w_4652 , w_4653 , w_4654 , w_4655 , 
		w_4656 , w_4657 , w_4658 , w_4659 , w_4660 , w_4661 , w_4662 , w_4663 , w_4664 , w_4665 , 
		w_4666 , w_4667 , w_4668 , w_4669 , w_4670 , w_4671 , w_4672 , w_4673 , w_4674 , w_4675 , 
		w_4676 , w_4677 , w_4678 , w_4679 , w_4680 , w_4681 , w_4682 , w_4683 , w_4684 , w_4685 , 
		w_4686 , w_4687 , w_4688 , w_4689 , w_4690 , w_4691 , w_4692 , w_4693 , w_4694 , w_4695 , 
		w_4696 , w_4697 , w_4698 , w_4699 , w_4700 , w_4701 , w_4702 , w_4703 , w_4704 , w_4705 , 
		w_4706 , w_4707 , w_4708 , w_4709 , w_4710 , w_4711 , w_4712 , w_4713 , w_4714 , w_4715 , 
		w_4716 , w_4717 , w_4718 , w_4719 , w_4720 , w_4721 , w_4722 , w_4723 , w_4724 , w_4725 , 
		w_4726 , w_4727 , w_4728 , w_4729 , w_4730 , w_4731 , w_4732 , w_4733 , w_4734 , w_4735 , 
		w_4736 , w_4737 , w_4738 , w_4739 , w_4740 , w_4741 , w_4742 , w_4743 , w_4744 , w_4745 , 
		w_4746 , w_4747 , w_4748 , w_4749 , w_4750 , w_4751 , w_4752 , w_4753 , w_4754 , w_4755 , 
		w_4756 , w_4757 , w_4758 , w_4759 , w_4760 , w_4761 , w_4762 , w_4763 , w_4764 , w_4765 , 
		w_4766 , w_4767 , w_4768 , w_4769 , w_4770 , w_4771 , w_4772 , w_4773 , w_4774 , w_4775 , 
		w_4776 , w_4777 , w_4778 , w_4779 , w_4780 , w_4781 , w_4782 , w_4783 , w_4784 , w_4785 , 
		w_4786 , w_4787 , w_4788 , w_4789 , w_4790 , w_4791 , w_4792 , w_4793 , w_4794 , w_4795 , 
		w_4796 , w_4797 , w_4798 , w_4799 , w_4800 , w_4801 , w_4802 , w_4803 , w_4804 , w_4805 , 
		w_4806 , w_4807 , w_4808 , w_4809 , w_4810 , w_4811 , w_4812 , w_4813 , w_4814 , w_4815 , 
		w_4816 , w_4817 , w_4818 , w_4819 , w_4820 , w_4821 , w_4822 , w_4823 , w_4824 , w_4825 , 
		w_4826 , w_4827 , w_4828 , w_4829 , w_4830 , w_4831 , w_4832 , w_4833 , w_4834 , w_4835 , 
		w_4836 , w_4837 , w_4838 , w_4839 , w_4840 , w_4841 , w_4842 , w_4843 , w_4844 , w_4845 , 
		w_4846 , w_4847 , w_4848 , w_4849 , w_4850 , w_4851 , w_4852 , w_4853 , w_4854 , w_4855 , 
		w_4856 , w_4857 , w_4858 , w_4859 , w_4860 , w_4861 , w_4862 , w_4863 , w_4864 , w_4865 , 
		w_4866 , w_4867 , w_4868 , w_4869 , w_4870 , w_4871 , w_4872 , w_4873 , w_4874 , w_4875 , 
		w_4876 , w_4877 , w_4878 , w_4879 , w_4880 , w_4881 , w_4882 , w_4883 , w_4884 , w_4885 , 
		w_4886 , w_4887 , w_4888 , w_4889 , w_4890 , w_4891 , w_4892 , w_4893 , w_4894 , w_4895 , 
		w_4896 , w_4897 , w_4898 , w_4899 , w_4900 , w_4901 , w_4902 , w_4903 , w_4904 , w_4905 , 
		w_4906 , w_4907 , w_4908 , w_4909 , w_4910 , w_4911 , w_4912 , w_4913 , w_4914 , w_4915 , 
		w_4916 , w_4917 , w_4918 , w_4919 , w_4920 , w_4921 , w_4922 , w_4923 , w_4924 , w_4925 , 
		w_4926 , w_4927 , w_4928 , w_4929 , w_4930 , w_4931 , w_4932 , w_4933 , w_4934 , w_4935 , 
		w_4936 , w_4937 , w_4938 , w_4939 , w_4940 , w_4941 , w_4942 , w_4943 , w_4944 , w_4945 , 
		w_4946 , w_4947 , w_4948 , w_4949 , w_4950 , w_4951 , w_4952 , w_4953 , w_4954 , w_4955 , 
		w_4956 , w_4957 , w_4958 , w_4959 , w_4960 , w_4961 , w_4962 , w_4963 , w_4964 , w_4965 , 
		w_4966 , w_4967 , w_4968 , w_4969 , w_4970 , w_4971 , w_4972 , w_4973 , w_4974 , w_4975 , 
		w_4976 , w_4977 , w_4978 , w_4979 , w_4980 , w_4981 , w_4982 , w_4983 , w_4984 , w_4985 , 
		w_4986 , w_4987 , w_4988 , w_4989 , w_4990 , w_4991 , w_4992 , w_4993 , w_4994 , w_4995 , 
		w_4996 , w_4997 , w_4998 , w_4999 , w_5000 , w_5001 , w_5002 , w_5003 , w_5004 , w_5005 , 
		w_5006 , w_5007 , w_5008 , w_5009 , w_5010 , w_5011 , w_5012 , w_5013 , w_5014 , w_5015 , 
		w_5016 , w_5017 , w_5018 , w_5019 , w_5020 , w_5021 , w_5022 , w_5023 , w_5024 , w_5025 , 
		w_5026 , w_5027 , w_5028 , w_5029 , w_5030 , w_5031 , w_5032 , w_5033 , w_5034 , w_5035 , 
		w_5036 , w_5037 , w_5038 , w_5039 , w_5040 , w_5041 , w_5042 , w_5043 , w_5044 , w_5045 , 
		w_5046 , w_5047 , w_5048 , w_5049 , w_5050 , w_5051 , w_5052 , w_5053 , w_5054 , w_5055 , 
		w_5056 , w_5057 , w_5058 , w_5059 , w_5060 , w_5061 , w_5062 , w_5063 , w_5064 , w_5065 , 
		w_5066 , w_5067 , w_5068 , w_5069 , w_5070 , w_5071 , w_5072 , w_5073 , w_5074 , w_5075 , 
		w_5076 , w_5077 , w_5078 , w_5079 , w_5080 , w_5081 , w_5082 , w_5083 , w_5084 , w_5085 , 
		w_5086 , w_5087 , w_5088 , w_5089 , w_5090 , w_5091 , w_5092 , w_5093 , w_5094 , w_5095 , 
		w_5096 , w_5097 , w_5098 , w_5099 , w_5100 , w_5101 , w_5102 , w_5103 , w_5104 , w_5105 , 
		w_5106 , w_5107 , w_5108 , w_5109 , w_5110 , w_5111 , w_5112 , w_5113 , w_5114 , w_5115 , 
		w_5116 , w_5117 , w_5118 , w_5119 , w_5120 , w_5121 , w_5122 , w_5123 , w_5124 , w_5125 , 
		w_5126 , w_5127 , w_5128 , w_5129 , w_5130 , w_5131 , w_5132 , w_5133 , w_5134 , w_5135 , 
		w_5136 , w_5137 , w_5138 , w_5139 , w_5140 , w_5141 , w_5142 , w_5143 , w_5144 , w_5145 , 
		w_5146 , w_5147 , w_5148 , w_5149 , w_5150 , w_5151 , w_5152 , w_5153 , w_5154 , w_5155 , 
		w_5156 , w_5157 , w_5158 , w_5159 , w_5160 , w_5161 , w_5162 , w_5163 , w_5164 , w_5165 , 
		w_5166 , w_5167 , w_5168 , w_5169 , w_5170 , w_5171 , w_5172 , w_5173 , w_5174 , w_5175 , 
		w_5176 , w_5177 , w_5178 , w_5179 , w_5180 , w_5181 , w_5182 , w_5183 , w_5184 , w_5185 , 
		w_5186 , w_5187 , w_5188 , w_5189 , w_5190 , w_5191 , w_5192 , w_5193 , w_5194 , w_5195 , 
		w_5196 , w_5197 , w_5198 , w_5199 , w_5200 , w_5201 , w_5202 , w_5203 , w_5204 , w_5205 , 
		w_5206 , w_5207 , w_5208 , w_5209 , w_5210 , w_5211 , w_5212 , w_5213 , w_5214 , w_5215 , 
		w_5216 , w_5217 , w_5218 , w_5219 , w_5220 , w_5221 , w_5222 , w_5223 , w_5224 , w_5225 , 
		w_5226 , w_5227 , w_5228 , w_5229 , w_5230 , w_5231 , w_5232 , w_5233 , w_5234 , w_5235 , 
		w_5236 , w_5237 , w_5238 , w_5239 , w_5240 , w_5241 , w_5242 , w_5243 , w_5244 , w_5245 , 
		w_5246 , w_5247 , w_5248 , w_5249 , w_5250 , w_5251 , w_5252 , w_5253 , w_5254 , w_5255 , 
		w_5256 , w_5257 , w_5258 , w_5259 , w_5260 , w_5261 , w_5262 , w_5263 , w_5264 , w_5265 , 
		w_5266 , w_5267 , w_5268 , w_5269 , w_5270 , w_5271 , w_5272 , w_5273 , w_5274 , w_5275 , 
		w_5276 , w_5277 , w_5278 , w_5279 , w_5280 , w_5281 , w_5282 , w_5283 , w_5284 , w_5285 , 
		w_5286 , w_5287 , w_5288 , w_5289 , w_5290 , w_5291 , w_5292 , w_5293 , w_5294 , w_5295 , 
		w_5296 , w_5297 , w_5298 , w_5299 , w_5300 , w_5301 , w_5302 , w_5303 , w_5304 , w_5305 , 
		w_5306 , w_5307 , w_5308 , w_5309 , w_5310 , w_5311 , w_5312 , w_5313 , w_5314 , w_5315 , 
		w_5316 , w_5317 , w_5318 , w_5319 , w_5320 , w_5321 , w_5322 , w_5323 , w_5324 , w_5325 , 
		w_5326 , w_5327 , w_5328 , w_5329 , w_5330 , w_5331 , w_5332 , w_5333 , w_5334 , w_5335 , 
		w_5336 , w_5337 , w_5338 , w_5339 , w_5340 , w_5341 , w_5342 , w_5343 , w_5344 , w_5345 , 
		w_5346 , w_5347 , w_5348 , w_5349 , w_5350 , w_5351 , w_5352 , w_5353 , w_5354 , w_5355 , 
		w_5356 , w_5357 , w_5358 , w_5359 , w_5360 , w_5361 , w_5362 , w_5363 , w_5364 , w_5365 , 
		w_5366 , w_5367 , w_5368 , w_5369 , w_5370 , w_5371 , w_5372 , w_5373 , w_5374 , w_5375 , 
		w_5376 , w_5377 , w_5378 , w_5379 , w_5380 , w_5381 , w_5382 , w_5383 , w_5384 , w_5385 , 
		w_5386 , w_5387 , w_5388 , w_5389 , w_5390 , w_5391 , w_5392 , w_5393 , w_5394 , w_5395 , 
		w_5396 , w_5397 , w_5398 , w_5399 , w_5400 , w_5401 , w_5402 , w_5403 , w_5404 , w_5405 , 
		w_5406 , w_5407 , w_5408 , w_5409 , w_5410 , w_5411 , w_5412 , w_5413 , w_5414 , w_5415 , 
		w_5416 , w_5417 , w_5418 , w_5419 , w_5420 , w_5421 , w_5422 , w_5423 , w_5424 , w_5425 , 
		w_5426 , w_5427 , w_5428 , w_5429 , w_5430 , w_5431 , w_5432 , w_5433 , w_5434 , w_5435 , 
		w_5436 , w_5437 , w_5438 , w_5439 , w_5440 , w_5441 , w_5442 , w_5443 , w_5444 , w_5445 , 
		w_5446 , w_5447 , w_5448 , w_5449 , w_5450 , w_5451 , w_5452 , w_5453 , w_5454 , w_5455 , 
		w_5456 , w_5457 , w_5458 , w_5459 , w_5460 , w_5461 , w_5462 , w_5463 , w_5464 , w_5465 , 
		w_5466 , w_5467 , w_5468 , w_5469 , w_5470 , w_5471 , w_5472 , w_5473 , w_5474 , w_5475 , 
		w_5476 , w_5477 , w_5478 , w_5479 , w_5480 , w_5481 , w_5482 , w_5483 , w_5484 , w_5485 , 
		w_5486 , w_5487 , w_5488 , w_5489 , w_5490 , w_5491 , w_5492 , w_5493 , w_5494 , w_5495 , 
		w_5496 , w_5497 , w_5498 , w_5499 , w_5500 , w_5501 , w_5502 , w_5503 , w_5504 , w_5505 , 
		w_5506 , w_5507 , w_5508 , w_5509 , w_5510 , w_5511 , w_5512 , w_5513 , w_5514 , w_5515 , 
		w_5516 , w_5517 , w_5518 , w_5519 , w_5520 , w_5521 , w_5522 , w_5523 , w_5524 , w_5525 , 
		w_5526 , w_5527 , w_5528 , w_5529 , w_5530 , w_5531 , w_5532 , w_5533 , w_5534 , w_5535 , 
		w_5536 , w_5537 , w_5538 , w_5539 , w_5540 , w_5541 , w_5542 , w_5543 , w_5544 , w_5545 , 
		w_5546 , w_5547 , w_5548 , w_5549 , w_5550 , w_5551 , w_5552 , w_5553 , w_5554 , w_5555 , 
		w_5556 , w_5557 , w_5558 , w_5559 , w_5560 , w_5561 , w_5562 , w_5563 , w_5564 , w_5565 , 
		w_5566 , w_5567 , w_5568 , w_5569 , w_5570 , w_5571 , w_5572 , w_5573 , w_5574 , w_5575 , 
		w_5576 , w_5577 , w_5578 , w_5579 , w_5580 , w_5581 , w_5582 , w_5583 , w_5584 , w_5585 , 
		w_5586 , w_5587 , w_5588 , w_5589 , w_5590 , w_5591 , w_5592 , w_5593 , w_5594 , w_5595 , 
		w_5596 , w_5597 , w_5598 , w_5599 , w_5600 , w_5601 , w_5602 , w_5603 , w_5604 , w_5605 , 
		w_5606 , w_5607 , w_5608 , w_5609 , w_5610 , w_5611 , w_5612 , w_5613 , w_5614 , w_5615 , 
		w_5616 , w_5617 , w_5618 , w_5619 , w_5620 , w_5621 , w_5622 , w_5623 , w_5624 , w_5625 , 
		w_5626 , w_5627 , w_5628 , w_5629 , w_5630 , w_5631 , w_5632 , w_5633 , w_5634 , w_5635 , 
		w_5636 , w_5637 , w_5638 , w_5639 , w_5640 , w_5641 , w_5642 , w_5643 , w_5644 , w_5645 , 
		w_5646 , w_5647 , w_5648 , w_5649 , w_5650 , w_5651 , w_5652 , w_5653 , w_5654 , w_5655 , 
		w_5656 , w_5657 , w_5658 , w_5659 , w_5660 , w_5661 , w_5662 , w_5663 , w_5664 , w_5665 , 
		w_5666 , w_5667 , w_5668 , w_5669 , w_5670 , w_5671 , w_5672 , w_5673 , w_5674 , w_5675 , 
		w_5676 , w_5677 , w_5678 , w_5679 , w_5680 , w_5681 , w_5682 , w_5683 , w_5684 , w_5685 , 
		w_5686 , w_5687 , w_5688 , w_5689 , w_5690 , w_5691 , w_5692 , w_5693 , w_5694 , w_5695 , 
		w_5696 , w_5697 , w_5698 , w_5699 , w_5700 , w_5701 , w_5702 , w_5703 , w_5704 , w_5705 , 
		w_5706 , w_5707 , w_5708 , w_5709 , w_5710 , w_5711 , w_5712 , w_5713 , w_5714 , w_5715 , 
		w_5716 , w_5717 , w_5718 , w_5719 , w_5720 , w_5721 , w_5722 , w_5723 , w_5724 , w_5725 , 
		w_5726 , w_5727 , w_5728 , w_5729 , w_5730 , w_5731 , w_5732 , w_5733 , w_5734 , w_5735 , 
		w_5736 , w_5737 , w_5738 , w_5739 , w_5740 , w_5741 , w_5742 , w_5743 , w_5744 , w_5745 , 
		w_5746 , w_5747 , w_5748 , w_5749 , w_5750 , w_5751 , w_5752 , w_5753 , w_5754 , w_5755 , 
		w_5756 , w_5757 , w_5758 , w_5759 , w_5760 , w_5761 , w_5762 , w_5763 , w_5764 , w_5765 , 
		w_5766 , w_5767 , w_5768 , w_5769 , w_5770 , w_5771 , w_5772 , w_5773 , w_5774 , w_5775 , 
		w_5776 , w_5777 , w_5778 , w_5779 , w_5780 , w_5781 , w_5782 , w_5783 , w_5784 , w_5785 , 
		w_5786 , w_5787 , w_5788 , w_5789 , w_5790 , w_5791 , w_5792 , w_5793 , w_5794 , w_5795 , 
		w_5796 , w_5797 , w_5798 , w_5799 , w_5800 , w_5801 , w_5802 , w_5803 , w_5804 , w_5805 , 
		w_5806 , w_5807 , w_5808 , w_5809 , w_5810 , w_5811 , w_5812 , w_5813 , w_5814 , w_5815 , 
		w_5816 , w_5817 , w_5818 , w_5819 , w_5820 , w_5821 , w_5822 , w_5823 , w_5824 , w_5825 , 
		w_5826 , w_5827 , w_5828 , w_5829 , w_5830 , w_5831 , w_5832 , w_5833 , w_5834 , w_5835 , 
		w_5836 , w_5837 , w_5838 , w_5839 , w_5840 , w_5841 , w_5842 , w_5843 , w_5844 , w_5845 , 
		w_5846 , w_5847 , w_5848 , w_5849 , w_5850 , w_5851 , w_5852 , w_5853 , w_5854 , w_5855 , 
		w_5856 , w_5857 , w_5858 , w_5859 , w_5860 , w_5861 , w_5862 , w_5863 , w_5864 , w_5865 , 
		w_5866 , w_5867 , w_5868 , w_5869 , w_5870 , w_5871 , w_5872 , w_5873 , w_5874 , w_5875 , 
		w_5876 , w_5877 , w_5878 , w_5879 , w_5880 , w_5881 , w_5882 , w_5883 , w_5884 , w_5885 , 
		w_5886 , w_5887 , w_5888 , w_5889 , w_5890 , w_5891 , w_5892 , w_5893 , w_5894 , w_5895 , 
		w_5896 , w_5897 , w_5898 , w_5899 , w_5900 , w_5901 , w_5902 , w_5903 , w_5904 , w_5905 , 
		w_5906 , w_5907 , w_5908 , w_5909 , w_5910 , w_5911 , w_5912 , w_5913 , w_5914 , w_5915 , 
		w_5916 , w_5917 , w_5918 , w_5919 , w_5920 , w_5921 , w_5922 , w_5923 , w_5924 , w_5925 , 
		w_5926 , w_5927 , w_5928 , w_5929 , w_5930 , w_5931 , w_5932 , w_5933 , w_5934 , w_5935 , 
		w_5936 , w_5937 , w_5938 , w_5939 , w_5940 , w_5941 , w_5942 , w_5943 , w_5944 , w_5945 , 
		w_5946 , w_5947 , w_5948 , w_5949 , w_5950 , w_5951 , w_5952 , w_5953 , w_5954 , w_5955 , 
		w_5956 , w_5957 , w_5958 , w_5959 , w_5960 , w_5961 , w_5962 , w_5963 , w_5964 , w_5965 , 
		w_5966 , w_5967 , w_5968 , w_5969 , w_5970 , w_5971 , w_5972 , w_5973 , w_5974 , w_5975 , 
		w_5976 , w_5977 , w_5978 , w_5979 , w_5980 , w_5981 , w_5982 , w_5983 , w_5984 , w_5985 , 
		w_5986 , w_5987 , w_5988 , w_5989 , w_5990 , w_5991 , w_5992 , w_5993 , w_5994 , w_5995 , 
		w_5996 , w_5997 , w_5998 , w_5999 , w_6000 , w_6001 , w_6002 , w_6003 , w_6004 , w_6005 , 
		w_6006 , w_6007 , w_6008 , w_6009 , w_6010 , w_6011 , w_6012 , w_6013 , w_6014 , w_6015 , 
		w_6016 , w_6017 , w_6018 , w_6019 , w_6020 , w_6021 , w_6022 , w_6023 , w_6024 , w_6025 , 
		w_6026 , w_6027 , w_6028 , w_6029 , w_6030 , w_6031 , w_6032 , w_6033 , w_6034 , w_6035 , 
		w_6036 , w_6037 , w_6038 , w_6039 , w_6040 , w_6041 , w_6042 , w_6043 , w_6044 , w_6045 , 
		w_6046 , w_6047 , w_6048 , w_6049 , w_6050 , w_6051 , w_6052 , w_6053 , w_6054 , w_6055 , 
		w_6056 , w_6057 , w_6058 , w_6059 , w_6060 , w_6061 , w_6062 , w_6063 , w_6064 , w_6065 , 
		w_6066 , w_6067 , w_6068 , w_6069 , w_6070 , w_6071 , w_6072 , w_6073 , w_6074 , w_6075 , 
		w_6076 , w_6077 , w_6078 , w_6079 , w_6080 , w_6081 , w_6082 , w_6083 , w_6084 , w_6085 , 
		w_6086 , w_6087 , w_6088 , w_6089 , w_6090 , w_6091 , w_6092 , w_6093 , w_6094 , w_6095 , 
		w_6096 , w_6097 , w_6098 , w_6099 , w_6100 , w_6101 , w_6102 , w_6103 , w_6104 , w_6105 , 
		w_6106 , w_6107 , w_6108 , w_6109 , w_6110 , w_6111 , w_6112 , w_6113 , w_6114 , w_6115 , 
		w_6116 , w_6117 , w_6118 , w_6119 , w_6120 , w_6121 , w_6122 , w_6123 , w_6124 , w_6125 , 
		w_6126 , w_6127 , w_6128 , w_6129 , w_6130 , w_6131 , w_6132 , w_6133 , w_6134 , w_6135 , 
		w_6136 , w_6137 , w_6138 , w_6139 , w_6140 , w_6141 , w_6142 , w_6143 , w_6144 , w_6145 , 
		w_6146 , w_6147 , w_6148 , w_6149 , w_6150 , w_6151 , w_6152 , w_6153 , w_6154 , w_6155 , 
		w_6156 , w_6157 , w_6158 , w_6159 , w_6160 , w_6161 , w_6162 , w_6163 , w_6164 , w_6165 , 
		w_6166 , w_6167 , w_6168 , w_6169 , w_6170 , w_6171 , w_6172 , w_6173 , w_6174 , w_6175 , 
		w_6176 , w_6177 , w_6178 , w_6179 , w_6180 , w_6181 , w_6182 , w_6183 , w_6184 , w_6185 , 
		w_6186 , w_6187 , w_6188 , w_6189 , w_6190 , w_6191 , w_6192 , w_6193 , w_6194 , w_6195 , 
		w_6196 , w_6197 , w_6198 , w_6199 , w_6200 , w_6201 , w_6202 , w_6203 , w_6204 , w_6205 , 
		w_6206 , w_6207 , w_6208 , w_6209 , w_6210 , w_6211 , w_6212 , w_6213 , w_6214 , w_6215 , 
		w_6216 , w_6217 , w_6218 , w_6219 , w_6220 , w_6221 , w_6222 , w_6223 , w_6224 , w_6225 , 
		w_6226 , w_6227 , w_6228 , w_6229 , w_6230 , w_6231 , w_6232 , w_6233 , w_6234 , w_6235 , 
		w_6236 , w_6237 , w_6238 , w_6239 , w_6240 , w_6241 , w_6242 , w_6243 , w_6244 , w_6245 , 
		w_6246 , w_6247 , w_6248 , w_6249 , w_6250 , w_6251 , w_6252 , w_6253 , w_6254 , w_6255 , 
		w_6256 , w_6257 , w_6258 , w_6259 , w_6260 , w_6261 , w_6262 , w_6263 , w_6264 , w_6265 , 
		w_6266 , w_6267 , w_6268 , w_6269 , w_6270 , w_6271 , w_6272 , w_6273 , w_6274 , w_6275 , 
		w_6276 , w_6277 , w_6278 , w_6279 , w_6280 , w_6281 , w_6282 , w_6283 , w_6284 , w_6285 , 
		w_6286 , w_6287 , w_6288 , w_6289 , w_6290 , w_6291 , w_6292 , w_6293 , w_6294 , w_6295 , 
		w_6296 , w_6297 , w_6298 , w_6299 , w_6300 , w_6301 , w_6302 , w_6303 , w_6304 , w_6305 , 
		w_6306 , w_6307 , w_6308 , w_6309 , w_6310 , w_6311 , w_6312 , w_6313 , w_6314 , w_6315 , 
		w_6316 , w_6317 , w_6318 , w_6319 , w_6320 , w_6321 , w_6322 , w_6323 , w_6324 , w_6325 , 
		w_6326 , w_6327 , w_6328 , w_6329 , w_6330 , w_6331 , w_6332 , w_6333 , w_6334 , w_6335 , 
		w_6336 , w_6337 , w_6338 , w_6339 , w_6340 , w_6341 , w_6342 , w_6343 , w_6344 , w_6345 , 
		w_6346 , w_6347 , w_6348 , w_6349 , w_6350 , w_6351 , w_6352 , w_6353 , w_6354 , w_6355 , 
		w_6356 , w_6357 , w_6358 , w_6359 , w_6360 , w_6361 , w_6362 , w_6363 , w_6364 , w_6365 , 
		w_6366 , w_6367 , w_6368 , w_6369 , w_6370 , w_6371 , w_6372 , w_6373 , w_6374 , w_6375 , 
		w_6376 , w_6377 , w_6378 , w_6379 , w_6380 , w_6381 , w_6382 , w_6383 , w_6384 , w_6385 , 
		w_6386 , w_6387 , w_6388 , w_6389 , w_6390 , w_6391 , w_6392 , w_6393 , w_6394 , w_6395 , 
		w_6396 , w_6397 , w_6398 , w_6399 , w_6400 , w_6401 , w_6402 , w_6403 , w_6404 , w_6405 , 
		w_6406 , w_6407 , w_6408 , w_6409 , w_6410 , w_6411 , w_6412 , w_6413 , w_6414 , w_6415 , 
		w_6416 , w_6417 , w_6418 , w_6419 , w_6420 , w_6421 , w_6422 , w_6423 , w_6424 , w_6425 , 
		w_6426 , w_6427 , w_6428 , w_6429 , w_6430 , w_6431 , w_6432 , w_6433 , w_6434 , w_6435 , 
		w_6436 , w_6437 , w_6438 , w_6439 , w_6440 , w_6441 , w_6442 , w_6443 , w_6444 , w_6445 , 
		w_6446 , w_6447 , w_6448 , w_6449 , w_6450 , w_6451 , w_6452 , w_6453 , w_6454 , w_6455 , 
		w_6456 , w_6457 , w_6458 , w_6459 , w_6460 , w_6461 , w_6462 , w_6463 , w_6464 , w_6465 , 
		w_6466 , w_6467 , w_6468 , w_6469 , w_6470 , w_6471 , w_6472 , w_6473 , w_6474 , w_6475 , 
		w_6476 , w_6477 , w_6478 , w_6479 , w_6480 , w_6481 , w_6482 , w_6483 , w_6484 , w_6485 , 
		w_6486 , w_6487 , w_6488 , w_6489 , w_6490 , w_6491 , w_6492 , w_6493 , w_6494 , w_6495 , 
		w_6496 , w_6497 , w_6498 , w_6499 , w_6500 , w_6501 , w_6502 , w_6503 , w_6504 , w_6505 , 
		w_6506 , w_6507 , w_6508 , w_6509 , w_6510 , w_6511 , w_6512 , w_6513 , w_6514 , w_6515 , 
		w_6516 , w_6517 , w_6518 , w_6519 , w_6520 , w_6521 , w_6522 , w_6523 , w_6524 , w_6525 , 
		w_6526 , w_6527 , w_6528 , w_6529 , w_6530 , w_6531 , w_6532 , w_6533 , w_6534 , w_6535 , 
		w_6536 , w_6537 , w_6538 , w_6539 , w_6540 , w_6541 , w_6542 , w_6543 , w_6544 , w_6545 , 
		w_6546 , w_6547 , w_6548 , w_6549 , w_6550 , w_6551 , w_6552 , w_6553 , w_6554 , w_6555 , 
		w_6556 , w_6557 , w_6558 , w_6559 , w_6560 , w_6561 , w_6562 , w_6563 , w_6564 , w_6565 , 
		w_6566 , w_6567 , w_6568 , w_6569 , w_6570 , w_6571 , w_6572 , w_6573 , w_6574 , w_6575 , 
		w_6576 , w_6577 , w_6578 , w_6579 , w_6580 , w_6581 , w_6582 , w_6583 , w_6584 , w_6585 , 
		w_6586 , w_6587 , w_6588 , w_6589 , w_6590 , w_6591 , w_6592 , w_6593 , w_6594 , w_6595 , 
		w_6596 , w_6597 , w_6598 , w_6599 , w_6600 , w_6601 , w_6602 , w_6603 , w_6604 , w_6605 , 
		w_6606 , w_6607 , w_6608 , w_6609 , w_6610 , w_6611 , w_6612 , w_6613 , w_6614 , w_6615 , 
		w_6616 , w_6617 , w_6618 , w_6619 , w_6620 , w_6621 , w_6622 , w_6623 , w_6624 , w_6625 , 
		w_6626 , w_6627 , w_6628 , w_6629 , w_6630 , w_6631 , w_6632 , w_6633 , w_6634 , w_6635 , 
		w_6636 , w_6637 , w_6638 , w_6639 , w_6640 , w_6641 , w_6642 , w_6643 , w_6644 , w_6645 , 
		w_6646 , w_6647 , w_6648 , w_6649 , w_6650 , w_6651 , w_6652 , w_6653 , w_6654 , w_6655 , 
		w_6656 , w_6657 , w_6658 , w_6659 , w_6660 , w_6661 , w_6662 , w_6663 , w_6664 , w_6665 , 
		w_6666 , w_6667 , w_6668 , w_6669 , w_6670 , w_6671 , w_6672 , w_6673 , w_6674 , w_6675 , 
		w_6676 , w_6677 , w_6678 , w_6679 , w_6680 , w_6681 , w_6682 , w_6683 , w_6684 , w_6685 , 
		w_6686 , w_6687 , w_6688 , w_6689 , w_6690 , w_6691 , w_6692 , w_6693 , w_6694 , w_6695 , 
		w_6696 , w_6697 , w_6698 , w_6699 , w_6700 , w_6701 , w_6702 , w_6703 , w_6704 , w_6705 , 
		w_6706 , w_6707 , w_6708 , w_6709 , w_6710 , w_6711 , w_6712 , w_6713 , w_6714 , w_6715 , 
		w_6716 , w_6717 , w_6718 , w_6719 , w_6720 , w_6721 , w_6722 , w_6723 , w_6724 , w_6725 , 
		w_6726 , w_6727 , w_6728 , w_6729 , w_6730 , w_6731 , w_6732 , w_6733 , w_6734 , w_6735 , 
		w_6736 , w_6737 , w_6738 , w_6739 , w_6740 , w_6741 , w_6742 , w_6743 , w_6744 , w_6745 , 
		w_6746 , w_6747 , w_6748 , w_6749 , w_6750 , w_6751 , w_6752 , w_6753 , w_6754 , w_6755 , 
		w_6756 , w_6757 , w_6758 , w_6759 , w_6760 , w_6761 , w_6762 , w_6763 , w_6764 , w_6765 , 
		w_6766 , w_6767 , w_6768 , w_6769 , w_6770 , w_6771 , w_6772 , w_6773 , w_6774 , w_6775 , 
		w_6776 , w_6777 , w_6778 , w_6779 , w_6780 , w_6781 , w_6782 , w_6783 , w_6784 , w_6785 , 
		w_6786 , w_6787 , w_6788 , w_6789 , w_6790 , w_6791 , w_6792 , w_6793 , w_6794 , w_6795 , 
		w_6796 , w_6797 , w_6798 , w_6799 , w_6800 , w_6801 , w_6802 , w_6803 , w_6804 , w_6805 , 
		w_6806 , w_6807 , w_6808 , w_6809 , w_6810 , w_6811 , w_6812 , w_6813 , w_6814 , w_6815 , 
		w_6816 , w_6817 , w_6818 , w_6819 , w_6820 , w_6821 , w_6822 , w_6823 , w_6824 , w_6825 , 
		w_6826 , w_6827 , w_6828 , w_6829 , w_6830 , w_6831 , w_6832 , w_6833 , w_6834 , w_6835 , 
		w_6836 , w_6837 , w_6838 , w_6839 , w_6840 , w_6841 , w_6842 , w_6843 , w_6844 , w_6845 , 
		w_6846 , w_6847 , w_6848 , w_6849 , w_6850 , w_6851 , w_6852 , w_6853 , w_6854 , w_6855 , 
		w_6856 , w_6857 , w_6858 , w_6859 , w_6860 , w_6861 , w_6862 , w_6863 , w_6864 , w_6865 , 
		w_6866 , w_6867 , w_6868 , w_6869 , w_6870 , w_6871 , w_6872 , w_6873 , w_6874 , w_6875 , 
		w_6876 , w_6877 , w_6878 , w_6879 , w_6880 , w_6881 , w_6882 , w_6883 , w_6884 , w_6885 , 
		w_6886 , w_6887 , w_6888 , w_6889 , w_6890 , w_6891 , w_6892 , w_6893 , w_6894 , w_6895 , 
		w_6896 , w_6897 , w_6898 , w_6899 , w_6900 , w_6901 , w_6902 , w_6903 , w_6904 , w_6905 , 
		w_6906 , w_6907 , w_6908 , w_6909 , w_6910 , w_6911 , w_6912 , w_6913 , w_6914 , w_6915 , 
		w_6916 , w_6917 , w_6918 , w_6919 , w_6920 , w_6921 , w_6922 , w_6923 , w_6924 , w_6925 , 
		w_6926 , w_6927 , w_6928 , w_6929 , w_6930 , w_6931 , w_6932 , w_6933 , w_6934 , w_6935 , 
		w_6936 , w_6937 , w_6938 , w_6939 , w_6940 , w_6941 , w_6942 , w_6943 , w_6944 , w_6945 , 
		w_6946 , w_6947 , w_6948 , w_6949 , w_6950 , w_6951 , w_6952 , w_6953 , w_6954 , w_6955 , 
		w_6956 , w_6957 , w_6958 , w_6959 , w_6960 , w_6961 , w_6962 , w_6963 , w_6964 , w_6965 , 
		w_6966 , w_6967 , w_6968 , w_6969 , w_6970 , w_6971 , w_6972 , w_6973 , w_6974 , w_6975 , 
		w_6976 , w_6977 , w_6978 , w_6979 , w_6980 , w_6981 , w_6982 , w_6983 , w_6984 , w_6985 , 
		w_6986 , w_6987 , w_6988 , w_6989 , w_6990 , w_6991 , w_6992 , w_6993 , w_6994 , w_6995 , 
		w_6996 , w_6997 , w_6998 , w_6999 , w_7000 , w_7001 , w_7002 , w_7003 , w_7004 , w_7005 , 
		w_7006 , w_7007 , w_7008 , w_7009 , w_7010 , w_7011 , w_7012 , w_7013 , w_7014 , w_7015 , 
		w_7016 , w_7017 , w_7018 , w_7019 , w_7020 , w_7021 , w_7022 , w_7023 , w_7024 , w_7025 , 
		w_7026 , w_7027 , w_7028 , w_7029 , w_7030 , w_7031 , w_7032 , w_7033 , w_7034 , w_7035 , 
		w_7036 , w_7037 , w_7038 , w_7039 , w_7040 , w_7041 , w_7042 , w_7043 , w_7044 , w_7045 , 
		w_7046 , w_7047 , w_7048 , w_7049 , w_7050 , w_7051 , w_7052 , w_7053 , w_7054 , w_7055 , 
		w_7056 , w_7057 , w_7058 , w_7059 , w_7060 , w_7061 , w_7062 , w_7063 , w_7064 , w_7065 , 
		w_7066 , w_7067 , w_7068 , w_7069 , w_7070 , w_7071 , w_7072 , w_7073 , w_7074 , w_7075 , 
		w_7076 , w_7077 , w_7078 , w_7079 , w_7080 , w_7081 , w_7082 , w_7083 , w_7084 , w_7085 , 
		w_7086 , w_7087 , w_7088 , w_7089 , w_7090 , w_7091 , w_7092 , w_7093 , w_7094 , w_7095 , 
		w_7096 , w_7097 , w_7098 , w_7099 , w_7100 , w_7101 , w_7102 , w_7103 , w_7104 , w_7105 , 
		w_7106 , w_7107 , w_7108 , w_7109 , w_7110 , w_7111 , w_7112 , w_7113 , w_7114 , w_7115 , 
		w_7116 , w_7117 , w_7118 , w_7119 , w_7120 , w_7121 , w_7122 , w_7123 , w_7124 , w_7125 , 
		w_7126 , w_7127 , w_7128 , w_7129 , w_7130 , w_7131 , w_7132 , w_7133 , w_7134 , w_7135 , 
		w_7136 , w_7137 , w_7138 , w_7139 , w_7140 , w_7141 , w_7142 , w_7143 , w_7144 , w_7145 , 
		w_7146 , w_7147 , w_7148 , w_7149 , w_7150 , w_7151 , w_7152 , w_7153 , w_7154 , w_7155 , 
		w_7156 , w_7157 , w_7158 , w_7159 , w_7160 , w_7161 , w_7162 , w_7163 , w_7164 , w_7165 , 
		w_7166 , w_7167 , w_7168 , w_7169 , w_7170 , w_7171 , w_7172 , w_7173 , w_7174 , w_7175 , 
		w_7176 , w_7177 , w_7178 , w_7179 , w_7180 , w_7181 , w_7182 , w_7183 , w_7184 , w_7185 , 
		w_7186 , w_7187 , w_7188 , w_7189 , w_7190 , w_7191 , w_7192 , w_7193 , w_7194 , w_7195 , 
		w_7196 , w_7197 , w_7198 , w_7199 , w_7200 , w_7201 , w_7202 , w_7203 , w_7204 , w_7205 , 
		w_7206 , w_7207 , w_7208 , w_7209 , w_7210 , w_7211 , w_7212 , w_7213 , w_7214 , w_7215 , 
		w_7216 , w_7217 , w_7218 , w_7219 , w_7220 , w_7221 , w_7222 , w_7223 , w_7224 , w_7225 , 
		w_7226 , w_7227 , w_7228 , w_7229 , w_7230 , w_7231 , w_7232 , w_7233 , w_7234 , w_7235 , 
		w_7236 , w_7237 , w_7238 , w_7239 , w_7240 , w_7241 , w_7242 , w_7243 , w_7244 , w_7245 , 
		w_7246 , w_7247 , w_7248 , w_7249 , w_7250 , w_7251 , w_7252 , w_7253 , w_7254 , w_7255 , 
		w_7256 , w_7257 , w_7258 , w_7259 , w_7260 , w_7261 , w_7262 , w_7263 , w_7264 , w_7265 , 
		w_7266 , w_7267 , w_7268 , w_7269 , w_7270 , w_7271 , w_7272 , w_7273 , w_7274 , w_7275 , 
		w_7276 , w_7277 , w_7278 , w_7279 , w_7280 , w_7281 , w_7282 , w_7283 , w_7284 , w_7285 , 
		w_7286 , w_7287 , w_7288 , w_7289 , w_7290 , w_7291 , w_7292 , w_7293 , w_7294 , w_7295 , 
		w_7296 , w_7297 , w_7298 , w_7299 , w_7300 , w_7301 , w_7302 , w_7303 , w_7304 , w_7305 , 
		w_7306 , w_7307 , w_7308 , w_7309 , w_7310 , w_7311 , w_7312 , w_7313 , w_7314 , w_7315 , 
		w_7316 , w_7317 , w_7318 , w_7319 , w_7320 , w_7321 , w_7322 , w_7323 , w_7324 , w_7325 , 
		w_7326 , w_7327 , w_7328 , w_7329 , w_7330 , w_7331 , w_7332 , w_7333 , w_7334 , w_7335 , 
		w_7336 , w_7337 , w_7338 , w_7339 , w_7340 , w_7341 , w_7342 , w_7343 , w_7344 , w_7345 , 
		w_7346 , w_7347 , w_7348 , w_7349 , w_7350 , w_7351 , w_7352 , w_7353 , w_7354 , w_7355 , 
		w_7356 , w_7357 , w_7358 , w_7359 , w_7360 , w_7361 , w_7362 , w_7363 , w_7364 , w_7365 , 
		w_7366 , w_7367 , w_7368 , w_7369 , w_7370 , w_7371 , w_7372 , w_7373 , w_7374 , w_7375 , 
		w_7376 , w_7377 , w_7378 , w_7379 , w_7380 , w_7381 , w_7382 , w_7383 , w_7384 , w_7385 , 
		w_7386 , w_7387 , w_7388 , w_7389 , w_7390 , w_7391 , w_7392 , w_7393 , w_7394 , w_7395 , 
		w_7396 , w_7397 , w_7398 , w_7399 , w_7400 , w_7401 , w_7402 , w_7403 , w_7404 , w_7405 , 
		w_7406 , w_7407 , w_7408 , w_7409 , w_7410 , w_7411 , w_7412 , w_7413 , w_7414 , w_7415 , 
		w_7416 , w_7417 , w_7418 , w_7419 , w_7420 , w_7421 , w_7422 , w_7423 , w_7424 , w_7425 , 
		w_7426 , w_7427 , w_7428 , w_7429 , w_7430 , w_7431 , w_7432 , w_7433 , w_7434 , w_7435 , 
		w_7436 , w_7437 , w_7438 , w_7439 , w_7440 , w_7441 , w_7442 , w_7443 , w_7444 , w_7445 , 
		w_7446 , w_7447 , w_7448 , w_7449 , w_7450 , w_7451 , w_7452 , w_7453 , w_7454 , w_7455 , 
		w_7456 , w_7457 , w_7458 , w_7459 , w_7460 , w_7461 , w_7462 , w_7463 , w_7464 , w_7465 , 
		w_7466 , w_7467 , w_7468 , w_7469 , w_7470 , w_7471 , w_7472 , w_7473 , w_7474 , w_7475 , 
		w_7476 , w_7477 , w_7478 , w_7479 , w_7480 , w_7481 , w_7482 , w_7483 , w_7484 , w_7485 , 
		w_7486 , w_7487 , w_7488 , w_7489 , w_7490 , w_7491 , w_7492 , w_7493 , w_7494 , w_7495 , 
		w_7496 , w_7497 , w_7498 , w_7499 , w_7500 , w_7501 , w_7502 , w_7503 , w_7504 , w_7505 , 
		w_7506 , w_7507 , w_7508 , w_7509 , w_7510 , w_7511 , w_7512 , w_7513 , w_7514 , w_7515 , 
		w_7516 , w_7517 , w_7518 , w_7519 , w_7520 , w_7521 , w_7522 , w_7523 , w_7524 , w_7525 , 
		w_7526 , w_7527 , w_7528 , w_7529 , w_7530 , w_7531 , w_7532 , w_7533 , w_7534 , w_7535 , 
		w_7536 , w_7537 , w_7538 , w_7539 , w_7540 , w_7541 , w_7542 , w_7543 , w_7544 , w_7545 , 
		w_7546 , w_7547 , w_7548 , w_7549 , w_7550 , w_7551 , w_7552 , w_7553 , w_7554 , w_7555 , 
		w_7556 , w_7557 , w_7558 , w_7559 , w_7560 , w_7561 , w_7562 , w_7563 , w_7564 , w_7565 , 
		w_7566 , w_7567 , w_7568 , w_7569 , w_7570 , w_7571 , w_7572 , w_7573 , w_7574 , w_7575 , 
		w_7576 , w_7577 , w_7578 , w_7579 , w_7580 , w_7581 , w_7582 , w_7583 , w_7584 , w_7585 , 
		w_7586 , w_7587 , w_7588 , w_7589 , w_7590 , w_7591 , w_7592 , w_7593 , w_7594 , w_7595 , 
		w_7596 , w_7597 , w_7598 , w_7599 , w_7600 , w_7601 , w_7602 , w_7603 , w_7604 , w_7605 , 
		w_7606 , w_7607 , w_7608 , w_7609 , w_7610 , w_7611 , w_7612 , w_7613 , w_7614 , w_7615 , 
		w_7616 , w_7617 , w_7618 , w_7619 , w_7620 , w_7621 , w_7622 , w_7623 , w_7624 , w_7625 , 
		w_7626 , w_7627 , w_7628 , w_7629 , w_7630 , w_7631 , w_7632 , w_7633 , w_7634 , w_7635 , 
		w_7636 , w_7637 , w_7638 , w_7639 , w_7640 , w_7641 , w_7642 , w_7643 , w_7644 , w_7645 , 
		w_7646 , w_7647 , w_7648 , w_7649 , w_7650 , w_7651 , w_7652 , w_7653 , w_7654 , w_7655 , 
		w_7656 , w_7657 , w_7658 , w_7659 , w_7660 , w_7661 , w_7662 , w_7663 , w_7664 , w_7665 , 
		w_7666 , w_7667 , w_7668 , w_7669 , w_7670 , w_7671 , w_7672 , w_7673 , w_7674 , w_7675 , 
		w_7676 , w_7677 , w_7678 , w_7679 , w_7680 , w_7681 , w_7682 , w_7683 , w_7684 , w_7685 , 
		w_7686 , w_7687 , w_7688 , w_7689 , w_7690 , w_7691 , w_7692 , w_7693 , w_7694 , w_7695 , 
		w_7696 , w_7697 , w_7698 , w_7699 , w_7700 , w_7701 , w_7702 , w_7703 , w_7704 , w_7705 , 
		w_7706 , w_7707 , w_7708 , w_7709 , w_7710 , w_7711 , w_7712 , w_7713 , w_7714 , w_7715 , 
		w_7716 , w_7717 , w_7718 , w_7719 , w_7720 , w_7721 , w_7722 , w_7723 , w_7724 , w_7725 , 
		w_7726 , w_7727 , w_7728 , w_7729 , w_7730 , w_7731 , w_7732 , w_7733 , w_7734 , w_7735 , 
		w_7736 , w_7737 , w_7738 , w_7739 , w_7740 , w_7741 , w_7742 , w_7743 , w_7744 , w_7745 , 
		w_7746 , w_7747 , w_7748 , w_7749 , w_7750 , w_7751 , w_7752 , w_7753 , w_7754 , w_7755 , 
		w_7756 , w_7757 , w_7758 , w_7759 , w_7760 , w_7761 , w_7762 , w_7763 , w_7764 , w_7765 , 
		w_7766 , w_7767 , w_7768 , w_7769 , w_7770 , w_7771 , w_7772 , w_7773 , w_7774 , w_7775 , 
		w_7776 , w_7777 , w_7778 , w_7779 , w_7780 , w_7781 , w_7782 , w_7783 , w_7784 , w_7785 , 
		w_7786 , w_7787 , w_7788 , w_7789 , w_7790 , w_7791 , w_7792 , w_7793 , w_7794 , w_7795 , 
		w_7796 , w_7797 , w_7798 , w_7799 , w_7800 , w_7801 , w_7802 , w_7803 , w_7804 , w_7805 , 
		w_7806 , w_7807 , w_7808 , w_7809 , w_7810 , w_7811 , w_7812 , w_7813 , w_7814 , w_7815 , 
		w_7816 , w_7817 , w_7818 , w_7819 , w_7820 , w_7821 , w_7822 , w_7823 , w_7824 , w_7825 , 
		w_7826 , w_7827 , w_7828 , w_7829 , w_7830 , w_7831 , w_7832 , w_7833 , w_7834 , w_7835 , 
		w_7836 , w_7837 , w_7838 , w_7839 , w_7840 , w_7841 , w_7842 , w_7843 , w_7844 , w_7845 , 
		w_7846 , w_7847 , w_7848 , w_7849 , w_7850 , w_7851 , w_7852 , w_7853 , w_7854 , w_7855 , 
		w_7856 , w_7857 , w_7858 , w_7859 , w_7860 , w_7861 , w_7862 , w_7863 , w_7864 , w_7865 , 
		w_7866 , w_7867 , w_7868 , w_7869 , w_7870 , w_7871 , w_7872 , w_7873 , w_7874 , w_7875 , 
		w_7876 , w_7877 , w_7878 , w_7879 , w_7880 , w_7881 , w_7882 , w_7883 , w_7884 , w_7885 , 
		w_7886 , w_7887 , w_7888 , w_7889 , w_7890 , w_7891 , w_7892 , w_7893 , w_7894 , w_7895 , 
		w_7896 , w_7897 , w_7898 , w_7899 , w_7900 , w_7901 , w_7902 , w_7903 , w_7904 , w_7905 , 
		w_7906 , w_7907 , w_7908 , w_7909 , w_7910 , w_7911 , w_7912 , w_7913 , w_7914 , w_7915 , 
		w_7916 , w_7917 , w_7918 , w_7919 , w_7920 , w_7921 , w_7922 , w_7923 , w_7924 , w_7925 , 
		w_7926 , w_7927 , w_7928 , w_7929 , w_7930 , w_7931 , w_7932 , w_7933 , w_7934 , w_7935 , 
		w_7936 , w_7937 , w_7938 , w_7939 , w_7940 , w_7941 , w_7942 , w_7943 , w_7944 , w_7945 , 
		w_7946 , w_7947 , w_7948 , w_7949 , w_7950 , w_7951 , w_7952 , w_7953 , w_7954 , w_7955 , 
		w_7956 , w_7957 , w_7958 , w_7959 , w_7960 , w_7961 , w_7962 , w_7963 , w_7964 , w_7965 , 
		w_7966 , w_7967 , w_7968 , w_7969 , w_7970 , w_7971 , w_7972 , w_7973 , w_7974 , w_7975 , 
		w_7976 , w_7977 , w_7978 , w_7979 , w_7980 , w_7981 , w_7982 , w_7983 , w_7984 , w_7985 , 
		w_7986 , w_7987 , w_7988 , w_7989 , w_7990 , w_7991 , w_7992 , w_7993 , w_7994 , w_7995 , 
		w_7996 , w_7997 , w_7998 , w_7999 , w_8000 , w_8001 , w_8002 , w_8003 , w_8004 , w_8005 , 
		w_8006 , w_8007 , w_8008 , w_8009 , w_8010 , w_8011 , w_8012 , w_8013 , w_8014 , w_8015 , 
		w_8016 , w_8017 , w_8018 , w_8019 , w_8020 , w_8021 , w_8022 , w_8023 , w_8024 , w_8025 , 
		w_8026 , w_8027 , w_8028 , w_8029 , w_8030 , w_8031 , w_8032 , w_8033 , w_8034 , w_8035 , 
		w_8036 , w_8037 , w_8038 , w_8039 , w_8040 , w_8041 , w_8042 , w_8043 , w_8044 , w_8045 , 
		w_8046 , w_8047 , w_8048 , w_8049 , w_8050 , w_8051 , w_8052 , w_8053 , w_8054 , w_8055 , 
		w_8056 , w_8057 , w_8058 , w_8059 , w_8060 , w_8061 , w_8062 , w_8063 , w_8064 , w_8065 , 
		w_8066 , w_8067 , w_8068 , w_8069 , w_8070 , w_8071 , w_8072 , w_8073 , w_8074 , w_8075 , 
		w_8076 , w_8077 , w_8078 , w_8079 , w_8080 , w_8081 , w_8082 , w_8083 , w_8084 , w_8085 , 
		w_8086 , w_8087 , w_8088 , w_8089 , w_8090 , w_8091 , w_8092 , w_8093 , w_8094 , w_8095 , 
		w_8096 , w_8097 , w_8098 , w_8099 , w_8100 , w_8101 , w_8102 , w_8103 , w_8104 , w_8105 , 
		w_8106 , w_8107 , w_8108 , w_8109 , w_8110 , w_8111 , w_8112 , w_8113 , w_8114 , w_8115 , 
		w_8116 , w_8117 , w_8118 , w_8119 , w_8120 , w_8121 , w_8122 , w_8123 , w_8124 , w_8125 , 
		w_8126 , w_8127 , w_8128 , w_8129 , w_8130 , w_8131 , w_8132 , w_8133 , w_8134 , w_8135 , 
		w_8136 , w_8137 , w_8138 , w_8139 , w_8140 , w_8141 , w_8142 , w_8143 , w_8144 , w_8145 , 
		w_8146 , w_8147 , w_8148 , w_8149 , w_8150 , w_8151 , w_8152 , w_8153 , w_8154 , w_8155 , 
		w_8156 , w_8157 , w_8158 , w_8159 , w_8160 , w_8161 , w_8162 , w_8163 , w_8164 , w_8165 , 
		w_8166 , w_8167 , w_8168 , w_8169 , w_8170 , w_8171 , w_8172 , w_8173 , w_8174 , w_8175 , 
		w_8176 , w_8177 , w_8178 , w_8179 , w_8180 , w_8181 , w_8182 , w_8183 , w_8184 , w_8185 , 
		w_8186 , w_8187 , w_8188 , w_8189 , w_8190 , w_8191 , w_8192 , w_8193 , w_8194 , w_8195 , 
		w_8196 , w_8197 , w_8198 , w_8199 , w_8200 , w_8201 , w_8202 , w_8203 , w_8204 , w_8205 , 
		w_8206 , w_8207 , w_8208 , w_8209 , w_8210 , w_8211 , w_8212 , w_8213 , w_8214 , w_8215 , 
		w_8216 , w_8217 , w_8218 , w_8219 , w_8220 , w_8221 , w_8222 , w_8223 , w_8224 , w_8225 , 
		w_8226 , w_8227 , w_8228 , w_8229 , w_8230 , w_8231 , w_8232 , w_8233 , w_8234 , w_8235 , 
		w_8236 , w_8237 , w_8238 , w_8239 , w_8240 , w_8241 , w_8242 , w_8243 , w_8244 , w_8245 , 
		w_8246 , w_8247 , w_8248 , w_8249 , w_8250 , w_8251 , w_8252 , w_8253 , w_8254 , w_8255 , 
		w_8256 , w_8257 , w_8258 , w_8259 , w_8260 , w_8261 , w_8262 , w_8263 , w_8264 , w_8265 , 
		w_8266 , w_8267 , w_8268 , w_8269 , w_8270 , w_8271 , w_8272 , w_8273 , w_8274 , w_8275 , 
		w_8276 , w_8277 , w_8278 , w_8279 , w_8280 , w_8281 , w_8282 , w_8283 , w_8284 , w_8285 , 
		w_8286 , w_8287 , w_8288 , w_8289 , w_8290 , w_8291 , w_8292 , w_8293 , w_8294 , w_8295 , 
		w_8296 , w_8297 , w_8298 , w_8299 , w_8300 , w_8301 , w_8302 , w_8303 , w_8304 , w_8305 , 
		w_8306 , w_8307 , w_8308 , w_8309 , w_8310 , w_8311 , w_8312 , w_8313 , w_8314 , w_8315 , 
		w_8316 , w_8317 , w_8318 , w_8319 , w_8320 , w_8321 , w_8322 , w_8323 , w_8324 , w_8325 , 
		w_8326 , w_8327 , w_8328 , w_8329 , w_8330 , w_8331 , w_8332 , w_8333 , w_8334 , w_8335 , 
		w_8336 , w_8337 , w_8338 , w_8339 , w_8340 , w_8341 , w_8342 , w_8343 , w_8344 , w_8345 , 
		w_8346 , w_8347 , w_8348 , w_8349 , w_8350 , w_8351 , w_8352 , w_8353 , w_8354 , w_8355 , 
		w_8356 , w_8357 , w_8358 , w_8359 , w_8360 , w_8361 , w_8362 , w_8363 , w_8364 , w_8365 , 
		w_8366 , w_8367 , w_8368 , w_8369 , w_8370 , w_8371 , w_8372 , w_8373 , w_8374 , w_8375 , 
		w_8376 , w_8377 , w_8378 , w_8379 , w_8380 , w_8381 , w_8382 , w_8383 , w_8384 , w_8385 , 
		w_8386 , w_8387 , w_8388 , w_8389 , w_8390 , w_8391 , w_8392 , w_8393 , w_8394 , w_8395 , 
		w_8396 , w_8397 , w_8398 , w_8399 , w_8400 , w_8401 , w_8402 , w_8403 , w_8404 , w_8405 , 
		w_8406 , w_8407 , w_8408 , w_8409 , w_8410 , w_8411 , w_8412 , w_8413 , w_8414 , w_8415 , 
		w_8416 , w_8417 , w_8418 , w_8419 , w_8420 , w_8421 , w_8422 , w_8423 , w_8424 , w_8425 , 
		w_8426 , w_8427 , w_8428 , w_8429 , w_8430 , w_8431 , w_8432 , w_8433 , w_8434 , w_8435 , 
		w_8436 , w_8437 , w_8438 , w_8439 , w_8440 , w_8441 , w_8442 , w_8443 , w_8444 , w_8445 , 
		w_8446 , w_8447 , w_8448 , w_8449 , w_8450 , w_8451 , w_8452 , w_8453 , w_8454 , w_8455 , 
		w_8456 , w_8457 , w_8458 , w_8459 , w_8460 , w_8461 , w_8462 , w_8463 , w_8464 , w_8465 , 
		w_8466 , w_8467 , w_8468 , w_8469 , w_8470 , w_8471 , w_8472 , w_8473 , w_8474 , w_8475 , 
		w_8476 , w_8477 , w_8478 , w_8479 , w_8480 , w_8481 , w_8482 , w_8483 , w_8484 , w_8485 , 
		w_8486 , w_8487 , w_8488 , w_8489 , w_8490 , w_8491 , w_8492 , w_8493 , w_8494 , w_8495 , 
		w_8496 , w_8497 , w_8498 , w_8499 , w_8500 , w_8501 , w_8502 , w_8503 , w_8504 , w_8505 , 
		w_8506 , w_8507 , w_8508 , w_8509 , w_8510 , w_8511 , w_8512 , w_8513 , w_8514 , w_8515 , 
		w_8516 , w_8517 , w_8518 , w_8519 , w_8520 , w_8521 , w_8522 , w_8523 , w_8524 , w_8525 , 
		w_8526 , w_8527 , w_8528 , w_8529 , w_8530 , w_8531 , w_8532 , w_8533 , w_8534 , w_8535 , 
		w_8536 , w_8537 , w_8538 , w_8539 , w_8540 , w_8541 , w_8542 , w_8543 , w_8544 , w_8545 , 
		w_8546 , w_8547 , w_8548 , w_8549 , w_8550 , w_8551 , w_8552 , w_8553 , w_8554 , w_8555 , 
		w_8556 , w_8557 , w_8558 , w_8559 , w_8560 , w_8561 , w_8562 , w_8563 , w_8564 , w_8565 , 
		w_8566 , w_8567 , w_8568 , w_8569 , w_8570 , w_8571 , w_8572 , w_8573 , w_8574 , w_8575 , 
		w_8576 , w_8577 , w_8578 , w_8579 , w_8580 , w_8581 , w_8582 , w_8583 , w_8584 , w_8585 , 
		w_8586 , w_8587 , w_8588 , w_8589 , w_8590 , w_8591 , w_8592 , w_8593 , w_8594 , w_8595 , 
		w_8596 , w_8597 , w_8598 , w_8599 , w_8600 , w_8601 , w_8602 , w_8603 , w_8604 , w_8605 , 
		w_8606 , w_8607 , w_8608 , w_8609 , w_8610 , w_8611 , w_8612 , w_8613 , w_8614 , w_8615 , 
		w_8616 , w_8617 , w_8618 , w_8619 , w_8620 , w_8621 , w_8622 , w_8623 , w_8624 , w_8625 , 
		w_8626 , w_8627 , w_8628 , w_8629 , w_8630 , w_8631 , w_8632 , w_8633 , w_8634 , w_8635 , 
		w_8636 , w_8637 , w_8638 , w_8639 , w_8640 , w_8641 , w_8642 , w_8643 , w_8644 , w_8645 , 
		w_8646 , w_8647 , w_8648 , w_8649 , w_8650 , w_8651 , w_8652 , w_8653 , w_8654 , w_8655 , 
		w_8656 , w_8657 , w_8658 , w_8659 , w_8660 , w_8661 , w_8662 , w_8663 , w_8664 , w_8665 , 
		w_8666 , w_8667 , w_8668 , w_8669 , w_8670 , w_8671 , w_8672 , w_8673 , w_8674 , w_8675 , 
		w_8676 , w_8677 , w_8678 , w_8679 , w_8680 , w_8681 , w_8682 , w_8683 , w_8684 , w_8685 , 
		w_8686 , w_8687 , w_8688 , w_8689 , w_8690 , w_8691 , w_8692 , w_8693 , w_8694 , w_8695 , 
		w_8696 , w_8697 , w_8698 , w_8699 , w_8700 , w_8701 , w_8702 , w_8703 , w_8704 , w_8705 , 
		w_8706 , w_8707 , w_8708 , w_8709 , w_8710 , w_8711 , w_8712 , w_8713 , w_8714 , w_8715 , 
		w_8716 , w_8717 , w_8718 , w_8719 , w_8720 , w_8721 , w_8722 , w_8723 , w_8724 , w_8725 , 
		w_8726 , w_8727 , w_8728 , w_8729 , w_8730 , w_8731 , w_8732 , w_8733 , w_8734 , w_8735 , 
		w_8736 , w_8737 , w_8738 , w_8739 , w_8740 , w_8741 , w_8742 , w_8743 , w_8744 , w_8745 , 
		w_8746 , w_8747 , w_8748 , w_8749 , w_8750 , w_8751 , w_8752 , w_8753 , w_8754 , w_8755 , 
		w_8756 , w_8757 , w_8758 , w_8759 , w_8760 , w_8761 , w_8762 , w_8763 , w_8764 , w_8765 , 
		w_8766 , w_8767 , w_8768 , w_8769 , w_8770 , w_8771 , w_8772 , w_8773 , w_8774 , w_8775 , 
		w_8776 , w_8777 , w_8778 , w_8779 , w_8780 , w_8781 , w_8782 , w_8783 , w_8784 , w_8785 , 
		w_8786 , w_8787 , w_8788 , w_8789 , w_8790 , w_8791 , w_8792 , w_8793 , w_8794 , w_8795 , 
		w_8796 , w_8797 , w_8798 , w_8799 , w_8800 , w_8801 , w_8802 , w_8803 , w_8804 , w_8805 , 
		w_8806 , w_8807 , w_8808 , w_8809 , w_8810 , w_8811 , w_8812 , w_8813 , w_8814 , w_8815 , 
		w_8816 , w_8817 , w_8818 , w_8819 , w_8820 , w_8821 , w_8822 , w_8823 , w_8824 , w_8825 , 
		w_8826 , w_8827 , w_8828 , w_8829 , w_8830 , w_8831 , w_8832 , w_8833 , w_8834 , w_8835 , 
		w_8836 , w_8837 , w_8838 , w_8839 , w_8840 , w_8841 , w_8842 , w_8843 , w_8844 , w_8845 , 
		w_8846 , w_8847 , w_8848 , w_8849 , w_8850 , w_8851 , w_8852 , w_8853 , w_8854 , w_8855 , 
		w_8856 , w_8857 , w_8858 , w_8859 , w_8860 , w_8861 , w_8862 , w_8863 , w_8864 , w_8865 , 
		w_8866 , w_8867 , w_8868 , w_8869 , w_8870 , w_8871 , w_8872 , w_8873 , w_8874 , w_8875 , 
		w_8876 , w_8877 , w_8878 , w_8879 , w_8880 , w_8881 , w_8882 , w_8883 , w_8884 , w_8885 , 
		w_8886 , w_8887 , w_8888 , w_8889 , w_8890 , w_8891 , w_8892 , w_8893 , w_8894 , w_8895 , 
		w_8896 , w_8897 , w_8898 , w_8899 , w_8900 , w_8901 , w_8902 , w_8903 , w_8904 , w_8905 , 
		w_8906 , w_8907 , w_8908 , w_8909 , w_8910 , w_8911 , w_8912 , w_8913 , w_8914 , w_8915 , 
		w_8916 , w_8917 , w_8918 , w_8919 , w_8920 , w_8921 , w_8922 , w_8923 , w_8924 , w_8925 , 
		w_8926 , w_8927 , w_8928 , w_8929 , w_8930 , w_8931 , w_8932 , w_8933 , w_8934 , w_8935 , 
		w_8936 , w_8937 , w_8938 , w_8939 , w_8940 , w_8941 , w_8942 , w_8943 , w_8944 , w_8945 , 
		w_8946 , w_8947 , w_8948 , w_8949 , w_8950 , w_8951 , w_8952 , w_8953 , w_8954 , w_8955 , 
		w_8956 , w_8957 , w_8958 , w_8959 , w_8960 , w_8961 , w_8962 , w_8963 , w_8964 , w_8965 , 
		w_8966 , w_8967 , w_8968 , w_8969 , w_8970 , w_8971 , w_8972 , w_8973 , w_8974 , w_8975 , 
		w_8976 , w_8977 , w_8978 , w_8979 , w_8980 , w_8981 , w_8982 , w_8983 , w_8984 , w_8985 , 
		w_8986 , w_8987 , w_8988 , w_8989 , w_8990 , w_8991 , w_8992 , w_8993 , w_8994 , w_8995 , 
		w_8996 , w_8997 , w_8998 , w_8999 , w_9000 , w_9001 , w_9002 , w_9003 , w_9004 , w_9005 , 
		w_9006 , w_9007 , w_9008 , w_9009 , w_9010 , w_9011 , w_9012 , w_9013 , w_9014 , w_9015 , 
		w_9016 , w_9017 , w_9018 , w_9019 , w_9020 , w_9021 , w_9022 , w_9023 , w_9024 , w_9025 , 
		w_9026 , w_9027 , w_9028 , w_9029 , w_9030 , w_9031 , w_9032 , w_9033 , w_9034 , w_9035 , 
		w_9036 , w_9037 , w_9038 , w_9039 , w_9040 , w_9041 , w_9042 , w_9043 , w_9044 , w_9045 , 
		w_9046 , w_9047 , w_9048 , w_9049 , w_9050 , w_9051 , w_9052 , w_9053 , w_9054 , w_9055 , 
		w_9056 , w_9057 , w_9058 , w_9059 , w_9060 , w_9061 , w_9062 , w_9063 , w_9064 , w_9065 , 
		w_9066 , w_9067 , w_9068 , w_9069 , w_9070 , w_9071 , w_9072 , w_9073 , w_9074 , w_9075 , 
		w_9076 , w_9077 , w_9078 , w_9079 , w_9080 , w_9081 , w_9082 , w_9083 , w_9084 , w_9085 , 
		w_9086 , w_9087 , w_9088 , w_9089 , w_9090 , w_9091 , w_9092 , w_9093 , w_9094 , w_9095 , 
		w_9096 , w_9097 , w_9098 , w_9099 , w_9100 , w_9101 , w_9102 , w_9103 , w_9104 , w_9105 , 
		w_9106 , w_9107 , w_9108 , w_9109 , w_9110 , w_9111 , w_9112 , w_9113 , w_9114 , w_9115 , 
		w_9116 , w_9117 , w_9118 , w_9119 , w_9120 , w_9121 , w_9122 , w_9123 , w_9124 , w_9125 , 
		w_9126 , w_9127 , w_9128 , w_9129 , w_9130 , w_9131 , w_9132 , w_9133 , w_9134 , w_9135 , 
		w_9136 , w_9137 , w_9138 , w_9139 , w_9140 , w_9141 , w_9142 , w_9143 , w_9144 , w_9145 , 
		w_9146 , w_9147 , w_9148 , w_9149 , w_9150 , w_9151 , w_9152 , w_9153 , w_9154 , w_9155 , 
		w_9156 , w_9157 , w_9158 , w_9159 , w_9160 , w_9161 , w_9162 , w_9163 , w_9164 , w_9165 , 
		w_9166 , w_9167 , w_9168 , w_9169 , w_9170 , w_9171 , w_9172 , w_9173 , w_9174 , w_9175 , 
		w_9176 , w_9177 , w_9178 , w_9179 , w_9180 , w_9181 , w_9182 , w_9183 , w_9184 , w_9185 , 
		w_9186 , w_9187 , w_9188 , w_9189 , w_9190 , w_9191 , w_9192 , w_9193 , w_9194 , w_9195 , 
		w_9196 , w_9197 , w_9198 , w_9199 , w_9200 , w_9201 , w_9202 , w_9203 , w_9204 , w_9205 , 
		w_9206 , w_9207 , w_9208 , w_9209 , w_9210 , w_9211 , w_9212 , w_9213 , w_9214 , w_9215 , 
		w_9216 , w_9217 , w_9218 , w_9219 , w_9220 , w_9221 , w_9222 , w_9223 , w_9224 , w_9225 , 
		w_9226 , w_9227 , w_9228 , w_9229 , w_9230 , w_9231 , w_9232 , w_9233 , w_9234 , w_9235 , 
		w_9236 , w_9237 , w_9238 , w_9239 , w_9240 , w_9241 , w_9242 , w_9243 , w_9244 , w_9245 , 
		w_9246 , w_9247 , w_9248 , w_9249 , w_9250 , w_9251 , w_9252 , w_9253 , w_9254 , w_9255 , 
		w_9256 , w_9257 , w_9258 , w_9259 , w_9260 , w_9261 , w_9262 , w_9263 , w_9264 , w_9265 , 
		w_9266 , w_9267 , w_9268 , w_9269 , w_9270 , w_9271 , w_9272 , w_9273 , w_9274 , w_9275 , 
		w_9276 , w_9277 , w_9278 , w_9279 , w_9280 , w_9281 , w_9282 , w_9283 , w_9284 , w_9285 , 
		w_9286 , w_9287 , w_9288 , w_9289 , w_9290 , w_9291 , w_9292 , w_9293 , w_9294 , w_9295 , 
		w_9296 , w_9297 , w_9298 , w_9299 , w_9300 , w_9301 , w_9302 , w_9303 , w_9304 , w_9305 , 
		w_9306 , w_9307 , w_9308 , w_9309 , w_9310 , w_9311 , w_9312 , w_9313 , w_9314 , w_9315 , 
		w_9316 , w_9317 , w_9318 , w_9319 , w_9320 , w_9321 , w_9322 , w_9323 , w_9324 , w_9325 , 
		w_9326 , w_9327 , w_9328 , w_9329 , w_9330 , w_9331 , w_9332 , w_9333 , w_9334 , w_9335 , 
		w_9336 , w_9337 , w_9338 , w_9339 , w_9340 , w_9341 , w_9342 , w_9343 , w_9344 , w_9345 , 
		w_9346 , w_9347 , w_9348 , w_9349 , w_9350 , w_9351 , w_9352 , w_9353 , w_9354 , w_9355 , 
		w_9356 , w_9357 , w_9358 , w_9359 , w_9360 , w_9361 , w_9362 , w_9363 , w_9364 , w_9365 , 
		w_9366 , w_9367 , w_9368 , w_9369 , w_9370 , w_9371 , w_9372 , w_9373 , w_9374 , w_9375 , 
		w_9376 , w_9377 , w_9378 , w_9379 , w_9380 , w_9381 , w_9382 , w_9383 , w_9384 , w_9385 , 
		w_9386 , w_9387 , w_9388 , w_9389 , w_9390 , w_9391 , w_9392 , w_9393 , w_9394 , w_9395 , 
		w_9396 , w_9397 , w_9398 , w_9399 , w_9400 , w_9401 , w_9402 , w_9403 , w_9404 , w_9405 , 
		w_9406 , w_9407 , w_9408 , w_9409 , w_9410 , w_9411 , w_9412 , w_9413 , w_9414 , w_9415 , 
		w_9416 , w_9417 , w_9418 , w_9419 , w_9420 , w_9421 , w_9422 , w_9423 , w_9424 , w_9425 , 
		w_9426 , w_9427 , w_9428 , w_9429 , w_9430 , w_9431 , w_9432 , w_9433 , w_9434 , w_9435 , 
		w_9436 , w_9437 , w_9438 , w_9439 , w_9440 , w_9441 , w_9442 , w_9443 , w_9444 , w_9445 , 
		w_9446 , w_9447 , w_9448 , w_9449 , w_9450 , w_9451 , w_9452 , w_9453 , w_9454 , w_9455 , 
		w_9456 , w_9457 , w_9458 , w_9459 , w_9460 , w_9461 , w_9462 , w_9463 , w_9464 , w_9465 , 
		w_9466 , w_9467 , w_9468 , w_9469 , w_9470 , w_9471 , w_9472 , w_9473 , w_9474 , w_9475 , 
		w_9476 , w_9477 , w_9478 , w_9479 , w_9480 , w_9481 , w_9482 , w_9483 , w_9484 , w_9485 , 
		w_9486 , w_9487 , w_9488 , w_9489 , w_9490 , w_9491 , w_9492 , w_9493 , w_9494 , w_9495 , 
		w_9496 , w_9497 , w_9498 , w_9499 , w_9500 , w_9501 , w_9502 , w_9503 , w_9504 , w_9505 , 
		w_9506 , w_9507 , w_9508 , w_9509 , w_9510 , w_9511 , w_9512 , w_9513 , w_9514 , w_9515 , 
		w_9516 , w_9517 , w_9518 , w_9519 , w_9520 , w_9521 , w_9522 , w_9523 , w_9524 , w_9525 , 
		w_9526 , w_9527 , w_9528 , w_9529 , w_9530 , w_9531 , w_9532 , w_9533 , w_9534 , w_9535 , 
		w_9536 , w_9537 , w_9538 , w_9539 , w_9540 , w_9541 , w_9542 , w_9543 , w_9544 , w_9545 , 
		w_9546 , w_9547 , w_9548 , w_9549 , w_9550 , w_9551 , w_9552 , w_9553 , w_9554 , w_9555 , 
		w_9556 , w_9557 , w_9558 , w_9559 , w_9560 , w_9561 , w_9562 , w_9563 , w_9564 , w_9565 , 
		w_9566 , w_9567 , w_9568 , w_9569 , w_9570 , w_9571 , w_9572 , w_9573 , w_9574 , w_9575 , 
		w_9576 , w_9577 , w_9578 , w_9579 , w_9580 , w_9581 , w_9582 , w_9583 , w_9584 , w_9585 , 
		w_9586 , w_9587 , w_9588 , w_9589 , w_9590 , w_9591 , w_9592 , w_9593 , w_9594 , w_9595 , 
		w_9596 , w_9597 , w_9598 , w_9599 , w_9600 , w_9601 , w_9602 , w_9603 , w_9604 , w_9605 , 
		w_9606 , w_9607 , w_9608 , w_9609 , w_9610 , w_9611 , w_9612 , w_9613 , w_9614 , w_9615 , 
		w_9616 , w_9617 , w_9618 , w_9619 , w_9620 , w_9621 , w_9622 , w_9623 , w_9624 , w_9625 , 
		w_9626 , w_9627 , w_9628 , w_9629 , w_9630 , w_9631 , w_9632 , w_9633 , w_9634 , w_9635 , 
		w_9636 , w_9637 , w_9638 , w_9639 , w_9640 , w_9641 , w_9642 , w_9643 , w_9644 , w_9645 , 
		w_9646 , w_9647 , w_9648 , w_9649 , w_9650 , w_9651 , w_9652 , w_9653 , w_9654 , w_9655 , 
		w_9656 , w_9657 , w_9658 , w_9659 , w_9660 , w_9661 , w_9662 , w_9663 , w_9664 , w_9665 , 
		w_9666 , w_9667 , w_9668 , w_9669 , w_9670 , w_9671 , w_9672 , w_9673 , w_9674 , w_9675 , 
		w_9676 , w_9677 , w_9678 , w_9679 , w_9680 , w_9681 , w_9682 , w_9683 , w_9684 , w_9685 , 
		w_9686 , w_9687 , w_9688 , w_9689 , w_9690 , w_9691 , w_9692 , w_9693 , w_9694 , w_9695 , 
		w_9696 , w_9697 , w_9698 , w_9699 , w_9700 , w_9701 , w_9702 , w_9703 , w_9704 , w_9705 , 
		w_9706 , w_9707 , w_9708 , w_9709 , w_9710 , w_9711 , w_9712 , w_9713 , w_9714 , w_9715 , 
		w_9716 , w_9717 , w_9718 , w_9719 , w_9720 , w_9721 , w_9722 , w_9723 , w_9724 , w_9725 , 
		w_9726 , w_9727 , w_9728 , w_9729 , w_9730 , w_9731 , w_9732 , w_9733 , w_9734 , w_9735 , 
		w_9736 , w_9737 , w_9738 , w_9739 , w_9740 , w_9741 , w_9742 , w_9743 , w_9744 , w_9745 , 
		w_9746 , w_9747 , w_9748 , w_9749 , w_9750 , w_9751 , w_9752 , w_9753 , w_9754 , w_9755 , 
		w_9756 , w_9757 , w_9758 , w_9759 , w_9760 , w_9761 , w_9762 , w_9763 , w_9764 , w_9765 , 
		w_9766 , w_9767 , w_9768 , w_9769 , w_9770 , w_9771 , w_9772 , w_9773 , w_9774 , w_9775 , 
		w_9776 , w_9777 , w_9778 , w_9779 , w_9780 , w_9781 , w_9782 , w_9783 , w_9784 , w_9785 , 
		w_9786 , w_9787 , w_9788 , w_9789 , w_9790 , w_9791 , w_9792 , w_9793 , w_9794 , w_9795 , 
		w_9796 , w_9797 , w_9798 , w_9799 , w_9800 , w_9801 , w_9802 , w_9803 , w_9804 , w_9805 , 
		w_9806 , w_9807 , w_9808 , w_9809 , w_9810 , w_9811 , w_9812 , w_9813 , w_9814 , w_9815 , 
		w_9816 , w_9817 , w_9818 , w_9819 , w_9820 , w_9821 , w_9822 , w_9823 , w_9824 , w_9825 , 
		w_9826 , w_9827 , w_9828 , w_9829 , w_9830 , w_9831 , w_9832 , w_9833 , w_9834 , w_9835 , 
		w_9836 , w_9837 , w_9838 , w_9839 , w_9840 , w_9841 , w_9842 , w_9843 , w_9844 , w_9845 , 
		w_9846 , w_9847 , w_9848 , w_9849 , w_9850 , w_9851 , w_9852 , w_9853 , w_9854 , w_9855 , 
		w_9856 , w_9857 , w_9858 , w_9859 , w_9860 , w_9861 , w_9862 , w_9863 , w_9864 , w_9865 , 
		w_9866 , w_9867 , w_9868 , w_9869 , w_9870 , w_9871 , w_9872 , w_9873 , w_9874 , w_9875 , 
		w_9876 , w_9877 , w_9878 , w_9879 , w_9880 , w_9881 , w_9882 , w_9883 , w_9884 , w_9885 , 
		w_9886 , w_9887 , w_9888 , w_9889 , w_9890 , w_9891 , w_9892 , w_9893 , w_9894 , w_9895 , 
		w_9896 , w_9897 , w_9898 , w_9899 , w_9900 , w_9901 , w_9902 , w_9903 , w_9904 , w_9905 , 
		w_9906 , w_9907 , w_9908 , w_9909 , w_9910 , w_9911 , w_9912 , w_9913 , w_9914 , w_9915 , 
		w_9916 , w_9917 , w_9918 , w_9919 , w_9920 , w_9921 , w_9922 , w_9923 , w_9924 , w_9925 , 
		w_9926 , w_9927 , w_9928 , w_9929 , w_9930 , w_9931 , w_9932 , w_9933 , w_9934 , w_9935 , 
		w_9936 , w_9937 , w_9938 , w_9939 , w_9940 , w_9941 , w_9942 , w_9943 , w_9944 , w_9945 , 
		w_9946 , w_9947 , w_9948 , w_9949 , w_9950 , w_9951 , w_9952 , w_9953 , w_9954 , w_9955 , 
		w_9956 , w_9957 , w_9958 , w_9959 , w_9960 , w_9961 , w_9962 , w_9963 , w_9964 , w_9965 , 
		w_9966 , w_9967 , w_9968 , w_9969 , w_9970 , w_9971 , w_9972 , w_9973 , w_9974 , w_9975 , 
		w_9976 , w_9977 , w_9978 , w_9979 , w_9980 , w_9981 , w_9982 , w_9983 , w_9984 , w_9985 , 
		w_9986 , w_9987 , w_9988 , w_9989 , w_9990 , w_9991 , w_9992 , w_9993 , w_9994 , w_9995 , 
		w_9996 , w_9997 , w_9998 , w_9999 , w_10000 , w_10001 , w_10002 , w_10003 , w_10004 , w_10005 , 
		w_10006 , w_10007 , w_10008 , w_10009 , w_10010 , w_10011 , w_10012 , w_10013 , w_10014 , w_10015 , 
		w_10016 , w_10017 , w_10018 , w_10019 , w_10020 , w_10021 , w_10022 , w_10023 , w_10024 , w_10025 , 
		w_10026 , w_10027 , w_10028 , w_10029 , w_10030 , w_10031 , w_10032 , w_10033 , w_10034 , w_10035 , 
		w_10036 , w_10037 , w_10038 , w_10039 , w_10040 , w_10041 , w_10042 , w_10043 , w_10044 , w_10045 , 
		w_10046 , w_10047 , w_10048 , w_10049 , w_10050 , w_10051 , w_10052 , w_10053 , w_10054 , w_10055 , 
		w_10056 , w_10057 , w_10058 , w_10059 , w_10060 , w_10061 , w_10062 , w_10063 , w_10064 , w_10065 , 
		w_10066 , w_10067 , w_10068 , w_10069 , w_10070 , w_10071 , w_10072 , w_10073 , w_10074 , w_10075 , 
		w_10076 , w_10077 , w_10078 , w_10079 , w_10080 , w_10081 , w_10082 , w_10083 , w_10084 , w_10085 , 
		w_10086 , w_10087 , w_10088 , w_10089 , w_10090 , w_10091 , w_10092 , w_10093 , w_10094 , w_10095 , 
		w_10096 , w_10097 , w_10098 , w_10099 , w_10100 , w_10101 , w_10102 , w_10103 , w_10104 , w_10105 , 
		w_10106 , w_10107 , w_10108 , w_10109 , w_10110 , w_10111 , w_10112 , w_10113 , w_10114 , w_10115 , 
		w_10116 , w_10117 , w_10118 , w_10119 , w_10120 , w_10121 , w_10122 , w_10123 , w_10124 , w_10125 , 
		w_10126 , w_10127 , w_10128 , w_10129 , w_10130 , w_10131 , w_10132 , w_10133 , w_10134 , w_10135 , 
		w_10136 , w_10137 , w_10138 , w_10139 , w_10140 , w_10141 , w_10142 , w_10143 , w_10144 , w_10145 , 
		w_10146 , w_10147 , w_10148 , w_10149 , w_10150 , w_10151 , w_10152 , w_10153 , w_10154 , w_10155 , 
		w_10156 , w_10157 , w_10158 , w_10159 , w_10160 , w_10161 , w_10162 , w_10163 , w_10164 , w_10165 , 
		w_10166 , w_10167 , w_10168 , w_10169 , w_10170 , w_10171 , w_10172 , w_10173 , w_10174 , w_10175 , 
		w_10176 , w_10177 , w_10178 , w_10179 , w_10180 , w_10181 , w_10182 , w_10183 , w_10184 , w_10185 , 
		w_10186 , w_10187 , w_10188 , w_10189 , w_10190 , w_10191 , w_10192 , w_10193 , w_10194 , w_10195 , 
		w_10196 , w_10197 , w_10198 , w_10199 , w_10200 , w_10201 , w_10202 , w_10203 , w_10204 , w_10205 , 
		w_10206 , w_10207 , w_10208 , w_10209 , w_10210 , w_10211 , w_10212 , w_10213 , w_10214 , w_10215 , 
		w_10216 , w_10217 , w_10218 , w_10219 , w_10220 , w_10221 , w_10222 , w_10223 , w_10224 , w_10225 , 
		w_10226 , w_10227 , w_10228 , w_10229 , w_10230 , w_10231 , w_10232 , w_10233 , w_10234 , w_10235 , 
		w_10236 , w_10237 , w_10238 , w_10239 , w_10240 , w_10241 , w_10242 , w_10243 , w_10244 , w_10245 , 
		w_10246 , w_10247 , w_10248 , w_10249 , w_10250 , w_10251 , w_10252 , w_10253 , w_10254 , w_10255 , 
		w_10256 , w_10257 , w_10258 , w_10259 , w_10260 , w_10261 , w_10262 , w_10263 , w_10264 , w_10265 , 
		w_10266 , w_10267 , w_10268 , w_10269 , w_10270 , w_10271 , w_10272 , w_10273 , w_10274 , w_10275 , 
		w_10276 , w_10277 , w_10278 , w_10279 , w_10280 , w_10281 , w_10282 , w_10283 , w_10284 , w_10285 , 
		w_10286 , w_10287 , w_10288 , w_10289 , w_10290 , w_10291 , w_10292 , w_10293 , w_10294 , w_10295 , 
		w_10296 , w_10297 , w_10298 , w_10299 , w_10300 , w_10301 , w_10302 , w_10303 , w_10304 , w_10305 , 
		w_10306 , w_10307 , w_10308 , w_10309 , w_10310 , w_10311 , w_10312 , w_10313 , w_10314 , w_10315 , 
		w_10316 , w_10317 , w_10318 , w_10319 , w_10320 , w_10321 , w_10322 , w_10323 , w_10324 , w_10325 , 
		w_10326 , w_10327 , w_10328 , w_10329 , w_10330 , w_10331 , w_10332 , w_10333 , w_10334 , w_10335 , 
		w_10336 , w_10337 , w_10338 , w_10339 , w_10340 , w_10341 , w_10342 , w_10343 , w_10344 , w_10345 , 
		w_10346 , w_10347 , w_10348 , w_10349 , w_10350 , w_10351 , w_10352 , w_10353 , w_10354 , w_10355 , 
		w_10356 , w_10357 , w_10358 , w_10359 , w_10360 , w_10361 , w_10362 , w_10363 , w_10364 , w_10365 , 
		w_10366 , w_10367 , w_10368 , w_10369 , w_10370 , w_10371 , w_10372 , w_10373 , w_10374 , w_10375 , 
		w_10376 , w_10377 , w_10378 , w_10379 , w_10380 , w_10381 , w_10382 , w_10383 , w_10384 , w_10385 , 
		w_10386 , w_10387 , w_10388 , w_10389 , w_10390 , w_10391 , w_10392 , w_10393 , w_10394 , w_10395 , 
		w_10396 , w_10397 , w_10398 , w_10399 , w_10400 , w_10401 , w_10402 , w_10403 , w_10404 , w_10405 , 
		w_10406 , w_10407 , w_10408 , w_10409 , w_10410 , w_10411 , w_10412 , w_10413 , w_10414 , w_10415 , 
		w_10416 , w_10417 , w_10418 , w_10419 , w_10420 , w_10421 , w_10422 , w_10423 , w_10424 , w_10425 , 
		w_10426 , w_10427 , w_10428 , w_10429 , w_10430 , w_10431 , w_10432 , w_10433 , w_10434 , w_10435 , 
		w_10436 , w_10437 , w_10438 , w_10439 , w_10440 , w_10441 , w_10442 , w_10443 , w_10444 , w_10445 , 
		w_10446 , w_10447 , w_10448 , w_10449 , w_10450 , w_10451 , w_10452 , w_10453 , w_10454 , w_10455 , 
		w_10456 , w_10457 , w_10458 , w_10459 , w_10460 , w_10461 , w_10462 , w_10463 , w_10464 , w_10465 , 
		w_10466 , w_10467 , w_10468 , w_10469 , w_10470 , w_10471 , w_10472 , w_10473 , w_10474 , w_10475 , 
		w_10476 , w_10477 , w_10478 , w_10479 , w_10480 , w_10481 , w_10482 , w_10483 , w_10484 , w_10485 , 
		w_10486 , w_10487 , w_10488 , w_10489 , w_10490 , w_10491 , w_10492 , w_10493 , w_10494 , w_10495 , 
		w_10496 , w_10497 , w_10498 , w_10499 , w_10500 , w_10501 , w_10502 , w_10503 , w_10504 , w_10505 , 
		w_10506 , w_10507 , w_10508 , w_10509 , w_10510 , w_10511 , w_10512 , w_10513 , w_10514 , w_10515 , 
		w_10516 , w_10517 , w_10518 , w_10519 , w_10520 , w_10521 , w_10522 , w_10523 , w_10524 , w_10525 , 
		w_10526 , w_10527 , w_10528 , w_10529 , w_10530 , w_10531 , w_10532 , w_10533 , w_10534 , w_10535 , 
		w_10536 , w_10537 , w_10538 , w_10539 , w_10540 , w_10541 , w_10542 , w_10543 , w_10544 , w_10545 , 
		w_10546 , w_10547 , w_10548 , w_10549 , w_10550 , w_10551 , w_10552 , w_10553 , w_10554 , w_10555 , 
		w_10556 , w_10557 , w_10558 , w_10559 , w_10560 , w_10561 , w_10562 , w_10563 , w_10564 , w_10565 , 
		w_10566 , w_10567 , w_10568 , w_10569 , w_10570 , w_10571 , w_10572 , w_10573 , w_10574 , w_10575 , 
		w_10576 , w_10577 , w_10578 , w_10579 , w_10580 , w_10581 , w_10582 , w_10583 , w_10584 , w_10585 , 
		w_10586 , w_10587 , w_10588 , w_10589 , w_10590 , w_10591 , w_10592 , w_10593 , w_10594 , w_10595 , 
		w_10596 , w_10597 , w_10598 , w_10599 , w_10600 , w_10601 , w_10602 , w_10603 , w_10604 , w_10605 , 
		w_10606 , w_10607 , w_10608 , w_10609 , w_10610 , w_10611 , w_10612 , w_10613 , w_10614 , w_10615 , 
		w_10616 , w_10617 , w_10618 , w_10619 , w_10620 , w_10621 , w_10622 , w_10623 , w_10624 , w_10625 , 
		w_10626 , w_10627 , w_10628 , w_10629 , w_10630 , w_10631 , w_10632 , w_10633 , w_10634 , w_10635 , 
		w_10636 , w_10637 , w_10638 , w_10639 , w_10640 , w_10641 , w_10642 , w_10643 , w_10644 , w_10645 , 
		w_10646 , w_10647 , w_10648 , w_10649 , w_10650 , w_10651 , w_10652 , w_10653 , w_10654 , w_10655 , 
		w_10656 , w_10657 , w_10658 , w_10659 , w_10660 , w_10661 , w_10662 , w_10663 , w_10664 , w_10665 , 
		w_10666 , w_10667 , w_10668 , w_10669 , w_10670 , w_10671 , w_10672 , w_10673 , w_10674 , w_10675 , 
		w_10676 , w_10677 , w_10678 , w_10679 , w_10680 , w_10681 , w_10682 , w_10683 , w_10684 , w_10685 , 
		w_10686 , w_10687 , w_10688 , w_10689 , w_10690 , w_10691 , w_10692 , w_10693 , w_10694 , w_10695 , 
		w_10696 , w_10697 , w_10698 , w_10699 , w_10700 , w_10701 , w_10702 , w_10703 , w_10704 , w_10705 , 
		w_10706 , w_10707 , w_10708 , w_10709 , w_10710 , w_10711 , w_10712 , w_10713 , w_10714 , w_10715 , 
		w_10716 , w_10717 , w_10718 , w_10719 , w_10720 , w_10721 , w_10722 , w_10723 , w_10724 , w_10725 , 
		w_10726 , w_10727 , w_10728 , w_10729 , w_10730 , w_10731 , w_10732 , w_10733 , w_10734 , w_10735 , 
		w_10736 , w_10737 , w_10738 , w_10739 , w_10740 , w_10741 , w_10742 , w_10743 , w_10744 , w_10745 , 
		w_10746 , w_10747 , w_10748 , w_10749 , w_10750 , w_10751 , w_10752 , w_10753 , w_10754 , w_10755 , 
		w_10756 , w_10757 , w_10758 , w_10759 , w_10760 , w_10761 , w_10762 , w_10763 , w_10764 , w_10765 , 
		w_10766 , w_10767 , w_10768 , w_10769 , w_10770 , w_10771 , w_10772 , w_10773 , w_10774 , w_10775 , 
		w_10776 , w_10777 , w_10778 , w_10779 , w_10780 , w_10781 , w_10782 , w_10783 , w_10784 , w_10785 , 
		w_10786 , w_10787 , w_10788 , w_10789 , w_10790 , w_10791 , w_10792 , w_10793 , w_10794 , w_10795 , 
		w_10796 , w_10797 , w_10798 , w_10799 , w_10800 , w_10801 , w_10802 , w_10803 , w_10804 , w_10805 , 
		w_10806 , w_10807 , w_10808 , w_10809 , w_10810 , w_10811 , w_10812 , w_10813 , w_10814 , w_10815 , 
		w_10816 , w_10817 , w_10818 , w_10819 , w_10820 , w_10821 , w_10822 , w_10823 , w_10824 , w_10825 , 
		w_10826 , w_10827 , w_10828 , w_10829 , w_10830 , w_10831 , w_10832 , w_10833 , w_10834 , w_10835 , 
		w_10836 , w_10837 , w_10838 , w_10839 , w_10840 , w_10841 , w_10842 , w_10843 , w_10844 , w_10845 , 
		w_10846 , w_10847 , w_10848 , w_10849 , w_10850 , w_10851 , w_10852 , w_10853 , w_10854 , w_10855 , 
		w_10856 , w_10857 , w_10858 , w_10859 , w_10860 , w_10861 , w_10862 , w_10863 , w_10864 , w_10865 , 
		w_10866 , w_10867 , w_10868 , w_10869 , w_10870 , w_10871 , w_10872 , w_10873 , w_10874 , w_10875 , 
		w_10876 , w_10877 , w_10878 , w_10879 , w_10880 , w_10881 , w_10882 , w_10883 , w_10884 , w_10885 , 
		w_10886 , w_10887 , w_10888 , w_10889 , w_10890 , w_10891 , w_10892 , w_10893 , w_10894 , w_10895 , 
		w_10896 , w_10897 , w_10898 , w_10899 , w_10900 , w_10901 , w_10902 , w_10903 , w_10904 , w_10905 , 
		w_10906 , w_10907 , w_10908 , w_10909 , w_10910 , w_10911 , w_10912 , w_10913 , w_10914 , w_10915 , 
		w_10916 , w_10917 , w_10918 , w_10919 , w_10920 , w_10921 , w_10922 , w_10923 , w_10924 , w_10925 , 
		w_10926 , w_10927 , w_10928 , w_10929 , w_10930 , w_10931 , w_10932 , w_10933 , w_10934 , w_10935 , 
		w_10936 , w_10937 , w_10938 , w_10939 , w_10940 , w_10941 , w_10942 , w_10943 , w_10944 , w_10945 , 
		w_10946 , w_10947 , w_10948 , w_10949 , w_10950 , w_10951 , w_10952 , w_10953 , w_10954 , w_10955 , 
		w_10956 , w_10957 , w_10958 , w_10959 , w_10960 , w_10961 , w_10962 , w_10963 , w_10964 , w_10965 , 
		w_10966 , w_10967 , w_10968 , w_10969 , w_10970 , w_10971 , w_10972 , w_10973 , w_10974 , w_10975 , 
		w_10976 , w_10977 , w_10978 , w_10979 , w_10980 , w_10981 , w_10982 , w_10983 , w_10984 , w_10985 , 
		w_10986 , w_10987 , w_10988 , w_10989 , w_10990 , w_10991 , w_10992 , w_10993 , w_10994 , w_10995 , 
		w_10996 , w_10997 , w_10998 , w_10999 , w_11000 , w_11001 , w_11002 , w_11003 , w_11004 , w_11005 , 
		w_11006 , w_11007 , w_11008 , w_11009 , w_11010 , w_11011 , w_11012 , w_11013 , w_11014 , w_11015 , 
		w_11016 , w_11017 , w_11018 , w_11019 , w_11020 , w_11021 , w_11022 , w_11023 , w_11024 , w_11025 , 
		w_11026 , w_11027 , w_11028 , w_11029 , w_11030 , w_11031 , w_11032 , w_11033 , w_11034 , w_11035 , 
		w_11036 , w_11037 , w_11038 , w_11039 , w_11040 , w_11041 , w_11042 , w_11043 , w_11044 , w_11045 , 
		w_11046 , w_11047 , w_11048 , w_11049 , w_11050 , w_11051 , w_11052 , w_11053 , w_11054 , w_11055 , 
		w_11056 , w_11057 , w_11058 , w_11059 , w_11060 , w_11061 , w_11062 , w_11063 , w_11064 , w_11065 , 
		w_11066 , w_11067 , w_11068 , w_11069 , w_11070 , w_11071 , w_11072 , w_11073 , w_11074 , w_11075 , 
		w_11076 , w_11077 , w_11078 , w_11079 , w_11080 , w_11081 , w_11082 , w_11083 , w_11084 , w_11085 , 
		w_11086 , w_11087 , w_11088 , w_11089 , w_11090 , w_11091 , w_11092 , w_11093 , w_11094 , w_11095 , 
		w_11096 , w_11097 , w_11098 , w_11099 , w_11100 , w_11101 , w_11102 , w_11103 , w_11104 , w_11105 , 
		w_11106 , w_11107 , w_11108 , w_11109 , w_11110 , w_11111 , w_11112 , w_11113 , w_11114 , w_11115 , 
		w_11116 , w_11117 , w_11118 , w_11119 , w_11120 , w_11121 , w_11122 , w_11123 , w_11124 , w_11125 , 
		w_11126 , w_11127 , w_11128 , w_11129 , w_11130 , w_11131 , w_11132 , w_11133 , w_11134 , w_11135 , 
		w_11136 , w_11137 , w_11138 , w_11139 , w_11140 , w_11141 , w_11142 , w_11143 , w_11144 , w_11145 , 
		w_11146 , w_11147 , w_11148 , w_11149 , w_11150 , w_11151 , w_11152 , w_11153 , w_11154 , w_11155 , 
		w_11156 , w_11157 , w_11158 , w_11159 , w_11160 , w_11161 , w_11162 , w_11163 , w_11164 , w_11165 , 
		w_11166 , w_11167 , w_11168 , w_11169 , w_11170 , w_11171 , w_11172 , w_11173 , w_11174 , w_11175 , 
		w_11176 , w_11177 , w_11178 , w_11179 , w_11180 , w_11181 , w_11182 , w_11183 , w_11184 , w_11185 , 
		w_11186 , w_11187 , w_11188 , w_11189 , w_11190 , w_11191 , w_11192 , w_11193 , w_11194 , w_11195 , 
		w_11196 , w_11197 , w_11198 , w_11199 , w_11200 , w_11201 , w_11202 , w_11203 , w_11204 , w_11205 , 
		w_11206 , w_11207 , w_11208 , w_11209 , w_11210 , w_11211 , w_11212 , w_11213 , w_11214 , w_11215 , 
		w_11216 , w_11217 , w_11218 , w_11219 , w_11220 , w_11221 , w_11222 , w_11223 , w_11224 , w_11225 , 
		w_11226 , w_11227 , w_11228 , w_11229 , w_11230 , w_11231 , w_11232 , w_11233 , w_11234 , w_11235 , 
		w_11236 , w_11237 , w_11238 , w_11239 , w_11240 , w_11241 , w_11242 , w_11243 , w_11244 , w_11245 , 
		w_11246 , w_11247 , w_11248 , w_11249 , w_11250 , w_11251 , w_11252 , w_11253 , w_11254 , w_11255 , 
		w_11256 , w_11257 , w_11258 , w_11259 , w_11260 , w_11261 , w_11262 , w_11263 , w_11264 , w_11265 , 
		w_11266 , w_11267 , w_11268 , w_11269 , w_11270 , w_11271 , w_11272 , w_11273 , w_11274 , w_11275 , 
		w_11276 , w_11277 , w_11278 , w_11279 , w_11280 , w_11281 , w_11282 , w_11283 , w_11284 , w_11285 , 
		w_11286 , w_11287 , w_11288 , w_11289 , w_11290 , w_11291 , w_11292 , w_11293 , w_11294 , w_11295 , 
		w_11296 , w_11297 , w_11298 , w_11299 , w_11300 , w_11301 , w_11302 , w_11303 , w_11304 , w_11305 , 
		w_11306 , w_11307 , w_11308 , w_11309 , w_11310 , w_11311 , w_11312 , w_11313 , w_11314 , w_11315 , 
		w_11316 , w_11317 , w_11318 , w_11319 , w_11320 , w_11321 , w_11322 , w_11323 , w_11324 , w_11325 , 
		w_11326 , w_11327 , w_11328 , w_11329 , w_11330 , w_11331 , w_11332 , w_11333 , w_11334 , w_11335 , 
		w_11336 , w_11337 , w_11338 , w_11339 , w_11340 , w_11341 , w_11342 , w_11343 , w_11344 , w_11345 , 
		w_11346 , w_11347 , w_11348 , w_11349 , w_11350 , w_11351 , w_11352 , w_11353 , w_11354 , w_11355 , 
		w_11356 , w_11357 , w_11358 , w_11359 , w_11360 , w_11361 , w_11362 , w_11363 , w_11364 , w_11365 , 
		w_11366 , w_11367 , w_11368 , w_11369 , w_11370 , w_11371 , w_11372 , w_11373 , w_11374 , w_11375 , 
		w_11376 , w_11377 , w_11378 , w_11379 , w_11380 , w_11381 , w_11382 , w_11383 , w_11384 , w_11385 , 
		w_11386 , w_11387 , w_11388 , w_11389 , w_11390 , w_11391 , w_11392 , w_11393 , w_11394 , w_11395 , 
		w_11396 , w_11397 , w_11398 , w_11399 , w_11400 , w_11401 , w_11402 , w_11403 , w_11404 , w_11405 , 
		w_11406 , w_11407 , w_11408 , w_11409 , w_11410 , w_11411 , w_11412 , w_11413 , w_11414 , w_11415 , 
		w_11416 , w_11417 , w_11418 , w_11419 , w_11420 , w_11421 , w_11422 , w_11423 , w_11424 , w_11425 , 
		w_11426 , w_11427 , w_11428 , w_11429 , w_11430 , w_11431 , w_11432 , w_11433 , w_11434 , w_11435 , 
		w_11436 , w_11437 , w_11438 , w_11439 , w_11440 , w_11441 , w_11442 , w_11443 , w_11444 , w_11445 , 
		w_11446 , w_11447 , w_11448 , w_11449 , w_11450 , w_11451 , w_11452 , w_11453 , w_11454 , w_11455 , 
		w_11456 , w_11457 , w_11458 , w_11459 , w_11460 , w_11461 , w_11462 , w_11463 , w_11464 , w_11465 , 
		w_11466 , w_11467 , w_11468 , w_11469 , w_11470 , w_11471 , w_11472 , w_11473 , w_11474 , w_11475 , 
		w_11476 , w_11477 , w_11478 , w_11479 , w_11480 , w_11481 , w_11482 , w_11483 , w_11484 , w_11485 , 
		w_11486 , w_11487 , w_11488 , w_11489 , w_11490 , w_11491 , w_11492 , w_11493 , w_11494 , w_11495 , 
		w_11496 , w_11497 , w_11498 , w_11499 , w_11500 , w_11501 , w_11502 , w_11503 , w_11504 , w_11505 , 
		w_11506 , w_11507 , w_11508 , w_11509 , w_11510 , w_11511 , w_11512 , w_11513 , w_11514 , w_11515 , 
		w_11516 , w_11517 , w_11518 , w_11519 , w_11520 , w_11521 , w_11522 , w_11523 , w_11524 , w_11525 , 
		w_11526 , w_11527 , w_11528 , w_11529 , w_11530 , w_11531 , w_11532 , w_11533 , w_11534 , w_11535 , 
		w_11536 , w_11537 , w_11538 , w_11539 , w_11540 , w_11541 , w_11542 , w_11543 , w_11544 , w_11545 , 
		w_11546 , w_11547 , w_11548 , w_11549 , w_11550 , w_11551 , w_11552 , w_11553 , w_11554 , w_11555 , 
		w_11556 , w_11557 , w_11558 , w_11559 , w_11560 , w_11561 , w_11562 , w_11563 , w_11564 , w_11565 , 
		w_11566 , w_11567 , w_11568 , w_11569 , w_11570 , w_11571 , w_11572 , w_11573 , w_11574 , w_11575 , 
		w_11576 , w_11577 , w_11578 , w_11579 , w_11580 , w_11581 , w_11582 , w_11583 , w_11584 , w_11585 , 
		w_11586 , w_11587 , w_11588 , w_11589 , w_11590 , w_11591 , w_11592 , w_11593 , w_11594 , w_11595 , 
		w_11596 , w_11597 , w_11598 , w_11599 , w_11600 , w_11601 , w_11602 , w_11603 , w_11604 , w_11605 , 
		w_11606 , w_11607 , w_11608 , w_11609 , w_11610 , w_11611 , w_11612 , w_11613 , w_11614 , w_11615 , 
		w_11616 , w_11617 , w_11618 , w_11619 , w_11620 , w_11621 , w_11622 , w_11623 , w_11624 , w_11625 , 
		w_11626 , w_11627 , w_11628 , w_11629 , w_11630 , w_11631 , w_11632 , w_11633 , w_11634 , w_11635 , 
		w_11636 , w_11637 , w_11638 , w_11639 , w_11640 , w_11641 , w_11642 , w_11643 , w_11644 , w_11645 , 
		w_11646 , w_11647 , w_11648 , w_11649 , w_11650 , w_11651 , w_11652 , w_11653 , w_11654 , w_11655 , 
		w_11656 , w_11657 , w_11658 , w_11659 , w_11660 , w_11661 , w_11662 , w_11663 , w_11664 , w_11665 , 
		w_11666 , w_11667 , w_11668 , w_11669 , w_11670 , w_11671 , w_11672 , w_11673 , w_11674 , w_11675 , 
		w_11676 , w_11677 , w_11678 , w_11679 , w_11680 , w_11681 , w_11682 , w_11683 , w_11684 , w_11685 , 
		w_11686 , w_11687 , w_11688 , w_11689 , w_11690 , w_11691 , w_11692 , w_11693 , w_11694 , w_11695 , 
		w_11696 , w_11697 , w_11698 , w_11699 , w_11700 , w_11701 , w_11702 , w_11703 , w_11704 , w_11705 , 
		w_11706 , w_11707 , w_11708 , w_11709 , w_11710 , w_11711 , w_11712 , w_11713 , w_11714 , w_11715 , 
		w_11716 , w_11717 , w_11718 , w_11719 , w_11720 , w_11721 , w_11722 , w_11723 , w_11724 , w_11725 , 
		w_11726 , w_11727 , w_11728 , w_11729 , w_11730 , w_11731 , w_11732 , w_11733 , w_11734 , w_11735 , 
		w_11736 , w_11737 , w_11738 , w_11739 , w_11740 , w_11741 , w_11742 , w_11743 , w_11744 , w_11745 , 
		w_11746 , w_11747 , w_11748 , w_11749 , w_11750 , w_11751 , w_11752 , w_11753 , w_11754 , w_11755 , 
		w_11756 , w_11757 , w_11758 , w_11759 , w_11760 , w_11761 , w_11762 , w_11763 , w_11764 , w_11765 , 
		w_11766 , w_11767 , w_11768 , w_11769 , w_11770 , w_11771 , w_11772 , w_11773 , w_11774 , w_11775 , 
		w_11776 , w_11777 , w_11778 , w_11779 , w_11780 , w_11781 , w_11782 , w_11783 , w_11784 , w_11785 , 
		w_11786 , w_11787 , w_11788 , w_11789 , w_11790 , w_11791 , w_11792 , w_11793 , w_11794 , w_11795 , 
		w_11796 , w_11797 , w_11798 , w_11799 , w_11800 , w_11801 , w_11802 , w_11803 , w_11804 , w_11805 , 
		w_11806 , w_11807 , w_11808 , w_11809 , w_11810 , w_11811 , w_11812 , w_11813 , w_11814 , w_11815 , 
		w_11816 , w_11817 , w_11818 , w_11819 , w_11820 , w_11821 , w_11822 , w_11823 , w_11824 , w_11825 , 
		w_11826 , w_11827 , w_11828 , w_11829 , w_11830 , w_11831 , w_11832 , w_11833 , w_11834 , w_11835 , 
		w_11836 , w_11837 , w_11838 , w_11839 , w_11840 , w_11841 , w_11842 , w_11843 , w_11844 , w_11845 , 
		w_11846 , w_11847 , w_11848 , w_11849 , w_11850 , w_11851 , w_11852 , w_11853 , w_11854 , w_11855 , 
		w_11856 , w_11857 , w_11858 , w_11859 , w_11860 , w_11861 , w_11862 , w_11863 , w_11864 , w_11865 , 
		w_11866 , w_11867 , w_11868 , w_11869 , w_11870 , w_11871 , w_11872 , w_11873 , w_11874 , w_11875 , 
		w_11876 , w_11877 , w_11878 , w_11879 , w_11880 , w_11881 , w_11882 , w_11883 , w_11884 , w_11885 , 
		w_11886 , w_11887 , w_11888 , w_11889 , w_11890 , w_11891 , w_11892 , w_11893 , w_11894 , w_11895 , 
		w_11896 , w_11897 , w_11898 , w_11899 , w_11900 , w_11901 , w_11902 , w_11903 , w_11904 , w_11905 , 
		w_11906 , w_11907 , w_11908 , w_11909 , w_11910 , w_11911 , w_11912 , w_11913 , w_11914 , w_11915 , 
		w_11916 , w_11917 , w_11918 , w_11919 , w_11920 , w_11921 , w_11922 , w_11923 , w_11924 , w_11925 , 
		w_11926 , w_11927 , w_11928 , w_11929 , w_11930 , w_11931 , w_11932 , w_11933 , w_11934 , w_11935 , 
		w_11936 , w_11937 , w_11938 , w_11939 , w_11940 , w_11941 , w_11942 , w_11943 , w_11944 , w_11945 , 
		w_11946 , w_11947 , w_11948 , w_11949 , w_11950 , w_11951 , w_11952 , w_11953 , w_11954 , w_11955 , 
		w_11956 , w_11957 , w_11958 , w_11959 , w_11960 , w_11961 , w_11962 , w_11963 , w_11964 , w_11965 , 
		w_11966 , w_11967 , w_11968 , w_11969 , w_11970 , w_11971 , w_11972 , w_11973 , w_11974 , w_11975 , 
		w_11976 , w_11977 , w_11978 , w_11979 , w_11980 , w_11981 , w_11982 , w_11983 , w_11984 , w_11985 , 
		w_11986 , w_11987 , w_11988 , w_11989 , w_11990 , w_11991 , w_11992 , w_11993 , w_11994 , w_11995 , 
		w_11996 , w_11997 , w_11998 , w_11999 , w_12000 , w_12001 , w_12002 , w_12003 , w_12004 , w_12005 , 
		w_12006 , w_12007 , w_12008 , w_12009 , w_12010 , w_12011 , w_12012 , w_12013 , w_12014 , w_12015 , 
		w_12016 , w_12017 , w_12018 , w_12019 , w_12020 , w_12021 , w_12022 , w_12023 , w_12024 , w_12025 , 
		w_12026 , w_12027 , w_12028 , w_12029 , w_12030 , w_12031 , w_12032 , w_12033 , w_12034 , w_12035 , 
		w_12036 , w_12037 , w_12038 , w_12039 , w_12040 , w_12041 , w_12042 , w_12043 , w_12044 , w_12045 , 
		w_12046 , w_12047 , w_12048 , w_12049 , w_12050 , w_12051 , w_12052 , w_12053 , w_12054 , w_12055 , 
		w_12056 , w_12057 , w_12058 , w_12059 , w_12060 , w_12061 , w_12062 , w_12063 , w_12064 , w_12065 , 
		w_12066 , w_12067 , w_12068 , w_12069 , w_12070 , w_12071 , w_12072 , w_12073 , w_12074 , w_12075 , 
		w_12076 , w_12077 , w_12078 , w_12079 , w_12080 , w_12081 , w_12082 , w_12083 , w_12084 , w_12085 , 
		w_12086 , w_12087 , w_12088 , w_12089 , w_12090 , w_12091 , w_12092 , w_12093 , w_12094 , w_12095 , 
		w_12096 , w_12097 , w_12098 , w_12099 , w_12100 , w_12101 , w_12102 , w_12103 , w_12104 , w_12105 , 
		w_12106 , w_12107 , w_12108 , w_12109 , w_12110 , w_12111 , w_12112 , w_12113 , w_12114 , w_12115 , 
		w_12116 , w_12117 , w_12118 , w_12119 , w_12120 , w_12121 , w_12122 , w_12123 , w_12124 , w_12125 , 
		w_12126 , w_12127 , w_12128 , w_12129 , w_12130 , w_12131 , w_12132 , w_12133 , w_12134 , w_12135 , 
		w_12136 , w_12137 , w_12138 , w_12139 , w_12140 , w_12141 , w_12142 , w_12143 , w_12144 , w_12145 , 
		w_12146 , w_12147 , w_12148 , w_12149 , w_12150 , w_12151 , w_12152 , w_12153 , w_12154 , w_12155 , 
		w_12156 , w_12157 , w_12158 , w_12159 , w_12160 , w_12161 , w_12162 , w_12163 , w_12164 , w_12165 , 
		w_12166 , w_12167 , w_12168 , w_12169 , w_12170 , w_12171 , w_12172 , w_12173 , w_12174 , w_12175 , 
		w_12176 , w_12177 , w_12178 , w_12179 , w_12180 , w_12181 , w_12182 , w_12183 , w_12184 , w_12185 , 
		w_12186 , w_12187 , w_12188 , w_12189 , w_12190 , w_12191 , w_12192 , w_12193 , w_12194 , w_12195 , 
		w_12196 , w_12197 , w_12198 , w_12199 , w_12200 , w_12201 , w_12202 , w_12203 , w_12204 , w_12205 , 
		w_12206 , w_12207 , w_12208 , w_12209 , w_12210 , w_12211 , w_12212 , w_12213 , w_12214 , w_12215 , 
		w_12216 , w_12217 , w_12218 , w_12219 , w_12220 , w_12221 , w_12222 , w_12223 , w_12224 , w_12225 , 
		w_12226 , w_12227 , w_12228 , w_12229 , w_12230 , w_12231 , w_12232 , w_12233 , w_12234 , w_12235 , 
		w_12236 , w_12237 , w_12238 , w_12239 , w_12240 , w_12241 , w_12242 , w_12243 , w_12244 , w_12245 , 
		w_12246 , w_12247 , w_12248 , w_12249 , w_12250 , w_12251 , w_12252 , w_12253 , w_12254 , w_12255 , 
		w_12256 , w_12257 , w_12258 , w_12259 , w_12260 , w_12261 , w_12262 , w_12263 , w_12264 , w_12265 , 
		w_12266 , w_12267 , w_12268 , w_12269 , w_12270 , w_12271 , w_12272 , w_12273 , w_12274 , w_12275 , 
		w_12276 , w_12277 , w_12278 , w_12279 , w_12280 , w_12281 , w_12282 , w_12283 , w_12284 , w_12285 , 
		w_12286 , w_12287 , w_12288 , w_12289 , w_12290 , w_12291 , w_12292 , w_12293 , w_12294 , w_12295 , 
		w_12296 , w_12297 , w_12298 , w_12299 , w_12300 , w_12301 , w_12302 , w_12303 , w_12304 , w_12305 , 
		w_12306 , w_12307 , w_12308 , w_12309 , w_12310 , w_12311 , w_12312 , w_12313 , w_12314 , w_12315 , 
		w_12316 , w_12317 , w_12318 , w_12319 , w_12320 , w_12321 , w_12322 , w_12323 , w_12324 , w_12325 , 
		w_12326 , w_12327 , w_12328 , w_12329 , w_12330 , w_12331 , w_12332 , w_12333 , w_12334 , w_12335 , 
		w_12336 , w_12337 , w_12338 , w_12339 , w_12340 , w_12341 , w_12342 , w_12343 , w_12344 , w_12345 , 
		w_12346 , w_12347 , w_12348 , w_12349 , w_12350 , w_12351 , w_12352 , w_12353 , w_12354 , w_12355 , 
		w_12356 , w_12357 , w_12358 , w_12359 , w_12360 , w_12361 , w_12362 , w_12363 , w_12364 , w_12365 , 
		w_12366 , w_12367 , w_12368 , w_12369 , w_12370 , w_12371 , w_12372 , w_12373 , w_12374 , w_12375 , 
		w_12376 , w_12377 , w_12378 , w_12379 , w_12380 , w_12381 , w_12382 , w_12383 , w_12384 , w_12385 , 
		w_12386 , w_12387 , w_12388 , w_12389 , w_12390 , w_12391 , w_12392 , w_12393 , w_12394 , w_12395 , 
		w_12396 , w_12397 , w_12398 , w_12399 , w_12400 , w_12401 , w_12402 , w_12403 , w_12404 , w_12405 , 
		w_12406 , w_12407 , w_12408 , w_12409 , w_12410 , w_12411 , w_12412 , w_12413 , w_12414 , w_12415 , 
		w_12416 , w_12417 , w_12418 , w_12419 , w_12420 , w_12421 , w_12422 , w_12423 , w_12424 , w_12425 , 
		w_12426 , w_12427 , w_12428 , w_12429 , w_12430 , w_12431 , w_12432 , w_12433 , w_12434 , w_12435 , 
		w_12436 , w_12437 , w_12438 , w_12439 , w_12440 , w_12441 , w_12442 , w_12443 , w_12444 , w_12445 , 
		w_12446 , w_12447 , w_12448 , w_12449 , w_12450 , w_12451 , w_12452 , w_12453 , w_12454 , w_12455 , 
		w_12456 , w_12457 , w_12458 , w_12459 , w_12460 , w_12461 , w_12462 , w_12463 , w_12464 , w_12465 , 
		w_12466 , w_12467 , w_12468 , w_12469 , w_12470 , w_12471 , w_12472 , w_12473 , w_12474 , w_12475 , 
		w_12476 , w_12477 , w_12478 , w_12479 , w_12480 , w_12481 , w_12482 , w_12483 , w_12484 , w_12485 , 
		w_12486 , w_12487 , w_12488 , w_12489 , w_12490 , w_12491 , w_12492 , w_12493 , w_12494 , w_12495 , 
		w_12496 , w_12497 , w_12498 , w_12499 , w_12500 , w_12501 , w_12502 , w_12503 , w_12504 , w_12505 , 
		w_12506 , w_12507 , w_12508 , w_12509 , w_12510 , w_12511 , w_12512 , w_12513 , w_12514 , w_12515 , 
		w_12516 , w_12517 , w_12518 , w_12519 , w_12520 , w_12521 , w_12522 , w_12523 , w_12524 , w_12525 , 
		w_12526 , w_12527 , w_12528 , w_12529 , w_12530 , w_12531 , w_12532 , w_12533 , w_12534 , w_12535 , 
		w_12536 , w_12537 , w_12538 , w_12539 , w_12540 , w_12541 , w_12542 , w_12543 , w_12544 , w_12545 , 
		w_12546 , w_12547 , w_12548 , w_12549 , w_12550 , w_12551 , w_12552 , w_12553 , w_12554 , w_12555 , 
		w_12556 , w_12557 , w_12558 , w_12559 , w_12560 , w_12561 , w_12562 , w_12563 , w_12564 , w_12565 , 
		w_12566 , w_12567 , w_12568 , w_12569 , w_12570 , w_12571 , w_12572 , w_12573 , w_12574 , w_12575 , 
		w_12576 , w_12577 , w_12578 , w_12579 , w_12580 , w_12581 , w_12582 , w_12583 , w_12584 , w_12585 , 
		w_12586 , w_12587 , w_12588 , w_12589 , w_12590 , w_12591 , w_12592 , w_12593 , w_12594 , w_12595 , 
		w_12596 , w_12597 , w_12598 , w_12599 , w_12600 , w_12601 , w_12602 , w_12603 , w_12604 , w_12605 , 
		w_12606 , w_12607 , w_12608 , w_12609 , w_12610 , w_12611 , w_12612 , w_12613 , w_12614 , w_12615 , 
		w_12616 , w_12617 , w_12618 , w_12619 , w_12620 , w_12621 , w_12622 , w_12623 , w_12624 , w_12625 , 
		w_12626 , w_12627 , w_12628 , w_12629 , w_12630 , w_12631 , w_12632 , w_12633 , w_12634 , w_12635 , 
		w_12636 , w_12637 , w_12638 , w_12639 , w_12640 , w_12641 , w_12642 , w_12643 , w_12644 , w_12645 , 
		w_12646 , w_12647 , w_12648 , w_12649 , w_12650 , w_12651 , w_12652 , w_12653 , w_12654 , w_12655 , 
		w_12656 , w_12657 , w_12658 , w_12659 , w_12660 , w_12661 , w_12662 , w_12663 , w_12664 , w_12665 , 
		w_12666 , w_12667 , w_12668 , w_12669 , w_12670 , w_12671 , w_12672 , w_12673 , w_12674 , w_12675 , 
		w_12676 , w_12677 , w_12678 , w_12679 , w_12680 , w_12681 , w_12682 , w_12683 , w_12684 , w_12685 , 
		w_12686 , w_12687 , w_12688 , w_12689 , w_12690 , w_12691 , w_12692 , w_12693 , w_12694 , w_12695 , 
		w_12696 , w_12697 , w_12698 , w_12699 , w_12700 , w_12701 , w_12702 , w_12703 , w_12704 , w_12705 , 
		w_12706 , w_12707 , w_12708 , w_12709 , w_12710 , w_12711 , w_12712 , w_12713 , w_12714 , w_12715 , 
		w_12716 , w_12717 , w_12718 , w_12719 , w_12720 , w_12721 , w_12722 , w_12723 , w_12724 , w_12725 , 
		w_12726 , w_12727 , w_12728 , w_12729 , w_12730 , w_12731 , w_12732 , w_12733 , w_12734 , w_12735 , 
		w_12736 , w_12737 , w_12738 , w_12739 , w_12740 , w_12741 , w_12742 , w_12743 , w_12744 , w_12745 , 
		w_12746 , w_12747 , w_12748 , w_12749 , w_12750 , w_12751 , w_12752 , w_12753 , w_12754 , w_12755 , 
		w_12756 , w_12757 , w_12758 , w_12759 , w_12760 , w_12761 , w_12762 , w_12763 , w_12764 , w_12765 , 
		w_12766 , w_12767 , w_12768 , w_12769 , w_12770 , w_12771 , w_12772 , w_12773 , w_12774 , w_12775 , 
		w_12776 , w_12777 , w_12778 , w_12779 , w_12780 , w_12781 , w_12782 , w_12783 , w_12784 , w_12785 , 
		w_12786 , w_12787 , w_12788 , w_12789 , w_12790 , w_12791 , w_12792 , w_12793 , w_12794 , w_12795 , 
		w_12796 , w_12797 , w_12798 , w_12799 , w_12800 , w_12801 , w_12802 , w_12803 , w_12804 , w_12805 , 
		w_12806 , w_12807 , w_12808 , w_12809 , w_12810 , w_12811 , w_12812 , w_12813 , w_12814 , w_12815 , 
		w_12816 , w_12817 , w_12818 , w_12819 , w_12820 , w_12821 , w_12822 , w_12823 , w_12824 , w_12825 , 
		w_12826 , w_12827 , w_12828 , w_12829 , w_12830 , w_12831 , w_12832 , w_12833 , w_12834 , w_12835 , 
		w_12836 , w_12837 , w_12838 , w_12839 , w_12840 , w_12841 , w_12842 , w_12843 , w_12844 , w_12845 , 
		w_12846 , w_12847 , w_12848 , w_12849 , w_12850 , w_12851 , w_12852 , w_12853 , w_12854 , w_12855 , 
		w_12856 , w_12857 , w_12858 , w_12859 , w_12860 , w_12861 , w_12862 , w_12863 , w_12864 , w_12865 , 
		w_12866 , w_12867 , w_12868 , w_12869 , w_12870 , w_12871 , w_12872 , w_12873 , w_12874 , w_12875 , 
		w_12876 , w_12877 , w_12878 , w_12879 , w_12880 , w_12881 , w_12882 , w_12883 , w_12884 , w_12885 , 
		w_12886 , w_12887 , w_12888 , w_12889 , w_12890 , w_12891 , w_12892 , w_12893 , w_12894 , w_12895 , 
		w_12896 , w_12897 , w_12898 , w_12899 , w_12900 , w_12901 , w_12902 , w_12903 , w_12904 , w_12905 , 
		w_12906 , w_12907 , w_12908 , w_12909 , w_12910 , w_12911 , w_12912 , w_12913 , w_12914 , w_12915 , 
		w_12916 , w_12917 , w_12918 , w_12919 , w_12920 , w_12921 , w_12922 , w_12923 , w_12924 , w_12925 , 
		w_12926 , w_12927 , w_12928 , w_12929 , w_12930 , w_12931 , w_12932 , w_12933 , w_12934 , w_12935 , 
		w_12936 , w_12937 , w_12938 , w_12939 , w_12940 , w_12941 , w_12942 , w_12943 , w_12944 , w_12945 , 
		w_12946 , w_12947 , w_12948 , w_12949 , w_12950 , w_12951 , w_12952 , w_12953 , w_12954 , w_12955 , 
		w_12956 , w_12957 , w_12958 , w_12959 , w_12960 , w_12961 , w_12962 , w_12963 , w_12964 , w_12965 , 
		w_12966 , w_12967 , w_12968 , w_12969 , w_12970 , w_12971 , w_12972 , w_12973 , w_12974 , w_12975 , 
		w_12976 , w_12977 , w_12978 , w_12979 , w_12980 , w_12981 , w_12982 , w_12983 , w_12984 , w_12985 , 
		w_12986 , w_12987 , w_12988 , w_12989 , w_12990 , w_12991 , w_12992 , w_12993 , w_12994 , w_12995 , 
		w_12996 , w_12997 , w_12998 , w_12999 , w_13000 , w_13001 , w_13002 , w_13003 , w_13004 , w_13005 , 
		w_13006 , w_13007 , w_13008 , w_13009 , w_13010 , w_13011 , w_13012 , w_13013 , w_13014 , w_13015 , 
		w_13016 , w_13017 , w_13018 , w_13019 , w_13020 , w_13021 , w_13022 , w_13023 , w_13024 , w_13025 , 
		w_13026 , w_13027 , w_13028 , w_13029 , w_13030 , w_13031 , w_13032 , w_13033 , w_13034 , w_13035 , 
		w_13036 , w_13037 , w_13038 , w_13039 , w_13040 , w_13041 , w_13042 , w_13043 , w_13044 , w_13045 , 
		w_13046 , w_13047 , w_13048 , w_13049 , w_13050 , w_13051 , w_13052 , w_13053 , w_13054 , w_13055 , 
		w_13056 , w_13057 , w_13058 , w_13059 , w_13060 , w_13061 , w_13062 , w_13063 , w_13064 , w_13065 , 
		w_13066 , w_13067 , w_13068 , w_13069 , w_13070 , w_13071 , w_13072 , w_13073 , w_13074 , w_13075 , 
		w_13076 , w_13077 , w_13078 , w_13079 , w_13080 , w_13081 , w_13082 , w_13083 , w_13084 , w_13085 , 
		w_13086 , w_13087 , w_13088 , w_13089 , w_13090 , w_13091 , w_13092 , w_13093 , w_13094 , w_13095 , 
		w_13096 , w_13097 , w_13098 , w_13099 , w_13100 , w_13101 , w_13102 , w_13103 , w_13104 , w_13105 , 
		w_13106 , w_13107 , w_13108 , w_13109 , w_13110 , w_13111 , w_13112 , w_13113 , w_13114 , w_13115 , 
		w_13116 , w_13117 , w_13118 , w_13119 , w_13120 , w_13121 , w_13122 , w_13123 , w_13124 , w_13125 , 
		w_13126 , w_13127 , w_13128 , w_13129 , w_13130 , w_13131 , w_13132 , w_13133 , w_13134 , w_13135 , 
		w_13136 , w_13137 , w_13138 , w_13139 , w_13140 , w_13141 , w_13142 , w_13143 , w_13144 , w_13145 , 
		w_13146 , w_13147 , w_13148 , w_13149 , w_13150 , w_13151 , w_13152 , w_13153 , w_13154 , w_13155 , 
		w_13156 , w_13157 , w_13158 , w_13159 , w_13160 , w_13161 , w_13162 , w_13163 , w_13164 , w_13165 , 
		w_13166 , w_13167 , w_13168 , w_13169 , w_13170 , w_13171 , w_13172 , w_13173 , w_13174 , w_13175 , 
		w_13176 , w_13177 , w_13178 , w_13179 , w_13180 , w_13181 , w_13182 , w_13183 , w_13184 , w_13185 , 
		w_13186 , w_13187 , w_13188 , w_13189 , w_13190 , w_13191 , w_13192 , w_13193 , w_13194 , w_13195 , 
		w_13196 , w_13197 , w_13198 , w_13199 , w_13200 , w_13201 , w_13202 , w_13203 , w_13204 , w_13205 , 
		w_13206 , w_13207 , w_13208 , w_13209 , w_13210 , w_13211 , w_13212 , w_13213 , w_13214 , w_13215 , 
		w_13216 , w_13217 , w_13218 , w_13219 , w_13220 , w_13221 , w_13222 , w_13223 , w_13224 , w_13225 , 
		w_13226 , w_13227 , w_13228 , w_13229 , w_13230 , w_13231 , w_13232 , w_13233 , w_13234 , w_13235 , 
		w_13236 , w_13237 , w_13238 , w_13239 , w_13240 , w_13241 , w_13242 , w_13243 , w_13244 , w_13245 , 
		w_13246 , w_13247 , w_13248 , w_13249 , w_13250 , w_13251 , w_13252 , w_13253 , w_13254 , w_13255 , 
		w_13256 , w_13257 , w_13258 , w_13259 , w_13260 , w_13261 , w_13262 , w_13263 , w_13264 , w_13265 , 
		w_13266 , w_13267 , w_13268 , w_13269 , w_13270 , w_13271 , w_13272 , w_13273 , w_13274 , w_13275 , 
		w_13276 , w_13277 , w_13278 , w_13279 , w_13280 , w_13281 , w_13282 , w_13283 , w_13284 , w_13285 , 
		w_13286 , w_13287 , w_13288 , w_13289 , w_13290 , w_13291 , w_13292 , w_13293 , w_13294 , w_13295 , 
		w_13296 , w_13297 , w_13298 , w_13299 , w_13300 , w_13301 , w_13302 , w_13303 , w_13304 , w_13305 , 
		w_13306 , w_13307 , w_13308 , w_13309 , w_13310 , w_13311 , w_13312 , w_13313 , w_13314 , w_13315 , 
		w_13316 , w_13317 , w_13318 , w_13319 , w_13320 , w_13321 , w_13322 , w_13323 , w_13324 , w_13325 , 
		w_13326 , w_13327 , w_13328 , w_13329 , w_13330 , w_13331 , w_13332 , w_13333 , w_13334 , w_13335 , 
		w_13336 , w_13337 , w_13338 , w_13339 , w_13340 , w_13341 , w_13342 , w_13343 , w_13344 , w_13345 , 
		w_13346 , w_13347 , w_13348 , w_13349 , w_13350 , w_13351 , w_13352 , w_13353 , w_13354 , w_13355 , 
		w_13356 , w_13357 , w_13358 , w_13359 , w_13360 , w_13361 , w_13362 , w_13363 , w_13364 , w_13365 , 
		w_13366 , w_13367 , w_13368 , w_13369 , w_13370 , w_13371 , w_13372 , w_13373 , w_13374 , w_13375 , 
		w_13376 , w_13377 , w_13378 , w_13379 , w_13380 , w_13381 , w_13382 , w_13383 , w_13384 , w_13385 , 
		w_13386 , w_13387 , w_13388 , w_13389 , w_13390 , w_13391 , w_13392 , w_13393 , w_13394 , w_13395 , 
		w_13396 , w_13397 , w_13398 , w_13399 , w_13400 , w_13401 , w_13402 , w_13403 , w_13404 , w_13405 , 
		w_13406 , w_13407 , w_13408 , w_13409 , w_13410 , w_13411 , w_13412 , w_13413 , w_13414 , w_13415 , 
		w_13416 , w_13417 , w_13418 , w_13419 , w_13420 , w_13421 , w_13422 , w_13423 , w_13424 , w_13425 , 
		w_13426 , w_13427 , w_13428 , w_13429 , w_13430 , w_13431 , w_13432 , w_13433 , w_13434 , w_13435 , 
		w_13436 , w_13437 , w_13438 , w_13439 , w_13440 , w_13441 , w_13442 , w_13443 , w_13444 , w_13445 , 
		w_13446 , w_13447 , w_13448 , w_13449 , w_13450 , w_13451 , w_13452 , w_13453 , w_13454 , w_13455 , 
		w_13456 , w_13457 , w_13458 , w_13459 , w_13460 , w_13461 , w_13462 , w_13463 , w_13464 , w_13465 , 
		w_13466 , w_13467 , w_13468 , w_13469 , w_13470 , w_13471 , w_13472 , w_13473 , w_13474 , w_13475 , 
		w_13476 , w_13477 , w_13478 , w_13479 , w_13480 , w_13481 , w_13482 , w_13483 , w_13484 , w_13485 , 
		w_13486 , w_13487 , w_13488 , w_13489 , w_13490 , w_13491 , w_13492 , w_13493 , w_13494 , w_13495 , 
		w_13496 , w_13497 , w_13498 , w_13499 , w_13500 , w_13501 , w_13502 , w_13503 , w_13504 , w_13505 , 
		w_13506 , w_13507 , w_13508 , w_13509 , w_13510 , w_13511 , w_13512 , w_13513 , w_13514 , w_13515 , 
		w_13516 , w_13517 , w_13518 , w_13519 , w_13520 , w_13521 , w_13522 , w_13523 , w_13524 , w_13525 , 
		w_13526 , w_13527 , w_13528 , w_13529 , w_13530 , w_13531 , w_13532 , w_13533 , w_13534 , w_13535 , 
		w_13536 , w_13537 , w_13538 , w_13539 , w_13540 , w_13541 , w_13542 , w_13543 , w_13544 , w_13545 , 
		w_13546 , w_13547 , w_13548 , w_13549 , w_13550 , w_13551 , w_13552 , w_13553 , w_13554 , w_13555 , 
		w_13556 , w_13557 , w_13558 , w_13559 , w_13560 , w_13561 , w_13562 , w_13563 , w_13564 , w_13565 , 
		w_13566 , w_13567 , w_13568 , w_13569 , w_13570 , w_13571 , w_13572 , w_13573 , w_13574 , w_13575 , 
		w_13576 , w_13577 , w_13578 , w_13579 , w_13580 , w_13581 , w_13582 , w_13583 , w_13584 , w_13585 , 
		w_13586 , w_13587 , w_13588 , w_13589 , w_13590 , w_13591 , w_13592 , w_13593 , w_13594 , w_13595 , 
		w_13596 , w_13597 , w_13598 , w_13599 , w_13600 , w_13601 , w_13602 , w_13603 , w_13604 , w_13605 , 
		w_13606 , w_13607 , w_13608 , w_13609 , w_13610 , w_13611 , w_13612 , w_13613 , w_13614 , w_13615 , 
		w_13616 , w_13617 , w_13618 , w_13619 , w_13620 , w_13621 , w_13622 , w_13623 , w_13624 , w_13625 , 
		w_13626 , w_13627 , w_13628 , w_13629 , w_13630 , w_13631 , w_13632 , w_13633 , w_13634 , w_13635 , 
		w_13636 , w_13637 , w_13638 , w_13639 , w_13640 , w_13641 , w_13642 , w_13643 , w_13644 , w_13645 , 
		w_13646 , w_13647 , w_13648 , w_13649 , w_13650 , w_13651 , w_13652 , w_13653 , w_13654 , w_13655 , 
		w_13656 , w_13657 , w_13658 , w_13659 , w_13660 , w_13661 , w_13662 , w_13663 , w_13664 , w_13665 , 
		w_13666 , w_13667 , w_13668 , w_13669 , w_13670 , w_13671 , w_13672 , w_13673 , w_13674 , w_13675 , 
		w_13676 , w_13677 , w_13678 , w_13679 , w_13680 , w_13681 , w_13682 , w_13683 , w_13684 , w_13685 , 
		w_13686 , w_13687 , w_13688 , w_13689 , w_13690 , w_13691 , w_13692 , w_13693 , w_13694 , w_13695 , 
		w_13696 , w_13697 , w_13698 , w_13699 , w_13700 , w_13701 , w_13702 , w_13703 , w_13704 , w_13705 , 
		w_13706 , w_13707 , w_13708 , w_13709 , w_13710 , w_13711 , w_13712 , w_13713 , w_13714 , w_13715 , 
		w_13716 , w_13717 , w_13718 , w_13719 , w_13720 , w_13721 , w_13722 , w_13723 , w_13724 , w_13725 , 
		w_13726 , w_13727 , w_13728 , w_13729 , w_13730 , w_13731 , w_13732 , w_13733 , w_13734 , w_13735 , 
		w_13736 , w_13737 , w_13738 , w_13739 , w_13740 , w_13741 , w_13742 , w_13743 , w_13744 , w_13745 , 
		w_13746 , w_13747 , w_13748 , w_13749 , w_13750 , w_13751 , w_13752 , w_13753 , w_13754 , w_13755 , 
		w_13756 , w_13757 , w_13758 , w_13759 , w_13760 , w_13761 , w_13762 , w_13763 , w_13764 , w_13765 , 
		w_13766 , w_13767 , w_13768 , w_13769 , w_13770 , w_13771 , w_13772 , w_13773 , w_13774 , w_13775 , 
		w_13776 , w_13777 , w_13778 , w_13779 , w_13780 , w_13781 , w_13782 , w_13783 , w_13784 , w_13785 , 
		w_13786 , w_13787 , w_13788 , w_13789 , w_13790 , w_13791 , w_13792 , w_13793 , w_13794 , w_13795 , 
		w_13796 , w_13797 , w_13798 , w_13799 , w_13800 , w_13801 , w_13802 , w_13803 , w_13804 , w_13805 , 
		w_13806 , w_13807 , w_13808 , w_13809 , w_13810 , w_13811 , w_13812 , w_13813 , w_13814 , w_13815 , 
		w_13816 , w_13817 , w_13818 , w_13819 , w_13820 , w_13821 , w_13822 , w_13823 , w_13824 , w_13825 , 
		w_13826 , w_13827 , w_13828 , w_13829 , w_13830 , w_13831 , w_13832 , w_13833 , w_13834 , w_13835 , 
		w_13836 , w_13837 , w_13838 , w_13839 , w_13840 , w_13841 , w_13842 , w_13843 , w_13844 , w_13845 , 
		w_13846 , w_13847 , w_13848 , w_13849 , w_13850 , w_13851 , w_13852 , w_13853 , w_13854 , w_13855 , 
		w_13856 , w_13857 , w_13858 , w_13859 , w_13860 , w_13861 , w_13862 , w_13863 , w_13864 , w_13865 , 
		w_13866 , w_13867 , w_13868 , w_13869 , w_13870 , w_13871 , w_13872 , w_13873 , w_13874 , w_13875 , 
		w_13876 , w_13877 , w_13878 , w_13879 , w_13880 , w_13881 , w_13882 , w_13883 , w_13884 , w_13885 , 
		w_13886 , w_13887 , w_13888 , w_13889 , w_13890 , w_13891 , w_13892 , w_13893 , w_13894 , w_13895 , 
		w_13896 , w_13897 , w_13898 , w_13899 , w_13900 , w_13901 , w_13902 , w_13903 , w_13904 , w_13905 , 
		w_13906 , w_13907 , w_13908 , w_13909 , w_13910 , w_13911 , w_13912 , w_13913 , w_13914 , w_13915 , 
		w_13916 , w_13917 , w_13918 , w_13919 , w_13920 , w_13921 , w_13922 , w_13923 , w_13924 , w_13925 , 
		w_13926 , w_13927 , w_13928 , w_13929 , w_13930 , w_13931 , w_13932 , w_13933 , w_13934 , w_13935 , 
		w_13936 , w_13937 , w_13938 , w_13939 , w_13940 , w_13941 , w_13942 , w_13943 , w_13944 , w_13945 , 
		w_13946 , w_13947 , w_13948 , w_13949 , w_13950 , w_13951 , w_13952 , w_13953 , w_13954 , w_13955 , 
		w_13956 , w_13957 , w_13958 , w_13959 , w_13960 , w_13961 , w_13962 , w_13963 , w_13964 , w_13965 , 
		w_13966 , w_13967 , w_13968 , w_13969 , w_13970 , w_13971 , w_13972 , w_13973 , w_13974 , w_13975 , 
		w_13976 , w_13977 , w_13978 , w_13979 , w_13980 , w_13981 , w_13982 , w_13983 , w_13984 , w_13985 , 
		w_13986 , w_13987 , w_13988 , w_13989 , w_13990 , w_13991 , w_13992 , w_13993 , w_13994 , w_13995 , 
		w_13996 , w_13997 , w_13998 , w_13999 , w_14000 , w_14001 , w_14002 , w_14003 , w_14004 , w_14005 , 
		w_14006 , w_14007 , w_14008 , w_14009 , w_14010 , w_14011 , w_14012 , w_14013 , w_14014 , w_14015 , 
		w_14016 , w_14017 , w_14018 , w_14019 , w_14020 , w_14021 , w_14022 , w_14023 , w_14024 , w_14025 , 
		w_14026 , w_14027 , w_14028 , w_14029 , w_14030 , w_14031 , w_14032 , w_14033 , w_14034 , w_14035 , 
		w_14036 , w_14037 , w_14038 , w_14039 , w_14040 , w_14041 , w_14042 , w_14043 , w_14044 , w_14045 , 
		w_14046 , w_14047 , w_14048 , w_14049 , w_14050 , w_14051 , w_14052 , w_14053 , w_14054 , w_14055 , 
		w_14056 , w_14057 , w_14058 , w_14059 , w_14060 , w_14061 , w_14062 , w_14063 , w_14064 , w_14065 , 
		w_14066 , w_14067 , w_14068 , w_14069 , w_14070 , w_14071 , w_14072 , w_14073 , w_14074 , w_14075 , 
		w_14076 , w_14077 , w_14078 , w_14079 , w_14080 , w_14081 , w_14082 , w_14083 , w_14084 , w_14085 , 
		w_14086 , w_14087 , w_14088 , w_14089 , w_14090 , w_14091 , w_14092 , w_14093 , w_14094 , w_14095 , 
		w_14096 , w_14097 , w_14098 , w_14099 , w_14100 , w_14101 , w_14102 , w_14103 , w_14104 , w_14105 , 
		w_14106 , w_14107 , w_14108 , w_14109 , w_14110 , w_14111 , w_14112 , w_14113 , w_14114 , w_14115 , 
		w_14116 , w_14117 , w_14118 , w_14119 , w_14120 , w_14121 , w_14122 , w_14123 , w_14124 , w_14125 , 
		w_14126 , w_14127 , w_14128 , w_14129 , w_14130 , w_14131 , w_14132 , w_14133 , w_14134 , w_14135 , 
		w_14136 , w_14137 , w_14138 , w_14139 , w_14140 , w_14141 , w_14142 , w_14143 , w_14144 , w_14145 , 
		w_14146 , w_14147 , w_14148 , w_14149 , w_14150 , w_14151 , w_14152 , w_14153 , w_14154 , w_14155 , 
		w_14156 , w_14157 , w_14158 , w_14159 , w_14160 , w_14161 , w_14162 , w_14163 , w_14164 , w_14165 , 
		w_14166 , w_14167 , w_14168 , w_14169 , w_14170 , w_14171 , w_14172 , w_14173 , w_14174 , w_14175 , 
		w_14176 , w_14177 , w_14178 , w_14179 , w_14180 , w_14181 , w_14182 , w_14183 , w_14184 , w_14185 , 
		w_14186 , w_14187 , w_14188 , w_14189 , w_14190 , w_14191 , w_14192 , w_14193 , w_14194 , w_14195 , 
		w_14196 , w_14197 , w_14198 , w_14199 , w_14200 , w_14201 , w_14202 , w_14203 , w_14204 , w_14205 , 
		w_14206 , w_14207 , w_14208 , w_14209 , w_14210 , w_14211 , w_14212 , w_14213 , w_14214 , w_14215 , 
		w_14216 , w_14217 , w_14218 , w_14219 , w_14220 , w_14221 , w_14222 , w_14223 , w_14224 , w_14225 , 
		w_14226 , w_14227 , w_14228 , w_14229 , w_14230 , w_14231 , w_14232 , w_14233 , w_14234 , w_14235 , 
		w_14236 , w_14237 , w_14238 , w_14239 , w_14240 , w_14241 , w_14242 , w_14243 , w_14244 , w_14245 , 
		w_14246 , w_14247 , w_14248 , w_14249 , w_14250 , w_14251 , w_14252 , w_14253 , w_14254 , w_14255 , 
		w_14256 , w_14257 , w_14258 , w_14259 , w_14260 , w_14261 , w_14262 , w_14263 , w_14264 , w_14265 , 
		w_14266 , w_14267 , w_14268 , w_14269 , w_14270 , w_14271 , w_14272 , w_14273 , w_14274 , w_14275 , 
		w_14276 , w_14277 , w_14278 , w_14279 , w_14280 , w_14281 , w_14282 , w_14283 , w_14284 , w_14285 , 
		w_14286 , w_14287 , w_14288 , w_14289 , w_14290 , w_14291 , w_14292 , w_14293 , w_14294 , w_14295 , 
		w_14296 , w_14297 , w_14298 , w_14299 , w_14300 , w_14301 , w_14302 , w_14303 , w_14304 , w_14305 , 
		w_14306 , w_14307 , w_14308 , w_14309 , w_14310 , w_14311 , w_14312 , w_14313 , w_14314 , w_14315 , 
		w_14316 , w_14317 , w_14318 , w_14319 , w_14320 , w_14321 , w_14322 , w_14323 , w_14324 , w_14325 , 
		w_14326 , w_14327 , w_14328 , w_14329 , w_14330 , w_14331 , w_14332 , w_14333 , w_14334 , w_14335 , 
		w_14336 , w_14337 , w_14338 , w_14339 , w_14340 , w_14341 , w_14342 , w_14343 , w_14344 , w_14345 , 
		w_14346 , w_14347 , w_14348 , w_14349 , w_14350 , w_14351 , w_14352 , w_14353 , w_14354 , w_14355 , 
		w_14356 , w_14357 , w_14358 , w_14359 , w_14360 , w_14361 , w_14362 , w_14363 , w_14364 , w_14365 , 
		w_14366 , w_14367 , w_14368 , w_14369 , w_14370 , w_14371 , w_14372 , w_14373 , w_14374 , w_14375 , 
		w_14376 , w_14377 , w_14378 , w_14379 , w_14380 , w_14381 , w_14382 , w_14383 , w_14384 , w_14385 , 
		w_14386 , w_14387 , w_14388 , w_14389 , w_14390 , w_14391 , w_14392 , w_14393 , w_14394 , w_14395 , 
		w_14396 , w_14397 , w_14398 , w_14399 , w_14400 , w_14401 , w_14402 , w_14403 , w_14404 , w_14405 , 
		w_14406 , w_14407 , w_14408 , w_14409 , w_14410 , w_14411 , w_14412 , w_14413 , w_14414 , w_14415 , 
		w_14416 , w_14417 , w_14418 , w_14419 , w_14420 , w_14421 , w_14422 , w_14423 , w_14424 , w_14425 , 
		w_14426 , w_14427 , w_14428 , w_14429 , w_14430 , w_14431 , w_14432 , w_14433 , w_14434 , w_14435 , 
		w_14436 , w_14437 , w_14438 , w_14439 , w_14440 , w_14441 , w_14442 , w_14443 , w_14444 , w_14445 , 
		w_14446 , w_14447 , w_14448 , w_14449 , w_14450 , w_14451 , w_14452 , w_14453 , w_14454 , w_14455 , 
		w_14456 , w_14457 , w_14458 , w_14459 , w_14460 , w_14461 , w_14462 , w_14463 , w_14464 , w_14465 , 
		w_14466 , w_14467 , w_14468 , w_14469 , w_14470 , w_14471 , w_14472 , w_14473 , w_14474 , w_14475 , 
		w_14476 , w_14477 , w_14478 , w_14479 , w_14480 , w_14481 , w_14482 , w_14483 , w_14484 , w_14485 , 
		w_14486 , w_14487 , w_14488 , w_14489 , w_14490 , w_14491 , w_14492 , w_14493 , w_14494 , w_14495 , 
		w_14496 , w_14497 , w_14498 , w_14499 , w_14500 , w_14501 , w_14502 , w_14503 , w_14504 , w_14505 , 
		w_14506 , w_14507 , w_14508 , w_14509 , w_14510 , w_14511 , w_14512 , w_14513 , w_14514 , w_14515 , 
		w_14516 , w_14517 , w_14518 , w_14519 , w_14520 , w_14521 , w_14522 , w_14523 , w_14524 , w_14525 , 
		w_14526 , w_14527 , w_14528 , w_14529 , w_14530 , w_14531 , w_14532 , w_14533 , w_14534 , w_14535 , 
		w_14536 , w_14537 , w_14538 , w_14539 , w_14540 , w_14541 , w_14542 , w_14543 , w_14544 , w_14545 , 
		w_14546 , w_14547 , w_14548 , w_14549 , w_14550 , w_14551 , w_14552 , w_14553 , w_14554 , w_14555 , 
		w_14556 , w_14557 , w_14558 , w_14559 , w_14560 , w_14561 , w_14562 , w_14563 , w_14564 , w_14565 , 
		w_14566 , w_14567 , w_14568 , w_14569 , w_14570 , w_14571 , w_14572 , w_14573 , w_14574 , w_14575 , 
		w_14576 , w_14577 , w_14578 , w_14579 , w_14580 , w_14581 , w_14582 , w_14583 , w_14584 , w_14585 , 
		w_14586 , w_14587 , w_14588 , w_14589 , w_14590 , w_14591 , w_14592 , w_14593 , w_14594 , w_14595 , 
		w_14596 , w_14597 , w_14598 , w_14599 , w_14600 , w_14601 , w_14602 , w_14603 , w_14604 , w_14605 , 
		w_14606 , w_14607 , w_14608 , w_14609 , w_14610 , w_14611 , w_14612 , w_14613 , w_14614 , w_14615 , 
		w_14616 , w_14617 , w_14618 , w_14619 , w_14620 , w_14621 , w_14622 , w_14623 , w_14624 , w_14625 , 
		w_14626 , w_14627 , w_14628 , w_14629 , w_14630 , w_14631 , w_14632 , w_14633 , w_14634 , w_14635 , 
		w_14636 , w_14637 , w_14638 , w_14639 , w_14640 , w_14641 , w_14642 , w_14643 , w_14644 , w_14645 , 
		w_14646 , w_14647 , w_14648 , w_14649 , w_14650 , w_14651 , w_14652 , w_14653 , w_14654 , w_14655 , 
		w_14656 , w_14657 , w_14658 , w_14659 , w_14660 , w_14661 , w_14662 , w_14663 , w_14664 , w_14665 , 
		w_14666 , w_14667 , w_14668 , w_14669 , w_14670 , w_14671 , w_14672 , w_14673 , w_14674 , w_14675 , 
		w_14676 , w_14677 , w_14678 , w_14679 , w_14680 , w_14681 , w_14682 , w_14683 , w_14684 , w_14685 , 
		w_14686 , w_14687 , w_14688 , w_14689 , w_14690 , w_14691 , w_14692 , w_14693 , w_14694 , w_14695 , 
		w_14696 , w_14697 , w_14698 , w_14699 , w_14700 , w_14701 , w_14702 , w_14703 , w_14704 , w_14705 , 
		w_14706 , w_14707 , w_14708 , w_14709 , w_14710 , w_14711 , w_14712 , w_14713 , w_14714 , w_14715 , 
		w_14716 , w_14717 , w_14718 , w_14719 , w_14720 , w_14721 , w_14722 , w_14723 , w_14724 , w_14725 , 
		w_14726 , w_14727 , w_14728 , w_14729 , w_14730 , w_14731 , w_14732 , w_14733 , w_14734 , w_14735 , 
		w_14736 , w_14737 , w_14738 , w_14739 , w_14740 , w_14741 , w_14742 , w_14743 , w_14744 , w_14745 , 
		w_14746 , w_14747 , w_14748 , w_14749 , w_14750 , w_14751 , w_14752 , w_14753 , w_14754 , w_14755 , 
		w_14756 , w_14757 , w_14758 , w_14759 , w_14760 , w_14761 , w_14762 , w_14763 , w_14764 , w_14765 , 
		w_14766 , w_14767 , w_14768 , w_14769 , w_14770 , w_14771 , w_14772 , w_14773 , w_14774 , w_14775 , 
		w_14776 , w_14777 , w_14778 , w_14779 , w_14780 , w_14781 , w_14782 , w_14783 , w_14784 , w_14785 , 
		w_14786 , w_14787 , w_14788 , w_14789 , w_14790 , w_14791 , w_14792 , w_14793 , w_14794 , w_14795 , 
		w_14796 , w_14797 , w_14798 , w_14799 , w_14800 , w_14801 , w_14802 , w_14803 , w_14804 , w_14805 , 
		w_14806 , w_14807 , w_14808 , w_14809 , w_14810 , w_14811 , w_14812 , w_14813 , w_14814 , w_14815 , 
		w_14816 , w_14817 , w_14818 , w_14819 , w_14820 , w_14821 , w_14822 , w_14823 , w_14824 , w_14825 , 
		w_14826 , w_14827 , w_14828 , w_14829 , w_14830 , w_14831 , w_14832 , w_14833 , w_14834 , w_14835 , 
		w_14836 , w_14837 , w_14838 , w_14839 , w_14840 , w_14841 , w_14842 , w_14843 , w_14844 , w_14845 , 
		w_14846 , w_14847 , w_14848 , w_14849 , w_14850 , w_14851 , w_14852 , w_14853 , w_14854 , w_14855 , 
		w_14856 , w_14857 , w_14858 , w_14859 , w_14860 , w_14861 , w_14862 , w_14863 , w_14864 , w_14865 , 
		w_14866 , w_14867 , w_14868 , w_14869 , w_14870 , w_14871 , w_14872 , w_14873 , w_14874 , w_14875 , 
		w_14876 , w_14877 , w_14878 , w_14879 , w_14880 , w_14881 , w_14882 , w_14883 , w_14884 , w_14885 , 
		w_14886 , w_14887 , w_14888 , w_14889 , w_14890 , w_14891 , w_14892 , w_14893 , w_14894 , w_14895 , 
		w_14896 , w_14897 , w_14898 , w_14899 , w_14900 , w_14901 , w_14902 , w_14903 , w_14904 , w_14905 , 
		w_14906 , w_14907 , w_14908 , w_14909 , w_14910 , w_14911 , w_14912 , w_14913 , w_14914 , w_14915 , 
		w_14916 , w_14917 , w_14918 , w_14919 , w_14920 , w_14921 , w_14922 , w_14923 , w_14924 , w_14925 , 
		w_14926 , w_14927 , w_14928 , w_14929 , w_14930 , w_14931 , w_14932 , w_14933 , w_14934 , w_14935 , 
		w_14936 , w_14937 , w_14938 , w_14939 , w_14940 , w_14941 , w_14942 , w_14943 , w_14944 , w_14945 , 
		w_14946 , w_14947 , w_14948 , w_14949 , w_14950 , w_14951 , w_14952 , w_14953 , w_14954 , w_14955 , 
		w_14956 , w_14957 , w_14958 , w_14959 , w_14960 , w_14961 , w_14962 , w_14963 , w_14964 , w_14965 , 
		w_14966 , w_14967 , w_14968 , w_14969 , w_14970 , w_14971 , w_14972 , w_14973 , w_14974 , w_14975 , 
		w_14976 , w_14977 , w_14978 , w_14979 , w_14980 , w_14981 , w_14982 , w_14983 , w_14984 , w_14985 , 
		w_14986 , w_14987 , w_14988 , w_14989 , w_14990 , w_14991 , w_14992 , w_14993 , w_14994 , w_14995 , 
		w_14996 , w_14997 , w_14998 , w_14999 , w_15000 , w_15001 , w_15002 , w_15003 , w_15004 , w_15005 , 
		w_15006 , w_15007 , w_15008 , w_15009 , w_15010 , w_15011 , w_15012 , w_15013 , w_15014 , w_15015 , 
		w_15016 , w_15017 , w_15018 , w_15019 , w_15020 , w_15021 , w_15022 , w_15023 , w_15024 , w_15025 , 
		w_15026 , w_15027 , w_15028 , w_15029 , w_15030 , w_15031 , w_15032 , w_15033 , w_15034 , w_15035 , 
		w_15036 , w_15037 , w_15038 , w_15039 , w_15040 , w_15041 , w_15042 , w_15043 , w_15044 , w_15045 , 
		w_15046 , w_15047 , w_15048 , w_15049 , w_15050 , w_15051 , w_15052 , w_15053 , w_15054 , w_15055 , 
		w_15056 , w_15057 , w_15058 , w_15059 , w_15060 , w_15061 , w_15062 , w_15063 , w_15064 , w_15065 , 
		w_15066 , w_15067 , w_15068 , w_15069 , w_15070 , w_15071 , w_15072 , w_15073 , w_15074 , w_15075 , 
		w_15076 , w_15077 , w_15078 , w_15079 , w_15080 , w_15081 , w_15082 , w_15083 , w_15084 , w_15085 , 
		w_15086 , w_15087 , w_15088 , w_15089 , w_15090 , w_15091 , w_15092 , w_15093 , w_15094 , w_15095 , 
		w_15096 , w_15097 , w_15098 , w_15099 , w_15100 , w_15101 , w_15102 , w_15103 , w_15104 , w_15105 , 
		w_15106 , w_15107 , w_15108 , w_15109 , w_15110 , w_15111 , w_15112 , w_15113 , w_15114 , w_15115 , 
		w_15116 , w_15117 , w_15118 , w_15119 , w_15120 , w_15121 , w_15122 , w_15123 , w_15124 , w_15125 , 
		w_15126 , w_15127 , w_15128 , w_15129 , w_15130 , w_15131 , w_15132 , w_15133 , w_15134 , w_15135 , 
		w_15136 , w_15137 , w_15138 , w_15139 , w_15140 , w_15141 , w_15142 , w_15143 , w_15144 , w_15145 , 
		w_15146 , w_15147 , w_15148 , w_15149 , w_15150 , w_15151 , w_15152 , w_15153 , w_15154 , w_15155 , 
		w_15156 , w_15157 , w_15158 , w_15159 , w_15160 , w_15161 , w_15162 , w_15163 , w_15164 , w_15165 , 
		w_15166 , w_15167 , w_15168 , w_15169 , w_15170 , w_15171 , w_15172 , w_15173 , w_15174 , w_15175 , 
		w_15176 , w_15177 , w_15178 , w_15179 , w_15180 , w_15181 , w_15182 , w_15183 , w_15184 , w_15185 , 
		w_15186 , w_15187 , w_15188 , w_15189 , w_15190 , w_15191 , w_15192 , w_15193 , w_15194 , w_15195 , 
		w_15196 , w_15197 , w_15198 , w_15199 , w_15200 , w_15201 , w_15202 , w_15203 , w_15204 , w_15205 , 
		w_15206 , w_15207 , w_15208 , w_15209 , w_15210 , w_15211 , w_15212 , w_15213 , w_15214 , w_15215 , 
		w_15216 , w_15217 , w_15218 , w_15219 , w_15220 , w_15221 , w_15222 , w_15223 , w_15224 , w_15225 , 
		w_15226 , w_15227 , w_15228 , w_15229 , w_15230 , w_15231 , w_15232 , w_15233 , w_15234 , w_15235 , 
		w_15236 , w_15237 , w_15238 , w_15239 , w_15240 , w_15241 , w_15242 , w_15243 , w_15244 , w_15245 , 
		w_15246 , w_15247 , w_15248 , w_15249 , w_15250 , w_15251 , w_15252 , w_15253 , w_15254 , w_15255 , 
		w_15256 , w_15257 , w_15258 , w_15259 , w_15260 , w_15261 , w_15262 , w_15263 , w_15264 , w_15265 , 
		w_15266 , w_15267 , w_15268 , w_15269 , w_15270 , w_15271 , w_15272 , w_15273 , w_15274 , w_15275 , 
		w_15276 , w_15277 , w_15278 , w_15279 , w_15280 , w_15281 , w_15282 , w_15283 , w_15284 , w_15285 , 
		w_15286 , w_15287 , w_15288 , w_15289 , w_15290 , w_15291 , w_15292 , w_15293 , w_15294 , w_15295 , 
		w_15296 , w_15297 , w_15298 , w_15299 , w_15300 , w_15301 , w_15302 , w_15303 , w_15304 , w_15305 , 
		w_15306 , w_15307 , w_15308 , w_15309 , w_15310 , w_15311 , w_15312 , w_15313 , w_15314 , w_15315 , 
		w_15316 , w_15317 , w_15318 , w_15319 , w_15320 , w_15321 , w_15322 , w_15323 , w_15324 , w_15325 , 
		w_15326 , w_15327 , w_15328 , w_15329 , w_15330 , w_15331 , w_15332 , w_15333 , w_15334 , w_15335 , 
		w_15336 , w_15337 , w_15338 , w_15339 , w_15340 , w_15341 , w_15342 , w_15343 , w_15344 , w_15345 , 
		w_15346 , w_15347 , w_15348 , w_15349 , w_15350 , w_15351 , w_15352 , w_15353 , w_15354 , w_15355 , 
		w_15356 , w_15357 , w_15358 , w_15359 , w_15360 , w_15361 , w_15362 , w_15363 , w_15364 , w_15365 , 
		w_15366 , w_15367 , w_15368 , w_15369 , w_15370 , w_15371 , w_15372 , w_15373 , w_15374 , w_15375 , 
		w_15376 , w_15377 , w_15378 , w_15379 , w_15380 , w_15381 , w_15382 , w_15383 , w_15384 , w_15385 , 
		w_15386 , w_15387 , w_15388 , w_15389 , w_15390 , w_15391 , w_15392 , w_15393 , w_15394 , w_15395 , 
		w_15396 , w_15397 , w_15398 , w_15399 , w_15400 , w_15401 , w_15402 , w_15403 , w_15404 , w_15405 , 
		w_15406 , w_15407 , w_15408 , w_15409 , w_15410 , w_15411 , w_15412 , w_15413 , w_15414 , w_15415 , 
		w_15416 , w_15417 , w_15418 , w_15419 , w_15420 , w_15421 , w_15422 , w_15423 , w_15424 , w_15425 , 
		w_15426 , w_15427 , w_15428 , w_15429 , w_15430 , w_15431 , w_15432 , w_15433 , w_15434 , w_15435 , 
		w_15436 , w_15437 , w_15438 , w_15439 , w_15440 , w_15441 , w_15442 , w_15443 , w_15444 , w_15445 , 
		w_15446 , w_15447 , w_15448 , w_15449 , w_15450 , w_15451 , w_15452 , w_15453 , w_15454 , w_15455 , 
		w_15456 , w_15457 , w_15458 , w_15459 , w_15460 , w_15461 , w_15462 , w_15463 , w_15464 , w_15465 , 
		w_15466 , w_15467 , w_15468 , w_15469 , w_15470 , w_15471 , w_15472 , w_15473 , w_15474 , w_15475 , 
		w_15476 , w_15477 , w_15478 , w_15479 , w_15480 , w_15481 , w_15482 , w_15483 , w_15484 , w_15485 , 
		w_15486 , w_15487 , w_15488 , w_15489 , w_15490 , w_15491 , w_15492 , w_15493 , w_15494 , w_15495 , 
		w_15496 , w_15497 , w_15498 , w_15499 , w_15500 , w_15501 , w_15502 , w_15503 , w_15504 , w_15505 , 
		w_15506 , w_15507 , w_15508 , w_15509 , w_15510 , w_15511 , w_15512 , w_15513 , w_15514 , w_15515 , 
		w_15516 , w_15517 , w_15518 , w_15519 , w_15520 , w_15521 , w_15522 , w_15523 , w_15524 , w_15525 , 
		w_15526 , w_15527 , w_15528 , w_15529 , w_15530 , w_15531 , w_15532 , w_15533 , w_15534 , w_15535 , 
		w_15536 , w_15537 , w_15538 , w_15539 , w_15540 , w_15541 , w_15542 , w_15543 , w_15544 , w_15545 , 
		w_15546 , w_15547 , w_15548 , w_15549 , w_15550 , w_15551 , w_15552 , w_15553 , w_15554 , w_15555 , 
		w_15556 , w_15557 , w_15558 , w_15559 , w_15560 , w_15561 , w_15562 , w_15563 , w_15564 , w_15565 , 
		w_15566 , w_15567 , w_15568 , w_15569 , w_15570 , w_15571 , w_15572 , w_15573 , w_15574 , w_15575 , 
		w_15576 , w_15577 , w_15578 , w_15579 , w_15580 , w_15581 , w_15582 , w_15583 , w_15584 , w_15585 , 
		w_15586 , w_15587 , w_15588 , w_15589 , w_15590 , w_15591 , w_15592 , w_15593 , w_15594 , w_15595 , 
		w_15596 , w_15597 , w_15598 , w_15599 , w_15600 , w_15601 , w_15602 , w_15603 , w_15604 , w_15605 , 
		w_15606 , w_15607 , w_15608 , w_15609 , w_15610 , w_15611 , w_15612 , w_15613 , w_15614 , w_15615 , 
		w_15616 , w_15617 , w_15618 , w_15619 , w_15620 , w_15621 , w_15622 , w_15623 , w_15624 , w_15625 , 
		w_15626 , w_15627 , w_15628 , w_15629 , w_15630 , w_15631 , w_15632 , w_15633 , w_15634 , w_15635 , 
		w_15636 , w_15637 , w_15638 , w_15639 , w_15640 , w_15641 , w_15642 , w_15643 , w_15644 , w_15645 , 
		w_15646 , w_15647 , w_15648 , w_15649 , w_15650 , w_15651 , w_15652 , w_15653 , w_15654 , w_15655 , 
		w_15656 , w_15657 , w_15658 , w_15659 , w_15660 , w_15661 , w_15662 , w_15663 , w_15664 , w_15665 , 
		w_15666 , w_15667 , w_15668 , w_15669 , w_15670 , w_15671 , w_15672 , w_15673 , w_15674 , w_15675 , 
		w_15676 , w_15677 , w_15678 , w_15679 , w_15680 , w_15681 , w_15682 , w_15683 , w_15684 , w_15685 , 
		w_15686 , w_15687 , w_15688 , w_15689 , w_15690 , w_15691 , w_15692 , w_15693 , w_15694 , w_15695 , 
		w_15696 , w_15697 , w_15698 , w_15699 , w_15700 , w_15701 , w_15702 , w_15703 , w_15704 , w_15705 , 
		w_15706 , w_15707 , w_15708 , w_15709 , w_15710 , w_15711 , w_15712 , w_15713 , w_15714 , w_15715 , 
		w_15716 , w_15717 , w_15718 , w_15719 , w_15720 , w_15721 , w_15722 , w_15723 , w_15724 , w_15725 , 
		w_15726 , w_15727 , w_15728 , w_15729 , w_15730 , w_15731 , w_15732 , w_15733 , w_15734 , w_15735 , 
		w_15736 , w_15737 , w_15738 , w_15739 , w_15740 , w_15741 , w_15742 , w_15743 , w_15744 , w_15745 , 
		w_15746 , w_15747 , w_15748 , w_15749 , w_15750 , w_15751 , w_15752 , w_15753 , w_15754 , w_15755 , 
		w_15756 , w_15757 , w_15758 , w_15759 , w_15760 , w_15761 , w_15762 , w_15763 , w_15764 , w_15765 , 
		w_15766 , w_15767 , w_15768 , w_15769 , w_15770 , w_15771 , w_15772 , w_15773 , w_15774 , w_15775 , 
		w_15776 , w_15777 , w_15778 , w_15779 , w_15780 , w_15781 , w_15782 , w_15783 , w_15784 , w_15785 , 
		w_15786 , w_15787 , w_15788 , w_15789 , w_15790 , w_15791 , w_15792 , w_15793 , w_15794 , w_15795 , 
		w_15796 , w_15797 , w_15798 , w_15799 , w_15800 , w_15801 , w_15802 , w_15803 , w_15804 , w_15805 , 
		w_15806 , w_15807 , w_15808 , w_15809 , w_15810 , w_15811 , w_15812 , w_15813 , w_15814 , w_15815 , 
		w_15816 , w_15817 , w_15818 , w_15819 , w_15820 , w_15821 , w_15822 , w_15823 , w_15824 , w_15825 , 
		w_15826 , w_15827 , w_15828 , w_15829 , w_15830 , w_15831 , w_15832 , w_15833 , w_15834 , w_15835 , 
		w_15836 , w_15837 , w_15838 , w_15839 , w_15840 , w_15841 , w_15842 , w_15843 , w_15844 , w_15845 , 
		w_15846 , w_15847 , w_15848 , w_15849 , w_15850 , w_15851 , w_15852 , w_15853 , w_15854 , w_15855 , 
		w_15856 , w_15857 , w_15858 , w_15859 , w_15860 , w_15861 , w_15862 , w_15863 , w_15864 , w_15865 , 
		w_15866 , w_15867 , w_15868 , w_15869 , w_15870 , w_15871 , w_15872 , w_15873 , w_15874 , w_15875 , 
		w_15876 , w_15877 , w_15878 , w_15879 , w_15880 , w_15881 , w_15882 , w_15883 , w_15884 , w_15885 , 
		w_15886 , w_15887 , w_15888 , w_15889 , w_15890 , w_15891 , w_15892 , w_15893 , w_15894 , w_15895 , 
		w_15896 , w_15897 , w_15898 , w_15899 , w_15900 , w_15901 , w_15902 , w_15903 , w_15904 , w_15905 , 
		w_15906 , w_15907 , w_15908 , w_15909 , w_15910 , w_15911 , w_15912 , w_15913 , w_15914 , w_15915 , 
		w_15916 , w_15917 , w_15918 , w_15919 , w_15920 , w_15921 , w_15922 , w_15923 , w_15924 , w_15925 , 
		w_15926 , w_15927 , w_15928 , w_15929 , w_15930 , w_15931 , w_15932 , w_15933 , w_15934 , w_15935 , 
		w_15936 , w_15937 , w_15938 , w_15939 , w_15940 , w_15941 , w_15942 , w_15943 , w_15944 , w_15945 , 
		w_15946 , w_15947 , w_15948 , w_15949 , w_15950 , w_15951 , w_15952 , w_15953 , w_15954 , w_15955 , 
		w_15956 , w_15957 , w_15958 , w_15959 , w_15960 , w_15961 , w_15962 , w_15963 , w_15964 , w_15965 , 
		w_15966 , w_15967 , w_15968 , w_15969 , w_15970 , w_15971 , w_15972 , w_15973 , w_15974 , w_15975 , 
		w_15976 , w_15977 , w_15978 , w_15979 , w_15980 , w_15981 , w_15982 , w_15983 , w_15984 , w_15985 , 
		w_15986 , w_15987 , w_15988 , w_15989 , w_15990 , w_15991 , w_15992 , w_15993 , w_15994 , w_15995 , 
		w_15996 , w_15997 , w_15998 , w_15999 , w_16000 , w_16001 , w_16002 , w_16003 , w_16004 , w_16005 , 
		w_16006 , w_16007 , w_16008 , w_16009 , w_16010 , w_16011 , w_16012 , w_16013 , w_16014 , w_16015 , 
		w_16016 , w_16017 , w_16018 , w_16019 , w_16020 , w_16021 , w_16022 , w_16023 , w_16024 , w_16025 , 
		w_16026 , w_16027 , w_16028 , w_16029 , w_16030 , w_16031 , w_16032 , w_16033 , w_16034 , w_16035 , 
		w_16036 , w_16037 , w_16038 , w_16039 , w_16040 , w_16041 , w_16042 , w_16043 , w_16044 , w_16045 , 
		w_16046 , w_16047 , w_16048 , w_16049 , w_16050 , w_16051 , w_16052 , w_16053 , w_16054 , w_16055 , 
		w_16056 , w_16057 , w_16058 , w_16059 , w_16060 , w_16061 , w_16062 , w_16063 , w_16064 , w_16065 , 
		w_16066 , w_16067 , w_16068 , w_16069 , w_16070 , w_16071 , w_16072 , w_16073 , w_16074 , w_16075 , 
		w_16076 , w_16077 , w_16078 , w_16079 , w_16080 , w_16081 , w_16082 , w_16083 , w_16084 , w_16085 , 
		w_16086 , w_16087 , w_16088 , w_16089 , w_16090 , w_16091 , w_16092 , w_16093 , w_16094 , w_16095 , 
		w_16096 , w_16097 , w_16098 , w_16099 , w_16100 , w_16101 , w_16102 , w_16103 , w_16104 , w_16105 , 
		w_16106 , w_16107 , w_16108 , w_16109 , w_16110 , w_16111 , w_16112 , w_16113 , w_16114 , w_16115 , 
		w_16116 , w_16117 , w_16118 , w_16119 , w_16120 , w_16121 , w_16122 , w_16123 , w_16124 , w_16125 , 
		w_16126 , w_16127 , w_16128 , w_16129 , w_16130 , w_16131 , w_16132 , w_16133 , w_16134 , w_16135 , 
		w_16136 , w_16137 , w_16138 , w_16139 , w_16140 , w_16141 , w_16142 , w_16143 , w_16144 , w_16145 , 
		w_16146 , w_16147 , w_16148 , w_16149 , w_16150 , w_16151 , w_16152 , w_16153 , w_16154 , w_16155 , 
		w_16156 , w_16157 , w_16158 , w_16159 , w_16160 , w_16161 , w_16162 , w_16163 , w_16164 , w_16165 , 
		w_16166 , w_16167 , w_16168 , w_16169 , w_16170 , w_16171 , w_16172 , w_16173 , w_16174 , w_16175 , 
		w_16176 , w_16177 , w_16178 , w_16179 , w_16180 , w_16181 , w_16182 , w_16183 , w_16184 , w_16185 , 
		w_16186 , w_16187 , w_16188 , w_16189 , w_16190 , w_16191 , w_16192 , w_16193 , w_16194 , w_16195 , 
		w_16196 , w_16197 , w_16198 , w_16199 , w_16200 , w_16201 , w_16202 , w_16203 , w_16204 , w_16205 , 
		w_16206 , w_16207 , w_16208 , w_16209 , w_16210 , w_16211 , w_16212 , w_16213 , w_16214 , w_16215 , 
		w_16216 , w_16217 , w_16218 , w_16219 , w_16220 , w_16221 , w_16222 , w_16223 , w_16224 , w_16225 , 
		w_16226 , w_16227 , w_16228 , w_16229 , w_16230 , w_16231 , w_16232 , w_16233 , w_16234 , w_16235 , 
		w_16236 , w_16237 , w_16238 , w_16239 , w_16240 , w_16241 , w_16242 , w_16243 , w_16244 , w_16245 , 
		w_16246 , w_16247 , w_16248 , w_16249 , w_16250 , w_16251 , w_16252 , w_16253 , w_16254 , w_16255 , 
		w_16256 , w_16257 , w_16258 , w_16259 , w_16260 , w_16261 , w_16262 , w_16263 , w_16264 , w_16265 , 
		w_16266 , w_16267 , w_16268 , w_16269 , w_16270 , w_16271 , w_16272 , w_16273 , w_16274 , w_16275 , 
		w_16276 , w_16277 , w_16278 , w_16279 , w_16280 , w_16281 , w_16282 , w_16283 , w_16284 , w_16285 , 
		w_16286 , w_16287 , w_16288 , w_16289 , w_16290 , w_16291 , w_16292 , w_16293 , w_16294 , w_16295 , 
		w_16296 , w_16297 , w_16298 , w_16299 , w_16300 , w_16301 , w_16302 , w_16303 , w_16304 , w_16305 , 
		w_16306 , w_16307 , w_16308 , w_16309 , w_16310 , w_16311 , w_16312 , w_16313 , w_16314 , w_16315 , 
		w_16316 , w_16317 , w_16318 , w_16319 , w_16320 , w_16321 , w_16322 , w_16323 , w_16324 , w_16325 , 
		w_16326 , w_16327 , w_16328 , w_16329 , w_16330 , w_16331 , w_16332 , w_16333 , w_16334 , w_16335 , 
		w_16336 , w_16337 , w_16338 , w_16339 , w_16340 , w_16341 , w_16342 , w_16343 , w_16344 , w_16345 , 
		w_16346 , w_16347 , w_16348 , w_16349 , w_16350 , w_16351 , w_16352 , w_16353 , w_16354 , w_16355 , 
		w_16356 , w_16357 , w_16358 , w_16359 , w_16360 , w_16361 , w_16362 , w_16363 , w_16364 , w_16365 , 
		w_16366 , w_16367 , w_16368 , w_16369 , w_16370 , w_16371 , w_16372 , w_16373 , w_16374 , w_16375 , 
		w_16376 , w_16377 , w_16378 , w_16379 , w_16380 , w_16381 , w_16382 , w_16383 , w_16384 , w_16385 , 
		w_16386 , w_16387 , w_16388 , w_16389 , w_16390 , w_16391 , w_16392 , w_16393 , w_16394 , w_16395 , 
		w_16396 , w_16397 , w_16398 , w_16399 , w_16400 , w_16401 , w_16402 , w_16403 , w_16404 , w_16405 , 
		w_16406 , w_16407 , w_16408 , w_16409 , w_16410 , w_16411 , w_16412 , w_16413 , w_16414 , w_16415 , 
		w_16416 , w_16417 , w_16418 , w_16419 , w_16420 , w_16421 , w_16422 , w_16423 , w_16424 , w_16425 , 
		w_16426 , w_16427 , w_16428 , w_16429 , w_16430 , w_16431 , w_16432 , w_16433 , w_16434 , w_16435 , 
		w_16436 , w_16437 , w_16438 , w_16439 , w_16440 , w_16441 , w_16442 , w_16443 , w_16444 , w_16445 , 
		w_16446 , w_16447 , w_16448 , w_16449 , w_16450 , w_16451 , w_16452 , w_16453 , w_16454 , w_16455 , 
		w_16456 , w_16457 , w_16458 , w_16459 , w_16460 , w_16461 , w_16462 , w_16463 , w_16464 , w_16465 , 
		w_16466 , w_16467 , w_16468 , w_16469 , w_16470 , w_16471 , w_16472 , w_16473 , w_16474 , w_16475 , 
		w_16476 , w_16477 , w_16478 , w_16479 , w_16480 , w_16481 , w_16482 , w_16483 , w_16484 , w_16485 , 
		w_16486 , w_16487 , w_16488 , w_16489 , w_16490 , w_16491 , w_16492 , w_16493 , w_16494 , w_16495 , 
		w_16496 , w_16497 , w_16498 , w_16499 , w_16500 , w_16501 , w_16502 , w_16503 , w_16504 , w_16505 , 
		w_16506 , w_16507 , w_16508 , w_16509 , w_16510 , w_16511 , w_16512 , w_16513 , w_16514 , w_16515 , 
		w_16516 , w_16517 , w_16518 , w_16519 , w_16520 , w_16521 , w_16522 , w_16523 , w_16524 , w_16525 , 
		w_16526 , w_16527 , w_16528 , w_16529 , w_16530 , w_16531 , w_16532 , w_16533 , w_16534 , w_16535 , 
		w_16536 , w_16537 , w_16538 , w_16539 , w_16540 , w_16541 , w_16542 , w_16543 , w_16544 , w_16545 , 
		w_16546 , w_16547 , w_16548 , w_16549 , w_16550 , w_16551 , w_16552 , w_16553 , w_16554 , w_16555 , 
		w_16556 , w_16557 , w_16558 , w_16559 , w_16560 , w_16561 , w_16562 , w_16563 , w_16564 , w_16565 , 
		w_16566 , w_16567 , w_16568 , w_16569 , w_16570 , w_16571 , w_16572 , w_16573 , w_16574 , w_16575 , 
		w_16576 , w_16577 , w_16578 , w_16579 , w_16580 , w_16581 , w_16582 , w_16583 , w_16584 , w_16585 , 
		w_16586 , w_16587 , w_16588 , w_16589 , w_16590 , w_16591 , w_16592 , w_16593 , w_16594 , w_16595 , 
		w_16596 , w_16597 , w_16598 , w_16599 , w_16600 , w_16601 , w_16602 , w_16603 , w_16604 , w_16605 , 
		w_16606 , w_16607 , w_16608 , w_16609 , w_16610 , w_16611 , w_16612 , w_16613 , w_16614 , w_16615 , 
		w_16616 , w_16617 , w_16618 , w_16619 , w_16620 , w_16621 , w_16622 , w_16623 , w_16624 , w_16625 , 
		w_16626 , w_16627 , w_16628 , w_16629 , w_16630 , w_16631 , w_16632 , w_16633 , w_16634 , w_16635 , 
		w_16636 , w_16637 , w_16638 , w_16639 , w_16640 , w_16641 , w_16642 , w_16643 , w_16644 , w_16645 , 
		w_16646 , w_16647 , w_16648 , w_16649 , w_16650 , w_16651 , w_16652 , w_16653 , w_16654 , w_16655 , 
		w_16656 , w_16657 , w_16658 , w_16659 , w_16660 , w_16661 , w_16662 , w_16663 , w_16664 , w_16665 , 
		w_16666 , w_16667 , w_16668 , w_16669 , w_16670 , w_16671 , w_16672 , w_16673 , w_16674 , w_16675 , 
		w_16676 , w_16677 , w_16678 , w_16679 , w_16680 , w_16681 , w_16682 , w_16683 , w_16684 , w_16685 , 
		w_16686 , w_16687 , w_16688 , w_16689 , w_16690 , w_16691 , w_16692 , w_16693 , w_16694 , w_16695 , 
		w_16696 , w_16697 , w_16698 , w_16699 , w_16700 , w_16701 , w_16702 , w_16703 , w_16704 , w_16705 , 
		w_16706 , w_16707 , w_16708 , w_16709 , w_16710 , w_16711 , w_16712 , w_16713 , w_16714 , w_16715 , 
		w_16716 , w_16717 , w_16718 , w_16719 , w_16720 , w_16721 , w_16722 , w_16723 , w_16724 , w_16725 , 
		w_16726 , w_16727 , w_16728 , w_16729 , w_16730 , w_16731 , w_16732 , w_16733 , w_16734 , w_16735 , 
		w_16736 , w_16737 , w_16738 , w_16739 , w_16740 , w_16741 , w_16742 , w_16743 , w_16744 , w_16745 , 
		w_16746 , w_16747 , w_16748 , w_16749 , w_16750 , w_16751 , w_16752 , w_16753 , w_16754 , w_16755 , 
		w_16756 , w_16757 , w_16758 , w_16759 , w_16760 , w_16761 , w_16762 , w_16763 , w_16764 , w_16765 , 
		w_16766 , w_16767 , w_16768 , w_16769 , w_16770 , w_16771 , w_16772 , w_16773 , w_16774 , w_16775 , 
		w_16776 , w_16777 , w_16778 , w_16779 , w_16780 , w_16781 , w_16782 , w_16783 , w_16784 , w_16785 , 
		w_16786 , w_16787 , w_16788 , w_16789 , w_16790 , w_16791 , w_16792 , w_16793 , w_16794 , w_16795 , 
		w_16796 , w_16797 , w_16798 , w_16799 , w_16800 , w_16801 , w_16802 , w_16803 , w_16804 , w_16805 , 
		w_16806 , w_16807 , w_16808 , w_16809 , w_16810 , w_16811 , w_16812 , w_16813 , w_16814 , w_16815 , 
		w_16816 , w_16817 , w_16818 , w_16819 , w_16820 , w_16821 , w_16822 , w_16823 , w_16824 , w_16825 , 
		w_16826 , w_16827 , w_16828 , w_16829 , w_16830 , w_16831 , w_16832 , w_16833 , w_16834 , w_16835 , 
		w_16836 , w_16837 , w_16838 , w_16839 , w_16840 , w_16841 , w_16842 , w_16843 , w_16844 , w_16845 , 
		w_16846 , w_16847 , w_16848 , w_16849 , w_16850 , w_16851 , w_16852 , w_16853 , w_16854 , w_16855 , 
		w_16856 , w_16857 , w_16858 , w_16859 , w_16860 , w_16861 , w_16862 , w_16863 , w_16864 , w_16865 , 
		w_16866 , w_16867 , w_16868 , w_16869 , w_16870 , w_16871 , w_16872 , w_16873 , w_16874 , w_16875 , 
		w_16876 , w_16877 , w_16878 , w_16879 , w_16880 , w_16881 , w_16882 , w_16883 , w_16884 , w_16885 , 
		w_16886 , w_16887 , w_16888 , w_16889 , w_16890 , w_16891 , w_16892 , w_16893 , w_16894 , w_16895 , 
		w_16896 , w_16897 , w_16898 , w_16899 , w_16900 , w_16901 , w_16902 , w_16903 , w_16904 , w_16905 , 
		w_16906 , w_16907 , w_16908 , w_16909 , w_16910 , w_16911 , w_16912 , w_16913 , w_16914 , w_16915 , 
		w_16916 , w_16917 , w_16918 , w_16919 , w_16920 , w_16921 , w_16922 , w_16923 , w_16924 , w_16925 , 
		w_16926 , w_16927 , w_16928 , w_16929 , w_16930 , w_16931 , w_16932 , w_16933 , w_16934 , w_16935 , 
		w_16936 , w_16937 , w_16938 , w_16939 , w_16940 , w_16941 , w_16942 , w_16943 , w_16944 , w_16945 , 
		w_16946 , w_16947 , w_16948 , w_16949 , w_16950 , w_16951 , w_16952 , w_16953 , w_16954 , w_16955 , 
		w_16956 , w_16957 , w_16958 , w_16959 , w_16960 , w_16961 , w_16962 , w_16963 , w_16964 , w_16965 , 
		w_16966 , w_16967 , w_16968 , w_16969 , w_16970 , w_16971 , w_16972 , w_16973 , w_16974 , w_16975 , 
		w_16976 , w_16977 , w_16978 , w_16979 , w_16980 , w_16981 , w_16982 , w_16983 , w_16984 , w_16985 , 
		w_16986 , w_16987 , w_16988 , w_16989 , w_16990 , w_16991 , w_16992 , w_16993 , w_16994 , w_16995 , 
		w_16996 , w_16997 , w_16998 , w_16999 , w_17000 , w_17001 , w_17002 , w_17003 , w_17004 , w_17005 , 
		w_17006 , w_17007 , w_17008 , w_17009 , w_17010 , w_17011 , w_17012 , w_17013 , w_17014 , w_17015 , 
		w_17016 , w_17017 , w_17018 , w_17019 , w_17020 , w_17021 , w_17022 , w_17023 , w_17024 , w_17025 , 
		w_17026 , w_17027 , w_17028 , w_17029 , w_17030 , w_17031 , w_17032 , w_17033 , w_17034 , w_17035 , 
		w_17036 , w_17037 , w_17038 , w_17039 , w_17040 , w_17041 , w_17042 , w_17043 , w_17044 , w_17045 , 
		w_17046 , w_17047 , w_17048 , w_17049 , w_17050 , w_17051 , w_17052 , w_17053 , w_17054 , w_17055 , 
		w_17056 , w_17057 , w_17058 , w_17059 , w_17060 , w_17061 , w_17062 , w_17063 , w_17064 , w_17065 , 
		w_17066 , w_17067 , w_17068 , w_17069 , w_17070 , w_17071 , w_17072 , w_17073 , w_17074 , w_17075 , 
		w_17076 , w_17077 , w_17078 , w_17079 , w_17080 , w_17081 , w_17082 , w_17083 , w_17084 , w_17085 , 
		w_17086 , w_17087 , w_17088 , w_17089 , w_17090 , w_17091 , w_17092 , w_17093 , w_17094 , w_17095 , 
		w_17096 , w_17097 , w_17098 , w_17099 , w_17100 , w_17101 , w_17102 , w_17103 , w_17104 , w_17105 , 
		w_17106 , w_17107 , w_17108 , w_17109 , w_17110 , w_17111 , w_17112 , w_17113 , w_17114 , w_17115 , 
		w_17116 , w_17117 , w_17118 , w_17119 , w_17120 , w_17121 , w_17122 , w_17123 , w_17124 , w_17125 , 
		w_17126 , w_17127 , w_17128 , w_17129 , w_17130 , w_17131 , w_17132 , w_17133 , w_17134 , w_17135 , 
		w_17136 , w_17137 , w_17138 , w_17139 , w_17140 , w_17141 , w_17142 , w_17143 , w_17144 , w_17145 , 
		w_17146 , w_17147 , w_17148 , w_17149 , w_17150 , w_17151 , w_17152 , w_17153 , w_17154 , w_17155 , 
		w_17156 , w_17157 , w_17158 , w_17159 , w_17160 , w_17161 , w_17162 , w_17163 , w_17164 , w_17165 , 
		w_17166 , w_17167 , w_17168 , w_17169 , w_17170 , w_17171 , w_17172 , w_17173 , w_17174 , w_17175 , 
		w_17176 , w_17177 , w_17178 , w_17179 , w_17180 , w_17181 , w_17182 , w_17183 , w_17184 , w_17185 , 
		w_17186 , w_17187 , w_17188 , w_17189 , w_17190 , w_17191 , w_17192 , w_17193 , w_17194 , w_17195 , 
		w_17196 , w_17197 , w_17198 , w_17199 , w_17200 , w_17201 , w_17202 , w_17203 , w_17204 , w_17205 , 
		w_17206 , w_17207 , w_17208 , w_17209 , w_17210 , w_17211 , w_17212 , w_17213 , w_17214 , w_17215 , 
		w_17216 , w_17217 , w_17218 , w_17219 , w_17220 , w_17221 , w_17222 , w_17223 , w_17224 , w_17225 , 
		w_17226 , w_17227 , w_17228 , w_17229 , w_17230 , w_17231 , w_17232 , w_17233 , w_17234 , w_17235 , 
		w_17236 , w_17237 , w_17238 , w_17239 , w_17240 , w_17241 , w_17242 , w_17243 , w_17244 , w_17245 , 
		w_17246 , w_17247 , w_17248 , w_17249 , w_17250 , w_17251 , w_17252 , w_17253 , w_17254 , w_17255 , 
		w_17256 , w_17257 , w_17258 , w_17259 , w_17260 , w_17261 , w_17262 , w_17263 , w_17264 , w_17265 , 
		w_17266 , w_17267 , w_17268 , w_17269 , w_17270 , w_17271 , w_17272 , w_17273 , w_17274 , w_17275 , 
		w_17276 , w_17277 , w_17278 , w_17279 , w_17280 , w_17281 , w_17282 , w_17283 , w_17284 , w_17285 , 
		w_17286 , w_17287 , w_17288 , w_17289 , w_17290 , w_17291 , w_17292 , w_17293 , w_17294 , w_17295 , 
		w_17296 , w_17297 , w_17298 , w_17299 , w_17300 , w_17301 , w_17302 , w_17303 , w_17304 , w_17305 , 
		w_17306 , w_17307 , w_17308 , w_17309 , w_17310 , w_17311 , w_17312 , w_17313 , w_17314 , w_17315 , 
		w_17316 , w_17317 , w_17318 , w_17319 , w_17320 , w_17321 , w_17322 , w_17323 , w_17324 , w_17325 , 
		w_17326 , w_17327 , w_17328 , w_17329 , w_17330 , w_17331 , w_17332 , w_17333 , w_17334 , w_17335 , 
		w_17336 , w_17337 , w_17338 , w_17339 , w_17340 , w_17341 , w_17342 , w_17343 , w_17344 , w_17345 , 
		w_17346 , w_17347 , w_17348 , w_17349 , w_17350 , w_17351 , w_17352 , w_17353 , w_17354 , w_17355 , 
		w_17356 , w_17357 , w_17358 , w_17359 , w_17360 , w_17361 , w_17362 , w_17363 , w_17364 , w_17365 , 
		w_17366 , w_17367 , w_17368 , w_17369 , w_17370 , w_17371 , w_17372 , w_17373 , w_17374 , w_17375 , 
		w_17376 , w_17377 , w_17378 , w_17379 , w_17380 , w_17381 , w_17382 , w_17383 , w_17384 , w_17385 , 
		w_17386 , w_17387 , w_17388 , w_17389 , w_17390 , w_17391 , w_17392 , w_17393 , w_17394 , w_17395 , 
		w_17396 , w_17397 , w_17398 , w_17399 , w_17400 , w_17401 , w_17402 , w_17403 , w_17404 , w_17405 , 
		w_17406 , w_17407 , w_17408 , w_17409 , w_17410 , w_17411 , w_17412 , w_17413 , w_17414 , w_17415 , 
		w_17416 , w_17417 , w_17418 , w_17419 , w_17420 , w_17421 , w_17422 , w_17423 , w_17424 , w_17425 , 
		w_17426 , w_17427 , w_17428 , w_17429 , w_17430 , w_17431 , w_17432 , w_17433 , w_17434 , w_17435 , 
		w_17436 , w_17437 , w_17438 , w_17439 , w_17440 , w_17441 , w_17442 , w_17443 , w_17444 , w_17445 , 
		w_17446 , w_17447 , w_17448 , w_17449 , w_17450 , w_17451 , w_17452 , w_17453 , w_17454 , w_17455 , 
		w_17456 , w_17457 , w_17458 , w_17459 , w_17460 , w_17461 , w_17462 , w_17463 , w_17464 , w_17465 , 
		w_17466 , w_17467 , w_17468 , w_17469 , w_17470 , w_17471 , w_17472 , w_17473 , w_17474 , w_17475 , 
		w_17476 , w_17477 , w_17478 , w_17479 , w_17480 , w_17481 , w_17482 , w_17483 , w_17484 , w_17485 , 
		w_17486 , w_17487 , w_17488 , w_17489 , w_17490 , w_17491 , w_17492 , w_17493 , w_17494 , w_17495 , 
		w_17496 , w_17497 , w_17498 , w_17499 , w_17500 , w_17501 , w_17502 , w_17503 , w_17504 , w_17505 , 
		w_17506 , w_17507 , w_17508 , w_17509 , w_17510 , w_17511 , w_17512 , w_17513 , w_17514 , w_17515 , 
		w_17516 , w_17517 , w_17518 , w_17519 , w_17520 , w_17521 , w_17522 , w_17523 , w_17524 , w_17525 , 
		w_17526 , w_17527 , w_17528 , w_17529 , w_17530 , w_17531 , w_17532 , w_17533 , w_17534 , w_17535 , 
		w_17536 , w_17537 , w_17538 , w_17539 , w_17540 , w_17541 , w_17542 , w_17543 , w_17544 , w_17545 , 
		w_17546 , w_17547 , w_17548 , w_17549 , w_17550 , w_17551 , w_17552 , w_17553 , w_17554 , w_17555 , 
		w_17556 , w_17557 , w_17558 , w_17559 , w_17560 , w_17561 , w_17562 , w_17563 , w_17564 , w_17565 , 
		w_17566 , w_17567 , w_17568 , w_17569 , w_17570 , w_17571 , w_17572 , w_17573 , w_17574 , w_17575 , 
		w_17576 , w_17577 , w_17578 , w_17579 , w_17580 , w_17581 , w_17582 , w_17583 , w_17584 , w_17585 , 
		w_17586 , w_17587 , w_17588 , w_17589 , w_17590 , w_17591 , w_17592 , w_17593 , w_17594 , w_17595 , 
		w_17596 , w_17597 , w_17598 , w_17599 , w_17600 , w_17601 , w_17602 , w_17603 , w_17604 , w_17605 , 
		w_17606 , w_17607 , w_17608 , w_17609 , w_17610 , w_17611 , w_17612 , w_17613 , w_17614 , w_17615 , 
		w_17616 , w_17617 , w_17618 , w_17619 , w_17620 , w_17621 , w_17622 , w_17623 , w_17624 , w_17625 , 
		w_17626 , w_17627 , w_17628 , w_17629 , w_17630 , w_17631 , w_17632 , w_17633 , w_17634 , w_17635 , 
		w_17636 , w_17637 , w_17638 , w_17639 , w_17640 , w_17641 , w_17642 , w_17643 , w_17644 , w_17645 , 
		w_17646 , w_17647 , w_17648 , w_17649 , w_17650 , w_17651 , w_17652 , w_17653 , w_17654 , w_17655 , 
		w_17656 , w_17657 , w_17658 , w_17659 , w_17660 , w_17661 , w_17662 , w_17663 , w_17664 , w_17665 , 
		w_17666 , w_17667 , w_17668 , w_17669 , w_17670 , w_17671 , w_17672 , w_17673 , w_17674 , w_17675 , 
		w_17676 , w_17677 , w_17678 , w_17679 , w_17680 , w_17681 , w_17682 , w_17683 , w_17684 , w_17685 , 
		w_17686 , w_17687 , w_17688 , w_17689 , w_17690 , w_17691 , w_17692 , w_17693 , w_17694 , w_17695 , 
		w_17696 , w_17697 , w_17698 , w_17699 , w_17700 , w_17701 , w_17702 , w_17703 , w_17704 , w_17705 , 
		w_17706 , w_17707 , w_17708 , w_17709 , w_17710 , w_17711 , w_17712 , w_17713 , w_17714 , w_17715 , 
		w_17716 , w_17717 , w_17718 , w_17719 , w_17720 , w_17721 , w_17722 , w_17723 , w_17724 , w_17725 , 
		w_17726 , w_17727 , w_17728 , w_17729 , w_17730 , w_17731 , w_17732 , w_17733 , w_17734 , w_17735 , 
		w_17736 , w_17737 , w_17738 , w_17739 , w_17740 , w_17741 , w_17742 , w_17743 , w_17744 , w_17745 , 
		w_17746 , w_17747 , w_17748 , w_17749 , w_17750 , w_17751 , w_17752 , w_17753 , w_17754 , w_17755 , 
		w_17756 , w_17757 , w_17758 , w_17759 , w_17760 , w_17761 , w_17762 , w_17763 , w_17764 , w_17765 , 
		w_17766 , w_17767 , w_17768 , w_17769 , w_17770 , w_17771 , w_17772 , w_17773 , w_17774 , w_17775 , 
		w_17776 , w_17777 , w_17778 , w_17779 , w_17780 , w_17781 , w_17782 , w_17783 , w_17784 , w_17785 , 
		w_17786 , w_17787 , w_17788 , w_17789 , w_17790 , w_17791 , w_17792 , w_17793 , w_17794 , w_17795 , 
		w_17796 , w_17797 , w_17798 , w_17799 , w_17800 , w_17801 , w_17802 , w_17803 , w_17804 , w_17805 , 
		w_17806 , w_17807 , w_17808 , w_17809 , w_17810 , w_17811 , w_17812 , w_17813 , w_17814 , w_17815 , 
		w_17816 , w_17817 , w_17818 , w_17819 , w_17820 , w_17821 , w_17822 , w_17823 , w_17824 , w_17825 , 
		w_17826 , w_17827 , w_17828 , w_17829 , w_17830 , w_17831 , w_17832 , w_17833 , w_17834 , w_17835 , 
		w_17836 , w_17837 , w_17838 , w_17839 , w_17840 , w_17841 , w_17842 , w_17843 , w_17844 , w_17845 , 
		w_17846 , w_17847 , w_17848 , w_17849 , w_17850 , w_17851 , w_17852 , w_17853 , w_17854 , w_17855 , 
		w_17856 , w_17857 , w_17858 , w_17859 , w_17860 , w_17861 , w_17862 , w_17863 , w_17864 , w_17865 , 
		w_17866 , w_17867 , w_17868 , w_17869 , w_17870 , w_17871 , w_17872 , w_17873 , w_17874 , w_17875 , 
		w_17876 , w_17877 , w_17878 , w_17879 , w_17880 , w_17881 , w_17882 , w_17883 , w_17884 , w_17885 , 
		w_17886 , w_17887 , w_17888 , w_17889 , w_17890 , w_17891 , w_17892 , w_17893 , w_17894 , w_17895 , 
		w_17896 , w_17897 , w_17898 , w_17899 , w_17900 , w_17901 , w_17902 , w_17903 , w_17904 , w_17905 , 
		w_17906 , w_17907 , w_17908 , w_17909 , w_17910 , w_17911 , w_17912 , w_17913 , w_17914 , w_17915 , 
		w_17916 , w_17917 , w_17918 , w_17919 , w_17920 , w_17921 , w_17922 , w_17923 , w_17924 , w_17925 , 
		w_17926 , w_17927 , w_17928 , w_17929 , w_17930 , w_17931 , w_17932 , w_17933 , w_17934 , w_17935 , 
		w_17936 , w_17937 , w_17938 , w_17939 , w_17940 , w_17941 , w_17942 , w_17943 , w_17944 , w_17945 , 
		w_17946 , w_17947 , w_17948 , w_17949 , w_17950 , w_17951 , w_17952 , w_17953 , w_17954 , w_17955 , 
		w_17956 , w_17957 , w_17958 , w_17959 , w_17960 , w_17961 , w_17962 , w_17963 , w_17964 , w_17965 , 
		w_17966 , w_17967 , w_17968 , w_17969 , w_17970 , w_17971 , w_17972 , w_17973 , w_17974 , w_17975 , 
		w_17976 , w_17977 , w_17978 , w_17979 , w_17980 , w_17981 , w_17982 , w_17983 , w_17984 , w_17985 , 
		w_17986 , w_17987 , w_17988 , w_17989 , w_17990 , w_17991 , w_17992 , w_17993 , w_17994 , w_17995 , 
		w_17996 , w_17997 , w_17998 , w_17999 , w_18000 , w_18001 , w_18002 , w_18003 , w_18004 , w_18005 , 
		w_18006 , w_18007 , w_18008 , w_18009 , w_18010 , w_18011 , w_18012 , w_18013 , w_18014 , w_18015 , 
		w_18016 , w_18017 , w_18018 , w_18019 , w_18020 , w_18021 , w_18022 , w_18023 , w_18024 , w_18025 , 
		w_18026 , w_18027 , w_18028 , w_18029 , w_18030 , w_18031 , w_18032 , w_18033 , w_18034 , w_18035 , 
		w_18036 , w_18037 , w_18038 , w_18039 , w_18040 , w_18041 , w_18042 , w_18043 , w_18044 , w_18045 , 
		w_18046 , w_18047 , w_18048 , w_18049 , w_18050 , w_18051 , w_18052 , w_18053 , w_18054 , w_18055 , 
		w_18056 , w_18057 , w_18058 , w_18059 , w_18060 , w_18061 , w_18062 , w_18063 , w_18064 , w_18065 , 
		w_18066 , w_18067 , w_18068 , w_18069 , w_18070 , w_18071 , w_18072 , w_18073 , w_18074 , w_18075 , 
		w_18076 , w_18077 , w_18078 , w_18079 , w_18080 , w_18081 , w_18082 , w_18083 , w_18084 , w_18085 , 
		w_18086 , w_18087 , w_18088 , w_18089 , w_18090 , w_18091 , w_18092 , w_18093 , w_18094 , w_18095 , 
		w_18096 , w_18097 , w_18098 , w_18099 , w_18100 , w_18101 , w_18102 , w_18103 , w_18104 , w_18105 , 
		w_18106 , w_18107 , w_18108 , w_18109 , w_18110 , w_18111 , w_18112 , w_18113 , w_18114 , w_18115 , 
		w_18116 , w_18117 , w_18118 , w_18119 , w_18120 , w_18121 , w_18122 , w_18123 , w_18124 , w_18125 , 
		w_18126 , w_18127 , w_18128 , w_18129 , w_18130 , w_18131 , w_18132 , w_18133 , w_18134 , w_18135 , 
		w_18136 , w_18137 , w_18138 , w_18139 , w_18140 , w_18141 , w_18142 , w_18143 , w_18144 , w_18145 , 
		w_18146 , w_18147 , w_18148 , w_18149 , w_18150 , w_18151 , w_18152 , w_18153 , w_18154 , w_18155 , 
		w_18156 , w_18157 , w_18158 , w_18159 , w_18160 , w_18161 , w_18162 , w_18163 , w_18164 , w_18165 , 
		w_18166 , w_18167 , w_18168 , w_18169 , w_18170 , w_18171 , w_18172 , w_18173 , w_18174 , w_18175 , 
		w_18176 , w_18177 , w_18178 , w_18179 , w_18180 , w_18181 , w_18182 , w_18183 , w_18184 , w_18185 , 
		w_18186 , w_18187 , w_18188 , w_18189 , w_18190 , w_18191 , w_18192 , w_18193 , w_18194 , w_18195 , 
		w_18196 , w_18197 , w_18198 , w_18199 , w_18200 , w_18201 , w_18202 , w_18203 , w_18204 , w_18205 , 
		w_18206 , w_18207 , w_18208 , w_18209 , w_18210 , w_18211 , w_18212 , w_18213 , w_18214 , w_18215 , 
		w_18216 , w_18217 , w_18218 , w_18219 , w_18220 , w_18221 , w_18222 , w_18223 , w_18224 , w_18225 , 
		w_18226 , w_18227 , w_18228 , w_18229 , w_18230 , w_18231 , w_18232 , w_18233 , w_18234 , w_18235 , 
		w_18236 , w_18237 , w_18238 , w_18239 , w_18240 , w_18241 , w_18242 , w_18243 , w_18244 , w_18245 , 
		w_18246 , w_18247 , w_18248 , w_18249 , w_18250 , w_18251 , w_18252 , w_18253 , w_18254 , w_18255 , 
		w_18256 , w_18257 , w_18258 , w_18259 , w_18260 , w_18261 , w_18262 , w_18263 , w_18264 , w_18265 , 
		w_18266 , w_18267 , w_18268 , w_18269 , w_18270 , w_18271 , w_18272 , w_18273 , w_18274 , w_18275 , 
		w_18276 , w_18277 , w_18278 , w_18279 , w_18280 , w_18281 , w_18282 , w_18283 , w_18284 , w_18285 , 
		w_18286 , w_18287 , w_18288 , w_18289 , w_18290 , w_18291 , w_18292 , w_18293 , w_18294 , w_18295 , 
		w_18296 , w_18297 , w_18298 , w_18299 , w_18300 , w_18301 , w_18302 , w_18303 , w_18304 , w_18305 , 
		w_18306 , w_18307 , w_18308 , w_18309 , w_18310 , w_18311 , w_18312 , w_18313 , w_18314 , w_18315 , 
		w_18316 , w_18317 , w_18318 , w_18319 , w_18320 , w_18321 , w_18322 , w_18323 , w_18324 , w_18325 , 
		w_18326 , w_18327 , w_18328 , w_18329 , w_18330 , w_18331 , w_18332 , w_18333 , w_18334 , w_18335 , 
		w_18336 , w_18337 , w_18338 , w_18339 , w_18340 , w_18341 , w_18342 , w_18343 , w_18344 , w_18345 , 
		w_18346 , w_18347 , w_18348 , w_18349 , w_18350 , w_18351 , w_18352 , w_18353 , w_18354 , w_18355 , 
		w_18356 , w_18357 , w_18358 , w_18359 , w_18360 , w_18361 , w_18362 , w_18363 , w_18364 , w_18365 , 
		w_18366 , w_18367 , w_18368 , w_18369 , w_18370 , w_18371 , w_18372 , w_18373 , w_18374 , w_18375 , 
		w_18376 , w_18377 , w_18378 , w_18379 , w_18380 , w_18381 , w_18382 , w_18383 , w_18384 , w_18385 , 
		w_18386 , w_18387 , w_18388 , w_18389 , w_18390 , w_18391 , w_18392 , w_18393 , w_18394 , w_18395 , 
		w_18396 , w_18397 , w_18398 , w_18399 , w_18400 , w_18401 , w_18402 , w_18403 , w_18404 , w_18405 , 
		w_18406 , w_18407 , w_18408 , w_18409 , w_18410 , w_18411 , w_18412 , w_18413 , w_18414 , w_18415 , 
		w_18416 , w_18417 , w_18418 , w_18419 , w_18420 , w_18421 , w_18422 , w_18423 , w_18424 , w_18425 , 
		w_18426 , w_18427 , w_18428 , w_18429 , w_18430 , w_18431 , w_18432 , w_18433 , w_18434 , w_18435 , 
		w_18436 , w_18437 , w_18438 , w_18439 , w_18440 , w_18441 , w_18442 , w_18443 , w_18444 , w_18445 , 
		w_18446 , w_18447 , w_18448 , w_18449 , w_18450 , w_18451 , w_18452 , w_18453 , w_18454 , w_18455 , 
		w_18456 , w_18457 , w_18458 , w_18459 , w_18460 , w_18461 , w_18462 , w_18463 , w_18464 , w_18465 , 
		w_18466 , w_18467 , w_18468 , w_18469 , w_18470 , w_18471 , w_18472 , w_18473 , w_18474 , w_18475 , 
		w_18476 , w_18477 , w_18478 , w_18479 , w_18480 , w_18481 , w_18482 , w_18483 , w_18484 , w_18485 , 
		w_18486 , w_18487 , w_18488 , w_18489 , w_18490 , w_18491 , w_18492 , w_18493 , w_18494 , w_18495 , 
		w_18496 , w_18497 , w_18498 , w_18499 , w_18500 , w_18501 , w_18502 , w_18503 , w_18504 , w_18505 , 
		w_18506 , w_18507 , w_18508 , w_18509 , w_18510 , w_18511 , w_18512 , w_18513 , w_18514 , w_18515 , 
		w_18516 , w_18517 , w_18518 , w_18519 , w_18520 , w_18521 , w_18522 , w_18523 , w_18524 , w_18525 , 
		w_18526 , w_18527 , w_18528 , w_18529 , w_18530 , w_18531 , w_18532 , w_18533 , w_18534 , w_18535 , 
		w_18536 , w_18537 , w_18538 , w_18539 , w_18540 , w_18541 , w_18542 , w_18543 , w_18544 , w_18545 , 
		w_18546 , w_18547 , w_18548 , w_18549 , w_18550 , w_18551 , w_18552 , w_18553 , w_18554 , w_18555 , 
		w_18556 , w_18557 , w_18558 , w_18559 , w_18560 , w_18561 , w_18562 , w_18563 , w_18564 , w_18565 , 
		w_18566 , w_18567 , w_18568 , w_18569 , w_18570 , w_18571 , w_18572 , w_18573 , w_18574 , w_18575 , 
		w_18576 , w_18577 , w_18578 , w_18579 , w_18580 , w_18581 , w_18582 , w_18583 , w_18584 , w_18585 , 
		w_18586 , w_18587 , w_18588 , w_18589 , w_18590 , w_18591 , w_18592 , w_18593 , w_18594 , w_18595 , 
		w_18596 , w_18597 , w_18598 , w_18599 , w_18600 , w_18601 , w_18602 , w_18603 , w_18604 , w_18605 , 
		w_18606 , w_18607 , w_18608 , w_18609 , w_18610 , w_18611 , w_18612 , w_18613 , w_18614 , w_18615 , 
		w_18616 , w_18617 , w_18618 , w_18619 , w_18620 , w_18621 , w_18622 , w_18623 , w_18624 , w_18625 , 
		w_18626 , w_18627 , w_18628 , w_18629 , w_18630 , w_18631 , w_18632 , w_18633 , w_18634 , w_18635 , 
		w_18636 , w_18637 , w_18638 , w_18639 , w_18640 , w_18641 , w_18642 , w_18643 , w_18644 , w_18645 , 
		w_18646 , w_18647 , w_18648 , w_18649 , w_18650 , w_18651 , w_18652 , w_18653 , w_18654 , w_18655 , 
		w_18656 , w_18657 , w_18658 , w_18659 , w_18660 , w_18661 , w_18662 , w_18663 , w_18664 , w_18665 , 
		w_18666 , w_18667 , w_18668 , w_18669 , w_18670 , w_18671 , w_18672 , w_18673 , w_18674 , w_18675 , 
		w_18676 , w_18677 , w_18678 , w_18679 , w_18680 , w_18681 , w_18682 , w_18683 , w_18684 , w_18685 , 
		w_18686 , w_18687 , w_18688 , w_18689 , w_18690 , w_18691 , w_18692 , w_18693 , w_18694 , w_18695 , 
		w_18696 , w_18697 , w_18698 , w_18699 , w_18700 , w_18701 , w_18702 , w_18703 , w_18704 , w_18705 , 
		w_18706 , w_18707 , w_18708 , w_18709 , w_18710 , w_18711 , w_18712 , w_18713 , w_18714 , w_18715 , 
		w_18716 , w_18717 , w_18718 , w_18719 , w_18720 , w_18721 , w_18722 , w_18723 , w_18724 , w_18725 , 
		w_18726 , w_18727 , w_18728 , w_18729 , w_18730 , w_18731 , w_18732 , w_18733 , w_18734 , w_18735 , 
		w_18736 , w_18737 , w_18738 , w_18739 , w_18740 , w_18741 , w_18742 , w_18743 , w_18744 , w_18745 , 
		w_18746 , w_18747 , w_18748 , w_18749 , w_18750 , w_18751 , w_18752 , w_18753 , w_18754 , w_18755 , 
		w_18756 , w_18757 , w_18758 , w_18759 , w_18760 , w_18761 , w_18762 , w_18763 , w_18764 , w_18765 , 
		w_18766 , w_18767 , w_18768 , w_18769 , w_18770 , w_18771 , w_18772 , w_18773 , w_18774 , w_18775 , 
		w_18776 , w_18777 , w_18778 , w_18779 , w_18780 , w_18781 , w_18782 , w_18783 , w_18784 , w_18785 , 
		w_18786 , w_18787 , w_18788 , w_18789 , w_18790 , w_18791 , w_18792 , w_18793 , w_18794 , w_18795 , 
		w_18796 , w_18797 , w_18798 , w_18799 , w_18800 , w_18801 , w_18802 , w_18803 , w_18804 , w_18805 , 
		w_18806 , w_18807 , w_18808 , w_18809 , w_18810 , w_18811 , w_18812 , w_18813 , w_18814 , w_18815 , 
		w_18816 , w_18817 , w_18818 , w_18819 , w_18820 , w_18821 , w_18822 , w_18823 , w_18824 , w_18825 , 
		w_18826 , w_18827 , w_18828 , w_18829 , w_18830 , w_18831 , w_18832 , w_18833 , w_18834 , w_18835 , 
		w_18836 , w_18837 , w_18838 , w_18839 , w_18840 , w_18841 , w_18842 , w_18843 , w_18844 , w_18845 , 
		w_18846 , w_18847 , w_18848 , w_18849 , w_18850 , w_18851 , w_18852 , w_18853 , w_18854 , w_18855 , 
		w_18856 , w_18857 , w_18858 , w_18859 , w_18860 , w_18861 , w_18862 , w_18863 , w_18864 , w_18865 , 
		w_18866 , w_18867 , w_18868 , w_18869 , w_18870 , w_18871 , w_18872 , w_18873 , w_18874 , w_18875 , 
		w_18876 , w_18877 , w_18878 , w_18879 , w_18880 , w_18881 , w_18882 , w_18883 , w_18884 , w_18885 , 
		w_18886 , w_18887 , w_18888 , w_18889 , w_18890 , w_18891 , w_18892 , w_18893 , w_18894 , w_18895 , 
		w_18896 , w_18897 , w_18898 , w_18899 , w_18900 , w_18901 , w_18902 , w_18903 , w_18904 , w_18905 , 
		w_18906 , w_18907 , w_18908 , w_18909 , w_18910 , w_18911 , w_18912 , w_18913 , w_18914 , w_18915 , 
		w_18916 , w_18917 , w_18918 , w_18919 , w_18920 , w_18921 , w_18922 , w_18923 , w_18924 , w_18925 , 
		w_18926 , w_18927 , w_18928 , w_18929 , w_18930 , w_18931 , w_18932 , w_18933 , w_18934 , w_18935 , 
		w_18936 , w_18937 , w_18938 , w_18939 , w_18940 , w_18941 , w_18942 , w_18943 , w_18944 , w_18945 , 
		w_18946 , w_18947 , w_18948 , w_18949 , w_18950 , w_18951 , w_18952 , w_18953 , w_18954 , w_18955 , 
		w_18956 , w_18957 , w_18958 , w_18959 , w_18960 , w_18961 , w_18962 , w_18963 , w_18964 , w_18965 , 
		w_18966 , w_18967 , w_18968 , w_18969 , w_18970 , w_18971 , w_18972 , w_18973 , w_18974 , w_18975 , 
		w_18976 , w_18977 , w_18978 , w_18979 , w_18980 , w_18981 , w_18982 , w_18983 , w_18984 , w_18985 , 
		w_18986 , w_18987 , w_18988 , w_18989 , w_18990 , w_18991 , w_18992 , w_18993 , w_18994 , w_18995 , 
		w_18996 , w_18997 , w_18998 , w_18999 , w_19000 , w_19001 , w_19002 , w_19003 , w_19004 , w_19005 , 
		w_19006 , w_19007 , w_19008 , w_19009 , w_19010 , w_19011 , w_19012 , w_19013 , w_19014 , w_19015 , 
		w_19016 , w_19017 , w_19018 , w_19019 , w_19020 , w_19021 , w_19022 , w_19023 , w_19024 , w_19025 , 
		w_19026 , w_19027 , w_19028 , w_19029 , w_19030 , w_19031 , w_19032 , w_19033 , w_19034 , w_19035 , 
		w_19036 , w_19037 , w_19038 , w_19039 , w_19040 , w_19041 , w_19042 , w_19043 , w_19044 , w_19045 , 
		w_19046 , w_19047 , w_19048 , w_19049 , w_19050 , w_19051 , w_19052 , w_19053 , w_19054 , w_19055 , 
		w_19056 , w_19057 , w_19058 , w_19059 , w_19060 , w_19061 , w_19062 , w_19063 , w_19064 , w_19065 , 
		w_19066 , w_19067 , w_19068 , w_19069 , w_19070 , w_19071 , w_19072 , w_19073 , w_19074 , w_19075 , 
		w_19076 , w_19077 , w_19078 , w_19079 , w_19080 , w_19081 , w_19082 , w_19083 , w_19084 , w_19085 , 
		w_19086 , w_19087 , w_19088 , w_19089 , w_19090 , w_19091 , w_19092 , w_19093 , w_19094 , w_19095 , 
		w_19096 , w_19097 , w_19098 , w_19099 , w_19100 , w_19101 , w_19102 , w_19103 , w_19104 , w_19105 , 
		w_19106 , w_19107 , w_19108 , w_19109 , w_19110 , w_19111 , w_19112 , w_19113 , w_19114 , w_19115 , 
		w_19116 , w_19117 , w_19118 , w_19119 , w_19120 , w_19121 , w_19122 , w_19123 , w_19124 , w_19125 , 
		w_19126 , w_19127 , w_19128 , w_19129 , w_19130 , w_19131 , w_19132 , w_19133 , w_19134 , w_19135 , 
		w_19136 , w_19137 , w_19138 , w_19139 , w_19140 , w_19141 , w_19142 , w_19143 , w_19144 , w_19145 , 
		w_19146 , w_19147 , w_19148 , w_19149 , w_19150 , w_19151 , w_19152 , w_19153 , w_19154 , w_19155 , 
		w_19156 , w_19157 , w_19158 , w_19159 , w_19160 , w_19161 , w_19162 , w_19163 , w_19164 , w_19165 , 
		w_19166 , w_19167 , w_19168 , w_19169 , w_19170 , w_19171 , w_19172 , w_19173 , w_19174 , w_19175 , 
		w_19176 , w_19177 , w_19178 , w_19179 , w_19180 , w_19181 , w_19182 , w_19183 , w_19184 , w_19185 , 
		w_19186 , w_19187 , w_19188 , w_19189 , w_19190 , w_19191 , w_19192 , w_19193 , w_19194 , w_19195 , 
		w_19196 , w_19197 , w_19198 , w_19199 , w_19200 , w_19201 , w_19202 , w_19203 , w_19204 , w_19205 , 
		w_19206 , w_19207 , w_19208 , w_19209 , w_19210 , w_19211 , w_19212 , w_19213 , w_19214 , w_19215 , 
		w_19216 , w_19217 , w_19218 , w_19219 , w_19220 , w_19221 , w_19222 , w_19223 , w_19224 , w_19225 , 
		w_19226 , w_19227 , w_19228 , w_19229 , w_19230 , w_19231 , w_19232 , w_19233 , w_19234 , w_19235 , 
		w_19236 , w_19237 , w_19238 , w_19239 , w_19240 , w_19241 , w_19242 , w_19243 , w_19244 , w_19245 , 
		w_19246 , w_19247 , w_19248 , w_19249 , w_19250 , w_19251 , w_19252 , w_19253 , w_19254 , w_19255 , 
		w_19256 , w_19257 , w_19258 , w_19259 , w_19260 , w_19261 , w_19262 , w_19263 , w_19264 , w_19265 , 
		w_19266 , w_19267 , w_19268 , w_19269 , w_19270 , w_19271 , w_19272 , w_19273 , w_19274 , w_19275 , 
		w_19276 , w_19277 , w_19278 , w_19279 , w_19280 , w_19281 , w_19282 , w_19283 , w_19284 , w_19285 , 
		w_19286 , w_19287 , w_19288 , w_19289 , w_19290 , w_19291 , w_19292 , w_19293 , w_19294 , w_19295 , 
		w_19296 , w_19297 , w_19298 , w_19299 , w_19300 , w_19301 , w_19302 , w_19303 , w_19304 , w_19305 , 
		w_19306 , w_19307 , w_19308 , w_19309 , w_19310 , w_19311 , w_19312 , w_19313 , w_19314 , w_19315 , 
		w_19316 , w_19317 , w_19318 , w_19319 , w_19320 , w_19321 , w_19322 , w_19323 , w_19324 , w_19325 , 
		w_19326 , w_19327 , w_19328 , w_19329 , w_19330 , w_19331 , w_19332 , w_19333 , w_19334 , w_19335 , 
		w_19336 , w_19337 , w_19338 , w_19339 , w_19340 , w_19341 , w_19342 , w_19343 , w_19344 , w_19345 , 
		w_19346 , w_19347 , w_19348 , w_19349 , w_19350 , w_19351 , w_19352 , w_19353 , w_19354 , w_19355 , 
		w_19356 , w_19357 , w_19358 , w_19359 , w_19360 , w_19361 , w_19362 , w_19363 , w_19364 , w_19365 , 
		w_19366 , w_19367 , w_19368 , w_19369 , w_19370 , w_19371 , w_19372 , w_19373 , w_19374 , w_19375 , 
		w_19376 , w_19377 , w_19378 , w_19379 , w_19380 , w_19381 , w_19382 , w_19383 , w_19384 , w_19385 , 
		w_19386 , w_19387 , w_19388 , w_19389 , w_19390 , w_19391 , w_19392 , w_19393 , w_19394 , w_19395 , 
		w_19396 , w_19397 , w_19398 , w_19399 , w_19400 , w_19401 , w_19402 , w_19403 , w_19404 , w_19405 , 
		w_19406 , w_19407 , w_19408 , w_19409 , w_19410 , w_19411 , w_19412 , w_19413 , w_19414 , w_19415 , 
		w_19416 , w_19417 , w_19418 , w_19419 , w_19420 , w_19421 , w_19422 , w_19423 , w_19424 , w_19425 , 
		w_19426 , w_19427 , w_19428 , w_19429 , w_19430 , w_19431 , w_19432 , w_19433 , w_19434 , w_19435 , 
		w_19436 , w_19437 , w_19438 , w_19439 , w_19440 , w_19441 , w_19442 , w_19443 , w_19444 , w_19445 , 
		w_19446 , w_19447 , w_19448 , w_19449 , w_19450 , w_19451 , w_19452 , w_19453 , w_19454 , w_19455 , 
		w_19456 , w_19457 , w_19458 , w_19459 , w_19460 , w_19461 , w_19462 , w_19463 , w_19464 , w_19465 , 
		w_19466 , w_19467 , w_19468 , w_19469 , w_19470 , w_19471 , w_19472 , w_19473 , w_19474 , w_19475 , 
		w_19476 , w_19477 , w_19478 , w_19479 , w_19480 , w_19481 , w_19482 , w_19483 , w_19484 , w_19485 , 
		w_19486 , w_19487 , w_19488 , w_19489 , w_19490 , w_19491 , w_19492 , w_19493 , w_19494 , w_19495 , 
		w_19496 , w_19497 , w_19498 , w_19499 , w_19500 , w_19501 , w_19502 , w_19503 , w_19504 , w_19505 , 
		w_19506 , w_19507 , w_19508 , w_19509 , w_19510 , w_19511 , w_19512 , w_19513 , w_19514 , w_19515 , 
		w_19516 , w_19517 , w_19518 , w_19519 , w_19520 , w_19521 , w_19522 , w_19523 , w_19524 , w_19525 , 
		w_19526 , w_19527 , w_19528 , w_19529 , w_19530 , w_19531 , w_19532 , w_19533 , w_19534 , w_19535 , 
		w_19536 , w_19537 , w_19538 , w_19539 , w_19540 , w_19541 , w_19542 , w_19543 , w_19544 , w_19545 , 
		w_19546 , w_19547 , w_19548 , w_19549 , w_19550 , w_19551 , w_19552 , w_19553 , w_19554 , w_19555 , 
		w_19556 , w_19557 , w_19558 , w_19559 , w_19560 , w_19561 , w_19562 , w_19563 , w_19564 , w_19565 , 
		w_19566 , w_19567 , w_19568 , w_19569 , w_19570 , w_19571 , w_19572 , w_19573 , w_19574 , w_19575 , 
		w_19576 , w_19577 , w_19578 , w_19579 , w_19580 , w_19581 , w_19582 , w_19583 , w_19584 , w_19585 , 
		w_19586 , w_19587 , w_19588 , w_19589 , w_19590 , w_19591 , w_19592 , w_19593 , w_19594 , w_19595 , 
		w_19596 , w_19597 , w_19598 , w_19599 , w_19600 , w_19601 , w_19602 , w_19603 , w_19604 , w_19605 , 
		w_19606 , w_19607 , w_19608 , w_19609 , w_19610 , w_19611 , w_19612 , w_19613 , w_19614 , w_19615 , 
		w_19616 , w_19617 , w_19618 , w_19619 , w_19620 , w_19621 , w_19622 , w_19623 , w_19624 , w_19625 , 
		w_19626 , w_19627 , w_19628 , w_19629 , w_19630 , w_19631 , w_19632 , w_19633 , w_19634 , w_19635 , 
		w_19636 , w_19637 , w_19638 , w_19639 , w_19640 , w_19641 , w_19642 , w_19643 , w_19644 , w_19645 , 
		w_19646 , w_19647 , w_19648 , w_19649 , w_19650 , w_19651 , w_19652 , w_19653 , w_19654 , w_19655 , 
		w_19656 , w_19657 , w_19658 , w_19659 , w_19660 , w_19661 , w_19662 , w_19663 , w_19664 , w_19665 , 
		w_19666 , w_19667 , w_19668 , w_19669 , w_19670 , w_19671 , w_19672 , w_19673 , w_19674 , w_19675 , 
		w_19676 , w_19677 , w_19678 , w_19679 , w_19680 , w_19681 , w_19682 , w_19683 , w_19684 , w_19685 , 
		w_19686 , w_19687 , w_19688 , w_19689 , w_19690 , w_19691 , w_19692 , w_19693 , w_19694 , w_19695 , 
		w_19696 , w_19697 , w_19698 , w_19699 , w_19700 , w_19701 , w_19702 , w_19703 , w_19704 , w_19705 , 
		w_19706 , w_19707 , w_19708 , w_19709 , w_19710 , w_19711 , w_19712 , w_19713 , w_19714 , w_19715 , 
		w_19716 , w_19717 , w_19718 , w_19719 , w_19720 , w_19721 , w_19722 , w_19723 , w_19724 , w_19725 , 
		w_19726 , w_19727 , w_19728 , w_19729 , w_19730 , w_19731 , w_19732 , w_19733 , w_19734 , w_19735 , 
		w_19736 , w_19737 , w_19738 , w_19739 , w_19740 , w_19741 , w_19742 , w_19743 , w_19744 , w_19745 , 
		w_19746 , w_19747 , w_19748 , w_19749 , w_19750 , w_19751 , w_19752 , w_19753 , w_19754 , w_19755 , 
		w_19756 , w_19757 , w_19758 , w_19759 , w_19760 , w_19761 , w_19762 , w_19763 , w_19764 , w_19765 , 
		w_19766 , w_19767 , w_19768 , w_19769 , w_19770 , w_19771 , w_19772 , w_19773 , w_19774 , w_19775 , 
		w_19776 , w_19777 , w_19778 , w_19779 , w_19780 , w_19781 , w_19782 , w_19783 , w_19784 , w_19785 , 
		w_19786 , w_19787 , w_19788 , w_19789 , w_19790 , w_19791 , w_19792 , w_19793 , w_19794 , w_19795 , 
		w_19796 , w_19797 , w_19798 , w_19799 , w_19800 , w_19801 , w_19802 , w_19803 , w_19804 , w_19805 , 
		w_19806 , w_19807 , w_19808 , w_19809 , w_19810 , w_19811 , w_19812 , w_19813 , w_19814 , w_19815 , 
		w_19816 , w_19817 , w_19818 , w_19819 , w_19820 , w_19821 , w_19822 , w_19823 , w_19824 , w_19825 , 
		w_19826 , w_19827 , w_19828 , w_19829 , w_19830 , w_19831 , w_19832 , w_19833 , w_19834 , w_19835 , 
		w_19836 , w_19837 , w_19838 , w_19839 , w_19840 , w_19841 , w_19842 , w_19843 , w_19844 , w_19845 , 
		w_19846 , w_19847 , w_19848 , w_19849 , w_19850 , w_19851 , w_19852 , w_19853 , w_19854 , w_19855 , 
		w_19856 , w_19857 , w_19858 , w_19859 , w_19860 , w_19861 , w_19862 , w_19863 , w_19864 , w_19865 , 
		w_19866 , w_19867 , w_19868 , w_19869 , w_19870 , w_19871 , w_19872 , w_19873 , w_19874 , w_19875 , 
		w_19876 , w_19877 , w_19878 , w_19879 , w_19880 , w_19881 , w_19882 , w_19883 , w_19884 , w_19885 , 
		w_19886 , w_19887 , w_19888 , w_19889 , w_19890 , w_19891 , w_19892 , w_19893 , w_19894 , w_19895 , 
		w_19896 , w_19897 , w_19898 , w_19899 , w_19900 , w_19901 , w_19902 , w_19903 , w_19904 , w_19905 , 
		w_19906 , w_19907 , w_19908 , w_19909 , w_19910 , w_19911 , w_19912 , w_19913 , w_19914 , w_19915 , 
		w_19916 , w_19917 , w_19918 , w_19919 , w_19920 , w_19921 , w_19922 , w_19923 , w_19924 , w_19925 , 
		w_19926 , w_19927 , w_19928 , w_19929 , w_19930 , w_19931 , w_19932 , w_19933 , w_19934 , w_19935 , 
		w_19936 , w_19937 , w_19938 , w_19939 , w_19940 , w_19941 , w_19942 , w_19943 , w_19944 , w_19945 , 
		w_19946 , w_19947 , w_19948 , w_19949 , w_19950 , w_19951 , w_19952 , w_19953 , w_19954 , w_19955 , 
		w_19956 , w_19957 , w_19958 , w_19959 , w_19960 , w_19961 , w_19962 , w_19963 , w_19964 , w_19965 , 
		w_19966 , w_19967 , w_19968 , w_19969 , w_19970 , w_19971 , w_19972 , w_19973 , w_19974 , w_19975 , 
		w_19976 , w_19977 , w_19978 , w_19979 , w_19980 , w_19981 , w_19982 , w_19983 , w_19984 , w_19985 , 
		w_19986 , w_19987 , w_19988 , w_19989 , w_19990 , w_19991 , w_19992 , w_19993 , w_19994 , w_19995 , 
		w_19996 , w_19997 , w_19998 , w_19999 , w_20000 , w_20001 , w_20002 , w_20003 , w_20004 , w_20005 , 
		w_20006 , w_20007 , w_20008 , w_20009 , w_20010 , w_20011 , w_20012 , w_20013 , w_20014 , w_20015 , 
		w_20016 , w_20017 , w_20018 , w_20019 , w_20020 , w_20021 , w_20022 , w_20023 , w_20024 , w_20025 , 
		w_20026 , w_20027 , w_20028 , w_20029 , w_20030 , w_20031 , w_20032 , w_20033 , w_20034 , w_20035 , 
		w_20036 , w_20037 , w_20038 , w_20039 , w_20040 , w_20041 , w_20042 , w_20043 , w_20044 , w_20045 , 
		w_20046 , w_20047 , w_20048 , w_20049 , w_20050 , w_20051 , w_20052 , w_20053 , w_20054 , w_20055 , 
		w_20056 , w_20057 , w_20058 , w_20059 , w_20060 , w_20061 , w_20062 , w_20063 , w_20064 , w_20065 , 
		w_20066 , w_20067 , w_20068 , w_20069 , w_20070 , w_20071 , w_20072 , w_20073 , w_20074 , w_20075 , 
		w_20076 , w_20077 , w_20078 , w_20079 , w_20080 , w_20081 , w_20082 , w_20083 , w_20084 , w_20085 , 
		w_20086 , w_20087 , w_20088 , w_20089 , w_20090 , w_20091 , w_20092 , w_20093 , w_20094 , w_20095 , 
		w_20096 , w_20097 , w_20098 , w_20099 , w_20100 , w_20101 , w_20102 , w_20103 , w_20104 , w_20105 , 
		w_20106 , w_20107 , w_20108 , w_20109 , w_20110 , w_20111 , w_20112 , w_20113 , w_20114 , w_20115 , 
		w_20116 , w_20117 , w_20118 , w_20119 , w_20120 , w_20121 , w_20122 , w_20123 , w_20124 , w_20125 , 
		w_20126 , w_20127 , w_20128 , w_20129 , w_20130 , w_20131 , w_20132 , w_20133 , w_20134 , w_20135 , 
		w_20136 , w_20137 , w_20138 , w_20139 , w_20140 , w_20141 , w_20142 , w_20143 , w_20144 , w_20145 , 
		w_20146 , w_20147 , w_20148 , w_20149 , w_20150 , w_20151 , w_20152 , w_20153 , w_20154 , w_20155 , 
		w_20156 , w_20157 , w_20158 , w_20159 , w_20160 , w_20161 , w_20162 , w_20163 , w_20164 , w_20165 , 
		w_20166 , w_20167 , w_20168 , w_20169 , w_20170 , w_20171 , w_20172 , w_20173 , w_20174 , w_20175 , 
		w_20176 , w_20177 , w_20178 , w_20179 , w_20180 , w_20181 , w_20182 , w_20183 , w_20184 , w_20185 , 
		w_20186 , w_20187 , w_20188 , w_20189 , w_20190 , w_20191 , w_20192 , w_20193 , w_20194 , w_20195 , 
		w_20196 , w_20197 , w_20198 , w_20199 , w_20200 , w_20201 , w_20202 , w_20203 , w_20204 , w_20205 , 
		w_20206 , w_20207 , w_20208 , w_20209 , w_20210 , w_20211 , w_20212 , w_20213 , w_20214 , w_20215 , 
		w_20216 , w_20217 , w_20218 , w_20219 , w_20220 , w_20221 , w_20222 , w_20223 , w_20224 , w_20225 , 
		w_20226 , w_20227 , w_20228 , w_20229 , w_20230 , w_20231 , w_20232 , w_20233 , w_20234 , w_20235 , 
		w_20236 , w_20237 , w_20238 , w_20239 , w_20240 , w_20241 , w_20242 , w_20243 , w_20244 , w_20245 , 
		w_20246 , w_20247 , w_20248 , w_20249 , w_20250 , w_20251 , w_20252 , w_20253 , w_20254 , w_20255 , 
		w_20256 , w_20257 , w_20258 , w_20259 , w_20260 , w_20261 , w_20262 , w_20263 , w_20264 , w_20265 , 
		w_20266 , w_20267 , w_20268 , w_20269 , w_20270 , w_20271 , w_20272 , w_20273 , w_20274 , w_20275 , 
		w_20276 , w_20277 , w_20278 , w_20279 , w_20280 , w_20281 , w_20282 , w_20283 , w_20284 , w_20285 , 
		w_20286 , w_20287 , w_20288 , w_20289 , w_20290 , w_20291 , w_20292 , w_20293 , w_20294 , w_20295 , 
		w_20296 , w_20297 , w_20298 , w_20299 , w_20300 , w_20301 , w_20302 , w_20303 , w_20304 , w_20305 , 
		w_20306 , w_20307 , w_20308 , w_20309 , w_20310 , w_20311 , w_20312 , w_20313 , w_20314 , w_20315 , 
		w_20316 , w_20317 , w_20318 , w_20319 , w_20320 , w_20321 , w_20322 , w_20323 , w_20324 , w_20325 , 
		w_20326 , w_20327 , w_20328 , w_20329 , w_20330 , w_20331 , w_20332 , w_20333 , w_20334 , w_20335 , 
		w_20336 , w_20337 , w_20338 , w_20339 , w_20340 , w_20341 , w_20342 , w_20343 , w_20344 , w_20345 , 
		w_20346 , w_20347 , w_20348 , w_20349 , w_20350 , w_20351 , w_20352 , w_20353 , w_20354 , w_20355 , 
		w_20356 , w_20357 , w_20358 , w_20359 , w_20360 , w_20361 , w_20362 , w_20363 , w_20364 , w_20365 , 
		w_20366 , w_20367 , w_20368 , w_20369 , w_20370 , w_20371 , w_20372 , w_20373 , w_20374 , w_20375 , 
		w_20376 , w_20377 , w_20378 , w_20379 , w_20380 , w_20381 , w_20382 , w_20383 , w_20384 , w_20385 , 
		w_20386 , w_20387 , w_20388 , w_20389 , w_20390 , w_20391 , w_20392 , w_20393 , w_20394 , w_20395 , 
		w_20396 , w_20397 , w_20398 , w_20399 , w_20400 , w_20401 , w_20402 , w_20403 , w_20404 , w_20405 , 
		w_20406 , w_20407 , w_20408 , w_20409 , w_20410 , w_20411 , w_20412 , w_20413 , w_20414 , w_20415 , 
		w_20416 , w_20417 , w_20418 , w_20419 , w_20420 , w_20421 , w_20422 , w_20423 , w_20424 , w_20425 , 
		w_20426 , w_20427 , w_20428 , w_20429 , w_20430 , w_20431 , w_20432 , w_20433 , w_20434 , w_20435 , 
		w_20436 , w_20437 , w_20438 , w_20439 , w_20440 , w_20441 , w_20442 , w_20443 , w_20444 , w_20445 , 
		w_20446 , w_20447 , w_20448 , w_20449 , w_20450 , w_20451 , w_20452 , w_20453 , w_20454 , w_20455 , 
		w_20456 , w_20457 , w_20458 , w_20459 , w_20460 , w_20461 , w_20462 , w_20463 , w_20464 , w_20465 , 
		w_20466 , w_20467 , w_20468 , w_20469 , w_20470 , w_20471 , w_20472 , w_20473 , w_20474 , w_20475 , 
		w_20476 , w_20477 , w_20478 , w_20479 , w_20480 , w_20481 , w_20482 , w_20483 , w_20484 , w_20485 , 
		w_20486 , w_20487 , w_20488 , w_20489 , w_20490 , w_20491 , w_20492 , w_20493 , w_20494 , w_20495 , 
		w_20496 , w_20497 , w_20498 , w_20499 , w_20500 , w_20501 , w_20502 , w_20503 , w_20504 , w_20505 , 
		w_20506 , w_20507 , w_20508 , w_20509 , w_20510 , w_20511 , w_20512 , w_20513 , w_20514 , w_20515 , 
		w_20516 , w_20517 , w_20518 , w_20519 , w_20520 , w_20521 , w_20522 , w_20523 , w_20524 , w_20525 , 
		w_20526 , w_20527 , w_20528 , w_20529 , w_20530 , w_20531 , w_20532 , w_20533 , w_20534 , w_20535 , 
		w_20536 , w_20537 , w_20538 , w_20539 , w_20540 , w_20541 , w_20542 , w_20543 , w_20544 , w_20545 , 
		w_20546 , w_20547 , w_20548 , w_20549 , w_20550 , w_20551 , w_20552 , w_20553 , w_20554 , w_20555 , 
		w_20556 , w_20557 , w_20558 , w_20559 , w_20560 , w_20561 , w_20562 , w_20563 , w_20564 , w_20565 , 
		w_20566 , w_20567 , w_20568 , w_20569 , w_20570 , w_20571 , w_20572 , w_20573 , w_20574 , w_20575 , 
		w_20576 , w_20577 , w_20578 , w_20579 , w_20580 , w_20581 , w_20582 , w_20583 , w_20584 , w_20585 , 
		w_20586 , w_20587 , w_20588 , w_20589 , w_20590 , w_20591 , w_20592 , w_20593 , w_20594 , w_20595 , 
		w_20596 , w_20597 , w_20598 , w_20599 , w_20600 , w_20601 , w_20602 , w_20603 , w_20604 , w_20605 , 
		w_20606 , w_20607 , w_20608 , w_20609 , w_20610 , w_20611 , w_20612 , w_20613 , w_20614 , w_20615 , 
		w_20616 , w_20617 , w_20618 , w_20619 , w_20620 , w_20621 , w_20622 , w_20623 , w_20624 , w_20625 , 
		w_20626 , w_20627 , w_20628 , w_20629 , w_20630 , w_20631 , w_20632 , w_20633 , w_20634 , w_20635 , 
		w_20636 , w_20637 , w_20638 , w_20639 , w_20640 , w_20641 , w_20642 , w_20643 , w_20644 , w_20645 , 
		w_20646 , w_20647 , w_20648 , w_20649 , w_20650 , w_20651 , w_20652 , w_20653 , w_20654 , w_20655 , 
		w_20656 , w_20657 , w_20658 , w_20659 , w_20660 , w_20661 , w_20662 , w_20663 , w_20664 , w_20665 , 
		w_20666 , w_20667 , w_20668 , w_20669 , w_20670 , w_20671 , w_20672 , w_20673 , w_20674 , w_20675 , 
		w_20676 , w_20677 , w_20678 , w_20679 , w_20680 , w_20681 , w_20682 , w_20683 , w_20684 , w_20685 , 
		w_20686 , w_20687 , w_20688 , w_20689 , w_20690 , w_20691 , w_20692 , w_20693 , w_20694 , w_20695 , 
		w_20696 , w_20697 , w_20698 , w_20699 , w_20700 , w_20701 , w_20702 , w_20703 , w_20704 , w_20705 , 
		w_20706 , w_20707 , w_20708 , w_20709 , w_20710 , w_20711 , w_20712 , w_20713 , w_20714 , w_20715 , 
		w_20716 , w_20717 , w_20718 , w_20719 , w_20720 , w_20721 , w_20722 , w_20723 , w_20724 , w_20725 , 
		w_20726 , w_20727 , w_20728 , w_20729 , w_20730 , w_20731 , w_20732 , w_20733 , w_20734 , w_20735 , 
		w_20736 , w_20737 , w_20738 , w_20739 , w_20740 , w_20741 , w_20742 , w_20743 , w_20744 , w_20745 , 
		w_20746 , w_20747 , w_20748 , w_20749 , w_20750 , w_20751 , w_20752 , w_20753 , w_20754 , w_20755 , 
		w_20756 , w_20757 , w_20758 , w_20759 , w_20760 , w_20761 , w_20762 , w_20763 , w_20764 , w_20765 , 
		w_20766 , w_20767 , w_20768 , w_20769 , w_20770 , w_20771 , w_20772 , w_20773 , w_20774 , w_20775 , 
		w_20776 , w_20777 , w_20778 , w_20779 , w_20780 , w_20781 , w_20782 , w_20783 , w_20784 , w_20785 , 
		w_20786 , w_20787 , w_20788 , w_20789 , w_20790 , w_20791 , w_20792 , w_20793 , w_20794 , w_20795 , 
		w_20796 , w_20797 , w_20798 , w_20799 , w_20800 , w_20801 , w_20802 , w_20803 , w_20804 , w_20805 , 
		w_20806 , w_20807 , w_20808 , w_20809 , w_20810 , w_20811 , w_20812 , w_20813 , w_20814 , w_20815 , 
		w_20816 , w_20817 , w_20818 , w_20819 , w_20820 , w_20821 , w_20822 , w_20823 , w_20824 , w_20825 , 
		w_20826 , w_20827 , w_20828 , w_20829 , w_20830 , w_20831 , w_20832 , w_20833 , w_20834 , w_20835 , 
		w_20836 , w_20837 , w_20838 , w_20839 , w_20840 , w_20841 , w_20842 , w_20843 , w_20844 , w_20845 , 
		w_20846 , w_20847 , w_20848 , w_20849 , w_20850 , w_20851 , w_20852 , w_20853 , w_20854 , w_20855 , 
		w_20856 , w_20857 , w_20858 , w_20859 , w_20860 , w_20861 , w_20862 , w_20863 , w_20864 , w_20865 , 
		w_20866 , w_20867 , w_20868 , w_20869 , w_20870 , w_20871 , w_20872 , w_20873 , w_20874 , w_20875 , 
		w_20876 , w_20877 , w_20878 , w_20879 , w_20880 , w_20881 , w_20882 , w_20883 , w_20884 , w_20885 , 
		w_20886 , w_20887 , w_20888 , w_20889 , w_20890 , w_20891 , w_20892 , w_20893 , w_20894 , w_20895 , 
		w_20896 , w_20897 , w_20898 , w_20899 , w_20900 , w_20901 , w_20902 , w_20903 , w_20904 , w_20905 , 
		w_20906 , w_20907 , w_20908 , w_20909 , w_20910 , w_20911 , w_20912 , w_20913 , w_20914 , w_20915 , 
		w_20916 , w_20917 , w_20918 , w_20919 , w_20920 , w_20921 , w_20922 , w_20923 , w_20924 , w_20925 , 
		w_20926 , w_20927 , w_20928 , w_20929 , w_20930 , w_20931 , w_20932 , w_20933 , w_20934 , w_20935 , 
		w_20936 , w_20937 , w_20938 , w_20939 , w_20940 , w_20941 , w_20942 , w_20943 , w_20944 , w_20945 , 
		w_20946 , w_20947 , w_20948 , w_20949 , w_20950 , w_20951 , w_20952 , w_20953 , w_20954 , w_20955 , 
		w_20956 , w_20957 , w_20958 , w_20959 , w_20960 , w_20961 , w_20962 , w_20963 , w_20964 , w_20965 , 
		w_20966 , w_20967 , w_20968 , w_20969 , w_20970 , w_20971 , w_20972 , w_20973 , w_20974 , w_20975 , 
		w_20976 , w_20977 , w_20978 , w_20979 , w_20980 , w_20981 , w_20982 , w_20983 , w_20984 , w_20985 , 
		w_20986 , w_20987 , w_20988 , w_20989 , w_20990 , w_20991 , w_20992 , w_20993 , w_20994 , w_20995 , 
		w_20996 , w_20997 , w_20998 , w_20999 , w_21000 , w_21001 , w_21002 , w_21003 , w_21004 , w_21005 , 
		w_21006 , w_21007 , w_21008 , w_21009 , w_21010 , w_21011 , w_21012 , w_21013 , w_21014 , w_21015 , 
		w_21016 , w_21017 , w_21018 , w_21019 , w_21020 , w_21021 , w_21022 , w_21023 , w_21024 , w_21025 , 
		w_21026 , w_21027 , w_21028 , w_21029 , w_21030 , w_21031 , w_21032 , w_21033 , w_21034 , w_21035 , 
		w_21036 , w_21037 , w_21038 , w_21039 , w_21040 , w_21041 , w_21042 , w_21043 , w_21044 , w_21045 , 
		w_21046 , w_21047 , w_21048 , w_21049 , w_21050 , w_21051 , w_21052 , w_21053 , w_21054 , w_21055 , 
		w_21056 , w_21057 , w_21058 , w_21059 , w_21060 , w_21061 , w_21062 , w_21063 , w_21064 , w_21065 , 
		w_21066 , w_21067 , w_21068 , w_21069 , w_21070 , w_21071 , w_21072 , w_21073 , w_21074 , w_21075 , 
		w_21076 , w_21077 , w_21078 , w_21079 , w_21080 , w_21081 , w_21082 , w_21083 , w_21084 , w_21085 , 
		w_21086 , w_21087 , w_21088 , w_21089 , w_21090 , w_21091 , w_21092 , w_21093 , w_21094 , w_21095 , 
		w_21096 , w_21097 , w_21098 , w_21099 , w_21100 , w_21101 , w_21102 , w_21103 , w_21104 , w_21105 , 
		w_21106 , w_21107 , w_21108 , w_21109 , w_21110 , w_21111 , w_21112 , w_21113 , w_21114 , w_21115 , 
		w_21116 , w_21117 , w_21118 , w_21119 , w_21120 , w_21121 , w_21122 , w_21123 , w_21124 , w_21125 , 
		w_21126 , w_21127 , w_21128 , w_21129 , w_21130 , w_21131 , w_21132 , w_21133 , w_21134 , w_21135 , 
		w_21136 , w_21137 , w_21138 , w_21139 , w_21140 , w_21141 , w_21142 , w_21143 , w_21144 , w_21145 , 
		w_21146 , w_21147 , w_21148 , w_21149 , w_21150 , w_21151 , w_21152 , w_21153 , w_21154 , w_21155 , 
		w_21156 , w_21157 , w_21158 , w_21159 , w_21160 , w_21161 , w_21162 , w_21163 , w_21164 , w_21165 , 
		w_21166 , w_21167 , w_21168 , w_21169 , w_21170 , w_21171 , w_21172 , w_21173 , w_21174 , w_21175 , 
		w_21176 , w_21177 , w_21178 , w_21179 , w_21180 , w_21181 , w_21182 , w_21183 , w_21184 , w_21185 , 
		w_21186 , w_21187 , w_21188 , w_21189 , w_21190 , w_21191 , w_21192 , w_21193 , w_21194 , w_21195 , 
		w_21196 , w_21197 , w_21198 , w_21199 , w_21200 , w_21201 , w_21202 , w_21203 , w_21204 , w_21205 , 
		w_21206 , w_21207 , w_21208 , w_21209 , w_21210 , w_21211 , w_21212 , w_21213 , w_21214 , w_21215 , 
		w_21216 , w_21217 , w_21218 , w_21219 , w_21220 , w_21221 , w_21222 , w_21223 , w_21224 , w_21225 , 
		w_21226 , w_21227 , w_21228 , w_21229 , w_21230 , w_21231 , w_21232 , w_21233 , w_21234 , w_21235 , 
		w_21236 , w_21237 , w_21238 , w_21239 , w_21240 , w_21241 , w_21242 , w_21243 , w_21244 , w_21245 , 
		w_21246 , w_21247 , w_21248 , w_21249 , w_21250 , w_21251 , w_21252 , w_21253 , w_21254 , w_21255 , 
		w_21256 , w_21257 , w_21258 , w_21259 , w_21260 , w_21261 , w_21262 , w_21263 , w_21264 , w_21265 , 
		w_21266 , w_21267 , w_21268 , w_21269 , w_21270 , w_21271 , w_21272 , w_21273 , w_21274 , w_21275 , 
		w_21276 , w_21277 , w_21278 , w_21279 , w_21280 , w_21281 , w_21282 , w_21283 , w_21284 , w_21285 , 
		w_21286 , w_21287 , w_21288 , w_21289 , w_21290 , w_21291 , w_21292 , w_21293 , w_21294 , w_21295 , 
		w_21296 , w_21297 , w_21298 , w_21299 , w_21300 , w_21301 , w_21302 , w_21303 , w_21304 , w_21305 , 
		w_21306 , w_21307 , w_21308 , w_21309 , w_21310 , w_21311 , w_21312 , w_21313 , w_21314 , w_21315 , 
		w_21316 , w_21317 , w_21318 , w_21319 , w_21320 , w_21321 , w_21322 , w_21323 , w_21324 , w_21325 , 
		w_21326 , w_21327 , w_21328 , w_21329 , w_21330 , w_21331 , w_21332 , w_21333 , w_21334 , w_21335 , 
		w_21336 , w_21337 , w_21338 , w_21339 , w_21340 , w_21341 , w_21342 , w_21343 , w_21344 , w_21345 , 
		w_21346 , w_21347 , w_21348 , w_21349 , w_21350 , w_21351 , w_21352 , w_21353 , w_21354 , w_21355 , 
		w_21356 , w_21357 , w_21358 , w_21359 , w_21360 , w_21361 , w_21362 , w_21363 , w_21364 , w_21365 , 
		w_21366 , w_21367 , w_21368 , w_21369 , w_21370 , w_21371 , w_21372 , w_21373 , w_21374 , w_21375 , 
		w_21376 , w_21377 , w_21378 , w_21379 , w_21380 , w_21381 , w_21382 , w_21383 , w_21384 , w_21385 , 
		w_21386 , w_21387 , w_21388 , w_21389 , w_21390 , w_21391 , w_21392 , w_21393 , w_21394 , w_21395 , 
		w_21396 , w_21397 , w_21398 , w_21399 , w_21400 , w_21401 , w_21402 , w_21403 , w_21404 , w_21405 , 
		w_21406 , w_21407 , w_21408 , w_21409 , w_21410 , w_21411 , w_21412 , w_21413 , w_21414 , w_21415 , 
		w_21416 , w_21417 , w_21418 , w_21419 , w_21420 , w_21421 , w_21422 , w_21423 , w_21424 , w_21425 , 
		w_21426 , w_21427 , w_21428 , w_21429 , w_21430 , w_21431 , w_21432 , w_21433 , w_21434 , w_21435 , 
		w_21436 , w_21437 , w_21438 , w_21439 , w_21440 , w_21441 , w_21442 , w_21443 , w_21444 , w_21445 , 
		w_21446 , w_21447 , w_21448 , w_21449 , w_21450 , w_21451 , w_21452 , w_21453 , w_21454 , w_21455 , 
		w_21456 , w_21457 , w_21458 , w_21459 , w_21460 , w_21461 , w_21462 , w_21463 , w_21464 , w_21465 , 
		w_21466 , w_21467 , w_21468 , w_21469 , w_21470 , w_21471 , w_21472 , w_21473 , w_21474 , w_21475 , 
		w_21476 , w_21477 , w_21478 , w_21479 , w_21480 , w_21481 , w_21482 , w_21483 , w_21484 , w_21485 , 
		w_21486 , w_21487 , w_21488 , w_21489 , w_21490 , w_21491 , w_21492 , w_21493 , w_21494 , w_21495 , 
		w_21496 , w_21497 , w_21498 , w_21499 , w_21500 , w_21501 , w_21502 , w_21503 , w_21504 , w_21505 , 
		w_21506 , w_21507 , w_21508 , w_21509 , w_21510 , w_21511 , w_21512 , w_21513 , w_21514 , w_21515 , 
		w_21516 , w_21517 , w_21518 , w_21519 , w_21520 , w_21521 , w_21522 , w_21523 , w_21524 , w_21525 , 
		w_21526 , w_21527 , w_21528 , w_21529 , w_21530 , w_21531 , w_21532 , w_21533 , w_21534 , w_21535 , 
		w_21536 , w_21537 , w_21538 , w_21539 , w_21540 , w_21541 , w_21542 , w_21543 , w_21544 , w_21545 , 
		w_21546 , w_21547 , w_21548 , w_21549 , w_21550 , w_21551 , w_21552 , w_21553 , w_21554 , w_21555 , 
		w_21556 , w_21557 , w_21558 , w_21559 , w_21560 , w_21561 , w_21562 , w_21563 , w_21564 , w_21565 , 
		w_21566 , w_21567 , w_21568 , w_21569 , w_21570 , w_21571 , w_21572 , w_21573 , w_21574 , w_21575 , 
		w_21576 , w_21577 , w_21578 , w_21579 , w_21580 , w_21581 , w_21582 , w_21583 , w_21584 , w_21585 , 
		w_21586 , w_21587 , w_21588 , w_21589 , w_21590 , w_21591 , w_21592 , w_21593 , w_21594 , w_21595 , 
		w_21596 , w_21597 , w_21598 , w_21599 , w_21600 , w_21601 , w_21602 , w_21603 , w_21604 , w_21605 , 
		w_21606 , w_21607 , w_21608 , w_21609 , w_21610 , w_21611 , w_21612 , w_21613 , w_21614 , w_21615 , 
		w_21616 , w_21617 , w_21618 , w_21619 , w_21620 , w_21621 , w_21622 , w_21623 , w_21624 , w_21625 , 
		w_21626 , w_21627 , w_21628 , w_21629 , w_21630 , w_21631 , w_21632 , w_21633 , w_21634 , w_21635 , 
		w_21636 , w_21637 , w_21638 , w_21639 , w_21640 , w_21641 , w_21642 , w_21643 , w_21644 , w_21645 , 
		w_21646 , w_21647 , w_21648 , w_21649 , w_21650 , w_21651 , w_21652 , w_21653 , w_21654 , w_21655 , 
		w_21656 , w_21657 , w_21658 , w_21659 , w_21660 , w_21661 , w_21662 , w_21663 , w_21664 , w_21665 , 
		w_21666 , w_21667 , w_21668 , w_21669 , w_21670 , w_21671 , w_21672 , w_21673 , w_21674 , w_21675 , 
		w_21676 , w_21677 , w_21678 , w_21679 , w_21680 , w_21681 , w_21682 , w_21683 , w_21684 , w_21685 , 
		w_21686 , w_21687 , w_21688 , w_21689 , w_21690 , w_21691 , w_21692 , w_21693 , w_21694 , w_21695 , 
		w_21696 , w_21697 , w_21698 , w_21699 , w_21700 , w_21701 , w_21702 , w_21703 , w_21704 , w_21705 , 
		w_21706 , w_21707 , w_21708 , w_21709 , w_21710 , w_21711 , w_21712 , w_21713 , w_21714 , w_21715 , 
		w_21716 , w_21717 , w_21718 , w_21719 , w_21720 , w_21721 , w_21722 , w_21723 , w_21724 , w_21725 , 
		w_21726 , w_21727 , w_21728 , w_21729 , w_21730 , w_21731 , w_21732 , w_21733 , w_21734 , w_21735 , 
		w_21736 , w_21737 , w_21738 , w_21739 , w_21740 , w_21741 , w_21742 , w_21743 , w_21744 , w_21745 , 
		w_21746 , w_21747 , w_21748 , w_21749 , w_21750 , w_21751 , w_21752 , w_21753 , w_21754 , w_21755 , 
		w_21756 , w_21757 , w_21758 , w_21759 , w_21760 , w_21761 , w_21762 , w_21763 , w_21764 , w_21765 , 
		w_21766 , w_21767 , w_21768 , w_21769 , w_21770 , w_21771 , w_21772 , w_21773 , w_21774 , w_21775 , 
		w_21776 , w_21777 , w_21778 , w_21779 , w_21780 , w_21781 , w_21782 , w_21783 , w_21784 , w_21785 , 
		w_21786 , w_21787 , w_21788 , w_21789 , w_21790 , w_21791 , w_21792 , w_21793 , w_21794 , w_21795 , 
		w_21796 , w_21797 , w_21798 , w_21799 , w_21800 , w_21801 , w_21802 , w_21803 , w_21804 , w_21805 , 
		w_21806 , w_21807 , w_21808 , w_21809 , w_21810 , w_21811 , w_21812 , w_21813 , w_21814 , w_21815 , 
		w_21816 , w_21817 , w_21818 , w_21819 , w_21820 , w_21821 , w_21822 , w_21823 , w_21824 , w_21825 , 
		w_21826 , w_21827 , w_21828 , w_21829 , w_21830 , w_21831 , w_21832 , w_21833 , w_21834 , w_21835 , 
		w_21836 , w_21837 , w_21838 , w_21839 , w_21840 , w_21841 , w_21842 , w_21843 , w_21844 , w_21845 , 
		w_21846 , w_21847 , w_21848 , w_21849 , w_21850 , w_21851 , w_21852 , w_21853 , w_21854 , w_21855 , 
		w_21856 , w_21857 , w_21858 , w_21859 , w_21860 , w_21861 , w_21862 , w_21863 , w_21864 , w_21865 , 
		w_21866 , w_21867 , w_21868 , w_21869 , w_21870 , w_21871 , w_21872 , w_21873 , w_21874 , w_21875 , 
		w_21876 , w_21877 , w_21878 , w_21879 , w_21880 , w_21881 , w_21882 , w_21883 , w_21884 , w_21885 , 
		w_21886 , w_21887 , w_21888 , w_21889 , w_21890 , w_21891 , w_21892 , w_21893 , w_21894 , w_21895 , 
		w_21896 , w_21897 , w_21898 , w_21899 , w_21900 , w_21901 , w_21902 , w_21903 , w_21904 , w_21905 , 
		w_21906 , w_21907 , w_21908 , w_21909 , w_21910 , w_21911 , w_21912 , w_21913 , w_21914 , w_21915 , 
		w_21916 , w_21917 , w_21918 , w_21919 , w_21920 , w_21921 , w_21922 , w_21923 , w_21924 , w_21925 , 
		w_21926 , w_21927 , w_21928 , w_21929 , w_21930 , w_21931 , w_21932 , w_21933 , w_21934 , w_21935 , 
		w_21936 , w_21937 , w_21938 , w_21939 , w_21940 , w_21941 , w_21942 , w_21943 , w_21944 , w_21945 , 
		w_21946 , w_21947 , w_21948 , w_21949 , w_21950 , w_21951 , w_21952 , w_21953 , w_21954 , w_21955 , 
		w_21956 , w_21957 , w_21958 , w_21959 , w_21960 , w_21961 , w_21962 , w_21963 , w_21964 , w_21965 , 
		w_21966 , w_21967 , w_21968 , w_21969 , w_21970 , w_21971 , w_21972 , w_21973 , w_21974 , w_21975 , 
		w_21976 , w_21977 , w_21978 , w_21979 , w_21980 , w_21981 , w_21982 , w_21983 , w_21984 , w_21985 , 
		w_21986 , w_21987 , w_21988 , w_21989 , w_21990 , w_21991 , w_21992 , w_21993 , w_21994 , w_21995 , 
		w_21996 , w_21997 , w_21998 , w_21999 , w_22000 , w_22001 , w_22002 , w_22003 , w_22004 , w_22005 , 
		w_22006 , w_22007 , w_22008 , w_22009 , w_22010 , w_22011 , w_22012 , w_22013 , w_22014 , w_22015 , 
		w_22016 , w_22017 , w_22018 , w_22019 , w_22020 , w_22021 , w_22022 , w_22023 , w_22024 , w_22025 , 
		w_22026 , w_22027 , w_22028 , w_22029 , w_22030 , w_22031 , w_22032 , w_22033 , w_22034 , w_22035 , 
		w_22036 , w_22037 , w_22038 , w_22039 , w_22040 , w_22041 , w_22042 , w_22043 , w_22044 , w_22045 , 
		w_22046 , w_22047 , w_22048 , w_22049 , w_22050 , w_22051 , w_22052 , w_22053 , w_22054 , w_22055 , 
		w_22056 , w_22057 , w_22058 , w_22059 , w_22060 , w_22061 , w_22062 , w_22063 , w_22064 , w_22065 , 
		w_22066 , w_22067 , w_22068 , w_22069 , w_22070 , w_22071 , w_22072 , w_22073 , w_22074 , w_22075 , 
		w_22076 , w_22077 , w_22078 , w_22079 , w_22080 , w_22081 , w_22082 , w_22083 , w_22084 , w_22085 , 
		w_22086 , w_22087 , w_22088 , w_22089 , w_22090 , w_22091 , w_22092 , w_22093 , w_22094 , w_22095 , 
		w_22096 , w_22097 , w_22098 , w_22099 , w_22100 , w_22101 , w_22102 , w_22103 , w_22104 , w_22105 , 
		w_22106 , w_22107 , w_22108 , w_22109 , w_22110 , w_22111 , w_22112 , w_22113 , w_22114 , w_22115 , 
		w_22116 , w_22117 , w_22118 , w_22119 , w_22120 , w_22121 , w_22122 , w_22123 , w_22124 , w_22125 , 
		w_22126 , w_22127 , w_22128 , w_22129 , w_22130 , w_22131 , w_22132 , w_22133 , w_22134 , w_22135 , 
		w_22136 , w_22137 , w_22138 , w_22139 , w_22140 , w_22141 , w_22142 , w_22143 , w_22144 , w_22145 , 
		w_22146 , w_22147 , w_22148 , w_22149 , w_22150 , w_22151 , w_22152 , w_22153 , w_22154 , w_22155 , 
		w_22156 , w_22157 , w_22158 , w_22159 , w_22160 , w_22161 , w_22162 , w_22163 , w_22164 , w_22165 , 
		w_22166 , w_22167 , w_22168 , w_22169 , w_22170 , w_22171 , w_22172 , w_22173 , w_22174 , w_22175 , 
		w_22176 , w_22177 , w_22178 , w_22179 , w_22180 , w_22181 , w_22182 , w_22183 , w_22184 , w_22185 , 
		w_22186 , w_22187 , w_22188 , w_22189 , w_22190 , w_22191 , w_22192 , w_22193 , w_22194 , w_22195 , 
		w_22196 , w_22197 , w_22198 , w_22199 , w_22200 , w_22201 , w_22202 , w_22203 , w_22204 , w_22205 , 
		w_22206 , w_22207 , w_22208 , w_22209 , w_22210 , w_22211 , w_22212 , w_22213 , w_22214 , w_22215 , 
		w_22216 , w_22217 , w_22218 , w_22219 , w_22220 , w_22221 , w_22222 , w_22223 , w_22224 , w_22225 , 
		w_22226 , w_22227 , w_22228 , w_22229 , w_22230 , w_22231 , w_22232 , w_22233 , w_22234 , w_22235 , 
		w_22236 , w_22237 , w_22238 , w_22239 , w_22240 , w_22241 , w_22242 , w_22243 , w_22244 , w_22245 , 
		w_22246 , w_22247 , w_22248 , w_22249 , w_22250 , w_22251 , w_22252 , w_22253 , w_22254 , w_22255 , 
		w_22256 , w_22257 , w_22258 , w_22259 , w_22260 , w_22261 , w_22262 , w_22263 , w_22264 , w_22265 , 
		w_22266 , w_22267 , w_22268 , w_22269 , w_22270 , w_22271 , w_22272 , w_22273 , w_22274 , w_22275 , 
		w_22276 , w_22277 , w_22278 , w_22279 , w_22280 , w_22281 , w_22282 , w_22283 , w_22284 , w_22285 , 
		w_22286 , w_22287 , w_22288 , w_22289 , w_22290 , w_22291 , w_22292 , w_22293 , w_22294 , w_22295 , 
		w_22296 , w_22297 , w_22298 , w_22299 , w_22300 , w_22301 , w_22302 , w_22303 , w_22304 , w_22305 , 
		w_22306 , w_22307 , w_22308 , w_22309 , w_22310 , w_22311 , w_22312 , w_22313 , w_22314 , w_22315 , 
		w_22316 , w_22317 , w_22318 , w_22319 , w_22320 , w_22321 , w_22322 , w_22323 , w_22324 , w_22325 , 
		w_22326 , w_22327 , w_22328 , w_22329 , w_22330 , w_22331 , w_22332 , w_22333 , w_22334 , w_22335 , 
		w_22336 , w_22337 , w_22338 , w_22339 , w_22340 , w_22341 , w_22342 , w_22343 , w_22344 , w_22345 , 
		w_22346 , w_22347 , w_22348 , w_22349 , w_22350 , w_22351 , w_22352 , w_22353 , w_22354 , w_22355 , 
		w_22356 , w_22357 , w_22358 , w_22359 , w_22360 , w_22361 , w_22362 , w_22363 , w_22364 , w_22365 , 
		w_22366 , w_22367 , w_22368 , w_22369 , w_22370 , w_22371 , w_22372 , w_22373 , w_22374 , w_22375 , 
		w_22376 , w_22377 , w_22378 , w_22379 , w_22380 , w_22381 , w_22382 , w_22383 , w_22384 , w_22385 , 
		w_22386 , w_22387 , w_22388 , w_22389 , w_22390 , w_22391 , w_22392 , w_22393 , w_22394 , w_22395 , 
		w_22396 , w_22397 , w_22398 , w_22399 , w_22400 , w_22401 , w_22402 , w_22403 , w_22404 , w_22405 , 
		w_22406 , w_22407 , w_22408 , w_22409 , w_22410 , w_22411 , w_22412 , w_22413 , w_22414 , w_22415 , 
		w_22416 , w_22417 , w_22418 , w_22419 , w_22420 , w_22421 , w_22422 , w_22423 , w_22424 , w_22425 , 
		w_22426 , w_22427 , w_22428 , w_22429 , w_22430 , w_22431 , w_22432 , w_22433 , w_22434 , w_22435 , 
		w_22436 , w_22437 , w_22438 , w_22439 , w_22440 , w_22441 , w_22442 , w_22443 , w_22444 , w_22445 , 
		w_22446 , w_22447 , w_22448 , w_22449 , w_22450 , w_22451 , w_22452 , w_22453 , w_22454 , w_22455 , 
		w_22456 , w_22457 , w_22458 , w_22459 , w_22460 , w_22461 , w_22462 , w_22463 , w_22464 , w_22465 , 
		w_22466 , w_22467 , w_22468 , w_22469 , w_22470 , w_22471 , w_22472 , w_22473 , w_22474 , w_22475 , 
		w_22476 , w_22477 , w_22478 , w_22479 , w_22480 , w_22481 , w_22482 , w_22483 , w_22484 , w_22485 , 
		w_22486 , w_22487 , w_22488 , w_22489 , w_22490 , w_22491 , w_22492 , w_22493 , w_22494 , w_22495 , 
		w_22496 , w_22497 , w_22498 , w_22499 , w_22500 , w_22501 , w_22502 , w_22503 , w_22504 , w_22505 , 
		w_22506 , w_22507 , w_22508 , w_22509 , w_22510 , w_22511 , w_22512 , w_22513 , w_22514 , w_22515 , 
		w_22516 , w_22517 , w_22518 , w_22519 , w_22520 , w_22521 , w_22522 , w_22523 , w_22524 , w_22525 , 
		w_22526 , w_22527 , w_22528 , w_22529 , w_22530 , w_22531 , w_22532 , w_22533 , w_22534 , w_22535 , 
		w_22536 , w_22537 , w_22538 , w_22539 , w_22540 , w_22541 , w_22542 , w_22543 , w_22544 , w_22545 , 
		w_22546 , w_22547 , w_22548 , w_22549 , w_22550 , w_22551 , w_22552 , w_22553 , w_22554 , w_22555 , 
		w_22556 , w_22557 , w_22558 , w_22559 , w_22560 , w_22561 , w_22562 , w_22563 , w_22564 , w_22565 , 
		w_22566 , w_22567 , w_22568 , w_22569 , w_22570 , w_22571 , w_22572 , w_22573 , w_22574 , w_22575 , 
		w_22576 , w_22577 , w_22578 , w_22579 , w_22580 , w_22581 , w_22582 , w_22583 , w_22584 , w_22585 , 
		w_22586 , w_22587 , w_22588 , w_22589 , w_22590 , w_22591 , w_22592 , w_22593 , w_22594 , w_22595 , 
		w_22596 , w_22597 , w_22598 , w_22599 , w_22600 , w_22601 , w_22602 , w_22603 , w_22604 , w_22605 , 
		w_22606 , w_22607 , w_22608 , w_22609 , w_22610 , w_22611 , w_22612 , w_22613 , w_22614 , w_22615 , 
		w_22616 , w_22617 , w_22618 , w_22619 , w_22620 , w_22621 , w_22622 , w_22623 , w_22624 , w_22625 , 
		w_22626 , w_22627 , w_22628 , w_22629 , w_22630 , w_22631 , w_22632 , w_22633 , w_22634 , w_22635 , 
		w_22636 , w_22637 , w_22638 , w_22639 , w_22640 , w_22641 , w_22642 , w_22643 , w_22644 , w_22645 , 
		w_22646 , w_22647 , w_22648 , w_22649 , w_22650 , w_22651 , w_22652 , w_22653 , w_22654 , w_22655 , 
		w_22656 , w_22657 , w_22658 , w_22659 , w_22660 , w_22661 , w_22662 , w_22663 , w_22664 , w_22665 , 
		w_22666 , w_22667 , w_22668 , w_22669 , w_22670 , w_22671 , w_22672 , w_22673 , w_22674 , w_22675 , 
		w_22676 , w_22677 , w_22678 , w_22679 , w_22680 , w_22681 , w_22682 , w_22683 , w_22684 , w_22685 , 
		w_22686 , w_22687 , w_22688 , w_22689 , w_22690 , w_22691 , w_22692 , w_22693 , w_22694 , w_22695 , 
		w_22696 , w_22697 , w_22698 , w_22699 , w_22700 , w_22701 , w_22702 , w_22703 , w_22704 , w_22705 , 
		w_22706 , w_22707 , w_22708 , w_22709 , w_22710 , w_22711 , w_22712 , w_22713 , w_22714 , w_22715 , 
		w_22716 , w_22717 , w_22718 , w_22719 , w_22720 , w_22721 , w_22722 , w_22723 , w_22724 , w_22725 , 
		w_22726 , w_22727 , w_22728 , w_22729 , w_22730 , w_22731 , w_22732 , w_22733 , w_22734 , w_22735 , 
		w_22736 , w_22737 , w_22738 , w_22739 , w_22740 , w_22741 , w_22742 , w_22743 , w_22744 , w_22745 , 
		w_22746 , w_22747 , w_22748 , w_22749 , w_22750 , w_22751 , w_22752 , w_22753 , w_22754 , w_22755 , 
		w_22756 , w_22757 , w_22758 , w_22759 , w_22760 , w_22761 , w_22762 , w_22763 , w_22764 , w_22765 , 
		w_22766 , w_22767 , w_22768 , w_22769 , w_22770 , w_22771 , w_22772 , w_22773 , w_22774 , w_22775 , 
		w_22776 , w_22777 , w_22778 , w_22779 , w_22780 , w_22781 , w_22782 , w_22783 , w_22784 , w_22785 , 
		w_22786 , w_22787 , w_22788 , w_22789 , w_22790 , w_22791 , w_22792 , w_22793 , w_22794 , w_22795 , 
		w_22796 , w_22797 , w_22798 , w_22799 , w_22800 , w_22801 , w_22802 , w_22803 , w_22804 , w_22805 , 
		w_22806 , w_22807 , w_22808 , w_22809 , w_22810 , w_22811 , w_22812 , w_22813 , w_22814 , w_22815 , 
		w_22816 , w_22817 , w_22818 , w_22819 , w_22820 , w_22821 , w_22822 , w_22823 , w_22824 , w_22825 , 
		w_22826 , w_22827 , w_22828 , w_22829 , w_22830 , w_22831 , w_22832 , w_22833 , w_22834 , w_22835 , 
		w_22836 , w_22837 , w_22838 , w_22839 , w_22840 , w_22841 , w_22842 , w_22843 , w_22844 , w_22845 , 
		w_22846 , w_22847 , w_22848 , w_22849 , w_22850 , w_22851 , w_22852 , w_22853 , w_22854 , w_22855 , 
		w_22856 , w_22857 , w_22858 , w_22859 , w_22860 , w_22861 , w_22862 , w_22863 , w_22864 , w_22865 , 
		w_22866 , w_22867 , w_22868 , w_22869 , w_22870 , w_22871 , w_22872 , w_22873 , w_22874 , w_22875 , 
		w_22876 , w_22877 , w_22878 , w_22879 , w_22880 , w_22881 , w_22882 , w_22883 , w_22884 , w_22885 , 
		w_22886 , w_22887 , w_22888 , w_22889 , w_22890 , w_22891 , w_22892 , w_22893 , w_22894 , w_22895 , 
		w_22896 , w_22897 , w_22898 , w_22899 , w_22900 , w_22901 , w_22902 , w_22903 , w_22904 , w_22905 , 
		w_22906 , w_22907 , w_22908 , w_22909 , w_22910 , w_22911 , w_22912 , w_22913 , w_22914 , w_22915 , 
		w_22916 , w_22917 , w_22918 , w_22919 , w_22920 , w_22921 , w_22922 , w_22923 , w_22924 , w_22925 , 
		w_22926 , w_22927 , w_22928 , w_22929 , w_22930 , w_22931 , w_22932 , w_22933 , w_22934 , w_22935 , 
		w_22936 , w_22937 , w_22938 , w_22939 , w_22940 , w_22941 , w_22942 , w_22943 , w_22944 , w_22945 , 
		w_22946 , w_22947 , w_22948 , w_22949 , w_22950 , w_22951 , w_22952 , w_22953 , w_22954 , w_22955 , 
		w_22956 , w_22957 , w_22958 , w_22959 , w_22960 , w_22961 , w_22962 , w_22963 , w_22964 , w_22965 , 
		w_22966 , w_22967 , w_22968 , w_22969 , w_22970 , w_22971 , w_22972 , w_22973 , w_22974 , w_22975 , 
		w_22976 , w_22977 , w_22978 , w_22979 , w_22980 , w_22981 , w_22982 , w_22983 , w_22984 , w_22985 , 
		w_22986 , w_22987 , w_22988 , w_22989 , w_22990 , w_22991 , w_22992 , w_22993 , w_22994 , w_22995 , 
		w_22996 , w_22997 , w_22998 , w_22999 , w_23000 , w_23001 , w_23002 , w_23003 , w_23004 , w_23005 , 
		w_23006 , w_23007 , w_23008 , w_23009 , w_23010 , w_23011 , w_23012 , w_23013 , w_23014 , w_23015 , 
		w_23016 , w_23017 , w_23018 , w_23019 , w_23020 , w_23021 , w_23022 , w_23023 , w_23024 , w_23025 , 
		w_23026 , w_23027 , w_23028 , w_23029 , w_23030 , w_23031 , w_23032 , w_23033 , w_23034 , w_23035 , 
		w_23036 , w_23037 , w_23038 , w_23039 , w_23040 , w_23041 , w_23042 , w_23043 , w_23044 , w_23045 , 
		w_23046 , w_23047 , w_23048 , w_23049 , w_23050 , w_23051 , w_23052 , w_23053 , w_23054 , w_23055 , 
		w_23056 , w_23057 , w_23058 , w_23059 , w_23060 , w_23061 , w_23062 , w_23063 , w_23064 , w_23065 , 
		w_23066 , w_23067 , w_23068 , w_23069 , w_23070 , w_23071 , w_23072 , w_23073 , w_23074 , w_23075 , 
		w_23076 , w_23077 , w_23078 , w_23079 , w_23080 , w_23081 , w_23082 , w_23083 , w_23084 , w_23085 , 
		w_23086 , w_23087 , w_23088 , w_23089 , w_23090 , w_23091 , w_23092 , w_23093 , w_23094 , w_23095 , 
		w_23096 , w_23097 , w_23098 , w_23099 , w_23100 , w_23101 , w_23102 , w_23103 , w_23104 , w_23105 , 
		w_23106 , w_23107 , w_23108 , w_23109 , w_23110 , w_23111 , w_23112 , w_23113 , w_23114 , w_23115 , 
		w_23116 , w_23117 , w_23118 , w_23119 , w_23120 , w_23121 , w_23122 , w_23123 , w_23124 , w_23125 , 
		w_23126 , w_23127 , w_23128 , w_23129 , w_23130 , w_23131 , w_23132 , w_23133 , w_23134 , w_23135 , 
		w_23136 , w_23137 , w_23138 , w_23139 , w_23140 , w_23141 , w_23142 , w_23143 , w_23144 , w_23145 , 
		w_23146 , w_23147 , w_23148 , w_23149 , w_23150 , w_23151 , w_23152 , w_23153 , w_23154 , w_23155 , 
		w_23156 , w_23157 , w_23158 , w_23159 , w_23160 , w_23161 , w_23162 , w_23163 , w_23164 , w_23165 , 
		w_23166 , w_23167 , w_23168 , w_23169 , w_23170 , w_23171 , w_23172 , w_23173 , w_23174 , w_23175 , 
		w_23176 , w_23177 , w_23178 , w_23179 , w_23180 , w_23181 , w_23182 , w_23183 , w_23184 , w_23185 , 
		w_23186 , w_23187 , w_23188 , w_23189 , w_23190 , w_23191 , w_23192 , w_23193 , w_23194 , w_23195 , 
		w_23196 , w_23197 , w_23198 , w_23199 , w_23200 , w_23201 , w_23202 , w_23203 , w_23204 , w_23205 , 
		w_23206 , w_23207 , w_23208 , w_23209 , w_23210 , w_23211 , w_23212 , w_23213 , w_23214 , w_23215 , 
		w_23216 , w_23217 , w_23218 , w_23219 , w_23220 , w_23221 , w_23222 , w_23223 , w_23224 , w_23225 , 
		w_23226 , w_23227 , w_23228 , w_23229 , w_23230 , w_23231 , w_23232 , w_23233 , w_23234 , w_23235 , 
		w_23236 , w_23237 , w_23238 , w_23239 , w_23240 , w_23241 , w_23242 , w_23243 , w_23244 , w_23245 , 
		w_23246 , w_23247 , w_23248 , w_23249 , w_23250 , w_23251 , w_23252 , w_23253 , w_23254 , w_23255 , 
		w_23256 , w_23257 , w_23258 , w_23259 , w_23260 , w_23261 , w_23262 , w_23263 , w_23264 , w_23265 , 
		w_23266 , w_23267 , w_23268 , w_23269 , w_23270 , w_23271 , w_23272 , w_23273 , w_23274 , w_23275 , 
		w_23276 , w_23277 , w_23278 , w_23279 , w_23280 , w_23281 , w_23282 , w_23283 , w_23284 , w_23285 , 
		w_23286 , w_23287 , w_23288 , w_23289 , w_23290 , w_23291 , w_23292 , w_23293 , w_23294 , w_23295 , 
		w_23296 , w_23297 , w_23298 , w_23299 , w_23300 , w_23301 , w_23302 , w_23303 , w_23304 , w_23305 , 
		w_23306 , w_23307 , w_23308 , w_23309 , w_23310 , w_23311 , w_23312 , w_23313 , w_23314 , w_23315 , 
		w_23316 , w_23317 , w_23318 , w_23319 , w_23320 , w_23321 , w_23322 , w_23323 , w_23324 , w_23325 , 
		w_23326 , w_23327 , w_23328 , w_23329 , w_23330 , w_23331 , w_23332 , w_23333 , w_23334 , w_23335 , 
		w_23336 , w_23337 , w_23338 , w_23339 , w_23340 , w_23341 , w_23342 , w_23343 , w_23344 , w_23345 , 
		w_23346 , w_23347 , w_23348 , w_23349 , w_23350 , w_23351 , w_23352 , w_23353 , w_23354 , w_23355 , 
		w_23356 , w_23357 , w_23358 , w_23359 , w_23360 , w_23361 , w_23362 , w_23363 , w_23364 , w_23365 , 
		w_23366 , w_23367 , w_23368 , w_23369 , w_23370 , w_23371 , w_23372 , w_23373 , w_23374 , w_23375 , 
		w_23376 , w_23377 , w_23378 , w_23379 , w_23380 , w_23381 , w_23382 , w_23383 , w_23384 , w_23385 , 
		w_23386 , w_23387 , w_23388 , w_23389 , w_23390 , w_23391 , w_23392 , w_23393 , w_23394 , w_23395 , 
		w_23396 , w_23397 , w_23398 , w_23399 , w_23400 , w_23401 , w_23402 , w_23403 , w_23404 , w_23405 , 
		w_23406 , w_23407 , w_23408 , w_23409 , w_23410 , w_23411 , w_23412 , w_23413 , w_23414 , w_23415 , 
		w_23416 , w_23417 , w_23418 , w_23419 , w_23420 , w_23421 , w_23422 , w_23423 , w_23424 , w_23425 , 
		w_23426 , w_23427 , w_23428 , w_23429 , w_23430 , w_23431 , w_23432 , w_23433 , w_23434 , w_23435 , 
		w_23436 , w_23437 , w_23438 , w_23439 , w_23440 , w_23441 , w_23442 , w_23443 , w_23444 , w_23445 , 
		w_23446 , w_23447 , w_23448 , w_23449 , w_23450 , w_23451 , w_23452 , w_23453 , w_23454 , w_23455 , 
		w_23456 , w_23457 , w_23458 , w_23459 , w_23460 , w_23461 , w_23462 , w_23463 , w_23464 , w_23465 , 
		w_23466 , w_23467 , w_23468 , w_23469 , w_23470 , w_23471 , w_23472 , w_23473 , w_23474 , w_23475 , 
		w_23476 , w_23477 , w_23478 , w_23479 , w_23480 , w_23481 , w_23482 , w_23483 , w_23484 , w_23485 , 
		w_23486 , w_23487 , w_23488 , w_23489 , w_23490 , w_23491 , w_23492 , w_23493 , w_23494 , w_23495 , 
		w_23496 , w_23497 , w_23498 , w_23499 , w_23500 , w_23501 , w_23502 , w_23503 , w_23504 , w_23505 , 
		w_23506 , w_23507 , w_23508 , w_23509 , w_23510 , w_23511 , w_23512 , w_23513 , w_23514 , w_23515 , 
		w_23516 , w_23517 , w_23518 , w_23519 , w_23520 , w_23521 , w_23522 , w_23523 , w_23524 , w_23525 , 
		w_23526 , w_23527 , w_23528 , w_23529 , w_23530 , w_23531 , w_23532 , w_23533 , w_23534 , w_23535 , 
		w_23536 , w_23537 , w_23538 , w_23539 , w_23540 , w_23541 , w_23542 , w_23543 , w_23544 , w_23545 , 
		w_23546 , w_23547 , w_23548 , w_23549 , w_23550 , w_23551 , w_23552 , w_23553 , w_23554 , w_23555 , 
		w_23556 , w_23557 , w_23558 , w_23559 , w_23560 , w_23561 , w_23562 , w_23563 , w_23564 , w_23565 , 
		w_23566 , w_23567 , w_23568 , w_23569 , w_23570 , w_23571 , w_23572 , w_23573 , w_23574 , w_23575 , 
		w_23576 , w_23577 , w_23578 , w_23579 , w_23580 , w_23581 , w_23582 , w_23583 , w_23584 , w_23585 , 
		w_23586 , w_23587 , w_23588 , w_23589 , w_23590 , w_23591 , w_23592 , w_23593 , w_23594 , w_23595 , 
		w_23596 , w_23597 , w_23598 , w_23599 , w_23600 , w_23601 , w_23602 , w_23603 , w_23604 , w_23605 , 
		w_23606 , w_23607 , w_23608 , w_23609 , w_23610 , w_23611 , w_23612 , w_23613 , w_23614 , w_23615 , 
		w_23616 , w_23617 , w_23618 , w_23619 , w_23620 , w_23621 , w_23622 , w_23623 , w_23624 , w_23625 , 
		w_23626 , w_23627 , w_23628 , w_23629 , w_23630 , w_23631 , w_23632 , w_23633 , w_23634 , w_23635 , 
		w_23636 , w_23637 , w_23638 , w_23639 , w_23640 , w_23641 , w_23642 , w_23643 , w_23644 , w_23645 , 
		w_23646 , w_23647 , w_23648 , w_23649 , w_23650 , w_23651 , w_23652 , w_23653 , w_23654 , w_23655 , 
		w_23656 , w_23657 , w_23658 , w_23659 , w_23660 , w_23661 , w_23662 , w_23663 , w_23664 , w_23665 , 
		w_23666 , w_23667 , w_23668 , w_23669 , w_23670 , w_23671 , w_23672 , w_23673 , w_23674 , w_23675 , 
		w_23676 , w_23677 , w_23678 , w_23679 , w_23680 , w_23681 , w_23682 , w_23683 , w_23684 , w_23685 , 
		w_23686 , w_23687 , w_23688 , w_23689 , w_23690 , w_23691 , w_23692 , w_23693 , w_23694 , w_23695 , 
		w_23696 , w_23697 , w_23698 , w_23699 , w_23700 , w_23701 , w_23702 , w_23703 , w_23704 , w_23705 , 
		w_23706 , w_23707 , w_23708 , w_23709 , w_23710 , w_23711 , w_23712 , w_23713 , w_23714 , w_23715 , 
		w_23716 , w_23717 , w_23718 , w_23719 , w_23720 , w_23721 , w_23722 , w_23723 , w_23724 , w_23725 , 
		w_23726 , w_23727 , w_23728 , w_23729 , w_23730 , w_23731 , w_23732 , w_23733 , w_23734 , w_23735 , 
		w_23736 , w_23737 , w_23738 , w_23739 , w_23740 , w_23741 , w_23742 , w_23743 , w_23744 , w_23745 , 
		w_23746 , w_23747 , w_23748 , w_23749 , w_23750 , w_23751 , w_23752 , w_23753 , w_23754 , w_23755 , 
		w_23756 , w_23757 , w_23758 , w_23759 , w_23760 , w_23761 , w_23762 , w_23763 , w_23764 , w_23765 , 
		w_23766 , w_23767 , w_23768 , w_23769 , w_23770 , w_23771 , w_23772 , w_23773 , w_23774 , w_23775 , 
		w_23776 , w_23777 , w_23778 , w_23779 , w_23780 , w_23781 , w_23782 , w_23783 , w_23784 , w_23785 , 
		w_23786 , w_23787 , w_23788 , w_23789 , w_23790 , w_23791 , w_23792 , w_23793 , w_23794 , w_23795 , 
		w_23796 , w_23797 , w_23798 , w_23799 , w_23800 , w_23801 , w_23802 , w_23803 , w_23804 , w_23805 , 
		w_23806 , w_23807 , w_23808 , w_23809 , w_23810 , w_23811 , w_23812 , w_23813 , w_23814 , w_23815 , 
		w_23816 , w_23817 , w_23818 , w_23819 , w_23820 , w_23821 , w_23822 , w_23823 , w_23824 , w_23825 , 
		w_23826 , w_23827 , w_23828 , w_23829 , w_23830 , w_23831 , w_23832 , w_23833 , w_23834 , w_23835 , 
		w_23836 , w_23837 , w_23838 , w_23839 , w_23840 , w_23841 , w_23842 , w_23843 , w_23844 , w_23845 , 
		w_23846 , w_23847 , w_23848 , w_23849 , w_23850 , w_23851 , w_23852 , w_23853 , w_23854 , w_23855 , 
		w_23856 , w_23857 , w_23858 , w_23859 , w_23860 , w_23861 , w_23862 , w_23863 , w_23864 , w_23865 , 
		w_23866 , w_23867 , w_23868 , w_23869 , w_23870 , w_23871 , w_23872 , w_23873 , w_23874 , w_23875 , 
		w_23876 , w_23877 , w_23878 , w_23879 , w_23880 , w_23881 , w_23882 , w_23883 , w_23884 , w_23885 , 
		w_23886 , w_23887 , w_23888 , w_23889 , w_23890 , w_23891 , w_23892 , w_23893 , w_23894 , w_23895 , 
		w_23896 , w_23897 , w_23898 , w_23899 , w_23900 , w_23901 , w_23902 , w_23903 , w_23904 , w_23905 , 
		w_23906 , w_23907 , w_23908 , w_23909 , w_23910 , w_23911 , w_23912 , w_23913 , w_23914 , w_23915 , 
		w_23916 , w_23917 , w_23918 , w_23919 , w_23920 , w_23921 , w_23922 , w_23923 , w_23924 , w_23925 , 
		w_23926 , w_23927 , w_23928 , w_23929 , w_23930 , w_23931 , w_23932 , w_23933 , w_23934 , w_23935 , 
		w_23936 , w_23937 , w_23938 , w_23939 , w_23940 , w_23941 , w_23942 , w_23943 , w_23944 , w_23945 , 
		w_23946 , w_23947 , w_23948 , w_23949 , w_23950 , w_23951 , w_23952 , w_23953 , w_23954 , w_23955 , 
		w_23956 , w_23957 , w_23958 , w_23959 , w_23960 , w_23961 , w_23962 , w_23963 , w_23964 , w_23965 , 
		w_23966 , w_23967 , w_23968 , w_23969 , w_23970 , w_23971 , w_23972 , w_23973 , w_23974 , w_23975 , 
		w_23976 , w_23977 , w_23978 , w_23979 , w_23980 , w_23981 , w_23982 , w_23983 , w_23984 , w_23985 , 
		w_23986 , w_23987 , w_23988 , w_23989 , w_23990 , w_23991 , w_23992 , w_23993 , w_23994 , w_23995 , 
		w_23996 , w_23997 , w_23998 , w_23999 , w_24000 , w_24001 , w_24002 , w_24003 , w_24004 , w_24005 , 
		w_24006 , w_24007 , w_24008 , w_24009 , w_24010 , w_24011 , w_24012 , w_24013 , w_24014 , w_24015 , 
		w_24016 , w_24017 , w_24018 , w_24019 , w_24020 , w_24021 , w_24022 , w_24023 , w_24024 , w_24025 , 
		w_24026 , w_24027 , w_24028 , w_24029 , w_24030 , w_24031 , w_24032 , w_24033 , w_24034 , w_24035 , 
		w_24036 , w_24037 , w_24038 , w_24039 , w_24040 , w_24041 , w_24042 , w_24043 , w_24044 , w_24045 , 
		w_24046 , w_24047 , w_24048 , w_24049 , w_24050 , w_24051 , w_24052 , w_24053 , w_24054 , w_24055 , 
		w_24056 , w_24057 , w_24058 , w_24059 , w_24060 , w_24061 , w_24062 , w_24063 , w_24064 , w_24065 , 
		w_24066 , w_24067 , w_24068 , w_24069 , w_24070 , w_24071 , w_24072 , w_24073 , w_24074 , w_24075 , 
		w_24076 , w_24077 , w_24078 , w_24079 , w_24080 , w_24081 , w_24082 , w_24083 , w_24084 , w_24085 , 
		w_24086 , w_24087 , w_24088 , w_24089 , w_24090 , w_24091 , w_24092 , w_24093 , w_24094 , w_24095 , 
		w_24096 , w_24097 , w_24098 , w_24099 , w_24100 , w_24101 , w_24102 , w_24103 , w_24104 , w_24105 , 
		w_24106 , w_24107 , w_24108 , w_24109 , w_24110 , w_24111 , w_24112 , w_24113 , w_24114 , w_24115 , 
		w_24116 , w_24117 , w_24118 , w_24119 , w_24120 , w_24121 , w_24122 , w_24123 , w_24124 , w_24125 , 
		w_24126 , w_24127 , w_24128 , w_24129 , w_24130 , w_24131 , w_24132 , w_24133 , w_24134 , w_24135 , 
		w_24136 , w_24137 , w_24138 , w_24139 , w_24140 , w_24141 , w_24142 , w_24143 , w_24144 , w_24145 , 
		w_24146 , w_24147 , w_24148 , w_24149 , w_24150 , w_24151 , w_24152 , w_24153 , w_24154 , w_24155 , 
		w_24156 , w_24157 , w_24158 , w_24159 , w_24160 , w_24161 , w_24162 , w_24163 , w_24164 , w_24165 , 
		w_24166 , w_24167 , w_24168 , w_24169 , w_24170 , w_24171 , w_24172 , w_24173 , w_24174 , w_24175 , 
		w_24176 , w_24177 , w_24178 , w_24179 , w_24180 , w_24181 , w_24182 , w_24183 , w_24184 , w_24185 , 
		w_24186 , w_24187 , w_24188 , w_24189 , w_24190 , w_24191 , w_24192 , w_24193 , w_24194 , w_24195 , 
		w_24196 , w_24197 , w_24198 , w_24199 , w_24200 , w_24201 , w_24202 , w_24203 , w_24204 , w_24205 , 
		w_24206 , w_24207 , w_24208 , w_24209 , w_24210 , w_24211 , w_24212 , w_24213 , w_24214 , w_24215 , 
		w_24216 , w_24217 , w_24218 , w_24219 , w_24220 , w_24221 , w_24222 , w_24223 , w_24224 , w_24225 , 
		w_24226 , w_24227 , w_24228 , w_24229 , w_24230 , w_24231 , w_24232 , w_24233 , w_24234 , w_24235 , 
		w_24236 , w_24237 , w_24238 , w_24239 , w_24240 , w_24241 , w_24242 , w_24243 , w_24244 , w_24245 , 
		w_24246 , w_24247 , w_24248 , w_24249 , w_24250 , w_24251 , w_24252 , w_24253 , w_24254 , w_24255 , 
		w_24256 , w_24257 , w_24258 , w_24259 , w_24260 , w_24261 , w_24262 , w_24263 , w_24264 , w_24265 , 
		w_24266 , w_24267 , w_24268 , w_24269 , w_24270 , w_24271 , w_24272 , w_24273 , w_24274 , w_24275 , 
		w_24276 , w_24277 , w_24278 , w_24279 , w_24280 , w_24281 , w_24282 , w_24283 , w_24284 , w_24285 , 
		w_24286 , w_24287 , w_24288 , w_24289 , w_24290 , w_24291 , w_24292 , w_24293 , w_24294 , w_24295 , 
		w_24296 , w_24297 , w_24298 , w_24299 , w_24300 , w_24301 , w_24302 , w_24303 , w_24304 , w_24305 , 
		w_24306 , w_24307 , w_24308 , w_24309 , w_24310 , w_24311 , w_24312 , w_24313 , w_24314 , w_24315 , 
		w_24316 , w_24317 , w_24318 , w_24319 , w_24320 , w_24321 , w_24322 , w_24323 , w_24324 , w_24325 , 
		w_24326 , w_24327 , w_24328 , w_24329 , w_24330 , w_24331 , w_24332 , w_24333 , w_24334 , w_24335 , 
		w_24336 , w_24337 , w_24338 , w_24339 , w_24340 , w_24341 , w_24342 , w_24343 , w_24344 , w_24345 , 
		w_24346 , w_24347 , w_24348 , w_24349 , w_24350 , w_24351 , w_24352 , w_24353 , w_24354 , w_24355 , 
		w_24356 , w_24357 , w_24358 , w_24359 , w_24360 , w_24361 , w_24362 , w_24363 , w_24364 , w_24365 , 
		w_24366 , w_24367 , w_24368 , w_24369 , w_24370 , w_24371 , w_24372 , w_24373 , w_24374 , w_24375 , 
		w_24376 , w_24377 , w_24378 , w_24379 , w_24380 , w_24381 , w_24382 , w_24383 , w_24384 , w_24385 , 
		w_24386 , w_24387 , w_24388 , w_24389 , w_24390 , w_24391 , w_24392 , w_24393 , w_24394 , w_24395 , 
		w_24396 , w_24397 , w_24398 , w_24399 , w_24400 , w_24401 , w_24402 , w_24403 , w_24404 , w_24405 , 
		w_24406 , w_24407 , w_24408 , w_24409 , w_24410 , w_24411 , w_24412 , w_24413 , w_24414 , w_24415 , 
		w_24416 , w_24417 , w_24418 , w_24419 , w_24420 , w_24421 , w_24422 , w_24423 , w_24424 , w_24425 , 
		w_24426 , w_24427 , w_24428 , w_24429 , w_24430 , w_24431 , w_24432 , w_24433 , w_24434 , w_24435 , 
		w_24436 , w_24437 , w_24438 , w_24439 , w_24440 , w_24441 , w_24442 , w_24443 , w_24444 , w_24445 , 
		w_24446 , w_24447 , w_24448 , w_24449 , w_24450 , w_24451 , w_24452 , w_24453 , w_24454 , w_24455 , 
		w_24456 , w_24457 , w_24458 , w_24459 , w_24460 , w_24461 , w_24462 , w_24463 , w_24464 , w_24465 , 
		w_24466 , w_24467 , w_24468 , w_24469 , w_24470 , w_24471 , w_24472 , w_24473 , w_24474 , w_24475 , 
		w_24476 , w_24477 , w_24478 , w_24479 , w_24480 , w_24481 , w_24482 , w_24483 , w_24484 , w_24485 , 
		w_24486 , w_24487 , w_24488 , w_24489 , w_24490 , w_24491 , w_24492 , w_24493 , w_24494 , w_24495 , 
		w_24496 , w_24497 , w_24498 , w_24499 , w_24500 , w_24501 , w_24502 , w_24503 , w_24504 , w_24505 , 
		w_24506 , w_24507 , w_24508 , w_24509 , w_24510 , w_24511 , w_24512 , w_24513 , w_24514 , w_24515 , 
		w_24516 , w_24517 , w_24518 , w_24519 , w_24520 , w_24521 , w_24522 , w_24523 , w_24524 , w_24525 , 
		w_24526 , w_24527 , w_24528 , w_24529 , w_24530 , w_24531 , w_24532 , w_24533 , w_24534 , w_24535 , 
		w_24536 , w_24537 , w_24538 , w_24539 , w_24540 , w_24541 , w_24542 , w_24543 , w_24544 , w_24545 , 
		w_24546 , w_24547 , w_24548 , w_24549 , w_24550 , w_24551 , w_24552 , w_24553 , w_24554 , w_24555 , 
		w_24556 , w_24557 , w_24558 , w_24559 , w_24560 , w_24561 , w_24562 , w_24563 , w_24564 , w_24565 , 
		w_24566 , w_24567 , w_24568 , w_24569 , w_24570 , w_24571 , w_24572 , w_24573 , w_24574 , w_24575 , 
		w_24576 , w_24577 , w_24578 , w_24579 , w_24580 , w_24581 , w_24582 , w_24583 , w_24584 , w_24585 , 
		w_24586 , w_24587 , w_24588 , w_24589 , w_24590 , w_24591 , w_24592 , w_24593 , w_24594 , w_24595 , 
		w_24596 , w_24597 , w_24598 , w_24599 , w_24600 , w_24601 , w_24602 , w_24603 , w_24604 , w_24605 , 
		w_24606 , w_24607 , w_24608 , w_24609 , w_24610 , w_24611 , w_24612 , w_24613 , w_24614 , w_24615 , 
		w_24616 , w_24617 , w_24618 , w_24619 , w_24620 , w_24621 , w_24622 , w_24623 , w_24624 , w_24625 , 
		w_24626 , w_24627 , w_24628 , w_24629 , w_24630 , w_24631 , w_24632 , w_24633 , w_24634 , w_24635 , 
		w_24636 , w_24637 , w_24638 , w_24639 , w_24640 , w_24641 , w_24642 , w_24643 , w_24644 , w_24645 , 
		w_24646 , w_24647 , w_24648 , w_24649 , w_24650 , w_24651 , w_24652 , w_24653 , w_24654 , w_24655 , 
		w_24656 , w_24657 , w_24658 , w_24659 , w_24660 , w_24661 , w_24662 , w_24663 , w_24664 , w_24665 , 
		w_24666 , w_24667 , w_24668 , w_24669 , w_24670 , w_24671 , w_24672 , w_24673 , w_24674 , w_24675 , 
		w_24676 , w_24677 , w_24678 , w_24679 , w_24680 , w_24681 , w_24682 , w_24683 , w_24684 , w_24685 , 
		w_24686 , w_24687 , w_24688 , w_24689 , w_24690 , w_24691 , w_24692 , w_24693 , w_24694 , w_24695 , 
		w_24696 , w_24697 , w_24698 , w_24699 , w_24700 , w_24701 , w_24702 , w_24703 , w_24704 , w_24705 , 
		w_24706 , w_24707 , w_24708 , w_24709 , w_24710 , w_24711 , w_24712 , w_24713 , w_24714 , w_24715 , 
		w_24716 , w_24717 , w_24718 , w_24719 , w_24720 , w_24721 , w_24722 , w_24723 , w_24724 , w_24725 , 
		w_24726 , w_24727 , w_24728 , w_24729 , w_24730 , w_24731 , w_24732 , w_24733 , w_24734 , w_24735 , 
		w_24736 , w_24737 , w_24738 , w_24739 , w_24740 , w_24741 , w_24742 , w_24743 , w_24744 , w_24745 , 
		w_24746 , w_24747 , w_24748 , w_24749 , w_24750 , w_24751 , w_24752 , w_24753 , w_24754 , w_24755 , 
		w_24756 , w_24757 , w_24758 , w_24759 , w_24760 , w_24761 , w_24762 , w_24763 , w_24764 , w_24765 , 
		w_24766 , w_24767 , w_24768 , w_24769 , w_24770 , w_24771 , w_24772 , w_24773 , w_24774 , w_24775 , 
		w_24776 , w_24777 , w_24778 , w_24779 , w_24780 , w_24781 , w_24782 , w_24783 , w_24784 , w_24785 , 
		w_24786 , w_24787 , w_24788 , w_24789 , w_24790 , w_24791 , w_24792 , w_24793 , w_24794 , w_24795 , 
		w_24796 , w_24797 , w_24798 , w_24799 , w_24800 , w_24801 , w_24802 , w_24803 , w_24804 , w_24805 , 
		w_24806 , w_24807 , w_24808 , w_24809 , w_24810 , w_24811 , w_24812 , w_24813 , w_24814 , w_24815 , 
		w_24816 , w_24817 , w_24818 , w_24819 , w_24820 , w_24821 , w_24822 , w_24823 , w_24824 , w_24825 , 
		w_24826 , w_24827 , w_24828 , w_24829 , w_24830 , w_24831 , w_24832 , w_24833 , w_24834 , w_24835 , 
		w_24836 , w_24837 , w_24838 , w_24839 , w_24840 , w_24841 , w_24842 , w_24843 , w_24844 , w_24845 , 
		w_24846 , w_24847 , w_24848 , w_24849 , w_24850 , w_24851 , w_24852 , w_24853 , w_24854 , w_24855 , 
		w_24856 , w_24857 , w_24858 , w_24859 , w_24860 , w_24861 , w_24862 , w_24863 , w_24864 , w_24865 , 
		w_24866 , w_24867 , w_24868 , w_24869 , w_24870 , w_24871 , w_24872 , w_24873 , w_24874 , w_24875 , 
		w_24876 , w_24877 , w_24878 , w_24879 , w_24880 , w_24881 , w_24882 , w_24883 , w_24884 , w_24885 , 
		w_24886 , w_24887 , w_24888 , w_24889 , w_24890 , w_24891 , w_24892 , w_24893 , w_24894 , w_24895 , 
		w_24896 , w_24897 , w_24898 , w_24899 , w_24900 , w_24901 , w_24902 , w_24903 , w_24904 , w_24905 , 
		w_24906 , w_24907 , w_24908 , w_24909 , w_24910 , w_24911 , w_24912 , w_24913 , w_24914 , w_24915 , 
		w_24916 , w_24917 , w_24918 , w_24919 , w_24920 , w_24921 , w_24922 , w_24923 , w_24924 , w_24925 , 
		w_24926 , w_24927 , w_24928 , w_24929 , w_24930 , w_24931 , w_24932 , w_24933 , w_24934 , w_24935 , 
		w_24936 , w_24937 , w_24938 , w_24939 , w_24940 , w_24941 , w_24942 , w_24943 , w_24944 , w_24945 , 
		w_24946 , w_24947 , w_24948 , w_24949 , w_24950 , w_24951 , w_24952 , w_24953 , w_24954 , w_24955 , 
		w_24956 , w_24957 , w_24958 , w_24959 , w_24960 , w_24961 , w_24962 , w_24963 , w_24964 , w_24965 , 
		w_24966 , w_24967 , w_24968 , w_24969 , w_24970 , w_24971 , w_24972 , w_24973 , w_24974 , w_24975 , 
		w_24976 , w_24977 , w_24978 , w_24979 , w_24980 , w_24981 , w_24982 , w_24983 , w_24984 , w_24985 , 
		w_24986 , w_24987 , w_24988 , w_24989 , w_24990 , w_24991 , w_24992 , w_24993 , w_24994 , w_24995 , 
		w_24996 , w_24997 , w_24998 , w_24999 , w_25000 , w_25001 , w_25002 , w_25003 , w_25004 , w_25005 , 
		w_25006 , w_25007 , w_25008 , w_25009 , w_25010 , w_25011 , w_25012 , w_25013 , w_25014 , w_25015 , 
		w_25016 , w_25017 , w_25018 , w_25019 , w_25020 , w_25021 , w_25022 , w_25023 , w_25024 , w_25025 , 
		w_25026 , w_25027 , w_25028 , w_25029 , w_25030 , w_25031 , w_25032 , w_25033 , w_25034 , w_25035 , 
		w_25036 , w_25037 , w_25038 , w_25039 , w_25040 , w_25041 , w_25042 , w_25043 , w_25044 , w_25045 , 
		w_25046 , w_25047 , w_25048 , w_25049 , w_25050 , w_25051 , w_25052 , w_25053 , w_25054 , w_25055 , 
		w_25056 , w_25057 , w_25058 , w_25059 , w_25060 , w_25061 , w_25062 , w_25063 , w_25064 , w_25065 , 
		w_25066 , w_25067 , w_25068 , w_25069 , w_25070 , w_25071 , w_25072 , w_25073 , w_25074 , w_25075 , 
		w_25076 , w_25077 , w_25078 , w_25079 , w_25080 , w_25081 , w_25082 , w_25083 , w_25084 , w_25085 , 
		w_25086 , w_25087 , w_25088 , w_25089 , w_25090 , w_25091 , w_25092 , w_25093 , w_25094 , w_25095 , 
		w_25096 , w_25097 , w_25098 , w_25099 , w_25100 , w_25101 , w_25102 , w_25103 , w_25104 , w_25105 , 
		w_25106 , w_25107 , w_25108 , w_25109 , w_25110 , w_25111 , w_25112 , w_25113 , w_25114 , w_25115 , 
		w_25116 , w_25117 , w_25118 , w_25119 , w_25120 , w_25121 , w_25122 , w_25123 , w_25124 , w_25125 , 
		w_25126 , w_25127 , w_25128 , w_25129 , w_25130 , w_25131 , w_25132 , w_25133 , w_25134 , w_25135 , 
		w_25136 , w_25137 , w_25138 , w_25139 , w_25140 , w_25141 , w_25142 , w_25143 , w_25144 , w_25145 , 
		w_25146 , w_25147 , w_25148 , w_25149 , w_25150 , w_25151 , w_25152 , w_25153 , w_25154 , w_25155 , 
		w_25156 , w_25157 , w_25158 , w_25159 , w_25160 , w_25161 , w_25162 , w_25163 , w_25164 , w_25165 , 
		w_25166 , w_25167 , w_25168 , w_25169 , w_25170 , w_25171 , w_25172 , w_25173 , w_25174 , w_25175 , 
		w_25176 , w_25177 , w_25178 , w_25179 , w_25180 , w_25181 , w_25182 , w_25183 , w_25184 , w_25185 , 
		w_25186 , w_25187 , w_25188 , w_25189 , w_25190 , w_25191 , w_25192 , w_25193 , w_25194 , w_25195 , 
		w_25196 , w_25197 , w_25198 , w_25199 , w_25200 , w_25201 , w_25202 , w_25203 , w_25204 , w_25205 , 
		w_25206 , w_25207 , w_25208 , w_25209 , w_25210 , w_25211 , w_25212 , w_25213 , w_25214 , w_25215 , 
		w_25216 , w_25217 , w_25218 , w_25219 , w_25220 , w_25221 , w_25222 , w_25223 , w_25224 , w_25225 , 
		w_25226 , w_25227 , w_25228 , w_25229 , w_25230 , w_25231 , w_25232 , w_25233 , w_25234 , w_25235 , 
		w_25236 , w_25237 , w_25238 , w_25239 , w_25240 , w_25241 , w_25242 , w_25243 , w_25244 , w_25245 , 
		w_25246 , w_25247 , w_25248 , w_25249 , w_25250 , w_25251 , w_25252 , w_25253 , w_25254 , w_25255 , 
		w_25256 , w_25257 , w_25258 , w_25259 , w_25260 , w_25261 , w_25262 , w_25263 , w_25264 , w_25265 , 
		w_25266 , w_25267 , w_25268 , w_25269 , w_25270 , w_25271 , w_25272 , w_25273 , w_25274 , w_25275 , 
		w_25276 , w_25277 , w_25278 , w_25279 , w_25280 , w_25281 , w_25282 , w_25283 , w_25284 , w_25285 , 
		w_25286 , w_25287 , w_25288 , w_25289 , w_25290 , w_25291 , w_25292 , w_25293 , w_25294 , w_25295 , 
		w_25296 , w_25297 , w_25298 , w_25299 , w_25300 , w_25301 , w_25302 , w_25303 , w_25304 , w_25305 , 
		w_25306 , w_25307 , w_25308 , w_25309 , w_25310 , w_25311 , w_25312 , w_25313 , w_25314 , w_25315 , 
		w_25316 , w_25317 , w_25318 , w_25319 , w_25320 , w_25321 , w_25322 , w_25323 , w_25324 , w_25325 , 
		w_25326 , w_25327 , w_25328 , w_25329 , w_25330 , w_25331 , w_25332 , w_25333 , w_25334 , w_25335 , 
		w_25336 , w_25337 , w_25338 , w_25339 , w_25340 , w_25341 , w_25342 , w_25343 , w_25344 , w_25345 , 
		w_25346 , w_25347 , w_25348 , w_25349 , w_25350 , w_25351 , w_25352 , w_25353 , w_25354 , w_25355 , 
		w_25356 , w_25357 , w_25358 , w_25359 , w_25360 , w_25361 , w_25362 , w_25363 , w_25364 , w_25365 , 
		w_25366 , w_25367 , w_25368 , w_25369 , w_25370 , w_25371 , w_25372 , w_25373 , w_25374 , w_25375 , 
		w_25376 , w_25377 , w_25378 , w_25379 , w_25380 , w_25381 , w_25382 , w_25383 , w_25384 , w_25385 , 
		w_25386 , w_25387 , w_25388 , w_25389 , w_25390 , w_25391 , w_25392 , w_25393 , w_25394 , w_25395 , 
		w_25396 , w_25397 , w_25398 , w_25399 , w_25400 , w_25401 , w_25402 , w_25403 , w_25404 , w_25405 , 
		w_25406 , w_25407 , w_25408 , w_25409 , w_25410 , w_25411 , w_25412 , w_25413 , w_25414 , w_25415 , 
		w_25416 , w_25417 , w_25418 , w_25419 , w_25420 , w_25421 , w_25422 , w_25423 , w_25424 , w_25425 , 
		w_25426 , w_25427 , w_25428 , w_25429 , w_25430 , w_25431 , w_25432 , w_25433 , w_25434 , w_25435 , 
		w_25436 , w_25437 , w_25438 , w_25439 , w_25440 , w_25441 , w_25442 , w_25443 , w_25444 , w_25445 , 
		w_25446 , w_25447 , w_25448 , w_25449 , w_25450 , w_25451 , w_25452 , w_25453 , w_25454 , w_25455 , 
		w_25456 , w_25457 , w_25458 , w_25459 , w_25460 , w_25461 , w_25462 , w_25463 , w_25464 , w_25465 , 
		w_25466 , w_25467 , w_25468 , w_25469 , w_25470 , w_25471 , w_25472 , w_25473 , w_25474 , w_25475 , 
		w_25476 , w_25477 , w_25478 , w_25479 , w_25480 , w_25481 , w_25482 , w_25483 , w_25484 , w_25485 , 
		w_25486 , w_25487 , w_25488 , w_25489 , w_25490 , w_25491 , w_25492 , w_25493 , w_25494 , w_25495 , 
		w_25496 , w_25497 , w_25498 , w_25499 , w_25500 , w_25501 , w_25502 , w_25503 , w_25504 , w_25505 , 
		w_25506 , w_25507 , w_25508 , w_25509 , w_25510 , w_25511 , w_25512 , w_25513 , w_25514 , w_25515 , 
		w_25516 , w_25517 , w_25518 , w_25519 , w_25520 , w_25521 , w_25522 , w_25523 , w_25524 , w_25525 , 
		w_25526 , w_25527 , w_25528 , w_25529 , w_25530 , w_25531 , w_25532 , w_25533 , w_25534 , w_25535 , 
		w_25536 , w_25537 , w_25538 , w_25539 , w_25540 , w_25541 , w_25542 , w_25543 , w_25544 , w_25545 , 
		w_25546 , w_25547 , w_25548 , w_25549 , w_25550 , w_25551 , w_25552 , w_25553 , w_25554 , w_25555 , 
		w_25556 , w_25557 , w_25558 , w_25559 , w_25560 , w_25561 , w_25562 , w_25563 , w_25564 , w_25565 , 
		w_25566 , w_25567 , w_25568 , w_25569 , w_25570 , w_25571 , w_25572 , w_25573 , w_25574 , w_25575 , 
		w_25576 , w_25577 , w_25578 , w_25579 , w_25580 , w_25581 , w_25582 , w_25583 , w_25584 , w_25585 , 
		w_25586 , w_25587 , w_25588 , w_25589 , w_25590 , w_25591 , w_25592 , w_25593 , w_25594 , w_25595 , 
		w_25596 , w_25597 , w_25598 , w_25599 , w_25600 , w_25601 , w_25602 , w_25603 , w_25604 , w_25605 , 
		w_25606 , w_25607 , w_25608 , w_25609 , w_25610 , w_25611 , w_25612 , w_25613 , w_25614 , w_25615 , 
		w_25616 , w_25617 , w_25618 , w_25619 , w_25620 , w_25621 , w_25622 , w_25623 , w_25624 , w_25625 , 
		w_25626 , w_25627 , w_25628 , w_25629 , w_25630 , w_25631 , w_25632 , w_25633 , w_25634 , w_25635 , 
		w_25636 , w_25637 , w_25638 , w_25639 , w_25640 , w_25641 , w_25642 , w_25643 , w_25644 , w_25645 , 
		w_25646 , w_25647 , w_25648 , w_25649 , w_25650 , w_25651 , w_25652 , w_25653 , w_25654 , w_25655 , 
		w_25656 , w_25657 , w_25658 , w_25659 , w_25660 , w_25661 , w_25662 , w_25663 , w_25664 , w_25665 , 
		w_25666 , w_25667 , w_25668 , w_25669 , w_25670 , w_25671 , w_25672 , w_25673 , w_25674 , w_25675 , 
		w_25676 , w_25677 , w_25678 , w_25679 , w_25680 , w_25681 , w_25682 , w_25683 , w_25684 , w_25685 , 
		w_25686 , w_25687 , w_25688 , w_25689 , w_25690 , w_25691 , w_25692 , w_25693 , w_25694 , w_25695 , 
		w_25696 , w_25697 , w_25698 , w_25699 , w_25700 , w_25701 , w_25702 , w_25703 , w_25704 , w_25705 , 
		w_25706 , w_25707 , w_25708 , w_25709 , w_25710 , w_25711 , w_25712 , w_25713 , w_25714 , w_25715 , 
		w_25716 , w_25717 , w_25718 , w_25719 , w_25720 , w_25721 , w_25722 , w_25723 , w_25724 , w_25725 , 
		w_25726 , w_25727 , w_25728 , w_25729 , w_25730 , w_25731 , w_25732 , w_25733 , w_25734 , w_25735 , 
		w_25736 , w_25737 , w_25738 , w_25739 , w_25740 , w_25741 , w_25742 , w_25743 , w_25744 , w_25745 , 
		w_25746 , w_25747 , w_25748 , w_25749 , w_25750 , w_25751 , w_25752 , w_25753 , w_25754 , w_25755 , 
		w_25756 , w_25757 , w_25758 , w_25759 , w_25760 , w_25761 , w_25762 , w_25763 , w_25764 , w_25765 , 
		w_25766 , w_25767 , w_25768 , w_25769 , w_25770 , w_25771 , w_25772 , w_25773 , w_25774 , w_25775 , 
		w_25776 , w_25777 , w_25778 , w_25779 , w_25780 , w_25781 , w_25782 , w_25783 , w_25784 , w_25785 , 
		w_25786 , w_25787 , w_25788 , w_25789 , w_25790 , w_25791 , w_25792 , w_25793 , w_25794 , w_25795 , 
		w_25796 , w_25797 , w_25798 , w_25799 , w_25800 , w_25801 , w_25802 , w_25803 , w_25804 , w_25805 , 
		w_25806 , w_25807 , w_25808 , w_25809 , w_25810 , w_25811 , w_25812 , w_25813 , w_25814 , w_25815 , 
		w_25816 , w_25817 , w_25818 , w_25819 , w_25820 , w_25821 , w_25822 , w_25823 , w_25824 , w_25825 , 
		w_25826 , w_25827 , w_25828 , w_25829 , w_25830 , w_25831 , w_25832 , w_25833 , w_25834 , w_25835 , 
		w_25836 , w_25837 , w_25838 , w_25839 , w_25840 , w_25841 , w_25842 , w_25843 , w_25844 , w_25845 , 
		w_25846 , w_25847 , w_25848 , w_25849 , w_25850 , w_25851 , w_25852 , w_25853 , w_25854 , w_25855 , 
		w_25856 , w_25857 , w_25858 , w_25859 , w_25860 , w_25861 , w_25862 , w_25863 , w_25864 , w_25865 , 
		w_25866 , w_25867 , w_25868 , w_25869 , w_25870 , w_25871 , w_25872 , w_25873 , w_25874 , w_25875 , 
		w_25876 , w_25877 , w_25878 , w_25879 , w_25880 , w_25881 , w_25882 , w_25883 , w_25884 , w_25885 , 
		w_25886 , w_25887 , w_25888 , w_25889 , w_25890 , w_25891 , w_25892 , w_25893 , w_25894 , w_25895 , 
		w_25896 , w_25897 , w_25898 , w_25899 , w_25900 , w_25901 , w_25902 , w_25903 , w_25904 , w_25905 , 
		w_25906 , w_25907 , w_25908 , w_25909 , w_25910 , w_25911 , w_25912 , w_25913 , w_25914 , w_25915 , 
		w_25916 , w_25917 , w_25918 , w_25919 , w_25920 , w_25921 , w_25922 , w_25923 , w_25924 , w_25925 , 
		w_25926 , w_25927 , w_25928 , w_25929 , w_25930 , w_25931 , w_25932 , w_25933 , w_25934 , w_25935 , 
		w_25936 , w_25937 , w_25938 , w_25939 , w_25940 , w_25941 , w_25942 , w_25943 , w_25944 , w_25945 , 
		w_25946 , w_25947 , w_25948 , w_25949 , w_25950 , w_25951 , w_25952 , w_25953 , w_25954 , w_25955 , 
		w_25956 , w_25957 , w_25958 , w_25959 , w_25960 , w_25961 , w_25962 , w_25963 , w_25964 , w_25965 , 
		w_25966 , w_25967 , w_25968 , w_25969 , w_25970 , w_25971 , w_25972 , w_25973 , w_25974 , w_25975 , 
		w_25976 , w_25977 , w_25978 , w_25979 , w_25980 , w_25981 , w_25982 , w_25983 , w_25984 , w_25985 , 
		w_25986 , w_25987 , w_25988 , w_25989 , w_25990 , w_25991 , w_25992 , w_25993 , w_25994 , w_25995 , 
		w_25996 , w_25997 , w_25998 , w_25999 , w_26000 , w_26001 , w_26002 , w_26003 , w_26004 , w_26005 , 
		w_26006 , w_26007 , w_26008 , w_26009 , w_26010 , w_26011 , w_26012 , w_26013 , w_26014 , w_26015 , 
		w_26016 , w_26017 , w_26018 , w_26019 , w_26020 , w_26021 , w_26022 , w_26023 , w_26024 , w_26025 , 
		w_26026 , w_26027 , w_26028 , w_26029 , w_26030 , w_26031 , w_26032 , w_26033 , w_26034 , w_26035 , 
		w_26036 , w_26037 , w_26038 , w_26039 , w_26040 , w_26041 , w_26042 , w_26043 , w_26044 , w_26045 , 
		w_26046 , w_26047 , w_26048 , w_26049 , w_26050 , w_26051 , w_26052 , w_26053 , w_26054 , w_26055 , 
		w_26056 , w_26057 , w_26058 , w_26059 , w_26060 , w_26061 , w_26062 , w_26063 , w_26064 , w_26065 , 
		w_26066 , w_26067 , w_26068 , w_26069 , w_26070 , w_26071 , w_26072 , w_26073 , w_26074 , w_26075 , 
		w_26076 , w_26077 , w_26078 , w_26079 , w_26080 , w_26081 , w_26082 , w_26083 , w_26084 , w_26085 , 
		w_26086 , w_26087 , w_26088 , w_26089 , w_26090 , w_26091 , w_26092 , w_26093 , w_26094 , w_26095 , 
		w_26096 , w_26097 , w_26098 , w_26099 , w_26100 , w_26101 , w_26102 , w_26103 , w_26104 , w_26105 , 
		w_26106 , w_26107 , w_26108 , w_26109 , w_26110 , w_26111 , w_26112 , w_26113 , w_26114 , w_26115 , 
		w_26116 , w_26117 , w_26118 , w_26119 , w_26120 , w_26121 , w_26122 , w_26123 , w_26124 , w_26125 , 
		w_26126 , w_26127 , w_26128 , w_26129 , w_26130 , w_26131 , w_26132 , w_26133 , w_26134 , w_26135 , 
		w_26136 , w_26137 , w_26138 , w_26139 , w_26140 , w_26141 , w_26142 , w_26143 , w_26144 , w_26145 , 
		w_26146 , w_26147 , w_26148 , w_26149 , w_26150 , w_26151 , w_26152 , w_26153 , w_26154 , w_26155 , 
		w_26156 , w_26157 , w_26158 , w_26159 , w_26160 , w_26161 , w_26162 , w_26163 , w_26164 , w_26165 , 
		w_26166 , w_26167 , w_26168 , w_26169 , w_26170 , w_26171 , w_26172 , w_26173 , w_26174 , w_26175 , 
		w_26176 , w_26177 , w_26178 , w_26179 , w_26180 , w_26181 , w_26182 , w_26183 , w_26184 , w_26185 , 
		w_26186 , w_26187 , w_26188 , w_26189 , w_26190 , w_26191 , w_26192 , w_26193 , w_26194 , w_26195 , 
		w_26196 , w_26197 , w_26198 , w_26199 , w_26200 , w_26201 , w_26202 , w_26203 , w_26204 , w_26205 , 
		w_26206 , w_26207 , w_26208 , w_26209 , w_26210 , w_26211 , w_26212 , w_26213 , w_26214 , w_26215 , 
		w_26216 , w_26217 , w_26218 , w_26219 , w_26220 , w_26221 , w_26222 , w_26223 , w_26224 , w_26225 , 
		w_26226 , w_26227 , w_26228 , w_26229 , w_26230 , w_26231 , w_26232 , w_26233 , w_26234 , w_26235 , 
		w_26236 , w_26237 , w_26238 , w_26239 , w_26240 , w_26241 , w_26242 , w_26243 , w_26244 , w_26245 , 
		w_26246 , w_26247 , w_26248 , w_26249 , w_26250 , w_26251 , w_26252 , w_26253 , w_26254 , w_26255 , 
		w_26256 , w_26257 , w_26258 , w_26259 , w_26260 , w_26261 , w_26262 , w_26263 , w_26264 , w_26265 , 
		w_26266 , w_26267 , w_26268 , w_26269 , w_26270 , w_26271 , w_26272 , w_26273 , w_26274 , w_26275 , 
		w_26276 , w_26277 , w_26278 , w_26279 , w_26280 , w_26281 , w_26282 , w_26283 , w_26284 , w_26285 , 
		w_26286 , w_26287 , w_26288 , w_26289 , w_26290 , w_26291 , w_26292 , w_26293 , w_26294 , w_26295 , 
		w_26296 , w_26297 , w_26298 , w_26299 , w_26300 , w_26301 , w_26302 , w_26303 , w_26304 , w_26305 , 
		w_26306 , w_26307 , w_26308 , w_26309 , w_26310 , w_26311 , w_26312 , w_26313 , w_26314 , w_26315 , 
		w_26316 , w_26317 , w_26318 , w_26319 , w_26320 , w_26321 , w_26322 , w_26323 , w_26324 , w_26325 , 
		w_26326 , w_26327 , w_26328 , w_26329 , w_26330 , w_26331 , w_26332 , w_26333 , w_26334 , w_26335 , 
		w_26336 , w_26337 , w_26338 , w_26339 , w_26340 , w_26341 , w_26342 , w_26343 , w_26344 , w_26345 , 
		w_26346 , w_26347 , w_26348 , w_26349 , w_26350 , w_26351 , w_26352 , w_26353 , w_26354 , w_26355 , 
		w_26356 , w_26357 , w_26358 , w_26359 , w_26360 , w_26361 , w_26362 , w_26363 , w_26364 , w_26365 , 
		w_26366 , w_26367 , w_26368 , w_26369 , w_26370 , w_26371 , w_26372 , w_26373 , w_26374 , w_26375 , 
		w_26376 , w_26377 , w_26378 , w_26379 , w_26380 , w_26381 , w_26382 , w_26383 , w_26384 , w_26385 , 
		w_26386 , w_26387 , w_26388 , w_26389 , w_26390 , w_26391 , w_26392 , w_26393 , w_26394 , w_26395 , 
		w_26396 , w_26397 , w_26398 , w_26399 , w_26400 , w_26401 , w_26402 , w_26403 , w_26404 , w_26405 , 
		w_26406 , w_26407 , w_26408 , w_26409 , w_26410 , w_26411 , w_26412 , w_26413 , w_26414 , w_26415 , 
		w_26416 , w_26417 , w_26418 , w_26419 , w_26420 , w_26421 , w_26422 , w_26423 , w_26424 , w_26425 , 
		w_26426 , w_26427 , w_26428 , w_26429 , w_26430 , w_26431 , w_26432 , w_26433 , w_26434 , w_26435 , 
		w_26436 , w_26437 , w_26438 , w_26439 , w_26440 , w_26441 , w_26442 , w_26443 , w_26444 , w_26445 , 
		w_26446 , w_26447 , w_26448 , w_26449 , w_26450 , w_26451 , w_26452 , w_26453 , w_26454 , w_26455 , 
		w_26456 , w_26457 , w_26458 , w_26459 , w_26460 , w_26461 , w_26462 , w_26463 , w_26464 , w_26465 , 
		w_26466 , w_26467 , w_26468 , w_26469 , w_26470 , w_26471 , w_26472 , w_26473 , w_26474 , w_26475 , 
		w_26476 , w_26477 , w_26478 , w_26479 , w_26480 , w_26481 , w_26482 , w_26483 , w_26484 , w_26485 , 
		w_26486 , w_26487 , w_26488 , w_26489 , w_26490 , w_26491 , w_26492 , w_26493 , w_26494 , w_26495 , 
		w_26496 , w_26497 , w_26498 , w_26499 , w_26500 , w_26501 , w_26502 , w_26503 , w_26504 , w_26505 , 
		w_26506 , w_26507 , w_26508 , w_26509 , w_26510 , w_26511 , w_26512 , w_26513 , w_26514 , w_26515 , 
		w_26516 , w_26517 , w_26518 , w_26519 , w_26520 , w_26521 , w_26522 , w_26523 , w_26524 , w_26525 , 
		w_26526 , w_26527 , w_26528 , w_26529 , w_26530 , w_26531 , w_26532 , w_26533 , w_26534 , w_26535 , 
		w_26536 , w_26537 , w_26538 , w_26539 , w_26540 , w_26541 , w_26542 , w_26543 , w_26544 , w_26545 , 
		w_26546 , w_26547 , w_26548 , w_26549 , w_26550 , w_26551 , w_26552 , w_26553 , w_26554 , w_26555 , 
		w_26556 , w_26557 , w_26558 , w_26559 , w_26560 , w_26561 , w_26562 , w_26563 , w_26564 , w_26565 , 
		w_26566 , w_26567 , w_26568 , w_26569 , w_26570 , w_26571 , w_26572 , w_26573 , w_26574 , w_26575 , 
		w_26576 , w_26577 , w_26578 , w_26579 , w_26580 , w_26581 , w_26582 , w_26583 , w_26584 , w_26585 , 
		w_26586 , w_26587 , w_26588 , w_26589 , w_26590 , w_26591 , w_26592 , w_26593 , w_26594 , w_26595 , 
		w_26596 , w_26597 , w_26598 , w_26599 , w_26600 , w_26601 , w_26602 , w_26603 , w_26604 , w_26605 , 
		w_26606 , w_26607 , w_26608 , w_26609 , w_26610 , w_26611 , w_26612 , w_26613 , w_26614 , w_26615 , 
		w_26616 , w_26617 , w_26618 , w_26619 , w_26620 , w_26621 , w_26622 , w_26623 , w_26624 , w_26625 , 
		w_26626 , w_26627 , w_26628 , w_26629 , w_26630 , w_26631 , w_26632 , w_26633 , w_26634 , w_26635 , 
		w_26636 , w_26637 , w_26638 , w_26639 , w_26640 , w_26641 , w_26642 , w_26643 , w_26644 , w_26645 , 
		w_26646 , w_26647 , w_26648 , w_26649 , w_26650 , w_26651 , w_26652 , w_26653 , w_26654 , w_26655 , 
		w_26656 , w_26657 , w_26658 , w_26659 , w_26660 , w_26661 , w_26662 , w_26663 , w_26664 , w_26665 , 
		w_26666 , w_26667 , w_26668 , w_26669 , w_26670 , w_26671 , w_26672 , w_26673 , w_26674 , w_26675 , 
		w_26676 , w_26677 , w_26678 , w_26679 , w_26680 , w_26681 , w_26682 , w_26683 , w_26684 , w_26685 , 
		w_26686 , w_26687 , w_26688 , w_26689 , w_26690 , w_26691 , w_26692 , w_26693 , w_26694 , w_26695 , 
		w_26696 , w_26697 , w_26698 , w_26699 , w_26700 , w_26701 , w_26702 , w_26703 , w_26704 , w_26705 , 
		w_26706 , w_26707 , w_26708 , w_26709 , w_26710 , w_26711 , w_26712 , w_26713 , w_26714 , w_26715 , 
		w_26716 , w_26717 , w_26718 , w_26719 , w_26720 , w_26721 , w_26722 , w_26723 , w_26724 , w_26725 , 
		w_26726 , w_26727 , w_26728 , w_26729 , w_26730 , w_26731 , w_26732 , w_26733 , w_26734 , w_26735 , 
		w_26736 , w_26737 , w_26738 , w_26739 , w_26740 , w_26741 , w_26742 , w_26743 , w_26744 , w_26745 , 
		w_26746 , w_26747 , w_26748 , w_26749 , w_26750 , w_26751 , w_26752 , w_26753 , w_26754 , w_26755 , 
		w_26756 , w_26757 , w_26758 , w_26759 , w_26760 , w_26761 , w_26762 , w_26763 , w_26764 , w_26765 , 
		w_26766 , w_26767 , w_26768 , w_26769 , w_26770 , w_26771 , w_26772 , w_26773 , w_26774 , w_26775 , 
		w_26776 , w_26777 , w_26778 , w_26779 , w_26780 , w_26781 , w_26782 , w_26783 , w_26784 , w_26785 , 
		w_26786 , w_26787 , w_26788 , w_26789 , w_26790 , w_26791 , w_26792 , w_26793 , w_26794 , w_26795 , 
		w_26796 , w_26797 , w_26798 , w_26799 , w_26800 , w_26801 , w_26802 , w_26803 , w_26804 , w_26805 , 
		w_26806 , w_26807 , w_26808 , w_26809 , w_26810 , w_26811 , w_26812 , w_26813 , w_26814 , w_26815 , 
		w_26816 , w_26817 , w_26818 , w_26819 , w_26820 , w_26821 , w_26822 , w_26823 , w_26824 , w_26825 , 
		w_26826 , w_26827 , w_26828 , w_26829 , w_26830 , w_26831 , w_26832 , w_26833 , w_26834 , w_26835 , 
		w_26836 , w_26837 , w_26838 , w_26839 , w_26840 , w_26841 , w_26842 , w_26843 , w_26844 , w_26845 , 
		w_26846 , w_26847 , w_26848 , w_26849 , w_26850 , w_26851 , w_26852 , w_26853 , w_26854 , w_26855 , 
		w_26856 , w_26857 , w_26858 , w_26859 , w_26860 , w_26861 , w_26862 , w_26863 , w_26864 , w_26865 , 
		w_26866 , w_26867 , w_26868 , w_26869 , w_26870 , w_26871 , w_26872 , w_26873 , w_26874 , w_26875 , 
		w_26876 , w_26877 , w_26878 , w_26879 , w_26880 , w_26881 , w_26882 , w_26883 , w_26884 , w_26885 , 
		w_26886 , w_26887 , w_26888 , w_26889 , w_26890 , w_26891 , w_26892 , w_26893 , w_26894 , w_26895 , 
		w_26896 , w_26897 , w_26898 , w_26899 , w_26900 , w_26901 , w_26902 , w_26903 , w_26904 , w_26905 , 
		w_26906 , w_26907 , w_26908 , w_26909 , w_26910 , w_26911 , w_26912 , w_26913 , w_26914 , w_26915 , 
		w_26916 , w_26917 , w_26918 , w_26919 , w_26920 , w_26921 , w_26922 , w_26923 , w_26924 , w_26925 , 
		w_26926 , w_26927 , w_26928 , w_26929 , w_26930 , w_26931 , w_26932 , w_26933 , w_26934 , w_26935 , 
		w_26936 , w_26937 , w_26938 , w_26939 , w_26940 , w_26941 , w_26942 , w_26943 , w_26944 , w_26945 , 
		w_26946 , w_26947 , w_26948 , w_26949 , w_26950 , w_26951 , w_26952 , w_26953 , w_26954 , w_26955 , 
		w_26956 , w_26957 , w_26958 , w_26959 , w_26960 , w_26961 , w_26962 , w_26963 , w_26964 , w_26965 , 
		w_26966 , w_26967 , w_26968 , w_26969 , w_26970 , w_26971 , w_26972 , w_26973 , w_26974 , w_26975 , 
		w_26976 , w_26977 , w_26978 , w_26979 , w_26980 , w_26981 , w_26982 , w_26983 , w_26984 , w_26985 , 
		w_26986 , w_26987 , w_26988 , w_26989 , w_26990 , w_26991 , w_26992 , w_26993 , w_26994 , w_26995 , 
		w_26996 , w_26997 , w_26998 , w_26999 , w_27000 , w_27001 , w_27002 , w_27003 , w_27004 , w_27005 , 
		w_27006 , w_27007 , w_27008 , w_27009 , w_27010 , w_27011 , w_27012 , w_27013 , w_27014 , w_27015 , 
		w_27016 , w_27017 , w_27018 , w_27019 , w_27020 , w_27021 , w_27022 , w_27023 , w_27024 , w_27025 , 
		w_27026 , w_27027 , w_27028 , w_27029 , w_27030 , w_27031 , w_27032 , w_27033 , w_27034 , w_27035 , 
		w_27036 , w_27037 , w_27038 , w_27039 , w_27040 , w_27041 , w_27042 , w_27043 , w_27044 , w_27045 , 
		w_27046 , w_27047 , w_27048 , w_27049 , w_27050 , w_27051 , w_27052 , w_27053 , w_27054 , w_27055 , 
		w_27056 , w_27057 , w_27058 , w_27059 , w_27060 , w_27061 , w_27062 , w_27063 , w_27064 , w_27065 , 
		w_27066 , w_27067 , w_27068 , w_27069 , w_27070 , w_27071 , w_27072 , w_27073 , w_27074 , w_27075 , 
		w_27076 , w_27077 , w_27078 , w_27079 , w_27080 , w_27081 , w_27082 , w_27083 , w_27084 , w_27085 , 
		w_27086 , w_27087 , w_27088 , w_27089 , w_27090 , w_27091 , w_27092 , w_27093 , w_27094 , w_27095 , 
		w_27096 , w_27097 , w_27098 , w_27099 , w_27100 , w_27101 , w_27102 , w_27103 , w_27104 , w_27105 , 
		w_27106 , w_27107 , w_27108 , w_27109 , w_27110 , w_27111 , w_27112 , w_27113 , w_27114 , w_27115 , 
		w_27116 , w_27117 , w_27118 , w_27119 , w_27120 , w_27121 , w_27122 , w_27123 , w_27124 , w_27125 , 
		w_27126 , w_27127 , w_27128 , w_27129 , w_27130 , w_27131 , w_27132 , w_27133 , w_27134 , w_27135 , 
		w_27136 , w_27137 , w_27138 , w_27139 , w_27140 , w_27141 , w_27142 , w_27143 , w_27144 , w_27145 , 
		w_27146 , w_27147 , w_27148 , w_27149 , w_27150 , w_27151 , w_27152 , w_27153 , w_27154 , w_27155 , 
		w_27156 , w_27157 , w_27158 , w_27159 , w_27160 , w_27161 , w_27162 , w_27163 , w_27164 , w_27165 , 
		w_27166 , w_27167 , w_27168 , w_27169 , w_27170 , w_27171 , w_27172 , w_27173 , w_27174 , w_27175 , 
		w_27176 , w_27177 , w_27178 , w_27179 , w_27180 , w_27181 , w_27182 , w_27183 , w_27184 , w_27185 , 
		w_27186 , w_27187 , w_27188 , w_27189 , w_27190 , w_27191 , w_27192 , w_27193 , w_27194 , w_27195 , 
		w_27196 , w_27197 , w_27198 , w_27199 , w_27200 , w_27201 , w_27202 , w_27203 , w_27204 , w_27205 , 
		w_27206 , w_27207 , w_27208 , w_27209 , w_27210 , w_27211 , w_27212 , w_27213 , w_27214 , w_27215 , 
		w_27216 , w_27217 , w_27218 , w_27219 , w_27220 , w_27221 , w_27222 , w_27223 , w_27224 , w_27225 , 
		w_27226 , w_27227 , w_27228 , w_27229 , w_27230 , w_27231 , w_27232 , w_27233 , w_27234 , w_27235 , 
		w_27236 , w_27237 , w_27238 , w_27239 , w_27240 , w_27241 , w_27242 , w_27243 , w_27244 , w_27245 , 
		w_27246 , w_27247 , w_27248 , w_27249 , w_27250 , w_27251 , w_27252 , w_27253 , w_27254 , w_27255 , 
		w_27256 , w_27257 , w_27258 , w_27259 , w_27260 , w_27261 , w_27262 , w_27263 , w_27264 , w_27265 , 
		w_27266 , w_27267 , w_27268 , w_27269 , w_27270 , w_27271 , w_27272 , w_27273 , w_27274 , w_27275 , 
		w_27276 , w_27277 , w_27278 , w_27279 , w_27280 , w_27281 , w_27282 , w_27283 , w_27284 , w_27285 , 
		w_27286 , w_27287 , w_27288 , w_27289 , w_27290 , w_27291 , w_27292 , w_27293 , w_27294 , w_27295 , 
		w_27296 , w_27297 , w_27298 , w_27299 , w_27300 , w_27301 , w_27302 , w_27303 , w_27304 , w_27305 , 
		w_27306 , w_27307 , w_27308 , w_27309 , w_27310 , w_27311 , w_27312 , w_27313 , w_27314 , w_27315 , 
		w_27316 , w_27317 , w_27318 , w_27319 , w_27320 , w_27321 , w_27322 , w_27323 , w_27324 , w_27325 , 
		w_27326 , w_27327 , w_27328 , w_27329 , w_27330 , w_27331 , w_27332 , w_27333 , w_27334 , w_27335 , 
		w_27336 , w_27337 , w_27338 , w_27339 , w_27340 , w_27341 , w_27342 , w_27343 , w_27344 , w_27345 , 
		w_27346 , w_27347 , w_27348 , w_27349 , w_27350 , w_27351 , w_27352 , w_27353 , w_27354 , w_27355 , 
		w_27356 , w_27357 , w_27358 , w_27359 , w_27360 , w_27361 , w_27362 , w_27363 , w_27364 , w_27365 , 
		w_27366 , w_27367 , w_27368 , w_27369 , w_27370 , w_27371 , w_27372 , w_27373 , w_27374 , w_27375 , 
		w_27376 , w_27377 , w_27378 , w_27379 , w_27380 , w_27381 , w_27382 , w_27383 , w_27384 , w_27385 , 
		w_27386 , w_27387 , w_27388 , w_27389 , w_27390 , w_27391 , w_27392 , w_27393 , w_27394 , w_27395 , 
		w_27396 , w_27397 , w_27398 , w_27399 , w_27400 , w_27401 , w_27402 , w_27403 , w_27404 , w_27405 , 
		w_27406 , w_27407 , w_27408 , w_27409 , w_27410 , w_27411 , w_27412 , w_27413 , w_27414 , w_27415 , 
		w_27416 , w_27417 , w_27418 , w_27419 , w_27420 , w_27421 , w_27422 , w_27423 , w_27424 , w_27425 , 
		w_27426 , w_27427 , w_27428 , w_27429 , w_27430 , w_27431 , w_27432 , w_27433 , w_27434 , w_27435 , 
		w_27436 , w_27437 , w_27438 , w_27439 , w_27440 , w_27441 , w_27442 , w_27443 , w_27444 , w_27445 , 
		w_27446 , w_27447 , w_27448 , w_27449 , w_27450 , w_27451 , w_27452 , w_27453 , w_27454 , w_27455 , 
		w_27456 , w_27457 , w_27458 , w_27459 , w_27460 , w_27461 , w_27462 , w_27463 , w_27464 , w_27465 , 
		w_27466 , w_27467 , w_27468 , w_27469 , w_27470 , w_27471 , w_27472 , w_27473 , w_27474 , w_27475 , 
		w_27476 , w_27477 , w_27478 , w_27479 , w_27480 , w_27481 , w_27482 , w_27483 , w_27484 , w_27485 , 
		w_27486 , w_27487 , w_27488 , w_27489 , w_27490 , w_27491 , w_27492 , w_27493 , w_27494 , w_27495 , 
		w_27496 , w_27497 , w_27498 , w_27499 , w_27500 , w_27501 , w_27502 , w_27503 , w_27504 , w_27505 , 
		w_27506 , w_27507 , w_27508 , w_27509 , w_27510 , w_27511 , w_27512 , w_27513 , w_27514 , w_27515 , 
		w_27516 , w_27517 , w_27518 , w_27519 , w_27520 , w_27521 , w_27522 , w_27523 , w_27524 , w_27525 , 
		w_27526 , w_27527 , w_27528 , w_27529 , w_27530 , w_27531 , w_27532 , w_27533 , w_27534 , w_27535 , 
		w_27536 , w_27537 , w_27538 , w_27539 , w_27540 , w_27541 , w_27542 , w_27543 , w_27544 , w_27545 , 
		w_27546 , w_27547 , w_27548 , w_27549 , w_27550 , w_27551 , w_27552 , w_27553 , w_27554 , w_27555 , 
		w_27556 , w_27557 , w_27558 , w_27559 , w_27560 , w_27561 , w_27562 , w_27563 , w_27564 , w_27565 , 
		w_27566 , w_27567 , w_27568 , w_27569 , w_27570 , w_27571 , w_27572 , w_27573 , w_27574 , w_27575 , 
		w_27576 , w_27577 , w_27578 , w_27579 , w_27580 , w_27581 , w_27582 , w_27583 , w_27584 , w_27585 , 
		w_27586 , w_27587 , w_27588 , w_27589 , w_27590 , w_27591 , w_27592 , w_27593 , w_27594 , w_27595 , 
		w_27596 , w_27597 , w_27598 , w_27599 , w_27600 , w_27601 , w_27602 , w_27603 , w_27604 , w_27605 , 
		w_27606 , w_27607 , w_27608 , w_27609 , w_27610 , w_27611 , w_27612 , w_27613 , w_27614 , w_27615 , 
		w_27616 , w_27617 , w_27618 , w_27619 , w_27620 , w_27621 , w_27622 , w_27623 , w_27624 , w_27625 , 
		w_27626 , w_27627 , w_27628 , w_27629 , w_27630 , w_27631 , w_27632 , w_27633 , w_27634 , w_27635 , 
		w_27636 , w_27637 , w_27638 , w_27639 , w_27640 , w_27641 , w_27642 , w_27643 , w_27644 , w_27645 , 
		w_27646 , w_27647 , w_27648 , w_27649 , w_27650 , w_27651 , w_27652 , w_27653 , w_27654 , w_27655 , 
		w_27656 , w_27657 , w_27658 , w_27659 , w_27660 , w_27661 , w_27662 , w_27663 , w_27664 , w_27665 , 
		w_27666 , w_27667 , w_27668 , w_27669 , w_27670 , w_27671 , w_27672 , w_27673 , w_27674 , w_27675 , 
		w_27676 , w_27677 , w_27678 , w_27679 , w_27680 , w_27681 , w_27682 , w_27683 , w_27684 , w_27685 , 
		w_27686 , w_27687 , w_27688 , w_27689 , w_27690 , w_27691 , w_27692 , w_27693 , w_27694 , w_27695 , 
		w_27696 , w_27697 , w_27698 , w_27699 , w_27700 , w_27701 , w_27702 , w_27703 , w_27704 , w_27705 , 
		w_27706 , w_27707 , w_27708 , w_27709 , w_27710 , w_27711 , w_27712 , w_27713 , w_27714 , w_27715 , 
		w_27716 , w_27717 , w_27718 , w_27719 , w_27720 , w_27721 , w_27722 , w_27723 , w_27724 , w_27725 , 
		w_27726 , w_27727 , w_27728 , w_27729 , w_27730 , w_27731 , w_27732 , w_27733 , w_27734 , w_27735 , 
		w_27736 , w_27737 , w_27738 , w_27739 , w_27740 , w_27741 , w_27742 , w_27743 , w_27744 , w_27745 , 
		w_27746 , w_27747 , w_27748 , w_27749 , w_27750 , w_27751 , w_27752 , w_27753 , w_27754 , w_27755 , 
		w_27756 , w_27757 , w_27758 , w_27759 , w_27760 , w_27761 , w_27762 , w_27763 , w_27764 , w_27765 , 
		w_27766 , w_27767 , w_27768 , w_27769 , w_27770 , w_27771 , w_27772 , w_27773 , w_27774 , w_27775 , 
		w_27776 , w_27777 , w_27778 , w_27779 , w_27780 , w_27781 , w_27782 , w_27783 , w_27784 , w_27785 , 
		w_27786 , w_27787 , w_27788 , w_27789 , w_27790 , w_27791 , w_27792 , w_27793 , w_27794 , w_27795 , 
		w_27796 , w_27797 , w_27798 , w_27799 , w_27800 , w_27801 , w_27802 , w_27803 , w_27804 , w_27805 , 
		w_27806 , w_27807 , w_27808 , w_27809 , w_27810 , w_27811 , w_27812 , w_27813 , w_27814 , w_27815 , 
		w_27816 , w_27817 , w_27818 , w_27819 , w_27820 , w_27821 , w_27822 , w_27823 , w_27824 , w_27825 , 
		w_27826 , w_27827 , w_27828 , w_27829 , w_27830 , w_27831 , w_27832 , w_27833 , w_27834 , w_27835 , 
		w_27836 , w_27837 , w_27838 , w_27839 , w_27840 , w_27841 , w_27842 , w_27843 , w_27844 , w_27845 , 
		w_27846 , w_27847 , w_27848 , w_27849 , w_27850 , w_27851 , w_27852 , w_27853 , w_27854 , w_27855 , 
		w_27856 , w_27857 , w_27858 , w_27859 , w_27860 , w_27861 , w_27862 , w_27863 , w_27864 , w_27865 , 
		w_27866 , w_27867 , w_27868 , w_27869 , w_27870 , w_27871 , w_27872 , w_27873 , w_27874 , w_27875 , 
		w_27876 , w_27877 , w_27878 , w_27879 , w_27880 , w_27881 , w_27882 , w_27883 , w_27884 , w_27885 , 
		w_27886 , w_27887 , w_27888 , w_27889 , w_27890 , w_27891 , w_27892 , w_27893 , w_27894 , w_27895 , 
		w_27896 , w_27897 , w_27898 , w_27899 , w_27900 , w_27901 , w_27902 , w_27903 , w_27904 , w_27905 , 
		w_27906 , w_27907 , w_27908 , w_27909 , w_27910 , w_27911 , w_27912 , w_27913 , w_27914 , w_27915 , 
		w_27916 , w_27917 , w_27918 , w_27919 , w_27920 , w_27921 , w_27922 , w_27923 , w_27924 , w_27925 , 
		w_27926 , w_27927 , w_27928 , w_27929 , w_27930 , w_27931 , w_27932 , w_27933 , w_27934 , w_27935 , 
		w_27936 , w_27937 , w_27938 , w_27939 , w_27940 , w_27941 , w_27942 , w_27943 , w_27944 , w_27945 , 
		w_27946 , w_27947 , w_27948 , w_27949 , w_27950 , w_27951 , w_27952 , w_27953 , w_27954 , w_27955 , 
		w_27956 , w_27957 , w_27958 , w_27959 , w_27960 , w_27961 , w_27962 , w_27963 , w_27964 , w_27965 , 
		w_27966 , w_27967 , w_27968 , w_27969 , w_27970 , w_27971 , w_27972 , w_27973 , w_27974 , w_27975 , 
		w_27976 , w_27977 , w_27978 , w_27979 , w_27980 , w_27981 , w_27982 , w_27983 , w_27984 , w_27985 , 
		w_27986 , w_27987 , w_27988 , w_27989 , w_27990 , w_27991 , w_27992 , w_27993 , w_27994 , w_27995 , 
		w_27996 , w_27997 , w_27998 , w_27999 , w_28000 , w_28001 , w_28002 , w_28003 , w_28004 , w_28005 , 
		w_28006 , w_28007 , w_28008 , w_28009 , w_28010 , w_28011 , w_28012 , w_28013 , w_28014 , w_28015 , 
		w_28016 , w_28017 , w_28018 , w_28019 , w_28020 , w_28021 , w_28022 , w_28023 , w_28024 , w_28025 , 
		w_28026 , w_28027 , w_28028 , w_28029 , w_28030 , w_28031 , w_28032 , w_28033 , w_28034 , w_28035 , 
		w_28036 , w_28037 , w_28038 , w_28039 , w_28040 , w_28041 , w_28042 , w_28043 , w_28044 , w_28045 , 
		w_28046 , w_28047 , w_28048 , w_28049 , w_28050 , w_28051 , w_28052 , w_28053 , w_28054 , w_28055 , 
		w_28056 , w_28057 , w_28058 , w_28059 , w_28060 , w_28061 , w_28062 , w_28063 , w_28064 , w_28065 , 
		w_28066 , w_28067 , w_28068 , w_28069 , w_28070 , w_28071 , w_28072 , w_28073 , w_28074 , w_28075 , 
		w_28076 , w_28077 , w_28078 , w_28079 , w_28080 , w_28081 , w_28082 , w_28083 , w_28084 , w_28085 , 
		w_28086 , w_28087 , w_28088 , w_28089 , w_28090 , w_28091 , w_28092 , w_28093 , w_28094 , w_28095 , 
		w_28096 , w_28097 , w_28098 , w_28099 , w_28100 , w_28101 , w_28102 , w_28103 , w_28104 , w_28105 , 
		w_28106 , w_28107 , w_28108 , w_28109 , w_28110 , w_28111 , w_28112 , w_28113 , w_28114 , w_28115 , 
		w_28116 , w_28117 , w_28118 , w_28119 , w_28120 , w_28121 , w_28122 , w_28123 , w_28124 , w_28125 , 
		w_28126 , w_28127 , w_28128 , w_28129 , w_28130 , w_28131 , w_28132 , w_28133 , w_28134 , w_28135 , 
		w_28136 , w_28137 , w_28138 , w_28139 , w_28140 , w_28141 , w_28142 , w_28143 , w_28144 , w_28145 , 
		w_28146 , w_28147 , w_28148 , w_28149 , w_28150 , w_28151 , w_28152 , w_28153 , w_28154 , w_28155 , 
		w_28156 , w_28157 , w_28158 , w_28159 , w_28160 , w_28161 , w_28162 , w_28163 , w_28164 , w_28165 , 
		w_28166 , w_28167 , w_28168 , w_28169 , w_28170 , w_28171 , w_28172 , w_28173 , w_28174 , w_28175 , 
		w_28176 , w_28177 , w_28178 , w_28179 , w_28180 , w_28181 , w_28182 , w_28183 , w_28184 , w_28185 , 
		w_28186 , w_28187 , w_28188 , w_28189 , w_28190 , w_28191 , w_28192 , w_28193 , w_28194 , w_28195 , 
		w_28196 , w_28197 , w_28198 , w_28199 , w_28200 , w_28201 , w_28202 , w_28203 , w_28204 , w_28205 , 
		w_28206 , w_28207 , w_28208 , w_28209 , w_28210 , w_28211 , w_28212 , w_28213 , w_28214 , w_28215 , 
		w_28216 , w_28217 , w_28218 , w_28219 , w_28220 , w_28221 , w_28222 , w_28223 , w_28224 , w_28225 , 
		w_28226 , w_28227 , w_28228 , w_28229 , w_28230 , w_28231 , w_28232 , w_28233 , w_28234 , w_28235 , 
		w_28236 , w_28237 , w_28238 , w_28239 , w_28240 , w_28241 , w_28242 , w_28243 , w_28244 , w_28245 , 
		w_28246 , w_28247 , w_28248 , w_28249 , w_28250 , w_28251 , w_28252 , w_28253 , w_28254 , w_28255 , 
		w_28256 , w_28257 , w_28258 , w_28259 , w_28260 , w_28261 , w_28262 , w_28263 , w_28264 , w_28265 , 
		w_28266 , w_28267 , w_28268 , w_28269 , w_28270 , w_28271 , w_28272 , w_28273 , w_28274 , w_28275 , 
		w_28276 , w_28277 , w_28278 , w_28279 , w_28280 , w_28281 , w_28282 , w_28283 , w_28284 , w_28285 , 
		w_28286 , w_28287 , w_28288 , w_28289 , w_28290 , w_28291 , w_28292 , w_28293 , w_28294 , w_28295 , 
		w_28296 , w_28297 , w_28298 , w_28299 , w_28300 , w_28301 , w_28302 , w_28303 , w_28304 , w_28305 , 
		w_28306 , w_28307 , w_28308 , w_28309 , w_28310 , w_28311 , w_28312 , w_28313 , w_28314 , w_28315 , 
		w_28316 , w_28317 , w_28318 , w_28319 , w_28320 , w_28321 , w_28322 , w_28323 , w_28324 , w_28325 , 
		w_28326 , w_28327 , w_28328 , w_28329 , w_28330 , w_28331 , w_28332 , w_28333 , w_28334 , w_28335 , 
		w_28336 , w_28337 , w_28338 , w_28339 , w_28340 , w_28341 , w_28342 , w_28343 , w_28344 , w_28345 , 
		w_28346 , w_28347 , w_28348 , w_28349 , w_28350 , w_28351 , w_28352 , w_28353 , w_28354 , w_28355 , 
		w_28356 , w_28357 , w_28358 , w_28359 , w_28360 , w_28361 , w_28362 , w_28363 , w_28364 , w_28365 , 
		w_28366 , w_28367 , w_28368 , w_28369 , w_28370 , w_28371 , w_28372 , w_28373 , w_28374 , w_28375 , 
		w_28376 , w_28377 , w_28378 , w_28379 , w_28380 , w_28381 , w_28382 , w_28383 , w_28384 , w_28385 , 
		w_28386 , w_28387 , w_28388 , w_28389 , w_28390 , w_28391 , w_28392 , w_28393 , w_28394 , w_28395 , 
		w_28396 , w_28397 , w_28398 , w_28399 , w_28400 , w_28401 , w_28402 , w_28403 , w_28404 , w_28405 , 
		w_28406 , w_28407 , w_28408 , w_28409 , w_28410 , w_28411 , w_28412 , w_28413 , w_28414 , w_28415 , 
		w_28416 , w_28417 , w_28418 , w_28419 , w_28420 , w_28421 , w_28422 , w_28423 , w_28424 , w_28425 , 
		w_28426 , w_28427 , w_28428 , w_28429 , w_28430 , w_28431 , w_28432 , w_28433 , w_28434 , w_28435 , 
		w_28436 , w_28437 , w_28438 , w_28439 , w_28440 , w_28441 , w_28442 , w_28443 , w_28444 , w_28445 , 
		w_28446 , w_28447 , w_28448 , w_28449 , w_28450 , w_28451 , w_28452 , w_28453 , w_28454 , w_28455 , 
		w_28456 , w_28457 , w_28458 , w_28459 , w_28460 , w_28461 , w_28462 , w_28463 , w_28464 , w_28465 , 
		w_28466 , w_28467 , w_28468 , w_28469 , w_28470 , w_28471 , w_28472 , w_28473 , w_28474 , w_28475 , 
		w_28476 , w_28477 , w_28478 , w_28479 , w_28480 , w_28481 , w_28482 , w_28483 , w_28484 , w_28485 , 
		w_28486 , w_28487 , w_28488 , w_28489 , w_28490 , w_28491 , w_28492 , w_28493 , w_28494 , w_28495 , 
		w_28496 , w_28497 , w_28498 , w_28499 , w_28500 , w_28501 , w_28502 , w_28503 , w_28504 , w_28505 , 
		w_28506 , w_28507 , w_28508 , w_28509 , w_28510 , w_28511 , w_28512 , w_28513 , w_28514 , w_28515 , 
		w_28516 , w_28517 , w_28518 , w_28519 , w_28520 , w_28521 , w_28522 , w_28523 , w_28524 , w_28525 , 
		w_28526 , w_28527 , w_28528 , w_28529 , w_28530 , w_28531 , w_28532 , w_28533 , w_28534 , w_28535 , 
		w_28536 , w_28537 , w_28538 , w_28539 , w_28540 , w_28541 , w_28542 , w_28543 , w_28544 , w_28545 , 
		w_28546 , w_28547 , w_28548 , w_28549 , w_28550 , w_28551 , w_28552 , w_28553 , w_28554 , w_28555 , 
		w_28556 , w_28557 , w_28558 , w_28559 , w_28560 , w_28561 , w_28562 , w_28563 , w_28564 , w_28565 , 
		w_28566 , w_28567 , w_28568 , w_28569 , w_28570 , w_28571 , w_28572 , w_28573 , w_28574 , w_28575 , 
		w_28576 , w_28577 , w_28578 , w_28579 , w_28580 , w_28581 , w_28582 , w_28583 , w_28584 , w_28585 , 
		w_28586 , w_28587 , w_28588 , w_28589 , w_28590 , w_28591 , w_28592 , w_28593 , w_28594 , w_28595 , 
		w_28596 , w_28597 , w_28598 , w_28599 , w_28600 , w_28601 , w_28602 , w_28603 , w_28604 , w_28605 , 
		w_28606 , w_28607 , w_28608 , w_28609 , w_28610 , w_28611 , w_28612 , w_28613 , w_28614 , w_28615 , 
		w_28616 , w_28617 , w_28618 , w_28619 , w_28620 , w_28621 , w_28622 , w_28623 , w_28624 , w_28625 , 
		w_28626 , w_28627 , w_28628 , w_28629 , w_28630 , w_28631 , w_28632 , w_28633 , w_28634 , w_28635 , 
		w_28636 , w_28637 , w_28638 , w_28639 , w_28640 , w_28641 , w_28642 , w_28643 , w_28644 , w_28645 , 
		w_28646 , w_28647 , w_28648 , w_28649 , w_28650 , w_28651 , w_28652 , w_28653 , w_28654 , w_28655 , 
		w_28656 , w_28657 , w_28658 , w_28659 , w_28660 , w_28661 , w_28662 , w_28663 , w_28664 , w_28665 , 
		w_28666 , w_28667 , w_28668 , w_28669 , w_28670 , w_28671 , w_28672 , w_28673 , w_28674 , w_28675 , 
		w_28676 , w_28677 , w_28678 , w_28679 , w_28680 , w_28681 , w_28682 , w_28683 , w_28684 , w_28685 , 
		w_28686 , w_28687 , w_28688 , w_28689 , w_28690 , w_28691 , w_28692 , w_28693 , w_28694 , w_28695 , 
		w_28696 , w_28697 , w_28698 , w_28699 , w_28700 , w_28701 , w_28702 , w_28703 , w_28704 , w_28705 , 
		w_28706 , w_28707 , w_28708 , w_28709 , w_28710 , w_28711 , w_28712 , w_28713 , w_28714 , w_28715 , 
		w_28716 , w_28717 , w_28718 , w_28719 , w_28720 , w_28721 , w_28722 , w_28723 , w_28724 , w_28725 , 
		w_28726 , w_28727 , w_28728 , w_28729 , w_28730 , w_28731 , w_28732 , w_28733 , w_28734 , w_28735 , 
		w_28736 , w_28737 , w_28738 , w_28739 , w_28740 , w_28741 , w_28742 , w_28743 , w_28744 , w_28745 , 
		w_28746 , w_28747 , w_28748 , w_28749 , w_28750 , w_28751 , w_28752 , w_28753 , w_28754 , w_28755 , 
		w_28756 , w_28757 , w_28758 , w_28759 , w_28760 , w_28761 , w_28762 , w_28763 , w_28764 , w_28765 , 
		w_28766 , w_28767 , w_28768 , w_28769 , w_28770 , w_28771 , w_28772 , w_28773 , w_28774 , w_28775 , 
		w_28776 , w_28777 , w_28778 , w_28779 , w_28780 , w_28781 , w_28782 , w_28783 , w_28784 , w_28785 , 
		w_28786 , w_28787 , w_28788 , w_28789 , w_28790 , w_28791 , w_28792 , w_28793 , w_28794 , w_28795 , 
		w_28796 , w_28797 , w_28798 , w_28799 , w_28800 , w_28801 , w_28802 , w_28803 , w_28804 , w_28805 , 
		w_28806 , w_28807 , w_28808 , w_28809 , w_28810 , w_28811 , w_28812 , w_28813 , w_28814 , w_28815 , 
		w_28816 , w_28817 , w_28818 , w_28819 , w_28820 , w_28821 , w_28822 , w_28823 , w_28824 , w_28825 , 
		w_28826 , w_28827 , w_28828 , w_28829 , w_28830 , w_28831 , w_28832 , w_28833 , w_28834 , w_28835 , 
		w_28836 , w_28837 , w_28838 , w_28839 , w_28840 , w_28841 , w_28842 , w_28843 , w_28844 , w_28845 , 
		w_28846 , w_28847 , w_28848 , w_28849 , w_28850 , w_28851 , w_28852 , w_28853 , w_28854 , w_28855 , 
		w_28856 , w_28857 , w_28858 , w_28859 , w_28860 , w_28861 , w_28862 , w_28863 , w_28864 , w_28865 , 
		w_28866 , w_28867 , w_28868 , w_28869 , w_28870 , w_28871 , w_28872 , w_28873 , w_28874 , w_28875 , 
		w_28876 , w_28877 , w_28878 , w_28879 , w_28880 , w_28881 , w_28882 , w_28883 , w_28884 , w_28885 , 
		w_28886 , w_28887 , w_28888 , w_28889 , w_28890 , w_28891 , w_28892 , w_28893 , w_28894 , w_28895 , 
		w_28896 , w_28897 , w_28898 , w_28899 , w_28900 , w_28901 , w_28902 , w_28903 , w_28904 , w_28905 , 
		w_28906 , w_28907 , w_28908 , w_28909 , w_28910 , w_28911 , w_28912 , w_28913 , w_28914 , w_28915 , 
		w_28916 , w_28917 , w_28918 , w_28919 , w_28920 , w_28921 , w_28922 , w_28923 , w_28924 , w_28925 , 
		w_28926 , w_28927 , w_28928 , w_28929 , w_28930 , w_28931 , w_28932 , w_28933 , w_28934 , w_28935 , 
		w_28936 , w_28937 , w_28938 , w_28939 , w_28940 , w_28941 , w_28942 , w_28943 , w_28944 , w_28945 , 
		w_28946 , w_28947 , w_28948 , w_28949 , w_28950 , w_28951 , w_28952 , w_28953 , w_28954 , w_28955 , 
		w_28956 , w_28957 , w_28958 , w_28959 , w_28960 , w_28961 , w_28962 , w_28963 , w_28964 , w_28965 , 
		w_28966 , w_28967 , w_28968 , w_28969 , w_28970 , w_28971 , w_28972 , w_28973 , w_28974 , w_28975 , 
		w_28976 , w_28977 , w_28978 , w_28979 , w_28980 , w_28981 , w_28982 , w_28983 , w_28984 , w_28985 , 
		w_28986 , w_28987 , w_28988 , w_28989 , w_28990 , w_28991 , w_28992 , w_28993 , w_28994 , w_28995 , 
		w_28996 , w_28997 , w_28998 , w_28999 , w_29000 , w_29001 , w_29002 , w_29003 , w_29004 , w_29005 , 
		w_29006 , w_29007 , w_29008 , w_29009 , w_29010 , w_29011 , w_29012 , w_29013 , w_29014 , w_29015 , 
		w_29016 , w_29017 , w_29018 , w_29019 , w_29020 , w_29021 , w_29022 , w_29023 , w_29024 , w_29025 , 
		w_29026 , w_29027 , w_29028 , w_29029 , w_29030 , w_29031 , w_29032 , w_29033 , w_29034 , w_29035 , 
		w_29036 , w_29037 , w_29038 , w_29039 , w_29040 , w_29041 , w_29042 , w_29043 , w_29044 , w_29045 , 
		w_29046 , w_29047 , w_29048 , w_29049 , w_29050 , w_29051 , w_29052 , w_29053 , w_29054 , w_29055 , 
		w_29056 , w_29057 , w_29058 , w_29059 , w_29060 , w_29061 , w_29062 , w_29063 , w_29064 , w_29065 , 
		w_29066 , w_29067 , w_29068 , w_29069 , w_29070 , w_29071 , w_29072 , w_29073 , w_29074 , w_29075 , 
		w_29076 , w_29077 , w_29078 , w_29079 , w_29080 , w_29081 , w_29082 , w_29083 , w_29084 , w_29085 , 
		w_29086 , w_29087 , w_29088 , w_29089 , w_29090 , w_29091 , w_29092 , w_29093 , w_29094 , w_29095 , 
		w_29096 , w_29097 , w_29098 , w_29099 , w_29100 , w_29101 , w_29102 , w_29103 , w_29104 , w_29105 , 
		w_29106 , w_29107 , w_29108 , w_29109 , w_29110 , w_29111 , w_29112 , w_29113 , w_29114 , w_29115 , 
		w_29116 , w_29117 , w_29118 , w_29119 , w_29120 , w_29121 , w_29122 , w_29123 , w_29124 , w_29125 , 
		w_29126 , w_29127 , w_29128 , w_29129 , w_29130 , w_29131 , w_29132 , w_29133 , w_29134 , w_29135 , 
		w_29136 , w_29137 , w_29138 , w_29139 , w_29140 , w_29141 , w_29142 , w_29143 , w_29144 , w_29145 , 
		w_29146 , w_29147 , w_29148 , w_29149 , w_29150 , w_29151 , w_29152 , w_29153 , w_29154 , w_29155 , 
		w_29156 , w_29157 , w_29158 , w_29159 , w_29160 , w_29161 , w_29162 , w_29163 , w_29164 , w_29165 , 
		w_29166 , w_29167 , w_29168 , w_29169 , w_29170 , w_29171 , w_29172 , w_29173 , w_29174 , w_29175 , 
		w_29176 , w_29177 , w_29178 , w_29179 , w_29180 , w_29181 , w_29182 , w_29183 , w_29184 , w_29185 , 
		w_29186 , w_29187 , w_29188 , w_29189 , w_29190 , w_29191 , w_29192 , w_29193 , w_29194 , w_29195 , 
		w_29196 , w_29197 , w_29198 , w_29199 , w_29200 , w_29201 , w_29202 , w_29203 , w_29204 , w_29205 , 
		w_29206 , w_29207 , w_29208 , w_29209 , w_29210 , w_29211 , w_29212 , w_29213 , w_29214 , w_29215 , 
		w_29216 , w_29217 , w_29218 , w_29219 , w_29220 , w_29221 , w_29222 , w_29223 , w_29224 , w_29225 , 
		w_29226 , w_29227 , w_29228 , w_29229 , w_29230 , w_29231 , w_29232 , w_29233 , w_29234 , w_29235 , 
		w_29236 , w_29237 , w_29238 , w_29239 , w_29240 , w_29241 , w_29242 , w_29243 , w_29244 , w_29245 , 
		w_29246 , w_29247 , w_29248 , w_29249 , w_29250 , w_29251 , w_29252 , w_29253 , w_29254 , w_29255 , 
		w_29256 , w_29257 , w_29258 , w_29259 , w_29260 , w_29261 , w_29262 , w_29263 , w_29264 , w_29265 , 
		w_29266 , w_29267 , w_29268 , w_29269 , w_29270 , w_29271 , w_29272 , w_29273 , w_29274 , w_29275 , 
		w_29276 , w_29277 , w_29278 , w_29279 , w_29280 , w_29281 , w_29282 , w_29283 , w_29284 , w_29285 , 
		w_29286 , w_29287 , w_29288 , w_29289 , w_29290 , w_29291 , w_29292 , w_29293 , w_29294 , w_29295 , 
		w_29296 , w_29297 , w_29298 , w_29299 , w_29300 , w_29301 , w_29302 , w_29303 , w_29304 , w_29305 , 
		w_29306 , w_29307 , w_29308 , w_29309 , w_29310 , w_29311 , w_29312 , w_29313 , w_29314 , w_29315 , 
		w_29316 , w_29317 , w_29318 , w_29319 , w_29320 , w_29321 , w_29322 , w_29323 , w_29324 , w_29325 , 
		w_29326 , w_29327 , w_29328 , w_29329 , w_29330 , w_29331 , w_29332 , w_29333 , w_29334 , w_29335 , 
		w_29336 , w_29337 , w_29338 , w_29339 , w_29340 , w_29341 , w_29342 , w_29343 , w_29344 , w_29345 , 
		w_29346 , w_29347 , w_29348 , w_29349 , w_29350 , w_29351 , w_29352 , w_29353 , w_29354 , w_29355 , 
		w_29356 , w_29357 , w_29358 , w_29359 , w_29360 , w_29361 , w_29362 , w_29363 , w_29364 , w_29365 , 
		w_29366 , w_29367 , w_29368 , w_29369 , w_29370 , w_29371 , w_29372 , w_29373 , w_29374 , w_29375 , 
		w_29376 , w_29377 , w_29378 , w_29379 , w_29380 , w_29381 , w_29382 , w_29383 , w_29384 , w_29385 , 
		w_29386 , w_29387 , w_29388 , w_29389 , w_29390 , w_29391 , w_29392 , w_29393 , w_29394 , w_29395 , 
		w_29396 , w_29397 , w_29398 , w_29399 , w_29400 , w_29401 , w_29402 , w_29403 , w_29404 , w_29405 , 
		w_29406 , w_29407 , w_29408 , w_29409 , w_29410 , w_29411 , w_29412 , w_29413 , w_29414 , w_29415 , 
		w_29416 , w_29417 , w_29418 , w_29419 , w_29420 , w_29421 , w_29422 , w_29423 , w_29424 , w_29425 , 
		w_29426 , w_29427 , w_29428 , w_29429 , w_29430 , w_29431 , w_29432 , w_29433 , w_29434 , w_29435 , 
		w_29436 , w_29437 , w_29438 , w_29439 , w_29440 , w_29441 , w_29442 , w_29443 , w_29444 , w_29445 , 
		w_29446 , w_29447 , w_29448 , w_29449 , w_29450 , w_29451 , w_29452 , w_29453 , w_29454 , w_29455 , 
		w_29456 , w_29457 , w_29458 , w_29459 , w_29460 , w_29461 , w_29462 , w_29463 , w_29464 , w_29465 , 
		w_29466 , w_29467 , w_29468 , w_29469 , w_29470 , w_29471 , w_29472 , w_29473 , w_29474 , w_29475 , 
		w_29476 , w_29477 , w_29478 , w_29479 , w_29480 , w_29481 , w_29482 , w_29483 , w_29484 , w_29485 , 
		w_29486 , w_29487 , w_29488 , w_29489 , w_29490 , w_29491 , w_29492 , w_29493 , w_29494 , w_29495 , 
		w_29496 , w_29497 , w_29498 , w_29499 , w_29500 , w_29501 , w_29502 , w_29503 , w_29504 , w_29505 , 
		w_29506 , w_29507 , w_29508 , w_29509 , w_29510 , w_29511 , w_29512 , w_29513 , w_29514 , w_29515 , 
		w_29516 , w_29517 , w_29518 , w_29519 , w_29520 , w_29521 , w_29522 , w_29523 , w_29524 , w_29525 , 
		w_29526 , w_29527 , w_29528 , w_29529 , w_29530 , w_29531 , w_29532 , w_29533 , w_29534 , w_29535 , 
		w_29536 , w_29537 , w_29538 , w_29539 , w_29540 , w_29541 , w_29542 , w_29543 , w_29544 , w_29545 , 
		w_29546 , w_29547 , w_29548 , w_29549 , w_29550 , w_29551 , w_29552 , w_29553 , w_29554 , w_29555 , 
		w_29556 , w_29557 , w_29558 , w_29559 , w_29560 , w_29561 , w_29562 , w_29563 , w_29564 , w_29565 , 
		w_29566 , w_29567 , w_29568 , w_29569 , w_29570 , w_29571 , w_29572 , w_29573 , w_29574 , w_29575 , 
		w_29576 , w_29577 , w_29578 , w_29579 , w_29580 , w_29581 , w_29582 , w_29583 , w_29584 , w_29585 , 
		w_29586 , w_29587 , w_29588 , w_29589 , w_29590 , w_29591 , w_29592 , w_29593 , w_29594 , w_29595 , 
		w_29596 , w_29597 , w_29598 , w_29599 , w_29600 , w_29601 , w_29602 , w_29603 , w_29604 , w_29605 , 
		w_29606 , w_29607 , w_29608 , w_29609 , w_29610 , w_29611 , w_29612 , w_29613 , w_29614 , w_29615 , 
		w_29616 , w_29617 , w_29618 , w_29619 , w_29620 , w_29621 , w_29622 , w_29623 , w_29624 , w_29625 , 
		w_29626 , w_29627 , w_29628 , w_29629 , w_29630 , w_29631 , w_29632 , w_29633 , w_29634 , w_29635 , 
		w_29636 , w_29637 , w_29638 , w_29639 , w_29640 , w_29641 , w_29642 , w_29643 , w_29644 , w_29645 , 
		w_29646 , w_29647 , w_29648 , w_29649 , w_29650 , w_29651 , w_29652 , w_29653 , w_29654 , w_29655 , 
		w_29656 , w_29657 , w_29658 , w_29659 , w_29660 , w_29661 , w_29662 , w_29663 , w_29664 , w_29665 , 
		w_29666 , w_29667 , w_29668 , w_29669 , w_29670 , w_29671 , w_29672 , w_29673 , w_29674 , w_29675 , 
		w_29676 , w_29677 , w_29678 , w_29679 , w_29680 , w_29681 , w_29682 , w_29683 , w_29684 , w_29685 , 
		w_29686 , w_29687 , w_29688 , w_29689 , w_29690 , w_29691 , w_29692 , w_29693 , w_29694 , w_29695 , 
		w_29696 , w_29697 , w_29698 , w_29699 , w_29700 , w_29701 , w_29702 , w_29703 , w_29704 , w_29705 , 
		w_29706 , w_29707 , w_29708 , w_29709 , w_29710 , w_29711 , w_29712 , w_29713 , w_29714 , w_29715 , 
		w_29716 , w_29717 , w_29718 , w_29719 , w_29720 , w_29721 , w_29722 , w_29723 , w_29724 , w_29725 , 
		w_29726 , w_29727 , w_29728 , w_29729 , w_29730 , w_29731 , w_29732 , w_29733 , w_29734 , w_29735 , 
		w_29736 , w_29737 , w_29738 , w_29739 , w_29740 , w_29741 , w_29742 , w_29743 , w_29744 , w_29745 , 
		w_29746 , w_29747 , w_29748 , w_29749 , w_29750 , w_29751 , w_29752 , w_29753 , w_29754 , w_29755 , 
		w_29756 , w_29757 , w_29758 , w_29759 , w_29760 , w_29761 , w_29762 , w_29763 , w_29764 , w_29765 , 
		w_29766 , w_29767 , w_29768 , w_29769 , w_29770 , w_29771 , w_29772 , w_29773 , w_29774 , w_29775 , 
		w_29776 , w_29777 , w_29778 , w_29779 , w_29780 , w_29781 , w_29782 , w_29783 , w_29784 , w_29785 , 
		w_29786 , w_29787 , w_29788 , w_29789 , w_29790 , w_29791 , w_29792 , w_29793 , w_29794 , w_29795 , 
		w_29796 , w_29797 , w_29798 , w_29799 , w_29800 , w_29801 , w_29802 , w_29803 , w_29804 , w_29805 , 
		w_29806 , w_29807 , w_29808 , w_29809 , w_29810 , w_29811 , w_29812 , w_29813 , w_29814 , w_29815 , 
		w_29816 , w_29817 , w_29818 , w_29819 , w_29820 , w_29821 , w_29822 , w_29823 , w_29824 , w_29825 , 
		w_29826 , w_29827 , w_29828 , w_29829 , w_29830 , w_29831 , w_29832 , w_29833 , w_29834 , w_29835 , 
		w_29836 , w_29837 , w_29838 , w_29839 , w_29840 , w_29841 , w_29842 , w_29843 , w_29844 , w_29845 , 
		w_29846 , w_29847 , w_29848 , w_29849 , w_29850 , w_29851 , w_29852 , w_29853 , w_29854 , w_29855 , 
		w_29856 , w_29857 , w_29858 , w_29859 , w_29860 , w_29861 , w_29862 , w_29863 , w_29864 , w_29865 , 
		w_29866 , w_29867 , w_29868 , w_29869 , w_29870 , w_29871 , w_29872 , w_29873 , w_29874 , w_29875 , 
		w_29876 , w_29877 , w_29878 , w_29879 , w_29880 , w_29881 , w_29882 , w_29883 , w_29884 , w_29885 , 
		w_29886 , w_29887 , w_29888 , w_29889 , w_29890 , w_29891 , w_29892 , w_29893 , w_29894 , w_29895 , 
		w_29896 , w_29897 , w_29898 , w_29899 , w_29900 , w_29901 , w_29902 , w_29903 , w_29904 , w_29905 , 
		w_29906 , w_29907 , w_29908 , w_29909 , w_29910 , w_29911 , w_29912 , w_29913 , w_29914 , w_29915 , 
		w_29916 , w_29917 , w_29918 , w_29919 , w_29920 , w_29921 , w_29922 , w_29923 , w_29924 , w_29925 , 
		w_29926 , w_29927 , w_29928 , w_29929 , w_29930 , w_29931 , w_29932 , w_29933 , w_29934 , w_29935 , 
		w_29936 , w_29937 , w_29938 , w_29939 , w_29940 , w_29941 , w_29942 , w_29943 , w_29944 , w_29945 , 
		w_29946 , w_29947 , w_29948 , w_29949 , w_29950 , w_29951 , w_29952 , w_29953 , w_29954 , w_29955 , 
		w_29956 , w_29957 , w_29958 , w_29959 , w_29960 , w_29961 , w_29962 , w_29963 , w_29964 , w_29965 , 
		w_29966 , w_29967 , w_29968 , w_29969 , w_29970 , w_29971 , w_29972 , w_29973 , w_29974 , w_29975 , 
		w_29976 , w_29977 , w_29978 , w_29979 , w_29980 , w_29981 , w_29982 , w_29983 , w_29984 , w_29985 , 
		w_29986 , w_29987 , w_29988 , w_29989 , w_29990 , w_29991 , w_29992 , w_29993 , w_29994 , w_29995 , 
		w_29996 , w_29997 , w_29998 , w_29999 , w_30000 , w_30001 , w_30002 , w_30003 , w_30004 , w_30005 , 
		w_30006 , w_30007 , w_30008 , w_30009 , w_30010 , w_30011 , w_30012 , w_30013 , w_30014 , w_30015 , 
		w_30016 , w_30017 , w_30018 , w_30019 , w_30020 , w_30021 , w_30022 , w_30023 , w_30024 , w_30025 , 
		w_30026 , w_30027 , w_30028 , w_30029 , w_30030 , w_30031 , w_30032 , w_30033 , w_30034 , w_30035 , 
		w_30036 , w_30037 , w_30038 , w_30039 , w_30040 , w_30041 , w_30042 , w_30043 , w_30044 , w_30045 , 
		w_30046 , w_30047 , w_30048 , w_30049 , w_30050 , w_30051 , w_30052 , w_30053 , w_30054 , w_30055 , 
		w_30056 , w_30057 , w_30058 , w_30059 , w_30060 , w_30061 , w_30062 , w_30063 , w_30064 , w_30065 , 
		w_30066 , w_30067 , w_30068 , w_30069 , w_30070 , w_30071 , w_30072 , w_30073 , w_30074 , w_30075 , 
		w_30076 , w_30077 , w_30078 , w_30079 , w_30080 , w_30081 , w_30082 , w_30083 , w_30084 , w_30085 , 
		w_30086 , w_30087 , w_30088 , w_30089 , w_30090 , w_30091 , w_30092 , w_30093 , w_30094 , w_30095 , 
		w_30096 , w_30097 , w_30098 , w_30099 , w_30100 , w_30101 , w_30102 , w_30103 , w_30104 , w_30105 , 
		w_30106 , w_30107 , w_30108 , w_30109 , w_30110 , w_30111 , w_30112 , w_30113 , w_30114 , w_30115 , 
		w_30116 , w_30117 , w_30118 , w_30119 , w_30120 , w_30121 , w_30122 , w_30123 , w_30124 , w_30125 , 
		w_30126 , w_30127 , w_30128 , w_30129 , w_30130 , w_30131 , w_30132 , w_30133 , w_30134 , w_30135 , 
		w_30136 , w_30137 , w_30138 , w_30139 , w_30140 , w_30141 , w_30142 , w_30143 , w_30144 , w_30145 , 
		w_30146 , w_30147 , w_30148 , w_30149 , w_30150 , w_30151 , w_30152 , w_30153 , w_30154 , w_30155 , 
		w_30156 , w_30157 , w_30158 , w_30159 , w_30160 , w_30161 , w_30162 , w_30163 , w_30164 , w_30165 , 
		w_30166 , w_30167 , w_30168 , w_30169 , w_30170 , w_30171 , w_30172 , w_30173 , w_30174 , w_30175 , 
		w_30176 , w_30177 , w_30178 , w_30179 , w_30180 , w_30181 , w_30182 , w_30183 , w_30184 , w_30185 , 
		w_30186 , w_30187 , w_30188 , w_30189 , w_30190 , w_30191 , w_30192 , w_30193 , w_30194 , w_30195 , 
		w_30196 , w_30197 , w_30198 , w_30199 , w_30200 , w_30201 , w_30202 , w_30203 , w_30204 , w_30205 , 
		w_30206 , w_30207 , w_30208 , w_30209 , w_30210 , w_30211 , w_30212 , w_30213 , w_30214 , w_30215 , 
		w_30216 , w_30217 , w_30218 , w_30219 , w_30220 , w_30221 , w_30222 , w_30223 , w_30224 , w_30225 , 
		w_30226 , w_30227 , w_30228 , w_30229 , w_30230 , w_30231 , w_30232 , w_30233 , w_30234 , w_30235 , 
		w_30236 , w_30237 , w_30238 , w_30239 , w_30240 , w_30241 , w_30242 , w_30243 , w_30244 , w_30245 , 
		w_30246 , w_30247 , w_30248 , w_30249 , w_30250 , w_30251 , w_30252 , w_30253 , w_30254 , w_30255 , 
		w_30256 , w_30257 , w_30258 , w_30259 , w_30260 , w_30261 , w_30262 , w_30263 , w_30264 , w_30265 , 
		w_30266 , w_30267 , w_30268 , w_30269 , w_30270 , w_30271 , w_30272 , w_30273 , w_30274 , w_30275 , 
		w_30276 , w_30277 , w_30278 , w_30279 , w_30280 , w_30281 , w_30282 , w_30283 , w_30284 , w_30285 , 
		w_30286 , w_30287 , w_30288 , w_30289 , w_30290 , w_30291 , w_30292 , w_30293 , w_30294 , w_30295 , 
		w_30296 , w_30297 , w_30298 , w_30299 , w_30300 , w_30301 , w_30302 , w_30303 , w_30304 , w_30305 , 
		w_30306 , w_30307 , w_30308 , w_30309 , w_30310 , w_30311 , w_30312 , w_30313 , w_30314 , w_30315 , 
		w_30316 , w_30317 , w_30318 , w_30319 , w_30320 , w_30321 , w_30322 , w_30323 , w_30324 , w_30325 , 
		w_30326 , w_30327 , w_30328 , w_30329 , w_30330 , w_30331 , w_30332 , w_30333 , w_30334 , w_30335 , 
		w_30336 , w_30337 , w_30338 , w_30339 , w_30340 , w_30341 , w_30342 , w_30343 , w_30344 , w_30345 , 
		w_30346 , w_30347 , w_30348 , w_30349 , w_30350 , w_30351 , w_30352 , w_30353 , w_30354 , w_30355 , 
		w_30356 , w_30357 , w_30358 , w_30359 , w_30360 , w_30361 , w_30362 , w_30363 , w_30364 , w_30365 , 
		w_30366 , w_30367 , w_30368 , w_30369 , w_30370 , w_30371 , w_30372 , w_30373 , w_30374 , w_30375 , 
		w_30376 , w_30377 , w_30378 , w_30379 , w_30380 , w_30381 , w_30382 , w_30383 , w_30384 , w_30385 , 
		w_30386 , w_30387 , w_30388 , w_30389 , w_30390 , w_30391 , w_30392 , w_30393 , w_30394 , w_30395 , 
		w_30396 , w_30397 , w_30398 , w_30399 , w_30400 , w_30401 , w_30402 , w_30403 , w_30404 , w_30405 , 
		w_30406 , w_30407 , w_30408 , w_30409 , w_30410 , w_30411 , w_30412 , w_30413 , w_30414 , w_30415 , 
		w_30416 , w_30417 , w_30418 , w_30419 , w_30420 , w_30421 , w_30422 , w_30423 , w_30424 , w_30425 , 
		w_30426 , w_30427 , w_30428 , w_30429 , w_30430 , w_30431 , w_30432 , w_30433 , w_30434 , w_30435 , 
		w_30436 , w_30437 , w_30438 , w_30439 , w_30440 , w_30441 , w_30442 , w_30443 , w_30444 , w_30445 , 
		w_30446 , w_30447 , w_30448 , w_30449 , w_30450 , w_30451 , w_30452 , w_30453 , w_30454 , w_30455 , 
		w_30456 , w_30457 , w_30458 , w_30459 , w_30460 , w_30461 , w_30462 , w_30463 , w_30464 , w_30465 , 
		w_30466 , w_30467 , w_30468 , w_30469 , w_30470 , w_30471 , w_30472 , w_30473 , w_30474 , w_30475 , 
		w_30476 , w_30477 , w_30478 , w_30479 , w_30480 , w_30481 , w_30482 , w_30483 , w_30484 , w_30485 , 
		w_30486 , w_30487 , w_30488 , w_30489 , w_30490 , w_30491 , w_30492 , w_30493 , w_30494 , w_30495 , 
		w_30496 , w_30497 , w_30498 , w_30499 , w_30500 , w_30501 , w_30502 , w_30503 , w_30504 , w_30505 , 
		w_30506 , w_30507 , w_30508 , w_30509 , w_30510 , w_30511 , w_30512 , w_30513 , w_30514 , w_30515 , 
		w_30516 , w_30517 , w_30518 , w_30519 , w_30520 , w_30521 , w_30522 , w_30523 , w_30524 , w_30525 , 
		w_30526 , w_30527 , w_30528 , w_30529 , w_30530 , w_30531 , w_30532 , w_30533 , w_30534 , w_30535 , 
		w_30536 , w_30537 , w_30538 , w_30539 , w_30540 , w_30541 , w_30542 , w_30543 , w_30544 , w_30545 , 
		w_30546 , w_30547 , w_30548 , w_30549 , w_30550 , w_30551 , w_30552 , w_30553 , w_30554 , w_30555 , 
		w_30556 , w_30557 , w_30558 , w_30559 , w_30560 , w_30561 , w_30562 , w_30563 , w_30564 , w_30565 , 
		w_30566 , w_30567 , w_30568 , w_30569 , w_30570 , w_30571 , w_30572 , w_30573 , w_30574 , w_30575 , 
		w_30576 , w_30577 , w_30578 , w_30579 , w_30580 , w_30581 , w_30582 , w_30583 , w_30584 , w_30585 , 
		w_30586 , w_30587 , w_30588 , w_30589 , w_30590 , w_30591 , w_30592 , w_30593 , w_30594 , w_30595 , 
		w_30596 , w_30597 , w_30598 , w_30599 , w_30600 , w_30601 , w_30602 , w_30603 , w_30604 , w_30605 , 
		w_30606 , w_30607 , w_30608 , w_30609 , w_30610 , w_30611 , w_30612 , w_30613 , w_30614 , w_30615 , 
		w_30616 , w_30617 , w_30618 , w_30619 , w_30620 , w_30621 , w_30622 , w_30623 , w_30624 , w_30625 , 
		w_30626 , w_30627 , w_30628 , w_30629 , w_30630 , w_30631 , w_30632 , w_30633 , w_30634 , w_30635 , 
		w_30636 , w_30637 , w_30638 , w_30639 , w_30640 , w_30641 , w_30642 , w_30643 , w_30644 , w_30645 , 
		w_30646 , w_30647 , w_30648 , w_30649 , w_30650 , w_30651 , w_30652 , w_30653 , w_30654 , w_30655 , 
		w_30656 , w_30657 , w_30658 , w_30659 , w_30660 , w_30661 , w_30662 , w_30663 , w_30664 , w_30665 , 
		w_30666 , w_30667 , w_30668 , w_30669 , w_30670 , w_30671 , w_30672 , w_30673 , w_30674 , w_30675 , 
		w_30676 , w_30677 , w_30678 , w_30679 , w_30680 , w_30681 , w_30682 , w_30683 , w_30684 , w_30685 , 
		w_30686 , w_30687 , w_30688 , w_30689 , w_30690 , w_30691 , w_30692 , w_30693 , w_30694 , w_30695 , 
		w_30696 , w_30697 , w_30698 , w_30699 , w_30700 , w_30701 , w_30702 , w_30703 , w_30704 , w_30705 , 
		w_30706 , w_30707 , w_30708 , w_30709 , w_30710 , w_30711 , w_30712 , w_30713 , w_30714 , w_30715 , 
		w_30716 , w_30717 , w_30718 , w_30719 , w_30720 , w_30721 , w_30722 , w_30723 , w_30724 , w_30725 , 
		w_30726 , w_30727 , w_30728 , w_30729 , w_30730 , w_30731 , w_30732 , w_30733 , w_30734 , w_30735 , 
		w_30736 , w_30737 , w_30738 , w_30739 , w_30740 , w_30741 , w_30742 , w_30743 , w_30744 , w_30745 , 
		w_30746 , w_30747 , w_30748 , w_30749 , w_30750 , w_30751 , w_30752 , w_30753 , w_30754 , w_30755 , 
		w_30756 , w_30757 , w_30758 , w_30759 , w_30760 , w_30761 , w_30762 , w_30763 , w_30764 , w_30765 , 
		w_30766 , w_30767 , w_30768 , w_30769 , w_30770 , w_30771 , w_30772 , w_30773 , w_30774 , w_30775 , 
		w_30776 , w_30777 , w_30778 , w_30779 , w_30780 , w_30781 , w_30782 , w_30783 , w_30784 , w_30785 , 
		w_30786 , w_30787 , w_30788 , w_30789 , w_30790 , w_30791 , w_30792 , w_30793 , w_30794 , w_30795 , 
		w_30796 , w_30797 , w_30798 , w_30799 , w_30800 , w_30801 , w_30802 , w_30803 , w_30804 , w_30805 , 
		w_30806 , w_30807 , w_30808 , w_30809 , w_30810 , w_30811 , w_30812 , w_30813 , w_30814 , w_30815 , 
		w_30816 , w_30817 , w_30818 , w_30819 , w_30820 , w_30821 , w_30822 , w_30823 , w_30824 , w_30825 , 
		w_30826 , w_30827 , w_30828 , w_30829 , w_30830 , w_30831 , w_30832 , w_30833 , w_30834 , w_30835 , 
		w_30836 , w_30837 , w_30838 , w_30839 , w_30840 , w_30841 , w_30842 , w_30843 , w_30844 , w_30845 , 
		w_30846 , w_30847 , w_30848 , w_30849 , w_30850 , w_30851 , w_30852 , w_30853 , w_30854 , w_30855 , 
		w_30856 , w_30857 , w_30858 , w_30859 , w_30860 , w_30861 , w_30862 , w_30863 , w_30864 , w_30865 , 
		w_30866 , w_30867 , w_30868 , w_30869 , w_30870 , w_30871 , w_30872 , w_30873 , w_30874 , w_30875 , 
		w_30876 , w_30877 , w_30878 , w_30879 , w_30880 , w_30881 , w_30882 , w_30883 , w_30884 , w_30885 , 
		w_30886 , w_30887 , w_30888 , w_30889 , w_30890 , w_30891 , w_30892 , w_30893 , w_30894 , w_30895 , 
		w_30896 , w_30897 , w_30898 , w_30899 , w_30900 , w_30901 , w_30902 , w_30903 , w_30904 , w_30905 , 
		w_30906 , w_30907 , w_30908 , w_30909 , w_30910 , w_30911 , w_30912 , w_30913 , w_30914 , w_30915 , 
		w_30916 , w_30917 , w_30918 , w_30919 , w_30920 , w_30921 , w_30922 , w_30923 , w_30924 , w_30925 , 
		w_30926 , w_30927 , w_30928 , w_30929 , w_30930 , w_30931 , w_30932 , w_30933 , w_30934 , w_30935 , 
		w_30936 , w_30937 , w_30938 , w_30939 , w_30940 , w_30941 , w_30942 , w_30943 , w_30944 , w_30945 , 
		w_30946 , w_30947 , w_30948 , w_30949 , w_30950 , w_30951 , w_30952 , w_30953 , w_30954 , w_30955 , 
		w_30956 , w_30957 , w_30958 , w_30959 , w_30960 , w_30961 , w_30962 , w_30963 , w_30964 , w_30965 , 
		w_30966 , w_30967 , w_30968 , w_30969 , w_30970 , w_30971 , w_30972 , w_30973 , w_30974 , w_30975 , 
		w_30976 , w_30977 , w_30978 , w_30979 , w_30980 , w_30981 , w_30982 , w_30983 , w_30984 , w_30985 , 
		w_30986 , w_30987 , w_30988 , w_30989 , w_30990 , w_30991 , w_30992 , w_30993 , w_30994 , w_30995 , 
		w_30996 , w_30997 , w_30998 , w_30999 , w_31000 , w_31001 , w_31002 , w_31003 , w_31004 , w_31005 , 
		w_31006 , w_31007 , w_31008 , w_31009 , w_31010 , w_31011 , w_31012 , w_31013 , w_31014 , w_31015 , 
		w_31016 , w_31017 , w_31018 , w_31019 , w_31020 , w_31021 , w_31022 , w_31023 , w_31024 , w_31025 , 
		w_31026 , w_31027 , w_31028 , w_31029 , w_31030 , w_31031 , w_31032 , w_31033 , w_31034 , w_31035 , 
		w_31036 , w_31037 , w_31038 , w_31039 , w_31040 , w_31041 , w_31042 , w_31043 , w_31044 , w_31045 , 
		w_31046 , w_31047 , w_31048 , w_31049 , w_31050 , w_31051 , w_31052 , w_31053 , w_31054 , w_31055 , 
		w_31056 , w_31057 , w_31058 , w_31059 , w_31060 , w_31061 , w_31062 , w_31063 , w_31064 , w_31065 , 
		w_31066 , w_31067 , w_31068 , w_31069 , w_31070 , w_31071 , w_31072 , w_31073 , w_31074 , w_31075 , 
		w_31076 , w_31077 , w_31078 , w_31079 , w_31080 , w_31081 , w_31082 , w_31083 , w_31084 , w_31085 , 
		w_31086 , w_31087 , w_31088 , w_31089 , w_31090 , w_31091 , w_31092 , w_31093 , w_31094 , w_31095 , 
		w_31096 , w_31097 , w_31098 , w_31099 , w_31100 , w_31101 , w_31102 , w_31103 , w_31104 , w_31105 , 
		w_31106 , w_31107 , w_31108 , w_31109 , w_31110 , w_31111 , w_31112 , w_31113 , w_31114 , w_31115 , 
		w_31116 , w_31117 , w_31118 , w_31119 , w_31120 , w_31121 , w_31122 , w_31123 , w_31124 , w_31125 , 
		w_31126 , w_31127 , w_31128 , w_31129 , w_31130 , w_31131 , w_31132 , w_31133 , w_31134 , w_31135 , 
		w_31136 , w_31137 , w_31138 , w_31139 , w_31140 , w_31141 , w_31142 , w_31143 , w_31144 , w_31145 , 
		w_31146 , w_31147 , w_31148 , w_31149 , w_31150 , w_31151 , w_31152 , w_31153 , w_31154 , w_31155 , 
		w_31156 , w_31157 , w_31158 , w_31159 , w_31160 , w_31161 , w_31162 , w_31163 , w_31164 , w_31165 , 
		w_31166 , w_31167 , w_31168 , w_31169 , w_31170 , w_31171 , w_31172 , w_31173 , w_31174 , w_31175 , 
		w_31176 , w_31177 , w_31178 , w_31179 , w_31180 , w_31181 , w_31182 , w_31183 , w_31184 , w_31185 , 
		w_31186 , w_31187 , w_31188 , w_31189 , w_31190 , w_31191 , w_31192 , w_31193 , w_31194 , w_31195 , 
		w_31196 , w_31197 , w_31198 , w_31199 , w_31200 , w_31201 , w_31202 , w_31203 , w_31204 , w_31205 , 
		w_31206 , w_31207 , w_31208 , w_31209 , w_31210 , w_31211 , w_31212 , w_31213 , w_31214 , w_31215 , 
		w_31216 , w_31217 , w_31218 , w_31219 , w_31220 , w_31221 , w_31222 , w_31223 , w_31224 , w_31225 , 
		w_31226 , w_31227 , w_31228 , w_31229 , w_31230 , w_31231 , w_31232 , w_31233 , w_31234 , w_31235 , 
		w_31236 , w_31237 , w_31238 , w_31239 , w_31240 , w_31241 , w_31242 , w_31243 , w_31244 , w_31245 , 
		w_31246 , w_31247 , w_31248 , w_31249 , w_31250 , w_31251 , w_31252 , w_31253 , w_31254 , w_31255 , 
		w_31256 , w_31257 , w_31258 , w_31259 , w_31260 , w_31261 , w_31262 , w_31263 , w_31264 , w_31265 , 
		w_31266 , w_31267 , w_31268 , w_31269 , w_31270 , w_31271 , w_31272 , w_31273 , w_31274 , w_31275 , 
		w_31276 , w_31277 , w_31278 , w_31279 , w_31280 , w_31281 , w_31282 , w_31283 , w_31284 , w_31285 , 
		w_31286 , w_31287 , w_31288 , w_31289 , w_31290 , w_31291 , w_31292 , w_31293 , w_31294 , w_31295 , 
		w_31296 , w_31297 , w_31298 , w_31299 , w_31300 , w_31301 , w_31302 , w_31303 , w_31304 , w_31305 , 
		w_31306 , w_31307 , w_31308 , w_31309 , w_31310 , w_31311 , w_31312 , w_31313 , w_31314 , w_31315 , 
		w_31316 , w_31317 , w_31318 , w_31319 , w_31320 , w_31321 , w_31322 , w_31323 , w_31324 , w_31325 , 
		w_31326 , w_31327 , w_31328 , w_31329 , w_31330 , w_31331 , w_31332 , w_31333 , w_31334 , w_31335 , 
		w_31336 , w_31337 , w_31338 , w_31339 , w_31340 , w_31341 , w_31342 , w_31343 , w_31344 , w_31345 , 
		w_31346 , w_31347 , w_31348 , w_31349 , w_31350 , w_31351 , w_31352 , w_31353 , w_31354 , w_31355 , 
		w_31356 , w_31357 , w_31358 , w_31359 , w_31360 , w_31361 , w_31362 , w_31363 , w_31364 , w_31365 , 
		w_31366 , w_31367 , w_31368 , w_31369 , w_31370 , w_31371 , w_31372 , w_31373 , w_31374 , w_31375 , 
		w_31376 , w_31377 , w_31378 , w_31379 , w_31380 , w_31381 , w_31382 , w_31383 , w_31384 , w_31385 , 
		w_31386 , w_31387 , w_31388 , w_31389 , w_31390 , w_31391 , w_31392 , w_31393 , w_31394 , w_31395 , 
		w_31396 , w_31397 , w_31398 , w_31399 , w_31400 , w_31401 , w_31402 , w_31403 , w_31404 , w_31405 , 
		w_31406 , w_31407 , w_31408 , w_31409 , w_31410 , w_31411 , w_31412 , w_31413 , w_31414 , w_31415 , 
		w_31416 , w_31417 , w_31418 , w_31419 , w_31420 , w_31421 , w_31422 , w_31423 , w_31424 , w_31425 , 
		w_31426 , w_31427 , w_31428 , w_31429 , w_31430 , w_31431 , w_31432 , w_31433 , w_31434 , w_31435 , 
		w_31436 , w_31437 , w_31438 , w_31439 , w_31440 , w_31441 , w_31442 , w_31443 , w_31444 , w_31445 , 
		w_31446 , w_31447 , w_31448 , w_31449 , w_31450 , w_31451 , w_31452 , w_31453 , w_31454 , w_31455 , 
		w_31456 , w_31457 , w_31458 , w_31459 , w_31460 , w_31461 , w_31462 , w_31463 , w_31464 , w_31465 , 
		w_31466 , w_31467 , w_31468 , w_31469 , w_31470 , w_31471 , w_31472 , w_31473 , w_31474 , w_31475 , 
		w_31476 , w_31477 , w_31478 , w_31479 , w_31480 , w_31481 , w_31482 , w_31483 , w_31484 , w_31485 , 
		w_31486 , w_31487 , w_31488 , w_31489 , w_31490 , w_31491 , w_31492 , w_31493 , w_31494 , w_31495 , 
		w_31496 , w_31497 , w_31498 , w_31499 , w_31500 , w_31501 , w_31502 , w_31503 , w_31504 , w_31505 , 
		w_31506 , w_31507 , w_31508 , w_31509 , w_31510 , w_31511 , w_31512 , w_31513 , w_31514 , w_31515 , 
		w_31516 , w_31517 , w_31518 , w_31519 , w_31520 , w_31521 , w_31522 , w_31523 , w_31524 , w_31525 , 
		w_31526 , w_31527 , w_31528 , w_31529 , w_31530 , w_31531 , w_31532 , w_31533 , w_31534 , w_31535 , 
		w_31536 , w_31537 , w_31538 , w_31539 , w_31540 , w_31541 , w_31542 , w_31543 , w_31544 , w_31545 , 
		w_31546 , w_31547 , w_31548 , w_31549 , w_31550 , w_31551 , w_31552 , w_31553 , w_31554 , w_31555 , 
		w_31556 , w_31557 , w_31558 , w_31559 , w_31560 , w_31561 , w_31562 , w_31563 , w_31564 , w_31565 , 
		w_31566 , w_31567 , w_31568 , w_31569 , w_31570 , w_31571 , w_31572 , w_31573 , w_31574 , w_31575 , 
		w_31576 , w_31577 , w_31578 , w_31579 , w_31580 , w_31581 , w_31582 , w_31583 , w_31584 , w_31585 , 
		w_31586 , w_31587 , w_31588 , w_31589 , w_31590 , w_31591 , w_31592 , w_31593 , w_31594 , w_31595 , 
		w_31596 , w_31597 , w_31598 , w_31599 , w_31600 , w_31601 , w_31602 , w_31603 , w_31604 , w_31605 , 
		w_31606 , w_31607 , w_31608 , w_31609 , w_31610 , w_31611 , w_31612 , w_31613 , w_31614 , w_31615 , 
		w_31616 , w_31617 , w_31618 , w_31619 , w_31620 , w_31621 , w_31622 , w_31623 , w_31624 , w_31625 , 
		w_31626 , w_31627 , w_31628 , w_31629 , w_31630 , w_31631 , w_31632 , w_31633 , w_31634 , w_31635 , 
		w_31636 , w_31637 , w_31638 , w_31639 , w_31640 , w_31641 , w_31642 , w_31643 , w_31644 , w_31645 , 
		w_31646 , w_31647 , w_31648 , w_31649 , w_31650 , w_31651 , w_31652 , w_31653 , w_31654 , w_31655 , 
		w_31656 , w_31657 , w_31658 , w_31659 , w_31660 , w_31661 , w_31662 , w_31663 , w_31664 , w_31665 , 
		w_31666 , w_31667 , w_31668 , w_31669 , w_31670 , w_31671 , w_31672 , w_31673 , w_31674 , w_31675 , 
		w_31676 , w_31677 , w_31678 , w_31679 , w_31680 , w_31681 , w_31682 , w_31683 , w_31684 , w_31685 , 
		w_31686 , w_31687 , w_31688 , w_31689 , w_31690 , w_31691 , w_31692 , w_31693 , w_31694 , w_31695 , 
		w_31696 , w_31697 , w_31698 , w_31699 , w_31700 , w_31701 , w_31702 , w_31703 , w_31704 , w_31705 , 
		w_31706 , w_31707 , w_31708 , w_31709 , w_31710 , w_31711 , w_31712 , w_31713 , w_31714 , w_31715 , 
		w_31716 , w_31717 , w_31718 , w_31719 , w_31720 , w_31721 , w_31722 , w_31723 , w_31724 , w_31725 , 
		w_31726 , w_31727 , w_31728 , w_31729 , w_31730 , w_31731 , w_31732 , w_31733 , w_31734 , w_31735 , 
		w_31736 , w_31737 , w_31738 , w_31739 , w_31740 , w_31741 , w_31742 , w_31743 , w_31744 , w_31745 , 
		w_31746 , w_31747 , w_31748 , w_31749 , w_31750 , w_31751 , w_31752 , w_31753 , w_31754 , w_31755 , 
		w_31756 , w_31757 , w_31758 , w_31759 , w_31760 , w_31761 , w_31762 , w_31763 , w_31764 , w_31765 , 
		w_31766 , w_31767 , w_31768 , w_31769 , w_31770 , w_31771 , w_31772 , w_31773 , w_31774 , w_31775 , 
		w_31776 , w_31777 , w_31778 , w_31779 , w_31780 , w_31781 , w_31782 , w_31783 , w_31784 , w_31785 , 
		w_31786 , w_31787 , w_31788 , w_31789 , w_31790 , w_31791 , w_31792 , w_31793 , w_31794 , w_31795 , 
		w_31796 , w_31797 , w_31798 , w_31799 , w_31800 , w_31801 , w_31802 , w_31803 , w_31804 , w_31805 , 
		w_31806 , w_31807 , w_31808 , w_31809 , w_31810 , w_31811 , w_31812 , w_31813 , w_31814 , w_31815 , 
		w_31816 , w_31817 , w_31818 , w_31819 , w_31820 , w_31821 , w_31822 , w_31823 , w_31824 , w_31825 , 
		w_31826 , w_31827 , w_31828 , w_31829 , w_31830 , w_31831 , w_31832 , w_31833 , w_31834 , w_31835 , 
		w_31836 , w_31837 , w_31838 , w_31839 , w_31840 , w_31841 , w_31842 , w_31843 , w_31844 , w_31845 , 
		w_31846 , w_31847 , w_31848 , w_31849 , w_31850 , w_31851 , w_31852 , w_31853 , w_31854 , w_31855 , 
		w_31856 , w_31857 , w_31858 , w_31859 , w_31860 , w_31861 , w_31862 , w_31863 , w_31864 , w_31865 , 
		w_31866 , w_31867 , w_31868 , w_31869 , w_31870 , w_31871 , w_31872 , w_31873 , w_31874 , w_31875 , 
		w_31876 , w_31877 , w_31878 , w_31879 , w_31880 , w_31881 , w_31882 , w_31883 , w_31884 , w_31885 , 
		w_31886 , w_31887 , w_31888 , w_31889 , w_31890 , w_31891 , w_31892 , w_31893 , w_31894 , w_31895 , 
		w_31896 , w_31897 , w_31898 , w_31899 , w_31900 , w_31901 , w_31902 , w_31903 , w_31904 , w_31905 , 
		w_31906 , w_31907 , w_31908 , w_31909 , w_31910 , w_31911 , w_31912 , w_31913 , w_31914 , w_31915 , 
		w_31916 , w_31917 , w_31918 , w_31919 , w_31920 , w_31921 , w_31922 , w_31923 , w_31924 , w_31925 , 
		w_31926 , w_31927 , w_31928 , w_31929 , w_31930 , w_31931 , w_31932 , w_31933 , w_31934 , w_31935 , 
		w_31936 , w_31937 , w_31938 , w_31939 , w_31940 , w_31941 , w_31942 , w_31943 , w_31944 , w_31945 , 
		w_31946 , w_31947 , w_31948 , w_31949 , w_31950 , w_31951 , w_31952 , w_31953 , w_31954 , w_31955 , 
		w_31956 , w_31957 , w_31958 , w_31959 , w_31960 , w_31961 , w_31962 , w_31963 , w_31964 , w_31965 , 
		w_31966 , w_31967 , w_31968 , w_31969 , w_31970 , w_31971 , w_31972 , w_31973 , w_31974 , w_31975 , 
		w_31976 , w_31977 , w_31978 , w_31979 , w_31980 , w_31981 , w_31982 , w_31983 , w_31984 , w_31985 , 
		w_31986 , w_31987 , w_31988 , w_31989 , w_31990 , w_31991 , w_31992 , w_31993 , w_31994 , w_31995 , 
		w_31996 , w_31997 , w_31998 , w_31999 , w_32000 , w_32001 , w_32002 , w_32003 , w_32004 , w_32005 , 
		w_32006 , w_32007 , w_32008 , w_32009 , w_32010 , w_32011 , w_32012 , w_32013 , w_32014 , w_32015 , 
		w_32016 , w_32017 , w_32018 , w_32019 , w_32020 , w_32021 , w_32022 , w_32023 , w_32024 , w_32025 , 
		w_32026 , w_32027 , w_32028 , w_32029 , w_32030 , w_32031 , w_32032 , w_32033 , w_32034 , w_32035 , 
		w_32036 , w_32037 , w_32038 , w_32039 , w_32040 , w_32041 , w_32042 , w_32043 , w_32044 , w_32045 , 
		w_32046 , w_32047 , w_32048 , w_32049 , w_32050 , w_32051 , w_32052 , w_32053 , w_32054 , w_32055 , 
		w_32056 , w_32057 , w_32058 , w_32059 , w_32060 , w_32061 , w_32062 , w_32063 , w_32064 , w_32065 , 
		w_32066 , w_32067 , w_32068 , w_32069 , w_32070 , w_32071 , w_32072 , w_32073 , w_32074 , w_32075 , 
		w_32076 , w_32077 , w_32078 , w_32079 , w_32080 , w_32081 , w_32082 , w_32083 , w_32084 , w_32085 , 
		w_32086 , w_32087 , w_32088 , w_32089 , w_32090 , w_32091 , w_32092 , w_32093 , w_32094 , w_32095 , 
		w_32096 , w_32097 , w_32098 , w_32099 , w_32100 , w_32101 , w_32102 , w_32103 , w_32104 , w_32105 , 
		w_32106 , w_32107 , w_32108 , w_32109 , w_32110 , w_32111 , w_32112 , w_32113 , w_32114 , w_32115 , 
		w_32116 , w_32117 , w_32118 , w_32119 , w_32120 , w_32121 , w_32122 , w_32123 , w_32124 , w_32125 , 
		w_32126 , w_32127 , w_32128 , w_32129 , w_32130 , w_32131 , w_32132 , w_32133 , w_32134 , w_32135 , 
		w_32136 , w_32137 , w_32138 , w_32139 , w_32140 , w_32141 , w_32142 , w_32143 , w_32144 , w_32145 , 
		w_32146 , w_32147 , w_32148 , w_32149 , w_32150 , w_32151 , w_32152 , w_32153 , w_32154 , w_32155 , 
		w_32156 , w_32157 , w_32158 , w_32159 , w_32160 , w_32161 , w_32162 , w_32163 , w_32164 , w_32165 , 
		w_32166 , w_32167 , w_32168 , w_32169 , w_32170 , w_32171 , w_32172 , w_32173 , w_32174 , w_32175 , 
		w_32176 , w_32177 , w_32178 , w_32179 , w_32180 , w_32181 , w_32182 , w_32183 , w_32184 , w_32185 , 
		w_32186 , w_32187 , w_32188 , w_32189 , w_32190 , w_32191 , w_32192 , w_32193 , w_32194 , w_32195 , 
		w_32196 , w_32197 , w_32198 , w_32199 , w_32200 , w_32201 , w_32202 , w_32203 , w_32204 , w_32205 , 
		w_32206 , w_32207 , w_32208 , w_32209 , w_32210 , w_32211 , w_32212 , w_32213 , w_32214 , w_32215 , 
		w_32216 , w_32217 , w_32218 , w_32219 , w_32220 , w_32221 , w_32222 , w_32223 , w_32224 , w_32225 , 
		w_32226 , w_32227 , w_32228 , w_32229 , w_32230 , w_32231 , w_32232 , w_32233 , w_32234 , w_32235 , 
		w_32236 , w_32237 , w_32238 , w_32239 , w_32240 , w_32241 , w_32242 , w_32243 , w_32244 , w_32245 , 
		w_32246 , w_32247 , w_32248 , w_32249 , w_32250 , w_32251 , w_32252 , w_32253 , w_32254 , w_32255 , 
		w_32256 , w_32257 , w_32258 , w_32259 , w_32260 , w_32261 , w_32262 , w_32263 , w_32264 , w_32265 , 
		w_32266 , w_32267 , w_32268 , w_32269 , w_32270 , w_32271 , w_32272 , w_32273 , w_32274 , w_32275 , 
		w_32276 , w_32277 , w_32278 , w_32279 , w_32280 , w_32281 , w_32282 , w_32283 , w_32284 , w_32285 , 
		w_32286 , w_32287 , w_32288 , w_32289 , w_32290 , w_32291 , w_32292 , w_32293 , w_32294 , w_32295 , 
		w_32296 , w_32297 , w_32298 , w_32299 , w_32300 , w_32301 , w_32302 , w_32303 , w_32304 , w_32305 , 
		w_32306 , w_32307 , w_32308 , w_32309 , w_32310 , w_32311 , w_32312 , w_32313 , w_32314 , w_32315 , 
		w_32316 , w_32317 , w_32318 , w_32319 , w_32320 , w_32321 , w_32322 , w_32323 , w_32324 , w_32325 , 
		w_32326 , w_32327 , w_32328 , w_32329 , w_32330 , w_32331 , w_32332 , w_32333 , w_32334 , w_32335 , 
		w_32336 , w_32337 , w_32338 , w_32339 , w_32340 , w_32341 , w_32342 , w_32343 , w_32344 , w_32345 , 
		w_32346 , w_32347 , w_32348 , w_32349 , w_32350 , w_32351 , w_32352 , w_32353 , w_32354 , w_32355 , 
		w_32356 , w_32357 , w_32358 , w_32359 , w_32360 , w_32361 , w_32362 , w_32363 , w_32364 , w_32365 , 
		w_32366 , w_32367 , w_32368 , w_32369 , w_32370 , w_32371 , w_32372 , w_32373 , w_32374 , w_32375 , 
		w_32376 , w_32377 , w_32378 , w_32379 , w_32380 , w_32381 , w_32382 , w_32383 , w_32384 , w_32385 , 
		w_32386 , w_32387 , w_32388 , w_32389 , w_32390 , w_32391 , w_32392 , w_32393 , w_32394 , w_32395 , 
		w_32396 , w_32397 , w_32398 , w_32399 , w_32400 , w_32401 , w_32402 , w_32403 , w_32404 , w_32405 , 
		w_32406 , w_32407 , w_32408 , w_32409 , w_32410 , w_32411 , w_32412 , w_32413 , w_32414 , w_32415 , 
		w_32416 , w_32417 , w_32418 , w_32419 , w_32420 , w_32421 , w_32422 , w_32423 , w_32424 , w_32425 , 
		w_32426 , w_32427 , w_32428 , w_32429 , w_32430 , w_32431 , w_32432 , w_32433 , w_32434 , w_32435 , 
		w_32436 , w_32437 , w_32438 , w_32439 , w_32440 , w_32441 , w_32442 , w_32443 , w_32444 , w_32445 , 
		w_32446 , w_32447 , w_32448 , w_32449 , w_32450 , w_32451 , w_32452 , w_32453 , w_32454 , w_32455 , 
		w_32456 , w_32457 , w_32458 , w_32459 , w_32460 , w_32461 , w_32462 , w_32463 , w_32464 , w_32465 , 
		w_32466 , w_32467 , w_32468 , w_32469 , w_32470 , w_32471 , w_32472 , w_32473 , w_32474 , w_32475 , 
		w_32476 , w_32477 , w_32478 , w_32479 , w_32480 , w_32481 , w_32482 , w_32483 , w_32484 , w_32485 , 
		w_32486 , w_32487 , w_32488 , w_32489 , w_32490 , w_32491 , w_32492 , w_32493 , w_32494 , w_32495 , 
		w_32496 , w_32497 , w_32498 , w_32499 , w_32500 , w_32501 , w_32502 , w_32503 , w_32504 , w_32505 , 
		w_32506 , w_32507 , w_32508 , w_32509 , w_32510 , w_32511 , w_32512 , w_32513 , w_32514 , w_32515 , 
		w_32516 , w_32517 , w_32518 , w_32519 , w_32520 , w_32521 , w_32522 , w_32523 , w_32524 , w_32525 , 
		w_32526 , w_32527 , w_32528 , w_32529 , w_32530 , w_32531 , w_32532 , w_32533 , w_32534 , w_32535 , 
		w_32536 , w_32537 , w_32538 , w_32539 , w_32540 , w_32541 , w_32542 , w_32543 , w_32544 , w_32545 , 
		w_32546 , w_32547 , w_32548 , w_32549 , w_32550 , w_32551 , w_32552 , w_32553 , w_32554 , w_32555 , 
		w_32556 , w_32557 , w_32558 , w_32559 , w_32560 , w_32561 , w_32562 , w_32563 , w_32564 , w_32565 , 
		w_32566 , w_32567 , w_32568 , w_32569 , w_32570 , w_32571 , w_32572 , w_32573 , w_32574 , w_32575 , 
		w_32576 , w_32577 , w_32578 , w_32579 , w_32580 , w_32581 , w_32582 , w_32583 , w_32584 , w_32585 , 
		w_32586 , w_32587 , w_32588 , w_32589 , w_32590 , w_32591 , w_32592 , w_32593 , w_32594 , w_32595 , 
		w_32596 , w_32597 , w_32598 , w_32599 , w_32600 , w_32601 , w_32602 , w_32603 , w_32604 , w_32605 , 
		w_32606 , w_32607 , w_32608 , w_32609 , w_32610 , w_32611 , w_32612 , w_32613 , w_32614 , w_32615 , 
		w_32616 , w_32617 , w_32618 , w_32619 , w_32620 , w_32621 , w_32622 , w_32623 , w_32624 , w_32625 , 
		w_32626 , w_32627 , w_32628 , w_32629 , w_32630 , w_32631 , w_32632 , w_32633 , w_32634 , w_32635 , 
		w_32636 , w_32637 , w_32638 , w_32639 , w_32640 , w_32641 , w_32642 , w_32643 , w_32644 , w_32645 , 
		w_32646 , w_32647 , w_32648 , w_32649 , w_32650 , w_32651 , w_32652 , w_32653 , w_32654 , w_32655 , 
		w_32656 , w_32657 , w_32658 , w_32659 , w_32660 , w_32661 , w_32662 , w_32663 , w_32664 , w_32665 , 
		w_32666 , w_32667 , w_32668 , w_32669 , w_32670 , w_32671 , w_32672 , w_32673 , w_32674 , w_32675 , 
		w_32676 , w_32677 , w_32678 , w_32679 , w_32680 , w_32681 , w_32682 , w_32683 , w_32684 , w_32685 , 
		w_32686 , w_32687 , w_32688 , w_32689 , w_32690 , w_32691 , w_32692 , w_32693 , w_32694 , w_32695 , 
		w_32696 , w_32697 , w_32698 , w_32699 , w_32700 , w_32701 , w_32702 , w_32703 , w_32704 , w_32705 , 
		w_32706 , w_32707 , w_32708 , w_32709 , w_32710 , w_32711 , w_32712 , w_32713 , w_32714 , w_32715 , 
		w_32716 , w_32717 , w_32718 , w_32719 , w_32720 , w_32721 , w_32722 , w_32723 , w_32724 , w_32725 , 
		w_32726 , w_32727 , w_32728 , w_32729 , w_32730 , w_32731 , w_32732 , w_32733 , w_32734 , w_32735 , 
		w_32736 , w_32737 , w_32738 , w_32739 , w_32740 , w_32741 , w_32742 , w_32743 , w_32744 , w_32745 , 
		w_32746 , w_32747 , w_32748 , w_32749 , w_32750 , w_32751 , w_32752 , w_32753 , w_32754 , w_32755 , 
		w_32756 , w_32757 , w_32758 , w_32759 , w_32760 , w_32761 , w_32762 , w_32763 , w_32764 , w_32765 , 
		w_32766 , w_32767 , w_32768 , w_32769 , w_32770 , w_32771 , w_32772 , w_32773 , w_32774 , w_32775 , 
		w_32776 , w_32777 , w_32778 , w_32779 , w_32780 , w_32781 , w_32782 , w_32783 , w_32784 , w_32785 , 
		w_32786 , w_32787 , w_32788 , w_32789 , w_32790 , w_32791 , w_32792 , w_32793 , w_32794 , w_32795 , 
		w_32796 , w_32797 , w_32798 , w_32799 , w_32800 , w_32801 , w_32802 , w_32803 , w_32804 , w_32805 , 
		w_32806 , w_32807 , w_32808 , w_32809 , w_32810 , w_32811 , w_32812 , w_32813 , w_32814 , w_32815 , 
		w_32816 , w_32817 , w_32818 , w_32819 , w_32820 , w_32821 , w_32822 , w_32823 , w_32824 , w_32825 , 
		w_32826 , w_32827 , w_32828 , w_32829 , w_32830 , w_32831 , w_32832 , w_32833 , w_32834 , w_32835 , 
		w_32836 , w_32837 , w_32838 , w_32839 , w_32840 , w_32841 , w_32842 , w_32843 , w_32844 , w_32845 , 
		w_32846 , w_32847 , w_32848 , w_32849 , w_32850 , w_32851 , w_32852 , w_32853 , w_32854 , w_32855 , 
		w_32856 , w_32857 , w_32858 , w_32859 , w_32860 , w_32861 , w_32862 , w_32863 , w_32864 , w_32865 , 
		w_32866 , w_32867 , w_32868 , w_32869 , w_32870 , w_32871 , w_32872 , w_32873 , w_32874 , w_32875 , 
		w_32876 , w_32877 , w_32878 , w_32879 , w_32880 , w_32881 , w_32882 , w_32883 , w_32884 , w_32885 , 
		w_32886 , w_32887 , w_32888 , w_32889 , w_32890 , w_32891 , w_32892 , w_32893 , w_32894 , w_32895 , 
		w_32896 , w_32897 , w_32898 , w_32899 , w_32900 , w_32901 , w_32902 , w_32903 , w_32904 , w_32905 , 
		w_32906 , w_32907 , w_32908 , w_32909 , w_32910 , w_32911 , w_32912 , w_32913 , w_32914 , w_32915 , 
		w_32916 , w_32917 , w_32918 , w_32919 , w_32920 , w_32921 , w_32922 , w_32923 , w_32924 , w_32925 , 
		w_32926 , w_32927 , w_32928 , w_32929 , w_32930 , w_32931 , w_32932 , w_32933 , w_32934 , w_32935 , 
		w_32936 , w_32937 , w_32938 , w_32939 , w_32940 , w_32941 , w_32942 , w_32943 , w_32944 , w_32945 , 
		w_32946 , w_32947 , w_32948 , w_32949 , w_32950 , w_32951 , w_32952 , w_32953 , w_32954 , w_32955 , 
		w_32956 , w_32957 , w_32958 , w_32959 , w_32960 , w_32961 , w_32962 , w_32963 , w_32964 , w_32965 , 
		w_32966 , w_32967 , w_32968 , w_32969 , w_32970 , w_32971 , w_32972 , w_32973 , w_32974 , w_32975 , 
		w_32976 , w_32977 , w_32978 , w_32979 , w_32980 , w_32981 , w_32982 , w_32983 , w_32984 , w_32985 , 
		w_32986 , w_32987 , w_32988 , w_32989 , w_32990 , w_32991 , w_32992 , w_32993 , w_32994 , w_32995 , 
		w_32996 , w_32997 , w_32998 , w_32999 , w_33000 , w_33001 , w_33002 , w_33003 , w_33004 , w_33005 , 
		w_33006 , w_33007 , w_33008 , w_33009 , w_33010 , w_33011 , w_33012 , w_33013 , w_33014 , w_33015 , 
		w_33016 , w_33017 , w_33018 , w_33019 , w_33020 , w_33021 , w_33022 , w_33023 , w_33024 , w_33025 , 
		w_33026 , w_33027 , w_33028 , w_33029 , w_33030 , w_33031 , w_33032 , w_33033 , w_33034 , w_33035 , 
		w_33036 , w_33037 , w_33038 , w_33039 , w_33040 , w_33041 , w_33042 , w_33043 , w_33044 , w_33045 , 
		w_33046 , w_33047 , w_33048 , w_33049 , w_33050 , w_33051 , w_33052 , w_33053 , w_33054 , w_33055 , 
		w_33056 , w_33057 , w_33058 , w_33059 , w_33060 , w_33061 , w_33062 , w_33063 , w_33064 , w_33065 , 
		w_33066 , w_33067 , w_33068 , w_33069 , w_33070 , w_33071 , w_33072 , w_33073 , w_33074 , w_33075 , 
		w_33076 , w_33077 , w_33078 , w_33079 , w_33080 , w_33081 , w_33082 , w_33083 , w_33084 , w_33085 , 
		w_33086 , w_33087 , w_33088 , w_33089 , w_33090 , w_33091 , w_33092 , w_33093 , w_33094 , w_33095 , 
		w_33096 , w_33097 , w_33098 , w_33099 , w_33100 , w_33101 , w_33102 , w_33103 , w_33104 , w_33105 , 
		w_33106 , w_33107 , w_33108 , w_33109 , w_33110 , w_33111 , w_33112 , w_33113 , w_33114 , w_33115 , 
		w_33116 , w_33117 , w_33118 , w_33119 , w_33120 , w_33121 , w_33122 , w_33123 , w_33124 , w_33125 , 
		w_33126 , w_33127 , w_33128 , w_33129 , w_33130 , w_33131 , w_33132 , w_33133 , w_33134 , w_33135 , 
		w_33136 , w_33137 , w_33138 , w_33139 , w_33140 , w_33141 , w_33142 , w_33143 , w_33144 , w_33145 , 
		w_33146 , w_33147 , w_33148 , w_33149 , w_33150 , w_33151 , w_33152 , w_33153 , w_33154 , w_33155 , 
		w_33156 , w_33157 , w_33158 , w_33159 , w_33160 , w_33161 , w_33162 , w_33163 , w_33164 , w_33165 , 
		w_33166 , w_33167 , w_33168 , w_33169 , w_33170 , w_33171 , w_33172 , w_33173 , w_33174 , w_33175 , 
		w_33176 , w_33177 , w_33178 , w_33179 , w_33180 , w_33181 , w_33182 , w_33183 , w_33184 , w_33185 , 
		w_33186 , w_33187 , w_33188 , w_33189 , w_33190 , w_33191 , w_33192 , w_33193 , w_33194 , w_33195 , 
		w_33196 , w_33197 , w_33198 , w_33199 , w_33200 , w_33201 , w_33202 , w_33203 , w_33204 , w_33205 , 
		w_33206 , w_33207 , w_33208 , w_33209 , w_33210 , w_33211 , w_33212 , w_33213 , w_33214 , w_33215 , 
		w_33216 , w_33217 , w_33218 , w_33219 , w_33220 , w_33221 , w_33222 , w_33223 , w_33224 , w_33225 , 
		w_33226 , w_33227 , w_33228 , w_33229 , w_33230 , w_33231 , w_33232 , w_33233 , w_33234 , w_33235 , 
		w_33236 , w_33237 , w_33238 , w_33239 , w_33240 , w_33241 , w_33242 , w_33243 , w_33244 , w_33245 , 
		w_33246 , w_33247 , w_33248 , w_33249 , w_33250 , w_33251 , w_33252 , w_33253 , w_33254 , w_33255 , 
		w_33256 , w_33257 , w_33258 , w_33259 , w_33260 , w_33261 , w_33262 , w_33263 , w_33264 , w_33265 , 
		w_33266 , w_33267 , w_33268 , w_33269 , w_33270 , w_33271 , w_33272 , w_33273 , w_33274 , w_33275 , 
		w_33276 , w_33277 , w_33278 , w_33279 , w_33280 , w_33281 , w_33282 , w_33283 , w_33284 , w_33285 , 
		w_33286 , w_33287 , w_33288 , w_33289 , w_33290 , w_33291 , w_33292 , w_33293 , w_33294 , w_33295 , 
		w_33296 , w_33297 , w_33298 , w_33299 , w_33300 , w_33301 , w_33302 , w_33303 , w_33304 , w_33305 , 
		w_33306 , w_33307 , w_33308 , w_33309 , w_33310 , w_33311 , w_33312 , w_33313 , w_33314 , w_33315 , 
		w_33316 , w_33317 , w_33318 , w_33319 , w_33320 , w_33321 , w_33322 , w_33323 , w_33324 , w_33325 , 
		w_33326 , w_33327 , w_33328 , w_33329 , w_33330 , w_33331 , w_33332 , w_33333 , w_33334 , w_33335 , 
		w_33336 , w_33337 , w_33338 , w_33339 , w_33340 , w_33341 , w_33342 , w_33343 , w_33344 , w_33345 , 
		w_33346 , w_33347 , w_33348 , w_33349 , w_33350 , w_33351 , w_33352 , w_33353 , w_33354 , w_33355 , 
		w_33356 , w_33357 , w_33358 , w_33359 , w_33360 , w_33361 , w_33362 , w_33363 , w_33364 , w_33365 , 
		w_33366 , w_33367 , w_33368 , w_33369 , w_33370 , w_33371 , w_33372 , w_33373 , w_33374 , w_33375 , 
		w_33376 , w_33377 , w_33378 , w_33379 , w_33380 , w_33381 , w_33382 , w_33383 , w_33384 , w_33385 , 
		w_33386 , w_33387 , w_33388 , w_33389 , w_33390 , w_33391 , w_33392 , w_33393 , w_33394 , w_33395 , 
		w_33396 , w_33397 , w_33398 , w_33399 , w_33400 , w_33401 , w_33402 , w_33403 , w_33404 , w_33405 , 
		w_33406 , w_33407 , w_33408 , w_33409 , w_33410 , w_33411 , w_33412 , w_33413 , w_33414 , w_33415 , 
		w_33416 , w_33417 , w_33418 , w_33419 , w_33420 , w_33421 , w_33422 , w_33423 , w_33424 , w_33425 , 
		w_33426 , w_33427 , w_33428 , w_33429 , w_33430 , w_33431 , w_33432 , w_33433 , w_33434 , w_33435 , 
		w_33436 , w_33437 , w_33438 , w_33439 , w_33440 , w_33441 , w_33442 , w_33443 , w_33444 , w_33445 , 
		w_33446 , w_33447 , w_33448 , w_33449 , w_33450 , w_33451 , w_33452 , w_33453 , w_33454 , w_33455 , 
		w_33456 , w_33457 , w_33458 , w_33459 , w_33460 , w_33461 , w_33462 , w_33463 , w_33464 , w_33465 , 
		w_33466 , w_33467 , w_33468 , w_33469 , w_33470 , w_33471 , w_33472 , w_33473 , w_33474 , w_33475 , 
		w_33476 , w_33477 , w_33478 , w_33479 , w_33480 , w_33481 , w_33482 , w_33483 , w_33484 , w_33485 , 
		w_33486 , w_33487 , w_33488 , w_33489 , w_33490 , w_33491 , w_33492 , w_33493 , w_33494 , w_33495 , 
		w_33496 , w_33497 , w_33498 , w_33499 , w_33500 , w_33501 , w_33502 , w_33503 , w_33504 , w_33505 , 
		w_33506 , w_33507 , w_33508 , w_33509 , w_33510 , w_33511 , w_33512 , w_33513 , w_33514 , w_33515 , 
		w_33516 , w_33517 , w_33518 , w_33519 , w_33520 , w_33521 , w_33522 , w_33523 , w_33524 , w_33525 , 
		w_33526 , w_33527 , w_33528 , w_33529 , w_33530 , w_33531 , w_33532 , w_33533 , w_33534 , w_33535 , 
		w_33536 , w_33537 , w_33538 , w_33539 , w_33540 , w_33541 , w_33542 , w_33543 , w_33544 , w_33545 , 
		w_33546 , w_33547 , w_33548 , w_33549 , w_33550 , w_33551 , w_33552 , w_33553 , w_33554 , w_33555 , 
		w_33556 , w_33557 , w_33558 , w_33559 , w_33560 , w_33561 , w_33562 , w_33563 , w_33564 , w_33565 , 
		w_33566 , w_33567 , w_33568 , w_33569 , w_33570 , w_33571 , w_33572 , w_33573 , w_33574 , w_33575 , 
		w_33576 , w_33577 , w_33578 , w_33579 , w_33580 , w_33581 , w_33582 , w_33583 , w_33584 , w_33585 , 
		w_33586 , w_33587 , w_33588 , w_33589 , w_33590 , w_33591 , w_33592 , w_33593 , w_33594 , w_33595 , 
		w_33596 , w_33597 , w_33598 , w_33599 , w_33600 , w_33601 , w_33602 , w_33603 , w_33604 , w_33605 , 
		w_33606 , w_33607 , w_33608 , w_33609 , w_33610 , w_33611 , w_33612 , w_33613 , w_33614 , w_33615 , 
		w_33616 , w_33617 , w_33618 , w_33619 , w_33620 , w_33621 , w_33622 , w_33623 , w_33624 , w_33625 , 
		w_33626 , w_33627 , w_33628 , w_33629 , w_33630 , w_33631 , w_33632 , w_33633 , w_33634 , w_33635 , 
		w_33636 , w_33637 , w_33638 , w_33639 , w_33640 , w_33641 , w_33642 , w_33643 , w_33644 , w_33645 , 
		w_33646 , w_33647 , w_33648 , w_33649 , w_33650 , w_33651 , w_33652 , w_33653 , w_33654 , w_33655 , 
		w_33656 , w_33657 , w_33658 , w_33659 , w_33660 , w_33661 , w_33662 , w_33663 , w_33664 , w_33665 , 
		w_33666 , w_33667 , w_33668 , w_33669 , w_33670 , w_33671 , w_33672 , w_33673 , w_33674 , w_33675 , 
		w_33676 , w_33677 , w_33678 , w_33679 , w_33680 , w_33681 , w_33682 , w_33683 , w_33684 , w_33685 , 
		w_33686 , w_33687 , w_33688 , w_33689 , w_33690 , w_33691 , w_33692 , w_33693 , w_33694 , w_33695 , 
		w_33696 , w_33697 , w_33698 , w_33699 , w_33700 , w_33701 , w_33702 , w_33703 , w_33704 , w_33705 , 
		w_33706 , w_33707 , w_33708 , w_33709 , w_33710 , w_33711 , w_33712 , w_33713 , w_33714 , w_33715 , 
		w_33716 , w_33717 , w_33718 , w_33719 , w_33720 , w_33721 , w_33722 , w_33723 , w_33724 , w_33725 , 
		w_33726 , w_33727 , w_33728 , w_33729 , w_33730 , w_33731 , w_33732 , w_33733 , w_33734 , w_33735 , 
		w_33736 , w_33737 , w_33738 , w_33739 , w_33740 , w_33741 , w_33742 , w_33743 , w_33744 , w_33745 , 
		w_33746 , w_33747 , w_33748 , w_33749 , w_33750 , w_33751 , w_33752 , w_33753 , w_33754 , w_33755 , 
		w_33756 , w_33757 , w_33758 , w_33759 , w_33760 , w_33761 , w_33762 , w_33763 , w_33764 , w_33765 , 
		w_33766 , w_33767 , w_33768 , w_33769 , w_33770 , w_33771 , w_33772 , w_33773 , w_33774 , w_33775 , 
		w_33776 , w_33777 , w_33778 , w_33779 , w_33780 , w_33781 , w_33782 , w_33783 , w_33784 , w_33785 , 
		w_33786 , w_33787 , w_33788 , w_33789 , w_33790 , w_33791 , w_33792 , w_33793 , w_33794 , w_33795 , 
		w_33796 , w_33797 , w_33798 , w_33799 , w_33800 , w_33801 , w_33802 , w_33803 , w_33804 , w_33805 , 
		w_33806 , w_33807 , w_33808 , w_33809 , w_33810 , w_33811 , w_33812 , w_33813 , w_33814 , w_33815 , 
		w_33816 , w_33817 , w_33818 , w_33819 , w_33820 , w_33821 , w_33822 , w_33823 , w_33824 , w_33825 , 
		w_33826 , w_33827 , w_33828 , w_33829 , w_33830 , w_33831 , w_33832 , w_33833 , w_33834 , w_33835 , 
		w_33836 , w_33837 , w_33838 , w_33839 , w_33840 , w_33841 , w_33842 , w_33843 , w_33844 , w_33845 , 
		w_33846 , w_33847 , w_33848 , w_33849 , w_33850 , w_33851 , w_33852 , w_33853 , w_33854 , w_33855 , 
		w_33856 , w_33857 , w_33858 , w_33859 , w_33860 , w_33861 , w_33862 , w_33863 , w_33864 , w_33865 , 
		w_33866 , w_33867 , w_33868 , w_33869 , w_33870 , w_33871 , w_33872 , w_33873 , w_33874 , w_33875 , 
		w_33876 , w_33877 , w_33878 , w_33879 , w_33880 , w_33881 , w_33882 , w_33883 , w_33884 , w_33885 , 
		w_33886 , w_33887 , w_33888 , w_33889 , w_33890 , w_33891 , w_33892 , w_33893 , w_33894 , w_33895 , 
		w_33896 , w_33897 , w_33898 , w_33899 , w_33900 , w_33901 , w_33902 , w_33903 , w_33904 , w_33905 , 
		w_33906 , w_33907 , w_33908 , w_33909 , w_33910 , w_33911 , w_33912 , w_33913 , w_33914 , w_33915 , 
		w_33916 , w_33917 , w_33918 , w_33919 , w_33920 , w_33921 , w_33922 , w_33923 , w_33924 , w_33925 , 
		w_33926 , w_33927 , w_33928 , w_33929 , w_33930 , w_33931 , w_33932 , w_33933 , w_33934 , w_33935 , 
		w_33936 , w_33937 , w_33938 , w_33939 , w_33940 , w_33941 , w_33942 , w_33943 , w_33944 , w_33945 , 
		w_33946 , w_33947 , w_33948 , w_33949 , w_33950 , w_33951 , w_33952 , w_33953 , w_33954 , w_33955 , 
		w_33956 , w_33957 , w_33958 , w_33959 , w_33960 , w_33961 , w_33962 , w_33963 , w_33964 , w_33965 , 
		w_33966 , w_33967 , w_33968 , w_33969 , w_33970 , w_33971 , w_33972 , w_33973 , w_33974 , w_33975 , 
		w_33976 , w_33977 , w_33978 , w_33979 , w_33980 , w_33981 , w_33982 , w_33983 , w_33984 , w_33985 , 
		w_33986 , w_33987 , w_33988 , w_33989 , w_33990 , w_33991 , w_33992 , w_33993 , w_33994 , w_33995 , 
		w_33996 , w_33997 , w_33998 , w_33999 , w_34000 , w_34001 , w_34002 , w_34003 , w_34004 , w_34005 , 
		w_34006 , w_34007 , w_34008 , w_34009 , w_34010 , w_34011 , w_34012 , w_34013 , w_34014 , w_34015 , 
		w_34016 , w_34017 , w_34018 , w_34019 , w_34020 , w_34021 , w_34022 , w_34023 , w_34024 , w_34025 , 
		w_34026 , w_34027 , w_34028 , w_34029 , w_34030 , w_34031 , w_34032 , w_34033 , w_34034 , w_34035 , 
		w_34036 , w_34037 , w_34038 , w_34039 , w_34040 , w_34041 , w_34042 , w_34043 , w_34044 , w_34045 , 
		w_34046 , w_34047 , w_34048 , w_34049 , w_34050 , w_34051 , w_34052 , w_34053 , w_34054 , w_34055 , 
		w_34056 , w_34057 , w_34058 , w_34059 , w_34060 , w_34061 , w_34062 , w_34063 , w_34064 , w_34065 , 
		w_34066 , w_34067 , w_34068 , w_34069 , w_34070 , w_34071 , w_34072 , w_34073 , w_34074 , w_34075 , 
		w_34076 , w_34077 , w_34078 , w_34079 , w_34080 , w_34081 , w_34082 , w_34083 , w_34084 , w_34085 , 
		w_34086 , w_34087 , w_34088 , w_34089 , w_34090 , w_34091 , w_34092 , w_34093 , w_34094 , w_34095 , 
		w_34096 , w_34097 , w_34098 , w_34099 , w_34100 , w_34101 , w_34102 , w_34103 , w_34104 , w_34105 , 
		w_34106 , w_34107 , w_34108 , w_34109 , w_34110 , w_34111 , w_34112 , w_34113 , w_34114 , w_34115 , 
		w_34116 , w_34117 , w_34118 , w_34119 , w_34120 , w_34121 , w_34122 , w_34123 , w_34124 , w_34125 , 
		w_34126 , w_34127 , w_34128 , w_34129 , w_34130 , w_34131 , w_34132 , w_34133 , w_34134 , w_34135 , 
		w_34136 , w_34137 , w_34138 , w_34139 , w_34140 , w_34141 , w_34142 , w_34143 , w_34144 , w_34145 , 
		w_34146 , w_34147 , w_34148 , w_34149 , w_34150 , w_34151 , w_34152 , w_34153 , w_34154 , w_34155 , 
		w_34156 , w_34157 , w_34158 , w_34159 , w_34160 , w_34161 , w_34162 , w_34163 , w_34164 , w_34165 , 
		w_34166 , w_34167 , w_34168 , w_34169 , w_34170 , w_34171 , w_34172 , w_34173 , w_34174 , w_34175 , 
		w_34176 , w_34177 , w_34178 , w_34179 , w_34180 , w_34181 , w_34182 , w_34183 , w_34184 , w_34185 , 
		w_34186 , w_34187 , w_34188 , w_34189 , w_34190 , w_34191 , w_34192 , w_34193 , w_34194 , w_34195 , 
		w_34196 , w_34197 , w_34198 , w_34199 , w_34200 , w_34201 , w_34202 , w_34203 , w_34204 , w_34205 , 
		w_34206 , w_34207 , w_34208 , w_34209 , w_34210 , w_34211 , w_34212 , w_34213 , w_34214 , w_34215 , 
		w_34216 , w_34217 , w_34218 , w_34219 , w_34220 , w_34221 , w_34222 , w_34223 , w_34224 , w_34225 , 
		w_34226 , w_34227 , w_34228 , w_34229 , w_34230 , w_34231 , w_34232 , w_34233 , w_34234 , w_34235 , 
		w_34236 , w_34237 , w_34238 , w_34239 , w_34240 , w_34241 , w_34242 , w_34243 , w_34244 , w_34245 , 
		w_34246 , w_34247 , w_34248 , w_34249 , w_34250 , w_34251 , w_34252 , w_34253 , w_34254 , w_34255 , 
		w_34256 , w_34257 , w_34258 , w_34259 , w_34260 , w_34261 , w_34262 , w_34263 , w_34264 , w_34265 , 
		w_34266 , w_34267 , w_34268 , w_34269 , w_34270 , w_34271 , w_34272 , w_34273 , w_34274 , w_34275 , 
		w_34276 , w_34277 , w_34278 , w_34279 , w_34280 , w_34281 , w_34282 , w_34283 , w_34284 , w_34285 , 
		w_34286 , w_34287 , w_34288 , w_34289 , w_34290 , w_34291 , w_34292 , w_34293 , w_34294 , w_34295 , 
		w_34296 , w_34297 , w_34298 , w_34299 , w_34300 , w_34301 , w_34302 , w_34303 , w_34304 , w_34305 , 
		w_34306 , w_34307 , w_34308 , w_34309 , w_34310 , w_34311 , w_34312 , w_34313 , w_34314 , w_34315 , 
		w_34316 , w_34317 , w_34318 , w_34319 , w_34320 , w_34321 , w_34322 , w_34323 , w_34324 , w_34325 , 
		w_34326 , w_34327 , w_34328 , w_34329 , w_34330 , w_34331 , w_34332 , w_34333 , w_34334 , w_34335 , 
		w_34336 , w_34337 , w_34338 , w_34339 , w_34340 , w_34341 , w_34342 , w_34343 , w_34344 , w_34345 , 
		w_34346 , w_34347 , w_34348 , w_34349 , w_34350 , w_34351 , w_34352 , w_34353 , w_34354 , w_34355 , 
		w_34356 , w_34357 , w_34358 , w_34359 , w_34360 , w_34361 , w_34362 , w_34363 , w_34364 , w_34365 , 
		w_34366 , w_34367 , w_34368 , w_34369 , w_34370 , w_34371 , w_34372 , w_34373 , w_34374 , w_34375 , 
		w_34376 , w_34377 , w_34378 , w_34379 , w_34380 , w_34381 , w_34382 , w_34383 , w_34384 , w_34385 , 
		w_34386 , w_34387 , w_34388 , w_34389 , w_34390 , w_34391 , w_34392 , w_34393 , w_34394 , w_34395 , 
		w_34396 , w_34397 , w_34398 , w_34399 , w_34400 , w_34401 , w_34402 , w_34403 , w_34404 , w_34405 , 
		w_34406 , w_34407 , w_34408 , w_34409 , w_34410 , w_34411 , w_34412 , w_34413 , w_34414 , w_34415 , 
		w_34416 , w_34417 , w_34418 , w_34419 , w_34420 , w_34421 , w_34422 , w_34423 , w_34424 , w_34425 , 
		w_34426 , w_34427 , w_34428 , w_34429 , w_34430 , w_34431 , w_34432 , w_34433 , w_34434 , w_34435 , 
		w_34436 , w_34437 , w_34438 , w_34439 , w_34440 , w_34441 , w_34442 , w_34443 , w_34444 , w_34445 , 
		w_34446 , w_34447 , w_34448 , w_34449 , w_34450 , w_34451 , w_34452 , w_34453 , w_34454 , w_34455 , 
		w_34456 , w_34457 , w_34458 , w_34459 , w_34460 , w_34461 , w_34462 , w_34463 , w_34464 , w_34465 , 
		w_34466 , w_34467 , w_34468 , w_34469 , w_34470 , w_34471 , w_34472 , w_34473 , w_34474 , w_34475 , 
		w_34476 , w_34477 , w_34478 , w_34479 , w_34480 , w_34481 , w_34482 , w_34483 , w_34484 , w_34485 , 
		w_34486 , w_34487 , w_34488 , w_34489 , w_34490 , w_34491 , w_34492 , w_34493 , w_34494 , w_34495 , 
		w_34496 , w_34497 , w_34498 , w_34499 , w_34500 , w_34501 , w_34502 , w_34503 , w_34504 , w_34505 , 
		w_34506 , w_34507 , w_34508 , w_34509 , w_34510 , w_34511 , w_34512 , w_34513 , w_34514 , w_34515 , 
		w_34516 , w_34517 , w_34518 , w_34519 , w_34520 , w_34521 , w_34522 , w_34523 , w_34524 , w_34525 , 
		w_34526 , w_34527 , w_34528 , w_34529 , w_34530 , w_34531 , w_34532 , w_34533 , w_34534 , w_34535 , 
		w_34536 , w_34537 , w_34538 , w_34539 , w_34540 , w_34541 , w_34542 , w_34543 , w_34544 , w_34545 , 
		w_34546 , w_34547 , w_34548 , w_34549 , w_34550 , w_34551 , w_34552 , w_34553 , w_34554 , w_34555 , 
		w_34556 , w_34557 , w_34558 , w_34559 , w_34560 , w_34561 , w_34562 , w_34563 , w_34564 , w_34565 , 
		w_34566 , w_34567 , w_34568 , w_34569 , w_34570 , w_34571 , w_34572 , w_34573 , w_34574 , w_34575 , 
		w_34576 , w_34577 , w_34578 , w_34579 , w_34580 , w_34581 , w_34582 , w_34583 , w_34584 , w_34585 , 
		w_34586 , w_34587 , w_34588 , w_34589 , w_34590 , w_34591 , w_34592 , w_34593 , w_34594 , w_34595 , 
		w_34596 , w_34597 , w_34598 , w_34599 , w_34600 , w_34601 , w_34602 , w_34603 , w_34604 , w_34605 , 
		w_34606 , w_34607 , w_34608 , w_34609 , w_34610 , w_34611 , w_34612 , w_34613 , w_34614 , w_34615 , 
		w_34616 , w_34617 , w_34618 , w_34619 , w_34620 , w_34621 , w_34622 , w_34623 , w_34624 , w_34625 , 
		w_34626 , w_34627 , w_34628 , w_34629 , w_34630 , w_34631 , w_34632 , w_34633 , w_34634 , w_34635 , 
		w_34636 , w_34637 , w_34638 , w_34639 , w_34640 , w_34641 , w_34642 , w_34643 , w_34644 , w_34645 , 
		w_34646 , w_34647 , w_34648 , w_34649 , w_34650 , w_34651 , w_34652 , w_34653 , w_34654 , w_34655 , 
		w_34656 , w_34657 , w_34658 , w_34659 , w_34660 , w_34661 , w_34662 , w_34663 , w_34664 , w_34665 , 
		w_34666 , w_34667 , w_34668 , w_34669 , w_34670 , w_34671 , w_34672 , w_34673 , w_34674 , w_34675 , 
		w_34676 , w_34677 , w_34678 , w_34679 , w_34680 , w_34681 , w_34682 , w_34683 , w_34684 , w_34685 , 
		w_34686 , w_34687 , w_34688 , w_34689 , w_34690 , w_34691 , w_34692 , w_34693 , w_34694 , w_34695 , 
		w_34696 , w_34697 , w_34698 , w_34699 , w_34700 , w_34701 , w_34702 , w_34703 , w_34704 , w_34705 , 
		w_34706 , w_34707 , w_34708 , w_34709 , w_34710 , w_34711 , w_34712 , w_34713 , w_34714 , w_34715 , 
		w_34716 , w_34717 , w_34718 , w_34719 , w_34720 , w_34721 , w_34722 , w_34723 , w_34724 , w_34725 , 
		w_34726 , w_34727 , w_34728 , w_34729 , w_34730 , w_34731 , w_34732 , w_34733 , w_34734 , w_34735 , 
		w_34736 , w_34737 , w_34738 , w_34739 , w_34740 , w_34741 , w_34742 , w_34743 , w_34744 , w_34745 , 
		w_34746 , w_34747 , w_34748 , w_34749 , w_34750 , w_34751 , w_34752 , w_34753 , w_34754 , w_34755 , 
		w_34756 , w_34757 , w_34758 , w_34759 , w_34760 , w_34761 , w_34762 , w_34763 , w_34764 , w_34765 , 
		w_34766 , w_34767 , w_34768 , w_34769 , w_34770 , w_34771 , w_34772 , w_34773 , w_34774 , w_34775 , 
		w_34776 , w_34777 , w_34778 , w_34779 , w_34780 , w_34781 , w_34782 , w_34783 , w_34784 , w_34785 , 
		w_34786 , w_34787 , w_34788 , w_34789 , w_34790 , w_34791 , w_34792 , w_34793 , w_34794 , w_34795 , 
		w_34796 , w_34797 , w_34798 , w_34799 , w_34800 , w_34801 , w_34802 , w_34803 , w_34804 , w_34805 , 
		w_34806 , w_34807 , w_34808 , w_34809 , w_34810 , w_34811 , w_34812 , w_34813 , w_34814 , w_34815 , 
		w_34816 , w_34817 , w_34818 , w_34819 , w_34820 , w_34821 , w_34822 , w_34823 , w_34824 , w_34825 , 
		w_34826 , w_34827 , w_34828 , w_34829 , w_34830 , w_34831 , w_34832 , w_34833 , w_34834 , w_34835 , 
		w_34836 , w_34837 , w_34838 , w_34839 , w_34840 , w_34841 , w_34842 , w_34843 , w_34844 , w_34845 , 
		w_34846 , w_34847 , w_34848 , w_34849 , w_34850 , w_34851 , w_34852 , w_34853 , w_34854 , w_34855 , 
		w_34856 , w_34857 , w_34858 , w_34859 , w_34860 , w_34861 , w_34862 , w_34863 , w_34864 , w_34865 , 
		w_34866 , w_34867 , w_34868 , w_34869 , w_34870 , w_34871 , w_34872 , w_34873 , w_34874 , w_34875 , 
		w_34876 , w_34877 , w_34878 , w_34879 , w_34880 , w_34881 , w_34882 , w_34883 , w_34884 , w_34885 , 
		w_34886 , w_34887 , w_34888 , w_34889 , w_34890 , w_34891 , w_34892 , w_34893 , w_34894 , w_34895 , 
		w_34896 , w_34897 , w_34898 , w_34899 , w_34900 , w_34901 , w_34902 , w_34903 , w_34904 , w_34905 , 
		w_34906 , w_34907 , w_34908 , w_34909 , w_34910 , w_34911 , w_34912 , w_34913 , w_34914 , w_34915 , 
		w_34916 , w_34917 , w_34918 , w_34919 , w_34920 , w_34921 , w_34922 , w_34923 , w_34924 , w_34925 , 
		w_34926 , w_34927 , w_34928 , w_34929 , w_34930 , w_34931 , w_34932 , w_34933 , w_34934 , w_34935 , 
		w_34936 , w_34937 , w_34938 , w_34939 , w_34940 , w_34941 , w_34942 , w_34943 , w_34944 , w_34945 , 
		w_34946 , w_34947 , w_34948 , w_34949 , w_34950 , w_34951 , w_34952 , w_34953 , w_34954 , w_34955 , 
		w_34956 , w_34957 , w_34958 , w_34959 , w_34960 , w_34961 , w_34962 , w_34963 , w_34964 , w_34965 , 
		w_34966 , w_34967 , w_34968 , w_34969 , w_34970 , w_34971 , w_34972 , w_34973 , w_34974 , w_34975 , 
		w_34976 , w_34977 , w_34978 , w_34979 , w_34980 , w_34981 , w_34982 , w_34983 , w_34984 , w_34985 , 
		w_34986 , w_34987 , w_34988 , w_34989 , w_34990 , w_34991 , w_34992 , w_34993 , w_34994 , w_34995 , 
		w_34996 , w_34997 , w_34998 , w_34999 , w_35000 , w_35001 , w_35002 , w_35003 , w_35004 , w_35005 , 
		w_35006 , w_35007 , w_35008 , w_35009 , w_35010 , w_35011 , w_35012 , w_35013 , w_35014 , w_35015 , 
		w_35016 , w_35017 , w_35018 , w_35019 , w_35020 , w_35021 , w_35022 , w_35023 , w_35024 , w_35025 , 
		w_35026 , w_35027 , w_35028 , w_35029 , w_35030 , w_35031 , w_35032 , w_35033 , w_35034 , w_35035 , 
		w_35036 , w_35037 , w_35038 , w_35039 , w_35040 , w_35041 , w_35042 , w_35043 , w_35044 , w_35045 , 
		w_35046 , w_35047 , w_35048 , w_35049 , w_35050 , w_35051 , w_35052 , w_35053 , w_35054 , w_35055 , 
		w_35056 , w_35057 , w_35058 , w_35059 , w_35060 , w_35061 , w_35062 , w_35063 , w_35064 , w_35065 , 
		w_35066 , w_35067 , w_35068 , w_35069 , w_35070 , w_35071 , w_35072 , w_35073 , w_35074 , w_35075 , 
		w_35076 , w_35077 , w_35078 , w_35079 , w_35080 , w_35081 , w_35082 , w_35083 , w_35084 , w_35085 , 
		w_35086 , w_35087 , w_35088 , w_35089 , w_35090 , w_35091 , w_35092 , w_35093 , w_35094 , w_35095 , 
		w_35096 , w_35097 , w_35098 , w_35099 , w_35100 , w_35101 , w_35102 , w_35103 , w_35104 , w_35105 , 
		w_35106 , w_35107 , w_35108 , w_35109 , w_35110 , w_35111 , w_35112 , w_35113 , w_35114 , w_35115 , 
		w_35116 , w_35117 , w_35118 , w_35119 , w_35120 , w_35121 , w_35122 , w_35123 , w_35124 , w_35125 , 
		w_35126 , w_35127 , w_35128 , w_35129 , w_35130 , w_35131 , w_35132 , w_35133 , w_35134 , w_35135 , 
		w_35136 , w_35137 , w_35138 , w_35139 , w_35140 , w_35141 , w_35142 , w_35143 , w_35144 , w_35145 , 
		w_35146 , w_35147 , w_35148 , w_35149 , w_35150 , w_35151 , w_35152 , w_35153 , w_35154 , w_35155 , 
		w_35156 , w_35157 , w_35158 , w_35159 , w_35160 , w_35161 , w_35162 , w_35163 , w_35164 , w_35165 , 
		w_35166 , w_35167 , w_35168 , w_35169 , w_35170 , w_35171 , w_35172 , w_35173 , w_35174 , w_35175 , 
		w_35176 , w_35177 , w_35178 , w_35179 , w_35180 , w_35181 , w_35182 , w_35183 , w_35184 , w_35185 , 
		w_35186 , w_35187 , w_35188 , w_35189 , w_35190 , w_35191 , w_35192 , w_35193 , w_35194 , w_35195 , 
		w_35196 , w_35197 , w_35198 , w_35199 , w_35200 , w_35201 , w_35202 , w_35203 , w_35204 , w_35205 , 
		w_35206 , w_35207 , w_35208 , w_35209 , w_35210 , w_35211 , w_35212 , w_35213 , w_35214 , w_35215 , 
		w_35216 , w_35217 , w_35218 , w_35219 , w_35220 , w_35221 , w_35222 , w_35223 , w_35224 , w_35225 , 
		w_35226 , w_35227 , w_35228 , w_35229 , w_35230 , w_35231 , w_35232 , w_35233 , w_35234 , w_35235 , 
		w_35236 , w_35237 , w_35238 , w_35239 , w_35240 , w_35241 , w_35242 , w_35243 , w_35244 , w_35245 , 
		w_35246 , w_35247 , w_35248 , w_35249 , w_35250 , w_35251 , w_35252 , w_35253 , w_35254 , w_35255 , 
		w_35256 , w_35257 , w_35258 , w_35259 , w_35260 , w_35261 , w_35262 , w_35263 , w_35264 , w_35265 , 
		w_35266 , w_35267 , w_35268 , w_35269 , w_35270 , w_35271 , w_35272 , w_35273 , w_35274 , w_35275 , 
		w_35276 , w_35277 , w_35278 , w_35279 , w_35280 , w_35281 , w_35282 , w_35283 , w_35284 , w_35285 , 
		w_35286 , w_35287 , w_35288 , w_35289 , w_35290 , w_35291 , w_35292 , w_35293 , w_35294 , w_35295 , 
		w_35296 , w_35297 , w_35298 , w_35299 , w_35300 , w_35301 , w_35302 , w_35303 , w_35304 , w_35305 , 
		w_35306 , w_35307 , w_35308 , w_35309 , w_35310 , w_35311 , w_35312 , w_35313 , w_35314 , w_35315 , 
		w_35316 , w_35317 , w_35318 , w_35319 , w_35320 , w_35321 , w_35322 , w_35323 , w_35324 , w_35325 , 
		w_35326 , w_35327 , w_35328 , w_35329 , w_35330 , w_35331 , w_35332 , w_35333 , w_35334 , w_35335 , 
		w_35336 , w_35337 , w_35338 , w_35339 , w_35340 , w_35341 , w_35342 , w_35343 , w_35344 , w_35345 , 
		w_35346 , w_35347 , w_35348 , w_35349 , w_35350 , w_35351 , w_35352 , w_35353 , w_35354 , w_35355 , 
		w_35356 , w_35357 , w_35358 , w_35359 , w_35360 , w_35361 , w_35362 , w_35363 , w_35364 , w_35365 , 
		w_35366 , w_35367 , w_35368 , w_35369 , w_35370 , w_35371 , w_35372 , w_35373 , w_35374 , w_35375 , 
		w_35376 , w_35377 , w_35378 , w_35379 , w_35380 , w_35381 , w_35382 , w_35383 , w_35384 , w_35385 , 
		w_35386 , w_35387 , w_35388 , w_35389 , w_35390 , w_35391 , w_35392 , w_35393 , w_35394 , w_35395 , 
		w_35396 , w_35397 , w_35398 , w_35399 , w_35400 , w_35401 , w_35402 , w_35403 , w_35404 , w_35405 , 
		w_35406 , w_35407 , w_35408 , w_35409 , w_35410 , w_35411 , w_35412 , w_35413 , w_35414 , w_35415 , 
		w_35416 , w_35417 , w_35418 , w_35419 , w_35420 , w_35421 , w_35422 , w_35423 , w_35424 , w_35425 , 
		w_35426 , w_35427 , w_35428 , w_35429 , w_35430 , w_35431 , w_35432 , w_35433 , w_35434 , w_35435 , 
		w_35436 , w_35437 , w_35438 , w_35439 , w_35440 , w_35441 , w_35442 , w_35443 , w_35444 , w_35445 , 
		w_35446 , w_35447 , w_35448 , w_35449 , w_35450 , w_35451 , w_35452 , w_35453 , w_35454 , w_35455 , 
		w_35456 , w_35457 , w_35458 , w_35459 , w_35460 , w_35461 , w_35462 , w_35463 , w_35464 , w_35465 , 
		w_35466 , w_35467 , w_35468 , w_35469 , w_35470 , w_35471 , w_35472 , w_35473 , w_35474 , w_35475 , 
		w_35476 , w_35477 , w_35478 , w_35479 , w_35480 , w_35481 , w_35482 , w_35483 , w_35484 , w_35485 , 
		w_35486 , w_35487 , w_35488 , w_35489 , w_35490 , w_35491 , w_35492 , w_35493 , w_35494 , w_35495 , 
		w_35496 , w_35497 , w_35498 , w_35499 , w_35500 , w_35501 , w_35502 , w_35503 , w_35504 , w_35505 , 
		w_35506 , w_35507 , w_35508 , w_35509 , w_35510 , w_35511 , w_35512 , w_35513 , w_35514 , w_35515 , 
		w_35516 , w_35517 , w_35518 , w_35519 , w_35520 , w_35521 , w_35522 , w_35523 , w_35524 , w_35525 , 
		w_35526 , w_35527 , w_35528 , w_35529 , w_35530 , w_35531 , w_35532 , w_35533 , w_35534 , w_35535 , 
		w_35536 , w_35537 , w_35538 , w_35539 , w_35540 , w_35541 , w_35542 , w_35543 , w_35544 , w_35545 , 
		w_35546 , w_35547 , w_35548 , w_35549 , w_35550 , w_35551 , w_35552 , w_35553 , w_35554 , w_35555 , 
		w_35556 , w_35557 , w_35558 , w_35559 , w_35560 , w_35561 , w_35562 , w_35563 , w_35564 , w_35565 , 
		w_35566 , w_35567 , w_35568 , w_35569 , w_35570 , w_35571 , w_35572 , w_35573 , w_35574 , w_35575 , 
		w_35576 , w_35577 , w_35578 , w_35579 , w_35580 , w_35581 , w_35582 , w_35583 , w_35584 , w_35585 , 
		w_35586 , w_35587 , w_35588 , w_35589 , w_35590 , w_35591 , w_35592 , w_35593 , w_35594 , w_35595 , 
		w_35596 , w_35597 , w_35598 , w_35599 , w_35600 , w_35601 , w_35602 , w_35603 , w_35604 , w_35605 , 
		w_35606 , w_35607 , w_35608 , w_35609 , w_35610 , w_35611 , w_35612 , w_35613 , w_35614 , w_35615 , 
		w_35616 , w_35617 , w_35618 , w_35619 , w_35620 , w_35621 , w_35622 , w_35623 , w_35624 , w_35625 , 
		w_35626 , w_35627 , w_35628 , w_35629 , w_35630 , w_35631 , w_35632 , w_35633 , w_35634 , w_35635 , 
		w_35636 , w_35637 , w_35638 , w_35639 , w_35640 , w_35641 , w_35642 , w_35643 , w_35644 , w_35645 , 
		w_35646 , w_35647 , w_35648 , w_35649 , w_35650 , w_35651 , w_35652 , w_35653 , w_35654 , w_35655 , 
		w_35656 , w_35657 , w_35658 , w_35659 , w_35660 , w_35661 , w_35662 , w_35663 , w_35664 , w_35665 , 
		w_35666 , w_35667 , w_35668 , w_35669 , w_35670 , w_35671 , w_35672 , w_35673 , w_35674 , w_35675 , 
		w_35676 , w_35677 , w_35678 , w_35679 , w_35680 , w_35681 , w_35682 , w_35683 , w_35684 , w_35685 , 
		w_35686 , w_35687 , w_35688 , w_35689 , w_35690 , w_35691 , w_35692 , w_35693 , w_35694 , w_35695 , 
		w_35696 , w_35697 , w_35698 , w_35699 , w_35700 , w_35701 , w_35702 , w_35703 , w_35704 , w_35705 , 
		w_35706 , w_35707 , w_35708 , w_35709 , w_35710 , w_35711 , w_35712 , w_35713 , w_35714 , w_35715 , 
		w_35716 , w_35717 , w_35718 , w_35719 , w_35720 , w_35721 , w_35722 , w_35723 , w_35724 , w_35725 , 
		w_35726 , w_35727 , w_35728 , w_35729 , w_35730 , w_35731 , w_35732 , w_35733 , w_35734 , w_35735 , 
		w_35736 , w_35737 , w_35738 , w_35739 , w_35740 , w_35741 , w_35742 , w_35743 , w_35744 , w_35745 , 
		w_35746 , w_35747 , w_35748 , w_35749 , w_35750 , w_35751 , w_35752 , w_35753 , w_35754 , w_35755 , 
		w_35756 , w_35757 , w_35758 , w_35759 , w_35760 , w_35761 , w_35762 , w_35763 , w_35764 , w_35765 , 
		w_35766 , w_35767 , w_35768 , w_35769 , w_35770 , w_35771 , w_35772 , w_35773 , w_35774 , w_35775 , 
		w_35776 , w_35777 , w_35778 , w_35779 , w_35780 , w_35781 , w_35782 , w_35783 , w_35784 , w_35785 , 
		w_35786 , w_35787 , w_35788 , w_35789 , w_35790 , w_35791 , w_35792 , w_35793 , w_35794 , w_35795 , 
		w_35796 , w_35797 , w_35798 , w_35799 , w_35800 , w_35801 , w_35802 , w_35803 , w_35804 , w_35805 , 
		w_35806 , w_35807 , w_35808 , w_35809 , w_35810 , w_35811 , w_35812 , w_35813 , w_35814 , w_35815 , 
		w_35816 , w_35817 , w_35818 , w_35819 , w_35820 , w_35821 , w_35822 , w_35823 , w_35824 , w_35825 , 
		w_35826 , w_35827 , w_35828 , w_35829 , w_35830 , w_35831 , w_35832 , w_35833 , w_35834 , w_35835 , 
		w_35836 , w_35837 , w_35838 , w_35839 , w_35840 , w_35841 , w_35842 , w_35843 , w_35844 , w_35845 , 
		w_35846 , w_35847 , w_35848 , w_35849 , w_35850 , w_35851 , w_35852 , w_35853 , w_35854 , w_35855 , 
		w_35856 , w_35857 , w_35858 , w_35859 , w_35860 , w_35861 , w_35862 , w_35863 , w_35864 , w_35865 , 
		w_35866 , w_35867 , w_35868 , w_35869 , w_35870 , w_35871 , w_35872 , w_35873 , w_35874 , w_35875 , 
		w_35876 , w_35877 , w_35878 , w_35879 , w_35880 , w_35881 , w_35882 , w_35883 , w_35884 , w_35885 , 
		w_35886 , w_35887 , w_35888 , w_35889 , w_35890 , w_35891 , w_35892 , w_35893 , w_35894 , w_35895 , 
		w_35896 , w_35897 , w_35898 , w_35899 , w_35900 , w_35901 , w_35902 , w_35903 , w_35904 , w_35905 , 
		w_35906 , w_35907 , w_35908 , w_35909 , w_35910 , w_35911 , w_35912 , w_35913 , w_35914 , w_35915 , 
		w_35916 , w_35917 , w_35918 , w_35919 , w_35920 , w_35921 , w_35922 , w_35923 , w_35924 , w_35925 , 
		w_35926 , w_35927 , w_35928 , w_35929 , w_35930 , w_35931 , w_35932 , w_35933 , w_35934 , w_35935 , 
		w_35936 , w_35937 , w_35938 , w_35939 , w_35940 , w_35941 , w_35942 , w_35943 , w_35944 , w_35945 , 
		w_35946 , w_35947 , w_35948 , w_35949 , w_35950 , w_35951 , w_35952 , w_35953 , w_35954 , w_35955 , 
		w_35956 , w_35957 , w_35958 , w_35959 , w_35960 , w_35961 , w_35962 , w_35963 , w_35964 , w_35965 , 
		w_35966 , w_35967 , w_35968 , w_35969 , w_35970 , w_35971 , w_35972 , w_35973 , w_35974 , w_35975 , 
		w_35976 , w_35977 , w_35978 , w_35979 , w_35980 , w_35981 , w_35982 , w_35983 , w_35984 , w_35985 , 
		w_35986 , w_35987 , w_35988 , w_35989 , w_35990 , w_35991 , w_35992 , w_35993 , w_35994 , w_35995 , 
		w_35996 , w_35997 , w_35998 , w_35999 , w_36000 , w_36001 , w_36002 , w_36003 , w_36004 , w_36005 , 
		w_36006 , w_36007 , w_36008 , w_36009 , w_36010 , w_36011 , w_36012 , w_36013 , w_36014 , w_36015 , 
		w_36016 , w_36017 , w_36018 , w_36019 , w_36020 , w_36021 , w_36022 , w_36023 , w_36024 , w_36025 , 
		w_36026 , w_36027 , w_36028 , w_36029 , w_36030 , w_36031 , w_36032 , w_36033 , w_36034 , w_36035 , 
		w_36036 , w_36037 , w_36038 , w_36039 , w_36040 , w_36041 , w_36042 , w_36043 , w_36044 , w_36045 , 
		w_36046 , w_36047 , w_36048 , w_36049 , w_36050 , w_36051 , w_36052 , w_36053 , w_36054 , w_36055 , 
		w_36056 , w_36057 , w_36058 , w_36059 , w_36060 , w_36061 , w_36062 , w_36063 , w_36064 , w_36065 , 
		w_36066 , w_36067 , w_36068 , w_36069 , w_36070 , w_36071 , w_36072 , w_36073 , w_36074 , w_36075 , 
		w_36076 , w_36077 , w_36078 , w_36079 , w_36080 , w_36081 , w_36082 , w_36083 , w_36084 , w_36085 , 
		w_36086 , w_36087 , w_36088 , w_36089 , w_36090 , w_36091 , w_36092 , w_36093 , w_36094 , w_36095 , 
		w_36096 , w_36097 , w_36098 , w_36099 , w_36100 , w_36101 , w_36102 , w_36103 , w_36104 , w_36105 , 
		w_36106 , w_36107 , w_36108 , w_36109 , w_36110 , w_36111 , w_36112 , w_36113 , w_36114 , w_36115 , 
		w_36116 , w_36117 , w_36118 , w_36119 , w_36120 , w_36121 , w_36122 , w_36123 , w_36124 , w_36125 , 
		w_36126 , w_36127 , w_36128 , w_36129 , w_36130 , w_36131 , w_36132 , w_36133 , w_36134 , w_36135 , 
		w_36136 , w_36137 , w_36138 , w_36139 , w_36140 , w_36141 , w_36142 , w_36143 , w_36144 , w_36145 , 
		w_36146 , w_36147 , w_36148 , w_36149 , w_36150 , w_36151 , w_36152 , w_36153 , w_36154 , w_36155 , 
		w_36156 , w_36157 , w_36158 , w_36159 , w_36160 , w_36161 , w_36162 , w_36163 , w_36164 , w_36165 , 
		w_36166 , w_36167 , w_36168 , w_36169 , w_36170 , w_36171 , w_36172 , w_36173 , w_36174 , w_36175 , 
		w_36176 , w_36177 , w_36178 , w_36179 , w_36180 , w_36181 , w_36182 , w_36183 , w_36184 , w_36185 , 
		w_36186 , w_36187 , w_36188 , w_36189 , w_36190 , w_36191 , w_36192 , w_36193 , w_36194 , w_36195 , 
		w_36196 , w_36197 , w_36198 , w_36199 , w_36200 , w_36201 , w_36202 , w_36203 , w_36204 , w_36205 , 
		w_36206 , w_36207 , w_36208 , w_36209 , w_36210 , w_36211 , w_36212 , w_36213 , w_36214 , w_36215 , 
		w_36216 , w_36217 , w_36218 , w_36219 , w_36220 , w_36221 , w_36222 , w_36223 , w_36224 , w_36225 , 
		w_36226 , w_36227 , w_36228 , w_36229 , w_36230 , w_36231 , w_36232 , w_36233 , w_36234 , w_36235 , 
		w_36236 , w_36237 , w_36238 , w_36239 , w_36240 , w_36241 , w_36242 , w_36243 , w_36244 , w_36245 , 
		w_36246 , w_36247 , w_36248 , w_36249 , w_36250 , w_36251 , w_36252 , w_36253 , w_36254 , w_36255 , 
		w_36256 , w_36257 , w_36258 , w_36259 , w_36260 , w_36261 , w_36262 , w_36263 , w_36264 , w_36265 , 
		w_36266 , w_36267 , w_36268 , w_36269 , w_36270 , w_36271 , w_36272 , w_36273 , w_36274 , w_36275 , 
		w_36276 , w_36277 , w_36278 , w_36279 , w_36280 , w_36281 , w_36282 , w_36283 , w_36284 , w_36285 , 
		w_36286 , w_36287 , w_36288 , w_36289 , w_36290 , w_36291 , w_36292 , w_36293 , w_36294 , w_36295 , 
		w_36296 , w_36297 , w_36298 , w_36299 , w_36300 , w_36301 , w_36302 , w_36303 , w_36304 , w_36305 , 
		w_36306 , w_36307 , w_36308 , w_36309 , w_36310 , w_36311 , w_36312 , w_36313 , w_36314 , w_36315 , 
		w_36316 , w_36317 , w_36318 , w_36319 , w_36320 , w_36321 , w_36322 , w_36323 , w_36324 , w_36325 , 
		w_36326 , w_36327 , w_36328 , w_36329 , w_36330 , w_36331 , w_36332 , w_36333 , w_36334 , w_36335 , 
		w_36336 , w_36337 , w_36338 , w_36339 , w_36340 , w_36341 , w_36342 , w_36343 , w_36344 , w_36345 , 
		w_36346 , w_36347 , w_36348 , w_36349 , w_36350 , w_36351 , w_36352 , w_36353 , w_36354 , w_36355 , 
		w_36356 , w_36357 , w_36358 , w_36359 , w_36360 , w_36361 , w_36362 , w_36363 , w_36364 , w_36365 , 
		w_36366 , w_36367 , w_36368 , w_36369 , w_36370 , w_36371 , w_36372 , w_36373 , w_36374 , w_36375 , 
		w_36376 , w_36377 , w_36378 , w_36379 , w_36380 , w_36381 , w_36382 , w_36383 , w_36384 , w_36385 , 
		w_36386 , w_36387 , w_36388 , w_36389 , w_36390 , w_36391 , w_36392 , w_36393 , w_36394 , w_36395 , 
		w_36396 , w_36397 , w_36398 , w_36399 , w_36400 , w_36401 , w_36402 , w_36403 , w_36404 , w_36405 , 
		w_36406 , w_36407 , w_36408 , w_36409 , w_36410 , w_36411 , w_36412 , w_36413 , w_36414 , w_36415 , 
		w_36416 , w_36417 , w_36418 , w_36419 , w_36420 , w_36421 , w_36422 , w_36423 , w_36424 , w_36425 , 
		w_36426 , w_36427 , w_36428 , w_36429 , w_36430 , w_36431 , w_36432 , w_36433 , w_36434 , w_36435 , 
		w_36436 , w_36437 , w_36438 , w_36439 , w_36440 , w_36441 , w_36442 , w_36443 , w_36444 , w_36445 , 
		w_36446 , w_36447 , w_36448 , w_36449 , w_36450 , w_36451 , w_36452 , w_36453 , w_36454 , w_36455 , 
		w_36456 , w_36457 , w_36458 , w_36459 , w_36460 , w_36461 , w_36462 , w_36463 , w_36464 , w_36465 , 
		w_36466 , w_36467 , w_36468 , w_36469 , w_36470 , w_36471 , w_36472 , w_36473 , w_36474 , w_36475 , 
		w_36476 , w_36477 , w_36478 , w_36479 , w_36480 , w_36481 , w_36482 , w_36483 , w_36484 , w_36485 , 
		w_36486 , w_36487 , w_36488 , w_36489 , w_36490 , w_36491 , w_36492 , w_36493 , w_36494 , w_36495 , 
		w_36496 , w_36497 , w_36498 , w_36499 , w_36500 , w_36501 , w_36502 , w_36503 , w_36504 , w_36505 , 
		w_36506 , w_36507 , w_36508 , w_36509 , w_36510 , w_36511 , w_36512 , w_36513 , w_36514 , w_36515 , 
		w_36516 , w_36517 , w_36518 , w_36519 , w_36520 , w_36521 , w_36522 , w_36523 , w_36524 , w_36525 , 
		w_36526 , w_36527 , w_36528 , w_36529 , w_36530 , w_36531 , w_36532 , w_36533 , w_36534 , w_36535 , 
		w_36536 , w_36537 , w_36538 , w_36539 , w_36540 , w_36541 , w_36542 , w_36543 , w_36544 , w_36545 , 
		w_36546 , w_36547 , w_36548 , w_36549 , w_36550 , w_36551 , w_36552 , w_36553 , w_36554 , w_36555 , 
		w_36556 , w_36557 , w_36558 , w_36559 , w_36560 , w_36561 , w_36562 , w_36563 , w_36564 , w_36565 , 
		w_36566 , w_36567 , w_36568 , w_36569 , w_36570 , w_36571 , w_36572 , w_36573 , w_36574 , w_36575 , 
		w_36576 , w_36577 , w_36578 , w_36579 , w_36580 , w_36581 , w_36582 , w_36583 , w_36584 , w_36585 , 
		w_36586 , w_36587 , w_36588 , w_36589 , w_36590 , w_36591 , w_36592 , w_36593 , w_36594 , w_36595 , 
		w_36596 , w_36597 , w_36598 , w_36599 , w_36600 , w_36601 , w_36602 , w_36603 , w_36604 , w_36605 , 
		w_36606 , w_36607 , w_36608 , w_36609 , w_36610 , w_36611 , w_36612 , w_36613 , w_36614 , w_36615 , 
		w_36616 , w_36617 , w_36618 , w_36619 , w_36620 , w_36621 , w_36622 , w_36623 , w_36624 , w_36625 , 
		w_36626 , w_36627 , w_36628 , w_36629 , w_36630 , w_36631 , w_36632 , w_36633 , w_36634 , w_36635 , 
		w_36636 , w_36637 , w_36638 , w_36639 , w_36640 , w_36641 , w_36642 , w_36643 , w_36644 , w_36645 , 
		w_36646 , w_36647 , w_36648 , w_36649 , w_36650 , w_36651 , w_36652 , w_36653 , w_36654 , w_36655 , 
		w_36656 , w_36657 , w_36658 , w_36659 , w_36660 , w_36661 , w_36662 , w_36663 , w_36664 , w_36665 , 
		w_36666 , w_36667 , w_36668 , w_36669 , w_36670 , w_36671 , w_36672 , w_36673 , w_36674 , w_36675 , 
		w_36676 , w_36677 , w_36678 , w_36679 , w_36680 , w_36681 , w_36682 , w_36683 , w_36684 , w_36685 , 
		w_36686 , w_36687 , w_36688 , w_36689 , w_36690 , w_36691 , w_36692 , w_36693 , w_36694 , w_36695 , 
		w_36696 , w_36697 , w_36698 , w_36699 , w_36700 , w_36701 , w_36702 , w_36703 , w_36704 , w_36705 , 
		w_36706 , w_36707 , w_36708 , w_36709 , w_36710 , w_36711 , w_36712 , w_36713 , w_36714 , w_36715 , 
		w_36716 , w_36717 , w_36718 , w_36719 , w_36720 , w_36721 , w_36722 , w_36723 , w_36724 , w_36725 , 
		w_36726 , w_36727 , w_36728 , w_36729 , w_36730 , w_36731 , w_36732 , w_36733 , w_36734 , w_36735 , 
		w_36736 , w_36737 , w_36738 , w_36739 , w_36740 , w_36741 , w_36742 , w_36743 , w_36744 , w_36745 , 
		w_36746 , w_36747 , w_36748 , w_36749 , w_36750 , w_36751 , w_36752 , w_36753 , w_36754 , w_36755 , 
		w_36756 , w_36757 , w_36758 , w_36759 , w_36760 , w_36761 , w_36762 , w_36763 , w_36764 , w_36765 , 
		w_36766 , w_36767 , w_36768 , w_36769 , w_36770 , w_36771 , w_36772 , w_36773 , w_36774 , w_36775 , 
		w_36776 , w_36777 , w_36778 , w_36779 , w_36780 , w_36781 , w_36782 , w_36783 , w_36784 , w_36785 , 
		w_36786 , w_36787 , w_36788 , w_36789 , w_36790 , w_36791 , w_36792 , w_36793 , w_36794 , w_36795 , 
		w_36796 , w_36797 , w_36798 , w_36799 , w_36800 , w_36801 , w_36802 , w_36803 , w_36804 , w_36805 , 
		w_36806 , w_36807 , w_36808 , w_36809 , w_36810 , w_36811 , w_36812 , w_36813 , w_36814 , w_36815 , 
		w_36816 , w_36817 , w_36818 , w_36819 , w_36820 , w_36821 , w_36822 , w_36823 , w_36824 , w_36825 , 
		w_36826 , w_36827 , w_36828 , w_36829 , w_36830 , w_36831 , w_36832 , w_36833 , w_36834 , w_36835 , 
		w_36836 , w_36837 , w_36838 , w_36839 , w_36840 , w_36841 , w_36842 , w_36843 , w_36844 , w_36845 , 
		w_36846 , w_36847 , w_36848 , w_36849 , w_36850 , w_36851 , w_36852 , w_36853 , w_36854 , w_36855 , 
		w_36856 , w_36857 , w_36858 , w_36859 , w_36860 , w_36861 , w_36862 , w_36863 , w_36864 , w_36865 , 
		w_36866 , w_36867 , w_36868 , w_36869 , w_36870 , w_36871 , w_36872 , w_36873 , w_36874 , w_36875 , 
		w_36876 , w_36877 , w_36878 , w_36879 , w_36880 , w_36881 , w_36882 , w_36883 , w_36884 , w_36885 , 
		w_36886 , w_36887 , w_36888 , w_36889 , w_36890 , w_36891 , w_36892 , w_36893 , w_36894 , w_36895 , 
		w_36896 , w_36897 , w_36898 , w_36899 , w_36900 , w_36901 , w_36902 , w_36903 , w_36904 , w_36905 , 
		w_36906 , w_36907 , w_36908 , w_36909 , w_36910 , w_36911 , w_36912 , w_36913 , w_36914 , w_36915 , 
		w_36916 , w_36917 , w_36918 , w_36919 , w_36920 , w_36921 , w_36922 , w_36923 , w_36924 , w_36925 , 
		w_36926 , w_36927 , w_36928 , w_36929 , w_36930 , w_36931 , w_36932 , w_36933 , w_36934 , w_36935 , 
		w_36936 , w_36937 , w_36938 , w_36939 , w_36940 , w_36941 , w_36942 , w_36943 , w_36944 , w_36945 , 
		w_36946 , w_36947 , w_36948 , w_36949 , w_36950 , w_36951 , w_36952 , w_36953 , w_36954 , w_36955 , 
		w_36956 , w_36957 , w_36958 , w_36959 , w_36960 , w_36961 , w_36962 , w_36963 , w_36964 , w_36965 , 
		w_36966 , w_36967 , w_36968 , w_36969 , w_36970 , w_36971 , w_36972 , w_36973 , w_36974 , w_36975 , 
		w_36976 , w_36977 , w_36978 , w_36979 , w_36980 , w_36981 , w_36982 , w_36983 , w_36984 , w_36985 , 
		w_36986 , w_36987 , w_36988 , w_36989 , w_36990 , w_36991 , w_36992 , w_36993 , w_36994 , w_36995 , 
		w_36996 , w_36997 , w_36998 , w_36999 , w_37000 , w_37001 , w_37002 , w_37003 , w_37004 , w_37005 , 
		w_37006 , w_37007 , w_37008 , w_37009 , w_37010 , w_37011 , w_37012 , w_37013 , w_37014 , w_37015 , 
		w_37016 , w_37017 , w_37018 , w_37019 , w_37020 , w_37021 , w_37022 , w_37023 , w_37024 , w_37025 , 
		w_37026 , w_37027 , w_37028 , w_37029 , w_37030 , w_37031 , w_37032 , w_37033 , w_37034 , w_37035 , 
		w_37036 , w_37037 , w_37038 , w_37039 , w_37040 , w_37041 , w_37042 , w_37043 , w_37044 , w_37045 , 
		w_37046 , w_37047 , w_37048 , w_37049 , w_37050 , w_37051 , w_37052 , w_37053 , w_37054 , w_37055 , 
		w_37056 , w_37057 , w_37058 , w_37059 , w_37060 , w_37061 , w_37062 , w_37063 , w_37064 , w_37065 , 
		w_37066 , w_37067 , w_37068 , w_37069 , w_37070 , w_37071 , w_37072 , w_37073 , w_37074 , w_37075 , 
		w_37076 , w_37077 , w_37078 , w_37079 , w_37080 , w_37081 , w_37082 , w_37083 , w_37084 , w_37085 , 
		w_37086 , w_37087 , w_37088 , w_37089 , w_37090 , w_37091 , w_37092 , w_37093 , w_37094 , w_37095 , 
		w_37096 , w_37097 , w_37098 , w_37099 , w_37100 , w_37101 , w_37102 , w_37103 , w_37104 , w_37105 , 
		w_37106 , w_37107 , w_37108 , w_37109 , w_37110 , w_37111 , w_37112 , w_37113 , w_37114 , w_37115 , 
		w_37116 , w_37117 , w_37118 , w_37119 , w_37120 , w_37121 , w_37122 , w_37123 , w_37124 , w_37125 , 
		w_37126 , w_37127 , w_37128 , w_37129 , w_37130 , w_37131 , w_37132 , w_37133 , w_37134 , w_37135 , 
		w_37136 , w_37137 , w_37138 , w_37139 , w_37140 , w_37141 , w_37142 , w_37143 , w_37144 , w_37145 , 
		w_37146 , w_37147 , w_37148 , w_37149 , w_37150 , w_37151 , w_37152 , w_37153 , w_37154 , w_37155 , 
		w_37156 , w_37157 , w_37158 , w_37159 , w_37160 , w_37161 , w_37162 , w_37163 , w_37164 , w_37165 , 
		w_37166 , w_37167 , w_37168 , w_37169 , w_37170 , w_37171 , w_37172 , w_37173 , w_37174 , w_37175 , 
		w_37176 , w_37177 , w_37178 , w_37179 , w_37180 , w_37181 , w_37182 , w_37183 , w_37184 , w_37185 , 
		w_37186 , w_37187 , w_37188 , w_37189 , w_37190 , w_37191 , w_37192 , w_37193 , w_37194 , w_37195 , 
		w_37196 , w_37197 , w_37198 , w_37199 , w_37200 , w_37201 , w_37202 , w_37203 , w_37204 , w_37205 , 
		w_37206 , w_37207 , w_37208 , w_37209 , w_37210 , w_37211 , w_37212 , w_37213 , w_37214 , w_37215 , 
		w_37216 , w_37217 , w_37218 , w_37219 , w_37220 , w_37221 , w_37222 , w_37223 , w_37224 , w_37225 , 
		w_37226 , w_37227 , w_37228 , w_37229 , w_37230 , w_37231 , w_37232 , w_37233 , w_37234 , w_37235 , 
		w_37236 , w_37237 , w_37238 , w_37239 , w_37240 , w_37241 , w_37242 , w_37243 , w_37244 , w_37245 , 
		w_37246 , w_37247 , w_37248 , w_37249 , w_37250 , w_37251 , w_37252 , w_37253 , w_37254 , w_37255 , 
		w_37256 , w_37257 , w_37258 , w_37259 , w_37260 , w_37261 , w_37262 , w_37263 , w_37264 , w_37265 , 
		w_37266 , w_37267 , w_37268 , w_37269 , w_37270 , w_37271 , w_37272 , w_37273 , w_37274 , w_37275 , 
		w_37276 , w_37277 , w_37278 , w_37279 , w_37280 , w_37281 , w_37282 , w_37283 , w_37284 , w_37285 , 
		w_37286 , w_37287 , w_37288 , w_37289 , w_37290 , w_37291 , w_37292 , w_37293 , w_37294 , w_37295 , 
		w_37296 , w_37297 , w_37298 , w_37299 , w_37300 , w_37301 , w_37302 , w_37303 , w_37304 , w_37305 , 
		w_37306 , w_37307 , w_37308 , w_37309 , w_37310 , w_37311 , w_37312 , w_37313 , w_37314 , w_37315 , 
		w_37316 , w_37317 , w_37318 , w_37319 , w_37320 , w_37321 , w_37322 , w_37323 , w_37324 , w_37325 , 
		w_37326 , w_37327 , w_37328 , w_37329 , w_37330 , w_37331 , w_37332 , w_37333 , w_37334 , w_37335 , 
		w_37336 , w_37337 , w_37338 , w_37339 , w_37340 , w_37341 , w_37342 , w_37343 , w_37344 , w_37345 , 
		w_37346 , w_37347 , w_37348 , w_37349 , w_37350 , w_37351 , w_37352 , w_37353 , w_37354 , w_37355 , 
		w_37356 , w_37357 , w_37358 , w_37359 , w_37360 , w_37361 , w_37362 , w_37363 , w_37364 , w_37365 , 
		w_37366 , w_37367 , w_37368 , w_37369 , w_37370 , w_37371 , w_37372 , w_37373 , w_37374 , w_37375 , 
		w_37376 , w_37377 , w_37378 , w_37379 , w_37380 , w_37381 , w_37382 , w_37383 , w_37384 , w_37385 , 
		w_37386 , w_37387 , w_37388 , w_37389 , w_37390 , w_37391 , w_37392 , w_37393 , w_37394 , w_37395 , 
		w_37396 , w_37397 , w_37398 , w_37399 , w_37400 , w_37401 , w_37402 , w_37403 , w_37404 , w_37405 , 
		w_37406 , w_37407 , w_37408 , w_37409 , w_37410 , w_37411 , w_37412 , w_37413 , w_37414 , w_37415 , 
		w_37416 , w_37417 , w_37418 , w_37419 , w_37420 , w_37421 , w_37422 , w_37423 , w_37424 , w_37425 , 
		w_37426 , w_37427 , w_37428 , w_37429 , w_37430 , w_37431 , w_37432 , w_37433 , w_37434 , w_37435 , 
		w_37436 , w_37437 , w_37438 , w_37439 , w_37440 , w_37441 , w_37442 , w_37443 , w_37444 , w_37445 , 
		w_37446 , w_37447 , w_37448 , w_37449 , w_37450 , w_37451 , w_37452 , w_37453 , w_37454 , w_37455 , 
		w_37456 , w_37457 , w_37458 , w_37459 , w_37460 , w_37461 , w_37462 , w_37463 , w_37464 , w_37465 , 
		w_37466 , w_37467 , w_37468 , w_37469 , w_37470 , w_37471 , w_37472 , w_37473 , w_37474 , w_37475 , 
		w_37476 , w_37477 , w_37478 , w_37479 , w_37480 , w_37481 , w_37482 , w_37483 , w_37484 , w_37485 , 
		w_37486 , w_37487 , w_37488 , w_37489 , w_37490 , w_37491 , w_37492 , w_37493 , w_37494 , w_37495 , 
		w_37496 , w_37497 , w_37498 , w_37499 , w_37500 , w_37501 , w_37502 , w_37503 , w_37504 , w_37505 , 
		w_37506 , w_37507 , w_37508 , w_37509 , w_37510 , w_37511 , w_37512 , w_37513 , w_37514 , w_37515 , 
		w_37516 , w_37517 , w_37518 , w_37519 , w_37520 , w_37521 , w_37522 , w_37523 , w_37524 , w_37525 , 
		w_37526 , w_37527 , w_37528 , w_37529 , w_37530 , w_37531 , w_37532 , w_37533 , w_37534 , w_37535 , 
		w_37536 , w_37537 , w_37538 , w_37539 , w_37540 , w_37541 , w_37542 , w_37543 , w_37544 , w_37545 , 
		w_37546 , w_37547 , w_37548 , w_37549 , w_37550 , w_37551 , w_37552 , w_37553 , w_37554 , w_37555 , 
		w_37556 , w_37557 , w_37558 , w_37559 , w_37560 , w_37561 , w_37562 , w_37563 , w_37564 , w_37565 , 
		w_37566 , w_37567 , w_37568 , w_37569 , w_37570 , w_37571 , w_37572 , w_37573 , w_37574 , w_37575 , 
		w_37576 , w_37577 , w_37578 , w_37579 , w_37580 , w_37581 , w_37582 , w_37583 , w_37584 , w_37585 , 
		w_37586 , w_37587 , w_37588 , w_37589 , w_37590 , w_37591 , w_37592 , w_37593 , w_37594 , w_37595 , 
		w_37596 , w_37597 , w_37598 , w_37599 , w_37600 , w_37601 , w_37602 , w_37603 , w_37604 , w_37605 , 
		w_37606 , w_37607 , w_37608 , w_37609 , w_37610 , w_37611 , w_37612 , w_37613 , w_37614 , w_37615 , 
		w_37616 , w_37617 , w_37618 , w_37619 , w_37620 , w_37621 , w_37622 , w_37623 , w_37624 , w_37625 , 
		w_37626 , w_37627 , w_37628 , w_37629 , w_37630 , w_37631 , w_37632 , w_37633 , w_37634 , w_37635 , 
		w_37636 , w_37637 , w_37638 , w_37639 , w_37640 , w_37641 , w_37642 , w_37643 , w_37644 , w_37645 , 
		w_37646 , w_37647 , w_37648 , w_37649 , w_37650 , w_37651 , w_37652 , w_37653 , w_37654 , w_37655 , 
		w_37656 , w_37657 , w_37658 , w_37659 , w_37660 , w_37661 , w_37662 , w_37663 , w_37664 , w_37665 , 
		w_37666 , w_37667 , w_37668 , w_37669 , w_37670 , w_37671 , w_37672 , w_37673 , w_37674 , w_37675 , 
		w_37676 , w_37677 , w_37678 , w_37679 , w_37680 , w_37681 , w_37682 , w_37683 , w_37684 , w_37685 , 
		w_37686 , w_37687 , w_37688 , w_37689 , w_37690 , w_37691 , w_37692 , w_37693 , w_37694 , w_37695 , 
		w_37696 , w_37697 , w_37698 , w_37699 , w_37700 , w_37701 , w_37702 , w_37703 , w_37704 , w_37705 , 
		w_37706 , w_37707 , w_37708 , w_37709 , w_37710 , w_37711 , w_37712 , w_37713 , w_37714 , w_37715 , 
		w_37716 , w_37717 , w_37718 , w_37719 , w_37720 , w_37721 , w_37722 , w_37723 , w_37724 , w_37725 , 
		w_37726 , w_37727 , w_37728 , w_37729 , w_37730 , w_37731 , w_37732 , w_37733 , w_37734 , w_37735 , 
		w_37736 , w_37737 , w_37738 , w_37739 , w_37740 , w_37741 , w_37742 , w_37743 , w_37744 , w_37745 , 
		w_37746 , w_37747 , w_37748 , w_37749 , w_37750 , w_37751 , w_37752 , w_37753 , w_37754 , w_37755 , 
		w_37756 , w_37757 , w_37758 , w_37759 , w_37760 , w_37761 , w_37762 , w_37763 , w_37764 , w_37765 , 
		w_37766 , w_37767 , w_37768 , w_37769 , w_37770 , w_37771 , w_37772 , w_37773 , w_37774 , w_37775 , 
		w_37776 , w_37777 , w_37778 , w_37779 , w_37780 , w_37781 , w_37782 , w_37783 , w_37784 , w_37785 , 
		w_37786 , w_37787 , w_37788 , w_37789 , w_37790 , w_37791 , w_37792 , w_37793 , w_37794 , w_37795 , 
		w_37796 , w_37797 , w_37798 , w_37799 , w_37800 , w_37801 , w_37802 , w_37803 , w_37804 , w_37805 , 
		w_37806 , w_37807 , w_37808 , w_37809 , w_37810 , w_37811 , w_37812 , w_37813 , w_37814 , w_37815 , 
		w_37816 , w_37817 , w_37818 , w_37819 , w_37820 , w_37821 , w_37822 , w_37823 , w_37824 , w_37825 , 
		w_37826 , w_37827 , w_37828 , w_37829 , w_37830 , w_37831 , w_37832 , w_37833 , w_37834 , w_37835 , 
		w_37836 , w_37837 , w_37838 , w_37839 , w_37840 , w_37841 , w_37842 , w_37843 , w_37844 , w_37845 , 
		w_37846 , w_37847 , w_37848 , w_37849 , w_37850 , w_37851 , w_37852 , w_37853 , w_37854 , w_37855 , 
		w_37856 , w_37857 , w_37858 , w_37859 , w_37860 , w_37861 , w_37862 , w_37863 , w_37864 , w_37865 , 
		w_37866 , w_37867 , w_37868 , w_37869 , w_37870 , w_37871 , w_37872 , w_37873 , w_37874 , w_37875 , 
		w_37876 , w_37877 , w_37878 , w_37879 , w_37880 , w_37881 , w_37882 , w_37883 , w_37884 , w_37885 , 
		w_37886 , w_37887 , w_37888 , w_37889 , w_37890 , w_37891 , w_37892 , w_37893 , w_37894 , w_37895 , 
		w_37896 , w_37897 , w_37898 , w_37899 , w_37900 , w_37901 , w_37902 , w_37903 , w_37904 , w_37905 , 
		w_37906 , w_37907 , w_37908 , w_37909 , w_37910 , w_37911 , w_37912 , w_37913 , w_37914 , w_37915 , 
		w_37916 , w_37917 , w_37918 , w_37919 , w_37920 , w_37921 , w_37922 , w_37923 , w_37924 , w_37925 , 
		w_37926 , w_37927 , w_37928 , w_37929 , w_37930 , w_37931 , w_37932 , w_37933 , w_37934 , w_37935 , 
		w_37936 , w_37937 , w_37938 , w_37939 , w_37940 , w_37941 , w_37942 , w_37943 , w_37944 , w_37945 , 
		w_37946 , w_37947 , w_37948 , w_37949 , w_37950 , w_37951 , w_37952 , w_37953 , w_37954 , w_37955 , 
		w_37956 , w_37957 , w_37958 , w_37959 , w_37960 , w_37961 , w_37962 , w_37963 , w_37964 , w_37965 , 
		w_37966 , w_37967 , w_37968 , w_37969 , w_37970 , w_37971 , w_37972 , w_37973 , w_37974 , w_37975 , 
		w_37976 , w_37977 , w_37978 , w_37979 , w_37980 , w_37981 , w_37982 , w_37983 , w_37984 , w_37985 , 
		w_37986 , w_37987 , w_37988 , w_37989 , w_37990 , w_37991 , w_37992 , w_37993 , w_37994 , w_37995 , 
		w_37996 , w_37997 , w_37998 , w_37999 , w_38000 , w_38001 , w_38002 , w_38003 , w_38004 , w_38005 , 
		w_38006 , w_38007 , w_38008 , w_38009 , w_38010 , w_38011 , w_38012 , w_38013 , w_38014 , w_38015 , 
		w_38016 , w_38017 , w_38018 , w_38019 , w_38020 , w_38021 , w_38022 , w_38023 , w_38024 , w_38025 , 
		w_38026 , w_38027 , w_38028 , w_38029 , w_38030 , w_38031 , w_38032 , w_38033 , w_38034 , w_38035 , 
		w_38036 , w_38037 , w_38038 , w_38039 , w_38040 , w_38041 , w_38042 , w_38043 , w_38044 , w_38045 , 
		w_38046 , w_38047 , w_38048 , w_38049 , w_38050 , w_38051 , w_38052 , w_38053 , w_38054 , w_38055 , 
		w_38056 , w_38057 , w_38058 , w_38059 , w_38060 , w_38061 , w_38062 , w_38063 , w_38064 , w_38065 , 
		w_38066 , w_38067 , w_38068 , w_38069 , w_38070 , w_38071 , w_38072 , w_38073 , w_38074 , w_38075 , 
		w_38076 , w_38077 , w_38078 , w_38079 , w_38080 , w_38081 , w_38082 , w_38083 , w_38084 , w_38085 , 
		w_38086 , w_38087 , w_38088 , w_38089 , w_38090 , w_38091 , w_38092 , w_38093 , w_38094 , w_38095 , 
		w_38096 , w_38097 , w_38098 , w_38099 , w_38100 , w_38101 , w_38102 , w_38103 , w_38104 , w_38105 , 
		w_38106 , w_38107 , w_38108 , w_38109 , w_38110 , w_38111 , w_38112 , w_38113 , w_38114 , w_38115 , 
		w_38116 , w_38117 , w_38118 , w_38119 , w_38120 , w_38121 , w_38122 , w_38123 , w_38124 , w_38125 , 
		w_38126 , w_38127 , w_38128 , w_38129 , w_38130 , w_38131 , w_38132 , w_38133 , w_38134 , w_38135 , 
		w_38136 , w_38137 , w_38138 , w_38139 , w_38140 , w_38141 , w_38142 , w_38143 , w_38144 , w_38145 , 
		w_38146 , w_38147 , w_38148 , w_38149 , w_38150 , w_38151 , w_38152 , w_38153 , w_38154 , w_38155 , 
		w_38156 , w_38157 , w_38158 , w_38159 , w_38160 , w_38161 , w_38162 , w_38163 , w_38164 , w_38165 , 
		w_38166 , w_38167 , w_38168 , w_38169 , w_38170 , w_38171 , w_38172 , w_38173 , w_38174 , w_38175 , 
		w_38176 , w_38177 , w_38178 , w_38179 , w_38180 , w_38181 , w_38182 , w_38183 , w_38184 , w_38185 , 
		w_38186 , w_38187 , w_38188 , w_38189 , w_38190 , w_38191 , w_38192 , w_38193 , w_38194 , w_38195 , 
		w_38196 , w_38197 , w_38198 , w_38199 , w_38200 , w_38201 , w_38202 , w_38203 , w_38204 , w_38205 , 
		w_38206 , w_38207 , w_38208 , w_38209 , w_38210 , w_38211 , w_38212 , w_38213 , w_38214 , w_38215 , 
		w_38216 , w_38217 , w_38218 , w_38219 , w_38220 , w_38221 , w_38222 , w_38223 , w_38224 , w_38225 , 
		w_38226 , w_38227 , w_38228 , w_38229 , w_38230 , w_38231 , w_38232 , w_38233 , w_38234 , w_38235 , 
		w_38236 , w_38237 , w_38238 , w_38239 , w_38240 , w_38241 , w_38242 , w_38243 , w_38244 , w_38245 , 
		w_38246 , w_38247 , w_38248 , w_38249 , w_38250 , w_38251 , w_38252 , w_38253 , w_38254 , w_38255 , 
		w_38256 , w_38257 , w_38258 , w_38259 , w_38260 , w_38261 , w_38262 , w_38263 , w_38264 , w_38265 , 
		w_38266 , w_38267 , w_38268 , w_38269 , w_38270 , w_38271 , w_38272 , w_38273 , w_38274 , w_38275 , 
		w_38276 , w_38277 , w_38278 , w_38279 , w_38280 , w_38281 , w_38282 , w_38283 , w_38284 , w_38285 , 
		w_38286 , w_38287 , w_38288 , w_38289 , w_38290 , w_38291 , w_38292 , w_38293 , w_38294 , w_38295 , 
		w_38296 , w_38297 , w_38298 , w_38299 , w_38300 , w_38301 , w_38302 , w_38303 , w_38304 , w_38305 , 
		w_38306 , w_38307 , w_38308 , w_38309 , w_38310 , w_38311 , w_38312 , w_38313 , w_38314 , w_38315 , 
		w_38316 , w_38317 , w_38318 , w_38319 , w_38320 , w_38321 , w_38322 , w_38323 , w_38324 , w_38325 , 
		w_38326 , w_38327 , w_38328 , w_38329 , w_38330 , w_38331 , w_38332 , w_38333 , w_38334 , w_38335 , 
		w_38336 , w_38337 , w_38338 , w_38339 , w_38340 , w_38341 , w_38342 , w_38343 , w_38344 , w_38345 , 
		w_38346 , w_38347 , w_38348 , w_38349 , w_38350 , w_38351 , w_38352 , w_38353 , w_38354 , w_38355 , 
		w_38356 , w_38357 , w_38358 , w_38359 , w_38360 , w_38361 , w_38362 , w_38363 , w_38364 , w_38365 , 
		w_38366 , w_38367 , w_38368 , w_38369 , w_38370 , w_38371 , w_38372 , w_38373 , w_38374 , w_38375 , 
		w_38376 , w_38377 , w_38378 , w_38379 , w_38380 , w_38381 , w_38382 , w_38383 , w_38384 , w_38385 , 
		w_38386 , w_38387 , w_38388 , w_38389 , w_38390 , w_38391 , w_38392 , w_38393 , w_38394 , w_38395 , 
		w_38396 , w_38397 , w_38398 , w_38399 , w_38400 , w_38401 , w_38402 , w_38403 , w_38404 , w_38405 , 
		w_38406 , w_38407 , w_38408 , w_38409 , w_38410 , w_38411 , w_38412 , w_38413 , w_38414 , w_38415 , 
		w_38416 , w_38417 , w_38418 , w_38419 , w_38420 , w_38421 , w_38422 , w_38423 , w_38424 , w_38425 , 
		w_38426 , w_38427 , w_38428 , w_38429 , w_38430 , w_38431 , w_38432 , w_38433 , w_38434 , w_38435 , 
		w_38436 , w_38437 , w_38438 , w_38439 , w_38440 , w_38441 , w_38442 , w_38443 , w_38444 , w_38445 , 
		w_38446 , w_38447 , w_38448 , w_38449 , w_38450 , w_38451 , w_38452 , w_38453 , w_38454 , w_38455 , 
		w_38456 , w_38457 , w_38458 , w_38459 , w_38460 , w_38461 , w_38462 , w_38463 , w_38464 , w_38465 , 
		w_38466 , w_38467 , w_38468 , w_38469 , w_38470 , w_38471 , w_38472 , w_38473 , w_38474 , w_38475 , 
		w_38476 , w_38477 , w_38478 , w_38479 , w_38480 , w_38481 , w_38482 , w_38483 , w_38484 , w_38485 , 
		w_38486 , w_38487 , w_38488 , w_38489 , w_38490 , w_38491 , w_38492 , w_38493 , w_38494 , w_38495 , 
		w_38496 , w_38497 , w_38498 , w_38499 , w_38500 , w_38501 , w_38502 , w_38503 , w_38504 , w_38505 , 
		w_38506 , w_38507 , w_38508 , w_38509 , w_38510 , w_38511 , w_38512 , w_38513 , w_38514 , w_38515 , 
		w_38516 , w_38517 , w_38518 , w_38519 , w_38520 , w_38521 , w_38522 , w_38523 , w_38524 , w_38525 , 
		w_38526 , w_38527 , w_38528 , w_38529 , w_38530 , w_38531 , w_38532 , w_38533 , w_38534 , w_38535 , 
		w_38536 , w_38537 , w_38538 , w_38539 , w_38540 , w_38541 , w_38542 , w_38543 , w_38544 , w_38545 , 
		w_38546 , w_38547 , w_38548 , w_38549 , w_38550 , w_38551 , w_38552 , w_38553 , w_38554 , w_38555 , 
		w_38556 , w_38557 , w_38558 , w_38559 , w_38560 , w_38561 , w_38562 , w_38563 , w_38564 , w_38565 , 
		w_38566 , w_38567 , w_38568 , w_38569 , w_38570 , w_38571 , w_38572 , w_38573 , w_38574 , w_38575 , 
		w_38576 , w_38577 , w_38578 , w_38579 , w_38580 , w_38581 , w_38582 , w_38583 , w_38584 , w_38585 , 
		w_38586 , w_38587 , w_38588 , w_38589 , w_38590 , w_38591 , w_38592 , w_38593 , w_38594 , w_38595 , 
		w_38596 , w_38597 , w_38598 , w_38599 , w_38600 , w_38601 , w_38602 , w_38603 , w_38604 , w_38605 , 
		w_38606 , w_38607 , w_38608 , w_38609 , w_38610 , w_38611 , w_38612 , w_38613 , w_38614 , w_38615 , 
		w_38616 , w_38617 , w_38618 , w_38619 , w_38620 , w_38621 , w_38622 , w_38623 , w_38624 , w_38625 , 
		w_38626 , w_38627 , w_38628 , w_38629 , w_38630 , w_38631 , w_38632 , w_38633 , w_38634 , w_38635 , 
		w_38636 , w_38637 , w_38638 , w_38639 , w_38640 , w_38641 , w_38642 , w_38643 , w_38644 , w_38645 , 
		w_38646 , w_38647 , w_38648 , w_38649 , w_38650 , w_38651 , w_38652 , w_38653 , w_38654 , w_38655 , 
		w_38656 , w_38657 , w_38658 , w_38659 , w_38660 , w_38661 , w_38662 , w_38663 , w_38664 , w_38665 , 
		w_38666 , w_38667 , w_38668 , w_38669 , w_38670 , w_38671 , w_38672 , w_38673 , w_38674 , w_38675 , 
		w_38676 , w_38677 , w_38678 , w_38679 , w_38680 , w_38681 , w_38682 , w_38683 , w_38684 , w_38685 , 
		w_38686 , w_38687 , w_38688 , w_38689 , w_38690 , w_38691 , w_38692 , w_38693 , w_38694 , w_38695 , 
		w_38696 , w_38697 , w_38698 , w_38699 , w_38700 , w_38701 , w_38702 , w_38703 , w_38704 , w_38705 , 
		w_38706 , w_38707 , w_38708 , w_38709 , w_38710 , w_38711 , w_38712 , w_38713 , w_38714 , w_38715 , 
		w_38716 , w_38717 , w_38718 , w_38719 , w_38720 , w_38721 , w_38722 , w_38723 , w_38724 , w_38725 , 
		w_38726 , w_38727 , w_38728 , w_38729 , w_38730 , w_38731 , w_38732 , w_38733 , w_38734 , w_38735 , 
		w_38736 , w_38737 , w_38738 , w_38739 , w_38740 , w_38741 , w_38742 , w_38743 , w_38744 , w_38745 , 
		w_38746 , w_38747 , w_38748 , w_38749 , w_38750 , w_38751 , w_38752 , w_38753 , w_38754 , w_38755 , 
		w_38756 , w_38757 , w_38758 , w_38759 , w_38760 , w_38761 , w_38762 , w_38763 , w_38764 , w_38765 , 
		w_38766 , w_38767 , w_38768 , w_38769 , w_38770 , w_38771 , w_38772 , w_38773 , w_38774 , w_38775 , 
		w_38776 , w_38777 , w_38778 , w_38779 , w_38780 , w_38781 , w_38782 , w_38783 , w_38784 , w_38785 , 
		w_38786 , w_38787 , w_38788 , w_38789 , w_38790 , w_38791 , w_38792 , w_38793 , w_38794 , w_38795 , 
		w_38796 , w_38797 , w_38798 , w_38799 , w_38800 , w_38801 , w_38802 , w_38803 , w_38804 , w_38805 , 
		w_38806 , w_38807 , w_38808 , w_38809 , w_38810 , w_38811 , w_38812 , w_38813 , w_38814 , w_38815 , 
		w_38816 , w_38817 , w_38818 , w_38819 , w_38820 , w_38821 , w_38822 , w_38823 , w_38824 , w_38825 , 
		w_38826 , w_38827 , w_38828 , w_38829 , w_38830 , w_38831 , w_38832 , w_38833 , w_38834 , w_38835 , 
		w_38836 , w_38837 , w_38838 , w_38839 , w_38840 , w_38841 , w_38842 , w_38843 , w_38844 , w_38845 , 
		w_38846 , w_38847 , w_38848 , w_38849 , w_38850 , w_38851 , w_38852 , w_38853 , w_38854 , w_38855 , 
		w_38856 , w_38857 , w_38858 , w_38859 , w_38860 , w_38861 , w_38862 , w_38863 , w_38864 , w_38865 , 
		w_38866 , w_38867 , w_38868 , w_38869 , w_38870 , w_38871 , w_38872 , w_38873 , w_38874 , w_38875 , 
		w_38876 , w_38877 , w_38878 , w_38879 , w_38880 , w_38881 , w_38882 , w_38883 , w_38884 , w_38885 , 
		w_38886 , w_38887 , w_38888 , w_38889 , w_38890 , w_38891 , w_38892 , w_38893 , w_38894 , w_38895 , 
		w_38896 , w_38897 , w_38898 , w_38899 , w_38900 , w_38901 , w_38902 , w_38903 , w_38904 , w_38905 , 
		w_38906 , w_38907 , w_38908 , w_38909 , w_38910 , w_38911 , w_38912 , w_38913 , w_38914 , w_38915 , 
		w_38916 , w_38917 , w_38918 , w_38919 , w_38920 , w_38921 , w_38922 , w_38923 , w_38924 , w_38925 , 
		w_38926 , w_38927 , w_38928 , w_38929 , w_38930 , w_38931 , w_38932 , w_38933 , w_38934 , w_38935 , 
		w_38936 , w_38937 , w_38938 , w_38939 , w_38940 , w_38941 , w_38942 , w_38943 , w_38944 , w_38945 , 
		w_38946 , w_38947 , w_38948 , w_38949 , w_38950 , w_38951 , w_38952 , w_38953 , w_38954 , w_38955 , 
		w_38956 , w_38957 , w_38958 , w_38959 , w_38960 , w_38961 , w_38962 , w_38963 , w_38964 , w_38965 , 
		w_38966 , w_38967 , w_38968 , w_38969 , w_38970 , w_38971 , w_38972 , w_38973 , w_38974 , w_38975 , 
		w_38976 , w_38977 , w_38978 , w_38979 , w_38980 , w_38981 , w_38982 , w_38983 , w_38984 , w_38985 , 
		w_38986 , w_38987 , w_38988 , w_38989 , w_38990 , w_38991 , w_38992 , w_38993 , w_38994 , w_38995 , 
		w_38996 , w_38997 , w_38998 , w_38999 , w_39000 , w_39001 , w_39002 , w_39003 , w_39004 , w_39005 , 
		w_39006 , w_39007 , w_39008 , w_39009 , w_39010 , w_39011 , w_39012 , w_39013 , w_39014 , w_39015 , 
		w_39016 , w_39017 , w_39018 , w_39019 , w_39020 , w_39021 , w_39022 , w_39023 , w_39024 , w_39025 , 
		w_39026 , w_39027 , w_39028 , w_39029 , w_39030 , w_39031 , w_39032 , w_39033 , w_39034 , w_39035 , 
		w_39036 , w_39037 , w_39038 , w_39039 , w_39040 , w_39041 , w_39042 , w_39043 , w_39044 , w_39045 , 
		w_39046 , w_39047 , w_39048 , w_39049 , w_39050 , w_39051 , w_39052 , w_39053 , w_39054 , w_39055 , 
		w_39056 , w_39057 , w_39058 , w_39059 , w_39060 , w_39061 , w_39062 , w_39063 , w_39064 , w_39065 , 
		w_39066 , w_39067 , w_39068 , w_39069 , w_39070 , w_39071 , w_39072 , w_39073 , w_39074 , w_39075 , 
		w_39076 , w_39077 , w_39078 , w_39079 , w_39080 , w_39081 , w_39082 , w_39083 , w_39084 , w_39085 , 
		w_39086 , w_39087 , w_39088 , w_39089 , w_39090 , w_39091 , w_39092 , w_39093 , w_39094 , w_39095 , 
		w_39096 , w_39097 , w_39098 , w_39099 , w_39100 , w_39101 , w_39102 , w_39103 , w_39104 , w_39105 , 
		w_39106 , w_39107 , w_39108 , w_39109 , w_39110 , w_39111 , w_39112 , w_39113 , w_39114 , w_39115 , 
		w_39116 , w_39117 , w_39118 , w_39119 , w_39120 , w_39121 , w_39122 , w_39123 , w_39124 , w_39125 , 
		w_39126 , w_39127 , w_39128 , w_39129 , w_39130 , w_39131 , w_39132 , w_39133 , w_39134 , w_39135 , 
		w_39136 , w_39137 , w_39138 , w_39139 , w_39140 , w_39141 , w_39142 , w_39143 , w_39144 , w_39145 , 
		w_39146 , w_39147 , w_39148 , w_39149 , w_39150 , w_39151 , w_39152 , w_39153 , w_39154 , w_39155 , 
		w_39156 , w_39157 , w_39158 , w_39159 , w_39160 , w_39161 , w_39162 , w_39163 , w_39164 , w_39165 , 
		w_39166 , w_39167 , w_39168 , w_39169 , w_39170 , w_39171 , w_39172 , w_39173 , w_39174 , w_39175 , 
		w_39176 , w_39177 , w_39178 , w_39179 , w_39180 , w_39181 , w_39182 , w_39183 , w_39184 , w_39185 , 
		w_39186 , w_39187 , w_39188 , w_39189 , w_39190 , w_39191 , w_39192 , w_39193 , w_39194 , w_39195 , 
		w_39196 , w_39197 , w_39198 , w_39199 , w_39200 , w_39201 , w_39202 , w_39203 , w_39204 , w_39205 , 
		w_39206 , w_39207 , w_39208 , w_39209 , w_39210 , w_39211 , w_39212 , w_39213 , w_39214 , w_39215 , 
		w_39216 , w_39217 , w_39218 , w_39219 , w_39220 , w_39221 , w_39222 , w_39223 , w_39224 , w_39225 , 
		w_39226 , w_39227 , w_39228 , w_39229 , w_39230 , w_39231 , w_39232 , w_39233 , w_39234 , w_39235 , 
		w_39236 , w_39237 , w_39238 , w_39239 , w_39240 , w_39241 , w_39242 , w_39243 , w_39244 , w_39245 , 
		w_39246 , w_39247 , w_39248 , w_39249 , w_39250 , w_39251 , w_39252 , w_39253 , w_39254 , w_39255 , 
		w_39256 , w_39257 , w_39258 , w_39259 , w_39260 , w_39261 , w_39262 , w_39263 , w_39264 , w_39265 , 
		w_39266 , w_39267 , w_39268 , w_39269 , w_39270 , w_39271 , w_39272 , w_39273 , w_39274 , w_39275 , 
		w_39276 , w_39277 , w_39278 , w_39279 , w_39280 , w_39281 , w_39282 , w_39283 , w_39284 , w_39285 , 
		w_39286 , w_39287 , w_39288 , w_39289 , w_39290 , w_39291 , w_39292 , w_39293 , w_39294 , w_39295 , 
		w_39296 , w_39297 , w_39298 , w_39299 , w_39300 , w_39301 , w_39302 , w_39303 , w_39304 , w_39305 , 
		w_39306 , w_39307 , w_39308 , w_39309 , w_39310 , w_39311 , w_39312 , w_39313 , w_39314 , w_39315 , 
		w_39316 , w_39317 , w_39318 , w_39319 , w_39320 , w_39321 , w_39322 , w_39323 , w_39324 , w_39325 , 
		w_39326 , w_39327 , w_39328 , w_39329 , w_39330 , w_39331 , w_39332 , w_39333 , w_39334 , w_39335 , 
		w_39336 , w_39337 , w_39338 , w_39339 , w_39340 , w_39341 , w_39342 , w_39343 , w_39344 , w_39345 , 
		w_39346 , w_39347 , w_39348 , w_39349 , w_39350 , w_39351 , w_39352 , w_39353 , w_39354 , w_39355 , 
		w_39356 , w_39357 , w_39358 , w_39359 , w_39360 , w_39361 , w_39362 , w_39363 , w_39364 , w_39365 , 
		w_39366 , w_39367 , w_39368 , w_39369 , w_39370 , w_39371 , w_39372 , w_39373 , w_39374 , w_39375 , 
		w_39376 , w_39377 , w_39378 , w_39379 , w_39380 , w_39381 , w_39382 , w_39383 , w_39384 , w_39385 , 
		w_39386 , w_39387 , w_39388 , w_39389 , w_39390 , w_39391 , w_39392 , w_39393 , w_39394 , w_39395 , 
		w_39396 , w_39397 , w_39398 , w_39399 , w_39400 , w_39401 , w_39402 , w_39403 , w_39404 , w_39405 , 
		w_39406 , w_39407 , w_39408 , w_39409 , w_39410 , w_39411 , w_39412 , w_39413 , w_39414 , w_39415 , 
		w_39416 , w_39417 , w_39418 , w_39419 , w_39420 , w_39421 , w_39422 , w_39423 , w_39424 , w_39425 , 
		w_39426 , w_39427 , w_39428 , w_39429 , w_39430 , w_39431 , w_39432 , w_39433 , w_39434 , w_39435 , 
		w_39436 , w_39437 , w_39438 , w_39439 , w_39440 , w_39441 , w_39442 , w_39443 , w_39444 , w_39445 , 
		w_39446 , w_39447 , w_39448 , w_39449 , w_39450 , w_39451 , w_39452 , w_39453 , w_39454 , w_39455 , 
		w_39456 , w_39457 , w_39458 , w_39459 , w_39460 , w_39461 , w_39462 , w_39463 , w_39464 , w_39465 , 
		w_39466 , w_39467 , w_39468 , w_39469 , w_39470 , w_39471 , w_39472 , w_39473 , w_39474 , w_39475 , 
		w_39476 , w_39477 , w_39478 , w_39479 , w_39480 , w_39481 , w_39482 , w_39483 , w_39484 , w_39485 , 
		w_39486 , w_39487 , w_39488 , w_39489 , w_39490 , w_39491 , w_39492 , w_39493 , w_39494 , w_39495 , 
		w_39496 , w_39497 , w_39498 , w_39499 , w_39500 , w_39501 , w_39502 , w_39503 , w_39504 , w_39505 , 
		w_39506 , w_39507 , w_39508 , w_39509 , w_39510 , w_39511 , w_39512 , w_39513 , w_39514 , w_39515 , 
		w_39516 , w_39517 , w_39518 , w_39519 , w_39520 , w_39521 , w_39522 , w_39523 , w_39524 , w_39525 , 
		w_39526 , w_39527 , w_39528 , w_39529 , w_39530 , w_39531 , w_39532 , w_39533 , w_39534 , w_39535 , 
		w_39536 , w_39537 , w_39538 , w_39539 , w_39540 , w_39541 , w_39542 , w_39543 , w_39544 , w_39545 , 
		w_39546 , w_39547 , w_39548 , w_39549 , w_39550 , w_39551 , w_39552 , w_39553 , w_39554 , w_39555 , 
		w_39556 , w_39557 , w_39558 , w_39559 , w_39560 , w_39561 , w_39562 , w_39563 , w_39564 , w_39565 , 
		w_39566 , w_39567 , w_39568 , w_39569 , w_39570 , w_39571 , w_39572 , w_39573 , w_39574 , w_39575 , 
		w_39576 , w_39577 , w_39578 , w_39579 , w_39580 , w_39581 , w_39582 , w_39583 , w_39584 , w_39585 , 
		w_39586 , w_39587 , w_39588 , w_39589 , w_39590 , w_39591 , w_39592 , w_39593 , w_39594 , w_39595 , 
		w_39596 , w_39597 , w_39598 , w_39599 , w_39600 , w_39601 , w_39602 , w_39603 , w_39604 , w_39605 , 
		w_39606 , w_39607 , w_39608 , w_39609 , w_39610 , w_39611 , w_39612 , w_39613 , w_39614 , w_39615 , 
		w_39616 , w_39617 , w_39618 , w_39619 , w_39620 , w_39621 , w_39622 , w_39623 , w_39624 , w_39625 , 
		w_39626 , w_39627 , w_39628 , w_39629 , w_39630 , w_39631 , w_39632 , w_39633 , w_39634 , w_39635 , 
		w_39636 , w_39637 , w_39638 , w_39639 , w_39640 , w_39641 , w_39642 , w_39643 , w_39644 , w_39645 , 
		w_39646 , w_39647 , w_39648 , w_39649 , w_39650 , w_39651 , w_39652 , w_39653 , w_39654 , w_39655 , 
		w_39656 , w_39657 , w_39658 , w_39659 , w_39660 , w_39661 , w_39662 , w_39663 , w_39664 , w_39665 , 
		w_39666 , w_39667 , w_39668 , w_39669 , w_39670 , w_39671 , w_39672 , w_39673 , w_39674 , w_39675 , 
		w_39676 , w_39677 , w_39678 , w_39679 , w_39680 , w_39681 , w_39682 , w_39683 , w_39684 , w_39685 , 
		w_39686 , w_39687 , w_39688 , w_39689 , w_39690 , w_39691 , w_39692 , w_39693 , w_39694 , w_39695 , 
		w_39696 , w_39697 , w_39698 , w_39699 , w_39700 , w_39701 , w_39702 , w_39703 , w_39704 , w_39705 , 
		w_39706 , w_39707 , w_39708 , w_39709 , w_39710 , w_39711 , w_39712 , w_39713 , w_39714 , w_39715 , 
		w_39716 , w_39717 , w_39718 , w_39719 , w_39720 , w_39721 , w_39722 , w_39723 , w_39724 , w_39725 , 
		w_39726 , w_39727 , w_39728 , w_39729 , w_39730 , w_39731 , w_39732 , w_39733 , w_39734 , w_39735 , 
		w_39736 , w_39737 , w_39738 , w_39739 , w_39740 , w_39741 , w_39742 , w_39743 , w_39744 , w_39745 , 
		w_39746 , w_39747 , w_39748 , w_39749 , w_39750 , w_39751 , w_39752 , w_39753 , w_39754 , w_39755 , 
		w_39756 , w_39757 , w_39758 , w_39759 , w_39760 , w_39761 , w_39762 , w_39763 , w_39764 , w_39765 , 
		w_39766 , w_39767 , w_39768 , w_39769 , w_39770 , w_39771 , w_39772 , w_39773 , w_39774 , w_39775 , 
		w_39776 , w_39777 , w_39778 , w_39779 , w_39780 , w_39781 , w_39782 , w_39783 , w_39784 , w_39785 , 
		w_39786 , w_39787 , w_39788 , w_39789 , w_39790 , w_39791 , w_39792 , w_39793 , w_39794 , w_39795 , 
		w_39796 , w_39797 , w_39798 , w_39799 , w_39800 , w_39801 , w_39802 , w_39803 , w_39804 , w_39805 , 
		w_39806 , w_39807 , w_39808 , w_39809 , w_39810 , w_39811 , w_39812 , w_39813 , w_39814 , w_39815 , 
		w_39816 , w_39817 , w_39818 , w_39819 , w_39820 , w_39821 , w_39822 , w_39823 , w_39824 , w_39825 , 
		w_39826 , w_39827 , w_39828 , w_39829 , w_39830 , w_39831 , w_39832 , w_39833 , w_39834 , w_39835 , 
		w_39836 , w_39837 , w_39838 , w_39839 , w_39840 , w_39841 , w_39842 , w_39843 , w_39844 , w_39845 , 
		w_39846 , w_39847 , w_39848 , w_39849 , w_39850 , w_39851 , w_39852 , w_39853 , w_39854 , w_39855 , 
		w_39856 , w_39857 , w_39858 , w_39859 , w_39860 , w_39861 , w_39862 , w_39863 , w_39864 , w_39865 , 
		w_39866 , w_39867 , w_39868 , w_39869 , w_39870 , w_39871 , w_39872 , w_39873 , w_39874 , w_39875 , 
		w_39876 , w_39877 , w_39878 , w_39879 , w_39880 , w_39881 , w_39882 , w_39883 , w_39884 , w_39885 , 
		w_39886 , w_39887 , w_39888 , w_39889 , w_39890 , w_39891 , w_39892 , w_39893 , w_39894 , w_39895 , 
		w_39896 , w_39897 , w_39898 , w_39899 , w_39900 , w_39901 , w_39902 , w_39903 , w_39904 , w_39905 , 
		w_39906 , w_39907 , w_39908 , w_39909 , w_39910 , w_39911 , w_39912 , w_39913 , w_39914 , w_39915 , 
		w_39916 , w_39917 , w_39918 , w_39919 , w_39920 , w_39921 , w_39922 , w_39923 , w_39924 , w_39925 , 
		w_39926 , w_39927 , w_39928 , w_39929 , w_39930 , w_39931 , w_39932 , w_39933 , w_39934 , w_39935 , 
		w_39936 , w_39937 , w_39938 , w_39939 , w_39940 , w_39941 , w_39942 , w_39943 , w_39944 , w_39945 , 
		w_39946 , w_39947 , w_39948 , w_39949 , w_39950 , w_39951 , w_39952 , w_39953 , w_39954 , w_39955 , 
		w_39956 , w_39957 , w_39958 , w_39959 , w_39960 , w_39961 , w_39962 , w_39963 , w_39964 , w_39965 , 
		w_39966 , w_39967 , w_39968 , w_39969 , w_39970 , w_39971 , w_39972 , w_39973 , w_39974 , w_39975 , 
		w_39976 , w_39977 , w_39978 , w_39979 , w_39980 , w_39981 , w_39982 , w_39983 , w_39984 , w_39985 , 
		w_39986 , w_39987 , w_39988 , w_39989 , w_39990 , w_39991 , w_39992 , w_39993 , w_39994 , w_39995 , 
		w_39996 , w_39997 , w_39998 , w_39999 , w_40000 , w_40001 , w_40002 , w_40003 , w_40004 , w_40005 , 
		w_40006 , w_40007 , w_40008 , w_40009 , w_40010 , w_40011 , w_40012 , w_40013 , w_40014 , w_40015 , 
		w_40016 , w_40017 , w_40018 , w_40019 , w_40020 , w_40021 , w_40022 , w_40023 , w_40024 , w_40025 , 
		w_40026 , w_40027 , w_40028 , w_40029 , w_40030 , w_40031 , w_40032 , w_40033 , w_40034 , w_40035 , 
		w_40036 , w_40037 , w_40038 , w_40039 , w_40040 , w_40041 , w_40042 , w_40043 , w_40044 , w_40045 , 
		w_40046 , w_40047 , w_40048 , w_40049 , w_40050 , w_40051 , w_40052 , w_40053 , w_40054 , w_40055 , 
		w_40056 , w_40057 , w_40058 , w_40059 , w_40060 , w_40061 , w_40062 , w_40063 , w_40064 , w_40065 , 
		w_40066 , w_40067 , w_40068 , w_40069 , w_40070 , w_40071 , w_40072 , w_40073 , w_40074 , w_40075 , 
		w_40076 , w_40077 , w_40078 , w_40079 , w_40080 , w_40081 , w_40082 , w_40083 , w_40084 , w_40085 , 
		w_40086 , w_40087 , w_40088 , w_40089 , w_40090 , w_40091 , w_40092 , w_40093 , w_40094 , w_40095 , 
		w_40096 , w_40097 , w_40098 , w_40099 , w_40100 , w_40101 , w_40102 , w_40103 , w_40104 , w_40105 , 
		w_40106 , w_40107 , w_40108 , w_40109 , w_40110 , w_40111 , w_40112 , w_40113 , w_40114 , w_40115 , 
		w_40116 , w_40117 , w_40118 , w_40119 , w_40120 , w_40121 , w_40122 , w_40123 , w_40124 , w_40125 , 
		w_40126 , w_40127 , w_40128 , w_40129 , w_40130 , w_40131 , w_40132 , w_40133 , w_40134 , w_40135 , 
		w_40136 , w_40137 , w_40138 , w_40139 , w_40140 , w_40141 , w_40142 , w_40143 , w_40144 , w_40145 , 
		w_40146 , w_40147 , w_40148 , w_40149 , w_40150 , w_40151 , w_40152 , w_40153 , w_40154 , w_40155 , 
		w_40156 , w_40157 , w_40158 , w_40159 , w_40160 , w_40161 , w_40162 , w_40163 , w_40164 , w_40165 , 
		w_40166 , w_40167 , w_40168 , w_40169 , w_40170 , w_40171 , w_40172 , w_40173 , w_40174 , w_40175 , 
		w_40176 , w_40177 , w_40178 , w_40179 , w_40180 , w_40181 , w_40182 , w_40183 , w_40184 , w_40185 , 
		w_40186 , w_40187 , w_40188 , w_40189 , w_40190 , w_40191 , w_40192 , w_40193 , w_40194 , w_40195 , 
		w_40196 , w_40197 , w_40198 , w_40199 , w_40200 , w_40201 , w_40202 , w_40203 , w_40204 , w_40205 , 
		w_40206 , w_40207 , w_40208 , w_40209 , w_40210 , w_40211 , w_40212 , w_40213 , w_40214 , w_40215 , 
		w_40216 , w_40217 , w_40218 , w_40219 , w_40220 , w_40221 , w_40222 , w_40223 , w_40224 , w_40225 , 
		w_40226 , w_40227 , w_40228 , w_40229 , w_40230 , w_40231 , w_40232 , w_40233 , w_40234 , w_40235 , 
		w_40236 , w_40237 , w_40238 , w_40239 , w_40240 , w_40241 , w_40242 , w_40243 , w_40244 , w_40245 , 
		w_40246 , w_40247 , w_40248 , w_40249 , w_40250 , w_40251 , w_40252 , w_40253 , w_40254 , w_40255 , 
		w_40256 , w_40257 , w_40258 , w_40259 , w_40260 , w_40261 , w_40262 , w_40263 , w_40264 , w_40265 , 
		w_40266 , w_40267 , w_40268 , w_40269 , w_40270 , w_40271 , w_40272 , w_40273 , w_40274 , w_40275 , 
		w_40276 , w_40277 , w_40278 , w_40279 , w_40280 , w_40281 , w_40282 , w_40283 , w_40284 , w_40285 , 
		w_40286 , w_40287 , w_40288 , w_40289 , w_40290 , w_40291 , w_40292 , w_40293 , w_40294 , w_40295 , 
		w_40296 , w_40297 , w_40298 , w_40299 , w_40300 , w_40301 , w_40302 , w_40303 , w_40304 , w_40305 , 
		w_40306 , w_40307 , w_40308 , w_40309 , w_40310 , w_40311 , w_40312 , w_40313 , w_40314 , w_40315 , 
		w_40316 , w_40317 , w_40318 , w_40319 , w_40320 , w_40321 , w_40322 , w_40323 , w_40324 , w_40325 , 
		w_40326 , w_40327 , w_40328 , w_40329 , w_40330 , w_40331 , w_40332 , w_40333 , w_40334 , w_40335 , 
		w_40336 , w_40337 , w_40338 , w_40339 , w_40340 , w_40341 , w_40342 , w_40343 , w_40344 , w_40345 , 
		w_40346 , w_40347 , w_40348 , w_40349 , w_40350 , w_40351 , w_40352 , w_40353 , w_40354 , w_40355 , 
		w_40356 , w_40357 , w_40358 , w_40359 , w_40360 , w_40361 , w_40362 , w_40363 , w_40364 , w_40365 , 
		w_40366 , w_40367 , w_40368 , w_40369 , w_40370 , w_40371 , w_40372 , w_40373 , w_40374 , w_40375 , 
		w_40376 , w_40377 , w_40378 , w_40379 , w_40380 , w_40381 , w_40382 , w_40383 , w_40384 , w_40385 , 
		w_40386 , w_40387 , w_40388 , w_40389 , w_40390 , w_40391 , w_40392 , w_40393 , w_40394 , w_40395 , 
		w_40396 , w_40397 , w_40398 , w_40399 , w_40400 , w_40401 , w_40402 , w_40403 , w_40404 , w_40405 , 
		w_40406 , w_40407 , w_40408 , w_40409 , w_40410 , w_40411 , w_40412 , w_40413 , w_40414 , w_40415 , 
		w_40416 , w_40417 , w_40418 , w_40419 , w_40420 , w_40421 , w_40422 , w_40423 , w_40424 , w_40425 , 
		w_40426 , w_40427 , w_40428 , w_40429 , w_40430 , w_40431 , w_40432 , w_40433 , w_40434 , w_40435 , 
		w_40436 , w_40437 , w_40438 , w_40439 , w_40440 , w_40441 , w_40442 , w_40443 , w_40444 , w_40445 , 
		w_40446 , w_40447 , w_40448 , w_40449 , w_40450 , w_40451 , w_40452 , w_40453 , w_40454 , w_40455 , 
		w_40456 , w_40457 , w_40458 , w_40459 , w_40460 , w_40461 , w_40462 , w_40463 , w_40464 , w_40465 , 
		w_40466 , w_40467 , w_40468 , w_40469 , w_40470 , w_40471 , w_40472 , w_40473 , w_40474 , w_40475 , 
		w_40476 , w_40477 , w_40478 , w_40479 , w_40480 , w_40481 , w_40482 , w_40483 , w_40484 , w_40485 , 
		w_40486 , w_40487 , w_40488 , w_40489 , w_40490 , w_40491 , w_40492 , w_40493 , w_40494 , w_40495 , 
		w_40496 , w_40497 , w_40498 , w_40499 , w_40500 , w_40501 , w_40502 , w_40503 , w_40504 , w_40505 , 
		w_40506 , w_40507 , w_40508 , w_40509 , w_40510 , w_40511 , w_40512 , w_40513 , w_40514 , w_40515 , 
		w_40516 , w_40517 , w_40518 , w_40519 , w_40520 , w_40521 , w_40522 , w_40523 , w_40524 , w_40525 , 
		w_40526 , w_40527 , w_40528 , w_40529 , w_40530 , w_40531 , w_40532 , w_40533 , w_40534 , w_40535 , 
		w_40536 , w_40537 , w_40538 , w_40539 , w_40540 , w_40541 , w_40542 , w_40543 , w_40544 , w_40545 , 
		w_40546 , w_40547 , w_40548 , w_40549 , w_40550 , w_40551 , w_40552 , w_40553 , w_40554 , w_40555 , 
		w_40556 , w_40557 , w_40558 , w_40559 , w_40560 , w_40561 , w_40562 , w_40563 , w_40564 , w_40565 , 
		w_40566 , w_40567 , w_40568 , w_40569 , w_40570 , w_40571 , w_40572 , w_40573 , w_40574 , w_40575 , 
		w_40576 , w_40577 , w_40578 , w_40579 , w_40580 , w_40581 , w_40582 , w_40583 , w_40584 , w_40585 , 
		w_40586 , w_40587 , w_40588 , w_40589 , w_40590 , w_40591 , w_40592 , w_40593 , w_40594 , w_40595 , 
		w_40596 , w_40597 , w_40598 , w_40599 , w_40600 , w_40601 , w_40602 , w_40603 , w_40604 , w_40605 , 
		w_40606 , w_40607 , w_40608 , w_40609 , w_40610 , w_40611 , w_40612 , w_40613 , w_40614 , w_40615 , 
		w_40616 , w_40617 , w_40618 , w_40619 , w_40620 , w_40621 , w_40622 , w_40623 , w_40624 , w_40625 , 
		w_40626 , w_40627 , w_40628 , w_40629 , w_40630 , w_40631 , w_40632 , w_40633 , w_40634 , w_40635 , 
		w_40636 , w_40637 , w_40638 , w_40639 , w_40640 , w_40641 , w_40642 , w_40643 , w_40644 , w_40645 , 
		w_40646 , w_40647 , w_40648 , w_40649 , w_40650 , w_40651 , w_40652 , w_40653 , w_40654 , w_40655 , 
		w_40656 , w_40657 , w_40658 , w_40659 , w_40660 , w_40661 , w_40662 , w_40663 , w_40664 , w_40665 , 
		w_40666 , w_40667 , w_40668 , w_40669 , w_40670 , w_40671 , w_40672 , w_40673 , w_40674 , w_40675 , 
		w_40676 , w_40677 , w_40678 , w_40679 , w_40680 , w_40681 , w_40682 , w_40683 , w_40684 , w_40685 , 
		w_40686 , w_40687 , w_40688 , w_40689 , w_40690 , w_40691 , w_40692 , w_40693 , w_40694 , w_40695 , 
		w_40696 , w_40697 , w_40698 , w_40699 , w_40700 , w_40701 , w_40702 , w_40703 , w_40704 , w_40705 , 
		w_40706 , w_40707 , w_40708 , w_40709 , w_40710 , w_40711 , w_40712 , w_40713 , w_40714 , w_40715 , 
		w_40716 , w_40717 , w_40718 , w_40719 , w_40720 , w_40721 , w_40722 , w_40723 , w_40724 , w_40725 , 
		w_40726 , w_40727 , w_40728 , w_40729 , w_40730 , w_40731 , w_40732 , w_40733 , w_40734 , w_40735 , 
		w_40736 , w_40737 , w_40738 , w_40739 , w_40740 , w_40741 , w_40742 , w_40743 , w_40744 , w_40745 , 
		w_40746 , w_40747 , w_40748 , w_40749 , w_40750 , w_40751 , w_40752 , w_40753 , w_40754 , w_40755 , 
		w_40756 , w_40757 , w_40758 , w_40759 , w_40760 , w_40761 , w_40762 , w_40763 , w_40764 , w_40765 , 
		w_40766 , w_40767 , w_40768 , w_40769 , w_40770 , w_40771 , w_40772 , w_40773 , w_40774 , w_40775 , 
		w_40776 , w_40777 , w_40778 , w_40779 , w_40780 , w_40781 , w_40782 , w_40783 , w_40784 , w_40785 , 
		w_40786 , w_40787 , w_40788 , w_40789 , w_40790 , w_40791 , w_40792 , w_40793 , w_40794 , w_40795 , 
		w_40796 , w_40797 , w_40798 , w_40799 , w_40800 , w_40801 , w_40802 , w_40803 , w_40804 , w_40805 , 
		w_40806 , w_40807 , w_40808 , w_40809 , w_40810 , w_40811 , w_40812 , w_40813 , w_40814 , w_40815 , 
		w_40816 , w_40817 , w_40818 , w_40819 , w_40820 , w_40821 , w_40822 , w_40823 , w_40824 , w_40825 , 
		w_40826 , w_40827 , w_40828 , w_40829 , w_40830 , w_40831 , w_40832 , w_40833 , w_40834 , w_40835 , 
		w_40836 , w_40837 , w_40838 , w_40839 , w_40840 , w_40841 , w_40842 , w_40843 , w_40844 , w_40845 , 
		w_40846 , w_40847 , w_40848 , w_40849 , w_40850 , w_40851 , w_40852 , w_40853 , w_40854 , w_40855 , 
		w_40856 , w_40857 , w_40858 , w_40859 , w_40860 , w_40861 , w_40862 , w_40863 , w_40864 , w_40865 , 
		w_40866 , w_40867 , w_40868 , w_40869 , w_40870 , w_40871 , w_40872 , w_40873 , w_40874 , w_40875 , 
		w_40876 , w_40877 , w_40878 , w_40879 , w_40880 , w_40881 , w_40882 , w_40883 , w_40884 , w_40885 , 
		w_40886 , w_40887 , w_40888 , w_40889 , w_40890 , w_40891 , w_40892 , w_40893 , w_40894 , w_40895 , 
		w_40896 , w_40897 , w_40898 , w_40899 , w_40900 , w_40901 , w_40902 , w_40903 , w_40904 , w_40905 , 
		w_40906 , w_40907 , w_40908 , w_40909 , w_40910 , w_40911 , w_40912 , w_40913 , w_40914 , w_40915 , 
		w_40916 , w_40917 , w_40918 , w_40919 , w_40920 , w_40921 , w_40922 , w_40923 , w_40924 , w_40925 , 
		w_40926 , w_40927 , w_40928 , w_40929 , w_40930 , w_40931 , w_40932 , w_40933 , w_40934 , w_40935 , 
		w_40936 , w_40937 , w_40938 , w_40939 , w_40940 , w_40941 , w_40942 , w_40943 , w_40944 , w_40945 , 
		w_40946 , w_40947 , w_40948 , w_40949 , w_40950 , w_40951 , w_40952 , w_40953 , w_40954 , w_40955 , 
		w_40956 , w_40957 , w_40958 , w_40959 , w_40960 , w_40961 , w_40962 , w_40963 , w_40964 , w_40965 , 
		w_40966 , w_40967 , w_40968 , w_40969 , w_40970 , w_40971 , w_40972 , w_40973 , w_40974 , w_40975 , 
		w_40976 , w_40977 , w_40978 , w_40979 , w_40980 , w_40981 , w_40982 , w_40983 , w_40984 , w_40985 , 
		w_40986 , w_40987 , w_40988 , w_40989 , w_40990 , w_40991 , w_40992 , w_40993 , w_40994 , w_40995 , 
		w_40996 , w_40997 , w_40998 , w_40999 , w_41000 , w_41001 , w_41002 , w_41003 , w_41004 , w_41005 , 
		w_41006 , w_41007 , w_41008 , w_41009 , w_41010 , w_41011 , w_41012 , w_41013 , w_41014 , w_41015 , 
		w_41016 , w_41017 , w_41018 , w_41019 , w_41020 , w_41021 , w_41022 , w_41023 , w_41024 , w_41025 , 
		w_41026 , w_41027 , w_41028 , w_41029 , w_41030 , w_41031 , w_41032 , w_41033 , w_41034 , w_41035 , 
		w_41036 , w_41037 , w_41038 , w_41039 , w_41040 , w_41041 , w_41042 , w_41043 , w_41044 , w_41045 , 
		w_41046 , w_41047 , w_41048 , w_41049 , w_41050 , w_41051 , w_41052 , w_41053 , w_41054 , w_41055 , 
		w_41056 , w_41057 , w_41058 , w_41059 , w_41060 , w_41061 , w_41062 , w_41063 , w_41064 , w_41065 , 
		w_41066 , w_41067 , w_41068 , w_41069 , w_41070 , w_41071 , w_41072 , w_41073 , w_41074 , w_41075 , 
		w_41076 , w_41077 , w_41078 , w_41079 , w_41080 , w_41081 , w_41082 , w_41083 , w_41084 , w_41085 , 
		w_41086 , w_41087 , w_41088 , w_41089 , w_41090 , w_41091 , w_41092 , w_41093 , w_41094 , w_41095 , 
		w_41096 , w_41097 , w_41098 , w_41099 , w_41100 , w_41101 , w_41102 , w_41103 , w_41104 , w_41105 , 
		w_41106 , w_41107 , w_41108 , w_41109 , w_41110 , w_41111 , w_41112 , w_41113 , w_41114 , w_41115 , 
		w_41116 , w_41117 , w_41118 , w_41119 , w_41120 , w_41121 , w_41122 , w_41123 , w_41124 , w_41125 , 
		w_41126 , w_41127 , w_41128 , w_41129 , w_41130 , w_41131 , w_41132 , w_41133 , w_41134 , w_41135 , 
		w_41136 , w_41137 , w_41138 , w_41139 , w_41140 , w_41141 , w_41142 , w_41143 , w_41144 , w_41145 , 
		w_41146 , w_41147 , w_41148 , w_41149 , w_41150 , w_41151 , w_41152 , w_41153 , w_41154 , w_41155 , 
		w_41156 , w_41157 , w_41158 , w_41159 , w_41160 , w_41161 , w_41162 , w_41163 , w_41164 , w_41165 , 
		w_41166 , w_41167 , w_41168 , w_41169 , w_41170 , w_41171 , w_41172 , w_41173 , w_41174 , w_41175 , 
		w_41176 , w_41177 , w_41178 , w_41179 , w_41180 , w_41181 , w_41182 , w_41183 , w_41184 , w_41185 , 
		w_41186 , w_41187 , w_41188 , w_41189 , w_41190 , w_41191 , w_41192 , w_41193 , w_41194 , w_41195 , 
		w_41196 , w_41197 , w_41198 , w_41199 , w_41200 , w_41201 , w_41202 , w_41203 , w_41204 , w_41205 , 
		w_41206 , w_41207 , w_41208 , w_41209 , w_41210 , w_41211 , w_41212 , w_41213 , w_41214 , w_41215 , 
		w_41216 , w_41217 , w_41218 , w_41219 , w_41220 , w_41221 , w_41222 , w_41223 , w_41224 , w_41225 , 
		w_41226 , w_41227 , w_41228 , w_41229 , w_41230 , w_41231 , w_41232 , w_41233 , w_41234 , w_41235 , 
		w_41236 , w_41237 , w_41238 , w_41239 , w_41240 , w_41241 , w_41242 , w_41243 , w_41244 , w_41245 , 
		w_41246 , w_41247 , w_41248 , w_41249 , w_41250 , w_41251 , w_41252 , w_41253 , w_41254 , w_41255 , 
		w_41256 , w_41257 , w_41258 , w_41259 , w_41260 , w_41261 , w_41262 , w_41263 , w_41264 , w_41265 , 
		w_41266 , w_41267 , w_41268 , w_41269 , w_41270 , w_41271 , w_41272 , w_41273 , w_41274 , w_41275 , 
		w_41276 , w_41277 , w_41278 , w_41279 , w_41280 , w_41281 , w_41282 , w_41283 , w_41284 , w_41285 , 
		w_41286 , w_41287 , w_41288 , w_41289 , w_41290 , w_41291 , w_41292 , w_41293 , w_41294 , w_41295 , 
		w_41296 , w_41297 , w_41298 , w_41299 , w_41300 , w_41301 , w_41302 , w_41303 , w_41304 , w_41305 , 
		w_41306 , w_41307 , w_41308 , w_41309 , w_41310 , w_41311 , w_41312 , w_41313 , w_41314 , w_41315 , 
		w_41316 , w_41317 , w_41318 , w_41319 , w_41320 , w_41321 , w_41322 , w_41323 , w_41324 , w_41325 , 
		w_41326 , w_41327 , w_41328 , w_41329 , w_41330 , w_41331 , w_41332 , w_41333 , w_41334 , w_41335 , 
		w_41336 , w_41337 , w_41338 , w_41339 , w_41340 , w_41341 , w_41342 , w_41343 , w_41344 , w_41345 , 
		w_41346 , w_41347 , w_41348 , w_41349 , w_41350 , w_41351 , w_41352 , w_41353 , w_41354 , w_41355 , 
		w_41356 , w_41357 , w_41358 , w_41359 , w_41360 , w_41361 , w_41362 , w_41363 , w_41364 , w_41365 , 
		w_41366 , w_41367 , w_41368 , w_41369 , w_41370 , w_41371 , w_41372 , w_41373 , w_41374 , w_41375 , 
		w_41376 , w_41377 , w_41378 , w_41379 , w_41380 , w_41381 , w_41382 , w_41383 , w_41384 , w_41385 , 
		w_41386 , w_41387 , w_41388 , w_41389 , w_41390 , w_41391 , w_41392 , w_41393 , w_41394 , w_41395 , 
		w_41396 , w_41397 , w_41398 , w_41399 , w_41400 , w_41401 , w_41402 , w_41403 , w_41404 , w_41405 , 
		w_41406 , w_41407 , w_41408 , w_41409 , w_41410 , w_41411 , w_41412 , w_41413 , w_41414 , w_41415 , 
		w_41416 , w_41417 , w_41418 , w_41419 , w_41420 , w_41421 , w_41422 , w_41423 , w_41424 , w_41425 , 
		w_41426 , w_41427 , w_41428 , w_41429 , w_41430 , w_41431 , w_41432 , w_41433 , w_41434 , w_41435 , 
		w_41436 , w_41437 , w_41438 , w_41439 , w_41440 , w_41441 , w_41442 , w_41443 , w_41444 , w_41445 , 
		w_41446 , w_41447 , w_41448 , w_41449 , w_41450 , w_41451 , w_41452 , w_41453 , w_41454 , w_41455 , 
		w_41456 , w_41457 , w_41458 , w_41459 , w_41460 , w_41461 , w_41462 , w_41463 , w_41464 , w_41465 , 
		w_41466 , w_41467 , w_41468 , w_41469 , w_41470 , w_41471 , w_41472 , w_41473 , w_41474 , w_41475 , 
		w_41476 , w_41477 , w_41478 , w_41479 , w_41480 , w_41481 , w_41482 , w_41483 , w_41484 , w_41485 , 
		w_41486 , w_41487 , w_41488 , w_41489 , w_41490 , w_41491 , w_41492 , w_41493 , w_41494 , w_41495 , 
		w_41496 , w_41497 , w_41498 , w_41499 , w_41500 , w_41501 , w_41502 , w_41503 , w_41504 , w_41505 , 
		w_41506 , w_41507 , w_41508 , w_41509 , w_41510 , w_41511 , w_41512 , w_41513 , w_41514 , w_41515 , 
		w_41516 , w_41517 , w_41518 , w_41519 , w_41520 , w_41521 , w_41522 , w_41523 , w_41524 , w_41525 , 
		w_41526 , w_41527 , w_41528 , w_41529 , w_41530 , w_41531 , w_41532 , w_41533 , w_41534 , w_41535 , 
		w_41536 , w_41537 , w_41538 , w_41539 , w_41540 , w_41541 , w_41542 , w_41543 , w_41544 , w_41545 , 
		w_41546 , w_41547 , w_41548 , w_41549 , w_41550 , w_41551 , w_41552 , w_41553 , w_41554 , w_41555 , 
		w_41556 , w_41557 , w_41558 , w_41559 , w_41560 , w_41561 , w_41562 , w_41563 , w_41564 , w_41565 , 
		w_41566 , w_41567 , w_41568 , w_41569 , w_41570 , w_41571 , w_41572 , w_41573 , w_41574 , w_41575 , 
		w_41576 , w_41577 , w_41578 , w_41579 , w_41580 , w_41581 , w_41582 , w_41583 , w_41584 , w_41585 , 
		w_41586 , w_41587 , w_41588 , w_41589 , w_41590 , w_41591 , w_41592 , w_41593 , w_41594 , w_41595 , 
		w_41596 , w_41597 , w_41598 , w_41599 , w_41600 , w_41601 , w_41602 , w_41603 , w_41604 , w_41605 , 
		w_41606 , w_41607 , w_41608 , w_41609 , w_41610 , w_41611 , w_41612 , w_41613 , w_41614 , w_41615 , 
		w_41616 , w_41617 , w_41618 , w_41619 , w_41620 , w_41621 , w_41622 , w_41623 , w_41624 , w_41625 , 
		w_41626 , w_41627 , w_41628 , w_41629 , w_41630 , w_41631 , w_41632 , w_41633 , w_41634 , w_41635 , 
		w_41636 , w_41637 , w_41638 , w_41639 , w_41640 , w_41641 , w_41642 , w_41643 , w_41644 , w_41645 , 
		w_41646 , w_41647 , w_41648 , w_41649 , w_41650 , w_41651 , w_41652 , w_41653 , w_41654 , w_41655 , 
		w_41656 , w_41657 , w_41658 , w_41659 , w_41660 , w_41661 , w_41662 , w_41663 , w_41664 , w_41665 , 
		w_41666 , w_41667 , w_41668 , w_41669 , w_41670 , w_41671 , w_41672 , w_41673 , w_41674 , w_41675 , 
		w_41676 , w_41677 , w_41678 , w_41679 , w_41680 , w_41681 , w_41682 , w_41683 , w_41684 , w_41685 , 
		w_41686 , w_41687 , w_41688 , w_41689 , w_41690 , w_41691 , w_41692 , w_41693 , w_41694 , w_41695 , 
		w_41696 , w_41697 , w_41698 , w_41699 , w_41700 , w_41701 , w_41702 , w_41703 , w_41704 , w_41705 , 
		w_41706 , w_41707 , w_41708 , w_41709 , w_41710 , w_41711 , w_41712 , w_41713 , w_41714 , w_41715 , 
		w_41716 , w_41717 , w_41718 , w_41719 , w_41720 , w_41721 , w_41722 , w_41723 , w_41724 , w_41725 , 
		w_41726 , w_41727 , w_41728 , w_41729 , w_41730 , w_41731 , w_41732 , w_41733 , w_41734 , w_41735 , 
		w_41736 , w_41737 , w_41738 , w_41739 , w_41740 , w_41741 , w_41742 , w_41743 , w_41744 , w_41745 , 
		w_41746 , w_41747 , w_41748 , w_41749 , w_41750 , w_41751 , w_41752 , w_41753 , w_41754 , w_41755 , 
		w_41756 , w_41757 , w_41758 , w_41759 , w_41760 , w_41761 , w_41762 , w_41763 , w_41764 , w_41765 , 
		w_41766 , w_41767 , w_41768 , w_41769 , w_41770 , w_41771 , w_41772 , w_41773 , w_41774 , w_41775 , 
		w_41776 , w_41777 , w_41778 , w_41779 , w_41780 , w_41781 , w_41782 , w_41783 , w_41784 , w_41785 , 
		w_41786 , w_41787 , w_41788 , w_41789 , w_41790 , w_41791 , w_41792 , w_41793 , w_41794 , w_41795 , 
		w_41796 , w_41797 , w_41798 , w_41799 , w_41800 , w_41801 , w_41802 , w_41803 , w_41804 , w_41805 , 
		w_41806 , w_41807 , w_41808 , w_41809 , w_41810 , w_41811 , w_41812 , w_41813 , w_41814 , w_41815 , 
		w_41816 , w_41817 , w_41818 , w_41819 , w_41820 , w_41821 , w_41822 , w_41823 , w_41824 , w_41825 , 
		w_41826 , w_41827 , w_41828 , w_41829 , w_41830 , w_41831 , w_41832 , w_41833 , w_41834 , w_41835 , 
		w_41836 , w_41837 , w_41838 , w_41839 , w_41840 , w_41841 , w_41842 , w_41843 , w_41844 , w_41845 , 
		w_41846 , w_41847 , w_41848 , w_41849 , w_41850 , w_41851 , w_41852 , w_41853 , w_41854 , w_41855 , 
		w_41856 , w_41857 , w_41858 , w_41859 , w_41860 , w_41861 , w_41862 , w_41863 , w_41864 , w_41865 , 
		w_41866 , w_41867 , w_41868 , w_41869 , w_41870 , w_41871 , w_41872 , w_41873 , w_41874 , w_41875 , 
		w_41876 , w_41877 , w_41878 , w_41879 , w_41880 , w_41881 , w_41882 , w_41883 , w_41884 , w_41885 , 
		w_41886 , w_41887 , w_41888 , w_41889 , w_41890 , w_41891 , w_41892 , w_41893 , w_41894 , w_41895 , 
		w_41896 , w_41897 , w_41898 , w_41899 , w_41900 , w_41901 , w_41902 , w_41903 , w_41904 , w_41905 , 
		w_41906 , w_41907 , w_41908 , w_41909 , w_41910 , w_41911 , w_41912 , w_41913 , w_41914 , w_41915 , 
		w_41916 , w_41917 , w_41918 , w_41919 , w_41920 , w_41921 , w_41922 , w_41923 , w_41924 , w_41925 , 
		w_41926 , w_41927 , w_41928 , w_41929 , w_41930 , w_41931 , w_41932 , w_41933 , w_41934 , w_41935 , 
		w_41936 , w_41937 , w_41938 , w_41939 , w_41940 , w_41941 , w_41942 , w_41943 , w_41944 , w_41945 , 
		w_41946 , w_41947 , w_41948 , w_41949 , w_41950 , w_41951 , w_41952 , w_41953 , w_41954 , w_41955 , 
		w_41956 , w_41957 , w_41958 , w_41959 , w_41960 , w_41961 , w_41962 , w_41963 , w_41964 , w_41965 , 
		w_41966 , w_41967 , w_41968 , w_41969 , w_41970 , w_41971 , w_41972 , w_41973 , w_41974 , w_41975 , 
		w_41976 , w_41977 , w_41978 , w_41979 , w_41980 , w_41981 , w_41982 , w_41983 , w_41984 , w_41985 , 
		w_41986 , w_41987 , w_41988 , w_41989 , w_41990 , w_41991 , w_41992 , w_41993 , w_41994 , w_41995 , 
		w_41996 , w_41997 , w_41998 , w_41999 , w_42000 , w_42001 , w_42002 , w_42003 , w_42004 , w_42005 , 
		w_42006 , w_42007 , w_42008 , w_42009 , w_42010 , w_42011 , w_42012 , w_42013 , w_42014 , w_42015 , 
		w_42016 , w_42017 , w_42018 , w_42019 , w_42020 , w_42021 , w_42022 , w_42023 , w_42024 , w_42025 , 
		w_42026 , w_42027 , w_42028 , w_42029 , w_42030 , w_42031 , w_42032 , w_42033 , w_42034 , w_42035 , 
		w_42036 , w_42037 , w_42038 , w_42039 , w_42040 , w_42041 , w_42042 , w_42043 , w_42044 , w_42045 , 
		w_42046 , w_42047 , w_42048 , w_42049 , w_42050 , w_42051 , w_42052 , w_42053 , w_42054 , w_42055 , 
		w_42056 , w_42057 , w_42058 , w_42059 , w_42060 , w_42061 , w_42062 , w_42063 , w_42064 , w_42065 , 
		w_42066 , w_42067 , w_42068 , w_42069 , w_42070 , w_42071 , w_42072 , w_42073 , w_42074 , w_42075 , 
		w_42076 , w_42077 , w_42078 , w_42079 , w_42080 , w_42081 , w_42082 , w_42083 , w_42084 , w_42085 , 
		w_42086 , w_42087 , w_42088 , w_42089 , w_42090 , w_42091 , w_42092 , w_42093 , w_42094 , w_42095 , 
		w_42096 , w_42097 , w_42098 , w_42099 , w_42100 , w_42101 , w_42102 , w_42103 , w_42104 , w_42105 , 
		w_42106 , w_42107 , w_42108 , w_42109 , w_42110 , w_42111 , w_42112 , w_42113 , w_42114 , w_42115 , 
		w_42116 , w_42117 , w_42118 , w_42119 , w_42120 , w_42121 , w_42122 , w_42123 , w_42124 , w_42125 , 
		w_42126 , w_42127 , w_42128 , w_42129 , w_42130 , w_42131 , w_42132 , w_42133 , w_42134 , w_42135 , 
		w_42136 , w_42137 , w_42138 , w_42139 , w_42140 , w_42141 , w_42142 , w_42143 , w_42144 , w_42145 , 
		w_42146 , w_42147 , w_42148 , w_42149 , w_42150 , w_42151 , w_42152 , w_42153 , w_42154 , w_42155 , 
		w_42156 , w_42157 , w_42158 , w_42159 , w_42160 , w_42161 , w_42162 , w_42163 , w_42164 , w_42165 , 
		w_42166 , w_42167 , w_42168 , w_42169 , w_42170 , w_42171 , w_42172 , w_42173 , w_42174 , w_42175 , 
		w_42176 , w_42177 , w_42178 , w_42179 , w_42180 , w_42181 , w_42182 , w_42183 , w_42184 , w_42185 , 
		w_42186 , w_42187 , w_42188 , w_42189 , w_42190 , w_42191 , w_42192 , w_42193 , w_42194 , w_42195 , 
		w_42196 , w_42197 , w_42198 , w_42199 , w_42200 , w_42201 , w_42202 , w_42203 , w_42204 , w_42205 , 
		w_42206 , w_42207 , w_42208 , w_42209 , w_42210 , w_42211 , w_42212 , w_42213 , w_42214 , w_42215 , 
		w_42216 , w_42217 , w_42218 , w_42219 , w_42220 , w_42221 , w_42222 , w_42223 , w_42224 , w_42225 , 
		w_42226 , w_42227 , w_42228 , w_42229 , w_42230 , w_42231 , w_42232 , w_42233 , w_42234 , w_42235 , 
		w_42236 , w_42237 , w_42238 , w_42239 , w_42240 , w_42241 , w_42242 , w_42243 , w_42244 , w_42245 , 
		w_42246 , w_42247 , w_42248 , w_42249 , w_42250 , w_42251 , w_42252 , w_42253 , w_42254 , w_42255 , 
		w_42256 , w_42257 , w_42258 , w_42259 , w_42260 , w_42261 , w_42262 , w_42263 , w_42264 , w_42265 , 
		w_42266 , w_42267 , w_42268 , w_42269 , w_42270 , w_42271 , w_42272 , w_42273 , w_42274 , w_42275 , 
		w_42276 , w_42277 , w_42278 , w_42279 , w_42280 , w_42281 , w_42282 , w_42283 , w_42284 , w_42285 , 
		w_42286 , w_42287 , w_42288 , w_42289 , w_42290 , w_42291 , w_42292 , w_42293 , w_42294 , w_42295 , 
		w_42296 , w_42297 , w_42298 , w_42299 , w_42300 , w_42301 , w_42302 , w_42303 , w_42304 , w_42305 , 
		w_42306 , w_42307 , w_42308 , w_42309 , w_42310 , w_42311 , w_42312 , w_42313 , w_42314 , w_42315 , 
		w_42316 , w_42317 , w_42318 , w_42319 , w_42320 , w_42321 , w_42322 , w_42323 , w_42324 , w_42325 , 
		w_42326 , w_42327 , w_42328 , w_42329 , w_42330 , w_42331 , w_42332 , w_42333 , w_42334 , w_42335 , 
		w_42336 , w_42337 , w_42338 , w_42339 , w_42340 , w_42341 , w_42342 , w_42343 , w_42344 , w_42345 , 
		w_42346 , w_42347 , w_42348 , w_42349 , w_42350 , w_42351 , w_42352 , w_42353 , w_42354 , w_42355 , 
		w_42356 , w_42357 , w_42358 , w_42359 , w_42360 , w_42361 , w_42362 , w_42363 , w_42364 , w_42365 , 
		w_42366 , w_42367 , w_42368 , w_42369 , w_42370 , w_42371 , w_42372 , w_42373 , w_42374 , w_42375 , 
		w_42376 , w_42377 , w_42378 , w_42379 , w_42380 , w_42381 , w_42382 , w_42383 , w_42384 , w_42385 , 
		w_42386 , w_42387 , w_42388 , w_42389 , w_42390 , w_42391 , w_42392 , w_42393 , w_42394 , w_42395 , 
		w_42396 , w_42397 , w_42398 , w_42399 , w_42400 , w_42401 , w_42402 , w_42403 , w_42404 , w_42405 , 
		w_42406 , w_42407 , w_42408 , w_42409 , w_42410 , w_42411 , w_42412 , w_42413 , w_42414 , w_42415 , 
		w_42416 , w_42417 , w_42418 , w_42419 , w_42420 , w_42421 , w_42422 , w_42423 , w_42424 , w_42425 , 
		w_42426 , w_42427 , w_42428 , w_42429 , w_42430 , w_42431 , w_42432 , w_42433 , w_42434 , w_42435 , 
		w_42436 , w_42437 , w_42438 , w_42439 , w_42440 , w_42441 , w_42442 , w_42443 , w_42444 , w_42445 , 
		w_42446 , w_42447 , w_42448 , w_42449 , w_42450 , w_42451 , w_42452 , w_42453 , w_42454 , w_42455 , 
		w_42456 , w_42457 , w_42458 , w_42459 , w_42460 , w_42461 , w_42462 , w_42463 , w_42464 , w_42465 , 
		w_42466 , w_42467 , w_42468 , w_42469 , w_42470 , w_42471 , w_42472 , w_42473 , w_42474 , w_42475 , 
		w_42476 , w_42477 , w_42478 , w_42479 , w_42480 , w_42481 , w_42482 , w_42483 , w_42484 , w_42485 , 
		w_42486 , w_42487 , w_42488 , w_42489 , w_42490 , w_42491 , w_42492 , w_42493 , w_42494 , w_42495 , 
		w_42496 , w_42497 , w_42498 , w_42499 , w_42500 , w_42501 , w_42502 , w_42503 , w_42504 , w_42505 , 
		w_42506 , w_42507 , w_42508 , w_42509 , w_42510 , w_42511 , w_42512 , w_42513 , w_42514 , w_42515 , 
		w_42516 , w_42517 , w_42518 , w_42519 , w_42520 , w_42521 , w_42522 , w_42523 , w_42524 , w_42525 , 
		w_42526 , w_42527 , w_42528 , w_42529 , w_42530 , w_42531 , w_42532 , w_42533 , w_42534 , w_42535 , 
		w_42536 , w_42537 , w_42538 , w_42539 , w_42540 , w_42541 , w_42542 , w_42543 , w_42544 , w_42545 , 
		w_42546 , w_42547 , w_42548 , w_42549 , w_42550 , w_42551 , w_42552 , w_42553 , w_42554 , w_42555 , 
		w_42556 , w_42557 , w_42558 , w_42559 , w_42560 , w_42561 , w_42562 , w_42563 , w_42564 , w_42565 , 
		w_42566 , w_42567 , w_42568 , w_42569 , w_42570 , w_42571 , w_42572 , w_42573 , w_42574 , w_42575 , 
		w_42576 , w_42577 , w_42578 , w_42579 , w_42580 , w_42581 , w_42582 , w_42583 , w_42584 , w_42585 , 
		w_42586 , w_42587 , w_42588 , w_42589 , w_42590 , w_42591 , w_42592 , w_42593 , w_42594 , w_42595 , 
		w_42596 , w_42597 , w_42598 , w_42599 , w_42600 , w_42601 , w_42602 , w_42603 , w_42604 , w_42605 , 
		w_42606 , w_42607 , w_42608 , w_42609 , w_42610 , w_42611 , w_42612 , w_42613 , w_42614 , w_42615 , 
		w_42616 , w_42617 , w_42618 , w_42619 , w_42620 , w_42621 , w_42622 , w_42623 , w_42624 , w_42625 , 
		w_42626 , w_42627 , w_42628 , w_42629 , w_42630 , w_42631 , w_42632 , w_42633 , w_42634 , w_42635 , 
		w_42636 , w_42637 , w_42638 , w_42639 , w_42640 , w_42641 , w_42642 , w_42643 , w_42644 , w_42645 , 
		w_42646 , w_42647 , w_42648 , w_42649 , w_42650 , w_42651 , w_42652 , w_42653 , w_42654 , w_42655 , 
		w_42656 , w_42657 , w_42658 , w_42659 , w_42660 , w_42661 , w_42662 , w_42663 , w_42664 , w_42665 , 
		w_42666 , w_42667 , w_42668 , w_42669 , w_42670 , w_42671 , w_42672 , w_42673 , w_42674 , w_42675 , 
		w_42676 , w_42677 , w_42678 , w_42679 , w_42680 , w_42681 , w_42682 , w_42683 , w_42684 , w_42685 , 
		w_42686 , w_42687 , w_42688 , w_42689 , w_42690 , w_42691 , w_42692 , w_42693 , w_42694 , w_42695 , 
		w_42696 , w_42697 , w_42698 , w_42699 , w_42700 , w_42701 , w_42702 , w_42703 , w_42704 , w_42705 , 
		w_42706 , w_42707 , w_42708 , w_42709 , w_42710 , w_42711 , w_42712 , w_42713 , w_42714 , w_42715 , 
		w_42716 , w_42717 , w_42718 , w_42719 , w_42720 , w_42721 , w_42722 , w_42723 , w_42724 , w_42725 , 
		w_42726 , w_42727 , w_42728 , w_42729 , w_42730 , w_42731 , w_42732 , w_42733 , w_42734 , w_42735 , 
		w_42736 , w_42737 , w_42738 , w_42739 , w_42740 , w_42741 , w_42742 , w_42743 , w_42744 , w_42745 , 
		w_42746 , w_42747 , w_42748 , w_42749 , w_42750 , w_42751 , w_42752 , w_42753 , w_42754 , w_42755 , 
		w_42756 , w_42757 , w_42758 , w_42759 , w_42760 , w_42761 , w_42762 , w_42763 , w_42764 , w_42765 , 
		w_42766 , w_42767 , w_42768 , w_42769 , w_42770 , w_42771 , w_42772 , w_42773 , w_42774 , w_42775 , 
		w_42776 , w_42777 , w_42778 , w_42779 , w_42780 , w_42781 , w_42782 , w_42783 , w_42784 , w_42785 , 
		w_42786 , w_42787 , w_42788 , w_42789 , w_42790 , w_42791 , w_42792 , w_42793 , w_42794 , w_42795 , 
		w_42796 , w_42797 , w_42798 , w_42799 , w_42800 , w_42801 , w_42802 , w_42803 , w_42804 , w_42805 , 
		w_42806 , w_42807 , w_42808 , w_42809 , w_42810 , w_42811 , w_42812 , w_42813 , w_42814 , w_42815 , 
		w_42816 , w_42817 , w_42818 , w_42819 , w_42820 , w_42821 , w_42822 , w_42823 , w_42824 , w_42825 , 
		w_42826 , w_42827 , w_42828 , w_42829 , w_42830 , w_42831 , w_42832 , w_42833 , w_42834 , w_42835 , 
		w_42836 , w_42837 , w_42838 , w_42839 , w_42840 , w_42841 , w_42842 , w_42843 , w_42844 , w_42845 , 
		w_42846 , w_42847 , w_42848 , w_42849 , w_42850 , w_42851 , w_42852 , w_42853 , w_42854 , w_42855 , 
		w_42856 , w_42857 , w_42858 , w_42859 , w_42860 , w_42861 , w_42862 , w_42863 , w_42864 , w_42865 , 
		w_42866 , w_42867 , w_42868 , w_42869 , w_42870 , w_42871 , w_42872 , w_42873 , w_42874 , w_42875 , 
		w_42876 , w_42877 , w_42878 , w_42879 , w_42880 , w_42881 , w_42882 , w_42883 , w_42884 , w_42885 , 
		w_42886 , w_42887 , w_42888 , w_42889 , w_42890 , w_42891 , w_42892 , w_42893 , w_42894 , w_42895 , 
		w_42896 , w_42897 , w_42898 , w_42899 , w_42900 , w_42901 , w_42902 , w_42903 , w_42904 , w_42905 , 
		w_42906 , w_42907 , w_42908 , w_42909 , w_42910 , w_42911 , w_42912 , w_42913 , w_42914 , w_42915 , 
		w_42916 , w_42917 , w_42918 , w_42919 , w_42920 , w_42921 , w_42922 , w_42923 , w_42924 , w_42925 , 
		w_42926 , w_42927 , w_42928 , w_42929 , w_42930 , w_42931 , w_42932 , w_42933 , w_42934 , w_42935 , 
		w_42936 , w_42937 , w_42938 , w_42939 , w_42940 , w_42941 , w_42942 , w_42943 , w_42944 , w_42945 , 
		w_42946 , w_42947 , w_42948 , w_42949 , w_42950 , w_42951 , w_42952 , w_42953 , w_42954 , w_42955 , 
		w_42956 , w_42957 , w_42958 , w_42959 , w_42960 , w_42961 , w_42962 , w_42963 , w_42964 , w_42965 , 
		w_42966 , w_42967 , w_42968 , w_42969 , w_42970 , w_42971 , w_42972 , w_42973 , w_42974 , w_42975 , 
		w_42976 , w_42977 , w_42978 , w_42979 , w_42980 , w_42981 , w_42982 , w_42983 , w_42984 , w_42985 , 
		w_42986 , w_42987 , w_42988 , w_42989 , w_42990 , w_42991 , w_42992 , w_42993 , w_42994 , w_42995 , 
		w_42996 , w_42997 , w_42998 , w_42999 , w_43000 , w_43001 , w_43002 , w_43003 , w_43004 , w_43005 , 
		w_43006 , w_43007 , w_43008 , w_43009 , w_43010 , w_43011 , w_43012 , w_43013 , w_43014 , w_43015 , 
		w_43016 , w_43017 , w_43018 , w_43019 , w_43020 , w_43021 , w_43022 , w_43023 , w_43024 , w_43025 , 
		w_43026 , w_43027 , w_43028 , w_43029 , w_43030 , w_43031 , w_43032 , w_43033 , w_43034 , w_43035 , 
		w_43036 , w_43037 , w_43038 , w_43039 , w_43040 , w_43041 , w_43042 , w_43043 , w_43044 , w_43045 , 
		w_43046 , w_43047 , w_43048 , w_43049 , w_43050 , w_43051 , w_43052 , w_43053 , w_43054 , w_43055 , 
		w_43056 , w_43057 , w_43058 , w_43059 , w_43060 , w_43061 , w_43062 , w_43063 , w_43064 , w_43065 , 
		w_43066 , w_43067 , w_43068 , w_43069 , w_43070 , w_43071 , w_43072 , w_43073 , w_43074 , w_43075 , 
		w_43076 , w_43077 , w_43078 , w_43079 , w_43080 , w_43081 , w_43082 , w_43083 , w_43084 , w_43085 , 
		w_43086 , w_43087 , w_43088 , w_43089 , w_43090 , w_43091 , w_43092 , w_43093 , w_43094 , w_43095 , 
		w_43096 , w_43097 , w_43098 , w_43099 , w_43100 , w_43101 , w_43102 , w_43103 , w_43104 , w_43105 , 
		w_43106 , w_43107 , w_43108 , w_43109 , w_43110 , w_43111 , w_43112 , w_43113 , w_43114 , w_43115 , 
		w_43116 , w_43117 , w_43118 , w_43119 , w_43120 , w_43121 , w_43122 , w_43123 , w_43124 , w_43125 , 
		w_43126 , w_43127 , w_43128 , w_43129 , w_43130 , w_43131 , w_43132 , w_43133 , w_43134 , w_43135 , 
		w_43136 , w_43137 , w_43138 , w_43139 , w_43140 , w_43141 , w_43142 , w_43143 , w_43144 , w_43145 , 
		w_43146 , w_43147 , w_43148 , w_43149 , w_43150 , w_43151 , w_43152 , w_43153 , w_43154 , w_43155 , 
		w_43156 , w_43157 , w_43158 , w_43159 , w_43160 , w_43161 , w_43162 , w_43163 , w_43164 , w_43165 , 
		w_43166 , w_43167 , w_43168 , w_43169 , w_43170 , w_43171 , w_43172 , w_43173 , w_43174 , w_43175 , 
		w_43176 , w_43177 , w_43178 , w_43179 , w_43180 , w_43181 , w_43182 , w_43183 , w_43184 , w_43185 , 
		w_43186 , w_43187 , w_43188 , w_43189 , w_43190 , w_43191 , w_43192 , w_43193 , w_43194 , w_43195 , 
		w_43196 , w_43197 , w_43198 , w_43199 , w_43200 , w_43201 , w_43202 , w_43203 , w_43204 , w_43205 , 
		w_43206 , w_43207 , w_43208 , w_43209 , w_43210 , w_43211 , w_43212 , w_43213 , w_43214 , w_43215 , 
		w_43216 , w_43217 , w_43218 , w_43219 , w_43220 , w_43221 , w_43222 , w_43223 , w_43224 , w_43225 , 
		w_43226 , w_43227 , w_43228 , w_43229 , w_43230 , w_43231 , w_43232 , w_43233 , w_43234 , w_43235 , 
		w_43236 , w_43237 , w_43238 , w_43239 , w_43240 , w_43241 , w_43242 , w_43243 , w_43244 , w_43245 , 
		w_43246 , w_43247 , w_43248 , w_43249 , w_43250 , w_43251 , w_43252 , w_43253 , w_43254 , w_43255 , 
		w_43256 , w_43257 , w_43258 , w_43259 , w_43260 , w_43261 , w_43262 , w_43263 , w_43264 , w_43265 , 
		w_43266 , w_43267 , w_43268 , w_43269 , w_43270 , w_43271 , w_43272 , w_43273 , w_43274 , w_43275 , 
		w_43276 , w_43277 , w_43278 , w_43279 , w_43280 , w_43281 , w_43282 , w_43283 , w_43284 , w_43285 , 
		w_43286 , w_43287 , w_43288 , w_43289 , w_43290 , w_43291 , w_43292 , w_43293 , w_43294 , w_43295 , 
		w_43296 , w_43297 , w_43298 , w_43299 , w_43300 , w_43301 , w_43302 , w_43303 , w_43304 , w_43305 , 
		w_43306 , w_43307 , w_43308 , w_43309 , w_43310 , w_43311 , w_43312 , w_43313 , w_43314 , w_43315 , 
		w_43316 , w_43317 , w_43318 , w_43319 , w_43320 , w_43321 , w_43322 , w_43323 , w_43324 , w_43325 , 
		w_43326 , w_43327 , w_43328 , w_43329 , w_43330 , w_43331 , w_43332 , w_43333 , w_43334 , w_43335 , 
		w_43336 , w_43337 , w_43338 , w_43339 , w_43340 , w_43341 , w_43342 , w_43343 , w_43344 , w_43345 , 
		w_43346 , w_43347 , w_43348 , w_43349 , w_43350 , w_43351 , w_43352 , w_43353 , w_43354 , w_43355 , 
		w_43356 , w_43357 , w_43358 , w_43359 , w_43360 , w_43361 , w_43362 , w_43363 , w_43364 , w_43365 , 
		w_43366 , w_43367 , w_43368 , w_43369 , w_43370 , w_43371 , w_43372 , w_43373 , w_43374 , w_43375 , 
		w_43376 , w_43377 , w_43378 , w_43379 , w_43380 , w_43381 , w_43382 , w_43383 , w_43384 , w_43385 , 
		w_43386 , w_43387 , w_43388 , w_43389 , w_43390 , w_43391 , w_43392 , w_43393 , w_43394 , w_43395 , 
		w_43396 , w_43397 , w_43398 , w_43399 , w_43400 , w_43401 , w_43402 , w_43403 , w_43404 , w_43405 , 
		w_43406 , w_43407 , w_43408 , w_43409 , w_43410 , w_43411 , w_43412 , w_43413 , w_43414 , w_43415 , 
		w_43416 , w_43417 , w_43418 , w_43419 , w_43420 , w_43421 , w_43422 , w_43423 , w_43424 , w_43425 , 
		w_43426 , w_43427 , w_43428 , w_43429 , w_43430 , w_43431 , w_43432 , w_43433 , w_43434 , w_43435 , 
		w_43436 , w_43437 , w_43438 , w_43439 , w_43440 , w_43441 , w_43442 , w_43443 , w_43444 , w_43445 , 
		w_43446 , w_43447 , w_43448 , w_43449 , w_43450 , w_43451 , w_43452 , w_43453 , w_43454 , w_43455 , 
		w_43456 , w_43457 , w_43458 , w_43459 , w_43460 , w_43461 , w_43462 , w_43463 , w_43464 , w_43465 , 
		w_43466 , w_43467 , w_43468 , w_43469 , w_43470 , w_43471 , w_43472 , w_43473 , w_43474 , w_43475 , 
		w_43476 , w_43477 , w_43478 , w_43479 , w_43480 , w_43481 , w_43482 , w_43483 , w_43484 , w_43485 , 
		w_43486 , w_43487 , w_43488 , w_43489 , w_43490 , w_43491 , w_43492 , w_43493 , w_43494 , w_43495 , 
		w_43496 , w_43497 , w_43498 , w_43499 , w_43500 , w_43501 , w_43502 , w_43503 , w_43504 , w_43505 , 
		w_43506 , w_43507 , w_43508 , w_43509 , w_43510 , w_43511 , w_43512 , w_43513 , w_43514 , w_43515 , 
		w_43516 , w_43517 , w_43518 , w_43519 , w_43520 , w_43521 , w_43522 , w_43523 , w_43524 , w_43525 , 
		w_43526 , w_43527 , w_43528 , w_43529 , w_43530 , w_43531 , w_43532 , w_43533 , w_43534 , w_43535 , 
		w_43536 , w_43537 , w_43538 , w_43539 , w_43540 , w_43541 , w_43542 , w_43543 , w_43544 , w_43545 , 
		w_43546 , w_43547 , w_43548 , w_43549 , w_43550 , w_43551 , w_43552 , w_43553 , w_43554 , w_43555 , 
		w_43556 , w_43557 , w_43558 , w_43559 , w_43560 , w_43561 , w_43562 , w_43563 , w_43564 , w_43565 , 
		w_43566 , w_43567 , w_43568 , w_43569 , w_43570 , w_43571 , w_43572 , w_43573 , w_43574 , w_43575 , 
		w_43576 , w_43577 , w_43578 , w_43579 , w_43580 , w_43581 , w_43582 , w_43583 , w_43584 , w_43585 , 
		w_43586 , w_43587 , w_43588 , w_43589 , w_43590 , w_43591 , w_43592 , w_43593 , w_43594 , w_43595 , 
		w_43596 , w_43597 , w_43598 , w_43599 , w_43600 , w_43601 , w_43602 , w_43603 , w_43604 , w_43605 , 
		w_43606 , w_43607 , w_43608 , w_43609 , w_43610 , w_43611 , w_43612 , w_43613 , w_43614 , w_43615 , 
		w_43616 , w_43617 , w_43618 , w_43619 , w_43620 , w_43621 , w_43622 , w_43623 , w_43624 , w_43625 , 
		w_43626 , w_43627 , w_43628 , w_43629 , w_43630 , w_43631 , w_43632 , w_43633 , w_43634 , w_43635 , 
		w_43636 , w_43637 , w_43638 , w_43639 , w_43640 , w_43641 , w_43642 , w_43643 , w_43644 , w_43645 , 
		w_43646 , w_43647 , w_43648 , w_43649 , w_43650 , w_43651 , w_43652 , w_43653 , w_43654 , w_43655 , 
		w_43656 , w_43657 , w_43658 , w_43659 , w_43660 , w_43661 , w_43662 , w_43663 , w_43664 , w_43665 , 
		w_43666 , w_43667 , w_43668 , w_43669 , w_43670 , w_43671 , w_43672 , w_43673 , w_43674 , w_43675 , 
		w_43676 , w_43677 , w_43678 , w_43679 , w_43680 , w_43681 , w_43682 , w_43683 , w_43684 , w_43685 , 
		w_43686 , w_43687 , w_43688 , w_43689 , w_43690 , w_43691 , w_43692 , w_43693 , w_43694 , w_43695 , 
		w_43696 , w_43697 , w_43698 , w_43699 , w_43700 , w_43701 , w_43702 , w_43703 , w_43704 , w_43705 , 
		w_43706 , w_43707 , w_43708 , w_43709 , w_43710 , w_43711 , w_43712 , w_43713 , w_43714 , w_43715 , 
		w_43716 , w_43717 , w_43718 , w_43719 , w_43720 , w_43721 , w_43722 , w_43723 , w_43724 , w_43725 , 
		w_43726 , w_43727 , w_43728 , w_43729 , w_43730 , w_43731 , w_43732 , w_43733 , w_43734 , w_43735 , 
		w_43736 , w_43737 , w_43738 , w_43739 , w_43740 , w_43741 , w_43742 , w_43743 , w_43744 , w_43745 , 
		w_43746 , w_43747 , w_43748 , w_43749 , w_43750 , w_43751 , w_43752 , w_43753 , w_43754 , w_43755 , 
		w_43756 , w_43757 , w_43758 , w_43759 , w_43760 , w_43761 , w_43762 , w_43763 , w_43764 , w_43765 , 
		w_43766 , w_43767 , w_43768 , w_43769 , w_43770 , w_43771 , w_43772 , w_43773 , w_43774 , w_43775 , 
		w_43776 , w_43777 , w_43778 , w_43779 , w_43780 , w_43781 , w_43782 , w_43783 , w_43784 , w_43785 , 
		w_43786 , w_43787 , w_43788 , w_43789 , w_43790 , w_43791 , w_43792 , w_43793 , w_43794 , w_43795 , 
		w_43796 , w_43797 , w_43798 , w_43799 , w_43800 , w_43801 , w_43802 , w_43803 , w_43804 , w_43805 , 
		w_43806 , w_43807 , w_43808 , w_43809 , w_43810 , w_43811 , w_43812 , w_43813 , w_43814 , w_43815 , 
		w_43816 , w_43817 , w_43818 , w_43819 , w_43820 , w_43821 , w_43822 , w_43823 , w_43824 , w_43825 , 
		w_43826 , w_43827 , w_43828 , w_43829 , w_43830 , w_43831 , w_43832 , w_43833 , w_43834 , w_43835 , 
		w_43836 , w_43837 , w_43838 , w_43839 , w_43840 , w_43841 , w_43842 , w_43843 , w_43844 , w_43845 , 
		w_43846 , w_43847 , w_43848 , w_43849 , w_43850 , w_43851 , w_43852 , w_43853 , w_43854 , w_43855 , 
		w_43856 , w_43857 , w_43858 , w_43859 , w_43860 , w_43861 , w_43862 , w_43863 , w_43864 , w_43865 , 
		w_43866 , w_43867 , w_43868 , w_43869 , w_43870 , w_43871 , w_43872 , w_43873 , w_43874 , w_43875 , 
		w_43876 , w_43877 , w_43878 , w_43879 , w_43880 , w_43881 , w_43882 , w_43883 , w_43884 , w_43885 , 
		w_43886 , w_43887 , w_43888 , w_43889 , w_43890 , w_43891 , w_43892 , w_43893 , w_43894 , w_43895 , 
		w_43896 , w_43897 , w_43898 , w_43899 , w_43900 , w_43901 , w_43902 , w_43903 , w_43904 , w_43905 , 
		w_43906 , w_43907 , w_43908 , w_43909 , w_43910 , w_43911 , w_43912 , w_43913 , w_43914 , w_43915 , 
		w_43916 , w_43917 , w_43918 , w_43919 , w_43920 , w_43921 , w_43922 , w_43923 , w_43924 , w_43925 , 
		w_43926 , w_43927 , w_43928 , w_43929 , w_43930 , w_43931 , w_43932 , w_43933 , w_43934 , w_43935 , 
		w_43936 , w_43937 , w_43938 , w_43939 , w_43940 , w_43941 , w_43942 , w_43943 , w_43944 , w_43945 , 
		w_43946 , w_43947 , w_43948 , w_43949 , w_43950 , w_43951 , w_43952 , w_43953 , w_43954 , w_43955 , 
		w_43956 , w_43957 , w_43958 , w_43959 , w_43960 , w_43961 , w_43962 , w_43963 , w_43964 , w_43965 , 
		w_43966 , w_43967 , w_43968 , w_43969 , w_43970 , w_43971 , w_43972 , w_43973 , w_43974 , w_43975 , 
		w_43976 , w_43977 , w_43978 , w_43979 , w_43980 , w_43981 , w_43982 , w_43983 , w_43984 , w_43985 , 
		w_43986 , w_43987 , w_43988 , w_43989 , w_43990 , w_43991 , w_43992 , w_43993 , w_43994 , w_43995 , 
		w_43996 , w_43997 , w_43998 , w_43999 , w_44000 , w_44001 , w_44002 , w_44003 , w_44004 , w_44005 , 
		w_44006 , w_44007 , w_44008 , w_44009 , w_44010 , w_44011 , w_44012 , w_44013 , w_44014 , w_44015 , 
		w_44016 , w_44017 , w_44018 , w_44019 , w_44020 , w_44021 , w_44022 , w_44023 , w_44024 , w_44025 , 
		w_44026 , w_44027 , w_44028 , w_44029 , w_44030 , w_44031 , w_44032 , w_44033 , w_44034 , w_44035 , 
		w_44036 , w_44037 , w_44038 , w_44039 , w_44040 , w_44041 , w_44042 , w_44043 , w_44044 , w_44045 , 
		w_44046 , w_44047 , w_44048 , w_44049 , w_44050 , w_44051 , w_44052 , w_44053 , w_44054 , w_44055 , 
		w_44056 , w_44057 , w_44058 , w_44059 , w_44060 , w_44061 , w_44062 , w_44063 , w_44064 , w_44065 , 
		w_44066 , w_44067 , w_44068 , w_44069 , w_44070 , w_44071 , w_44072 , w_44073 , w_44074 , w_44075 , 
		w_44076 , w_44077 , w_44078 , w_44079 , w_44080 , w_44081 , w_44082 , w_44083 , w_44084 , w_44085 , 
		w_44086 , w_44087 , w_44088 , w_44089 , w_44090 , w_44091 , w_44092 , w_44093 , w_44094 , w_44095 , 
		w_44096 , w_44097 , w_44098 , w_44099 , w_44100 , w_44101 , w_44102 , w_44103 , w_44104 , w_44105 , 
		w_44106 , w_44107 , w_44108 , w_44109 , w_44110 , w_44111 , w_44112 , w_44113 , w_44114 , w_44115 , 
		w_44116 , w_44117 , w_44118 , w_44119 , w_44120 , w_44121 , w_44122 , w_44123 , w_44124 , w_44125 , 
		w_44126 , w_44127 , w_44128 , w_44129 , w_44130 , w_44131 , w_44132 , w_44133 , w_44134 , w_44135 , 
		w_44136 , w_44137 , w_44138 , w_44139 , w_44140 , w_44141 , w_44142 , w_44143 , w_44144 , w_44145 , 
		w_44146 , w_44147 , w_44148 , w_44149 , w_44150 , w_44151 , w_44152 , w_44153 , w_44154 , w_44155 , 
		w_44156 , w_44157 , w_44158 , w_44159 , w_44160 , w_44161 , w_44162 , w_44163 , w_44164 , w_44165 , 
		w_44166 , w_44167 , w_44168 , w_44169 , w_44170 , w_44171 , w_44172 , w_44173 , w_44174 , w_44175 , 
		w_44176 , w_44177 , w_44178 , w_44179 , w_44180 , w_44181 , w_44182 , w_44183 , w_44184 , w_44185 , 
		w_44186 , w_44187 , w_44188 , w_44189 , w_44190 , w_44191 , w_44192 , w_44193 , w_44194 , w_44195 , 
		w_44196 , w_44197 , w_44198 , w_44199 , w_44200 , w_44201 , w_44202 , w_44203 , w_44204 , w_44205 , 
		w_44206 , w_44207 , w_44208 , w_44209 , w_44210 , w_44211 , w_44212 , w_44213 , w_44214 , w_44215 , 
		w_44216 , w_44217 , w_44218 , w_44219 , w_44220 , w_44221 , w_44222 , w_44223 , w_44224 , w_44225 , 
		w_44226 , w_44227 , w_44228 , w_44229 , w_44230 , w_44231 , w_44232 , w_44233 , w_44234 , w_44235 , 
		w_44236 , w_44237 , w_44238 , w_44239 , w_44240 , w_44241 , w_44242 , w_44243 , w_44244 , w_44245 , 
		w_44246 , w_44247 , w_44248 , w_44249 , w_44250 , w_44251 , w_44252 , w_44253 , w_44254 , w_44255 , 
		w_44256 , w_44257 , w_44258 , w_44259 , w_44260 , w_44261 , w_44262 , w_44263 , w_44264 , w_44265 , 
		w_44266 , w_44267 , w_44268 , w_44269 , w_44270 , w_44271 , w_44272 , w_44273 , w_44274 , w_44275 , 
		w_44276 , w_44277 , w_44278 , w_44279 , w_44280 , w_44281 , w_44282 , w_44283 , w_44284 , w_44285 , 
		w_44286 , w_44287 , w_44288 , w_44289 , w_44290 , w_44291 , w_44292 , w_44293 , w_44294 , w_44295 , 
		w_44296 , w_44297 , w_44298 , w_44299 , w_44300 , w_44301 , w_44302 , w_44303 , w_44304 , w_44305 , 
		w_44306 , w_44307 , w_44308 , w_44309 , w_44310 , w_44311 , w_44312 , w_44313 , w_44314 , w_44315 , 
		w_44316 , w_44317 , w_44318 , w_44319 , w_44320 , w_44321 , w_44322 , w_44323 , w_44324 , w_44325 , 
		w_44326 , w_44327 , w_44328 , w_44329 , w_44330 , w_44331 , w_44332 , w_44333 , w_44334 , w_44335 , 
		w_44336 , w_44337 , w_44338 , w_44339 , w_44340 , w_44341 , w_44342 , w_44343 , w_44344 , w_44345 , 
		w_44346 , w_44347 , w_44348 , w_44349 , w_44350 , w_44351 , w_44352 , w_44353 , w_44354 , w_44355 , 
		w_44356 , w_44357 , w_44358 , w_44359 , w_44360 , w_44361 , w_44362 , w_44363 , w_44364 , w_44365 , 
		w_44366 , w_44367 , w_44368 , w_44369 , w_44370 , w_44371 , w_44372 , w_44373 , w_44374 , w_44375 , 
		w_44376 , w_44377 , w_44378 , w_44379 , w_44380 , w_44381 , w_44382 , w_44383 , w_44384 , w_44385 , 
		w_44386 , w_44387 , w_44388 , w_44389 , w_44390 , w_44391 , w_44392 , w_44393 , w_44394 , w_44395 , 
		w_44396 , w_44397 , w_44398 , w_44399 , w_44400 , w_44401 , w_44402 , w_44403 , w_44404 , w_44405 , 
		w_44406 , w_44407 , w_44408 , w_44409 , w_44410 , w_44411 , w_44412 , w_44413 , w_44414 , w_44415 , 
		w_44416 , w_44417 , w_44418 , w_44419 , w_44420 , w_44421 , w_44422 , w_44423 , w_44424 , w_44425 , 
		w_44426 , w_44427 , w_44428 , w_44429 , w_44430 , w_44431 , w_44432 , w_44433 , w_44434 , w_44435 , 
		w_44436 , w_44437 , w_44438 , w_44439 , w_44440 , w_44441 , w_44442 , w_44443 , w_44444 , w_44445 , 
		w_44446 , w_44447 , w_44448 , w_44449 , w_44450 , w_44451 , w_44452 , w_44453 , w_44454 , w_44455 , 
		w_44456 , w_44457 , w_44458 , w_44459 , w_44460 , w_44461 , w_44462 , w_44463 , w_44464 , w_44465 , 
		w_44466 , w_44467 , w_44468 , w_44469 , w_44470 , w_44471 , w_44472 , w_44473 , w_44474 , w_44475 , 
		w_44476 , w_44477 , w_44478 , w_44479 , w_44480 , w_44481 , w_44482 , w_44483 , w_44484 , w_44485 , 
		w_44486 , w_44487 , w_44488 , w_44489 , w_44490 , w_44491 , w_44492 , w_44493 , w_44494 , w_44495 , 
		w_44496 , w_44497 , w_44498 , w_44499 , w_44500 , w_44501 , w_44502 , w_44503 , w_44504 , w_44505 , 
		w_44506 , w_44507 , w_44508 , w_44509 , w_44510 , w_44511 , w_44512 , w_44513 , w_44514 , w_44515 , 
		w_44516 , w_44517 , w_44518 , w_44519 , w_44520 , w_44521 , w_44522 , w_44523 , w_44524 , w_44525 , 
		w_44526 , w_44527 , w_44528 , w_44529 , w_44530 , w_44531 , w_44532 , w_44533 , w_44534 , w_44535 , 
		w_44536 , w_44537 , w_44538 , w_44539 , w_44540 , w_44541 , w_44542 , w_44543 , w_44544 , w_44545 , 
		w_44546 , w_44547 , w_44548 , w_44549 , w_44550 , w_44551 , w_44552 , w_44553 , w_44554 , w_44555 , 
		w_44556 , w_44557 , w_44558 , w_44559 , w_44560 , w_44561 , w_44562 , w_44563 , w_44564 , w_44565 , 
		w_44566 , w_44567 , w_44568 , w_44569 , w_44570 , w_44571 , w_44572 , w_44573 , w_44574 , w_44575 , 
		w_44576 , w_44577 , w_44578 , w_44579 , w_44580 , w_44581 , w_44582 , w_44583 , w_44584 , w_44585 , 
		w_44586 , w_44587 , w_44588 , w_44589 , w_44590 , w_44591 , w_44592 , w_44593 , w_44594 , w_44595 , 
		w_44596 , w_44597 , w_44598 , w_44599 , w_44600 , w_44601 , w_44602 , w_44603 , w_44604 , w_44605 , 
		w_44606 , w_44607 , w_44608 , w_44609 , w_44610 , w_44611 , w_44612 , w_44613 , w_44614 , w_44615 , 
		w_44616 , w_44617 , w_44618 , w_44619 , w_44620 , w_44621 , w_44622 , w_44623 , w_44624 , w_44625 , 
		w_44626 , w_44627 , w_44628 , w_44629 , w_44630 , w_44631 , w_44632 , w_44633 , w_44634 , w_44635 , 
		w_44636 , w_44637 , w_44638 , w_44639 , w_44640 , w_44641 , w_44642 , w_44643 , w_44644 , w_44645 , 
		w_44646 , w_44647 , w_44648 , w_44649 , w_44650 , w_44651 , w_44652 , w_44653 , w_44654 , w_44655 , 
		w_44656 , w_44657 , w_44658 , w_44659 , w_44660 , w_44661 , w_44662 , w_44663 , w_44664 , w_44665 , 
		w_44666 , w_44667 , w_44668 , w_44669 , w_44670 , w_44671 , w_44672 , w_44673 , w_44674 , w_44675 , 
		w_44676 , w_44677 , w_44678 , w_44679 , w_44680 , w_44681 , w_44682 , w_44683 , w_44684 , w_44685 , 
		w_44686 , w_44687 , w_44688 , w_44689 , w_44690 , w_44691 , w_44692 , w_44693 , w_44694 , w_44695 , 
		w_44696 , w_44697 , w_44698 , w_44699 , w_44700 , w_44701 , w_44702 , w_44703 , w_44704 , w_44705 , 
		w_44706 , w_44707 , w_44708 , w_44709 , w_44710 , w_44711 , w_44712 , w_44713 , w_44714 , w_44715 , 
		w_44716 , w_44717 , w_44718 , w_44719 , w_44720 , w_44721 , w_44722 , w_44723 , w_44724 , w_44725 , 
		w_44726 , w_44727 , w_44728 , w_44729 , w_44730 , w_44731 , w_44732 , w_44733 , w_44734 , w_44735 , 
		w_44736 , w_44737 , w_44738 , w_44739 , w_44740 , w_44741 , w_44742 , w_44743 , w_44744 , w_44745 , 
		w_44746 , w_44747 , w_44748 , w_44749 , w_44750 , w_44751 , w_44752 , w_44753 , w_44754 , w_44755 , 
		w_44756 , w_44757 , w_44758 , w_44759 , w_44760 , w_44761 , w_44762 , w_44763 , w_44764 , w_44765 , 
		w_44766 , w_44767 , w_44768 , w_44769 , w_44770 , w_44771 , w_44772 , w_44773 , w_44774 , w_44775 , 
		w_44776 , w_44777 , w_44778 , w_44779 , w_44780 , w_44781 , w_44782 , w_44783 , w_44784 , w_44785 , 
		w_44786 , w_44787 , w_44788 , w_44789 , w_44790 , w_44791 , w_44792 , w_44793 , w_44794 , w_44795 , 
		w_44796 , w_44797 , w_44798 , w_44799 , w_44800 , w_44801 , w_44802 , w_44803 , w_44804 , w_44805 , 
		w_44806 , w_44807 , w_44808 , w_44809 , w_44810 , w_44811 , w_44812 , w_44813 , w_44814 , w_44815 , 
		w_44816 , w_44817 , w_44818 , w_44819 , w_44820 , w_44821 , w_44822 , w_44823 , w_44824 , w_44825 , 
		w_44826 , w_44827 , w_44828 , w_44829 , w_44830 , w_44831 , w_44832 , w_44833 , w_44834 , w_44835 , 
		w_44836 , w_44837 , w_44838 , w_44839 , w_44840 , w_44841 , w_44842 , w_44843 , w_44844 , w_44845 , 
		w_44846 , w_44847 , w_44848 , w_44849 , w_44850 , w_44851 , w_44852 , w_44853 , w_44854 , w_44855 , 
		w_44856 , w_44857 , w_44858 , w_44859 , w_44860 , w_44861 , w_44862 , w_44863 , w_44864 , w_44865 , 
		w_44866 , w_44867 , w_44868 , w_44869 , w_44870 , w_44871 , w_44872 , w_44873 , w_44874 , w_44875 , 
		w_44876 , w_44877 , w_44878 , w_44879 , w_44880 , w_44881 , w_44882 , w_44883 , w_44884 , w_44885 , 
		w_44886 , w_44887 , w_44888 , w_44889 , w_44890 , w_44891 , w_44892 , w_44893 , w_44894 , w_44895 , 
		w_44896 , w_44897 , w_44898 , w_44899 , w_44900 , w_44901 , w_44902 , w_44903 , w_44904 , w_44905 , 
		w_44906 , w_44907 , w_44908 , w_44909 , w_44910 , w_44911 , w_44912 , w_44913 , w_44914 , w_44915 , 
		w_44916 , w_44917 , w_44918 , w_44919 , w_44920 , w_44921 , w_44922 , w_44923 , w_44924 , w_44925 , 
		w_44926 , w_44927 , w_44928 , w_44929 , w_44930 , w_44931 , w_44932 , w_44933 , w_44934 , w_44935 , 
		w_44936 , w_44937 , w_44938 , w_44939 , w_44940 , w_44941 , w_44942 , w_44943 , w_44944 , w_44945 , 
		w_44946 , w_44947 , w_44948 , w_44949 , w_44950 , w_44951 , w_44952 , w_44953 , w_44954 , w_44955 , 
		w_44956 , w_44957 , w_44958 , w_44959 , w_44960 , w_44961 , w_44962 , w_44963 , w_44964 , w_44965 , 
		w_44966 , w_44967 , w_44968 , w_44969 , w_44970 , w_44971 , w_44972 , w_44973 , w_44974 , w_44975 , 
		w_44976 , w_44977 , w_44978 , w_44979 , w_44980 , w_44981 , w_44982 , w_44983 , w_44984 , w_44985 , 
		w_44986 , w_44987 , w_44988 , w_44989 , w_44990 , w_44991 , w_44992 , w_44993 , w_44994 , w_44995 , 
		w_44996 , w_44997 , w_44998 , w_44999 , w_45000 , w_45001 , w_45002 , w_45003 , w_45004 , w_45005 , 
		w_45006 , w_45007 , w_45008 , w_45009 , w_45010 , w_45011 , w_45012 , w_45013 , w_45014 , w_45015 , 
		w_45016 , w_45017 , w_45018 , w_45019 , w_45020 , w_45021 , w_45022 , w_45023 , w_45024 , w_45025 , 
		w_45026 , w_45027 , w_45028 , w_45029 , w_45030 , w_45031 , w_45032 , w_45033 , w_45034 , w_45035 , 
		w_45036 , w_45037 , w_45038 , w_45039 , w_45040 , w_45041 , w_45042 , w_45043 , w_45044 , w_45045 , 
		w_45046 , w_45047 , w_45048 , w_45049 , w_45050 , w_45051 , w_45052 , w_45053 , w_45054 , w_45055 , 
		w_45056 , w_45057 , w_45058 , w_45059 , w_45060 , w_45061 , w_45062 , w_45063 , w_45064 , w_45065 , 
		w_45066 , w_45067 , w_45068 , w_45069 , w_45070 , w_45071 , w_45072 , w_45073 , w_45074 , w_45075 , 
		w_45076 , w_45077 , w_45078 , w_45079 , w_45080 , w_45081 , w_45082 , w_45083 , w_45084 , w_45085 , 
		w_45086 , w_45087 , w_45088 , w_45089 , w_45090 , w_45091 , w_45092 , w_45093 , w_45094 , w_45095 , 
		w_45096 , w_45097 , w_45098 , w_45099 , w_45100 , w_45101 , w_45102 , w_45103 , w_45104 , w_45105 , 
		w_45106 , w_45107 , w_45108 , w_45109 , w_45110 , w_45111 , w_45112 , w_45113 , w_45114 , w_45115 , 
		w_45116 , w_45117 , w_45118 , w_45119 , w_45120 , w_45121 , w_45122 , w_45123 , w_45124 , w_45125 , 
		w_45126 , w_45127 , w_45128 , w_45129 , w_45130 , w_45131 , w_45132 , w_45133 , w_45134 , w_45135 , 
		w_45136 , w_45137 , w_45138 , w_45139 , w_45140 , w_45141 , w_45142 , w_45143 , w_45144 , w_45145 , 
		w_45146 , w_45147 , w_45148 , w_45149 , w_45150 , w_45151 , w_45152 , w_45153 , w_45154 , w_45155 , 
		w_45156 , w_45157 , w_45158 , w_45159 , w_45160 , w_45161 , w_45162 , w_45163 , w_45164 , w_45165 , 
		w_45166 , w_45167 , w_45168 , w_45169 , w_45170 , w_45171 , w_45172 , w_45173 , w_45174 , w_45175 , 
		w_45176 , w_45177 , w_45178 , w_45179 , w_45180 , w_45181 , w_45182 , w_45183 , w_45184 , w_45185 , 
		w_45186 , w_45187 , w_45188 , w_45189 , w_45190 , w_45191 , w_45192 , w_45193 , w_45194 , w_45195 , 
		w_45196 , w_45197 , w_45198 , w_45199 , w_45200 , w_45201 , w_45202 , w_45203 , w_45204 , w_45205 , 
		w_45206 , w_45207 , w_45208 , w_45209 , w_45210 , w_45211 , w_45212 , w_45213 , w_45214 , w_45215 , 
		w_45216 , w_45217 , w_45218 , w_45219 , w_45220 , w_45221 , w_45222 , w_45223 , w_45224 , w_45225 , 
		w_45226 , w_45227 , w_45228 , w_45229 , w_45230 , w_45231 , w_45232 , w_45233 , w_45234 , w_45235 , 
		w_45236 , w_45237 , w_45238 , w_45239 , w_45240 , w_45241 , w_45242 , w_45243 , w_45244 , w_45245 , 
		w_45246 , w_45247 , w_45248 , w_45249 , w_45250 , w_45251 , w_45252 , w_45253 , w_45254 , w_45255 , 
		w_45256 , w_45257 , w_45258 , w_45259 , w_45260 , w_45261 , w_45262 , w_45263 , w_45264 , w_45265 , 
		w_45266 , w_45267 , w_45268 , w_45269 , w_45270 , w_45271 , w_45272 , w_45273 , w_45274 , w_45275 , 
		w_45276 , w_45277 , w_45278 , w_45279 , w_45280 , w_45281 , w_45282 , w_45283 , w_45284 , w_45285 , 
		w_45286 , w_45287 , w_45288 , w_45289 , w_45290 , w_45291 , w_45292 , w_45293 , w_45294 , w_45295 , 
		w_45296 , w_45297 , w_45298 , w_45299 , w_45300 , w_45301 , w_45302 , w_45303 , w_45304 , w_45305 , 
		w_45306 , w_45307 , w_45308 , w_45309 , w_45310 , w_45311 , w_45312 , w_45313 , w_45314 , w_45315 , 
		w_45316 , w_45317 , w_45318 , w_45319 , w_45320 , w_45321 , w_45322 , w_45323 , w_45324 , w_45325 , 
		w_45326 , w_45327 , w_45328 , w_45329 , w_45330 , w_45331 , w_45332 , w_45333 , w_45334 , w_45335 , 
		w_45336 , w_45337 , w_45338 , w_45339 , w_45340 , w_45341 , w_45342 , w_45343 , w_45344 , w_45345 , 
		w_45346 , w_45347 , w_45348 , w_45349 , w_45350 , w_45351 , w_45352 , w_45353 , w_45354 , w_45355 , 
		w_45356 , w_45357 , w_45358 , w_45359 , w_45360 , w_45361 , w_45362 , w_45363 , w_45364 , w_45365 , 
		w_45366 , w_45367 , w_45368 , w_45369 , w_45370 , w_45371 , w_45372 , w_45373 , w_45374 , w_45375 , 
		w_45376 , w_45377 , w_45378 , w_45379 , w_45380 , w_45381 , w_45382 , w_45383 , w_45384 , w_45385 , 
		w_45386 , w_45387 , w_45388 , w_45389 , w_45390 , w_45391 , w_45392 , w_45393 , w_45394 , w_45395 , 
		w_45396 , w_45397 , w_45398 , w_45399 , w_45400 , w_45401 , w_45402 , w_45403 , w_45404 , w_45405 , 
		w_45406 , w_45407 , w_45408 , w_45409 , w_45410 , w_45411 , w_45412 , w_45413 , w_45414 , w_45415 , 
		w_45416 , w_45417 , w_45418 , w_45419 , w_45420 , w_45421 , w_45422 , w_45423 , w_45424 , w_45425 , 
		w_45426 , w_45427 , w_45428 , w_45429 , w_45430 , w_45431 , w_45432 , w_45433 , w_45434 , w_45435 , 
		w_45436 , w_45437 , w_45438 , w_45439 , w_45440 , w_45441 , w_45442 , w_45443 , w_45444 , w_45445 , 
		w_45446 , w_45447 , w_45448 , w_45449 , w_45450 , w_45451 , w_45452 , w_45453 , w_45454 , w_45455 , 
		w_45456 , w_45457 , w_45458 , w_45459 , w_45460 , w_45461 , w_45462 , w_45463 , w_45464 , w_45465 , 
		w_45466 , w_45467 , w_45468 , w_45469 , w_45470 , w_45471 , w_45472 , w_45473 , w_45474 , w_45475 , 
		w_45476 , w_45477 , w_45478 , w_45479 , w_45480 , w_45481 , w_45482 , w_45483 , w_45484 , w_45485 , 
		w_45486 , w_45487 , w_45488 , w_45489 , w_45490 , w_45491 , w_45492 , w_45493 , w_45494 , w_45495 , 
		w_45496 , w_45497 , w_45498 , w_45499 , w_45500 , w_45501 , w_45502 , w_45503 , w_45504 , w_45505 , 
		w_45506 , w_45507 , w_45508 , w_45509 , w_45510 , w_45511 , w_45512 , w_45513 , w_45514 , w_45515 , 
		w_45516 , w_45517 , w_45518 , w_45519 , w_45520 , w_45521 , w_45522 , w_45523 , w_45524 , w_45525 , 
		w_45526 , w_45527 , w_45528 , w_45529 , w_45530 , w_45531 , w_45532 , w_45533 , w_45534 , w_45535 , 
		w_45536 , w_45537 , w_45538 , w_45539 , w_45540 , w_45541 , w_45542 , w_45543 , w_45544 , w_45545 , 
		w_45546 , w_45547 , w_45548 , w_45549 , w_45550 , w_45551 , w_45552 , w_45553 , w_45554 , w_45555 , 
		w_45556 , w_45557 , w_45558 , w_45559 , w_45560 , w_45561 , w_45562 , w_45563 , w_45564 , w_45565 , 
		w_45566 , w_45567 , w_45568 , w_45569 , w_45570 , w_45571 , w_45572 , w_45573 , w_45574 , w_45575 , 
		w_45576 , w_45577 , w_45578 , w_45579 , w_45580 , w_45581 , w_45582 , w_45583 , w_45584 , w_45585 , 
		w_45586 , w_45587 , w_45588 , w_45589 , w_45590 , w_45591 , w_45592 , w_45593 , w_45594 , w_45595 , 
		w_45596 , w_45597 , w_45598 , w_45599 , w_45600 , w_45601 , w_45602 , w_45603 , w_45604 , w_45605 , 
		w_45606 , w_45607 , w_45608 , w_45609 , w_45610 , w_45611 , w_45612 , w_45613 , w_45614 , w_45615 , 
		w_45616 , w_45617 , w_45618 , w_45619 , w_45620 , w_45621 , w_45622 , w_45623 , w_45624 , w_45625 , 
		w_45626 , w_45627 , w_45628 , w_45629 , w_45630 , w_45631 , w_45632 , w_45633 , w_45634 , w_45635 , 
		w_45636 , w_45637 , w_45638 , w_45639 , w_45640 , w_45641 , w_45642 , w_45643 , w_45644 , w_45645 , 
		w_45646 , w_45647 , w_45648 , w_45649 , w_45650 , w_45651 , w_45652 , w_45653 , w_45654 , w_45655 , 
		w_45656 , w_45657 , w_45658 , w_45659 , w_45660 , w_45661 , w_45662 , w_45663 , w_45664 , w_45665 , 
		w_45666 , w_45667 , w_45668 , w_45669 , w_45670 , w_45671 , w_45672 , w_45673 , w_45674 , w_45675 , 
		w_45676 , w_45677 , w_45678 , w_45679 , w_45680 , w_45681 , w_45682 , w_45683 , w_45684 , w_45685 , 
		w_45686 , w_45687 , w_45688 , w_45689 , w_45690 , w_45691 , w_45692 , w_45693 , w_45694 , w_45695 , 
		w_45696 , w_45697 , w_45698 , w_45699 , w_45700 , w_45701 , w_45702 , w_45703 , w_45704 , w_45705 , 
		w_45706 , w_45707 , w_45708 , w_45709 , w_45710 , w_45711 , w_45712 , w_45713 , w_45714 , w_45715 , 
		w_45716 , w_45717 , w_45718 , w_45719 , w_45720 , w_45721 , w_45722 , w_45723 , w_45724 , w_45725 , 
		w_45726 , w_45727 , w_45728 , w_45729 , w_45730 , w_45731 , w_45732 , w_45733 , w_45734 , w_45735 , 
		w_45736 , w_45737 , w_45738 , w_45739 , w_45740 , w_45741 , w_45742 , w_45743 , w_45744 , w_45745 , 
		w_45746 , w_45747 , w_45748 , w_45749 , w_45750 , w_45751 , w_45752 , w_45753 , w_45754 , w_45755 , 
		w_45756 , w_45757 , w_45758 , w_45759 , w_45760 , w_45761 , w_45762 , w_45763 , w_45764 , w_45765 , 
		w_45766 , w_45767 , w_45768 , w_45769 , w_45770 , w_45771 , w_45772 , w_45773 , w_45774 , w_45775 , 
		w_45776 , w_45777 , w_45778 , w_45779 , w_45780 , w_45781 , w_45782 , w_45783 , w_45784 , w_45785 , 
		w_45786 , w_45787 , w_45788 , w_45789 , w_45790 , w_45791 , w_45792 , w_45793 , w_45794 , w_45795 , 
		w_45796 , w_45797 , w_45798 , w_45799 , w_45800 , w_45801 , w_45802 , w_45803 , w_45804 , w_45805 , 
		w_45806 , w_45807 , w_45808 , w_45809 , w_45810 , w_45811 , w_45812 , w_45813 , w_45814 , w_45815 , 
		w_45816 , w_45817 , w_45818 , w_45819 , w_45820 , w_45821 , w_45822 , w_45823 , w_45824 , w_45825 , 
		w_45826 , w_45827 , w_45828 , w_45829 , w_45830 , w_45831 , w_45832 , w_45833 , w_45834 , w_45835 , 
		w_45836 , w_45837 , w_45838 , w_45839 , w_45840 , w_45841 , w_45842 , w_45843 , w_45844 , w_45845 , 
		w_45846 , w_45847 , w_45848 , w_45849 , w_45850 , w_45851 , w_45852 , w_45853 , w_45854 , w_45855 , 
		w_45856 , w_45857 , w_45858 , w_45859 , w_45860 , w_45861 , w_45862 , w_45863 , w_45864 , w_45865 , 
		w_45866 , w_45867 , w_45868 , w_45869 , w_45870 , w_45871 , w_45872 , w_45873 , w_45874 , w_45875 , 
		w_45876 , w_45877 , w_45878 , w_45879 , w_45880 , w_45881 , w_45882 , w_45883 , w_45884 , w_45885 , 
		w_45886 , w_45887 , w_45888 , w_45889 , w_45890 , w_45891 , w_45892 , w_45893 , w_45894 , w_45895 , 
		w_45896 , w_45897 , w_45898 , w_45899 , w_45900 , w_45901 , w_45902 , w_45903 , w_45904 , w_45905 , 
		w_45906 , w_45907 , w_45908 , w_45909 , w_45910 , w_45911 , w_45912 , w_45913 , w_45914 , w_45915 , 
		w_45916 , w_45917 , w_45918 , w_45919 , w_45920 , w_45921 , w_45922 , w_45923 , w_45924 , w_45925 , 
		w_45926 , w_45927 , w_45928 , w_45929 , w_45930 , w_45931 , w_45932 , w_45933 , w_45934 , w_45935 , 
		w_45936 , w_45937 , w_45938 , w_45939 , w_45940 , w_45941 , w_45942 , w_45943 , w_45944 , w_45945 , 
		w_45946 , w_45947 , w_45948 , w_45949 , w_45950 , w_45951 , w_45952 , w_45953 , w_45954 , w_45955 , 
		w_45956 , w_45957 , w_45958 , w_45959 , w_45960 , w_45961 , w_45962 , w_45963 , w_45964 , w_45965 , 
		w_45966 , w_45967 , w_45968 , w_45969 , w_45970 , w_45971 , w_45972 , w_45973 , w_45974 , w_45975 , 
		w_45976 , w_45977 , w_45978 , w_45979 , w_45980 , w_45981 , w_45982 , w_45983 , w_45984 , w_45985 , 
		w_45986 , w_45987 , w_45988 , w_45989 , w_45990 , w_45991 , w_45992 , w_45993 , w_45994 , w_45995 , 
		w_45996 , w_45997 , w_45998 , w_45999 , w_46000 , w_46001 , w_46002 , w_46003 , w_46004 , w_46005 , 
		w_46006 , w_46007 , w_46008 , w_46009 , w_46010 , w_46011 , w_46012 , w_46013 , w_46014 , w_46015 , 
		w_46016 , w_46017 , w_46018 , w_46019 , w_46020 , w_46021 , w_46022 , w_46023 , w_46024 , w_46025 , 
		w_46026 , w_46027 , w_46028 , w_46029 , w_46030 , w_46031 , w_46032 , w_46033 , w_46034 , w_46035 , 
		w_46036 , w_46037 , w_46038 , w_46039 , w_46040 , w_46041 , w_46042 , w_46043 , w_46044 , w_46045 , 
		w_46046 , w_46047 , w_46048 , w_46049 , w_46050 , w_46051 , w_46052 , w_46053 , w_46054 , w_46055 , 
		w_46056 , w_46057 , w_46058 , w_46059 , w_46060 , w_46061 , w_46062 , w_46063 , w_46064 , w_46065 , 
		w_46066 , w_46067 , w_46068 , w_46069 , w_46070 , w_46071 , w_46072 , w_46073 , w_46074 , w_46075 , 
		w_46076 , w_46077 , w_46078 , w_46079 , w_46080 , w_46081 , w_46082 , w_46083 , w_46084 , w_46085 , 
		w_46086 , w_46087 , w_46088 , w_46089 , w_46090 , w_46091 , w_46092 , w_46093 , w_46094 , w_46095 , 
		w_46096 , w_46097 , w_46098 , w_46099 , w_46100 , w_46101 , w_46102 , w_46103 , w_46104 , w_46105 , 
		w_46106 , w_46107 , w_46108 , w_46109 , w_46110 , w_46111 , w_46112 , w_46113 , w_46114 , w_46115 , 
		w_46116 , w_46117 , w_46118 , w_46119 , w_46120 , w_46121 , w_46122 , w_46123 , w_46124 , w_46125 , 
		w_46126 , w_46127 , w_46128 , w_46129 , w_46130 , w_46131 , w_46132 , w_46133 , w_46134 , w_46135 , 
		w_46136 , w_46137 , w_46138 , w_46139 , w_46140 , w_46141 , w_46142 , w_46143 , w_46144 , w_46145 , 
		w_46146 , w_46147 , w_46148 , w_46149 , w_46150 , w_46151 , w_46152 , w_46153 , w_46154 , w_46155 , 
		w_46156 , w_46157 , w_46158 , w_46159 , w_46160 , w_46161 , w_46162 , w_46163 , w_46164 , w_46165 , 
		w_46166 , w_46167 , w_46168 , w_46169 , w_46170 , w_46171 , w_46172 , w_46173 , w_46174 , w_46175 , 
		w_46176 , w_46177 , w_46178 , w_46179 , w_46180 , w_46181 , w_46182 , w_46183 , w_46184 , w_46185 , 
		w_46186 , w_46187 , w_46188 , w_46189 , w_46190 , w_46191 , w_46192 , w_46193 , w_46194 , w_46195 , 
		w_46196 , w_46197 , w_46198 , w_46199 , w_46200 , w_46201 , w_46202 , w_46203 , w_46204 , w_46205 , 
		w_46206 , w_46207 , w_46208 , w_46209 , w_46210 , w_46211 , w_46212 , w_46213 , w_46214 , w_46215 , 
		w_46216 , w_46217 , w_46218 , w_46219 , w_46220 , w_46221 , w_46222 , w_46223 , w_46224 , w_46225 , 
		w_46226 , w_46227 , w_46228 , w_46229 , w_46230 , w_46231 , w_46232 , w_46233 , w_46234 , w_46235 , 
		w_46236 , w_46237 , w_46238 , w_46239 , w_46240 , w_46241 , w_46242 , w_46243 , w_46244 , w_46245 , 
		w_46246 , w_46247 , w_46248 , w_46249 , w_46250 , w_46251 , w_46252 , w_46253 , w_46254 , w_46255 , 
		w_46256 , w_46257 , w_46258 , w_46259 , w_46260 , w_46261 , w_46262 , w_46263 , w_46264 , w_46265 , 
		w_46266 , w_46267 , w_46268 , w_46269 , w_46270 , w_46271 , w_46272 , w_46273 , w_46274 , w_46275 , 
		w_46276 , w_46277 , w_46278 , w_46279 , w_46280 , w_46281 , w_46282 , w_46283 , w_46284 , w_46285 , 
		w_46286 , w_46287 , w_46288 , w_46289 , w_46290 , w_46291 , w_46292 , w_46293 , w_46294 , w_46295 , 
		w_46296 , w_46297 , w_46298 , w_46299 , w_46300 , w_46301 , w_46302 , w_46303 , w_46304 , w_46305 , 
		w_46306 , w_46307 , w_46308 , w_46309 , w_46310 , w_46311 , w_46312 , w_46313 , w_46314 , w_46315 , 
		w_46316 , w_46317 , w_46318 , w_46319 , w_46320 , w_46321 , w_46322 , w_46323 , w_46324 , w_46325 , 
		w_46326 , w_46327 , w_46328 , w_46329 , w_46330 , w_46331 , w_46332 , w_46333 , w_46334 , w_46335 , 
		w_46336 , w_46337 , w_46338 , w_46339 , w_46340 , w_46341 , w_46342 , w_46343 , w_46344 , w_46345 , 
		w_46346 , w_46347 , w_46348 , w_46349 , w_46350 , w_46351 , w_46352 , w_46353 , w_46354 , w_46355 , 
		w_46356 , w_46357 , w_46358 , w_46359 , w_46360 , w_46361 , w_46362 , w_46363 , w_46364 , w_46365 , 
		w_46366 , w_46367 , w_46368 , w_46369 , w_46370 , w_46371 , w_46372 , w_46373 , w_46374 , w_46375 , 
		w_46376 , w_46377 , w_46378 , w_46379 , w_46380 , w_46381 , w_46382 , w_46383 , w_46384 , w_46385 , 
		w_46386 , w_46387 , w_46388 , w_46389 , w_46390 , w_46391 , w_46392 , w_46393 , w_46394 , w_46395 , 
		w_46396 , w_46397 , w_46398 , w_46399 , w_46400 , w_46401 , w_46402 , w_46403 , w_46404 , w_46405 , 
		w_46406 , w_46407 , w_46408 , w_46409 , w_46410 , w_46411 , w_46412 , w_46413 , w_46414 , w_46415 , 
		w_46416 , w_46417 , w_46418 , w_46419 , w_46420 , w_46421 , w_46422 , w_46423 , w_46424 , w_46425 , 
		w_46426 , w_46427 , w_46428 , w_46429 , w_46430 , w_46431 , w_46432 , w_46433 , w_46434 , w_46435 , 
		w_46436 , w_46437 , w_46438 , w_46439 , w_46440 , w_46441 , w_46442 , w_46443 , w_46444 , w_46445 , 
		w_46446 , w_46447 , w_46448 , w_46449 , w_46450 , w_46451 , w_46452 , w_46453 , w_46454 , w_46455 , 
		w_46456 , w_46457 , w_46458 , w_46459 , w_46460 , w_46461 , w_46462 , w_46463 , w_46464 , w_46465 , 
		w_46466 , w_46467 , w_46468 , w_46469 , w_46470 , w_46471 , w_46472 , w_46473 , w_46474 , w_46475 , 
		w_46476 , w_46477 , w_46478 , w_46479 , w_46480 , w_46481 , w_46482 , w_46483 , w_46484 , w_46485 , 
		w_46486 , w_46487 , w_46488 , w_46489 , w_46490 , w_46491 , w_46492 , w_46493 , w_46494 , w_46495 , 
		w_46496 , w_46497 , w_46498 , w_46499 , w_46500 , w_46501 , w_46502 , w_46503 , w_46504 , w_46505 , 
		w_46506 , w_46507 , w_46508 , w_46509 , w_46510 , w_46511 , w_46512 , w_46513 , w_46514 , w_46515 , 
		w_46516 , w_46517 , w_46518 , w_46519 , w_46520 , w_46521 , w_46522 , w_46523 , w_46524 , w_46525 , 
		w_46526 , w_46527 , w_46528 , w_46529 , w_46530 , w_46531 , w_46532 , w_46533 , w_46534 , w_46535 , 
		w_46536 , w_46537 , w_46538 , w_46539 , w_46540 , w_46541 , w_46542 , w_46543 , w_46544 , w_46545 , 
		w_46546 , w_46547 , w_46548 , w_46549 , w_46550 , w_46551 , w_46552 , w_46553 , w_46554 , w_46555 , 
		w_46556 , w_46557 , w_46558 , w_46559 , w_46560 , w_46561 , w_46562 , w_46563 , w_46564 , w_46565 , 
		w_46566 , w_46567 , w_46568 , w_46569 , w_46570 , w_46571 , w_46572 , w_46573 , w_46574 , w_46575 , 
		w_46576 , w_46577 , w_46578 , w_46579 , w_46580 , w_46581 , w_46582 , w_46583 , w_46584 , w_46585 , 
		w_46586 , w_46587 , w_46588 , w_46589 , w_46590 , w_46591 , w_46592 , w_46593 , w_46594 , w_46595 , 
		w_46596 , w_46597 , w_46598 , w_46599 , w_46600 , w_46601 , w_46602 , w_46603 , w_46604 , w_46605 , 
		w_46606 , w_46607 , w_46608 , w_46609 , w_46610 , w_46611 , w_46612 , w_46613 , w_46614 , w_46615 , 
		w_46616 , w_46617 , w_46618 , w_46619 , w_46620 , w_46621 , w_46622 , w_46623 , w_46624 , w_46625 , 
		w_46626 , w_46627 , w_46628 , w_46629 , w_46630 , w_46631 , w_46632 , w_46633 , w_46634 , w_46635 , 
		w_46636 , w_46637 , w_46638 , w_46639 , w_46640 , w_46641 , w_46642 , w_46643 , w_46644 , w_46645 , 
		w_46646 , w_46647 , w_46648 , w_46649 , w_46650 , w_46651 , w_46652 , w_46653 , w_46654 , w_46655 , 
		w_46656 , w_46657 , w_46658 , w_46659 , w_46660 , w_46661 , w_46662 , w_46663 , w_46664 , w_46665 , 
		w_46666 , w_46667 , w_46668 , w_46669 , w_46670 , w_46671 , w_46672 , w_46673 , w_46674 , w_46675 , 
		w_46676 , w_46677 , w_46678 , w_46679 , w_46680 , w_46681 , w_46682 , w_46683 , w_46684 , w_46685 , 
		w_46686 , w_46687 , w_46688 , w_46689 , w_46690 , w_46691 , w_46692 , w_46693 , w_46694 , w_46695 , 
		w_46696 , w_46697 , w_46698 , w_46699 , w_46700 , w_46701 , w_46702 , w_46703 , w_46704 , w_46705 , 
		w_46706 , w_46707 , w_46708 , w_46709 , w_46710 , w_46711 , w_46712 , w_46713 , w_46714 , w_46715 , 
		w_46716 , w_46717 , w_46718 , w_46719 , w_46720 , w_46721 , w_46722 , w_46723 , w_46724 , w_46725 , 
		w_46726 , w_46727 , w_46728 , w_46729 , w_46730 , w_46731 , w_46732 , w_46733 , w_46734 , w_46735 , 
		w_46736 , w_46737 , w_46738 , w_46739 , w_46740 , w_46741 , w_46742 , w_46743 , w_46744 , w_46745 , 
		w_46746 , w_46747 , w_46748 , w_46749 , w_46750 , w_46751 , w_46752 , w_46753 , w_46754 , w_46755 , 
		w_46756 , w_46757 , w_46758 , w_46759 , w_46760 , w_46761 , w_46762 , w_46763 , w_46764 , w_46765 , 
		w_46766 , w_46767 , w_46768 , w_46769 , w_46770 , w_46771 , w_46772 , w_46773 , w_46774 , w_46775 , 
		w_46776 , w_46777 , w_46778 , w_46779 , w_46780 , w_46781 , w_46782 , w_46783 , w_46784 , w_46785 , 
		w_46786 , w_46787 , w_46788 , w_46789 , w_46790 , w_46791 , w_46792 , w_46793 , w_46794 , w_46795 , 
		w_46796 , w_46797 , w_46798 , w_46799 , w_46800 , w_46801 , w_46802 , w_46803 , w_46804 , w_46805 , 
		w_46806 , w_46807 , w_46808 , w_46809 , w_46810 , w_46811 , w_46812 , w_46813 , w_46814 , w_46815 , 
		w_46816 , w_46817 , w_46818 , w_46819 , w_46820 , w_46821 , w_46822 , w_46823 , w_46824 , w_46825 , 
		w_46826 , w_46827 , w_46828 , w_46829 , w_46830 , w_46831 , w_46832 , w_46833 , w_46834 , w_46835 , 
		w_46836 , w_46837 , w_46838 , w_46839 , w_46840 , w_46841 , w_46842 , w_46843 , w_46844 , w_46845 , 
		w_46846 , w_46847 , w_46848 , w_46849 , w_46850 , w_46851 , w_46852 , w_46853 , w_46854 , w_46855 , 
		w_46856 , w_46857 , w_46858 , w_46859 , w_46860 , w_46861 , w_46862 , w_46863 , w_46864 , w_46865 , 
		w_46866 , w_46867 , w_46868 , w_46869 , w_46870 , w_46871 , w_46872 , w_46873 , w_46874 , w_46875 , 
		w_46876 , w_46877 , w_46878 , w_46879 , w_46880 , w_46881 , w_46882 , w_46883 , w_46884 , w_46885 , 
		w_46886 , w_46887 , w_46888 , w_46889 , w_46890 , w_46891 , w_46892 , w_46893 , w_46894 , w_46895 , 
		w_46896 , w_46897 , w_46898 , w_46899 , w_46900 , w_46901 , w_46902 , w_46903 , w_46904 , w_46905 , 
		w_46906 , w_46907 , w_46908 , w_46909 , w_46910 , w_46911 , w_46912 , w_46913 , w_46914 , w_46915 , 
		w_46916 , w_46917 , w_46918 , w_46919 , w_46920 , w_46921 , w_46922 , w_46923 , w_46924 , w_46925 , 
		w_46926 , w_46927 , w_46928 , w_46929 , w_46930 , w_46931 , w_46932 , w_46933 , w_46934 , w_46935 , 
		w_46936 , w_46937 , w_46938 , w_46939 , w_46940 , w_46941 , w_46942 , w_46943 , w_46944 , w_46945 , 
		w_46946 , w_46947 , w_46948 , w_46949 , w_46950 , w_46951 , w_46952 , w_46953 , w_46954 , w_46955 , 
		w_46956 , w_46957 , w_46958 , w_46959 , w_46960 , w_46961 , w_46962 , w_46963 , w_46964 , w_46965 , 
		w_46966 , w_46967 , w_46968 , w_46969 , w_46970 , w_46971 , w_46972 , w_46973 , w_46974 , w_46975 , 
		w_46976 , w_46977 , w_46978 , w_46979 , w_46980 , w_46981 , w_46982 , w_46983 , w_46984 , w_46985 , 
		w_46986 , w_46987 , w_46988 , w_46989 , w_46990 , w_46991 , w_46992 , w_46993 , w_46994 , w_46995 , 
		w_46996 , w_46997 , w_46998 , w_46999 , w_47000 , w_47001 , w_47002 , w_47003 , w_47004 , w_47005 , 
		w_47006 , w_47007 , w_47008 , w_47009 , w_47010 , w_47011 , w_47012 , w_47013 , w_47014 , w_47015 , 
		w_47016 , w_47017 , w_47018 , w_47019 , w_47020 , w_47021 , w_47022 , w_47023 , w_47024 , w_47025 , 
		w_47026 , w_47027 , w_47028 , w_47029 , w_47030 , w_47031 , w_47032 , w_47033 , w_47034 , w_47035 , 
		w_47036 , w_47037 , w_47038 , w_47039 , w_47040 , w_47041 , w_47042 , w_47043 , w_47044 , w_47045 , 
		w_47046 , w_47047 , w_47048 , w_47049 , w_47050 , w_47051 , w_47052 , w_47053 , w_47054 , w_47055 , 
		w_47056 , w_47057 , w_47058 , w_47059 , w_47060 , w_47061 , w_47062 , w_47063 , w_47064 , w_47065 , 
		w_47066 , w_47067 , w_47068 , w_47069 , w_47070 , w_47071 , w_47072 , w_47073 , w_47074 , w_47075 , 
		w_47076 , w_47077 , w_47078 , w_47079 , w_47080 , w_47081 , w_47082 , w_47083 , w_47084 , w_47085 , 
		w_47086 , w_47087 , w_47088 , w_47089 , w_47090 , w_47091 , w_47092 , w_47093 , w_47094 , w_47095 , 
		w_47096 , w_47097 , w_47098 , w_47099 , w_47100 , w_47101 , w_47102 , w_47103 , w_47104 , w_47105 , 
		w_47106 , w_47107 , w_47108 , w_47109 , w_47110 , w_47111 , w_47112 , w_47113 , w_47114 , w_47115 , 
		w_47116 , w_47117 , w_47118 , w_47119 , w_47120 , w_47121 , w_47122 , w_47123 , w_47124 , w_47125 , 
		w_47126 , w_47127 , w_47128 , w_47129 , w_47130 , w_47131 , w_47132 , w_47133 , w_47134 , w_47135 , 
		w_47136 , w_47137 , w_47138 , w_47139 , w_47140 , w_47141 , w_47142 , w_47143 , w_47144 , w_47145 , 
		w_47146 , w_47147 , w_47148 , w_47149 , w_47150 , w_47151 , w_47152 , w_47153 , w_47154 , w_47155 , 
		w_47156 , w_47157 , w_47158 , w_47159 , w_47160 , w_47161 , w_47162 , w_47163 , w_47164 , w_47165 , 
		w_47166 , w_47167 , w_47168 , w_47169 , w_47170 , w_47171 , w_47172 , w_47173 , w_47174 , w_47175 , 
		w_47176 , w_47177 , w_47178 , w_47179 , w_47180 , w_47181 , w_47182 , w_47183 , w_47184 , w_47185 , 
		w_47186 , w_47187 , w_47188 , w_47189 , w_47190 , w_47191 , w_47192 , w_47193 , w_47194 , w_47195 , 
		w_47196 , w_47197 , w_47198 , w_47199 , w_47200 , w_47201 , w_47202 , w_47203 , w_47204 , w_47205 , 
		w_47206 , w_47207 , w_47208 , w_47209 , w_47210 , w_47211 , w_47212 , w_47213 , w_47214 , w_47215 , 
		w_47216 , w_47217 , w_47218 , w_47219 , w_47220 , w_47221 , w_47222 , w_47223 , w_47224 , w_47225 , 
		w_47226 , w_47227 , w_47228 , w_47229 , w_47230 , w_47231 , w_47232 , w_47233 , w_47234 , w_47235 , 
		w_47236 , w_47237 , w_47238 , w_47239 , w_47240 , w_47241 , w_47242 , w_47243 , w_47244 , w_47245 , 
		w_47246 , w_47247 , w_47248 , w_47249 , w_47250 , w_47251 , w_47252 , w_47253 , w_47254 , w_47255 , 
		w_47256 , w_47257 , w_47258 , w_47259 , w_47260 , w_47261 , w_47262 , w_47263 , w_47264 , w_47265 , 
		w_47266 , w_47267 , w_47268 , w_47269 , w_47270 , w_47271 , w_47272 , w_47273 , w_47274 , w_47275 , 
		w_47276 , w_47277 , w_47278 , w_47279 , w_47280 , w_47281 , w_47282 , w_47283 , w_47284 , w_47285 , 
		w_47286 , w_47287 , w_47288 , w_47289 , w_47290 , w_47291 , w_47292 , w_47293 , w_47294 , w_47295 , 
		w_47296 , w_47297 , w_47298 , w_47299 , w_47300 , w_47301 , w_47302 , w_47303 , w_47304 , w_47305 , 
		w_47306 , w_47307 , w_47308 , w_47309 , w_47310 , w_47311 , w_47312 , w_47313 , w_47314 , w_47315 , 
		w_47316 , w_47317 , w_47318 , w_47319 , w_47320 , w_47321 , w_47322 , w_47323 , w_47324 , w_47325 , 
		w_47326 , w_47327 , w_47328 , w_47329 , w_47330 , w_47331 , w_47332 , w_47333 , w_47334 , w_47335 , 
		w_47336 , w_47337 , w_47338 , w_47339 , w_47340 , w_47341 , w_47342 , w_47343 , w_47344 , w_47345 , 
		w_47346 , w_47347 , w_47348 , w_47349 , w_47350 , w_47351 , w_47352 , w_47353 , w_47354 , w_47355 , 
		w_47356 , w_47357 , w_47358 , w_47359 , w_47360 , w_47361 , w_47362 , w_47363 , w_47364 , w_47365 , 
		w_47366 , w_47367 , w_47368 , w_47369 , w_47370 , w_47371 ;
buf ( R_61_85b54e8_b1 , \14014_b1 );
buf ( R_61_85b54e8_b0 , \14014_b0 );
buf ( R_62_85b5590_b1 , \14196_b1 );
buf ( R_62_85b5590_b0 , \14196_b0 );
buf ( R_63_85b5638_b1 , \14286_b1 );
buf ( R_63_85b5638_b0 , \14286_b0 );
buf ( R_64_85b56e0_b1 , \14377_b1 );
buf ( R_64_85b56e0_b0 , \14377_b0 );
buf ( R_65_85b5788_b1 , \14422_b1 );
buf ( R_65_85b5788_b0 , \14422_b0 );
buf ( R_66_85b5830_b1 , \14467_b1 );
buf ( R_66_85b5830_b0 , \14467_b0 );
buf ( R_67_85b58d8_b1 , \14510_b1 );
buf ( R_67_85b58d8_b0 , \14510_b0 );
buf ( R_68_85b5980_b1 , \14553_b1 );
buf ( R_68_85b5980_b0 , \14553_b0 );
buf ( R_69_85b5a28_b1 , \14576_b1 );
buf ( R_69_85b5a28_b0 , \14576_b0 );
buf ( R_6a_85b5ad0_b1 , \14599_b1 );
buf ( R_6a_85b5ad0_b0 , \14599_b0 );
buf ( R_6b_85b5b78_b1 , \14621_b1 );
buf ( R_6b_85b5b78_b0 , \14621_b0 );
buf ( R_6c_85b5c20_b1 , \14643_b1 );
buf ( R_6c_85b5c20_b0 , \14643_b0 );
buf ( R_6d_85b5cc8_b1 , \14665_b1 );
buf ( R_6d_85b5cc8_b0 , \14665_b0 );
buf ( R_6e_85b5d70_b1 , \14687_b1 );
buf ( R_6e_85b5d70_b0 , \14687_b0 );
buf ( R_6f_85b5e18_b1 , \14707_b1 );
buf ( R_6f_85b5e18_b0 , \14707_b0 );
buf ( R_70_85b5ec0_b1 , \14727_b1 );
buf ( R_70_85b5ec0_b0 , \14727_b0 );
buf ( R_71_85b5f68_b1 , \14739_b1 );
buf ( R_71_85b5f68_b0 , \14739_b0 );
buf ( R_72_85b6010_b1 , \14751_b1 );
buf ( R_72_85b6010_b0 , \14751_b0 );
buf ( R_73_85b60b8_b1 , \14763_b1 );
buf ( R_73_85b60b8_b0 , \14763_b0 );
buf ( R_74_85b6160_b1 , \14775_b1 );
buf ( R_74_85b6160_b0 , \14775_b0 );
buf ( R_75_85b6208_b1 , \14787_b1 );
buf ( R_75_85b6208_b0 , \14787_b0 );
buf ( R_76_85b62b0_b1 , \14799_b1 );
buf ( R_76_85b62b0_b0 , \14799_b0 );
buf ( R_77_85b6358_b1 , \14810_b1 );
buf ( R_77_85b6358_b0 , \14810_b0 );
buf ( R_78_85b6400_b1 , \14821_b1 );
buf ( R_78_85b6400_b0 , \14821_b0 );
buf ( R_79_85b64a8_b1 , \14832_b1 );
buf ( R_79_85b64a8_b0 , \14832_b0 );
buf ( R_7a_85b6550_b1 , \14843_b1 );
buf ( R_7a_85b6550_b0 , \14843_b0 );
buf ( R_7b_85b65f8_b1 , \14854_b1 );
buf ( R_7b_85b65f8_b0 , \14854_b0 );
buf ( R_7c_85b66a0_b1 , \14865_b1 );
buf ( R_7c_85b66a0_b0 , \14865_b0 );
buf ( R_7d_85b6748_b1 , \14876_b1 );
buf ( R_7d_85b6748_b0 , \14876_b0 );
buf ( R_7e_85b67f0_b1 , \14887_b1 );
buf ( R_7e_85b67f0_b0 , \14887_b0 );
buf ( R_7f_85b6898_b1 , \14894_b1 );
buf ( R_7f_85b6898_b0 , \14894_b0 );
buf ( R_80_85b6940_b1 , \14901_b1 );
buf ( R_80_85b6940_b0 , \14901_b0 );
buf ( R_81_85b69e8_b1 , \14906_b1 );
buf ( R_81_85b69e8_b0 , \14906_b0 );
buf ( R_82_85b6a90_b1 , \14911_b1 );
buf ( R_82_85b6a90_b0 , \14911_b0 );
buf ( R_83_85b6b38_b1 , \14916_b1 );
buf ( R_83_85b6b38_b0 , \14916_b0 );
buf ( R_84_85b6be0_b1 , \14921_b1 );
buf ( R_84_85b6be0_b0 , \14921_b0 );
buf ( R_85_85b6c88_b1 , \14926_b1 );
buf ( R_85_85b6c88_b0 , \14926_b0 );
buf ( R_86_85b6d30_b1 , \14931_b1 );
buf ( R_86_85b6d30_b0 , \14931_b0 );
buf ( R_87_85b6dd8_b1 , \14936_b1 );
buf ( R_87_85b6dd8_b0 , \14936_b0 );
buf ( R_88_85b6e80_b1 , \14941_b1 );
buf ( R_88_85b6e80_b0 , \14941_b0 );
buf ( R_89_85b6f28_b1 , \14946_b1 );
buf ( R_89_85b6f28_b0 , \14946_b0 );
buf ( R_8a_85b6fd0_b1 , \14951_b1 );
buf ( R_8a_85b6fd0_b0 , \14951_b0 );
buf ( R_8b_85b7078_b1 , \14956_b1 );
buf ( R_8b_85b7078_b0 , \14956_b0 );
buf ( R_8c_85b7120_b1 , \14961_b1 );
buf ( R_8c_85b7120_b0 , \14961_b0 );
buf ( R_8d_85b71c8_b1 , \14966_b1 );
buf ( R_8d_85b71c8_b0 , \14966_b0 );
buf ( R_8e_85b7270_b1 , \14971_b1 );
buf ( R_8e_85b7270_b0 , \14971_b0 );
buf ( R_8f_85b7318_b1 , \14976_b1 );
buf ( R_8f_85b7318_b0 , \14976_b0 );
buf ( R_90_85b73c0_b1 , \14981_b1 );
buf ( R_90_85b73c0_b0 , \14981_b0 );
buf ( R_91_85b7468_b1 , \14986_b1 );
buf ( R_91_85b7468_b0 , \14986_b0 );
buf ( R_92_85b7510_b1 , \14991_b1 );
buf ( R_92_85b7510_b0 , \14991_b0 );
buf ( R_93_85b75b8_b1 , \14996_b1 );
buf ( R_93_85b75b8_b0 , \14996_b0 );
buf ( R_94_85b7660_b1 , \15001_b1 );
buf ( R_94_85b7660_b0 , \15001_b0 );
buf ( R_95_85b7708_b1 , \15006_b1 );
buf ( R_95_85b7708_b0 , \15006_b0 );
buf ( R_96_85b77b0_b1 , \15011_b1 );
buf ( R_96_85b77b0_b0 , \15011_b0 );
buf ( R_97_85b7858_b1 , \15016_b1 );
buf ( R_97_85b7858_b0 , \15016_b0 );
buf ( R_98_85b7900_b1 , \15021_b1 );
buf ( R_98_85b7900_b0 , \15021_b0 );
buf ( R_99_85b79a8_b1 , \15026_b1 );
buf ( R_99_85b79a8_b0 , \15026_b0 );
buf ( R_9a_85b7a50_b1 , \15031_b1 );
buf ( R_9a_85b7a50_b0 , \15031_b0 );
buf ( \159_b1 , RIb4bfa38_65_b1 );
buf ( \159_b0 , RIb4bfa38_65_b0 );
buf ( \160_b1 , RIa167a08_1_b1 );
buf ( \160_b0 , RIa167a08_1_b0 );
buf ( \161_b1 , RIb4ca3e8_33_b1 );
buf ( \161_b0 , RIb4ca3e8_33_b0 );
or ( \162_b1 , \160_b1 , \161_b1 );
xor ( \162_b0 , \160_b0 , w_0 );
not ( w_0 , w_1 );
and ( w_1 , \161_b1 , \161_b0 );
buf ( \163_b1 , RIa167990_2_b1 );
buf ( \163_b0 , RIa167990_2_b0 );
buf ( \164_b1 , RIb4c6c20_34_b1 );
buf ( \164_b0 , RIb4c6c20_34_b0 );
or ( \165_b1 , \163_b1 , \164_b1 );
xor ( \165_b0 , \163_b0 , w_2 );
not ( w_2 , w_3 );
and ( w_3 , \164_b1 , \164_b0 );
or ( \166_b1 , \162_b1 , w_4 );
or ( \166_b0 , \162_b0 , \165_b0 );
not ( \165_b0 , w_5 );
and ( w_5 , w_4 , \165_b1 );
buf ( \167_b1 , RIa167918_3_b1 );
buf ( \167_b0 , RIa167918_3_b0 );
buf ( \168_b1 , RIb4c6ba8_35_b1 );
buf ( \168_b0 , RIb4c6ba8_35_b0 );
or ( \169_b1 , \167_b1 , \168_b1 );
xor ( \169_b0 , \167_b0 , w_6 );
not ( w_6 , w_7 );
and ( w_7 , \168_b1 , \168_b0 );
or ( \170_b1 , \166_b1 , w_8 );
or ( \170_b0 , \166_b0 , \169_b0 );
not ( \169_b0 , w_9 );
and ( w_9 , w_8 , \169_b1 );
buf ( \171_b1 , RIa1678a0_4_b1 );
buf ( \171_b0 , RIa1678a0_4_b0 );
buf ( \172_b1 , RIb4c6b30_36_b1 );
buf ( \172_b0 , RIb4c6b30_36_b0 );
or ( \173_b1 , \171_b1 , \172_b1 );
xor ( \173_b0 , \171_b0 , w_10 );
not ( w_10 , w_11 );
and ( w_11 , \172_b1 , \172_b0 );
or ( \174_b1 , \170_b1 , w_12 );
or ( \174_b0 , \170_b0 , \173_b0 );
not ( \173_b0 , w_13 );
and ( w_13 , w_12 , \173_b1 );
buf ( \175_b1 , RIa167828_5_b1 );
buf ( \175_b0 , RIa167828_5_b0 );
buf ( \176_b1 , RIb4c6ab8_37_b1 );
buf ( \176_b0 , RIb4c6ab8_37_b0 );
or ( \177_b1 , \175_b1 , \176_b1 );
xor ( \177_b0 , \175_b0 , w_14 );
not ( w_14 , w_15 );
and ( w_15 , \176_b1 , \176_b0 );
or ( \178_b1 , \174_b1 , w_16 );
or ( \178_b0 , \174_b0 , \177_b0 );
not ( \177_b0 , w_17 );
and ( w_17 , w_16 , \177_b1 );
buf ( \179_b1 , RIa1677b0_6_b1 );
buf ( \179_b0 , RIa1677b0_6_b0 );
buf ( \180_b1 , RIb4c6a40_38_b1 );
buf ( \180_b0 , RIb4c6a40_38_b0 );
or ( \181_b1 , \179_b1 , \180_b1 );
xor ( \181_b0 , \179_b0 , w_18 );
not ( w_18 , w_19 );
and ( w_19 , \180_b1 , \180_b0 );
or ( \182_b1 , \178_b1 , w_20 );
or ( \182_b0 , \178_b0 , \181_b0 );
not ( \181_b0 , w_21 );
and ( w_21 , w_20 , \181_b1 );
buf ( \183_b1 , RIa167738_7_b1 );
buf ( \183_b0 , RIa167738_7_b0 );
buf ( \184_b1 , RIb4c69c8_39_b1 );
buf ( \184_b0 , RIb4c69c8_39_b0 );
or ( \185_b1 , \183_b1 , \184_b1 );
xor ( \185_b0 , \183_b0 , w_22 );
not ( w_22 , w_23 );
and ( w_23 , \184_b1 , \184_b0 );
or ( \186_b1 , \182_b1 , w_24 );
or ( \186_b0 , \182_b0 , \185_b0 );
not ( \185_b0 , w_25 );
and ( w_25 , w_24 , \185_b1 );
buf ( \187_b1 , RIa1676c0_8_b1 );
buf ( \187_b0 , RIa1676c0_8_b0 );
buf ( \188_b1 , RIb4c6950_40_b1 );
buf ( \188_b0 , RIb4c6950_40_b0 );
or ( \189_b1 , \187_b1 , \188_b1 );
xor ( \189_b0 , \187_b0 , w_26 );
not ( w_26 , w_27 );
and ( w_27 , \188_b1 , \188_b0 );
or ( \190_b1 , \186_b1 , w_28 );
or ( \190_b0 , \186_b0 , \189_b0 );
not ( \189_b0 , w_29 );
and ( w_29 , w_28 , \189_b1 );
buf ( \191_b1 , RIa167648_9_b1 );
buf ( \191_b0 , RIa167648_9_b0 );
buf ( \192_b1 , RIb4c68d8_41_b1 );
buf ( \192_b0 , RIb4c68d8_41_b0 );
or ( \193_b1 , \191_b1 , \192_b1 );
xor ( \193_b0 , \191_b0 , w_30 );
not ( w_30 , w_31 );
and ( w_31 , \192_b1 , \192_b0 );
or ( \194_b1 , \190_b1 , w_32 );
or ( \194_b0 , \190_b0 , \193_b0 );
not ( \193_b0 , w_33 );
and ( w_33 , w_32 , \193_b1 );
buf ( \195_b1 , RIa1675d0_10_b1 );
buf ( \195_b0 , RIa1675d0_10_b0 );
buf ( \196_b1 , RIb4c6860_42_b1 );
buf ( \196_b0 , RIb4c6860_42_b0 );
or ( \197_b1 , \195_b1 , \196_b1 );
xor ( \197_b0 , \195_b0 , w_34 );
not ( w_34 , w_35 );
and ( w_35 , \196_b1 , \196_b0 );
or ( \198_b1 , \194_b1 , w_36 );
or ( \198_b0 , \194_b0 , \197_b0 );
not ( \197_b0 , w_37 );
and ( w_37 , w_36 , \197_b1 );
buf ( \199_b1 , RIa167558_11_b1 );
buf ( \199_b0 , RIa167558_11_b0 );
buf ( \200_b1 , RIb4c67e8_43_b1 );
buf ( \200_b0 , RIb4c67e8_43_b0 );
or ( \201_b1 , \199_b1 , \200_b1 );
xor ( \201_b0 , \199_b0 , w_38 );
not ( w_38 , w_39 );
and ( w_39 , \200_b1 , \200_b0 );
or ( \202_b1 , \198_b1 , w_40 );
or ( \202_b0 , \198_b0 , \201_b0 );
not ( \201_b0 , w_41 );
and ( w_41 , w_40 , \201_b1 );
buf ( \203_b1 , RIa1674e0_12_b1 );
buf ( \203_b0 , RIa1674e0_12_b0 );
buf ( \204_b1 , RIb4c6770_44_b1 );
buf ( \204_b0 , RIb4c6770_44_b0 );
or ( \205_b1 , \203_b1 , \204_b1 );
xor ( \205_b0 , \203_b0 , w_42 );
not ( w_42 , w_43 );
and ( w_43 , \204_b1 , \204_b0 );
or ( \206_b1 , \202_b1 , w_44 );
or ( \206_b0 , \202_b0 , \205_b0 );
not ( \205_b0 , w_45 );
and ( w_45 , w_44 , \205_b1 );
buf ( \207_b1 , RIa167468_13_b1 );
buf ( \207_b0 , RIa167468_13_b0 );
buf ( \208_b1 , RIb4c3368_45_b1 );
buf ( \208_b0 , RIb4c3368_45_b0 );
or ( \209_b1 , \207_b1 , \208_b1 );
xor ( \209_b0 , \207_b0 , w_46 );
not ( w_46 , w_47 );
and ( w_47 , \208_b1 , \208_b0 );
or ( \210_b1 , \206_b1 , w_48 );
or ( \210_b0 , \206_b0 , \209_b0 );
not ( \209_b0 , w_49 );
and ( w_49 , w_48 , \209_b1 );
buf ( \211_b1 , RIa1673f0_14_b1 );
buf ( \211_b0 , RIa1673f0_14_b0 );
buf ( \212_b1 , RIb4c32f0_46_b1 );
buf ( \212_b0 , RIb4c32f0_46_b0 );
or ( \213_b1 , \211_b1 , \212_b1 );
xor ( \213_b0 , \211_b0 , w_50 );
not ( w_50 , w_51 );
and ( w_51 , \212_b1 , \212_b0 );
or ( \214_b1 , \210_b1 , w_52 );
or ( \214_b0 , \210_b0 , \213_b0 );
not ( \213_b0 , w_53 );
and ( w_53 , w_52 , \213_b1 );
buf ( \215_b1 , RIa167378_15_b1 );
buf ( \215_b0 , RIa167378_15_b0 );
buf ( \216_b1 , RIb4c3278_47_b1 );
buf ( \216_b0 , RIb4c3278_47_b0 );
or ( \217_b1 , \215_b1 , \216_b1 );
xor ( \217_b0 , \215_b0 , w_54 );
not ( w_54 , w_55 );
and ( w_55 , \216_b1 , \216_b0 );
or ( \218_b1 , \214_b1 , w_56 );
or ( \218_b0 , \214_b0 , \217_b0 );
not ( \217_b0 , w_57 );
and ( w_57 , w_56 , \217_b1 );
buf ( \219_b1 , RIa167300_16_b1 );
buf ( \219_b0 , RIa167300_16_b0 );
buf ( \220_b1 , RIb4c3200_48_b1 );
buf ( \220_b0 , RIb4c3200_48_b0 );
or ( \221_b1 , \219_b1 , \220_b1 );
xor ( \221_b0 , \219_b0 , w_58 );
not ( w_58 , w_59 );
and ( w_59 , \220_b1 , \220_b0 );
or ( \222_b1 , \218_b1 , w_60 );
or ( \222_b0 , \218_b0 , \221_b0 );
not ( \221_b0 , w_61 );
and ( w_61 , w_60 , \221_b1 );
buf ( \223_b1 , RIa167288_17_b1 );
buf ( \223_b0 , RIa167288_17_b0 );
buf ( \224_b1 , RIb4c3188_49_b1 );
buf ( \224_b0 , RIb4c3188_49_b0 );
or ( \225_b1 , \223_b1 , \224_b1 );
xor ( \225_b0 , \223_b0 , w_62 );
not ( w_62 , w_63 );
and ( w_63 , \224_b1 , \224_b0 );
or ( \226_b1 , \222_b1 , w_64 );
or ( \226_b0 , \222_b0 , \225_b0 );
not ( \225_b0 , w_65 );
and ( w_65 , w_64 , \225_b1 );
buf ( \227_b1 , RIa167210_18_b1 );
buf ( \227_b0 , RIa167210_18_b0 );
buf ( \228_b1 , RIb4c3110_50_b1 );
buf ( \228_b0 , RIb4c3110_50_b0 );
or ( \229_b1 , \227_b1 , \228_b1 );
xor ( \229_b0 , \227_b0 , w_66 );
not ( w_66 , w_67 );
and ( w_67 , \228_b1 , \228_b0 );
or ( \230_b1 , \226_b1 , w_68 );
or ( \230_b0 , \226_b0 , \229_b0 );
not ( \229_b0 , w_69 );
and ( w_69 , w_68 , \229_b1 );
buf ( \231_b1 , RIa167198_19_b1 );
buf ( \231_b0 , RIa167198_19_b0 );
buf ( \232_b1 , RIb4c3098_51_b1 );
buf ( \232_b0 , RIb4c3098_51_b0 );
or ( \233_b1 , \231_b1 , \232_b1 );
xor ( \233_b0 , \231_b0 , w_70 );
not ( w_70 , w_71 );
and ( w_71 , \232_b1 , \232_b0 );
or ( \234_b1 , \230_b1 , w_72 );
or ( \234_b0 , \230_b0 , \233_b0 );
not ( \233_b0 , w_73 );
and ( w_73 , w_72 , \233_b1 );
buf ( \235_b1 , RIa167120_20_b1 );
buf ( \235_b0 , RIa167120_20_b0 );
buf ( \236_b1 , RIb4c3020_52_b1 );
buf ( \236_b0 , RIb4c3020_52_b0 );
or ( \237_b1 , \235_b1 , \236_b1 );
xor ( \237_b0 , \235_b0 , w_74 );
not ( w_74 , w_75 );
and ( w_75 , \236_b1 , \236_b0 );
or ( \238_b1 , \234_b1 , w_76 );
or ( \238_b0 , \234_b0 , \237_b0 );
not ( \237_b0 , w_77 );
and ( w_77 , w_76 , \237_b1 );
buf ( \239_b1 , RIa1670a8_21_b1 );
buf ( \239_b0 , RIa1670a8_21_b0 );
buf ( \240_b1 , RIb4c2fa8_53_b1 );
buf ( \240_b0 , RIb4c2fa8_53_b0 );
or ( \241_b1 , \239_b1 , \240_b1 );
xor ( \241_b0 , \239_b0 , w_78 );
not ( w_78 , w_79 );
and ( w_79 , \240_b1 , \240_b0 );
or ( \242_b1 , \238_b1 , w_80 );
or ( \242_b0 , \238_b0 , \241_b0 );
not ( \241_b0 , w_81 );
and ( w_81 , w_80 , \241_b1 );
buf ( \243_b1 , RIa167030_22_b1 );
buf ( \243_b0 , RIa167030_22_b0 );
buf ( \244_b1 , RIb4c2f30_54_b1 );
buf ( \244_b0 , RIb4c2f30_54_b0 );
or ( \245_b1 , \243_b1 , \244_b1 );
xor ( \245_b0 , \243_b0 , w_82 );
not ( w_82 , w_83 );
and ( w_83 , \244_b1 , \244_b0 );
or ( \246_b1 , \242_b1 , w_84 );
or ( \246_b0 , \242_b0 , \245_b0 );
not ( \245_b0 , w_85 );
and ( w_85 , w_84 , \245_b1 );
buf ( \247_b1 , RIa166fb8_23_b1 );
buf ( \247_b0 , RIa166fb8_23_b0 );
buf ( \248_b1 , RIb4c2eb8_55_b1 );
buf ( \248_b0 , RIb4c2eb8_55_b0 );
or ( \249_b1 , \247_b1 , \248_b1 );
xor ( \249_b0 , \247_b0 , w_86 );
not ( w_86 , w_87 );
and ( w_87 , \248_b1 , \248_b0 );
or ( \250_b1 , \246_b1 , w_88 );
or ( \250_b0 , \246_b0 , \249_b0 );
not ( \249_b0 , w_89 );
and ( w_89 , w_88 , \249_b1 );
buf ( \251_b1 , RIa166f40_24_b1 );
buf ( \251_b0 , RIa166f40_24_b0 );
buf ( \252_b1 , RIb4c2e40_56_b1 );
buf ( \252_b0 , RIb4c2e40_56_b0 );
or ( \253_b1 , \251_b1 , \252_b1 );
xor ( \253_b0 , \251_b0 , w_90 );
not ( w_90 , w_91 );
and ( w_91 , \252_b1 , \252_b0 );
or ( \254_b1 , \250_b1 , w_92 );
or ( \254_b0 , \250_b0 , \253_b0 );
not ( \253_b0 , w_93 );
and ( w_93 , w_92 , \253_b1 );
buf ( \255_b1 , RIa166ec8_25_b1 );
buf ( \255_b0 , RIa166ec8_25_b0 );
buf ( \256_b1 , RIb4c2dc8_57_b1 );
buf ( \256_b0 , RIb4c2dc8_57_b0 );
or ( \257_b1 , \255_b1 , \256_b1 );
xor ( \257_b0 , \255_b0 , w_94 );
not ( w_94 , w_95 );
and ( w_95 , \256_b1 , \256_b0 );
or ( \258_b1 , \254_b1 , w_96 );
or ( \258_b0 , \254_b0 , \257_b0 );
not ( \257_b0 , w_97 );
and ( w_97 , w_96 , \257_b1 );
buf ( \259_b1 , RIa166e50_26_b1 );
buf ( \259_b0 , RIa166e50_26_b0 );
buf ( \260_b1 , RIb4c2d50_58_b1 );
buf ( \260_b0 , RIb4c2d50_58_b0 );
or ( \261_b1 , \259_b1 , \260_b1 );
xor ( \261_b0 , \259_b0 , w_98 );
not ( w_98 , w_99 );
and ( w_99 , \260_b1 , \260_b0 );
or ( \262_b1 , \258_b1 , w_100 );
or ( \262_b0 , \258_b0 , \261_b0 );
not ( \261_b0 , w_101 );
and ( w_101 , w_100 , \261_b1 );
buf ( \263_b1 , RIa166dd8_27_b1 );
buf ( \263_b0 , RIa166dd8_27_b0 );
buf ( \264_b1 , RIb4c2cd8_59_b1 );
buf ( \264_b0 , RIb4c2cd8_59_b0 );
or ( \265_b1 , \263_b1 , \264_b1 );
xor ( \265_b0 , \263_b0 , w_102 );
not ( w_102 , w_103 );
and ( w_103 , \264_b1 , \264_b0 );
or ( \266_b1 , \262_b1 , w_104 );
or ( \266_b0 , \262_b0 , \265_b0 );
not ( \265_b0 , w_105 );
and ( w_105 , w_104 , \265_b1 );
buf ( \267_b1 , RIa166d60_28_b1 );
buf ( \267_b0 , RIa166d60_28_b0 );
buf ( \268_b1 , RIb4c2c60_60_b1 );
buf ( \268_b0 , RIb4c2c60_60_b0 );
or ( \269_b1 , \267_b1 , \268_b1 );
xor ( \269_b0 , \267_b0 , w_106 );
not ( w_106 , w_107 );
and ( w_107 , \268_b1 , \268_b0 );
or ( \270_b1 , \266_b1 , w_108 );
or ( \270_b0 , \266_b0 , \269_b0 );
not ( \269_b0 , w_109 );
and ( w_109 , w_108 , \269_b1 );
buf ( \271_b1 , RIa166ce8_29_b1 );
buf ( \271_b0 , RIa166ce8_29_b0 );
buf ( \272_b1 , RIb4c2be8_61_b1 );
buf ( \272_b0 , RIb4c2be8_61_b0 );
or ( \273_b1 , \271_b1 , \272_b1 );
xor ( \273_b0 , \271_b0 , w_110 );
not ( w_110 , w_111 );
and ( w_111 , \272_b1 , \272_b0 );
or ( \274_b1 , \270_b1 , w_112 );
or ( \274_b0 , \270_b0 , \273_b0 );
not ( \273_b0 , w_113 );
and ( w_113 , w_112 , \273_b1 );
buf ( \275_b1 , RIa166c70_30_b1 );
buf ( \275_b0 , RIa166c70_30_b0 );
buf ( \276_b1 , RIb4c2b70_62_b1 );
buf ( \276_b0 , RIb4c2b70_62_b0 );
or ( \277_b1 , \275_b1 , \276_b1 );
xor ( \277_b0 , \275_b0 , w_114 );
not ( w_114 , w_115 );
and ( w_115 , \276_b1 , \276_b0 );
or ( \278_b1 , \274_b1 , w_116 );
or ( \278_b0 , \274_b0 , \277_b0 );
not ( \277_b0 , w_117 );
and ( w_117 , w_116 , \277_b1 );
buf ( \279_b1 , RIb4ca4d8_31_b1 );
buf ( \279_b0 , RIb4ca4d8_31_b0 );
buf ( \280_b1 , RIb4c2af8_63_b1 );
buf ( \280_b0 , RIb4c2af8_63_b0 );
or ( \281_b1 , \279_b1 , \280_b1 );
xor ( \281_b0 , \279_b0 , w_118 );
not ( w_118 , w_119 );
and ( w_119 , \280_b1 , \280_b0 );
or ( \282_b1 , \278_b1 , w_120 );
or ( \282_b0 , \278_b0 , \281_b0 );
not ( \281_b0 , w_121 );
and ( w_121 , w_120 , \281_b1 );
buf ( \283_b1 , RIb4ca460_32_b1 );
buf ( \283_b0 , RIb4ca460_32_b0 );
buf ( \284_b1 , RIb4bfab0_64_b1 );
buf ( \284_b0 , RIb4bfab0_64_b0 );
or ( \285_b1 , \283_b1 , \284_b1 );
xor ( \285_b0 , \283_b0 , w_122 );
not ( w_122 , w_123 );
and ( w_123 , \284_b1 , \284_b0 );
or ( \286_b1 , \282_b1 , w_124 );
or ( \286_b0 , \282_b0 , \285_b0 );
not ( \285_b0 , w_125 );
and ( w_125 , w_124 , \285_b1 );
buf ( \287_b1 , \286_b1 );
buf ( \287_b0 , \286_b0 );
buf ( \288_b1 , \287_b1 );
not ( \288_b1 , w_126 );
not ( \288_b0 , w_127 );
and ( w_126 , w_127 , \287_b0 );
and ( \289_nR13d_b1 , RIb4c69c8_39_b1 , w_128 );
xor ( w_128 , RIb4c69c8_39_b0 , \288_b1 );
not ( \288_b1 , w_129 );
and ( \289_nR13d_b0 , w_129 , \288_b0 );
buf ( \290_b1 , \289_nR13d_b1 );
buf ( \290_b0 , \289_nR13d_b0 );
and ( \291_nR13c_b1 , RIb4c6950_40_b1 , w_130 );
xor ( w_130 , RIb4c6950_40_b0 , \288_b1 );
not ( \288_b1 , w_131 );
and ( \291_nR13c_b0 , w_131 , \288_b0 );
buf ( \292_b1 , \291_nR13c_b1 );
buf ( \292_b0 , \291_nR13c_b0 );
or ( \293_b1 , \290_b1 , \292_b1 );
xor ( \293_b0 , \290_b0 , w_132 );
not ( w_132 , w_133 );
and ( w_133 , \292_b1 , \292_b0 );
and ( \294_nR13b_b1 , RIb4c68d8_41_b1 , w_134 );
xor ( w_134 , RIb4c68d8_41_b0 , \288_b1 );
not ( \288_b1 , w_135 );
and ( \294_nR13b_b0 , w_135 , \288_b0 );
buf ( \295_b1 , \294_nR13b_b1 );
buf ( \295_b0 , \294_nR13b_b0 );
or ( \296_b1 , \292_b1 , \295_b1 );
xor ( \296_b0 , \292_b0 , w_136 );
not ( w_136 , w_137 );
and ( w_137 , \295_b1 , \295_b0 );
buf ( \297_b1 , \296_b1 );
not ( \297_b1 , w_138 );
not ( \297_b0 , w_139 );
and ( w_138 , w_139 , \296_b0 );
or ( \298_b1 , \293_b1 , \297_b1 );
not ( \297_b1 , w_140 );
and ( \298_b0 , \293_b0 , w_141 );
and ( w_140 , w_141 , \297_b0 );
or ( \299_b1 , \159_b1 , \298_b1 );
not ( \298_b1 , w_142 );
and ( \299_b0 , \159_b0 , w_143 );
and ( w_142 , w_143 , \298_b0 );
buf ( \300_b1 , \299_b1 );
not ( \300_b1 , w_144 );
not ( \300_b0 , w_145 );
and ( w_144 , w_145 , \299_b0 );
or ( \301_b1 , \292_b1 , \295_b1 );
not ( \295_b1 , w_146 );
and ( \301_b0 , \292_b0 , w_147 );
and ( w_146 , w_147 , \295_b0 );
buf ( \302_b1 , \301_b1 );
not ( \302_b1 , w_148 );
not ( \302_b0 , w_149 );
and ( w_148 , w_149 , \301_b0 );
or ( \303_b1 , \290_b1 , \302_b1 );
not ( \302_b1 , w_150 );
and ( \303_b0 , \290_b0 , w_151 );
and ( w_150 , w_151 , \302_b0 );
or ( \304_b1 , \300_b1 , w_152 );
xor ( \304_b0 , \300_b0 , w_154 );
not ( w_154 , w_155 );
and ( w_155 , w_152 , w_153 );
buf ( w_152 , \303_b1 );
not ( w_152 , w_156 );
not ( w_153 , w_157 );
and ( w_156 , w_157 , \303_b0 );
buf ( \305_b1 , RIb4bf948_67_b1 );
buf ( \305_b0 , RIb4bf948_67_b0 );
and ( \306_nR13f_b1 , RIb4c6ab8_37_b1 , w_158 );
xor ( w_158 , RIb4c6ab8_37_b0 , \288_b1 );
not ( \288_b1 , w_159 );
and ( \306_nR13f_b0 , w_159 , \288_b0 );
buf ( \307_b1 , \306_nR13f_b1 );
buf ( \307_b0 , \306_nR13f_b0 );
and ( \308_nR13e_b1 , RIb4c6a40_38_b1 , w_160 );
xor ( w_160 , RIb4c6a40_38_b0 , \288_b1 );
not ( \288_b1 , w_161 );
and ( \308_nR13e_b0 , w_161 , \288_b0 );
buf ( \309_b1 , \308_nR13e_b1 );
buf ( \309_b0 , \308_nR13e_b0 );
or ( \310_b1 , \307_b1 , \309_b1 );
xor ( \310_b0 , \307_b0 , w_162 );
not ( w_162 , w_163 );
and ( w_163 , \309_b1 , \309_b0 );
or ( \311_b1 , \309_b1 , \290_b1 );
xor ( \311_b0 , \309_b0 , w_164 );
not ( w_164 , w_165 );
and ( w_165 , \290_b1 , \290_b0 );
buf ( \312_b1 , \311_b1 );
not ( \312_b1 , w_166 );
not ( \312_b0 , w_167 );
and ( w_166 , w_167 , \311_b0 );
or ( \313_b1 , \310_b1 , \312_b1 );
not ( \312_b1 , w_168 );
and ( \313_b0 , \310_b0 , w_169 );
and ( w_168 , w_169 , \312_b0 );
or ( \314_b1 , \305_b1 , \313_b1 );
not ( \313_b1 , w_170 );
and ( \314_b0 , \305_b0 , w_171 );
and ( w_170 , w_171 , \313_b0 );
buf ( \315_b1 , RIb4bf9c0_66_b1 );
buf ( \315_b0 , RIb4bf9c0_66_b0 );
or ( \316_b1 , \315_b1 , \311_b1 );
not ( \311_b1 , w_172 );
and ( \316_b0 , \315_b0 , w_173 );
and ( w_172 , w_173 , \311_b0 );
or ( \317_b1 , \314_b1 , w_175 );
not ( w_175 , w_176 );
and ( \317_b0 , \314_b0 , w_177 );
and ( w_176 ,  , w_177 );
buf ( w_175 , \316_b1 );
not ( w_175 , w_178 );
not (  , w_179 );
and ( w_178 , w_179 , \316_b0 );
or ( \318_b1 , \309_b1 , \290_b1 );
not ( \290_b1 , w_180 );
and ( \318_b0 , \309_b0 , w_181 );
and ( w_180 , w_181 , \290_b0 );
buf ( \319_b1 , \318_b1 );
not ( \319_b1 , w_182 );
not ( \319_b0 , w_183 );
and ( w_182 , w_183 , \318_b0 );
or ( \320_b1 , \307_b1 , \319_b1 );
not ( \319_b1 , w_184 );
and ( \320_b0 , \307_b0 , w_185 );
and ( w_184 , w_185 , \319_b0 );
or ( \321_b1 , \317_b1 , w_186 );
xor ( \321_b0 , \317_b0 , w_188 );
not ( w_188 , w_189 );
and ( w_189 , w_186 , w_187 );
buf ( w_186 , \320_b1 );
not ( w_186 , w_190 );
not ( w_187 , w_191 );
and ( w_190 , w_191 , \320_b0 );
or ( \322_b1 , \304_b1 , \321_b1 );
not ( \321_b1 , w_192 );
and ( \322_b0 , \304_b0 , w_193 );
and ( w_192 , w_193 , \321_b0 );
buf ( \323_b1 , RIb4bf858_69_b1 );
buf ( \323_b0 , RIb4bf858_69_b0 );
and ( \324_nR141_b1 , RIb4c6ba8_35_b1 , w_194 );
xor ( w_194 , RIb4c6ba8_35_b0 , \288_b1 );
not ( \288_b1 , w_195 );
and ( \324_nR141_b0 , w_195 , \288_b0 );
buf ( \325_b1 , \324_nR141_b1 );
buf ( \325_b0 , \324_nR141_b0 );
and ( \326_nR140_b1 , RIb4c6b30_36_b1 , w_196 );
xor ( w_196 , RIb4c6b30_36_b0 , \288_b1 );
not ( \288_b1 , w_197 );
and ( \326_nR140_b0 , w_197 , \288_b0 );
buf ( \327_b1 , \326_nR140_b1 );
buf ( \327_b0 , \326_nR140_b0 );
or ( \328_b1 , \325_b1 , \327_b1 );
xor ( \328_b0 , \325_b0 , w_198 );
not ( w_198 , w_199 );
and ( w_199 , \327_b1 , \327_b0 );
or ( \329_b1 , \327_b1 , \307_b1 );
xor ( \329_b0 , \327_b0 , w_200 );
not ( w_200 , w_201 );
and ( w_201 , \307_b1 , \307_b0 );
buf ( \330_b1 , \329_b1 );
not ( \330_b1 , w_202 );
not ( \330_b0 , w_203 );
and ( w_202 , w_203 , \329_b0 );
or ( \331_b1 , \328_b1 , \330_b1 );
not ( \330_b1 , w_204 );
and ( \331_b0 , \328_b0 , w_205 );
and ( w_204 , w_205 , \330_b0 );
or ( \332_b1 , \323_b1 , \331_b1 );
not ( \331_b1 , w_206 );
and ( \332_b0 , \323_b0 , w_207 );
and ( w_206 , w_207 , \331_b0 );
buf ( \333_b1 , RIb4bf8d0_68_b1 );
buf ( \333_b0 , RIb4bf8d0_68_b0 );
or ( \334_b1 , \333_b1 , \329_b1 );
not ( \329_b1 , w_208 );
and ( \334_b0 , \333_b0 , w_209 );
and ( w_208 , w_209 , \329_b0 );
or ( \335_b1 , \332_b1 , w_211 );
not ( w_211 , w_212 );
and ( \335_b0 , \332_b0 , w_213 );
and ( w_212 ,  , w_213 );
buf ( w_211 , \334_b1 );
not ( w_211 , w_214 );
not (  , w_215 );
and ( w_214 , w_215 , \334_b0 );
or ( \336_b1 , \327_b1 , \307_b1 );
not ( \307_b1 , w_216 );
and ( \336_b0 , \327_b0 , w_217 );
and ( w_216 , w_217 , \307_b0 );
buf ( \337_b1 , \336_b1 );
not ( \337_b1 , w_218 );
not ( \337_b0 , w_219 );
and ( w_218 , w_219 , \336_b0 );
or ( \338_b1 , \325_b1 , \337_b1 );
not ( \337_b1 , w_220 );
and ( \338_b0 , \325_b0 , w_221 );
and ( w_220 , w_221 , \337_b0 );
or ( \339_b1 , \335_b1 , w_222 );
xor ( \339_b0 , \335_b0 , w_224 );
not ( w_224 , w_225 );
and ( w_225 , w_222 , w_223 );
buf ( w_222 , \338_b1 );
not ( w_222 , w_226 );
not ( w_223 , w_227 );
and ( w_226 , w_227 , \338_b0 );
or ( \340_b1 , \321_b1 , \339_b1 );
not ( \339_b1 , w_228 );
and ( \340_b0 , \321_b0 , w_229 );
and ( w_228 , w_229 , \339_b0 );
or ( \341_b1 , \304_b1 , \339_b1 );
not ( \339_b1 , w_230 );
and ( \341_b0 , \304_b0 , w_231 );
and ( w_230 , w_231 , \339_b0 );
buf ( \343_b1 , RIb4bf768_71_b1 );
buf ( \343_b0 , RIb4bf768_71_b0 );
and ( \344_nR143_b1 , RIb4ca3e8_33_b1 , w_232 );
xor ( w_232 , RIb4ca3e8_33_b0 , \288_b1 );
not ( \288_b1 , w_233 );
and ( \344_nR143_b0 , w_233 , \288_b0 );
buf ( \345_b1 , \344_nR143_b1 );
buf ( \345_b0 , \344_nR143_b0 );
and ( \346_nR142_b1 , RIb4c6c20_34_b1 , w_234 );
xor ( w_234 , RIb4c6c20_34_b0 , \288_b1 );
not ( \288_b1 , w_235 );
and ( \346_nR142_b0 , w_235 , \288_b0 );
buf ( \347_b1 , \346_nR142_b1 );
buf ( \347_b0 , \346_nR142_b0 );
or ( \348_b1 , \345_b1 , \347_b1 );
xor ( \348_b0 , \345_b0 , w_236 );
not ( w_236 , w_237 );
and ( w_237 , \347_b1 , \347_b0 );
or ( \349_b1 , \347_b1 , \325_b1 );
xor ( \349_b0 , \347_b0 , w_238 );
not ( w_238 , w_239 );
and ( w_239 , \325_b1 , \325_b0 );
buf ( \350_b1 , \349_b1 );
not ( \350_b1 , w_240 );
not ( \350_b0 , w_241 );
and ( w_240 , w_241 , \349_b0 );
or ( \351_b1 , \348_b1 , \350_b1 );
not ( \350_b1 , w_242 );
and ( \351_b0 , \348_b0 , w_243 );
and ( w_242 , w_243 , \350_b0 );
or ( \352_b1 , \343_b1 , \351_b1 );
not ( \351_b1 , w_244 );
and ( \352_b0 , \343_b0 , w_245 );
and ( w_244 , w_245 , \351_b0 );
buf ( \353_b1 , RIb4bf7e0_70_b1 );
buf ( \353_b0 , RIb4bf7e0_70_b0 );
or ( \354_b1 , \353_b1 , \349_b1 );
not ( \349_b1 , w_246 );
and ( \354_b0 , \353_b0 , w_247 );
and ( w_246 , w_247 , \349_b0 );
or ( \355_b1 , \352_b1 , w_249 );
not ( w_249 , w_250 );
and ( \355_b0 , \352_b0 , w_251 );
and ( w_250 ,  , w_251 );
buf ( w_249 , \354_b1 );
not ( w_249 , w_252 );
not (  , w_253 );
and ( w_252 , w_253 , \354_b0 );
or ( \356_b1 , \347_b1 , \325_b1 );
not ( \325_b1 , w_254 );
and ( \356_b0 , \347_b0 , w_255 );
and ( w_254 , w_255 , \325_b0 );
buf ( \357_b1 , \356_b1 );
not ( \357_b1 , w_256 );
not ( \357_b0 , w_257 );
and ( w_256 , w_257 , \356_b0 );
or ( \358_b1 , \345_b1 , \357_b1 );
not ( \357_b1 , w_258 );
and ( \358_b0 , \345_b0 , w_259 );
and ( w_258 , w_259 , \357_b0 );
or ( \359_b1 , \355_b1 , w_260 );
xor ( \359_b0 , \355_b0 , w_262 );
not ( w_262 , w_263 );
and ( w_263 , w_260 , w_261 );
buf ( w_260 , \358_b1 );
not ( w_260 , w_264 );
not ( w_261 , w_265 );
and ( w_264 , w_265 , \358_b0 );
buf ( \360_b1 , RIb4bf6f0_72_b1 );
buf ( \360_b0 , RIb4bf6f0_72_b0 );
or ( \361_b1 , \360_b1 , \345_b1 );
not ( \345_b1 , w_266 );
and ( \361_b0 , \360_b0 , w_267 );
and ( w_266 , w_267 , \345_b0 );
or ( \362_b1 , \359_b1 , w_268 );
or ( \362_b0 , \359_b0 , \361_b0 );
not ( \361_b0 , w_269 );
and ( w_269 , w_268 , \361_b1 );
or ( \363_b1 , \342_b1 , \362_b1 );
not ( \362_b1 , w_270 );
and ( \363_b0 , \342_b0 , w_271 );
and ( w_270 , w_271 , \362_b0 );
or ( \364_b1 , \353_b1 , \351_b1 );
not ( \351_b1 , w_272 );
and ( \364_b0 , \353_b0 , w_273 );
and ( w_272 , w_273 , \351_b0 );
or ( \365_b1 , \323_b1 , \349_b1 );
not ( \349_b1 , w_274 );
and ( \365_b0 , \323_b0 , w_275 );
and ( w_274 , w_275 , \349_b0 );
or ( \366_b1 , \364_b1 , w_277 );
not ( w_277 , w_278 );
and ( \366_b0 , \364_b0 , w_279 );
and ( w_278 ,  , w_279 );
buf ( w_277 , \365_b1 );
not ( w_277 , w_280 );
not (  , w_281 );
and ( w_280 , w_281 , \365_b0 );
or ( \367_b1 , \366_b1 , w_282 );
xor ( \367_b0 , \366_b0 , w_284 );
not ( w_284 , w_285 );
and ( w_285 , w_282 , w_283 );
buf ( w_282 , \358_b1 );
not ( w_282 , w_286 );
not ( w_283 , w_287 );
and ( w_286 , w_287 , \358_b0 );
or ( \368_b1 , \362_b1 , \367_b1 );
not ( \367_b1 , w_288 );
and ( \368_b0 , \362_b0 , w_289 );
and ( w_288 , w_289 , \367_b0 );
or ( \369_b1 , \342_b1 , \367_b1 );
not ( \367_b1 , w_290 );
and ( \369_b0 , \342_b0 , w_291 );
and ( w_290 , w_291 , \367_b0 );
or ( \371_b1 , \343_b1 , \345_b1 );
not ( \345_b1 , w_292 );
and ( \371_b0 , \343_b0 , w_293 );
and ( w_292 , w_293 , \345_b0 );
buf ( \372_b1 , \303_b1 );
not ( \372_b1 , w_294 );
not ( \372_b0 , w_295 );
and ( w_294 , w_295 , \303_b0 );
or ( \373_b1 , \315_b1 , \313_b1 );
not ( \313_b1 , w_296 );
and ( \373_b0 , \315_b0 , w_297 );
and ( w_296 , w_297 , \313_b0 );
or ( \374_b1 , \159_b1 , \311_b1 );
not ( \311_b1 , w_298 );
and ( \374_b0 , \159_b0 , w_299 );
and ( w_298 , w_299 , \311_b0 );
or ( \375_b1 , \373_b1 , w_301 );
not ( w_301 , w_302 );
and ( \375_b0 , \373_b0 , w_303 );
and ( w_302 ,  , w_303 );
buf ( w_301 , \374_b1 );
not ( w_301 , w_304 );
not (  , w_305 );
and ( w_304 , w_305 , \374_b0 );
or ( \376_b1 , \375_b1 , w_306 );
xor ( \376_b0 , \375_b0 , w_308 );
not ( w_308 , w_309 );
and ( w_309 , w_306 , w_307 );
buf ( w_306 , \320_b1 );
not ( w_306 , w_310 );
not ( w_307 , w_311 );
and ( w_310 , w_311 , \320_b0 );
or ( \377_b1 , \372_b1 , \376_b1 );
xor ( \377_b0 , \372_b0 , w_312 );
not ( w_312 , w_313 );
and ( w_313 , \376_b1 , \376_b0 );
or ( \378_b1 , \333_b1 , \331_b1 );
not ( \331_b1 , w_314 );
and ( \378_b0 , \333_b0 , w_315 );
and ( w_314 , w_315 , \331_b0 );
or ( \379_b1 , \305_b1 , \329_b1 );
not ( \329_b1 , w_316 );
and ( \379_b0 , \305_b0 , w_317 );
and ( w_316 , w_317 , \329_b0 );
or ( \380_b1 , \378_b1 , w_319 );
not ( w_319 , w_320 );
and ( \380_b0 , \378_b0 , w_321 );
and ( w_320 ,  , w_321 );
buf ( w_319 , \379_b1 );
not ( w_319 , w_322 );
not (  , w_323 );
and ( w_322 , w_323 , \379_b0 );
or ( \381_b1 , \380_b1 , w_324 );
xor ( \381_b0 , \380_b0 , w_326 );
not ( w_326 , w_327 );
and ( w_327 , w_324 , w_325 );
buf ( w_324 , \338_b1 );
not ( w_324 , w_328 );
not ( w_325 , w_329 );
and ( w_328 , w_329 , \338_b0 );
or ( \382_b1 , \377_b1 , \381_b1 );
xor ( \382_b0 , \377_b0 , w_330 );
not ( w_330 , w_331 );
and ( w_331 , \381_b1 , \381_b0 );
or ( \383_b1 , \371_b1 , \382_b1 );
not ( \382_b1 , w_332 );
and ( \383_b0 , \371_b0 , w_333 );
and ( w_332 , w_333 , \382_b0 );
or ( \384_b1 , \370_b1 , \383_b1 );
not ( \383_b1 , w_334 );
and ( \384_b0 , \370_b0 , w_335 );
and ( w_334 , w_335 , \383_b0 );
or ( \385_b1 , \372_b1 , \376_b1 );
not ( \376_b1 , w_336 );
and ( \385_b0 , \372_b0 , w_337 );
and ( w_336 , w_337 , \376_b0 );
or ( \386_b1 , \376_b1 , \381_b1 );
not ( \381_b1 , w_338 );
and ( \386_b0 , \376_b0 , w_339 );
and ( w_338 , w_339 , \381_b0 );
or ( \387_b1 , \372_b1 , \381_b1 );
not ( \381_b1 , w_340 );
and ( \387_b0 , \372_b0 , w_341 );
and ( w_340 , w_341 , \381_b0 );
or ( \389_b1 , \159_b1 , \313_b1 );
not ( \313_b1 , w_342 );
and ( \389_b0 , \159_b0 , w_343 );
and ( w_342 , w_343 , \313_b0 );
buf ( \390_b1 , \389_b1 );
not ( \390_b1 , w_344 );
not ( \390_b0 , w_345 );
and ( w_344 , w_345 , \389_b0 );
or ( \391_b1 , \390_b1 , w_346 );
xor ( \391_b0 , \390_b0 , w_348 );
not ( w_348 , w_349 );
and ( w_349 , w_346 , w_347 );
buf ( w_346 , \320_b1 );
not ( w_346 , w_350 );
not ( w_347 , w_351 );
and ( w_350 , w_351 , \320_b0 );
or ( \392_b1 , \305_b1 , \331_b1 );
not ( \331_b1 , w_352 );
and ( \392_b0 , \305_b0 , w_353 );
and ( w_352 , w_353 , \331_b0 );
or ( \393_b1 , \315_b1 , \329_b1 );
not ( \329_b1 , w_354 );
and ( \393_b0 , \315_b0 , w_355 );
and ( w_354 , w_355 , \329_b0 );
or ( \394_b1 , \392_b1 , w_357 );
not ( w_357 , w_358 );
and ( \394_b0 , \392_b0 , w_359 );
and ( w_358 ,  , w_359 );
buf ( w_357 , \393_b1 );
not ( w_357 , w_360 );
not (  , w_361 );
and ( w_360 , w_361 , \393_b0 );
or ( \395_b1 , \394_b1 , w_362 );
xor ( \395_b0 , \394_b0 , w_364 );
not ( w_364 , w_365 );
and ( w_365 , w_362 , w_363 );
buf ( w_362 , \338_b1 );
not ( w_362 , w_366 );
not ( w_363 , w_367 );
and ( w_366 , w_367 , \338_b0 );
or ( \396_b1 , \391_b1 , \395_b1 );
xor ( \396_b0 , \391_b0 , w_368 );
not ( w_368 , w_369 );
and ( w_369 , \395_b1 , \395_b0 );
or ( \397_b1 , \323_b1 , \351_b1 );
not ( \351_b1 , w_370 );
and ( \397_b0 , \323_b0 , w_371 );
and ( w_370 , w_371 , \351_b0 );
or ( \398_b1 , \333_b1 , \349_b1 );
not ( \349_b1 , w_372 );
and ( \398_b0 , \333_b0 , w_373 );
and ( w_372 , w_373 , \349_b0 );
or ( \399_b1 , \397_b1 , w_375 );
not ( w_375 , w_376 );
and ( \399_b0 , \397_b0 , w_377 );
and ( w_376 ,  , w_377 );
buf ( w_375 , \398_b1 );
not ( w_375 , w_378 );
not (  , w_379 );
and ( w_378 , w_379 , \398_b0 );
or ( \400_b1 , \399_b1 , w_380 );
xor ( \400_b0 , \399_b0 , w_382 );
not ( w_382 , w_383 );
and ( w_383 , w_380 , w_381 );
buf ( w_380 , \358_b1 );
not ( w_380 , w_384 );
not ( w_381 , w_385 );
and ( w_384 , w_385 , \358_b0 );
or ( \401_b1 , \396_b1 , \400_b1 );
xor ( \401_b0 , \396_b0 , w_386 );
not ( w_386 , w_387 );
and ( w_387 , \400_b1 , \400_b0 );
or ( \402_b1 , \388_b1 , \401_b1 );
xor ( \402_b0 , \388_b0 , w_388 );
not ( w_388 , w_389 );
and ( w_389 , \401_b1 , \401_b0 );
or ( \403_b1 , \353_b1 , \345_b1 );
not ( \345_b1 , w_390 );
and ( \403_b0 , \353_b0 , w_391 );
and ( w_390 , w_391 , \345_b0 );
buf ( \404_b1 , \403_b1 );
not ( \404_b1 , w_392 );
not ( \404_b0 , w_393 );
and ( w_392 , w_393 , \403_b0 );
or ( \405_b1 , \402_b1 , \404_b1 );
xor ( \405_b0 , \402_b0 , w_394 );
not ( w_394 , w_395 );
and ( w_395 , \404_b1 , \404_b0 );
or ( \406_b1 , \383_b1 , \405_b1 );
not ( \405_b1 , w_396 );
and ( \406_b0 , \383_b0 , w_397 );
and ( w_396 , w_397 , \405_b0 );
or ( \407_b1 , \370_b1 , \405_b1 );
not ( \405_b1 , w_398 );
and ( \407_b0 , \370_b0 , w_399 );
and ( w_398 , w_399 , \405_b0 );
or ( \409_b1 , \388_b1 , \401_b1 );
not ( \401_b1 , w_400 );
and ( \409_b0 , \388_b0 , w_401 );
and ( w_400 , w_401 , \401_b0 );
or ( \410_b1 , \401_b1 , \404_b1 );
not ( \404_b1 , w_402 );
and ( \410_b0 , \401_b0 , w_403 );
and ( w_402 , w_403 , \404_b0 );
or ( \411_b1 , \388_b1 , \404_b1 );
not ( \404_b1 , w_404 );
and ( \411_b0 , \388_b0 , w_405 );
and ( w_404 , w_405 , \404_b0 );
buf ( \413_b1 , \320_b1 );
not ( \413_b1 , w_406 );
not ( \413_b0 , w_407 );
and ( w_406 , w_407 , \320_b0 );
or ( \414_b1 , \315_b1 , \331_b1 );
not ( \331_b1 , w_408 );
and ( \414_b0 , \315_b0 , w_409 );
and ( w_408 , w_409 , \331_b0 );
or ( \415_b1 , \159_b1 , \329_b1 );
not ( \329_b1 , w_410 );
and ( \415_b0 , \159_b0 , w_411 );
and ( w_410 , w_411 , \329_b0 );
or ( \416_b1 , \414_b1 , w_413 );
not ( w_413 , w_414 );
and ( \416_b0 , \414_b0 , w_415 );
and ( w_414 ,  , w_415 );
buf ( w_413 , \415_b1 );
not ( w_413 , w_416 );
not (  , w_417 );
and ( w_416 , w_417 , \415_b0 );
or ( \417_b1 , \416_b1 , w_418 );
xor ( \417_b0 , \416_b0 , w_420 );
not ( w_420 , w_421 );
and ( w_421 , w_418 , w_419 );
buf ( w_418 , \338_b1 );
not ( w_418 , w_422 );
not ( w_419 , w_423 );
and ( w_422 , w_423 , \338_b0 );
or ( \418_b1 , \413_b1 , \417_b1 );
xor ( \418_b0 , \413_b0 , w_424 );
not ( w_424 , w_425 );
and ( w_425 , \417_b1 , \417_b0 );
or ( \419_b1 , \333_b1 , \351_b1 );
not ( \351_b1 , w_426 );
and ( \419_b0 , \333_b0 , w_427 );
and ( w_426 , w_427 , \351_b0 );
or ( \420_b1 , \305_b1 , \349_b1 );
not ( \349_b1 , w_428 );
and ( \420_b0 , \305_b0 , w_429 );
and ( w_428 , w_429 , \349_b0 );
or ( \421_b1 , \419_b1 , w_431 );
not ( w_431 , w_432 );
and ( \421_b0 , \419_b0 , w_433 );
and ( w_432 ,  , w_433 );
buf ( w_431 , \420_b1 );
not ( w_431 , w_434 );
not (  , w_435 );
and ( w_434 , w_435 , \420_b0 );
or ( \422_b1 , \421_b1 , w_436 );
xor ( \422_b0 , \421_b0 , w_438 );
not ( w_438 , w_439 );
and ( w_439 , w_436 , w_437 );
buf ( w_436 , \358_b1 );
not ( w_436 , w_440 );
not ( w_437 , w_441 );
and ( w_440 , w_441 , \358_b0 );
or ( \423_b1 , \418_b1 , \422_b1 );
xor ( \423_b0 , \418_b0 , w_442 );
not ( w_442 , w_443 );
and ( w_443 , \422_b1 , \422_b0 );
or ( \424_b1 , \412_b1 , \423_b1 );
xor ( \424_b0 , \412_b0 , w_444 );
not ( w_444 , w_445 );
and ( w_445 , \423_b1 , \423_b0 );
or ( \425_b1 , \391_b1 , \395_b1 );
not ( \395_b1 , w_446 );
and ( \425_b0 , \391_b0 , w_447 );
and ( w_446 , w_447 , \395_b0 );
or ( \426_b1 , \395_b1 , \400_b1 );
not ( \400_b1 , w_448 );
and ( \426_b0 , \395_b0 , w_449 );
and ( w_448 , w_449 , \400_b0 );
or ( \427_b1 , \391_b1 , \400_b1 );
not ( \400_b1 , w_450 );
and ( \427_b0 , \391_b0 , w_451 );
and ( w_450 , w_451 , \400_b0 );
buf ( \429_b1 , \403_b1 );
buf ( \429_b0 , \403_b0 );
or ( \430_b1 , \428_b1 , \429_b1 );
xor ( \430_b0 , \428_b0 , w_452 );
not ( w_452 , w_453 );
and ( w_453 , \429_b1 , \429_b0 );
or ( \431_b1 , \323_b1 , \345_b1 );
not ( \345_b1 , w_454 );
and ( \431_b0 , \323_b0 , w_455 );
and ( w_454 , w_455 , \345_b0 );
or ( \432_b1 , \430_b1 , \431_b1 );
xor ( \432_b0 , \430_b0 , w_456 );
not ( w_456 , w_457 );
and ( w_457 , \431_b1 , \431_b0 );
or ( \433_b1 , \424_b1 , \432_b1 );
xor ( \433_b0 , \424_b0 , w_458 );
not ( w_458 , w_459 );
and ( w_459 , \432_b1 , \432_b0 );
or ( \434_b1 , \408_b1 , \433_b1 );
xor ( \434_b0 , \408_b0 , w_460 );
not ( w_460 , w_461 );
and ( w_461 , \433_b1 , \433_b0 );
or ( \435_b1 , \353_b1 , \331_b1 );
not ( \331_b1 , w_462 );
and ( \435_b0 , \353_b0 , w_463 );
and ( w_462 , w_463 , \331_b0 );
or ( \436_b1 , \323_b1 , \329_b1 );
not ( \329_b1 , w_464 );
and ( \436_b0 , \323_b0 , w_465 );
and ( w_464 , w_465 , \329_b0 );
or ( \437_b1 , \435_b1 , w_467 );
not ( w_467 , w_468 );
and ( \437_b0 , \435_b0 , w_469 );
and ( w_468 ,  , w_469 );
buf ( w_467 , \436_b1 );
not ( w_467 , w_470 );
not (  , w_471 );
and ( w_470 , w_471 , \436_b0 );
or ( \438_b1 , \437_b1 , w_472 );
xor ( \438_b0 , \437_b0 , w_474 );
not ( w_474 , w_475 );
and ( w_475 , w_472 , w_473 );
buf ( w_472 , \338_b1 );
not ( w_472 , w_476 );
not ( w_473 , w_477 );
and ( w_476 , w_477 , \338_b0 );
or ( \439_b1 , \360_b1 , \351_b1 );
not ( \351_b1 , w_478 );
and ( \439_b0 , \360_b0 , w_479 );
and ( w_478 , w_479 , \351_b0 );
or ( \440_b1 , \343_b1 , \349_b1 );
not ( \349_b1 , w_480 );
and ( \440_b0 , \343_b0 , w_481 );
and ( w_480 , w_481 , \349_b0 );
or ( \441_b1 , \439_b1 , w_483 );
not ( w_483 , w_484 );
and ( \441_b0 , \439_b0 , w_485 );
and ( w_484 ,  , w_485 );
buf ( w_483 , \440_b1 );
not ( w_483 , w_486 );
not (  , w_487 );
and ( w_486 , w_487 , \440_b0 );
or ( \442_b1 , \441_b1 , w_488 );
xor ( \442_b0 , \441_b0 , w_490 );
not ( w_490 , w_491 );
and ( w_491 , w_488 , w_489 );
buf ( w_488 , \358_b1 );
not ( w_488 , w_492 );
not ( w_489 , w_493 );
and ( w_492 , w_493 , \358_b0 );
or ( \443_b1 , \438_b1 , \442_b1 );
not ( \442_b1 , w_494 );
and ( \443_b0 , \438_b0 , w_495 );
and ( w_494 , w_495 , \442_b0 );
buf ( \444_b1 , RIb4bf678_73_b1 );
buf ( \444_b0 , RIb4bf678_73_b0 );
or ( \445_b1 , \444_b1 , \345_b1 );
not ( \345_b1 , w_496 );
and ( \445_b0 , \444_b0 , w_497 );
and ( w_496 , w_497 , \345_b0 );
or ( \446_b1 , \442_b1 , \445_b1 );
not ( \445_b1 , w_498 );
and ( \446_b0 , \442_b0 , w_499 );
and ( w_498 , w_499 , \445_b0 );
or ( \447_b1 , \438_b1 , \445_b1 );
not ( \445_b1 , w_500 );
and ( \447_b0 , \438_b0 , w_501 );
and ( w_500 , w_501 , \445_b0 );
and ( \449_nR13a_b1 , RIb4c6860_42_b1 , w_502 );
xor ( w_502 , RIb4c6860_42_b0 , \288_b1 );
not ( \288_b1 , w_503 );
and ( \449_nR13a_b0 , w_503 , \288_b0 );
buf ( \450_b1 , \449_nR13a_b1 );
buf ( \450_b0 , \449_nR13a_b0 );
and ( \451_nR139_b1 , RIb4c67e8_43_b1 , w_504 );
xor ( w_504 , RIb4c67e8_43_b0 , \288_b1 );
not ( \288_b1 , w_505 );
and ( \451_nR139_b0 , w_505 , \288_b0 );
buf ( \452_b1 , \451_nR139_b1 );
buf ( \452_b0 , \451_nR139_b0 );
or ( \453_b1 , \450_b1 , \452_b1 );
not ( \452_b1 , w_506 );
and ( \453_b0 , \450_b0 , w_507 );
and ( w_506 , w_507 , \452_b0 );
buf ( \454_b1 , \453_b1 );
not ( \454_b1 , w_508 );
not ( \454_b0 , w_509 );
and ( w_508 , w_509 , \453_b0 );
or ( \455_b1 , \295_b1 , \454_b1 );
not ( \454_b1 , w_510 );
and ( \455_b0 , \295_b0 , w_511 );
and ( w_510 , w_511 , \454_b0 );
buf ( \456_b1 , \455_b1 );
not ( \456_b1 , w_512 );
not ( \456_b0 , w_513 );
and ( w_512 , w_513 , \455_b0 );
or ( \457_b1 , \315_b1 , \298_b1 );
not ( \298_b1 , w_514 );
and ( \457_b0 , \315_b0 , w_515 );
and ( w_514 , w_515 , \298_b0 );
or ( \458_b1 , \159_b1 , \296_b1 );
not ( \296_b1 , w_516 );
and ( \458_b0 , \159_b0 , w_517 );
and ( w_516 , w_517 , \296_b0 );
or ( \459_b1 , \457_b1 , w_519 );
not ( w_519 , w_520 );
and ( \459_b0 , \457_b0 , w_521 );
and ( w_520 ,  , w_521 );
buf ( w_519 , \458_b1 );
not ( w_519 , w_522 );
not (  , w_523 );
and ( w_522 , w_523 , \458_b0 );
or ( \460_b1 , \459_b1 , w_524 );
xor ( \460_b0 , \459_b0 , w_526 );
not ( w_526 , w_527 );
and ( w_527 , w_524 , w_525 );
buf ( w_524 , \303_b1 );
not ( w_524 , w_528 );
not ( w_525 , w_529 );
and ( w_528 , w_529 , \303_b0 );
or ( \461_b1 , \456_b1 , \460_b1 );
not ( \460_b1 , w_530 );
and ( \461_b0 , \456_b0 , w_531 );
and ( w_530 , w_531 , \460_b0 );
or ( \462_b1 , \333_b1 , \313_b1 );
not ( \313_b1 , w_532 );
and ( \462_b0 , \333_b0 , w_533 );
and ( w_532 , w_533 , \313_b0 );
or ( \463_b1 , \305_b1 , \311_b1 );
not ( \311_b1 , w_534 );
and ( \463_b0 , \305_b0 , w_535 );
and ( w_534 , w_535 , \311_b0 );
or ( \464_b1 , \462_b1 , w_537 );
not ( w_537 , w_538 );
and ( \464_b0 , \462_b0 , w_539 );
and ( w_538 ,  , w_539 );
buf ( w_537 , \463_b1 );
not ( w_537 , w_540 );
not (  , w_541 );
and ( w_540 , w_541 , \463_b0 );
or ( \465_b1 , \464_b1 , w_542 );
xor ( \465_b0 , \464_b0 , w_544 );
not ( w_544 , w_545 );
and ( w_545 , w_542 , w_543 );
buf ( w_542 , \320_b1 );
not ( w_542 , w_546 );
not ( w_543 , w_547 );
and ( w_546 , w_547 , \320_b0 );
or ( \466_b1 , \460_b1 , \465_b1 );
not ( \465_b1 , w_548 );
and ( \466_b0 , \460_b0 , w_549 );
and ( w_548 , w_549 , \465_b0 );
or ( \467_b1 , \456_b1 , \465_b1 );
not ( \465_b1 , w_550 );
and ( \467_b0 , \456_b0 , w_551 );
and ( w_550 , w_551 , \465_b0 );
or ( \469_b1 , \448_b1 , \468_b1 );
not ( \468_b1 , w_552 );
and ( \469_b0 , \448_b0 , w_553 );
and ( w_552 , w_553 , \468_b0 );
or ( \470_b1 , \359_b1 , w_554 );
xor ( \470_b0 , \359_b0 , w_556 );
not ( w_556 , w_557 );
and ( w_557 , w_554 , w_555 );
buf ( w_554 , \361_b1 );
not ( w_554 , w_558 );
not ( w_555 , w_559 );
and ( w_558 , w_559 , \361_b0 );
or ( \471_b1 , \468_b1 , \470_b1 );
not ( \470_b1 , w_560 );
and ( \471_b0 , \468_b0 , w_561 );
and ( w_560 , w_561 , \470_b0 );
or ( \472_b1 , \448_b1 , \470_b1 );
not ( \470_b1 , w_562 );
and ( \472_b0 , \448_b0 , w_563 );
and ( w_562 , w_563 , \470_b0 );
or ( \474_b1 , \342_b1 , \362_b1 );
xor ( \474_b0 , \342_b0 , w_564 );
not ( w_564 , w_565 );
and ( w_565 , \362_b1 , \362_b0 );
or ( \475_b1 , \474_b1 , \367_b1 );
xor ( \475_b0 , \474_b0 , w_566 );
not ( w_566 , w_567 );
and ( w_567 , \367_b1 , \367_b0 );
or ( \476_b1 , \473_b1 , \475_b1 );
not ( \475_b1 , w_568 );
and ( \476_b0 , \473_b0 , w_569 );
and ( w_568 , w_569 , \475_b0 );
or ( \477_b1 , \371_b1 , \382_b1 );
xor ( \477_b0 , \371_b0 , w_570 );
not ( w_570 , w_571 );
and ( w_571 , \382_b1 , \382_b0 );
or ( \478_b1 , \475_b1 , \477_b1 );
not ( \477_b1 , w_572 );
and ( \478_b0 , \475_b0 , w_573 );
and ( w_572 , w_573 , \477_b0 );
or ( \479_b1 , \473_b1 , \477_b1 );
not ( \477_b1 , w_574 );
and ( \479_b0 , \473_b0 , w_575 );
and ( w_574 , w_575 , \477_b0 );
or ( \481_b1 , \370_b1 , \383_b1 );
xor ( \481_b0 , \370_b0 , w_576 );
not ( w_576 , w_577 );
and ( w_577 , \383_b1 , \383_b0 );
or ( \482_b1 , \481_b1 , \405_b1 );
xor ( \482_b0 , \481_b0 , w_578 );
not ( w_578 , w_579 );
and ( w_579 , \405_b1 , \405_b0 );
or ( \483_b1 , \480_b1 , \482_b1 );
not ( \482_b1 , w_580 );
and ( \483_b0 , \480_b0 , w_581 );
and ( w_580 , w_581 , \482_b0 );
or ( \484_b1 , \434_b1 , \483_b1 );
xor ( \484_b0 , \434_b0 , w_582 );
not ( w_582 , w_583 );
and ( w_583 , \483_b1 , \483_b0 );
or ( \485_b1 , \480_b1 , \482_b1 );
xor ( \485_b0 , \480_b0 , w_584 );
not ( w_584 , w_585 );
and ( w_585 , \482_b1 , \482_b0 );
or ( \486_b1 , \343_b1 , \331_b1 );
not ( \331_b1 , w_586 );
and ( \486_b0 , \343_b0 , w_587 );
and ( w_586 , w_587 , \331_b0 );
or ( \487_b1 , \353_b1 , \329_b1 );
not ( \329_b1 , w_588 );
and ( \487_b0 , \353_b0 , w_589 );
and ( w_588 , w_589 , \329_b0 );
or ( \488_b1 , \486_b1 , w_591 );
not ( w_591 , w_592 );
and ( \488_b0 , \486_b0 , w_593 );
and ( w_592 ,  , w_593 );
buf ( w_591 , \487_b1 );
not ( w_591 , w_594 );
not (  , w_595 );
and ( w_594 , w_595 , \487_b0 );
or ( \489_b1 , \488_b1 , w_596 );
xor ( \489_b0 , \488_b0 , w_598 );
not ( w_598 , w_599 );
and ( w_599 , w_596 , w_597 );
buf ( w_596 , \338_b1 );
not ( w_596 , w_600 );
not ( w_597 , w_601 );
and ( w_600 , w_601 , \338_b0 );
or ( \490_b1 , \444_b1 , \351_b1 );
not ( \351_b1 , w_602 );
and ( \490_b0 , \444_b0 , w_603 );
and ( w_602 , w_603 , \351_b0 );
or ( \491_b1 , \360_b1 , \349_b1 );
not ( \349_b1 , w_604 );
and ( \491_b0 , \360_b0 , w_605 );
and ( w_604 , w_605 , \349_b0 );
or ( \492_b1 , \490_b1 , w_607 );
not ( w_607 , w_608 );
and ( \492_b0 , \490_b0 , w_609 );
and ( w_608 ,  , w_609 );
buf ( w_607 , \491_b1 );
not ( w_607 , w_610 );
not (  , w_611 );
and ( w_610 , w_611 , \491_b0 );
or ( \493_b1 , \492_b1 , w_612 );
xor ( \493_b0 , \492_b0 , w_614 );
not ( w_614 , w_615 );
and ( w_615 , w_612 , w_613 );
buf ( w_612 , \358_b1 );
not ( w_612 , w_616 );
not ( w_613 , w_617 );
and ( w_616 , w_617 , \358_b0 );
or ( \494_b1 , \489_b1 , \493_b1 );
not ( \493_b1 , w_618 );
and ( \494_b0 , \489_b0 , w_619 );
and ( w_618 , w_619 , \493_b0 );
buf ( \495_b1 , RIb4bf600_74_b1 );
buf ( \495_b0 , RIb4bf600_74_b0 );
or ( \496_b1 , \495_b1 , \345_b1 );
not ( \345_b1 , w_620 );
and ( \496_b0 , \495_b0 , w_621 );
and ( w_620 , w_621 , \345_b0 );
or ( \497_b1 , \493_b1 , \496_b1 );
not ( \496_b1 , w_622 );
and ( \497_b0 , \493_b0 , w_623 );
and ( w_622 , w_623 , \496_b0 );
or ( \498_b1 , \489_b1 , \496_b1 );
not ( \496_b1 , w_624 );
and ( \498_b0 , \489_b0 , w_625 );
and ( w_624 , w_625 , \496_b0 );
or ( \500_b1 , \295_b1 , \450_b1 );
xor ( \500_b0 , \295_b0 , w_626 );
not ( w_626 , w_627 );
and ( w_627 , \450_b1 , \450_b0 );
or ( \501_b1 , \450_b1 , \452_b1 );
xor ( \501_b0 , \450_b0 , w_628 );
not ( w_628 , w_629 );
and ( w_629 , \452_b1 , \452_b0 );
buf ( \502_b1 , \501_b1 );
not ( \502_b1 , w_630 );
not ( \502_b0 , w_631 );
and ( w_630 , w_631 , \501_b0 );
or ( \503_b1 , \500_b1 , \502_b1 );
not ( \502_b1 , w_632 );
and ( \503_b0 , \500_b0 , w_633 );
and ( w_632 , w_633 , \502_b0 );
or ( \504_b1 , \159_b1 , \503_b1 );
not ( \503_b1 , w_634 );
and ( \504_b0 , \159_b0 , w_635 );
and ( w_634 , w_635 , \503_b0 );
buf ( \505_b1 , \504_b1 );
not ( \505_b1 , w_636 );
not ( \505_b0 , w_637 );
and ( w_636 , w_637 , \504_b0 );
or ( \506_b1 , \505_b1 , w_638 );
xor ( \506_b0 , \505_b0 , w_640 );
not ( w_640 , w_641 );
and ( w_641 , w_638 , w_639 );
buf ( w_638 , \455_b1 );
not ( w_638 , w_642 );
not ( w_639 , w_643 );
and ( w_642 , w_643 , \455_b0 );
or ( \507_b1 , \305_b1 , \298_b1 );
not ( \298_b1 , w_644 );
and ( \507_b0 , \305_b0 , w_645 );
and ( w_644 , w_645 , \298_b0 );
or ( \508_b1 , \315_b1 , \296_b1 );
not ( \296_b1 , w_646 );
and ( \508_b0 , \315_b0 , w_647 );
and ( w_646 , w_647 , \296_b0 );
or ( \509_b1 , \507_b1 , w_649 );
not ( w_649 , w_650 );
and ( \509_b0 , \507_b0 , w_651 );
and ( w_650 ,  , w_651 );
buf ( w_649 , \508_b1 );
not ( w_649 , w_652 );
not (  , w_653 );
and ( w_652 , w_653 , \508_b0 );
or ( \510_b1 , \509_b1 , w_654 );
xor ( \510_b0 , \509_b0 , w_656 );
not ( w_656 , w_657 );
and ( w_657 , w_654 , w_655 );
buf ( w_654 , \303_b1 );
not ( w_654 , w_658 );
not ( w_655 , w_659 );
and ( w_658 , w_659 , \303_b0 );
or ( \511_b1 , \506_b1 , \510_b1 );
not ( \510_b1 , w_660 );
and ( \511_b0 , \506_b0 , w_661 );
and ( w_660 , w_661 , \510_b0 );
or ( \512_b1 , \323_b1 , \313_b1 );
not ( \313_b1 , w_662 );
and ( \512_b0 , \323_b0 , w_663 );
and ( w_662 , w_663 , \313_b0 );
or ( \513_b1 , \333_b1 , \311_b1 );
not ( \311_b1 , w_664 );
and ( \513_b0 , \333_b0 , w_665 );
and ( w_664 , w_665 , \311_b0 );
or ( \514_b1 , \512_b1 , w_667 );
not ( w_667 , w_668 );
and ( \514_b0 , \512_b0 , w_669 );
and ( w_668 ,  , w_669 );
buf ( w_667 , \513_b1 );
not ( w_667 , w_670 );
not (  , w_671 );
and ( w_670 , w_671 , \513_b0 );
or ( \515_b1 , \514_b1 , w_672 );
xor ( \515_b0 , \514_b0 , w_674 );
not ( w_674 , w_675 );
and ( w_675 , w_672 , w_673 );
buf ( w_672 , \320_b1 );
not ( w_672 , w_676 );
not ( w_673 , w_677 );
and ( w_676 , w_677 , \320_b0 );
or ( \516_b1 , \510_b1 , \515_b1 );
not ( \515_b1 , w_678 );
and ( \516_b0 , \510_b0 , w_679 );
and ( w_678 , w_679 , \515_b0 );
or ( \517_b1 , \506_b1 , \515_b1 );
not ( \515_b1 , w_680 );
and ( \517_b0 , \506_b0 , w_681 );
and ( w_680 , w_681 , \515_b0 );
or ( \519_b1 , \499_b1 , \518_b1 );
not ( \518_b1 , w_682 );
and ( \519_b0 , \499_b0 , w_683 );
and ( w_682 , w_683 , \518_b0 );
or ( \520_b1 , \438_b1 , \442_b1 );
xor ( \520_b0 , \438_b0 , w_684 );
not ( w_684 , w_685 );
and ( w_685 , \442_b1 , \442_b0 );
or ( \521_b1 , \520_b1 , \445_b1 );
xor ( \521_b0 , \520_b0 , w_686 );
not ( w_686 , w_687 );
and ( w_687 , \445_b1 , \445_b0 );
or ( \522_b1 , \518_b1 , \521_b1 );
not ( \521_b1 , w_688 );
and ( \522_b0 , \518_b0 , w_689 );
and ( w_688 , w_689 , \521_b0 );
or ( \523_b1 , \499_b1 , \521_b1 );
not ( \521_b1 , w_690 );
and ( \523_b0 , \499_b0 , w_691 );
and ( w_690 , w_691 , \521_b0 );
or ( \525_b1 , \304_b1 , \321_b1 );
xor ( \525_b0 , \304_b0 , w_692 );
not ( w_692 , w_693 );
and ( w_693 , \321_b1 , \321_b0 );
or ( \526_b1 , \525_b1 , \339_b1 );
xor ( \526_b0 , \525_b0 , w_694 );
not ( w_694 , w_695 );
and ( w_695 , \339_b1 , \339_b0 );
or ( \527_b1 , \524_b1 , \526_b1 );
not ( \526_b1 , w_696 );
and ( \527_b0 , \524_b0 , w_697 );
and ( w_696 , w_697 , \526_b0 );
or ( \528_b1 , \448_b1 , \468_b1 );
xor ( \528_b0 , \448_b0 , w_698 );
not ( w_698 , w_699 );
and ( w_699 , \468_b1 , \468_b0 );
or ( \529_b1 , \528_b1 , \470_b1 );
xor ( \529_b0 , \528_b0 , w_700 );
not ( w_700 , w_701 );
and ( w_701 , \470_b1 , \470_b0 );
or ( \530_b1 , \526_b1 , \529_b1 );
not ( \529_b1 , w_702 );
and ( \530_b0 , \526_b0 , w_703 );
and ( w_702 , w_703 , \529_b0 );
or ( \531_b1 , \524_b1 , \529_b1 );
not ( \529_b1 , w_704 );
and ( \531_b0 , \524_b0 , w_705 );
and ( w_704 , w_705 , \529_b0 );
or ( \533_b1 , \473_b1 , \475_b1 );
xor ( \533_b0 , \473_b0 , w_706 );
not ( w_706 , w_707 );
and ( w_707 , \475_b1 , \475_b0 );
or ( \534_b1 , \533_b1 , \477_b1 );
xor ( \534_b0 , \533_b0 , w_708 );
not ( w_708 , w_709 );
and ( w_709 , \477_b1 , \477_b0 );
or ( \535_b1 , \532_b1 , \534_b1 );
not ( \534_b1 , w_710 );
and ( \535_b0 , \532_b0 , w_711 );
and ( w_710 , w_711 , \534_b0 );
or ( \536_b1 , \485_b1 , \535_b1 );
not ( \535_b1 , w_712 );
and ( \536_b0 , \485_b0 , w_713 );
and ( w_712 , w_713 , \535_b0 );
or ( \537_b1 , \485_b1 , \535_b1 );
xor ( \537_b0 , \485_b0 , w_714 );
not ( w_714 , w_715 );
and ( w_715 , \535_b1 , \535_b0 );
or ( \538_b1 , \532_b1 , \534_b1 );
xor ( \538_b0 , \532_b0 , w_716 );
not ( w_716 , w_717 );
and ( w_717 , \534_b1 , \534_b0 );
or ( \539_b1 , \353_b1 , \313_b1 );
not ( \313_b1 , w_718 );
and ( \539_b0 , \353_b0 , w_719 );
and ( w_718 , w_719 , \313_b0 );
or ( \540_b1 , \323_b1 , \311_b1 );
not ( \311_b1 , w_720 );
and ( \540_b0 , \323_b0 , w_721 );
and ( w_720 , w_721 , \311_b0 );
or ( \541_b1 , \539_b1 , w_723 );
not ( w_723 , w_724 );
and ( \541_b0 , \539_b0 , w_725 );
and ( w_724 ,  , w_725 );
buf ( w_723 , \540_b1 );
not ( w_723 , w_726 );
not (  , w_727 );
and ( w_726 , w_727 , \540_b0 );
or ( \542_b1 , \541_b1 , w_728 );
xor ( \542_b0 , \541_b0 , w_730 );
not ( w_730 , w_731 );
and ( w_731 , w_728 , w_729 );
buf ( w_728 , \320_b1 );
not ( w_728 , w_732 );
not ( w_729 , w_733 );
and ( w_732 , w_733 , \320_b0 );
or ( \543_b1 , \360_b1 , \331_b1 );
not ( \331_b1 , w_734 );
and ( \543_b0 , \360_b0 , w_735 );
and ( w_734 , w_735 , \331_b0 );
or ( \544_b1 , \343_b1 , \329_b1 );
not ( \329_b1 , w_736 );
and ( \544_b0 , \343_b0 , w_737 );
and ( w_736 , w_737 , \329_b0 );
or ( \545_b1 , \543_b1 , w_739 );
not ( w_739 , w_740 );
and ( \545_b0 , \543_b0 , w_741 );
and ( w_740 ,  , w_741 );
buf ( w_739 , \544_b1 );
not ( w_739 , w_742 );
not (  , w_743 );
and ( w_742 , w_743 , \544_b0 );
or ( \546_b1 , \545_b1 , w_744 );
xor ( \546_b0 , \545_b0 , w_746 );
not ( w_746 , w_747 );
and ( w_747 , w_744 , w_745 );
buf ( w_744 , \338_b1 );
not ( w_744 , w_748 );
not ( w_745 , w_749 );
and ( w_748 , w_749 , \338_b0 );
or ( \547_b1 , \542_b1 , \546_b1 );
not ( \546_b1 , w_750 );
and ( \547_b0 , \542_b0 , w_751 );
and ( w_750 , w_751 , \546_b0 );
or ( \548_b1 , \495_b1 , \351_b1 );
not ( \351_b1 , w_752 );
and ( \548_b0 , \495_b0 , w_753 );
and ( w_752 , w_753 , \351_b0 );
or ( \549_b1 , \444_b1 , \349_b1 );
not ( \349_b1 , w_754 );
and ( \549_b0 , \444_b0 , w_755 );
and ( w_754 , w_755 , \349_b0 );
or ( \550_b1 , \548_b1 , w_757 );
not ( w_757 , w_758 );
and ( \550_b0 , \548_b0 , w_759 );
and ( w_758 ,  , w_759 );
buf ( w_757 , \549_b1 );
not ( w_757 , w_760 );
not (  , w_761 );
and ( w_760 , w_761 , \549_b0 );
or ( \551_b1 , \550_b1 , w_762 );
xor ( \551_b0 , \550_b0 , w_764 );
not ( w_764 , w_765 );
and ( w_765 , w_762 , w_763 );
buf ( w_762 , \358_b1 );
not ( w_762 , w_766 );
not ( w_763 , w_767 );
and ( w_766 , w_767 , \358_b0 );
or ( \552_b1 , \546_b1 , \551_b1 );
not ( \551_b1 , w_768 );
and ( \552_b0 , \546_b0 , w_769 );
and ( w_768 , w_769 , \551_b0 );
or ( \553_b1 , \542_b1 , \551_b1 );
not ( \551_b1 , w_770 );
and ( \553_b0 , \542_b0 , w_771 );
and ( w_770 , w_771 , \551_b0 );
and ( \555_nR138_b1 , RIb4c6770_44_b1 , w_772 );
xor ( w_772 , RIb4c6770_44_b0 , \288_b1 );
not ( \288_b1 , w_773 );
and ( \555_nR138_b0 , w_773 , \288_b0 );
buf ( \556_b1 , \555_nR138_b1 );
buf ( \556_b0 , \555_nR138_b0 );
and ( \557_nR137_b1 , RIb4c3368_45_b1 , w_774 );
xor ( w_774 , RIb4c3368_45_b0 , \288_b1 );
not ( \288_b1 , w_775 );
and ( \557_nR137_b0 , w_775 , \288_b0 );
buf ( \558_b1 , \557_nR137_b1 );
buf ( \558_b0 , \557_nR137_b0 );
or ( \559_b1 , \556_b1 , \558_b1 );
not ( \558_b1 , w_776 );
and ( \559_b0 , \556_b0 , w_777 );
and ( w_776 , w_777 , \558_b0 );
buf ( \560_b1 , \559_b1 );
not ( \560_b1 , w_778 );
not ( \560_b0 , w_779 );
and ( w_778 , w_779 , \559_b0 );
or ( \561_b1 , \452_b1 , \560_b1 );
not ( \560_b1 , w_780 );
and ( \561_b0 , \452_b0 , w_781 );
and ( w_780 , w_781 , \560_b0 );
buf ( \562_b1 , \561_b1 );
not ( \562_b1 , w_782 );
not ( \562_b0 , w_783 );
and ( w_782 , w_783 , \561_b0 );
or ( \563_b1 , \315_b1 , \503_b1 );
not ( \503_b1 , w_784 );
and ( \563_b0 , \315_b0 , w_785 );
and ( w_784 , w_785 , \503_b0 );
or ( \564_b1 , \159_b1 , \501_b1 );
not ( \501_b1 , w_786 );
and ( \564_b0 , \159_b0 , w_787 );
and ( w_786 , w_787 , \501_b0 );
or ( \565_b1 , \563_b1 , w_789 );
not ( w_789 , w_790 );
and ( \565_b0 , \563_b0 , w_791 );
and ( w_790 ,  , w_791 );
buf ( w_789 , \564_b1 );
not ( w_789 , w_792 );
not (  , w_793 );
and ( w_792 , w_793 , \564_b0 );
or ( \566_b1 , \565_b1 , w_794 );
xor ( \566_b0 , \565_b0 , w_796 );
not ( w_796 , w_797 );
and ( w_797 , w_794 , w_795 );
buf ( w_794 , \455_b1 );
not ( w_794 , w_798 );
not ( w_795 , w_799 );
and ( w_798 , w_799 , \455_b0 );
or ( \567_b1 , \562_b1 , \566_b1 );
not ( \566_b1 , w_800 );
and ( \567_b0 , \562_b0 , w_801 );
and ( w_800 , w_801 , \566_b0 );
or ( \568_b1 , \333_b1 , \298_b1 );
not ( \298_b1 , w_802 );
and ( \568_b0 , \333_b0 , w_803 );
and ( w_802 , w_803 , \298_b0 );
or ( \569_b1 , \305_b1 , \296_b1 );
not ( \296_b1 , w_804 );
and ( \569_b0 , \305_b0 , w_805 );
and ( w_804 , w_805 , \296_b0 );
or ( \570_b1 , \568_b1 , w_807 );
not ( w_807 , w_808 );
and ( \570_b0 , \568_b0 , w_809 );
and ( w_808 ,  , w_809 );
buf ( w_807 , \569_b1 );
not ( w_807 , w_810 );
not (  , w_811 );
and ( w_810 , w_811 , \569_b0 );
or ( \571_b1 , \570_b1 , w_812 );
xor ( \571_b0 , \570_b0 , w_814 );
not ( w_814 , w_815 );
and ( w_815 , w_812 , w_813 );
buf ( w_812 , \303_b1 );
not ( w_812 , w_816 );
not ( w_813 , w_817 );
and ( w_816 , w_817 , \303_b0 );
or ( \572_b1 , \566_b1 , \571_b1 );
not ( \571_b1 , w_818 );
and ( \572_b0 , \566_b0 , w_819 );
and ( w_818 , w_819 , \571_b0 );
or ( \573_b1 , \562_b1 , \571_b1 );
not ( \571_b1 , w_820 );
and ( \573_b0 , \562_b0 , w_821 );
and ( w_820 , w_821 , \571_b0 );
or ( \575_b1 , \554_b1 , w_822 );
or ( \575_b0 , \554_b0 , \574_b0 );
not ( \574_b0 , w_823 );
and ( w_823 , w_822 , \574_b1 );
or ( \576_b1 , \456_b1 , \460_b1 );
xor ( \576_b0 , \456_b0 , w_824 );
not ( w_824 , w_825 );
and ( w_825 , \460_b1 , \460_b0 );
or ( \577_b1 , \576_b1 , \465_b1 );
xor ( \577_b0 , \576_b0 , w_826 );
not ( w_826 , w_827 );
and ( w_827 , \465_b1 , \465_b0 );
or ( \578_b1 , \575_b1 , \577_b1 );
not ( \577_b1 , w_828 );
and ( \578_b0 , \575_b0 , w_829 );
and ( w_828 , w_829 , \577_b0 );
or ( \579_b1 , \499_b1 , \518_b1 );
xor ( \579_b0 , \499_b0 , w_830 );
not ( w_830 , w_831 );
and ( w_831 , \518_b1 , \518_b0 );
or ( \580_b1 , \579_b1 , \521_b1 );
xor ( \580_b0 , \579_b0 , w_832 );
not ( w_832 , w_833 );
and ( w_833 , \521_b1 , \521_b0 );
or ( \581_b1 , \577_b1 , \580_b1 );
not ( \580_b1 , w_834 );
and ( \581_b0 , \577_b0 , w_835 );
and ( w_834 , w_835 , \580_b0 );
or ( \582_b1 , \575_b1 , \580_b1 );
not ( \580_b1 , w_836 );
and ( \582_b0 , \575_b0 , w_837 );
and ( w_836 , w_837 , \580_b0 );
or ( \584_b1 , \343_b1 , \313_b1 );
not ( \313_b1 , w_838 );
and ( \584_b0 , \343_b0 , w_839 );
and ( w_838 , w_839 , \313_b0 );
or ( \585_b1 , \353_b1 , \311_b1 );
not ( \311_b1 , w_840 );
and ( \585_b0 , \353_b0 , w_841 );
and ( w_840 , w_841 , \311_b0 );
or ( \586_b1 , \584_b1 , w_843 );
not ( w_843 , w_844 );
and ( \586_b0 , \584_b0 , w_845 );
and ( w_844 ,  , w_845 );
buf ( w_843 , \585_b1 );
not ( w_843 , w_846 );
not (  , w_847 );
and ( w_846 , w_847 , \585_b0 );
or ( \587_b1 , \586_b1 , w_848 );
xor ( \587_b0 , \586_b0 , w_850 );
not ( w_850 , w_851 );
and ( w_851 , w_848 , w_849 );
buf ( w_848 , \320_b1 );
not ( w_848 , w_852 );
not ( w_849 , w_853 );
and ( w_852 , w_853 , \320_b0 );
or ( \588_b1 , \444_b1 , \331_b1 );
not ( \331_b1 , w_854 );
and ( \588_b0 , \444_b0 , w_855 );
and ( w_854 , w_855 , \331_b0 );
or ( \589_b1 , \360_b1 , \329_b1 );
not ( \329_b1 , w_856 );
and ( \589_b0 , \360_b0 , w_857 );
and ( w_856 , w_857 , \329_b0 );
or ( \590_b1 , \588_b1 , w_859 );
not ( w_859 , w_860 );
and ( \590_b0 , \588_b0 , w_861 );
and ( w_860 ,  , w_861 );
buf ( w_859 , \589_b1 );
not ( w_859 , w_862 );
not (  , w_863 );
and ( w_862 , w_863 , \589_b0 );
or ( \591_b1 , \590_b1 , w_864 );
xor ( \591_b0 , \590_b0 , w_866 );
not ( w_866 , w_867 );
and ( w_867 , w_864 , w_865 );
buf ( w_864 , \338_b1 );
not ( w_864 , w_868 );
not ( w_865 , w_869 );
and ( w_868 , w_869 , \338_b0 );
or ( \592_b1 , \587_b1 , \591_b1 );
not ( \591_b1 , w_870 );
and ( \592_b0 , \587_b0 , w_871 );
and ( w_870 , w_871 , \591_b0 );
buf ( \593_b1 , RIb4bf588_75_b1 );
buf ( \593_b0 , RIb4bf588_75_b0 );
or ( \594_b1 , \593_b1 , \351_b1 );
not ( \351_b1 , w_872 );
and ( \594_b0 , \593_b0 , w_873 );
and ( w_872 , w_873 , \351_b0 );
or ( \595_b1 , \495_b1 , \349_b1 );
not ( \349_b1 , w_874 );
and ( \595_b0 , \495_b0 , w_875 );
and ( w_874 , w_875 , \349_b0 );
or ( \596_b1 , \594_b1 , w_877 );
not ( w_877 , w_878 );
and ( \596_b0 , \594_b0 , w_879 );
and ( w_878 ,  , w_879 );
buf ( w_877 , \595_b1 );
not ( w_877 , w_880 );
not (  , w_881 );
and ( w_880 , w_881 , \595_b0 );
or ( \597_b1 , \596_b1 , w_882 );
xor ( \597_b0 , \596_b0 , w_884 );
not ( w_884 , w_885 );
and ( w_885 , w_882 , w_883 );
buf ( w_882 , \358_b1 );
not ( w_882 , w_886 );
not ( w_883 , w_887 );
and ( w_886 , w_887 , \358_b0 );
or ( \598_b1 , \591_b1 , \597_b1 );
not ( \597_b1 , w_888 );
and ( \598_b0 , \591_b0 , w_889 );
and ( w_888 , w_889 , \597_b0 );
or ( \599_b1 , \587_b1 , \597_b1 );
not ( \597_b1 , w_890 );
and ( \599_b0 , \587_b0 , w_891 );
and ( w_890 , w_891 , \597_b0 );
or ( \601_b1 , \452_b1 , \556_b1 );
xor ( \601_b0 , \452_b0 , w_892 );
not ( w_892 , w_893 );
and ( w_893 , \556_b1 , \556_b0 );
or ( \602_b1 , \556_b1 , \558_b1 );
xor ( \602_b0 , \556_b0 , w_894 );
not ( w_894 , w_895 );
and ( w_895 , \558_b1 , \558_b0 );
buf ( \603_b1 , \602_b1 );
not ( \603_b1 , w_896 );
not ( \603_b0 , w_897 );
and ( w_896 , w_897 , \602_b0 );
or ( \604_b1 , \601_b1 , \603_b1 );
not ( \603_b1 , w_898 );
and ( \604_b0 , \601_b0 , w_899 );
and ( w_898 , w_899 , \603_b0 );
or ( \605_b1 , \159_b1 , \604_b1 );
not ( \604_b1 , w_900 );
and ( \605_b0 , \159_b0 , w_901 );
and ( w_900 , w_901 , \604_b0 );
buf ( \606_b1 , \605_b1 );
not ( \606_b1 , w_902 );
not ( \606_b0 , w_903 );
and ( w_902 , w_903 , \605_b0 );
or ( \607_b1 , \606_b1 , w_904 );
xor ( \607_b0 , \606_b0 , w_906 );
not ( w_906 , w_907 );
and ( w_907 , w_904 , w_905 );
buf ( w_904 , \561_b1 );
not ( w_904 , w_908 );
not ( w_905 , w_909 );
and ( w_908 , w_909 , \561_b0 );
or ( \608_b1 , \305_b1 , \503_b1 );
not ( \503_b1 , w_910 );
and ( \608_b0 , \305_b0 , w_911 );
and ( w_910 , w_911 , \503_b0 );
or ( \609_b1 , \315_b1 , \501_b1 );
not ( \501_b1 , w_912 );
and ( \609_b0 , \315_b0 , w_913 );
and ( w_912 , w_913 , \501_b0 );
or ( \610_b1 , \608_b1 , w_915 );
not ( w_915 , w_916 );
and ( \610_b0 , \608_b0 , w_917 );
and ( w_916 ,  , w_917 );
buf ( w_915 , \609_b1 );
not ( w_915 , w_918 );
not (  , w_919 );
and ( w_918 , w_919 , \609_b0 );
or ( \611_b1 , \610_b1 , w_920 );
xor ( \611_b0 , \610_b0 , w_922 );
not ( w_922 , w_923 );
and ( w_923 , w_920 , w_921 );
buf ( w_920 , \455_b1 );
not ( w_920 , w_924 );
not ( w_921 , w_925 );
and ( w_924 , w_925 , \455_b0 );
or ( \612_b1 , \607_b1 , \611_b1 );
not ( \611_b1 , w_926 );
and ( \612_b0 , \607_b0 , w_927 );
and ( w_926 , w_927 , \611_b0 );
or ( \613_b1 , \323_b1 , \298_b1 );
not ( \298_b1 , w_928 );
and ( \613_b0 , \323_b0 , w_929 );
and ( w_928 , w_929 , \298_b0 );
or ( \614_b1 , \333_b1 , \296_b1 );
not ( \296_b1 , w_930 );
and ( \614_b0 , \333_b0 , w_931 );
and ( w_930 , w_931 , \296_b0 );
or ( \615_b1 , \613_b1 , w_933 );
not ( w_933 , w_934 );
and ( \615_b0 , \613_b0 , w_935 );
and ( w_934 ,  , w_935 );
buf ( w_933 , \614_b1 );
not ( w_933 , w_936 );
not (  , w_937 );
and ( w_936 , w_937 , \614_b0 );
or ( \616_b1 , \615_b1 , w_938 );
xor ( \616_b0 , \615_b0 , w_940 );
not ( w_940 , w_941 );
and ( w_941 , w_938 , w_939 );
buf ( w_938 , \303_b1 );
not ( w_938 , w_942 );
not ( w_939 , w_943 );
and ( w_942 , w_943 , \303_b0 );
or ( \617_b1 , \611_b1 , \616_b1 );
not ( \616_b1 , w_944 );
and ( \617_b0 , \611_b0 , w_945 );
and ( w_944 , w_945 , \616_b0 );
or ( \618_b1 , \607_b1 , \616_b1 );
not ( \616_b1 , w_946 );
and ( \618_b0 , \607_b0 , w_947 );
and ( w_946 , w_947 , \616_b0 );
or ( \620_b1 , \600_b1 , \619_b1 );
not ( \619_b1 , w_948 );
and ( \620_b0 , \600_b0 , w_949 );
and ( w_948 , w_949 , \619_b0 );
buf ( \621_b1 , RIb4bf510_76_b1 );
buf ( \621_b0 , RIb4bf510_76_b0 );
or ( \622_b1 , \621_b1 , \345_b1 );
not ( \345_b1 , w_950 );
and ( \622_b0 , \621_b0 , w_951 );
and ( w_950 , w_951 , \345_b0 );
buf ( \623_b1 , \622_b1 );
buf ( \623_b0 , \622_b0 );
or ( \624_b1 , \619_b1 , \623_b1 );
not ( \623_b1 , w_952 );
and ( \624_b0 , \619_b0 , w_953 );
and ( w_952 , w_953 , \623_b0 );
or ( \625_b1 , \600_b1 , \623_b1 );
not ( \623_b1 , w_954 );
and ( \625_b0 , \600_b0 , w_955 );
and ( w_954 , w_955 , \623_b0 );
or ( \627_b1 , \593_b1 , \345_b1 );
not ( \345_b1 , w_956 );
and ( \627_b0 , \593_b0 , w_957 );
and ( w_956 , w_957 , \345_b0 );
or ( \628_b1 , \542_b1 , \546_b1 );
xor ( \628_b0 , \542_b0 , w_958 );
not ( w_958 , w_959 );
and ( w_959 , \546_b1 , \546_b0 );
or ( \629_b1 , \628_b1 , \551_b1 );
xor ( \629_b0 , \628_b0 , w_960 );
not ( w_960 , w_961 );
and ( w_961 , \551_b1 , \551_b0 );
or ( \630_b1 , \627_b1 , \629_b1 );
not ( \629_b1 , w_962 );
and ( \630_b0 , \627_b0 , w_963 );
and ( w_962 , w_963 , \629_b0 );
or ( \631_b1 , \562_b1 , \566_b1 );
xor ( \631_b0 , \562_b0 , w_964 );
not ( w_964 , w_965 );
and ( w_965 , \566_b1 , \566_b0 );
or ( \632_b1 , \631_b1 , \571_b1 );
xor ( \632_b0 , \631_b0 , w_966 );
not ( w_966 , w_967 );
and ( w_967 , \571_b1 , \571_b0 );
or ( \633_b1 , \629_b1 , \632_b1 );
not ( \632_b1 , w_968 );
and ( \633_b0 , \629_b0 , w_969 );
and ( w_968 , w_969 , \632_b0 );
or ( \634_b1 , \627_b1 , \632_b1 );
not ( \632_b1 , w_970 );
and ( \634_b0 , \627_b0 , w_971 );
and ( w_970 , w_971 , \632_b0 );
or ( \636_b1 , \626_b1 , \635_b1 );
not ( \635_b1 , w_972 );
and ( \636_b0 , \626_b0 , w_973 );
and ( w_972 , w_973 , \635_b0 );
or ( \637_b1 , \489_b1 , \493_b1 );
xor ( \637_b0 , \489_b0 , w_974 );
not ( w_974 , w_975 );
and ( w_975 , \493_b1 , \493_b0 );
or ( \638_b1 , \637_b1 , \496_b1 );
xor ( \638_b0 , \637_b0 , w_976 );
not ( w_976 , w_977 );
and ( w_977 , \496_b1 , \496_b0 );
or ( \639_b1 , \635_b1 , \638_b1 );
not ( \638_b1 , w_978 );
and ( \639_b0 , \635_b0 , w_979 );
and ( w_978 , w_979 , \638_b0 );
or ( \640_b1 , \626_b1 , \638_b1 );
not ( \638_b1 , w_980 );
and ( \640_b0 , \626_b0 , w_981 );
and ( w_980 , w_981 , \638_b0 );
or ( \642_b1 , \506_b1 , \510_b1 );
xor ( \642_b0 , \506_b0 , w_982 );
not ( w_982 , w_983 );
and ( w_983 , \510_b1 , \510_b0 );
or ( \643_b1 , \642_b1 , \515_b1 );
xor ( \643_b0 , \642_b0 , w_984 );
not ( w_984 , w_985 );
and ( w_985 , \515_b1 , \515_b0 );
or ( \644_b1 , \554_b1 , w_986 );
xor ( \644_b0 , \554_b0 , w_988 );
not ( w_988 , w_989 );
and ( w_989 , w_986 , w_987 );
buf ( w_986 , \574_b1 );
not ( w_986 , w_990 );
not ( w_987 , w_991 );
and ( w_990 , w_991 , \574_b0 );
or ( \645_b1 , \643_b1 , \644_b1 );
not ( \644_b1 , w_992 );
and ( \645_b0 , \643_b0 , w_993 );
and ( w_992 , w_993 , \644_b0 );
or ( \646_b1 , \641_b1 , \645_b1 );
not ( \645_b1 , w_994 );
and ( \646_b0 , \641_b0 , w_995 );
and ( w_994 , w_995 , \645_b0 );
or ( \647_b1 , \575_b1 , \577_b1 );
xor ( \647_b0 , \575_b0 , w_996 );
not ( w_996 , w_997 );
and ( w_997 , \577_b1 , \577_b0 );
or ( \648_b1 , \647_b1 , \580_b1 );
xor ( \648_b0 , \647_b0 , w_998 );
not ( w_998 , w_999 );
and ( w_999 , \580_b1 , \580_b0 );
or ( \649_b1 , \645_b1 , \648_b1 );
not ( \648_b1 , w_1000 );
and ( \649_b0 , \645_b0 , w_1001 );
and ( w_1000 , w_1001 , \648_b0 );
or ( \650_b1 , \641_b1 , \648_b1 );
not ( \648_b1 , w_1002 );
and ( \650_b0 , \641_b0 , w_1003 );
and ( w_1002 , w_1003 , \648_b0 );
or ( \652_b1 , \583_b1 , \651_b1 );
not ( \651_b1 , w_1004 );
and ( \652_b0 , \583_b0 , w_1005 );
and ( w_1004 , w_1005 , \651_b0 );
or ( \653_b1 , \524_b1 , \526_b1 );
xor ( \653_b0 , \524_b0 , w_1006 );
not ( w_1006 , w_1007 );
and ( w_1007 , \526_b1 , \526_b0 );
or ( \654_b1 , \653_b1 , \529_b1 );
xor ( \654_b0 , \653_b0 , w_1008 );
not ( w_1008 , w_1009 );
and ( w_1009 , \529_b1 , \529_b0 );
or ( \655_b1 , \651_b1 , \654_b1 );
not ( \654_b1 , w_1010 );
and ( \655_b0 , \651_b0 , w_1011 );
and ( w_1010 , w_1011 , \654_b0 );
or ( \656_b1 , \583_b1 , \654_b1 );
not ( \654_b1 , w_1012 );
and ( \656_b0 , \583_b0 , w_1013 );
and ( w_1012 , w_1013 , \654_b0 );
or ( \658_b1 , \538_b1 , \657_b1 );
not ( \657_b1 , w_1014 );
and ( \658_b0 , \538_b0 , w_1015 );
and ( w_1014 , w_1015 , \657_b0 );
or ( \659_b1 , \538_b1 , \657_b1 );
xor ( \659_b0 , \538_b0 , w_1016 );
not ( w_1016 , w_1017 );
and ( w_1017 , \657_b1 , \657_b0 );
or ( \660_b1 , \583_b1 , \651_b1 );
xor ( \660_b0 , \583_b0 , w_1018 );
not ( w_1018 , w_1019 );
and ( w_1019 , \651_b1 , \651_b0 );
or ( \661_b1 , \660_b1 , \654_b1 );
xor ( \661_b0 , \660_b0 , w_1020 );
not ( w_1020 , w_1021 );
and ( w_1021 , \654_b1 , \654_b0 );
and ( \662_nR136_b1 , RIb4c32f0_46_b1 , w_1022 );
xor ( w_1022 , RIb4c32f0_46_b0 , \288_b1 );
not ( \288_b1 , w_1023 );
and ( \662_nR136_b0 , w_1023 , \288_b0 );
buf ( \663_b1 , \662_nR136_b1 );
buf ( \663_b0 , \662_nR136_b0 );
and ( \664_nR135_b1 , RIb4c3278_47_b1 , w_1024 );
xor ( w_1024 , RIb4c3278_47_b0 , \288_b1 );
not ( \288_b1 , w_1025 );
and ( \664_nR135_b0 , w_1025 , \288_b0 );
buf ( \665_b1 , \664_nR135_b1 );
buf ( \665_b0 , \664_nR135_b0 );
or ( \666_b1 , \663_b1 , \665_b1 );
not ( \665_b1 , w_1026 );
and ( \666_b0 , \663_b0 , w_1027 );
and ( w_1026 , w_1027 , \665_b0 );
buf ( \667_b1 , \666_b1 );
not ( \667_b1 , w_1028 );
not ( \667_b0 , w_1029 );
and ( w_1028 , w_1029 , \666_b0 );
or ( \668_b1 , \558_b1 , \667_b1 );
not ( \667_b1 , w_1030 );
and ( \668_b0 , \558_b0 , w_1031 );
and ( w_1030 , w_1031 , \667_b0 );
buf ( \669_b1 , \668_b1 );
not ( \669_b1 , w_1032 );
not ( \669_b0 , w_1033 );
and ( w_1032 , w_1033 , \668_b0 );
or ( \670_b1 , \315_b1 , \604_b1 );
not ( \604_b1 , w_1034 );
and ( \670_b0 , \315_b0 , w_1035 );
and ( w_1034 , w_1035 , \604_b0 );
or ( \671_b1 , \159_b1 , \602_b1 );
not ( \602_b1 , w_1036 );
and ( \671_b0 , \159_b0 , w_1037 );
and ( w_1036 , w_1037 , \602_b0 );
or ( \672_b1 , \670_b1 , w_1039 );
not ( w_1039 , w_1040 );
and ( \672_b0 , \670_b0 , w_1041 );
and ( w_1040 ,  , w_1041 );
buf ( w_1039 , \671_b1 );
not ( w_1039 , w_1042 );
not (  , w_1043 );
and ( w_1042 , w_1043 , \671_b0 );
or ( \673_b1 , \672_b1 , w_1044 );
xor ( \673_b0 , \672_b0 , w_1046 );
not ( w_1046 , w_1047 );
and ( w_1047 , w_1044 , w_1045 );
buf ( w_1044 , \561_b1 );
not ( w_1044 , w_1048 );
not ( w_1045 , w_1049 );
and ( w_1048 , w_1049 , \561_b0 );
or ( \674_b1 , \669_b1 , \673_b1 );
not ( \673_b1 , w_1050 );
and ( \674_b0 , \669_b0 , w_1051 );
and ( w_1050 , w_1051 , \673_b0 );
or ( \675_b1 , \333_b1 , \503_b1 );
not ( \503_b1 , w_1052 );
and ( \675_b0 , \333_b0 , w_1053 );
and ( w_1052 , w_1053 , \503_b0 );
or ( \676_b1 , \305_b1 , \501_b1 );
not ( \501_b1 , w_1054 );
and ( \676_b0 , \305_b0 , w_1055 );
and ( w_1054 , w_1055 , \501_b0 );
or ( \677_b1 , \675_b1 , w_1057 );
not ( w_1057 , w_1058 );
and ( \677_b0 , \675_b0 , w_1059 );
and ( w_1058 ,  , w_1059 );
buf ( w_1057 , \676_b1 );
not ( w_1057 , w_1060 );
not (  , w_1061 );
and ( w_1060 , w_1061 , \676_b0 );
or ( \678_b1 , \677_b1 , w_1062 );
xor ( \678_b0 , \677_b0 , w_1064 );
not ( w_1064 , w_1065 );
and ( w_1065 , w_1062 , w_1063 );
buf ( w_1062 , \455_b1 );
not ( w_1062 , w_1066 );
not ( w_1063 , w_1067 );
and ( w_1066 , w_1067 , \455_b0 );
or ( \679_b1 , \673_b1 , \678_b1 );
not ( \678_b1 , w_1068 );
and ( \679_b0 , \673_b0 , w_1069 );
and ( w_1068 , w_1069 , \678_b0 );
or ( \680_b1 , \669_b1 , \678_b1 );
not ( \678_b1 , w_1070 );
and ( \680_b0 , \669_b0 , w_1071 );
and ( w_1070 , w_1071 , \678_b0 );
or ( \682_b1 , \353_b1 , \298_b1 );
not ( \298_b1 , w_1072 );
and ( \682_b0 , \353_b0 , w_1073 );
and ( w_1072 , w_1073 , \298_b0 );
or ( \683_b1 , \323_b1 , \296_b1 );
not ( \296_b1 , w_1074 );
and ( \683_b0 , \323_b0 , w_1075 );
and ( w_1074 , w_1075 , \296_b0 );
or ( \684_b1 , \682_b1 , w_1077 );
not ( w_1077 , w_1078 );
and ( \684_b0 , \682_b0 , w_1079 );
and ( w_1078 ,  , w_1079 );
buf ( w_1077 , \683_b1 );
not ( w_1077 , w_1080 );
not (  , w_1081 );
and ( w_1080 , w_1081 , \683_b0 );
or ( \685_b1 , \684_b1 , w_1082 );
xor ( \685_b0 , \684_b0 , w_1084 );
not ( w_1084 , w_1085 );
and ( w_1085 , w_1082 , w_1083 );
buf ( w_1082 , \303_b1 );
not ( w_1082 , w_1086 );
not ( w_1083 , w_1087 );
and ( w_1086 , w_1087 , \303_b0 );
or ( \686_b1 , \360_b1 , \313_b1 );
not ( \313_b1 , w_1088 );
and ( \686_b0 , \360_b0 , w_1089 );
and ( w_1088 , w_1089 , \313_b0 );
or ( \687_b1 , \343_b1 , \311_b1 );
not ( \311_b1 , w_1090 );
and ( \687_b0 , \343_b0 , w_1091 );
and ( w_1090 , w_1091 , \311_b0 );
or ( \688_b1 , \686_b1 , w_1093 );
not ( w_1093 , w_1094 );
and ( \688_b0 , \686_b0 , w_1095 );
and ( w_1094 ,  , w_1095 );
buf ( w_1093 , \687_b1 );
not ( w_1093 , w_1096 );
not (  , w_1097 );
and ( w_1096 , w_1097 , \687_b0 );
or ( \689_b1 , \688_b1 , w_1098 );
xor ( \689_b0 , \688_b0 , w_1100 );
not ( w_1100 , w_1101 );
and ( w_1101 , w_1098 , w_1099 );
buf ( w_1098 , \320_b1 );
not ( w_1098 , w_1102 );
not ( w_1099 , w_1103 );
and ( w_1102 , w_1103 , \320_b0 );
or ( \690_b1 , \685_b1 , \689_b1 );
not ( \689_b1 , w_1104 );
and ( \690_b0 , \685_b0 , w_1105 );
and ( w_1104 , w_1105 , \689_b0 );
or ( \691_b1 , \495_b1 , \331_b1 );
not ( \331_b1 , w_1106 );
and ( \691_b0 , \495_b0 , w_1107 );
and ( w_1106 , w_1107 , \331_b0 );
or ( \692_b1 , \444_b1 , \329_b1 );
not ( \329_b1 , w_1108 );
and ( \692_b0 , \444_b0 , w_1109 );
and ( w_1108 , w_1109 , \329_b0 );
or ( \693_b1 , \691_b1 , w_1111 );
not ( w_1111 , w_1112 );
and ( \693_b0 , \691_b0 , w_1113 );
and ( w_1112 ,  , w_1113 );
buf ( w_1111 , \692_b1 );
not ( w_1111 , w_1114 );
not (  , w_1115 );
and ( w_1114 , w_1115 , \692_b0 );
or ( \694_b1 , \693_b1 , w_1116 );
xor ( \694_b0 , \693_b0 , w_1118 );
not ( w_1118 , w_1119 );
and ( w_1119 , w_1116 , w_1117 );
buf ( w_1116 , \338_b1 );
not ( w_1116 , w_1120 );
not ( w_1117 , w_1121 );
and ( w_1120 , w_1121 , \338_b0 );
or ( \695_b1 , \689_b1 , \694_b1 );
not ( \694_b1 , w_1122 );
and ( \695_b0 , \689_b0 , w_1123 );
and ( w_1122 , w_1123 , \694_b0 );
or ( \696_b1 , \685_b1 , \694_b1 );
not ( \694_b1 , w_1124 );
and ( \696_b0 , \685_b0 , w_1125 );
and ( w_1124 , w_1125 , \694_b0 );
or ( \698_b1 , \681_b1 , \697_b1 );
not ( \697_b1 , w_1126 );
and ( \698_b0 , \681_b0 , w_1127 );
and ( w_1126 , w_1127 , \697_b0 );
or ( \699_b1 , \621_b1 , \351_b1 );
not ( \351_b1 , w_1128 );
and ( \699_b0 , \621_b0 , w_1129 );
and ( w_1128 , w_1129 , \351_b0 );
or ( \700_b1 , \593_b1 , \349_b1 );
not ( \349_b1 , w_1130 );
and ( \700_b0 , \593_b0 , w_1131 );
and ( w_1130 , w_1131 , \349_b0 );
or ( \701_b1 , \699_b1 , w_1133 );
not ( w_1133 , w_1134 );
and ( \701_b0 , \699_b0 , w_1135 );
and ( w_1134 ,  , w_1135 );
buf ( w_1133 , \700_b1 );
not ( w_1133 , w_1136 );
not (  , w_1137 );
and ( w_1136 , w_1137 , \700_b0 );
or ( \702_b1 , \701_b1 , w_1138 );
xor ( \702_b0 , \701_b0 , w_1140 );
not ( w_1140 , w_1141 );
and ( w_1141 , w_1138 , w_1139 );
buf ( w_1138 , \358_b1 );
not ( w_1138 , w_1142 );
not ( w_1139 , w_1143 );
and ( w_1142 , w_1143 , \358_b0 );
buf ( \703_b1 , RIb4bf498_77_b1 );
buf ( \703_b0 , RIb4bf498_77_b0 );
or ( \704_b1 , \703_b1 , \345_b1 );
not ( \345_b1 , w_1144 );
and ( \704_b0 , \703_b0 , w_1145 );
and ( w_1144 , w_1145 , \345_b0 );
or ( \705_b1 , \702_b1 , \704_b1 );
not ( \704_b1 , w_1146 );
and ( \705_b0 , \702_b0 , w_1147 );
and ( w_1146 , w_1147 , \704_b0 );
or ( \706_b1 , \697_b1 , \705_b1 );
not ( \705_b1 , w_1148 );
and ( \706_b0 , \697_b0 , w_1149 );
and ( w_1148 , w_1149 , \705_b0 );
or ( \707_b1 , \681_b1 , \705_b1 );
not ( \705_b1 , w_1150 );
and ( \707_b0 , \681_b0 , w_1151 );
and ( w_1150 , w_1151 , \705_b0 );
or ( \709_b1 , \587_b1 , \591_b1 );
xor ( \709_b0 , \587_b0 , w_1152 );
not ( w_1152 , w_1153 );
and ( w_1153 , \591_b1 , \591_b0 );
or ( \710_b1 , \709_b1 , \597_b1 );
xor ( \710_b0 , \709_b0 , w_1154 );
not ( w_1154 , w_1155 );
and ( w_1155 , \597_b1 , \597_b0 );
or ( \711_b1 , \607_b1 , \611_b1 );
xor ( \711_b0 , \607_b0 , w_1156 );
not ( w_1156 , w_1157 );
and ( w_1157 , \611_b1 , \611_b0 );
or ( \712_b1 , \711_b1 , \616_b1 );
xor ( \712_b0 , \711_b0 , w_1158 );
not ( w_1158 , w_1159 );
and ( w_1159 , \616_b1 , \616_b0 );
or ( \713_b1 , \710_b1 , \712_b1 );
not ( \712_b1 , w_1160 );
and ( \713_b0 , \710_b0 , w_1161 );
and ( w_1160 , w_1161 , \712_b0 );
buf ( \714_b1 , \622_b1 );
not ( \714_b1 , w_1162 );
not ( \714_b0 , w_1163 );
and ( w_1162 , w_1163 , \622_b0 );
or ( \715_b1 , \712_b1 , \714_b1 );
not ( \714_b1 , w_1164 );
and ( \715_b0 , \712_b0 , w_1165 );
and ( w_1164 , w_1165 , \714_b0 );
or ( \716_b1 , \710_b1 , \714_b1 );
not ( \714_b1 , w_1166 );
and ( \716_b0 , \710_b0 , w_1167 );
and ( w_1166 , w_1167 , \714_b0 );
or ( \718_b1 , \708_b1 , \717_b1 );
not ( \717_b1 , w_1168 );
and ( \718_b0 , \708_b0 , w_1169 );
and ( w_1168 , w_1169 , \717_b0 );
or ( \719_b1 , \627_b1 , \629_b1 );
xor ( \719_b0 , \627_b0 , w_1170 );
not ( w_1170 , w_1171 );
and ( w_1171 , \629_b1 , \629_b0 );
or ( \720_b1 , \719_b1 , \632_b1 );
xor ( \720_b0 , \719_b0 , w_1172 );
not ( w_1172 , w_1173 );
and ( w_1173 , \632_b1 , \632_b0 );
or ( \721_b1 , \717_b1 , \720_b1 );
not ( \720_b1 , w_1174 );
and ( \721_b0 , \717_b0 , w_1175 );
and ( w_1174 , w_1175 , \720_b0 );
or ( \722_b1 , \708_b1 , \720_b1 );
not ( \720_b1 , w_1176 );
and ( \722_b0 , \708_b0 , w_1177 );
and ( w_1176 , w_1177 , \720_b0 );
or ( \724_b1 , \626_b1 , \635_b1 );
xor ( \724_b0 , \626_b0 , w_1178 );
not ( w_1178 , w_1179 );
and ( w_1179 , \635_b1 , \635_b0 );
or ( \725_b1 , \724_b1 , \638_b1 );
xor ( \725_b0 , \724_b0 , w_1180 );
not ( w_1180 , w_1181 );
and ( w_1181 , \638_b1 , \638_b0 );
or ( \726_b1 , \723_b1 , \725_b1 );
not ( \725_b1 , w_1182 );
and ( \726_b0 , \723_b0 , w_1183 );
and ( w_1182 , w_1183 , \725_b0 );
or ( \727_b1 , \643_b1 , \644_b1 );
xor ( \727_b0 , \643_b0 , w_1184 );
not ( w_1184 , w_1185 );
and ( w_1185 , \644_b1 , \644_b0 );
or ( \728_b1 , \725_b1 , \727_b1 );
not ( \727_b1 , w_1186 );
and ( \728_b0 , \725_b0 , w_1187 );
and ( w_1186 , w_1187 , \727_b0 );
or ( \729_b1 , \723_b1 , \727_b1 );
not ( \727_b1 , w_1188 );
and ( \729_b0 , \723_b0 , w_1189 );
and ( w_1188 , w_1189 , \727_b0 );
or ( \731_b1 , \641_b1 , \645_b1 );
xor ( \731_b0 , \641_b0 , w_1190 );
not ( w_1190 , w_1191 );
and ( w_1191 , \645_b1 , \645_b0 );
or ( \732_b1 , \731_b1 , \648_b1 );
xor ( \732_b0 , \731_b0 , w_1192 );
not ( w_1192 , w_1193 );
and ( w_1193 , \648_b1 , \648_b0 );
or ( \733_b1 , \730_b1 , \732_b1 );
not ( \732_b1 , w_1194 );
and ( \733_b0 , \730_b0 , w_1195 );
and ( w_1194 , w_1195 , \732_b0 );
or ( \734_b1 , \661_b1 , \733_b1 );
not ( \733_b1 , w_1196 );
and ( \734_b0 , \661_b0 , w_1197 );
and ( w_1196 , w_1197 , \733_b0 );
or ( \735_b1 , \661_b1 , \733_b1 );
xor ( \735_b0 , \661_b0 , w_1198 );
not ( w_1198 , w_1199 );
and ( w_1199 , \733_b1 , \733_b0 );
or ( \736_b1 , \730_b1 , \732_b1 );
xor ( \736_b0 , \730_b0 , w_1200 );
not ( w_1200 , w_1201 );
and ( w_1201 , \732_b1 , \732_b0 );
or ( \737_b1 , \558_b1 , \663_b1 );
xor ( \737_b0 , \558_b0 , w_1202 );
not ( w_1202 , w_1203 );
and ( w_1203 , \663_b1 , \663_b0 );
or ( \738_b1 , \663_b1 , \665_b1 );
xor ( \738_b0 , \663_b0 , w_1204 );
not ( w_1204 , w_1205 );
and ( w_1205 , \665_b1 , \665_b0 );
buf ( \739_b1 , \738_b1 );
not ( \739_b1 , w_1206 );
not ( \739_b0 , w_1207 );
and ( w_1206 , w_1207 , \738_b0 );
or ( \740_b1 , \737_b1 , \739_b1 );
not ( \739_b1 , w_1208 );
and ( \740_b0 , \737_b0 , w_1209 );
and ( w_1208 , w_1209 , \739_b0 );
or ( \741_b1 , \159_b1 , \740_b1 );
not ( \740_b1 , w_1210 );
and ( \741_b0 , \159_b0 , w_1211 );
and ( w_1210 , w_1211 , \740_b0 );
buf ( \742_b1 , \741_b1 );
not ( \742_b1 , w_1212 );
not ( \742_b0 , w_1213 );
and ( w_1212 , w_1213 , \741_b0 );
or ( \743_b1 , \742_b1 , w_1214 );
xor ( \743_b0 , \742_b0 , w_1216 );
not ( w_1216 , w_1217 );
and ( w_1217 , w_1214 , w_1215 );
buf ( w_1214 , \668_b1 );
not ( w_1214 , w_1218 );
not ( w_1215 , w_1219 );
and ( w_1218 , w_1219 , \668_b0 );
or ( \744_b1 , \305_b1 , \604_b1 );
not ( \604_b1 , w_1220 );
and ( \744_b0 , \305_b0 , w_1221 );
and ( w_1220 , w_1221 , \604_b0 );
or ( \745_b1 , \315_b1 , \602_b1 );
not ( \602_b1 , w_1222 );
and ( \745_b0 , \315_b0 , w_1223 );
and ( w_1222 , w_1223 , \602_b0 );
or ( \746_b1 , \744_b1 , w_1225 );
not ( w_1225 , w_1226 );
and ( \746_b0 , \744_b0 , w_1227 );
and ( w_1226 ,  , w_1227 );
buf ( w_1225 , \745_b1 );
not ( w_1225 , w_1228 );
not (  , w_1229 );
and ( w_1228 , w_1229 , \745_b0 );
or ( \747_b1 , \746_b1 , w_1230 );
xor ( \747_b0 , \746_b0 , w_1232 );
not ( w_1232 , w_1233 );
and ( w_1233 , w_1230 , w_1231 );
buf ( w_1230 , \561_b1 );
not ( w_1230 , w_1234 );
not ( w_1231 , w_1235 );
and ( w_1234 , w_1235 , \561_b0 );
or ( \748_b1 , \743_b1 , \747_b1 );
not ( \747_b1 , w_1236 );
and ( \748_b0 , \743_b0 , w_1237 );
and ( w_1236 , w_1237 , \747_b0 );
or ( \749_b1 , \323_b1 , \503_b1 );
not ( \503_b1 , w_1238 );
and ( \749_b0 , \323_b0 , w_1239 );
and ( w_1238 , w_1239 , \503_b0 );
or ( \750_b1 , \333_b1 , \501_b1 );
not ( \501_b1 , w_1240 );
and ( \750_b0 , \333_b0 , w_1241 );
and ( w_1240 , w_1241 , \501_b0 );
or ( \751_b1 , \749_b1 , w_1243 );
not ( w_1243 , w_1244 );
and ( \751_b0 , \749_b0 , w_1245 );
and ( w_1244 ,  , w_1245 );
buf ( w_1243 , \750_b1 );
not ( w_1243 , w_1246 );
not (  , w_1247 );
and ( w_1246 , w_1247 , \750_b0 );
or ( \752_b1 , \751_b1 , w_1248 );
xor ( \752_b0 , \751_b0 , w_1250 );
not ( w_1250 , w_1251 );
and ( w_1251 , w_1248 , w_1249 );
buf ( w_1248 , \455_b1 );
not ( w_1248 , w_1252 );
not ( w_1249 , w_1253 );
and ( w_1252 , w_1253 , \455_b0 );
or ( \753_b1 , \747_b1 , \752_b1 );
not ( \752_b1 , w_1254 );
and ( \753_b0 , \747_b0 , w_1255 );
and ( w_1254 , w_1255 , \752_b0 );
or ( \754_b1 , \743_b1 , \752_b1 );
not ( \752_b1 , w_1256 );
and ( \754_b0 , \743_b0 , w_1257 );
and ( w_1256 , w_1257 , \752_b0 );
or ( \756_b1 , \343_b1 , \298_b1 );
not ( \298_b1 , w_1258 );
and ( \756_b0 , \343_b0 , w_1259 );
and ( w_1258 , w_1259 , \298_b0 );
or ( \757_b1 , \353_b1 , \296_b1 );
not ( \296_b1 , w_1260 );
and ( \757_b0 , \353_b0 , w_1261 );
and ( w_1260 , w_1261 , \296_b0 );
or ( \758_b1 , \756_b1 , w_1263 );
not ( w_1263 , w_1264 );
and ( \758_b0 , \756_b0 , w_1265 );
and ( w_1264 ,  , w_1265 );
buf ( w_1263 , \757_b1 );
not ( w_1263 , w_1266 );
not (  , w_1267 );
and ( w_1266 , w_1267 , \757_b0 );
or ( \759_b1 , \758_b1 , w_1268 );
xor ( \759_b0 , \758_b0 , w_1270 );
not ( w_1270 , w_1271 );
and ( w_1271 , w_1268 , w_1269 );
buf ( w_1268 , \303_b1 );
not ( w_1268 , w_1272 );
not ( w_1269 , w_1273 );
and ( w_1272 , w_1273 , \303_b0 );
or ( \760_b1 , \444_b1 , \313_b1 );
not ( \313_b1 , w_1274 );
and ( \760_b0 , \444_b0 , w_1275 );
and ( w_1274 , w_1275 , \313_b0 );
or ( \761_b1 , \360_b1 , \311_b1 );
not ( \311_b1 , w_1276 );
and ( \761_b0 , \360_b0 , w_1277 );
and ( w_1276 , w_1277 , \311_b0 );
or ( \762_b1 , \760_b1 , w_1279 );
not ( w_1279 , w_1280 );
and ( \762_b0 , \760_b0 , w_1281 );
and ( w_1280 ,  , w_1281 );
buf ( w_1279 , \761_b1 );
not ( w_1279 , w_1282 );
not (  , w_1283 );
and ( w_1282 , w_1283 , \761_b0 );
or ( \763_b1 , \762_b1 , w_1284 );
xor ( \763_b0 , \762_b0 , w_1286 );
not ( w_1286 , w_1287 );
and ( w_1287 , w_1284 , w_1285 );
buf ( w_1284 , \320_b1 );
not ( w_1284 , w_1288 );
not ( w_1285 , w_1289 );
and ( w_1288 , w_1289 , \320_b0 );
or ( \764_b1 , \759_b1 , \763_b1 );
not ( \763_b1 , w_1290 );
and ( \764_b0 , \759_b0 , w_1291 );
and ( w_1290 , w_1291 , \763_b0 );
or ( \765_b1 , \593_b1 , \331_b1 );
not ( \331_b1 , w_1292 );
and ( \765_b0 , \593_b0 , w_1293 );
and ( w_1292 , w_1293 , \331_b0 );
or ( \766_b1 , \495_b1 , \329_b1 );
not ( \329_b1 , w_1294 );
and ( \766_b0 , \495_b0 , w_1295 );
and ( w_1294 , w_1295 , \329_b0 );
or ( \767_b1 , \765_b1 , w_1297 );
not ( w_1297 , w_1298 );
and ( \767_b0 , \765_b0 , w_1299 );
and ( w_1298 ,  , w_1299 );
buf ( w_1297 , \766_b1 );
not ( w_1297 , w_1300 );
not (  , w_1301 );
and ( w_1300 , w_1301 , \766_b0 );
or ( \768_b1 , \767_b1 , w_1302 );
xor ( \768_b0 , \767_b0 , w_1304 );
not ( w_1304 , w_1305 );
and ( w_1305 , w_1302 , w_1303 );
buf ( w_1302 , \338_b1 );
not ( w_1302 , w_1306 );
not ( w_1303 , w_1307 );
and ( w_1306 , w_1307 , \338_b0 );
or ( \769_b1 , \763_b1 , \768_b1 );
not ( \768_b1 , w_1308 );
and ( \769_b0 , \763_b0 , w_1309 );
and ( w_1308 , w_1309 , \768_b0 );
or ( \770_b1 , \759_b1 , \768_b1 );
not ( \768_b1 , w_1310 );
and ( \770_b0 , \759_b0 , w_1311 );
and ( w_1310 , w_1311 , \768_b0 );
or ( \772_b1 , \755_b1 , \771_b1 );
not ( \771_b1 , w_1312 );
and ( \772_b0 , \755_b0 , w_1313 );
and ( w_1312 , w_1313 , \771_b0 );
or ( \773_b1 , \703_b1 , \351_b1 );
not ( \351_b1 , w_1314 );
and ( \773_b0 , \703_b0 , w_1315 );
and ( w_1314 , w_1315 , \351_b0 );
or ( \774_b1 , \621_b1 , \349_b1 );
not ( \349_b1 , w_1316 );
and ( \774_b0 , \621_b0 , w_1317 );
and ( w_1316 , w_1317 , \349_b0 );
or ( \775_b1 , \773_b1 , w_1319 );
not ( w_1319 , w_1320 );
and ( \775_b0 , \773_b0 , w_1321 );
and ( w_1320 ,  , w_1321 );
buf ( w_1319 , \774_b1 );
not ( w_1319 , w_1322 );
not (  , w_1323 );
and ( w_1322 , w_1323 , \774_b0 );
or ( \776_b1 , \775_b1 , w_1324 );
xor ( \776_b0 , \775_b0 , w_1326 );
not ( w_1326 , w_1327 );
and ( w_1327 , w_1324 , w_1325 );
buf ( w_1324 , \358_b1 );
not ( w_1324 , w_1328 );
not ( w_1325 , w_1329 );
and ( w_1328 , w_1329 , \358_b0 );
buf ( \777_b1 , RIb4bf420_78_b1 );
buf ( \777_b0 , RIb4bf420_78_b0 );
or ( \778_b1 , \777_b1 , \345_b1 );
not ( \345_b1 , w_1330 );
and ( \778_b0 , \777_b0 , w_1331 );
and ( w_1330 , w_1331 , \345_b0 );
or ( \779_b1 , \776_b1 , w_1332 );
or ( \779_b0 , \776_b0 , \778_b0 );
not ( \778_b0 , w_1333 );
and ( w_1333 , w_1332 , \778_b1 );
or ( \780_b1 , \771_b1 , \779_b1 );
not ( \779_b1 , w_1334 );
and ( \780_b0 , \771_b0 , w_1335 );
and ( w_1334 , w_1335 , \779_b0 );
or ( \781_b1 , \755_b1 , \779_b1 );
not ( \779_b1 , w_1336 );
and ( \781_b0 , \755_b0 , w_1337 );
and ( w_1336 , w_1337 , \779_b0 );
or ( \783_b1 , \669_b1 , \673_b1 );
xor ( \783_b0 , \669_b0 , w_1338 );
not ( w_1338 , w_1339 );
and ( w_1339 , \673_b1 , \673_b0 );
or ( \784_b1 , \783_b1 , \678_b1 );
xor ( \784_b0 , \783_b0 , w_1340 );
not ( w_1340 , w_1341 );
and ( w_1341 , \678_b1 , \678_b0 );
or ( \785_b1 , \685_b1 , \689_b1 );
xor ( \785_b0 , \685_b0 , w_1342 );
not ( w_1342 , w_1343 );
and ( w_1343 , \689_b1 , \689_b0 );
or ( \786_b1 , \785_b1 , \694_b1 );
xor ( \786_b0 , \785_b0 , w_1344 );
not ( w_1344 , w_1345 );
and ( w_1345 , \694_b1 , \694_b0 );
or ( \787_b1 , \784_b1 , \786_b1 );
not ( \786_b1 , w_1346 );
and ( \787_b0 , \784_b0 , w_1347 );
and ( w_1346 , w_1347 , \786_b0 );
or ( \788_b1 , \702_b1 , \704_b1 );
xor ( \788_b0 , \702_b0 , w_1348 );
not ( w_1348 , w_1349 );
and ( w_1349 , \704_b1 , \704_b0 );
or ( \789_b1 , \786_b1 , \788_b1 );
not ( \788_b1 , w_1350 );
and ( \789_b0 , \786_b0 , w_1351 );
and ( w_1350 , w_1351 , \788_b0 );
or ( \790_b1 , \784_b1 , \788_b1 );
not ( \788_b1 , w_1352 );
and ( \790_b0 , \784_b0 , w_1353 );
and ( w_1352 , w_1353 , \788_b0 );
or ( \792_b1 , \782_b1 , \791_b1 );
not ( \791_b1 , w_1354 );
and ( \792_b0 , \782_b0 , w_1355 );
and ( w_1354 , w_1355 , \791_b0 );
or ( \793_b1 , \710_b1 , \712_b1 );
xor ( \793_b0 , \710_b0 , w_1356 );
not ( w_1356 , w_1357 );
and ( w_1357 , \712_b1 , \712_b0 );
or ( \794_b1 , \793_b1 , \714_b1 );
xor ( \794_b0 , \793_b0 , w_1358 );
not ( w_1358 , w_1359 );
and ( w_1359 , \714_b1 , \714_b0 );
or ( \795_b1 , \791_b1 , \794_b1 );
not ( \794_b1 , w_1360 );
and ( \795_b0 , \791_b0 , w_1361 );
and ( w_1360 , w_1361 , \794_b0 );
or ( \796_b1 , \782_b1 , \794_b1 );
not ( \794_b1 , w_1362 );
and ( \796_b0 , \782_b0 , w_1363 );
and ( w_1362 , w_1363 , \794_b0 );
or ( \798_b1 , \600_b1 , \619_b1 );
xor ( \798_b0 , \600_b0 , w_1364 );
not ( w_1364 , w_1365 );
and ( w_1365 , \619_b1 , \619_b0 );
or ( \799_b1 , \798_b1 , \623_b1 );
xor ( \799_b0 , \798_b0 , w_1366 );
not ( w_1366 , w_1367 );
and ( w_1367 , \623_b1 , \623_b0 );
or ( \800_b1 , \797_b1 , \799_b1 );
not ( \799_b1 , w_1368 );
and ( \800_b0 , \797_b0 , w_1369 );
and ( w_1368 , w_1369 , \799_b0 );
or ( \801_b1 , \708_b1 , \717_b1 );
xor ( \801_b0 , \708_b0 , w_1370 );
not ( w_1370 , w_1371 );
and ( w_1371 , \717_b1 , \717_b0 );
or ( \802_b1 , \801_b1 , \720_b1 );
xor ( \802_b0 , \801_b0 , w_1372 );
not ( w_1372 , w_1373 );
and ( w_1373 , \720_b1 , \720_b0 );
or ( \803_b1 , \799_b1 , \802_b1 );
not ( \802_b1 , w_1374 );
and ( \803_b0 , \799_b0 , w_1375 );
and ( w_1374 , w_1375 , \802_b0 );
or ( \804_b1 , \797_b1 , \802_b1 );
not ( \802_b1 , w_1376 );
and ( \804_b0 , \797_b0 , w_1377 );
and ( w_1376 , w_1377 , \802_b0 );
or ( \806_b1 , \723_b1 , \725_b1 );
xor ( \806_b0 , \723_b0 , w_1378 );
not ( w_1378 , w_1379 );
and ( w_1379 , \725_b1 , \725_b0 );
or ( \807_b1 , \806_b1 , \727_b1 );
xor ( \807_b0 , \806_b0 , w_1380 );
not ( w_1380 , w_1381 );
and ( w_1381 , \727_b1 , \727_b0 );
or ( \808_b1 , \805_b1 , \807_b1 );
not ( \807_b1 , w_1382 );
and ( \808_b0 , \805_b0 , w_1383 );
and ( w_1382 , w_1383 , \807_b0 );
or ( \809_b1 , \736_b1 , \808_b1 );
not ( \808_b1 , w_1384 );
and ( \809_b0 , \736_b0 , w_1385 );
and ( w_1384 , w_1385 , \808_b0 );
or ( \810_b1 , \736_b1 , \808_b1 );
xor ( \810_b0 , \736_b0 , w_1386 );
not ( w_1386 , w_1387 );
and ( w_1387 , \808_b1 , \808_b0 );
or ( \811_b1 , \805_b1 , \807_b1 );
xor ( \811_b0 , \805_b0 , w_1388 );
not ( w_1388 , w_1389 );
and ( w_1389 , \807_b1 , \807_b0 );
and ( \812_nR134_b1 , RIb4c3200_48_b1 , w_1390 );
xor ( w_1390 , RIb4c3200_48_b0 , \288_b1 );
not ( \288_b1 , w_1391 );
and ( \812_nR134_b0 , w_1391 , \288_b0 );
buf ( \813_b1 , \812_nR134_b1 );
buf ( \813_b0 , \812_nR134_b0 );
and ( \814_nR133_b1 , RIb4c3188_49_b1 , w_1392 );
xor ( w_1392 , RIb4c3188_49_b0 , \288_b1 );
not ( \288_b1 , w_1393 );
and ( \814_nR133_b0 , w_1393 , \288_b0 );
buf ( \815_b1 , \814_nR133_b1 );
buf ( \815_b0 , \814_nR133_b0 );
or ( \816_b1 , \813_b1 , \815_b1 );
not ( \815_b1 , w_1394 );
and ( \816_b0 , \813_b0 , w_1395 );
and ( w_1394 , w_1395 , \815_b0 );
buf ( \817_b1 , \816_b1 );
not ( \817_b1 , w_1396 );
not ( \817_b0 , w_1397 );
and ( w_1396 , w_1397 , \816_b0 );
or ( \818_b1 , \665_b1 , \817_b1 );
not ( \817_b1 , w_1398 );
and ( \818_b0 , \665_b0 , w_1399 );
and ( w_1398 , w_1399 , \817_b0 );
buf ( \819_b1 , \818_b1 );
not ( \819_b1 , w_1400 );
not ( \819_b0 , w_1401 );
and ( w_1400 , w_1401 , \818_b0 );
or ( \820_b1 , \315_b1 , \740_b1 );
not ( \740_b1 , w_1402 );
and ( \820_b0 , \315_b0 , w_1403 );
and ( w_1402 , w_1403 , \740_b0 );
or ( \821_b1 , \159_b1 , \738_b1 );
not ( \738_b1 , w_1404 );
and ( \821_b0 , \159_b0 , w_1405 );
and ( w_1404 , w_1405 , \738_b0 );
or ( \822_b1 , \820_b1 , w_1407 );
not ( w_1407 , w_1408 );
and ( \822_b0 , \820_b0 , w_1409 );
and ( w_1408 ,  , w_1409 );
buf ( w_1407 , \821_b1 );
not ( w_1407 , w_1410 );
not (  , w_1411 );
and ( w_1410 , w_1411 , \821_b0 );
or ( \823_b1 , \822_b1 , w_1412 );
xor ( \823_b0 , \822_b0 , w_1414 );
not ( w_1414 , w_1415 );
and ( w_1415 , w_1412 , w_1413 );
buf ( w_1412 , \668_b1 );
not ( w_1412 , w_1416 );
not ( w_1413 , w_1417 );
and ( w_1416 , w_1417 , \668_b0 );
or ( \824_b1 , \819_b1 , \823_b1 );
not ( \823_b1 , w_1418 );
and ( \824_b0 , \819_b0 , w_1419 );
and ( w_1418 , w_1419 , \823_b0 );
or ( \825_b1 , \333_b1 , \604_b1 );
not ( \604_b1 , w_1420 );
and ( \825_b0 , \333_b0 , w_1421 );
and ( w_1420 , w_1421 , \604_b0 );
or ( \826_b1 , \305_b1 , \602_b1 );
not ( \602_b1 , w_1422 );
and ( \826_b0 , \305_b0 , w_1423 );
and ( w_1422 , w_1423 , \602_b0 );
or ( \827_b1 , \825_b1 , w_1425 );
not ( w_1425 , w_1426 );
and ( \827_b0 , \825_b0 , w_1427 );
and ( w_1426 ,  , w_1427 );
buf ( w_1425 , \826_b1 );
not ( w_1425 , w_1428 );
not (  , w_1429 );
and ( w_1428 , w_1429 , \826_b0 );
or ( \828_b1 , \827_b1 , w_1430 );
xor ( \828_b0 , \827_b0 , w_1432 );
not ( w_1432 , w_1433 );
and ( w_1433 , w_1430 , w_1431 );
buf ( w_1430 , \561_b1 );
not ( w_1430 , w_1434 );
not ( w_1431 , w_1435 );
and ( w_1434 , w_1435 , \561_b0 );
or ( \829_b1 , \823_b1 , \828_b1 );
not ( \828_b1 , w_1436 );
and ( \829_b0 , \823_b0 , w_1437 );
and ( w_1436 , w_1437 , \828_b0 );
or ( \830_b1 , \819_b1 , \828_b1 );
not ( \828_b1 , w_1438 );
and ( \830_b0 , \819_b0 , w_1439 );
and ( w_1438 , w_1439 , \828_b0 );
or ( \832_b1 , \621_b1 , \331_b1 );
not ( \331_b1 , w_1440 );
and ( \832_b0 , \621_b0 , w_1441 );
and ( w_1440 , w_1441 , \331_b0 );
or ( \833_b1 , \593_b1 , \329_b1 );
not ( \329_b1 , w_1442 );
and ( \833_b0 , \593_b0 , w_1443 );
and ( w_1442 , w_1443 , \329_b0 );
or ( \834_b1 , \832_b1 , w_1445 );
not ( w_1445 , w_1446 );
and ( \834_b0 , \832_b0 , w_1447 );
and ( w_1446 ,  , w_1447 );
buf ( w_1445 , \833_b1 );
not ( w_1445 , w_1448 );
not (  , w_1449 );
and ( w_1448 , w_1449 , \833_b0 );
or ( \835_b1 , \834_b1 , w_1450 );
xor ( \835_b0 , \834_b0 , w_1452 );
not ( w_1452 , w_1453 );
and ( w_1453 , w_1450 , w_1451 );
buf ( w_1450 , \338_b1 );
not ( w_1450 , w_1454 );
not ( w_1451 , w_1455 );
and ( w_1454 , w_1455 , \338_b0 );
or ( \836_b1 , \777_b1 , \351_b1 );
not ( \351_b1 , w_1456 );
and ( \836_b0 , \777_b0 , w_1457 );
and ( w_1456 , w_1457 , \351_b0 );
or ( \837_b1 , \703_b1 , \349_b1 );
not ( \349_b1 , w_1458 );
and ( \837_b0 , \703_b0 , w_1459 );
and ( w_1458 , w_1459 , \349_b0 );
or ( \838_b1 , \836_b1 , w_1461 );
not ( w_1461 , w_1462 );
and ( \838_b0 , \836_b0 , w_1463 );
and ( w_1462 ,  , w_1463 );
buf ( w_1461 , \837_b1 );
not ( w_1461 , w_1464 );
not (  , w_1465 );
and ( w_1464 , w_1465 , \837_b0 );
or ( \839_b1 , \838_b1 , w_1466 );
xor ( \839_b0 , \838_b0 , w_1468 );
not ( w_1468 , w_1469 );
and ( w_1469 , w_1466 , w_1467 );
buf ( w_1466 , \358_b1 );
not ( w_1466 , w_1470 );
not ( w_1467 , w_1471 );
and ( w_1470 , w_1471 , \358_b0 );
or ( \840_b1 , \835_b1 , \839_b1 );
not ( \839_b1 , w_1472 );
and ( \840_b0 , \835_b0 , w_1473 );
and ( w_1472 , w_1473 , \839_b0 );
buf ( \841_b1 , RIb4bf3a8_79_b1 );
buf ( \841_b0 , RIb4bf3a8_79_b0 );
or ( \842_b1 , \841_b1 , \345_b1 );
not ( \345_b1 , w_1474 );
and ( \842_b0 , \841_b0 , w_1475 );
and ( w_1474 , w_1475 , \345_b0 );
or ( \843_b1 , \839_b1 , \842_b1 );
not ( \842_b1 , w_1476 );
and ( \843_b0 , \839_b0 , w_1477 );
and ( w_1476 , w_1477 , \842_b0 );
or ( \844_b1 , \835_b1 , \842_b1 );
not ( \842_b1 , w_1478 );
and ( \844_b0 , \835_b0 , w_1479 );
and ( w_1478 , w_1479 , \842_b0 );
or ( \846_b1 , \831_b1 , \845_b1 );
not ( \845_b1 , w_1480 );
and ( \846_b0 , \831_b0 , w_1481 );
and ( w_1480 , w_1481 , \845_b0 );
or ( \847_b1 , \353_b1 , \503_b1 );
not ( \503_b1 , w_1482 );
and ( \847_b0 , \353_b0 , w_1483 );
and ( w_1482 , w_1483 , \503_b0 );
or ( \848_b1 , \323_b1 , \501_b1 );
not ( \501_b1 , w_1484 );
and ( \848_b0 , \323_b0 , w_1485 );
and ( w_1484 , w_1485 , \501_b0 );
or ( \849_b1 , \847_b1 , w_1487 );
not ( w_1487 , w_1488 );
and ( \849_b0 , \847_b0 , w_1489 );
and ( w_1488 ,  , w_1489 );
buf ( w_1487 , \848_b1 );
not ( w_1487 , w_1490 );
not (  , w_1491 );
and ( w_1490 , w_1491 , \848_b0 );
or ( \850_b1 , \849_b1 , w_1492 );
xor ( \850_b0 , \849_b0 , w_1494 );
not ( w_1494 , w_1495 );
and ( w_1495 , w_1492 , w_1493 );
buf ( w_1492 , \455_b1 );
not ( w_1492 , w_1496 );
not ( w_1493 , w_1497 );
and ( w_1496 , w_1497 , \455_b0 );
or ( \851_b1 , \360_b1 , \298_b1 );
not ( \298_b1 , w_1498 );
and ( \851_b0 , \360_b0 , w_1499 );
and ( w_1498 , w_1499 , \298_b0 );
or ( \852_b1 , \343_b1 , \296_b1 );
not ( \296_b1 , w_1500 );
and ( \852_b0 , \343_b0 , w_1501 );
and ( w_1500 , w_1501 , \296_b0 );
or ( \853_b1 , \851_b1 , w_1503 );
not ( w_1503 , w_1504 );
and ( \853_b0 , \851_b0 , w_1505 );
and ( w_1504 ,  , w_1505 );
buf ( w_1503 , \852_b1 );
not ( w_1503 , w_1506 );
not (  , w_1507 );
and ( w_1506 , w_1507 , \852_b0 );
or ( \854_b1 , \853_b1 , w_1508 );
xor ( \854_b0 , \853_b0 , w_1510 );
not ( w_1510 , w_1511 );
and ( w_1511 , w_1508 , w_1509 );
buf ( w_1508 , \303_b1 );
not ( w_1508 , w_1512 );
not ( w_1509 , w_1513 );
and ( w_1512 , w_1513 , \303_b0 );
or ( \855_b1 , \850_b1 , \854_b1 );
not ( \854_b1 , w_1514 );
and ( \855_b0 , \850_b0 , w_1515 );
and ( w_1514 , w_1515 , \854_b0 );
or ( \856_b1 , \495_b1 , \313_b1 );
not ( \313_b1 , w_1516 );
and ( \856_b0 , \495_b0 , w_1517 );
and ( w_1516 , w_1517 , \313_b0 );
or ( \857_b1 , \444_b1 , \311_b1 );
not ( \311_b1 , w_1518 );
and ( \857_b0 , \444_b0 , w_1519 );
and ( w_1518 , w_1519 , \311_b0 );
or ( \858_b1 , \856_b1 , w_1521 );
not ( w_1521 , w_1522 );
and ( \858_b0 , \856_b0 , w_1523 );
and ( w_1522 ,  , w_1523 );
buf ( w_1521 , \857_b1 );
not ( w_1521 , w_1524 );
not (  , w_1525 );
and ( w_1524 , w_1525 , \857_b0 );
or ( \859_b1 , \858_b1 , w_1526 );
xor ( \859_b0 , \858_b0 , w_1528 );
not ( w_1528 , w_1529 );
and ( w_1529 , w_1526 , w_1527 );
buf ( w_1526 , \320_b1 );
not ( w_1526 , w_1530 );
not ( w_1527 , w_1531 );
and ( w_1530 , w_1531 , \320_b0 );
or ( \860_b1 , \854_b1 , \859_b1 );
not ( \859_b1 , w_1532 );
and ( \860_b0 , \854_b0 , w_1533 );
and ( w_1532 , w_1533 , \859_b0 );
or ( \861_b1 , \850_b1 , \859_b1 );
not ( \859_b1 , w_1534 );
and ( \861_b0 , \850_b0 , w_1535 );
and ( w_1534 , w_1535 , \859_b0 );
or ( \863_b1 , \845_b1 , \862_b1 );
not ( \862_b1 , w_1536 );
and ( \863_b0 , \845_b0 , w_1537 );
and ( w_1536 , w_1537 , \862_b0 );
or ( \864_b1 , \831_b1 , \862_b1 );
not ( \862_b1 , w_1538 );
and ( \864_b0 , \831_b0 , w_1539 );
and ( w_1538 , w_1539 , \862_b0 );
or ( \866_b1 , \743_b1 , \747_b1 );
xor ( \866_b0 , \743_b0 , w_1540 );
not ( w_1540 , w_1541 );
and ( w_1541 , \747_b1 , \747_b0 );
or ( \867_b1 , \866_b1 , \752_b1 );
xor ( \867_b0 , \866_b0 , w_1542 );
not ( w_1542 , w_1543 );
and ( w_1543 , \752_b1 , \752_b0 );
or ( \868_b1 , \759_b1 , \763_b1 );
xor ( \868_b0 , \759_b0 , w_1544 );
not ( w_1544 , w_1545 );
and ( w_1545 , \763_b1 , \763_b0 );
or ( \869_b1 , \868_b1 , \768_b1 );
xor ( \869_b0 , \868_b0 , w_1546 );
not ( w_1546 , w_1547 );
and ( w_1547 , \768_b1 , \768_b0 );
or ( \870_b1 , \867_b1 , \869_b1 );
not ( \869_b1 , w_1548 );
and ( \870_b0 , \867_b0 , w_1549 );
and ( w_1548 , w_1549 , \869_b0 );
or ( \871_b1 , \776_b1 , w_1550 );
xor ( \871_b0 , \776_b0 , w_1552 );
not ( w_1552 , w_1553 );
and ( w_1553 , w_1550 , w_1551 );
buf ( w_1550 , \778_b1 );
not ( w_1550 , w_1554 );
not ( w_1551 , w_1555 );
and ( w_1554 , w_1555 , \778_b0 );
or ( \872_b1 , \869_b1 , \871_b1 );
not ( \871_b1 , w_1556 );
and ( \872_b0 , \869_b0 , w_1557 );
and ( w_1556 , w_1557 , \871_b0 );
or ( \873_b1 , \867_b1 , \871_b1 );
not ( \871_b1 , w_1558 );
and ( \873_b0 , \867_b0 , w_1559 );
and ( w_1558 , w_1559 , \871_b0 );
or ( \875_b1 , \865_b1 , \874_b1 );
not ( \874_b1 , w_1560 );
and ( \875_b0 , \865_b0 , w_1561 );
and ( w_1560 , w_1561 , \874_b0 );
or ( \876_b1 , \784_b1 , \786_b1 );
xor ( \876_b0 , \784_b0 , w_1562 );
not ( w_1562 , w_1563 );
and ( w_1563 , \786_b1 , \786_b0 );
or ( \877_b1 , \876_b1 , \788_b1 );
xor ( \877_b0 , \876_b0 , w_1564 );
not ( w_1564 , w_1565 );
and ( w_1565 , \788_b1 , \788_b0 );
or ( \878_b1 , \874_b1 , \877_b1 );
not ( \877_b1 , w_1566 );
and ( \878_b0 , \874_b0 , w_1567 );
and ( w_1566 , w_1567 , \877_b0 );
or ( \879_b1 , \865_b1 , \877_b1 );
not ( \877_b1 , w_1568 );
and ( \879_b0 , \865_b0 , w_1569 );
and ( w_1568 , w_1569 , \877_b0 );
or ( \881_b1 , \681_b1 , \697_b1 );
xor ( \881_b0 , \681_b0 , w_1570 );
not ( w_1570 , w_1571 );
and ( w_1571 , \697_b1 , \697_b0 );
or ( \882_b1 , \881_b1 , \705_b1 );
xor ( \882_b0 , \881_b0 , w_1572 );
not ( w_1572 , w_1573 );
and ( w_1573 , \705_b1 , \705_b0 );
or ( \883_b1 , \880_b1 , \882_b1 );
not ( \882_b1 , w_1574 );
and ( \883_b0 , \880_b0 , w_1575 );
and ( w_1574 , w_1575 , \882_b0 );
or ( \884_b1 , \782_b1 , \791_b1 );
xor ( \884_b0 , \782_b0 , w_1576 );
not ( w_1576 , w_1577 );
and ( w_1577 , \791_b1 , \791_b0 );
or ( \885_b1 , \884_b1 , \794_b1 );
xor ( \885_b0 , \884_b0 , w_1578 );
not ( w_1578 , w_1579 );
and ( w_1579 , \794_b1 , \794_b0 );
or ( \886_b1 , \882_b1 , \885_b1 );
not ( \885_b1 , w_1580 );
and ( \886_b0 , \882_b0 , w_1581 );
and ( w_1580 , w_1581 , \885_b0 );
or ( \887_b1 , \880_b1 , \885_b1 );
not ( \885_b1 , w_1582 );
and ( \887_b0 , \880_b0 , w_1583 );
and ( w_1582 , w_1583 , \885_b0 );
or ( \889_b1 , \797_b1 , \799_b1 );
xor ( \889_b0 , \797_b0 , w_1584 );
not ( w_1584 , w_1585 );
and ( w_1585 , \799_b1 , \799_b0 );
or ( \890_b1 , \889_b1 , \802_b1 );
xor ( \890_b0 , \889_b0 , w_1586 );
not ( w_1586 , w_1587 );
and ( w_1587 , \802_b1 , \802_b0 );
or ( \891_b1 , \888_b1 , \890_b1 );
not ( \890_b1 , w_1588 );
and ( \891_b0 , \888_b0 , w_1589 );
and ( w_1588 , w_1589 , \890_b0 );
or ( \892_b1 , \811_b1 , \891_b1 );
not ( \891_b1 , w_1590 );
and ( \892_b0 , \811_b0 , w_1591 );
and ( w_1590 , w_1591 , \891_b0 );
or ( \893_b1 , \811_b1 , \891_b1 );
xor ( \893_b0 , \811_b0 , w_1592 );
not ( w_1592 , w_1593 );
and ( w_1593 , \891_b1 , \891_b0 );
or ( \894_b1 , \888_b1 , \890_b1 );
xor ( \894_b0 , \888_b0 , w_1594 );
not ( w_1594 , w_1595 );
and ( w_1595 , \890_b1 , \890_b0 );
or ( \895_b1 , \703_b1 , \331_b1 );
not ( \331_b1 , w_1596 );
and ( \895_b0 , \703_b0 , w_1597 );
and ( w_1596 , w_1597 , \331_b0 );
or ( \896_b1 , \621_b1 , \329_b1 );
not ( \329_b1 , w_1598 );
and ( \896_b0 , \621_b0 , w_1599 );
and ( w_1598 , w_1599 , \329_b0 );
or ( \897_b1 , \895_b1 , w_1601 );
not ( w_1601 , w_1602 );
and ( \897_b0 , \895_b0 , w_1603 );
and ( w_1602 ,  , w_1603 );
buf ( w_1601 , \896_b1 );
not ( w_1601 , w_1604 );
not (  , w_1605 );
and ( w_1604 , w_1605 , \896_b0 );
or ( \898_b1 , \897_b1 , w_1606 );
xor ( \898_b0 , \897_b0 , w_1608 );
not ( w_1608 , w_1609 );
and ( w_1609 , w_1606 , w_1607 );
buf ( w_1606 , \338_b1 );
not ( w_1606 , w_1610 );
not ( w_1607 , w_1611 );
and ( w_1610 , w_1611 , \338_b0 );
or ( \899_b1 , \841_b1 , \351_b1 );
not ( \351_b1 , w_1612 );
and ( \899_b0 , \841_b0 , w_1613 );
and ( w_1612 , w_1613 , \351_b0 );
or ( \900_b1 , \777_b1 , \349_b1 );
not ( \349_b1 , w_1614 );
and ( \900_b0 , \777_b0 , w_1615 );
and ( w_1614 , w_1615 , \349_b0 );
or ( \901_b1 , \899_b1 , w_1617 );
not ( w_1617 , w_1618 );
and ( \901_b0 , \899_b0 , w_1619 );
and ( w_1618 ,  , w_1619 );
buf ( w_1617 , \900_b1 );
not ( w_1617 , w_1620 );
not (  , w_1621 );
and ( w_1620 , w_1621 , \900_b0 );
or ( \902_b1 , \901_b1 , w_1622 );
xor ( \902_b0 , \901_b0 , w_1624 );
not ( w_1624 , w_1625 );
and ( w_1625 , w_1622 , w_1623 );
buf ( w_1622 , \358_b1 );
not ( w_1622 , w_1626 );
not ( w_1623 , w_1627 );
and ( w_1626 , w_1627 , \358_b0 );
or ( \903_b1 , \898_b1 , \902_b1 );
not ( \902_b1 , w_1628 );
and ( \903_b0 , \898_b0 , w_1629 );
and ( w_1628 , w_1629 , \902_b0 );
buf ( \904_b1 , RIb4bf330_80_b1 );
buf ( \904_b0 , RIb4bf330_80_b0 );
or ( \905_b1 , \904_b1 , \345_b1 );
not ( \345_b1 , w_1630 );
and ( \905_b0 , \904_b0 , w_1631 );
and ( w_1630 , w_1631 , \345_b0 );
or ( \906_b1 , \902_b1 , \905_b1 );
not ( \905_b1 , w_1632 );
and ( \906_b0 , \902_b0 , w_1633 );
and ( w_1632 , w_1633 , \905_b0 );
or ( \907_b1 , \898_b1 , \905_b1 );
not ( \905_b1 , w_1634 );
and ( \907_b0 , \898_b0 , w_1635 );
and ( w_1634 , w_1635 , \905_b0 );
or ( \909_b1 , \665_b1 , \813_b1 );
xor ( \909_b0 , \665_b0 , w_1636 );
not ( w_1636 , w_1637 );
and ( w_1637 , \813_b1 , \813_b0 );
or ( \910_b1 , \813_b1 , \815_b1 );
xor ( \910_b0 , \813_b0 , w_1638 );
not ( w_1638 , w_1639 );
and ( w_1639 , \815_b1 , \815_b0 );
buf ( \911_b1 , \910_b1 );
not ( \911_b1 , w_1640 );
not ( \911_b0 , w_1641 );
and ( w_1640 , w_1641 , \910_b0 );
or ( \912_b1 , \909_b1 , \911_b1 );
not ( \911_b1 , w_1642 );
and ( \912_b0 , \909_b0 , w_1643 );
and ( w_1642 , w_1643 , \911_b0 );
or ( \913_b1 , \159_b1 , \912_b1 );
not ( \912_b1 , w_1644 );
and ( \913_b0 , \159_b0 , w_1645 );
and ( w_1644 , w_1645 , \912_b0 );
buf ( \914_b1 , \913_b1 );
not ( \914_b1 , w_1646 );
not ( \914_b0 , w_1647 );
and ( w_1646 , w_1647 , \913_b0 );
or ( \915_b1 , \914_b1 , w_1648 );
xor ( \915_b0 , \914_b0 , w_1650 );
not ( w_1650 , w_1651 );
and ( w_1651 , w_1648 , w_1649 );
buf ( w_1648 , \818_b1 );
not ( w_1648 , w_1652 );
not ( w_1649 , w_1653 );
and ( w_1652 , w_1653 , \818_b0 );
or ( \916_b1 , \305_b1 , \740_b1 );
not ( \740_b1 , w_1654 );
and ( \916_b0 , \305_b0 , w_1655 );
and ( w_1654 , w_1655 , \740_b0 );
or ( \917_b1 , \315_b1 , \738_b1 );
not ( \738_b1 , w_1656 );
and ( \917_b0 , \315_b0 , w_1657 );
and ( w_1656 , w_1657 , \738_b0 );
or ( \918_b1 , \916_b1 , w_1659 );
not ( w_1659 , w_1660 );
and ( \918_b0 , \916_b0 , w_1661 );
and ( w_1660 ,  , w_1661 );
buf ( w_1659 , \917_b1 );
not ( w_1659 , w_1662 );
not (  , w_1663 );
and ( w_1662 , w_1663 , \917_b0 );
or ( \919_b1 , \918_b1 , w_1664 );
xor ( \919_b0 , \918_b0 , w_1666 );
not ( w_1666 , w_1667 );
and ( w_1667 , w_1664 , w_1665 );
buf ( w_1664 , \668_b1 );
not ( w_1664 , w_1668 );
not ( w_1665 , w_1669 );
and ( w_1668 , w_1669 , \668_b0 );
or ( \920_b1 , \915_b1 , \919_b1 );
not ( \919_b1 , w_1670 );
and ( \920_b0 , \915_b0 , w_1671 );
and ( w_1670 , w_1671 , \919_b0 );
or ( \921_b1 , \323_b1 , \604_b1 );
not ( \604_b1 , w_1672 );
and ( \921_b0 , \323_b0 , w_1673 );
and ( w_1672 , w_1673 , \604_b0 );
or ( \922_b1 , \333_b1 , \602_b1 );
not ( \602_b1 , w_1674 );
and ( \922_b0 , \333_b0 , w_1675 );
and ( w_1674 , w_1675 , \602_b0 );
or ( \923_b1 , \921_b1 , w_1677 );
not ( w_1677 , w_1678 );
and ( \923_b0 , \921_b0 , w_1679 );
and ( w_1678 ,  , w_1679 );
buf ( w_1677 , \922_b1 );
not ( w_1677 , w_1680 );
not (  , w_1681 );
and ( w_1680 , w_1681 , \922_b0 );
or ( \924_b1 , \923_b1 , w_1682 );
xor ( \924_b0 , \923_b0 , w_1684 );
not ( w_1684 , w_1685 );
and ( w_1685 , w_1682 , w_1683 );
buf ( w_1682 , \561_b1 );
not ( w_1682 , w_1686 );
not ( w_1683 , w_1687 );
and ( w_1686 , w_1687 , \561_b0 );
or ( \925_b1 , \919_b1 , \924_b1 );
not ( \924_b1 , w_1688 );
and ( \925_b0 , \919_b0 , w_1689 );
and ( w_1688 , w_1689 , \924_b0 );
or ( \926_b1 , \915_b1 , \924_b1 );
not ( \924_b1 , w_1690 );
and ( \926_b0 , \915_b0 , w_1691 );
and ( w_1690 , w_1691 , \924_b0 );
or ( \928_b1 , \908_b1 , \927_b1 );
not ( \927_b1 , w_1692 );
and ( \928_b0 , \908_b0 , w_1693 );
and ( w_1692 , w_1693 , \927_b0 );
or ( \929_b1 , \343_b1 , \503_b1 );
not ( \503_b1 , w_1694 );
and ( \929_b0 , \343_b0 , w_1695 );
and ( w_1694 , w_1695 , \503_b0 );
or ( \930_b1 , \353_b1 , \501_b1 );
not ( \501_b1 , w_1696 );
and ( \930_b0 , \353_b0 , w_1697 );
and ( w_1696 , w_1697 , \501_b0 );
or ( \931_b1 , \929_b1 , w_1699 );
not ( w_1699 , w_1700 );
and ( \931_b0 , \929_b0 , w_1701 );
and ( w_1700 ,  , w_1701 );
buf ( w_1699 , \930_b1 );
not ( w_1699 , w_1702 );
not (  , w_1703 );
and ( w_1702 , w_1703 , \930_b0 );
or ( \932_b1 , \931_b1 , w_1704 );
xor ( \932_b0 , \931_b0 , w_1706 );
not ( w_1706 , w_1707 );
and ( w_1707 , w_1704 , w_1705 );
buf ( w_1704 , \455_b1 );
not ( w_1704 , w_1708 );
not ( w_1705 , w_1709 );
and ( w_1708 , w_1709 , \455_b0 );
or ( \933_b1 , \444_b1 , \298_b1 );
not ( \298_b1 , w_1710 );
and ( \933_b0 , \444_b0 , w_1711 );
and ( w_1710 , w_1711 , \298_b0 );
or ( \934_b1 , \360_b1 , \296_b1 );
not ( \296_b1 , w_1712 );
and ( \934_b0 , \360_b0 , w_1713 );
and ( w_1712 , w_1713 , \296_b0 );
or ( \935_b1 , \933_b1 , w_1715 );
not ( w_1715 , w_1716 );
and ( \935_b0 , \933_b0 , w_1717 );
and ( w_1716 ,  , w_1717 );
buf ( w_1715 , \934_b1 );
not ( w_1715 , w_1718 );
not (  , w_1719 );
and ( w_1718 , w_1719 , \934_b0 );
or ( \936_b1 , \935_b1 , w_1720 );
xor ( \936_b0 , \935_b0 , w_1722 );
not ( w_1722 , w_1723 );
and ( w_1723 , w_1720 , w_1721 );
buf ( w_1720 , \303_b1 );
not ( w_1720 , w_1724 );
not ( w_1721 , w_1725 );
and ( w_1724 , w_1725 , \303_b0 );
or ( \937_b1 , \932_b1 , \936_b1 );
not ( \936_b1 , w_1726 );
and ( \937_b0 , \932_b0 , w_1727 );
and ( w_1726 , w_1727 , \936_b0 );
or ( \938_b1 , \593_b1 , \313_b1 );
not ( \313_b1 , w_1728 );
and ( \938_b0 , \593_b0 , w_1729 );
and ( w_1728 , w_1729 , \313_b0 );
or ( \939_b1 , \495_b1 , \311_b1 );
not ( \311_b1 , w_1730 );
and ( \939_b0 , \495_b0 , w_1731 );
and ( w_1730 , w_1731 , \311_b0 );
or ( \940_b1 , \938_b1 , w_1733 );
not ( w_1733 , w_1734 );
and ( \940_b0 , \938_b0 , w_1735 );
and ( w_1734 ,  , w_1735 );
buf ( w_1733 , \939_b1 );
not ( w_1733 , w_1736 );
not (  , w_1737 );
and ( w_1736 , w_1737 , \939_b0 );
or ( \941_b1 , \940_b1 , w_1738 );
xor ( \941_b0 , \940_b0 , w_1740 );
not ( w_1740 , w_1741 );
and ( w_1741 , w_1738 , w_1739 );
buf ( w_1738 , \320_b1 );
not ( w_1738 , w_1742 );
not ( w_1739 , w_1743 );
and ( w_1742 , w_1743 , \320_b0 );
or ( \942_b1 , \936_b1 , \941_b1 );
not ( \941_b1 , w_1744 );
and ( \942_b0 , \936_b0 , w_1745 );
and ( w_1744 , w_1745 , \941_b0 );
or ( \943_b1 , \932_b1 , \941_b1 );
not ( \941_b1 , w_1746 );
and ( \943_b0 , \932_b0 , w_1747 );
and ( w_1746 , w_1747 , \941_b0 );
or ( \945_b1 , \927_b1 , \944_b1 );
not ( \944_b1 , w_1748 );
and ( \945_b0 , \927_b0 , w_1749 );
and ( w_1748 , w_1749 , \944_b0 );
or ( \946_b1 , \908_b1 , \944_b1 );
not ( \944_b1 , w_1750 );
and ( \946_b0 , \908_b0 , w_1751 );
and ( w_1750 , w_1751 , \944_b0 );
or ( \948_b1 , \819_b1 , \823_b1 );
xor ( \948_b0 , \819_b0 , w_1752 );
not ( w_1752 , w_1753 );
and ( w_1753 , \823_b1 , \823_b0 );
or ( \949_b1 , \948_b1 , \828_b1 );
xor ( \949_b0 , \948_b0 , w_1754 );
not ( w_1754 , w_1755 );
and ( w_1755 , \828_b1 , \828_b0 );
or ( \950_b1 , \835_b1 , \839_b1 );
xor ( \950_b0 , \835_b0 , w_1756 );
not ( w_1756 , w_1757 );
and ( w_1757 , \839_b1 , \839_b0 );
or ( \951_b1 , \950_b1 , \842_b1 );
xor ( \951_b0 , \950_b0 , w_1758 );
not ( w_1758 , w_1759 );
and ( w_1759 , \842_b1 , \842_b0 );
or ( \952_b1 , \949_b1 , \951_b1 );
not ( \951_b1 , w_1760 );
and ( \952_b0 , \949_b0 , w_1761 );
and ( w_1760 , w_1761 , \951_b0 );
or ( \953_b1 , \850_b1 , \854_b1 );
xor ( \953_b0 , \850_b0 , w_1762 );
not ( w_1762 , w_1763 );
and ( w_1763 , \854_b1 , \854_b0 );
or ( \954_b1 , \953_b1 , \859_b1 );
xor ( \954_b0 , \953_b0 , w_1764 );
not ( w_1764 , w_1765 );
and ( w_1765 , \859_b1 , \859_b0 );
or ( \955_b1 , \951_b1 , \954_b1 );
not ( \954_b1 , w_1766 );
and ( \955_b0 , \951_b0 , w_1767 );
and ( w_1766 , w_1767 , \954_b0 );
or ( \956_b1 , \949_b1 , \954_b1 );
not ( \954_b1 , w_1768 );
and ( \956_b0 , \949_b0 , w_1769 );
and ( w_1768 , w_1769 , \954_b0 );
or ( \958_b1 , \947_b1 , \957_b1 );
not ( \957_b1 , w_1770 );
and ( \958_b0 , \947_b0 , w_1771 );
and ( w_1770 , w_1771 , \957_b0 );
or ( \959_b1 , \867_b1 , \869_b1 );
xor ( \959_b0 , \867_b0 , w_1772 );
not ( w_1772 , w_1773 );
and ( w_1773 , \869_b1 , \869_b0 );
or ( \960_b1 , \959_b1 , \871_b1 );
xor ( \960_b0 , \959_b0 , w_1774 );
not ( w_1774 , w_1775 );
and ( w_1775 , \871_b1 , \871_b0 );
or ( \961_b1 , \957_b1 , \960_b1 );
not ( \960_b1 , w_1776 );
and ( \961_b0 , \957_b0 , w_1777 );
and ( w_1776 , w_1777 , \960_b0 );
or ( \962_b1 , \947_b1 , \960_b1 );
not ( \960_b1 , w_1778 );
and ( \962_b0 , \947_b0 , w_1779 );
and ( w_1778 , w_1779 , \960_b0 );
or ( \964_b1 , \755_b1 , \771_b1 );
xor ( \964_b0 , \755_b0 , w_1780 );
not ( w_1780 , w_1781 );
and ( w_1781 , \771_b1 , \771_b0 );
or ( \965_b1 , \964_b1 , \779_b1 );
xor ( \965_b0 , \964_b0 , w_1782 );
not ( w_1782 , w_1783 );
and ( w_1783 , \779_b1 , \779_b0 );
or ( \966_b1 , \963_b1 , \965_b1 );
not ( \965_b1 , w_1784 );
and ( \966_b0 , \963_b0 , w_1785 );
and ( w_1784 , w_1785 , \965_b0 );
or ( \967_b1 , \865_b1 , \874_b1 );
xor ( \967_b0 , \865_b0 , w_1786 );
not ( w_1786 , w_1787 );
and ( w_1787 , \874_b1 , \874_b0 );
or ( \968_b1 , \967_b1 , \877_b1 );
xor ( \968_b0 , \967_b0 , w_1788 );
not ( w_1788 , w_1789 );
and ( w_1789 , \877_b1 , \877_b0 );
or ( \969_b1 , \965_b1 , \968_b1 );
not ( \968_b1 , w_1790 );
and ( \969_b0 , \965_b0 , w_1791 );
and ( w_1790 , w_1791 , \968_b0 );
or ( \970_b1 , \963_b1 , \968_b1 );
not ( \968_b1 , w_1792 );
and ( \970_b0 , \963_b0 , w_1793 );
and ( w_1792 , w_1793 , \968_b0 );
or ( \972_b1 , \880_b1 , \882_b1 );
xor ( \972_b0 , \880_b0 , w_1794 );
not ( w_1794 , w_1795 );
and ( w_1795 , \882_b1 , \882_b0 );
or ( \973_b1 , \972_b1 , \885_b1 );
xor ( \973_b0 , \972_b0 , w_1796 );
not ( w_1796 , w_1797 );
and ( w_1797 , \885_b1 , \885_b0 );
or ( \974_b1 , \971_b1 , \973_b1 );
not ( \973_b1 , w_1798 );
and ( \974_b0 , \971_b0 , w_1799 );
and ( w_1798 , w_1799 , \973_b0 );
or ( \975_b1 , \894_b1 , \974_b1 );
not ( \974_b1 , w_1800 );
and ( \975_b0 , \894_b0 , w_1801 );
and ( w_1800 , w_1801 , \974_b0 );
or ( \976_b1 , \894_b1 , \974_b1 );
xor ( \976_b0 , \894_b0 , w_1802 );
not ( w_1802 , w_1803 );
and ( w_1803 , \974_b1 , \974_b0 );
or ( \977_b1 , \971_b1 , \973_b1 );
xor ( \977_b0 , \971_b0 , w_1804 );
not ( w_1804 , w_1805 );
and ( w_1805 , \973_b1 , \973_b0 );
and ( \978_nR132_b1 , RIb4c3110_50_b1 , w_1806 );
xor ( w_1806 , RIb4c3110_50_b0 , \288_b1 );
not ( \288_b1 , w_1807 );
and ( \978_nR132_b0 , w_1807 , \288_b0 );
buf ( \979_b1 , \978_nR132_b1 );
buf ( \979_b0 , \978_nR132_b0 );
and ( \980_nR131_b1 , RIb4c3098_51_b1 , w_1808 );
xor ( w_1808 , RIb4c3098_51_b0 , \288_b1 );
not ( \288_b1 , w_1809 );
and ( \980_nR131_b0 , w_1809 , \288_b0 );
buf ( \981_b1 , \980_nR131_b1 );
buf ( \981_b0 , \980_nR131_b0 );
or ( \982_b1 , \979_b1 , \981_b1 );
not ( \981_b1 , w_1810 );
and ( \982_b0 , \979_b0 , w_1811 );
and ( w_1810 , w_1811 , \981_b0 );
buf ( \983_b1 , \982_b1 );
not ( \983_b1 , w_1812 );
not ( \983_b0 , w_1813 );
and ( w_1812 , w_1813 , \982_b0 );
or ( \984_b1 , \815_b1 , \983_b1 );
not ( \983_b1 , w_1814 );
and ( \984_b0 , \815_b0 , w_1815 );
and ( w_1814 , w_1815 , \983_b0 );
buf ( \985_b1 , \984_b1 );
not ( \985_b1 , w_1816 );
not ( \985_b0 , w_1817 );
and ( w_1816 , w_1817 , \984_b0 );
or ( \986_b1 , \315_b1 , \912_b1 );
not ( \912_b1 , w_1818 );
and ( \986_b0 , \315_b0 , w_1819 );
and ( w_1818 , w_1819 , \912_b0 );
or ( \987_b1 , \159_b1 , \910_b1 );
not ( \910_b1 , w_1820 );
and ( \987_b0 , \159_b0 , w_1821 );
and ( w_1820 , w_1821 , \910_b0 );
or ( \988_b1 , \986_b1 , w_1823 );
not ( w_1823 , w_1824 );
and ( \988_b0 , \986_b0 , w_1825 );
and ( w_1824 ,  , w_1825 );
buf ( w_1823 , \987_b1 );
not ( w_1823 , w_1826 );
not (  , w_1827 );
and ( w_1826 , w_1827 , \987_b0 );
or ( \989_b1 , \988_b1 , w_1828 );
xor ( \989_b0 , \988_b0 , w_1830 );
not ( w_1830 , w_1831 );
and ( w_1831 , w_1828 , w_1829 );
buf ( w_1828 , \818_b1 );
not ( w_1828 , w_1832 );
not ( w_1829 , w_1833 );
and ( w_1832 , w_1833 , \818_b0 );
or ( \990_b1 , \985_b1 , \989_b1 );
not ( \989_b1 , w_1834 );
and ( \990_b0 , \985_b0 , w_1835 );
and ( w_1834 , w_1835 , \989_b0 );
or ( \991_b1 , \333_b1 , \740_b1 );
not ( \740_b1 , w_1836 );
and ( \991_b0 , \333_b0 , w_1837 );
and ( w_1836 , w_1837 , \740_b0 );
or ( \992_b1 , \305_b1 , \738_b1 );
not ( \738_b1 , w_1838 );
and ( \992_b0 , \305_b0 , w_1839 );
and ( w_1838 , w_1839 , \738_b0 );
or ( \993_b1 , \991_b1 , w_1841 );
not ( w_1841 , w_1842 );
and ( \993_b0 , \991_b0 , w_1843 );
and ( w_1842 ,  , w_1843 );
buf ( w_1841 , \992_b1 );
not ( w_1841 , w_1844 );
not (  , w_1845 );
and ( w_1844 , w_1845 , \992_b0 );
or ( \994_b1 , \993_b1 , w_1846 );
xor ( \994_b0 , \993_b0 , w_1848 );
not ( w_1848 , w_1849 );
and ( w_1849 , w_1846 , w_1847 );
buf ( w_1846 , \668_b1 );
not ( w_1846 , w_1850 );
not ( w_1847 , w_1851 );
and ( w_1850 , w_1851 , \668_b0 );
or ( \995_b1 , \989_b1 , \994_b1 );
not ( \994_b1 , w_1852 );
and ( \995_b0 , \989_b0 , w_1853 );
and ( w_1852 , w_1853 , \994_b0 );
or ( \996_b1 , \985_b1 , \994_b1 );
not ( \994_b1 , w_1854 );
and ( \996_b0 , \985_b0 , w_1855 );
and ( w_1854 , w_1855 , \994_b0 );
or ( \998_b1 , \353_b1 , \604_b1 );
not ( \604_b1 , w_1856 );
and ( \998_b0 , \353_b0 , w_1857 );
and ( w_1856 , w_1857 , \604_b0 );
or ( \999_b1 , \323_b1 , \602_b1 );
not ( \602_b1 , w_1858 );
and ( \999_b0 , \323_b0 , w_1859 );
and ( w_1858 , w_1859 , \602_b0 );
or ( \1000_b1 , \998_b1 , w_1861 );
not ( w_1861 , w_1862 );
and ( \1000_b0 , \998_b0 , w_1863 );
and ( w_1862 ,  , w_1863 );
buf ( w_1861 , \999_b1 );
not ( w_1861 , w_1864 );
not (  , w_1865 );
and ( w_1864 , w_1865 , \999_b0 );
or ( \1001_b1 , \1000_b1 , w_1866 );
xor ( \1001_b0 , \1000_b0 , w_1868 );
not ( w_1868 , w_1869 );
and ( w_1869 , w_1866 , w_1867 );
buf ( w_1866 , \561_b1 );
not ( w_1866 , w_1870 );
not ( w_1867 , w_1871 );
and ( w_1870 , w_1871 , \561_b0 );
or ( \1002_b1 , \360_b1 , \503_b1 );
not ( \503_b1 , w_1872 );
and ( \1002_b0 , \360_b0 , w_1873 );
and ( w_1872 , w_1873 , \503_b0 );
or ( \1003_b1 , \343_b1 , \501_b1 );
not ( \501_b1 , w_1874 );
and ( \1003_b0 , \343_b0 , w_1875 );
and ( w_1874 , w_1875 , \501_b0 );
or ( \1004_b1 , \1002_b1 , w_1877 );
not ( w_1877 , w_1878 );
and ( \1004_b0 , \1002_b0 , w_1879 );
and ( w_1878 ,  , w_1879 );
buf ( w_1877 , \1003_b1 );
not ( w_1877 , w_1880 );
not (  , w_1881 );
and ( w_1880 , w_1881 , \1003_b0 );
or ( \1005_b1 , \1004_b1 , w_1882 );
xor ( \1005_b0 , \1004_b0 , w_1884 );
not ( w_1884 , w_1885 );
and ( w_1885 , w_1882 , w_1883 );
buf ( w_1882 , \455_b1 );
not ( w_1882 , w_1886 );
not ( w_1883 , w_1887 );
and ( w_1886 , w_1887 , \455_b0 );
or ( \1006_b1 , \1001_b1 , \1005_b1 );
not ( \1005_b1 , w_1888 );
and ( \1006_b0 , \1001_b0 , w_1889 );
and ( w_1888 , w_1889 , \1005_b0 );
or ( \1007_b1 , \495_b1 , \298_b1 );
not ( \298_b1 , w_1890 );
and ( \1007_b0 , \495_b0 , w_1891 );
and ( w_1890 , w_1891 , \298_b0 );
or ( \1008_b1 , \444_b1 , \296_b1 );
not ( \296_b1 , w_1892 );
and ( \1008_b0 , \444_b0 , w_1893 );
and ( w_1892 , w_1893 , \296_b0 );
or ( \1009_b1 , \1007_b1 , w_1895 );
not ( w_1895 , w_1896 );
and ( \1009_b0 , \1007_b0 , w_1897 );
and ( w_1896 ,  , w_1897 );
buf ( w_1895 , \1008_b1 );
not ( w_1895 , w_1898 );
not (  , w_1899 );
and ( w_1898 , w_1899 , \1008_b0 );
or ( \1010_b1 , \1009_b1 , w_1900 );
xor ( \1010_b0 , \1009_b0 , w_1902 );
not ( w_1902 , w_1903 );
and ( w_1903 , w_1900 , w_1901 );
buf ( w_1900 , \303_b1 );
not ( w_1900 , w_1904 );
not ( w_1901 , w_1905 );
and ( w_1904 , w_1905 , \303_b0 );
or ( \1011_b1 , \1005_b1 , \1010_b1 );
not ( \1010_b1 , w_1906 );
and ( \1011_b0 , \1005_b0 , w_1907 );
and ( w_1906 , w_1907 , \1010_b0 );
or ( \1012_b1 , \1001_b1 , \1010_b1 );
not ( \1010_b1 , w_1908 );
and ( \1012_b0 , \1001_b0 , w_1909 );
and ( w_1908 , w_1909 , \1010_b0 );
or ( \1014_b1 , \997_b1 , \1013_b1 );
not ( \1013_b1 , w_1910 );
and ( \1014_b0 , \997_b0 , w_1911 );
and ( w_1910 , w_1911 , \1013_b0 );
or ( \1015_b1 , \621_b1 , \313_b1 );
not ( \313_b1 , w_1912 );
and ( \1015_b0 , \621_b0 , w_1913 );
and ( w_1912 , w_1913 , \313_b0 );
or ( \1016_b1 , \593_b1 , \311_b1 );
not ( \311_b1 , w_1914 );
and ( \1016_b0 , \593_b0 , w_1915 );
and ( w_1914 , w_1915 , \311_b0 );
or ( \1017_b1 , \1015_b1 , w_1917 );
not ( w_1917 , w_1918 );
and ( \1017_b0 , \1015_b0 , w_1919 );
and ( w_1918 ,  , w_1919 );
buf ( w_1917 , \1016_b1 );
not ( w_1917 , w_1920 );
not (  , w_1921 );
and ( w_1920 , w_1921 , \1016_b0 );
or ( \1018_b1 , \1017_b1 , w_1922 );
xor ( \1018_b0 , \1017_b0 , w_1924 );
not ( w_1924 , w_1925 );
and ( w_1925 , w_1922 , w_1923 );
buf ( w_1922 , \320_b1 );
not ( w_1922 , w_1926 );
not ( w_1923 , w_1927 );
and ( w_1926 , w_1927 , \320_b0 );
or ( \1019_b1 , \777_b1 , \331_b1 );
not ( \331_b1 , w_1928 );
and ( \1019_b0 , \777_b0 , w_1929 );
and ( w_1928 , w_1929 , \331_b0 );
or ( \1020_b1 , \703_b1 , \329_b1 );
not ( \329_b1 , w_1930 );
and ( \1020_b0 , \703_b0 , w_1931 );
and ( w_1930 , w_1931 , \329_b0 );
or ( \1021_b1 , \1019_b1 , w_1933 );
not ( w_1933 , w_1934 );
and ( \1021_b0 , \1019_b0 , w_1935 );
and ( w_1934 ,  , w_1935 );
buf ( w_1933 , \1020_b1 );
not ( w_1933 , w_1936 );
not (  , w_1937 );
and ( w_1936 , w_1937 , \1020_b0 );
or ( \1022_b1 , \1021_b1 , w_1938 );
xor ( \1022_b0 , \1021_b0 , w_1940 );
not ( w_1940 , w_1941 );
and ( w_1941 , w_1938 , w_1939 );
buf ( w_1938 , \338_b1 );
not ( w_1938 , w_1942 );
not ( w_1939 , w_1943 );
and ( w_1942 , w_1943 , \338_b0 );
or ( \1023_b1 , \1018_b1 , \1022_b1 );
not ( \1022_b1 , w_1944 );
and ( \1023_b0 , \1018_b0 , w_1945 );
and ( w_1944 , w_1945 , \1022_b0 );
or ( \1024_b1 , \904_b1 , \351_b1 );
not ( \351_b1 , w_1946 );
and ( \1024_b0 , \904_b0 , w_1947 );
and ( w_1946 , w_1947 , \351_b0 );
or ( \1025_b1 , \841_b1 , \349_b1 );
not ( \349_b1 , w_1948 );
and ( \1025_b0 , \841_b0 , w_1949 );
and ( w_1948 , w_1949 , \349_b0 );
or ( \1026_b1 , \1024_b1 , w_1951 );
not ( w_1951 , w_1952 );
and ( \1026_b0 , \1024_b0 , w_1953 );
and ( w_1952 ,  , w_1953 );
buf ( w_1951 , \1025_b1 );
not ( w_1951 , w_1954 );
not (  , w_1955 );
and ( w_1954 , w_1955 , \1025_b0 );
or ( \1027_b1 , \1026_b1 , w_1956 );
xor ( \1027_b0 , \1026_b0 , w_1958 );
not ( w_1958 , w_1959 );
and ( w_1959 , w_1956 , w_1957 );
buf ( w_1956 , \358_b1 );
not ( w_1956 , w_1960 );
not ( w_1957 , w_1961 );
and ( w_1960 , w_1961 , \358_b0 );
or ( \1028_b1 , \1022_b1 , \1027_b1 );
not ( \1027_b1 , w_1962 );
and ( \1028_b0 , \1022_b0 , w_1963 );
and ( w_1962 , w_1963 , \1027_b0 );
or ( \1029_b1 , \1018_b1 , \1027_b1 );
not ( \1027_b1 , w_1964 );
and ( \1029_b0 , \1018_b0 , w_1965 );
and ( w_1964 , w_1965 , \1027_b0 );
or ( \1031_b1 , \1013_b1 , \1030_b1 );
not ( \1030_b1 , w_1966 );
and ( \1031_b0 , \1013_b0 , w_1967 );
and ( w_1966 , w_1967 , \1030_b0 );
or ( \1032_b1 , \997_b1 , \1030_b1 );
not ( \1030_b1 , w_1968 );
and ( \1032_b0 , \997_b0 , w_1969 );
and ( w_1968 , w_1969 , \1030_b0 );
or ( \1034_b1 , \898_b1 , \902_b1 );
xor ( \1034_b0 , \898_b0 , w_1970 );
not ( w_1970 , w_1971 );
and ( w_1971 , \902_b1 , \902_b0 );
or ( \1035_b1 , \1034_b1 , \905_b1 );
xor ( \1035_b0 , \1034_b0 , w_1972 );
not ( w_1972 , w_1973 );
and ( w_1973 , \905_b1 , \905_b0 );
or ( \1036_b1 , \932_b1 , \936_b1 );
xor ( \1036_b0 , \932_b0 , w_1974 );
not ( w_1974 , w_1975 );
and ( w_1975 , \936_b1 , \936_b0 );
or ( \1037_b1 , \1036_b1 , \941_b1 );
xor ( \1037_b0 , \1036_b0 , w_1976 );
not ( w_1976 , w_1977 );
and ( w_1977 , \941_b1 , \941_b0 );
or ( \1038_b1 , \1035_b1 , w_1978 );
or ( \1038_b0 , \1035_b0 , \1037_b0 );
not ( \1037_b0 , w_1979 );
and ( w_1979 , w_1978 , \1037_b1 );
or ( \1039_b1 , \1033_b1 , \1038_b1 );
not ( \1038_b1 , w_1980 );
and ( \1039_b0 , \1033_b0 , w_1981 );
and ( w_1980 , w_1981 , \1038_b0 );
or ( \1040_b1 , \949_b1 , \951_b1 );
xor ( \1040_b0 , \949_b0 , w_1982 );
not ( w_1982 , w_1983 );
and ( w_1983 , \951_b1 , \951_b0 );
or ( \1041_b1 , \1040_b1 , \954_b1 );
xor ( \1041_b0 , \1040_b0 , w_1984 );
not ( w_1984 , w_1985 );
and ( w_1985 , \954_b1 , \954_b0 );
or ( \1042_b1 , \1038_b1 , \1041_b1 );
not ( \1041_b1 , w_1986 );
and ( \1042_b0 , \1038_b0 , w_1987 );
and ( w_1986 , w_1987 , \1041_b0 );
or ( \1043_b1 , \1033_b1 , \1041_b1 );
not ( \1041_b1 , w_1988 );
and ( \1043_b0 , \1033_b0 , w_1989 );
and ( w_1988 , w_1989 , \1041_b0 );
or ( \1045_b1 , \831_b1 , \845_b1 );
xor ( \1045_b0 , \831_b0 , w_1990 );
not ( w_1990 , w_1991 );
and ( w_1991 , \845_b1 , \845_b0 );
or ( \1046_b1 , \1045_b1 , \862_b1 );
xor ( \1046_b0 , \1045_b0 , w_1992 );
not ( w_1992 , w_1993 );
and ( w_1993 , \862_b1 , \862_b0 );
or ( \1047_b1 , \1044_b1 , \1046_b1 );
not ( \1046_b1 , w_1994 );
and ( \1047_b0 , \1044_b0 , w_1995 );
and ( w_1994 , w_1995 , \1046_b0 );
or ( \1048_b1 , \947_b1 , \957_b1 );
xor ( \1048_b0 , \947_b0 , w_1996 );
not ( w_1996 , w_1997 );
and ( w_1997 , \957_b1 , \957_b0 );
or ( \1049_b1 , \1048_b1 , \960_b1 );
xor ( \1049_b0 , \1048_b0 , w_1998 );
not ( w_1998 , w_1999 );
and ( w_1999 , \960_b1 , \960_b0 );
or ( \1050_b1 , \1046_b1 , \1049_b1 );
not ( \1049_b1 , w_2000 );
and ( \1050_b0 , \1046_b0 , w_2001 );
and ( w_2000 , w_2001 , \1049_b0 );
or ( \1051_b1 , \1044_b1 , \1049_b1 );
not ( \1049_b1 , w_2002 );
and ( \1051_b0 , \1044_b0 , w_2003 );
and ( w_2002 , w_2003 , \1049_b0 );
or ( \1053_b1 , \963_b1 , \965_b1 );
xor ( \1053_b0 , \963_b0 , w_2004 );
not ( w_2004 , w_2005 );
and ( w_2005 , \965_b1 , \965_b0 );
or ( \1054_b1 , \1053_b1 , \968_b1 );
xor ( \1054_b0 , \1053_b0 , w_2006 );
not ( w_2006 , w_2007 );
and ( w_2007 , \968_b1 , \968_b0 );
or ( \1055_b1 , \1052_b1 , \1054_b1 );
not ( \1054_b1 , w_2008 );
and ( \1055_b0 , \1052_b0 , w_2009 );
and ( w_2008 , w_2009 , \1054_b0 );
or ( \1056_b1 , \977_b1 , \1055_b1 );
not ( \1055_b1 , w_2010 );
and ( \1056_b0 , \977_b0 , w_2011 );
and ( w_2010 , w_2011 , \1055_b0 );
or ( \1057_b1 , \977_b1 , \1055_b1 );
xor ( \1057_b0 , \977_b0 , w_2012 );
not ( w_2012 , w_2013 );
and ( w_2013 , \1055_b1 , \1055_b0 );
or ( \1058_b1 , \1052_b1 , \1054_b1 );
xor ( \1058_b0 , \1052_b0 , w_2014 );
not ( w_2014 , w_2015 );
and ( w_2015 , \1054_b1 , \1054_b0 );
or ( \1059_b1 , \815_b1 , \979_b1 );
xor ( \1059_b0 , \815_b0 , w_2016 );
not ( w_2016 , w_2017 );
and ( w_2017 , \979_b1 , \979_b0 );
or ( \1060_b1 , \979_b1 , \981_b1 );
xor ( \1060_b0 , \979_b0 , w_2018 );
not ( w_2018 , w_2019 );
and ( w_2019 , \981_b1 , \981_b0 );
buf ( \1061_b1 , \1060_b1 );
not ( \1061_b1 , w_2020 );
not ( \1061_b0 , w_2021 );
and ( w_2020 , w_2021 , \1060_b0 );
or ( \1062_b1 , \1059_b1 , \1061_b1 );
not ( \1061_b1 , w_2022 );
and ( \1062_b0 , \1059_b0 , w_2023 );
and ( w_2022 , w_2023 , \1061_b0 );
or ( \1063_b1 , \159_b1 , \1062_b1 );
not ( \1062_b1 , w_2024 );
and ( \1063_b0 , \159_b0 , w_2025 );
and ( w_2024 , w_2025 , \1062_b0 );
buf ( \1064_b1 , \1063_b1 );
not ( \1064_b1 , w_2026 );
not ( \1064_b0 , w_2027 );
and ( w_2026 , w_2027 , \1063_b0 );
or ( \1065_b1 , \1064_b1 , w_2028 );
xor ( \1065_b0 , \1064_b0 , w_2030 );
not ( w_2030 , w_2031 );
and ( w_2031 , w_2028 , w_2029 );
buf ( w_2028 , \984_b1 );
not ( w_2028 , w_2032 );
not ( w_2029 , w_2033 );
and ( w_2032 , w_2033 , \984_b0 );
or ( \1066_b1 , \305_b1 , \912_b1 );
not ( \912_b1 , w_2034 );
and ( \1066_b0 , \305_b0 , w_2035 );
and ( w_2034 , w_2035 , \912_b0 );
or ( \1067_b1 , \315_b1 , \910_b1 );
not ( \910_b1 , w_2036 );
and ( \1067_b0 , \315_b0 , w_2037 );
and ( w_2036 , w_2037 , \910_b0 );
or ( \1068_b1 , \1066_b1 , w_2039 );
not ( w_2039 , w_2040 );
and ( \1068_b0 , \1066_b0 , w_2041 );
and ( w_2040 ,  , w_2041 );
buf ( w_2039 , \1067_b1 );
not ( w_2039 , w_2042 );
not (  , w_2043 );
and ( w_2042 , w_2043 , \1067_b0 );
or ( \1069_b1 , \1068_b1 , w_2044 );
xor ( \1069_b0 , \1068_b0 , w_2046 );
not ( w_2046 , w_2047 );
and ( w_2047 , w_2044 , w_2045 );
buf ( w_2044 , \818_b1 );
not ( w_2044 , w_2048 );
not ( w_2045 , w_2049 );
and ( w_2048 , w_2049 , \818_b0 );
or ( \1070_b1 , \1065_b1 , \1069_b1 );
not ( \1069_b1 , w_2050 );
and ( \1070_b0 , \1065_b0 , w_2051 );
and ( w_2050 , w_2051 , \1069_b0 );
or ( \1071_b1 , \323_b1 , \740_b1 );
not ( \740_b1 , w_2052 );
and ( \1071_b0 , \323_b0 , w_2053 );
and ( w_2052 , w_2053 , \740_b0 );
or ( \1072_b1 , \333_b1 , \738_b1 );
not ( \738_b1 , w_2054 );
and ( \1072_b0 , \333_b0 , w_2055 );
and ( w_2054 , w_2055 , \738_b0 );
or ( \1073_b1 , \1071_b1 , w_2057 );
not ( w_2057 , w_2058 );
and ( \1073_b0 , \1071_b0 , w_2059 );
and ( w_2058 ,  , w_2059 );
buf ( w_2057 , \1072_b1 );
not ( w_2057 , w_2060 );
not (  , w_2061 );
and ( w_2060 , w_2061 , \1072_b0 );
or ( \1074_b1 , \1073_b1 , w_2062 );
xor ( \1074_b0 , \1073_b0 , w_2064 );
not ( w_2064 , w_2065 );
and ( w_2065 , w_2062 , w_2063 );
buf ( w_2062 , \668_b1 );
not ( w_2062 , w_2066 );
not ( w_2063 , w_2067 );
and ( w_2066 , w_2067 , \668_b0 );
or ( \1075_b1 , \1069_b1 , \1074_b1 );
not ( \1074_b1 , w_2068 );
and ( \1075_b0 , \1069_b0 , w_2069 );
and ( w_2068 , w_2069 , \1074_b0 );
or ( \1076_b1 , \1065_b1 , \1074_b1 );
not ( \1074_b1 , w_2070 );
and ( \1076_b0 , \1065_b0 , w_2071 );
and ( w_2070 , w_2071 , \1074_b0 );
or ( \1078_b1 , \343_b1 , \604_b1 );
not ( \604_b1 , w_2072 );
and ( \1078_b0 , \343_b0 , w_2073 );
and ( w_2072 , w_2073 , \604_b0 );
or ( \1079_b1 , \353_b1 , \602_b1 );
not ( \602_b1 , w_2074 );
and ( \1079_b0 , \353_b0 , w_2075 );
and ( w_2074 , w_2075 , \602_b0 );
or ( \1080_b1 , \1078_b1 , w_2077 );
not ( w_2077 , w_2078 );
and ( \1080_b0 , \1078_b0 , w_2079 );
and ( w_2078 ,  , w_2079 );
buf ( w_2077 , \1079_b1 );
not ( w_2077 , w_2080 );
not (  , w_2081 );
and ( w_2080 , w_2081 , \1079_b0 );
or ( \1081_b1 , \1080_b1 , w_2082 );
xor ( \1081_b0 , \1080_b0 , w_2084 );
not ( w_2084 , w_2085 );
and ( w_2085 , w_2082 , w_2083 );
buf ( w_2082 , \561_b1 );
not ( w_2082 , w_2086 );
not ( w_2083 , w_2087 );
and ( w_2086 , w_2087 , \561_b0 );
or ( \1082_b1 , \444_b1 , \503_b1 );
not ( \503_b1 , w_2088 );
and ( \1082_b0 , \444_b0 , w_2089 );
and ( w_2088 , w_2089 , \503_b0 );
or ( \1083_b1 , \360_b1 , \501_b1 );
not ( \501_b1 , w_2090 );
and ( \1083_b0 , \360_b0 , w_2091 );
and ( w_2090 , w_2091 , \501_b0 );
or ( \1084_b1 , \1082_b1 , w_2093 );
not ( w_2093 , w_2094 );
and ( \1084_b0 , \1082_b0 , w_2095 );
and ( w_2094 ,  , w_2095 );
buf ( w_2093 , \1083_b1 );
not ( w_2093 , w_2096 );
not (  , w_2097 );
and ( w_2096 , w_2097 , \1083_b0 );
or ( \1085_b1 , \1084_b1 , w_2098 );
xor ( \1085_b0 , \1084_b0 , w_2100 );
not ( w_2100 , w_2101 );
and ( w_2101 , w_2098 , w_2099 );
buf ( w_2098 , \455_b1 );
not ( w_2098 , w_2102 );
not ( w_2099 , w_2103 );
and ( w_2102 , w_2103 , \455_b0 );
or ( \1086_b1 , \1081_b1 , \1085_b1 );
not ( \1085_b1 , w_2104 );
and ( \1086_b0 , \1081_b0 , w_2105 );
and ( w_2104 , w_2105 , \1085_b0 );
or ( \1087_b1 , \593_b1 , \298_b1 );
not ( \298_b1 , w_2106 );
and ( \1087_b0 , \593_b0 , w_2107 );
and ( w_2106 , w_2107 , \298_b0 );
or ( \1088_b1 , \495_b1 , \296_b1 );
not ( \296_b1 , w_2108 );
and ( \1088_b0 , \495_b0 , w_2109 );
and ( w_2108 , w_2109 , \296_b0 );
or ( \1089_b1 , \1087_b1 , w_2111 );
not ( w_2111 , w_2112 );
and ( \1089_b0 , \1087_b0 , w_2113 );
and ( w_2112 ,  , w_2113 );
buf ( w_2111 , \1088_b1 );
not ( w_2111 , w_2114 );
not (  , w_2115 );
and ( w_2114 , w_2115 , \1088_b0 );
or ( \1090_b1 , \1089_b1 , w_2116 );
xor ( \1090_b0 , \1089_b0 , w_2118 );
not ( w_2118 , w_2119 );
and ( w_2119 , w_2116 , w_2117 );
buf ( w_2116 , \303_b1 );
not ( w_2116 , w_2120 );
not ( w_2117 , w_2121 );
and ( w_2120 , w_2121 , \303_b0 );
or ( \1091_b1 , \1085_b1 , \1090_b1 );
not ( \1090_b1 , w_2122 );
and ( \1091_b0 , \1085_b0 , w_2123 );
and ( w_2122 , w_2123 , \1090_b0 );
or ( \1092_b1 , \1081_b1 , \1090_b1 );
not ( \1090_b1 , w_2124 );
and ( \1092_b0 , \1081_b0 , w_2125 );
and ( w_2124 , w_2125 , \1090_b0 );
or ( \1094_b1 , \1077_b1 , \1093_b1 );
not ( \1093_b1 , w_2126 );
and ( \1094_b0 , \1077_b0 , w_2127 );
and ( w_2126 , w_2127 , \1093_b0 );
or ( \1095_b1 , \703_b1 , \313_b1 );
not ( \313_b1 , w_2128 );
and ( \1095_b0 , \703_b0 , w_2129 );
and ( w_2128 , w_2129 , \313_b0 );
or ( \1096_b1 , \621_b1 , \311_b1 );
not ( \311_b1 , w_2130 );
and ( \1096_b0 , \621_b0 , w_2131 );
and ( w_2130 , w_2131 , \311_b0 );
or ( \1097_b1 , \1095_b1 , w_2133 );
not ( w_2133 , w_2134 );
and ( \1097_b0 , \1095_b0 , w_2135 );
and ( w_2134 ,  , w_2135 );
buf ( w_2133 , \1096_b1 );
not ( w_2133 , w_2136 );
not (  , w_2137 );
and ( w_2136 , w_2137 , \1096_b0 );
or ( \1098_b1 , \1097_b1 , w_2138 );
xor ( \1098_b0 , \1097_b0 , w_2140 );
not ( w_2140 , w_2141 );
and ( w_2141 , w_2138 , w_2139 );
buf ( w_2138 , \320_b1 );
not ( w_2138 , w_2142 );
not ( w_2139 , w_2143 );
and ( w_2142 , w_2143 , \320_b0 );
or ( \1099_b1 , \841_b1 , \331_b1 );
not ( \331_b1 , w_2144 );
and ( \1099_b0 , \841_b0 , w_2145 );
and ( w_2144 , w_2145 , \331_b0 );
or ( \1100_b1 , \777_b1 , \329_b1 );
not ( \329_b1 , w_2146 );
and ( \1100_b0 , \777_b0 , w_2147 );
and ( w_2146 , w_2147 , \329_b0 );
or ( \1101_b1 , \1099_b1 , w_2149 );
not ( w_2149 , w_2150 );
and ( \1101_b0 , \1099_b0 , w_2151 );
and ( w_2150 ,  , w_2151 );
buf ( w_2149 , \1100_b1 );
not ( w_2149 , w_2152 );
not (  , w_2153 );
and ( w_2152 , w_2153 , \1100_b0 );
or ( \1102_b1 , \1101_b1 , w_2154 );
xor ( \1102_b0 , \1101_b0 , w_2156 );
not ( w_2156 , w_2157 );
and ( w_2157 , w_2154 , w_2155 );
buf ( w_2154 , \338_b1 );
not ( w_2154 , w_2158 );
not ( w_2155 , w_2159 );
and ( w_2158 , w_2159 , \338_b0 );
or ( \1103_b1 , \1098_b1 , \1102_b1 );
not ( \1102_b1 , w_2160 );
and ( \1103_b0 , \1098_b0 , w_2161 );
and ( w_2160 , w_2161 , \1102_b0 );
buf ( \1104_b1 , RIb4bf2b8_81_b1 );
buf ( \1104_b0 , RIb4bf2b8_81_b0 );
or ( \1105_b1 , \1104_b1 , \351_b1 );
not ( \351_b1 , w_2162 );
and ( \1105_b0 , \1104_b0 , w_2163 );
and ( w_2162 , w_2163 , \351_b0 );
or ( \1106_b1 , \904_b1 , \349_b1 );
not ( \349_b1 , w_2164 );
and ( \1106_b0 , \904_b0 , w_2165 );
and ( w_2164 , w_2165 , \349_b0 );
or ( \1107_b1 , \1105_b1 , w_2167 );
not ( w_2167 , w_2168 );
and ( \1107_b0 , \1105_b0 , w_2169 );
and ( w_2168 ,  , w_2169 );
buf ( w_2167 , \1106_b1 );
not ( w_2167 , w_2170 );
not (  , w_2171 );
and ( w_2170 , w_2171 , \1106_b0 );
or ( \1108_b1 , \1107_b1 , w_2172 );
xor ( \1108_b0 , \1107_b0 , w_2174 );
not ( w_2174 , w_2175 );
and ( w_2175 , w_2172 , w_2173 );
buf ( w_2172 , \358_b1 );
not ( w_2172 , w_2176 );
not ( w_2173 , w_2177 );
and ( w_2176 , w_2177 , \358_b0 );
or ( \1109_b1 , \1102_b1 , \1108_b1 );
not ( \1108_b1 , w_2178 );
and ( \1109_b0 , \1102_b0 , w_2179 );
and ( w_2178 , w_2179 , \1108_b0 );
or ( \1110_b1 , \1098_b1 , \1108_b1 );
not ( \1108_b1 , w_2180 );
and ( \1110_b0 , \1098_b0 , w_2181 );
and ( w_2180 , w_2181 , \1108_b0 );
or ( \1112_b1 , \1093_b1 , \1111_b1 );
not ( \1111_b1 , w_2182 );
and ( \1112_b0 , \1093_b0 , w_2183 );
and ( w_2182 , w_2183 , \1111_b0 );
or ( \1113_b1 , \1077_b1 , \1111_b1 );
not ( \1111_b1 , w_2184 );
and ( \1113_b0 , \1077_b0 , w_2185 );
and ( w_2184 , w_2185 , \1111_b0 );
or ( \1115_b1 , \1104_b1 , \345_b1 );
not ( \345_b1 , w_2186 );
and ( \1115_b0 , \1104_b0 , w_2187 );
and ( w_2186 , w_2187 , \345_b0 );
or ( \1116_b1 , \1001_b1 , \1005_b1 );
xor ( \1116_b0 , \1001_b0 , w_2188 );
not ( w_2188 , w_2189 );
and ( w_2189 , \1005_b1 , \1005_b0 );
or ( \1117_b1 , \1116_b1 , \1010_b1 );
xor ( \1117_b0 , \1116_b0 , w_2190 );
not ( w_2190 , w_2191 );
and ( w_2191 , \1010_b1 , \1010_b0 );
or ( \1118_b1 , \1115_b1 , \1117_b1 );
not ( \1117_b1 , w_2192 );
and ( \1118_b0 , \1115_b0 , w_2193 );
and ( w_2192 , w_2193 , \1117_b0 );
or ( \1119_b1 , \1018_b1 , \1022_b1 );
xor ( \1119_b0 , \1018_b0 , w_2194 );
not ( w_2194 , w_2195 );
and ( w_2195 , \1022_b1 , \1022_b0 );
or ( \1120_b1 , \1119_b1 , \1027_b1 );
xor ( \1120_b0 , \1119_b0 , w_2196 );
not ( w_2196 , w_2197 );
and ( w_2197 , \1027_b1 , \1027_b0 );
or ( \1121_b1 , \1117_b1 , \1120_b1 );
not ( \1120_b1 , w_2198 );
and ( \1121_b0 , \1117_b0 , w_2199 );
and ( w_2198 , w_2199 , \1120_b0 );
or ( \1122_b1 , \1115_b1 , \1120_b1 );
not ( \1120_b1 , w_2200 );
and ( \1122_b0 , \1115_b0 , w_2201 );
and ( w_2200 , w_2201 , \1120_b0 );
or ( \1124_b1 , \1114_b1 , \1123_b1 );
not ( \1123_b1 , w_2202 );
and ( \1124_b0 , \1114_b0 , w_2203 );
and ( w_2202 , w_2203 , \1123_b0 );
or ( \1125_b1 , \915_b1 , \919_b1 );
xor ( \1125_b0 , \915_b0 , w_2204 );
not ( w_2204 , w_2205 );
and ( w_2205 , \919_b1 , \919_b0 );
or ( \1126_b1 , \1125_b1 , \924_b1 );
xor ( \1126_b0 , \1125_b0 , w_2206 );
not ( w_2206 , w_2207 );
and ( w_2207 , \924_b1 , \924_b0 );
or ( \1127_b1 , \1123_b1 , \1126_b1 );
not ( \1126_b1 , w_2208 );
and ( \1127_b0 , \1123_b0 , w_2209 );
and ( w_2208 , w_2209 , \1126_b0 );
or ( \1128_b1 , \1114_b1 , \1126_b1 );
not ( \1126_b1 , w_2210 );
and ( \1128_b0 , \1114_b0 , w_2211 );
and ( w_2210 , w_2211 , \1126_b0 );
or ( \1130_b1 , \908_b1 , \927_b1 );
xor ( \1130_b0 , \908_b0 , w_2212 );
not ( w_2212 , w_2213 );
and ( w_2213 , \927_b1 , \927_b0 );
or ( \1131_b1 , \1130_b1 , \944_b1 );
xor ( \1131_b0 , \1130_b0 , w_2214 );
not ( w_2214 , w_2215 );
and ( w_2215 , \944_b1 , \944_b0 );
or ( \1132_b1 , \1129_b1 , \1131_b1 );
not ( \1131_b1 , w_2216 );
and ( \1132_b0 , \1129_b0 , w_2217 );
and ( w_2216 , w_2217 , \1131_b0 );
or ( \1133_b1 , \1033_b1 , \1038_b1 );
xor ( \1133_b0 , \1033_b0 , w_2218 );
not ( w_2218 , w_2219 );
and ( w_2219 , \1038_b1 , \1038_b0 );
or ( \1134_b1 , \1133_b1 , \1041_b1 );
xor ( \1134_b0 , \1133_b0 , w_2220 );
not ( w_2220 , w_2221 );
and ( w_2221 , \1041_b1 , \1041_b0 );
or ( \1135_b1 , \1131_b1 , \1134_b1 );
not ( \1134_b1 , w_2222 );
and ( \1135_b0 , \1131_b0 , w_2223 );
and ( w_2222 , w_2223 , \1134_b0 );
or ( \1136_b1 , \1129_b1 , \1134_b1 );
not ( \1134_b1 , w_2224 );
and ( \1136_b0 , \1129_b0 , w_2225 );
and ( w_2224 , w_2225 , \1134_b0 );
or ( \1138_b1 , \353_b1 , \740_b1 );
not ( \740_b1 , w_2226 );
and ( \1138_b0 , \353_b0 , w_2227 );
and ( w_2226 , w_2227 , \740_b0 );
or ( \1139_b1 , \323_b1 , \738_b1 );
not ( \738_b1 , w_2228 );
and ( \1139_b0 , \323_b0 , w_2229 );
and ( w_2228 , w_2229 , \738_b0 );
or ( \1140_b1 , \1138_b1 , w_2231 );
not ( w_2231 , w_2232 );
and ( \1140_b0 , \1138_b0 , w_2233 );
and ( w_2232 ,  , w_2233 );
buf ( w_2231 , \1139_b1 );
not ( w_2231 , w_2234 );
not (  , w_2235 );
and ( w_2234 , w_2235 , \1139_b0 );
or ( \1141_b1 , \1140_b1 , w_2236 );
xor ( \1141_b0 , \1140_b0 , w_2238 );
not ( w_2238 , w_2239 );
and ( w_2239 , w_2236 , w_2237 );
buf ( w_2236 , \668_b1 );
not ( w_2236 , w_2240 );
not ( w_2237 , w_2241 );
and ( w_2240 , w_2241 , \668_b0 );
or ( \1142_b1 , \360_b1 , \604_b1 );
not ( \604_b1 , w_2242 );
and ( \1142_b0 , \360_b0 , w_2243 );
and ( w_2242 , w_2243 , \604_b0 );
or ( \1143_b1 , \343_b1 , \602_b1 );
not ( \602_b1 , w_2244 );
and ( \1143_b0 , \343_b0 , w_2245 );
and ( w_2244 , w_2245 , \602_b0 );
or ( \1144_b1 , \1142_b1 , w_2247 );
not ( w_2247 , w_2248 );
and ( \1144_b0 , \1142_b0 , w_2249 );
and ( w_2248 ,  , w_2249 );
buf ( w_2247 , \1143_b1 );
not ( w_2247 , w_2250 );
not (  , w_2251 );
and ( w_2250 , w_2251 , \1143_b0 );
or ( \1145_b1 , \1144_b1 , w_2252 );
xor ( \1145_b0 , \1144_b0 , w_2254 );
not ( w_2254 , w_2255 );
and ( w_2255 , w_2252 , w_2253 );
buf ( w_2252 , \561_b1 );
not ( w_2252 , w_2256 );
not ( w_2253 , w_2257 );
and ( w_2256 , w_2257 , \561_b0 );
or ( \1146_b1 , \1141_b1 , \1145_b1 );
not ( \1145_b1 , w_2258 );
and ( \1146_b0 , \1141_b0 , w_2259 );
and ( w_2258 , w_2259 , \1145_b0 );
or ( \1147_b1 , \495_b1 , \503_b1 );
not ( \503_b1 , w_2260 );
and ( \1147_b0 , \495_b0 , w_2261 );
and ( w_2260 , w_2261 , \503_b0 );
or ( \1148_b1 , \444_b1 , \501_b1 );
not ( \501_b1 , w_2262 );
and ( \1148_b0 , \444_b0 , w_2263 );
and ( w_2262 , w_2263 , \501_b0 );
or ( \1149_b1 , \1147_b1 , w_2265 );
not ( w_2265 , w_2266 );
and ( \1149_b0 , \1147_b0 , w_2267 );
and ( w_2266 ,  , w_2267 );
buf ( w_2265 , \1148_b1 );
not ( w_2265 , w_2268 );
not (  , w_2269 );
and ( w_2268 , w_2269 , \1148_b0 );
or ( \1150_b1 , \1149_b1 , w_2270 );
xor ( \1150_b0 , \1149_b0 , w_2272 );
not ( w_2272 , w_2273 );
and ( w_2273 , w_2270 , w_2271 );
buf ( w_2270 , \455_b1 );
not ( w_2270 , w_2274 );
not ( w_2271 , w_2275 );
and ( w_2274 , w_2275 , \455_b0 );
or ( \1151_b1 , \1145_b1 , \1150_b1 );
not ( \1150_b1 , w_2276 );
and ( \1151_b0 , \1145_b0 , w_2277 );
and ( w_2276 , w_2277 , \1150_b0 );
or ( \1152_b1 , \1141_b1 , \1150_b1 );
not ( \1150_b1 , w_2278 );
and ( \1152_b0 , \1141_b0 , w_2279 );
and ( w_2278 , w_2279 , \1150_b0 );
or ( \1154_b1 , \621_b1 , \298_b1 );
not ( \298_b1 , w_2280 );
and ( \1154_b0 , \621_b0 , w_2281 );
and ( w_2280 , w_2281 , \298_b0 );
or ( \1155_b1 , \593_b1 , \296_b1 );
not ( \296_b1 , w_2282 );
and ( \1155_b0 , \593_b0 , w_2283 );
and ( w_2282 , w_2283 , \296_b0 );
or ( \1156_b1 , \1154_b1 , w_2285 );
not ( w_2285 , w_2286 );
and ( \1156_b0 , \1154_b0 , w_2287 );
and ( w_2286 ,  , w_2287 );
buf ( w_2285 , \1155_b1 );
not ( w_2285 , w_2288 );
not (  , w_2289 );
and ( w_2288 , w_2289 , \1155_b0 );
or ( \1157_b1 , \1156_b1 , w_2290 );
xor ( \1157_b0 , \1156_b0 , w_2292 );
not ( w_2292 , w_2293 );
and ( w_2293 , w_2290 , w_2291 );
buf ( w_2290 , \303_b1 );
not ( w_2290 , w_2294 );
not ( w_2291 , w_2295 );
and ( w_2294 , w_2295 , \303_b0 );
or ( \1158_b1 , \777_b1 , \313_b1 );
not ( \313_b1 , w_2296 );
and ( \1158_b0 , \777_b0 , w_2297 );
and ( w_2296 , w_2297 , \313_b0 );
or ( \1159_b1 , \703_b1 , \311_b1 );
not ( \311_b1 , w_2298 );
and ( \1159_b0 , \703_b0 , w_2299 );
and ( w_2298 , w_2299 , \311_b0 );
or ( \1160_b1 , \1158_b1 , w_2301 );
not ( w_2301 , w_2302 );
and ( \1160_b0 , \1158_b0 , w_2303 );
and ( w_2302 ,  , w_2303 );
buf ( w_2301 , \1159_b1 );
not ( w_2301 , w_2304 );
not (  , w_2305 );
and ( w_2304 , w_2305 , \1159_b0 );
or ( \1161_b1 , \1160_b1 , w_2306 );
xor ( \1161_b0 , \1160_b0 , w_2308 );
not ( w_2308 , w_2309 );
and ( w_2309 , w_2306 , w_2307 );
buf ( w_2306 , \320_b1 );
not ( w_2306 , w_2310 );
not ( w_2307 , w_2311 );
and ( w_2310 , w_2311 , \320_b0 );
or ( \1162_b1 , \1157_b1 , \1161_b1 );
not ( \1161_b1 , w_2312 );
and ( \1162_b0 , \1157_b0 , w_2313 );
and ( w_2312 , w_2313 , \1161_b0 );
or ( \1163_b1 , \904_b1 , \331_b1 );
not ( \331_b1 , w_2314 );
and ( \1163_b0 , \904_b0 , w_2315 );
and ( w_2314 , w_2315 , \331_b0 );
or ( \1164_b1 , \841_b1 , \329_b1 );
not ( \329_b1 , w_2316 );
and ( \1164_b0 , \841_b0 , w_2317 );
and ( w_2316 , w_2317 , \329_b0 );
or ( \1165_b1 , \1163_b1 , w_2319 );
not ( w_2319 , w_2320 );
and ( \1165_b0 , \1163_b0 , w_2321 );
and ( w_2320 ,  , w_2321 );
buf ( w_2319 , \1164_b1 );
not ( w_2319 , w_2322 );
not (  , w_2323 );
and ( w_2322 , w_2323 , \1164_b0 );
or ( \1166_b1 , \1165_b1 , w_2324 );
xor ( \1166_b0 , \1165_b0 , w_2326 );
not ( w_2326 , w_2327 );
and ( w_2327 , w_2324 , w_2325 );
buf ( w_2324 , \338_b1 );
not ( w_2324 , w_2328 );
not ( w_2325 , w_2329 );
and ( w_2328 , w_2329 , \338_b0 );
or ( \1167_b1 , \1161_b1 , \1166_b1 );
not ( \1166_b1 , w_2330 );
and ( \1167_b0 , \1161_b0 , w_2331 );
and ( w_2330 , w_2331 , \1166_b0 );
or ( \1168_b1 , \1157_b1 , \1166_b1 );
not ( \1166_b1 , w_2332 );
and ( \1168_b0 , \1157_b0 , w_2333 );
and ( w_2332 , w_2333 , \1166_b0 );
or ( \1170_b1 , \1153_b1 , \1169_b1 );
not ( \1169_b1 , w_2334 );
and ( \1170_b0 , \1153_b0 , w_2335 );
and ( w_2334 , w_2335 , \1169_b0 );
and ( \1171_nR130_b1 , RIb4c3020_52_b1 , w_2336 );
xor ( w_2336 , RIb4c3020_52_b0 , \288_b1 );
not ( \288_b1 , w_2337 );
and ( \1171_nR130_b0 , w_2337 , \288_b0 );
buf ( \1172_b1 , \1171_nR130_b1 );
buf ( \1172_b0 , \1171_nR130_b0 );
and ( \1173_nR12f_b1 , RIb4c2fa8_53_b1 , w_2338 );
xor ( w_2338 , RIb4c2fa8_53_b0 , \288_b1 );
not ( \288_b1 , w_2339 );
and ( \1173_nR12f_b0 , w_2339 , \288_b0 );
buf ( \1174_b1 , \1173_nR12f_b1 );
buf ( \1174_b0 , \1173_nR12f_b0 );
or ( \1175_b1 , \1172_b1 , \1174_b1 );
not ( \1174_b1 , w_2340 );
and ( \1175_b0 , \1172_b0 , w_2341 );
and ( w_2340 , w_2341 , \1174_b0 );
buf ( \1176_b1 , \1175_b1 );
not ( \1176_b1 , w_2342 );
not ( \1176_b0 , w_2343 );
and ( w_2342 , w_2343 , \1175_b0 );
or ( \1177_b1 , \981_b1 , \1176_b1 );
not ( \1176_b1 , w_2344 );
and ( \1177_b0 , \981_b0 , w_2345 );
and ( w_2344 , w_2345 , \1176_b0 );
buf ( \1178_b1 , \1177_b1 );
not ( \1178_b1 , w_2346 );
not ( \1178_b0 , w_2347 );
and ( w_2346 , w_2347 , \1177_b0 );
or ( \1179_b1 , \315_b1 , \1062_b1 );
not ( \1062_b1 , w_2348 );
and ( \1179_b0 , \315_b0 , w_2349 );
and ( w_2348 , w_2349 , \1062_b0 );
or ( \1180_b1 , \159_b1 , \1060_b1 );
not ( \1060_b1 , w_2350 );
and ( \1180_b0 , \159_b0 , w_2351 );
and ( w_2350 , w_2351 , \1060_b0 );
or ( \1181_b1 , \1179_b1 , w_2353 );
not ( w_2353 , w_2354 );
and ( \1181_b0 , \1179_b0 , w_2355 );
and ( w_2354 ,  , w_2355 );
buf ( w_2353 , \1180_b1 );
not ( w_2353 , w_2356 );
not (  , w_2357 );
and ( w_2356 , w_2357 , \1180_b0 );
or ( \1182_b1 , \1181_b1 , w_2358 );
xor ( \1182_b0 , \1181_b0 , w_2360 );
not ( w_2360 , w_2361 );
and ( w_2361 , w_2358 , w_2359 );
buf ( w_2358 , \984_b1 );
not ( w_2358 , w_2362 );
not ( w_2359 , w_2363 );
and ( w_2362 , w_2363 , \984_b0 );
or ( \1183_b1 , \1178_b1 , \1182_b1 );
not ( \1182_b1 , w_2364 );
and ( \1183_b0 , \1178_b0 , w_2365 );
and ( w_2364 , w_2365 , \1182_b0 );
or ( \1184_b1 , \333_b1 , \912_b1 );
not ( \912_b1 , w_2366 );
and ( \1184_b0 , \333_b0 , w_2367 );
and ( w_2366 , w_2367 , \912_b0 );
or ( \1185_b1 , \305_b1 , \910_b1 );
not ( \910_b1 , w_2368 );
and ( \1185_b0 , \305_b0 , w_2369 );
and ( w_2368 , w_2369 , \910_b0 );
or ( \1186_b1 , \1184_b1 , w_2371 );
not ( w_2371 , w_2372 );
and ( \1186_b0 , \1184_b0 , w_2373 );
and ( w_2372 ,  , w_2373 );
buf ( w_2371 , \1185_b1 );
not ( w_2371 , w_2374 );
not (  , w_2375 );
and ( w_2374 , w_2375 , \1185_b0 );
or ( \1187_b1 , \1186_b1 , w_2376 );
xor ( \1187_b0 , \1186_b0 , w_2378 );
not ( w_2378 , w_2379 );
and ( w_2379 , w_2376 , w_2377 );
buf ( w_2376 , \818_b1 );
not ( w_2376 , w_2380 );
not ( w_2377 , w_2381 );
and ( w_2380 , w_2381 , \818_b0 );
or ( \1188_b1 , \1182_b1 , \1187_b1 );
not ( \1187_b1 , w_2382 );
and ( \1188_b0 , \1182_b0 , w_2383 );
and ( w_2382 , w_2383 , \1187_b0 );
or ( \1189_b1 , \1178_b1 , \1187_b1 );
not ( \1187_b1 , w_2384 );
and ( \1189_b0 , \1178_b0 , w_2385 );
and ( w_2384 , w_2385 , \1187_b0 );
or ( \1191_b1 , \1169_b1 , \1190_b1 );
not ( \1190_b1 , w_2386 );
and ( \1191_b0 , \1169_b0 , w_2387 );
and ( w_2386 , w_2387 , \1190_b0 );
or ( \1192_b1 , \1153_b1 , \1190_b1 );
not ( \1190_b1 , w_2388 );
and ( \1192_b0 , \1153_b0 , w_2389 );
and ( w_2388 , w_2389 , \1190_b0 );
buf ( \1194_b1 , RIb4bf240_82_b1 );
buf ( \1194_b0 , RIb4bf240_82_b0 );
or ( \1195_b1 , \1194_b1 , \345_b1 );
not ( \345_b1 , w_2390 );
and ( \1195_b0 , \1194_b0 , w_2391 );
and ( w_2390 , w_2391 , \345_b0 );
or ( \1196_b1 , \1098_b1 , \1102_b1 );
xor ( \1196_b0 , \1098_b0 , w_2392 );
not ( w_2392 , w_2393 );
and ( w_2393 , \1102_b1 , \1102_b0 );
or ( \1197_b1 , \1196_b1 , \1108_b1 );
xor ( \1197_b0 , \1196_b0 , w_2394 );
not ( w_2394 , w_2395 );
and ( w_2395 , \1108_b1 , \1108_b0 );
or ( \1198_b1 , \1195_b1 , w_2396 );
or ( \1198_b0 , \1195_b0 , \1197_b0 );
not ( \1197_b0 , w_2397 );
and ( w_2397 , w_2396 , \1197_b1 );
or ( \1199_b1 , \1193_b1 , \1198_b1 );
not ( \1198_b1 , w_2398 );
and ( \1199_b0 , \1193_b0 , w_2399 );
and ( w_2398 , w_2399 , \1198_b0 );
or ( \1200_b1 , \1065_b1 , \1069_b1 );
xor ( \1200_b0 , \1065_b0 , w_2400 );
not ( w_2400 , w_2401 );
and ( w_2401 , \1069_b1 , \1069_b0 );
or ( \1201_b1 , \1200_b1 , \1074_b1 );
xor ( \1201_b0 , \1200_b0 , w_2402 );
not ( w_2402 , w_2403 );
and ( w_2403 , \1074_b1 , \1074_b0 );
or ( \1202_b1 , \1081_b1 , \1085_b1 );
xor ( \1202_b0 , \1081_b0 , w_2404 );
not ( w_2404 , w_2405 );
and ( w_2405 , \1085_b1 , \1085_b0 );
or ( \1203_b1 , \1202_b1 , \1090_b1 );
xor ( \1203_b0 , \1202_b0 , w_2406 );
not ( w_2406 , w_2407 );
and ( w_2407 , \1090_b1 , \1090_b0 );
or ( \1204_b1 , \1201_b1 , \1203_b1 );
not ( \1203_b1 , w_2408 );
and ( \1204_b0 , \1201_b0 , w_2409 );
and ( w_2408 , w_2409 , \1203_b0 );
or ( \1205_b1 , \1198_b1 , \1204_b1 );
not ( \1204_b1 , w_2410 );
and ( \1205_b0 , \1198_b0 , w_2411 );
and ( w_2410 , w_2411 , \1204_b0 );
or ( \1206_b1 , \1193_b1 , \1204_b1 );
not ( \1204_b1 , w_2412 );
and ( \1206_b0 , \1193_b0 , w_2413 );
and ( w_2412 , w_2413 , \1204_b0 );
or ( \1208_b1 , \985_b1 , \989_b1 );
xor ( \1208_b0 , \985_b0 , w_2414 );
not ( w_2414 , w_2415 );
and ( w_2415 , \989_b1 , \989_b0 );
or ( \1209_b1 , \1208_b1 , \994_b1 );
xor ( \1209_b0 , \1208_b0 , w_2416 );
not ( w_2416 , w_2417 );
and ( w_2417 , \994_b1 , \994_b0 );
or ( \1210_b1 , \1077_b1 , \1093_b1 );
xor ( \1210_b0 , \1077_b0 , w_2418 );
not ( w_2418 , w_2419 );
and ( w_2419 , \1093_b1 , \1093_b0 );
or ( \1211_b1 , \1210_b1 , \1111_b1 );
xor ( \1211_b0 , \1210_b0 , w_2420 );
not ( w_2420 , w_2421 );
and ( w_2421 , \1111_b1 , \1111_b0 );
or ( \1212_b1 , \1209_b1 , \1211_b1 );
not ( \1211_b1 , w_2422 );
and ( \1212_b0 , \1209_b0 , w_2423 );
and ( w_2422 , w_2423 , \1211_b0 );
or ( \1213_b1 , \1115_b1 , \1117_b1 );
xor ( \1213_b0 , \1115_b0 , w_2424 );
not ( w_2424 , w_2425 );
and ( w_2425 , \1117_b1 , \1117_b0 );
or ( \1214_b1 , \1213_b1 , \1120_b1 );
xor ( \1214_b0 , \1213_b0 , w_2426 );
not ( w_2426 , w_2427 );
and ( w_2427 , \1120_b1 , \1120_b0 );
or ( \1215_b1 , \1211_b1 , \1214_b1 );
not ( \1214_b1 , w_2428 );
and ( \1215_b0 , \1211_b0 , w_2429 );
and ( w_2428 , w_2429 , \1214_b0 );
or ( \1216_b1 , \1209_b1 , \1214_b1 );
not ( \1214_b1 , w_2430 );
and ( \1216_b0 , \1209_b0 , w_2431 );
and ( w_2430 , w_2431 , \1214_b0 );
or ( \1218_b1 , \1207_b1 , \1217_b1 );
not ( \1217_b1 , w_2432 );
and ( \1218_b0 , \1207_b0 , w_2433 );
and ( w_2432 , w_2433 , \1217_b0 );
or ( \1219_b1 , \1035_b1 , w_2434 );
xor ( \1219_b0 , \1035_b0 , w_2436 );
not ( w_2436 , w_2437 );
and ( w_2437 , w_2434 , w_2435 );
buf ( w_2434 , \1037_b1 );
not ( w_2434 , w_2438 );
not ( w_2435 , w_2439 );
and ( w_2438 , w_2439 , \1037_b0 );
or ( \1220_b1 , \1217_b1 , \1219_b1 );
not ( \1219_b1 , w_2440 );
and ( \1220_b0 , \1217_b0 , w_2441 );
and ( w_2440 , w_2441 , \1219_b0 );
or ( \1221_b1 , \1207_b1 , \1219_b1 );
not ( \1219_b1 , w_2442 );
and ( \1221_b0 , \1207_b0 , w_2443 );
and ( w_2442 , w_2443 , \1219_b0 );
or ( \1223_b1 , \997_b1 , \1013_b1 );
xor ( \1223_b0 , \997_b0 , w_2444 );
not ( w_2444 , w_2445 );
and ( w_2445 , \1013_b1 , \1013_b0 );
or ( \1224_b1 , \1223_b1 , \1030_b1 );
xor ( \1224_b0 , \1223_b0 , w_2446 );
not ( w_2446 , w_2447 );
and ( w_2447 , \1030_b1 , \1030_b0 );
or ( \1225_b1 , \1114_b1 , \1123_b1 );
xor ( \1225_b0 , \1114_b0 , w_2448 );
not ( w_2448 , w_2449 );
and ( w_2449 , \1123_b1 , \1123_b0 );
or ( \1226_b1 , \1225_b1 , \1126_b1 );
xor ( \1226_b0 , \1225_b0 , w_2450 );
not ( w_2450 , w_2451 );
and ( w_2451 , \1126_b1 , \1126_b0 );
or ( \1227_b1 , \1224_b1 , \1226_b1 );
not ( \1226_b1 , w_2452 );
and ( \1227_b0 , \1224_b0 , w_2453 );
and ( w_2452 , w_2453 , \1226_b0 );
or ( \1228_b1 , \1222_b1 , \1227_b1 );
not ( \1227_b1 , w_2454 );
and ( \1228_b0 , \1222_b0 , w_2455 );
and ( w_2454 , w_2455 , \1227_b0 );
or ( \1229_b1 , \1129_b1 , \1131_b1 );
xor ( \1229_b0 , \1129_b0 , w_2456 );
not ( w_2456 , w_2457 );
and ( w_2457 , \1131_b1 , \1131_b0 );
or ( \1230_b1 , \1229_b1 , \1134_b1 );
xor ( \1230_b0 , \1229_b0 , w_2458 );
not ( w_2458 , w_2459 );
and ( w_2459 , \1134_b1 , \1134_b0 );
or ( \1231_b1 , \1227_b1 , \1230_b1 );
not ( \1230_b1 , w_2460 );
and ( \1231_b0 , \1227_b0 , w_2461 );
and ( w_2460 , w_2461 , \1230_b0 );
or ( \1232_b1 , \1222_b1 , \1230_b1 );
not ( \1230_b1 , w_2462 );
and ( \1232_b0 , \1222_b0 , w_2463 );
and ( w_2462 , w_2463 , \1230_b0 );
or ( \1234_b1 , \1137_b1 , \1233_b1 );
not ( \1233_b1 , w_2464 );
and ( \1234_b0 , \1137_b0 , w_2465 );
and ( w_2464 , w_2465 , \1233_b0 );
or ( \1235_b1 , \1044_b1 , \1046_b1 );
xor ( \1235_b0 , \1044_b0 , w_2466 );
not ( w_2466 , w_2467 );
and ( w_2467 , \1046_b1 , \1046_b0 );
or ( \1236_b1 , \1235_b1 , \1049_b1 );
xor ( \1236_b0 , \1235_b0 , w_2468 );
not ( w_2468 , w_2469 );
and ( w_2469 , \1049_b1 , \1049_b0 );
or ( \1237_b1 , \1233_b1 , \1236_b1 );
not ( \1236_b1 , w_2470 );
and ( \1237_b0 , \1233_b0 , w_2471 );
and ( w_2470 , w_2471 , \1236_b0 );
or ( \1238_b1 , \1137_b1 , \1236_b1 );
not ( \1236_b1 , w_2472 );
and ( \1238_b0 , \1137_b0 , w_2473 );
and ( w_2472 , w_2473 , \1236_b0 );
or ( \1240_b1 , \1058_b1 , \1239_b1 );
not ( \1239_b1 , w_2474 );
and ( \1240_b0 , \1058_b0 , w_2475 );
and ( w_2474 , w_2475 , \1239_b0 );
or ( \1241_b1 , \1058_b1 , \1239_b1 );
xor ( \1241_b0 , \1058_b0 , w_2476 );
not ( w_2476 , w_2477 );
and ( w_2477 , \1239_b1 , \1239_b0 );
or ( \1242_b1 , \1137_b1 , \1233_b1 );
xor ( \1242_b0 , \1137_b0 , w_2478 );
not ( w_2478 , w_2479 );
and ( w_2479 , \1233_b1 , \1233_b0 );
or ( \1243_b1 , \1242_b1 , \1236_b1 );
xor ( \1243_b0 , \1242_b0 , w_2480 );
not ( w_2480 , w_2481 );
and ( w_2481 , \1236_b1 , \1236_b0 );
or ( \1244_b1 , \343_b1 , \740_b1 );
not ( \740_b1 , w_2482 );
and ( \1244_b0 , \343_b0 , w_2483 );
and ( w_2482 , w_2483 , \740_b0 );
or ( \1245_b1 , \353_b1 , \738_b1 );
not ( \738_b1 , w_2484 );
and ( \1245_b0 , \353_b0 , w_2485 );
and ( w_2484 , w_2485 , \738_b0 );
or ( \1246_b1 , \1244_b1 , w_2487 );
not ( w_2487 , w_2488 );
and ( \1246_b0 , \1244_b0 , w_2489 );
and ( w_2488 ,  , w_2489 );
buf ( w_2487 , \1245_b1 );
not ( w_2487 , w_2490 );
not (  , w_2491 );
and ( w_2490 , w_2491 , \1245_b0 );
or ( \1247_b1 , \1246_b1 , w_2492 );
xor ( \1247_b0 , \1246_b0 , w_2494 );
not ( w_2494 , w_2495 );
and ( w_2495 , w_2492 , w_2493 );
buf ( w_2492 , \668_b1 );
not ( w_2492 , w_2496 );
not ( w_2493 , w_2497 );
and ( w_2496 , w_2497 , \668_b0 );
or ( \1248_b1 , \444_b1 , \604_b1 );
not ( \604_b1 , w_2498 );
and ( \1248_b0 , \444_b0 , w_2499 );
and ( w_2498 , w_2499 , \604_b0 );
or ( \1249_b1 , \360_b1 , \602_b1 );
not ( \602_b1 , w_2500 );
and ( \1249_b0 , \360_b0 , w_2501 );
and ( w_2500 , w_2501 , \602_b0 );
or ( \1250_b1 , \1248_b1 , w_2503 );
not ( w_2503 , w_2504 );
and ( \1250_b0 , \1248_b0 , w_2505 );
and ( w_2504 ,  , w_2505 );
buf ( w_2503 , \1249_b1 );
not ( w_2503 , w_2506 );
not (  , w_2507 );
and ( w_2506 , w_2507 , \1249_b0 );
or ( \1251_b1 , \1250_b1 , w_2508 );
xor ( \1251_b0 , \1250_b0 , w_2510 );
not ( w_2510 , w_2511 );
and ( w_2511 , w_2508 , w_2509 );
buf ( w_2508 , \561_b1 );
not ( w_2508 , w_2512 );
not ( w_2509 , w_2513 );
and ( w_2512 , w_2513 , \561_b0 );
or ( \1252_b1 , \1247_b1 , \1251_b1 );
not ( \1251_b1 , w_2514 );
and ( \1252_b0 , \1247_b0 , w_2515 );
and ( w_2514 , w_2515 , \1251_b0 );
or ( \1253_b1 , \593_b1 , \503_b1 );
not ( \503_b1 , w_2516 );
and ( \1253_b0 , \593_b0 , w_2517 );
and ( w_2516 , w_2517 , \503_b0 );
or ( \1254_b1 , \495_b1 , \501_b1 );
not ( \501_b1 , w_2518 );
and ( \1254_b0 , \495_b0 , w_2519 );
and ( w_2518 , w_2519 , \501_b0 );
or ( \1255_b1 , \1253_b1 , w_2521 );
not ( w_2521 , w_2522 );
and ( \1255_b0 , \1253_b0 , w_2523 );
and ( w_2522 ,  , w_2523 );
buf ( w_2521 , \1254_b1 );
not ( w_2521 , w_2524 );
not (  , w_2525 );
and ( w_2524 , w_2525 , \1254_b0 );
or ( \1256_b1 , \1255_b1 , w_2526 );
xor ( \1256_b0 , \1255_b0 , w_2528 );
not ( w_2528 , w_2529 );
and ( w_2529 , w_2526 , w_2527 );
buf ( w_2526 , \455_b1 );
not ( w_2526 , w_2530 );
not ( w_2527 , w_2531 );
and ( w_2530 , w_2531 , \455_b0 );
or ( \1257_b1 , \1251_b1 , \1256_b1 );
not ( \1256_b1 , w_2532 );
and ( \1257_b0 , \1251_b0 , w_2533 );
and ( w_2532 , w_2533 , \1256_b0 );
or ( \1258_b1 , \1247_b1 , \1256_b1 );
not ( \1256_b1 , w_2534 );
and ( \1258_b0 , \1247_b0 , w_2535 );
and ( w_2534 , w_2535 , \1256_b0 );
or ( \1260_b1 , \703_b1 , \298_b1 );
not ( \298_b1 , w_2536 );
and ( \1260_b0 , \703_b0 , w_2537 );
and ( w_2536 , w_2537 , \298_b0 );
or ( \1261_b1 , \621_b1 , \296_b1 );
not ( \296_b1 , w_2538 );
and ( \1261_b0 , \621_b0 , w_2539 );
and ( w_2538 , w_2539 , \296_b0 );
or ( \1262_b1 , \1260_b1 , w_2541 );
not ( w_2541 , w_2542 );
and ( \1262_b0 , \1260_b0 , w_2543 );
and ( w_2542 ,  , w_2543 );
buf ( w_2541 , \1261_b1 );
not ( w_2541 , w_2544 );
not (  , w_2545 );
and ( w_2544 , w_2545 , \1261_b0 );
or ( \1263_b1 , \1262_b1 , w_2546 );
xor ( \1263_b0 , \1262_b0 , w_2548 );
not ( w_2548 , w_2549 );
and ( w_2549 , w_2546 , w_2547 );
buf ( w_2546 , \303_b1 );
not ( w_2546 , w_2550 );
not ( w_2547 , w_2551 );
and ( w_2550 , w_2551 , \303_b0 );
or ( \1264_b1 , \841_b1 , \313_b1 );
not ( \313_b1 , w_2552 );
and ( \1264_b0 , \841_b0 , w_2553 );
and ( w_2552 , w_2553 , \313_b0 );
or ( \1265_b1 , \777_b1 , \311_b1 );
not ( \311_b1 , w_2554 );
and ( \1265_b0 , \777_b0 , w_2555 );
and ( w_2554 , w_2555 , \311_b0 );
or ( \1266_b1 , \1264_b1 , w_2557 );
not ( w_2557 , w_2558 );
and ( \1266_b0 , \1264_b0 , w_2559 );
and ( w_2558 ,  , w_2559 );
buf ( w_2557 , \1265_b1 );
not ( w_2557 , w_2560 );
not (  , w_2561 );
and ( w_2560 , w_2561 , \1265_b0 );
or ( \1267_b1 , \1266_b1 , w_2562 );
xor ( \1267_b0 , \1266_b0 , w_2564 );
not ( w_2564 , w_2565 );
and ( w_2565 , w_2562 , w_2563 );
buf ( w_2562 , \320_b1 );
not ( w_2562 , w_2566 );
not ( w_2563 , w_2567 );
and ( w_2566 , w_2567 , \320_b0 );
or ( \1268_b1 , \1263_b1 , \1267_b1 );
not ( \1267_b1 , w_2568 );
and ( \1268_b0 , \1263_b0 , w_2569 );
and ( w_2568 , w_2569 , \1267_b0 );
or ( \1269_b1 , \1104_b1 , \331_b1 );
not ( \331_b1 , w_2570 );
and ( \1269_b0 , \1104_b0 , w_2571 );
and ( w_2570 , w_2571 , \331_b0 );
or ( \1270_b1 , \904_b1 , \329_b1 );
not ( \329_b1 , w_2572 );
and ( \1270_b0 , \904_b0 , w_2573 );
and ( w_2572 , w_2573 , \329_b0 );
or ( \1271_b1 , \1269_b1 , w_2575 );
not ( w_2575 , w_2576 );
and ( \1271_b0 , \1269_b0 , w_2577 );
and ( w_2576 ,  , w_2577 );
buf ( w_2575 , \1270_b1 );
not ( w_2575 , w_2578 );
not (  , w_2579 );
and ( w_2578 , w_2579 , \1270_b0 );
or ( \1272_b1 , \1271_b1 , w_2580 );
xor ( \1272_b0 , \1271_b0 , w_2582 );
not ( w_2582 , w_2583 );
and ( w_2583 , w_2580 , w_2581 );
buf ( w_2580 , \338_b1 );
not ( w_2580 , w_2584 );
not ( w_2581 , w_2585 );
and ( w_2584 , w_2585 , \338_b0 );
or ( \1273_b1 , \1267_b1 , \1272_b1 );
not ( \1272_b1 , w_2586 );
and ( \1273_b0 , \1267_b0 , w_2587 );
and ( w_2586 , w_2587 , \1272_b0 );
or ( \1274_b1 , \1263_b1 , \1272_b1 );
not ( \1272_b1 , w_2588 );
and ( \1274_b0 , \1263_b0 , w_2589 );
and ( w_2588 , w_2589 , \1272_b0 );
or ( \1276_b1 , \1259_b1 , \1275_b1 );
not ( \1275_b1 , w_2590 );
and ( \1276_b0 , \1259_b0 , w_2591 );
and ( w_2590 , w_2591 , \1275_b0 );
or ( \1277_b1 , \981_b1 , \1172_b1 );
xor ( \1277_b0 , \981_b0 , w_2592 );
not ( w_2592 , w_2593 );
and ( w_2593 , \1172_b1 , \1172_b0 );
or ( \1278_b1 , \1172_b1 , \1174_b1 );
xor ( \1278_b0 , \1172_b0 , w_2594 );
not ( w_2594 , w_2595 );
and ( w_2595 , \1174_b1 , \1174_b0 );
buf ( \1279_b1 , \1278_b1 );
not ( \1279_b1 , w_2596 );
not ( \1279_b0 , w_2597 );
and ( w_2596 , w_2597 , \1278_b0 );
or ( \1280_b1 , \1277_b1 , \1279_b1 );
not ( \1279_b1 , w_2598 );
and ( \1280_b0 , \1277_b0 , w_2599 );
and ( w_2598 , w_2599 , \1279_b0 );
or ( \1281_b1 , \159_b1 , \1280_b1 );
not ( \1280_b1 , w_2600 );
and ( \1281_b0 , \159_b0 , w_2601 );
and ( w_2600 , w_2601 , \1280_b0 );
buf ( \1282_b1 , \1281_b1 );
not ( \1282_b1 , w_2602 );
not ( \1282_b0 , w_2603 );
and ( w_2602 , w_2603 , \1281_b0 );
or ( \1283_b1 , \1282_b1 , w_2604 );
xor ( \1283_b0 , \1282_b0 , w_2606 );
not ( w_2606 , w_2607 );
and ( w_2607 , w_2604 , w_2605 );
buf ( w_2604 , \1177_b1 );
not ( w_2604 , w_2608 );
not ( w_2605 , w_2609 );
and ( w_2608 , w_2609 , \1177_b0 );
or ( \1284_b1 , \305_b1 , \1062_b1 );
not ( \1062_b1 , w_2610 );
and ( \1284_b0 , \305_b0 , w_2611 );
and ( w_2610 , w_2611 , \1062_b0 );
or ( \1285_b1 , \315_b1 , \1060_b1 );
not ( \1060_b1 , w_2612 );
and ( \1285_b0 , \315_b0 , w_2613 );
and ( w_2612 , w_2613 , \1060_b0 );
or ( \1286_b1 , \1284_b1 , w_2615 );
not ( w_2615 , w_2616 );
and ( \1286_b0 , \1284_b0 , w_2617 );
and ( w_2616 ,  , w_2617 );
buf ( w_2615 , \1285_b1 );
not ( w_2615 , w_2618 );
not (  , w_2619 );
and ( w_2618 , w_2619 , \1285_b0 );
or ( \1287_b1 , \1286_b1 , w_2620 );
xor ( \1287_b0 , \1286_b0 , w_2622 );
not ( w_2622 , w_2623 );
and ( w_2623 , w_2620 , w_2621 );
buf ( w_2620 , \984_b1 );
not ( w_2620 , w_2624 );
not ( w_2621 , w_2625 );
and ( w_2624 , w_2625 , \984_b0 );
or ( \1288_b1 , \1283_b1 , \1287_b1 );
not ( \1287_b1 , w_2626 );
and ( \1288_b0 , \1283_b0 , w_2627 );
and ( w_2626 , w_2627 , \1287_b0 );
or ( \1289_b1 , \323_b1 , \912_b1 );
not ( \912_b1 , w_2628 );
and ( \1289_b0 , \323_b0 , w_2629 );
and ( w_2628 , w_2629 , \912_b0 );
or ( \1290_b1 , \333_b1 , \910_b1 );
not ( \910_b1 , w_2630 );
and ( \1290_b0 , \333_b0 , w_2631 );
and ( w_2630 , w_2631 , \910_b0 );
or ( \1291_b1 , \1289_b1 , w_2633 );
not ( w_2633 , w_2634 );
and ( \1291_b0 , \1289_b0 , w_2635 );
and ( w_2634 ,  , w_2635 );
buf ( w_2633 , \1290_b1 );
not ( w_2633 , w_2636 );
not (  , w_2637 );
and ( w_2636 , w_2637 , \1290_b0 );
or ( \1292_b1 , \1291_b1 , w_2638 );
xor ( \1292_b0 , \1291_b0 , w_2640 );
not ( w_2640 , w_2641 );
and ( w_2641 , w_2638 , w_2639 );
buf ( w_2638 , \818_b1 );
not ( w_2638 , w_2642 );
not ( w_2639 , w_2643 );
and ( w_2642 , w_2643 , \818_b0 );
or ( \1293_b1 , \1287_b1 , \1292_b1 );
not ( \1292_b1 , w_2644 );
and ( \1293_b0 , \1287_b0 , w_2645 );
and ( w_2644 , w_2645 , \1292_b0 );
or ( \1294_b1 , \1283_b1 , \1292_b1 );
not ( \1292_b1 , w_2646 );
and ( \1294_b0 , \1283_b0 , w_2647 );
and ( w_2646 , w_2647 , \1292_b0 );
or ( \1296_b1 , \1275_b1 , \1295_b1 );
not ( \1295_b1 , w_2648 );
and ( \1296_b0 , \1275_b0 , w_2649 );
and ( w_2648 , w_2649 , \1295_b0 );
or ( \1297_b1 , \1259_b1 , \1295_b1 );
not ( \1295_b1 , w_2650 );
and ( \1297_b0 , \1259_b0 , w_2651 );
and ( w_2650 , w_2651 , \1295_b0 );
buf ( \1299_b1 , RIb4bf1c8_83_b1 );
buf ( \1299_b0 , RIb4bf1c8_83_b0 );
or ( \1300_b1 , \1299_b1 , \351_b1 );
not ( \351_b1 , w_2652 );
and ( \1300_b0 , \1299_b0 , w_2653 );
and ( w_2652 , w_2653 , \351_b0 );
or ( \1301_b1 , \1194_b1 , \349_b1 );
not ( \349_b1 , w_2654 );
and ( \1301_b0 , \1194_b0 , w_2655 );
and ( w_2654 , w_2655 , \349_b0 );
or ( \1302_b1 , \1300_b1 , w_2657 );
not ( w_2657 , w_2658 );
and ( \1302_b0 , \1300_b0 , w_2659 );
and ( w_2658 ,  , w_2659 );
buf ( w_2657 , \1301_b1 );
not ( w_2657 , w_2660 );
not (  , w_2661 );
and ( w_2660 , w_2661 , \1301_b0 );
or ( \1303_b1 , \1302_b1 , w_2662 );
xor ( \1303_b0 , \1302_b0 , w_2664 );
not ( w_2664 , w_2665 );
and ( w_2665 , w_2662 , w_2663 );
buf ( w_2662 , \358_b1 );
not ( w_2662 , w_2666 );
not ( w_2663 , w_2667 );
and ( w_2666 , w_2667 , \358_b0 );
buf ( \1304_b1 , RIb4bf150_84_b1 );
buf ( \1304_b0 , RIb4bf150_84_b0 );
or ( \1305_b1 , \1304_b1 , \345_b1 );
not ( \345_b1 , w_2668 );
and ( \1305_b0 , \1304_b0 , w_2669 );
and ( w_2668 , w_2669 , \345_b0 );
or ( \1306_b1 , \1303_b1 , w_2670 );
or ( \1306_b0 , \1303_b0 , \1305_b0 );
not ( \1305_b0 , w_2671 );
and ( w_2671 , w_2670 , \1305_b1 );
or ( \1307_b1 , \1194_b1 , \351_b1 );
not ( \351_b1 , w_2672 );
and ( \1307_b0 , \1194_b0 , w_2673 );
and ( w_2672 , w_2673 , \351_b0 );
or ( \1308_b1 , \1104_b1 , \349_b1 );
not ( \349_b1 , w_2674 );
and ( \1308_b0 , \1104_b0 , w_2675 );
and ( w_2674 , w_2675 , \349_b0 );
or ( \1309_b1 , \1307_b1 , w_2677 );
not ( w_2677 , w_2678 );
and ( \1309_b0 , \1307_b0 , w_2679 );
and ( w_2678 ,  , w_2679 );
buf ( w_2677 , \1308_b1 );
not ( w_2677 , w_2680 );
not (  , w_2681 );
and ( w_2680 , w_2681 , \1308_b0 );
or ( \1310_b1 , \1309_b1 , w_2682 );
xor ( \1310_b0 , \1309_b0 , w_2684 );
not ( w_2684 , w_2685 );
and ( w_2685 , w_2682 , w_2683 );
buf ( w_2682 , \358_b1 );
not ( w_2682 , w_2686 );
not ( w_2683 , w_2687 );
and ( w_2686 , w_2687 , \358_b0 );
or ( \1311_b1 , \1306_b1 , \1310_b1 );
not ( \1310_b1 , w_2688 );
and ( \1311_b0 , \1306_b0 , w_2689 );
and ( w_2688 , w_2689 , \1310_b0 );
or ( \1312_b1 , \1299_b1 , \345_b1 );
not ( \345_b1 , w_2690 );
and ( \1312_b0 , \1299_b0 , w_2691 );
and ( w_2690 , w_2691 , \345_b0 );
or ( \1313_b1 , \1310_b1 , \1312_b1 );
not ( \1312_b1 , w_2692 );
and ( \1313_b0 , \1310_b0 , w_2693 );
and ( w_2692 , w_2693 , \1312_b0 );
or ( \1314_b1 , \1306_b1 , \1312_b1 );
not ( \1312_b1 , w_2694 );
and ( \1314_b0 , \1306_b0 , w_2695 );
and ( w_2694 , w_2695 , \1312_b0 );
or ( \1316_b1 , \1298_b1 , \1315_b1 );
not ( \1315_b1 , w_2696 );
and ( \1316_b0 , \1298_b0 , w_2697 );
and ( w_2696 , w_2697 , \1315_b0 );
or ( \1317_b1 , \1141_b1 , \1145_b1 );
xor ( \1317_b0 , \1141_b0 , w_2698 );
not ( w_2698 , w_2699 );
and ( w_2699 , \1145_b1 , \1145_b0 );
or ( \1318_b1 , \1317_b1 , \1150_b1 );
xor ( \1318_b0 , \1317_b0 , w_2700 );
not ( w_2700 , w_2701 );
and ( w_2701 , \1150_b1 , \1150_b0 );
or ( \1319_b1 , \1157_b1 , \1161_b1 );
xor ( \1319_b0 , \1157_b0 , w_2702 );
not ( w_2702 , w_2703 );
and ( w_2703 , \1161_b1 , \1161_b0 );
or ( \1320_b1 , \1319_b1 , \1166_b1 );
xor ( \1320_b0 , \1319_b0 , w_2704 );
not ( w_2704 , w_2705 );
and ( w_2705 , \1166_b1 , \1166_b0 );
or ( \1321_b1 , \1318_b1 , \1320_b1 );
not ( \1320_b1 , w_2706 );
and ( \1321_b0 , \1318_b0 , w_2707 );
and ( w_2706 , w_2707 , \1320_b0 );
or ( \1322_b1 , \1178_b1 , \1182_b1 );
xor ( \1322_b0 , \1178_b0 , w_2708 );
not ( w_2708 , w_2709 );
and ( w_2709 , \1182_b1 , \1182_b0 );
or ( \1323_b1 , \1322_b1 , \1187_b1 );
xor ( \1323_b0 , \1322_b0 , w_2710 );
not ( w_2710 , w_2711 );
and ( w_2711 , \1187_b1 , \1187_b0 );
or ( \1324_b1 , \1320_b1 , \1323_b1 );
not ( \1323_b1 , w_2712 );
and ( \1324_b0 , \1320_b0 , w_2713 );
and ( w_2712 , w_2713 , \1323_b0 );
or ( \1325_b1 , \1318_b1 , \1323_b1 );
not ( \1323_b1 , w_2714 );
and ( \1325_b0 , \1318_b0 , w_2715 );
and ( w_2714 , w_2715 , \1323_b0 );
or ( \1327_b1 , \1315_b1 , \1326_b1 );
not ( \1326_b1 , w_2716 );
and ( \1327_b0 , \1315_b0 , w_2717 );
and ( w_2716 , w_2717 , \1326_b0 );
or ( \1328_b1 , \1298_b1 , \1326_b1 );
not ( \1326_b1 , w_2718 );
and ( \1328_b0 , \1298_b0 , w_2719 );
and ( w_2718 , w_2719 , \1326_b0 );
or ( \1330_b1 , \1153_b1 , \1169_b1 );
xor ( \1330_b0 , \1153_b0 , w_2720 );
not ( w_2720 , w_2721 );
and ( w_2721 , \1169_b1 , \1169_b0 );
or ( \1331_b1 , \1330_b1 , \1190_b1 );
xor ( \1331_b0 , \1330_b0 , w_2722 );
not ( w_2722 , w_2723 );
and ( w_2723 , \1190_b1 , \1190_b0 );
or ( \1332_b1 , \1195_b1 , w_2724 );
xor ( \1332_b0 , \1195_b0 , w_2726 );
not ( w_2726 , w_2727 );
and ( w_2727 , w_2724 , w_2725 );
buf ( w_2724 , \1197_b1 );
not ( w_2724 , w_2728 );
not ( w_2725 , w_2729 );
and ( w_2728 , w_2729 , \1197_b0 );
or ( \1333_b1 , \1331_b1 , \1332_b1 );
not ( \1332_b1 , w_2730 );
and ( \1333_b0 , \1331_b0 , w_2731 );
and ( w_2730 , w_2731 , \1332_b0 );
or ( \1334_b1 , \1201_b1 , \1203_b1 );
xor ( \1334_b0 , \1201_b0 , w_2732 );
not ( w_2732 , w_2733 );
and ( w_2733 , \1203_b1 , \1203_b0 );
or ( \1335_b1 , \1332_b1 , \1334_b1 );
not ( \1334_b1 , w_2734 );
and ( \1335_b0 , \1332_b0 , w_2735 );
and ( w_2734 , w_2735 , \1334_b0 );
or ( \1336_b1 , \1331_b1 , \1334_b1 );
not ( \1334_b1 , w_2736 );
and ( \1336_b0 , \1331_b0 , w_2737 );
and ( w_2736 , w_2737 , \1334_b0 );
or ( \1338_b1 , \1329_b1 , \1337_b1 );
not ( \1337_b1 , w_2738 );
and ( \1338_b0 , \1329_b0 , w_2739 );
and ( w_2738 , w_2739 , \1337_b0 );
or ( \1339_b1 , \1209_b1 , \1211_b1 );
xor ( \1339_b0 , \1209_b0 , w_2740 );
not ( w_2740 , w_2741 );
and ( w_2741 , \1211_b1 , \1211_b0 );
or ( \1340_b1 , \1339_b1 , \1214_b1 );
xor ( \1340_b0 , \1339_b0 , w_2742 );
not ( w_2742 , w_2743 );
and ( w_2743 , \1214_b1 , \1214_b0 );
or ( \1341_b1 , \1337_b1 , \1340_b1 );
not ( \1340_b1 , w_2744 );
and ( \1341_b0 , \1337_b0 , w_2745 );
and ( w_2744 , w_2745 , \1340_b0 );
or ( \1342_b1 , \1329_b1 , \1340_b1 );
not ( \1340_b1 , w_2746 );
and ( \1342_b0 , \1329_b0 , w_2747 );
and ( w_2746 , w_2747 , \1340_b0 );
or ( \1344_b1 , \1207_b1 , \1217_b1 );
xor ( \1344_b0 , \1207_b0 , w_2748 );
not ( w_2748 , w_2749 );
and ( w_2749 , \1217_b1 , \1217_b0 );
or ( \1345_b1 , \1344_b1 , \1219_b1 );
xor ( \1345_b0 , \1344_b0 , w_2750 );
not ( w_2750 , w_2751 );
and ( w_2751 , \1219_b1 , \1219_b0 );
or ( \1346_b1 , \1343_b1 , \1345_b1 );
not ( \1345_b1 , w_2752 );
and ( \1346_b0 , \1343_b0 , w_2753 );
and ( w_2752 , w_2753 , \1345_b0 );
or ( \1347_b1 , \1224_b1 , \1226_b1 );
xor ( \1347_b0 , \1224_b0 , w_2754 );
not ( w_2754 , w_2755 );
and ( w_2755 , \1226_b1 , \1226_b0 );
or ( \1348_b1 , \1345_b1 , \1347_b1 );
not ( \1347_b1 , w_2756 );
and ( \1348_b0 , \1345_b0 , w_2757 );
and ( w_2756 , w_2757 , \1347_b0 );
or ( \1349_b1 , \1343_b1 , \1347_b1 );
not ( \1347_b1 , w_2758 );
and ( \1349_b0 , \1343_b0 , w_2759 );
and ( w_2758 , w_2759 , \1347_b0 );
or ( \1351_b1 , \1222_b1 , \1227_b1 );
xor ( \1351_b0 , \1222_b0 , w_2760 );
not ( w_2760 , w_2761 );
and ( w_2761 , \1227_b1 , \1227_b0 );
or ( \1352_b1 , \1351_b1 , \1230_b1 );
xor ( \1352_b0 , \1351_b0 , w_2762 );
not ( w_2762 , w_2763 );
and ( w_2763 , \1230_b1 , \1230_b0 );
or ( \1353_b1 , \1350_b1 , \1352_b1 );
not ( \1352_b1 , w_2764 );
and ( \1353_b0 , \1350_b0 , w_2765 );
and ( w_2764 , w_2765 , \1352_b0 );
or ( \1354_b1 , \1243_b1 , \1353_b1 );
not ( \1353_b1 , w_2766 );
and ( \1354_b0 , \1243_b0 , w_2767 );
and ( w_2766 , w_2767 , \1353_b0 );
or ( \1355_b1 , \1243_b1 , \1353_b1 );
xor ( \1355_b0 , \1243_b0 , w_2768 );
not ( w_2768 , w_2769 );
and ( w_2769 , \1353_b1 , \1353_b0 );
or ( \1356_b1 , \1350_b1 , \1352_b1 );
xor ( \1356_b0 , \1350_b0 , w_2770 );
not ( w_2770 , w_2771 );
and ( w_2771 , \1352_b1 , \1352_b0 );
and ( \1357_nR12e_b1 , RIb4c2f30_54_b1 , w_2772 );
xor ( w_2772 , RIb4c2f30_54_b0 , \288_b1 );
not ( \288_b1 , w_2773 );
and ( \1357_nR12e_b0 , w_2773 , \288_b0 );
buf ( \1358_b1 , \1357_nR12e_b1 );
buf ( \1358_b0 , \1357_nR12e_b0 );
and ( \1359_nR12d_b1 , RIb4c2eb8_55_b1 , w_2774 );
xor ( w_2774 , RIb4c2eb8_55_b0 , \288_b1 );
not ( \288_b1 , w_2775 );
and ( \1359_nR12d_b0 , w_2775 , \288_b0 );
buf ( \1360_b1 , \1359_nR12d_b1 );
buf ( \1360_b0 , \1359_nR12d_b0 );
or ( \1361_b1 , \1358_b1 , \1360_b1 );
not ( \1360_b1 , w_2776 );
and ( \1361_b0 , \1358_b0 , w_2777 );
and ( w_2776 , w_2777 , \1360_b0 );
buf ( \1362_b1 , \1361_b1 );
not ( \1362_b1 , w_2778 );
not ( \1362_b0 , w_2779 );
and ( w_2778 , w_2779 , \1361_b0 );
or ( \1363_b1 , \1174_b1 , \1362_b1 );
not ( \1362_b1 , w_2780 );
and ( \1363_b0 , \1174_b0 , w_2781 );
and ( w_2780 , w_2781 , \1362_b0 );
buf ( \1364_b1 , \1363_b1 );
not ( \1364_b1 , w_2782 );
not ( \1364_b0 , w_2783 );
and ( w_2782 , w_2783 , \1363_b0 );
or ( \1365_b1 , \315_b1 , \1280_b1 );
not ( \1280_b1 , w_2784 );
and ( \1365_b0 , \315_b0 , w_2785 );
and ( w_2784 , w_2785 , \1280_b0 );
or ( \1366_b1 , \159_b1 , \1278_b1 );
not ( \1278_b1 , w_2786 );
and ( \1366_b0 , \159_b0 , w_2787 );
and ( w_2786 , w_2787 , \1278_b0 );
or ( \1367_b1 , \1365_b1 , w_2789 );
not ( w_2789 , w_2790 );
and ( \1367_b0 , \1365_b0 , w_2791 );
and ( w_2790 ,  , w_2791 );
buf ( w_2789 , \1366_b1 );
not ( w_2789 , w_2792 );
not (  , w_2793 );
and ( w_2792 , w_2793 , \1366_b0 );
or ( \1368_b1 , \1367_b1 , w_2794 );
xor ( \1368_b0 , \1367_b0 , w_2796 );
not ( w_2796 , w_2797 );
and ( w_2797 , w_2794 , w_2795 );
buf ( w_2794 , \1177_b1 );
not ( w_2794 , w_2798 );
not ( w_2795 , w_2799 );
and ( w_2798 , w_2799 , \1177_b0 );
or ( \1369_b1 , \1364_b1 , \1368_b1 );
not ( \1368_b1 , w_2800 );
and ( \1369_b0 , \1364_b0 , w_2801 );
and ( w_2800 , w_2801 , \1368_b0 );
or ( \1370_b1 , \333_b1 , \1062_b1 );
not ( \1062_b1 , w_2802 );
and ( \1370_b0 , \333_b0 , w_2803 );
and ( w_2802 , w_2803 , \1062_b0 );
or ( \1371_b1 , \305_b1 , \1060_b1 );
not ( \1060_b1 , w_2804 );
and ( \1371_b0 , \305_b0 , w_2805 );
and ( w_2804 , w_2805 , \1060_b0 );
or ( \1372_b1 , \1370_b1 , w_2807 );
not ( w_2807 , w_2808 );
and ( \1372_b0 , \1370_b0 , w_2809 );
and ( w_2808 ,  , w_2809 );
buf ( w_2807 , \1371_b1 );
not ( w_2807 , w_2810 );
not (  , w_2811 );
and ( w_2810 , w_2811 , \1371_b0 );
or ( \1373_b1 , \1372_b1 , w_2812 );
xor ( \1373_b0 , \1372_b0 , w_2814 );
not ( w_2814 , w_2815 );
and ( w_2815 , w_2812 , w_2813 );
buf ( w_2812 , \984_b1 );
not ( w_2812 , w_2816 );
not ( w_2813 , w_2817 );
and ( w_2816 , w_2817 , \984_b0 );
or ( \1374_b1 , \1368_b1 , \1373_b1 );
not ( \1373_b1 , w_2818 );
and ( \1374_b0 , \1368_b0 , w_2819 );
and ( w_2818 , w_2819 , \1373_b0 );
or ( \1375_b1 , \1364_b1 , \1373_b1 );
not ( \1373_b1 , w_2820 );
and ( \1375_b0 , \1364_b0 , w_2821 );
and ( w_2820 , w_2821 , \1373_b0 );
or ( \1377_b1 , \353_b1 , \912_b1 );
not ( \912_b1 , w_2822 );
and ( \1377_b0 , \353_b0 , w_2823 );
and ( w_2822 , w_2823 , \912_b0 );
or ( \1378_b1 , \323_b1 , \910_b1 );
not ( \910_b1 , w_2824 );
and ( \1378_b0 , \323_b0 , w_2825 );
and ( w_2824 , w_2825 , \910_b0 );
or ( \1379_b1 , \1377_b1 , w_2827 );
not ( w_2827 , w_2828 );
and ( \1379_b0 , \1377_b0 , w_2829 );
and ( w_2828 ,  , w_2829 );
buf ( w_2827 , \1378_b1 );
not ( w_2827 , w_2830 );
not (  , w_2831 );
and ( w_2830 , w_2831 , \1378_b0 );
or ( \1380_b1 , \1379_b1 , w_2832 );
xor ( \1380_b0 , \1379_b0 , w_2834 );
not ( w_2834 , w_2835 );
and ( w_2835 , w_2832 , w_2833 );
buf ( w_2832 , \818_b1 );
not ( w_2832 , w_2836 );
not ( w_2833 , w_2837 );
and ( w_2836 , w_2837 , \818_b0 );
or ( \1381_b1 , \360_b1 , \740_b1 );
not ( \740_b1 , w_2838 );
and ( \1381_b0 , \360_b0 , w_2839 );
and ( w_2838 , w_2839 , \740_b0 );
or ( \1382_b1 , \343_b1 , \738_b1 );
not ( \738_b1 , w_2840 );
and ( \1382_b0 , \343_b0 , w_2841 );
and ( w_2840 , w_2841 , \738_b0 );
or ( \1383_b1 , \1381_b1 , w_2843 );
not ( w_2843 , w_2844 );
and ( \1383_b0 , \1381_b0 , w_2845 );
and ( w_2844 ,  , w_2845 );
buf ( w_2843 , \1382_b1 );
not ( w_2843 , w_2846 );
not (  , w_2847 );
and ( w_2846 , w_2847 , \1382_b0 );
or ( \1384_b1 , \1383_b1 , w_2848 );
xor ( \1384_b0 , \1383_b0 , w_2850 );
not ( w_2850 , w_2851 );
and ( w_2851 , w_2848 , w_2849 );
buf ( w_2848 , \668_b1 );
not ( w_2848 , w_2852 );
not ( w_2849 , w_2853 );
and ( w_2852 , w_2853 , \668_b0 );
or ( \1385_b1 , \1380_b1 , \1384_b1 );
not ( \1384_b1 , w_2854 );
and ( \1385_b0 , \1380_b0 , w_2855 );
and ( w_2854 , w_2855 , \1384_b0 );
or ( \1386_b1 , \495_b1 , \604_b1 );
not ( \604_b1 , w_2856 );
and ( \1386_b0 , \495_b0 , w_2857 );
and ( w_2856 , w_2857 , \604_b0 );
or ( \1387_b1 , \444_b1 , \602_b1 );
not ( \602_b1 , w_2858 );
and ( \1387_b0 , \444_b0 , w_2859 );
and ( w_2858 , w_2859 , \602_b0 );
or ( \1388_b1 , \1386_b1 , w_2861 );
not ( w_2861 , w_2862 );
and ( \1388_b0 , \1386_b0 , w_2863 );
and ( w_2862 ,  , w_2863 );
buf ( w_2861 , \1387_b1 );
not ( w_2861 , w_2864 );
not (  , w_2865 );
and ( w_2864 , w_2865 , \1387_b0 );
or ( \1389_b1 , \1388_b1 , w_2866 );
xor ( \1389_b0 , \1388_b0 , w_2868 );
not ( w_2868 , w_2869 );
and ( w_2869 , w_2866 , w_2867 );
buf ( w_2866 , \561_b1 );
not ( w_2866 , w_2870 );
not ( w_2867 , w_2871 );
and ( w_2870 , w_2871 , \561_b0 );
or ( \1390_b1 , \1384_b1 , \1389_b1 );
not ( \1389_b1 , w_2872 );
and ( \1390_b0 , \1384_b0 , w_2873 );
and ( w_2872 , w_2873 , \1389_b0 );
or ( \1391_b1 , \1380_b1 , \1389_b1 );
not ( \1389_b1 , w_2874 );
and ( \1391_b0 , \1380_b0 , w_2875 );
and ( w_2874 , w_2875 , \1389_b0 );
or ( \1393_b1 , \1376_b1 , \1392_b1 );
not ( \1392_b1 , w_2876 );
and ( \1393_b0 , \1376_b0 , w_2877 );
and ( w_2876 , w_2877 , \1392_b0 );
or ( \1394_b1 , \621_b1 , \503_b1 );
not ( \503_b1 , w_2878 );
and ( \1394_b0 , \621_b0 , w_2879 );
and ( w_2878 , w_2879 , \503_b0 );
or ( \1395_b1 , \593_b1 , \501_b1 );
not ( \501_b1 , w_2880 );
and ( \1395_b0 , \593_b0 , w_2881 );
and ( w_2880 , w_2881 , \501_b0 );
or ( \1396_b1 , \1394_b1 , w_2883 );
not ( w_2883 , w_2884 );
and ( \1396_b0 , \1394_b0 , w_2885 );
and ( w_2884 ,  , w_2885 );
buf ( w_2883 , \1395_b1 );
not ( w_2883 , w_2886 );
not (  , w_2887 );
and ( w_2886 , w_2887 , \1395_b0 );
or ( \1397_b1 , \1396_b1 , w_2888 );
xor ( \1397_b0 , \1396_b0 , w_2890 );
not ( w_2890 , w_2891 );
and ( w_2891 , w_2888 , w_2889 );
buf ( w_2888 , \455_b1 );
not ( w_2888 , w_2892 );
not ( w_2889 , w_2893 );
and ( w_2892 , w_2893 , \455_b0 );
or ( \1398_b1 , \777_b1 , \298_b1 );
not ( \298_b1 , w_2894 );
and ( \1398_b0 , \777_b0 , w_2895 );
and ( w_2894 , w_2895 , \298_b0 );
or ( \1399_b1 , \703_b1 , \296_b1 );
not ( \296_b1 , w_2896 );
and ( \1399_b0 , \703_b0 , w_2897 );
and ( w_2896 , w_2897 , \296_b0 );
or ( \1400_b1 , \1398_b1 , w_2899 );
not ( w_2899 , w_2900 );
and ( \1400_b0 , \1398_b0 , w_2901 );
and ( w_2900 ,  , w_2901 );
buf ( w_2899 , \1399_b1 );
not ( w_2899 , w_2902 );
not (  , w_2903 );
and ( w_2902 , w_2903 , \1399_b0 );
or ( \1401_b1 , \1400_b1 , w_2904 );
xor ( \1401_b0 , \1400_b0 , w_2906 );
not ( w_2906 , w_2907 );
and ( w_2907 , w_2904 , w_2905 );
buf ( w_2904 , \303_b1 );
not ( w_2904 , w_2908 );
not ( w_2905 , w_2909 );
and ( w_2908 , w_2909 , \303_b0 );
or ( \1402_b1 , \1397_b1 , \1401_b1 );
not ( \1401_b1 , w_2910 );
and ( \1402_b0 , \1397_b0 , w_2911 );
and ( w_2910 , w_2911 , \1401_b0 );
or ( \1403_b1 , \904_b1 , \313_b1 );
not ( \313_b1 , w_2912 );
and ( \1403_b0 , \904_b0 , w_2913 );
and ( w_2912 , w_2913 , \313_b0 );
or ( \1404_b1 , \841_b1 , \311_b1 );
not ( \311_b1 , w_2914 );
and ( \1404_b0 , \841_b0 , w_2915 );
and ( w_2914 , w_2915 , \311_b0 );
or ( \1405_b1 , \1403_b1 , w_2917 );
not ( w_2917 , w_2918 );
and ( \1405_b0 , \1403_b0 , w_2919 );
and ( w_2918 ,  , w_2919 );
buf ( w_2917 , \1404_b1 );
not ( w_2917 , w_2920 );
not (  , w_2921 );
and ( w_2920 , w_2921 , \1404_b0 );
or ( \1406_b1 , \1405_b1 , w_2922 );
xor ( \1406_b0 , \1405_b0 , w_2924 );
not ( w_2924 , w_2925 );
and ( w_2925 , w_2922 , w_2923 );
buf ( w_2922 , \320_b1 );
not ( w_2922 , w_2926 );
not ( w_2923 , w_2927 );
and ( w_2926 , w_2927 , \320_b0 );
or ( \1407_b1 , \1401_b1 , \1406_b1 );
not ( \1406_b1 , w_2928 );
and ( \1407_b0 , \1401_b0 , w_2929 );
and ( w_2928 , w_2929 , \1406_b0 );
or ( \1408_b1 , \1397_b1 , \1406_b1 );
not ( \1406_b1 , w_2930 );
and ( \1408_b0 , \1397_b0 , w_2931 );
and ( w_2930 , w_2931 , \1406_b0 );
or ( \1410_b1 , \1392_b1 , \1409_b1 );
not ( \1409_b1 , w_2932 );
and ( \1410_b0 , \1392_b0 , w_2933 );
and ( w_2932 , w_2933 , \1409_b0 );
or ( \1411_b1 , \1376_b1 , \1409_b1 );
not ( \1409_b1 , w_2934 );
and ( \1411_b0 , \1376_b0 , w_2935 );
and ( w_2934 , w_2935 , \1409_b0 );
or ( \1413_b1 , \1194_b1 , \331_b1 );
not ( \331_b1 , w_2936 );
and ( \1413_b0 , \1194_b0 , w_2937 );
and ( w_2936 , w_2937 , \331_b0 );
or ( \1414_b1 , \1104_b1 , \329_b1 );
not ( \329_b1 , w_2938 );
and ( \1414_b0 , \1104_b0 , w_2939 );
and ( w_2938 , w_2939 , \329_b0 );
or ( \1415_b1 , \1413_b1 , w_2941 );
not ( w_2941 , w_2942 );
and ( \1415_b0 , \1413_b0 , w_2943 );
and ( w_2942 ,  , w_2943 );
buf ( w_2941 , \1414_b1 );
not ( w_2941 , w_2944 );
not (  , w_2945 );
and ( w_2944 , w_2945 , \1414_b0 );
or ( \1416_b1 , \1415_b1 , w_2946 );
xor ( \1416_b0 , \1415_b0 , w_2948 );
not ( w_2948 , w_2949 );
and ( w_2949 , w_2946 , w_2947 );
buf ( w_2946 , \338_b1 );
not ( w_2946 , w_2950 );
not ( w_2947 , w_2951 );
and ( w_2950 , w_2951 , \338_b0 );
or ( \1417_b1 , \1304_b1 , \351_b1 );
not ( \351_b1 , w_2952 );
and ( \1417_b0 , \1304_b0 , w_2953 );
and ( w_2952 , w_2953 , \351_b0 );
or ( \1418_b1 , \1299_b1 , \349_b1 );
not ( \349_b1 , w_2954 );
and ( \1418_b0 , \1299_b0 , w_2955 );
and ( w_2954 , w_2955 , \349_b0 );
or ( \1419_b1 , \1417_b1 , w_2957 );
not ( w_2957 , w_2958 );
and ( \1419_b0 , \1417_b0 , w_2959 );
and ( w_2958 ,  , w_2959 );
buf ( w_2957 , \1418_b1 );
not ( w_2957 , w_2960 );
not (  , w_2961 );
and ( w_2960 , w_2961 , \1418_b0 );
or ( \1420_b1 , \1419_b1 , w_2962 );
xor ( \1420_b0 , \1419_b0 , w_2964 );
not ( w_2964 , w_2965 );
and ( w_2965 , w_2962 , w_2963 );
buf ( w_2962 , \358_b1 );
not ( w_2962 , w_2966 );
not ( w_2963 , w_2967 );
and ( w_2966 , w_2967 , \358_b0 );
or ( \1421_b1 , \1416_b1 , \1420_b1 );
not ( \1420_b1 , w_2968 );
and ( \1421_b0 , \1416_b0 , w_2969 );
and ( w_2968 , w_2969 , \1420_b0 );
buf ( \1422_b1 , RIb4bf0d8_85_b1 );
buf ( \1422_b0 , RIb4bf0d8_85_b0 );
or ( \1423_b1 , \1422_b1 , \345_b1 );
not ( \345_b1 , w_2970 );
and ( \1423_b0 , \1422_b0 , w_2971 );
and ( w_2970 , w_2971 , \345_b0 );
or ( \1424_b1 , \1420_b1 , \1423_b1 );
not ( \1423_b1 , w_2972 );
and ( \1424_b0 , \1420_b0 , w_2973 );
and ( w_2972 , w_2973 , \1423_b0 );
or ( \1425_b1 , \1416_b1 , \1423_b1 );
not ( \1423_b1 , w_2974 );
and ( \1425_b0 , \1416_b0 , w_2975 );
and ( w_2974 , w_2975 , \1423_b0 );
or ( \1427_b1 , \1263_b1 , \1267_b1 );
xor ( \1427_b0 , \1263_b0 , w_2976 );
not ( w_2976 , w_2977 );
and ( w_2977 , \1267_b1 , \1267_b0 );
or ( \1428_b1 , \1427_b1 , \1272_b1 );
xor ( \1428_b0 , \1427_b0 , w_2978 );
not ( w_2978 , w_2979 );
and ( w_2979 , \1272_b1 , \1272_b0 );
or ( \1429_b1 , \1426_b1 , \1428_b1 );
not ( \1428_b1 , w_2980 );
and ( \1429_b0 , \1426_b0 , w_2981 );
and ( w_2980 , w_2981 , \1428_b0 );
or ( \1430_b1 , \1303_b1 , w_2982 );
xor ( \1430_b0 , \1303_b0 , w_2984 );
not ( w_2984 , w_2985 );
and ( w_2985 , w_2982 , w_2983 );
buf ( w_2982 , \1305_b1 );
not ( w_2982 , w_2986 );
not ( w_2983 , w_2987 );
and ( w_2986 , w_2987 , \1305_b0 );
or ( \1431_b1 , \1428_b1 , \1430_b1 );
not ( \1430_b1 , w_2988 );
and ( \1431_b0 , \1428_b0 , w_2989 );
and ( w_2988 , w_2989 , \1430_b0 );
or ( \1432_b1 , \1426_b1 , \1430_b1 );
not ( \1430_b1 , w_2990 );
and ( \1432_b0 , \1426_b0 , w_2991 );
and ( w_2990 , w_2991 , \1430_b0 );
or ( \1434_b1 , \1412_b1 , \1433_b1 );
not ( \1433_b1 , w_2992 );
and ( \1434_b0 , \1412_b0 , w_2993 );
and ( w_2992 , w_2993 , \1433_b0 );
or ( \1435_b1 , \1247_b1 , \1251_b1 );
xor ( \1435_b0 , \1247_b0 , w_2994 );
not ( w_2994 , w_2995 );
and ( w_2995 , \1251_b1 , \1251_b0 );
or ( \1436_b1 , \1435_b1 , \1256_b1 );
xor ( \1436_b0 , \1435_b0 , w_2996 );
not ( w_2996 , w_2997 );
and ( w_2997 , \1256_b1 , \1256_b0 );
or ( \1437_b1 , \1283_b1 , \1287_b1 );
xor ( \1437_b0 , \1283_b0 , w_2998 );
not ( w_2998 , w_2999 );
and ( w_2999 , \1287_b1 , \1287_b0 );
or ( \1438_b1 , \1437_b1 , \1292_b1 );
xor ( \1438_b0 , \1437_b0 , w_3000 );
not ( w_3000 , w_3001 );
and ( w_3001 , \1292_b1 , \1292_b0 );
or ( \1439_b1 , \1436_b1 , \1438_b1 );
not ( \1438_b1 , w_3002 );
and ( \1439_b0 , \1436_b0 , w_3003 );
and ( w_3002 , w_3003 , \1438_b0 );
or ( \1440_b1 , \1433_b1 , \1439_b1 );
not ( \1439_b1 , w_3004 );
and ( \1440_b0 , \1433_b0 , w_3005 );
and ( w_3004 , w_3005 , \1439_b0 );
or ( \1441_b1 , \1412_b1 , \1439_b1 );
not ( \1439_b1 , w_3006 );
and ( \1441_b0 , \1412_b0 , w_3007 );
and ( w_3006 , w_3007 , \1439_b0 );
or ( \1443_b1 , \1259_b1 , \1275_b1 );
xor ( \1443_b0 , \1259_b0 , w_3008 );
not ( w_3008 , w_3009 );
and ( w_3009 , \1275_b1 , \1275_b0 );
or ( \1444_b1 , \1443_b1 , \1295_b1 );
xor ( \1444_b0 , \1443_b0 , w_3010 );
not ( w_3010 , w_3011 );
and ( w_3011 , \1295_b1 , \1295_b0 );
or ( \1445_b1 , \1306_b1 , \1310_b1 );
xor ( \1445_b0 , \1306_b0 , w_3012 );
not ( w_3012 , w_3013 );
and ( w_3013 , \1310_b1 , \1310_b0 );
or ( \1446_b1 , \1445_b1 , \1312_b1 );
xor ( \1446_b0 , \1445_b0 , w_3014 );
not ( w_3014 , w_3015 );
and ( w_3015 , \1312_b1 , \1312_b0 );
or ( \1447_b1 , \1444_b1 , \1446_b1 );
not ( \1446_b1 , w_3016 );
and ( \1447_b0 , \1444_b0 , w_3017 );
and ( w_3016 , w_3017 , \1446_b0 );
or ( \1448_b1 , \1318_b1 , \1320_b1 );
xor ( \1448_b0 , \1318_b0 , w_3018 );
not ( w_3018 , w_3019 );
and ( w_3019 , \1320_b1 , \1320_b0 );
or ( \1449_b1 , \1448_b1 , \1323_b1 );
xor ( \1449_b0 , \1448_b0 , w_3020 );
not ( w_3020 , w_3021 );
and ( w_3021 , \1323_b1 , \1323_b0 );
or ( \1450_b1 , \1446_b1 , \1449_b1 );
not ( \1449_b1 , w_3022 );
and ( \1450_b0 , \1446_b0 , w_3023 );
and ( w_3022 , w_3023 , \1449_b0 );
or ( \1451_b1 , \1444_b1 , \1449_b1 );
not ( \1449_b1 , w_3024 );
and ( \1451_b0 , \1444_b0 , w_3025 );
and ( w_3024 , w_3025 , \1449_b0 );
or ( \1453_b1 , \1442_b1 , \1452_b1 );
not ( \1452_b1 , w_3026 );
and ( \1453_b0 , \1442_b0 , w_3027 );
and ( w_3026 , w_3027 , \1452_b0 );
or ( \1454_b1 , \1331_b1 , \1332_b1 );
xor ( \1454_b0 , \1331_b0 , w_3028 );
not ( w_3028 , w_3029 );
and ( w_3029 , \1332_b1 , \1332_b0 );
or ( \1455_b1 , \1454_b1 , \1334_b1 );
xor ( \1455_b0 , \1454_b0 , w_3030 );
not ( w_3030 , w_3031 );
and ( w_3031 , \1334_b1 , \1334_b0 );
or ( \1456_b1 , \1452_b1 , \1455_b1 );
not ( \1455_b1 , w_3032 );
and ( \1456_b0 , \1452_b0 , w_3033 );
and ( w_3032 , w_3033 , \1455_b0 );
or ( \1457_b1 , \1442_b1 , \1455_b1 );
not ( \1455_b1 , w_3034 );
and ( \1457_b0 , \1442_b0 , w_3035 );
and ( w_3034 , w_3035 , \1455_b0 );
or ( \1459_b1 , \1193_b1 , \1198_b1 );
xor ( \1459_b0 , \1193_b0 , w_3036 );
not ( w_3036 , w_3037 );
and ( w_3037 , \1198_b1 , \1198_b0 );
or ( \1460_b1 , \1459_b1 , \1204_b1 );
xor ( \1460_b0 , \1459_b0 , w_3038 );
not ( w_3038 , w_3039 );
and ( w_3039 , \1204_b1 , \1204_b0 );
or ( \1461_b1 , \1458_b1 , \1460_b1 );
not ( \1460_b1 , w_3040 );
and ( \1461_b0 , \1458_b0 , w_3041 );
and ( w_3040 , w_3041 , \1460_b0 );
or ( \1462_b1 , \1329_b1 , \1337_b1 );
xor ( \1462_b0 , \1329_b0 , w_3042 );
not ( w_3042 , w_3043 );
and ( w_3043 , \1337_b1 , \1337_b0 );
or ( \1463_b1 , \1462_b1 , \1340_b1 );
xor ( \1463_b0 , \1462_b0 , w_3044 );
not ( w_3044 , w_3045 );
and ( w_3045 , \1340_b1 , \1340_b0 );
or ( \1464_b1 , \1460_b1 , \1463_b1 );
not ( \1463_b1 , w_3046 );
and ( \1464_b0 , \1460_b0 , w_3047 );
and ( w_3046 , w_3047 , \1463_b0 );
or ( \1465_b1 , \1458_b1 , \1463_b1 );
not ( \1463_b1 , w_3048 );
and ( \1465_b0 , \1458_b0 , w_3049 );
and ( w_3048 , w_3049 , \1463_b0 );
or ( \1467_b1 , \1343_b1 , \1345_b1 );
xor ( \1467_b0 , \1343_b0 , w_3050 );
not ( w_3050 , w_3051 );
and ( w_3051 , \1345_b1 , \1345_b0 );
or ( \1468_b1 , \1467_b1 , \1347_b1 );
xor ( \1468_b0 , \1467_b0 , w_3052 );
not ( w_3052 , w_3053 );
and ( w_3053 , \1347_b1 , \1347_b0 );
or ( \1469_b1 , \1466_b1 , \1468_b1 );
not ( \1468_b1 , w_3054 );
and ( \1469_b0 , \1466_b0 , w_3055 );
and ( w_3054 , w_3055 , \1468_b0 );
or ( \1470_b1 , \1356_b1 , \1469_b1 );
not ( \1469_b1 , w_3056 );
and ( \1470_b0 , \1356_b0 , w_3057 );
and ( w_3056 , w_3057 , \1469_b0 );
or ( \1471_b1 , \1356_b1 , \1469_b1 );
xor ( \1471_b0 , \1356_b0 , w_3058 );
not ( w_3058 , w_3059 );
and ( w_3059 , \1469_b1 , \1469_b0 );
or ( \1472_b1 , \1466_b1 , \1468_b1 );
xor ( \1472_b0 , \1466_b0 , w_3060 );
not ( w_3060 , w_3061 );
and ( w_3061 , \1468_b1 , \1468_b0 );
or ( \1473_b1 , \1174_b1 , \1358_b1 );
xor ( \1473_b0 , \1174_b0 , w_3062 );
not ( w_3062 , w_3063 );
and ( w_3063 , \1358_b1 , \1358_b0 );
or ( \1474_b1 , \1358_b1 , \1360_b1 );
xor ( \1474_b0 , \1358_b0 , w_3064 );
not ( w_3064 , w_3065 );
and ( w_3065 , \1360_b1 , \1360_b0 );
buf ( \1475_b1 , \1474_b1 );
not ( \1475_b1 , w_3066 );
not ( \1475_b0 , w_3067 );
and ( w_3066 , w_3067 , \1474_b0 );
or ( \1476_b1 , \1473_b1 , \1475_b1 );
not ( \1475_b1 , w_3068 );
and ( \1476_b0 , \1473_b0 , w_3069 );
and ( w_3068 , w_3069 , \1475_b0 );
or ( \1477_b1 , \159_b1 , \1476_b1 );
not ( \1476_b1 , w_3070 );
and ( \1477_b0 , \159_b0 , w_3071 );
and ( w_3070 , w_3071 , \1476_b0 );
buf ( \1478_b1 , \1477_b1 );
not ( \1478_b1 , w_3072 );
not ( \1478_b0 , w_3073 );
and ( w_3072 , w_3073 , \1477_b0 );
or ( \1479_b1 , \1478_b1 , w_3074 );
xor ( \1479_b0 , \1478_b0 , w_3076 );
not ( w_3076 , w_3077 );
and ( w_3077 , w_3074 , w_3075 );
buf ( w_3074 , \1363_b1 );
not ( w_3074 , w_3078 );
not ( w_3075 , w_3079 );
and ( w_3078 , w_3079 , \1363_b0 );
or ( \1480_b1 , \305_b1 , \1280_b1 );
not ( \1280_b1 , w_3080 );
and ( \1480_b0 , \305_b0 , w_3081 );
and ( w_3080 , w_3081 , \1280_b0 );
or ( \1481_b1 , \315_b1 , \1278_b1 );
not ( \1278_b1 , w_3082 );
and ( \1481_b0 , \315_b0 , w_3083 );
and ( w_3082 , w_3083 , \1278_b0 );
or ( \1482_b1 , \1480_b1 , w_3085 );
not ( w_3085 , w_3086 );
and ( \1482_b0 , \1480_b0 , w_3087 );
and ( w_3086 ,  , w_3087 );
buf ( w_3085 , \1481_b1 );
not ( w_3085 , w_3088 );
not (  , w_3089 );
and ( w_3088 , w_3089 , \1481_b0 );
or ( \1483_b1 , \1482_b1 , w_3090 );
xor ( \1483_b0 , \1482_b0 , w_3092 );
not ( w_3092 , w_3093 );
and ( w_3093 , w_3090 , w_3091 );
buf ( w_3090 , \1177_b1 );
not ( w_3090 , w_3094 );
not ( w_3091 , w_3095 );
and ( w_3094 , w_3095 , \1177_b0 );
or ( \1484_b1 , \1479_b1 , \1483_b1 );
not ( \1483_b1 , w_3096 );
and ( \1484_b0 , \1479_b0 , w_3097 );
and ( w_3096 , w_3097 , \1483_b0 );
or ( \1485_b1 , \323_b1 , \1062_b1 );
not ( \1062_b1 , w_3098 );
and ( \1485_b0 , \323_b0 , w_3099 );
and ( w_3098 , w_3099 , \1062_b0 );
or ( \1486_b1 , \333_b1 , \1060_b1 );
not ( \1060_b1 , w_3100 );
and ( \1486_b0 , \333_b0 , w_3101 );
and ( w_3100 , w_3101 , \1060_b0 );
or ( \1487_b1 , \1485_b1 , w_3103 );
not ( w_3103 , w_3104 );
and ( \1487_b0 , \1485_b0 , w_3105 );
and ( w_3104 ,  , w_3105 );
buf ( w_3103 , \1486_b1 );
not ( w_3103 , w_3106 );
not (  , w_3107 );
and ( w_3106 , w_3107 , \1486_b0 );
or ( \1488_b1 , \1487_b1 , w_3108 );
xor ( \1488_b0 , \1487_b0 , w_3110 );
not ( w_3110 , w_3111 );
and ( w_3111 , w_3108 , w_3109 );
buf ( w_3108 , \984_b1 );
not ( w_3108 , w_3112 );
not ( w_3109 , w_3113 );
and ( w_3112 , w_3113 , \984_b0 );
or ( \1489_b1 , \1483_b1 , \1488_b1 );
not ( \1488_b1 , w_3114 );
and ( \1489_b0 , \1483_b0 , w_3115 );
and ( w_3114 , w_3115 , \1488_b0 );
or ( \1490_b1 , \1479_b1 , \1488_b1 );
not ( \1488_b1 , w_3116 );
and ( \1490_b0 , \1479_b0 , w_3117 );
and ( w_3116 , w_3117 , \1488_b0 );
or ( \1492_b1 , \343_b1 , \912_b1 );
not ( \912_b1 , w_3118 );
and ( \1492_b0 , \343_b0 , w_3119 );
and ( w_3118 , w_3119 , \912_b0 );
or ( \1493_b1 , \353_b1 , \910_b1 );
not ( \910_b1 , w_3120 );
and ( \1493_b0 , \353_b0 , w_3121 );
and ( w_3120 , w_3121 , \910_b0 );
or ( \1494_b1 , \1492_b1 , w_3123 );
not ( w_3123 , w_3124 );
and ( \1494_b0 , \1492_b0 , w_3125 );
and ( w_3124 ,  , w_3125 );
buf ( w_3123 , \1493_b1 );
not ( w_3123 , w_3126 );
not (  , w_3127 );
and ( w_3126 , w_3127 , \1493_b0 );
or ( \1495_b1 , \1494_b1 , w_3128 );
xor ( \1495_b0 , \1494_b0 , w_3130 );
not ( w_3130 , w_3131 );
and ( w_3131 , w_3128 , w_3129 );
buf ( w_3128 , \818_b1 );
not ( w_3128 , w_3132 );
not ( w_3129 , w_3133 );
and ( w_3132 , w_3133 , \818_b0 );
or ( \1496_b1 , \444_b1 , \740_b1 );
not ( \740_b1 , w_3134 );
and ( \1496_b0 , \444_b0 , w_3135 );
and ( w_3134 , w_3135 , \740_b0 );
or ( \1497_b1 , \360_b1 , \738_b1 );
not ( \738_b1 , w_3136 );
and ( \1497_b0 , \360_b0 , w_3137 );
and ( w_3136 , w_3137 , \738_b0 );
or ( \1498_b1 , \1496_b1 , w_3139 );
not ( w_3139 , w_3140 );
and ( \1498_b0 , \1496_b0 , w_3141 );
and ( w_3140 ,  , w_3141 );
buf ( w_3139 , \1497_b1 );
not ( w_3139 , w_3142 );
not (  , w_3143 );
and ( w_3142 , w_3143 , \1497_b0 );
or ( \1499_b1 , \1498_b1 , w_3144 );
xor ( \1499_b0 , \1498_b0 , w_3146 );
not ( w_3146 , w_3147 );
and ( w_3147 , w_3144 , w_3145 );
buf ( w_3144 , \668_b1 );
not ( w_3144 , w_3148 );
not ( w_3145 , w_3149 );
and ( w_3148 , w_3149 , \668_b0 );
or ( \1500_b1 , \1495_b1 , \1499_b1 );
not ( \1499_b1 , w_3150 );
and ( \1500_b0 , \1495_b0 , w_3151 );
and ( w_3150 , w_3151 , \1499_b0 );
or ( \1501_b1 , \593_b1 , \604_b1 );
not ( \604_b1 , w_3152 );
and ( \1501_b0 , \593_b0 , w_3153 );
and ( w_3152 , w_3153 , \604_b0 );
or ( \1502_b1 , \495_b1 , \602_b1 );
not ( \602_b1 , w_3154 );
and ( \1502_b0 , \495_b0 , w_3155 );
and ( w_3154 , w_3155 , \602_b0 );
or ( \1503_b1 , \1501_b1 , w_3157 );
not ( w_3157 , w_3158 );
and ( \1503_b0 , \1501_b0 , w_3159 );
and ( w_3158 ,  , w_3159 );
buf ( w_3157 , \1502_b1 );
not ( w_3157 , w_3160 );
not (  , w_3161 );
and ( w_3160 , w_3161 , \1502_b0 );
or ( \1504_b1 , \1503_b1 , w_3162 );
xor ( \1504_b0 , \1503_b0 , w_3164 );
not ( w_3164 , w_3165 );
and ( w_3165 , w_3162 , w_3163 );
buf ( w_3162 , \561_b1 );
not ( w_3162 , w_3166 );
not ( w_3163 , w_3167 );
and ( w_3166 , w_3167 , \561_b0 );
or ( \1505_b1 , \1499_b1 , \1504_b1 );
not ( \1504_b1 , w_3168 );
and ( \1505_b0 , \1499_b0 , w_3169 );
and ( w_3168 , w_3169 , \1504_b0 );
or ( \1506_b1 , \1495_b1 , \1504_b1 );
not ( \1504_b1 , w_3170 );
and ( \1506_b0 , \1495_b0 , w_3171 );
and ( w_3170 , w_3171 , \1504_b0 );
or ( \1508_b1 , \1491_b1 , \1507_b1 );
not ( \1507_b1 , w_3172 );
and ( \1508_b0 , \1491_b0 , w_3173 );
and ( w_3172 , w_3173 , \1507_b0 );
or ( \1509_b1 , \703_b1 , \503_b1 );
not ( \503_b1 , w_3174 );
and ( \1509_b0 , \703_b0 , w_3175 );
and ( w_3174 , w_3175 , \503_b0 );
or ( \1510_b1 , \621_b1 , \501_b1 );
not ( \501_b1 , w_3176 );
and ( \1510_b0 , \621_b0 , w_3177 );
and ( w_3176 , w_3177 , \501_b0 );
or ( \1511_b1 , \1509_b1 , w_3179 );
not ( w_3179 , w_3180 );
and ( \1511_b0 , \1509_b0 , w_3181 );
and ( w_3180 ,  , w_3181 );
buf ( w_3179 , \1510_b1 );
not ( w_3179 , w_3182 );
not (  , w_3183 );
and ( w_3182 , w_3183 , \1510_b0 );
or ( \1512_b1 , \1511_b1 , w_3184 );
xor ( \1512_b0 , \1511_b0 , w_3186 );
not ( w_3186 , w_3187 );
and ( w_3187 , w_3184 , w_3185 );
buf ( w_3184 , \455_b1 );
not ( w_3184 , w_3188 );
not ( w_3185 , w_3189 );
and ( w_3188 , w_3189 , \455_b0 );
or ( \1513_b1 , \841_b1 , \298_b1 );
not ( \298_b1 , w_3190 );
and ( \1513_b0 , \841_b0 , w_3191 );
and ( w_3190 , w_3191 , \298_b0 );
or ( \1514_b1 , \777_b1 , \296_b1 );
not ( \296_b1 , w_3192 );
and ( \1514_b0 , \777_b0 , w_3193 );
and ( w_3192 , w_3193 , \296_b0 );
or ( \1515_b1 , \1513_b1 , w_3195 );
not ( w_3195 , w_3196 );
and ( \1515_b0 , \1513_b0 , w_3197 );
and ( w_3196 ,  , w_3197 );
buf ( w_3195 , \1514_b1 );
not ( w_3195 , w_3198 );
not (  , w_3199 );
and ( w_3198 , w_3199 , \1514_b0 );
or ( \1516_b1 , \1515_b1 , w_3200 );
xor ( \1516_b0 , \1515_b0 , w_3202 );
not ( w_3202 , w_3203 );
and ( w_3203 , w_3200 , w_3201 );
buf ( w_3200 , \303_b1 );
not ( w_3200 , w_3204 );
not ( w_3201 , w_3205 );
and ( w_3204 , w_3205 , \303_b0 );
or ( \1517_b1 , \1512_b1 , \1516_b1 );
not ( \1516_b1 , w_3206 );
and ( \1517_b0 , \1512_b0 , w_3207 );
and ( w_3206 , w_3207 , \1516_b0 );
or ( \1518_b1 , \1104_b1 , \313_b1 );
not ( \313_b1 , w_3208 );
and ( \1518_b0 , \1104_b0 , w_3209 );
and ( w_3208 , w_3209 , \313_b0 );
or ( \1519_b1 , \904_b1 , \311_b1 );
not ( \311_b1 , w_3210 );
and ( \1519_b0 , \904_b0 , w_3211 );
and ( w_3210 , w_3211 , \311_b0 );
or ( \1520_b1 , \1518_b1 , w_3213 );
not ( w_3213 , w_3214 );
and ( \1520_b0 , \1518_b0 , w_3215 );
and ( w_3214 ,  , w_3215 );
buf ( w_3213 , \1519_b1 );
not ( w_3213 , w_3216 );
not (  , w_3217 );
and ( w_3216 , w_3217 , \1519_b0 );
or ( \1521_b1 , \1520_b1 , w_3218 );
xor ( \1521_b0 , \1520_b0 , w_3220 );
not ( w_3220 , w_3221 );
and ( w_3221 , w_3218 , w_3219 );
buf ( w_3218 , \320_b1 );
not ( w_3218 , w_3222 );
not ( w_3219 , w_3223 );
and ( w_3222 , w_3223 , \320_b0 );
or ( \1522_b1 , \1516_b1 , \1521_b1 );
not ( \1521_b1 , w_3224 );
and ( \1522_b0 , \1516_b0 , w_3225 );
and ( w_3224 , w_3225 , \1521_b0 );
or ( \1523_b1 , \1512_b1 , \1521_b1 );
not ( \1521_b1 , w_3226 );
and ( \1523_b0 , \1512_b0 , w_3227 );
and ( w_3226 , w_3227 , \1521_b0 );
or ( \1525_b1 , \1507_b1 , \1524_b1 );
not ( \1524_b1 , w_3228 );
and ( \1525_b0 , \1507_b0 , w_3229 );
and ( w_3228 , w_3229 , \1524_b0 );
or ( \1526_b1 , \1491_b1 , \1524_b1 );
not ( \1524_b1 , w_3230 );
and ( \1526_b0 , \1491_b0 , w_3231 );
and ( w_3230 , w_3231 , \1524_b0 );
or ( \1528_b1 , \1299_b1 , \331_b1 );
not ( \331_b1 , w_3232 );
and ( \1528_b0 , \1299_b0 , w_3233 );
and ( w_3232 , w_3233 , \331_b0 );
or ( \1529_b1 , \1194_b1 , \329_b1 );
not ( \329_b1 , w_3234 );
and ( \1529_b0 , \1194_b0 , w_3235 );
and ( w_3234 , w_3235 , \329_b0 );
or ( \1530_b1 , \1528_b1 , w_3237 );
not ( w_3237 , w_3238 );
and ( \1530_b0 , \1528_b0 , w_3239 );
and ( w_3238 ,  , w_3239 );
buf ( w_3237 , \1529_b1 );
not ( w_3237 , w_3240 );
not (  , w_3241 );
and ( w_3240 , w_3241 , \1529_b0 );
or ( \1531_b1 , \1530_b1 , w_3242 );
xor ( \1531_b0 , \1530_b0 , w_3244 );
not ( w_3244 , w_3245 );
and ( w_3245 , w_3242 , w_3243 );
buf ( w_3242 , \338_b1 );
not ( w_3242 , w_3246 );
not ( w_3243 , w_3247 );
and ( w_3246 , w_3247 , \338_b0 );
or ( \1532_b1 , \1422_b1 , \351_b1 );
not ( \351_b1 , w_3248 );
and ( \1532_b0 , \1422_b0 , w_3249 );
and ( w_3248 , w_3249 , \351_b0 );
or ( \1533_b1 , \1304_b1 , \349_b1 );
not ( \349_b1 , w_3250 );
and ( \1533_b0 , \1304_b0 , w_3251 );
and ( w_3250 , w_3251 , \349_b0 );
or ( \1534_b1 , \1532_b1 , w_3253 );
not ( w_3253 , w_3254 );
and ( \1534_b0 , \1532_b0 , w_3255 );
and ( w_3254 ,  , w_3255 );
buf ( w_3253 , \1533_b1 );
not ( w_3253 , w_3256 );
not (  , w_3257 );
and ( w_3256 , w_3257 , \1533_b0 );
or ( \1535_b1 , \1534_b1 , w_3258 );
xor ( \1535_b0 , \1534_b0 , w_3260 );
not ( w_3260 , w_3261 );
and ( w_3261 , w_3258 , w_3259 );
buf ( w_3258 , \358_b1 );
not ( w_3258 , w_3262 );
not ( w_3259 , w_3263 );
and ( w_3262 , w_3263 , \358_b0 );
or ( \1536_b1 , \1531_b1 , \1535_b1 );
not ( \1535_b1 , w_3264 );
and ( \1536_b0 , \1531_b0 , w_3265 );
and ( w_3264 , w_3265 , \1535_b0 );
buf ( \1537_b1 , RIb4bf060_86_b1 );
buf ( \1537_b0 , RIb4bf060_86_b0 );
or ( \1538_b1 , \1537_b1 , \345_b1 );
not ( \345_b1 , w_3266 );
and ( \1538_b0 , \1537_b0 , w_3267 );
and ( w_3266 , w_3267 , \345_b0 );
or ( \1539_b1 , \1535_b1 , \1538_b1 );
not ( \1538_b1 , w_3268 );
and ( \1539_b0 , \1535_b0 , w_3269 );
and ( w_3268 , w_3269 , \1538_b0 );
or ( \1540_b1 , \1531_b1 , \1538_b1 );
not ( \1538_b1 , w_3270 );
and ( \1540_b0 , \1531_b0 , w_3271 );
and ( w_3270 , w_3271 , \1538_b0 );
or ( \1542_b1 , \1416_b1 , \1420_b1 );
xor ( \1542_b0 , \1416_b0 , w_3272 );
not ( w_3272 , w_3273 );
and ( w_3273 , \1420_b1 , \1420_b0 );
or ( \1543_b1 , \1542_b1 , \1423_b1 );
xor ( \1543_b0 , \1542_b0 , w_3274 );
not ( w_3274 , w_3275 );
and ( w_3275 , \1423_b1 , \1423_b0 );
or ( \1544_b1 , \1541_b1 , \1543_b1 );
not ( \1543_b1 , w_3276 );
and ( \1544_b0 , \1541_b0 , w_3277 );
and ( w_3276 , w_3277 , \1543_b0 );
or ( \1545_b1 , \1397_b1 , \1401_b1 );
xor ( \1545_b0 , \1397_b0 , w_3278 );
not ( w_3278 , w_3279 );
and ( w_3279 , \1401_b1 , \1401_b0 );
or ( \1546_b1 , \1545_b1 , \1406_b1 );
xor ( \1546_b0 , \1545_b0 , w_3280 );
not ( w_3280 , w_3281 );
and ( w_3281 , \1406_b1 , \1406_b0 );
or ( \1547_b1 , \1543_b1 , \1546_b1 );
not ( \1546_b1 , w_3282 );
and ( \1547_b0 , \1543_b0 , w_3283 );
and ( w_3282 , w_3283 , \1546_b0 );
or ( \1548_b1 , \1541_b1 , \1546_b1 );
not ( \1546_b1 , w_3284 );
and ( \1548_b0 , \1541_b0 , w_3285 );
and ( w_3284 , w_3285 , \1546_b0 );
or ( \1550_b1 , \1527_b1 , \1549_b1 );
not ( \1549_b1 , w_3286 );
and ( \1550_b0 , \1527_b0 , w_3287 );
and ( w_3286 , w_3287 , \1549_b0 );
or ( \1551_b1 , \1364_b1 , \1368_b1 );
xor ( \1551_b0 , \1364_b0 , w_3288 );
not ( w_3288 , w_3289 );
and ( w_3289 , \1368_b1 , \1368_b0 );
or ( \1552_b1 , \1551_b1 , \1373_b1 );
xor ( \1552_b0 , \1551_b0 , w_3290 );
not ( w_3290 , w_3291 );
and ( w_3291 , \1373_b1 , \1373_b0 );
or ( \1553_b1 , \1380_b1 , \1384_b1 );
xor ( \1553_b0 , \1380_b0 , w_3292 );
not ( w_3292 , w_3293 );
and ( w_3293 , \1384_b1 , \1384_b0 );
or ( \1554_b1 , \1553_b1 , \1389_b1 );
xor ( \1554_b0 , \1553_b0 , w_3294 );
not ( w_3294 , w_3295 );
and ( w_3295 , \1389_b1 , \1389_b0 );
or ( \1555_b1 , \1552_b1 , \1554_b1 );
not ( \1554_b1 , w_3296 );
and ( \1555_b0 , \1552_b0 , w_3297 );
and ( w_3296 , w_3297 , \1554_b0 );
or ( \1556_b1 , \1549_b1 , \1555_b1 );
not ( \1555_b1 , w_3298 );
and ( \1556_b0 , \1549_b0 , w_3299 );
and ( w_3298 , w_3299 , \1555_b0 );
or ( \1557_b1 , \1527_b1 , \1555_b1 );
not ( \1555_b1 , w_3300 );
and ( \1557_b0 , \1527_b0 , w_3301 );
and ( w_3300 , w_3301 , \1555_b0 );
or ( \1559_b1 , \1376_b1 , \1392_b1 );
xor ( \1559_b0 , \1376_b0 , w_3302 );
not ( w_3302 , w_3303 );
and ( w_3303 , \1392_b1 , \1392_b0 );
or ( \1560_b1 , \1559_b1 , \1409_b1 );
xor ( \1560_b0 , \1559_b0 , w_3304 );
not ( w_3304 , w_3305 );
and ( w_3305 , \1409_b1 , \1409_b0 );
or ( \1561_b1 , \1426_b1 , \1428_b1 );
xor ( \1561_b0 , \1426_b0 , w_3306 );
not ( w_3306 , w_3307 );
and ( w_3307 , \1428_b1 , \1428_b0 );
or ( \1562_b1 , \1561_b1 , \1430_b1 );
xor ( \1562_b0 , \1561_b0 , w_3308 );
not ( w_3308 , w_3309 );
and ( w_3309 , \1430_b1 , \1430_b0 );
or ( \1563_b1 , \1560_b1 , \1562_b1 );
not ( \1562_b1 , w_3310 );
and ( \1563_b0 , \1560_b0 , w_3311 );
and ( w_3310 , w_3311 , \1562_b0 );
or ( \1564_b1 , \1436_b1 , \1438_b1 );
xor ( \1564_b0 , \1436_b0 , w_3312 );
not ( w_3312 , w_3313 );
and ( w_3313 , \1438_b1 , \1438_b0 );
or ( \1565_b1 , \1562_b1 , \1564_b1 );
not ( \1564_b1 , w_3314 );
and ( \1565_b0 , \1562_b0 , w_3315 );
and ( w_3314 , w_3315 , \1564_b0 );
or ( \1566_b1 , \1560_b1 , \1564_b1 );
not ( \1564_b1 , w_3316 );
and ( \1566_b0 , \1560_b0 , w_3317 );
and ( w_3316 , w_3317 , \1564_b0 );
or ( \1568_b1 , \1558_b1 , \1567_b1 );
not ( \1567_b1 , w_3318 );
and ( \1568_b0 , \1558_b0 , w_3319 );
and ( w_3318 , w_3319 , \1567_b0 );
or ( \1569_b1 , \1444_b1 , \1446_b1 );
xor ( \1569_b0 , \1444_b0 , w_3320 );
not ( w_3320 , w_3321 );
and ( w_3321 , \1446_b1 , \1446_b0 );
or ( \1570_b1 , \1569_b1 , \1449_b1 );
xor ( \1570_b0 , \1569_b0 , w_3322 );
not ( w_3322 , w_3323 );
and ( w_3323 , \1449_b1 , \1449_b0 );
or ( \1571_b1 , \1567_b1 , \1570_b1 );
not ( \1570_b1 , w_3324 );
and ( \1571_b0 , \1567_b0 , w_3325 );
and ( w_3324 , w_3325 , \1570_b0 );
or ( \1572_b1 , \1558_b1 , \1570_b1 );
not ( \1570_b1 , w_3326 );
and ( \1572_b0 , \1558_b0 , w_3327 );
and ( w_3326 , w_3327 , \1570_b0 );
or ( \1574_b1 , \1298_b1 , \1315_b1 );
xor ( \1574_b0 , \1298_b0 , w_3328 );
not ( w_3328 , w_3329 );
and ( w_3329 , \1315_b1 , \1315_b0 );
or ( \1575_b1 , \1574_b1 , \1326_b1 );
xor ( \1575_b0 , \1574_b0 , w_3330 );
not ( w_3330 , w_3331 );
and ( w_3331 , \1326_b1 , \1326_b0 );
or ( \1576_b1 , \1573_b1 , \1575_b1 );
not ( \1575_b1 , w_3332 );
and ( \1576_b0 , \1573_b0 , w_3333 );
and ( w_3332 , w_3333 , \1575_b0 );
or ( \1577_b1 , \1442_b1 , \1452_b1 );
xor ( \1577_b0 , \1442_b0 , w_3334 );
not ( w_3334 , w_3335 );
and ( w_3335 , \1452_b1 , \1452_b0 );
or ( \1578_b1 , \1577_b1 , \1455_b1 );
xor ( \1578_b0 , \1577_b0 , w_3336 );
not ( w_3336 , w_3337 );
and ( w_3337 , \1455_b1 , \1455_b0 );
or ( \1579_b1 , \1575_b1 , \1578_b1 );
not ( \1578_b1 , w_3338 );
and ( \1579_b0 , \1575_b0 , w_3339 );
and ( w_3338 , w_3339 , \1578_b0 );
or ( \1580_b1 , \1573_b1 , \1578_b1 );
not ( \1578_b1 , w_3340 );
and ( \1580_b0 , \1573_b0 , w_3341 );
and ( w_3340 , w_3341 , \1578_b0 );
or ( \1582_b1 , \1458_b1 , \1460_b1 );
xor ( \1582_b0 , \1458_b0 , w_3342 );
not ( w_3342 , w_3343 );
and ( w_3343 , \1460_b1 , \1460_b0 );
or ( \1583_b1 , \1582_b1 , \1463_b1 );
xor ( \1583_b0 , \1582_b0 , w_3344 );
not ( w_3344 , w_3345 );
and ( w_3345 , \1463_b1 , \1463_b0 );
or ( \1584_b1 , \1581_b1 , \1583_b1 );
not ( \1583_b1 , w_3346 );
and ( \1584_b0 , \1581_b0 , w_3347 );
and ( w_3346 , w_3347 , \1583_b0 );
or ( \1585_b1 , \1472_b1 , \1584_b1 );
not ( \1584_b1 , w_3348 );
and ( \1585_b0 , \1472_b0 , w_3349 );
and ( w_3348 , w_3349 , \1584_b0 );
or ( \1586_b1 , \1472_b1 , \1584_b1 );
xor ( \1586_b0 , \1472_b0 , w_3350 );
not ( w_3350 , w_3351 );
and ( w_3351 , \1584_b1 , \1584_b0 );
or ( \1587_b1 , \1581_b1 , \1583_b1 );
xor ( \1587_b0 , \1581_b0 , w_3352 );
not ( w_3352 , w_3353 );
and ( w_3353 , \1583_b1 , \1583_b0 );
or ( \1588_b1 , \621_b1 , \604_b1 );
not ( \604_b1 , w_3354 );
and ( \1588_b0 , \621_b0 , w_3355 );
and ( w_3354 , w_3355 , \604_b0 );
or ( \1589_b1 , \593_b1 , \602_b1 );
not ( \602_b1 , w_3356 );
and ( \1589_b0 , \593_b0 , w_3357 );
and ( w_3356 , w_3357 , \602_b0 );
or ( \1590_b1 , \1588_b1 , w_3359 );
not ( w_3359 , w_3360 );
and ( \1590_b0 , \1588_b0 , w_3361 );
and ( w_3360 ,  , w_3361 );
buf ( w_3359 , \1589_b1 );
not ( w_3359 , w_3362 );
not (  , w_3363 );
and ( w_3362 , w_3363 , \1589_b0 );
or ( \1591_b1 , \1590_b1 , w_3364 );
xor ( \1591_b0 , \1590_b0 , w_3366 );
not ( w_3366 , w_3367 );
and ( w_3367 , w_3364 , w_3365 );
buf ( w_3364 , \561_b1 );
not ( w_3364 , w_3368 );
not ( w_3365 , w_3369 );
and ( w_3368 , w_3369 , \561_b0 );
or ( \1592_b1 , \777_b1 , \503_b1 );
not ( \503_b1 , w_3370 );
and ( \1592_b0 , \777_b0 , w_3371 );
and ( w_3370 , w_3371 , \503_b0 );
or ( \1593_b1 , \703_b1 , \501_b1 );
not ( \501_b1 , w_3372 );
and ( \1593_b0 , \703_b0 , w_3373 );
and ( w_3372 , w_3373 , \501_b0 );
or ( \1594_b1 , \1592_b1 , w_3375 );
not ( w_3375 , w_3376 );
and ( \1594_b0 , \1592_b0 , w_3377 );
and ( w_3376 ,  , w_3377 );
buf ( w_3375 , \1593_b1 );
not ( w_3375 , w_3378 );
not (  , w_3379 );
and ( w_3378 , w_3379 , \1593_b0 );
or ( \1595_b1 , \1594_b1 , w_3380 );
xor ( \1595_b0 , \1594_b0 , w_3382 );
not ( w_3382 , w_3383 );
and ( w_3383 , w_3380 , w_3381 );
buf ( w_3380 , \455_b1 );
not ( w_3380 , w_3384 );
not ( w_3381 , w_3385 );
and ( w_3384 , w_3385 , \455_b0 );
or ( \1596_b1 , \1591_b1 , \1595_b1 );
not ( \1595_b1 , w_3386 );
and ( \1596_b0 , \1591_b0 , w_3387 );
and ( w_3386 , w_3387 , \1595_b0 );
or ( \1597_b1 , \904_b1 , \298_b1 );
not ( \298_b1 , w_3388 );
and ( \1597_b0 , \904_b0 , w_3389 );
and ( w_3388 , w_3389 , \298_b0 );
or ( \1598_b1 , \841_b1 , \296_b1 );
not ( \296_b1 , w_3390 );
and ( \1598_b0 , \841_b0 , w_3391 );
and ( w_3390 , w_3391 , \296_b0 );
or ( \1599_b1 , \1597_b1 , w_3393 );
not ( w_3393 , w_3394 );
and ( \1599_b0 , \1597_b0 , w_3395 );
and ( w_3394 ,  , w_3395 );
buf ( w_3393 , \1598_b1 );
not ( w_3393 , w_3396 );
not (  , w_3397 );
and ( w_3396 , w_3397 , \1598_b0 );
or ( \1600_b1 , \1599_b1 , w_3398 );
xor ( \1600_b0 , \1599_b0 , w_3400 );
not ( w_3400 , w_3401 );
and ( w_3401 , w_3398 , w_3399 );
buf ( w_3398 , \303_b1 );
not ( w_3398 , w_3402 );
not ( w_3399 , w_3403 );
and ( w_3402 , w_3403 , \303_b0 );
or ( \1601_b1 , \1595_b1 , \1600_b1 );
not ( \1600_b1 , w_3404 );
and ( \1601_b0 , \1595_b0 , w_3405 );
and ( w_3404 , w_3405 , \1600_b0 );
or ( \1602_b1 , \1591_b1 , \1600_b1 );
not ( \1600_b1 , w_3406 );
and ( \1602_b0 , \1591_b0 , w_3407 );
and ( w_3406 , w_3407 , \1600_b0 );
and ( \1604_nR12c_b1 , RIb4c2e40_56_b1 , w_3408 );
xor ( w_3408 , RIb4c2e40_56_b0 , \288_b1 );
not ( \288_b1 , w_3409 );
and ( \1604_nR12c_b0 , w_3409 , \288_b0 );
buf ( \1605_b1 , \1604_nR12c_b1 );
buf ( \1605_b0 , \1604_nR12c_b0 );
and ( \1606_nR12b_b1 , RIb4c2dc8_57_b1 , w_3410 );
xor ( w_3410 , RIb4c2dc8_57_b0 , \288_b1 );
not ( \288_b1 , w_3411 );
and ( \1606_nR12b_b0 , w_3411 , \288_b0 );
buf ( \1607_b1 , \1606_nR12b_b1 );
buf ( \1607_b0 , \1606_nR12b_b0 );
or ( \1608_b1 , \1605_b1 , \1607_b1 );
not ( \1607_b1 , w_3412 );
and ( \1608_b0 , \1605_b0 , w_3413 );
and ( w_3412 , w_3413 , \1607_b0 );
buf ( \1609_b1 , \1608_b1 );
not ( \1609_b1 , w_3414 );
not ( \1609_b0 , w_3415 );
and ( w_3414 , w_3415 , \1608_b0 );
or ( \1610_b1 , \1360_b1 , \1609_b1 );
not ( \1609_b1 , w_3416 );
and ( \1610_b0 , \1360_b0 , w_3417 );
and ( w_3416 , w_3417 , \1609_b0 );
buf ( \1611_b1 , \1610_b1 );
not ( \1611_b1 , w_3418 );
not ( \1611_b0 , w_3419 );
and ( w_3418 , w_3419 , \1610_b0 );
or ( \1612_b1 , \315_b1 , \1476_b1 );
not ( \1476_b1 , w_3420 );
and ( \1612_b0 , \315_b0 , w_3421 );
and ( w_3420 , w_3421 , \1476_b0 );
or ( \1613_b1 , \159_b1 , \1474_b1 );
not ( \1474_b1 , w_3422 );
and ( \1613_b0 , \159_b0 , w_3423 );
and ( w_3422 , w_3423 , \1474_b0 );
or ( \1614_b1 , \1612_b1 , w_3425 );
not ( w_3425 , w_3426 );
and ( \1614_b0 , \1612_b0 , w_3427 );
and ( w_3426 ,  , w_3427 );
buf ( w_3425 , \1613_b1 );
not ( w_3425 , w_3428 );
not (  , w_3429 );
and ( w_3428 , w_3429 , \1613_b0 );
or ( \1615_b1 , \1614_b1 , w_3430 );
xor ( \1615_b0 , \1614_b0 , w_3432 );
not ( w_3432 , w_3433 );
and ( w_3433 , w_3430 , w_3431 );
buf ( w_3430 , \1363_b1 );
not ( w_3430 , w_3434 );
not ( w_3431 , w_3435 );
and ( w_3434 , w_3435 , \1363_b0 );
or ( \1616_b1 , \1611_b1 , \1615_b1 );
not ( \1615_b1 , w_3436 );
and ( \1616_b0 , \1611_b0 , w_3437 );
and ( w_3436 , w_3437 , \1615_b0 );
or ( \1617_b1 , \333_b1 , \1280_b1 );
not ( \1280_b1 , w_3438 );
and ( \1617_b0 , \333_b0 , w_3439 );
and ( w_3438 , w_3439 , \1280_b0 );
or ( \1618_b1 , \305_b1 , \1278_b1 );
not ( \1278_b1 , w_3440 );
and ( \1618_b0 , \305_b0 , w_3441 );
and ( w_3440 , w_3441 , \1278_b0 );
or ( \1619_b1 , \1617_b1 , w_3443 );
not ( w_3443 , w_3444 );
and ( \1619_b0 , \1617_b0 , w_3445 );
and ( w_3444 ,  , w_3445 );
buf ( w_3443 , \1618_b1 );
not ( w_3443 , w_3446 );
not (  , w_3447 );
and ( w_3446 , w_3447 , \1618_b0 );
or ( \1620_b1 , \1619_b1 , w_3448 );
xor ( \1620_b0 , \1619_b0 , w_3450 );
not ( w_3450 , w_3451 );
and ( w_3451 , w_3448 , w_3449 );
buf ( w_3448 , \1177_b1 );
not ( w_3448 , w_3452 );
not ( w_3449 , w_3453 );
and ( w_3452 , w_3453 , \1177_b0 );
or ( \1621_b1 , \1615_b1 , \1620_b1 );
not ( \1620_b1 , w_3454 );
and ( \1621_b0 , \1615_b0 , w_3455 );
and ( w_3454 , w_3455 , \1620_b0 );
or ( \1622_b1 , \1611_b1 , \1620_b1 );
not ( \1620_b1 , w_3456 );
and ( \1622_b0 , \1611_b0 , w_3457 );
and ( w_3456 , w_3457 , \1620_b0 );
or ( \1624_b1 , \1603_b1 , \1623_b1 );
not ( \1623_b1 , w_3458 );
and ( \1624_b0 , \1603_b0 , w_3459 );
and ( w_3458 , w_3459 , \1623_b0 );
or ( \1625_b1 , \353_b1 , \1062_b1 );
not ( \1062_b1 , w_3460 );
and ( \1625_b0 , \353_b0 , w_3461 );
and ( w_3460 , w_3461 , \1062_b0 );
or ( \1626_b1 , \323_b1 , \1060_b1 );
not ( \1060_b1 , w_3462 );
and ( \1626_b0 , \323_b0 , w_3463 );
and ( w_3462 , w_3463 , \1060_b0 );
or ( \1627_b1 , \1625_b1 , w_3465 );
not ( w_3465 , w_3466 );
and ( \1627_b0 , \1625_b0 , w_3467 );
and ( w_3466 ,  , w_3467 );
buf ( w_3465 , \1626_b1 );
not ( w_3465 , w_3468 );
not (  , w_3469 );
and ( w_3468 , w_3469 , \1626_b0 );
or ( \1628_b1 , \1627_b1 , w_3470 );
xor ( \1628_b0 , \1627_b0 , w_3472 );
not ( w_3472 , w_3473 );
and ( w_3473 , w_3470 , w_3471 );
buf ( w_3470 , \984_b1 );
not ( w_3470 , w_3474 );
not ( w_3471 , w_3475 );
and ( w_3474 , w_3475 , \984_b0 );
or ( \1629_b1 , \360_b1 , \912_b1 );
not ( \912_b1 , w_3476 );
and ( \1629_b0 , \360_b0 , w_3477 );
and ( w_3476 , w_3477 , \912_b0 );
or ( \1630_b1 , \343_b1 , \910_b1 );
not ( \910_b1 , w_3478 );
and ( \1630_b0 , \343_b0 , w_3479 );
and ( w_3478 , w_3479 , \910_b0 );
or ( \1631_b1 , \1629_b1 , w_3481 );
not ( w_3481 , w_3482 );
and ( \1631_b0 , \1629_b0 , w_3483 );
and ( w_3482 ,  , w_3483 );
buf ( w_3481 , \1630_b1 );
not ( w_3481 , w_3484 );
not (  , w_3485 );
and ( w_3484 , w_3485 , \1630_b0 );
or ( \1632_b1 , \1631_b1 , w_3486 );
xor ( \1632_b0 , \1631_b0 , w_3488 );
not ( w_3488 , w_3489 );
and ( w_3489 , w_3486 , w_3487 );
buf ( w_3486 , \818_b1 );
not ( w_3486 , w_3490 );
not ( w_3487 , w_3491 );
and ( w_3490 , w_3491 , \818_b0 );
or ( \1633_b1 , \1628_b1 , \1632_b1 );
not ( \1632_b1 , w_3492 );
and ( \1633_b0 , \1628_b0 , w_3493 );
and ( w_3492 , w_3493 , \1632_b0 );
or ( \1634_b1 , \495_b1 , \740_b1 );
not ( \740_b1 , w_3494 );
and ( \1634_b0 , \495_b0 , w_3495 );
and ( w_3494 , w_3495 , \740_b0 );
or ( \1635_b1 , \444_b1 , \738_b1 );
not ( \738_b1 , w_3496 );
and ( \1635_b0 , \444_b0 , w_3497 );
and ( w_3496 , w_3497 , \738_b0 );
or ( \1636_b1 , \1634_b1 , w_3499 );
not ( w_3499 , w_3500 );
and ( \1636_b0 , \1634_b0 , w_3501 );
and ( w_3500 ,  , w_3501 );
buf ( w_3499 , \1635_b1 );
not ( w_3499 , w_3502 );
not (  , w_3503 );
and ( w_3502 , w_3503 , \1635_b0 );
or ( \1637_b1 , \1636_b1 , w_3504 );
xor ( \1637_b0 , \1636_b0 , w_3506 );
not ( w_3506 , w_3507 );
and ( w_3507 , w_3504 , w_3505 );
buf ( w_3504 , \668_b1 );
not ( w_3504 , w_3508 );
not ( w_3505 , w_3509 );
and ( w_3508 , w_3509 , \668_b0 );
or ( \1638_b1 , \1632_b1 , \1637_b1 );
not ( \1637_b1 , w_3510 );
and ( \1638_b0 , \1632_b0 , w_3511 );
and ( w_3510 , w_3511 , \1637_b0 );
or ( \1639_b1 , \1628_b1 , \1637_b1 );
not ( \1637_b1 , w_3512 );
and ( \1639_b0 , \1628_b0 , w_3513 );
and ( w_3512 , w_3513 , \1637_b0 );
or ( \1641_b1 , \1623_b1 , \1640_b1 );
not ( \1640_b1 , w_3514 );
and ( \1641_b0 , \1623_b0 , w_3515 );
and ( w_3514 , w_3515 , \1640_b0 );
or ( \1642_b1 , \1603_b1 , \1640_b1 );
not ( \1640_b1 , w_3516 );
and ( \1642_b0 , \1603_b0 , w_3517 );
and ( w_3516 , w_3517 , \1640_b0 );
or ( \1644_b1 , \1479_b1 , \1483_b1 );
xor ( \1644_b0 , \1479_b0 , w_3518 );
not ( w_3518 , w_3519 );
and ( w_3519 , \1483_b1 , \1483_b0 );
or ( \1645_b1 , \1644_b1 , \1488_b1 );
xor ( \1645_b0 , \1644_b0 , w_3520 );
not ( w_3520 , w_3521 );
and ( w_3521 , \1488_b1 , \1488_b0 );
or ( \1646_b1 , \1495_b1 , \1499_b1 );
xor ( \1646_b0 , \1495_b0 , w_3522 );
not ( w_3522 , w_3523 );
and ( w_3523 , \1499_b1 , \1499_b0 );
or ( \1647_b1 , \1646_b1 , \1504_b1 );
xor ( \1647_b0 , \1646_b0 , w_3524 );
not ( w_3524 , w_3525 );
and ( w_3525 , \1504_b1 , \1504_b0 );
or ( \1648_b1 , \1645_b1 , \1647_b1 );
not ( \1647_b1 , w_3526 );
and ( \1648_b0 , \1645_b0 , w_3527 );
and ( w_3526 , w_3527 , \1647_b0 );
or ( \1649_b1 , \1512_b1 , \1516_b1 );
xor ( \1649_b0 , \1512_b0 , w_3528 );
not ( w_3528 , w_3529 );
and ( w_3529 , \1516_b1 , \1516_b0 );
or ( \1650_b1 , \1649_b1 , \1521_b1 );
xor ( \1650_b0 , \1649_b0 , w_3530 );
not ( w_3530 , w_3531 );
and ( w_3531 , \1521_b1 , \1521_b0 );
or ( \1651_b1 , \1647_b1 , \1650_b1 );
not ( \1650_b1 , w_3532 );
and ( \1651_b0 , \1647_b0 , w_3533 );
and ( w_3532 , w_3533 , \1650_b0 );
or ( \1652_b1 , \1645_b1 , \1650_b1 );
not ( \1650_b1 , w_3534 );
and ( \1652_b0 , \1645_b0 , w_3535 );
and ( w_3534 , w_3535 , \1650_b0 );
or ( \1654_b1 , \1643_b1 , \1653_b1 );
not ( \1653_b1 , w_3536 );
and ( \1654_b0 , \1643_b0 , w_3537 );
and ( w_3536 , w_3537 , \1653_b0 );
or ( \1655_b1 , \1194_b1 , \313_b1 );
not ( \313_b1 , w_3538 );
and ( \1655_b0 , \1194_b0 , w_3539 );
and ( w_3538 , w_3539 , \313_b0 );
or ( \1656_b1 , \1104_b1 , \311_b1 );
not ( \311_b1 , w_3540 );
and ( \1656_b0 , \1104_b0 , w_3541 );
and ( w_3540 , w_3541 , \311_b0 );
or ( \1657_b1 , \1655_b1 , w_3543 );
not ( w_3543 , w_3544 );
and ( \1657_b0 , \1655_b0 , w_3545 );
and ( w_3544 ,  , w_3545 );
buf ( w_3543 , \1656_b1 );
not ( w_3543 , w_3546 );
not (  , w_3547 );
and ( w_3546 , w_3547 , \1656_b0 );
or ( \1658_b1 , \1657_b1 , w_3548 );
xor ( \1658_b0 , \1657_b0 , w_3550 );
not ( w_3550 , w_3551 );
and ( w_3551 , w_3548 , w_3549 );
buf ( w_3548 , \320_b1 );
not ( w_3548 , w_3552 );
not ( w_3549 , w_3553 );
and ( w_3552 , w_3553 , \320_b0 );
or ( \1659_b1 , \1304_b1 , \331_b1 );
not ( \331_b1 , w_3554 );
and ( \1659_b0 , \1304_b0 , w_3555 );
and ( w_3554 , w_3555 , \331_b0 );
or ( \1660_b1 , \1299_b1 , \329_b1 );
not ( \329_b1 , w_3556 );
and ( \1660_b0 , \1299_b0 , w_3557 );
and ( w_3556 , w_3557 , \329_b0 );
or ( \1661_b1 , \1659_b1 , w_3559 );
not ( w_3559 , w_3560 );
and ( \1661_b0 , \1659_b0 , w_3561 );
and ( w_3560 ,  , w_3561 );
buf ( w_3559 , \1660_b1 );
not ( w_3559 , w_3562 );
not (  , w_3563 );
and ( w_3562 , w_3563 , \1660_b0 );
or ( \1662_b1 , \1661_b1 , w_3564 );
xor ( \1662_b0 , \1661_b0 , w_3566 );
not ( w_3566 , w_3567 );
and ( w_3567 , w_3564 , w_3565 );
buf ( w_3564 , \338_b1 );
not ( w_3564 , w_3568 );
not ( w_3565 , w_3569 );
and ( w_3568 , w_3569 , \338_b0 );
or ( \1663_b1 , \1658_b1 , \1662_b1 );
not ( \1662_b1 , w_3570 );
and ( \1663_b0 , \1658_b0 , w_3571 );
and ( w_3570 , w_3571 , \1662_b0 );
or ( \1664_b1 , \1537_b1 , \351_b1 );
not ( \351_b1 , w_3572 );
and ( \1664_b0 , \1537_b0 , w_3573 );
and ( w_3572 , w_3573 , \351_b0 );
or ( \1665_b1 , \1422_b1 , \349_b1 );
not ( \349_b1 , w_3574 );
and ( \1665_b0 , \1422_b0 , w_3575 );
and ( w_3574 , w_3575 , \349_b0 );
or ( \1666_b1 , \1664_b1 , w_3577 );
not ( w_3577 , w_3578 );
and ( \1666_b0 , \1664_b0 , w_3579 );
and ( w_3578 ,  , w_3579 );
buf ( w_3577 , \1665_b1 );
not ( w_3577 , w_3580 );
not (  , w_3581 );
and ( w_3580 , w_3581 , \1665_b0 );
or ( \1667_b1 , \1666_b1 , w_3582 );
xor ( \1667_b0 , \1666_b0 , w_3584 );
not ( w_3584 , w_3585 );
and ( w_3585 , w_3582 , w_3583 );
buf ( w_3582 , \358_b1 );
not ( w_3582 , w_3586 );
not ( w_3583 , w_3587 );
and ( w_3586 , w_3587 , \358_b0 );
or ( \1668_b1 , \1662_b1 , \1667_b1 );
not ( \1667_b1 , w_3588 );
and ( \1668_b0 , \1662_b0 , w_3589 );
and ( w_3588 , w_3589 , \1667_b0 );
or ( \1669_b1 , \1658_b1 , \1667_b1 );
not ( \1667_b1 , w_3590 );
and ( \1669_b0 , \1658_b0 , w_3591 );
and ( w_3590 , w_3591 , \1667_b0 );
or ( \1671_b1 , \1531_b1 , \1535_b1 );
xor ( \1671_b0 , \1531_b0 , w_3592 );
not ( w_3592 , w_3593 );
and ( w_3593 , \1535_b1 , \1535_b0 );
or ( \1672_b1 , \1671_b1 , \1538_b1 );
xor ( \1672_b0 , \1671_b0 , w_3594 );
not ( w_3594 , w_3595 );
and ( w_3595 , \1538_b1 , \1538_b0 );
or ( \1673_b1 , \1670_b1 , w_3596 );
or ( \1673_b0 , \1670_b0 , \1672_b0 );
not ( \1672_b0 , w_3597 );
and ( w_3597 , w_3596 , \1672_b1 );
or ( \1674_b1 , \1653_b1 , \1673_b1 );
not ( \1673_b1 , w_3598 );
and ( \1674_b0 , \1653_b0 , w_3599 );
and ( w_3598 , w_3599 , \1673_b0 );
or ( \1675_b1 , \1643_b1 , \1673_b1 );
not ( \1673_b1 , w_3600 );
and ( \1675_b0 , \1643_b0 , w_3601 );
and ( w_3600 , w_3601 , \1673_b0 );
or ( \1677_b1 , \1491_b1 , \1507_b1 );
xor ( \1677_b0 , \1491_b0 , w_3602 );
not ( w_3602 , w_3603 );
and ( w_3603 , \1507_b1 , \1507_b0 );
or ( \1678_b1 , \1677_b1 , \1524_b1 );
xor ( \1678_b0 , \1677_b0 , w_3604 );
not ( w_3604 , w_3605 );
and ( w_3605 , \1524_b1 , \1524_b0 );
or ( \1679_b1 , \1541_b1 , \1543_b1 );
xor ( \1679_b0 , \1541_b0 , w_3606 );
not ( w_3606 , w_3607 );
and ( w_3607 , \1543_b1 , \1543_b0 );
or ( \1680_b1 , \1679_b1 , \1546_b1 );
xor ( \1680_b0 , \1679_b0 , w_3608 );
not ( w_3608 , w_3609 );
and ( w_3609 , \1546_b1 , \1546_b0 );
or ( \1681_b1 , \1678_b1 , \1680_b1 );
not ( \1680_b1 , w_3610 );
and ( \1681_b0 , \1678_b0 , w_3611 );
and ( w_3610 , w_3611 , \1680_b0 );
or ( \1682_b1 , \1552_b1 , \1554_b1 );
xor ( \1682_b0 , \1552_b0 , w_3612 );
not ( w_3612 , w_3613 );
and ( w_3613 , \1554_b1 , \1554_b0 );
or ( \1683_b1 , \1680_b1 , \1682_b1 );
not ( \1682_b1 , w_3614 );
and ( \1683_b0 , \1680_b0 , w_3615 );
and ( w_3614 , w_3615 , \1682_b0 );
or ( \1684_b1 , \1678_b1 , \1682_b1 );
not ( \1682_b1 , w_3616 );
and ( \1684_b0 , \1678_b0 , w_3617 );
and ( w_3616 , w_3617 , \1682_b0 );
or ( \1686_b1 , \1676_b1 , \1685_b1 );
not ( \1685_b1 , w_3618 );
and ( \1686_b0 , \1676_b0 , w_3619 );
and ( w_3618 , w_3619 , \1685_b0 );
or ( \1687_b1 , \1560_b1 , \1562_b1 );
xor ( \1687_b0 , \1560_b0 , w_3620 );
not ( w_3620 , w_3621 );
and ( w_3621 , \1562_b1 , \1562_b0 );
or ( \1688_b1 , \1687_b1 , \1564_b1 );
xor ( \1688_b0 , \1687_b0 , w_3622 );
not ( w_3622 , w_3623 );
and ( w_3623 , \1564_b1 , \1564_b0 );
or ( \1689_b1 , \1685_b1 , \1688_b1 );
not ( \1688_b1 , w_3624 );
and ( \1689_b0 , \1685_b0 , w_3625 );
and ( w_3624 , w_3625 , \1688_b0 );
or ( \1690_b1 , \1676_b1 , \1688_b1 );
not ( \1688_b1 , w_3626 );
and ( \1690_b0 , \1676_b0 , w_3627 );
and ( w_3626 , w_3627 , \1688_b0 );
or ( \1692_b1 , \1412_b1 , \1433_b1 );
xor ( \1692_b0 , \1412_b0 , w_3628 );
not ( w_3628 , w_3629 );
and ( w_3629 , \1433_b1 , \1433_b0 );
or ( \1693_b1 , \1692_b1 , \1439_b1 );
xor ( \1693_b0 , \1692_b0 , w_3630 );
not ( w_3630 , w_3631 );
and ( w_3631 , \1439_b1 , \1439_b0 );
or ( \1694_b1 , \1691_b1 , \1693_b1 );
not ( \1693_b1 , w_3632 );
and ( \1694_b0 , \1691_b0 , w_3633 );
and ( w_3632 , w_3633 , \1693_b0 );
or ( \1695_b1 , \1558_b1 , \1567_b1 );
xor ( \1695_b0 , \1558_b0 , w_3634 );
not ( w_3634 , w_3635 );
and ( w_3635 , \1567_b1 , \1567_b0 );
or ( \1696_b1 , \1695_b1 , \1570_b1 );
xor ( \1696_b0 , \1695_b0 , w_3636 );
not ( w_3636 , w_3637 );
and ( w_3637 , \1570_b1 , \1570_b0 );
or ( \1697_b1 , \1693_b1 , \1696_b1 );
not ( \1696_b1 , w_3638 );
and ( \1697_b0 , \1693_b0 , w_3639 );
and ( w_3638 , w_3639 , \1696_b0 );
or ( \1698_b1 , \1691_b1 , \1696_b1 );
not ( \1696_b1 , w_3640 );
and ( \1698_b0 , \1691_b0 , w_3641 );
and ( w_3640 , w_3641 , \1696_b0 );
or ( \1700_b1 , \1573_b1 , \1575_b1 );
xor ( \1700_b0 , \1573_b0 , w_3642 );
not ( w_3642 , w_3643 );
and ( w_3643 , \1575_b1 , \1575_b0 );
or ( \1701_b1 , \1700_b1 , \1578_b1 );
xor ( \1701_b0 , \1700_b0 , w_3644 );
not ( w_3644 , w_3645 );
and ( w_3645 , \1578_b1 , \1578_b0 );
or ( \1702_b1 , \1699_b1 , \1701_b1 );
not ( \1701_b1 , w_3646 );
and ( \1702_b0 , \1699_b0 , w_3647 );
and ( w_3646 , w_3647 , \1701_b0 );
or ( \1703_b1 , \1587_b1 , \1702_b1 );
not ( \1702_b1 , w_3648 );
and ( \1703_b0 , \1587_b0 , w_3649 );
and ( w_3648 , w_3649 , \1702_b0 );
or ( \1704_b1 , \1587_b1 , \1702_b1 );
xor ( \1704_b0 , \1587_b0 , w_3650 );
not ( w_3650 , w_3651 );
and ( w_3651 , \1702_b1 , \1702_b0 );
or ( \1705_b1 , \1699_b1 , \1701_b1 );
xor ( \1705_b0 , \1699_b0 , w_3652 );
not ( w_3652 , w_3653 );
and ( w_3653 , \1701_b1 , \1701_b0 );
or ( \1706_b1 , \703_b1 , \604_b1 );
not ( \604_b1 , w_3654 );
and ( \1706_b0 , \703_b0 , w_3655 );
and ( w_3654 , w_3655 , \604_b0 );
or ( \1707_b1 , \621_b1 , \602_b1 );
not ( \602_b1 , w_3656 );
and ( \1707_b0 , \621_b0 , w_3657 );
and ( w_3656 , w_3657 , \602_b0 );
or ( \1708_b1 , \1706_b1 , w_3659 );
not ( w_3659 , w_3660 );
and ( \1708_b0 , \1706_b0 , w_3661 );
and ( w_3660 ,  , w_3661 );
buf ( w_3659 , \1707_b1 );
not ( w_3659 , w_3662 );
not (  , w_3663 );
and ( w_3662 , w_3663 , \1707_b0 );
or ( \1709_b1 , \1708_b1 , w_3664 );
xor ( \1709_b0 , \1708_b0 , w_3666 );
not ( w_3666 , w_3667 );
and ( w_3667 , w_3664 , w_3665 );
buf ( w_3664 , \561_b1 );
not ( w_3664 , w_3668 );
not ( w_3665 , w_3669 );
and ( w_3668 , w_3669 , \561_b0 );
or ( \1710_b1 , \841_b1 , \503_b1 );
not ( \503_b1 , w_3670 );
and ( \1710_b0 , \841_b0 , w_3671 );
and ( w_3670 , w_3671 , \503_b0 );
or ( \1711_b1 , \777_b1 , \501_b1 );
not ( \501_b1 , w_3672 );
and ( \1711_b0 , \777_b0 , w_3673 );
and ( w_3672 , w_3673 , \501_b0 );
or ( \1712_b1 , \1710_b1 , w_3675 );
not ( w_3675 , w_3676 );
and ( \1712_b0 , \1710_b0 , w_3677 );
and ( w_3676 ,  , w_3677 );
buf ( w_3675 , \1711_b1 );
not ( w_3675 , w_3678 );
not (  , w_3679 );
and ( w_3678 , w_3679 , \1711_b0 );
or ( \1713_b1 , \1712_b1 , w_3680 );
xor ( \1713_b0 , \1712_b0 , w_3682 );
not ( w_3682 , w_3683 );
and ( w_3683 , w_3680 , w_3681 );
buf ( w_3680 , \455_b1 );
not ( w_3680 , w_3684 );
not ( w_3681 , w_3685 );
and ( w_3684 , w_3685 , \455_b0 );
or ( \1714_b1 , \1709_b1 , \1713_b1 );
not ( \1713_b1 , w_3686 );
and ( \1714_b0 , \1709_b0 , w_3687 );
and ( w_3686 , w_3687 , \1713_b0 );
or ( \1715_b1 , \1104_b1 , \298_b1 );
not ( \298_b1 , w_3688 );
and ( \1715_b0 , \1104_b0 , w_3689 );
and ( w_3688 , w_3689 , \298_b0 );
or ( \1716_b1 , \904_b1 , \296_b1 );
not ( \296_b1 , w_3690 );
and ( \1716_b0 , \904_b0 , w_3691 );
and ( w_3690 , w_3691 , \296_b0 );
or ( \1717_b1 , \1715_b1 , w_3693 );
not ( w_3693 , w_3694 );
and ( \1717_b0 , \1715_b0 , w_3695 );
and ( w_3694 ,  , w_3695 );
buf ( w_3693 , \1716_b1 );
not ( w_3693 , w_3696 );
not (  , w_3697 );
and ( w_3696 , w_3697 , \1716_b0 );
or ( \1718_b1 , \1717_b1 , w_3698 );
xor ( \1718_b0 , \1717_b0 , w_3700 );
not ( w_3700 , w_3701 );
and ( w_3701 , w_3698 , w_3699 );
buf ( w_3698 , \303_b1 );
not ( w_3698 , w_3702 );
not ( w_3699 , w_3703 );
and ( w_3702 , w_3703 , \303_b0 );
or ( \1719_b1 , \1713_b1 , \1718_b1 );
not ( \1718_b1 , w_3704 );
and ( \1719_b0 , \1713_b0 , w_3705 );
and ( w_3704 , w_3705 , \1718_b0 );
or ( \1720_b1 , \1709_b1 , \1718_b1 );
not ( \1718_b1 , w_3706 );
and ( \1720_b0 , \1709_b0 , w_3707 );
and ( w_3706 , w_3707 , \1718_b0 );
or ( \1722_b1 , \343_b1 , \1062_b1 );
not ( \1062_b1 , w_3708 );
and ( \1722_b0 , \343_b0 , w_3709 );
and ( w_3708 , w_3709 , \1062_b0 );
or ( \1723_b1 , \353_b1 , \1060_b1 );
not ( \1060_b1 , w_3710 );
and ( \1723_b0 , \353_b0 , w_3711 );
and ( w_3710 , w_3711 , \1060_b0 );
or ( \1724_b1 , \1722_b1 , w_3713 );
not ( w_3713 , w_3714 );
and ( \1724_b0 , \1722_b0 , w_3715 );
and ( w_3714 ,  , w_3715 );
buf ( w_3713 , \1723_b1 );
not ( w_3713 , w_3716 );
not (  , w_3717 );
and ( w_3716 , w_3717 , \1723_b0 );
or ( \1725_b1 , \1724_b1 , w_3718 );
xor ( \1725_b0 , \1724_b0 , w_3720 );
not ( w_3720 , w_3721 );
and ( w_3721 , w_3718 , w_3719 );
buf ( w_3718 , \984_b1 );
not ( w_3718 , w_3722 );
not ( w_3719 , w_3723 );
and ( w_3722 , w_3723 , \984_b0 );
or ( \1726_b1 , \444_b1 , \912_b1 );
not ( \912_b1 , w_3724 );
and ( \1726_b0 , \444_b0 , w_3725 );
and ( w_3724 , w_3725 , \912_b0 );
or ( \1727_b1 , \360_b1 , \910_b1 );
not ( \910_b1 , w_3726 );
and ( \1727_b0 , \360_b0 , w_3727 );
and ( w_3726 , w_3727 , \910_b0 );
or ( \1728_b1 , \1726_b1 , w_3729 );
not ( w_3729 , w_3730 );
and ( \1728_b0 , \1726_b0 , w_3731 );
and ( w_3730 ,  , w_3731 );
buf ( w_3729 , \1727_b1 );
not ( w_3729 , w_3732 );
not (  , w_3733 );
and ( w_3732 , w_3733 , \1727_b0 );
or ( \1729_b1 , \1728_b1 , w_3734 );
xor ( \1729_b0 , \1728_b0 , w_3736 );
not ( w_3736 , w_3737 );
and ( w_3737 , w_3734 , w_3735 );
buf ( w_3734 , \818_b1 );
not ( w_3734 , w_3738 );
not ( w_3735 , w_3739 );
and ( w_3738 , w_3739 , \818_b0 );
or ( \1730_b1 , \1725_b1 , \1729_b1 );
not ( \1729_b1 , w_3740 );
and ( \1730_b0 , \1725_b0 , w_3741 );
and ( w_3740 , w_3741 , \1729_b0 );
or ( \1731_b1 , \593_b1 , \740_b1 );
not ( \740_b1 , w_3742 );
and ( \1731_b0 , \593_b0 , w_3743 );
and ( w_3742 , w_3743 , \740_b0 );
or ( \1732_b1 , \495_b1 , \738_b1 );
not ( \738_b1 , w_3744 );
and ( \1732_b0 , \495_b0 , w_3745 );
and ( w_3744 , w_3745 , \738_b0 );
or ( \1733_b1 , \1731_b1 , w_3747 );
not ( w_3747 , w_3748 );
and ( \1733_b0 , \1731_b0 , w_3749 );
and ( w_3748 ,  , w_3749 );
buf ( w_3747 , \1732_b1 );
not ( w_3747 , w_3750 );
not (  , w_3751 );
and ( w_3750 , w_3751 , \1732_b0 );
or ( \1734_b1 , \1733_b1 , w_3752 );
xor ( \1734_b0 , \1733_b0 , w_3754 );
not ( w_3754 , w_3755 );
and ( w_3755 , w_3752 , w_3753 );
buf ( w_3752 , \668_b1 );
not ( w_3752 , w_3756 );
not ( w_3753 , w_3757 );
and ( w_3756 , w_3757 , \668_b0 );
or ( \1735_b1 , \1729_b1 , \1734_b1 );
not ( \1734_b1 , w_3758 );
and ( \1735_b0 , \1729_b0 , w_3759 );
and ( w_3758 , w_3759 , \1734_b0 );
or ( \1736_b1 , \1725_b1 , \1734_b1 );
not ( \1734_b1 , w_3760 );
and ( \1736_b0 , \1725_b0 , w_3761 );
and ( w_3760 , w_3761 , \1734_b0 );
or ( \1738_b1 , \1721_b1 , \1737_b1 );
not ( \1737_b1 , w_3762 );
and ( \1738_b0 , \1721_b0 , w_3763 );
and ( w_3762 , w_3763 , \1737_b0 );
or ( \1739_b1 , \1360_b1 , \1605_b1 );
xor ( \1739_b0 , \1360_b0 , w_3764 );
not ( w_3764 , w_3765 );
and ( w_3765 , \1605_b1 , \1605_b0 );
or ( \1740_b1 , \1605_b1 , \1607_b1 );
xor ( \1740_b0 , \1605_b0 , w_3766 );
not ( w_3766 , w_3767 );
and ( w_3767 , \1607_b1 , \1607_b0 );
buf ( \1741_b1 , \1740_b1 );
not ( \1741_b1 , w_3768 );
not ( \1741_b0 , w_3769 );
and ( w_3768 , w_3769 , \1740_b0 );
or ( \1742_b1 , \1739_b1 , \1741_b1 );
not ( \1741_b1 , w_3770 );
and ( \1742_b0 , \1739_b0 , w_3771 );
and ( w_3770 , w_3771 , \1741_b0 );
or ( \1743_b1 , \159_b1 , \1742_b1 );
not ( \1742_b1 , w_3772 );
and ( \1743_b0 , \159_b0 , w_3773 );
and ( w_3772 , w_3773 , \1742_b0 );
buf ( \1744_b1 , \1743_b1 );
not ( \1744_b1 , w_3774 );
not ( \1744_b0 , w_3775 );
and ( w_3774 , w_3775 , \1743_b0 );
or ( \1745_b1 , \1744_b1 , w_3776 );
xor ( \1745_b0 , \1744_b0 , w_3778 );
not ( w_3778 , w_3779 );
and ( w_3779 , w_3776 , w_3777 );
buf ( w_3776 , \1610_b1 );
not ( w_3776 , w_3780 );
not ( w_3777 , w_3781 );
and ( w_3780 , w_3781 , \1610_b0 );
or ( \1746_b1 , \305_b1 , \1476_b1 );
not ( \1476_b1 , w_3782 );
and ( \1746_b0 , \305_b0 , w_3783 );
and ( w_3782 , w_3783 , \1476_b0 );
or ( \1747_b1 , \315_b1 , \1474_b1 );
not ( \1474_b1 , w_3784 );
and ( \1747_b0 , \315_b0 , w_3785 );
and ( w_3784 , w_3785 , \1474_b0 );
or ( \1748_b1 , \1746_b1 , w_3787 );
not ( w_3787 , w_3788 );
and ( \1748_b0 , \1746_b0 , w_3789 );
and ( w_3788 ,  , w_3789 );
buf ( w_3787 , \1747_b1 );
not ( w_3787 , w_3790 );
not (  , w_3791 );
and ( w_3790 , w_3791 , \1747_b0 );
or ( \1749_b1 , \1748_b1 , w_3792 );
xor ( \1749_b0 , \1748_b0 , w_3794 );
not ( w_3794 , w_3795 );
and ( w_3795 , w_3792 , w_3793 );
buf ( w_3792 , \1363_b1 );
not ( w_3792 , w_3796 );
not ( w_3793 , w_3797 );
and ( w_3796 , w_3797 , \1363_b0 );
or ( \1750_b1 , \1745_b1 , \1749_b1 );
not ( \1749_b1 , w_3798 );
and ( \1750_b0 , \1745_b0 , w_3799 );
and ( w_3798 , w_3799 , \1749_b0 );
or ( \1751_b1 , \323_b1 , \1280_b1 );
not ( \1280_b1 , w_3800 );
and ( \1751_b0 , \323_b0 , w_3801 );
and ( w_3800 , w_3801 , \1280_b0 );
or ( \1752_b1 , \333_b1 , \1278_b1 );
not ( \1278_b1 , w_3802 );
and ( \1752_b0 , \333_b0 , w_3803 );
and ( w_3802 , w_3803 , \1278_b0 );
or ( \1753_b1 , \1751_b1 , w_3805 );
not ( w_3805 , w_3806 );
and ( \1753_b0 , \1751_b0 , w_3807 );
and ( w_3806 ,  , w_3807 );
buf ( w_3805 , \1752_b1 );
not ( w_3805 , w_3808 );
not (  , w_3809 );
and ( w_3808 , w_3809 , \1752_b0 );
or ( \1754_b1 , \1753_b1 , w_3810 );
xor ( \1754_b0 , \1753_b0 , w_3812 );
not ( w_3812 , w_3813 );
and ( w_3813 , w_3810 , w_3811 );
buf ( w_3810 , \1177_b1 );
not ( w_3810 , w_3814 );
not ( w_3811 , w_3815 );
and ( w_3814 , w_3815 , \1177_b0 );
or ( \1755_b1 , \1749_b1 , \1754_b1 );
not ( \1754_b1 , w_3816 );
and ( \1755_b0 , \1749_b0 , w_3817 );
and ( w_3816 , w_3817 , \1754_b0 );
or ( \1756_b1 , \1745_b1 , \1754_b1 );
not ( \1754_b1 , w_3818 );
and ( \1756_b0 , \1745_b0 , w_3819 );
and ( w_3818 , w_3819 , \1754_b0 );
or ( \1758_b1 , \1737_b1 , \1757_b1 );
not ( \1757_b1 , w_3820 );
and ( \1758_b0 , \1737_b0 , w_3821 );
and ( w_3820 , w_3821 , \1757_b0 );
or ( \1759_b1 , \1721_b1 , \1757_b1 );
not ( \1757_b1 , w_3822 );
and ( \1759_b0 , \1721_b0 , w_3823 );
and ( w_3822 , w_3823 , \1757_b0 );
or ( \1761_b1 , \1299_b1 , \313_b1 );
not ( \313_b1 , w_3824 );
and ( \1761_b0 , \1299_b0 , w_3825 );
and ( w_3824 , w_3825 , \313_b0 );
or ( \1762_b1 , \1194_b1 , \311_b1 );
not ( \311_b1 , w_3826 );
and ( \1762_b0 , \1194_b0 , w_3827 );
and ( w_3826 , w_3827 , \311_b0 );
or ( \1763_b1 , \1761_b1 , w_3829 );
not ( w_3829 , w_3830 );
and ( \1763_b0 , \1761_b0 , w_3831 );
and ( w_3830 ,  , w_3831 );
buf ( w_3829 , \1762_b1 );
not ( w_3829 , w_3832 );
not (  , w_3833 );
and ( w_3832 , w_3833 , \1762_b0 );
or ( \1764_b1 , \1763_b1 , w_3834 );
xor ( \1764_b0 , \1763_b0 , w_3836 );
not ( w_3836 , w_3837 );
and ( w_3837 , w_3834 , w_3835 );
buf ( w_3834 , \320_b1 );
not ( w_3834 , w_3838 );
not ( w_3835 , w_3839 );
and ( w_3838 , w_3839 , \320_b0 );
or ( \1765_b1 , \1422_b1 , \331_b1 );
not ( \331_b1 , w_3840 );
and ( \1765_b0 , \1422_b0 , w_3841 );
and ( w_3840 , w_3841 , \331_b0 );
or ( \1766_b1 , \1304_b1 , \329_b1 );
not ( \329_b1 , w_3842 );
and ( \1766_b0 , \1304_b0 , w_3843 );
and ( w_3842 , w_3843 , \329_b0 );
or ( \1767_b1 , \1765_b1 , w_3845 );
not ( w_3845 , w_3846 );
and ( \1767_b0 , \1765_b0 , w_3847 );
and ( w_3846 ,  , w_3847 );
buf ( w_3845 , \1766_b1 );
not ( w_3845 , w_3848 );
not (  , w_3849 );
and ( w_3848 , w_3849 , \1766_b0 );
or ( \1768_b1 , \1767_b1 , w_3850 );
xor ( \1768_b0 , \1767_b0 , w_3852 );
not ( w_3852 , w_3853 );
and ( w_3853 , w_3850 , w_3851 );
buf ( w_3850 , \338_b1 );
not ( w_3850 , w_3854 );
not ( w_3851 , w_3855 );
and ( w_3854 , w_3855 , \338_b0 );
or ( \1769_b1 , \1764_b1 , \1768_b1 );
not ( \1768_b1 , w_3856 );
and ( \1769_b0 , \1764_b0 , w_3857 );
and ( w_3856 , w_3857 , \1768_b0 );
buf ( \1770_b1 , RIb4befe8_87_b1 );
buf ( \1770_b0 , RIb4befe8_87_b0 );
or ( \1771_b1 , \1770_b1 , \351_b1 );
not ( \351_b1 , w_3858 );
and ( \1771_b0 , \1770_b0 , w_3859 );
and ( w_3858 , w_3859 , \351_b0 );
or ( \1772_b1 , \1537_b1 , \349_b1 );
not ( \349_b1 , w_3860 );
and ( \1772_b0 , \1537_b0 , w_3861 );
and ( w_3860 , w_3861 , \349_b0 );
or ( \1773_b1 , \1771_b1 , w_3863 );
not ( w_3863 , w_3864 );
and ( \1773_b0 , \1771_b0 , w_3865 );
and ( w_3864 ,  , w_3865 );
buf ( w_3863 , \1772_b1 );
not ( w_3863 , w_3866 );
not (  , w_3867 );
and ( w_3866 , w_3867 , \1772_b0 );
or ( \1774_b1 , \1773_b1 , w_3868 );
xor ( \1774_b0 , \1773_b0 , w_3870 );
not ( w_3870 , w_3871 );
and ( w_3871 , w_3868 , w_3869 );
buf ( w_3868 , \358_b1 );
not ( w_3868 , w_3872 );
not ( w_3869 , w_3873 );
and ( w_3872 , w_3873 , \358_b0 );
or ( \1775_b1 , \1768_b1 , \1774_b1 );
not ( \1774_b1 , w_3874 );
and ( \1775_b0 , \1768_b0 , w_3875 );
and ( w_3874 , w_3875 , \1774_b0 );
or ( \1776_b1 , \1764_b1 , \1774_b1 );
not ( \1774_b1 , w_3876 );
and ( \1776_b0 , \1764_b0 , w_3877 );
and ( w_3876 , w_3877 , \1774_b0 );
buf ( \1778_b1 , RIb4bef70_88_b1 );
buf ( \1778_b0 , RIb4bef70_88_b0 );
or ( \1779_b1 , \1778_b1 , \345_b1 );
not ( \345_b1 , w_3878 );
and ( \1779_b0 , \1778_b0 , w_3879 );
and ( w_3878 , w_3879 , \345_b0 );
buf ( \1780_b1 , \1779_b1 );
buf ( \1780_b0 , \1779_b0 );
or ( \1781_b1 , \1777_b1 , \1780_b1 );
not ( \1780_b1 , w_3880 );
and ( \1781_b0 , \1777_b0 , w_3881 );
and ( w_3880 , w_3881 , \1780_b0 );
or ( \1782_b1 , \1770_b1 , \345_b1 );
not ( \345_b1 , w_3882 );
and ( \1782_b0 , \1770_b0 , w_3883 );
and ( w_3882 , w_3883 , \345_b0 );
or ( \1783_b1 , \1780_b1 , \1782_b1 );
not ( \1782_b1 , w_3884 );
and ( \1783_b0 , \1780_b0 , w_3885 );
and ( w_3884 , w_3885 , \1782_b0 );
or ( \1784_b1 , \1777_b1 , \1782_b1 );
not ( \1782_b1 , w_3886 );
and ( \1784_b0 , \1777_b0 , w_3887 );
and ( w_3886 , w_3887 , \1782_b0 );
or ( \1786_b1 , \1760_b1 , \1785_b1 );
not ( \1785_b1 , w_3888 );
and ( \1786_b0 , \1760_b0 , w_3889 );
and ( w_3888 , w_3889 , \1785_b0 );
or ( \1787_b1 , \1658_b1 , \1662_b1 );
xor ( \1787_b0 , \1658_b0 , w_3890 );
not ( w_3890 , w_3891 );
and ( w_3891 , \1662_b1 , \1662_b0 );
or ( \1788_b1 , \1787_b1 , \1667_b1 );
xor ( \1788_b0 , \1787_b0 , w_3892 );
not ( w_3892 , w_3893 );
and ( w_3893 , \1667_b1 , \1667_b0 );
or ( \1789_b1 , \1591_b1 , \1595_b1 );
xor ( \1789_b0 , \1591_b0 , w_3894 );
not ( w_3894 , w_3895 );
and ( w_3895 , \1595_b1 , \1595_b0 );
or ( \1790_b1 , \1789_b1 , \1600_b1 );
xor ( \1790_b0 , \1789_b0 , w_3896 );
not ( w_3896 , w_3897 );
and ( w_3897 , \1600_b1 , \1600_b0 );
or ( \1791_b1 , \1788_b1 , \1790_b1 );
not ( \1790_b1 , w_3898 );
and ( \1791_b0 , \1788_b0 , w_3899 );
and ( w_3898 , w_3899 , \1790_b0 );
or ( \1792_b1 , \1628_b1 , \1632_b1 );
xor ( \1792_b0 , \1628_b0 , w_3900 );
not ( w_3900 , w_3901 );
and ( w_3901 , \1632_b1 , \1632_b0 );
or ( \1793_b1 , \1792_b1 , \1637_b1 );
xor ( \1793_b0 , \1792_b0 , w_3902 );
not ( w_3902 , w_3903 );
and ( w_3903 , \1637_b1 , \1637_b0 );
or ( \1794_b1 , \1790_b1 , \1793_b1 );
not ( \1793_b1 , w_3904 );
and ( \1794_b0 , \1790_b0 , w_3905 );
and ( w_3904 , w_3905 , \1793_b0 );
or ( \1795_b1 , \1788_b1 , \1793_b1 );
not ( \1793_b1 , w_3906 );
and ( \1795_b0 , \1788_b0 , w_3907 );
and ( w_3906 , w_3907 , \1793_b0 );
or ( \1797_b1 , \1785_b1 , \1796_b1 );
not ( \1796_b1 , w_3908 );
and ( \1797_b0 , \1785_b0 , w_3909 );
and ( w_3908 , w_3909 , \1796_b0 );
or ( \1798_b1 , \1760_b1 , \1796_b1 );
not ( \1796_b1 , w_3910 );
and ( \1798_b0 , \1760_b0 , w_3911 );
and ( w_3910 , w_3911 , \1796_b0 );
or ( \1800_b1 , \1603_b1 , \1623_b1 );
xor ( \1800_b0 , \1603_b0 , w_3912 );
not ( w_3912 , w_3913 );
and ( w_3913 , \1623_b1 , \1623_b0 );
or ( \1801_b1 , \1800_b1 , \1640_b1 );
xor ( \1801_b0 , \1800_b0 , w_3914 );
not ( w_3914 , w_3915 );
and ( w_3915 , \1640_b1 , \1640_b0 );
or ( \1802_b1 , \1645_b1 , \1647_b1 );
xor ( \1802_b0 , \1645_b0 , w_3916 );
not ( w_3916 , w_3917 );
and ( w_3917 , \1647_b1 , \1647_b0 );
or ( \1803_b1 , \1802_b1 , \1650_b1 );
xor ( \1803_b0 , \1802_b0 , w_3918 );
not ( w_3918 , w_3919 );
and ( w_3919 , \1650_b1 , \1650_b0 );
or ( \1804_b1 , \1801_b1 , \1803_b1 );
not ( \1803_b1 , w_3920 );
and ( \1804_b0 , \1801_b0 , w_3921 );
and ( w_3920 , w_3921 , \1803_b0 );
or ( \1805_b1 , \1670_b1 , w_3922 );
xor ( \1805_b0 , \1670_b0 , w_3924 );
not ( w_3924 , w_3925 );
and ( w_3925 , w_3922 , w_3923 );
buf ( w_3922 , \1672_b1 );
not ( w_3922 , w_3926 );
not ( w_3923 , w_3927 );
and ( w_3926 , w_3927 , \1672_b0 );
or ( \1806_b1 , \1803_b1 , \1805_b1 );
not ( \1805_b1 , w_3928 );
and ( \1806_b0 , \1803_b0 , w_3929 );
and ( w_3928 , w_3929 , \1805_b0 );
or ( \1807_b1 , \1801_b1 , \1805_b1 );
not ( \1805_b1 , w_3930 );
and ( \1807_b0 , \1801_b0 , w_3931 );
and ( w_3930 , w_3931 , \1805_b0 );
or ( \1809_b1 , \1799_b1 , \1808_b1 );
not ( \1808_b1 , w_3932 );
and ( \1809_b0 , \1799_b0 , w_3933 );
and ( w_3932 , w_3933 , \1808_b0 );
or ( \1810_b1 , \1678_b1 , \1680_b1 );
xor ( \1810_b0 , \1678_b0 , w_3934 );
not ( w_3934 , w_3935 );
and ( w_3935 , \1680_b1 , \1680_b0 );
or ( \1811_b1 , \1810_b1 , \1682_b1 );
xor ( \1811_b0 , \1810_b0 , w_3936 );
not ( w_3936 , w_3937 );
and ( w_3937 , \1682_b1 , \1682_b0 );
or ( \1812_b1 , \1808_b1 , \1811_b1 );
not ( \1811_b1 , w_3938 );
and ( \1812_b0 , \1808_b0 , w_3939 );
and ( w_3938 , w_3939 , \1811_b0 );
or ( \1813_b1 , \1799_b1 , \1811_b1 );
not ( \1811_b1 , w_3940 );
and ( \1813_b0 , \1799_b0 , w_3941 );
and ( w_3940 , w_3941 , \1811_b0 );
or ( \1815_b1 , \1527_b1 , \1549_b1 );
xor ( \1815_b0 , \1527_b0 , w_3942 );
not ( w_3942 , w_3943 );
and ( w_3943 , \1549_b1 , \1549_b0 );
or ( \1816_b1 , \1815_b1 , \1555_b1 );
xor ( \1816_b0 , \1815_b0 , w_3944 );
not ( w_3944 , w_3945 );
and ( w_3945 , \1555_b1 , \1555_b0 );
or ( \1817_b1 , \1814_b1 , \1816_b1 );
not ( \1816_b1 , w_3946 );
and ( \1817_b0 , \1814_b0 , w_3947 );
and ( w_3946 , w_3947 , \1816_b0 );
or ( \1818_b1 , \1676_b1 , \1685_b1 );
xor ( \1818_b0 , \1676_b0 , w_3948 );
not ( w_3948 , w_3949 );
and ( w_3949 , \1685_b1 , \1685_b0 );
or ( \1819_b1 , \1818_b1 , \1688_b1 );
xor ( \1819_b0 , \1818_b0 , w_3950 );
not ( w_3950 , w_3951 );
and ( w_3951 , \1688_b1 , \1688_b0 );
or ( \1820_b1 , \1816_b1 , \1819_b1 );
not ( \1819_b1 , w_3952 );
and ( \1820_b0 , \1816_b0 , w_3953 );
and ( w_3952 , w_3953 , \1819_b0 );
or ( \1821_b1 , \1814_b1 , \1819_b1 );
not ( \1819_b1 , w_3954 );
and ( \1821_b0 , \1814_b0 , w_3955 );
and ( w_3954 , w_3955 , \1819_b0 );
or ( \1823_b1 , \1691_b1 , \1693_b1 );
xor ( \1823_b0 , \1691_b0 , w_3956 );
not ( w_3956 , w_3957 );
and ( w_3957 , \1693_b1 , \1693_b0 );
or ( \1824_b1 , \1823_b1 , \1696_b1 );
xor ( \1824_b0 , \1823_b0 , w_3958 );
not ( w_3958 , w_3959 );
and ( w_3959 , \1696_b1 , \1696_b0 );
or ( \1825_b1 , \1822_b1 , \1824_b1 );
not ( \1824_b1 , w_3960 );
and ( \1825_b0 , \1822_b0 , w_3961 );
and ( w_3960 , w_3961 , \1824_b0 );
or ( \1826_b1 , \1705_b1 , \1825_b1 );
not ( \1825_b1 , w_3962 );
and ( \1826_b0 , \1705_b0 , w_3963 );
and ( w_3962 , w_3963 , \1825_b0 );
or ( \1827_b1 , \1705_b1 , \1825_b1 );
xor ( \1827_b0 , \1705_b0 , w_3964 );
not ( w_3964 , w_3965 );
and ( w_3965 , \1825_b1 , \1825_b0 );
or ( \1828_b1 , \1822_b1 , \1824_b1 );
xor ( \1828_b0 , \1822_b0 , w_3966 );
not ( w_3966 , w_3967 );
and ( w_3967 , \1824_b1 , \1824_b0 );
and ( \1829_nR12a_b1 , RIb4c2d50_58_b1 , w_3968 );
xor ( w_3968 , RIb4c2d50_58_b0 , \288_b1 );
not ( \288_b1 , w_3969 );
and ( \1829_nR12a_b0 , w_3969 , \288_b0 );
buf ( \1830_b1 , \1829_nR12a_b1 );
buf ( \1830_b0 , \1829_nR12a_b0 );
and ( \1831_nR129_b1 , RIb4c2cd8_59_b1 , w_3970 );
xor ( w_3970 , RIb4c2cd8_59_b0 , \288_b1 );
not ( \288_b1 , w_3971 );
and ( \1831_nR129_b0 , w_3971 , \288_b0 );
buf ( \1832_b1 , \1831_nR129_b1 );
buf ( \1832_b0 , \1831_nR129_b0 );
or ( \1833_b1 , \1830_b1 , \1832_b1 );
not ( \1832_b1 , w_3972 );
and ( \1833_b0 , \1830_b0 , w_3973 );
and ( w_3972 , w_3973 , \1832_b0 );
buf ( \1834_b1 , \1833_b1 );
not ( \1834_b1 , w_3974 );
not ( \1834_b0 , w_3975 );
and ( w_3974 , w_3975 , \1833_b0 );
or ( \1835_b1 , \1607_b1 , \1834_b1 );
not ( \1834_b1 , w_3976 );
and ( \1835_b0 , \1607_b0 , w_3977 );
and ( w_3976 , w_3977 , \1834_b0 );
buf ( \1836_b1 , \1835_b1 );
not ( \1836_b1 , w_3978 );
not ( \1836_b0 , w_3979 );
and ( w_3978 , w_3979 , \1835_b0 );
or ( \1837_b1 , \315_b1 , \1742_b1 );
not ( \1742_b1 , w_3980 );
and ( \1837_b0 , \315_b0 , w_3981 );
and ( w_3980 , w_3981 , \1742_b0 );
or ( \1838_b1 , \159_b1 , \1740_b1 );
not ( \1740_b1 , w_3982 );
and ( \1838_b0 , \159_b0 , w_3983 );
and ( w_3982 , w_3983 , \1740_b0 );
or ( \1839_b1 , \1837_b1 , w_3985 );
not ( w_3985 , w_3986 );
and ( \1839_b0 , \1837_b0 , w_3987 );
and ( w_3986 ,  , w_3987 );
buf ( w_3985 , \1838_b1 );
not ( w_3985 , w_3988 );
not (  , w_3989 );
and ( w_3988 , w_3989 , \1838_b0 );
or ( \1840_b1 , \1839_b1 , w_3990 );
xor ( \1840_b0 , \1839_b0 , w_3992 );
not ( w_3992 , w_3993 );
and ( w_3993 , w_3990 , w_3991 );
buf ( w_3990 , \1610_b1 );
not ( w_3990 , w_3994 );
not ( w_3991 , w_3995 );
and ( w_3994 , w_3995 , \1610_b0 );
or ( \1841_b1 , \1836_b1 , \1840_b1 );
not ( \1840_b1 , w_3996 );
and ( \1841_b0 , \1836_b0 , w_3997 );
and ( w_3996 , w_3997 , \1840_b0 );
or ( \1842_b1 , \333_b1 , \1476_b1 );
not ( \1476_b1 , w_3998 );
and ( \1842_b0 , \333_b0 , w_3999 );
and ( w_3998 , w_3999 , \1476_b0 );
or ( \1843_b1 , \305_b1 , \1474_b1 );
not ( \1474_b1 , w_4000 );
and ( \1843_b0 , \305_b0 , w_4001 );
and ( w_4000 , w_4001 , \1474_b0 );
or ( \1844_b1 , \1842_b1 , w_4003 );
not ( w_4003 , w_4004 );
and ( \1844_b0 , \1842_b0 , w_4005 );
and ( w_4004 ,  , w_4005 );
buf ( w_4003 , \1843_b1 );
not ( w_4003 , w_4006 );
not (  , w_4007 );
and ( w_4006 , w_4007 , \1843_b0 );
or ( \1845_b1 , \1844_b1 , w_4008 );
xor ( \1845_b0 , \1844_b0 , w_4010 );
not ( w_4010 , w_4011 );
and ( w_4011 , w_4008 , w_4009 );
buf ( w_4008 , \1363_b1 );
not ( w_4008 , w_4012 );
not ( w_4009 , w_4013 );
and ( w_4012 , w_4013 , \1363_b0 );
or ( \1846_b1 , \1840_b1 , \1845_b1 );
not ( \1845_b1 , w_4014 );
and ( \1846_b0 , \1840_b0 , w_4015 );
and ( w_4014 , w_4015 , \1845_b0 );
or ( \1847_b1 , \1836_b1 , \1845_b1 );
not ( \1845_b1 , w_4016 );
and ( \1847_b0 , \1836_b0 , w_4017 );
and ( w_4016 , w_4017 , \1845_b0 );
or ( \1849_b1 , \353_b1 , \1280_b1 );
not ( \1280_b1 , w_4018 );
and ( \1849_b0 , \353_b0 , w_4019 );
and ( w_4018 , w_4019 , \1280_b0 );
or ( \1850_b1 , \323_b1 , \1278_b1 );
not ( \1278_b1 , w_4020 );
and ( \1850_b0 , \323_b0 , w_4021 );
and ( w_4020 , w_4021 , \1278_b0 );
or ( \1851_b1 , \1849_b1 , w_4023 );
not ( w_4023 , w_4024 );
and ( \1851_b0 , \1849_b0 , w_4025 );
and ( w_4024 ,  , w_4025 );
buf ( w_4023 , \1850_b1 );
not ( w_4023 , w_4026 );
not (  , w_4027 );
and ( w_4026 , w_4027 , \1850_b0 );
or ( \1852_b1 , \1851_b1 , w_4028 );
xor ( \1852_b0 , \1851_b0 , w_4030 );
not ( w_4030 , w_4031 );
and ( w_4031 , w_4028 , w_4029 );
buf ( w_4028 , \1177_b1 );
not ( w_4028 , w_4032 );
not ( w_4029 , w_4033 );
and ( w_4032 , w_4033 , \1177_b0 );
or ( \1853_b1 , \360_b1 , \1062_b1 );
not ( \1062_b1 , w_4034 );
and ( \1853_b0 , \360_b0 , w_4035 );
and ( w_4034 , w_4035 , \1062_b0 );
or ( \1854_b1 , \343_b1 , \1060_b1 );
not ( \1060_b1 , w_4036 );
and ( \1854_b0 , \343_b0 , w_4037 );
and ( w_4036 , w_4037 , \1060_b0 );
or ( \1855_b1 , \1853_b1 , w_4039 );
not ( w_4039 , w_4040 );
and ( \1855_b0 , \1853_b0 , w_4041 );
and ( w_4040 ,  , w_4041 );
buf ( w_4039 , \1854_b1 );
not ( w_4039 , w_4042 );
not (  , w_4043 );
and ( w_4042 , w_4043 , \1854_b0 );
or ( \1856_b1 , \1855_b1 , w_4044 );
xor ( \1856_b0 , \1855_b0 , w_4046 );
not ( w_4046 , w_4047 );
and ( w_4047 , w_4044 , w_4045 );
buf ( w_4044 , \984_b1 );
not ( w_4044 , w_4048 );
not ( w_4045 , w_4049 );
and ( w_4048 , w_4049 , \984_b0 );
or ( \1857_b1 , \1852_b1 , \1856_b1 );
not ( \1856_b1 , w_4050 );
and ( \1857_b0 , \1852_b0 , w_4051 );
and ( w_4050 , w_4051 , \1856_b0 );
or ( \1858_b1 , \495_b1 , \912_b1 );
not ( \912_b1 , w_4052 );
and ( \1858_b0 , \495_b0 , w_4053 );
and ( w_4052 , w_4053 , \912_b0 );
or ( \1859_b1 , \444_b1 , \910_b1 );
not ( \910_b1 , w_4054 );
and ( \1859_b0 , \444_b0 , w_4055 );
and ( w_4054 , w_4055 , \910_b0 );
or ( \1860_b1 , \1858_b1 , w_4057 );
not ( w_4057 , w_4058 );
and ( \1860_b0 , \1858_b0 , w_4059 );
and ( w_4058 ,  , w_4059 );
buf ( w_4057 , \1859_b1 );
not ( w_4057 , w_4060 );
not (  , w_4061 );
and ( w_4060 , w_4061 , \1859_b0 );
or ( \1861_b1 , \1860_b1 , w_4062 );
xor ( \1861_b0 , \1860_b0 , w_4064 );
not ( w_4064 , w_4065 );
and ( w_4065 , w_4062 , w_4063 );
buf ( w_4062 , \818_b1 );
not ( w_4062 , w_4066 );
not ( w_4063 , w_4067 );
and ( w_4066 , w_4067 , \818_b0 );
or ( \1862_b1 , \1856_b1 , \1861_b1 );
not ( \1861_b1 , w_4068 );
and ( \1862_b0 , \1856_b0 , w_4069 );
and ( w_4068 , w_4069 , \1861_b0 );
or ( \1863_b1 , \1852_b1 , \1861_b1 );
not ( \1861_b1 , w_4070 );
and ( \1863_b0 , \1852_b0 , w_4071 );
and ( w_4070 , w_4071 , \1861_b0 );
or ( \1865_b1 , \1848_b1 , \1864_b1 );
not ( \1864_b1 , w_4072 );
and ( \1865_b0 , \1848_b0 , w_4073 );
and ( w_4072 , w_4073 , \1864_b0 );
or ( \1866_b1 , \621_b1 , \740_b1 );
not ( \740_b1 , w_4074 );
and ( \1866_b0 , \621_b0 , w_4075 );
and ( w_4074 , w_4075 , \740_b0 );
or ( \1867_b1 , \593_b1 , \738_b1 );
not ( \738_b1 , w_4076 );
and ( \1867_b0 , \593_b0 , w_4077 );
and ( w_4076 , w_4077 , \738_b0 );
or ( \1868_b1 , \1866_b1 , w_4079 );
not ( w_4079 , w_4080 );
and ( \1868_b0 , \1866_b0 , w_4081 );
and ( w_4080 ,  , w_4081 );
buf ( w_4079 , \1867_b1 );
not ( w_4079 , w_4082 );
not (  , w_4083 );
and ( w_4082 , w_4083 , \1867_b0 );
or ( \1869_b1 , \1868_b1 , w_4084 );
xor ( \1869_b0 , \1868_b0 , w_4086 );
not ( w_4086 , w_4087 );
and ( w_4087 , w_4084 , w_4085 );
buf ( w_4084 , \668_b1 );
not ( w_4084 , w_4088 );
not ( w_4085 , w_4089 );
and ( w_4088 , w_4089 , \668_b0 );
or ( \1870_b1 , \777_b1 , \604_b1 );
not ( \604_b1 , w_4090 );
and ( \1870_b0 , \777_b0 , w_4091 );
and ( w_4090 , w_4091 , \604_b0 );
or ( \1871_b1 , \703_b1 , \602_b1 );
not ( \602_b1 , w_4092 );
and ( \1871_b0 , \703_b0 , w_4093 );
and ( w_4092 , w_4093 , \602_b0 );
or ( \1872_b1 , \1870_b1 , w_4095 );
not ( w_4095 , w_4096 );
and ( \1872_b0 , \1870_b0 , w_4097 );
and ( w_4096 ,  , w_4097 );
buf ( w_4095 , \1871_b1 );
not ( w_4095 , w_4098 );
not (  , w_4099 );
and ( w_4098 , w_4099 , \1871_b0 );
or ( \1873_b1 , \1872_b1 , w_4100 );
xor ( \1873_b0 , \1872_b0 , w_4102 );
not ( w_4102 , w_4103 );
and ( w_4103 , w_4100 , w_4101 );
buf ( w_4100 , \561_b1 );
not ( w_4100 , w_4104 );
not ( w_4101 , w_4105 );
and ( w_4104 , w_4105 , \561_b0 );
or ( \1874_b1 , \1869_b1 , \1873_b1 );
not ( \1873_b1 , w_4106 );
and ( \1874_b0 , \1869_b0 , w_4107 );
and ( w_4106 , w_4107 , \1873_b0 );
or ( \1875_b1 , \904_b1 , \503_b1 );
not ( \503_b1 , w_4108 );
and ( \1875_b0 , \904_b0 , w_4109 );
and ( w_4108 , w_4109 , \503_b0 );
or ( \1876_b1 , \841_b1 , \501_b1 );
not ( \501_b1 , w_4110 );
and ( \1876_b0 , \841_b0 , w_4111 );
and ( w_4110 , w_4111 , \501_b0 );
or ( \1877_b1 , \1875_b1 , w_4113 );
not ( w_4113 , w_4114 );
and ( \1877_b0 , \1875_b0 , w_4115 );
and ( w_4114 ,  , w_4115 );
buf ( w_4113 , \1876_b1 );
not ( w_4113 , w_4116 );
not (  , w_4117 );
and ( w_4116 , w_4117 , \1876_b0 );
or ( \1878_b1 , \1877_b1 , w_4118 );
xor ( \1878_b0 , \1877_b0 , w_4120 );
not ( w_4120 , w_4121 );
and ( w_4121 , w_4118 , w_4119 );
buf ( w_4118 , \455_b1 );
not ( w_4118 , w_4122 );
not ( w_4119 , w_4123 );
and ( w_4122 , w_4123 , \455_b0 );
or ( \1879_b1 , \1873_b1 , \1878_b1 );
not ( \1878_b1 , w_4124 );
and ( \1879_b0 , \1873_b0 , w_4125 );
and ( w_4124 , w_4125 , \1878_b0 );
or ( \1880_b1 , \1869_b1 , \1878_b1 );
not ( \1878_b1 , w_4126 );
and ( \1880_b0 , \1869_b0 , w_4127 );
and ( w_4126 , w_4127 , \1878_b0 );
or ( \1882_b1 , \1864_b1 , \1881_b1 );
not ( \1881_b1 , w_4128 );
and ( \1882_b0 , \1864_b0 , w_4129 );
and ( w_4128 , w_4129 , \1881_b0 );
or ( \1883_b1 , \1848_b1 , \1881_b1 );
not ( \1881_b1 , w_4130 );
and ( \1883_b0 , \1848_b0 , w_4131 );
and ( w_4130 , w_4131 , \1881_b0 );
or ( \1885_b1 , \1709_b1 , \1713_b1 );
xor ( \1885_b0 , \1709_b0 , w_4132 );
not ( w_4132 , w_4133 );
and ( w_4133 , \1713_b1 , \1713_b0 );
or ( \1886_b1 , \1885_b1 , \1718_b1 );
xor ( \1886_b0 , \1885_b0 , w_4134 );
not ( w_4134 , w_4135 );
and ( w_4135 , \1718_b1 , \1718_b0 );
or ( \1887_b1 , \1725_b1 , \1729_b1 );
xor ( \1887_b0 , \1725_b0 , w_4136 );
not ( w_4136 , w_4137 );
and ( w_4137 , \1729_b1 , \1729_b0 );
or ( \1888_b1 , \1887_b1 , \1734_b1 );
xor ( \1888_b0 , \1887_b0 , w_4138 );
not ( w_4138 , w_4139 );
and ( w_4139 , \1734_b1 , \1734_b0 );
or ( \1889_b1 , \1886_b1 , \1888_b1 );
not ( \1888_b1 , w_4140 );
and ( \1889_b0 , \1886_b0 , w_4141 );
and ( w_4140 , w_4141 , \1888_b0 );
or ( \1890_b1 , \1745_b1 , \1749_b1 );
xor ( \1890_b0 , \1745_b0 , w_4142 );
not ( w_4142 , w_4143 );
and ( w_4143 , \1749_b1 , \1749_b0 );
or ( \1891_b1 , \1890_b1 , \1754_b1 );
xor ( \1891_b0 , \1890_b0 , w_4144 );
not ( w_4144 , w_4145 );
and ( w_4145 , \1754_b1 , \1754_b0 );
or ( \1892_b1 , \1888_b1 , \1891_b1 );
not ( \1891_b1 , w_4146 );
and ( \1892_b0 , \1888_b0 , w_4147 );
and ( w_4146 , w_4147 , \1891_b0 );
or ( \1893_b1 , \1886_b1 , \1891_b1 );
not ( \1891_b1 , w_4148 );
and ( \1893_b0 , \1886_b0 , w_4149 );
and ( w_4148 , w_4149 , \1891_b0 );
or ( \1895_b1 , \1884_b1 , \1894_b1 );
not ( \1894_b1 , w_4150 );
and ( \1895_b0 , \1884_b0 , w_4151 );
and ( w_4150 , w_4151 , \1894_b0 );
or ( \1896_b1 , \1194_b1 , \298_b1 );
not ( \298_b1 , w_4152 );
and ( \1896_b0 , \1194_b0 , w_4153 );
and ( w_4152 , w_4153 , \298_b0 );
or ( \1897_b1 , \1104_b1 , \296_b1 );
not ( \296_b1 , w_4154 );
and ( \1897_b0 , \1104_b0 , w_4155 );
and ( w_4154 , w_4155 , \296_b0 );
or ( \1898_b1 , \1896_b1 , w_4157 );
not ( w_4157 , w_4158 );
and ( \1898_b0 , \1896_b0 , w_4159 );
and ( w_4158 ,  , w_4159 );
buf ( w_4157 , \1897_b1 );
not ( w_4157 , w_4160 );
not (  , w_4161 );
and ( w_4160 , w_4161 , \1897_b0 );
or ( \1899_b1 , \1898_b1 , w_4162 );
xor ( \1899_b0 , \1898_b0 , w_4164 );
not ( w_4164 , w_4165 );
and ( w_4165 , w_4162 , w_4163 );
buf ( w_4162 , \303_b1 );
not ( w_4162 , w_4166 );
not ( w_4163 , w_4167 );
and ( w_4166 , w_4167 , \303_b0 );
or ( \1900_b1 , \1304_b1 , \313_b1 );
not ( \313_b1 , w_4168 );
and ( \1900_b0 , \1304_b0 , w_4169 );
and ( w_4168 , w_4169 , \313_b0 );
or ( \1901_b1 , \1299_b1 , \311_b1 );
not ( \311_b1 , w_4170 );
and ( \1901_b0 , \1299_b0 , w_4171 );
and ( w_4170 , w_4171 , \311_b0 );
or ( \1902_b1 , \1900_b1 , w_4173 );
not ( w_4173 , w_4174 );
and ( \1902_b0 , \1900_b0 , w_4175 );
and ( w_4174 ,  , w_4175 );
buf ( w_4173 , \1901_b1 );
not ( w_4173 , w_4176 );
not (  , w_4177 );
and ( w_4176 , w_4177 , \1901_b0 );
or ( \1903_b1 , \1902_b1 , w_4178 );
xor ( \1903_b0 , \1902_b0 , w_4180 );
not ( w_4180 , w_4181 );
and ( w_4181 , w_4178 , w_4179 );
buf ( w_4178 , \320_b1 );
not ( w_4178 , w_4182 );
not ( w_4179 , w_4183 );
and ( w_4182 , w_4183 , \320_b0 );
or ( \1904_b1 , \1899_b1 , \1903_b1 );
not ( \1903_b1 , w_4184 );
and ( \1904_b0 , \1899_b0 , w_4185 );
and ( w_4184 , w_4185 , \1903_b0 );
or ( \1905_b1 , \1537_b1 , \331_b1 );
not ( \331_b1 , w_4186 );
and ( \1905_b0 , \1537_b0 , w_4187 );
and ( w_4186 , w_4187 , \331_b0 );
or ( \1906_b1 , \1422_b1 , \329_b1 );
not ( \329_b1 , w_4188 );
and ( \1906_b0 , \1422_b0 , w_4189 );
and ( w_4188 , w_4189 , \329_b0 );
or ( \1907_b1 , \1905_b1 , w_4191 );
not ( w_4191 , w_4192 );
and ( \1907_b0 , \1905_b0 , w_4193 );
and ( w_4192 ,  , w_4193 );
buf ( w_4191 , \1906_b1 );
not ( w_4191 , w_4194 );
not (  , w_4195 );
and ( w_4194 , w_4195 , \1906_b0 );
or ( \1908_b1 , \1907_b1 , w_4196 );
xor ( \1908_b0 , \1907_b0 , w_4198 );
not ( w_4198 , w_4199 );
and ( w_4199 , w_4196 , w_4197 );
buf ( w_4196 , \338_b1 );
not ( w_4196 , w_4200 );
not ( w_4197 , w_4201 );
and ( w_4200 , w_4201 , \338_b0 );
or ( \1909_b1 , \1903_b1 , \1908_b1 );
not ( \1908_b1 , w_4202 );
and ( \1909_b0 , \1903_b0 , w_4203 );
and ( w_4202 , w_4203 , \1908_b0 );
or ( \1910_b1 , \1899_b1 , \1908_b1 );
not ( \1908_b1 , w_4204 );
and ( \1910_b0 , \1899_b0 , w_4205 );
and ( w_4204 , w_4205 , \1908_b0 );
or ( \1912_b1 , \1764_b1 , \1768_b1 );
xor ( \1912_b0 , \1764_b0 , w_4206 );
not ( w_4206 , w_4207 );
and ( w_4207 , \1768_b1 , \1768_b0 );
or ( \1913_b1 , \1912_b1 , \1774_b1 );
xor ( \1913_b0 , \1912_b0 , w_4208 );
not ( w_4208 , w_4209 );
and ( w_4209 , \1774_b1 , \1774_b0 );
or ( \1914_b1 , \1911_b1 , \1913_b1 );
not ( \1913_b1 , w_4210 );
and ( \1914_b0 , \1911_b0 , w_4211 );
and ( w_4210 , w_4211 , \1913_b0 );
buf ( \1915_b1 , \1779_b1 );
not ( \1915_b1 , w_4212 );
not ( \1915_b0 , w_4213 );
and ( w_4212 , w_4213 , \1779_b0 );
or ( \1916_b1 , \1913_b1 , \1915_b1 );
not ( \1915_b1 , w_4214 );
and ( \1916_b0 , \1913_b0 , w_4215 );
and ( w_4214 , w_4215 , \1915_b0 );
or ( \1917_b1 , \1911_b1 , \1915_b1 );
not ( \1915_b1 , w_4216 );
and ( \1917_b0 , \1911_b0 , w_4217 );
and ( w_4216 , w_4217 , \1915_b0 );
or ( \1919_b1 , \1894_b1 , \1918_b1 );
not ( \1918_b1 , w_4218 );
and ( \1919_b0 , \1894_b0 , w_4219 );
and ( w_4218 , w_4219 , \1918_b0 );
or ( \1920_b1 , \1884_b1 , \1918_b1 );
not ( \1918_b1 , w_4220 );
and ( \1920_b0 , \1884_b0 , w_4221 );
and ( w_4220 , w_4221 , \1918_b0 );
or ( \1922_b1 , \1611_b1 , \1615_b1 );
xor ( \1922_b0 , \1611_b0 , w_4222 );
not ( w_4222 , w_4223 );
and ( w_4223 , \1615_b1 , \1615_b0 );
or ( \1923_b1 , \1922_b1 , \1620_b1 );
xor ( \1923_b0 , \1922_b0 , w_4224 );
not ( w_4224 , w_4225 );
and ( w_4225 , \1620_b1 , \1620_b0 );
or ( \1924_b1 , \1777_b1 , \1780_b1 );
xor ( \1924_b0 , \1777_b0 , w_4226 );
not ( w_4226 , w_4227 );
and ( w_4227 , \1780_b1 , \1780_b0 );
or ( \1925_b1 , \1924_b1 , \1782_b1 );
xor ( \1925_b0 , \1924_b0 , w_4228 );
not ( w_4228 , w_4229 );
and ( w_4229 , \1782_b1 , \1782_b0 );
or ( \1926_b1 , \1923_b1 , \1925_b1 );
not ( \1925_b1 , w_4230 );
and ( \1926_b0 , \1923_b0 , w_4231 );
and ( w_4230 , w_4231 , \1925_b0 );
or ( \1927_b1 , \1788_b1 , \1790_b1 );
xor ( \1927_b0 , \1788_b0 , w_4232 );
not ( w_4232 , w_4233 );
and ( w_4233 , \1790_b1 , \1790_b0 );
or ( \1928_b1 , \1927_b1 , \1793_b1 );
xor ( \1928_b0 , \1927_b0 , w_4234 );
not ( w_4234 , w_4235 );
and ( w_4235 , \1793_b1 , \1793_b0 );
or ( \1929_b1 , \1925_b1 , \1928_b1 );
not ( \1928_b1 , w_4236 );
and ( \1929_b0 , \1925_b0 , w_4237 );
and ( w_4236 , w_4237 , \1928_b0 );
or ( \1930_b1 , \1923_b1 , \1928_b1 );
not ( \1928_b1 , w_4238 );
and ( \1930_b0 , \1923_b0 , w_4239 );
and ( w_4238 , w_4239 , \1928_b0 );
or ( \1932_b1 , \1921_b1 , \1931_b1 );
not ( \1931_b1 , w_4240 );
and ( \1932_b0 , \1921_b0 , w_4241 );
and ( w_4240 , w_4241 , \1931_b0 );
or ( \1933_b1 , \1801_b1 , \1803_b1 );
xor ( \1933_b0 , \1801_b0 , w_4242 );
not ( w_4242 , w_4243 );
and ( w_4243 , \1803_b1 , \1803_b0 );
or ( \1934_b1 , \1933_b1 , \1805_b1 );
xor ( \1934_b0 , \1933_b0 , w_4244 );
not ( w_4244 , w_4245 );
and ( w_4245 , \1805_b1 , \1805_b0 );
or ( \1935_b1 , \1931_b1 , \1934_b1 );
not ( \1934_b1 , w_4246 );
and ( \1935_b0 , \1931_b0 , w_4247 );
and ( w_4246 , w_4247 , \1934_b0 );
or ( \1936_b1 , \1921_b1 , \1934_b1 );
not ( \1934_b1 , w_4248 );
and ( \1936_b0 , \1921_b0 , w_4249 );
and ( w_4248 , w_4249 , \1934_b0 );
or ( \1938_b1 , \1643_b1 , \1653_b1 );
xor ( \1938_b0 , \1643_b0 , w_4250 );
not ( w_4250 , w_4251 );
and ( w_4251 , \1653_b1 , \1653_b0 );
or ( \1939_b1 , \1938_b1 , \1673_b1 );
xor ( \1939_b0 , \1938_b0 , w_4252 );
not ( w_4252 , w_4253 );
and ( w_4253 , \1673_b1 , \1673_b0 );
or ( \1940_b1 , \1937_b1 , \1939_b1 );
not ( \1939_b1 , w_4254 );
and ( \1940_b0 , \1937_b0 , w_4255 );
and ( w_4254 , w_4255 , \1939_b0 );
or ( \1941_b1 , \1799_b1 , \1808_b1 );
xor ( \1941_b0 , \1799_b0 , w_4256 );
not ( w_4256 , w_4257 );
and ( w_4257 , \1808_b1 , \1808_b0 );
or ( \1942_b1 , \1941_b1 , \1811_b1 );
xor ( \1942_b0 , \1941_b0 , w_4258 );
not ( w_4258 , w_4259 );
and ( w_4259 , \1811_b1 , \1811_b0 );
or ( \1943_b1 , \1939_b1 , \1942_b1 );
not ( \1942_b1 , w_4260 );
and ( \1943_b0 , \1939_b0 , w_4261 );
and ( w_4260 , w_4261 , \1942_b0 );
or ( \1944_b1 , \1937_b1 , \1942_b1 );
not ( \1942_b1 , w_4262 );
and ( \1944_b0 , \1937_b0 , w_4263 );
and ( w_4262 , w_4263 , \1942_b0 );
or ( \1946_b1 , \1814_b1 , \1816_b1 );
xor ( \1946_b0 , \1814_b0 , w_4264 );
not ( w_4264 , w_4265 );
and ( w_4265 , \1816_b1 , \1816_b0 );
or ( \1947_b1 , \1946_b1 , \1819_b1 );
xor ( \1947_b0 , \1946_b0 , w_4266 );
not ( w_4266 , w_4267 );
and ( w_4267 , \1819_b1 , \1819_b0 );
or ( \1948_b1 , \1945_b1 , \1947_b1 );
not ( \1947_b1 , w_4268 );
and ( \1948_b0 , \1945_b0 , w_4269 );
and ( w_4268 , w_4269 , \1947_b0 );
or ( \1949_b1 , \1828_b1 , \1948_b1 );
not ( \1948_b1 , w_4270 );
and ( \1949_b0 , \1828_b0 , w_4271 );
and ( w_4270 , w_4271 , \1948_b0 );
or ( \1950_b1 , \1828_b1 , \1948_b1 );
xor ( \1950_b0 , \1828_b0 , w_4272 );
not ( w_4272 , w_4273 );
and ( w_4273 , \1948_b1 , \1948_b0 );
or ( \1951_b1 , \1945_b1 , \1947_b1 );
xor ( \1951_b0 , \1945_b0 , w_4274 );
not ( w_4274 , w_4275 );
and ( w_4275 , \1947_b1 , \1947_b0 );
or ( \1952_b1 , \1607_b1 , \1830_b1 );
xor ( \1952_b0 , \1607_b0 , w_4276 );
not ( w_4276 , w_4277 );
and ( w_4277 , \1830_b1 , \1830_b0 );
or ( \1953_b1 , \1830_b1 , \1832_b1 );
xor ( \1953_b0 , \1830_b0 , w_4278 );
not ( w_4278 , w_4279 );
and ( w_4279 , \1832_b1 , \1832_b0 );
buf ( \1954_b1 , \1953_b1 );
not ( \1954_b1 , w_4280 );
not ( \1954_b0 , w_4281 );
and ( w_4280 , w_4281 , \1953_b0 );
or ( \1955_b1 , \1952_b1 , \1954_b1 );
not ( \1954_b1 , w_4282 );
and ( \1955_b0 , \1952_b0 , w_4283 );
and ( w_4282 , w_4283 , \1954_b0 );
or ( \1956_b1 , \159_b1 , \1955_b1 );
not ( \1955_b1 , w_4284 );
and ( \1956_b0 , \159_b0 , w_4285 );
and ( w_4284 , w_4285 , \1955_b0 );
buf ( \1957_b1 , \1956_b1 );
not ( \1957_b1 , w_4286 );
not ( \1957_b0 , w_4287 );
and ( w_4286 , w_4287 , \1956_b0 );
or ( \1958_b1 , \1957_b1 , w_4288 );
xor ( \1958_b0 , \1957_b0 , w_4290 );
not ( w_4290 , w_4291 );
and ( w_4291 , w_4288 , w_4289 );
buf ( w_4288 , \1835_b1 );
not ( w_4288 , w_4292 );
not ( w_4289 , w_4293 );
and ( w_4292 , w_4293 , \1835_b0 );
or ( \1959_b1 , \305_b1 , \1742_b1 );
not ( \1742_b1 , w_4294 );
and ( \1959_b0 , \305_b0 , w_4295 );
and ( w_4294 , w_4295 , \1742_b0 );
or ( \1960_b1 , \315_b1 , \1740_b1 );
not ( \1740_b1 , w_4296 );
and ( \1960_b0 , \315_b0 , w_4297 );
and ( w_4296 , w_4297 , \1740_b0 );
or ( \1961_b1 , \1959_b1 , w_4299 );
not ( w_4299 , w_4300 );
and ( \1961_b0 , \1959_b0 , w_4301 );
and ( w_4300 ,  , w_4301 );
buf ( w_4299 , \1960_b1 );
not ( w_4299 , w_4302 );
not (  , w_4303 );
and ( w_4302 , w_4303 , \1960_b0 );
or ( \1962_b1 , \1961_b1 , w_4304 );
xor ( \1962_b0 , \1961_b0 , w_4306 );
not ( w_4306 , w_4307 );
and ( w_4307 , w_4304 , w_4305 );
buf ( w_4304 , \1610_b1 );
not ( w_4304 , w_4308 );
not ( w_4305 , w_4309 );
and ( w_4308 , w_4309 , \1610_b0 );
or ( \1963_b1 , \1958_b1 , \1962_b1 );
not ( \1962_b1 , w_4310 );
and ( \1963_b0 , \1958_b0 , w_4311 );
and ( w_4310 , w_4311 , \1962_b0 );
or ( \1964_b1 , \323_b1 , \1476_b1 );
not ( \1476_b1 , w_4312 );
and ( \1964_b0 , \323_b0 , w_4313 );
and ( w_4312 , w_4313 , \1476_b0 );
or ( \1965_b1 , \333_b1 , \1474_b1 );
not ( \1474_b1 , w_4314 );
and ( \1965_b0 , \333_b0 , w_4315 );
and ( w_4314 , w_4315 , \1474_b0 );
or ( \1966_b1 , \1964_b1 , w_4317 );
not ( w_4317 , w_4318 );
and ( \1966_b0 , \1964_b0 , w_4319 );
and ( w_4318 ,  , w_4319 );
buf ( w_4317 , \1965_b1 );
not ( w_4317 , w_4320 );
not (  , w_4321 );
and ( w_4320 , w_4321 , \1965_b0 );
or ( \1967_b1 , \1966_b1 , w_4322 );
xor ( \1967_b0 , \1966_b0 , w_4324 );
not ( w_4324 , w_4325 );
and ( w_4325 , w_4322 , w_4323 );
buf ( w_4322 , \1363_b1 );
not ( w_4322 , w_4326 );
not ( w_4323 , w_4327 );
and ( w_4326 , w_4327 , \1363_b0 );
or ( \1968_b1 , \1962_b1 , \1967_b1 );
not ( \1967_b1 , w_4328 );
and ( \1968_b0 , \1962_b0 , w_4329 );
and ( w_4328 , w_4329 , \1967_b0 );
or ( \1969_b1 , \1958_b1 , \1967_b1 );
not ( \1967_b1 , w_4330 );
and ( \1969_b0 , \1958_b0 , w_4331 );
and ( w_4330 , w_4331 , \1967_b0 );
or ( \1971_b1 , \343_b1 , \1280_b1 );
not ( \1280_b1 , w_4332 );
and ( \1971_b0 , \343_b0 , w_4333 );
and ( w_4332 , w_4333 , \1280_b0 );
or ( \1972_b1 , \353_b1 , \1278_b1 );
not ( \1278_b1 , w_4334 );
and ( \1972_b0 , \353_b0 , w_4335 );
and ( w_4334 , w_4335 , \1278_b0 );
or ( \1973_b1 , \1971_b1 , w_4337 );
not ( w_4337 , w_4338 );
and ( \1973_b0 , \1971_b0 , w_4339 );
and ( w_4338 ,  , w_4339 );
buf ( w_4337 , \1972_b1 );
not ( w_4337 , w_4340 );
not (  , w_4341 );
and ( w_4340 , w_4341 , \1972_b0 );
or ( \1974_b1 , \1973_b1 , w_4342 );
xor ( \1974_b0 , \1973_b0 , w_4344 );
not ( w_4344 , w_4345 );
and ( w_4345 , w_4342 , w_4343 );
buf ( w_4342 , \1177_b1 );
not ( w_4342 , w_4346 );
not ( w_4343 , w_4347 );
and ( w_4346 , w_4347 , \1177_b0 );
or ( \1975_b1 , \444_b1 , \1062_b1 );
not ( \1062_b1 , w_4348 );
and ( \1975_b0 , \444_b0 , w_4349 );
and ( w_4348 , w_4349 , \1062_b0 );
or ( \1976_b1 , \360_b1 , \1060_b1 );
not ( \1060_b1 , w_4350 );
and ( \1976_b0 , \360_b0 , w_4351 );
and ( w_4350 , w_4351 , \1060_b0 );
or ( \1977_b1 , \1975_b1 , w_4353 );
not ( w_4353 , w_4354 );
and ( \1977_b0 , \1975_b0 , w_4355 );
and ( w_4354 ,  , w_4355 );
buf ( w_4353 , \1976_b1 );
not ( w_4353 , w_4356 );
not (  , w_4357 );
and ( w_4356 , w_4357 , \1976_b0 );
or ( \1978_b1 , \1977_b1 , w_4358 );
xor ( \1978_b0 , \1977_b0 , w_4360 );
not ( w_4360 , w_4361 );
and ( w_4361 , w_4358 , w_4359 );
buf ( w_4358 , \984_b1 );
not ( w_4358 , w_4362 );
not ( w_4359 , w_4363 );
and ( w_4362 , w_4363 , \984_b0 );
or ( \1979_b1 , \1974_b1 , \1978_b1 );
not ( \1978_b1 , w_4364 );
and ( \1979_b0 , \1974_b0 , w_4365 );
and ( w_4364 , w_4365 , \1978_b0 );
or ( \1980_b1 , \593_b1 , \912_b1 );
not ( \912_b1 , w_4366 );
and ( \1980_b0 , \593_b0 , w_4367 );
and ( w_4366 , w_4367 , \912_b0 );
or ( \1981_b1 , \495_b1 , \910_b1 );
not ( \910_b1 , w_4368 );
and ( \1981_b0 , \495_b0 , w_4369 );
and ( w_4368 , w_4369 , \910_b0 );
or ( \1982_b1 , \1980_b1 , w_4371 );
not ( w_4371 , w_4372 );
and ( \1982_b0 , \1980_b0 , w_4373 );
and ( w_4372 ,  , w_4373 );
buf ( w_4371 , \1981_b1 );
not ( w_4371 , w_4374 );
not (  , w_4375 );
and ( w_4374 , w_4375 , \1981_b0 );
or ( \1983_b1 , \1982_b1 , w_4376 );
xor ( \1983_b0 , \1982_b0 , w_4378 );
not ( w_4378 , w_4379 );
and ( w_4379 , w_4376 , w_4377 );
buf ( w_4376 , \818_b1 );
not ( w_4376 , w_4380 );
not ( w_4377 , w_4381 );
and ( w_4380 , w_4381 , \818_b0 );
or ( \1984_b1 , \1978_b1 , \1983_b1 );
not ( \1983_b1 , w_4382 );
and ( \1984_b0 , \1978_b0 , w_4383 );
and ( w_4382 , w_4383 , \1983_b0 );
or ( \1985_b1 , \1974_b1 , \1983_b1 );
not ( \1983_b1 , w_4384 );
and ( \1985_b0 , \1974_b0 , w_4385 );
and ( w_4384 , w_4385 , \1983_b0 );
or ( \1987_b1 , \1970_b1 , \1986_b1 );
not ( \1986_b1 , w_4386 );
and ( \1987_b0 , \1970_b0 , w_4387 );
and ( w_4386 , w_4387 , \1986_b0 );
or ( \1988_b1 , \703_b1 , \740_b1 );
not ( \740_b1 , w_4388 );
and ( \1988_b0 , \703_b0 , w_4389 );
and ( w_4388 , w_4389 , \740_b0 );
or ( \1989_b1 , \621_b1 , \738_b1 );
not ( \738_b1 , w_4390 );
and ( \1989_b0 , \621_b0 , w_4391 );
and ( w_4390 , w_4391 , \738_b0 );
or ( \1990_b1 , \1988_b1 , w_4393 );
not ( w_4393 , w_4394 );
and ( \1990_b0 , \1988_b0 , w_4395 );
and ( w_4394 ,  , w_4395 );
buf ( w_4393 , \1989_b1 );
not ( w_4393 , w_4396 );
not (  , w_4397 );
and ( w_4396 , w_4397 , \1989_b0 );
or ( \1991_b1 , \1990_b1 , w_4398 );
xor ( \1991_b0 , \1990_b0 , w_4400 );
not ( w_4400 , w_4401 );
and ( w_4401 , w_4398 , w_4399 );
buf ( w_4398 , \668_b1 );
not ( w_4398 , w_4402 );
not ( w_4399 , w_4403 );
and ( w_4402 , w_4403 , \668_b0 );
or ( \1992_b1 , \841_b1 , \604_b1 );
not ( \604_b1 , w_4404 );
and ( \1992_b0 , \841_b0 , w_4405 );
and ( w_4404 , w_4405 , \604_b0 );
or ( \1993_b1 , \777_b1 , \602_b1 );
not ( \602_b1 , w_4406 );
and ( \1993_b0 , \777_b0 , w_4407 );
and ( w_4406 , w_4407 , \602_b0 );
or ( \1994_b1 , \1992_b1 , w_4409 );
not ( w_4409 , w_4410 );
and ( \1994_b0 , \1992_b0 , w_4411 );
and ( w_4410 ,  , w_4411 );
buf ( w_4409 , \1993_b1 );
not ( w_4409 , w_4412 );
not (  , w_4413 );
and ( w_4412 , w_4413 , \1993_b0 );
or ( \1995_b1 , \1994_b1 , w_4414 );
xor ( \1995_b0 , \1994_b0 , w_4416 );
not ( w_4416 , w_4417 );
and ( w_4417 , w_4414 , w_4415 );
buf ( w_4414 , \561_b1 );
not ( w_4414 , w_4418 );
not ( w_4415 , w_4419 );
and ( w_4418 , w_4419 , \561_b0 );
or ( \1996_b1 , \1991_b1 , \1995_b1 );
not ( \1995_b1 , w_4420 );
and ( \1996_b0 , \1991_b0 , w_4421 );
and ( w_4420 , w_4421 , \1995_b0 );
or ( \1997_b1 , \1104_b1 , \503_b1 );
not ( \503_b1 , w_4422 );
and ( \1997_b0 , \1104_b0 , w_4423 );
and ( w_4422 , w_4423 , \503_b0 );
or ( \1998_b1 , \904_b1 , \501_b1 );
not ( \501_b1 , w_4424 );
and ( \1998_b0 , \904_b0 , w_4425 );
and ( w_4424 , w_4425 , \501_b0 );
or ( \1999_b1 , \1997_b1 , w_4427 );
not ( w_4427 , w_4428 );
and ( \1999_b0 , \1997_b0 , w_4429 );
and ( w_4428 ,  , w_4429 );
buf ( w_4427 , \1998_b1 );
not ( w_4427 , w_4430 );
not (  , w_4431 );
and ( w_4430 , w_4431 , \1998_b0 );
or ( \2000_b1 , \1999_b1 , w_4432 );
xor ( \2000_b0 , \1999_b0 , w_4434 );
not ( w_4434 , w_4435 );
and ( w_4435 , w_4432 , w_4433 );
buf ( w_4432 , \455_b1 );
not ( w_4432 , w_4436 );
not ( w_4433 , w_4437 );
and ( w_4436 , w_4437 , \455_b0 );
or ( \2001_b1 , \1995_b1 , \2000_b1 );
not ( \2000_b1 , w_4438 );
and ( \2001_b0 , \1995_b0 , w_4439 );
and ( w_4438 , w_4439 , \2000_b0 );
or ( \2002_b1 , \1991_b1 , \2000_b1 );
not ( \2000_b1 , w_4440 );
and ( \2002_b0 , \1991_b0 , w_4441 );
and ( w_4440 , w_4441 , \2000_b0 );
or ( \2004_b1 , \1986_b1 , \2003_b1 );
not ( \2003_b1 , w_4442 );
and ( \2004_b0 , \1986_b0 , w_4443 );
and ( w_4442 , w_4443 , \2003_b0 );
or ( \2005_b1 , \1970_b1 , \2003_b1 );
not ( \2003_b1 , w_4444 );
and ( \2005_b0 , \1970_b0 , w_4445 );
and ( w_4444 , w_4445 , \2003_b0 );
or ( \2007_b1 , \1299_b1 , \298_b1 );
not ( \298_b1 , w_4446 );
and ( \2007_b0 , \1299_b0 , w_4447 );
and ( w_4446 , w_4447 , \298_b0 );
or ( \2008_b1 , \1194_b1 , \296_b1 );
not ( \296_b1 , w_4448 );
and ( \2008_b0 , \1194_b0 , w_4449 );
and ( w_4448 , w_4449 , \296_b0 );
or ( \2009_b1 , \2007_b1 , w_4451 );
not ( w_4451 , w_4452 );
and ( \2009_b0 , \2007_b0 , w_4453 );
and ( w_4452 ,  , w_4453 );
buf ( w_4451 , \2008_b1 );
not ( w_4451 , w_4454 );
not (  , w_4455 );
and ( w_4454 , w_4455 , \2008_b0 );
or ( \2010_b1 , \2009_b1 , w_4456 );
xor ( \2010_b0 , \2009_b0 , w_4458 );
not ( w_4458 , w_4459 );
and ( w_4459 , w_4456 , w_4457 );
buf ( w_4456 , \303_b1 );
not ( w_4456 , w_4460 );
not ( w_4457 , w_4461 );
and ( w_4460 , w_4461 , \303_b0 );
or ( \2011_b1 , \1422_b1 , \313_b1 );
not ( \313_b1 , w_4462 );
and ( \2011_b0 , \1422_b0 , w_4463 );
and ( w_4462 , w_4463 , \313_b0 );
or ( \2012_b1 , \1304_b1 , \311_b1 );
not ( \311_b1 , w_4464 );
and ( \2012_b0 , \1304_b0 , w_4465 );
and ( w_4464 , w_4465 , \311_b0 );
or ( \2013_b1 , \2011_b1 , w_4467 );
not ( w_4467 , w_4468 );
and ( \2013_b0 , \2011_b0 , w_4469 );
and ( w_4468 ,  , w_4469 );
buf ( w_4467 , \2012_b1 );
not ( w_4467 , w_4470 );
not (  , w_4471 );
and ( w_4470 , w_4471 , \2012_b0 );
or ( \2014_b1 , \2013_b1 , w_4472 );
xor ( \2014_b0 , \2013_b0 , w_4474 );
not ( w_4474 , w_4475 );
and ( w_4475 , w_4472 , w_4473 );
buf ( w_4472 , \320_b1 );
not ( w_4472 , w_4476 );
not ( w_4473 , w_4477 );
and ( w_4476 , w_4477 , \320_b0 );
or ( \2015_b1 , \2010_b1 , \2014_b1 );
not ( \2014_b1 , w_4478 );
and ( \2015_b0 , \2010_b0 , w_4479 );
and ( w_4478 , w_4479 , \2014_b0 );
or ( \2016_b1 , \1770_b1 , \331_b1 );
not ( \331_b1 , w_4480 );
and ( \2016_b0 , \1770_b0 , w_4481 );
and ( w_4480 , w_4481 , \331_b0 );
or ( \2017_b1 , \1537_b1 , \329_b1 );
not ( \329_b1 , w_4482 );
and ( \2017_b0 , \1537_b0 , w_4483 );
and ( w_4482 , w_4483 , \329_b0 );
or ( \2018_b1 , \2016_b1 , w_4485 );
not ( w_4485 , w_4486 );
and ( \2018_b0 , \2016_b0 , w_4487 );
and ( w_4486 ,  , w_4487 );
buf ( w_4485 , \2017_b1 );
not ( w_4485 , w_4488 );
not (  , w_4489 );
and ( w_4488 , w_4489 , \2017_b0 );
or ( \2019_b1 , \2018_b1 , w_4490 );
xor ( \2019_b0 , \2018_b0 , w_4492 );
not ( w_4492 , w_4493 );
and ( w_4493 , w_4490 , w_4491 );
buf ( w_4490 , \338_b1 );
not ( w_4490 , w_4494 );
not ( w_4491 , w_4495 );
and ( w_4494 , w_4495 , \338_b0 );
or ( \2020_b1 , \2014_b1 , \2019_b1 );
not ( \2019_b1 , w_4496 );
and ( \2020_b0 , \2014_b0 , w_4497 );
and ( w_4496 , w_4497 , \2019_b0 );
or ( \2021_b1 , \2010_b1 , \2019_b1 );
not ( \2019_b1 , w_4498 );
and ( \2021_b0 , \2010_b0 , w_4499 );
and ( w_4498 , w_4499 , \2019_b0 );
buf ( \2023_b1 , RIb4beef8_89_b1 );
buf ( \2023_b0 , RIb4beef8_89_b0 );
or ( \2024_b1 , \2023_b1 , \351_b1 );
not ( \351_b1 , w_4500 );
and ( \2024_b0 , \2023_b0 , w_4501 );
and ( w_4500 , w_4501 , \351_b0 );
or ( \2025_b1 , \1778_b1 , \349_b1 );
not ( \349_b1 , w_4502 );
and ( \2025_b0 , \1778_b0 , w_4503 );
and ( w_4502 , w_4503 , \349_b0 );
or ( \2026_b1 , \2024_b1 , w_4505 );
not ( w_4505 , w_4506 );
and ( \2026_b0 , \2024_b0 , w_4507 );
and ( w_4506 ,  , w_4507 );
buf ( w_4505 , \2025_b1 );
not ( w_4505 , w_4508 );
not (  , w_4509 );
and ( w_4508 , w_4509 , \2025_b0 );
or ( \2027_b1 , \2026_b1 , w_4510 );
xor ( \2027_b0 , \2026_b0 , w_4512 );
not ( w_4512 , w_4513 );
and ( w_4513 , w_4510 , w_4511 );
buf ( w_4510 , \358_b1 );
not ( w_4510 , w_4514 );
not ( w_4511 , w_4515 );
and ( w_4514 , w_4515 , \358_b0 );
buf ( \2028_b1 , RIb4bee80_90_b1 );
buf ( \2028_b0 , RIb4bee80_90_b0 );
or ( \2029_b1 , \2028_b1 , \345_b1 );
not ( \345_b1 , w_4516 );
and ( \2029_b0 , \2028_b0 , w_4517 );
and ( w_4516 , w_4517 , \345_b0 );
or ( \2030_b1 , \2027_b1 , w_4518 );
or ( \2030_b0 , \2027_b0 , \2029_b0 );
not ( \2029_b0 , w_4519 );
and ( w_4519 , w_4518 , \2029_b1 );
or ( \2031_b1 , \2022_b1 , \2030_b1 );
not ( \2030_b1 , w_4520 );
and ( \2031_b0 , \2022_b0 , w_4521 );
and ( w_4520 , w_4521 , \2030_b0 );
or ( \2032_b1 , \1778_b1 , \351_b1 );
not ( \351_b1 , w_4522 );
and ( \2032_b0 , \1778_b0 , w_4523 );
and ( w_4522 , w_4523 , \351_b0 );
or ( \2033_b1 , \1770_b1 , \349_b1 );
not ( \349_b1 , w_4524 );
and ( \2033_b0 , \1770_b0 , w_4525 );
and ( w_4524 , w_4525 , \349_b0 );
or ( \2034_b1 , \2032_b1 , w_4527 );
not ( w_4527 , w_4528 );
and ( \2034_b0 , \2032_b0 , w_4529 );
and ( w_4528 ,  , w_4529 );
buf ( w_4527 , \2033_b1 );
not ( w_4527 , w_4530 );
not (  , w_4531 );
and ( w_4530 , w_4531 , \2033_b0 );
or ( \2035_b1 , \2034_b1 , w_4532 );
xor ( \2035_b0 , \2034_b0 , w_4534 );
not ( w_4534 , w_4535 );
and ( w_4535 , w_4532 , w_4533 );
buf ( w_4532 , \358_b1 );
not ( w_4532 , w_4536 );
not ( w_4533 , w_4537 );
and ( w_4536 , w_4537 , \358_b0 );
or ( \2036_b1 , \2030_b1 , \2035_b1 );
not ( \2035_b1 , w_4538 );
and ( \2036_b0 , \2030_b0 , w_4539 );
and ( w_4538 , w_4539 , \2035_b0 );
or ( \2037_b1 , \2022_b1 , \2035_b1 );
not ( \2035_b1 , w_4540 );
and ( \2037_b0 , \2022_b0 , w_4541 );
and ( w_4540 , w_4541 , \2035_b0 );
or ( \2039_b1 , \2006_b1 , \2038_b1 );
not ( \2038_b1 , w_4542 );
and ( \2039_b0 , \2006_b0 , w_4543 );
and ( w_4542 , w_4543 , \2038_b0 );
or ( \2040_b1 , \2023_b1 , \345_b1 );
not ( \345_b1 , w_4544 );
and ( \2040_b0 , \2023_b0 , w_4545 );
and ( w_4544 , w_4545 , \345_b0 );
or ( \2041_b1 , \1899_b1 , \1903_b1 );
xor ( \2041_b0 , \1899_b0 , w_4546 );
not ( w_4546 , w_4547 );
and ( w_4547 , \1903_b1 , \1903_b0 );
or ( \2042_b1 , \2041_b1 , \1908_b1 );
xor ( \2042_b0 , \2041_b0 , w_4548 );
not ( w_4548 , w_4549 );
and ( w_4549 , \1908_b1 , \1908_b0 );
or ( \2043_b1 , \2040_b1 , \2042_b1 );
not ( \2042_b1 , w_4550 );
and ( \2043_b0 , \2040_b0 , w_4551 );
and ( w_4550 , w_4551 , \2042_b0 );
or ( \2044_b1 , \1869_b1 , \1873_b1 );
xor ( \2044_b0 , \1869_b0 , w_4552 );
not ( w_4552 , w_4553 );
and ( w_4553 , \1873_b1 , \1873_b0 );
or ( \2045_b1 , \2044_b1 , \1878_b1 );
xor ( \2045_b0 , \2044_b0 , w_4554 );
not ( w_4554 , w_4555 );
and ( w_4555 , \1878_b1 , \1878_b0 );
or ( \2046_b1 , \2042_b1 , \2045_b1 );
not ( \2045_b1 , w_4556 );
and ( \2046_b0 , \2042_b0 , w_4557 );
and ( w_4556 , w_4557 , \2045_b0 );
or ( \2047_b1 , \2040_b1 , \2045_b1 );
not ( \2045_b1 , w_4558 );
and ( \2047_b0 , \2040_b0 , w_4559 );
and ( w_4558 , w_4559 , \2045_b0 );
or ( \2049_b1 , \2038_b1 , \2048_b1 );
not ( \2048_b1 , w_4560 );
and ( \2049_b0 , \2038_b0 , w_4561 );
and ( w_4560 , w_4561 , \2048_b0 );
or ( \2050_b1 , \2006_b1 , \2048_b1 );
not ( \2048_b1 , w_4562 );
and ( \2050_b0 , \2006_b0 , w_4563 );
and ( w_4562 , w_4563 , \2048_b0 );
or ( \2052_b1 , \1848_b1 , \1864_b1 );
xor ( \2052_b0 , \1848_b0 , w_4564 );
not ( w_4564 , w_4565 );
and ( w_4565 , \1864_b1 , \1864_b0 );
or ( \2053_b1 , \2052_b1 , \1881_b1 );
xor ( \2053_b0 , \2052_b0 , w_4566 );
not ( w_4566 , w_4567 );
and ( w_4567 , \1881_b1 , \1881_b0 );
or ( \2054_b1 , \1886_b1 , \1888_b1 );
xor ( \2054_b0 , \1886_b0 , w_4568 );
not ( w_4568 , w_4569 );
and ( w_4569 , \1888_b1 , \1888_b0 );
or ( \2055_b1 , \2054_b1 , \1891_b1 );
xor ( \2055_b0 , \2054_b0 , w_4570 );
not ( w_4570 , w_4571 );
and ( w_4571 , \1891_b1 , \1891_b0 );
or ( \2056_b1 , \2053_b1 , \2055_b1 );
not ( \2055_b1 , w_4572 );
and ( \2056_b0 , \2053_b0 , w_4573 );
and ( w_4572 , w_4573 , \2055_b0 );
or ( \2057_b1 , \1911_b1 , \1913_b1 );
xor ( \2057_b0 , \1911_b0 , w_4574 );
not ( w_4574 , w_4575 );
and ( w_4575 , \1913_b1 , \1913_b0 );
or ( \2058_b1 , \2057_b1 , \1915_b1 );
xor ( \2058_b0 , \2057_b0 , w_4576 );
not ( w_4576 , w_4577 );
and ( w_4577 , \1915_b1 , \1915_b0 );
or ( \2059_b1 , \2055_b1 , \2058_b1 );
not ( \2058_b1 , w_4578 );
and ( \2059_b0 , \2055_b0 , w_4579 );
and ( w_4578 , w_4579 , \2058_b0 );
or ( \2060_b1 , \2053_b1 , \2058_b1 );
not ( \2058_b1 , w_4580 );
and ( \2060_b0 , \2053_b0 , w_4581 );
and ( w_4580 , w_4581 , \2058_b0 );
or ( \2062_b1 , \2051_b1 , \2061_b1 );
not ( \2061_b1 , w_4582 );
and ( \2062_b0 , \2051_b0 , w_4583 );
and ( w_4582 , w_4583 , \2061_b0 );
or ( \2063_b1 , \1721_b1 , \1737_b1 );
xor ( \2063_b0 , \1721_b0 , w_4584 );
not ( w_4584 , w_4585 );
and ( w_4585 , \1737_b1 , \1737_b0 );
or ( \2064_b1 , \2063_b1 , \1757_b1 );
xor ( \2064_b0 , \2063_b0 , w_4586 );
not ( w_4586 , w_4587 );
and ( w_4587 , \1757_b1 , \1757_b0 );
or ( \2065_b1 , \2061_b1 , \2064_b1 );
not ( \2064_b1 , w_4588 );
and ( \2065_b0 , \2061_b0 , w_4589 );
and ( w_4588 , w_4589 , \2064_b0 );
or ( \2066_b1 , \2051_b1 , \2064_b1 );
not ( \2064_b1 , w_4590 );
and ( \2066_b0 , \2051_b0 , w_4591 );
and ( w_4590 , w_4591 , \2064_b0 );
or ( \2068_b1 , \1884_b1 , \1894_b1 );
xor ( \2068_b0 , \1884_b0 , w_4592 );
not ( w_4592 , w_4593 );
and ( w_4593 , \1894_b1 , \1894_b0 );
or ( \2069_b1 , \2068_b1 , \1918_b1 );
xor ( \2069_b0 , \2068_b0 , w_4594 );
not ( w_4594 , w_4595 );
and ( w_4595 , \1918_b1 , \1918_b0 );
or ( \2070_b1 , \1923_b1 , \1925_b1 );
xor ( \2070_b0 , \1923_b0 , w_4596 );
not ( w_4596 , w_4597 );
and ( w_4597 , \1925_b1 , \1925_b0 );
or ( \2071_b1 , \2070_b1 , \1928_b1 );
xor ( \2071_b0 , \2070_b0 , w_4598 );
not ( w_4598 , w_4599 );
and ( w_4599 , \1928_b1 , \1928_b0 );
or ( \2072_b1 , \2069_b1 , \2071_b1 );
not ( \2071_b1 , w_4600 );
and ( \2072_b0 , \2069_b0 , w_4601 );
and ( w_4600 , w_4601 , \2071_b0 );
or ( \2073_b1 , \2067_b1 , \2072_b1 );
not ( \2072_b1 , w_4602 );
and ( \2073_b0 , \2067_b0 , w_4603 );
and ( w_4602 , w_4603 , \2072_b0 );
or ( \2074_b1 , \1760_b1 , \1785_b1 );
xor ( \2074_b0 , \1760_b0 , w_4604 );
not ( w_4604 , w_4605 );
and ( w_4605 , \1785_b1 , \1785_b0 );
or ( \2075_b1 , \2074_b1 , \1796_b1 );
xor ( \2075_b0 , \2074_b0 , w_4606 );
not ( w_4606 , w_4607 );
and ( w_4607 , \1796_b1 , \1796_b0 );
or ( \2076_b1 , \2072_b1 , \2075_b1 );
not ( \2075_b1 , w_4608 );
and ( \2076_b0 , \2072_b0 , w_4609 );
and ( w_4608 , w_4609 , \2075_b0 );
or ( \2077_b1 , \2067_b1 , \2075_b1 );
not ( \2075_b1 , w_4610 );
and ( \2077_b0 , \2067_b0 , w_4611 );
and ( w_4610 , w_4611 , \2075_b0 );
or ( \2079_b1 , \1937_b1 , \1939_b1 );
xor ( \2079_b0 , \1937_b0 , w_4612 );
not ( w_4612 , w_4613 );
and ( w_4613 , \1939_b1 , \1939_b0 );
or ( \2080_b1 , \2079_b1 , \1942_b1 );
xor ( \2080_b0 , \2079_b0 , w_4614 );
not ( w_4614 , w_4615 );
and ( w_4615 , \1942_b1 , \1942_b0 );
or ( \2081_b1 , \2078_b1 , \2080_b1 );
not ( \2080_b1 , w_4616 );
and ( \2081_b0 , \2078_b0 , w_4617 );
and ( w_4616 , w_4617 , \2080_b0 );
or ( \2082_b1 , \1951_b1 , \2081_b1 );
not ( \2081_b1 , w_4618 );
and ( \2082_b0 , \1951_b0 , w_4619 );
and ( w_4618 , w_4619 , \2081_b0 );
or ( \2083_b1 , \1951_b1 , \2081_b1 );
xor ( \2083_b0 , \1951_b0 , w_4620 );
not ( w_4620 , w_4621 );
and ( w_4621 , \2081_b1 , \2081_b0 );
or ( \2084_b1 , \2078_b1 , \2080_b1 );
xor ( \2084_b0 , \2078_b0 , w_4622 );
not ( w_4622 , w_4623 );
and ( w_4623 , \2080_b1 , \2080_b0 );
or ( \2085_b1 , \621_b1 , \912_b1 );
not ( \912_b1 , w_4624 );
and ( \2085_b0 , \621_b0 , w_4625 );
and ( w_4624 , w_4625 , \912_b0 );
or ( \2086_b1 , \593_b1 , \910_b1 );
not ( \910_b1 , w_4626 );
and ( \2086_b0 , \593_b0 , w_4627 );
and ( w_4626 , w_4627 , \910_b0 );
or ( \2087_b1 , \2085_b1 , w_4629 );
not ( w_4629 , w_4630 );
and ( \2087_b0 , \2085_b0 , w_4631 );
and ( w_4630 ,  , w_4631 );
buf ( w_4629 , \2086_b1 );
not ( w_4629 , w_4632 );
not (  , w_4633 );
and ( w_4632 , w_4633 , \2086_b0 );
or ( \2088_b1 , \2087_b1 , w_4634 );
xor ( \2088_b0 , \2087_b0 , w_4636 );
not ( w_4636 , w_4637 );
and ( w_4637 , w_4634 , w_4635 );
buf ( w_4634 , \818_b1 );
not ( w_4634 , w_4638 );
not ( w_4635 , w_4639 );
and ( w_4638 , w_4639 , \818_b0 );
or ( \2089_b1 , \777_b1 , \740_b1 );
not ( \740_b1 , w_4640 );
and ( \2089_b0 , \777_b0 , w_4641 );
and ( w_4640 , w_4641 , \740_b0 );
or ( \2090_b1 , \703_b1 , \738_b1 );
not ( \738_b1 , w_4642 );
and ( \2090_b0 , \703_b0 , w_4643 );
and ( w_4642 , w_4643 , \738_b0 );
or ( \2091_b1 , \2089_b1 , w_4645 );
not ( w_4645 , w_4646 );
and ( \2091_b0 , \2089_b0 , w_4647 );
and ( w_4646 ,  , w_4647 );
buf ( w_4645 , \2090_b1 );
not ( w_4645 , w_4648 );
not (  , w_4649 );
and ( w_4648 , w_4649 , \2090_b0 );
or ( \2092_b1 , \2091_b1 , w_4650 );
xor ( \2092_b0 , \2091_b0 , w_4652 );
not ( w_4652 , w_4653 );
and ( w_4653 , w_4650 , w_4651 );
buf ( w_4650 , \668_b1 );
not ( w_4650 , w_4654 );
not ( w_4651 , w_4655 );
and ( w_4654 , w_4655 , \668_b0 );
or ( \2093_b1 , \2088_b1 , \2092_b1 );
not ( \2092_b1 , w_4656 );
and ( \2093_b0 , \2088_b0 , w_4657 );
and ( w_4656 , w_4657 , \2092_b0 );
or ( \2094_b1 , \904_b1 , \604_b1 );
not ( \604_b1 , w_4658 );
and ( \2094_b0 , \904_b0 , w_4659 );
and ( w_4658 , w_4659 , \604_b0 );
or ( \2095_b1 , \841_b1 , \602_b1 );
not ( \602_b1 , w_4660 );
and ( \2095_b0 , \841_b0 , w_4661 );
and ( w_4660 , w_4661 , \602_b0 );
or ( \2096_b1 , \2094_b1 , w_4663 );
not ( w_4663 , w_4664 );
and ( \2096_b0 , \2094_b0 , w_4665 );
and ( w_4664 ,  , w_4665 );
buf ( w_4663 , \2095_b1 );
not ( w_4663 , w_4666 );
not (  , w_4667 );
and ( w_4666 , w_4667 , \2095_b0 );
or ( \2097_b1 , \2096_b1 , w_4668 );
xor ( \2097_b0 , \2096_b0 , w_4670 );
not ( w_4670 , w_4671 );
and ( w_4671 , w_4668 , w_4669 );
buf ( w_4668 , \561_b1 );
not ( w_4668 , w_4672 );
not ( w_4669 , w_4673 );
and ( w_4672 , w_4673 , \561_b0 );
or ( \2098_b1 , \2092_b1 , \2097_b1 );
not ( \2097_b1 , w_4674 );
and ( \2098_b0 , \2092_b0 , w_4675 );
and ( w_4674 , w_4675 , \2097_b0 );
or ( \2099_b1 , \2088_b1 , \2097_b1 );
not ( \2097_b1 , w_4676 );
and ( \2099_b0 , \2088_b0 , w_4677 );
and ( w_4676 , w_4677 , \2097_b0 );
or ( \2101_b1 , \353_b1 , \1476_b1 );
not ( \1476_b1 , w_4678 );
and ( \2101_b0 , \353_b0 , w_4679 );
and ( w_4678 , w_4679 , \1476_b0 );
or ( \2102_b1 , \323_b1 , \1474_b1 );
not ( \1474_b1 , w_4680 );
and ( \2102_b0 , \323_b0 , w_4681 );
and ( w_4680 , w_4681 , \1474_b0 );
or ( \2103_b1 , \2101_b1 , w_4683 );
not ( w_4683 , w_4684 );
and ( \2103_b0 , \2101_b0 , w_4685 );
and ( w_4684 ,  , w_4685 );
buf ( w_4683 , \2102_b1 );
not ( w_4683 , w_4686 );
not (  , w_4687 );
and ( w_4686 , w_4687 , \2102_b0 );
or ( \2104_b1 , \2103_b1 , w_4688 );
xor ( \2104_b0 , \2103_b0 , w_4690 );
not ( w_4690 , w_4691 );
and ( w_4691 , w_4688 , w_4689 );
buf ( w_4688 , \1363_b1 );
not ( w_4688 , w_4692 );
not ( w_4689 , w_4693 );
and ( w_4692 , w_4693 , \1363_b0 );
or ( \2105_b1 , \360_b1 , \1280_b1 );
not ( \1280_b1 , w_4694 );
and ( \2105_b0 , \360_b0 , w_4695 );
and ( w_4694 , w_4695 , \1280_b0 );
or ( \2106_b1 , \343_b1 , \1278_b1 );
not ( \1278_b1 , w_4696 );
and ( \2106_b0 , \343_b0 , w_4697 );
and ( w_4696 , w_4697 , \1278_b0 );
or ( \2107_b1 , \2105_b1 , w_4699 );
not ( w_4699 , w_4700 );
and ( \2107_b0 , \2105_b0 , w_4701 );
and ( w_4700 ,  , w_4701 );
buf ( w_4699 , \2106_b1 );
not ( w_4699 , w_4702 );
not (  , w_4703 );
and ( w_4702 , w_4703 , \2106_b0 );
or ( \2108_b1 , \2107_b1 , w_4704 );
xor ( \2108_b0 , \2107_b0 , w_4706 );
not ( w_4706 , w_4707 );
and ( w_4707 , w_4704 , w_4705 );
buf ( w_4704 , \1177_b1 );
not ( w_4704 , w_4708 );
not ( w_4705 , w_4709 );
and ( w_4708 , w_4709 , \1177_b0 );
or ( \2109_b1 , \2104_b1 , \2108_b1 );
not ( \2108_b1 , w_4710 );
and ( \2109_b0 , \2104_b0 , w_4711 );
and ( w_4710 , w_4711 , \2108_b0 );
or ( \2110_b1 , \495_b1 , \1062_b1 );
not ( \1062_b1 , w_4712 );
and ( \2110_b0 , \495_b0 , w_4713 );
and ( w_4712 , w_4713 , \1062_b0 );
or ( \2111_b1 , \444_b1 , \1060_b1 );
not ( \1060_b1 , w_4714 );
and ( \2111_b0 , \444_b0 , w_4715 );
and ( w_4714 , w_4715 , \1060_b0 );
or ( \2112_b1 , \2110_b1 , w_4717 );
not ( w_4717 , w_4718 );
and ( \2112_b0 , \2110_b0 , w_4719 );
and ( w_4718 ,  , w_4719 );
buf ( w_4717 , \2111_b1 );
not ( w_4717 , w_4720 );
not (  , w_4721 );
and ( w_4720 , w_4721 , \2111_b0 );
or ( \2113_b1 , \2112_b1 , w_4722 );
xor ( \2113_b0 , \2112_b0 , w_4724 );
not ( w_4724 , w_4725 );
and ( w_4725 , w_4722 , w_4723 );
buf ( w_4722 , \984_b1 );
not ( w_4722 , w_4726 );
not ( w_4723 , w_4727 );
and ( w_4726 , w_4727 , \984_b0 );
or ( \2114_b1 , \2108_b1 , \2113_b1 );
not ( \2113_b1 , w_4728 );
and ( \2114_b0 , \2108_b0 , w_4729 );
and ( w_4728 , w_4729 , \2113_b0 );
or ( \2115_b1 , \2104_b1 , \2113_b1 );
not ( \2113_b1 , w_4730 );
and ( \2115_b0 , \2104_b0 , w_4731 );
and ( w_4730 , w_4731 , \2113_b0 );
or ( \2117_b1 , \2100_b1 , \2116_b1 );
not ( \2116_b1 , w_4732 );
and ( \2117_b0 , \2100_b0 , w_4733 );
and ( w_4732 , w_4733 , \2116_b0 );
and ( \2118_nR128_b1 , RIb4c2c60_60_b1 , w_4734 );
xor ( w_4734 , RIb4c2c60_60_b0 , \288_b1 );
not ( \288_b1 , w_4735 );
and ( \2118_nR128_b0 , w_4735 , \288_b0 );
buf ( \2119_b1 , \2118_nR128_b1 );
buf ( \2119_b0 , \2118_nR128_b0 );
and ( \2120_nR127_b1 , RIb4c2be8_61_b1 , w_4736 );
xor ( w_4736 , RIb4c2be8_61_b0 , \288_b1 );
not ( \288_b1 , w_4737 );
and ( \2120_nR127_b0 , w_4737 , \288_b0 );
buf ( \2121_b1 , \2120_nR127_b1 );
buf ( \2121_b0 , \2120_nR127_b0 );
or ( \2122_b1 , \2119_b1 , \2121_b1 );
not ( \2121_b1 , w_4738 );
and ( \2122_b0 , \2119_b0 , w_4739 );
and ( w_4738 , w_4739 , \2121_b0 );
buf ( \2123_b1 , \2122_b1 );
not ( \2123_b1 , w_4740 );
not ( \2123_b0 , w_4741 );
and ( w_4740 , w_4741 , \2122_b0 );
or ( \2124_b1 , \1832_b1 , \2123_b1 );
not ( \2123_b1 , w_4742 );
and ( \2124_b0 , \1832_b0 , w_4743 );
and ( w_4742 , w_4743 , \2123_b0 );
buf ( \2125_b1 , \2124_b1 );
not ( \2125_b1 , w_4744 );
not ( \2125_b0 , w_4745 );
and ( w_4744 , w_4745 , \2124_b0 );
or ( \2126_b1 , \315_b1 , \1955_b1 );
not ( \1955_b1 , w_4746 );
and ( \2126_b0 , \315_b0 , w_4747 );
and ( w_4746 , w_4747 , \1955_b0 );
or ( \2127_b1 , \159_b1 , \1953_b1 );
not ( \1953_b1 , w_4748 );
and ( \2127_b0 , \159_b0 , w_4749 );
and ( w_4748 , w_4749 , \1953_b0 );
or ( \2128_b1 , \2126_b1 , w_4751 );
not ( w_4751 , w_4752 );
and ( \2128_b0 , \2126_b0 , w_4753 );
and ( w_4752 ,  , w_4753 );
buf ( w_4751 , \2127_b1 );
not ( w_4751 , w_4754 );
not (  , w_4755 );
and ( w_4754 , w_4755 , \2127_b0 );
or ( \2129_b1 , \2128_b1 , w_4756 );
xor ( \2129_b0 , \2128_b0 , w_4758 );
not ( w_4758 , w_4759 );
and ( w_4759 , w_4756 , w_4757 );
buf ( w_4756 , \1835_b1 );
not ( w_4756 , w_4760 );
not ( w_4757 , w_4761 );
and ( w_4760 , w_4761 , \1835_b0 );
or ( \2130_b1 , \2125_b1 , \2129_b1 );
not ( \2129_b1 , w_4762 );
and ( \2130_b0 , \2125_b0 , w_4763 );
and ( w_4762 , w_4763 , \2129_b0 );
or ( \2131_b1 , \333_b1 , \1742_b1 );
not ( \1742_b1 , w_4764 );
and ( \2131_b0 , \333_b0 , w_4765 );
and ( w_4764 , w_4765 , \1742_b0 );
or ( \2132_b1 , \305_b1 , \1740_b1 );
not ( \1740_b1 , w_4766 );
and ( \2132_b0 , \305_b0 , w_4767 );
and ( w_4766 , w_4767 , \1740_b0 );
or ( \2133_b1 , \2131_b1 , w_4769 );
not ( w_4769 , w_4770 );
and ( \2133_b0 , \2131_b0 , w_4771 );
and ( w_4770 ,  , w_4771 );
buf ( w_4769 , \2132_b1 );
not ( w_4769 , w_4772 );
not (  , w_4773 );
and ( w_4772 , w_4773 , \2132_b0 );
or ( \2134_b1 , \2133_b1 , w_4774 );
xor ( \2134_b0 , \2133_b0 , w_4776 );
not ( w_4776 , w_4777 );
and ( w_4777 , w_4774 , w_4775 );
buf ( w_4774 , \1610_b1 );
not ( w_4774 , w_4778 );
not ( w_4775 , w_4779 );
and ( w_4778 , w_4779 , \1610_b0 );
or ( \2135_b1 , \2129_b1 , \2134_b1 );
not ( \2134_b1 , w_4780 );
and ( \2135_b0 , \2129_b0 , w_4781 );
and ( w_4780 , w_4781 , \2134_b0 );
or ( \2136_b1 , \2125_b1 , \2134_b1 );
not ( \2134_b1 , w_4782 );
and ( \2136_b0 , \2125_b0 , w_4783 );
and ( w_4782 , w_4783 , \2134_b0 );
or ( \2138_b1 , \2116_b1 , \2137_b1 );
not ( \2137_b1 , w_4784 );
and ( \2138_b0 , \2116_b0 , w_4785 );
and ( w_4784 , w_4785 , \2137_b0 );
or ( \2139_b1 , \2100_b1 , \2137_b1 );
not ( \2137_b1 , w_4786 );
and ( \2139_b0 , \2100_b0 , w_4787 );
and ( w_4786 , w_4787 , \2137_b0 );
or ( \2141_b1 , \2010_b1 , \2014_b1 );
xor ( \2141_b0 , \2010_b0 , w_4788 );
not ( w_4788 , w_4789 );
and ( w_4789 , \2014_b1 , \2014_b0 );
or ( \2142_b1 , \2141_b1 , \2019_b1 );
xor ( \2142_b0 , \2141_b0 , w_4790 );
not ( w_4790 , w_4791 );
and ( w_4791 , \2019_b1 , \2019_b0 );
or ( \2143_b1 , \1974_b1 , \1978_b1 );
xor ( \2143_b0 , \1974_b0 , w_4792 );
not ( w_4792 , w_4793 );
and ( w_4793 , \1978_b1 , \1978_b0 );
or ( \2144_b1 , \2143_b1 , \1983_b1 );
xor ( \2144_b0 , \2143_b0 , w_4794 );
not ( w_4794 , w_4795 );
and ( w_4795 , \1983_b1 , \1983_b0 );
or ( \2145_b1 , \2142_b1 , \2144_b1 );
not ( \2144_b1 , w_4796 );
and ( \2145_b0 , \2142_b0 , w_4797 );
and ( w_4796 , w_4797 , \2144_b0 );
or ( \2146_b1 , \1991_b1 , \1995_b1 );
xor ( \2146_b0 , \1991_b0 , w_4798 );
not ( w_4798 , w_4799 );
and ( w_4799 , \1995_b1 , \1995_b0 );
or ( \2147_b1 , \2146_b1 , \2000_b1 );
xor ( \2147_b0 , \2146_b0 , w_4800 );
not ( w_4800 , w_4801 );
and ( w_4801 , \2000_b1 , \2000_b0 );
or ( \2148_b1 , \2144_b1 , \2147_b1 );
not ( \2147_b1 , w_4802 );
and ( \2148_b0 , \2144_b0 , w_4803 );
and ( w_4802 , w_4803 , \2147_b0 );
or ( \2149_b1 , \2142_b1 , \2147_b1 );
not ( \2147_b1 , w_4804 );
and ( \2149_b0 , \2142_b0 , w_4805 );
and ( w_4804 , w_4805 , \2147_b0 );
or ( \2151_b1 , \2140_b1 , \2150_b1 );
not ( \2150_b1 , w_4806 );
and ( \2151_b0 , \2140_b0 , w_4807 );
and ( w_4806 , w_4807 , \2150_b0 );
or ( \2152_b1 , \1778_b1 , \331_b1 );
not ( \331_b1 , w_4808 );
and ( \2152_b0 , \1778_b0 , w_4809 );
and ( w_4808 , w_4809 , \331_b0 );
or ( \2153_b1 , \1770_b1 , \329_b1 );
not ( \329_b1 , w_4810 );
and ( \2153_b0 , \1770_b0 , w_4811 );
and ( w_4810 , w_4811 , \329_b0 );
or ( \2154_b1 , \2152_b1 , w_4813 );
not ( w_4813 , w_4814 );
and ( \2154_b0 , \2152_b0 , w_4815 );
and ( w_4814 ,  , w_4815 );
buf ( w_4813 , \2153_b1 );
not ( w_4813 , w_4816 );
not (  , w_4817 );
and ( w_4816 , w_4817 , \2153_b0 );
or ( \2155_b1 , \2154_b1 , w_4818 );
xor ( \2155_b0 , \2154_b0 , w_4820 );
not ( w_4820 , w_4821 );
and ( w_4821 , w_4818 , w_4819 );
buf ( w_4818 , \338_b1 );
not ( w_4818 , w_4822 );
not ( w_4819 , w_4823 );
and ( w_4822 , w_4823 , \338_b0 );
or ( \2156_b1 , \2028_b1 , \351_b1 );
not ( \351_b1 , w_4824 );
and ( \2156_b0 , \2028_b0 , w_4825 );
and ( w_4824 , w_4825 , \351_b0 );
or ( \2157_b1 , \2023_b1 , \349_b1 );
not ( \349_b1 , w_4826 );
and ( \2157_b0 , \2023_b0 , w_4827 );
and ( w_4826 , w_4827 , \349_b0 );
or ( \2158_b1 , \2156_b1 , w_4829 );
not ( w_4829 , w_4830 );
and ( \2158_b0 , \2156_b0 , w_4831 );
and ( w_4830 ,  , w_4831 );
buf ( w_4829 , \2157_b1 );
not ( w_4829 , w_4832 );
not (  , w_4833 );
and ( w_4832 , w_4833 , \2157_b0 );
or ( \2159_b1 , \2158_b1 , w_4834 );
xor ( \2159_b0 , \2158_b0 , w_4836 );
not ( w_4836 , w_4837 );
and ( w_4837 , w_4834 , w_4835 );
buf ( w_4834 , \358_b1 );
not ( w_4834 , w_4838 );
not ( w_4835 , w_4839 );
and ( w_4838 , w_4839 , \358_b0 );
or ( \2160_b1 , \2155_b1 , \2159_b1 );
not ( \2159_b1 , w_4840 );
and ( \2160_b0 , \2155_b0 , w_4841 );
and ( w_4840 , w_4841 , \2159_b0 );
buf ( \2161_b1 , RIb4bc1f8_91_b1 );
buf ( \2161_b0 , RIb4bc1f8_91_b0 );
or ( \2162_b1 , \2161_b1 , \345_b1 );
not ( \345_b1 , w_4842 );
and ( \2162_b0 , \2161_b0 , w_4843 );
and ( w_4842 , w_4843 , \345_b0 );
or ( \2163_b1 , \2159_b1 , \2162_b1 );
not ( \2162_b1 , w_4844 );
and ( \2163_b0 , \2159_b0 , w_4845 );
and ( w_4844 , w_4845 , \2162_b0 );
or ( \2164_b1 , \2155_b1 , \2162_b1 );
not ( \2162_b1 , w_4846 );
and ( \2164_b0 , \2155_b0 , w_4847 );
and ( w_4846 , w_4847 , \2162_b0 );
or ( \2166_b1 , \1194_b1 , \503_b1 );
not ( \503_b1 , w_4848 );
and ( \2166_b0 , \1194_b0 , w_4849 );
and ( w_4848 , w_4849 , \503_b0 );
or ( \2167_b1 , \1104_b1 , \501_b1 );
not ( \501_b1 , w_4850 );
and ( \2167_b0 , \1104_b0 , w_4851 );
and ( w_4850 , w_4851 , \501_b0 );
or ( \2168_b1 , \2166_b1 , w_4853 );
not ( w_4853 , w_4854 );
and ( \2168_b0 , \2166_b0 , w_4855 );
and ( w_4854 ,  , w_4855 );
buf ( w_4853 , \2167_b1 );
not ( w_4853 , w_4856 );
not (  , w_4857 );
and ( w_4856 , w_4857 , \2167_b0 );
or ( \2169_b1 , \2168_b1 , w_4858 );
xor ( \2169_b0 , \2168_b0 , w_4860 );
not ( w_4860 , w_4861 );
and ( w_4861 , w_4858 , w_4859 );
buf ( w_4858 , \455_b1 );
not ( w_4858 , w_4862 );
not ( w_4859 , w_4863 );
and ( w_4862 , w_4863 , \455_b0 );
or ( \2170_b1 , \1304_b1 , \298_b1 );
not ( \298_b1 , w_4864 );
and ( \2170_b0 , \1304_b0 , w_4865 );
and ( w_4864 , w_4865 , \298_b0 );
or ( \2171_b1 , \1299_b1 , \296_b1 );
not ( \296_b1 , w_4866 );
and ( \2171_b0 , \1299_b0 , w_4867 );
and ( w_4866 , w_4867 , \296_b0 );
or ( \2172_b1 , \2170_b1 , w_4869 );
not ( w_4869 , w_4870 );
and ( \2172_b0 , \2170_b0 , w_4871 );
and ( w_4870 ,  , w_4871 );
buf ( w_4869 , \2171_b1 );
not ( w_4869 , w_4872 );
not (  , w_4873 );
and ( w_4872 , w_4873 , \2171_b0 );
or ( \2173_b1 , \2172_b1 , w_4874 );
xor ( \2173_b0 , \2172_b0 , w_4876 );
not ( w_4876 , w_4877 );
and ( w_4877 , w_4874 , w_4875 );
buf ( w_4874 , \303_b1 );
not ( w_4874 , w_4878 );
not ( w_4875 , w_4879 );
and ( w_4878 , w_4879 , \303_b0 );
or ( \2174_b1 , \2169_b1 , \2173_b1 );
not ( \2173_b1 , w_4880 );
and ( \2174_b0 , \2169_b0 , w_4881 );
and ( w_4880 , w_4881 , \2173_b0 );
or ( \2175_b1 , \1537_b1 , \313_b1 );
not ( \313_b1 , w_4882 );
and ( \2175_b0 , \1537_b0 , w_4883 );
and ( w_4882 , w_4883 , \313_b0 );
or ( \2176_b1 , \1422_b1 , \311_b1 );
not ( \311_b1 , w_4884 );
and ( \2176_b0 , \1422_b0 , w_4885 );
and ( w_4884 , w_4885 , \311_b0 );
or ( \2177_b1 , \2175_b1 , w_4887 );
not ( w_4887 , w_4888 );
and ( \2177_b0 , \2175_b0 , w_4889 );
and ( w_4888 ,  , w_4889 );
buf ( w_4887 , \2176_b1 );
not ( w_4887 , w_4890 );
not (  , w_4891 );
and ( w_4890 , w_4891 , \2176_b0 );
or ( \2178_b1 , \2177_b1 , w_4892 );
xor ( \2178_b0 , \2177_b0 , w_4894 );
not ( w_4894 , w_4895 );
and ( w_4895 , w_4892 , w_4893 );
buf ( w_4892 , \320_b1 );
not ( w_4892 , w_4896 );
not ( w_4893 , w_4897 );
and ( w_4896 , w_4897 , \320_b0 );
or ( \2179_b1 , \2173_b1 , \2178_b1 );
not ( \2178_b1 , w_4898 );
and ( \2179_b0 , \2173_b0 , w_4899 );
and ( w_4898 , w_4899 , \2178_b0 );
or ( \2180_b1 , \2169_b1 , \2178_b1 );
not ( \2178_b1 , w_4900 );
and ( \2180_b0 , \2169_b0 , w_4901 );
and ( w_4900 , w_4901 , \2178_b0 );
or ( \2182_b1 , \2165_b1 , \2181_b1 );
not ( \2181_b1 , w_4902 );
and ( \2182_b0 , \2165_b0 , w_4903 );
and ( w_4902 , w_4903 , \2181_b0 );
or ( \2183_b1 , \2027_b1 , w_4904 );
xor ( \2183_b0 , \2027_b0 , w_4906 );
not ( w_4906 , w_4907 );
and ( w_4907 , w_4904 , w_4905 );
buf ( w_4904 , \2029_b1 );
not ( w_4904 , w_4908 );
not ( w_4905 , w_4909 );
and ( w_4908 , w_4909 , \2029_b0 );
or ( \2184_b1 , \2181_b1 , \2183_b1 );
not ( \2183_b1 , w_4910 );
and ( \2184_b0 , \2181_b0 , w_4911 );
and ( w_4910 , w_4911 , \2183_b0 );
or ( \2185_b1 , \2165_b1 , \2183_b1 );
not ( \2183_b1 , w_4912 );
and ( \2185_b0 , \2165_b0 , w_4913 );
and ( w_4912 , w_4913 , \2183_b0 );
or ( \2187_b1 , \2150_b1 , \2186_b1 );
not ( \2186_b1 , w_4914 );
and ( \2187_b0 , \2150_b0 , w_4915 );
and ( w_4914 , w_4915 , \2186_b0 );
or ( \2188_b1 , \2140_b1 , \2186_b1 );
not ( \2186_b1 , w_4916 );
and ( \2188_b0 , \2140_b0 , w_4917 );
and ( w_4916 , w_4917 , \2186_b0 );
or ( \2190_b1 , \1836_b1 , \1840_b1 );
xor ( \2190_b0 , \1836_b0 , w_4918 );
not ( w_4918 , w_4919 );
and ( w_4919 , \1840_b1 , \1840_b0 );
or ( \2191_b1 , \2190_b1 , \1845_b1 );
xor ( \2191_b0 , \2190_b0 , w_4920 );
not ( w_4920 , w_4921 );
and ( w_4921 , \1845_b1 , \1845_b0 );
or ( \2192_b1 , \1852_b1 , \1856_b1 );
xor ( \2192_b0 , \1852_b0 , w_4922 );
not ( w_4922 , w_4923 );
and ( w_4923 , \1856_b1 , \1856_b0 );
or ( \2193_b1 , \2192_b1 , \1861_b1 );
xor ( \2193_b0 , \2192_b0 , w_4924 );
not ( w_4924 , w_4925 );
and ( w_4925 , \1861_b1 , \1861_b0 );
or ( \2194_b1 , \2191_b1 , \2193_b1 );
not ( \2193_b1 , w_4926 );
and ( \2194_b0 , \2191_b0 , w_4927 );
and ( w_4926 , w_4927 , \2193_b0 );
or ( \2195_b1 , \2040_b1 , \2042_b1 );
xor ( \2195_b0 , \2040_b0 , w_4928 );
not ( w_4928 , w_4929 );
and ( w_4929 , \2042_b1 , \2042_b0 );
or ( \2196_b1 , \2195_b1 , \2045_b1 );
xor ( \2196_b0 , \2195_b0 , w_4930 );
not ( w_4930 , w_4931 );
and ( w_4931 , \2045_b1 , \2045_b0 );
or ( \2197_b1 , \2193_b1 , \2196_b1 );
not ( \2196_b1 , w_4932 );
and ( \2197_b0 , \2193_b0 , w_4933 );
and ( w_4932 , w_4933 , \2196_b0 );
or ( \2198_b1 , \2191_b1 , \2196_b1 );
not ( \2196_b1 , w_4934 );
and ( \2198_b0 , \2191_b0 , w_4935 );
and ( w_4934 , w_4935 , \2196_b0 );
or ( \2200_b1 , \2189_b1 , \2199_b1 );
not ( \2199_b1 , w_4936 );
and ( \2200_b0 , \2189_b0 , w_4937 );
and ( w_4936 , w_4937 , \2199_b0 );
or ( \2201_b1 , \2053_b1 , \2055_b1 );
xor ( \2201_b0 , \2053_b0 , w_4938 );
not ( w_4938 , w_4939 );
and ( w_4939 , \2055_b1 , \2055_b0 );
or ( \2202_b1 , \2201_b1 , \2058_b1 );
xor ( \2202_b0 , \2201_b0 , w_4940 );
not ( w_4940 , w_4941 );
and ( w_4941 , \2058_b1 , \2058_b0 );
or ( \2203_b1 , \2199_b1 , \2202_b1 );
not ( \2202_b1 , w_4942 );
and ( \2203_b0 , \2199_b0 , w_4943 );
and ( w_4942 , w_4943 , \2202_b0 );
or ( \2204_b1 , \2189_b1 , \2202_b1 );
not ( \2202_b1 , w_4944 );
and ( \2204_b0 , \2189_b0 , w_4945 );
and ( w_4944 , w_4945 , \2202_b0 );
or ( \2206_b1 , \2051_b1 , \2061_b1 );
xor ( \2206_b0 , \2051_b0 , w_4946 );
not ( w_4946 , w_4947 );
and ( w_4947 , \2061_b1 , \2061_b0 );
or ( \2207_b1 , \2206_b1 , \2064_b1 );
xor ( \2207_b0 , \2206_b0 , w_4948 );
not ( w_4948 , w_4949 );
and ( w_4949 , \2064_b1 , \2064_b0 );
or ( \2208_b1 , \2205_b1 , \2207_b1 );
not ( \2207_b1 , w_4950 );
and ( \2208_b0 , \2205_b0 , w_4951 );
and ( w_4950 , w_4951 , \2207_b0 );
or ( \2209_b1 , \2069_b1 , \2071_b1 );
xor ( \2209_b0 , \2069_b0 , w_4952 );
not ( w_4952 , w_4953 );
and ( w_4953 , \2071_b1 , \2071_b0 );
or ( \2210_b1 , \2207_b1 , \2209_b1 );
not ( \2209_b1 , w_4954 );
and ( \2210_b0 , \2207_b0 , w_4955 );
and ( w_4954 , w_4955 , \2209_b0 );
or ( \2211_b1 , \2205_b1 , \2209_b1 );
not ( \2209_b1 , w_4956 );
and ( \2211_b0 , \2205_b0 , w_4957 );
and ( w_4956 , w_4957 , \2209_b0 );
or ( \2213_b1 , \2067_b1 , \2072_b1 );
xor ( \2213_b0 , \2067_b0 , w_4958 );
not ( w_4958 , w_4959 );
and ( w_4959 , \2072_b1 , \2072_b0 );
or ( \2214_b1 , \2213_b1 , \2075_b1 );
xor ( \2214_b0 , \2213_b0 , w_4960 );
not ( w_4960 , w_4961 );
and ( w_4961 , \2075_b1 , \2075_b0 );
or ( \2215_b1 , \2212_b1 , \2214_b1 );
not ( \2214_b1 , w_4962 );
and ( \2215_b0 , \2212_b0 , w_4963 );
and ( w_4962 , w_4963 , \2214_b0 );
or ( \2216_b1 , \1921_b1 , \1931_b1 );
xor ( \2216_b0 , \1921_b0 , w_4964 );
not ( w_4964 , w_4965 );
and ( w_4965 , \1931_b1 , \1931_b0 );
or ( \2217_b1 , \2216_b1 , \1934_b1 );
xor ( \2217_b0 , \2216_b0 , w_4966 );
not ( w_4966 , w_4967 );
and ( w_4967 , \1934_b1 , \1934_b0 );
or ( \2218_b1 , \2214_b1 , \2217_b1 );
not ( \2217_b1 , w_4968 );
and ( \2218_b0 , \2214_b0 , w_4969 );
and ( w_4968 , w_4969 , \2217_b0 );
or ( \2219_b1 , \2212_b1 , \2217_b1 );
not ( \2217_b1 , w_4970 );
and ( \2219_b0 , \2212_b0 , w_4971 );
and ( w_4970 , w_4971 , \2217_b0 );
or ( \2221_b1 , \2084_b1 , \2220_b1 );
not ( \2220_b1 , w_4972 );
and ( \2221_b0 , \2084_b0 , w_4973 );
and ( w_4972 , w_4973 , \2220_b0 );
or ( \2222_b1 , \2084_b1 , \2220_b1 );
xor ( \2222_b0 , \2084_b0 , w_4974 );
not ( w_4974 , w_4975 );
and ( w_4975 , \2220_b1 , \2220_b0 );
or ( \2223_b1 , \2212_b1 , \2214_b1 );
xor ( \2223_b0 , \2212_b0 , w_4976 );
not ( w_4976 , w_4977 );
and ( w_4977 , \2214_b1 , \2214_b0 );
or ( \2224_b1 , \2223_b1 , \2217_b1 );
xor ( \2224_b0 , \2223_b0 , w_4978 );
not ( w_4978 , w_4979 );
and ( w_4979 , \2217_b1 , \2217_b0 );
or ( \2225_b1 , \703_b1 , \912_b1 );
not ( \912_b1 , w_4980 );
and ( \2225_b0 , \703_b0 , w_4981 );
and ( w_4980 , w_4981 , \912_b0 );
or ( \2226_b1 , \621_b1 , \910_b1 );
not ( \910_b1 , w_4982 );
and ( \2226_b0 , \621_b0 , w_4983 );
and ( w_4982 , w_4983 , \910_b0 );
or ( \2227_b1 , \2225_b1 , w_4985 );
not ( w_4985 , w_4986 );
and ( \2227_b0 , \2225_b0 , w_4987 );
and ( w_4986 ,  , w_4987 );
buf ( w_4985 , \2226_b1 );
not ( w_4985 , w_4988 );
not (  , w_4989 );
and ( w_4988 , w_4989 , \2226_b0 );
or ( \2228_b1 , \2227_b1 , w_4990 );
xor ( \2228_b0 , \2227_b0 , w_4992 );
not ( w_4992 , w_4993 );
and ( w_4993 , w_4990 , w_4991 );
buf ( w_4990 , \818_b1 );
not ( w_4990 , w_4994 );
not ( w_4991 , w_4995 );
and ( w_4994 , w_4995 , \818_b0 );
or ( \2229_b1 , \841_b1 , \740_b1 );
not ( \740_b1 , w_4996 );
and ( \2229_b0 , \841_b0 , w_4997 );
and ( w_4996 , w_4997 , \740_b0 );
or ( \2230_b1 , \777_b1 , \738_b1 );
not ( \738_b1 , w_4998 );
and ( \2230_b0 , \777_b0 , w_4999 );
and ( w_4998 , w_4999 , \738_b0 );
or ( \2231_b1 , \2229_b1 , w_5001 );
not ( w_5001 , w_5002 );
and ( \2231_b0 , \2229_b0 , w_5003 );
and ( w_5002 ,  , w_5003 );
buf ( w_5001 , \2230_b1 );
not ( w_5001 , w_5004 );
not (  , w_5005 );
and ( w_5004 , w_5005 , \2230_b0 );
or ( \2232_b1 , \2231_b1 , w_5006 );
xor ( \2232_b0 , \2231_b0 , w_5008 );
not ( w_5008 , w_5009 );
and ( w_5009 , w_5006 , w_5007 );
buf ( w_5006 , \668_b1 );
not ( w_5006 , w_5010 );
not ( w_5007 , w_5011 );
and ( w_5010 , w_5011 , \668_b0 );
or ( \2233_b1 , \2228_b1 , \2232_b1 );
not ( \2232_b1 , w_5012 );
and ( \2233_b0 , \2228_b0 , w_5013 );
and ( w_5012 , w_5013 , \2232_b0 );
or ( \2234_b1 , \1104_b1 , \604_b1 );
not ( \604_b1 , w_5014 );
and ( \2234_b0 , \1104_b0 , w_5015 );
and ( w_5014 , w_5015 , \604_b0 );
or ( \2235_b1 , \904_b1 , \602_b1 );
not ( \602_b1 , w_5016 );
and ( \2235_b0 , \904_b0 , w_5017 );
and ( w_5016 , w_5017 , \602_b0 );
or ( \2236_b1 , \2234_b1 , w_5019 );
not ( w_5019 , w_5020 );
and ( \2236_b0 , \2234_b0 , w_5021 );
and ( w_5020 ,  , w_5021 );
buf ( w_5019 , \2235_b1 );
not ( w_5019 , w_5022 );
not (  , w_5023 );
and ( w_5022 , w_5023 , \2235_b0 );
or ( \2237_b1 , \2236_b1 , w_5024 );
xor ( \2237_b0 , \2236_b0 , w_5026 );
not ( w_5026 , w_5027 );
and ( w_5027 , w_5024 , w_5025 );
buf ( w_5024 , \561_b1 );
not ( w_5024 , w_5028 );
not ( w_5025 , w_5029 );
and ( w_5028 , w_5029 , \561_b0 );
or ( \2238_b1 , \2232_b1 , \2237_b1 );
not ( \2237_b1 , w_5030 );
and ( \2238_b0 , \2232_b0 , w_5031 );
and ( w_5030 , w_5031 , \2237_b0 );
or ( \2239_b1 , \2228_b1 , \2237_b1 );
not ( \2237_b1 , w_5032 );
and ( \2239_b0 , \2228_b0 , w_5033 );
and ( w_5032 , w_5033 , \2237_b0 );
or ( \2241_b1 , \343_b1 , \1476_b1 );
not ( \1476_b1 , w_5034 );
and ( \2241_b0 , \343_b0 , w_5035 );
and ( w_5034 , w_5035 , \1476_b0 );
or ( \2242_b1 , \353_b1 , \1474_b1 );
not ( \1474_b1 , w_5036 );
and ( \2242_b0 , \353_b0 , w_5037 );
and ( w_5036 , w_5037 , \1474_b0 );
or ( \2243_b1 , \2241_b1 , w_5039 );
not ( w_5039 , w_5040 );
and ( \2243_b0 , \2241_b0 , w_5041 );
and ( w_5040 ,  , w_5041 );
buf ( w_5039 , \2242_b1 );
not ( w_5039 , w_5042 );
not (  , w_5043 );
and ( w_5042 , w_5043 , \2242_b0 );
or ( \2244_b1 , \2243_b1 , w_5044 );
xor ( \2244_b0 , \2243_b0 , w_5046 );
not ( w_5046 , w_5047 );
and ( w_5047 , w_5044 , w_5045 );
buf ( w_5044 , \1363_b1 );
not ( w_5044 , w_5048 );
not ( w_5045 , w_5049 );
and ( w_5048 , w_5049 , \1363_b0 );
or ( \2245_b1 , \444_b1 , \1280_b1 );
not ( \1280_b1 , w_5050 );
and ( \2245_b0 , \444_b0 , w_5051 );
and ( w_5050 , w_5051 , \1280_b0 );
or ( \2246_b1 , \360_b1 , \1278_b1 );
not ( \1278_b1 , w_5052 );
and ( \2246_b0 , \360_b0 , w_5053 );
and ( w_5052 , w_5053 , \1278_b0 );
or ( \2247_b1 , \2245_b1 , w_5055 );
not ( w_5055 , w_5056 );
and ( \2247_b0 , \2245_b0 , w_5057 );
and ( w_5056 ,  , w_5057 );
buf ( w_5055 , \2246_b1 );
not ( w_5055 , w_5058 );
not (  , w_5059 );
and ( w_5058 , w_5059 , \2246_b0 );
or ( \2248_b1 , \2247_b1 , w_5060 );
xor ( \2248_b0 , \2247_b0 , w_5062 );
not ( w_5062 , w_5063 );
and ( w_5063 , w_5060 , w_5061 );
buf ( w_5060 , \1177_b1 );
not ( w_5060 , w_5064 );
not ( w_5061 , w_5065 );
and ( w_5064 , w_5065 , \1177_b0 );
or ( \2249_b1 , \2244_b1 , \2248_b1 );
not ( \2248_b1 , w_5066 );
and ( \2249_b0 , \2244_b0 , w_5067 );
and ( w_5066 , w_5067 , \2248_b0 );
or ( \2250_b1 , \593_b1 , \1062_b1 );
not ( \1062_b1 , w_5068 );
and ( \2250_b0 , \593_b0 , w_5069 );
and ( w_5068 , w_5069 , \1062_b0 );
or ( \2251_b1 , \495_b1 , \1060_b1 );
not ( \1060_b1 , w_5070 );
and ( \2251_b0 , \495_b0 , w_5071 );
and ( w_5070 , w_5071 , \1060_b0 );
or ( \2252_b1 , \2250_b1 , w_5073 );
not ( w_5073 , w_5074 );
and ( \2252_b0 , \2250_b0 , w_5075 );
and ( w_5074 ,  , w_5075 );
buf ( w_5073 , \2251_b1 );
not ( w_5073 , w_5076 );
not (  , w_5077 );
and ( w_5076 , w_5077 , \2251_b0 );
or ( \2253_b1 , \2252_b1 , w_5078 );
xor ( \2253_b0 , \2252_b0 , w_5080 );
not ( w_5080 , w_5081 );
and ( w_5081 , w_5078 , w_5079 );
buf ( w_5078 , \984_b1 );
not ( w_5078 , w_5082 );
not ( w_5079 , w_5083 );
and ( w_5082 , w_5083 , \984_b0 );
or ( \2254_b1 , \2248_b1 , \2253_b1 );
not ( \2253_b1 , w_5084 );
and ( \2254_b0 , \2248_b0 , w_5085 );
and ( w_5084 , w_5085 , \2253_b0 );
or ( \2255_b1 , \2244_b1 , \2253_b1 );
not ( \2253_b1 , w_5086 );
and ( \2255_b0 , \2244_b0 , w_5087 );
and ( w_5086 , w_5087 , \2253_b0 );
or ( \2257_b1 , \2240_b1 , \2256_b1 );
not ( \2256_b1 , w_5088 );
and ( \2257_b0 , \2240_b0 , w_5089 );
and ( w_5088 , w_5089 , \2256_b0 );
or ( \2258_b1 , \1832_b1 , \2119_b1 );
xor ( \2258_b0 , \1832_b0 , w_5090 );
not ( w_5090 , w_5091 );
and ( w_5091 , \2119_b1 , \2119_b0 );
or ( \2259_b1 , \2119_b1 , \2121_b1 );
xor ( \2259_b0 , \2119_b0 , w_5092 );
not ( w_5092 , w_5093 );
and ( w_5093 , \2121_b1 , \2121_b0 );
buf ( \2260_b1 , \2259_b1 );
not ( \2260_b1 , w_5094 );
not ( \2260_b0 , w_5095 );
and ( w_5094 , w_5095 , \2259_b0 );
or ( \2261_b1 , \2258_b1 , \2260_b1 );
not ( \2260_b1 , w_5096 );
and ( \2261_b0 , \2258_b0 , w_5097 );
and ( w_5096 , w_5097 , \2260_b0 );
or ( \2262_b1 , \159_b1 , \2261_b1 );
not ( \2261_b1 , w_5098 );
and ( \2262_b0 , \159_b0 , w_5099 );
and ( w_5098 , w_5099 , \2261_b0 );
buf ( \2263_b1 , \2262_b1 );
not ( \2263_b1 , w_5100 );
not ( \2263_b0 , w_5101 );
and ( w_5100 , w_5101 , \2262_b0 );
or ( \2264_b1 , \2263_b1 , w_5102 );
xor ( \2264_b0 , \2263_b0 , w_5104 );
not ( w_5104 , w_5105 );
and ( w_5105 , w_5102 , w_5103 );
buf ( w_5102 , \2124_b1 );
not ( w_5102 , w_5106 );
not ( w_5103 , w_5107 );
and ( w_5106 , w_5107 , \2124_b0 );
or ( \2265_b1 , \305_b1 , \1955_b1 );
not ( \1955_b1 , w_5108 );
and ( \2265_b0 , \305_b0 , w_5109 );
and ( w_5108 , w_5109 , \1955_b0 );
or ( \2266_b1 , \315_b1 , \1953_b1 );
not ( \1953_b1 , w_5110 );
and ( \2266_b0 , \315_b0 , w_5111 );
and ( w_5110 , w_5111 , \1953_b0 );
or ( \2267_b1 , \2265_b1 , w_5113 );
not ( w_5113 , w_5114 );
and ( \2267_b0 , \2265_b0 , w_5115 );
and ( w_5114 ,  , w_5115 );
buf ( w_5113 , \2266_b1 );
not ( w_5113 , w_5116 );
not (  , w_5117 );
and ( w_5116 , w_5117 , \2266_b0 );
or ( \2268_b1 , \2267_b1 , w_5118 );
xor ( \2268_b0 , \2267_b0 , w_5120 );
not ( w_5120 , w_5121 );
and ( w_5121 , w_5118 , w_5119 );
buf ( w_5118 , \1835_b1 );
not ( w_5118 , w_5122 );
not ( w_5119 , w_5123 );
and ( w_5122 , w_5123 , \1835_b0 );
or ( \2269_b1 , \2264_b1 , \2268_b1 );
not ( \2268_b1 , w_5124 );
and ( \2269_b0 , \2264_b0 , w_5125 );
and ( w_5124 , w_5125 , \2268_b0 );
or ( \2270_b1 , \323_b1 , \1742_b1 );
not ( \1742_b1 , w_5126 );
and ( \2270_b0 , \323_b0 , w_5127 );
and ( w_5126 , w_5127 , \1742_b0 );
or ( \2271_b1 , \333_b1 , \1740_b1 );
not ( \1740_b1 , w_5128 );
and ( \2271_b0 , \333_b0 , w_5129 );
and ( w_5128 , w_5129 , \1740_b0 );
or ( \2272_b1 , \2270_b1 , w_5131 );
not ( w_5131 , w_5132 );
and ( \2272_b0 , \2270_b0 , w_5133 );
and ( w_5132 ,  , w_5133 );
buf ( w_5131 , \2271_b1 );
not ( w_5131 , w_5134 );
not (  , w_5135 );
and ( w_5134 , w_5135 , \2271_b0 );
or ( \2273_b1 , \2272_b1 , w_5136 );
xor ( \2273_b0 , \2272_b0 , w_5138 );
not ( w_5138 , w_5139 );
and ( w_5139 , w_5136 , w_5137 );
buf ( w_5136 , \1610_b1 );
not ( w_5136 , w_5140 );
not ( w_5137 , w_5141 );
and ( w_5140 , w_5141 , \1610_b0 );
or ( \2274_b1 , \2268_b1 , \2273_b1 );
not ( \2273_b1 , w_5142 );
and ( \2274_b0 , \2268_b0 , w_5143 );
and ( w_5142 , w_5143 , \2273_b0 );
or ( \2275_b1 , \2264_b1 , \2273_b1 );
not ( \2273_b1 , w_5144 );
and ( \2275_b0 , \2264_b0 , w_5145 );
and ( w_5144 , w_5145 , \2273_b0 );
or ( \2277_b1 , \2256_b1 , \2276_b1 );
not ( \2276_b1 , w_5146 );
and ( \2277_b0 , \2256_b0 , w_5147 );
and ( w_5146 , w_5147 , \2276_b0 );
or ( \2278_b1 , \2240_b1 , \2276_b1 );
not ( \2276_b1 , w_5148 );
and ( \2278_b0 , \2240_b0 , w_5149 );
and ( w_5148 , w_5149 , \2276_b0 );
or ( \2280_b1 , \1299_b1 , \503_b1 );
not ( \503_b1 , w_5150 );
and ( \2280_b0 , \1299_b0 , w_5151 );
and ( w_5150 , w_5151 , \503_b0 );
or ( \2281_b1 , \1194_b1 , \501_b1 );
not ( \501_b1 , w_5152 );
and ( \2281_b0 , \1194_b0 , w_5153 );
and ( w_5152 , w_5153 , \501_b0 );
or ( \2282_b1 , \2280_b1 , w_5155 );
not ( w_5155 , w_5156 );
and ( \2282_b0 , \2280_b0 , w_5157 );
and ( w_5156 ,  , w_5157 );
buf ( w_5155 , \2281_b1 );
not ( w_5155 , w_5158 );
not (  , w_5159 );
and ( w_5158 , w_5159 , \2281_b0 );
or ( \2283_b1 , \2282_b1 , w_5160 );
xor ( \2283_b0 , \2282_b0 , w_5162 );
not ( w_5162 , w_5163 );
and ( w_5163 , w_5160 , w_5161 );
buf ( w_5160 , \455_b1 );
not ( w_5160 , w_5164 );
not ( w_5161 , w_5165 );
and ( w_5164 , w_5165 , \455_b0 );
or ( \2284_b1 , \1422_b1 , \298_b1 );
not ( \298_b1 , w_5166 );
and ( \2284_b0 , \1422_b0 , w_5167 );
and ( w_5166 , w_5167 , \298_b0 );
or ( \2285_b1 , \1304_b1 , \296_b1 );
not ( \296_b1 , w_5168 );
and ( \2285_b0 , \1304_b0 , w_5169 );
and ( w_5168 , w_5169 , \296_b0 );
or ( \2286_b1 , \2284_b1 , w_5171 );
not ( w_5171 , w_5172 );
and ( \2286_b0 , \2284_b0 , w_5173 );
and ( w_5172 ,  , w_5173 );
buf ( w_5171 , \2285_b1 );
not ( w_5171 , w_5174 );
not (  , w_5175 );
and ( w_5174 , w_5175 , \2285_b0 );
or ( \2287_b1 , \2286_b1 , w_5176 );
xor ( \2287_b0 , \2286_b0 , w_5178 );
not ( w_5178 , w_5179 );
and ( w_5179 , w_5176 , w_5177 );
buf ( w_5176 , \303_b1 );
not ( w_5176 , w_5180 );
not ( w_5177 , w_5181 );
and ( w_5180 , w_5181 , \303_b0 );
or ( \2288_b1 , \2283_b1 , \2287_b1 );
not ( \2287_b1 , w_5182 );
and ( \2288_b0 , \2283_b0 , w_5183 );
and ( w_5182 , w_5183 , \2287_b0 );
or ( \2289_b1 , \1770_b1 , \313_b1 );
not ( \313_b1 , w_5184 );
and ( \2289_b0 , \1770_b0 , w_5185 );
and ( w_5184 , w_5185 , \313_b0 );
or ( \2290_b1 , \1537_b1 , \311_b1 );
not ( \311_b1 , w_5186 );
and ( \2290_b0 , \1537_b0 , w_5187 );
and ( w_5186 , w_5187 , \311_b0 );
or ( \2291_b1 , \2289_b1 , w_5189 );
not ( w_5189 , w_5190 );
and ( \2291_b0 , \2289_b0 , w_5191 );
and ( w_5190 ,  , w_5191 );
buf ( w_5189 , \2290_b1 );
not ( w_5189 , w_5192 );
not (  , w_5193 );
and ( w_5192 , w_5193 , \2290_b0 );
or ( \2292_b1 , \2291_b1 , w_5194 );
xor ( \2292_b0 , \2291_b0 , w_5196 );
not ( w_5196 , w_5197 );
and ( w_5197 , w_5194 , w_5195 );
buf ( w_5194 , \320_b1 );
not ( w_5194 , w_5198 );
not ( w_5195 , w_5199 );
and ( w_5198 , w_5199 , \320_b0 );
or ( \2293_b1 , \2287_b1 , \2292_b1 );
not ( \2292_b1 , w_5200 );
and ( \2293_b0 , \2287_b0 , w_5201 );
and ( w_5200 , w_5201 , \2292_b0 );
or ( \2294_b1 , \2283_b1 , \2292_b1 );
not ( \2292_b1 , w_5202 );
and ( \2294_b0 , \2283_b0 , w_5203 );
and ( w_5202 , w_5203 , \2292_b0 );
or ( \2296_b1 , \2023_b1 , \331_b1 );
not ( \331_b1 , w_5204 );
and ( \2296_b0 , \2023_b0 , w_5205 );
and ( w_5204 , w_5205 , \331_b0 );
or ( \2297_b1 , \1778_b1 , \329_b1 );
not ( \329_b1 , w_5206 );
and ( \2297_b0 , \1778_b0 , w_5207 );
and ( w_5206 , w_5207 , \329_b0 );
or ( \2298_b1 , \2296_b1 , w_5209 );
not ( w_5209 , w_5210 );
and ( \2298_b0 , \2296_b0 , w_5211 );
and ( w_5210 ,  , w_5211 );
buf ( w_5209 , \2297_b1 );
not ( w_5209 , w_5212 );
not (  , w_5213 );
and ( w_5212 , w_5213 , \2297_b0 );
or ( \2299_b1 , \2298_b1 , w_5214 );
xor ( \2299_b0 , \2298_b0 , w_5216 );
not ( w_5216 , w_5217 );
and ( w_5217 , w_5214 , w_5215 );
buf ( w_5214 , \338_b1 );
not ( w_5214 , w_5218 );
not ( w_5215 , w_5219 );
and ( w_5218 , w_5219 , \338_b0 );
or ( \2300_b1 , \2161_b1 , \351_b1 );
not ( \351_b1 , w_5220 );
and ( \2300_b0 , \2161_b0 , w_5221 );
and ( w_5220 , w_5221 , \351_b0 );
or ( \2301_b1 , \2028_b1 , \349_b1 );
not ( \349_b1 , w_5222 );
and ( \2301_b0 , \2028_b0 , w_5223 );
and ( w_5222 , w_5223 , \349_b0 );
or ( \2302_b1 , \2300_b1 , w_5225 );
not ( w_5225 , w_5226 );
and ( \2302_b0 , \2300_b0 , w_5227 );
and ( w_5226 ,  , w_5227 );
buf ( w_5225 , \2301_b1 );
not ( w_5225 , w_5228 );
not (  , w_5229 );
and ( w_5228 , w_5229 , \2301_b0 );
or ( \2303_b1 , \2302_b1 , w_5230 );
xor ( \2303_b0 , \2302_b0 , w_5232 );
not ( w_5232 , w_5233 );
and ( w_5233 , w_5230 , w_5231 );
buf ( w_5230 , \358_b1 );
not ( w_5230 , w_5234 );
not ( w_5231 , w_5235 );
and ( w_5234 , w_5235 , \358_b0 );
or ( \2304_b1 , \2299_b1 , \2303_b1 );
not ( \2303_b1 , w_5236 );
and ( \2304_b0 , \2299_b0 , w_5237 );
and ( w_5236 , w_5237 , \2303_b0 );
buf ( \2305_b1 , RIb4bc180_92_b1 );
buf ( \2305_b0 , RIb4bc180_92_b0 );
or ( \2306_b1 , \2305_b1 , \345_b1 );
not ( \345_b1 , w_5238 );
and ( \2306_b0 , \2305_b0 , w_5239 );
and ( w_5238 , w_5239 , \345_b0 );
or ( \2307_b1 , \2303_b1 , \2306_b1 );
not ( \2306_b1 , w_5240 );
and ( \2307_b0 , \2303_b0 , w_5241 );
and ( w_5240 , w_5241 , \2306_b0 );
or ( \2308_b1 , \2299_b1 , \2306_b1 );
not ( \2306_b1 , w_5242 );
and ( \2308_b0 , \2299_b0 , w_5243 );
and ( w_5242 , w_5243 , \2306_b0 );
or ( \2310_b1 , \2295_b1 , \2309_b1 );
not ( \2309_b1 , w_5244 );
and ( \2310_b0 , \2295_b0 , w_5245 );
and ( w_5244 , w_5245 , \2309_b0 );
or ( \2311_b1 , \2155_b1 , \2159_b1 );
xor ( \2311_b0 , \2155_b0 , w_5246 );
not ( w_5246 , w_5247 );
and ( w_5247 , \2159_b1 , \2159_b0 );
or ( \2312_b1 , \2311_b1 , \2162_b1 );
xor ( \2312_b0 , \2311_b0 , w_5248 );
not ( w_5248 , w_5249 );
and ( w_5249 , \2162_b1 , \2162_b0 );
or ( \2313_b1 , \2309_b1 , \2312_b1 );
not ( \2312_b1 , w_5250 );
and ( \2313_b0 , \2309_b0 , w_5251 );
and ( w_5250 , w_5251 , \2312_b0 );
or ( \2314_b1 , \2295_b1 , \2312_b1 );
not ( \2312_b1 , w_5252 );
and ( \2314_b0 , \2295_b0 , w_5253 );
and ( w_5252 , w_5253 , \2312_b0 );
or ( \2316_b1 , \2279_b1 , \2315_b1 );
not ( \2315_b1 , w_5254 );
and ( \2316_b0 , \2279_b0 , w_5255 );
and ( w_5254 , w_5255 , \2315_b0 );
or ( \2317_b1 , \2088_b1 , \2092_b1 );
xor ( \2317_b0 , \2088_b0 , w_5256 );
not ( w_5256 , w_5257 );
and ( w_5257 , \2092_b1 , \2092_b0 );
or ( \2318_b1 , \2317_b1 , \2097_b1 );
xor ( \2318_b0 , \2317_b0 , w_5258 );
not ( w_5258 , w_5259 );
and ( w_5259 , \2097_b1 , \2097_b0 );
or ( \2319_b1 , \2104_b1 , \2108_b1 );
xor ( \2319_b0 , \2104_b0 , w_5260 );
not ( w_5260 , w_5261 );
and ( w_5261 , \2108_b1 , \2108_b0 );
or ( \2320_b1 , \2319_b1 , \2113_b1 );
xor ( \2320_b0 , \2319_b0 , w_5262 );
not ( w_5262 , w_5263 );
and ( w_5263 , \2113_b1 , \2113_b0 );
or ( \2321_b1 , \2318_b1 , \2320_b1 );
not ( \2320_b1 , w_5264 );
and ( \2321_b0 , \2318_b0 , w_5265 );
and ( w_5264 , w_5265 , \2320_b0 );
or ( \2322_b1 , \2169_b1 , \2173_b1 );
xor ( \2322_b0 , \2169_b0 , w_5266 );
not ( w_5266 , w_5267 );
and ( w_5267 , \2173_b1 , \2173_b0 );
or ( \2323_b1 , \2322_b1 , \2178_b1 );
xor ( \2323_b0 , \2322_b0 , w_5268 );
not ( w_5268 , w_5269 );
and ( w_5269 , \2178_b1 , \2178_b0 );
or ( \2324_b1 , \2320_b1 , \2323_b1 );
not ( \2323_b1 , w_5270 );
and ( \2324_b0 , \2320_b0 , w_5271 );
and ( w_5270 , w_5271 , \2323_b0 );
or ( \2325_b1 , \2318_b1 , \2323_b1 );
not ( \2323_b1 , w_5272 );
and ( \2325_b0 , \2318_b0 , w_5273 );
and ( w_5272 , w_5273 , \2323_b0 );
or ( \2327_b1 , \2315_b1 , \2326_b1 );
not ( \2326_b1 , w_5274 );
and ( \2327_b0 , \2315_b0 , w_5275 );
and ( w_5274 , w_5275 , \2326_b0 );
or ( \2328_b1 , \2279_b1 , \2326_b1 );
not ( \2326_b1 , w_5276 );
and ( \2328_b0 , \2279_b0 , w_5277 );
and ( w_5276 , w_5277 , \2326_b0 );
or ( \2330_b1 , \1958_b1 , \1962_b1 );
xor ( \2330_b0 , \1958_b0 , w_5278 );
not ( w_5278 , w_5279 );
and ( w_5279 , \1962_b1 , \1962_b0 );
or ( \2331_b1 , \2330_b1 , \1967_b1 );
xor ( \2331_b0 , \2330_b0 , w_5280 );
not ( w_5280 , w_5281 );
and ( w_5281 , \1967_b1 , \1967_b0 );
or ( \2332_b1 , \2142_b1 , \2144_b1 );
xor ( \2332_b0 , \2142_b0 , w_5282 );
not ( w_5282 , w_5283 );
and ( w_5283 , \2144_b1 , \2144_b0 );
or ( \2333_b1 , \2332_b1 , \2147_b1 );
xor ( \2333_b0 , \2332_b0 , w_5284 );
not ( w_5284 , w_5285 );
and ( w_5285 , \2147_b1 , \2147_b0 );
or ( \2334_b1 , \2331_b1 , \2333_b1 );
not ( \2333_b1 , w_5286 );
and ( \2334_b0 , \2331_b0 , w_5287 );
and ( w_5286 , w_5287 , \2333_b0 );
or ( \2335_b1 , \2165_b1 , \2181_b1 );
xor ( \2335_b0 , \2165_b0 , w_5288 );
not ( w_5288 , w_5289 );
and ( w_5289 , \2181_b1 , \2181_b0 );
or ( \2336_b1 , \2335_b1 , \2183_b1 );
xor ( \2336_b0 , \2335_b0 , w_5290 );
not ( w_5290 , w_5291 );
and ( w_5291 , \2183_b1 , \2183_b0 );
or ( \2337_b1 , \2333_b1 , \2336_b1 );
not ( \2336_b1 , w_5292 );
and ( \2337_b0 , \2333_b0 , w_5293 );
and ( w_5292 , w_5293 , \2336_b0 );
or ( \2338_b1 , \2331_b1 , \2336_b1 );
not ( \2336_b1 , w_5294 );
and ( \2338_b0 , \2331_b0 , w_5295 );
and ( w_5294 , w_5295 , \2336_b0 );
or ( \2340_b1 , \2329_b1 , \2339_b1 );
not ( \2339_b1 , w_5296 );
and ( \2340_b0 , \2329_b0 , w_5297 );
and ( w_5296 , w_5297 , \2339_b0 );
or ( \2341_b1 , \2022_b1 , \2030_b1 );
xor ( \2341_b0 , \2022_b0 , w_5298 );
not ( w_5298 , w_5299 );
and ( w_5299 , \2030_b1 , \2030_b0 );
or ( \2342_b1 , \2341_b1 , \2035_b1 );
xor ( \2342_b0 , \2341_b0 , w_5300 );
not ( w_5300 , w_5301 );
and ( w_5301 , \2035_b1 , \2035_b0 );
or ( \2343_b1 , \2339_b1 , \2342_b1 );
not ( \2342_b1 , w_5302 );
and ( \2343_b0 , \2339_b0 , w_5303 );
and ( w_5302 , w_5303 , \2342_b0 );
or ( \2344_b1 , \2329_b1 , \2342_b1 );
not ( \2342_b1 , w_5304 );
and ( \2344_b0 , \2329_b0 , w_5305 );
and ( w_5304 , w_5305 , \2342_b0 );
or ( \2346_b1 , \1970_b1 , \1986_b1 );
xor ( \2346_b0 , \1970_b0 , w_5306 );
not ( w_5306 , w_5307 );
and ( w_5307 , \1986_b1 , \1986_b0 );
or ( \2347_b1 , \2346_b1 , \2003_b1 );
xor ( \2347_b0 , \2346_b0 , w_5308 );
not ( w_5308 , w_5309 );
and ( w_5309 , \2003_b1 , \2003_b0 );
or ( \2348_b1 , \2140_b1 , \2150_b1 );
xor ( \2348_b0 , \2140_b0 , w_5310 );
not ( w_5310 , w_5311 );
and ( w_5311 , \2150_b1 , \2150_b0 );
or ( \2349_b1 , \2348_b1 , \2186_b1 );
xor ( \2349_b0 , \2348_b0 , w_5312 );
not ( w_5312 , w_5313 );
and ( w_5313 , \2186_b1 , \2186_b0 );
or ( \2350_b1 , \2347_b1 , \2349_b1 );
not ( \2349_b1 , w_5314 );
and ( \2350_b0 , \2347_b0 , w_5315 );
and ( w_5314 , w_5315 , \2349_b0 );
or ( \2351_b1 , \2191_b1 , \2193_b1 );
xor ( \2351_b0 , \2191_b0 , w_5316 );
not ( w_5316 , w_5317 );
and ( w_5317 , \2193_b1 , \2193_b0 );
or ( \2352_b1 , \2351_b1 , \2196_b1 );
xor ( \2352_b0 , \2351_b0 , w_5318 );
not ( w_5318 , w_5319 );
and ( w_5319 , \2196_b1 , \2196_b0 );
or ( \2353_b1 , \2349_b1 , \2352_b1 );
not ( \2352_b1 , w_5320 );
and ( \2353_b0 , \2349_b0 , w_5321 );
and ( w_5320 , w_5321 , \2352_b0 );
or ( \2354_b1 , \2347_b1 , \2352_b1 );
not ( \2352_b1 , w_5322 );
and ( \2354_b0 , \2347_b0 , w_5323 );
and ( w_5322 , w_5323 , \2352_b0 );
or ( \2356_b1 , \2345_b1 , \2355_b1 );
not ( \2355_b1 , w_5324 );
and ( \2356_b0 , \2345_b0 , w_5325 );
and ( w_5324 , w_5325 , \2355_b0 );
or ( \2357_b1 , \2006_b1 , \2038_b1 );
xor ( \2357_b0 , \2006_b0 , w_5326 );
not ( w_5326 , w_5327 );
and ( w_5327 , \2038_b1 , \2038_b0 );
or ( \2358_b1 , \2357_b1 , \2048_b1 );
xor ( \2358_b0 , \2357_b0 , w_5328 );
not ( w_5328 , w_5329 );
and ( w_5329 , \2048_b1 , \2048_b0 );
or ( \2359_b1 , \2355_b1 , \2358_b1 );
not ( \2358_b1 , w_5330 );
and ( \2359_b0 , \2355_b0 , w_5331 );
and ( w_5330 , w_5331 , \2358_b0 );
or ( \2360_b1 , \2345_b1 , \2358_b1 );
not ( \2358_b1 , w_5332 );
and ( \2360_b0 , \2345_b0 , w_5333 );
and ( w_5332 , w_5333 , \2358_b0 );
or ( \2362_b1 , \2205_b1 , \2207_b1 );
xor ( \2362_b0 , \2205_b0 , w_5334 );
not ( w_5334 , w_5335 );
and ( w_5335 , \2207_b1 , \2207_b0 );
or ( \2363_b1 , \2362_b1 , \2209_b1 );
xor ( \2363_b0 , \2362_b0 , w_5336 );
not ( w_5336 , w_5337 );
and ( w_5337 , \2209_b1 , \2209_b0 );
or ( \2364_b1 , \2361_b1 , \2363_b1 );
not ( \2363_b1 , w_5338 );
and ( \2364_b0 , \2361_b0 , w_5339 );
and ( w_5338 , w_5339 , \2363_b0 );
or ( \2365_b1 , \2224_b1 , \2364_b1 );
not ( \2364_b1 , w_5340 );
and ( \2365_b0 , \2224_b0 , w_5341 );
and ( w_5340 , w_5341 , \2364_b0 );
or ( \2366_b1 , \2224_b1 , \2364_b1 );
xor ( \2366_b0 , \2224_b0 , w_5342 );
not ( w_5342 , w_5343 );
and ( w_5343 , \2364_b1 , \2364_b0 );
or ( \2367_b1 , \2361_b1 , \2363_b1 );
xor ( \2367_b0 , \2361_b0 , w_5344 );
not ( w_5344 , w_5345 );
and ( w_5345 , \2363_b1 , \2363_b0 );
and ( \2368_nR126_b1 , RIb4c2b70_62_b1 , w_5346 );
xor ( w_5346 , RIb4c2b70_62_b0 , \288_b1 );
not ( \288_b1 , w_5347 );
and ( \2368_nR126_b0 , w_5347 , \288_b0 );
buf ( \2369_b1 , \2368_nR126_b1 );
buf ( \2369_b0 , \2368_nR126_b0 );
and ( \2370_nR125_b1 , RIb4c2af8_63_b1 , w_5348 );
xor ( w_5348 , RIb4c2af8_63_b0 , \288_b1 );
not ( \288_b1 , w_5349 );
and ( \2370_nR125_b0 , w_5349 , \288_b0 );
buf ( \2371_b1 , \2370_nR125_b1 );
buf ( \2371_b0 , \2370_nR125_b0 );
or ( \2372_b1 , \2369_b1 , \2371_b1 );
not ( \2371_b1 , w_5350 );
and ( \2372_b0 , \2369_b0 , w_5351 );
and ( w_5350 , w_5351 , \2371_b0 );
buf ( \2373_b1 , \2372_b1 );
not ( \2373_b1 , w_5352 );
not ( \2373_b0 , w_5353 );
and ( w_5352 , w_5353 , \2372_b0 );
or ( \2374_b1 , \2121_b1 , \2373_b1 );
not ( \2373_b1 , w_5354 );
and ( \2374_b0 , \2121_b0 , w_5355 );
and ( w_5354 , w_5355 , \2373_b0 );
buf ( \2375_b1 , \2374_b1 );
not ( \2375_b1 , w_5356 );
not ( \2375_b0 , w_5357 );
and ( w_5356 , w_5357 , \2374_b0 );
or ( \2376_b1 , \315_b1 , \2261_b1 );
not ( \2261_b1 , w_5358 );
and ( \2376_b0 , \315_b0 , w_5359 );
and ( w_5358 , w_5359 , \2261_b0 );
or ( \2377_b1 , \159_b1 , \2259_b1 );
not ( \2259_b1 , w_5360 );
and ( \2377_b0 , \159_b0 , w_5361 );
and ( w_5360 , w_5361 , \2259_b0 );
or ( \2378_b1 , \2376_b1 , w_5363 );
not ( w_5363 , w_5364 );
and ( \2378_b0 , \2376_b0 , w_5365 );
and ( w_5364 ,  , w_5365 );
buf ( w_5363 , \2377_b1 );
not ( w_5363 , w_5366 );
not (  , w_5367 );
and ( w_5366 , w_5367 , \2377_b0 );
or ( \2379_b1 , \2378_b1 , w_5368 );
xor ( \2379_b0 , \2378_b0 , w_5370 );
not ( w_5370 , w_5371 );
and ( w_5371 , w_5368 , w_5369 );
buf ( w_5368 , \2124_b1 );
not ( w_5368 , w_5372 );
not ( w_5369 , w_5373 );
and ( w_5372 , w_5373 , \2124_b0 );
or ( \2380_b1 , \2375_b1 , \2379_b1 );
not ( \2379_b1 , w_5374 );
and ( \2380_b0 , \2375_b0 , w_5375 );
and ( w_5374 , w_5375 , \2379_b0 );
or ( \2381_b1 , \333_b1 , \1955_b1 );
not ( \1955_b1 , w_5376 );
and ( \2381_b0 , \333_b0 , w_5377 );
and ( w_5376 , w_5377 , \1955_b0 );
or ( \2382_b1 , \305_b1 , \1953_b1 );
not ( \1953_b1 , w_5378 );
and ( \2382_b0 , \305_b0 , w_5379 );
and ( w_5378 , w_5379 , \1953_b0 );
or ( \2383_b1 , \2381_b1 , w_5381 );
not ( w_5381 , w_5382 );
and ( \2383_b0 , \2381_b0 , w_5383 );
and ( w_5382 ,  , w_5383 );
buf ( w_5381 , \2382_b1 );
not ( w_5381 , w_5384 );
not (  , w_5385 );
and ( w_5384 , w_5385 , \2382_b0 );
or ( \2384_b1 , \2383_b1 , w_5386 );
xor ( \2384_b0 , \2383_b0 , w_5388 );
not ( w_5388 , w_5389 );
and ( w_5389 , w_5386 , w_5387 );
buf ( w_5386 , \1835_b1 );
not ( w_5386 , w_5390 );
not ( w_5387 , w_5391 );
and ( w_5390 , w_5391 , \1835_b0 );
or ( \2385_b1 , \2379_b1 , \2384_b1 );
not ( \2384_b1 , w_5392 );
and ( \2385_b0 , \2379_b0 , w_5393 );
and ( w_5392 , w_5393 , \2384_b0 );
or ( \2386_b1 , \2375_b1 , \2384_b1 );
not ( \2384_b1 , w_5394 );
and ( \2386_b0 , \2375_b0 , w_5395 );
and ( w_5394 , w_5395 , \2384_b0 );
or ( \2388_b1 , \353_b1 , \1742_b1 );
not ( \1742_b1 , w_5396 );
and ( \2388_b0 , \353_b0 , w_5397 );
and ( w_5396 , w_5397 , \1742_b0 );
or ( \2389_b1 , \323_b1 , \1740_b1 );
not ( \1740_b1 , w_5398 );
and ( \2389_b0 , \323_b0 , w_5399 );
and ( w_5398 , w_5399 , \1740_b0 );
or ( \2390_b1 , \2388_b1 , w_5401 );
not ( w_5401 , w_5402 );
and ( \2390_b0 , \2388_b0 , w_5403 );
and ( w_5402 ,  , w_5403 );
buf ( w_5401 , \2389_b1 );
not ( w_5401 , w_5404 );
not (  , w_5405 );
and ( w_5404 , w_5405 , \2389_b0 );
or ( \2391_b1 , \2390_b1 , w_5406 );
xor ( \2391_b0 , \2390_b0 , w_5408 );
not ( w_5408 , w_5409 );
and ( w_5409 , w_5406 , w_5407 );
buf ( w_5406 , \1610_b1 );
not ( w_5406 , w_5410 );
not ( w_5407 , w_5411 );
and ( w_5410 , w_5411 , \1610_b0 );
or ( \2392_b1 , \360_b1 , \1476_b1 );
not ( \1476_b1 , w_5412 );
and ( \2392_b0 , \360_b0 , w_5413 );
and ( w_5412 , w_5413 , \1476_b0 );
or ( \2393_b1 , \343_b1 , \1474_b1 );
not ( \1474_b1 , w_5414 );
and ( \2393_b0 , \343_b0 , w_5415 );
and ( w_5414 , w_5415 , \1474_b0 );
or ( \2394_b1 , \2392_b1 , w_5417 );
not ( w_5417 , w_5418 );
and ( \2394_b0 , \2392_b0 , w_5419 );
and ( w_5418 ,  , w_5419 );
buf ( w_5417 , \2393_b1 );
not ( w_5417 , w_5420 );
not (  , w_5421 );
and ( w_5420 , w_5421 , \2393_b0 );
or ( \2395_b1 , \2394_b1 , w_5422 );
xor ( \2395_b0 , \2394_b0 , w_5424 );
not ( w_5424 , w_5425 );
and ( w_5425 , w_5422 , w_5423 );
buf ( w_5422 , \1363_b1 );
not ( w_5422 , w_5426 );
not ( w_5423 , w_5427 );
and ( w_5426 , w_5427 , \1363_b0 );
or ( \2396_b1 , \2391_b1 , \2395_b1 );
not ( \2395_b1 , w_5428 );
and ( \2396_b0 , \2391_b0 , w_5429 );
and ( w_5428 , w_5429 , \2395_b0 );
or ( \2397_b1 , \495_b1 , \1280_b1 );
not ( \1280_b1 , w_5430 );
and ( \2397_b0 , \495_b0 , w_5431 );
and ( w_5430 , w_5431 , \1280_b0 );
or ( \2398_b1 , \444_b1 , \1278_b1 );
not ( \1278_b1 , w_5432 );
and ( \2398_b0 , \444_b0 , w_5433 );
and ( w_5432 , w_5433 , \1278_b0 );
or ( \2399_b1 , \2397_b1 , w_5435 );
not ( w_5435 , w_5436 );
and ( \2399_b0 , \2397_b0 , w_5437 );
and ( w_5436 ,  , w_5437 );
buf ( w_5435 , \2398_b1 );
not ( w_5435 , w_5438 );
not (  , w_5439 );
and ( w_5438 , w_5439 , \2398_b0 );
or ( \2400_b1 , \2399_b1 , w_5440 );
xor ( \2400_b0 , \2399_b0 , w_5442 );
not ( w_5442 , w_5443 );
and ( w_5443 , w_5440 , w_5441 );
buf ( w_5440 , \1177_b1 );
not ( w_5440 , w_5444 );
not ( w_5441 , w_5445 );
and ( w_5444 , w_5445 , \1177_b0 );
or ( \2401_b1 , \2395_b1 , \2400_b1 );
not ( \2400_b1 , w_5446 );
and ( \2401_b0 , \2395_b0 , w_5447 );
and ( w_5446 , w_5447 , \2400_b0 );
or ( \2402_b1 , \2391_b1 , \2400_b1 );
not ( \2400_b1 , w_5448 );
and ( \2402_b0 , \2391_b0 , w_5449 );
and ( w_5448 , w_5449 , \2400_b0 );
or ( \2404_b1 , \2387_b1 , \2403_b1 );
not ( \2403_b1 , w_5450 );
and ( \2404_b0 , \2387_b0 , w_5451 );
and ( w_5450 , w_5451 , \2403_b0 );
or ( \2405_b1 , \621_b1 , \1062_b1 );
not ( \1062_b1 , w_5452 );
and ( \2405_b0 , \621_b0 , w_5453 );
and ( w_5452 , w_5453 , \1062_b0 );
or ( \2406_b1 , \593_b1 , \1060_b1 );
not ( \1060_b1 , w_5454 );
and ( \2406_b0 , \593_b0 , w_5455 );
and ( w_5454 , w_5455 , \1060_b0 );
or ( \2407_b1 , \2405_b1 , w_5457 );
not ( w_5457 , w_5458 );
and ( \2407_b0 , \2405_b0 , w_5459 );
and ( w_5458 ,  , w_5459 );
buf ( w_5457 , \2406_b1 );
not ( w_5457 , w_5460 );
not (  , w_5461 );
and ( w_5460 , w_5461 , \2406_b0 );
or ( \2408_b1 , \2407_b1 , w_5462 );
xor ( \2408_b0 , \2407_b0 , w_5464 );
not ( w_5464 , w_5465 );
and ( w_5465 , w_5462 , w_5463 );
buf ( w_5462 , \984_b1 );
not ( w_5462 , w_5466 );
not ( w_5463 , w_5467 );
and ( w_5466 , w_5467 , \984_b0 );
or ( \2409_b1 , \777_b1 , \912_b1 );
not ( \912_b1 , w_5468 );
and ( \2409_b0 , \777_b0 , w_5469 );
and ( w_5468 , w_5469 , \912_b0 );
or ( \2410_b1 , \703_b1 , \910_b1 );
not ( \910_b1 , w_5470 );
and ( \2410_b0 , \703_b0 , w_5471 );
and ( w_5470 , w_5471 , \910_b0 );
or ( \2411_b1 , \2409_b1 , w_5473 );
not ( w_5473 , w_5474 );
and ( \2411_b0 , \2409_b0 , w_5475 );
and ( w_5474 ,  , w_5475 );
buf ( w_5473 , \2410_b1 );
not ( w_5473 , w_5476 );
not (  , w_5477 );
and ( w_5476 , w_5477 , \2410_b0 );
or ( \2412_b1 , \2411_b1 , w_5478 );
xor ( \2412_b0 , \2411_b0 , w_5480 );
not ( w_5480 , w_5481 );
and ( w_5481 , w_5478 , w_5479 );
buf ( w_5478 , \818_b1 );
not ( w_5478 , w_5482 );
not ( w_5479 , w_5483 );
and ( w_5482 , w_5483 , \818_b0 );
or ( \2413_b1 , \2408_b1 , \2412_b1 );
not ( \2412_b1 , w_5484 );
and ( \2413_b0 , \2408_b0 , w_5485 );
and ( w_5484 , w_5485 , \2412_b0 );
or ( \2414_b1 , \904_b1 , \740_b1 );
not ( \740_b1 , w_5486 );
and ( \2414_b0 , \904_b0 , w_5487 );
and ( w_5486 , w_5487 , \740_b0 );
or ( \2415_b1 , \841_b1 , \738_b1 );
not ( \738_b1 , w_5488 );
and ( \2415_b0 , \841_b0 , w_5489 );
and ( w_5488 , w_5489 , \738_b0 );
or ( \2416_b1 , \2414_b1 , w_5491 );
not ( w_5491 , w_5492 );
and ( \2416_b0 , \2414_b0 , w_5493 );
and ( w_5492 ,  , w_5493 );
buf ( w_5491 , \2415_b1 );
not ( w_5491 , w_5494 );
not (  , w_5495 );
and ( w_5494 , w_5495 , \2415_b0 );
or ( \2417_b1 , \2416_b1 , w_5496 );
xor ( \2417_b0 , \2416_b0 , w_5498 );
not ( w_5498 , w_5499 );
and ( w_5499 , w_5496 , w_5497 );
buf ( w_5496 , \668_b1 );
not ( w_5496 , w_5500 );
not ( w_5497 , w_5501 );
and ( w_5500 , w_5501 , \668_b0 );
or ( \2418_b1 , \2412_b1 , \2417_b1 );
not ( \2417_b1 , w_5502 );
and ( \2418_b0 , \2412_b0 , w_5503 );
and ( w_5502 , w_5503 , \2417_b0 );
or ( \2419_b1 , \2408_b1 , \2417_b1 );
not ( \2417_b1 , w_5504 );
and ( \2419_b0 , \2408_b0 , w_5505 );
and ( w_5504 , w_5505 , \2417_b0 );
or ( \2421_b1 , \2403_b1 , \2420_b1 );
not ( \2420_b1 , w_5506 );
and ( \2421_b0 , \2403_b0 , w_5507 );
and ( w_5506 , w_5507 , \2420_b0 );
or ( \2422_b1 , \2387_b1 , \2420_b1 );
not ( \2420_b1 , w_5508 );
and ( \2422_b0 , \2387_b0 , w_5509 );
and ( w_5508 , w_5509 , \2420_b0 );
or ( \2424_b1 , \2228_b1 , \2232_b1 );
xor ( \2424_b0 , \2228_b0 , w_5510 );
not ( w_5510 , w_5511 );
and ( w_5511 , \2232_b1 , \2232_b0 );
or ( \2425_b1 , \2424_b1 , \2237_b1 );
xor ( \2425_b0 , \2424_b0 , w_5512 );
not ( w_5512 , w_5513 );
and ( w_5513 , \2237_b1 , \2237_b0 );
or ( \2426_b1 , \2283_b1 , \2287_b1 );
xor ( \2426_b0 , \2283_b0 , w_5514 );
not ( w_5514 , w_5515 );
and ( w_5515 , \2287_b1 , \2287_b0 );
or ( \2427_b1 , \2426_b1 , \2292_b1 );
xor ( \2427_b0 , \2426_b0 , w_5516 );
not ( w_5516 , w_5517 );
and ( w_5517 , \2292_b1 , \2292_b0 );
or ( \2428_b1 , \2425_b1 , \2427_b1 );
not ( \2427_b1 , w_5518 );
and ( \2428_b0 , \2425_b0 , w_5519 );
and ( w_5518 , w_5519 , \2427_b0 );
or ( \2429_b1 , \2299_b1 , \2303_b1 );
xor ( \2429_b0 , \2299_b0 , w_5520 );
not ( w_5520 , w_5521 );
and ( w_5521 , \2303_b1 , \2303_b0 );
or ( \2430_b1 , \2429_b1 , \2306_b1 );
xor ( \2430_b0 , \2429_b0 , w_5522 );
not ( w_5522 , w_5523 );
and ( w_5523 , \2306_b1 , \2306_b0 );
or ( \2431_b1 , \2427_b1 , \2430_b1 );
not ( \2430_b1 , w_5524 );
and ( \2431_b0 , \2427_b0 , w_5525 );
and ( w_5524 , w_5525 , \2430_b0 );
or ( \2432_b1 , \2425_b1 , \2430_b1 );
not ( \2430_b1 , w_5526 );
and ( \2432_b0 , \2425_b0 , w_5527 );
and ( w_5526 , w_5527 , \2430_b0 );
or ( \2434_b1 , \2423_b1 , \2433_b1 );
not ( \2433_b1 , w_5528 );
and ( \2434_b0 , \2423_b0 , w_5529 );
and ( w_5528 , w_5529 , \2433_b0 );
or ( \2435_b1 , \1778_b1 , \313_b1 );
not ( \313_b1 , w_5530 );
and ( \2435_b0 , \1778_b0 , w_5531 );
and ( w_5530 , w_5531 , \313_b0 );
or ( \2436_b1 , \1770_b1 , \311_b1 );
not ( \311_b1 , w_5532 );
and ( \2436_b0 , \1770_b0 , w_5533 );
and ( w_5532 , w_5533 , \311_b0 );
or ( \2437_b1 , \2435_b1 , w_5535 );
not ( w_5535 , w_5536 );
and ( \2437_b0 , \2435_b0 , w_5537 );
and ( w_5536 ,  , w_5537 );
buf ( w_5535 , \2436_b1 );
not ( w_5535 , w_5538 );
not (  , w_5539 );
and ( w_5538 , w_5539 , \2436_b0 );
or ( \2438_b1 , \2437_b1 , w_5540 );
xor ( \2438_b0 , \2437_b0 , w_5542 );
not ( w_5542 , w_5543 );
and ( w_5543 , w_5540 , w_5541 );
buf ( w_5540 , \320_b1 );
not ( w_5540 , w_5544 );
not ( w_5541 , w_5545 );
and ( w_5544 , w_5545 , \320_b0 );
or ( \2439_b1 , \2028_b1 , \331_b1 );
not ( \331_b1 , w_5546 );
and ( \2439_b0 , \2028_b0 , w_5547 );
and ( w_5546 , w_5547 , \331_b0 );
or ( \2440_b1 , \2023_b1 , \329_b1 );
not ( \329_b1 , w_5548 );
and ( \2440_b0 , \2023_b0 , w_5549 );
and ( w_5548 , w_5549 , \329_b0 );
or ( \2441_b1 , \2439_b1 , w_5551 );
not ( w_5551 , w_5552 );
and ( \2441_b0 , \2439_b0 , w_5553 );
and ( w_5552 ,  , w_5553 );
buf ( w_5551 , \2440_b1 );
not ( w_5551 , w_5554 );
not (  , w_5555 );
and ( w_5554 , w_5555 , \2440_b0 );
or ( \2442_b1 , \2441_b1 , w_5556 );
xor ( \2442_b0 , \2441_b0 , w_5558 );
not ( w_5558 , w_5559 );
and ( w_5559 , w_5556 , w_5557 );
buf ( w_5556 , \338_b1 );
not ( w_5556 , w_5560 );
not ( w_5557 , w_5561 );
and ( w_5560 , w_5561 , \338_b0 );
or ( \2443_b1 , \2438_b1 , \2442_b1 );
not ( \2442_b1 , w_5562 );
and ( \2443_b0 , \2438_b0 , w_5563 );
and ( w_5562 , w_5563 , \2442_b0 );
or ( \2444_b1 , \2305_b1 , \351_b1 );
not ( \351_b1 , w_5564 );
and ( \2444_b0 , \2305_b0 , w_5565 );
and ( w_5564 , w_5565 , \351_b0 );
or ( \2445_b1 , \2161_b1 , \349_b1 );
not ( \349_b1 , w_5566 );
and ( \2445_b0 , \2161_b0 , w_5567 );
and ( w_5566 , w_5567 , \349_b0 );
or ( \2446_b1 , \2444_b1 , w_5569 );
not ( w_5569 , w_5570 );
and ( \2446_b0 , \2444_b0 , w_5571 );
and ( w_5570 ,  , w_5571 );
buf ( w_5569 , \2445_b1 );
not ( w_5569 , w_5572 );
not (  , w_5573 );
and ( w_5572 , w_5573 , \2445_b0 );
or ( \2447_b1 , \2446_b1 , w_5574 );
xor ( \2447_b0 , \2446_b0 , w_5576 );
not ( w_5576 , w_5577 );
and ( w_5577 , w_5574 , w_5575 );
buf ( w_5574 , \358_b1 );
not ( w_5574 , w_5578 );
not ( w_5575 , w_5579 );
and ( w_5578 , w_5579 , \358_b0 );
or ( \2448_b1 , \2442_b1 , \2447_b1 );
not ( \2447_b1 , w_5580 );
and ( \2448_b0 , \2442_b0 , w_5581 );
and ( w_5580 , w_5581 , \2447_b0 );
or ( \2449_b1 , \2438_b1 , \2447_b1 );
not ( \2447_b1 , w_5582 );
and ( \2449_b0 , \2438_b0 , w_5583 );
and ( w_5582 , w_5583 , \2447_b0 );
or ( \2451_b1 , \1194_b1 , \604_b1 );
not ( \604_b1 , w_5584 );
and ( \2451_b0 , \1194_b0 , w_5585 );
and ( w_5584 , w_5585 , \604_b0 );
or ( \2452_b1 , \1104_b1 , \602_b1 );
not ( \602_b1 , w_5586 );
and ( \2452_b0 , \1104_b0 , w_5587 );
and ( w_5586 , w_5587 , \602_b0 );
or ( \2453_b1 , \2451_b1 , w_5589 );
not ( w_5589 , w_5590 );
and ( \2453_b0 , \2451_b0 , w_5591 );
and ( w_5590 ,  , w_5591 );
buf ( w_5589 , \2452_b1 );
not ( w_5589 , w_5592 );
not (  , w_5593 );
and ( w_5592 , w_5593 , \2452_b0 );
or ( \2454_b1 , \2453_b1 , w_5594 );
xor ( \2454_b0 , \2453_b0 , w_5596 );
not ( w_5596 , w_5597 );
and ( w_5597 , w_5594 , w_5595 );
buf ( w_5594 , \561_b1 );
not ( w_5594 , w_5598 );
not ( w_5595 , w_5599 );
and ( w_5598 , w_5599 , \561_b0 );
or ( \2455_b1 , \1304_b1 , \503_b1 );
not ( \503_b1 , w_5600 );
and ( \2455_b0 , \1304_b0 , w_5601 );
and ( w_5600 , w_5601 , \503_b0 );
or ( \2456_b1 , \1299_b1 , \501_b1 );
not ( \501_b1 , w_5602 );
and ( \2456_b0 , \1299_b0 , w_5603 );
and ( w_5602 , w_5603 , \501_b0 );
or ( \2457_b1 , \2455_b1 , w_5605 );
not ( w_5605 , w_5606 );
and ( \2457_b0 , \2455_b0 , w_5607 );
and ( w_5606 ,  , w_5607 );
buf ( w_5605 , \2456_b1 );
not ( w_5605 , w_5608 );
not (  , w_5609 );
and ( w_5608 , w_5609 , \2456_b0 );
or ( \2458_b1 , \2457_b1 , w_5610 );
xor ( \2458_b0 , \2457_b0 , w_5612 );
not ( w_5612 , w_5613 );
and ( w_5613 , w_5610 , w_5611 );
buf ( w_5610 , \455_b1 );
not ( w_5610 , w_5614 );
not ( w_5611 , w_5615 );
and ( w_5614 , w_5615 , \455_b0 );
or ( \2459_b1 , \2454_b1 , \2458_b1 );
not ( \2458_b1 , w_5616 );
and ( \2459_b0 , \2454_b0 , w_5617 );
and ( w_5616 , w_5617 , \2458_b0 );
or ( \2460_b1 , \1537_b1 , \298_b1 );
not ( \298_b1 , w_5618 );
and ( \2460_b0 , \1537_b0 , w_5619 );
and ( w_5618 , w_5619 , \298_b0 );
or ( \2461_b1 , \1422_b1 , \296_b1 );
not ( \296_b1 , w_5620 );
and ( \2461_b0 , \1422_b0 , w_5621 );
and ( w_5620 , w_5621 , \296_b0 );
or ( \2462_b1 , \2460_b1 , w_5623 );
not ( w_5623 , w_5624 );
and ( \2462_b0 , \2460_b0 , w_5625 );
and ( w_5624 ,  , w_5625 );
buf ( w_5623 , \2461_b1 );
not ( w_5623 , w_5626 );
not (  , w_5627 );
and ( w_5626 , w_5627 , \2461_b0 );
or ( \2463_b1 , \2462_b1 , w_5628 );
xor ( \2463_b0 , \2462_b0 , w_5630 );
not ( w_5630 , w_5631 );
and ( w_5631 , w_5628 , w_5629 );
buf ( w_5628 , \303_b1 );
not ( w_5628 , w_5632 );
not ( w_5629 , w_5633 );
and ( w_5632 , w_5633 , \303_b0 );
or ( \2464_b1 , \2458_b1 , \2463_b1 );
not ( \2463_b1 , w_5634 );
and ( \2464_b0 , \2458_b0 , w_5635 );
and ( w_5634 , w_5635 , \2463_b0 );
or ( \2465_b1 , \2454_b1 , \2463_b1 );
not ( \2463_b1 , w_5636 );
and ( \2465_b0 , \2454_b0 , w_5637 );
and ( w_5636 , w_5637 , \2463_b0 );
or ( \2467_b1 , \2450_b1 , w_5638 );
or ( \2467_b0 , \2450_b0 , \2466_b0 );
not ( \2466_b0 , w_5639 );
and ( w_5639 , w_5638 , \2466_b1 );
or ( \2468_b1 , \2433_b1 , \2467_b1 );
not ( \2467_b1 , w_5640 );
and ( \2468_b0 , \2433_b0 , w_5641 );
and ( w_5640 , w_5641 , \2467_b0 );
or ( \2469_b1 , \2423_b1 , \2467_b1 );
not ( \2467_b1 , w_5642 );
and ( \2469_b0 , \2423_b0 , w_5643 );
and ( w_5642 , w_5643 , \2467_b0 );
or ( \2471_b1 , \2125_b1 , \2129_b1 );
xor ( \2471_b0 , \2125_b0 , w_5644 );
not ( w_5644 , w_5645 );
and ( w_5645 , \2129_b1 , \2129_b0 );
or ( \2472_b1 , \2471_b1 , \2134_b1 );
xor ( \2472_b0 , \2471_b0 , w_5646 );
not ( w_5646 , w_5647 );
and ( w_5647 , \2134_b1 , \2134_b0 );
or ( \2473_b1 , \2295_b1 , \2309_b1 );
xor ( \2473_b0 , \2295_b0 , w_5648 );
not ( w_5648 , w_5649 );
and ( w_5649 , \2309_b1 , \2309_b0 );
or ( \2474_b1 , \2473_b1 , \2312_b1 );
xor ( \2474_b0 , \2473_b0 , w_5650 );
not ( w_5650 , w_5651 );
and ( w_5651 , \2312_b1 , \2312_b0 );
or ( \2475_b1 , \2472_b1 , \2474_b1 );
not ( \2474_b1 , w_5652 );
and ( \2475_b0 , \2472_b0 , w_5653 );
and ( w_5652 , w_5653 , \2474_b0 );
or ( \2476_b1 , \2318_b1 , \2320_b1 );
xor ( \2476_b0 , \2318_b0 , w_5654 );
not ( w_5654 , w_5655 );
and ( w_5655 , \2320_b1 , \2320_b0 );
or ( \2477_b1 , \2476_b1 , \2323_b1 );
xor ( \2477_b0 , \2476_b0 , w_5656 );
not ( w_5656 , w_5657 );
and ( w_5657 , \2323_b1 , \2323_b0 );
or ( \2478_b1 , \2474_b1 , \2477_b1 );
not ( \2477_b1 , w_5658 );
and ( \2478_b0 , \2474_b0 , w_5659 );
and ( w_5658 , w_5659 , \2477_b0 );
or ( \2479_b1 , \2472_b1 , \2477_b1 );
not ( \2477_b1 , w_5660 );
and ( \2479_b0 , \2472_b0 , w_5661 );
and ( w_5660 , w_5661 , \2477_b0 );
or ( \2481_b1 , \2470_b1 , \2480_b1 );
not ( \2480_b1 , w_5662 );
and ( \2481_b0 , \2470_b0 , w_5663 );
and ( w_5662 , w_5663 , \2480_b0 );
or ( \2482_b1 , \2100_b1 , \2116_b1 );
xor ( \2482_b0 , \2100_b0 , w_5664 );
not ( w_5664 , w_5665 );
and ( w_5665 , \2116_b1 , \2116_b0 );
or ( \2483_b1 , \2482_b1 , \2137_b1 );
xor ( \2483_b0 , \2482_b0 , w_5666 );
not ( w_5666 , w_5667 );
and ( w_5667 , \2137_b1 , \2137_b0 );
or ( \2484_b1 , \2480_b1 , \2483_b1 );
not ( \2483_b1 , w_5668 );
and ( \2484_b0 , \2480_b0 , w_5669 );
and ( w_5668 , w_5669 , \2483_b0 );
or ( \2485_b1 , \2470_b1 , \2483_b1 );
not ( \2483_b1 , w_5670 );
and ( \2485_b0 , \2470_b0 , w_5671 );
and ( w_5670 , w_5671 , \2483_b0 );
or ( \2487_b1 , \2329_b1 , \2339_b1 );
xor ( \2487_b0 , \2329_b0 , w_5672 );
not ( w_5672 , w_5673 );
and ( w_5673 , \2339_b1 , \2339_b0 );
or ( \2488_b1 , \2487_b1 , \2342_b1 );
xor ( \2488_b0 , \2487_b0 , w_5674 );
not ( w_5674 , w_5675 );
and ( w_5675 , \2342_b1 , \2342_b0 );
or ( \2489_b1 , \2486_b1 , \2488_b1 );
not ( \2488_b1 , w_5676 );
and ( \2489_b0 , \2486_b0 , w_5677 );
and ( w_5676 , w_5677 , \2488_b0 );
or ( \2490_b1 , \2347_b1 , \2349_b1 );
xor ( \2490_b0 , \2347_b0 , w_5678 );
not ( w_5678 , w_5679 );
and ( w_5679 , \2349_b1 , \2349_b0 );
or ( \2491_b1 , \2490_b1 , \2352_b1 );
xor ( \2491_b0 , \2490_b0 , w_5680 );
not ( w_5680 , w_5681 );
and ( w_5681 , \2352_b1 , \2352_b0 );
or ( \2492_b1 , \2488_b1 , \2491_b1 );
not ( \2491_b1 , w_5682 );
and ( \2492_b0 , \2488_b0 , w_5683 );
and ( w_5682 , w_5683 , \2491_b0 );
or ( \2493_b1 , \2486_b1 , \2491_b1 );
not ( \2491_b1 , w_5684 );
and ( \2493_b0 , \2486_b0 , w_5685 );
and ( w_5684 , w_5685 , \2491_b0 );
or ( \2495_b1 , \2345_b1 , \2355_b1 );
xor ( \2495_b0 , \2345_b0 , w_5686 );
not ( w_5686 , w_5687 );
and ( w_5687 , \2355_b1 , \2355_b0 );
or ( \2496_b1 , \2495_b1 , \2358_b1 );
xor ( \2496_b0 , \2495_b0 , w_5688 );
not ( w_5688 , w_5689 );
and ( w_5689 , \2358_b1 , \2358_b0 );
or ( \2497_b1 , \2494_b1 , \2496_b1 );
not ( \2496_b1 , w_5690 );
and ( \2497_b0 , \2494_b0 , w_5691 );
and ( w_5690 , w_5691 , \2496_b0 );
or ( \2498_b1 , \2189_b1 , \2199_b1 );
xor ( \2498_b0 , \2189_b0 , w_5692 );
not ( w_5692 , w_5693 );
and ( w_5693 , \2199_b1 , \2199_b0 );
or ( \2499_b1 , \2498_b1 , \2202_b1 );
xor ( \2499_b0 , \2498_b0 , w_5694 );
not ( w_5694 , w_5695 );
and ( w_5695 , \2202_b1 , \2202_b0 );
or ( \2500_b1 , \2496_b1 , \2499_b1 );
not ( \2499_b1 , w_5696 );
and ( \2500_b0 , \2496_b0 , w_5697 );
and ( w_5696 , w_5697 , \2499_b0 );
or ( \2501_b1 , \2494_b1 , \2499_b1 );
not ( \2499_b1 , w_5698 );
and ( \2501_b0 , \2494_b0 , w_5699 );
and ( w_5698 , w_5699 , \2499_b0 );
or ( \2503_b1 , \2367_b1 , \2502_b1 );
not ( \2502_b1 , w_5700 );
and ( \2503_b0 , \2367_b0 , w_5701 );
and ( w_5700 , w_5701 , \2502_b0 );
or ( \2504_b1 , \2367_b1 , \2502_b1 );
xor ( \2504_b0 , \2367_b0 , w_5702 );
not ( w_5702 , w_5703 );
and ( w_5703 , \2502_b1 , \2502_b0 );
or ( \2505_b1 , \2494_b1 , \2496_b1 );
xor ( \2505_b0 , \2494_b0 , w_5704 );
not ( w_5704 , w_5705 );
and ( w_5705 , \2496_b1 , \2496_b0 );
or ( \2506_b1 , \2505_b1 , \2499_b1 );
xor ( \2506_b0 , \2505_b0 , w_5706 );
not ( w_5706 , w_5707 );
and ( w_5707 , \2499_b1 , \2499_b0 );
or ( \2507_b1 , \1299_b1 , \604_b1 );
not ( \604_b1 , w_5708 );
and ( \2507_b0 , \1299_b0 , w_5709 );
and ( w_5708 , w_5709 , \604_b0 );
or ( \2508_b1 , \1194_b1 , \602_b1 );
not ( \602_b1 , w_5710 );
and ( \2508_b0 , \1194_b0 , w_5711 );
and ( w_5710 , w_5711 , \602_b0 );
or ( \2509_b1 , \2507_b1 , w_5713 );
not ( w_5713 , w_5714 );
and ( \2509_b0 , \2507_b0 , w_5715 );
and ( w_5714 ,  , w_5715 );
buf ( w_5713 , \2508_b1 );
not ( w_5713 , w_5716 );
not (  , w_5717 );
and ( w_5716 , w_5717 , \2508_b0 );
or ( \2510_b1 , \2509_b1 , w_5718 );
xor ( \2510_b0 , \2509_b0 , w_5720 );
not ( w_5720 , w_5721 );
and ( w_5721 , w_5718 , w_5719 );
buf ( w_5718 , \561_b1 );
not ( w_5718 , w_5722 );
not ( w_5719 , w_5723 );
and ( w_5722 , w_5723 , \561_b0 );
or ( \2511_b1 , \1422_b1 , \503_b1 );
not ( \503_b1 , w_5724 );
and ( \2511_b0 , \1422_b0 , w_5725 );
and ( w_5724 , w_5725 , \503_b0 );
or ( \2512_b1 , \1304_b1 , \501_b1 );
not ( \501_b1 , w_5726 );
and ( \2512_b0 , \1304_b0 , w_5727 );
and ( w_5726 , w_5727 , \501_b0 );
or ( \2513_b1 , \2511_b1 , w_5729 );
not ( w_5729 , w_5730 );
and ( \2513_b0 , \2511_b0 , w_5731 );
and ( w_5730 ,  , w_5731 );
buf ( w_5729 , \2512_b1 );
not ( w_5729 , w_5732 );
not (  , w_5733 );
and ( w_5732 , w_5733 , \2512_b0 );
or ( \2514_b1 , \2513_b1 , w_5734 );
xor ( \2514_b0 , \2513_b0 , w_5736 );
not ( w_5736 , w_5737 );
and ( w_5737 , w_5734 , w_5735 );
buf ( w_5734 , \455_b1 );
not ( w_5734 , w_5738 );
not ( w_5735 , w_5739 );
and ( w_5738 , w_5739 , \455_b0 );
or ( \2515_b1 , \2510_b1 , \2514_b1 );
not ( \2514_b1 , w_5740 );
and ( \2515_b0 , \2510_b0 , w_5741 );
and ( w_5740 , w_5741 , \2514_b0 );
or ( \2516_b1 , \1770_b1 , \298_b1 );
not ( \298_b1 , w_5742 );
and ( \2516_b0 , \1770_b0 , w_5743 );
and ( w_5742 , w_5743 , \298_b0 );
or ( \2517_b1 , \1537_b1 , \296_b1 );
not ( \296_b1 , w_5744 );
and ( \2517_b0 , \1537_b0 , w_5745 );
and ( w_5744 , w_5745 , \296_b0 );
or ( \2518_b1 , \2516_b1 , w_5747 );
not ( w_5747 , w_5748 );
and ( \2518_b0 , \2516_b0 , w_5749 );
and ( w_5748 ,  , w_5749 );
buf ( w_5747 , \2517_b1 );
not ( w_5747 , w_5750 );
not (  , w_5751 );
and ( w_5750 , w_5751 , \2517_b0 );
or ( \2519_b1 , \2518_b1 , w_5752 );
xor ( \2519_b0 , \2518_b0 , w_5754 );
not ( w_5754 , w_5755 );
and ( w_5755 , w_5752 , w_5753 );
buf ( w_5752 , \303_b1 );
not ( w_5752 , w_5756 );
not ( w_5753 , w_5757 );
and ( w_5756 , w_5757 , \303_b0 );
or ( \2520_b1 , \2514_b1 , \2519_b1 );
not ( \2519_b1 , w_5758 );
and ( \2520_b0 , \2514_b0 , w_5759 );
and ( w_5758 , w_5759 , \2519_b0 );
or ( \2521_b1 , \2510_b1 , \2519_b1 );
not ( \2519_b1 , w_5760 );
and ( \2521_b0 , \2510_b0 , w_5761 );
and ( w_5760 , w_5761 , \2519_b0 );
or ( \2523_b1 , \2023_b1 , \313_b1 );
not ( \313_b1 , w_5762 );
and ( \2523_b0 , \2023_b0 , w_5763 );
and ( w_5762 , w_5763 , \313_b0 );
or ( \2524_b1 , \1778_b1 , \311_b1 );
not ( \311_b1 , w_5764 );
and ( \2524_b0 , \1778_b0 , w_5765 );
and ( w_5764 , w_5765 , \311_b0 );
or ( \2525_b1 , \2523_b1 , w_5767 );
not ( w_5767 , w_5768 );
and ( \2525_b0 , \2523_b0 , w_5769 );
and ( w_5768 ,  , w_5769 );
buf ( w_5767 , \2524_b1 );
not ( w_5767 , w_5770 );
not (  , w_5771 );
and ( w_5770 , w_5771 , \2524_b0 );
or ( \2526_b1 , \2525_b1 , w_5772 );
xor ( \2526_b0 , \2525_b0 , w_5774 );
not ( w_5774 , w_5775 );
and ( w_5775 , w_5772 , w_5773 );
buf ( w_5772 , \320_b1 );
not ( w_5772 , w_5776 );
not ( w_5773 , w_5777 );
and ( w_5776 , w_5777 , \320_b0 );
or ( \2527_b1 , \2161_b1 , \331_b1 );
not ( \331_b1 , w_5778 );
and ( \2527_b0 , \2161_b0 , w_5779 );
and ( w_5778 , w_5779 , \331_b0 );
or ( \2528_b1 , \2028_b1 , \329_b1 );
not ( \329_b1 , w_5780 );
and ( \2528_b0 , \2028_b0 , w_5781 );
and ( w_5780 , w_5781 , \329_b0 );
or ( \2529_b1 , \2527_b1 , w_5783 );
not ( w_5783 , w_5784 );
and ( \2529_b0 , \2527_b0 , w_5785 );
and ( w_5784 ,  , w_5785 );
buf ( w_5783 , \2528_b1 );
not ( w_5783 , w_5786 );
not (  , w_5787 );
and ( w_5786 , w_5787 , \2528_b0 );
or ( \2530_b1 , \2529_b1 , w_5788 );
xor ( \2530_b0 , \2529_b0 , w_5790 );
not ( w_5790 , w_5791 );
and ( w_5791 , w_5788 , w_5789 );
buf ( w_5788 , \338_b1 );
not ( w_5788 , w_5792 );
not ( w_5789 , w_5793 );
and ( w_5792 , w_5793 , \338_b0 );
or ( \2531_b1 , \2526_b1 , \2530_b1 );
not ( \2530_b1 , w_5794 );
and ( \2531_b0 , \2526_b0 , w_5795 );
and ( w_5794 , w_5795 , \2530_b0 );
buf ( \2532_b1 , RIb4bc108_93_b1 );
buf ( \2532_b0 , RIb4bc108_93_b0 );
or ( \2533_b1 , \2532_b1 , \351_b1 );
not ( \351_b1 , w_5796 );
and ( \2533_b0 , \2532_b0 , w_5797 );
and ( w_5796 , w_5797 , \351_b0 );
or ( \2534_b1 , \2305_b1 , \349_b1 );
not ( \349_b1 , w_5798 );
and ( \2534_b0 , \2305_b0 , w_5799 );
and ( w_5798 , w_5799 , \349_b0 );
or ( \2535_b1 , \2533_b1 , w_5801 );
not ( w_5801 , w_5802 );
and ( \2535_b0 , \2533_b0 , w_5803 );
and ( w_5802 ,  , w_5803 );
buf ( w_5801 , \2534_b1 );
not ( w_5801 , w_5804 );
not (  , w_5805 );
and ( w_5804 , w_5805 , \2534_b0 );
or ( \2536_b1 , \2535_b1 , w_5806 );
xor ( \2536_b0 , \2535_b0 , w_5808 );
not ( w_5808 , w_5809 );
and ( w_5809 , w_5806 , w_5807 );
buf ( w_5806 , \358_b1 );
not ( w_5806 , w_5810 );
not ( w_5807 , w_5811 );
and ( w_5810 , w_5811 , \358_b0 );
or ( \2537_b1 , \2530_b1 , \2536_b1 );
not ( \2536_b1 , w_5812 );
and ( \2537_b0 , \2530_b0 , w_5813 );
and ( w_5812 , w_5813 , \2536_b0 );
or ( \2538_b1 , \2526_b1 , \2536_b1 );
not ( \2536_b1 , w_5814 );
and ( \2538_b0 , \2526_b0 , w_5815 );
and ( w_5814 , w_5815 , \2536_b0 );
or ( \2540_b1 , \2522_b1 , \2539_b1 );
not ( \2539_b1 , w_5816 );
and ( \2540_b0 , \2522_b0 , w_5817 );
and ( w_5816 , w_5817 , \2539_b0 );
buf ( \2541_b1 , RIb4bc090_94_b1 );
buf ( \2541_b0 , RIb4bc090_94_b0 );
or ( \2542_b1 , \2541_b1 , \345_b1 );
not ( \345_b1 , w_5818 );
and ( \2542_b0 , \2541_b0 , w_5819 );
and ( w_5818 , w_5819 , \345_b0 );
buf ( \2543_b1 , \2542_b1 );
buf ( \2543_b0 , \2542_b0 );
or ( \2544_b1 , \2539_b1 , \2543_b1 );
not ( \2543_b1 , w_5820 );
and ( \2544_b0 , \2539_b0 , w_5821 );
and ( w_5820 , w_5821 , \2543_b0 );
or ( \2545_b1 , \2522_b1 , \2543_b1 );
not ( \2543_b1 , w_5822 );
and ( \2545_b0 , \2522_b0 , w_5823 );
and ( w_5822 , w_5823 , \2543_b0 );
or ( \2547_b1 , \2121_b1 , \2369_b1 );
xor ( \2547_b0 , \2121_b0 , w_5824 );
not ( w_5824 , w_5825 );
and ( w_5825 , \2369_b1 , \2369_b0 );
or ( \2548_b1 , \2369_b1 , \2371_b1 );
xor ( \2548_b0 , \2369_b0 , w_5826 );
not ( w_5826 , w_5827 );
and ( w_5827 , \2371_b1 , \2371_b0 );
buf ( \2549_b1 , \2548_b1 );
not ( \2549_b1 , w_5828 );
not ( \2549_b0 , w_5829 );
and ( w_5828 , w_5829 , \2548_b0 );
or ( \2550_b1 , \2547_b1 , \2549_b1 );
not ( \2549_b1 , w_5830 );
and ( \2550_b0 , \2547_b0 , w_5831 );
and ( w_5830 , w_5831 , \2549_b0 );
or ( \2551_b1 , \159_b1 , \2550_b1 );
not ( \2550_b1 , w_5832 );
and ( \2551_b0 , \159_b0 , w_5833 );
and ( w_5832 , w_5833 , \2550_b0 );
buf ( \2552_b1 , \2551_b1 );
not ( \2552_b1 , w_5834 );
not ( \2552_b0 , w_5835 );
and ( w_5834 , w_5835 , \2551_b0 );
or ( \2553_b1 , \2552_b1 , w_5836 );
xor ( \2553_b0 , \2552_b0 , w_5838 );
not ( w_5838 , w_5839 );
and ( w_5839 , w_5836 , w_5837 );
buf ( w_5836 , \2374_b1 );
not ( w_5836 , w_5840 );
not ( w_5837 , w_5841 );
and ( w_5840 , w_5841 , \2374_b0 );
or ( \2554_b1 , \305_b1 , \2261_b1 );
not ( \2261_b1 , w_5842 );
and ( \2554_b0 , \305_b0 , w_5843 );
and ( w_5842 , w_5843 , \2261_b0 );
or ( \2555_b1 , \315_b1 , \2259_b1 );
not ( \2259_b1 , w_5844 );
and ( \2555_b0 , \315_b0 , w_5845 );
and ( w_5844 , w_5845 , \2259_b0 );
or ( \2556_b1 , \2554_b1 , w_5847 );
not ( w_5847 , w_5848 );
and ( \2556_b0 , \2554_b0 , w_5849 );
and ( w_5848 ,  , w_5849 );
buf ( w_5847 , \2555_b1 );
not ( w_5847 , w_5850 );
not (  , w_5851 );
and ( w_5850 , w_5851 , \2555_b0 );
or ( \2557_b1 , \2556_b1 , w_5852 );
xor ( \2557_b0 , \2556_b0 , w_5854 );
not ( w_5854 , w_5855 );
and ( w_5855 , w_5852 , w_5853 );
buf ( w_5852 , \2124_b1 );
not ( w_5852 , w_5856 );
not ( w_5853 , w_5857 );
and ( w_5856 , w_5857 , \2124_b0 );
or ( \2558_b1 , \2553_b1 , \2557_b1 );
not ( \2557_b1 , w_5858 );
and ( \2558_b0 , \2553_b0 , w_5859 );
and ( w_5858 , w_5859 , \2557_b0 );
or ( \2559_b1 , \323_b1 , \1955_b1 );
not ( \1955_b1 , w_5860 );
and ( \2559_b0 , \323_b0 , w_5861 );
and ( w_5860 , w_5861 , \1955_b0 );
or ( \2560_b1 , \333_b1 , \1953_b1 );
not ( \1953_b1 , w_5862 );
and ( \2560_b0 , \333_b0 , w_5863 );
and ( w_5862 , w_5863 , \1953_b0 );
or ( \2561_b1 , \2559_b1 , w_5865 );
not ( w_5865 , w_5866 );
and ( \2561_b0 , \2559_b0 , w_5867 );
and ( w_5866 ,  , w_5867 );
buf ( w_5865 , \2560_b1 );
not ( w_5865 , w_5868 );
not (  , w_5869 );
and ( w_5868 , w_5869 , \2560_b0 );
or ( \2562_b1 , \2561_b1 , w_5870 );
xor ( \2562_b0 , \2561_b0 , w_5872 );
not ( w_5872 , w_5873 );
and ( w_5873 , w_5870 , w_5871 );
buf ( w_5870 , \1835_b1 );
not ( w_5870 , w_5874 );
not ( w_5871 , w_5875 );
and ( w_5874 , w_5875 , \1835_b0 );
or ( \2563_b1 , \2557_b1 , \2562_b1 );
not ( \2562_b1 , w_5876 );
and ( \2563_b0 , \2557_b0 , w_5877 );
and ( w_5876 , w_5877 , \2562_b0 );
or ( \2564_b1 , \2553_b1 , \2562_b1 );
not ( \2562_b1 , w_5878 );
and ( \2564_b0 , \2553_b0 , w_5879 );
and ( w_5878 , w_5879 , \2562_b0 );
or ( \2566_b1 , \343_b1 , \1742_b1 );
not ( \1742_b1 , w_5880 );
and ( \2566_b0 , \343_b0 , w_5881 );
and ( w_5880 , w_5881 , \1742_b0 );
or ( \2567_b1 , \353_b1 , \1740_b1 );
not ( \1740_b1 , w_5882 );
and ( \2567_b0 , \353_b0 , w_5883 );
and ( w_5882 , w_5883 , \1740_b0 );
or ( \2568_b1 , \2566_b1 , w_5885 );
not ( w_5885 , w_5886 );
and ( \2568_b0 , \2566_b0 , w_5887 );
and ( w_5886 ,  , w_5887 );
buf ( w_5885 , \2567_b1 );
not ( w_5885 , w_5888 );
not (  , w_5889 );
and ( w_5888 , w_5889 , \2567_b0 );
or ( \2569_b1 , \2568_b1 , w_5890 );
xor ( \2569_b0 , \2568_b0 , w_5892 );
not ( w_5892 , w_5893 );
and ( w_5893 , w_5890 , w_5891 );
buf ( w_5890 , \1610_b1 );
not ( w_5890 , w_5894 );
not ( w_5891 , w_5895 );
and ( w_5894 , w_5895 , \1610_b0 );
or ( \2570_b1 , \444_b1 , \1476_b1 );
not ( \1476_b1 , w_5896 );
and ( \2570_b0 , \444_b0 , w_5897 );
and ( w_5896 , w_5897 , \1476_b0 );
or ( \2571_b1 , \360_b1 , \1474_b1 );
not ( \1474_b1 , w_5898 );
and ( \2571_b0 , \360_b0 , w_5899 );
and ( w_5898 , w_5899 , \1474_b0 );
or ( \2572_b1 , \2570_b1 , w_5901 );
not ( w_5901 , w_5902 );
and ( \2572_b0 , \2570_b0 , w_5903 );
and ( w_5902 ,  , w_5903 );
buf ( w_5901 , \2571_b1 );
not ( w_5901 , w_5904 );
not (  , w_5905 );
and ( w_5904 , w_5905 , \2571_b0 );
or ( \2573_b1 , \2572_b1 , w_5906 );
xor ( \2573_b0 , \2572_b0 , w_5908 );
not ( w_5908 , w_5909 );
and ( w_5909 , w_5906 , w_5907 );
buf ( w_5906 , \1363_b1 );
not ( w_5906 , w_5910 );
not ( w_5907 , w_5911 );
and ( w_5910 , w_5911 , \1363_b0 );
or ( \2574_b1 , \2569_b1 , \2573_b1 );
not ( \2573_b1 , w_5912 );
and ( \2574_b0 , \2569_b0 , w_5913 );
and ( w_5912 , w_5913 , \2573_b0 );
or ( \2575_b1 , \593_b1 , \1280_b1 );
not ( \1280_b1 , w_5914 );
and ( \2575_b0 , \593_b0 , w_5915 );
and ( w_5914 , w_5915 , \1280_b0 );
or ( \2576_b1 , \495_b1 , \1278_b1 );
not ( \1278_b1 , w_5916 );
and ( \2576_b0 , \495_b0 , w_5917 );
and ( w_5916 , w_5917 , \1278_b0 );
or ( \2577_b1 , \2575_b1 , w_5919 );
not ( w_5919 , w_5920 );
and ( \2577_b0 , \2575_b0 , w_5921 );
and ( w_5920 ,  , w_5921 );
buf ( w_5919 , \2576_b1 );
not ( w_5919 , w_5922 );
not (  , w_5923 );
and ( w_5922 , w_5923 , \2576_b0 );
or ( \2578_b1 , \2577_b1 , w_5924 );
xor ( \2578_b0 , \2577_b0 , w_5926 );
not ( w_5926 , w_5927 );
and ( w_5927 , w_5924 , w_5925 );
buf ( w_5924 , \1177_b1 );
not ( w_5924 , w_5928 );
not ( w_5925 , w_5929 );
and ( w_5928 , w_5929 , \1177_b0 );
or ( \2579_b1 , \2573_b1 , \2578_b1 );
not ( \2578_b1 , w_5930 );
and ( \2579_b0 , \2573_b0 , w_5931 );
and ( w_5930 , w_5931 , \2578_b0 );
or ( \2580_b1 , \2569_b1 , \2578_b1 );
not ( \2578_b1 , w_5932 );
and ( \2580_b0 , \2569_b0 , w_5933 );
and ( w_5932 , w_5933 , \2578_b0 );
or ( \2582_b1 , \2565_b1 , \2581_b1 );
not ( \2581_b1 , w_5934 );
and ( \2582_b0 , \2565_b0 , w_5935 );
and ( w_5934 , w_5935 , \2581_b0 );
or ( \2583_b1 , \703_b1 , \1062_b1 );
not ( \1062_b1 , w_5936 );
and ( \2583_b0 , \703_b0 , w_5937 );
and ( w_5936 , w_5937 , \1062_b0 );
or ( \2584_b1 , \621_b1 , \1060_b1 );
not ( \1060_b1 , w_5938 );
and ( \2584_b0 , \621_b0 , w_5939 );
and ( w_5938 , w_5939 , \1060_b0 );
or ( \2585_b1 , \2583_b1 , w_5941 );
not ( w_5941 , w_5942 );
and ( \2585_b0 , \2583_b0 , w_5943 );
and ( w_5942 ,  , w_5943 );
buf ( w_5941 , \2584_b1 );
not ( w_5941 , w_5944 );
not (  , w_5945 );
and ( w_5944 , w_5945 , \2584_b0 );
or ( \2586_b1 , \2585_b1 , w_5946 );
xor ( \2586_b0 , \2585_b0 , w_5948 );
not ( w_5948 , w_5949 );
and ( w_5949 , w_5946 , w_5947 );
buf ( w_5946 , \984_b1 );
not ( w_5946 , w_5950 );
not ( w_5947 , w_5951 );
and ( w_5950 , w_5951 , \984_b0 );
or ( \2587_b1 , \841_b1 , \912_b1 );
not ( \912_b1 , w_5952 );
and ( \2587_b0 , \841_b0 , w_5953 );
and ( w_5952 , w_5953 , \912_b0 );
or ( \2588_b1 , \777_b1 , \910_b1 );
not ( \910_b1 , w_5954 );
and ( \2588_b0 , \777_b0 , w_5955 );
and ( w_5954 , w_5955 , \910_b0 );
or ( \2589_b1 , \2587_b1 , w_5957 );
not ( w_5957 , w_5958 );
and ( \2589_b0 , \2587_b0 , w_5959 );
and ( w_5958 ,  , w_5959 );
buf ( w_5957 , \2588_b1 );
not ( w_5957 , w_5960 );
not (  , w_5961 );
and ( w_5960 , w_5961 , \2588_b0 );
or ( \2590_b1 , \2589_b1 , w_5962 );
xor ( \2590_b0 , \2589_b0 , w_5964 );
not ( w_5964 , w_5965 );
and ( w_5965 , w_5962 , w_5963 );
buf ( w_5962 , \818_b1 );
not ( w_5962 , w_5966 );
not ( w_5963 , w_5967 );
and ( w_5966 , w_5967 , \818_b0 );
or ( \2591_b1 , \2586_b1 , \2590_b1 );
not ( \2590_b1 , w_5968 );
and ( \2591_b0 , \2586_b0 , w_5969 );
and ( w_5968 , w_5969 , \2590_b0 );
or ( \2592_b1 , \1104_b1 , \740_b1 );
not ( \740_b1 , w_5970 );
and ( \2592_b0 , \1104_b0 , w_5971 );
and ( w_5970 , w_5971 , \740_b0 );
or ( \2593_b1 , \904_b1 , \738_b1 );
not ( \738_b1 , w_5972 );
and ( \2593_b0 , \904_b0 , w_5973 );
and ( w_5972 , w_5973 , \738_b0 );
or ( \2594_b1 , \2592_b1 , w_5975 );
not ( w_5975 , w_5976 );
and ( \2594_b0 , \2592_b0 , w_5977 );
and ( w_5976 ,  , w_5977 );
buf ( w_5975 , \2593_b1 );
not ( w_5975 , w_5978 );
not (  , w_5979 );
and ( w_5978 , w_5979 , \2593_b0 );
or ( \2595_b1 , \2594_b1 , w_5980 );
xor ( \2595_b0 , \2594_b0 , w_5982 );
not ( w_5982 , w_5983 );
and ( w_5983 , w_5980 , w_5981 );
buf ( w_5980 , \668_b1 );
not ( w_5980 , w_5984 );
not ( w_5981 , w_5985 );
and ( w_5984 , w_5985 , \668_b0 );
or ( \2596_b1 , \2590_b1 , \2595_b1 );
not ( \2595_b1 , w_5986 );
and ( \2596_b0 , \2590_b0 , w_5987 );
and ( w_5986 , w_5987 , \2595_b0 );
or ( \2597_b1 , \2586_b1 , \2595_b1 );
not ( \2595_b1 , w_5988 );
and ( \2597_b0 , \2586_b0 , w_5989 );
and ( w_5988 , w_5989 , \2595_b0 );
or ( \2599_b1 , \2581_b1 , \2598_b1 );
not ( \2598_b1 , w_5990 );
and ( \2599_b0 , \2581_b0 , w_5991 );
and ( w_5990 , w_5991 , \2598_b0 );
or ( \2600_b1 , \2565_b1 , \2598_b1 );
not ( \2598_b1 , w_5992 );
and ( \2600_b0 , \2565_b0 , w_5993 );
and ( w_5992 , w_5993 , \2598_b0 );
or ( \2602_b1 , \2546_b1 , \2601_b1 );
not ( \2601_b1 , w_5994 );
and ( \2602_b0 , \2546_b0 , w_5995 );
and ( w_5994 , w_5995 , \2601_b0 );
or ( \2603_b1 , \2532_b1 , \345_b1 );
not ( \345_b1 , w_5996 );
and ( \2603_b0 , \2532_b0 , w_5997 );
and ( w_5996 , w_5997 , \345_b0 );
or ( \2604_b1 , \2438_b1 , \2442_b1 );
xor ( \2604_b0 , \2438_b0 , w_5998 );
not ( w_5998 , w_5999 );
and ( w_5999 , \2442_b1 , \2442_b0 );
or ( \2605_b1 , \2604_b1 , \2447_b1 );
xor ( \2605_b0 , \2604_b0 , w_6000 );
not ( w_6000 , w_6001 );
and ( w_6001 , \2447_b1 , \2447_b0 );
or ( \2606_b1 , \2603_b1 , \2605_b1 );
not ( \2605_b1 , w_6002 );
and ( \2606_b0 , \2603_b0 , w_6003 );
and ( w_6002 , w_6003 , \2605_b0 );
or ( \2607_b1 , \2454_b1 , \2458_b1 );
xor ( \2607_b0 , \2454_b0 , w_6004 );
not ( w_6004 , w_6005 );
and ( w_6005 , \2458_b1 , \2458_b0 );
or ( \2608_b1 , \2607_b1 , \2463_b1 );
xor ( \2608_b0 , \2607_b0 , w_6006 );
not ( w_6006 , w_6007 );
and ( w_6007 , \2463_b1 , \2463_b0 );
or ( \2609_b1 , \2605_b1 , \2608_b1 );
not ( \2608_b1 , w_6008 );
and ( \2609_b0 , \2605_b0 , w_6009 );
and ( w_6008 , w_6009 , \2608_b0 );
or ( \2610_b1 , \2603_b1 , \2608_b1 );
not ( \2608_b1 , w_6010 );
and ( \2610_b0 , \2603_b0 , w_6011 );
and ( w_6010 , w_6011 , \2608_b0 );
or ( \2612_b1 , \2601_b1 , \2611_b1 );
not ( \2611_b1 , w_6012 );
and ( \2612_b0 , \2601_b0 , w_6013 );
and ( w_6012 , w_6013 , \2611_b0 );
or ( \2613_b1 , \2546_b1 , \2611_b1 );
not ( \2611_b1 , w_6014 );
and ( \2613_b0 , \2546_b0 , w_6015 );
and ( w_6014 , w_6015 , \2611_b0 );
or ( \2615_b1 , \2375_b1 , \2379_b1 );
xor ( \2615_b0 , \2375_b0 , w_6016 );
not ( w_6016 , w_6017 );
and ( w_6017 , \2379_b1 , \2379_b0 );
or ( \2616_b1 , \2615_b1 , \2384_b1 );
xor ( \2616_b0 , \2615_b0 , w_6018 );
not ( w_6018 , w_6019 );
and ( w_6019 , \2384_b1 , \2384_b0 );
or ( \2617_b1 , \2391_b1 , \2395_b1 );
xor ( \2617_b0 , \2391_b0 , w_6020 );
not ( w_6020 , w_6021 );
and ( w_6021 , \2395_b1 , \2395_b0 );
or ( \2618_b1 , \2617_b1 , \2400_b1 );
xor ( \2618_b0 , \2617_b0 , w_6022 );
not ( w_6022 , w_6023 );
and ( w_6023 , \2400_b1 , \2400_b0 );
or ( \2619_b1 , \2616_b1 , \2618_b1 );
not ( \2618_b1 , w_6024 );
and ( \2619_b0 , \2616_b0 , w_6025 );
and ( w_6024 , w_6025 , \2618_b0 );
or ( \2620_b1 , \2408_b1 , \2412_b1 );
xor ( \2620_b0 , \2408_b0 , w_6026 );
not ( w_6026 , w_6027 );
and ( w_6027 , \2412_b1 , \2412_b0 );
or ( \2621_b1 , \2620_b1 , \2417_b1 );
xor ( \2621_b0 , \2620_b0 , w_6028 );
not ( w_6028 , w_6029 );
and ( w_6029 , \2417_b1 , \2417_b0 );
or ( \2622_b1 , \2618_b1 , \2621_b1 );
not ( \2621_b1 , w_6030 );
and ( \2622_b0 , \2618_b0 , w_6031 );
and ( w_6030 , w_6031 , \2621_b0 );
or ( \2623_b1 , \2616_b1 , \2621_b1 );
not ( \2621_b1 , w_6032 );
and ( \2623_b0 , \2616_b0 , w_6033 );
and ( w_6032 , w_6033 , \2621_b0 );
or ( \2625_b1 , \2244_b1 , \2248_b1 );
xor ( \2625_b0 , \2244_b0 , w_6034 );
not ( w_6034 , w_6035 );
and ( w_6035 , \2248_b1 , \2248_b0 );
or ( \2626_b1 , \2625_b1 , \2253_b1 );
xor ( \2626_b0 , \2625_b0 , w_6036 );
not ( w_6036 , w_6037 );
and ( w_6037 , \2253_b1 , \2253_b0 );
or ( \2627_b1 , \2624_b1 , \2626_b1 );
not ( \2626_b1 , w_6038 );
and ( \2627_b0 , \2624_b0 , w_6039 );
and ( w_6038 , w_6039 , \2626_b0 );
or ( \2628_b1 , \2264_b1 , \2268_b1 );
xor ( \2628_b0 , \2264_b0 , w_6040 );
not ( w_6040 , w_6041 );
and ( w_6041 , \2268_b1 , \2268_b0 );
or ( \2629_b1 , \2628_b1 , \2273_b1 );
xor ( \2629_b0 , \2628_b0 , w_6042 );
not ( w_6042 , w_6043 );
and ( w_6043 , \2273_b1 , \2273_b0 );
or ( \2630_b1 , \2626_b1 , \2629_b1 );
not ( \2629_b1 , w_6044 );
and ( \2630_b0 , \2626_b0 , w_6045 );
and ( w_6044 , w_6045 , \2629_b0 );
or ( \2631_b1 , \2624_b1 , \2629_b1 );
not ( \2629_b1 , w_6046 );
and ( \2631_b0 , \2624_b0 , w_6047 );
and ( w_6046 , w_6047 , \2629_b0 );
or ( \2633_b1 , \2614_b1 , \2632_b1 );
not ( \2632_b1 , w_6048 );
and ( \2633_b0 , \2614_b0 , w_6049 );
and ( w_6048 , w_6049 , \2632_b0 );
or ( \2634_b1 , \2387_b1 , \2403_b1 );
xor ( \2634_b0 , \2387_b0 , w_6050 );
not ( w_6050 , w_6051 );
and ( w_6051 , \2403_b1 , \2403_b0 );
or ( \2635_b1 , \2634_b1 , \2420_b1 );
xor ( \2635_b0 , \2634_b0 , w_6052 );
not ( w_6052 , w_6053 );
and ( w_6053 , \2420_b1 , \2420_b0 );
or ( \2636_b1 , \2425_b1 , \2427_b1 );
xor ( \2636_b0 , \2425_b0 , w_6054 );
not ( w_6054 , w_6055 );
and ( w_6055 , \2427_b1 , \2427_b0 );
or ( \2637_b1 , \2636_b1 , \2430_b1 );
xor ( \2637_b0 , \2636_b0 , w_6056 );
not ( w_6056 , w_6057 );
and ( w_6057 , \2430_b1 , \2430_b0 );
or ( \2638_b1 , \2635_b1 , \2637_b1 );
not ( \2637_b1 , w_6058 );
and ( \2638_b0 , \2635_b0 , w_6059 );
and ( w_6058 , w_6059 , \2637_b0 );
or ( \2639_b1 , \2450_b1 , w_6060 );
xor ( \2639_b0 , \2450_b0 , w_6062 );
not ( w_6062 , w_6063 );
and ( w_6063 , w_6060 , w_6061 );
buf ( w_6060 , \2466_b1 );
not ( w_6060 , w_6064 );
not ( w_6061 , w_6065 );
and ( w_6064 , w_6065 , \2466_b0 );
or ( \2640_b1 , \2637_b1 , \2639_b1 );
not ( \2639_b1 , w_6066 );
and ( \2640_b0 , \2637_b0 , w_6067 );
and ( w_6066 , w_6067 , \2639_b0 );
or ( \2641_b1 , \2635_b1 , \2639_b1 );
not ( \2639_b1 , w_6068 );
and ( \2641_b0 , \2635_b0 , w_6069 );
and ( w_6068 , w_6069 , \2639_b0 );
or ( \2643_b1 , \2632_b1 , \2642_b1 );
not ( \2642_b1 , w_6070 );
and ( \2643_b0 , \2632_b0 , w_6071 );
and ( w_6070 , w_6071 , \2642_b0 );
or ( \2644_b1 , \2614_b1 , \2642_b1 );
not ( \2642_b1 , w_6072 );
and ( \2644_b0 , \2614_b0 , w_6073 );
and ( w_6072 , w_6073 , \2642_b0 );
or ( \2646_b1 , \2240_b1 , \2256_b1 );
xor ( \2646_b0 , \2240_b0 , w_6074 );
not ( w_6074 , w_6075 );
and ( w_6075 , \2256_b1 , \2256_b0 );
or ( \2647_b1 , \2646_b1 , \2276_b1 );
xor ( \2647_b0 , \2646_b0 , w_6076 );
not ( w_6076 , w_6077 );
and ( w_6077 , \2276_b1 , \2276_b0 );
or ( \2648_b1 , \2423_b1 , \2433_b1 );
xor ( \2648_b0 , \2423_b0 , w_6078 );
not ( w_6078 , w_6079 );
and ( w_6079 , \2433_b1 , \2433_b0 );
or ( \2649_b1 , \2648_b1 , \2467_b1 );
xor ( \2649_b0 , \2648_b0 , w_6080 );
not ( w_6080 , w_6081 );
and ( w_6081 , \2467_b1 , \2467_b0 );
or ( \2650_b1 , \2647_b1 , \2649_b1 );
not ( \2649_b1 , w_6082 );
and ( \2650_b0 , \2647_b0 , w_6083 );
and ( w_6082 , w_6083 , \2649_b0 );
or ( \2651_b1 , \2472_b1 , \2474_b1 );
xor ( \2651_b0 , \2472_b0 , w_6084 );
not ( w_6084 , w_6085 );
and ( w_6085 , \2474_b1 , \2474_b0 );
or ( \2652_b1 , \2651_b1 , \2477_b1 );
xor ( \2652_b0 , \2651_b0 , w_6086 );
not ( w_6086 , w_6087 );
and ( w_6087 , \2477_b1 , \2477_b0 );
or ( \2653_b1 , \2649_b1 , \2652_b1 );
not ( \2652_b1 , w_6088 );
and ( \2653_b0 , \2649_b0 , w_6089 );
and ( w_6088 , w_6089 , \2652_b0 );
or ( \2654_b1 , \2647_b1 , \2652_b1 );
not ( \2652_b1 , w_6090 );
and ( \2654_b0 , \2647_b0 , w_6091 );
and ( w_6090 , w_6091 , \2652_b0 );
or ( \2656_b1 , \2645_b1 , \2655_b1 );
not ( \2655_b1 , w_6092 );
and ( \2656_b0 , \2645_b0 , w_6093 );
and ( w_6092 , w_6093 , \2655_b0 );
or ( \2657_b1 , \2331_b1 , \2333_b1 );
xor ( \2657_b0 , \2331_b0 , w_6094 );
not ( w_6094 , w_6095 );
and ( w_6095 , \2333_b1 , \2333_b0 );
or ( \2658_b1 , \2657_b1 , \2336_b1 );
xor ( \2658_b0 , \2657_b0 , w_6096 );
not ( w_6096 , w_6097 );
and ( w_6097 , \2336_b1 , \2336_b0 );
or ( \2659_b1 , \2655_b1 , \2658_b1 );
not ( \2658_b1 , w_6098 );
and ( \2659_b0 , \2655_b0 , w_6099 );
and ( w_6098 , w_6099 , \2658_b0 );
or ( \2660_b1 , \2645_b1 , \2658_b1 );
not ( \2658_b1 , w_6100 );
and ( \2660_b0 , \2645_b0 , w_6101 );
and ( w_6100 , w_6101 , \2658_b0 );
or ( \2662_b1 , \2279_b1 , \2315_b1 );
xor ( \2662_b0 , \2279_b0 , w_6102 );
not ( w_6102 , w_6103 );
and ( w_6103 , \2315_b1 , \2315_b0 );
or ( \2663_b1 , \2662_b1 , \2326_b1 );
xor ( \2663_b0 , \2662_b0 , w_6104 );
not ( w_6104 , w_6105 );
and ( w_6105 , \2326_b1 , \2326_b0 );
or ( \2664_b1 , \2470_b1 , \2480_b1 );
xor ( \2664_b0 , \2470_b0 , w_6106 );
not ( w_6106 , w_6107 );
and ( w_6107 , \2480_b1 , \2480_b0 );
or ( \2665_b1 , \2664_b1 , \2483_b1 );
xor ( \2665_b0 , \2664_b0 , w_6108 );
not ( w_6108 , w_6109 );
and ( w_6109 , \2483_b1 , \2483_b0 );
or ( \2666_b1 , \2663_b1 , \2665_b1 );
not ( \2665_b1 , w_6110 );
and ( \2666_b0 , \2663_b0 , w_6111 );
and ( w_6110 , w_6111 , \2665_b0 );
or ( \2667_b1 , \2661_b1 , \2666_b1 );
not ( \2666_b1 , w_6112 );
and ( \2667_b0 , \2661_b0 , w_6113 );
and ( w_6112 , w_6113 , \2666_b0 );
or ( \2668_b1 , \2486_b1 , \2488_b1 );
xor ( \2668_b0 , \2486_b0 , w_6114 );
not ( w_6114 , w_6115 );
and ( w_6115 , \2488_b1 , \2488_b0 );
or ( \2669_b1 , \2668_b1 , \2491_b1 );
xor ( \2669_b0 , \2668_b0 , w_6116 );
not ( w_6116 , w_6117 );
and ( w_6117 , \2491_b1 , \2491_b0 );
or ( \2670_b1 , \2666_b1 , \2669_b1 );
not ( \2669_b1 , w_6118 );
and ( \2670_b0 , \2666_b0 , w_6119 );
and ( w_6118 , w_6119 , \2669_b0 );
or ( \2671_b1 , \2661_b1 , \2669_b1 );
not ( \2669_b1 , w_6120 );
and ( \2671_b0 , \2661_b0 , w_6121 );
and ( w_6120 , w_6121 , \2669_b0 );
or ( \2673_b1 , \2506_b1 , \2672_b1 );
not ( \2672_b1 , w_6122 );
and ( \2673_b0 , \2506_b0 , w_6123 );
and ( w_6122 , w_6123 , \2672_b0 );
or ( \2674_b1 , \2506_b1 , \2672_b1 );
xor ( \2674_b0 , \2506_b0 , w_6124 );
not ( w_6124 , w_6125 );
and ( w_6125 , \2672_b1 , \2672_b0 );
or ( \2675_b1 , \2661_b1 , \2666_b1 );
xor ( \2675_b0 , \2661_b0 , w_6126 );
not ( w_6126 , w_6127 );
and ( w_6127 , \2666_b1 , \2666_b0 );
or ( \2676_b1 , \2675_b1 , \2669_b1 );
xor ( \2676_b0 , \2675_b0 , w_6128 );
not ( w_6128 , w_6129 );
and ( w_6129 , \2669_b1 , \2669_b0 );
or ( \2677_b1 , \621_b1 , \1280_b1 );
not ( \1280_b1 , w_6130 );
and ( \2677_b0 , \621_b0 , w_6131 );
and ( w_6130 , w_6131 , \1280_b0 );
or ( \2678_b1 , \593_b1 , \1278_b1 );
not ( \1278_b1 , w_6132 );
and ( \2678_b0 , \593_b0 , w_6133 );
and ( w_6132 , w_6133 , \1278_b0 );
or ( \2679_b1 , \2677_b1 , w_6135 );
not ( w_6135 , w_6136 );
and ( \2679_b0 , \2677_b0 , w_6137 );
and ( w_6136 ,  , w_6137 );
buf ( w_6135 , \2678_b1 );
not ( w_6135 , w_6138 );
not (  , w_6139 );
and ( w_6138 , w_6139 , \2678_b0 );
or ( \2680_b1 , \2679_b1 , w_6140 );
xor ( \2680_b0 , \2679_b0 , w_6142 );
not ( w_6142 , w_6143 );
and ( w_6143 , w_6140 , w_6141 );
buf ( w_6140 , \1177_b1 );
not ( w_6140 , w_6144 );
not ( w_6141 , w_6145 );
and ( w_6144 , w_6145 , \1177_b0 );
or ( \2681_b1 , \777_b1 , \1062_b1 );
not ( \1062_b1 , w_6146 );
and ( \2681_b0 , \777_b0 , w_6147 );
and ( w_6146 , w_6147 , \1062_b0 );
or ( \2682_b1 , \703_b1 , \1060_b1 );
not ( \1060_b1 , w_6148 );
and ( \2682_b0 , \703_b0 , w_6149 );
and ( w_6148 , w_6149 , \1060_b0 );
or ( \2683_b1 , \2681_b1 , w_6151 );
not ( w_6151 , w_6152 );
and ( \2683_b0 , \2681_b0 , w_6153 );
and ( w_6152 ,  , w_6153 );
buf ( w_6151 , \2682_b1 );
not ( w_6151 , w_6154 );
not (  , w_6155 );
and ( w_6154 , w_6155 , \2682_b0 );
or ( \2684_b1 , \2683_b1 , w_6156 );
xor ( \2684_b0 , \2683_b0 , w_6158 );
not ( w_6158 , w_6159 );
and ( w_6159 , w_6156 , w_6157 );
buf ( w_6156 , \984_b1 );
not ( w_6156 , w_6160 );
not ( w_6157 , w_6161 );
and ( w_6160 , w_6161 , \984_b0 );
or ( \2685_b1 , \2680_b1 , \2684_b1 );
not ( \2684_b1 , w_6162 );
and ( \2685_b0 , \2680_b0 , w_6163 );
and ( w_6162 , w_6163 , \2684_b0 );
or ( \2686_b1 , \904_b1 , \912_b1 );
not ( \912_b1 , w_6164 );
and ( \2686_b0 , \904_b0 , w_6165 );
and ( w_6164 , w_6165 , \912_b0 );
or ( \2687_b1 , \841_b1 , \910_b1 );
not ( \910_b1 , w_6166 );
and ( \2687_b0 , \841_b0 , w_6167 );
and ( w_6166 , w_6167 , \910_b0 );
or ( \2688_b1 , \2686_b1 , w_6169 );
not ( w_6169 , w_6170 );
and ( \2688_b0 , \2686_b0 , w_6171 );
and ( w_6170 ,  , w_6171 );
buf ( w_6169 , \2687_b1 );
not ( w_6169 , w_6172 );
not (  , w_6173 );
and ( w_6172 , w_6173 , \2687_b0 );
or ( \2689_b1 , \2688_b1 , w_6174 );
xor ( \2689_b0 , \2688_b0 , w_6176 );
not ( w_6176 , w_6177 );
and ( w_6177 , w_6174 , w_6175 );
buf ( w_6174 , \818_b1 );
not ( w_6174 , w_6178 );
not ( w_6175 , w_6179 );
and ( w_6178 , w_6179 , \818_b0 );
or ( \2690_b1 , \2684_b1 , \2689_b1 );
not ( \2689_b1 , w_6180 );
and ( \2690_b0 , \2684_b0 , w_6181 );
and ( w_6180 , w_6181 , \2689_b0 );
or ( \2691_b1 , \2680_b1 , \2689_b1 );
not ( \2689_b1 , w_6182 );
and ( \2691_b0 , \2680_b0 , w_6183 );
and ( w_6182 , w_6183 , \2689_b0 );
buf ( \2693_b1 , \2371_b1 );
not ( \2693_b1 , w_6184 );
not ( \2693_b0 , w_6185 );
and ( w_6184 , w_6185 , \2371_b0 );
or ( \2694_b1 , \315_b1 , \2550_b1 );
not ( \2550_b1 , w_6186 );
and ( \2694_b0 , \315_b0 , w_6187 );
and ( w_6186 , w_6187 , \2550_b0 );
or ( \2695_b1 , \159_b1 , \2548_b1 );
not ( \2548_b1 , w_6188 );
and ( \2695_b0 , \159_b0 , w_6189 );
and ( w_6188 , w_6189 , \2548_b0 );
or ( \2696_b1 , \2694_b1 , w_6191 );
not ( w_6191 , w_6192 );
and ( \2696_b0 , \2694_b0 , w_6193 );
and ( w_6192 ,  , w_6193 );
buf ( w_6191 , \2695_b1 );
not ( w_6191 , w_6194 );
not (  , w_6195 );
and ( w_6194 , w_6195 , \2695_b0 );
or ( \2697_b1 , \2696_b1 , w_6196 );
xor ( \2697_b0 , \2696_b0 , w_6198 );
not ( w_6198 , w_6199 );
and ( w_6199 , w_6196 , w_6197 );
buf ( w_6196 , \2374_b1 );
not ( w_6196 , w_6200 );
not ( w_6197 , w_6201 );
and ( w_6200 , w_6201 , \2374_b0 );
or ( \2698_b1 , \2693_b1 , \2697_b1 );
not ( \2697_b1 , w_6202 );
and ( \2698_b0 , \2693_b0 , w_6203 );
and ( w_6202 , w_6203 , \2697_b0 );
or ( \2699_b1 , \333_b1 , \2261_b1 );
not ( \2261_b1 , w_6204 );
and ( \2699_b0 , \333_b0 , w_6205 );
and ( w_6204 , w_6205 , \2261_b0 );
or ( \2700_b1 , \305_b1 , \2259_b1 );
not ( \2259_b1 , w_6206 );
and ( \2700_b0 , \305_b0 , w_6207 );
and ( w_6206 , w_6207 , \2259_b0 );
or ( \2701_b1 , \2699_b1 , w_6209 );
not ( w_6209 , w_6210 );
and ( \2701_b0 , \2699_b0 , w_6211 );
and ( w_6210 ,  , w_6211 );
buf ( w_6209 , \2700_b1 );
not ( w_6209 , w_6212 );
not (  , w_6213 );
and ( w_6212 , w_6213 , \2700_b0 );
or ( \2702_b1 , \2701_b1 , w_6214 );
xor ( \2702_b0 , \2701_b0 , w_6216 );
not ( w_6216 , w_6217 );
and ( w_6217 , w_6214 , w_6215 );
buf ( w_6214 , \2124_b1 );
not ( w_6214 , w_6218 );
not ( w_6215 , w_6219 );
and ( w_6218 , w_6219 , \2124_b0 );
or ( \2703_b1 , \2697_b1 , \2702_b1 );
not ( \2702_b1 , w_6220 );
and ( \2703_b0 , \2697_b0 , w_6221 );
and ( w_6220 , w_6221 , \2702_b0 );
or ( \2704_b1 , \2693_b1 , \2702_b1 );
not ( \2702_b1 , w_6222 );
and ( \2704_b0 , \2693_b0 , w_6223 );
and ( w_6222 , w_6223 , \2702_b0 );
or ( \2706_b1 , \2692_b1 , \2705_b1 );
not ( \2705_b1 , w_6224 );
and ( \2706_b0 , \2692_b0 , w_6225 );
and ( w_6224 , w_6225 , \2705_b0 );
or ( \2707_b1 , \353_b1 , \1955_b1 );
not ( \1955_b1 , w_6226 );
and ( \2707_b0 , \353_b0 , w_6227 );
and ( w_6226 , w_6227 , \1955_b0 );
or ( \2708_b1 , \323_b1 , \1953_b1 );
not ( \1953_b1 , w_6228 );
and ( \2708_b0 , \323_b0 , w_6229 );
and ( w_6228 , w_6229 , \1953_b0 );
or ( \2709_b1 , \2707_b1 , w_6231 );
not ( w_6231 , w_6232 );
and ( \2709_b0 , \2707_b0 , w_6233 );
and ( w_6232 ,  , w_6233 );
buf ( w_6231 , \2708_b1 );
not ( w_6231 , w_6234 );
not (  , w_6235 );
and ( w_6234 , w_6235 , \2708_b0 );
or ( \2710_b1 , \2709_b1 , w_6236 );
xor ( \2710_b0 , \2709_b0 , w_6238 );
not ( w_6238 , w_6239 );
and ( w_6239 , w_6236 , w_6237 );
buf ( w_6236 , \1835_b1 );
not ( w_6236 , w_6240 );
not ( w_6237 , w_6241 );
and ( w_6240 , w_6241 , \1835_b0 );
or ( \2711_b1 , \360_b1 , \1742_b1 );
not ( \1742_b1 , w_6242 );
and ( \2711_b0 , \360_b0 , w_6243 );
and ( w_6242 , w_6243 , \1742_b0 );
or ( \2712_b1 , \343_b1 , \1740_b1 );
not ( \1740_b1 , w_6244 );
and ( \2712_b0 , \343_b0 , w_6245 );
and ( w_6244 , w_6245 , \1740_b0 );
or ( \2713_b1 , \2711_b1 , w_6247 );
not ( w_6247 , w_6248 );
and ( \2713_b0 , \2711_b0 , w_6249 );
and ( w_6248 ,  , w_6249 );
buf ( w_6247 , \2712_b1 );
not ( w_6247 , w_6250 );
not (  , w_6251 );
and ( w_6250 , w_6251 , \2712_b0 );
or ( \2714_b1 , \2713_b1 , w_6252 );
xor ( \2714_b0 , \2713_b0 , w_6254 );
not ( w_6254 , w_6255 );
and ( w_6255 , w_6252 , w_6253 );
buf ( w_6252 , \1610_b1 );
not ( w_6252 , w_6256 );
not ( w_6253 , w_6257 );
and ( w_6256 , w_6257 , \1610_b0 );
or ( \2715_b1 , \2710_b1 , \2714_b1 );
not ( \2714_b1 , w_6258 );
and ( \2715_b0 , \2710_b0 , w_6259 );
and ( w_6258 , w_6259 , \2714_b0 );
or ( \2716_b1 , \495_b1 , \1476_b1 );
not ( \1476_b1 , w_6260 );
and ( \2716_b0 , \495_b0 , w_6261 );
and ( w_6260 , w_6261 , \1476_b0 );
or ( \2717_b1 , \444_b1 , \1474_b1 );
not ( \1474_b1 , w_6262 );
and ( \2717_b0 , \444_b0 , w_6263 );
and ( w_6262 , w_6263 , \1474_b0 );
or ( \2718_b1 , \2716_b1 , w_6265 );
not ( w_6265 , w_6266 );
and ( \2718_b0 , \2716_b0 , w_6267 );
and ( w_6266 ,  , w_6267 );
buf ( w_6265 , \2717_b1 );
not ( w_6265 , w_6268 );
not (  , w_6269 );
and ( w_6268 , w_6269 , \2717_b0 );
or ( \2719_b1 , \2718_b1 , w_6270 );
xor ( \2719_b0 , \2718_b0 , w_6272 );
not ( w_6272 , w_6273 );
and ( w_6273 , w_6270 , w_6271 );
buf ( w_6270 , \1363_b1 );
not ( w_6270 , w_6274 );
not ( w_6271 , w_6275 );
and ( w_6274 , w_6275 , \1363_b0 );
or ( \2720_b1 , \2714_b1 , \2719_b1 );
not ( \2719_b1 , w_6276 );
and ( \2720_b0 , \2714_b0 , w_6277 );
and ( w_6276 , w_6277 , \2719_b0 );
or ( \2721_b1 , \2710_b1 , \2719_b1 );
not ( \2719_b1 , w_6278 );
and ( \2721_b0 , \2710_b0 , w_6279 );
and ( w_6278 , w_6279 , \2719_b0 );
or ( \2723_b1 , \2705_b1 , \2722_b1 );
not ( \2722_b1 , w_6280 );
and ( \2723_b0 , \2705_b0 , w_6281 );
and ( w_6280 , w_6281 , \2722_b0 );
or ( \2724_b1 , \2692_b1 , \2722_b1 );
not ( \2722_b1 , w_6282 );
and ( \2724_b0 , \2692_b0 , w_6283 );
and ( w_6282 , w_6283 , \2722_b0 );
or ( \2726_b1 , \1778_b1 , \298_b1 );
not ( \298_b1 , w_6284 );
and ( \2726_b0 , \1778_b0 , w_6285 );
and ( w_6284 , w_6285 , \298_b0 );
or ( \2727_b1 , \1770_b1 , \296_b1 );
not ( \296_b1 , w_6286 );
and ( \2727_b0 , \1770_b0 , w_6287 );
and ( w_6286 , w_6287 , \296_b0 );
or ( \2728_b1 , \2726_b1 , w_6289 );
not ( w_6289 , w_6290 );
and ( \2728_b0 , \2726_b0 , w_6291 );
and ( w_6290 ,  , w_6291 );
buf ( w_6289 , \2727_b1 );
not ( w_6289 , w_6292 );
not (  , w_6293 );
and ( w_6292 , w_6293 , \2727_b0 );
or ( \2729_b1 , \2728_b1 , w_6294 );
xor ( \2729_b0 , \2728_b0 , w_6296 );
not ( w_6296 , w_6297 );
and ( w_6297 , w_6294 , w_6295 );
buf ( w_6294 , \303_b1 );
not ( w_6294 , w_6298 );
not ( w_6295 , w_6299 );
and ( w_6298 , w_6299 , \303_b0 );
or ( \2730_b1 , \2028_b1 , \313_b1 );
not ( \313_b1 , w_6300 );
and ( \2730_b0 , \2028_b0 , w_6301 );
and ( w_6300 , w_6301 , \313_b0 );
or ( \2731_b1 , \2023_b1 , \311_b1 );
not ( \311_b1 , w_6302 );
and ( \2731_b0 , \2023_b0 , w_6303 );
and ( w_6302 , w_6303 , \311_b0 );
or ( \2732_b1 , \2730_b1 , w_6305 );
not ( w_6305 , w_6306 );
and ( \2732_b0 , \2730_b0 , w_6307 );
and ( w_6306 ,  , w_6307 );
buf ( w_6305 , \2731_b1 );
not ( w_6305 , w_6308 );
not (  , w_6309 );
and ( w_6308 , w_6309 , \2731_b0 );
or ( \2733_b1 , \2732_b1 , w_6310 );
xor ( \2733_b0 , \2732_b0 , w_6312 );
not ( w_6312 , w_6313 );
and ( w_6313 , w_6310 , w_6311 );
buf ( w_6310 , \320_b1 );
not ( w_6310 , w_6314 );
not ( w_6311 , w_6315 );
and ( w_6314 , w_6315 , \320_b0 );
or ( \2734_b1 , \2729_b1 , \2733_b1 );
not ( \2733_b1 , w_6316 );
and ( \2734_b0 , \2729_b0 , w_6317 );
and ( w_6316 , w_6317 , \2733_b0 );
or ( \2735_b1 , \2305_b1 , \331_b1 );
not ( \331_b1 , w_6318 );
and ( \2735_b0 , \2305_b0 , w_6319 );
and ( w_6318 , w_6319 , \331_b0 );
or ( \2736_b1 , \2161_b1 , \329_b1 );
not ( \329_b1 , w_6320 );
and ( \2736_b0 , \2161_b0 , w_6321 );
and ( w_6320 , w_6321 , \329_b0 );
or ( \2737_b1 , \2735_b1 , w_6323 );
not ( w_6323 , w_6324 );
and ( \2737_b0 , \2735_b0 , w_6325 );
and ( w_6324 ,  , w_6325 );
buf ( w_6323 , \2736_b1 );
not ( w_6323 , w_6326 );
not (  , w_6327 );
and ( w_6326 , w_6327 , \2736_b0 );
or ( \2738_b1 , \2737_b1 , w_6328 );
xor ( \2738_b0 , \2737_b0 , w_6330 );
not ( w_6330 , w_6331 );
and ( w_6331 , w_6328 , w_6329 );
buf ( w_6328 , \338_b1 );
not ( w_6328 , w_6332 );
not ( w_6329 , w_6333 );
and ( w_6332 , w_6333 , \338_b0 );
or ( \2739_b1 , \2733_b1 , \2738_b1 );
not ( \2738_b1 , w_6334 );
and ( \2739_b0 , \2733_b0 , w_6335 );
and ( w_6334 , w_6335 , \2738_b0 );
or ( \2740_b1 , \2729_b1 , \2738_b1 );
not ( \2738_b1 , w_6336 );
and ( \2740_b0 , \2729_b0 , w_6337 );
and ( w_6336 , w_6337 , \2738_b0 );
or ( \2742_b1 , \1194_b1 , \740_b1 );
not ( \740_b1 , w_6338 );
and ( \2742_b0 , \1194_b0 , w_6339 );
and ( w_6338 , w_6339 , \740_b0 );
or ( \2743_b1 , \1104_b1 , \738_b1 );
not ( \738_b1 , w_6340 );
and ( \2743_b0 , \1104_b0 , w_6341 );
and ( w_6340 , w_6341 , \738_b0 );
or ( \2744_b1 , \2742_b1 , w_6343 );
not ( w_6343 , w_6344 );
and ( \2744_b0 , \2742_b0 , w_6345 );
and ( w_6344 ,  , w_6345 );
buf ( w_6343 , \2743_b1 );
not ( w_6343 , w_6346 );
not (  , w_6347 );
and ( w_6346 , w_6347 , \2743_b0 );
or ( \2745_b1 , \2744_b1 , w_6348 );
xor ( \2745_b0 , \2744_b0 , w_6350 );
not ( w_6350 , w_6351 );
and ( w_6351 , w_6348 , w_6349 );
buf ( w_6348 , \668_b1 );
not ( w_6348 , w_6352 );
not ( w_6349 , w_6353 );
and ( w_6352 , w_6353 , \668_b0 );
or ( \2746_b1 , \1304_b1 , \604_b1 );
not ( \604_b1 , w_6354 );
and ( \2746_b0 , \1304_b0 , w_6355 );
and ( w_6354 , w_6355 , \604_b0 );
or ( \2747_b1 , \1299_b1 , \602_b1 );
not ( \602_b1 , w_6356 );
and ( \2747_b0 , \1299_b0 , w_6357 );
and ( w_6356 , w_6357 , \602_b0 );
or ( \2748_b1 , \2746_b1 , w_6359 );
not ( w_6359 , w_6360 );
and ( \2748_b0 , \2746_b0 , w_6361 );
and ( w_6360 ,  , w_6361 );
buf ( w_6359 , \2747_b1 );
not ( w_6359 , w_6362 );
not (  , w_6363 );
and ( w_6362 , w_6363 , \2747_b0 );
or ( \2749_b1 , \2748_b1 , w_6364 );
xor ( \2749_b0 , \2748_b0 , w_6366 );
not ( w_6366 , w_6367 );
and ( w_6367 , w_6364 , w_6365 );
buf ( w_6364 , \561_b1 );
not ( w_6364 , w_6368 );
not ( w_6365 , w_6369 );
and ( w_6368 , w_6369 , \561_b0 );
or ( \2750_b1 , \2745_b1 , \2749_b1 );
not ( \2749_b1 , w_6370 );
and ( \2750_b0 , \2745_b0 , w_6371 );
and ( w_6370 , w_6371 , \2749_b0 );
or ( \2751_b1 , \1537_b1 , \503_b1 );
not ( \503_b1 , w_6372 );
and ( \2751_b0 , \1537_b0 , w_6373 );
and ( w_6372 , w_6373 , \503_b0 );
or ( \2752_b1 , \1422_b1 , \501_b1 );
not ( \501_b1 , w_6374 );
and ( \2752_b0 , \1422_b0 , w_6375 );
and ( w_6374 , w_6375 , \501_b0 );
or ( \2753_b1 , \2751_b1 , w_6377 );
not ( w_6377 , w_6378 );
and ( \2753_b0 , \2751_b0 , w_6379 );
and ( w_6378 ,  , w_6379 );
buf ( w_6377 , \2752_b1 );
not ( w_6377 , w_6380 );
not (  , w_6381 );
and ( w_6380 , w_6381 , \2752_b0 );
or ( \2754_b1 , \2753_b1 , w_6382 );
xor ( \2754_b0 , \2753_b0 , w_6384 );
not ( w_6384 , w_6385 );
and ( w_6385 , w_6382 , w_6383 );
buf ( w_6382 , \455_b1 );
not ( w_6382 , w_6386 );
not ( w_6383 , w_6387 );
and ( w_6386 , w_6387 , \455_b0 );
or ( \2755_b1 , \2749_b1 , \2754_b1 );
not ( \2754_b1 , w_6388 );
and ( \2755_b0 , \2749_b0 , w_6389 );
and ( w_6388 , w_6389 , \2754_b0 );
or ( \2756_b1 , \2745_b1 , \2754_b1 );
not ( \2754_b1 , w_6390 );
and ( \2756_b0 , \2745_b0 , w_6391 );
and ( w_6390 , w_6391 , \2754_b0 );
or ( \2758_b1 , \2741_b1 , \2757_b1 );
not ( \2757_b1 , w_6392 );
and ( \2758_b0 , \2741_b0 , w_6393 );
and ( w_6392 , w_6393 , \2757_b0 );
or ( \2759_b1 , \2541_b1 , \351_b1 );
not ( \351_b1 , w_6394 );
and ( \2759_b0 , \2541_b0 , w_6395 );
and ( w_6394 , w_6395 , \351_b0 );
or ( \2760_b1 , \2532_b1 , \349_b1 );
not ( \349_b1 , w_6396 );
and ( \2760_b0 , \2532_b0 , w_6397 );
and ( w_6396 , w_6397 , \349_b0 );
or ( \2761_b1 , \2759_b1 , w_6399 );
not ( w_6399 , w_6400 );
and ( \2761_b0 , \2759_b0 , w_6401 );
and ( w_6400 ,  , w_6401 );
buf ( w_6399 , \2760_b1 );
not ( w_6399 , w_6402 );
not (  , w_6403 );
and ( w_6402 , w_6403 , \2760_b0 );
or ( \2762_b1 , \2761_b1 , w_6404 );
xor ( \2762_b0 , \2761_b0 , w_6406 );
not ( w_6406 , w_6407 );
and ( w_6407 , w_6404 , w_6405 );
buf ( w_6404 , \358_b1 );
not ( w_6404 , w_6408 );
not ( w_6405 , w_6409 );
and ( w_6408 , w_6409 , \358_b0 );
buf ( \2763_b1 , RIb4bc018_95_b1 );
buf ( \2763_b0 , RIb4bc018_95_b0 );
or ( \2764_b1 , \2763_b1 , \345_b1 );
not ( \345_b1 , w_6410 );
and ( \2764_b0 , \2763_b0 , w_6411 );
and ( w_6410 , w_6411 , \345_b0 );
or ( \2765_b1 , \2762_b1 , w_6412 );
or ( \2765_b0 , \2762_b0 , \2764_b0 );
not ( \2764_b0 , w_6413 );
and ( w_6413 , w_6412 , \2764_b1 );
or ( \2766_b1 , \2757_b1 , \2765_b1 );
not ( \2765_b1 , w_6414 );
and ( \2766_b0 , \2757_b0 , w_6415 );
and ( w_6414 , w_6415 , \2765_b0 );
or ( \2767_b1 , \2741_b1 , \2765_b1 );
not ( \2765_b1 , w_6416 );
and ( \2767_b0 , \2741_b0 , w_6417 );
and ( w_6416 , w_6417 , \2765_b0 );
or ( \2769_b1 , \2725_b1 , \2768_b1 );
not ( \2768_b1 , w_6418 );
and ( \2769_b0 , \2725_b0 , w_6419 );
and ( w_6418 , w_6419 , \2768_b0 );
or ( \2770_b1 , \2510_b1 , \2514_b1 );
xor ( \2770_b0 , \2510_b0 , w_6420 );
not ( w_6420 , w_6421 );
and ( w_6421 , \2514_b1 , \2514_b0 );
or ( \2771_b1 , \2770_b1 , \2519_b1 );
xor ( \2771_b0 , \2770_b0 , w_6422 );
not ( w_6422 , w_6423 );
and ( w_6423 , \2519_b1 , \2519_b0 );
or ( \2772_b1 , \2526_b1 , \2530_b1 );
xor ( \2772_b0 , \2526_b0 , w_6424 );
not ( w_6424 , w_6425 );
and ( w_6425 , \2530_b1 , \2530_b0 );
or ( \2773_b1 , \2772_b1 , \2536_b1 );
xor ( \2773_b0 , \2772_b0 , w_6426 );
not ( w_6426 , w_6427 );
and ( w_6427 , \2536_b1 , \2536_b0 );
or ( \2774_b1 , \2771_b1 , \2773_b1 );
not ( \2773_b1 , w_6428 );
and ( \2774_b0 , \2771_b0 , w_6429 );
and ( w_6428 , w_6429 , \2773_b0 );
buf ( \2775_b1 , \2542_b1 );
not ( \2775_b1 , w_6430 );
not ( \2775_b0 , w_6431 );
and ( w_6430 , w_6431 , \2542_b0 );
or ( \2776_b1 , \2773_b1 , \2775_b1 );
not ( \2775_b1 , w_6432 );
and ( \2776_b0 , \2773_b0 , w_6433 );
and ( w_6432 , w_6433 , \2775_b0 );
or ( \2777_b1 , \2771_b1 , \2775_b1 );
not ( \2775_b1 , w_6434 );
and ( \2777_b0 , \2771_b0 , w_6435 );
and ( w_6434 , w_6435 , \2775_b0 );
or ( \2779_b1 , \2768_b1 , \2778_b1 );
not ( \2778_b1 , w_6436 );
and ( \2779_b0 , \2768_b0 , w_6437 );
and ( w_6436 , w_6437 , \2778_b0 );
or ( \2780_b1 , \2725_b1 , \2778_b1 );
not ( \2778_b1 , w_6438 );
and ( \2780_b0 , \2725_b0 , w_6439 );
and ( w_6438 , w_6439 , \2778_b0 );
or ( \2782_b1 , \2553_b1 , \2557_b1 );
xor ( \2782_b0 , \2553_b0 , w_6440 );
not ( w_6440 , w_6441 );
and ( w_6441 , \2557_b1 , \2557_b0 );
or ( \2783_b1 , \2782_b1 , \2562_b1 );
xor ( \2783_b0 , \2782_b0 , w_6442 );
not ( w_6442 , w_6443 );
and ( w_6443 , \2562_b1 , \2562_b0 );
or ( \2784_b1 , \2569_b1 , \2573_b1 );
xor ( \2784_b0 , \2569_b0 , w_6444 );
not ( w_6444 , w_6445 );
and ( w_6445 , \2573_b1 , \2573_b0 );
or ( \2785_b1 , \2784_b1 , \2578_b1 );
xor ( \2785_b0 , \2784_b0 , w_6446 );
not ( w_6446 , w_6447 );
and ( w_6447 , \2578_b1 , \2578_b0 );
or ( \2786_b1 , \2783_b1 , \2785_b1 );
not ( \2785_b1 , w_6448 );
and ( \2786_b0 , \2783_b0 , w_6449 );
and ( w_6448 , w_6449 , \2785_b0 );
or ( \2787_b1 , \2586_b1 , \2590_b1 );
xor ( \2787_b0 , \2586_b0 , w_6450 );
not ( w_6450 , w_6451 );
and ( w_6451 , \2590_b1 , \2590_b0 );
or ( \2788_b1 , \2787_b1 , \2595_b1 );
xor ( \2788_b0 , \2787_b0 , w_6452 );
not ( w_6452 , w_6453 );
and ( w_6453 , \2595_b1 , \2595_b0 );
or ( \2789_b1 , \2785_b1 , \2788_b1 );
not ( \2788_b1 , w_6454 );
and ( \2789_b0 , \2785_b0 , w_6455 );
and ( w_6454 , w_6455 , \2788_b0 );
or ( \2790_b1 , \2783_b1 , \2788_b1 );
not ( \2788_b1 , w_6456 );
and ( \2790_b0 , \2783_b0 , w_6457 );
and ( w_6456 , w_6457 , \2788_b0 );
or ( \2792_b1 , \2603_b1 , \2605_b1 );
xor ( \2792_b0 , \2603_b0 , w_6458 );
not ( w_6458 , w_6459 );
and ( w_6459 , \2605_b1 , \2605_b0 );
or ( \2793_b1 , \2792_b1 , \2608_b1 );
xor ( \2793_b0 , \2792_b0 , w_6460 );
not ( w_6460 , w_6461 );
and ( w_6461 , \2608_b1 , \2608_b0 );
or ( \2794_b1 , \2791_b1 , \2793_b1 );
not ( \2793_b1 , w_6462 );
and ( \2794_b0 , \2791_b0 , w_6463 );
and ( w_6462 , w_6463 , \2793_b0 );
or ( \2795_b1 , \2616_b1 , \2618_b1 );
xor ( \2795_b0 , \2616_b0 , w_6464 );
not ( w_6464 , w_6465 );
and ( w_6465 , \2618_b1 , \2618_b0 );
or ( \2796_b1 , \2795_b1 , \2621_b1 );
xor ( \2796_b0 , \2795_b0 , w_6466 );
not ( w_6466 , w_6467 );
and ( w_6467 , \2621_b1 , \2621_b0 );
or ( \2797_b1 , \2793_b1 , \2796_b1 );
not ( \2796_b1 , w_6468 );
and ( \2797_b0 , \2793_b0 , w_6469 );
and ( w_6468 , w_6469 , \2796_b0 );
or ( \2798_b1 , \2791_b1 , \2796_b1 );
not ( \2796_b1 , w_6470 );
and ( \2798_b0 , \2791_b0 , w_6471 );
and ( w_6470 , w_6471 , \2796_b0 );
or ( \2800_b1 , \2781_b1 , \2799_b1 );
not ( \2799_b1 , w_6472 );
and ( \2800_b0 , \2781_b0 , w_6473 );
and ( w_6472 , w_6473 , \2799_b0 );
or ( \2801_b1 , \2635_b1 , \2637_b1 );
xor ( \2801_b0 , \2635_b0 , w_6474 );
not ( w_6474 , w_6475 );
and ( w_6475 , \2637_b1 , \2637_b0 );
or ( \2802_b1 , \2801_b1 , \2639_b1 );
xor ( \2802_b0 , \2801_b0 , w_6476 );
not ( w_6476 , w_6477 );
and ( w_6477 , \2639_b1 , \2639_b0 );
or ( \2803_b1 , \2799_b1 , \2802_b1 );
not ( \2802_b1 , w_6478 );
and ( \2803_b0 , \2799_b0 , w_6479 );
and ( w_6478 , w_6479 , \2802_b0 );
or ( \2804_b1 , \2781_b1 , \2802_b1 );
not ( \2802_b1 , w_6480 );
and ( \2804_b0 , \2781_b0 , w_6481 );
and ( w_6480 , w_6481 , \2802_b0 );
or ( \2806_b1 , \2614_b1 , \2632_b1 );
xor ( \2806_b0 , \2614_b0 , w_6482 );
not ( w_6482 , w_6483 );
and ( w_6483 , \2632_b1 , \2632_b0 );
or ( \2807_b1 , \2806_b1 , \2642_b1 );
xor ( \2807_b0 , \2806_b0 , w_6484 );
not ( w_6484 , w_6485 );
and ( w_6485 , \2642_b1 , \2642_b0 );
or ( \2808_b1 , \2805_b1 , \2807_b1 );
not ( \2807_b1 , w_6486 );
and ( \2808_b0 , \2805_b0 , w_6487 );
and ( w_6486 , w_6487 , \2807_b0 );
or ( \2809_b1 , \2647_b1 , \2649_b1 );
xor ( \2809_b0 , \2647_b0 , w_6488 );
not ( w_6488 , w_6489 );
and ( w_6489 , \2649_b1 , \2649_b0 );
or ( \2810_b1 , \2809_b1 , \2652_b1 );
xor ( \2810_b0 , \2809_b0 , w_6490 );
not ( w_6490 , w_6491 );
and ( w_6491 , \2652_b1 , \2652_b0 );
or ( \2811_b1 , \2807_b1 , \2810_b1 );
not ( \2810_b1 , w_6492 );
and ( \2811_b0 , \2807_b0 , w_6493 );
and ( w_6492 , w_6493 , \2810_b0 );
or ( \2812_b1 , \2805_b1 , \2810_b1 );
not ( \2810_b1 , w_6494 );
and ( \2812_b0 , \2805_b0 , w_6495 );
and ( w_6494 , w_6495 , \2810_b0 );
or ( \2814_b1 , \2645_b1 , \2655_b1 );
xor ( \2814_b0 , \2645_b0 , w_6496 );
not ( w_6496 , w_6497 );
and ( w_6497 , \2655_b1 , \2655_b0 );
or ( \2815_b1 , \2814_b1 , \2658_b1 );
xor ( \2815_b0 , \2814_b0 , w_6498 );
not ( w_6498 , w_6499 );
and ( w_6499 , \2658_b1 , \2658_b0 );
or ( \2816_b1 , \2813_b1 , \2815_b1 );
not ( \2815_b1 , w_6500 );
and ( \2816_b0 , \2813_b0 , w_6501 );
and ( w_6500 , w_6501 , \2815_b0 );
or ( \2817_b1 , \2663_b1 , \2665_b1 );
xor ( \2817_b0 , \2663_b0 , w_6502 );
not ( w_6502 , w_6503 );
and ( w_6503 , \2665_b1 , \2665_b0 );
or ( \2818_b1 , \2815_b1 , \2817_b1 );
not ( \2817_b1 , w_6504 );
and ( \2818_b0 , \2815_b0 , w_6505 );
and ( w_6504 , w_6505 , \2817_b0 );
or ( \2819_b1 , \2813_b1 , \2817_b1 );
not ( \2817_b1 , w_6506 );
and ( \2819_b0 , \2813_b0 , w_6507 );
and ( w_6506 , w_6507 , \2817_b0 );
or ( \2821_b1 , \2676_b1 , \2820_b1 );
not ( \2820_b1 , w_6508 );
and ( \2821_b0 , \2676_b0 , w_6509 );
and ( w_6508 , w_6509 , \2820_b0 );
or ( \2822_b1 , \2676_b1 , \2820_b1 );
xor ( \2822_b0 , \2676_b0 , w_6510 );
not ( w_6510 , w_6511 );
and ( w_6511 , \2820_b1 , \2820_b0 );
or ( \2823_b1 , \2813_b1 , \2815_b1 );
xor ( \2823_b0 , \2813_b0 , w_6512 );
not ( w_6512 , w_6513 );
and ( w_6513 , \2815_b1 , \2815_b0 );
or ( \2824_b1 , \2823_b1 , \2817_b1 );
xor ( \2824_b0 , \2823_b0 , w_6514 );
not ( w_6514 , w_6515 );
and ( w_6515 , \2817_b1 , \2817_b0 );
or ( \2825_b1 , \1770_b1 , \503_b1 );
not ( \503_b1 , w_6516 );
and ( \2825_b0 , \1770_b0 , w_6517 );
and ( w_6516 , w_6517 , \503_b0 );
or ( \2826_b1 , \1537_b1 , \501_b1 );
not ( \501_b1 , w_6518 );
and ( \2826_b0 , \1537_b0 , w_6519 );
and ( w_6518 , w_6519 , \501_b0 );
or ( \2827_b1 , \2825_b1 , w_6521 );
not ( w_6521 , w_6522 );
and ( \2827_b0 , \2825_b0 , w_6523 );
and ( w_6522 ,  , w_6523 );
buf ( w_6521 , \2826_b1 );
not ( w_6521 , w_6524 );
not (  , w_6525 );
and ( w_6524 , w_6525 , \2826_b0 );
or ( \2828_b1 , \2827_b1 , w_6526 );
xor ( \2828_b0 , \2827_b0 , w_6528 );
not ( w_6528 , w_6529 );
and ( w_6529 , w_6526 , w_6527 );
buf ( w_6526 , \455_b1 );
not ( w_6526 , w_6530 );
not ( w_6527 , w_6531 );
and ( w_6530 , w_6531 , \455_b0 );
or ( \2829_b1 , \2023_b1 , \298_b1 );
not ( \298_b1 , w_6532 );
and ( \2829_b0 , \2023_b0 , w_6533 );
and ( w_6532 , w_6533 , \298_b0 );
or ( \2830_b1 , \1778_b1 , \296_b1 );
not ( \296_b1 , w_6534 );
and ( \2830_b0 , \1778_b0 , w_6535 );
and ( w_6534 , w_6535 , \296_b0 );
or ( \2831_b1 , \2829_b1 , w_6537 );
not ( w_6537 , w_6538 );
and ( \2831_b0 , \2829_b0 , w_6539 );
and ( w_6538 ,  , w_6539 );
buf ( w_6537 , \2830_b1 );
not ( w_6537 , w_6540 );
not (  , w_6541 );
and ( w_6540 , w_6541 , \2830_b0 );
or ( \2832_b1 , \2831_b1 , w_6542 );
xor ( \2832_b0 , \2831_b0 , w_6544 );
not ( w_6544 , w_6545 );
and ( w_6545 , w_6542 , w_6543 );
buf ( w_6542 , \303_b1 );
not ( w_6542 , w_6546 );
not ( w_6543 , w_6547 );
and ( w_6546 , w_6547 , \303_b0 );
or ( \2833_b1 , \2828_b1 , \2832_b1 );
not ( \2832_b1 , w_6548 );
and ( \2833_b0 , \2828_b0 , w_6549 );
and ( w_6548 , w_6549 , \2832_b0 );
or ( \2834_b1 , \2161_b1 , \313_b1 );
not ( \313_b1 , w_6550 );
and ( \2834_b0 , \2161_b0 , w_6551 );
and ( w_6550 , w_6551 , \313_b0 );
or ( \2835_b1 , \2028_b1 , \311_b1 );
not ( \311_b1 , w_6552 );
and ( \2835_b0 , \2028_b0 , w_6553 );
and ( w_6552 , w_6553 , \311_b0 );
or ( \2836_b1 , \2834_b1 , w_6555 );
not ( w_6555 , w_6556 );
and ( \2836_b0 , \2834_b0 , w_6557 );
and ( w_6556 ,  , w_6557 );
buf ( w_6555 , \2835_b1 );
not ( w_6555 , w_6558 );
not (  , w_6559 );
and ( w_6558 , w_6559 , \2835_b0 );
or ( \2837_b1 , \2836_b1 , w_6560 );
xor ( \2837_b0 , \2836_b0 , w_6562 );
not ( w_6562 , w_6563 );
and ( w_6563 , w_6560 , w_6561 );
buf ( w_6560 , \320_b1 );
not ( w_6560 , w_6564 );
not ( w_6561 , w_6565 );
and ( w_6564 , w_6565 , \320_b0 );
or ( \2838_b1 , \2832_b1 , \2837_b1 );
not ( \2837_b1 , w_6566 );
and ( \2838_b0 , \2832_b0 , w_6567 );
and ( w_6566 , w_6567 , \2837_b0 );
or ( \2839_b1 , \2828_b1 , \2837_b1 );
not ( \2837_b1 , w_6568 );
and ( \2839_b0 , \2828_b0 , w_6569 );
and ( w_6568 , w_6569 , \2837_b0 );
or ( \2841_b1 , \2532_b1 , \331_b1 );
not ( \331_b1 , w_6570 );
and ( \2841_b0 , \2532_b0 , w_6571 );
and ( w_6570 , w_6571 , \331_b0 );
or ( \2842_b1 , \2305_b1 , \329_b1 );
not ( \329_b1 , w_6572 );
and ( \2842_b0 , \2305_b0 , w_6573 );
and ( w_6572 , w_6573 , \329_b0 );
or ( \2843_b1 , \2841_b1 , w_6575 );
not ( w_6575 , w_6576 );
and ( \2843_b0 , \2841_b0 , w_6577 );
and ( w_6576 ,  , w_6577 );
buf ( w_6575 , \2842_b1 );
not ( w_6575 , w_6578 );
not (  , w_6579 );
and ( w_6578 , w_6579 , \2842_b0 );
or ( \2844_b1 , \2843_b1 , w_6580 );
xor ( \2844_b0 , \2843_b0 , w_6582 );
not ( w_6582 , w_6583 );
and ( w_6583 , w_6580 , w_6581 );
buf ( w_6580 , \338_b1 );
not ( w_6580 , w_6584 );
not ( w_6581 , w_6585 );
and ( w_6584 , w_6585 , \338_b0 );
or ( \2845_b1 , \2763_b1 , \351_b1 );
not ( \351_b1 , w_6586 );
and ( \2845_b0 , \2763_b0 , w_6587 );
and ( w_6586 , w_6587 , \351_b0 );
or ( \2846_b1 , \2541_b1 , \349_b1 );
not ( \349_b1 , w_6588 );
and ( \2846_b0 , \2541_b0 , w_6589 );
and ( w_6588 , w_6589 , \349_b0 );
or ( \2847_b1 , \2845_b1 , w_6591 );
not ( w_6591 , w_6592 );
and ( \2847_b0 , \2845_b0 , w_6593 );
and ( w_6592 ,  , w_6593 );
buf ( w_6591 , \2846_b1 );
not ( w_6591 , w_6594 );
not (  , w_6595 );
and ( w_6594 , w_6595 , \2846_b0 );
or ( \2848_b1 , \2847_b1 , w_6596 );
xor ( \2848_b0 , \2847_b0 , w_6598 );
not ( w_6598 , w_6599 );
and ( w_6599 , w_6596 , w_6597 );
buf ( w_6596 , \358_b1 );
not ( w_6596 , w_6600 );
not ( w_6597 , w_6601 );
and ( w_6600 , w_6601 , \358_b0 );
or ( \2849_b1 , \2844_b1 , \2848_b1 );
not ( \2848_b1 , w_6602 );
and ( \2849_b0 , \2844_b0 , w_6603 );
and ( w_6602 , w_6603 , \2848_b0 );
buf ( \2850_b1 , RIb4bbfa0_96_b1 );
buf ( \2850_b0 , RIb4bbfa0_96_b0 );
or ( \2851_b1 , \2850_b1 , w_6605 );
not ( w_6605 , w_6606 );
and ( \2851_b0 , \2850_b0 , w_6607 );
and ( w_6606 ,  , w_6607 );
buf ( w_6605 , \345_b1 );
not ( w_6605 , w_6608 );
not (  , w_6609 );
and ( w_6608 , w_6609 , \345_b0 );
buf ( \2852_b1 , \2851_b1 );
not ( \2852_b1 , w_6610 );
not ( \2852_b0 , w_6611 );
and ( w_6610 , w_6611 , \2851_b0 );
or ( \2853_b1 , \2848_b1 , \2852_b1 );
not ( \2852_b1 , w_6612 );
and ( \2853_b0 , \2848_b0 , w_6613 );
and ( w_6612 , w_6613 , \2852_b0 );
or ( \2854_b1 , \2844_b1 , \2852_b1 );
not ( \2852_b1 , w_6614 );
and ( \2854_b0 , \2844_b0 , w_6615 );
and ( w_6614 , w_6615 , \2852_b0 );
or ( \2856_b1 , \2840_b1 , \2855_b1 );
not ( \2855_b1 , w_6616 );
and ( \2856_b0 , \2840_b0 , w_6617 );
and ( w_6616 , w_6617 , \2855_b0 );
or ( \2857_b1 , \1104_b1 , \912_b1 );
not ( \912_b1 , w_6618 );
and ( \2857_b0 , \1104_b0 , w_6619 );
and ( w_6618 , w_6619 , \912_b0 );
or ( \2858_b1 , \904_b1 , \910_b1 );
not ( \910_b1 , w_6620 );
and ( \2858_b0 , \904_b0 , w_6621 );
and ( w_6620 , w_6621 , \910_b0 );
or ( \2859_b1 , \2857_b1 , w_6623 );
not ( w_6623 , w_6624 );
and ( \2859_b0 , \2857_b0 , w_6625 );
and ( w_6624 ,  , w_6625 );
buf ( w_6623 , \2858_b1 );
not ( w_6623 , w_6626 );
not (  , w_6627 );
and ( w_6626 , w_6627 , \2858_b0 );
or ( \2860_b1 , \2859_b1 , w_6628 );
xor ( \2860_b0 , \2859_b0 , w_6630 );
not ( w_6630 , w_6631 );
and ( w_6631 , w_6628 , w_6629 );
buf ( w_6628 , \818_b1 );
not ( w_6628 , w_6632 );
not ( w_6629 , w_6633 );
and ( w_6632 , w_6633 , \818_b0 );
or ( \2861_b1 , \1299_b1 , \740_b1 );
not ( \740_b1 , w_6634 );
and ( \2861_b0 , \1299_b0 , w_6635 );
and ( w_6634 , w_6635 , \740_b0 );
or ( \2862_b1 , \1194_b1 , \738_b1 );
not ( \738_b1 , w_6636 );
and ( \2862_b0 , \1194_b0 , w_6637 );
and ( w_6636 , w_6637 , \738_b0 );
or ( \2863_b1 , \2861_b1 , w_6639 );
not ( w_6639 , w_6640 );
and ( \2863_b0 , \2861_b0 , w_6641 );
and ( w_6640 ,  , w_6641 );
buf ( w_6639 , \2862_b1 );
not ( w_6639 , w_6642 );
not (  , w_6643 );
and ( w_6642 , w_6643 , \2862_b0 );
or ( \2864_b1 , \2863_b1 , w_6644 );
xor ( \2864_b0 , \2863_b0 , w_6646 );
not ( w_6646 , w_6647 );
and ( w_6647 , w_6644 , w_6645 );
buf ( w_6644 , \668_b1 );
not ( w_6644 , w_6648 );
not ( w_6645 , w_6649 );
and ( w_6648 , w_6649 , \668_b0 );
or ( \2865_b1 , \2860_b1 , \2864_b1 );
not ( \2864_b1 , w_6650 );
and ( \2865_b0 , \2860_b0 , w_6651 );
and ( w_6650 , w_6651 , \2864_b0 );
or ( \2866_b1 , \1422_b1 , \604_b1 );
not ( \604_b1 , w_6652 );
and ( \2866_b0 , \1422_b0 , w_6653 );
and ( w_6652 , w_6653 , \604_b0 );
or ( \2867_b1 , \1304_b1 , \602_b1 );
not ( \602_b1 , w_6654 );
and ( \2867_b0 , \1304_b0 , w_6655 );
and ( w_6654 , w_6655 , \602_b0 );
or ( \2868_b1 , \2866_b1 , w_6657 );
not ( w_6657 , w_6658 );
and ( \2868_b0 , \2866_b0 , w_6659 );
and ( w_6658 ,  , w_6659 );
buf ( w_6657 , \2867_b1 );
not ( w_6657 , w_6660 );
not (  , w_6661 );
and ( w_6660 , w_6661 , \2867_b0 );
or ( \2869_b1 , \2868_b1 , w_6662 );
xor ( \2869_b0 , \2868_b0 , w_6664 );
not ( w_6664 , w_6665 );
and ( w_6665 , w_6662 , w_6663 );
buf ( w_6662 , \561_b1 );
not ( w_6662 , w_6666 );
not ( w_6663 , w_6667 );
and ( w_6666 , w_6667 , \561_b0 );
or ( \2870_b1 , \2864_b1 , \2869_b1 );
not ( \2869_b1 , w_6668 );
and ( \2870_b0 , \2864_b0 , w_6669 );
and ( w_6668 , w_6669 , \2869_b0 );
or ( \2871_b1 , \2860_b1 , \2869_b1 );
not ( \2869_b1 , w_6670 );
and ( \2871_b0 , \2860_b0 , w_6671 );
and ( w_6670 , w_6671 , \2869_b0 );
or ( \2873_b1 , \2855_b1 , \2872_b1 );
not ( \2872_b1 , w_6672 );
and ( \2873_b0 , \2855_b0 , w_6673 );
and ( w_6672 , w_6673 , \2872_b0 );
or ( \2874_b1 , \2840_b1 , \2872_b1 );
not ( \2872_b1 , w_6674 );
and ( \2874_b0 , \2840_b0 , w_6675 );
and ( w_6674 , w_6675 , \2872_b0 );
or ( \2876_b1 , \593_b1 , \1476_b1 );
not ( \1476_b1 , w_6676 );
and ( \2876_b0 , \593_b0 , w_6677 );
and ( w_6676 , w_6677 , \1476_b0 );
or ( \2877_b1 , \495_b1 , \1474_b1 );
not ( \1474_b1 , w_6678 );
and ( \2877_b0 , \495_b0 , w_6679 );
and ( w_6678 , w_6679 , \1474_b0 );
or ( \2878_b1 , \2876_b1 , w_6681 );
not ( w_6681 , w_6682 );
and ( \2878_b0 , \2876_b0 , w_6683 );
and ( w_6682 ,  , w_6683 );
buf ( w_6681 , \2877_b1 );
not ( w_6681 , w_6684 );
not (  , w_6685 );
and ( w_6684 , w_6685 , \2877_b0 );
or ( \2879_b1 , \2878_b1 , w_6686 );
xor ( \2879_b0 , \2878_b0 , w_6688 );
not ( w_6688 , w_6689 );
and ( w_6689 , w_6686 , w_6687 );
buf ( w_6686 , \1363_b1 );
not ( w_6686 , w_6690 );
not ( w_6687 , w_6691 );
and ( w_6690 , w_6691 , \1363_b0 );
or ( \2880_b1 , \703_b1 , \1280_b1 );
not ( \1280_b1 , w_6692 );
and ( \2880_b0 , \703_b0 , w_6693 );
and ( w_6692 , w_6693 , \1280_b0 );
or ( \2881_b1 , \621_b1 , \1278_b1 );
not ( \1278_b1 , w_6694 );
and ( \2881_b0 , \621_b0 , w_6695 );
and ( w_6694 , w_6695 , \1278_b0 );
or ( \2882_b1 , \2880_b1 , w_6697 );
not ( w_6697 , w_6698 );
and ( \2882_b0 , \2880_b0 , w_6699 );
and ( w_6698 ,  , w_6699 );
buf ( w_6697 , \2881_b1 );
not ( w_6697 , w_6700 );
not (  , w_6701 );
and ( w_6700 , w_6701 , \2881_b0 );
or ( \2883_b1 , \2882_b1 , w_6702 );
xor ( \2883_b0 , \2882_b0 , w_6704 );
not ( w_6704 , w_6705 );
and ( w_6705 , w_6702 , w_6703 );
buf ( w_6702 , \1177_b1 );
not ( w_6702 , w_6706 );
not ( w_6703 , w_6707 );
and ( w_6706 , w_6707 , \1177_b0 );
or ( \2884_b1 , \2879_b1 , \2883_b1 );
not ( \2883_b1 , w_6708 );
and ( \2884_b0 , \2879_b0 , w_6709 );
and ( w_6708 , w_6709 , \2883_b0 );
or ( \2885_b1 , \841_b1 , \1062_b1 );
not ( \1062_b1 , w_6710 );
and ( \2885_b0 , \841_b0 , w_6711 );
and ( w_6710 , w_6711 , \1062_b0 );
or ( \2886_b1 , \777_b1 , \1060_b1 );
not ( \1060_b1 , w_6712 );
and ( \2886_b0 , \777_b0 , w_6713 );
and ( w_6712 , w_6713 , \1060_b0 );
or ( \2887_b1 , \2885_b1 , w_6715 );
not ( w_6715 , w_6716 );
and ( \2887_b0 , \2885_b0 , w_6717 );
and ( w_6716 ,  , w_6717 );
buf ( w_6715 , \2886_b1 );
not ( w_6715 , w_6718 );
not (  , w_6719 );
and ( w_6718 , w_6719 , \2886_b0 );
or ( \2888_b1 , \2887_b1 , w_6720 );
xor ( \2888_b0 , \2887_b0 , w_6722 );
not ( w_6722 , w_6723 );
and ( w_6723 , w_6720 , w_6721 );
buf ( w_6720 , \984_b1 );
not ( w_6720 , w_6724 );
not ( w_6721 , w_6725 );
and ( w_6724 , w_6725 , \984_b0 );
or ( \2889_b1 , \2883_b1 , \2888_b1 );
not ( \2888_b1 , w_6726 );
and ( \2889_b0 , \2883_b0 , w_6727 );
and ( w_6726 , w_6727 , \2888_b0 );
or ( \2890_b1 , \2879_b1 , \2888_b1 );
not ( \2888_b1 , w_6728 );
and ( \2890_b0 , \2879_b0 , w_6729 );
and ( w_6728 , w_6729 , \2888_b0 );
or ( \2892_b1 , \323_b1 , \2261_b1 );
not ( \2261_b1 , w_6730 );
and ( \2892_b0 , \323_b0 , w_6731 );
and ( w_6730 , w_6731 , \2261_b0 );
or ( \2893_b1 , \333_b1 , \2259_b1 );
not ( \2259_b1 , w_6732 );
and ( \2893_b0 , \333_b0 , w_6733 );
and ( w_6732 , w_6733 , \2259_b0 );
or ( \2894_b1 , \2892_b1 , w_6735 );
not ( w_6735 , w_6736 );
and ( \2894_b0 , \2892_b0 , w_6737 );
and ( w_6736 ,  , w_6737 );
buf ( w_6735 , \2893_b1 );
not ( w_6735 , w_6738 );
not (  , w_6739 );
and ( w_6738 , w_6739 , \2893_b0 );
or ( \2895_b1 , \2894_b1 , w_6740 );
xor ( \2895_b0 , \2894_b0 , w_6742 );
not ( w_6742 , w_6743 );
and ( w_6743 , w_6740 , w_6741 );
buf ( w_6740 , \2124_b1 );
not ( w_6740 , w_6744 );
not ( w_6741 , w_6745 );
and ( w_6744 , w_6745 , \2124_b0 );
or ( \2896_b1 , \343_b1 , \1955_b1 );
not ( \1955_b1 , w_6746 );
and ( \2896_b0 , \343_b0 , w_6747 );
and ( w_6746 , w_6747 , \1955_b0 );
or ( \2897_b1 , \353_b1 , \1953_b1 );
not ( \1953_b1 , w_6748 );
and ( \2897_b0 , \353_b0 , w_6749 );
and ( w_6748 , w_6749 , \1953_b0 );
or ( \2898_b1 , \2896_b1 , w_6751 );
not ( w_6751 , w_6752 );
and ( \2898_b0 , \2896_b0 , w_6753 );
and ( w_6752 ,  , w_6753 );
buf ( w_6751 , \2897_b1 );
not ( w_6751 , w_6754 );
not (  , w_6755 );
and ( w_6754 , w_6755 , \2897_b0 );
or ( \2899_b1 , \2898_b1 , w_6756 );
xor ( \2899_b0 , \2898_b0 , w_6758 );
not ( w_6758 , w_6759 );
and ( w_6759 , w_6756 , w_6757 );
buf ( w_6756 , \1835_b1 );
not ( w_6756 , w_6760 );
not ( w_6757 , w_6761 );
and ( w_6760 , w_6761 , \1835_b0 );
or ( \2900_b1 , \2895_b1 , \2899_b1 );
not ( \2899_b1 , w_6762 );
and ( \2900_b0 , \2895_b0 , w_6763 );
and ( w_6762 , w_6763 , \2899_b0 );
or ( \2901_b1 , \444_b1 , \1742_b1 );
not ( \1742_b1 , w_6764 );
and ( \2901_b0 , \444_b0 , w_6765 );
and ( w_6764 , w_6765 , \1742_b0 );
or ( \2902_b1 , \360_b1 , \1740_b1 );
not ( \1740_b1 , w_6766 );
and ( \2902_b0 , \360_b0 , w_6767 );
and ( w_6766 , w_6767 , \1740_b0 );
or ( \2903_b1 , \2901_b1 , w_6769 );
not ( w_6769 , w_6770 );
and ( \2903_b0 , \2901_b0 , w_6771 );
and ( w_6770 ,  , w_6771 );
buf ( w_6769 , \2902_b1 );
not ( w_6769 , w_6772 );
not (  , w_6773 );
and ( w_6772 , w_6773 , \2902_b0 );
or ( \2904_b1 , \2903_b1 , w_6774 );
xor ( \2904_b0 , \2903_b0 , w_6776 );
not ( w_6776 , w_6777 );
and ( w_6777 , w_6774 , w_6775 );
buf ( w_6774 , \1610_b1 );
not ( w_6774 , w_6778 );
not ( w_6775 , w_6779 );
and ( w_6778 , w_6779 , \1610_b0 );
or ( \2905_b1 , \2899_b1 , \2904_b1 );
not ( \2904_b1 , w_6780 );
and ( \2905_b0 , \2899_b0 , w_6781 );
and ( w_6780 , w_6781 , \2904_b0 );
or ( \2906_b1 , \2895_b1 , \2904_b1 );
not ( \2904_b1 , w_6782 );
and ( \2906_b0 , \2895_b0 , w_6783 );
and ( w_6782 , w_6783 , \2904_b0 );
or ( \2908_b1 , \2891_b1 , \2907_b1 );
not ( \2907_b1 , w_6784 );
and ( \2908_b0 , \2891_b0 , w_6785 );
and ( w_6784 , w_6785 , \2907_b0 );
and ( \2909_nR123_b0 , RIb4bfab0_64_b0 , w_6786 );
and ( \2909_nR123_b0 , 1'b0_b0 , w_6787 );
and ( w_6800 , w_6801 , w_6788 );
and ( w_6788 , 1'b0_b0 , w_6789 );
and ( w_6801 , 1'b0_b1 , w_6790 );
and ( \2909_nR123_b1 , RIb4bfab0_64_b0 , w_6791 );
and ( RIb4bfab0_64_b1 , w_6802 , w_6792 );
and ( w_6801 , 1'b0_b0 , w_6793 );
and ( \2909_nR123_b1 , \2909_nR123_b0 , w_6794 );
and ( w_6799 , w_6803 , \287_b1 );
or ( w_6786 , w_6787 , w_6795 );
or ( w_6795 , w_6789 , \287_b0 );
or ( w_6790 , w_6791 , w_6796 );
or ( w_6796 , w_6792 , w_6797 );
or ( w_6797 , w_6793 , w_6798 );
or ( w_6798 , w_6794 , w_6799 );
not ( RIb4bfab0_64_b1 , w_6800 );
not ( RIb4bfab0_64_b0 , w_6801 );
not ( \2909_nR123_b1 , w_6802 );
not ( \287_b0 , w_6803 );
buf ( \2910_b1 , \2909_nR123_b1 );
buf ( \2910_b0 , \2909_nR123_b0 );
or ( \2911_b1 , \2371_b1 , \2910_b1 );
xor ( \2911_b0 , \2371_b0 , w_6804 );
not ( w_6804 , w_6805 );
and ( w_6805 , \2910_b1 , \2910_b0 );
buf ( \2912_b1 , \2910_b1 );
not ( \2912_b1 , w_6806 );
not ( \2912_b0 , w_6807 );
and ( w_6806 , w_6807 , \2910_b0 );
or ( \2913_b1 , \2911_b1 , \2912_b1 );
not ( \2912_b1 , w_6808 );
and ( \2913_b0 , \2911_b0 , w_6809 );
and ( w_6808 , w_6809 , \2912_b0 );
or ( \2914_b1 , \159_b1 , \2913_b1 );
not ( \2913_b1 , w_6810 );
and ( \2914_b0 , \159_b0 , w_6811 );
and ( w_6810 , w_6811 , \2913_b0 );
buf ( \2915_b1 , \2914_b1 );
not ( \2915_b1 , w_6812 );
not ( \2915_b0 , w_6813 );
and ( w_6812 , w_6813 , \2914_b0 );
or ( \2916_b1 , \2915_b1 , w_6814 );
xor ( \2916_b0 , \2915_b0 , w_6816 );
not ( w_6816 , w_6817 );
and ( w_6817 , w_6814 , w_6815 );
buf ( w_6814 , \2371_b1 );
not ( w_6814 , w_6818 );
not ( w_6815 , w_6819 );
and ( w_6818 , w_6819 , \2371_b0 );
or ( \2917_b1 , \305_b1 , \2550_b1 );
not ( \2550_b1 , w_6820 );
and ( \2917_b0 , \305_b0 , w_6821 );
and ( w_6820 , w_6821 , \2550_b0 );
or ( \2918_b1 , \315_b1 , \2548_b1 );
not ( \2548_b1 , w_6822 );
and ( \2918_b0 , \315_b0 , w_6823 );
and ( w_6822 , w_6823 , \2548_b0 );
or ( \2919_b1 , \2917_b1 , w_6825 );
not ( w_6825 , w_6826 );
and ( \2919_b0 , \2917_b0 , w_6827 );
and ( w_6826 ,  , w_6827 );
buf ( w_6825 , \2918_b1 );
not ( w_6825 , w_6828 );
not (  , w_6829 );
and ( w_6828 , w_6829 , \2918_b0 );
or ( \2920_b1 , \2919_b1 , w_6830 );
xor ( \2920_b0 , \2919_b0 , w_6832 );
not ( w_6832 , w_6833 );
and ( w_6833 , w_6830 , w_6831 );
buf ( w_6830 , \2374_b1 );
not ( w_6830 , w_6834 );
not ( w_6831 , w_6835 );
and ( w_6834 , w_6835 , \2374_b0 );
or ( \2921_b1 , \2916_b1 , \2920_b1 );
not ( \2920_b1 , w_6836 );
and ( \2921_b0 , \2916_b0 , w_6837 );
and ( w_6836 , w_6837 , \2920_b0 );
or ( \2922_b1 , \2907_b1 , \2921_b1 );
not ( \2921_b1 , w_6838 );
and ( \2922_b0 , \2907_b0 , w_6839 );
and ( w_6838 , w_6839 , \2921_b0 );
or ( \2923_b1 , \2891_b1 , \2921_b1 );
not ( \2921_b1 , w_6840 );
and ( \2923_b0 , \2891_b0 , w_6841 );
and ( w_6840 , w_6841 , \2921_b0 );
or ( \2925_b1 , \2875_b1 , \2924_b1 );
not ( \2924_b1 , w_6842 );
and ( \2925_b0 , \2875_b0 , w_6843 );
and ( w_6842 , w_6843 , \2924_b0 );
or ( \2926_b1 , \2729_b1 , \2733_b1 );
xor ( \2926_b0 , \2729_b0 , w_6844 );
not ( w_6844 , w_6845 );
and ( w_6845 , \2733_b1 , \2733_b0 );
or ( \2927_b1 , \2926_b1 , \2738_b1 );
xor ( \2927_b0 , \2926_b0 , w_6846 );
not ( w_6846 , w_6847 );
and ( w_6847 , \2738_b1 , \2738_b0 );
or ( \2928_b1 , \2745_b1 , \2749_b1 );
xor ( \2928_b0 , \2745_b0 , w_6848 );
not ( w_6848 , w_6849 );
and ( w_6849 , \2749_b1 , \2749_b0 );
or ( \2929_b1 , \2928_b1 , \2754_b1 );
xor ( \2929_b0 , \2928_b0 , w_6850 );
not ( w_6850 , w_6851 );
and ( w_6851 , \2754_b1 , \2754_b0 );
or ( \2930_b1 , \2927_b1 , \2929_b1 );
not ( \2929_b1 , w_6852 );
and ( \2930_b0 , \2927_b0 , w_6853 );
and ( w_6852 , w_6853 , \2929_b0 );
or ( \2931_b1 , \2762_b1 , w_6854 );
xor ( \2931_b0 , \2762_b0 , w_6856 );
not ( w_6856 , w_6857 );
and ( w_6857 , w_6854 , w_6855 );
buf ( w_6854 , \2764_b1 );
not ( w_6854 , w_6858 );
not ( w_6855 , w_6859 );
and ( w_6858 , w_6859 , \2764_b0 );
or ( \2932_b1 , \2929_b1 , \2931_b1 );
not ( \2931_b1 , w_6860 );
and ( \2932_b0 , \2929_b0 , w_6861 );
and ( w_6860 , w_6861 , \2931_b0 );
or ( \2933_b1 , \2927_b1 , \2931_b1 );
not ( \2931_b1 , w_6862 );
and ( \2933_b0 , \2927_b0 , w_6863 );
and ( w_6862 , w_6863 , \2931_b0 );
or ( \2935_b1 , \2924_b1 , \2934_b1 );
not ( \2934_b1 , w_6864 );
and ( \2935_b0 , \2924_b0 , w_6865 );
and ( w_6864 , w_6865 , \2934_b0 );
or ( \2936_b1 , \2875_b1 , \2934_b1 );
not ( \2934_b1 , w_6866 );
and ( \2936_b0 , \2875_b0 , w_6867 );
and ( w_6866 , w_6867 , \2934_b0 );
or ( \2938_b1 , \2680_b1 , \2684_b1 );
xor ( \2938_b0 , \2680_b0 , w_6868 );
not ( w_6868 , w_6869 );
and ( w_6869 , \2684_b1 , \2684_b0 );
or ( \2939_b1 , \2938_b1 , \2689_b1 );
xor ( \2939_b0 , \2938_b0 , w_6870 );
not ( w_6870 , w_6871 );
and ( w_6871 , \2689_b1 , \2689_b0 );
or ( \2940_b1 , \2693_b1 , \2697_b1 );
xor ( \2940_b0 , \2693_b0 , w_6872 );
not ( w_6872 , w_6873 );
and ( w_6873 , \2697_b1 , \2697_b0 );
or ( \2941_b1 , \2940_b1 , \2702_b1 );
xor ( \2941_b0 , \2940_b0 , w_6874 );
not ( w_6874 , w_6875 );
and ( w_6875 , \2702_b1 , \2702_b0 );
or ( \2942_b1 , \2939_b1 , \2941_b1 );
not ( \2941_b1 , w_6876 );
and ( \2942_b0 , \2939_b0 , w_6877 );
and ( w_6876 , w_6877 , \2941_b0 );
or ( \2943_b1 , \2710_b1 , \2714_b1 );
xor ( \2943_b0 , \2710_b0 , w_6878 );
not ( w_6878 , w_6879 );
and ( w_6879 , \2714_b1 , \2714_b0 );
or ( \2944_b1 , \2943_b1 , \2719_b1 );
xor ( \2944_b0 , \2943_b0 , w_6880 );
not ( w_6880 , w_6881 );
and ( w_6881 , \2719_b1 , \2719_b0 );
or ( \2945_b1 , \2941_b1 , \2944_b1 );
not ( \2944_b1 , w_6882 );
and ( \2945_b0 , \2941_b0 , w_6883 );
and ( w_6882 , w_6883 , \2944_b0 );
or ( \2946_b1 , \2939_b1 , \2944_b1 );
not ( \2944_b1 , w_6884 );
and ( \2946_b0 , \2939_b0 , w_6885 );
and ( w_6884 , w_6885 , \2944_b0 );
or ( \2948_b1 , \2783_b1 , \2785_b1 );
xor ( \2948_b0 , \2783_b0 , w_6886 );
not ( w_6886 , w_6887 );
and ( w_6887 , \2785_b1 , \2785_b0 );
or ( \2949_b1 , \2948_b1 , \2788_b1 );
xor ( \2949_b0 , \2948_b0 , w_6888 );
not ( w_6888 , w_6889 );
and ( w_6889 , \2788_b1 , \2788_b0 );
or ( \2950_b1 , \2947_b1 , \2949_b1 );
not ( \2949_b1 , w_6890 );
and ( \2950_b0 , \2947_b0 , w_6891 );
and ( w_6890 , w_6891 , \2949_b0 );
or ( \2951_b1 , \2771_b1 , \2773_b1 );
xor ( \2951_b0 , \2771_b0 , w_6892 );
not ( w_6892 , w_6893 );
and ( w_6893 , \2773_b1 , \2773_b0 );
or ( \2952_b1 , \2951_b1 , \2775_b1 );
xor ( \2952_b0 , \2951_b0 , w_6894 );
not ( w_6894 , w_6895 );
and ( w_6895 , \2775_b1 , \2775_b0 );
or ( \2953_b1 , \2949_b1 , \2952_b1 );
not ( \2952_b1 , w_6896 );
and ( \2953_b0 , \2949_b0 , w_6897 );
and ( w_6896 , w_6897 , \2952_b0 );
or ( \2954_b1 , \2947_b1 , \2952_b1 );
not ( \2952_b1 , w_6898 );
and ( \2954_b0 , \2947_b0 , w_6899 );
and ( w_6898 , w_6899 , \2952_b0 );
or ( \2956_b1 , \2937_b1 , \2955_b1 );
not ( \2955_b1 , w_6900 );
and ( \2956_b0 , \2937_b0 , w_6901 );
and ( w_6900 , w_6901 , \2955_b0 );
or ( \2957_b1 , \2522_b1 , \2539_b1 );
xor ( \2957_b0 , \2522_b0 , w_6902 );
not ( w_6902 , w_6903 );
and ( w_6903 , \2539_b1 , \2539_b0 );
or ( \2958_b1 , \2957_b1 , \2543_b1 );
xor ( \2958_b0 , \2957_b0 , w_6904 );
not ( w_6904 , w_6905 );
and ( w_6905 , \2543_b1 , \2543_b0 );
or ( \2959_b1 , \2955_b1 , \2958_b1 );
not ( \2958_b1 , w_6906 );
and ( \2959_b0 , \2955_b0 , w_6907 );
and ( w_6906 , w_6907 , \2958_b0 );
or ( \2960_b1 , \2937_b1 , \2958_b1 );
not ( \2958_b1 , w_6908 );
and ( \2960_b0 , \2937_b0 , w_6909 );
and ( w_6908 , w_6909 , \2958_b0 );
or ( \2962_b1 , \2565_b1 , \2581_b1 );
xor ( \2962_b0 , \2565_b0 , w_6910 );
not ( w_6910 , w_6911 );
and ( w_6911 , \2581_b1 , \2581_b0 );
or ( \2963_b1 , \2962_b1 , \2598_b1 );
xor ( \2963_b0 , \2962_b0 , w_6912 );
not ( w_6912 , w_6913 );
and ( w_6913 , \2598_b1 , \2598_b0 );
or ( \2964_b1 , \2725_b1 , \2768_b1 );
xor ( \2964_b0 , \2725_b0 , w_6914 );
not ( w_6914 , w_6915 );
and ( w_6915 , \2768_b1 , \2768_b0 );
or ( \2965_b1 , \2964_b1 , \2778_b1 );
xor ( \2965_b0 , \2964_b0 , w_6916 );
not ( w_6916 , w_6917 );
and ( w_6917 , \2778_b1 , \2778_b0 );
or ( \2966_b1 , \2963_b1 , \2965_b1 );
not ( \2965_b1 , w_6918 );
and ( \2966_b0 , \2963_b0 , w_6919 );
and ( w_6918 , w_6919 , \2965_b0 );
or ( \2967_b1 , \2791_b1 , \2793_b1 );
xor ( \2967_b0 , \2791_b0 , w_6920 );
not ( w_6920 , w_6921 );
and ( w_6921 , \2793_b1 , \2793_b0 );
or ( \2968_b1 , \2967_b1 , \2796_b1 );
xor ( \2968_b0 , \2967_b0 , w_6922 );
not ( w_6922 , w_6923 );
and ( w_6923 , \2796_b1 , \2796_b0 );
or ( \2969_b1 , \2965_b1 , \2968_b1 );
not ( \2968_b1 , w_6924 );
and ( \2969_b0 , \2965_b0 , w_6925 );
and ( w_6924 , w_6925 , \2968_b0 );
or ( \2970_b1 , \2963_b1 , \2968_b1 );
not ( \2968_b1 , w_6926 );
and ( \2970_b0 , \2963_b0 , w_6927 );
and ( w_6926 , w_6927 , \2968_b0 );
or ( \2972_b1 , \2961_b1 , \2971_b1 );
not ( \2971_b1 , w_6928 );
and ( \2972_b0 , \2961_b0 , w_6929 );
and ( w_6928 , w_6929 , \2971_b0 );
or ( \2973_b1 , \2624_b1 , \2626_b1 );
xor ( \2973_b0 , \2624_b0 , w_6930 );
not ( w_6930 , w_6931 );
and ( w_6931 , \2626_b1 , \2626_b0 );
or ( \2974_b1 , \2973_b1 , \2629_b1 );
xor ( \2974_b0 , \2973_b0 , w_6932 );
not ( w_6932 , w_6933 );
and ( w_6933 , \2629_b1 , \2629_b0 );
or ( \2975_b1 , \2971_b1 , \2974_b1 );
not ( \2974_b1 , w_6934 );
and ( \2975_b0 , \2971_b0 , w_6935 );
and ( w_6934 , w_6935 , \2974_b0 );
or ( \2976_b1 , \2961_b1 , \2974_b1 );
not ( \2974_b1 , w_6936 );
and ( \2976_b0 , \2961_b0 , w_6937 );
and ( w_6936 , w_6937 , \2974_b0 );
or ( \2978_b1 , \2546_b1 , \2601_b1 );
xor ( \2978_b0 , \2546_b0 , w_6938 );
not ( w_6938 , w_6939 );
and ( w_6939 , \2601_b1 , \2601_b0 );
or ( \2979_b1 , \2978_b1 , \2611_b1 );
xor ( \2979_b0 , \2978_b0 , w_6940 );
not ( w_6940 , w_6941 );
and ( w_6941 , \2611_b1 , \2611_b0 );
or ( \2980_b1 , \2781_b1 , \2799_b1 );
xor ( \2980_b0 , \2781_b0 , w_6942 );
not ( w_6942 , w_6943 );
and ( w_6943 , \2799_b1 , \2799_b0 );
or ( \2981_b1 , \2980_b1 , \2802_b1 );
xor ( \2981_b0 , \2980_b0 , w_6944 );
not ( w_6944 , w_6945 );
and ( w_6945 , \2802_b1 , \2802_b0 );
or ( \2982_b1 , \2979_b1 , \2981_b1 );
not ( \2981_b1 , w_6946 );
and ( \2982_b0 , \2979_b0 , w_6947 );
and ( w_6946 , w_6947 , \2981_b0 );
or ( \2983_b1 , \2977_b1 , \2982_b1 );
not ( \2982_b1 , w_6948 );
and ( \2983_b0 , \2977_b0 , w_6949 );
and ( w_6948 , w_6949 , \2982_b0 );
or ( \2984_b1 , \2805_b1 , \2807_b1 );
xor ( \2984_b0 , \2805_b0 , w_6950 );
not ( w_6950 , w_6951 );
and ( w_6951 , \2807_b1 , \2807_b0 );
or ( \2985_b1 , \2984_b1 , \2810_b1 );
xor ( \2985_b0 , \2984_b0 , w_6952 );
not ( w_6952 , w_6953 );
and ( w_6953 , \2810_b1 , \2810_b0 );
or ( \2986_b1 , \2982_b1 , \2985_b1 );
not ( \2985_b1 , w_6954 );
and ( \2986_b0 , \2982_b0 , w_6955 );
and ( w_6954 , w_6955 , \2985_b0 );
or ( \2987_b1 , \2977_b1 , \2985_b1 );
not ( \2985_b1 , w_6956 );
and ( \2987_b0 , \2977_b0 , w_6957 );
and ( w_6956 , w_6957 , \2985_b0 );
or ( \2989_b1 , \2824_b1 , \2988_b1 );
not ( \2988_b1 , w_6958 );
and ( \2989_b0 , \2824_b0 , w_6959 );
and ( w_6958 , w_6959 , \2988_b0 );
or ( \2990_b1 , \2824_b1 , \2988_b1 );
xor ( \2990_b0 , \2824_b0 , w_6960 );
not ( w_6960 , w_6961 );
and ( w_6961 , \2988_b1 , \2988_b0 );
or ( \2991_b1 , \2977_b1 , \2982_b1 );
xor ( \2991_b0 , \2977_b0 , w_6962 );
not ( w_6962 , w_6963 );
and ( w_6963 , \2982_b1 , \2982_b0 );
or ( \2992_b1 , \2991_b1 , \2985_b1 );
xor ( \2992_b0 , \2991_b0 , w_6964 );
not ( w_6964 , w_6965 );
and ( w_6965 , \2985_b1 , \2985_b0 );
or ( \2993_b1 , \360_b1 , \1955_b1 );
not ( \1955_b1 , w_6966 );
and ( \2993_b0 , \360_b0 , w_6967 );
and ( w_6966 , w_6967 , \1955_b0 );
or ( \2994_b1 , \343_b1 , \1953_b1 );
not ( \1953_b1 , w_6968 );
and ( \2994_b0 , \343_b0 , w_6969 );
and ( w_6968 , w_6969 , \1953_b0 );
or ( \2995_b1 , \2993_b1 , w_6971 );
not ( w_6971 , w_6972 );
and ( \2995_b0 , \2993_b0 , w_6973 );
and ( w_6972 ,  , w_6973 );
buf ( w_6971 , \2994_b1 );
not ( w_6971 , w_6974 );
not (  , w_6975 );
and ( w_6974 , w_6975 , \2994_b0 );
or ( \2996_b1 , \2995_b1 , w_6976 );
xor ( \2996_b0 , \2995_b0 , w_6978 );
not ( w_6978 , w_6979 );
and ( w_6979 , w_6976 , w_6977 );
buf ( w_6976 , \1835_b1 );
not ( w_6976 , w_6980 );
not ( w_6977 , w_6981 );
and ( w_6980 , w_6981 , \1835_b0 );
or ( \2997_b1 , \495_b1 , \1742_b1 );
not ( \1742_b1 , w_6982 );
and ( \2997_b0 , \495_b0 , w_6983 );
and ( w_6982 , w_6983 , \1742_b0 );
or ( \2998_b1 , \444_b1 , \1740_b1 );
not ( \1740_b1 , w_6984 );
and ( \2998_b0 , \444_b0 , w_6985 );
and ( w_6984 , w_6985 , \1740_b0 );
or ( \2999_b1 , \2997_b1 , w_6987 );
not ( w_6987 , w_6988 );
and ( \2999_b0 , \2997_b0 , w_6989 );
and ( w_6988 ,  , w_6989 );
buf ( w_6987 , \2998_b1 );
not ( w_6987 , w_6990 );
not (  , w_6991 );
and ( w_6990 , w_6991 , \2998_b0 );
or ( \3000_b1 , \2999_b1 , w_6992 );
xor ( \3000_b0 , \2999_b0 , w_6994 );
not ( w_6994 , w_6995 );
and ( w_6995 , w_6992 , w_6993 );
buf ( w_6992 , \1610_b1 );
not ( w_6992 , w_6996 );
not ( w_6993 , w_6997 );
and ( w_6996 , w_6997 , \1610_b0 );
or ( \3001_b1 , \2996_b1 , \3000_b1 );
not ( \3000_b1 , w_6998 );
and ( \3001_b0 , \2996_b0 , w_6999 );
and ( w_6998 , w_6999 , \3000_b0 );
or ( \3002_b1 , \621_b1 , \1476_b1 );
not ( \1476_b1 , w_7000 );
and ( \3002_b0 , \621_b0 , w_7001 );
and ( w_7000 , w_7001 , \1476_b0 );
or ( \3003_b1 , \593_b1 , \1474_b1 );
not ( \1474_b1 , w_7002 );
and ( \3003_b0 , \593_b0 , w_7003 );
and ( w_7002 , w_7003 , \1474_b0 );
or ( \3004_b1 , \3002_b1 , w_7005 );
not ( w_7005 , w_7006 );
and ( \3004_b0 , \3002_b0 , w_7007 );
and ( w_7006 ,  , w_7007 );
buf ( w_7005 , \3003_b1 );
not ( w_7005 , w_7008 );
not (  , w_7009 );
and ( w_7008 , w_7009 , \3003_b0 );
or ( \3005_b1 , \3004_b1 , w_7010 );
xor ( \3005_b0 , \3004_b0 , w_7012 );
not ( w_7012 , w_7013 );
and ( w_7013 , w_7010 , w_7011 );
buf ( w_7010 , \1363_b1 );
not ( w_7010 , w_7014 );
not ( w_7011 , w_7015 );
and ( w_7014 , w_7015 , \1363_b0 );
or ( \3006_b1 , \3000_b1 , \3005_b1 );
not ( \3005_b1 , w_7016 );
and ( \3006_b0 , \3000_b0 , w_7017 );
and ( w_7016 , w_7017 , \3005_b0 );
or ( \3007_b1 , \2996_b1 , \3005_b1 );
not ( \3005_b1 , w_7018 );
and ( \3007_b0 , \2996_b0 , w_7019 );
and ( w_7018 , w_7019 , \3005_b0 );
or ( \3009_b1 , \315_b1 , \2913_b1 );
not ( \2913_b1 , w_7020 );
and ( \3009_b0 , \315_b0 , w_7021 );
and ( w_7020 , w_7021 , \2913_b0 );
or ( \3010_b1 , \159_b1 , \2910_b1 );
not ( \2910_b1 , w_7022 );
and ( \3010_b0 , \159_b0 , w_7023 );
and ( w_7022 , w_7023 , \2910_b0 );
or ( \3011_b1 , \3009_b1 , w_7025 );
not ( w_7025 , w_7026 );
and ( \3011_b0 , \3009_b0 , w_7027 );
and ( w_7026 ,  , w_7027 );
buf ( w_7025 , \3010_b1 );
not ( w_7025 , w_7028 );
not (  , w_7029 );
and ( w_7028 , w_7029 , \3010_b0 );
or ( \3012_b1 , \3011_b1 , w_7030 );
xor ( \3012_b0 , \3011_b0 , w_7032 );
not ( w_7032 , w_7033 );
and ( w_7033 , w_7030 , w_7031 );
buf ( w_7030 , \2371_b1 );
not ( w_7030 , w_7034 );
not ( w_7031 , w_7035 );
and ( w_7034 , w_7035 , \2371_b0 );
or ( \3013_b1 , \333_b1 , \2550_b1 );
not ( \2550_b1 , w_7036 );
and ( \3013_b0 , \333_b0 , w_7037 );
and ( w_7036 , w_7037 , \2550_b0 );
or ( \3014_b1 , \305_b1 , \2548_b1 );
not ( \2548_b1 , w_7038 );
and ( \3014_b0 , \305_b0 , w_7039 );
and ( w_7038 , w_7039 , \2548_b0 );
or ( \3015_b1 , \3013_b1 , w_7041 );
not ( w_7041 , w_7042 );
and ( \3015_b0 , \3013_b0 , w_7043 );
and ( w_7042 ,  , w_7043 );
buf ( w_7041 , \3014_b1 );
not ( w_7041 , w_7044 );
not (  , w_7045 );
and ( w_7044 , w_7045 , \3014_b0 );
or ( \3016_b1 , \3015_b1 , w_7046 );
xor ( \3016_b0 , \3015_b0 , w_7048 );
not ( w_7048 , w_7049 );
and ( w_7049 , w_7046 , w_7047 );
buf ( w_7046 , \2374_b1 );
not ( w_7046 , w_7050 );
not ( w_7047 , w_7051 );
and ( w_7050 , w_7051 , \2374_b0 );
or ( \3017_b1 , \3012_b1 , \3016_b1 );
not ( \3016_b1 , w_7052 );
and ( \3017_b0 , \3012_b0 , w_7053 );
and ( w_7052 , w_7053 , \3016_b0 );
or ( \3018_b1 , \353_b1 , \2261_b1 );
not ( \2261_b1 , w_7054 );
and ( \3018_b0 , \353_b0 , w_7055 );
and ( w_7054 , w_7055 , \2261_b0 );
or ( \3019_b1 , \323_b1 , \2259_b1 );
not ( \2259_b1 , w_7056 );
and ( \3019_b0 , \323_b0 , w_7057 );
and ( w_7056 , w_7057 , \2259_b0 );
or ( \3020_b1 , \3018_b1 , w_7059 );
not ( w_7059 , w_7060 );
and ( \3020_b0 , \3018_b0 , w_7061 );
and ( w_7060 ,  , w_7061 );
buf ( w_7059 , \3019_b1 );
not ( w_7059 , w_7062 );
not (  , w_7063 );
and ( w_7062 , w_7063 , \3019_b0 );
or ( \3021_b1 , \3020_b1 , w_7064 );
xor ( \3021_b0 , \3020_b0 , w_7066 );
not ( w_7066 , w_7067 );
and ( w_7067 , w_7064 , w_7065 );
buf ( w_7064 , \2124_b1 );
not ( w_7064 , w_7068 );
not ( w_7065 , w_7069 );
and ( w_7068 , w_7069 , \2124_b0 );
or ( \3022_b1 , \3016_b1 , \3021_b1 );
not ( \3021_b1 , w_7070 );
and ( \3022_b0 , \3016_b0 , w_7071 );
and ( w_7070 , w_7071 , \3021_b0 );
or ( \3023_b1 , \3012_b1 , \3021_b1 );
not ( \3021_b1 , w_7072 );
and ( \3023_b0 , \3012_b0 , w_7073 );
and ( w_7072 , w_7073 , \3021_b0 );
or ( \3025_b1 , \3008_b1 , \3024_b1 );
not ( \3024_b1 , w_7074 );
and ( \3025_b0 , \3008_b0 , w_7075 );
and ( w_7074 , w_7075 , \3024_b0 );
or ( \3026_b1 , \777_b1 , \1280_b1 );
not ( \1280_b1 , w_7076 );
and ( \3026_b0 , \777_b0 , w_7077 );
and ( w_7076 , w_7077 , \1280_b0 );
or ( \3027_b1 , \703_b1 , \1278_b1 );
not ( \1278_b1 , w_7078 );
and ( \3027_b0 , \703_b0 , w_7079 );
and ( w_7078 , w_7079 , \1278_b0 );
or ( \3028_b1 , \3026_b1 , w_7081 );
not ( w_7081 , w_7082 );
and ( \3028_b0 , \3026_b0 , w_7083 );
and ( w_7082 ,  , w_7083 );
buf ( w_7081 , \3027_b1 );
not ( w_7081 , w_7084 );
not (  , w_7085 );
and ( w_7084 , w_7085 , \3027_b0 );
or ( \3029_b1 , \3028_b1 , w_7086 );
xor ( \3029_b0 , \3028_b0 , w_7088 );
not ( w_7088 , w_7089 );
and ( w_7089 , w_7086 , w_7087 );
buf ( w_7086 , \1177_b1 );
not ( w_7086 , w_7090 );
not ( w_7087 , w_7091 );
and ( w_7090 , w_7091 , \1177_b0 );
or ( \3030_b1 , \904_b1 , \1062_b1 );
not ( \1062_b1 , w_7092 );
and ( \3030_b0 , \904_b0 , w_7093 );
and ( w_7092 , w_7093 , \1062_b0 );
or ( \3031_b1 , \841_b1 , \1060_b1 );
not ( \1060_b1 , w_7094 );
and ( \3031_b0 , \841_b0 , w_7095 );
and ( w_7094 , w_7095 , \1060_b0 );
or ( \3032_b1 , \3030_b1 , w_7097 );
not ( w_7097 , w_7098 );
and ( \3032_b0 , \3030_b0 , w_7099 );
and ( w_7098 ,  , w_7099 );
buf ( w_7097 , \3031_b1 );
not ( w_7097 , w_7100 );
not (  , w_7101 );
and ( w_7100 , w_7101 , \3031_b0 );
or ( \3033_b1 , \3032_b1 , w_7102 );
xor ( \3033_b0 , \3032_b0 , w_7104 );
not ( w_7104 , w_7105 );
and ( w_7105 , w_7102 , w_7103 );
buf ( w_7102 , \984_b1 );
not ( w_7102 , w_7106 );
not ( w_7103 , w_7107 );
and ( w_7106 , w_7107 , \984_b0 );
or ( \3034_b1 , \3029_b1 , \3033_b1 );
not ( \3033_b1 , w_7108 );
and ( \3034_b0 , \3029_b0 , w_7109 );
and ( w_7108 , w_7109 , \3033_b0 );
or ( \3035_b1 , \1194_b1 , \912_b1 );
not ( \912_b1 , w_7110 );
and ( \3035_b0 , \1194_b0 , w_7111 );
and ( w_7110 , w_7111 , \912_b0 );
or ( \3036_b1 , \1104_b1 , \910_b1 );
not ( \910_b1 , w_7112 );
and ( \3036_b0 , \1104_b0 , w_7113 );
and ( w_7112 , w_7113 , \910_b0 );
or ( \3037_b1 , \3035_b1 , w_7115 );
not ( w_7115 , w_7116 );
and ( \3037_b0 , \3035_b0 , w_7117 );
and ( w_7116 ,  , w_7117 );
buf ( w_7115 , \3036_b1 );
not ( w_7115 , w_7118 );
not (  , w_7119 );
and ( w_7118 , w_7119 , \3036_b0 );
or ( \3038_b1 , \3037_b1 , w_7120 );
xor ( \3038_b0 , \3037_b0 , w_7122 );
not ( w_7122 , w_7123 );
and ( w_7123 , w_7120 , w_7121 );
buf ( w_7120 , \818_b1 );
not ( w_7120 , w_7124 );
not ( w_7121 , w_7125 );
and ( w_7124 , w_7125 , \818_b0 );
or ( \3039_b1 , \3033_b1 , \3038_b1 );
not ( \3038_b1 , w_7126 );
and ( \3039_b0 , \3033_b0 , w_7127 );
and ( w_7126 , w_7127 , \3038_b0 );
or ( \3040_b1 , \3029_b1 , \3038_b1 );
not ( \3038_b1 , w_7128 );
and ( \3040_b0 , \3029_b0 , w_7129 );
and ( w_7128 , w_7129 , \3038_b0 );
or ( \3042_b1 , \3024_b1 , \3041_b1 );
not ( \3041_b1 , w_7130 );
and ( \3042_b0 , \3024_b0 , w_7131 );
and ( w_7130 , w_7131 , \3041_b0 );
or ( \3043_b1 , \3008_b1 , \3041_b1 );
not ( \3041_b1 , w_7132 );
and ( \3043_b0 , \3008_b0 , w_7133 );
and ( w_7132 , w_7133 , \3041_b0 );
or ( \3045_b1 , \2828_b1 , \2832_b1 );
xor ( \3045_b0 , \2828_b0 , w_7134 );
not ( w_7134 , w_7135 );
and ( w_7135 , \2832_b1 , \2832_b0 );
or ( \3046_b1 , \3045_b1 , \2837_b1 );
xor ( \3046_b0 , \3045_b0 , w_7136 );
not ( w_7136 , w_7137 );
and ( w_7137 , \2837_b1 , \2837_b0 );
or ( \3047_b1 , \2879_b1 , \2883_b1 );
xor ( \3047_b0 , \2879_b0 , w_7138 );
not ( w_7138 , w_7139 );
and ( w_7139 , \2883_b1 , \2883_b0 );
or ( \3048_b1 , \3047_b1 , \2888_b1 );
xor ( \3048_b0 , \3047_b0 , w_7140 );
not ( w_7140 , w_7141 );
and ( w_7141 , \2888_b1 , \2888_b0 );
or ( \3049_b1 , \3046_b1 , \3048_b1 );
not ( \3048_b1 , w_7142 );
and ( \3049_b0 , \3046_b0 , w_7143 );
and ( w_7142 , w_7143 , \3048_b0 );
or ( \3050_b1 , \2860_b1 , \2864_b1 );
xor ( \3050_b0 , \2860_b0 , w_7144 );
not ( w_7144 , w_7145 );
and ( w_7145 , \2864_b1 , \2864_b0 );
or ( \3051_b1 , \3050_b1 , \2869_b1 );
xor ( \3051_b0 , \3050_b0 , w_7146 );
not ( w_7146 , w_7147 );
and ( w_7147 , \2869_b1 , \2869_b0 );
or ( \3052_b1 , \3048_b1 , \3051_b1 );
not ( \3051_b1 , w_7148 );
and ( \3052_b0 , \3048_b0 , w_7149 );
and ( w_7148 , w_7149 , \3051_b0 );
or ( \3053_b1 , \3046_b1 , \3051_b1 );
not ( \3051_b1 , w_7150 );
and ( \3053_b0 , \3046_b0 , w_7151 );
and ( w_7150 , w_7151 , \3051_b0 );
or ( \3055_b1 , \3044_b1 , \3054_b1 );
not ( \3054_b1 , w_7152 );
and ( \3055_b0 , \3044_b0 , w_7153 );
and ( w_7152 , w_7153 , \3054_b0 );
or ( \3056_b1 , \1304_b1 , \740_b1 );
not ( \740_b1 , w_7154 );
and ( \3056_b0 , \1304_b0 , w_7155 );
and ( w_7154 , w_7155 , \740_b0 );
or ( \3057_b1 , \1299_b1 , \738_b1 );
not ( \738_b1 , w_7156 );
and ( \3057_b0 , \1299_b0 , w_7157 );
and ( w_7156 , w_7157 , \738_b0 );
or ( \3058_b1 , \3056_b1 , w_7159 );
not ( w_7159 , w_7160 );
and ( \3058_b0 , \3056_b0 , w_7161 );
and ( w_7160 ,  , w_7161 );
buf ( w_7159 , \3057_b1 );
not ( w_7159 , w_7162 );
not (  , w_7163 );
and ( w_7162 , w_7163 , \3057_b0 );
or ( \3059_b1 , \3058_b1 , w_7164 );
xor ( \3059_b0 , \3058_b0 , w_7166 );
not ( w_7166 , w_7167 );
and ( w_7167 , w_7164 , w_7165 );
buf ( w_7164 , \668_b1 );
not ( w_7164 , w_7168 );
not ( w_7165 , w_7169 );
and ( w_7168 , w_7169 , \668_b0 );
or ( \3060_b1 , \1537_b1 , \604_b1 );
not ( \604_b1 , w_7170 );
and ( \3060_b0 , \1537_b0 , w_7171 );
and ( w_7170 , w_7171 , \604_b0 );
or ( \3061_b1 , \1422_b1 , \602_b1 );
not ( \602_b1 , w_7172 );
and ( \3061_b0 , \1422_b0 , w_7173 );
and ( w_7172 , w_7173 , \602_b0 );
or ( \3062_b1 , \3060_b1 , w_7175 );
not ( w_7175 , w_7176 );
and ( \3062_b0 , \3060_b0 , w_7177 );
and ( w_7176 ,  , w_7177 );
buf ( w_7175 , \3061_b1 );
not ( w_7175 , w_7178 );
not (  , w_7179 );
and ( w_7178 , w_7179 , \3061_b0 );
or ( \3063_b1 , \3062_b1 , w_7180 );
xor ( \3063_b0 , \3062_b0 , w_7182 );
not ( w_7182 , w_7183 );
and ( w_7183 , w_7180 , w_7181 );
buf ( w_7180 , \561_b1 );
not ( w_7180 , w_7184 );
not ( w_7181 , w_7185 );
and ( w_7184 , w_7185 , \561_b0 );
or ( \3064_b1 , \3059_b1 , \3063_b1 );
not ( \3063_b1 , w_7186 );
and ( \3064_b0 , \3059_b0 , w_7187 );
and ( w_7186 , w_7187 , \3063_b0 );
or ( \3065_b1 , \1778_b1 , \503_b1 );
not ( \503_b1 , w_7188 );
and ( \3065_b0 , \1778_b0 , w_7189 );
and ( w_7188 , w_7189 , \503_b0 );
or ( \3066_b1 , \1770_b1 , \501_b1 );
not ( \501_b1 , w_7190 );
and ( \3066_b0 , \1770_b0 , w_7191 );
and ( w_7190 , w_7191 , \501_b0 );
or ( \3067_b1 , \3065_b1 , w_7193 );
not ( w_7193 , w_7194 );
and ( \3067_b0 , \3065_b0 , w_7195 );
and ( w_7194 ,  , w_7195 );
buf ( w_7193 , \3066_b1 );
not ( w_7193 , w_7196 );
not (  , w_7197 );
and ( w_7196 , w_7197 , \3066_b0 );
or ( \3068_b1 , \3067_b1 , w_7198 );
xor ( \3068_b0 , \3067_b0 , w_7200 );
not ( w_7200 , w_7201 );
and ( w_7201 , w_7198 , w_7199 );
buf ( w_7198 , \455_b1 );
not ( w_7198 , w_7202 );
not ( w_7199 , w_7203 );
and ( w_7202 , w_7203 , \455_b0 );
or ( \3069_b1 , \3063_b1 , \3068_b1 );
not ( \3068_b1 , w_7204 );
and ( \3069_b0 , \3063_b0 , w_7205 );
and ( w_7204 , w_7205 , \3068_b0 );
or ( \3070_b1 , \3059_b1 , \3068_b1 );
not ( \3068_b1 , w_7206 );
and ( \3070_b0 , \3059_b0 , w_7207 );
and ( w_7206 , w_7207 , \3068_b0 );
or ( \3072_b1 , \2028_b1 , \298_b1 );
not ( \298_b1 , w_7208 );
and ( \3072_b0 , \2028_b0 , w_7209 );
and ( w_7208 , w_7209 , \298_b0 );
or ( \3073_b1 , \2023_b1 , \296_b1 );
not ( \296_b1 , w_7210 );
and ( \3073_b0 , \2023_b0 , w_7211 );
and ( w_7210 , w_7211 , \296_b0 );
or ( \3074_b1 , \3072_b1 , w_7213 );
not ( w_7213 , w_7214 );
and ( \3074_b0 , \3072_b0 , w_7215 );
and ( w_7214 ,  , w_7215 );
buf ( w_7213 , \3073_b1 );
not ( w_7213 , w_7216 );
not (  , w_7217 );
and ( w_7216 , w_7217 , \3073_b0 );
or ( \3075_b1 , \3074_b1 , w_7218 );
xor ( \3075_b0 , \3074_b0 , w_7220 );
not ( w_7220 , w_7221 );
and ( w_7221 , w_7218 , w_7219 );
buf ( w_7218 , \303_b1 );
not ( w_7218 , w_7222 );
not ( w_7219 , w_7223 );
and ( w_7222 , w_7223 , \303_b0 );
or ( \3076_b1 , \2305_b1 , \313_b1 );
not ( \313_b1 , w_7224 );
and ( \3076_b0 , \2305_b0 , w_7225 );
and ( w_7224 , w_7225 , \313_b0 );
or ( \3077_b1 , \2161_b1 , \311_b1 );
not ( \311_b1 , w_7226 );
and ( \3077_b0 , \2161_b0 , w_7227 );
and ( w_7226 , w_7227 , \311_b0 );
or ( \3078_b1 , \3076_b1 , w_7229 );
not ( w_7229 , w_7230 );
and ( \3078_b0 , \3076_b0 , w_7231 );
and ( w_7230 ,  , w_7231 );
buf ( w_7229 , \3077_b1 );
not ( w_7229 , w_7232 );
not (  , w_7233 );
and ( w_7232 , w_7233 , \3077_b0 );
or ( \3079_b1 , \3078_b1 , w_7234 );
xor ( \3079_b0 , \3078_b0 , w_7236 );
not ( w_7236 , w_7237 );
and ( w_7237 , w_7234 , w_7235 );
buf ( w_7234 , \320_b1 );
not ( w_7234 , w_7238 );
not ( w_7235 , w_7239 );
and ( w_7238 , w_7239 , \320_b0 );
or ( \3080_b1 , \3075_b1 , \3079_b1 );
not ( \3079_b1 , w_7240 );
and ( \3080_b0 , \3075_b0 , w_7241 );
and ( w_7240 , w_7241 , \3079_b0 );
or ( \3081_b1 , \2541_b1 , \331_b1 );
not ( \331_b1 , w_7242 );
and ( \3081_b0 , \2541_b0 , w_7243 );
and ( w_7242 , w_7243 , \331_b0 );
or ( \3082_b1 , \2532_b1 , \329_b1 );
not ( \329_b1 , w_7244 );
and ( \3082_b0 , \2532_b0 , w_7245 );
and ( w_7244 , w_7245 , \329_b0 );
or ( \3083_b1 , \3081_b1 , w_7247 );
not ( w_7247 , w_7248 );
and ( \3083_b0 , \3081_b0 , w_7249 );
and ( w_7248 ,  , w_7249 );
buf ( w_7247 , \3082_b1 );
not ( w_7247 , w_7250 );
not (  , w_7251 );
and ( w_7250 , w_7251 , \3082_b0 );
or ( \3084_b1 , \3083_b1 , w_7252 );
xor ( \3084_b0 , \3083_b0 , w_7254 );
not ( w_7254 , w_7255 );
and ( w_7255 , w_7252 , w_7253 );
buf ( w_7252 , \338_b1 );
not ( w_7252 , w_7256 );
not ( w_7253 , w_7257 );
and ( w_7256 , w_7257 , \338_b0 );
or ( \3085_b1 , \3079_b1 , \3084_b1 );
not ( \3084_b1 , w_7258 );
and ( \3085_b0 , \3079_b0 , w_7259 );
and ( w_7258 , w_7259 , \3084_b0 );
or ( \3086_b1 , \3075_b1 , \3084_b1 );
not ( \3084_b1 , w_7260 );
and ( \3086_b0 , \3075_b0 , w_7261 );
and ( w_7260 , w_7261 , \3084_b0 );
or ( \3088_b1 , \3071_b1 , \3087_b1 );
not ( \3087_b1 , w_7262 );
and ( \3088_b0 , \3071_b0 , w_7263 );
and ( w_7262 , w_7263 , \3087_b0 );
or ( \3089_b1 , \2844_b1 , \2848_b1 );
xor ( \3089_b0 , \2844_b0 , w_7264 );
not ( w_7264 , w_7265 );
and ( w_7265 , \2848_b1 , \2848_b0 );
or ( \3090_b1 , \3089_b1 , \2852_b1 );
xor ( \3090_b0 , \3089_b0 , w_7266 );
not ( w_7266 , w_7267 );
and ( w_7267 , \2852_b1 , \2852_b0 );
or ( \3091_b1 , \3087_b1 , \3090_b1 );
not ( \3090_b1 , w_7268 );
and ( \3091_b0 , \3087_b0 , w_7269 );
and ( w_7268 , w_7269 , \3090_b0 );
or ( \3092_b1 , \3071_b1 , \3090_b1 );
not ( \3090_b1 , w_7270 );
and ( \3092_b0 , \3071_b0 , w_7271 );
and ( w_7270 , w_7271 , \3090_b0 );
or ( \3094_b1 , \3054_b1 , \3093_b1 );
not ( \3093_b1 , w_7272 );
and ( \3094_b0 , \3054_b0 , w_7273 );
and ( w_7272 , w_7273 , \3093_b0 );
or ( \3095_b1 , \3044_b1 , \3093_b1 );
not ( \3093_b1 , w_7274 );
and ( \3095_b0 , \3044_b0 , w_7275 );
and ( w_7274 , w_7275 , \3093_b0 );
or ( \3097_b1 , \2840_b1 , \2855_b1 );
xor ( \3097_b0 , \2840_b0 , w_7276 );
not ( w_7276 , w_7277 );
and ( w_7277 , \2855_b1 , \2855_b0 );
or ( \3098_b1 , \3097_b1 , \2872_b1 );
xor ( \3098_b0 , \3097_b0 , w_7278 );
not ( w_7278 , w_7279 );
and ( w_7279 , \2872_b1 , \2872_b0 );
or ( \3099_b1 , \2939_b1 , \2941_b1 );
xor ( \3099_b0 , \2939_b0 , w_7280 );
not ( w_7280 , w_7281 );
and ( w_7281 , \2941_b1 , \2941_b0 );
or ( \3100_b1 , \3099_b1 , \2944_b1 );
xor ( \3100_b0 , \3099_b0 , w_7282 );
not ( w_7282 , w_7283 );
and ( w_7283 , \2944_b1 , \2944_b0 );
or ( \3101_b1 , \3098_b1 , \3100_b1 );
not ( \3100_b1 , w_7284 );
and ( \3101_b0 , \3098_b0 , w_7285 );
and ( w_7284 , w_7285 , \3100_b0 );
or ( \3102_b1 , \2927_b1 , \2929_b1 );
xor ( \3102_b0 , \2927_b0 , w_7286 );
not ( w_7286 , w_7287 );
and ( w_7287 , \2929_b1 , \2929_b0 );
or ( \3103_b1 , \3102_b1 , \2931_b1 );
xor ( \3103_b0 , \3102_b0 , w_7288 );
not ( w_7288 , w_7289 );
and ( w_7289 , \2931_b1 , \2931_b0 );
or ( \3104_b1 , \3100_b1 , \3103_b1 );
not ( \3103_b1 , w_7290 );
and ( \3104_b0 , \3100_b0 , w_7291 );
and ( w_7290 , w_7291 , \3103_b0 );
or ( \3105_b1 , \3098_b1 , \3103_b1 );
not ( \3103_b1 , w_7292 );
and ( \3105_b0 , \3098_b0 , w_7293 );
and ( w_7292 , w_7293 , \3103_b0 );
or ( \3107_b1 , \3096_b1 , \3106_b1 );
not ( \3106_b1 , w_7294 );
and ( \3107_b0 , \3096_b0 , w_7295 );
and ( w_7294 , w_7295 , \3106_b0 );
or ( \3108_b1 , \2741_b1 , \2757_b1 );
xor ( \3108_b0 , \2741_b0 , w_7296 );
not ( w_7296 , w_7297 );
and ( w_7297 , \2757_b1 , \2757_b0 );
or ( \3109_b1 , \3108_b1 , \2765_b1 );
xor ( \3109_b0 , \3108_b0 , w_7298 );
not ( w_7298 , w_7299 );
and ( w_7299 , \2765_b1 , \2765_b0 );
or ( \3110_b1 , \3106_b1 , \3109_b1 );
not ( \3109_b1 , w_7300 );
and ( \3110_b0 , \3106_b0 , w_7301 );
and ( w_7300 , w_7301 , \3109_b0 );
or ( \3111_b1 , \3096_b1 , \3109_b1 );
not ( \3109_b1 , w_7302 );
and ( \3111_b0 , \3096_b0 , w_7303 );
and ( w_7302 , w_7303 , \3109_b0 );
or ( \3113_b1 , \2692_b1 , \2705_b1 );
xor ( \3113_b0 , \2692_b0 , w_7304 );
not ( w_7304 , w_7305 );
and ( w_7305 , \2705_b1 , \2705_b0 );
or ( \3114_b1 , \3113_b1 , \2722_b1 );
xor ( \3114_b0 , \3113_b0 , w_7306 );
not ( w_7306 , w_7307 );
and ( w_7307 , \2722_b1 , \2722_b0 );
or ( \3115_b1 , \2875_b1 , \2924_b1 );
xor ( \3115_b0 , \2875_b0 , w_7308 );
not ( w_7308 , w_7309 );
and ( w_7309 , \2924_b1 , \2924_b0 );
or ( \3116_b1 , \3115_b1 , \2934_b1 );
xor ( \3116_b0 , \3115_b0 , w_7310 );
not ( w_7310 , w_7311 );
and ( w_7311 , \2934_b1 , \2934_b0 );
or ( \3117_b1 , \3114_b1 , \3116_b1 );
not ( \3116_b1 , w_7312 );
and ( \3117_b0 , \3114_b0 , w_7313 );
and ( w_7312 , w_7313 , \3116_b0 );
or ( \3118_b1 , \2947_b1 , \2949_b1 );
xor ( \3118_b0 , \2947_b0 , w_7314 );
not ( w_7314 , w_7315 );
and ( w_7315 , \2949_b1 , \2949_b0 );
or ( \3119_b1 , \3118_b1 , \2952_b1 );
xor ( \3119_b0 , \3118_b0 , w_7316 );
not ( w_7316 , w_7317 );
and ( w_7317 , \2952_b1 , \2952_b0 );
or ( \3120_b1 , \3116_b1 , \3119_b1 );
not ( \3119_b1 , w_7318 );
and ( \3120_b0 , \3116_b0 , w_7319 );
and ( w_7318 , w_7319 , \3119_b0 );
or ( \3121_b1 , \3114_b1 , \3119_b1 );
not ( \3119_b1 , w_7320 );
and ( \3121_b0 , \3114_b0 , w_7321 );
and ( w_7320 , w_7321 , \3119_b0 );
or ( \3123_b1 , \3112_b1 , \3122_b1 );
not ( \3122_b1 , w_7322 );
and ( \3123_b0 , \3112_b0 , w_7323 );
and ( w_7322 , w_7323 , \3122_b0 );
or ( \3124_b1 , \2963_b1 , \2965_b1 );
xor ( \3124_b0 , \2963_b0 , w_7324 );
not ( w_7324 , w_7325 );
and ( w_7325 , \2965_b1 , \2965_b0 );
or ( \3125_b1 , \3124_b1 , \2968_b1 );
xor ( \3125_b0 , \3124_b0 , w_7326 );
not ( w_7326 , w_7327 );
and ( w_7327 , \2968_b1 , \2968_b0 );
or ( \3126_b1 , \3122_b1 , \3125_b1 );
not ( \3125_b1 , w_7328 );
and ( \3126_b0 , \3122_b0 , w_7329 );
and ( w_7328 , w_7329 , \3125_b0 );
or ( \3127_b1 , \3112_b1 , \3125_b1 );
not ( \3125_b1 , w_7330 );
and ( \3127_b0 , \3112_b0 , w_7331 );
and ( w_7330 , w_7331 , \3125_b0 );
or ( \3129_b1 , \2961_b1 , \2971_b1 );
xor ( \3129_b0 , \2961_b0 , w_7332 );
not ( w_7332 , w_7333 );
and ( w_7333 , \2971_b1 , \2971_b0 );
or ( \3130_b1 , \3129_b1 , \2974_b1 );
xor ( \3130_b0 , \3129_b0 , w_7334 );
not ( w_7334 , w_7335 );
and ( w_7335 , \2974_b1 , \2974_b0 );
or ( \3131_b1 , \3128_b1 , \3130_b1 );
not ( \3130_b1 , w_7336 );
and ( \3131_b0 , \3128_b0 , w_7337 );
and ( w_7336 , w_7337 , \3130_b0 );
or ( \3132_b1 , \2979_b1 , \2981_b1 );
xor ( \3132_b0 , \2979_b0 , w_7338 );
not ( w_7338 , w_7339 );
and ( w_7339 , \2981_b1 , \2981_b0 );
or ( \3133_b1 , \3130_b1 , \3132_b1 );
not ( \3132_b1 , w_7340 );
and ( \3133_b0 , \3130_b0 , w_7341 );
and ( w_7340 , w_7341 , \3132_b0 );
or ( \3134_b1 , \3128_b1 , \3132_b1 );
not ( \3132_b1 , w_7342 );
and ( \3134_b0 , \3128_b0 , w_7343 );
and ( w_7342 , w_7343 , \3132_b0 );
or ( \3136_b1 , \2992_b1 , \3135_b1 );
not ( \3135_b1 , w_7344 );
and ( \3136_b0 , \2992_b0 , w_7345 );
and ( w_7344 , w_7345 , \3135_b0 );
or ( \3137_b1 , \2992_b1 , \3135_b1 );
xor ( \3137_b0 , \2992_b0 , w_7346 );
not ( w_7346 , w_7347 );
and ( w_7347 , \3135_b1 , \3135_b0 );
or ( \3138_b1 , \3128_b1 , \3130_b1 );
xor ( \3138_b0 , \3128_b0 , w_7348 );
not ( w_7348 , w_7349 );
and ( w_7349 , \3130_b1 , \3130_b0 );
or ( \3139_b1 , \3138_b1 , \3132_b1 );
xor ( \3139_b0 , \3138_b0 , w_7350 );
not ( w_7350 , w_7351 );
and ( w_7351 , \3132_b1 , \3132_b0 );
or ( \3140_b1 , \343_b1 , \2261_b1 );
not ( \2261_b1 , w_7352 );
and ( \3140_b0 , \343_b0 , w_7353 );
and ( w_7352 , w_7353 , \2261_b0 );
or ( \3141_b1 , \353_b1 , \2259_b1 );
not ( \2259_b1 , w_7354 );
and ( \3141_b0 , \353_b0 , w_7355 );
and ( w_7354 , w_7355 , \2259_b0 );
or ( \3142_b1 , \3140_b1 , w_7357 );
not ( w_7357 , w_7358 );
and ( \3142_b0 , \3140_b0 , w_7359 );
and ( w_7358 ,  , w_7359 );
buf ( w_7357 , \3141_b1 );
not ( w_7357 , w_7360 );
not (  , w_7361 );
and ( w_7360 , w_7361 , \3141_b0 );
or ( \3143_b1 , \3142_b1 , w_7362 );
xor ( \3143_b0 , \3142_b0 , w_7364 );
not ( w_7364 , w_7365 );
and ( w_7365 , w_7362 , w_7363 );
buf ( w_7362 , \2124_b1 );
not ( w_7362 , w_7366 );
not ( w_7363 , w_7367 );
and ( w_7366 , w_7367 , \2124_b0 );
or ( \3144_b1 , \444_b1 , \1955_b1 );
not ( \1955_b1 , w_7368 );
and ( \3144_b0 , \444_b0 , w_7369 );
and ( w_7368 , w_7369 , \1955_b0 );
or ( \3145_b1 , \360_b1 , \1953_b1 );
not ( \1953_b1 , w_7370 );
and ( \3145_b0 , \360_b0 , w_7371 );
and ( w_7370 , w_7371 , \1953_b0 );
or ( \3146_b1 , \3144_b1 , w_7373 );
not ( w_7373 , w_7374 );
and ( \3146_b0 , \3144_b0 , w_7375 );
and ( w_7374 ,  , w_7375 );
buf ( w_7373 , \3145_b1 );
not ( w_7373 , w_7376 );
not (  , w_7377 );
and ( w_7376 , w_7377 , \3145_b0 );
or ( \3147_b1 , \3146_b1 , w_7378 );
xor ( \3147_b0 , \3146_b0 , w_7380 );
not ( w_7380 , w_7381 );
and ( w_7381 , w_7378 , w_7379 );
buf ( w_7378 , \1835_b1 );
not ( w_7378 , w_7382 );
not ( w_7379 , w_7383 );
and ( w_7382 , w_7383 , \1835_b0 );
or ( \3148_b1 , \3143_b1 , \3147_b1 );
not ( \3147_b1 , w_7384 );
and ( \3148_b0 , \3143_b0 , w_7385 );
and ( w_7384 , w_7385 , \3147_b0 );
or ( \3149_b1 , \593_b1 , \1742_b1 );
not ( \1742_b1 , w_7386 );
and ( \3149_b0 , \593_b0 , w_7387 );
and ( w_7386 , w_7387 , \1742_b0 );
or ( \3150_b1 , \495_b1 , \1740_b1 );
not ( \1740_b1 , w_7388 );
and ( \3150_b0 , \495_b0 , w_7389 );
and ( w_7388 , w_7389 , \1740_b0 );
or ( \3151_b1 , \3149_b1 , w_7391 );
not ( w_7391 , w_7392 );
and ( \3151_b0 , \3149_b0 , w_7393 );
and ( w_7392 ,  , w_7393 );
buf ( w_7391 , \3150_b1 );
not ( w_7391 , w_7394 );
not (  , w_7395 );
and ( w_7394 , w_7395 , \3150_b0 );
or ( \3152_b1 , \3151_b1 , w_7396 );
xor ( \3152_b0 , \3151_b0 , w_7398 );
not ( w_7398 , w_7399 );
and ( w_7399 , w_7396 , w_7397 );
buf ( w_7396 , \1610_b1 );
not ( w_7396 , w_7400 );
not ( w_7397 , w_7401 );
and ( w_7400 , w_7401 , \1610_b0 );
or ( \3153_b1 , \3147_b1 , \3152_b1 );
not ( \3152_b1 , w_7402 );
and ( \3153_b0 , \3147_b0 , w_7403 );
and ( w_7402 , w_7403 , \3152_b0 );
or ( \3154_b1 , \3143_b1 , \3152_b1 );
not ( \3152_b1 , w_7404 );
and ( \3154_b0 , \3143_b0 , w_7405 );
and ( w_7404 , w_7405 , \3152_b0 );
or ( \3156_b1 , \703_b1 , \1476_b1 );
not ( \1476_b1 , w_7406 );
and ( \3156_b0 , \703_b0 , w_7407 );
and ( w_7406 , w_7407 , \1476_b0 );
or ( \3157_b1 , \621_b1 , \1474_b1 );
not ( \1474_b1 , w_7408 );
and ( \3157_b0 , \621_b0 , w_7409 );
and ( w_7408 , w_7409 , \1474_b0 );
or ( \3158_b1 , \3156_b1 , w_7411 );
not ( w_7411 , w_7412 );
and ( \3158_b0 , \3156_b0 , w_7413 );
and ( w_7412 ,  , w_7413 );
buf ( w_7411 , \3157_b1 );
not ( w_7411 , w_7414 );
not (  , w_7415 );
and ( w_7414 , w_7415 , \3157_b0 );
or ( \3159_b1 , \3158_b1 , w_7416 );
xor ( \3159_b0 , \3158_b0 , w_7418 );
not ( w_7418 , w_7419 );
and ( w_7419 , w_7416 , w_7417 );
buf ( w_7416 , \1363_b1 );
not ( w_7416 , w_7420 );
not ( w_7417 , w_7421 );
and ( w_7420 , w_7421 , \1363_b0 );
or ( \3160_b1 , \841_b1 , \1280_b1 );
not ( \1280_b1 , w_7422 );
and ( \3160_b0 , \841_b0 , w_7423 );
and ( w_7422 , w_7423 , \1280_b0 );
or ( \3161_b1 , \777_b1 , \1278_b1 );
not ( \1278_b1 , w_7424 );
and ( \3161_b0 , \777_b0 , w_7425 );
and ( w_7424 , w_7425 , \1278_b0 );
or ( \3162_b1 , \3160_b1 , w_7427 );
not ( w_7427 , w_7428 );
and ( \3162_b0 , \3160_b0 , w_7429 );
and ( w_7428 ,  , w_7429 );
buf ( w_7427 , \3161_b1 );
not ( w_7427 , w_7430 );
not (  , w_7431 );
and ( w_7430 , w_7431 , \3161_b0 );
or ( \3163_b1 , \3162_b1 , w_7432 );
xor ( \3163_b0 , \3162_b0 , w_7434 );
not ( w_7434 , w_7435 );
and ( w_7435 , w_7432 , w_7433 );
buf ( w_7432 , \1177_b1 );
not ( w_7432 , w_7436 );
not ( w_7433 , w_7437 );
and ( w_7436 , w_7437 , \1177_b0 );
or ( \3164_b1 , \3159_b1 , \3163_b1 );
not ( \3163_b1 , w_7438 );
and ( \3164_b0 , \3159_b0 , w_7439 );
and ( w_7438 , w_7439 , \3163_b0 );
or ( \3165_b1 , \1104_b1 , \1062_b1 );
not ( \1062_b1 , w_7440 );
and ( \3165_b0 , \1104_b0 , w_7441 );
and ( w_7440 , w_7441 , \1062_b0 );
or ( \3166_b1 , \904_b1 , \1060_b1 );
not ( \1060_b1 , w_7442 );
and ( \3166_b0 , \904_b0 , w_7443 );
and ( w_7442 , w_7443 , \1060_b0 );
or ( \3167_b1 , \3165_b1 , w_7445 );
not ( w_7445 , w_7446 );
and ( \3167_b0 , \3165_b0 , w_7447 );
and ( w_7446 ,  , w_7447 );
buf ( w_7445 , \3166_b1 );
not ( w_7445 , w_7448 );
not (  , w_7449 );
and ( w_7448 , w_7449 , \3166_b0 );
or ( \3168_b1 , \3167_b1 , w_7450 );
xor ( \3168_b0 , \3167_b0 , w_7452 );
not ( w_7452 , w_7453 );
and ( w_7453 , w_7450 , w_7451 );
buf ( w_7450 , \984_b1 );
not ( w_7450 , w_7454 );
not ( w_7451 , w_7455 );
and ( w_7454 , w_7455 , \984_b0 );
or ( \3169_b1 , \3163_b1 , \3168_b1 );
not ( \3168_b1 , w_7456 );
and ( \3169_b0 , \3163_b0 , w_7457 );
and ( w_7456 , w_7457 , \3168_b0 );
or ( \3170_b1 , \3159_b1 , \3168_b1 );
not ( \3168_b1 , w_7458 );
and ( \3170_b0 , \3159_b0 , w_7459 );
and ( w_7458 , w_7459 , \3168_b0 );
or ( \3172_b1 , \3155_b1 , \3171_b1 );
not ( \3171_b1 , w_7460 );
and ( \3172_b0 , \3155_b0 , w_7461 );
and ( w_7460 , w_7461 , \3171_b0 );
or ( \3173_b1 , \305_b1 , \2913_b1 );
not ( \2913_b1 , w_7462 );
and ( \3173_b0 , \305_b0 , w_7463 );
and ( w_7462 , w_7463 , \2913_b0 );
or ( \3174_b1 , \315_b1 , \2910_b1 );
not ( \2910_b1 , w_7464 );
and ( \3174_b0 , \315_b0 , w_7465 );
and ( w_7464 , w_7465 , \2910_b0 );
or ( \3175_b1 , \3173_b1 , w_7467 );
not ( w_7467 , w_7468 );
and ( \3175_b0 , \3173_b0 , w_7469 );
and ( w_7468 ,  , w_7469 );
buf ( w_7467 , \3174_b1 );
not ( w_7467 , w_7470 );
not (  , w_7471 );
and ( w_7470 , w_7471 , \3174_b0 );
or ( \3176_b1 , \3175_b1 , w_7472 );
xor ( \3176_b0 , \3175_b0 , w_7474 );
not ( w_7474 , w_7475 );
and ( w_7475 , w_7472 , w_7473 );
buf ( w_7472 , \2371_b1 );
not ( w_7472 , w_7476 );
not ( w_7473 , w_7477 );
and ( w_7476 , w_7477 , \2371_b0 );
or ( \3177_b1 , \323_b1 , \2550_b1 );
not ( \2550_b1 , w_7478 );
and ( \3177_b0 , \323_b0 , w_7479 );
and ( w_7478 , w_7479 , \2550_b0 );
or ( \3178_b1 , \333_b1 , \2548_b1 );
not ( \2548_b1 , w_7480 );
and ( \3178_b0 , \333_b0 , w_7481 );
and ( w_7480 , w_7481 , \2548_b0 );
or ( \3179_b1 , \3177_b1 , w_7483 );
not ( w_7483 , w_7484 );
and ( \3179_b0 , \3177_b0 , w_7485 );
and ( w_7484 ,  , w_7485 );
buf ( w_7483 , \3178_b1 );
not ( w_7483 , w_7486 );
not (  , w_7487 );
and ( w_7486 , w_7487 , \3178_b0 );
or ( \3180_b1 , \3179_b1 , w_7488 );
xor ( \3180_b0 , \3179_b0 , w_7490 );
not ( w_7490 , w_7491 );
and ( w_7491 , w_7488 , w_7489 );
buf ( w_7488 , \2374_b1 );
not ( w_7488 , w_7492 );
not ( w_7489 , w_7493 );
and ( w_7492 , w_7493 , \2374_b0 );
or ( \3181_b1 , \3176_b1 , \3180_b1 );
not ( \3180_b1 , w_7494 );
and ( \3181_b0 , \3176_b0 , w_7495 );
and ( w_7494 , w_7495 , \3180_b0 );
or ( \3182_b1 , \3180_b1 , \358_b1 );
not ( \358_b1 , w_7496 );
and ( \3182_b0 , \3180_b0 , w_7497 );
and ( w_7496 , w_7497 , \358_b0 );
or ( \3183_b1 , \3176_b1 , \358_b1 );
not ( \358_b1 , w_7498 );
and ( \3183_b0 , \3176_b0 , w_7499 );
and ( w_7498 , w_7499 , \358_b0 );
or ( \3185_b1 , \3171_b1 , \3184_b1 );
not ( \3184_b1 , w_7500 );
and ( \3185_b0 , \3171_b0 , w_7501 );
and ( w_7500 , w_7501 , \3184_b0 );
or ( \3186_b1 , \3155_b1 , \3184_b1 );
not ( \3184_b1 , w_7502 );
and ( \3186_b0 , \3155_b0 , w_7503 );
and ( w_7502 , w_7503 , \3184_b0 );
or ( \3188_b1 , \2023_b1 , \503_b1 );
not ( \503_b1 , w_7504 );
and ( \3188_b0 , \2023_b0 , w_7505 );
and ( w_7504 , w_7505 , \503_b0 );
or ( \3189_b1 , \1778_b1 , \501_b1 );
not ( \501_b1 , w_7506 );
and ( \3189_b0 , \1778_b0 , w_7507 );
and ( w_7506 , w_7507 , \501_b0 );
or ( \3190_b1 , \3188_b1 , w_7509 );
not ( w_7509 , w_7510 );
and ( \3190_b0 , \3188_b0 , w_7511 );
and ( w_7510 ,  , w_7511 );
buf ( w_7509 , \3189_b1 );
not ( w_7509 , w_7512 );
not (  , w_7513 );
and ( w_7512 , w_7513 , \3189_b0 );
or ( \3191_b1 , \3190_b1 , w_7514 );
xor ( \3191_b0 , \3190_b0 , w_7516 );
not ( w_7516 , w_7517 );
and ( w_7517 , w_7514 , w_7515 );
buf ( w_7514 , \455_b1 );
not ( w_7514 , w_7518 );
not ( w_7515 , w_7519 );
and ( w_7518 , w_7519 , \455_b0 );
or ( \3192_b1 , \2161_b1 , \298_b1 );
not ( \298_b1 , w_7520 );
and ( \3192_b0 , \2161_b0 , w_7521 );
and ( w_7520 , w_7521 , \298_b0 );
or ( \3193_b1 , \2028_b1 , \296_b1 );
not ( \296_b1 , w_7522 );
and ( \3193_b0 , \2028_b0 , w_7523 );
and ( w_7522 , w_7523 , \296_b0 );
or ( \3194_b1 , \3192_b1 , w_7525 );
not ( w_7525 , w_7526 );
and ( \3194_b0 , \3192_b0 , w_7527 );
and ( w_7526 ,  , w_7527 );
buf ( w_7525 , \3193_b1 );
not ( w_7525 , w_7528 );
not (  , w_7529 );
and ( w_7528 , w_7529 , \3193_b0 );
or ( \3195_b1 , \3194_b1 , w_7530 );
xor ( \3195_b0 , \3194_b0 , w_7532 );
not ( w_7532 , w_7533 );
and ( w_7533 , w_7530 , w_7531 );
buf ( w_7530 , \303_b1 );
not ( w_7530 , w_7534 );
not ( w_7531 , w_7535 );
and ( w_7534 , w_7535 , \303_b0 );
or ( \3196_b1 , \3191_b1 , \3195_b1 );
not ( \3195_b1 , w_7536 );
and ( \3196_b0 , \3191_b0 , w_7537 );
and ( w_7536 , w_7537 , \3195_b0 );
or ( \3197_b1 , \2532_b1 , \313_b1 );
not ( \313_b1 , w_7538 );
and ( \3197_b0 , \2532_b0 , w_7539 );
and ( w_7538 , w_7539 , \313_b0 );
or ( \3198_b1 , \2305_b1 , \311_b1 );
not ( \311_b1 , w_7540 );
and ( \3198_b0 , \2305_b0 , w_7541 );
and ( w_7540 , w_7541 , \311_b0 );
or ( \3199_b1 , \3197_b1 , w_7543 );
not ( w_7543 , w_7544 );
and ( \3199_b0 , \3197_b0 , w_7545 );
and ( w_7544 ,  , w_7545 );
buf ( w_7543 , \3198_b1 );
not ( w_7543 , w_7546 );
not (  , w_7547 );
and ( w_7546 , w_7547 , \3198_b0 );
or ( \3200_b1 , \3199_b1 , w_7548 );
xor ( \3200_b0 , \3199_b0 , w_7550 );
not ( w_7550 , w_7551 );
and ( w_7551 , w_7548 , w_7549 );
buf ( w_7548 , \320_b1 );
not ( w_7548 , w_7552 );
not ( w_7549 , w_7553 );
and ( w_7552 , w_7553 , \320_b0 );
or ( \3201_b1 , \3195_b1 , \3200_b1 );
not ( \3200_b1 , w_7554 );
and ( \3201_b0 , \3195_b0 , w_7555 );
and ( w_7554 , w_7555 , \3200_b0 );
or ( \3202_b1 , \3191_b1 , \3200_b1 );
not ( \3200_b1 , w_7556 );
and ( \3202_b0 , \3191_b0 , w_7557 );
and ( w_7556 , w_7557 , \3200_b0 );
or ( \3204_b1 , \1299_b1 , \912_b1 );
not ( \912_b1 , w_7558 );
and ( \3204_b0 , \1299_b0 , w_7559 );
and ( w_7558 , w_7559 , \912_b0 );
or ( \3205_b1 , \1194_b1 , \910_b1 );
not ( \910_b1 , w_7560 );
and ( \3205_b0 , \1194_b0 , w_7561 );
and ( w_7560 , w_7561 , \910_b0 );
or ( \3206_b1 , \3204_b1 , w_7563 );
not ( w_7563 , w_7564 );
and ( \3206_b0 , \3204_b0 , w_7565 );
and ( w_7564 ,  , w_7565 );
buf ( w_7563 , \3205_b1 );
not ( w_7563 , w_7566 );
not (  , w_7567 );
and ( w_7566 , w_7567 , \3205_b0 );
or ( \3207_b1 , \3206_b1 , w_7568 );
xor ( \3207_b0 , \3206_b0 , w_7570 );
not ( w_7570 , w_7571 );
and ( w_7571 , w_7568 , w_7569 );
buf ( w_7568 , \818_b1 );
not ( w_7568 , w_7572 );
not ( w_7569 , w_7573 );
and ( w_7572 , w_7573 , \818_b0 );
or ( \3208_b1 , \1422_b1 , \740_b1 );
not ( \740_b1 , w_7574 );
and ( \3208_b0 , \1422_b0 , w_7575 );
and ( w_7574 , w_7575 , \740_b0 );
or ( \3209_b1 , \1304_b1 , \738_b1 );
not ( \738_b1 , w_7576 );
and ( \3209_b0 , \1304_b0 , w_7577 );
and ( w_7576 , w_7577 , \738_b0 );
or ( \3210_b1 , \3208_b1 , w_7579 );
not ( w_7579 , w_7580 );
and ( \3210_b0 , \3208_b0 , w_7581 );
and ( w_7580 ,  , w_7581 );
buf ( w_7579 , \3209_b1 );
not ( w_7579 , w_7582 );
not (  , w_7583 );
and ( w_7582 , w_7583 , \3209_b0 );
or ( \3211_b1 , \3210_b1 , w_7584 );
xor ( \3211_b0 , \3210_b0 , w_7586 );
not ( w_7586 , w_7587 );
and ( w_7587 , w_7584 , w_7585 );
buf ( w_7584 , \668_b1 );
not ( w_7584 , w_7588 );
not ( w_7585 , w_7589 );
and ( w_7588 , w_7589 , \668_b0 );
or ( \3212_b1 , \3207_b1 , \3211_b1 );
not ( \3211_b1 , w_7590 );
and ( \3212_b0 , \3207_b0 , w_7591 );
and ( w_7590 , w_7591 , \3211_b0 );
or ( \3213_b1 , \1770_b1 , \604_b1 );
not ( \604_b1 , w_7592 );
and ( \3213_b0 , \1770_b0 , w_7593 );
and ( w_7592 , w_7593 , \604_b0 );
or ( \3214_b1 , \1537_b1 , \602_b1 );
not ( \602_b1 , w_7594 );
and ( \3214_b0 , \1537_b0 , w_7595 );
and ( w_7594 , w_7595 , \602_b0 );
or ( \3215_b1 , \3213_b1 , w_7597 );
not ( w_7597 , w_7598 );
and ( \3215_b0 , \3213_b0 , w_7599 );
and ( w_7598 ,  , w_7599 );
buf ( w_7597 , \3214_b1 );
not ( w_7597 , w_7600 );
not (  , w_7601 );
and ( w_7600 , w_7601 , \3214_b0 );
or ( \3216_b1 , \3215_b1 , w_7602 );
xor ( \3216_b0 , \3215_b0 , w_7604 );
not ( w_7604 , w_7605 );
and ( w_7605 , w_7602 , w_7603 );
buf ( w_7602 , \561_b1 );
not ( w_7602 , w_7606 );
not ( w_7603 , w_7607 );
and ( w_7606 , w_7607 , \561_b0 );
or ( \3217_b1 , \3211_b1 , \3216_b1 );
not ( \3216_b1 , w_7608 );
and ( \3217_b0 , \3211_b0 , w_7609 );
and ( w_7608 , w_7609 , \3216_b0 );
or ( \3218_b1 , \3207_b1 , \3216_b1 );
not ( \3216_b1 , w_7610 );
and ( \3218_b0 , \3207_b0 , w_7611 );
and ( w_7610 , w_7611 , \3216_b0 );
or ( \3220_b1 , \3203_b1 , \3219_b1 );
not ( \3219_b1 , w_7612 );
and ( \3220_b0 , \3203_b0 , w_7613 );
and ( w_7612 , w_7613 , \3219_b0 );
or ( \3221_b1 , \2850_b1 , \351_b1 );
not ( \351_b1 , w_7614 );
and ( \3221_b0 , \2850_b0 , w_7615 );
and ( w_7614 , w_7615 , \351_b0 );
or ( \3222_b1 , \2763_b1 , \349_b1 );
not ( \349_b1 , w_7616 );
and ( \3222_b0 , \2763_b0 , w_7617 );
and ( w_7616 , w_7617 , \349_b0 );
or ( \3223_b1 , \3221_b1 , w_7619 );
not ( w_7619 , w_7620 );
and ( \3223_b0 , \3221_b0 , w_7621 );
and ( w_7620 ,  , w_7621 );
buf ( w_7619 , \3222_b1 );
not ( w_7619 , w_7622 );
not (  , w_7623 );
and ( w_7622 , w_7623 , \3222_b0 );
or ( \3224_b1 , \3223_b1 , w_7624 );
xor ( \3224_b0 , \3223_b0 , w_7626 );
not ( w_7626 , w_7627 );
and ( w_7627 , w_7624 , w_7625 );
buf ( w_7624 , \358_b1 );
not ( w_7624 , w_7628 );
not ( w_7625 , w_7629 );
and ( w_7628 , w_7629 , \358_b0 );
or ( \3225_b1 , \3219_b1 , \3224_b1 );
not ( \3224_b1 , w_7630 );
and ( \3225_b0 , \3219_b0 , w_7631 );
and ( w_7630 , w_7631 , \3224_b0 );
or ( \3226_b1 , \3203_b1 , \3224_b1 );
not ( \3224_b1 , w_7632 );
and ( \3226_b0 , \3203_b0 , w_7633 );
and ( w_7632 , w_7633 , \3224_b0 );
or ( \3228_b1 , \3187_b1 , \3227_b1 );
not ( \3227_b1 , w_7634 );
and ( \3228_b0 , \3187_b0 , w_7635 );
and ( w_7634 , w_7635 , \3227_b0 );
or ( \3229_b1 , \3059_b1 , \3063_b1 );
xor ( \3229_b0 , \3059_b0 , w_7636 );
not ( w_7636 , w_7637 );
and ( w_7637 , \3063_b1 , \3063_b0 );
or ( \3230_b1 , \3229_b1 , \3068_b1 );
xor ( \3230_b0 , \3229_b0 , w_7638 );
not ( w_7638 , w_7639 );
and ( w_7639 , \3068_b1 , \3068_b0 );
or ( \3231_b1 , \3075_b1 , \3079_b1 );
xor ( \3231_b0 , \3075_b0 , w_7640 );
not ( w_7640 , w_7641 );
and ( w_7641 , \3079_b1 , \3079_b0 );
or ( \3232_b1 , \3231_b1 , \3084_b1 );
xor ( \3232_b0 , \3231_b0 , w_7642 );
not ( w_7642 , w_7643 );
and ( w_7643 , \3084_b1 , \3084_b0 );
or ( \3233_b1 , \3230_b1 , \3232_b1 );
not ( \3232_b1 , w_7644 );
and ( \3233_b0 , \3230_b0 , w_7645 );
and ( w_7644 , w_7645 , \3232_b0 );
or ( \3234_b1 , \3029_b1 , \3033_b1 );
xor ( \3234_b0 , \3029_b0 , w_7646 );
not ( w_7646 , w_7647 );
and ( w_7647 , \3033_b1 , \3033_b0 );
or ( \3235_b1 , \3234_b1 , \3038_b1 );
xor ( \3235_b0 , \3234_b0 , w_7648 );
not ( w_7648 , w_7649 );
and ( w_7649 , \3038_b1 , \3038_b0 );
or ( \3236_b1 , \3232_b1 , \3235_b1 );
not ( \3235_b1 , w_7650 );
and ( \3236_b0 , \3232_b0 , w_7651 );
and ( w_7650 , w_7651 , \3235_b0 );
or ( \3237_b1 , \3230_b1 , \3235_b1 );
not ( \3235_b1 , w_7652 );
and ( \3237_b0 , \3230_b0 , w_7653 );
and ( w_7652 , w_7653 , \3235_b0 );
or ( \3239_b1 , \3227_b1 , \3238_b1 );
not ( \3238_b1 , w_7654 );
and ( \3239_b0 , \3227_b0 , w_7655 );
and ( w_7654 , w_7655 , \3238_b0 );
or ( \3240_b1 , \3187_b1 , \3238_b1 );
not ( \3238_b1 , w_7656 );
and ( \3240_b0 , \3187_b0 , w_7657 );
and ( w_7656 , w_7657 , \3238_b0 );
or ( \3242_b1 , \2895_b1 , \2899_b1 );
xor ( \3242_b0 , \2895_b0 , w_7658 );
not ( w_7658 , w_7659 );
and ( w_7659 , \2899_b1 , \2899_b0 );
or ( \3243_b1 , \3242_b1 , \2904_b1 );
xor ( \3243_b0 , \3242_b0 , w_7660 );
not ( w_7660 , w_7661 );
and ( w_7661 , \2904_b1 , \2904_b0 );
or ( \3244_b1 , \3046_b1 , \3048_b1 );
xor ( \3244_b0 , \3046_b0 , w_7662 );
not ( w_7662 , w_7663 );
and ( w_7663 , \3048_b1 , \3048_b0 );
or ( \3245_b1 , \3244_b1 , \3051_b1 );
xor ( \3245_b0 , \3244_b0 , w_7664 );
not ( w_7664 , w_7665 );
and ( w_7665 , \3051_b1 , \3051_b0 );
or ( \3246_b1 , \3243_b1 , \3245_b1 );
not ( \3245_b1 , w_7666 );
and ( \3246_b0 , \3243_b0 , w_7667 );
and ( w_7666 , w_7667 , \3245_b0 );
or ( \3247_b1 , \2916_b1 , \2920_b1 );
xor ( \3247_b0 , \2916_b0 , w_7668 );
not ( w_7668 , w_7669 );
and ( w_7669 , \2920_b1 , \2920_b0 );
or ( \3248_b1 , \3245_b1 , \3247_b1 );
not ( \3247_b1 , w_7670 );
and ( \3248_b0 , \3245_b0 , w_7671 );
and ( w_7670 , w_7671 , \3247_b0 );
or ( \3249_b1 , \3243_b1 , \3247_b1 );
not ( \3247_b1 , w_7672 );
and ( \3249_b0 , \3243_b0 , w_7673 );
and ( w_7672 , w_7673 , \3247_b0 );
or ( \3251_b1 , \3241_b1 , \3250_b1 );
not ( \3250_b1 , w_7674 );
and ( \3251_b0 , \3241_b0 , w_7675 );
and ( w_7674 , w_7675 , \3250_b0 );
or ( \3252_b1 , \3008_b1 , \3024_b1 );
xor ( \3252_b0 , \3008_b0 , w_7676 );
not ( w_7676 , w_7677 );
and ( w_7677 , \3024_b1 , \3024_b0 );
or ( \3253_b1 , \3252_b1 , \3041_b1 );
xor ( \3253_b0 , \3252_b0 , w_7678 );
not ( w_7678 , w_7679 );
and ( w_7679 , \3041_b1 , \3041_b0 );
or ( \3254_b1 , \3071_b1 , \3087_b1 );
xor ( \3254_b0 , \3071_b0 , w_7680 );
not ( w_7680 , w_7681 );
and ( w_7681 , \3087_b1 , \3087_b0 );
or ( \3255_b1 , \3254_b1 , \3090_b1 );
xor ( \3255_b0 , \3254_b0 , w_7682 );
not ( w_7682 , w_7683 );
and ( w_7683 , \3090_b1 , \3090_b0 );
or ( \3256_b1 , \3253_b1 , \3255_b1 );
not ( \3255_b1 , w_7684 );
and ( \3256_b0 , \3253_b0 , w_7685 );
and ( w_7684 , w_7685 , \3255_b0 );
or ( \3257_b1 , \3250_b1 , \3256_b1 );
not ( \3256_b1 , w_7686 );
and ( \3257_b0 , \3250_b0 , w_7687 );
and ( w_7686 , w_7687 , \3256_b0 );
or ( \3258_b1 , \3241_b1 , \3256_b1 );
not ( \3256_b1 , w_7688 );
and ( \3258_b0 , \3241_b0 , w_7689 );
and ( w_7688 , w_7689 , \3256_b0 );
or ( \3260_b1 , \2891_b1 , \2907_b1 );
xor ( \3260_b0 , \2891_b0 , w_7690 );
not ( w_7690 , w_7691 );
and ( w_7691 , \2907_b1 , \2907_b0 );
or ( \3261_b1 , \3260_b1 , \2921_b1 );
xor ( \3261_b0 , \3260_b0 , w_7692 );
not ( w_7692 , w_7693 );
and ( w_7693 , \2921_b1 , \2921_b0 );
or ( \3262_b1 , \3044_b1 , \3054_b1 );
xor ( \3262_b0 , \3044_b0 , w_7694 );
not ( w_7694 , w_7695 );
and ( w_7695 , \3054_b1 , \3054_b0 );
or ( \3263_b1 , \3262_b1 , \3093_b1 );
xor ( \3263_b0 , \3262_b0 , w_7696 );
not ( w_7696 , w_7697 );
and ( w_7697 , \3093_b1 , \3093_b0 );
or ( \3264_b1 , \3261_b1 , \3263_b1 );
not ( \3263_b1 , w_7698 );
and ( \3264_b0 , \3261_b0 , w_7699 );
and ( w_7698 , w_7699 , \3263_b0 );
or ( \3265_b1 , \3098_b1 , \3100_b1 );
xor ( \3265_b0 , \3098_b0 , w_7700 );
not ( w_7700 , w_7701 );
and ( w_7701 , \3100_b1 , \3100_b0 );
or ( \3266_b1 , \3265_b1 , \3103_b1 );
xor ( \3266_b0 , \3265_b0 , w_7702 );
not ( w_7702 , w_7703 );
and ( w_7703 , \3103_b1 , \3103_b0 );
or ( \3267_b1 , \3263_b1 , \3266_b1 );
not ( \3266_b1 , w_7704 );
and ( \3267_b0 , \3263_b0 , w_7705 );
and ( w_7704 , w_7705 , \3266_b0 );
or ( \3268_b1 , \3261_b1 , \3266_b1 );
not ( \3266_b1 , w_7706 );
and ( \3268_b0 , \3261_b0 , w_7707 );
and ( w_7706 , w_7707 , \3266_b0 );
or ( \3270_b1 , \3259_b1 , \3269_b1 );
not ( \3269_b1 , w_7708 );
and ( \3270_b0 , \3259_b0 , w_7709 );
and ( w_7708 , w_7709 , \3269_b0 );
or ( \3271_b1 , \3114_b1 , \3116_b1 );
xor ( \3271_b0 , \3114_b0 , w_7710 );
not ( w_7710 , w_7711 );
and ( w_7711 , \3116_b1 , \3116_b0 );
or ( \3272_b1 , \3271_b1 , \3119_b1 );
xor ( \3272_b0 , \3271_b0 , w_7712 );
not ( w_7712 , w_7713 );
and ( w_7713 , \3119_b1 , \3119_b0 );
or ( \3273_b1 , \3269_b1 , \3272_b1 );
not ( \3272_b1 , w_7714 );
and ( \3273_b0 , \3269_b0 , w_7715 );
and ( w_7714 , w_7715 , \3272_b0 );
or ( \3274_b1 , \3259_b1 , \3272_b1 );
not ( \3272_b1 , w_7716 );
and ( \3274_b0 , \3259_b0 , w_7717 );
and ( w_7716 , w_7717 , \3272_b0 );
or ( \3276_b1 , \2937_b1 , \2955_b1 );
xor ( \3276_b0 , \2937_b0 , w_7718 );
not ( w_7718 , w_7719 );
and ( w_7719 , \2955_b1 , \2955_b0 );
or ( \3277_b1 , \3276_b1 , \2958_b1 );
xor ( \3277_b0 , \3276_b0 , w_7720 );
not ( w_7720 , w_7721 );
and ( w_7721 , \2958_b1 , \2958_b0 );
or ( \3278_b1 , \3275_b1 , \3277_b1 );
not ( \3277_b1 , w_7722 );
and ( \3278_b0 , \3275_b0 , w_7723 );
and ( w_7722 , w_7723 , \3277_b0 );
or ( \3279_b1 , \3112_b1 , \3122_b1 );
xor ( \3279_b0 , \3112_b0 , w_7724 );
not ( w_7724 , w_7725 );
and ( w_7725 , \3122_b1 , \3122_b0 );
or ( \3280_b1 , \3279_b1 , \3125_b1 );
xor ( \3280_b0 , \3279_b0 , w_7726 );
not ( w_7726 , w_7727 );
and ( w_7727 , \3125_b1 , \3125_b0 );
or ( \3281_b1 , \3277_b1 , \3280_b1 );
not ( \3280_b1 , w_7728 );
and ( \3281_b0 , \3277_b0 , w_7729 );
and ( w_7728 , w_7729 , \3280_b0 );
or ( \3282_b1 , \3275_b1 , \3280_b1 );
not ( \3280_b1 , w_7730 );
and ( \3282_b0 , \3275_b0 , w_7731 );
and ( w_7730 , w_7731 , \3280_b0 );
or ( \3284_b1 , \3139_b1 , \3283_b1 );
not ( \3283_b1 , w_7732 );
and ( \3284_b0 , \3139_b0 , w_7733 );
and ( w_7732 , w_7733 , \3283_b0 );
or ( \3285_b1 , \3139_b1 , \3283_b1 );
xor ( \3285_b0 , \3139_b0 , w_7734 );
not ( w_7734 , w_7735 );
and ( w_7735 , \3283_b1 , \3283_b0 );
or ( \3286_b1 , \3275_b1 , \3277_b1 );
xor ( \3286_b0 , \3275_b0 , w_7736 );
not ( w_7736 , w_7737 );
and ( w_7737 , \3277_b1 , \3277_b0 );
or ( \3287_b1 , \3286_b1 , \3280_b1 );
xor ( \3287_b0 , \3286_b0 , w_7738 );
not ( w_7738 , w_7739 );
and ( w_7739 , \3280_b1 , \3280_b0 );
or ( \3288_b1 , \904_b1 , \1280_b1 );
not ( \1280_b1 , w_7740 );
and ( \3288_b0 , \904_b0 , w_7741 );
and ( w_7740 , w_7741 , \1280_b0 );
or ( \3289_b1 , \841_b1 , \1278_b1 );
not ( \1278_b1 , w_7742 );
and ( \3289_b0 , \841_b0 , w_7743 );
and ( w_7742 , w_7743 , \1278_b0 );
or ( \3290_b1 , \3288_b1 , w_7745 );
not ( w_7745 , w_7746 );
and ( \3290_b0 , \3288_b0 , w_7747 );
and ( w_7746 ,  , w_7747 );
buf ( w_7745 , \3289_b1 );
not ( w_7745 , w_7748 );
not (  , w_7749 );
and ( w_7748 , w_7749 , \3289_b0 );
or ( \3291_b1 , \3290_b1 , w_7750 );
xor ( \3291_b0 , \3290_b0 , w_7752 );
not ( w_7752 , w_7753 );
and ( w_7753 , w_7750 , w_7751 );
buf ( w_7750 , \1177_b1 );
not ( w_7750 , w_7754 );
not ( w_7751 , w_7755 );
and ( w_7754 , w_7755 , \1177_b0 );
or ( \3292_b1 , \1194_b1 , \1062_b1 );
not ( \1062_b1 , w_7756 );
and ( \3292_b0 , \1194_b0 , w_7757 );
and ( w_7756 , w_7757 , \1062_b0 );
or ( \3293_b1 , \1104_b1 , \1060_b1 );
not ( \1060_b1 , w_7758 );
and ( \3293_b0 , \1104_b0 , w_7759 );
and ( w_7758 , w_7759 , \1060_b0 );
or ( \3294_b1 , \3292_b1 , w_7761 );
not ( w_7761 , w_7762 );
and ( \3294_b0 , \3292_b0 , w_7763 );
and ( w_7762 ,  , w_7763 );
buf ( w_7761 , \3293_b1 );
not ( w_7761 , w_7764 );
not (  , w_7765 );
and ( w_7764 , w_7765 , \3293_b0 );
or ( \3295_b1 , \3294_b1 , w_7766 );
xor ( \3295_b0 , \3294_b0 , w_7768 );
not ( w_7768 , w_7769 );
and ( w_7769 , w_7766 , w_7767 );
buf ( w_7766 , \984_b1 );
not ( w_7766 , w_7770 );
not ( w_7767 , w_7771 );
and ( w_7770 , w_7771 , \984_b0 );
or ( \3296_b1 , \3291_b1 , \3295_b1 );
not ( \3295_b1 , w_7772 );
and ( \3296_b0 , \3291_b0 , w_7773 );
and ( w_7772 , w_7773 , \3295_b0 );
or ( \3297_b1 , \1304_b1 , \912_b1 );
not ( \912_b1 , w_7774 );
and ( \3297_b0 , \1304_b0 , w_7775 );
and ( w_7774 , w_7775 , \912_b0 );
or ( \3298_b1 , \1299_b1 , \910_b1 );
not ( \910_b1 , w_7776 );
and ( \3298_b0 , \1299_b0 , w_7777 );
and ( w_7776 , w_7777 , \910_b0 );
or ( \3299_b1 , \3297_b1 , w_7779 );
not ( w_7779 , w_7780 );
and ( \3299_b0 , \3297_b0 , w_7781 );
and ( w_7780 ,  , w_7781 );
buf ( w_7779 , \3298_b1 );
not ( w_7779 , w_7782 );
not (  , w_7783 );
and ( w_7782 , w_7783 , \3298_b0 );
or ( \3300_b1 , \3299_b1 , w_7784 );
xor ( \3300_b0 , \3299_b0 , w_7786 );
not ( w_7786 , w_7787 );
and ( w_7787 , w_7784 , w_7785 );
buf ( w_7784 , \818_b1 );
not ( w_7784 , w_7788 );
not ( w_7785 , w_7789 );
and ( w_7788 , w_7789 , \818_b0 );
or ( \3301_b1 , \3295_b1 , \3300_b1 );
not ( \3300_b1 , w_7790 );
and ( \3301_b0 , \3295_b0 , w_7791 );
and ( w_7790 , w_7791 , \3300_b0 );
or ( \3302_b1 , \3291_b1 , \3300_b1 );
not ( \3300_b1 , w_7792 );
and ( \3302_b0 , \3291_b0 , w_7793 );
and ( w_7792 , w_7793 , \3300_b0 );
or ( \3304_b1 , \495_b1 , \1955_b1 );
not ( \1955_b1 , w_7794 );
and ( \3304_b0 , \495_b0 , w_7795 );
and ( w_7794 , w_7795 , \1955_b0 );
or ( \3305_b1 , \444_b1 , \1953_b1 );
not ( \1953_b1 , w_7796 );
and ( \3305_b0 , \444_b0 , w_7797 );
and ( w_7796 , w_7797 , \1953_b0 );
or ( \3306_b1 , \3304_b1 , w_7799 );
not ( w_7799 , w_7800 );
and ( \3306_b0 , \3304_b0 , w_7801 );
and ( w_7800 ,  , w_7801 );
buf ( w_7799 , \3305_b1 );
not ( w_7799 , w_7802 );
not (  , w_7803 );
and ( w_7802 , w_7803 , \3305_b0 );
or ( \3307_b1 , \3306_b1 , w_7804 );
xor ( \3307_b0 , \3306_b0 , w_7806 );
not ( w_7806 , w_7807 );
and ( w_7807 , w_7804 , w_7805 );
buf ( w_7804 , \1835_b1 );
not ( w_7804 , w_7808 );
not ( w_7805 , w_7809 );
and ( w_7808 , w_7809 , \1835_b0 );
or ( \3308_b1 , \621_b1 , \1742_b1 );
not ( \1742_b1 , w_7810 );
and ( \3308_b0 , \621_b0 , w_7811 );
and ( w_7810 , w_7811 , \1742_b0 );
or ( \3309_b1 , \593_b1 , \1740_b1 );
not ( \1740_b1 , w_7812 );
and ( \3309_b0 , \593_b0 , w_7813 );
and ( w_7812 , w_7813 , \1740_b0 );
or ( \3310_b1 , \3308_b1 , w_7815 );
not ( w_7815 , w_7816 );
and ( \3310_b0 , \3308_b0 , w_7817 );
and ( w_7816 ,  , w_7817 );
buf ( w_7815 , \3309_b1 );
not ( w_7815 , w_7818 );
not (  , w_7819 );
and ( w_7818 , w_7819 , \3309_b0 );
or ( \3311_b1 , \3310_b1 , w_7820 );
xor ( \3311_b0 , \3310_b0 , w_7822 );
not ( w_7822 , w_7823 );
and ( w_7823 , w_7820 , w_7821 );
buf ( w_7820 , \1610_b1 );
not ( w_7820 , w_7824 );
not ( w_7821 , w_7825 );
and ( w_7824 , w_7825 , \1610_b0 );
or ( \3312_b1 , \3307_b1 , \3311_b1 );
not ( \3311_b1 , w_7826 );
and ( \3312_b0 , \3307_b0 , w_7827 );
and ( w_7826 , w_7827 , \3311_b0 );
or ( \3313_b1 , \777_b1 , \1476_b1 );
not ( \1476_b1 , w_7828 );
and ( \3313_b0 , \777_b0 , w_7829 );
and ( w_7828 , w_7829 , \1476_b0 );
or ( \3314_b1 , \703_b1 , \1474_b1 );
not ( \1474_b1 , w_7830 );
and ( \3314_b0 , \703_b0 , w_7831 );
and ( w_7830 , w_7831 , \1474_b0 );
or ( \3315_b1 , \3313_b1 , w_7833 );
not ( w_7833 , w_7834 );
and ( \3315_b0 , \3313_b0 , w_7835 );
and ( w_7834 ,  , w_7835 );
buf ( w_7833 , \3314_b1 );
not ( w_7833 , w_7836 );
not (  , w_7837 );
and ( w_7836 , w_7837 , \3314_b0 );
or ( \3316_b1 , \3315_b1 , w_7838 );
xor ( \3316_b0 , \3315_b0 , w_7840 );
not ( w_7840 , w_7841 );
and ( w_7841 , w_7838 , w_7839 );
buf ( w_7838 , \1363_b1 );
not ( w_7838 , w_7842 );
not ( w_7839 , w_7843 );
and ( w_7842 , w_7843 , \1363_b0 );
or ( \3317_b1 , \3311_b1 , \3316_b1 );
not ( \3316_b1 , w_7844 );
and ( \3317_b0 , \3311_b0 , w_7845 );
and ( w_7844 , w_7845 , \3316_b0 );
or ( \3318_b1 , \3307_b1 , \3316_b1 );
not ( \3316_b1 , w_7846 );
and ( \3318_b0 , \3307_b0 , w_7847 );
and ( w_7846 , w_7847 , \3316_b0 );
or ( \3320_b1 , \3303_b1 , \3319_b1 );
not ( \3319_b1 , w_7848 );
and ( \3320_b0 , \3303_b0 , w_7849 );
and ( w_7848 , w_7849 , \3319_b0 );
or ( \3321_b1 , \333_b1 , \2913_b1 );
not ( \2913_b1 , w_7850 );
and ( \3321_b0 , \333_b0 , w_7851 );
and ( w_7850 , w_7851 , \2913_b0 );
or ( \3322_b1 , \305_b1 , \2910_b1 );
not ( \2910_b1 , w_7852 );
and ( \3322_b0 , \305_b0 , w_7853 );
and ( w_7852 , w_7853 , \2910_b0 );
or ( \3323_b1 , \3321_b1 , w_7855 );
not ( w_7855 , w_7856 );
and ( \3323_b0 , \3321_b0 , w_7857 );
and ( w_7856 ,  , w_7857 );
buf ( w_7855 , \3322_b1 );
not ( w_7855 , w_7858 );
not (  , w_7859 );
and ( w_7858 , w_7859 , \3322_b0 );
or ( \3324_b1 , \3323_b1 , w_7860 );
xor ( \3324_b0 , \3323_b0 , w_7862 );
not ( w_7862 , w_7863 );
and ( w_7863 , w_7860 , w_7861 );
buf ( w_7860 , \2371_b1 );
not ( w_7860 , w_7864 );
not ( w_7861 , w_7865 );
and ( w_7864 , w_7865 , \2371_b0 );
or ( \3325_b1 , \353_b1 , \2550_b1 );
not ( \2550_b1 , w_7866 );
and ( \3325_b0 , \353_b0 , w_7867 );
and ( w_7866 , w_7867 , \2550_b0 );
or ( \3326_b1 , \323_b1 , \2548_b1 );
not ( \2548_b1 , w_7868 );
and ( \3326_b0 , \323_b0 , w_7869 );
and ( w_7868 , w_7869 , \2548_b0 );
or ( \3327_b1 , \3325_b1 , w_7871 );
not ( w_7871 , w_7872 );
and ( \3327_b0 , \3325_b0 , w_7873 );
and ( w_7872 ,  , w_7873 );
buf ( w_7871 , \3326_b1 );
not ( w_7871 , w_7874 );
not (  , w_7875 );
and ( w_7874 , w_7875 , \3326_b0 );
or ( \3328_b1 , \3327_b1 , w_7876 );
xor ( \3328_b0 , \3327_b0 , w_7878 );
not ( w_7878 , w_7879 );
and ( w_7879 , w_7876 , w_7877 );
buf ( w_7876 , \2374_b1 );
not ( w_7876 , w_7880 );
not ( w_7877 , w_7881 );
and ( w_7880 , w_7881 , \2374_b0 );
or ( \3329_b1 , \3324_b1 , \3328_b1 );
not ( \3328_b1 , w_7882 );
and ( \3329_b0 , \3324_b0 , w_7883 );
and ( w_7882 , w_7883 , \3328_b0 );
or ( \3330_b1 , \360_b1 , \2261_b1 );
not ( \2261_b1 , w_7884 );
and ( \3330_b0 , \360_b0 , w_7885 );
and ( w_7884 , w_7885 , \2261_b0 );
or ( \3331_b1 , \343_b1 , \2259_b1 );
not ( \2259_b1 , w_7886 );
and ( \3331_b0 , \343_b0 , w_7887 );
and ( w_7886 , w_7887 , \2259_b0 );
or ( \3332_b1 , \3330_b1 , w_7889 );
not ( w_7889 , w_7890 );
and ( \3332_b0 , \3330_b0 , w_7891 );
and ( w_7890 ,  , w_7891 );
buf ( w_7889 , \3331_b1 );
not ( w_7889 , w_7892 );
not (  , w_7893 );
and ( w_7892 , w_7893 , \3331_b0 );
or ( \3333_b1 , \3332_b1 , w_7894 );
xor ( \3333_b0 , \3332_b0 , w_7896 );
not ( w_7896 , w_7897 );
and ( w_7897 , w_7894 , w_7895 );
buf ( w_7894 , \2124_b1 );
not ( w_7894 , w_7898 );
not ( w_7895 , w_7899 );
and ( w_7898 , w_7899 , \2124_b0 );
or ( \3334_b1 , \3328_b1 , \3333_b1 );
not ( \3333_b1 , w_7900 );
and ( \3334_b0 , \3328_b0 , w_7901 );
and ( w_7900 , w_7901 , \3333_b0 );
or ( \3335_b1 , \3324_b1 , \3333_b1 );
not ( \3333_b1 , w_7902 );
and ( \3335_b0 , \3324_b0 , w_7903 );
and ( w_7902 , w_7903 , \3333_b0 );
or ( \3337_b1 , \3319_b1 , \3336_b1 );
not ( \3336_b1 , w_7904 );
and ( \3337_b0 , \3319_b0 , w_7905 );
and ( w_7904 , w_7905 , \3336_b0 );
or ( \3338_b1 , \3303_b1 , \3336_b1 );
not ( \3336_b1 , w_7906 );
and ( \3338_b0 , \3303_b0 , w_7907 );
and ( w_7906 , w_7907 , \3336_b0 );
or ( \3340_b1 , \2305_b1 , \298_b1 );
not ( \298_b1 , w_7908 );
and ( \3340_b0 , \2305_b0 , w_7909 );
and ( w_7908 , w_7909 , \298_b0 );
or ( \3341_b1 , \2161_b1 , \296_b1 );
not ( \296_b1 , w_7910 );
and ( \3341_b0 , \2161_b0 , w_7911 );
and ( w_7910 , w_7911 , \296_b0 );
or ( \3342_b1 , \3340_b1 , w_7913 );
not ( w_7913 , w_7914 );
and ( \3342_b0 , \3340_b0 , w_7915 );
and ( w_7914 ,  , w_7915 );
buf ( w_7913 , \3341_b1 );
not ( w_7913 , w_7916 );
not (  , w_7917 );
and ( w_7916 , w_7917 , \3341_b0 );
or ( \3343_b1 , \3342_b1 , w_7918 );
xor ( \3343_b0 , \3342_b0 , w_7920 );
not ( w_7920 , w_7921 );
and ( w_7921 , w_7918 , w_7919 );
buf ( w_7918 , \303_b1 );
not ( w_7918 , w_7922 );
not ( w_7919 , w_7923 );
and ( w_7922 , w_7923 , \303_b0 );
or ( \3344_b1 , \2541_b1 , \313_b1 );
not ( \313_b1 , w_7924 );
and ( \3344_b0 , \2541_b0 , w_7925 );
and ( w_7924 , w_7925 , \313_b0 );
or ( \3345_b1 , \2532_b1 , \311_b1 );
not ( \311_b1 , w_7926 );
and ( \3345_b0 , \2532_b0 , w_7927 );
and ( w_7926 , w_7927 , \311_b0 );
or ( \3346_b1 , \3344_b1 , w_7929 );
not ( w_7929 , w_7930 );
and ( \3346_b0 , \3344_b0 , w_7931 );
and ( w_7930 ,  , w_7931 );
buf ( w_7929 , \3345_b1 );
not ( w_7929 , w_7932 );
not (  , w_7933 );
and ( w_7932 , w_7933 , \3345_b0 );
or ( \3347_b1 , \3346_b1 , w_7934 );
xor ( \3347_b0 , \3346_b0 , w_7936 );
not ( w_7936 , w_7937 );
and ( w_7937 , w_7934 , w_7935 );
buf ( w_7934 , \320_b1 );
not ( w_7934 , w_7938 );
not ( w_7935 , w_7939 );
and ( w_7938 , w_7939 , \320_b0 );
or ( \3348_b1 , \3343_b1 , \3347_b1 );
not ( \3347_b1 , w_7940 );
and ( \3348_b0 , \3343_b0 , w_7941 );
and ( w_7940 , w_7941 , \3347_b0 );
or ( \3349_b1 , \2850_b1 , \331_b1 );
not ( \331_b1 , w_7942 );
and ( \3349_b0 , \2850_b0 , w_7943 );
and ( w_7942 , w_7943 , \331_b0 );
or ( \3350_b1 , \2763_b1 , \329_b1 );
not ( \329_b1 , w_7944 );
and ( \3350_b0 , \2763_b0 , w_7945 );
and ( w_7944 , w_7945 , \329_b0 );
or ( \3351_b1 , \3349_b1 , w_7947 );
not ( w_7947 , w_7948 );
and ( \3351_b0 , \3349_b0 , w_7949 );
and ( w_7948 ,  , w_7949 );
buf ( w_7947 , \3350_b1 );
not ( w_7947 , w_7950 );
not (  , w_7951 );
and ( w_7950 , w_7951 , \3350_b0 );
or ( \3352_b1 , \3351_b1 , w_7952 );
xor ( \3352_b0 , \3351_b0 , w_7954 );
not ( w_7954 , w_7955 );
and ( w_7955 , w_7952 , w_7953 );
buf ( w_7952 , \338_b1 );
not ( w_7952 , w_7956 );
not ( w_7953 , w_7957 );
and ( w_7956 , w_7957 , \338_b0 );
or ( \3353_b1 , \3347_b1 , \3352_b1 );
not ( \3352_b1 , w_7958 );
and ( \3353_b0 , \3347_b0 , w_7959 );
and ( w_7958 , w_7959 , \3352_b0 );
or ( \3354_b1 , \3343_b1 , \3352_b1 );
not ( \3352_b1 , w_7960 );
and ( \3354_b0 , \3343_b0 , w_7961 );
and ( w_7960 , w_7961 , \3352_b0 );
or ( \3356_b1 , \1537_b1 , \740_b1 );
not ( \740_b1 , w_7962 );
and ( \3356_b0 , \1537_b0 , w_7963 );
and ( w_7962 , w_7963 , \740_b0 );
or ( \3357_b1 , \1422_b1 , \738_b1 );
not ( \738_b1 , w_7964 );
and ( \3357_b0 , \1422_b0 , w_7965 );
and ( w_7964 , w_7965 , \738_b0 );
or ( \3358_b1 , \3356_b1 , w_7967 );
not ( w_7967 , w_7968 );
and ( \3358_b0 , \3356_b0 , w_7969 );
and ( w_7968 ,  , w_7969 );
buf ( w_7967 , \3357_b1 );
not ( w_7967 , w_7970 );
not (  , w_7971 );
and ( w_7970 , w_7971 , \3357_b0 );
or ( \3359_b1 , \3358_b1 , w_7972 );
xor ( \3359_b0 , \3358_b0 , w_7974 );
not ( w_7974 , w_7975 );
and ( w_7975 , w_7972 , w_7973 );
buf ( w_7972 , \668_b1 );
not ( w_7972 , w_7976 );
not ( w_7973 , w_7977 );
and ( w_7976 , w_7977 , \668_b0 );
or ( \3360_b1 , \1778_b1 , \604_b1 );
not ( \604_b1 , w_7978 );
and ( \3360_b0 , \1778_b0 , w_7979 );
and ( w_7978 , w_7979 , \604_b0 );
or ( \3361_b1 , \1770_b1 , \602_b1 );
not ( \602_b1 , w_7980 );
and ( \3361_b0 , \1770_b0 , w_7981 );
and ( w_7980 , w_7981 , \602_b0 );
or ( \3362_b1 , \3360_b1 , w_7983 );
not ( w_7983 , w_7984 );
and ( \3362_b0 , \3360_b0 , w_7985 );
and ( w_7984 ,  , w_7985 );
buf ( w_7983 , \3361_b1 );
not ( w_7983 , w_7986 );
not (  , w_7987 );
and ( w_7986 , w_7987 , \3361_b0 );
or ( \3363_b1 , \3362_b1 , w_7988 );
xor ( \3363_b0 , \3362_b0 , w_7990 );
not ( w_7990 , w_7991 );
and ( w_7991 , w_7988 , w_7989 );
buf ( w_7988 , \561_b1 );
not ( w_7988 , w_7992 );
not ( w_7989 , w_7993 );
and ( w_7992 , w_7993 , \561_b0 );
or ( \3364_b1 , \3359_b1 , \3363_b1 );
not ( \3363_b1 , w_7994 );
and ( \3364_b0 , \3359_b0 , w_7995 );
and ( w_7994 , w_7995 , \3363_b0 );
or ( \3365_b1 , \2028_b1 , \503_b1 );
not ( \503_b1 , w_7996 );
and ( \3365_b0 , \2028_b0 , w_7997 );
and ( w_7996 , w_7997 , \503_b0 );
or ( \3366_b1 , \2023_b1 , \501_b1 );
not ( \501_b1 , w_7998 );
and ( \3366_b0 , \2023_b0 , w_7999 );
and ( w_7998 , w_7999 , \501_b0 );
or ( \3367_b1 , \3365_b1 , w_8001 );
not ( w_8001 , w_8002 );
and ( \3367_b0 , \3365_b0 , w_8003 );
and ( w_8002 ,  , w_8003 );
buf ( w_8001 , \3366_b1 );
not ( w_8001 , w_8004 );
not (  , w_8005 );
and ( w_8004 , w_8005 , \3366_b0 );
or ( \3368_b1 , \3367_b1 , w_8006 );
xor ( \3368_b0 , \3367_b0 , w_8008 );
not ( w_8008 , w_8009 );
and ( w_8009 , w_8006 , w_8007 );
buf ( w_8006 , \455_b1 );
not ( w_8006 , w_8010 );
not ( w_8007 , w_8011 );
and ( w_8010 , w_8011 , \455_b0 );
or ( \3369_b1 , \3363_b1 , \3368_b1 );
not ( \3368_b1 , w_8012 );
and ( \3369_b0 , \3363_b0 , w_8013 );
and ( w_8012 , w_8013 , \3368_b0 );
or ( \3370_b1 , \3359_b1 , \3368_b1 );
not ( \3368_b1 , w_8014 );
and ( \3370_b0 , \3359_b0 , w_8015 );
and ( w_8014 , w_8015 , \3368_b0 );
or ( \3372_b1 , \3355_b1 , \3371_b1 );
not ( \3371_b1 , w_8016 );
and ( \3372_b0 , \3355_b0 , w_8017 );
and ( w_8016 , w_8017 , \3371_b0 );
or ( \3373_b1 , \2763_b1 , \331_b1 );
not ( \331_b1 , w_8018 );
and ( \3373_b0 , \2763_b0 , w_8019 );
and ( w_8018 , w_8019 , \331_b0 );
or ( \3374_b1 , \2541_b1 , \329_b1 );
not ( \329_b1 , w_8020 );
and ( \3374_b0 , \2541_b0 , w_8021 );
and ( w_8020 , w_8021 , \329_b0 );
or ( \3375_b1 , \3373_b1 , w_8023 );
not ( w_8023 , w_8024 );
and ( \3375_b0 , \3373_b0 , w_8025 );
and ( w_8024 ,  , w_8025 );
buf ( w_8023 , \3374_b1 );
not ( w_8023 , w_8026 );
not (  , w_8027 );
and ( w_8026 , w_8027 , \3374_b0 );
or ( \3376_b1 , \3375_b1 , w_8028 );
xor ( \3376_b0 , \3375_b0 , w_8030 );
not ( w_8030 , w_8031 );
and ( w_8031 , w_8028 , w_8029 );
buf ( w_8028 , \338_b1 );
not ( w_8028 , w_8032 );
not ( w_8029 , w_8033 );
and ( w_8032 , w_8033 , \338_b0 );
or ( \3377_b1 , \3371_b1 , \3376_b1 );
not ( \3376_b1 , w_8034 );
and ( \3377_b0 , \3371_b0 , w_8035 );
and ( w_8034 , w_8035 , \3376_b0 );
or ( \3378_b1 , \3355_b1 , \3376_b1 );
not ( \3376_b1 , w_8036 );
and ( \3378_b0 , \3355_b0 , w_8037 );
and ( w_8036 , w_8037 , \3376_b0 );
or ( \3380_b1 , \3339_b1 , \3379_b1 );
not ( \3379_b1 , w_8038 );
and ( \3380_b0 , \3339_b0 , w_8039 );
and ( w_8038 , w_8039 , \3379_b0 );
or ( \3381_b1 , \2850_b1 , w_8041 );
not ( w_8041 , w_8042 );
and ( \3381_b0 , \2850_b0 , w_8043 );
and ( w_8042 ,  , w_8043 );
buf ( w_8041 , \349_b1 );
not ( w_8041 , w_8044 );
not (  , w_8045 );
and ( w_8044 , w_8045 , \349_b0 );
or ( \3382_b1 , \3381_b1 , w_8046 );
xor ( \3382_b0 , \3381_b0 , w_8048 );
not ( w_8048 , w_8049 );
and ( w_8049 , w_8046 , w_8047 );
buf ( w_8046 , \358_b1 );
not ( w_8046 , w_8050 );
not ( w_8047 , w_8051 );
and ( w_8050 , w_8051 , \358_b0 );
or ( \3383_b1 , \3191_b1 , \3195_b1 );
xor ( \3383_b0 , \3191_b0 , w_8052 );
not ( w_8052 , w_8053 );
and ( w_8053 , \3195_b1 , \3195_b0 );
or ( \3384_b1 , \3383_b1 , \3200_b1 );
xor ( \3384_b0 , \3383_b0 , w_8054 );
not ( w_8054 , w_8055 );
and ( w_8055 , \3200_b1 , \3200_b0 );
or ( \3385_b1 , \3382_b1 , \3384_b1 );
not ( \3384_b1 , w_8056 );
and ( \3385_b0 , \3382_b0 , w_8057 );
and ( w_8056 , w_8057 , \3384_b0 );
or ( \3386_b1 , \3207_b1 , \3211_b1 );
xor ( \3386_b0 , \3207_b0 , w_8058 );
not ( w_8058 , w_8059 );
and ( w_8059 , \3211_b1 , \3211_b0 );
or ( \3387_b1 , \3386_b1 , \3216_b1 );
xor ( \3387_b0 , \3386_b0 , w_8060 );
not ( w_8060 , w_8061 );
and ( w_8061 , \3216_b1 , \3216_b0 );
or ( \3388_b1 , \3384_b1 , \3387_b1 );
not ( \3387_b1 , w_8062 );
and ( \3388_b0 , \3384_b0 , w_8063 );
and ( w_8062 , w_8063 , \3387_b0 );
or ( \3389_b1 , \3382_b1 , \3387_b1 );
not ( \3387_b1 , w_8064 );
and ( \3389_b0 , \3382_b0 , w_8065 );
and ( w_8064 , w_8065 , \3387_b0 );
or ( \3391_b1 , \3379_b1 , \3390_b1 );
not ( \3390_b1 , w_8066 );
and ( \3391_b0 , \3379_b0 , w_8067 );
and ( w_8066 , w_8067 , \3390_b0 );
or ( \3392_b1 , \3339_b1 , \3390_b1 );
not ( \3390_b1 , w_8068 );
and ( \3392_b0 , \3339_b0 , w_8069 );
and ( w_8068 , w_8069 , \3390_b0 );
or ( \3394_b1 , \3143_b1 , \3147_b1 );
xor ( \3394_b0 , \3143_b0 , w_8070 );
not ( w_8070 , w_8071 );
and ( w_8071 , \3147_b1 , \3147_b0 );
or ( \3395_b1 , \3394_b1 , \3152_b1 );
xor ( \3395_b0 , \3394_b0 , w_8072 );
not ( w_8072 , w_8073 );
and ( w_8073 , \3152_b1 , \3152_b0 );
or ( \3396_b1 , \3159_b1 , \3163_b1 );
xor ( \3396_b0 , \3159_b0 , w_8074 );
not ( w_8074 , w_8075 );
and ( w_8075 , \3163_b1 , \3163_b0 );
or ( \3397_b1 , \3396_b1 , \3168_b1 );
xor ( \3397_b0 , \3396_b0 , w_8076 );
not ( w_8076 , w_8077 );
and ( w_8077 , \3168_b1 , \3168_b0 );
or ( \3398_b1 , \3395_b1 , \3397_b1 );
not ( \3397_b1 , w_8078 );
and ( \3398_b0 , \3395_b0 , w_8079 );
and ( w_8078 , w_8079 , \3397_b0 );
or ( \3399_b1 , \3176_b1 , \3180_b1 );
xor ( \3399_b0 , \3176_b0 , w_8080 );
not ( w_8080 , w_8081 );
and ( w_8081 , \3180_b1 , \3180_b0 );
or ( \3400_b1 , \3399_b1 , \358_b1 );
xor ( \3400_b0 , \3399_b0 , w_8082 );
not ( w_8082 , w_8083 );
and ( w_8083 , \358_b1 , \358_b0 );
or ( \3401_b1 , \3397_b1 , \3400_b1 );
not ( \3400_b1 , w_8084 );
and ( \3401_b0 , \3397_b0 , w_8085 );
and ( w_8084 , w_8085 , \3400_b0 );
or ( \3402_b1 , \3395_b1 , \3400_b1 );
not ( \3400_b1 , w_8086 );
and ( \3402_b0 , \3395_b0 , w_8087 );
and ( w_8086 , w_8087 , \3400_b0 );
or ( \3404_b1 , \2996_b1 , \3000_b1 );
xor ( \3404_b0 , \2996_b0 , w_8088 );
not ( w_8088 , w_8089 );
and ( w_8089 , \3000_b1 , \3000_b0 );
or ( \3405_b1 , \3404_b1 , \3005_b1 );
xor ( \3405_b0 , \3404_b0 , w_8090 );
not ( w_8090 , w_8091 );
and ( w_8091 , \3005_b1 , \3005_b0 );
or ( \3406_b1 , \3403_b1 , \3405_b1 );
not ( \3405_b1 , w_8092 );
and ( \3406_b0 , \3403_b0 , w_8093 );
and ( w_8092 , w_8093 , \3405_b0 );
or ( \3407_b1 , \3012_b1 , \3016_b1 );
xor ( \3407_b0 , \3012_b0 , w_8094 );
not ( w_8094 , w_8095 );
and ( w_8095 , \3016_b1 , \3016_b0 );
or ( \3408_b1 , \3407_b1 , \3021_b1 );
xor ( \3408_b0 , \3407_b0 , w_8096 );
not ( w_8096 , w_8097 );
and ( w_8097 , \3021_b1 , \3021_b0 );
or ( \3409_b1 , \3405_b1 , \3408_b1 );
not ( \3408_b1 , w_8098 );
and ( \3409_b0 , \3405_b0 , w_8099 );
and ( w_8098 , w_8099 , \3408_b0 );
or ( \3410_b1 , \3403_b1 , \3408_b1 );
not ( \3408_b1 , w_8100 );
and ( \3410_b0 , \3403_b0 , w_8101 );
and ( w_8100 , w_8101 , \3408_b0 );
or ( \3412_b1 , \3393_b1 , \3411_b1 );
not ( \3411_b1 , w_8102 );
and ( \3412_b0 , \3393_b0 , w_8103 );
and ( w_8102 , w_8103 , \3411_b0 );
or ( \3413_b1 , \3155_b1 , \3171_b1 );
xor ( \3413_b0 , \3155_b0 , w_8104 );
not ( w_8104 , w_8105 );
and ( w_8105 , \3171_b1 , \3171_b0 );
or ( \3414_b1 , \3413_b1 , \3184_b1 );
xor ( \3414_b0 , \3413_b0 , w_8106 );
not ( w_8106 , w_8107 );
and ( w_8107 , \3184_b1 , \3184_b0 );
or ( \3415_b1 , \3203_b1 , \3219_b1 );
xor ( \3415_b0 , \3203_b0 , w_8108 );
not ( w_8108 , w_8109 );
and ( w_8109 , \3219_b1 , \3219_b0 );
or ( \3416_b1 , \3415_b1 , \3224_b1 );
xor ( \3416_b0 , \3415_b0 , w_8110 );
not ( w_8110 , w_8111 );
and ( w_8111 , \3224_b1 , \3224_b0 );
or ( \3417_b1 , \3414_b1 , \3416_b1 );
not ( \3416_b1 , w_8112 );
and ( \3417_b0 , \3414_b0 , w_8113 );
and ( w_8112 , w_8113 , \3416_b0 );
or ( \3418_b1 , \3230_b1 , \3232_b1 );
xor ( \3418_b0 , \3230_b0 , w_8114 );
not ( w_8114 , w_8115 );
and ( w_8115 , \3232_b1 , \3232_b0 );
or ( \3419_b1 , \3418_b1 , \3235_b1 );
xor ( \3419_b0 , \3418_b0 , w_8116 );
not ( w_8116 , w_8117 );
and ( w_8117 , \3235_b1 , \3235_b0 );
or ( \3420_b1 , \3416_b1 , \3419_b1 );
not ( \3419_b1 , w_8118 );
and ( \3420_b0 , \3416_b0 , w_8119 );
and ( w_8118 , w_8119 , \3419_b0 );
or ( \3421_b1 , \3414_b1 , \3419_b1 );
not ( \3419_b1 , w_8120 );
and ( \3421_b0 , \3414_b0 , w_8121 );
and ( w_8120 , w_8121 , \3419_b0 );
or ( \3423_b1 , \3411_b1 , \3422_b1 );
not ( \3422_b1 , w_8122 );
and ( \3423_b0 , \3411_b0 , w_8123 );
and ( w_8122 , w_8123 , \3422_b0 );
or ( \3424_b1 , \3393_b1 , \3422_b1 );
not ( \3422_b1 , w_8124 );
and ( \3424_b0 , \3393_b0 , w_8125 );
and ( w_8124 , w_8125 , \3422_b0 );
or ( \3426_b1 , \3187_b1 , \3227_b1 );
xor ( \3426_b0 , \3187_b0 , w_8126 );
not ( w_8126 , w_8127 );
and ( w_8127 , \3227_b1 , \3227_b0 );
or ( \3427_b1 , \3426_b1 , \3238_b1 );
xor ( \3427_b0 , \3426_b0 , w_8128 );
not ( w_8128 , w_8129 );
and ( w_8129 , \3238_b1 , \3238_b0 );
or ( \3428_b1 , \3243_b1 , \3245_b1 );
xor ( \3428_b0 , \3243_b0 , w_8130 );
not ( w_8130 , w_8131 );
and ( w_8131 , \3245_b1 , \3245_b0 );
or ( \3429_b1 , \3428_b1 , \3247_b1 );
xor ( \3429_b0 , \3428_b0 , w_8132 );
not ( w_8132 , w_8133 );
and ( w_8133 , \3247_b1 , \3247_b0 );
or ( \3430_b1 , \3427_b1 , \3429_b1 );
not ( \3429_b1 , w_8134 );
and ( \3430_b0 , \3427_b0 , w_8135 );
and ( w_8134 , w_8135 , \3429_b0 );
or ( \3431_b1 , \3253_b1 , \3255_b1 );
xor ( \3431_b0 , \3253_b0 , w_8136 );
not ( w_8136 , w_8137 );
and ( w_8137 , \3255_b1 , \3255_b0 );
or ( \3432_b1 , \3429_b1 , \3431_b1 );
not ( \3431_b1 , w_8138 );
and ( \3432_b0 , \3429_b0 , w_8139 );
and ( w_8138 , w_8139 , \3431_b0 );
or ( \3433_b1 , \3427_b1 , \3431_b1 );
not ( \3431_b1 , w_8140 );
and ( \3433_b0 , \3427_b0 , w_8141 );
and ( w_8140 , w_8141 , \3431_b0 );
or ( \3435_b1 , \3425_b1 , \3434_b1 );
not ( \3434_b1 , w_8142 );
and ( \3435_b0 , \3425_b0 , w_8143 );
and ( w_8142 , w_8143 , \3434_b0 );
or ( \3436_b1 , \3261_b1 , \3263_b1 );
xor ( \3436_b0 , \3261_b0 , w_8144 );
not ( w_8144 , w_8145 );
and ( w_8145 , \3263_b1 , \3263_b0 );
or ( \3437_b1 , \3436_b1 , \3266_b1 );
xor ( \3437_b0 , \3436_b0 , w_8146 );
not ( w_8146 , w_8147 );
and ( w_8147 , \3266_b1 , \3266_b0 );
or ( \3438_b1 , \3434_b1 , \3437_b1 );
not ( \3437_b1 , w_8148 );
and ( \3438_b0 , \3434_b0 , w_8149 );
and ( w_8148 , w_8149 , \3437_b0 );
or ( \3439_b1 , \3425_b1 , \3437_b1 );
not ( \3437_b1 , w_8150 );
and ( \3439_b0 , \3425_b0 , w_8151 );
and ( w_8150 , w_8151 , \3437_b0 );
or ( \3441_b1 , \3096_b1 , \3106_b1 );
xor ( \3441_b0 , \3096_b0 , w_8152 );
not ( w_8152 , w_8153 );
and ( w_8153 , \3106_b1 , \3106_b0 );
or ( \3442_b1 , \3441_b1 , \3109_b1 );
xor ( \3442_b0 , \3441_b0 , w_8154 );
not ( w_8154 , w_8155 );
and ( w_8155 , \3109_b1 , \3109_b0 );
or ( \3443_b1 , \3440_b1 , \3442_b1 );
not ( \3442_b1 , w_8156 );
and ( \3443_b0 , \3440_b0 , w_8157 );
and ( w_8156 , w_8157 , \3442_b0 );
or ( \3444_b1 , \3259_b1 , \3269_b1 );
xor ( \3444_b0 , \3259_b0 , w_8158 );
not ( w_8158 , w_8159 );
and ( w_8159 , \3269_b1 , \3269_b0 );
or ( \3445_b1 , \3444_b1 , \3272_b1 );
xor ( \3445_b0 , \3444_b0 , w_8160 );
not ( w_8160 , w_8161 );
and ( w_8161 , \3272_b1 , \3272_b0 );
or ( \3446_b1 , \3442_b1 , \3445_b1 );
not ( \3445_b1 , w_8162 );
and ( \3446_b0 , \3442_b0 , w_8163 );
and ( w_8162 , w_8163 , \3445_b0 );
or ( \3447_b1 , \3440_b1 , \3445_b1 );
not ( \3445_b1 , w_8164 );
and ( \3447_b0 , \3440_b0 , w_8165 );
and ( w_8164 , w_8165 , \3445_b0 );
or ( \3449_b1 , \3287_b1 , \3448_b1 );
not ( \3448_b1 , w_8166 );
and ( \3449_b0 , \3287_b0 , w_8167 );
and ( w_8166 , w_8167 , \3448_b0 );
or ( \3450_b1 , \3287_b1 , \3448_b1 );
xor ( \3450_b0 , \3287_b0 , w_8168 );
not ( w_8168 , w_8169 );
and ( w_8169 , \3448_b1 , \3448_b0 );
or ( \3451_b1 , \3440_b1 , \3442_b1 );
xor ( \3451_b0 , \3440_b0 , w_8170 );
not ( w_8170 , w_8171 );
and ( w_8171 , \3442_b1 , \3442_b0 );
or ( \3452_b1 , \3451_b1 , \3445_b1 );
xor ( \3452_b0 , \3451_b0 , w_8172 );
not ( w_8172 , w_8173 );
and ( w_8173 , \3445_b1 , \3445_b0 );
or ( \3453_b1 , \841_b1 , \1476_b1 );
not ( \1476_b1 , w_8174 );
and ( \3453_b0 , \841_b0 , w_8175 );
and ( w_8174 , w_8175 , \1476_b0 );
or ( \3454_b1 , \777_b1 , \1474_b1 );
not ( \1474_b1 , w_8176 );
and ( \3454_b0 , \777_b0 , w_8177 );
and ( w_8176 , w_8177 , \1474_b0 );
or ( \3455_b1 , \3453_b1 , w_8179 );
not ( w_8179 , w_8180 );
and ( \3455_b0 , \3453_b0 , w_8181 );
and ( w_8180 ,  , w_8181 );
buf ( w_8179 , \3454_b1 );
not ( w_8179 , w_8182 );
not (  , w_8183 );
and ( w_8182 , w_8183 , \3454_b0 );
or ( \3456_b1 , \3455_b1 , w_8184 );
xor ( \3456_b0 , \3455_b0 , w_8186 );
not ( w_8186 , w_8187 );
and ( w_8187 , w_8184 , w_8185 );
buf ( w_8184 , \1363_b1 );
not ( w_8184 , w_8188 );
not ( w_8185 , w_8189 );
and ( w_8188 , w_8189 , \1363_b0 );
or ( \3457_b1 , \1104_b1 , \1280_b1 );
not ( \1280_b1 , w_8190 );
and ( \3457_b0 , \1104_b0 , w_8191 );
and ( w_8190 , w_8191 , \1280_b0 );
or ( \3458_b1 , \904_b1 , \1278_b1 );
not ( \1278_b1 , w_8192 );
and ( \3458_b0 , \904_b0 , w_8193 );
and ( w_8192 , w_8193 , \1278_b0 );
or ( \3459_b1 , \3457_b1 , w_8195 );
not ( w_8195 , w_8196 );
and ( \3459_b0 , \3457_b0 , w_8197 );
and ( w_8196 ,  , w_8197 );
buf ( w_8195 , \3458_b1 );
not ( w_8195 , w_8198 );
not (  , w_8199 );
and ( w_8198 , w_8199 , \3458_b0 );
or ( \3460_b1 , \3459_b1 , w_8200 );
xor ( \3460_b0 , \3459_b0 , w_8202 );
not ( w_8202 , w_8203 );
and ( w_8203 , w_8200 , w_8201 );
buf ( w_8200 , \1177_b1 );
not ( w_8200 , w_8204 );
not ( w_8201 , w_8205 );
and ( w_8204 , w_8205 , \1177_b0 );
or ( \3461_b1 , \3456_b1 , \3460_b1 );
not ( \3460_b1 , w_8206 );
and ( \3461_b0 , \3456_b0 , w_8207 );
and ( w_8206 , w_8207 , \3460_b0 );
or ( \3462_b1 , \1299_b1 , \1062_b1 );
not ( \1062_b1 , w_8208 );
and ( \3462_b0 , \1299_b0 , w_8209 );
and ( w_8208 , w_8209 , \1062_b0 );
or ( \3463_b1 , \1194_b1 , \1060_b1 );
not ( \1060_b1 , w_8210 );
and ( \3463_b0 , \1194_b0 , w_8211 );
and ( w_8210 , w_8211 , \1060_b0 );
or ( \3464_b1 , \3462_b1 , w_8213 );
not ( w_8213 , w_8214 );
and ( \3464_b0 , \3462_b0 , w_8215 );
and ( w_8214 ,  , w_8215 );
buf ( w_8213 , \3463_b1 );
not ( w_8213 , w_8216 );
not (  , w_8217 );
and ( w_8216 , w_8217 , \3463_b0 );
or ( \3465_b1 , \3464_b1 , w_8218 );
xor ( \3465_b0 , \3464_b0 , w_8220 );
not ( w_8220 , w_8221 );
and ( w_8221 , w_8218 , w_8219 );
buf ( w_8218 , \984_b1 );
not ( w_8218 , w_8222 );
not ( w_8219 , w_8223 );
and ( w_8222 , w_8223 , \984_b0 );
or ( \3466_b1 , \3460_b1 , \3465_b1 );
not ( \3465_b1 , w_8224 );
and ( \3466_b0 , \3460_b0 , w_8225 );
and ( w_8224 , w_8225 , \3465_b0 );
or ( \3467_b1 , \3456_b1 , \3465_b1 );
not ( \3465_b1 , w_8226 );
and ( \3467_b0 , \3456_b0 , w_8227 );
and ( w_8226 , w_8227 , \3465_b0 );
or ( \3469_b1 , \444_b1 , \2261_b1 );
not ( \2261_b1 , w_8228 );
and ( \3469_b0 , \444_b0 , w_8229 );
and ( w_8228 , w_8229 , \2261_b0 );
or ( \3470_b1 , \360_b1 , \2259_b1 );
not ( \2259_b1 , w_8230 );
and ( \3470_b0 , \360_b0 , w_8231 );
and ( w_8230 , w_8231 , \2259_b0 );
or ( \3471_b1 , \3469_b1 , w_8233 );
not ( w_8233 , w_8234 );
and ( \3471_b0 , \3469_b0 , w_8235 );
and ( w_8234 ,  , w_8235 );
buf ( w_8233 , \3470_b1 );
not ( w_8233 , w_8236 );
not (  , w_8237 );
and ( w_8236 , w_8237 , \3470_b0 );
or ( \3472_b1 , \3471_b1 , w_8238 );
xor ( \3472_b0 , \3471_b0 , w_8240 );
not ( w_8240 , w_8241 );
and ( w_8241 , w_8238 , w_8239 );
buf ( w_8238 , \2124_b1 );
not ( w_8238 , w_8242 );
not ( w_8239 , w_8243 );
and ( w_8242 , w_8243 , \2124_b0 );
or ( \3473_b1 , \593_b1 , \1955_b1 );
not ( \1955_b1 , w_8244 );
and ( \3473_b0 , \593_b0 , w_8245 );
and ( w_8244 , w_8245 , \1955_b0 );
or ( \3474_b1 , \495_b1 , \1953_b1 );
not ( \1953_b1 , w_8246 );
and ( \3474_b0 , \495_b0 , w_8247 );
and ( w_8246 , w_8247 , \1953_b0 );
or ( \3475_b1 , \3473_b1 , w_8249 );
not ( w_8249 , w_8250 );
and ( \3475_b0 , \3473_b0 , w_8251 );
and ( w_8250 ,  , w_8251 );
buf ( w_8249 , \3474_b1 );
not ( w_8249 , w_8252 );
not (  , w_8253 );
and ( w_8252 , w_8253 , \3474_b0 );
or ( \3476_b1 , \3475_b1 , w_8254 );
xor ( \3476_b0 , \3475_b0 , w_8256 );
not ( w_8256 , w_8257 );
and ( w_8257 , w_8254 , w_8255 );
buf ( w_8254 , \1835_b1 );
not ( w_8254 , w_8258 );
not ( w_8255 , w_8259 );
and ( w_8258 , w_8259 , \1835_b0 );
or ( \3477_b1 , \3472_b1 , \3476_b1 );
not ( \3476_b1 , w_8260 );
and ( \3477_b0 , \3472_b0 , w_8261 );
and ( w_8260 , w_8261 , \3476_b0 );
or ( \3478_b1 , \703_b1 , \1742_b1 );
not ( \1742_b1 , w_8262 );
and ( \3478_b0 , \703_b0 , w_8263 );
and ( w_8262 , w_8263 , \1742_b0 );
or ( \3479_b1 , \621_b1 , \1740_b1 );
not ( \1740_b1 , w_8264 );
and ( \3479_b0 , \621_b0 , w_8265 );
and ( w_8264 , w_8265 , \1740_b0 );
or ( \3480_b1 , \3478_b1 , w_8267 );
not ( w_8267 , w_8268 );
and ( \3480_b0 , \3478_b0 , w_8269 );
and ( w_8268 ,  , w_8269 );
buf ( w_8267 , \3479_b1 );
not ( w_8267 , w_8270 );
not (  , w_8271 );
and ( w_8270 , w_8271 , \3479_b0 );
or ( \3481_b1 , \3480_b1 , w_8272 );
xor ( \3481_b0 , \3480_b0 , w_8274 );
not ( w_8274 , w_8275 );
and ( w_8275 , w_8272 , w_8273 );
buf ( w_8272 , \1610_b1 );
not ( w_8272 , w_8276 );
not ( w_8273 , w_8277 );
and ( w_8276 , w_8277 , \1610_b0 );
or ( \3482_b1 , \3476_b1 , \3481_b1 );
not ( \3481_b1 , w_8278 );
and ( \3482_b0 , \3476_b0 , w_8279 );
and ( w_8278 , w_8279 , \3481_b0 );
or ( \3483_b1 , \3472_b1 , \3481_b1 );
not ( \3481_b1 , w_8280 );
and ( \3483_b0 , \3472_b0 , w_8281 );
and ( w_8280 , w_8281 , \3481_b0 );
or ( \3485_b1 , \3468_b1 , \3484_b1 );
not ( \3484_b1 , w_8282 );
and ( \3485_b0 , \3468_b0 , w_8283 );
and ( w_8282 , w_8283 , \3484_b0 );
or ( \3486_b1 , \323_b1 , \2913_b1 );
not ( \2913_b1 , w_8284 );
and ( \3486_b0 , \323_b0 , w_8285 );
and ( w_8284 , w_8285 , \2913_b0 );
or ( \3487_b1 , \333_b1 , \2910_b1 );
not ( \2910_b1 , w_8286 );
and ( \3487_b0 , \333_b0 , w_8287 );
and ( w_8286 , w_8287 , \2910_b0 );
or ( \3488_b1 , \3486_b1 , w_8289 );
not ( w_8289 , w_8290 );
and ( \3488_b0 , \3486_b0 , w_8291 );
and ( w_8290 ,  , w_8291 );
buf ( w_8289 , \3487_b1 );
not ( w_8289 , w_8292 );
not (  , w_8293 );
and ( w_8292 , w_8293 , \3487_b0 );
or ( \3489_b1 , \3488_b1 , w_8294 );
xor ( \3489_b0 , \3488_b0 , w_8296 );
not ( w_8296 , w_8297 );
and ( w_8297 , w_8294 , w_8295 );
buf ( w_8294 , \2371_b1 );
not ( w_8294 , w_8298 );
not ( w_8295 , w_8299 );
and ( w_8298 , w_8299 , \2371_b0 );
or ( \3490_b1 , \343_b1 , \2550_b1 );
not ( \2550_b1 , w_8300 );
and ( \3490_b0 , \343_b0 , w_8301 );
and ( w_8300 , w_8301 , \2550_b0 );
or ( \3491_b1 , \353_b1 , \2548_b1 );
not ( \2548_b1 , w_8302 );
and ( \3491_b0 , \353_b0 , w_8303 );
and ( w_8302 , w_8303 , \2548_b0 );
or ( \3492_b1 , \3490_b1 , w_8305 );
not ( w_8305 , w_8306 );
and ( \3492_b0 , \3490_b0 , w_8307 );
and ( w_8306 ,  , w_8307 );
buf ( w_8305 , \3491_b1 );
not ( w_8305 , w_8308 );
not (  , w_8309 );
and ( w_8308 , w_8309 , \3491_b0 );
or ( \3493_b1 , \3492_b1 , w_8310 );
xor ( \3493_b0 , \3492_b0 , w_8312 );
not ( w_8312 , w_8313 );
and ( w_8313 , w_8310 , w_8311 );
buf ( w_8310 , \2374_b1 );
not ( w_8310 , w_8314 );
not ( w_8311 , w_8315 );
and ( w_8314 , w_8315 , \2374_b0 );
or ( \3494_b1 , \3489_b1 , \3493_b1 );
not ( \3493_b1 , w_8316 );
and ( \3494_b0 , \3489_b0 , w_8317 );
and ( w_8316 , w_8317 , \3493_b0 );
or ( \3495_b1 , \3493_b1 , \338_b1 );
not ( \338_b1 , w_8318 );
and ( \3495_b0 , \3493_b0 , w_8319 );
and ( w_8318 , w_8319 , \338_b0 );
or ( \3496_b1 , \3489_b1 , \338_b1 );
not ( \338_b1 , w_8320 );
and ( \3496_b0 , \3489_b0 , w_8321 );
and ( w_8320 , w_8321 , \338_b0 );
or ( \3498_b1 , \3484_b1 , \3497_b1 );
not ( \3497_b1 , w_8322 );
and ( \3498_b0 , \3484_b0 , w_8323 );
and ( w_8322 , w_8323 , \3497_b0 );
or ( \3499_b1 , \3468_b1 , \3497_b1 );
not ( \3497_b1 , w_8324 );
and ( \3499_b0 , \3468_b0 , w_8325 );
and ( w_8324 , w_8325 , \3497_b0 );
or ( \3501_b1 , \1422_b1 , \912_b1 );
not ( \912_b1 , w_8326 );
and ( \3501_b0 , \1422_b0 , w_8327 );
and ( w_8326 , w_8327 , \912_b0 );
or ( \3502_b1 , \1304_b1 , \910_b1 );
not ( \910_b1 , w_8328 );
and ( \3502_b0 , \1304_b0 , w_8329 );
and ( w_8328 , w_8329 , \910_b0 );
or ( \3503_b1 , \3501_b1 , w_8331 );
not ( w_8331 , w_8332 );
and ( \3503_b0 , \3501_b0 , w_8333 );
and ( w_8332 ,  , w_8333 );
buf ( w_8331 , \3502_b1 );
not ( w_8331 , w_8334 );
not (  , w_8335 );
and ( w_8334 , w_8335 , \3502_b0 );
or ( \3504_b1 , \3503_b1 , w_8336 );
xor ( \3504_b0 , \3503_b0 , w_8338 );
not ( w_8338 , w_8339 );
and ( w_8339 , w_8336 , w_8337 );
buf ( w_8336 , \818_b1 );
not ( w_8336 , w_8340 );
not ( w_8337 , w_8341 );
and ( w_8340 , w_8341 , \818_b0 );
or ( \3505_b1 , \1770_b1 , \740_b1 );
not ( \740_b1 , w_8342 );
and ( \3505_b0 , \1770_b0 , w_8343 );
and ( w_8342 , w_8343 , \740_b0 );
or ( \3506_b1 , \1537_b1 , \738_b1 );
not ( \738_b1 , w_8344 );
and ( \3506_b0 , \1537_b0 , w_8345 );
and ( w_8344 , w_8345 , \738_b0 );
or ( \3507_b1 , \3505_b1 , w_8347 );
not ( w_8347 , w_8348 );
and ( \3507_b0 , \3505_b0 , w_8349 );
and ( w_8348 ,  , w_8349 );
buf ( w_8347 , \3506_b1 );
not ( w_8347 , w_8350 );
not (  , w_8351 );
and ( w_8350 , w_8351 , \3506_b0 );
or ( \3508_b1 , \3507_b1 , w_8352 );
xor ( \3508_b0 , \3507_b0 , w_8354 );
not ( w_8354 , w_8355 );
and ( w_8355 , w_8352 , w_8353 );
buf ( w_8352 , \668_b1 );
not ( w_8352 , w_8356 );
not ( w_8353 , w_8357 );
and ( w_8356 , w_8357 , \668_b0 );
or ( \3509_b1 , \3504_b1 , \3508_b1 );
not ( \3508_b1 , w_8358 );
and ( \3509_b0 , \3504_b0 , w_8359 );
and ( w_8358 , w_8359 , \3508_b0 );
or ( \3510_b1 , \2023_b1 , \604_b1 );
not ( \604_b1 , w_8360 );
and ( \3510_b0 , \2023_b0 , w_8361 );
and ( w_8360 , w_8361 , \604_b0 );
or ( \3511_b1 , \1778_b1 , \602_b1 );
not ( \602_b1 , w_8362 );
and ( \3511_b0 , \1778_b0 , w_8363 );
and ( w_8362 , w_8363 , \602_b0 );
or ( \3512_b1 , \3510_b1 , w_8365 );
not ( w_8365 , w_8366 );
and ( \3512_b0 , \3510_b0 , w_8367 );
and ( w_8366 ,  , w_8367 );
buf ( w_8365 , \3511_b1 );
not ( w_8365 , w_8368 );
not (  , w_8369 );
and ( w_8368 , w_8369 , \3511_b0 );
or ( \3513_b1 , \3512_b1 , w_8370 );
xor ( \3513_b0 , \3512_b0 , w_8372 );
not ( w_8372 , w_8373 );
and ( w_8373 , w_8370 , w_8371 );
buf ( w_8370 , \561_b1 );
not ( w_8370 , w_8374 );
not ( w_8371 , w_8375 );
and ( w_8374 , w_8375 , \561_b0 );
or ( \3514_b1 , \3508_b1 , \3513_b1 );
not ( \3513_b1 , w_8376 );
and ( \3514_b0 , \3508_b0 , w_8377 );
and ( w_8376 , w_8377 , \3513_b0 );
or ( \3515_b1 , \3504_b1 , \3513_b1 );
not ( \3513_b1 , w_8378 );
and ( \3515_b0 , \3504_b0 , w_8379 );
and ( w_8378 , w_8379 , \3513_b0 );
or ( \3517_b1 , \2161_b1 , \503_b1 );
not ( \503_b1 , w_8380 );
and ( \3517_b0 , \2161_b0 , w_8381 );
and ( w_8380 , w_8381 , \503_b0 );
or ( \3518_b1 , \2028_b1 , \501_b1 );
not ( \501_b1 , w_8382 );
and ( \3518_b0 , \2028_b0 , w_8383 );
and ( w_8382 , w_8383 , \501_b0 );
or ( \3519_b1 , \3517_b1 , w_8385 );
not ( w_8385 , w_8386 );
and ( \3519_b0 , \3517_b0 , w_8387 );
and ( w_8386 ,  , w_8387 );
buf ( w_8385 , \3518_b1 );
not ( w_8385 , w_8388 );
not (  , w_8389 );
and ( w_8388 , w_8389 , \3518_b0 );
or ( \3520_b1 , \3519_b1 , w_8390 );
xor ( \3520_b0 , \3519_b0 , w_8392 );
not ( w_8392 , w_8393 );
and ( w_8393 , w_8390 , w_8391 );
buf ( w_8390 , \455_b1 );
not ( w_8390 , w_8394 );
not ( w_8391 , w_8395 );
and ( w_8394 , w_8395 , \455_b0 );
or ( \3521_b1 , \2532_b1 , \298_b1 );
not ( \298_b1 , w_8396 );
and ( \3521_b0 , \2532_b0 , w_8397 );
and ( w_8396 , w_8397 , \298_b0 );
or ( \3522_b1 , \2305_b1 , \296_b1 );
not ( \296_b1 , w_8398 );
and ( \3522_b0 , \2305_b0 , w_8399 );
and ( w_8398 , w_8399 , \296_b0 );
or ( \3523_b1 , \3521_b1 , w_8401 );
not ( w_8401 , w_8402 );
and ( \3523_b0 , \3521_b0 , w_8403 );
and ( w_8402 ,  , w_8403 );
buf ( w_8401 , \3522_b1 );
not ( w_8401 , w_8404 );
not (  , w_8405 );
and ( w_8404 , w_8405 , \3522_b0 );
or ( \3524_b1 , \3523_b1 , w_8406 );
xor ( \3524_b0 , \3523_b0 , w_8408 );
not ( w_8408 , w_8409 );
and ( w_8409 , w_8406 , w_8407 );
buf ( w_8406 , \303_b1 );
not ( w_8406 , w_8410 );
not ( w_8407 , w_8411 );
and ( w_8410 , w_8411 , \303_b0 );
or ( \3525_b1 , \3520_b1 , \3524_b1 );
not ( \3524_b1 , w_8412 );
and ( \3525_b0 , \3520_b0 , w_8413 );
and ( w_8412 , w_8413 , \3524_b0 );
or ( \3526_b1 , \2763_b1 , \313_b1 );
not ( \313_b1 , w_8414 );
and ( \3526_b0 , \2763_b0 , w_8415 );
and ( w_8414 , w_8415 , \313_b0 );
or ( \3527_b1 , \2541_b1 , \311_b1 );
not ( \311_b1 , w_8416 );
and ( \3527_b0 , \2541_b0 , w_8417 );
and ( w_8416 , w_8417 , \311_b0 );
or ( \3528_b1 , \3526_b1 , w_8419 );
not ( w_8419 , w_8420 );
and ( \3528_b0 , \3526_b0 , w_8421 );
and ( w_8420 ,  , w_8421 );
buf ( w_8419 , \3527_b1 );
not ( w_8419 , w_8422 );
not (  , w_8423 );
and ( w_8422 , w_8423 , \3527_b0 );
or ( \3529_b1 , \3528_b1 , w_8424 );
xor ( \3529_b0 , \3528_b0 , w_8426 );
not ( w_8426 , w_8427 );
and ( w_8427 , w_8424 , w_8425 );
buf ( w_8424 , \320_b1 );
not ( w_8424 , w_8428 );
not ( w_8425 , w_8429 );
and ( w_8428 , w_8429 , \320_b0 );
or ( \3530_b1 , \3524_b1 , \3529_b1 );
not ( \3529_b1 , w_8430 );
and ( \3530_b0 , \3524_b0 , w_8431 );
and ( w_8430 , w_8431 , \3529_b0 );
or ( \3531_b1 , \3520_b1 , \3529_b1 );
not ( \3529_b1 , w_8432 );
and ( \3531_b0 , \3520_b0 , w_8433 );
and ( w_8432 , w_8433 , \3529_b0 );
or ( \3533_b1 , \3516_b1 , \3532_b1 );
not ( \3532_b1 , w_8434 );
and ( \3533_b0 , \3516_b0 , w_8435 );
and ( w_8434 , w_8435 , \3532_b0 );
or ( \3534_b1 , \3343_b1 , \3347_b1 );
xor ( \3534_b0 , \3343_b0 , w_8436 );
not ( w_8436 , w_8437 );
and ( w_8437 , \3347_b1 , \3347_b0 );
or ( \3535_b1 , \3534_b1 , \3352_b1 );
xor ( \3535_b0 , \3534_b0 , w_8438 );
not ( w_8438 , w_8439 );
and ( w_8439 , \3352_b1 , \3352_b0 );
or ( \3536_b1 , \3532_b1 , \3535_b1 );
not ( \3535_b1 , w_8440 );
and ( \3536_b0 , \3532_b0 , w_8441 );
and ( w_8440 , w_8441 , \3535_b0 );
or ( \3537_b1 , \3516_b1 , \3535_b1 );
not ( \3535_b1 , w_8442 );
and ( \3537_b0 , \3516_b0 , w_8443 );
and ( w_8442 , w_8443 , \3535_b0 );
or ( \3539_b1 , \3500_b1 , \3538_b1 );
not ( \3538_b1 , w_8444 );
and ( \3539_b0 , \3500_b0 , w_8445 );
and ( w_8444 , w_8445 , \3538_b0 );
or ( \3540_b1 , \3291_b1 , \3295_b1 );
xor ( \3540_b0 , \3291_b0 , w_8446 );
not ( w_8446 , w_8447 );
and ( w_8447 , \3295_b1 , \3295_b0 );
or ( \3541_b1 , \3540_b1 , \3300_b1 );
xor ( \3541_b0 , \3540_b0 , w_8448 );
not ( w_8448 , w_8449 );
and ( w_8449 , \3300_b1 , \3300_b0 );
or ( \3542_b1 , \3307_b1 , \3311_b1 );
xor ( \3542_b0 , \3307_b0 , w_8450 );
not ( w_8450 , w_8451 );
and ( w_8451 , \3311_b1 , \3311_b0 );
or ( \3543_b1 , \3542_b1 , \3316_b1 );
xor ( \3543_b0 , \3542_b0 , w_8452 );
not ( w_8452 , w_8453 );
and ( w_8453 , \3316_b1 , \3316_b0 );
or ( \3544_b1 , \3541_b1 , \3543_b1 );
not ( \3543_b1 , w_8454 );
and ( \3544_b0 , \3541_b0 , w_8455 );
and ( w_8454 , w_8455 , \3543_b0 );
or ( \3545_b1 , \3359_b1 , \3363_b1 );
xor ( \3545_b0 , \3359_b0 , w_8456 );
not ( w_8456 , w_8457 );
and ( w_8457 , \3363_b1 , \3363_b0 );
or ( \3546_b1 , \3545_b1 , \3368_b1 );
xor ( \3546_b0 , \3545_b0 , w_8458 );
not ( w_8458 , w_8459 );
and ( w_8459 , \3368_b1 , \3368_b0 );
or ( \3547_b1 , \3543_b1 , \3546_b1 );
not ( \3546_b1 , w_8460 );
and ( \3547_b0 , \3543_b0 , w_8461 );
and ( w_8460 , w_8461 , \3546_b0 );
or ( \3548_b1 , \3541_b1 , \3546_b1 );
not ( \3546_b1 , w_8462 );
and ( \3548_b0 , \3541_b0 , w_8463 );
and ( w_8462 , w_8463 , \3546_b0 );
or ( \3550_b1 , \3538_b1 , \3549_b1 );
not ( \3549_b1 , w_8464 );
and ( \3550_b0 , \3538_b0 , w_8465 );
and ( w_8464 , w_8465 , \3549_b0 );
or ( \3551_b1 , \3500_b1 , \3549_b1 );
not ( \3549_b1 , w_8466 );
and ( \3551_b0 , \3500_b0 , w_8467 );
and ( w_8466 , w_8467 , \3549_b0 );
or ( \3553_b1 , \3355_b1 , \3371_b1 );
xor ( \3553_b0 , \3355_b0 , w_8468 );
not ( w_8468 , w_8469 );
and ( w_8469 , \3371_b1 , \3371_b0 );
or ( \3554_b1 , \3553_b1 , \3376_b1 );
xor ( \3554_b0 , \3553_b0 , w_8470 );
not ( w_8470 , w_8471 );
and ( w_8471 , \3376_b1 , \3376_b0 );
or ( \3555_b1 , \3395_b1 , \3397_b1 );
xor ( \3555_b0 , \3395_b0 , w_8472 );
not ( w_8472 , w_8473 );
and ( w_8473 , \3397_b1 , \3397_b0 );
or ( \3556_b1 , \3555_b1 , \3400_b1 );
xor ( \3556_b0 , \3555_b0 , w_8474 );
not ( w_8474 , w_8475 );
and ( w_8475 , \3400_b1 , \3400_b0 );
or ( \3557_b1 , \3554_b1 , \3556_b1 );
not ( \3556_b1 , w_8476 );
and ( \3557_b0 , \3554_b0 , w_8477 );
and ( w_8476 , w_8477 , \3556_b0 );
or ( \3558_b1 , \3382_b1 , \3384_b1 );
xor ( \3558_b0 , \3382_b0 , w_8478 );
not ( w_8478 , w_8479 );
and ( w_8479 , \3384_b1 , \3384_b0 );
or ( \3559_b1 , \3558_b1 , \3387_b1 );
xor ( \3559_b0 , \3558_b0 , w_8480 );
not ( w_8480 , w_8481 );
and ( w_8481 , \3387_b1 , \3387_b0 );
or ( \3560_b1 , \3556_b1 , \3559_b1 );
not ( \3559_b1 , w_8482 );
and ( \3560_b0 , \3556_b0 , w_8483 );
and ( w_8482 , w_8483 , \3559_b0 );
or ( \3561_b1 , \3554_b1 , \3559_b1 );
not ( \3559_b1 , w_8484 );
and ( \3561_b0 , \3554_b0 , w_8485 );
and ( w_8484 , w_8485 , \3559_b0 );
or ( \3563_b1 , \3552_b1 , \3562_b1 );
not ( \3562_b1 , w_8486 );
and ( \3563_b0 , \3552_b0 , w_8487 );
and ( w_8486 , w_8487 , \3562_b0 );
or ( \3564_b1 , \3414_b1 , \3416_b1 );
xor ( \3564_b0 , \3414_b0 , w_8488 );
not ( w_8488 , w_8489 );
and ( w_8489 , \3416_b1 , \3416_b0 );
or ( \3565_b1 , \3564_b1 , \3419_b1 );
xor ( \3565_b0 , \3564_b0 , w_8490 );
not ( w_8490 , w_8491 );
and ( w_8491 , \3419_b1 , \3419_b0 );
or ( \3566_b1 , \3562_b1 , \3565_b1 );
not ( \3565_b1 , w_8492 );
and ( \3566_b0 , \3562_b0 , w_8493 );
and ( w_8492 , w_8493 , \3565_b0 );
or ( \3567_b1 , \3552_b1 , \3565_b1 );
not ( \3565_b1 , w_8494 );
and ( \3567_b0 , \3552_b0 , w_8495 );
and ( w_8494 , w_8495 , \3565_b0 );
or ( \3569_b1 , \3339_b1 , \3379_b1 );
xor ( \3569_b0 , \3339_b0 , w_8496 );
not ( w_8496 , w_8497 );
and ( w_8497 , \3379_b1 , \3379_b0 );
or ( \3570_b1 , \3569_b1 , \3390_b1 );
xor ( \3570_b0 , \3569_b0 , w_8498 );
not ( w_8498 , w_8499 );
and ( w_8499 , \3390_b1 , \3390_b0 );
or ( \3571_b1 , \3403_b1 , \3405_b1 );
xor ( \3571_b0 , \3403_b0 , w_8500 );
not ( w_8500 , w_8501 );
and ( w_8501 , \3405_b1 , \3405_b0 );
or ( \3572_b1 , \3571_b1 , \3408_b1 );
xor ( \3572_b0 , \3571_b0 , w_8502 );
not ( w_8502 , w_8503 );
and ( w_8503 , \3408_b1 , \3408_b0 );
or ( \3573_b1 , \3570_b1 , \3572_b1 );
not ( \3572_b1 , w_8504 );
and ( \3573_b0 , \3570_b0 , w_8505 );
and ( w_8504 , w_8505 , \3572_b0 );
or ( \3574_b1 , \3568_b1 , \3573_b1 );
not ( \3573_b1 , w_8506 );
and ( \3574_b0 , \3568_b0 , w_8507 );
and ( w_8506 , w_8507 , \3573_b0 );
or ( \3575_b1 , \3427_b1 , \3429_b1 );
xor ( \3575_b0 , \3427_b0 , w_8508 );
not ( w_8508 , w_8509 );
and ( w_8509 , \3429_b1 , \3429_b0 );
or ( \3576_b1 , \3575_b1 , \3431_b1 );
xor ( \3576_b0 , \3575_b0 , w_8510 );
not ( w_8510 , w_8511 );
and ( w_8511 , \3431_b1 , \3431_b0 );
or ( \3577_b1 , \3573_b1 , \3576_b1 );
not ( \3576_b1 , w_8512 );
and ( \3577_b0 , \3573_b0 , w_8513 );
and ( w_8512 , w_8513 , \3576_b0 );
or ( \3578_b1 , \3568_b1 , \3576_b1 );
not ( \3576_b1 , w_8514 );
and ( \3578_b0 , \3568_b0 , w_8515 );
and ( w_8514 , w_8515 , \3576_b0 );
or ( \3580_b1 , \3241_b1 , \3250_b1 );
xor ( \3580_b0 , \3241_b0 , w_8516 );
not ( w_8516 , w_8517 );
and ( w_8517 , \3250_b1 , \3250_b0 );
or ( \3581_b1 , \3580_b1 , \3256_b1 );
xor ( \3581_b0 , \3580_b0 , w_8518 );
not ( w_8518 , w_8519 );
and ( w_8519 , \3256_b1 , \3256_b0 );
or ( \3582_b1 , \3579_b1 , \3581_b1 );
not ( \3581_b1 , w_8520 );
and ( \3582_b0 , \3579_b0 , w_8521 );
and ( w_8520 , w_8521 , \3581_b0 );
or ( \3583_b1 , \3425_b1 , \3434_b1 );
xor ( \3583_b0 , \3425_b0 , w_8522 );
not ( w_8522 , w_8523 );
and ( w_8523 , \3434_b1 , \3434_b0 );
or ( \3584_b1 , \3583_b1 , \3437_b1 );
xor ( \3584_b0 , \3583_b0 , w_8524 );
not ( w_8524 , w_8525 );
and ( w_8525 , \3437_b1 , \3437_b0 );
or ( \3585_b1 , \3581_b1 , \3584_b1 );
not ( \3584_b1 , w_8526 );
and ( \3585_b0 , \3581_b0 , w_8527 );
and ( w_8526 , w_8527 , \3584_b0 );
or ( \3586_b1 , \3579_b1 , \3584_b1 );
not ( \3584_b1 , w_8528 );
and ( \3586_b0 , \3579_b0 , w_8529 );
and ( w_8528 , w_8529 , \3584_b0 );
or ( \3588_b1 , \3452_b1 , \3587_b1 );
not ( \3587_b1 , w_8530 );
and ( \3588_b0 , \3452_b0 , w_8531 );
and ( w_8530 , w_8531 , \3587_b0 );
or ( \3589_b1 , \3452_b1 , \3587_b1 );
xor ( \3589_b0 , \3452_b0 , w_8532 );
not ( w_8532 , w_8533 );
and ( w_8533 , \3587_b1 , \3587_b0 );
or ( \3590_b1 , \3579_b1 , \3581_b1 );
xor ( \3590_b0 , \3579_b0 , w_8534 );
not ( w_8534 , w_8535 );
and ( w_8535 , \3581_b1 , \3581_b0 );
or ( \3591_b1 , \3590_b1 , \3584_b1 );
xor ( \3591_b0 , \3590_b0 , w_8536 );
not ( w_8536 , w_8537 );
and ( w_8537 , \3584_b1 , \3584_b0 );
or ( \3592_b1 , \353_b1 , \2913_b1 );
not ( \2913_b1 , w_8538 );
and ( \3592_b0 , \353_b0 , w_8539 );
and ( w_8538 , w_8539 , \2913_b0 );
or ( \3593_b1 , \323_b1 , \2910_b1 );
not ( \2910_b1 , w_8540 );
and ( \3593_b0 , \323_b0 , w_8541 );
and ( w_8540 , w_8541 , \2910_b0 );
or ( \3594_b1 , \3592_b1 , w_8543 );
not ( w_8543 , w_8544 );
and ( \3594_b0 , \3592_b0 , w_8545 );
and ( w_8544 ,  , w_8545 );
buf ( w_8543 , \3593_b1 );
not ( w_8543 , w_8546 );
not (  , w_8547 );
and ( w_8546 , w_8547 , \3593_b0 );
or ( \3595_b1 , \3594_b1 , w_8548 );
xor ( \3595_b0 , \3594_b0 , w_8550 );
not ( w_8550 , w_8551 );
and ( w_8551 , w_8548 , w_8549 );
buf ( w_8548 , \2371_b1 );
not ( w_8548 , w_8552 );
not ( w_8549 , w_8553 );
and ( w_8552 , w_8553 , \2371_b0 );
or ( \3596_b1 , \360_b1 , \2550_b1 );
not ( \2550_b1 , w_8554 );
and ( \3596_b0 , \360_b0 , w_8555 );
and ( w_8554 , w_8555 , \2550_b0 );
or ( \3597_b1 , \343_b1 , \2548_b1 );
not ( \2548_b1 , w_8556 );
and ( \3597_b0 , \343_b0 , w_8557 );
and ( w_8556 , w_8557 , \2548_b0 );
or ( \3598_b1 , \3596_b1 , w_8559 );
not ( w_8559 , w_8560 );
and ( \3598_b0 , \3596_b0 , w_8561 );
and ( w_8560 ,  , w_8561 );
buf ( w_8559 , \3597_b1 );
not ( w_8559 , w_8562 );
not (  , w_8563 );
and ( w_8562 , w_8563 , \3597_b0 );
or ( \3599_b1 , \3598_b1 , w_8564 );
xor ( \3599_b0 , \3598_b0 , w_8566 );
not ( w_8566 , w_8567 );
and ( w_8567 , w_8564 , w_8565 );
buf ( w_8564 , \2374_b1 );
not ( w_8564 , w_8568 );
not ( w_8565 , w_8569 );
and ( w_8568 , w_8569 , \2374_b0 );
or ( \3600_b1 , \3595_b1 , \3599_b1 );
not ( \3599_b1 , w_8570 );
and ( \3600_b0 , \3595_b0 , w_8571 );
and ( w_8570 , w_8571 , \3599_b0 );
or ( \3601_b1 , \495_b1 , \2261_b1 );
not ( \2261_b1 , w_8572 );
and ( \3601_b0 , \495_b0 , w_8573 );
and ( w_8572 , w_8573 , \2261_b0 );
or ( \3602_b1 , \444_b1 , \2259_b1 );
not ( \2259_b1 , w_8574 );
and ( \3602_b0 , \444_b0 , w_8575 );
and ( w_8574 , w_8575 , \2259_b0 );
or ( \3603_b1 , \3601_b1 , w_8577 );
not ( w_8577 , w_8578 );
and ( \3603_b0 , \3601_b0 , w_8579 );
and ( w_8578 ,  , w_8579 );
buf ( w_8577 , \3602_b1 );
not ( w_8577 , w_8580 );
not (  , w_8581 );
and ( w_8580 , w_8581 , \3602_b0 );
or ( \3604_b1 , \3603_b1 , w_8582 );
xor ( \3604_b0 , \3603_b0 , w_8584 );
not ( w_8584 , w_8585 );
and ( w_8585 , w_8582 , w_8583 );
buf ( w_8582 , \2124_b1 );
not ( w_8582 , w_8586 );
not ( w_8583 , w_8587 );
and ( w_8586 , w_8587 , \2124_b0 );
or ( \3605_b1 , \3599_b1 , \3604_b1 );
not ( \3604_b1 , w_8588 );
and ( \3605_b0 , \3599_b0 , w_8589 );
and ( w_8588 , w_8589 , \3604_b0 );
or ( \3606_b1 , \3595_b1 , \3604_b1 );
not ( \3604_b1 , w_8590 );
and ( \3606_b0 , \3595_b0 , w_8591 );
and ( w_8590 , w_8591 , \3604_b0 );
or ( \3608_b1 , \1194_b1 , \1280_b1 );
not ( \1280_b1 , w_8592 );
and ( \3608_b0 , \1194_b0 , w_8593 );
and ( w_8592 , w_8593 , \1280_b0 );
or ( \3609_b1 , \1104_b1 , \1278_b1 );
not ( \1278_b1 , w_8594 );
and ( \3609_b0 , \1104_b0 , w_8595 );
and ( w_8594 , w_8595 , \1278_b0 );
or ( \3610_b1 , \3608_b1 , w_8597 );
not ( w_8597 , w_8598 );
and ( \3610_b0 , \3608_b0 , w_8599 );
and ( w_8598 ,  , w_8599 );
buf ( w_8597 , \3609_b1 );
not ( w_8597 , w_8600 );
not (  , w_8601 );
and ( w_8600 , w_8601 , \3609_b0 );
or ( \3611_b1 , \3610_b1 , w_8602 );
xor ( \3611_b0 , \3610_b0 , w_8604 );
not ( w_8604 , w_8605 );
and ( w_8605 , w_8602 , w_8603 );
buf ( w_8602 , \1177_b1 );
not ( w_8602 , w_8606 );
not ( w_8603 , w_8607 );
and ( w_8606 , w_8607 , \1177_b0 );
or ( \3612_b1 , \1304_b1 , \1062_b1 );
not ( \1062_b1 , w_8608 );
and ( \3612_b0 , \1304_b0 , w_8609 );
and ( w_8608 , w_8609 , \1062_b0 );
or ( \3613_b1 , \1299_b1 , \1060_b1 );
not ( \1060_b1 , w_8610 );
and ( \3613_b0 , \1299_b0 , w_8611 );
and ( w_8610 , w_8611 , \1060_b0 );
or ( \3614_b1 , \3612_b1 , w_8613 );
not ( w_8613 , w_8614 );
and ( \3614_b0 , \3612_b0 , w_8615 );
and ( w_8614 ,  , w_8615 );
buf ( w_8613 , \3613_b1 );
not ( w_8613 , w_8616 );
not (  , w_8617 );
and ( w_8616 , w_8617 , \3613_b0 );
or ( \3615_b1 , \3614_b1 , w_8618 );
xor ( \3615_b0 , \3614_b0 , w_8620 );
not ( w_8620 , w_8621 );
and ( w_8621 , w_8618 , w_8619 );
buf ( w_8618 , \984_b1 );
not ( w_8618 , w_8622 );
not ( w_8619 , w_8623 );
and ( w_8622 , w_8623 , \984_b0 );
or ( \3616_b1 , \3611_b1 , \3615_b1 );
not ( \3615_b1 , w_8624 );
and ( \3616_b0 , \3611_b0 , w_8625 );
and ( w_8624 , w_8625 , \3615_b0 );
or ( \3617_b1 , \1537_b1 , \912_b1 );
not ( \912_b1 , w_8626 );
and ( \3617_b0 , \1537_b0 , w_8627 );
and ( w_8626 , w_8627 , \912_b0 );
or ( \3618_b1 , \1422_b1 , \910_b1 );
not ( \910_b1 , w_8628 );
and ( \3618_b0 , \1422_b0 , w_8629 );
and ( w_8628 , w_8629 , \910_b0 );
or ( \3619_b1 , \3617_b1 , w_8631 );
not ( w_8631 , w_8632 );
and ( \3619_b0 , \3617_b0 , w_8633 );
and ( w_8632 ,  , w_8633 );
buf ( w_8631 , \3618_b1 );
not ( w_8631 , w_8634 );
not (  , w_8635 );
and ( w_8634 , w_8635 , \3618_b0 );
or ( \3620_b1 , \3619_b1 , w_8636 );
xor ( \3620_b0 , \3619_b0 , w_8638 );
not ( w_8638 , w_8639 );
and ( w_8639 , w_8636 , w_8637 );
buf ( w_8636 , \818_b1 );
not ( w_8636 , w_8640 );
not ( w_8637 , w_8641 );
and ( w_8640 , w_8641 , \818_b0 );
or ( \3621_b1 , \3615_b1 , \3620_b1 );
not ( \3620_b1 , w_8642 );
and ( \3621_b0 , \3615_b0 , w_8643 );
and ( w_8642 , w_8643 , \3620_b0 );
or ( \3622_b1 , \3611_b1 , \3620_b1 );
not ( \3620_b1 , w_8644 );
and ( \3622_b0 , \3611_b0 , w_8645 );
and ( w_8644 , w_8645 , \3620_b0 );
or ( \3624_b1 , \3607_b1 , \3623_b1 );
not ( \3623_b1 , w_8646 );
and ( \3624_b0 , \3607_b0 , w_8647 );
and ( w_8646 , w_8647 , \3623_b0 );
or ( \3625_b1 , \621_b1 , \1955_b1 );
not ( \1955_b1 , w_8648 );
and ( \3625_b0 , \621_b0 , w_8649 );
and ( w_8648 , w_8649 , \1955_b0 );
or ( \3626_b1 , \593_b1 , \1953_b1 );
not ( \1953_b1 , w_8650 );
and ( \3626_b0 , \593_b0 , w_8651 );
and ( w_8650 , w_8651 , \1953_b0 );
or ( \3627_b1 , \3625_b1 , w_8653 );
not ( w_8653 , w_8654 );
and ( \3627_b0 , \3625_b0 , w_8655 );
and ( w_8654 ,  , w_8655 );
buf ( w_8653 , \3626_b1 );
not ( w_8653 , w_8656 );
not (  , w_8657 );
and ( w_8656 , w_8657 , \3626_b0 );
or ( \3628_b1 , \3627_b1 , w_8658 );
xor ( \3628_b0 , \3627_b0 , w_8660 );
not ( w_8660 , w_8661 );
and ( w_8661 , w_8658 , w_8659 );
buf ( w_8658 , \1835_b1 );
not ( w_8658 , w_8662 );
not ( w_8659 , w_8663 );
and ( w_8662 , w_8663 , \1835_b0 );
or ( \3629_b1 , \777_b1 , \1742_b1 );
not ( \1742_b1 , w_8664 );
and ( \3629_b0 , \777_b0 , w_8665 );
and ( w_8664 , w_8665 , \1742_b0 );
or ( \3630_b1 , \703_b1 , \1740_b1 );
not ( \1740_b1 , w_8666 );
and ( \3630_b0 , \703_b0 , w_8667 );
and ( w_8666 , w_8667 , \1740_b0 );
or ( \3631_b1 , \3629_b1 , w_8669 );
not ( w_8669 , w_8670 );
and ( \3631_b0 , \3629_b0 , w_8671 );
and ( w_8670 ,  , w_8671 );
buf ( w_8669 , \3630_b1 );
not ( w_8669 , w_8672 );
not (  , w_8673 );
and ( w_8672 , w_8673 , \3630_b0 );
or ( \3632_b1 , \3631_b1 , w_8674 );
xor ( \3632_b0 , \3631_b0 , w_8676 );
not ( w_8676 , w_8677 );
and ( w_8677 , w_8674 , w_8675 );
buf ( w_8674 , \1610_b1 );
not ( w_8674 , w_8678 );
not ( w_8675 , w_8679 );
and ( w_8678 , w_8679 , \1610_b0 );
or ( \3633_b1 , \3628_b1 , \3632_b1 );
not ( \3632_b1 , w_8680 );
and ( \3633_b0 , \3628_b0 , w_8681 );
and ( w_8680 , w_8681 , \3632_b0 );
or ( \3634_b1 , \904_b1 , \1476_b1 );
not ( \1476_b1 , w_8682 );
and ( \3634_b0 , \904_b0 , w_8683 );
and ( w_8682 , w_8683 , \1476_b0 );
or ( \3635_b1 , \841_b1 , \1474_b1 );
not ( \1474_b1 , w_8684 );
and ( \3635_b0 , \841_b0 , w_8685 );
and ( w_8684 , w_8685 , \1474_b0 );
or ( \3636_b1 , \3634_b1 , w_8687 );
not ( w_8687 , w_8688 );
and ( \3636_b0 , \3634_b0 , w_8689 );
and ( w_8688 ,  , w_8689 );
buf ( w_8687 , \3635_b1 );
not ( w_8687 , w_8690 );
not (  , w_8691 );
and ( w_8690 , w_8691 , \3635_b0 );
or ( \3637_b1 , \3636_b1 , w_8692 );
xor ( \3637_b0 , \3636_b0 , w_8694 );
not ( w_8694 , w_8695 );
and ( w_8695 , w_8692 , w_8693 );
buf ( w_8692 , \1363_b1 );
not ( w_8692 , w_8696 );
not ( w_8693 , w_8697 );
and ( w_8696 , w_8697 , \1363_b0 );
or ( \3638_b1 , \3632_b1 , \3637_b1 );
not ( \3637_b1 , w_8698 );
and ( \3638_b0 , \3632_b0 , w_8699 );
and ( w_8698 , w_8699 , \3637_b0 );
or ( \3639_b1 , \3628_b1 , \3637_b1 );
not ( \3637_b1 , w_8700 );
and ( \3639_b0 , \3628_b0 , w_8701 );
and ( w_8700 , w_8701 , \3637_b0 );
or ( \3641_b1 , \3623_b1 , \3640_b1 );
not ( \3640_b1 , w_8702 );
and ( \3641_b0 , \3623_b0 , w_8703 );
and ( w_8702 , w_8703 , \3640_b0 );
or ( \3642_b1 , \3607_b1 , \3640_b1 );
not ( \3640_b1 , w_8704 );
and ( \3642_b0 , \3607_b0 , w_8705 );
and ( w_8704 , w_8705 , \3640_b0 );
or ( \3644_b1 , \3456_b1 , \3460_b1 );
xor ( \3644_b0 , \3456_b0 , w_8706 );
not ( w_8706 , w_8707 );
and ( w_8707 , \3460_b1 , \3460_b0 );
or ( \3645_b1 , \3644_b1 , \3465_b1 );
xor ( \3645_b0 , \3644_b0 , w_8708 );
not ( w_8708 , w_8709 );
and ( w_8709 , \3465_b1 , \3465_b0 );
or ( \3646_b1 , \3472_b1 , \3476_b1 );
xor ( \3646_b0 , \3472_b0 , w_8710 );
not ( w_8710 , w_8711 );
and ( w_8711 , \3476_b1 , \3476_b0 );
or ( \3647_b1 , \3646_b1 , \3481_b1 );
xor ( \3647_b0 , \3646_b0 , w_8712 );
not ( w_8712 , w_8713 );
and ( w_8713 , \3481_b1 , \3481_b0 );
or ( \3648_b1 , \3645_b1 , \3647_b1 );
not ( \3647_b1 , w_8714 );
and ( \3648_b0 , \3645_b0 , w_8715 );
and ( w_8714 , w_8715 , \3647_b0 );
or ( \3649_b1 , \3504_b1 , \3508_b1 );
xor ( \3649_b0 , \3504_b0 , w_8716 );
not ( w_8716 , w_8717 );
and ( w_8717 , \3508_b1 , \3508_b0 );
or ( \3650_b1 , \3649_b1 , \3513_b1 );
xor ( \3650_b0 , \3649_b0 , w_8718 );
not ( w_8718 , w_8719 );
and ( w_8719 , \3513_b1 , \3513_b0 );
or ( \3651_b1 , \3647_b1 , \3650_b1 );
not ( \3650_b1 , w_8720 );
and ( \3651_b0 , \3647_b0 , w_8721 );
and ( w_8720 , w_8721 , \3650_b0 );
or ( \3652_b1 , \3645_b1 , \3650_b1 );
not ( \3650_b1 , w_8722 );
and ( \3652_b0 , \3645_b0 , w_8723 );
and ( w_8722 , w_8723 , \3650_b0 );
or ( \3654_b1 , \3643_b1 , \3653_b1 );
not ( \3653_b1 , w_8724 );
and ( \3654_b0 , \3643_b0 , w_8725 );
and ( w_8724 , w_8725 , \3653_b0 );
or ( \3655_b1 , \1778_b1 , \740_b1 );
not ( \740_b1 , w_8726 );
and ( \3655_b0 , \1778_b0 , w_8727 );
and ( w_8726 , w_8727 , \740_b0 );
or ( \3656_b1 , \1770_b1 , \738_b1 );
not ( \738_b1 , w_8728 );
and ( \3656_b0 , \1770_b0 , w_8729 );
and ( w_8728 , w_8729 , \738_b0 );
or ( \3657_b1 , \3655_b1 , w_8731 );
not ( w_8731 , w_8732 );
and ( \3657_b0 , \3655_b0 , w_8733 );
and ( w_8732 ,  , w_8733 );
buf ( w_8731 , \3656_b1 );
not ( w_8731 , w_8734 );
not (  , w_8735 );
and ( w_8734 , w_8735 , \3656_b0 );
or ( \3658_b1 , \3657_b1 , w_8736 );
xor ( \3658_b0 , \3657_b0 , w_8738 );
not ( w_8738 , w_8739 );
and ( w_8739 , w_8736 , w_8737 );
buf ( w_8736 , \668_b1 );
not ( w_8736 , w_8740 );
not ( w_8737 , w_8741 );
and ( w_8740 , w_8741 , \668_b0 );
or ( \3659_b1 , \2028_b1 , \604_b1 );
not ( \604_b1 , w_8742 );
and ( \3659_b0 , \2028_b0 , w_8743 );
and ( w_8742 , w_8743 , \604_b0 );
or ( \3660_b1 , \2023_b1 , \602_b1 );
not ( \602_b1 , w_8744 );
and ( \3660_b0 , \2023_b0 , w_8745 );
and ( w_8744 , w_8745 , \602_b0 );
or ( \3661_b1 , \3659_b1 , w_8747 );
not ( w_8747 , w_8748 );
and ( \3661_b0 , \3659_b0 , w_8749 );
and ( w_8748 ,  , w_8749 );
buf ( w_8747 , \3660_b1 );
not ( w_8747 , w_8750 );
not (  , w_8751 );
and ( w_8750 , w_8751 , \3660_b0 );
or ( \3662_b1 , \3661_b1 , w_8752 );
xor ( \3662_b0 , \3661_b0 , w_8754 );
not ( w_8754 , w_8755 );
and ( w_8755 , w_8752 , w_8753 );
buf ( w_8752 , \561_b1 );
not ( w_8752 , w_8756 );
not ( w_8753 , w_8757 );
and ( w_8756 , w_8757 , \561_b0 );
or ( \3663_b1 , \3658_b1 , \3662_b1 );
not ( \3662_b1 , w_8758 );
and ( \3663_b0 , \3658_b0 , w_8759 );
and ( w_8758 , w_8759 , \3662_b0 );
or ( \3664_b1 , \2305_b1 , \503_b1 );
not ( \503_b1 , w_8760 );
and ( \3664_b0 , \2305_b0 , w_8761 );
and ( w_8760 , w_8761 , \503_b0 );
or ( \3665_b1 , \2161_b1 , \501_b1 );
not ( \501_b1 , w_8762 );
and ( \3665_b0 , \2161_b0 , w_8763 );
and ( w_8762 , w_8763 , \501_b0 );
or ( \3666_b1 , \3664_b1 , w_8765 );
not ( w_8765 , w_8766 );
and ( \3666_b0 , \3664_b0 , w_8767 );
and ( w_8766 ,  , w_8767 );
buf ( w_8765 , \3665_b1 );
not ( w_8765 , w_8768 );
not (  , w_8769 );
and ( w_8768 , w_8769 , \3665_b0 );
or ( \3667_b1 , \3666_b1 , w_8770 );
xor ( \3667_b0 , \3666_b0 , w_8772 );
not ( w_8772 , w_8773 );
and ( w_8773 , w_8770 , w_8771 );
buf ( w_8770 , \455_b1 );
not ( w_8770 , w_8774 );
not ( w_8771 , w_8775 );
and ( w_8774 , w_8775 , \455_b0 );
or ( \3668_b1 , \3662_b1 , \3667_b1 );
not ( \3667_b1 , w_8776 );
and ( \3668_b0 , \3662_b0 , w_8777 );
and ( w_8776 , w_8777 , \3667_b0 );
or ( \3669_b1 , \3658_b1 , \3667_b1 );
not ( \3667_b1 , w_8778 );
and ( \3669_b0 , \3658_b0 , w_8779 );
and ( w_8778 , w_8779 , \3667_b0 );
or ( \3671_b1 , \2850_b1 , w_8781 );
not ( w_8781 , w_8782 );
and ( \3671_b0 , \2850_b0 , w_8783 );
and ( w_8782 ,  , w_8783 );
buf ( w_8781 , \329_b1 );
not ( w_8781 , w_8784 );
not (  , w_8785 );
and ( w_8784 , w_8785 , \329_b0 );
or ( \3672_b1 , \3671_b1 , w_8786 );
xor ( \3672_b0 , \3671_b0 , w_8788 );
not ( w_8788 , w_8789 );
and ( w_8789 , w_8786 , w_8787 );
buf ( w_8786 , \338_b1 );
not ( w_8786 , w_8790 );
not ( w_8787 , w_8791 );
and ( w_8790 , w_8791 , \338_b0 );
or ( \3673_b1 , \3670_b1 , \3672_b1 );
not ( \3672_b1 , w_8792 );
and ( \3673_b0 , \3670_b0 , w_8793 );
and ( w_8792 , w_8793 , \3672_b0 );
or ( \3674_b1 , \3520_b1 , \3524_b1 );
xor ( \3674_b0 , \3520_b0 , w_8794 );
not ( w_8794 , w_8795 );
and ( w_8795 , \3524_b1 , \3524_b0 );
or ( \3675_b1 , \3674_b1 , \3529_b1 );
xor ( \3675_b0 , \3674_b0 , w_8796 );
not ( w_8796 , w_8797 );
and ( w_8797 , \3529_b1 , \3529_b0 );
or ( \3676_b1 , \3672_b1 , \3675_b1 );
not ( \3675_b1 , w_8798 );
and ( \3676_b0 , \3672_b0 , w_8799 );
and ( w_8798 , w_8799 , \3675_b0 );
or ( \3677_b1 , \3670_b1 , \3675_b1 );
not ( \3675_b1 , w_8800 );
and ( \3677_b0 , \3670_b0 , w_8801 );
and ( w_8800 , w_8801 , \3675_b0 );
or ( \3679_b1 , \3653_b1 , \3678_b1 );
not ( \3678_b1 , w_8802 );
and ( \3679_b0 , \3653_b0 , w_8803 );
and ( w_8802 , w_8803 , \3678_b0 );
or ( \3680_b1 , \3643_b1 , \3678_b1 );
not ( \3678_b1 , w_8804 );
and ( \3680_b0 , \3643_b0 , w_8805 );
and ( w_8804 , w_8805 , \3678_b0 );
or ( \3682_b1 , \3324_b1 , \3328_b1 );
xor ( \3682_b0 , \3324_b0 , w_8806 );
not ( w_8806 , w_8807 );
and ( w_8807 , \3328_b1 , \3328_b0 );
or ( \3683_b1 , \3682_b1 , \3333_b1 );
xor ( \3683_b0 , \3682_b0 , w_8808 );
not ( w_8808 , w_8809 );
and ( w_8809 , \3333_b1 , \3333_b0 );
or ( \3684_b1 , \3516_b1 , \3532_b1 );
xor ( \3684_b0 , \3516_b0 , w_8810 );
not ( w_8810 , w_8811 );
and ( w_8811 , \3532_b1 , \3532_b0 );
or ( \3685_b1 , \3684_b1 , \3535_b1 );
xor ( \3685_b0 , \3684_b0 , w_8812 );
not ( w_8812 , w_8813 );
and ( w_8813 , \3535_b1 , \3535_b0 );
or ( \3686_b1 , \3683_b1 , \3685_b1 );
not ( \3685_b1 , w_8814 );
and ( \3686_b0 , \3683_b0 , w_8815 );
and ( w_8814 , w_8815 , \3685_b0 );
or ( \3687_b1 , \3541_b1 , \3543_b1 );
xor ( \3687_b0 , \3541_b0 , w_8816 );
not ( w_8816 , w_8817 );
and ( w_8817 , \3543_b1 , \3543_b0 );
or ( \3688_b1 , \3687_b1 , \3546_b1 );
xor ( \3688_b0 , \3687_b0 , w_8818 );
not ( w_8818 , w_8819 );
and ( w_8819 , \3546_b1 , \3546_b0 );
or ( \3689_b1 , \3685_b1 , \3688_b1 );
not ( \3688_b1 , w_8820 );
and ( \3689_b0 , \3685_b0 , w_8821 );
and ( w_8820 , w_8821 , \3688_b0 );
or ( \3690_b1 , \3683_b1 , \3688_b1 );
not ( \3688_b1 , w_8822 );
and ( \3690_b0 , \3683_b0 , w_8823 );
and ( w_8822 , w_8823 , \3688_b0 );
or ( \3692_b1 , \3681_b1 , \3691_b1 );
not ( \3691_b1 , w_8824 );
and ( \3692_b0 , \3681_b0 , w_8825 );
and ( w_8824 , w_8825 , \3691_b0 );
or ( \3693_b1 , \3303_b1 , \3319_b1 );
xor ( \3693_b0 , \3303_b0 , w_8826 );
not ( w_8826 , w_8827 );
and ( w_8827 , \3319_b1 , \3319_b0 );
or ( \3694_b1 , \3693_b1 , \3336_b1 );
xor ( \3694_b0 , \3693_b0 , w_8828 );
not ( w_8828 , w_8829 );
and ( w_8829 , \3336_b1 , \3336_b0 );
or ( \3695_b1 , \3691_b1 , \3694_b1 );
not ( \3694_b1 , w_8830 );
and ( \3695_b0 , \3691_b0 , w_8831 );
and ( w_8830 , w_8831 , \3694_b0 );
or ( \3696_b1 , \3681_b1 , \3694_b1 );
not ( \3694_b1 , w_8832 );
and ( \3696_b0 , \3681_b0 , w_8833 );
and ( w_8832 , w_8833 , \3694_b0 );
or ( \3698_b1 , \3552_b1 , \3562_b1 );
xor ( \3698_b0 , \3552_b0 , w_8834 );
not ( w_8834 , w_8835 );
and ( w_8835 , \3562_b1 , \3562_b0 );
or ( \3699_b1 , \3698_b1 , \3565_b1 );
xor ( \3699_b0 , \3698_b0 , w_8836 );
not ( w_8836 , w_8837 );
and ( w_8837 , \3565_b1 , \3565_b0 );
or ( \3700_b1 , \3697_b1 , \3699_b1 );
not ( \3699_b1 , w_8838 );
and ( \3700_b0 , \3697_b0 , w_8839 );
and ( w_8838 , w_8839 , \3699_b0 );
or ( \3701_b1 , \3570_b1 , \3572_b1 );
xor ( \3701_b0 , \3570_b0 , w_8840 );
not ( w_8840 , w_8841 );
and ( w_8841 , \3572_b1 , \3572_b0 );
or ( \3702_b1 , \3699_b1 , \3701_b1 );
not ( \3701_b1 , w_8842 );
and ( \3702_b0 , \3699_b0 , w_8843 );
and ( w_8842 , w_8843 , \3701_b0 );
or ( \3703_b1 , \3697_b1 , \3701_b1 );
not ( \3701_b1 , w_8844 );
and ( \3703_b0 , \3697_b0 , w_8845 );
and ( w_8844 , w_8845 , \3701_b0 );
or ( \3705_b1 , \3393_b1 , \3411_b1 );
xor ( \3705_b0 , \3393_b0 , w_8846 );
not ( w_8846 , w_8847 );
and ( w_8847 , \3411_b1 , \3411_b0 );
or ( \3706_b1 , \3705_b1 , \3422_b1 );
xor ( \3706_b0 , \3705_b0 , w_8848 );
not ( w_8848 , w_8849 );
and ( w_8849 , \3422_b1 , \3422_b0 );
or ( \3707_b1 , \3704_b1 , \3706_b1 );
not ( \3706_b1 , w_8850 );
and ( \3707_b0 , \3704_b0 , w_8851 );
and ( w_8850 , w_8851 , \3706_b0 );
or ( \3708_b1 , \3568_b1 , \3573_b1 );
xor ( \3708_b0 , \3568_b0 , w_8852 );
not ( w_8852 , w_8853 );
and ( w_8853 , \3573_b1 , \3573_b0 );
or ( \3709_b1 , \3708_b1 , \3576_b1 );
xor ( \3709_b0 , \3708_b0 , w_8854 );
not ( w_8854 , w_8855 );
and ( w_8855 , \3576_b1 , \3576_b0 );
or ( \3710_b1 , \3706_b1 , \3709_b1 );
not ( \3709_b1 , w_8856 );
and ( \3710_b0 , \3706_b0 , w_8857 );
and ( w_8856 , w_8857 , \3709_b0 );
or ( \3711_b1 , \3704_b1 , \3709_b1 );
not ( \3709_b1 , w_8858 );
and ( \3711_b0 , \3704_b0 , w_8859 );
and ( w_8858 , w_8859 , \3709_b0 );
or ( \3713_b1 , \3591_b1 , \3712_b1 );
not ( \3712_b1 , w_8860 );
and ( \3713_b0 , \3591_b0 , w_8861 );
and ( w_8860 , w_8861 , \3712_b0 );
or ( \3714_b1 , \3591_b1 , \3712_b1 );
xor ( \3714_b0 , \3591_b0 , w_8862 );
not ( w_8862 , w_8863 );
and ( w_8863 , \3712_b1 , \3712_b0 );
or ( \3715_b1 , \3704_b1 , \3706_b1 );
xor ( \3715_b0 , \3704_b0 , w_8864 );
not ( w_8864 , w_8865 );
and ( w_8865 , \3706_b1 , \3706_b0 );
or ( \3716_b1 , \3715_b1 , \3709_b1 );
xor ( \3716_b0 , \3715_b0 , w_8866 );
not ( w_8866 , w_8867 );
and ( w_8867 , \3709_b1 , \3709_b0 );
or ( \3717_b1 , \1770_b1 , \912_b1 );
not ( \912_b1 , w_8868 );
and ( \3717_b0 , \1770_b0 , w_8869 );
and ( w_8868 , w_8869 , \912_b0 );
or ( \3718_b1 , \1537_b1 , \910_b1 );
not ( \910_b1 , w_8870 );
and ( \3718_b0 , \1537_b0 , w_8871 );
and ( w_8870 , w_8871 , \910_b0 );
or ( \3719_b1 , \3717_b1 , w_8873 );
not ( w_8873 , w_8874 );
and ( \3719_b0 , \3717_b0 , w_8875 );
and ( w_8874 ,  , w_8875 );
buf ( w_8873 , \3718_b1 );
not ( w_8873 , w_8876 );
not (  , w_8877 );
and ( w_8876 , w_8877 , \3718_b0 );
or ( \3720_b1 , \3719_b1 , w_8878 );
xor ( \3720_b0 , \3719_b0 , w_8880 );
not ( w_8880 , w_8881 );
and ( w_8881 , w_8878 , w_8879 );
buf ( w_8878 , \818_b1 );
not ( w_8878 , w_8882 );
not ( w_8879 , w_8883 );
and ( w_8882 , w_8883 , \818_b0 );
or ( \3721_b1 , \2023_b1 , \740_b1 );
not ( \740_b1 , w_8884 );
and ( \3721_b0 , \2023_b0 , w_8885 );
and ( w_8884 , w_8885 , \740_b0 );
or ( \3722_b1 , \1778_b1 , \738_b1 );
not ( \738_b1 , w_8886 );
and ( \3722_b0 , \1778_b0 , w_8887 );
and ( w_8886 , w_8887 , \738_b0 );
or ( \3723_b1 , \3721_b1 , w_8889 );
not ( w_8889 , w_8890 );
and ( \3723_b0 , \3721_b0 , w_8891 );
and ( w_8890 ,  , w_8891 );
buf ( w_8889 , \3722_b1 );
not ( w_8889 , w_8892 );
not (  , w_8893 );
and ( w_8892 , w_8893 , \3722_b0 );
or ( \3724_b1 , \3723_b1 , w_8894 );
xor ( \3724_b0 , \3723_b0 , w_8896 );
not ( w_8896 , w_8897 );
and ( w_8897 , w_8894 , w_8895 );
buf ( w_8894 , \668_b1 );
not ( w_8894 , w_8898 );
not ( w_8895 , w_8899 );
and ( w_8898 , w_8899 , \668_b0 );
or ( \3725_b1 , \3720_b1 , \3724_b1 );
not ( \3724_b1 , w_8900 );
and ( \3725_b0 , \3720_b0 , w_8901 );
and ( w_8900 , w_8901 , \3724_b0 );
or ( \3726_b1 , \2161_b1 , \604_b1 );
not ( \604_b1 , w_8902 );
and ( \3726_b0 , \2161_b0 , w_8903 );
and ( w_8902 , w_8903 , \604_b0 );
or ( \3727_b1 , \2028_b1 , \602_b1 );
not ( \602_b1 , w_8904 );
and ( \3727_b0 , \2028_b0 , w_8905 );
and ( w_8904 , w_8905 , \602_b0 );
or ( \3728_b1 , \3726_b1 , w_8907 );
not ( w_8907 , w_8908 );
and ( \3728_b0 , \3726_b0 , w_8909 );
and ( w_8908 ,  , w_8909 );
buf ( w_8907 , \3727_b1 );
not ( w_8907 , w_8910 );
not (  , w_8911 );
and ( w_8910 , w_8911 , \3727_b0 );
or ( \3729_b1 , \3728_b1 , w_8912 );
xor ( \3729_b0 , \3728_b0 , w_8914 );
not ( w_8914 , w_8915 );
and ( w_8915 , w_8912 , w_8913 );
buf ( w_8912 , \561_b1 );
not ( w_8912 , w_8916 );
not ( w_8913 , w_8917 );
and ( w_8916 , w_8917 , \561_b0 );
or ( \3730_b1 , \3724_b1 , \3729_b1 );
not ( \3729_b1 , w_8918 );
and ( \3730_b0 , \3724_b0 , w_8919 );
and ( w_8918 , w_8919 , \3729_b0 );
or ( \3731_b1 , \3720_b1 , \3729_b1 );
not ( \3729_b1 , w_8920 );
and ( \3731_b0 , \3720_b0 , w_8921 );
and ( w_8920 , w_8921 , \3729_b0 );
or ( \3733_b1 , \2532_b1 , \503_b1 );
not ( \503_b1 , w_8922 );
and ( \3733_b0 , \2532_b0 , w_8923 );
and ( w_8922 , w_8923 , \503_b0 );
or ( \3734_b1 , \2305_b1 , \501_b1 );
not ( \501_b1 , w_8924 );
and ( \3734_b0 , \2305_b0 , w_8925 );
and ( w_8924 , w_8925 , \501_b0 );
or ( \3735_b1 , \3733_b1 , w_8927 );
not ( w_8927 , w_8928 );
and ( \3735_b0 , \3733_b0 , w_8929 );
and ( w_8928 ,  , w_8929 );
buf ( w_8927 , \3734_b1 );
not ( w_8927 , w_8930 );
not (  , w_8931 );
and ( w_8930 , w_8931 , \3734_b0 );
or ( \3736_b1 , \3735_b1 , w_8932 );
xor ( \3736_b0 , \3735_b0 , w_8934 );
not ( w_8934 , w_8935 );
and ( w_8935 , w_8932 , w_8933 );
buf ( w_8932 , \455_b1 );
not ( w_8932 , w_8936 );
not ( w_8933 , w_8937 );
and ( w_8936 , w_8937 , \455_b0 );
or ( \3737_b1 , \2763_b1 , \298_b1 );
not ( \298_b1 , w_8938 );
and ( \3737_b0 , \2763_b0 , w_8939 );
and ( w_8938 , w_8939 , \298_b0 );
or ( \3738_b1 , \2541_b1 , \296_b1 );
not ( \296_b1 , w_8940 );
and ( \3738_b0 , \2541_b0 , w_8941 );
and ( w_8940 , w_8941 , \296_b0 );
or ( \3739_b1 , \3737_b1 , w_8943 );
not ( w_8943 , w_8944 );
and ( \3739_b0 , \3737_b0 , w_8945 );
and ( w_8944 ,  , w_8945 );
buf ( w_8943 , \3738_b1 );
not ( w_8943 , w_8946 );
not (  , w_8947 );
and ( w_8946 , w_8947 , \3738_b0 );
or ( \3740_b1 , \3739_b1 , w_8948 );
xor ( \3740_b0 , \3739_b0 , w_8950 );
not ( w_8950 , w_8951 );
and ( w_8951 , w_8948 , w_8949 );
buf ( w_8948 , \303_b1 );
not ( w_8948 , w_8952 );
not ( w_8949 , w_8953 );
and ( w_8952 , w_8953 , \303_b0 );
or ( \3741_b1 , \3736_b1 , \3740_b1 );
not ( \3740_b1 , w_8954 );
and ( \3741_b0 , \3736_b0 , w_8955 );
and ( w_8954 , w_8955 , \3740_b0 );
or ( \3742_b1 , \2850_b1 , w_8957 );
not ( w_8957 , w_8958 );
and ( \3742_b0 , \2850_b0 , w_8959 );
and ( w_8958 ,  , w_8959 );
buf ( w_8957 , \311_b1 );
not ( w_8957 , w_8960 );
not (  , w_8961 );
and ( w_8960 , w_8961 , \311_b0 );
or ( \3743_b1 , \3742_b1 , w_8962 );
xor ( \3743_b0 , \3742_b0 , w_8964 );
not ( w_8964 , w_8965 );
and ( w_8965 , w_8962 , w_8963 );
buf ( w_8962 , \320_b1 );
not ( w_8962 , w_8966 );
not ( w_8963 , w_8967 );
and ( w_8966 , w_8967 , \320_b0 );
or ( \3744_b1 , \3740_b1 , \3743_b1 );
not ( \3743_b1 , w_8968 );
and ( \3744_b0 , \3740_b0 , w_8969 );
and ( w_8968 , w_8969 , \3743_b0 );
or ( \3745_b1 , \3736_b1 , \3743_b1 );
not ( \3743_b1 , w_8970 );
and ( \3745_b0 , \3736_b0 , w_8971 );
and ( w_8970 , w_8971 , \3743_b0 );
or ( \3747_b1 , \3732_b1 , \3746_b1 );
not ( \3746_b1 , w_8972 );
and ( \3747_b0 , \3732_b0 , w_8973 );
and ( w_8972 , w_8973 , \3746_b0 );
or ( \3748_b1 , \2541_b1 , \298_b1 );
not ( \298_b1 , w_8974 );
and ( \3748_b0 , \2541_b0 , w_8975 );
and ( w_8974 , w_8975 , \298_b0 );
or ( \3749_b1 , \2532_b1 , \296_b1 );
not ( \296_b1 , w_8976 );
and ( \3749_b0 , \2532_b0 , w_8977 );
and ( w_8976 , w_8977 , \296_b0 );
or ( \3750_b1 , \3748_b1 , w_8979 );
not ( w_8979 , w_8980 );
and ( \3750_b0 , \3748_b0 , w_8981 );
and ( w_8980 ,  , w_8981 );
buf ( w_8979 , \3749_b1 );
not ( w_8979 , w_8982 );
not (  , w_8983 );
and ( w_8982 , w_8983 , \3749_b0 );
or ( \3751_b1 , \3750_b1 , w_8984 );
xor ( \3751_b0 , \3750_b0 , w_8986 );
not ( w_8986 , w_8987 );
and ( w_8987 , w_8984 , w_8985 );
buf ( w_8984 , \303_b1 );
not ( w_8984 , w_8988 );
not ( w_8985 , w_8989 );
and ( w_8988 , w_8989 , \303_b0 );
or ( \3752_b1 , \3746_b1 , \3751_b1 );
not ( \3751_b1 , w_8990 );
and ( \3752_b0 , \3746_b0 , w_8991 );
and ( w_8990 , w_8991 , \3751_b0 );
or ( \3753_b1 , \3732_b1 , \3751_b1 );
not ( \3751_b1 , w_8992 );
and ( \3753_b0 , \3732_b0 , w_8993 );
and ( w_8992 , w_8993 , \3751_b0 );
or ( \3755_b1 , \1104_b1 , \1476_b1 );
not ( \1476_b1 , w_8994 );
and ( \3755_b0 , \1104_b0 , w_8995 );
and ( w_8994 , w_8995 , \1476_b0 );
or ( \3756_b1 , \904_b1 , \1474_b1 );
not ( \1474_b1 , w_8996 );
and ( \3756_b0 , \904_b0 , w_8997 );
and ( w_8996 , w_8997 , \1474_b0 );
or ( \3757_b1 , \3755_b1 , w_8999 );
not ( w_8999 , w_9000 );
and ( \3757_b0 , \3755_b0 , w_9001 );
and ( w_9000 ,  , w_9001 );
buf ( w_8999 , \3756_b1 );
not ( w_8999 , w_9002 );
not (  , w_9003 );
and ( w_9002 , w_9003 , \3756_b0 );
or ( \3758_b1 , \3757_b1 , w_9004 );
xor ( \3758_b0 , \3757_b0 , w_9006 );
not ( w_9006 , w_9007 );
and ( w_9007 , w_9004 , w_9005 );
buf ( w_9004 , \1363_b1 );
not ( w_9004 , w_9008 );
not ( w_9005 , w_9009 );
and ( w_9008 , w_9009 , \1363_b0 );
or ( \3759_b1 , \1299_b1 , \1280_b1 );
not ( \1280_b1 , w_9010 );
and ( \3759_b0 , \1299_b0 , w_9011 );
and ( w_9010 , w_9011 , \1280_b0 );
or ( \3760_b1 , \1194_b1 , \1278_b1 );
not ( \1278_b1 , w_9012 );
and ( \3760_b0 , \1194_b0 , w_9013 );
and ( w_9012 , w_9013 , \1278_b0 );
or ( \3761_b1 , \3759_b1 , w_9015 );
not ( w_9015 , w_9016 );
and ( \3761_b0 , \3759_b0 , w_9017 );
and ( w_9016 ,  , w_9017 );
buf ( w_9015 , \3760_b1 );
not ( w_9015 , w_9018 );
not (  , w_9019 );
and ( w_9018 , w_9019 , \3760_b0 );
or ( \3762_b1 , \3761_b1 , w_9020 );
xor ( \3762_b0 , \3761_b0 , w_9022 );
not ( w_9022 , w_9023 );
and ( w_9023 , w_9020 , w_9021 );
buf ( w_9020 , \1177_b1 );
not ( w_9020 , w_9024 );
not ( w_9021 , w_9025 );
and ( w_9024 , w_9025 , \1177_b0 );
or ( \3763_b1 , \3758_b1 , \3762_b1 );
not ( \3762_b1 , w_9026 );
and ( \3763_b0 , \3758_b0 , w_9027 );
and ( w_9026 , w_9027 , \3762_b0 );
or ( \3764_b1 , \1422_b1 , \1062_b1 );
not ( \1062_b1 , w_9028 );
and ( \3764_b0 , \1422_b0 , w_9029 );
and ( w_9028 , w_9029 , \1062_b0 );
or ( \3765_b1 , \1304_b1 , \1060_b1 );
not ( \1060_b1 , w_9030 );
and ( \3765_b0 , \1304_b0 , w_9031 );
and ( w_9030 , w_9031 , \1060_b0 );
or ( \3766_b1 , \3764_b1 , w_9033 );
not ( w_9033 , w_9034 );
and ( \3766_b0 , \3764_b0 , w_9035 );
and ( w_9034 ,  , w_9035 );
buf ( w_9033 , \3765_b1 );
not ( w_9033 , w_9036 );
not (  , w_9037 );
and ( w_9036 , w_9037 , \3765_b0 );
or ( \3767_b1 , \3766_b1 , w_9038 );
xor ( \3767_b0 , \3766_b0 , w_9040 );
not ( w_9040 , w_9041 );
and ( w_9041 , w_9038 , w_9039 );
buf ( w_9038 , \984_b1 );
not ( w_9038 , w_9042 );
not ( w_9039 , w_9043 );
and ( w_9042 , w_9043 , \984_b0 );
or ( \3768_b1 , \3762_b1 , \3767_b1 );
not ( \3767_b1 , w_9044 );
and ( \3768_b0 , \3762_b0 , w_9045 );
and ( w_9044 , w_9045 , \3767_b0 );
or ( \3769_b1 , \3758_b1 , \3767_b1 );
not ( \3767_b1 , w_9046 );
and ( \3769_b0 , \3758_b0 , w_9047 );
and ( w_9046 , w_9047 , \3767_b0 );
or ( \3771_b1 , \343_b1 , \2913_b1 );
not ( \2913_b1 , w_9048 );
and ( \3771_b0 , \343_b0 , w_9049 );
and ( w_9048 , w_9049 , \2913_b0 );
or ( \3772_b1 , \353_b1 , \2910_b1 );
not ( \2910_b1 , w_9050 );
and ( \3772_b0 , \353_b0 , w_9051 );
and ( w_9050 , w_9051 , \2910_b0 );
or ( \3773_b1 , \3771_b1 , w_9053 );
not ( w_9053 , w_9054 );
and ( \3773_b0 , \3771_b0 , w_9055 );
and ( w_9054 ,  , w_9055 );
buf ( w_9053 , \3772_b1 );
not ( w_9053 , w_9056 );
not (  , w_9057 );
and ( w_9056 , w_9057 , \3772_b0 );
or ( \3774_b1 , \3773_b1 , w_9058 );
xor ( \3774_b0 , \3773_b0 , w_9060 );
not ( w_9060 , w_9061 );
and ( w_9061 , w_9058 , w_9059 );
buf ( w_9058 , \2371_b1 );
not ( w_9058 , w_9062 );
not ( w_9059 , w_9063 );
and ( w_9062 , w_9063 , \2371_b0 );
or ( \3775_b1 , \444_b1 , \2550_b1 );
not ( \2550_b1 , w_9064 );
and ( \3775_b0 , \444_b0 , w_9065 );
and ( w_9064 , w_9065 , \2550_b0 );
or ( \3776_b1 , \360_b1 , \2548_b1 );
not ( \2548_b1 , w_9066 );
and ( \3776_b0 , \360_b0 , w_9067 );
and ( w_9066 , w_9067 , \2548_b0 );
or ( \3777_b1 , \3775_b1 , w_9069 );
not ( w_9069 , w_9070 );
and ( \3777_b0 , \3775_b0 , w_9071 );
and ( w_9070 ,  , w_9071 );
buf ( w_9069 , \3776_b1 );
not ( w_9069 , w_9072 );
not (  , w_9073 );
and ( w_9072 , w_9073 , \3776_b0 );
or ( \3778_b1 , \3777_b1 , w_9074 );
xor ( \3778_b0 , \3777_b0 , w_9076 );
not ( w_9076 , w_9077 );
and ( w_9077 , w_9074 , w_9075 );
buf ( w_9074 , \2374_b1 );
not ( w_9074 , w_9078 );
not ( w_9075 , w_9079 );
and ( w_9078 , w_9079 , \2374_b0 );
or ( \3779_b1 , \3774_b1 , \3778_b1 );
not ( \3778_b1 , w_9080 );
and ( \3779_b0 , \3774_b0 , w_9081 );
and ( w_9080 , w_9081 , \3778_b0 );
or ( \3780_b1 , \3778_b1 , \320_b1 );
not ( \320_b1 , w_9082 );
and ( \3780_b0 , \3778_b0 , w_9083 );
and ( w_9082 , w_9083 , \320_b0 );
or ( \3781_b1 , \3774_b1 , \320_b1 );
not ( \320_b1 , w_9084 );
and ( \3781_b0 , \3774_b0 , w_9085 );
and ( w_9084 , w_9085 , \320_b0 );
or ( \3783_b1 , \3770_b1 , \3782_b1 );
not ( \3782_b1 , w_9086 );
and ( \3783_b0 , \3770_b0 , w_9087 );
and ( w_9086 , w_9087 , \3782_b0 );
or ( \3784_b1 , \593_b1 , \2261_b1 );
not ( \2261_b1 , w_9088 );
and ( \3784_b0 , \593_b0 , w_9089 );
and ( w_9088 , w_9089 , \2261_b0 );
or ( \3785_b1 , \495_b1 , \2259_b1 );
not ( \2259_b1 , w_9090 );
and ( \3785_b0 , \495_b0 , w_9091 );
and ( w_9090 , w_9091 , \2259_b0 );
or ( \3786_b1 , \3784_b1 , w_9093 );
not ( w_9093 , w_9094 );
and ( \3786_b0 , \3784_b0 , w_9095 );
and ( w_9094 ,  , w_9095 );
buf ( w_9093 , \3785_b1 );
not ( w_9093 , w_9096 );
not (  , w_9097 );
and ( w_9096 , w_9097 , \3785_b0 );
or ( \3787_b1 , \3786_b1 , w_9098 );
xor ( \3787_b0 , \3786_b0 , w_9100 );
not ( w_9100 , w_9101 );
and ( w_9101 , w_9098 , w_9099 );
buf ( w_9098 , \2124_b1 );
not ( w_9098 , w_9102 );
not ( w_9099 , w_9103 );
and ( w_9102 , w_9103 , \2124_b0 );
or ( \3788_b1 , \703_b1 , \1955_b1 );
not ( \1955_b1 , w_9104 );
and ( \3788_b0 , \703_b0 , w_9105 );
and ( w_9104 , w_9105 , \1955_b0 );
or ( \3789_b1 , \621_b1 , \1953_b1 );
not ( \1953_b1 , w_9106 );
and ( \3789_b0 , \621_b0 , w_9107 );
and ( w_9106 , w_9107 , \1953_b0 );
or ( \3790_b1 , \3788_b1 , w_9109 );
not ( w_9109 , w_9110 );
and ( \3790_b0 , \3788_b0 , w_9111 );
and ( w_9110 ,  , w_9111 );
buf ( w_9109 , \3789_b1 );
not ( w_9109 , w_9112 );
not (  , w_9113 );
and ( w_9112 , w_9113 , \3789_b0 );
or ( \3791_b1 , \3790_b1 , w_9114 );
xor ( \3791_b0 , \3790_b0 , w_9116 );
not ( w_9116 , w_9117 );
and ( w_9117 , w_9114 , w_9115 );
buf ( w_9114 , \1835_b1 );
not ( w_9114 , w_9118 );
not ( w_9115 , w_9119 );
and ( w_9118 , w_9119 , \1835_b0 );
or ( \3792_b1 , \3787_b1 , \3791_b1 );
not ( \3791_b1 , w_9120 );
and ( \3792_b0 , \3787_b0 , w_9121 );
and ( w_9120 , w_9121 , \3791_b0 );
or ( \3793_b1 , \841_b1 , \1742_b1 );
not ( \1742_b1 , w_9122 );
and ( \3793_b0 , \841_b0 , w_9123 );
and ( w_9122 , w_9123 , \1742_b0 );
or ( \3794_b1 , \777_b1 , \1740_b1 );
not ( \1740_b1 , w_9124 );
and ( \3794_b0 , \777_b0 , w_9125 );
and ( w_9124 , w_9125 , \1740_b0 );
or ( \3795_b1 , \3793_b1 , w_9127 );
not ( w_9127 , w_9128 );
and ( \3795_b0 , \3793_b0 , w_9129 );
and ( w_9128 ,  , w_9129 );
buf ( w_9127 , \3794_b1 );
not ( w_9127 , w_9130 );
not (  , w_9131 );
and ( w_9130 , w_9131 , \3794_b0 );
or ( \3796_b1 , \3795_b1 , w_9132 );
xor ( \3796_b0 , \3795_b0 , w_9134 );
not ( w_9134 , w_9135 );
and ( w_9135 , w_9132 , w_9133 );
buf ( w_9132 , \1610_b1 );
not ( w_9132 , w_9136 );
not ( w_9133 , w_9137 );
and ( w_9136 , w_9137 , \1610_b0 );
or ( \3797_b1 , \3791_b1 , \3796_b1 );
not ( \3796_b1 , w_9138 );
and ( \3797_b0 , \3791_b0 , w_9139 );
and ( w_9138 , w_9139 , \3796_b0 );
or ( \3798_b1 , \3787_b1 , \3796_b1 );
not ( \3796_b1 , w_9140 );
and ( \3798_b0 , \3787_b0 , w_9141 );
and ( w_9140 , w_9141 , \3796_b0 );
or ( \3800_b1 , \3782_b1 , \3799_b1 );
not ( \3799_b1 , w_9142 );
and ( \3800_b0 , \3782_b0 , w_9143 );
and ( w_9142 , w_9143 , \3799_b0 );
or ( \3801_b1 , \3770_b1 , \3799_b1 );
not ( \3799_b1 , w_9144 );
and ( \3801_b0 , \3770_b0 , w_9145 );
and ( w_9144 , w_9145 , \3799_b0 );
or ( \3803_b1 , \3754_b1 , \3802_b1 );
not ( \3802_b1 , w_9146 );
and ( \3803_b0 , \3754_b0 , w_9147 );
and ( w_9146 , w_9147 , \3802_b0 );
or ( \3804_b1 , \2850_b1 , \313_b1 );
not ( \313_b1 , w_9148 );
and ( \3804_b0 , \2850_b0 , w_9149 );
and ( w_9148 , w_9149 , \313_b0 );
or ( \3805_b1 , \2763_b1 , \311_b1 );
not ( \311_b1 , w_9150 );
and ( \3805_b0 , \2763_b0 , w_9151 );
and ( w_9150 , w_9151 , \311_b0 );
or ( \3806_b1 , \3804_b1 , w_9153 );
not ( w_9153 , w_9154 );
and ( \3806_b0 , \3804_b0 , w_9155 );
and ( w_9154 ,  , w_9155 );
buf ( w_9153 , \3805_b1 );
not ( w_9153 , w_9156 );
not (  , w_9157 );
and ( w_9156 , w_9157 , \3805_b0 );
or ( \3807_b1 , \3806_b1 , w_9158 );
xor ( \3807_b0 , \3806_b0 , w_9160 );
not ( w_9160 , w_9161 );
and ( w_9161 , w_9158 , w_9159 );
buf ( w_9158 , \320_b1 );
not ( w_9158 , w_9162 );
not ( w_9159 , w_9163 );
and ( w_9162 , w_9163 , \320_b0 );
or ( \3808_b1 , \3658_b1 , \3662_b1 );
xor ( \3808_b0 , \3658_b0 , w_9164 );
not ( w_9164 , w_9165 );
and ( w_9165 , \3662_b1 , \3662_b0 );
or ( \3809_b1 , \3808_b1 , \3667_b1 );
xor ( \3809_b0 , \3808_b0 , w_9166 );
not ( w_9166 , w_9167 );
and ( w_9167 , \3667_b1 , \3667_b0 );
or ( \3810_b1 , \3807_b1 , \3809_b1 );
not ( \3809_b1 , w_9168 );
and ( \3810_b0 , \3807_b0 , w_9169 );
and ( w_9168 , w_9169 , \3809_b0 );
or ( \3811_b1 , \3611_b1 , \3615_b1 );
xor ( \3811_b0 , \3611_b0 , w_9170 );
not ( w_9170 , w_9171 );
and ( w_9171 , \3615_b1 , \3615_b0 );
or ( \3812_b1 , \3811_b1 , \3620_b1 );
xor ( \3812_b0 , \3811_b0 , w_9172 );
not ( w_9172 , w_9173 );
and ( w_9173 , \3620_b1 , \3620_b0 );
or ( \3813_b1 , \3809_b1 , \3812_b1 );
not ( \3812_b1 , w_9174 );
and ( \3813_b0 , \3809_b0 , w_9175 );
and ( w_9174 , w_9175 , \3812_b0 );
or ( \3814_b1 , \3807_b1 , \3812_b1 );
not ( \3812_b1 , w_9176 );
and ( \3814_b0 , \3807_b0 , w_9177 );
and ( w_9176 , w_9177 , \3812_b0 );
or ( \3816_b1 , \3802_b1 , \3815_b1 );
not ( \3815_b1 , w_9178 );
and ( \3816_b0 , \3802_b0 , w_9179 );
and ( w_9178 , w_9179 , \3815_b0 );
or ( \3817_b1 , \3754_b1 , \3815_b1 );
not ( \3815_b1 , w_9180 );
and ( \3817_b0 , \3754_b0 , w_9181 );
and ( w_9180 , w_9181 , \3815_b0 );
or ( \3819_b1 , \3489_b1 , \3493_b1 );
xor ( \3819_b0 , \3489_b0 , w_9182 );
not ( w_9182 , w_9183 );
and ( w_9183 , \3493_b1 , \3493_b0 );
or ( \3820_b1 , \3819_b1 , \338_b1 );
xor ( \3820_b0 , \3819_b0 , w_9184 );
not ( w_9184 , w_9185 );
and ( w_9185 , \338_b1 , \338_b0 );
or ( \3821_b1 , \3645_b1 , \3647_b1 );
xor ( \3821_b0 , \3645_b0 , w_9186 );
not ( w_9186 , w_9187 );
and ( w_9187 , \3647_b1 , \3647_b0 );
or ( \3822_b1 , \3821_b1 , \3650_b1 );
xor ( \3822_b0 , \3821_b0 , w_9188 );
not ( w_9188 , w_9189 );
and ( w_9189 , \3650_b1 , \3650_b0 );
or ( \3823_b1 , \3820_b1 , \3822_b1 );
not ( \3822_b1 , w_9190 );
and ( \3823_b0 , \3820_b0 , w_9191 );
and ( w_9190 , w_9191 , \3822_b0 );
or ( \3824_b1 , \3670_b1 , \3672_b1 );
xor ( \3824_b0 , \3670_b0 , w_9192 );
not ( w_9192 , w_9193 );
and ( w_9193 , \3672_b1 , \3672_b0 );
or ( \3825_b1 , \3824_b1 , \3675_b1 );
xor ( \3825_b0 , \3824_b0 , w_9194 );
not ( w_9194 , w_9195 );
and ( w_9195 , \3675_b1 , \3675_b0 );
or ( \3826_b1 , \3822_b1 , \3825_b1 );
not ( \3825_b1 , w_9196 );
and ( \3826_b0 , \3822_b0 , w_9197 );
and ( w_9196 , w_9197 , \3825_b0 );
or ( \3827_b1 , \3820_b1 , \3825_b1 );
not ( \3825_b1 , w_9198 );
and ( \3827_b0 , \3820_b0 , w_9199 );
and ( w_9198 , w_9199 , \3825_b0 );
or ( \3829_b1 , \3818_b1 , \3828_b1 );
not ( \3828_b1 , w_9200 );
and ( \3829_b0 , \3818_b0 , w_9201 );
and ( w_9200 , w_9201 , \3828_b0 );
or ( \3830_b1 , \3468_b1 , \3484_b1 );
xor ( \3830_b0 , \3468_b0 , w_9202 );
not ( w_9202 , w_9203 );
and ( w_9203 , \3484_b1 , \3484_b0 );
or ( \3831_b1 , \3830_b1 , \3497_b1 );
xor ( \3831_b0 , \3830_b0 , w_9204 );
not ( w_9204 , w_9205 );
and ( w_9205 , \3497_b1 , \3497_b0 );
or ( \3832_b1 , \3828_b1 , \3831_b1 );
not ( \3831_b1 , w_9206 );
and ( \3832_b0 , \3828_b0 , w_9207 );
and ( w_9206 , w_9207 , \3831_b0 );
or ( \3833_b1 , \3818_b1 , \3831_b1 );
not ( \3831_b1 , w_9208 );
and ( \3833_b0 , \3818_b0 , w_9209 );
and ( w_9208 , w_9209 , \3831_b0 );
or ( \3835_b1 , \3643_b1 , \3653_b1 );
xor ( \3835_b0 , \3643_b0 , w_9210 );
not ( w_9210 , w_9211 );
and ( w_9211 , \3653_b1 , \3653_b0 );
or ( \3836_b1 , \3835_b1 , \3678_b1 );
xor ( \3836_b0 , \3835_b0 , w_9212 );
not ( w_9212 , w_9213 );
and ( w_9213 , \3678_b1 , \3678_b0 );
or ( \3837_b1 , \3683_b1 , \3685_b1 );
xor ( \3837_b0 , \3683_b0 , w_9214 );
not ( w_9214 , w_9215 );
and ( w_9215 , \3685_b1 , \3685_b0 );
or ( \3838_b1 , \3837_b1 , \3688_b1 );
xor ( \3838_b0 , \3837_b0 , w_9216 );
not ( w_9216 , w_9217 );
and ( w_9217 , \3688_b1 , \3688_b0 );
or ( \3839_b1 , \3836_b1 , \3838_b1 );
not ( \3838_b1 , w_9218 );
and ( \3839_b0 , \3836_b0 , w_9219 );
and ( w_9218 , w_9219 , \3838_b0 );
or ( \3840_b1 , \3834_b1 , \3839_b1 );
not ( \3839_b1 , w_9220 );
and ( \3840_b0 , \3834_b0 , w_9221 );
and ( w_9220 , w_9221 , \3839_b0 );
or ( \3841_b1 , \3554_b1 , \3556_b1 );
xor ( \3841_b0 , \3554_b0 , w_9222 );
not ( w_9222 , w_9223 );
and ( w_9223 , \3556_b1 , \3556_b0 );
or ( \3842_b1 , \3841_b1 , \3559_b1 );
xor ( \3842_b0 , \3841_b0 , w_9224 );
not ( w_9224 , w_9225 );
and ( w_9225 , \3559_b1 , \3559_b0 );
or ( \3843_b1 , \3839_b1 , \3842_b1 );
not ( \3842_b1 , w_9226 );
and ( \3843_b0 , \3839_b0 , w_9227 );
and ( w_9226 , w_9227 , \3842_b0 );
or ( \3844_b1 , \3834_b1 , \3842_b1 );
not ( \3842_b1 , w_9228 );
and ( \3844_b0 , \3834_b0 , w_9229 );
and ( w_9228 , w_9229 , \3842_b0 );
or ( \3846_b1 , \3500_b1 , \3538_b1 );
xor ( \3846_b0 , \3500_b0 , w_9230 );
not ( w_9230 , w_9231 );
and ( w_9231 , \3538_b1 , \3538_b0 );
or ( \3847_b1 , \3846_b1 , \3549_b1 );
xor ( \3847_b0 , \3846_b0 , w_9232 );
not ( w_9232 , w_9233 );
and ( w_9233 , \3549_b1 , \3549_b0 );
or ( \3848_b1 , \3681_b1 , \3691_b1 );
xor ( \3848_b0 , \3681_b0 , w_9234 );
not ( w_9234 , w_9235 );
and ( w_9235 , \3691_b1 , \3691_b0 );
or ( \3849_b1 , \3848_b1 , \3694_b1 );
xor ( \3849_b0 , \3848_b0 , w_9236 );
not ( w_9236 , w_9237 );
and ( w_9237 , \3694_b1 , \3694_b0 );
or ( \3850_b1 , \3847_b1 , \3849_b1 );
not ( \3849_b1 , w_9238 );
and ( \3850_b0 , \3847_b0 , w_9239 );
and ( w_9238 , w_9239 , \3849_b0 );
or ( \3851_b1 , \3845_b1 , \3850_b1 );
not ( \3850_b1 , w_9240 );
and ( \3851_b0 , \3845_b0 , w_9241 );
and ( w_9240 , w_9241 , \3850_b0 );
or ( \3852_b1 , \3697_b1 , \3699_b1 );
xor ( \3852_b0 , \3697_b0 , w_9242 );
not ( w_9242 , w_9243 );
and ( w_9243 , \3699_b1 , \3699_b0 );
or ( \3853_b1 , \3852_b1 , \3701_b1 );
xor ( \3853_b0 , \3852_b0 , w_9244 );
not ( w_9244 , w_9245 );
and ( w_9245 , \3701_b1 , \3701_b0 );
or ( \3854_b1 , \3850_b1 , \3853_b1 );
not ( \3853_b1 , w_9246 );
and ( \3854_b0 , \3850_b0 , w_9247 );
and ( w_9246 , w_9247 , \3853_b0 );
or ( \3855_b1 , \3845_b1 , \3853_b1 );
not ( \3853_b1 , w_9248 );
and ( \3855_b0 , \3845_b0 , w_9249 );
and ( w_9248 , w_9249 , \3853_b0 );
or ( \3857_b1 , \3716_b1 , \3856_b1 );
not ( \3856_b1 , w_9250 );
and ( \3857_b0 , \3716_b0 , w_9251 );
and ( w_9250 , w_9251 , \3856_b0 );
or ( \3858_b1 , \3716_b1 , \3856_b1 );
xor ( \3858_b0 , \3716_b0 , w_9252 );
not ( w_9252 , w_9253 );
and ( w_9253 , \3856_b1 , \3856_b0 );
or ( \3859_b1 , \3845_b1 , \3850_b1 );
xor ( \3859_b0 , \3845_b0 , w_9254 );
not ( w_9254 , w_9255 );
and ( w_9255 , \3850_b1 , \3850_b0 );
or ( \3860_b1 , \3859_b1 , \3853_b1 );
xor ( \3860_b0 , \3859_b0 , w_9256 );
not ( w_9256 , w_9257 );
and ( w_9257 , \3853_b1 , \3853_b0 );
or ( \3861_b1 , \777_b1 , \1955_b1 );
not ( \1955_b1 , w_9258 );
and ( \3861_b0 , \777_b0 , w_9259 );
and ( w_9258 , w_9259 , \1955_b0 );
or ( \3862_b1 , \703_b1 , \1953_b1 );
not ( \1953_b1 , w_9260 );
and ( \3862_b0 , \703_b0 , w_9261 );
and ( w_9260 , w_9261 , \1953_b0 );
or ( \3863_b1 , \3861_b1 , w_9263 );
not ( w_9263 , w_9264 );
and ( \3863_b0 , \3861_b0 , w_9265 );
and ( w_9264 ,  , w_9265 );
buf ( w_9263 , \3862_b1 );
not ( w_9263 , w_9266 );
not (  , w_9267 );
and ( w_9266 , w_9267 , \3862_b0 );
or ( \3864_b1 , \3863_b1 , w_9268 );
xor ( \3864_b0 , \3863_b0 , w_9270 );
not ( w_9270 , w_9271 );
and ( w_9271 , w_9268 , w_9269 );
buf ( w_9268 , \1835_b1 );
not ( w_9268 , w_9272 );
not ( w_9269 , w_9273 );
and ( w_9272 , w_9273 , \1835_b0 );
or ( \3865_b1 , \904_b1 , \1742_b1 );
not ( \1742_b1 , w_9274 );
and ( \3865_b0 , \904_b0 , w_9275 );
and ( w_9274 , w_9275 , \1742_b0 );
or ( \3866_b1 , \841_b1 , \1740_b1 );
not ( \1740_b1 , w_9276 );
and ( \3866_b0 , \841_b0 , w_9277 );
and ( w_9276 , w_9277 , \1740_b0 );
or ( \3867_b1 , \3865_b1 , w_9279 );
not ( w_9279 , w_9280 );
and ( \3867_b0 , \3865_b0 , w_9281 );
and ( w_9280 ,  , w_9281 );
buf ( w_9279 , \3866_b1 );
not ( w_9279 , w_9282 );
not (  , w_9283 );
and ( w_9282 , w_9283 , \3866_b0 );
or ( \3868_b1 , \3867_b1 , w_9284 );
xor ( \3868_b0 , \3867_b0 , w_9286 );
not ( w_9286 , w_9287 );
and ( w_9287 , w_9284 , w_9285 );
buf ( w_9284 , \1610_b1 );
not ( w_9284 , w_9288 );
not ( w_9285 , w_9289 );
and ( w_9288 , w_9289 , \1610_b0 );
or ( \3869_b1 , \3864_b1 , \3868_b1 );
not ( \3868_b1 , w_9290 );
and ( \3869_b0 , \3864_b0 , w_9291 );
and ( w_9290 , w_9291 , \3868_b0 );
or ( \3870_b1 , \1194_b1 , \1476_b1 );
not ( \1476_b1 , w_9292 );
and ( \3870_b0 , \1194_b0 , w_9293 );
and ( w_9292 , w_9293 , \1476_b0 );
or ( \3871_b1 , \1104_b1 , \1474_b1 );
not ( \1474_b1 , w_9294 );
and ( \3871_b0 , \1104_b0 , w_9295 );
and ( w_9294 , w_9295 , \1474_b0 );
or ( \3872_b1 , \3870_b1 , w_9297 );
not ( w_9297 , w_9298 );
and ( \3872_b0 , \3870_b0 , w_9299 );
and ( w_9298 ,  , w_9299 );
buf ( w_9297 , \3871_b1 );
not ( w_9297 , w_9300 );
not (  , w_9301 );
and ( w_9300 , w_9301 , \3871_b0 );
or ( \3873_b1 , \3872_b1 , w_9302 );
xor ( \3873_b0 , \3872_b0 , w_9304 );
not ( w_9304 , w_9305 );
and ( w_9305 , w_9302 , w_9303 );
buf ( w_9302 , \1363_b1 );
not ( w_9302 , w_9306 );
not ( w_9303 , w_9307 );
and ( w_9306 , w_9307 , \1363_b0 );
or ( \3874_b1 , \3868_b1 , \3873_b1 );
not ( \3873_b1 , w_9308 );
and ( \3874_b0 , \3868_b0 , w_9309 );
and ( w_9308 , w_9309 , \3873_b0 );
or ( \3875_b1 , \3864_b1 , \3873_b1 );
not ( \3873_b1 , w_9310 );
and ( \3875_b0 , \3864_b0 , w_9311 );
and ( w_9310 , w_9311 , \3873_b0 );
or ( \3877_b1 , \360_b1 , \2913_b1 );
not ( \2913_b1 , w_9312 );
and ( \3877_b0 , \360_b0 , w_9313 );
and ( w_9312 , w_9313 , \2913_b0 );
or ( \3878_b1 , \343_b1 , \2910_b1 );
not ( \2910_b1 , w_9314 );
and ( \3878_b0 , \343_b0 , w_9315 );
and ( w_9314 , w_9315 , \2910_b0 );
or ( \3879_b1 , \3877_b1 , w_9317 );
not ( w_9317 , w_9318 );
and ( \3879_b0 , \3877_b0 , w_9319 );
and ( w_9318 ,  , w_9319 );
buf ( w_9317 , \3878_b1 );
not ( w_9317 , w_9320 );
not (  , w_9321 );
and ( w_9320 , w_9321 , \3878_b0 );
or ( \3880_b1 , \3879_b1 , w_9322 );
xor ( \3880_b0 , \3879_b0 , w_9324 );
not ( w_9324 , w_9325 );
and ( w_9325 , w_9322 , w_9323 );
buf ( w_9322 , \2371_b1 );
not ( w_9322 , w_9326 );
not ( w_9323 , w_9327 );
and ( w_9326 , w_9327 , \2371_b0 );
or ( \3881_b1 , \495_b1 , \2550_b1 );
not ( \2550_b1 , w_9328 );
and ( \3881_b0 , \495_b0 , w_9329 );
and ( w_9328 , w_9329 , \2550_b0 );
or ( \3882_b1 , \444_b1 , \2548_b1 );
not ( \2548_b1 , w_9330 );
and ( \3882_b0 , \444_b0 , w_9331 );
and ( w_9330 , w_9331 , \2548_b0 );
or ( \3883_b1 , \3881_b1 , w_9333 );
not ( w_9333 , w_9334 );
and ( \3883_b0 , \3881_b0 , w_9335 );
and ( w_9334 ,  , w_9335 );
buf ( w_9333 , \3882_b1 );
not ( w_9333 , w_9336 );
not (  , w_9337 );
and ( w_9336 , w_9337 , \3882_b0 );
or ( \3884_b1 , \3883_b1 , w_9338 );
xor ( \3884_b0 , \3883_b0 , w_9340 );
not ( w_9340 , w_9341 );
and ( w_9341 , w_9338 , w_9339 );
buf ( w_9338 , \2374_b1 );
not ( w_9338 , w_9342 );
not ( w_9339 , w_9343 );
and ( w_9342 , w_9343 , \2374_b0 );
or ( \3885_b1 , \3880_b1 , \3884_b1 );
not ( \3884_b1 , w_9344 );
and ( \3885_b0 , \3880_b0 , w_9345 );
and ( w_9344 , w_9345 , \3884_b0 );
or ( \3886_b1 , \621_b1 , \2261_b1 );
not ( \2261_b1 , w_9346 );
and ( \3886_b0 , \621_b0 , w_9347 );
and ( w_9346 , w_9347 , \2261_b0 );
or ( \3887_b1 , \593_b1 , \2259_b1 );
not ( \2259_b1 , w_9348 );
and ( \3887_b0 , \593_b0 , w_9349 );
and ( w_9348 , w_9349 , \2259_b0 );
or ( \3888_b1 , \3886_b1 , w_9351 );
not ( w_9351 , w_9352 );
and ( \3888_b0 , \3886_b0 , w_9353 );
and ( w_9352 ,  , w_9353 );
buf ( w_9351 , \3887_b1 );
not ( w_9351 , w_9354 );
not (  , w_9355 );
and ( w_9354 , w_9355 , \3887_b0 );
or ( \3889_b1 , \3888_b1 , w_9356 );
xor ( \3889_b0 , \3888_b0 , w_9358 );
not ( w_9358 , w_9359 );
and ( w_9359 , w_9356 , w_9357 );
buf ( w_9356 , \2124_b1 );
not ( w_9356 , w_9360 );
not ( w_9357 , w_9361 );
and ( w_9360 , w_9361 , \2124_b0 );
or ( \3890_b1 , \3884_b1 , \3889_b1 );
not ( \3889_b1 , w_9362 );
and ( \3890_b0 , \3884_b0 , w_9363 );
and ( w_9362 , w_9363 , \3889_b0 );
or ( \3891_b1 , \3880_b1 , \3889_b1 );
not ( \3889_b1 , w_9364 );
and ( \3891_b0 , \3880_b0 , w_9365 );
and ( w_9364 , w_9365 , \3889_b0 );
or ( \3893_b1 , \3876_b1 , \3892_b1 );
not ( \3892_b1 , w_9366 );
and ( \3893_b0 , \3876_b0 , w_9367 );
and ( w_9366 , w_9367 , \3892_b0 );
or ( \3894_b1 , \1304_b1 , \1280_b1 );
not ( \1280_b1 , w_9368 );
and ( \3894_b0 , \1304_b0 , w_9369 );
and ( w_9368 , w_9369 , \1280_b0 );
or ( \3895_b1 , \1299_b1 , \1278_b1 );
not ( \1278_b1 , w_9370 );
and ( \3895_b0 , \1299_b0 , w_9371 );
and ( w_9370 , w_9371 , \1278_b0 );
or ( \3896_b1 , \3894_b1 , w_9373 );
not ( w_9373 , w_9374 );
and ( \3896_b0 , \3894_b0 , w_9375 );
and ( w_9374 ,  , w_9375 );
buf ( w_9373 , \3895_b1 );
not ( w_9373 , w_9376 );
not (  , w_9377 );
and ( w_9376 , w_9377 , \3895_b0 );
or ( \3897_b1 , \3896_b1 , w_9378 );
xor ( \3897_b0 , \3896_b0 , w_9380 );
not ( w_9380 , w_9381 );
and ( w_9381 , w_9378 , w_9379 );
buf ( w_9378 , \1177_b1 );
not ( w_9378 , w_9382 );
not ( w_9379 , w_9383 );
and ( w_9382 , w_9383 , \1177_b0 );
or ( \3898_b1 , \1537_b1 , \1062_b1 );
not ( \1062_b1 , w_9384 );
and ( \3898_b0 , \1537_b0 , w_9385 );
and ( w_9384 , w_9385 , \1062_b0 );
or ( \3899_b1 , \1422_b1 , \1060_b1 );
not ( \1060_b1 , w_9386 );
and ( \3899_b0 , \1422_b0 , w_9387 );
and ( w_9386 , w_9387 , \1060_b0 );
or ( \3900_b1 , \3898_b1 , w_9389 );
not ( w_9389 , w_9390 );
and ( \3900_b0 , \3898_b0 , w_9391 );
and ( w_9390 ,  , w_9391 );
buf ( w_9389 , \3899_b1 );
not ( w_9389 , w_9392 );
not (  , w_9393 );
and ( w_9392 , w_9393 , \3899_b0 );
or ( \3901_b1 , \3900_b1 , w_9394 );
xor ( \3901_b0 , \3900_b0 , w_9396 );
not ( w_9396 , w_9397 );
and ( w_9397 , w_9394 , w_9395 );
buf ( w_9394 , \984_b1 );
not ( w_9394 , w_9398 );
not ( w_9395 , w_9399 );
and ( w_9398 , w_9399 , \984_b0 );
or ( \3902_b1 , \3897_b1 , \3901_b1 );
not ( \3901_b1 , w_9400 );
and ( \3902_b0 , \3897_b0 , w_9401 );
and ( w_9400 , w_9401 , \3901_b0 );
or ( \3903_b1 , \1778_b1 , \912_b1 );
not ( \912_b1 , w_9402 );
and ( \3903_b0 , \1778_b0 , w_9403 );
and ( w_9402 , w_9403 , \912_b0 );
or ( \3904_b1 , \1770_b1 , \910_b1 );
not ( \910_b1 , w_9404 );
and ( \3904_b0 , \1770_b0 , w_9405 );
and ( w_9404 , w_9405 , \910_b0 );
or ( \3905_b1 , \3903_b1 , w_9407 );
not ( w_9407 , w_9408 );
and ( \3905_b0 , \3903_b0 , w_9409 );
and ( w_9408 ,  , w_9409 );
buf ( w_9407 , \3904_b1 );
not ( w_9407 , w_9410 );
not (  , w_9411 );
and ( w_9410 , w_9411 , \3904_b0 );
or ( \3906_b1 , \3905_b1 , w_9412 );
xor ( \3906_b0 , \3905_b0 , w_9414 );
not ( w_9414 , w_9415 );
and ( w_9415 , w_9412 , w_9413 );
buf ( w_9412 , \818_b1 );
not ( w_9412 , w_9416 );
not ( w_9413 , w_9417 );
and ( w_9416 , w_9417 , \818_b0 );
or ( \3907_b1 , \3901_b1 , \3906_b1 );
not ( \3906_b1 , w_9418 );
and ( \3907_b0 , \3901_b0 , w_9419 );
and ( w_9418 , w_9419 , \3906_b0 );
or ( \3908_b1 , \3897_b1 , \3906_b1 );
not ( \3906_b1 , w_9420 );
and ( \3908_b0 , \3897_b0 , w_9421 );
and ( w_9420 , w_9421 , \3906_b0 );
or ( \3910_b1 , \3892_b1 , \3909_b1 );
not ( \3909_b1 , w_9422 );
and ( \3910_b0 , \3892_b0 , w_9423 );
and ( w_9422 , w_9423 , \3909_b0 );
or ( \3911_b1 , \3876_b1 , \3909_b1 );
not ( \3909_b1 , w_9424 );
and ( \3911_b0 , \3876_b0 , w_9425 );
and ( w_9424 , w_9425 , \3909_b0 );
or ( \3913_b1 , \3758_b1 , \3762_b1 );
xor ( \3913_b0 , \3758_b0 , w_9426 );
not ( w_9426 , w_9427 );
and ( w_9427 , \3762_b1 , \3762_b0 );
or ( \3914_b1 , \3913_b1 , \3767_b1 );
xor ( \3914_b0 , \3913_b0 , w_9428 );
not ( w_9428 , w_9429 );
and ( w_9429 , \3767_b1 , \3767_b0 );
or ( \3915_b1 , \3774_b1 , \3778_b1 );
xor ( \3915_b0 , \3774_b0 , w_9430 );
not ( w_9430 , w_9431 );
and ( w_9431 , \3778_b1 , \3778_b0 );
or ( \3916_b1 , \3915_b1 , \320_b1 );
xor ( \3916_b0 , \3915_b0 , w_9432 );
not ( w_9432 , w_9433 );
and ( w_9433 , \320_b1 , \320_b0 );
or ( \3917_b1 , \3914_b1 , \3916_b1 );
not ( \3916_b1 , w_9434 );
and ( \3917_b0 , \3914_b0 , w_9435 );
and ( w_9434 , w_9435 , \3916_b0 );
or ( \3918_b1 , \3787_b1 , \3791_b1 );
xor ( \3918_b0 , \3787_b0 , w_9436 );
not ( w_9436 , w_9437 );
and ( w_9437 , \3791_b1 , \3791_b0 );
or ( \3919_b1 , \3918_b1 , \3796_b1 );
xor ( \3919_b0 , \3918_b0 , w_9438 );
not ( w_9438 , w_9439 );
and ( w_9439 , \3796_b1 , \3796_b0 );
or ( \3920_b1 , \3916_b1 , \3919_b1 );
not ( \3919_b1 , w_9440 );
and ( \3920_b0 , \3916_b0 , w_9441 );
and ( w_9440 , w_9441 , \3919_b0 );
or ( \3921_b1 , \3914_b1 , \3919_b1 );
not ( \3919_b1 , w_9442 );
and ( \3921_b0 , \3914_b0 , w_9443 );
and ( w_9442 , w_9443 , \3919_b0 );
or ( \3923_b1 , \3912_b1 , \3922_b1 );
not ( \3922_b1 , w_9444 );
and ( \3923_b0 , \3912_b0 , w_9445 );
and ( w_9444 , w_9445 , \3922_b0 );
or ( \3924_b1 , \2028_b1 , \740_b1 );
not ( \740_b1 , w_9446 );
and ( \3924_b0 , \2028_b0 , w_9447 );
and ( w_9446 , w_9447 , \740_b0 );
or ( \3925_b1 , \2023_b1 , \738_b1 );
not ( \738_b1 , w_9448 );
and ( \3925_b0 , \2023_b0 , w_9449 );
and ( w_9448 , w_9449 , \738_b0 );
or ( \3926_b1 , \3924_b1 , w_9451 );
not ( w_9451 , w_9452 );
and ( \3926_b0 , \3924_b0 , w_9453 );
and ( w_9452 ,  , w_9453 );
buf ( w_9451 , \3925_b1 );
not ( w_9451 , w_9454 );
not (  , w_9455 );
and ( w_9454 , w_9455 , \3925_b0 );
or ( \3927_b1 , \3926_b1 , w_9456 );
xor ( \3927_b0 , \3926_b0 , w_9458 );
not ( w_9458 , w_9459 );
and ( w_9459 , w_9456 , w_9457 );
buf ( w_9456 , \668_b1 );
not ( w_9456 , w_9460 );
not ( w_9457 , w_9461 );
and ( w_9460 , w_9461 , \668_b0 );
or ( \3928_b1 , \2305_b1 , \604_b1 );
not ( \604_b1 , w_9462 );
and ( \3928_b0 , \2305_b0 , w_9463 );
and ( w_9462 , w_9463 , \604_b0 );
or ( \3929_b1 , \2161_b1 , \602_b1 );
not ( \602_b1 , w_9464 );
and ( \3929_b0 , \2161_b0 , w_9465 );
and ( w_9464 , w_9465 , \602_b0 );
or ( \3930_b1 , \3928_b1 , w_9467 );
not ( w_9467 , w_9468 );
and ( \3930_b0 , \3928_b0 , w_9469 );
and ( w_9468 ,  , w_9469 );
buf ( w_9467 , \3929_b1 );
not ( w_9467 , w_9470 );
not (  , w_9471 );
and ( w_9470 , w_9471 , \3929_b0 );
or ( \3931_b1 , \3930_b1 , w_9472 );
xor ( \3931_b0 , \3930_b0 , w_9474 );
not ( w_9474 , w_9475 );
and ( w_9475 , w_9472 , w_9473 );
buf ( w_9472 , \561_b1 );
not ( w_9472 , w_9476 );
not ( w_9473 , w_9477 );
and ( w_9476 , w_9477 , \561_b0 );
or ( \3932_b1 , \3927_b1 , \3931_b1 );
not ( \3931_b1 , w_9478 );
and ( \3932_b0 , \3927_b0 , w_9479 );
and ( w_9478 , w_9479 , \3931_b0 );
or ( \3933_b1 , \2541_b1 , \503_b1 );
not ( \503_b1 , w_9480 );
and ( \3933_b0 , \2541_b0 , w_9481 );
and ( w_9480 , w_9481 , \503_b0 );
or ( \3934_b1 , \2532_b1 , \501_b1 );
not ( \501_b1 , w_9482 );
and ( \3934_b0 , \2532_b0 , w_9483 );
and ( w_9482 , w_9483 , \501_b0 );
or ( \3935_b1 , \3933_b1 , w_9485 );
not ( w_9485 , w_9486 );
and ( \3935_b0 , \3933_b0 , w_9487 );
and ( w_9486 ,  , w_9487 );
buf ( w_9485 , \3934_b1 );
not ( w_9485 , w_9488 );
not (  , w_9489 );
and ( w_9488 , w_9489 , \3934_b0 );
or ( \3936_b1 , \3935_b1 , w_9490 );
xor ( \3936_b0 , \3935_b0 , w_9492 );
not ( w_9492 , w_9493 );
and ( w_9493 , w_9490 , w_9491 );
buf ( w_9490 , \455_b1 );
not ( w_9490 , w_9494 );
not ( w_9491 , w_9495 );
and ( w_9494 , w_9495 , \455_b0 );
or ( \3937_b1 , \3931_b1 , \3936_b1 );
not ( \3936_b1 , w_9496 );
and ( \3937_b0 , \3931_b0 , w_9497 );
and ( w_9496 , w_9497 , \3936_b0 );
or ( \3938_b1 , \3927_b1 , \3936_b1 );
not ( \3936_b1 , w_9498 );
and ( \3938_b0 , \3927_b0 , w_9499 );
and ( w_9498 , w_9499 , \3936_b0 );
or ( \3940_b1 , \3720_b1 , \3724_b1 );
xor ( \3940_b0 , \3720_b0 , w_9500 );
not ( w_9500 , w_9501 );
and ( w_9501 , \3724_b1 , \3724_b0 );
or ( \3941_b1 , \3940_b1 , \3729_b1 );
xor ( \3941_b0 , \3940_b0 , w_9502 );
not ( w_9502 , w_9503 );
and ( w_9503 , \3729_b1 , \3729_b0 );
or ( \3942_b1 , \3939_b1 , \3941_b1 );
not ( \3941_b1 , w_9504 );
and ( \3942_b0 , \3939_b0 , w_9505 );
and ( w_9504 , w_9505 , \3941_b0 );
or ( \3943_b1 , \3736_b1 , \3740_b1 );
xor ( \3943_b0 , \3736_b0 , w_9506 );
not ( w_9506 , w_9507 );
and ( w_9507 , \3740_b1 , \3740_b0 );
or ( \3944_b1 , \3943_b1 , \3743_b1 );
xor ( \3944_b0 , \3943_b0 , w_9508 );
not ( w_9508 , w_9509 );
and ( w_9509 , \3743_b1 , \3743_b0 );
or ( \3945_b1 , \3941_b1 , \3944_b1 );
not ( \3944_b1 , w_9510 );
and ( \3945_b0 , \3941_b0 , w_9511 );
and ( w_9510 , w_9511 , \3944_b0 );
or ( \3946_b1 , \3939_b1 , \3944_b1 );
not ( \3944_b1 , w_9512 );
and ( \3946_b0 , \3939_b0 , w_9513 );
and ( w_9512 , w_9513 , \3944_b0 );
or ( \3948_b1 , \3922_b1 , \3947_b1 );
not ( \3947_b1 , w_9514 );
and ( \3948_b0 , \3922_b0 , w_9515 );
and ( w_9514 , w_9515 , \3947_b0 );
or ( \3949_b1 , \3912_b1 , \3947_b1 );
not ( \3947_b1 , w_9516 );
and ( \3949_b0 , \3912_b0 , w_9517 );
and ( w_9516 , w_9517 , \3947_b0 );
or ( \3951_b1 , \3595_b1 , \3599_b1 );
xor ( \3951_b0 , \3595_b0 , w_9518 );
not ( w_9518 , w_9519 );
and ( w_9519 , \3599_b1 , \3599_b0 );
or ( \3952_b1 , \3951_b1 , \3604_b1 );
xor ( \3952_b0 , \3951_b0 , w_9520 );
not ( w_9520 , w_9521 );
and ( w_9521 , \3604_b1 , \3604_b0 );
or ( \3953_b1 , \3628_b1 , \3632_b1 );
xor ( \3953_b0 , \3628_b0 , w_9522 );
not ( w_9522 , w_9523 );
and ( w_9523 , \3632_b1 , \3632_b0 );
or ( \3954_b1 , \3953_b1 , \3637_b1 );
xor ( \3954_b0 , \3953_b0 , w_9524 );
not ( w_9524 , w_9525 );
and ( w_9525 , \3637_b1 , \3637_b0 );
or ( \3955_b1 , \3952_b1 , \3954_b1 );
not ( \3954_b1 , w_9526 );
and ( \3955_b0 , \3952_b0 , w_9527 );
and ( w_9526 , w_9527 , \3954_b0 );
or ( \3956_b1 , \3807_b1 , \3809_b1 );
xor ( \3956_b0 , \3807_b0 , w_9528 );
not ( w_9528 , w_9529 );
and ( w_9529 , \3809_b1 , \3809_b0 );
or ( \3957_b1 , \3956_b1 , \3812_b1 );
xor ( \3957_b0 , \3956_b0 , w_9530 );
not ( w_9530 , w_9531 );
and ( w_9531 , \3812_b1 , \3812_b0 );
or ( \3958_b1 , \3954_b1 , \3957_b1 );
not ( \3957_b1 , w_9532 );
and ( \3958_b0 , \3954_b0 , w_9533 );
and ( w_9532 , w_9533 , \3957_b0 );
or ( \3959_b1 , \3952_b1 , \3957_b1 );
not ( \3957_b1 , w_9534 );
and ( \3959_b0 , \3952_b0 , w_9535 );
and ( w_9534 , w_9535 , \3957_b0 );
or ( \3961_b1 , \3950_b1 , \3960_b1 );
not ( \3960_b1 , w_9536 );
and ( \3961_b0 , \3950_b0 , w_9537 );
and ( w_9536 , w_9537 , \3960_b0 );
or ( \3962_b1 , \3607_b1 , \3623_b1 );
xor ( \3962_b0 , \3607_b0 , w_9538 );
not ( w_9538 , w_9539 );
and ( w_9539 , \3623_b1 , \3623_b0 );
or ( \3963_b1 , \3962_b1 , \3640_b1 );
xor ( \3963_b0 , \3962_b0 , w_9540 );
not ( w_9540 , w_9541 );
and ( w_9541 , \3640_b1 , \3640_b0 );
or ( \3964_b1 , \3960_b1 , \3963_b1 );
not ( \3963_b1 , w_9542 );
and ( \3964_b0 , \3960_b0 , w_9543 );
and ( w_9542 , w_9543 , \3963_b0 );
or ( \3965_b1 , \3950_b1 , \3963_b1 );
not ( \3963_b1 , w_9544 );
and ( \3965_b0 , \3950_b0 , w_9545 );
and ( w_9544 , w_9545 , \3963_b0 );
or ( \3967_b1 , \3818_b1 , \3828_b1 );
xor ( \3967_b0 , \3818_b0 , w_9546 );
not ( w_9546 , w_9547 );
and ( w_9547 , \3828_b1 , \3828_b0 );
or ( \3968_b1 , \3967_b1 , \3831_b1 );
xor ( \3968_b0 , \3967_b0 , w_9548 );
not ( w_9548 , w_9549 );
and ( w_9549 , \3831_b1 , \3831_b0 );
or ( \3969_b1 , \3966_b1 , \3968_b1 );
not ( \3968_b1 , w_9550 );
and ( \3969_b0 , \3966_b0 , w_9551 );
and ( w_9550 , w_9551 , \3968_b0 );
or ( \3970_b1 , \3836_b1 , \3838_b1 );
xor ( \3970_b0 , \3836_b0 , w_9552 );
not ( w_9552 , w_9553 );
and ( w_9553 , \3838_b1 , \3838_b0 );
or ( \3971_b1 , \3968_b1 , \3970_b1 );
not ( \3970_b1 , w_9554 );
and ( \3971_b0 , \3968_b0 , w_9555 );
and ( w_9554 , w_9555 , \3970_b0 );
or ( \3972_b1 , \3966_b1 , \3970_b1 );
not ( \3970_b1 , w_9556 );
and ( \3972_b0 , \3966_b0 , w_9557 );
and ( w_9556 , w_9557 , \3970_b0 );
or ( \3974_b1 , \3834_b1 , \3839_b1 );
xor ( \3974_b0 , \3834_b0 , w_9558 );
not ( w_9558 , w_9559 );
and ( w_9559 , \3839_b1 , \3839_b0 );
or ( \3975_b1 , \3974_b1 , \3842_b1 );
xor ( \3975_b0 , \3974_b0 , w_9560 );
not ( w_9560 , w_9561 );
and ( w_9561 , \3842_b1 , \3842_b0 );
or ( \3976_b1 , \3973_b1 , \3975_b1 );
not ( \3975_b1 , w_9562 );
and ( \3976_b0 , \3973_b0 , w_9563 );
and ( w_9562 , w_9563 , \3975_b0 );
or ( \3977_b1 , \3847_b1 , \3849_b1 );
xor ( \3977_b0 , \3847_b0 , w_9564 );
not ( w_9564 , w_9565 );
and ( w_9565 , \3849_b1 , \3849_b0 );
or ( \3978_b1 , \3975_b1 , \3977_b1 );
not ( \3977_b1 , w_9566 );
and ( \3978_b0 , \3975_b0 , w_9567 );
and ( w_9566 , w_9567 , \3977_b0 );
or ( \3979_b1 , \3973_b1 , \3977_b1 );
not ( \3977_b1 , w_9568 );
and ( \3979_b0 , \3973_b0 , w_9569 );
and ( w_9568 , w_9569 , \3977_b0 );
or ( \3981_b1 , \3860_b1 , \3980_b1 );
not ( \3980_b1 , w_9570 );
and ( \3981_b0 , \3860_b0 , w_9571 );
and ( w_9570 , w_9571 , \3980_b0 );
or ( \3982_b1 , \3860_b1 , \3980_b1 );
xor ( \3982_b0 , \3860_b0 , w_9572 );
not ( w_9572 , w_9573 );
and ( w_9573 , \3980_b1 , \3980_b0 );
or ( \3983_b1 , \3973_b1 , \3975_b1 );
xor ( \3983_b0 , \3973_b0 , w_9574 );
not ( w_9574 , w_9575 );
and ( w_9575 , \3975_b1 , \3975_b0 );
or ( \3984_b1 , \3983_b1 , \3977_b1 );
xor ( \3984_b0 , \3983_b0 , w_9576 );
not ( w_9576 , w_9577 );
and ( w_9577 , \3977_b1 , \3977_b0 );
or ( \3985_b1 , \703_b1 , \2261_b1 );
not ( \2261_b1 , w_9578 );
and ( \3985_b0 , \703_b0 , w_9579 );
and ( w_9578 , w_9579 , \2261_b0 );
or ( \3986_b1 , \621_b1 , \2259_b1 );
not ( \2259_b1 , w_9580 );
and ( \3986_b0 , \621_b0 , w_9581 );
and ( w_9580 , w_9581 , \2259_b0 );
or ( \3987_b1 , \3985_b1 , w_9583 );
not ( w_9583 , w_9584 );
and ( \3987_b0 , \3985_b0 , w_9585 );
and ( w_9584 ,  , w_9585 );
buf ( w_9583 , \3986_b1 );
not ( w_9583 , w_9586 );
not (  , w_9587 );
and ( w_9586 , w_9587 , \3986_b0 );
or ( \3988_b1 , \3987_b1 , w_9588 );
xor ( \3988_b0 , \3987_b0 , w_9590 );
not ( w_9590 , w_9591 );
and ( w_9591 , w_9588 , w_9589 );
buf ( w_9588 , \2124_b1 );
not ( w_9588 , w_9592 );
not ( w_9589 , w_9593 );
and ( w_9592 , w_9593 , \2124_b0 );
or ( \3989_b1 , \841_b1 , \1955_b1 );
not ( \1955_b1 , w_9594 );
and ( \3989_b0 , \841_b0 , w_9595 );
and ( w_9594 , w_9595 , \1955_b0 );
or ( \3990_b1 , \777_b1 , \1953_b1 );
not ( \1953_b1 , w_9596 );
and ( \3990_b0 , \777_b0 , w_9597 );
and ( w_9596 , w_9597 , \1953_b0 );
or ( \3991_b1 , \3989_b1 , w_9599 );
not ( w_9599 , w_9600 );
and ( \3991_b0 , \3989_b0 , w_9601 );
and ( w_9600 ,  , w_9601 );
buf ( w_9599 , \3990_b1 );
not ( w_9599 , w_9602 );
not (  , w_9603 );
and ( w_9602 , w_9603 , \3990_b0 );
or ( \3992_b1 , \3991_b1 , w_9604 );
xor ( \3992_b0 , \3991_b0 , w_9606 );
not ( w_9606 , w_9607 );
and ( w_9607 , w_9604 , w_9605 );
buf ( w_9604 , \1835_b1 );
not ( w_9604 , w_9608 );
not ( w_9605 , w_9609 );
and ( w_9608 , w_9609 , \1835_b0 );
or ( \3993_b1 , \3988_b1 , \3992_b1 );
not ( \3992_b1 , w_9610 );
and ( \3993_b0 , \3988_b0 , w_9611 );
and ( w_9610 , w_9611 , \3992_b0 );
or ( \3994_b1 , \1104_b1 , \1742_b1 );
not ( \1742_b1 , w_9612 );
and ( \3994_b0 , \1104_b0 , w_9613 );
and ( w_9612 , w_9613 , \1742_b0 );
or ( \3995_b1 , \904_b1 , \1740_b1 );
not ( \1740_b1 , w_9614 );
and ( \3995_b0 , \904_b0 , w_9615 );
and ( w_9614 , w_9615 , \1740_b0 );
or ( \3996_b1 , \3994_b1 , w_9617 );
not ( w_9617 , w_9618 );
and ( \3996_b0 , \3994_b0 , w_9619 );
and ( w_9618 ,  , w_9619 );
buf ( w_9617 , \3995_b1 );
not ( w_9617 , w_9620 );
not (  , w_9621 );
and ( w_9620 , w_9621 , \3995_b0 );
or ( \3997_b1 , \3996_b1 , w_9622 );
xor ( \3997_b0 , \3996_b0 , w_9624 );
not ( w_9624 , w_9625 );
and ( w_9625 , w_9622 , w_9623 );
buf ( w_9622 , \1610_b1 );
not ( w_9622 , w_9626 );
not ( w_9623 , w_9627 );
and ( w_9626 , w_9627 , \1610_b0 );
or ( \3998_b1 , \3992_b1 , \3997_b1 );
not ( \3997_b1 , w_9628 );
and ( \3998_b0 , \3992_b0 , w_9629 );
and ( w_9628 , w_9629 , \3997_b0 );
or ( \3999_b1 , \3988_b1 , \3997_b1 );
not ( \3997_b1 , w_9630 );
and ( \3999_b0 , \3988_b0 , w_9631 );
and ( w_9630 , w_9631 , \3997_b0 );
or ( \4001_b1 , \444_b1 , \2913_b1 );
not ( \2913_b1 , w_9632 );
and ( \4001_b0 , \444_b0 , w_9633 );
and ( w_9632 , w_9633 , \2913_b0 );
or ( \4002_b1 , \360_b1 , \2910_b1 );
not ( \2910_b1 , w_9634 );
and ( \4002_b0 , \360_b0 , w_9635 );
and ( w_9634 , w_9635 , \2910_b0 );
or ( \4003_b1 , \4001_b1 , w_9637 );
not ( w_9637 , w_9638 );
and ( \4003_b0 , \4001_b0 , w_9639 );
and ( w_9638 ,  , w_9639 );
buf ( w_9637 , \4002_b1 );
not ( w_9637 , w_9640 );
not (  , w_9641 );
and ( w_9640 , w_9641 , \4002_b0 );
or ( \4004_b1 , \4003_b1 , w_9642 );
xor ( \4004_b0 , \4003_b0 , w_9644 );
not ( w_9644 , w_9645 );
and ( w_9645 , w_9642 , w_9643 );
buf ( w_9642 , \2371_b1 );
not ( w_9642 , w_9646 );
not ( w_9643 , w_9647 );
and ( w_9646 , w_9647 , \2371_b0 );
or ( \4005_b1 , \593_b1 , \2550_b1 );
not ( \2550_b1 , w_9648 );
and ( \4005_b0 , \593_b0 , w_9649 );
and ( w_9648 , w_9649 , \2550_b0 );
or ( \4006_b1 , \495_b1 , \2548_b1 );
not ( \2548_b1 , w_9650 );
and ( \4006_b0 , \495_b0 , w_9651 );
and ( w_9650 , w_9651 , \2548_b0 );
or ( \4007_b1 , \4005_b1 , w_9653 );
not ( w_9653 , w_9654 );
and ( \4007_b0 , \4005_b0 , w_9655 );
and ( w_9654 ,  , w_9655 );
buf ( w_9653 , \4006_b1 );
not ( w_9653 , w_9656 );
not (  , w_9657 );
and ( w_9656 , w_9657 , \4006_b0 );
or ( \4008_b1 , \4007_b1 , w_9658 );
xor ( \4008_b0 , \4007_b0 , w_9660 );
not ( w_9660 , w_9661 );
and ( w_9661 , w_9658 , w_9659 );
buf ( w_9658 , \2374_b1 );
not ( w_9658 , w_9662 );
not ( w_9659 , w_9663 );
and ( w_9662 , w_9663 , \2374_b0 );
or ( \4009_b1 , \4004_b1 , \4008_b1 );
not ( \4008_b1 , w_9664 );
and ( \4009_b0 , \4004_b0 , w_9665 );
and ( w_9664 , w_9665 , \4008_b0 );
or ( \4010_b1 , \4008_b1 , \303_b1 );
not ( \303_b1 , w_9666 );
and ( \4010_b0 , \4008_b0 , w_9667 );
and ( w_9666 , w_9667 , \303_b0 );
or ( \4011_b1 , \4004_b1 , \303_b1 );
not ( \303_b1 , w_9668 );
and ( \4011_b0 , \4004_b0 , w_9669 );
and ( w_9668 , w_9669 , \303_b0 );
or ( \4013_b1 , \4000_b1 , \4012_b1 );
not ( \4012_b1 , w_9670 );
and ( \4013_b0 , \4000_b0 , w_9671 );
and ( w_9670 , w_9671 , \4012_b0 );
or ( \4014_b1 , \1299_b1 , \1476_b1 );
not ( \1476_b1 , w_9672 );
and ( \4014_b0 , \1299_b0 , w_9673 );
and ( w_9672 , w_9673 , \1476_b0 );
or ( \4015_b1 , \1194_b1 , \1474_b1 );
not ( \1474_b1 , w_9674 );
and ( \4015_b0 , \1194_b0 , w_9675 );
and ( w_9674 , w_9675 , \1474_b0 );
or ( \4016_b1 , \4014_b1 , w_9677 );
not ( w_9677 , w_9678 );
and ( \4016_b0 , \4014_b0 , w_9679 );
and ( w_9678 ,  , w_9679 );
buf ( w_9677 , \4015_b1 );
not ( w_9677 , w_9680 );
not (  , w_9681 );
and ( w_9680 , w_9681 , \4015_b0 );
or ( \4017_b1 , \4016_b1 , w_9682 );
xor ( \4017_b0 , \4016_b0 , w_9684 );
not ( w_9684 , w_9685 );
and ( w_9685 , w_9682 , w_9683 );
buf ( w_9682 , \1363_b1 );
not ( w_9682 , w_9686 );
not ( w_9683 , w_9687 );
and ( w_9686 , w_9687 , \1363_b0 );
or ( \4018_b1 , \1422_b1 , \1280_b1 );
not ( \1280_b1 , w_9688 );
and ( \4018_b0 , \1422_b0 , w_9689 );
and ( w_9688 , w_9689 , \1280_b0 );
or ( \4019_b1 , \1304_b1 , \1278_b1 );
not ( \1278_b1 , w_9690 );
and ( \4019_b0 , \1304_b0 , w_9691 );
and ( w_9690 , w_9691 , \1278_b0 );
or ( \4020_b1 , \4018_b1 , w_9693 );
not ( w_9693 , w_9694 );
and ( \4020_b0 , \4018_b0 , w_9695 );
and ( w_9694 ,  , w_9695 );
buf ( w_9693 , \4019_b1 );
not ( w_9693 , w_9696 );
not (  , w_9697 );
and ( w_9696 , w_9697 , \4019_b0 );
or ( \4021_b1 , \4020_b1 , w_9698 );
xor ( \4021_b0 , \4020_b0 , w_9700 );
not ( w_9700 , w_9701 );
and ( w_9701 , w_9698 , w_9699 );
buf ( w_9698 , \1177_b1 );
not ( w_9698 , w_9702 );
not ( w_9699 , w_9703 );
and ( w_9702 , w_9703 , \1177_b0 );
or ( \4022_b1 , \4017_b1 , \4021_b1 );
not ( \4021_b1 , w_9704 );
and ( \4022_b0 , \4017_b0 , w_9705 );
and ( w_9704 , w_9705 , \4021_b0 );
or ( \4023_b1 , \1770_b1 , \1062_b1 );
not ( \1062_b1 , w_9706 );
and ( \4023_b0 , \1770_b0 , w_9707 );
and ( w_9706 , w_9707 , \1062_b0 );
or ( \4024_b1 , \1537_b1 , \1060_b1 );
not ( \1060_b1 , w_9708 );
and ( \4024_b0 , \1537_b0 , w_9709 );
and ( w_9708 , w_9709 , \1060_b0 );
or ( \4025_b1 , \4023_b1 , w_9711 );
not ( w_9711 , w_9712 );
and ( \4025_b0 , \4023_b0 , w_9713 );
and ( w_9712 ,  , w_9713 );
buf ( w_9711 , \4024_b1 );
not ( w_9711 , w_9714 );
not (  , w_9715 );
and ( w_9714 , w_9715 , \4024_b0 );
or ( \4026_b1 , \4025_b1 , w_9716 );
xor ( \4026_b0 , \4025_b0 , w_9718 );
not ( w_9718 , w_9719 );
and ( w_9719 , w_9716 , w_9717 );
buf ( w_9716 , \984_b1 );
not ( w_9716 , w_9720 );
not ( w_9717 , w_9721 );
and ( w_9720 , w_9721 , \984_b0 );
or ( \4027_b1 , \4021_b1 , \4026_b1 );
not ( \4026_b1 , w_9722 );
and ( \4027_b0 , \4021_b0 , w_9723 );
and ( w_9722 , w_9723 , \4026_b0 );
or ( \4028_b1 , \4017_b1 , \4026_b1 );
not ( \4026_b1 , w_9724 );
and ( \4028_b0 , \4017_b0 , w_9725 );
and ( w_9724 , w_9725 , \4026_b0 );
or ( \4030_b1 , \4012_b1 , \4029_b1 );
not ( \4029_b1 , w_9726 );
and ( \4030_b0 , \4012_b0 , w_9727 );
and ( w_9726 , w_9727 , \4029_b0 );
or ( \4031_b1 , \4000_b1 , \4029_b1 );
not ( \4029_b1 , w_9728 );
and ( \4031_b0 , \4000_b0 , w_9729 );
and ( w_9728 , w_9729 , \4029_b0 );
or ( \4033_b1 , \2023_b1 , \912_b1 );
not ( \912_b1 , w_9730 );
and ( \4033_b0 , \2023_b0 , w_9731 );
and ( w_9730 , w_9731 , \912_b0 );
or ( \4034_b1 , \1778_b1 , \910_b1 );
not ( \910_b1 , w_9732 );
and ( \4034_b0 , \1778_b0 , w_9733 );
and ( w_9732 , w_9733 , \910_b0 );
or ( \4035_b1 , \4033_b1 , w_9735 );
not ( w_9735 , w_9736 );
and ( \4035_b0 , \4033_b0 , w_9737 );
and ( w_9736 ,  , w_9737 );
buf ( w_9735 , \4034_b1 );
not ( w_9735 , w_9738 );
not (  , w_9739 );
and ( w_9738 , w_9739 , \4034_b0 );
or ( \4036_b1 , \4035_b1 , w_9740 );
xor ( \4036_b0 , \4035_b0 , w_9742 );
not ( w_9742 , w_9743 );
and ( w_9743 , w_9740 , w_9741 );
buf ( w_9740 , \818_b1 );
not ( w_9740 , w_9744 );
not ( w_9741 , w_9745 );
and ( w_9744 , w_9745 , \818_b0 );
or ( \4037_b1 , \2161_b1 , \740_b1 );
not ( \740_b1 , w_9746 );
and ( \4037_b0 , \2161_b0 , w_9747 );
and ( w_9746 , w_9747 , \740_b0 );
or ( \4038_b1 , \2028_b1 , \738_b1 );
not ( \738_b1 , w_9748 );
and ( \4038_b0 , \2028_b0 , w_9749 );
and ( w_9748 , w_9749 , \738_b0 );
or ( \4039_b1 , \4037_b1 , w_9751 );
not ( w_9751 , w_9752 );
and ( \4039_b0 , \4037_b0 , w_9753 );
and ( w_9752 ,  , w_9753 );
buf ( w_9751 , \4038_b1 );
not ( w_9751 , w_9754 );
not (  , w_9755 );
and ( w_9754 , w_9755 , \4038_b0 );
or ( \4040_b1 , \4039_b1 , w_9756 );
xor ( \4040_b0 , \4039_b0 , w_9758 );
not ( w_9758 , w_9759 );
and ( w_9759 , w_9756 , w_9757 );
buf ( w_9756 , \668_b1 );
not ( w_9756 , w_9760 );
not ( w_9757 , w_9761 );
and ( w_9760 , w_9761 , \668_b0 );
or ( \4041_b1 , \4036_b1 , \4040_b1 );
not ( \4040_b1 , w_9762 );
and ( \4041_b0 , \4036_b0 , w_9763 );
and ( w_9762 , w_9763 , \4040_b0 );
or ( \4042_b1 , \2532_b1 , \604_b1 );
not ( \604_b1 , w_9764 );
and ( \4042_b0 , \2532_b0 , w_9765 );
and ( w_9764 , w_9765 , \604_b0 );
or ( \4043_b1 , \2305_b1 , \602_b1 );
not ( \602_b1 , w_9766 );
and ( \4043_b0 , \2305_b0 , w_9767 );
and ( w_9766 , w_9767 , \602_b0 );
or ( \4044_b1 , \4042_b1 , w_9769 );
not ( w_9769 , w_9770 );
and ( \4044_b0 , \4042_b0 , w_9771 );
and ( w_9770 ,  , w_9771 );
buf ( w_9769 , \4043_b1 );
not ( w_9769 , w_9772 );
not (  , w_9773 );
and ( w_9772 , w_9773 , \4043_b0 );
or ( \4045_b1 , \4044_b1 , w_9774 );
xor ( \4045_b0 , \4044_b0 , w_9776 );
not ( w_9776 , w_9777 );
and ( w_9777 , w_9774 , w_9775 );
buf ( w_9774 , \561_b1 );
not ( w_9774 , w_9778 );
not ( w_9775 , w_9779 );
and ( w_9778 , w_9779 , \561_b0 );
or ( \4046_b1 , \4040_b1 , \4045_b1 );
not ( \4045_b1 , w_9780 );
and ( \4046_b0 , \4040_b0 , w_9781 );
and ( w_9780 , w_9781 , \4045_b0 );
or ( \4047_b1 , \4036_b1 , \4045_b1 );
not ( \4045_b1 , w_9782 );
and ( \4047_b0 , \4036_b0 , w_9783 );
and ( w_9782 , w_9783 , \4045_b0 );
or ( \4049_b1 , \2763_b1 , \503_b1 );
not ( \503_b1 , w_9784 );
and ( \4049_b0 , \2763_b0 , w_9785 );
and ( w_9784 , w_9785 , \503_b0 );
or ( \4050_b1 , \2541_b1 , \501_b1 );
not ( \501_b1 , w_9786 );
and ( \4050_b0 , \2541_b0 , w_9787 );
and ( w_9786 , w_9787 , \501_b0 );
or ( \4051_b1 , \4049_b1 , w_9789 );
not ( w_9789 , w_9790 );
and ( \4051_b0 , \4049_b0 , w_9791 );
and ( w_9790 ,  , w_9791 );
buf ( w_9789 , \4050_b1 );
not ( w_9789 , w_9792 );
not (  , w_9793 );
and ( w_9792 , w_9793 , \4050_b0 );
or ( \4052_b1 , \4051_b1 , w_9794 );
xor ( \4052_b0 , \4051_b0 , w_9796 );
not ( w_9796 , w_9797 );
and ( w_9797 , w_9794 , w_9795 );
buf ( w_9794 , \455_b1 );
not ( w_9794 , w_9798 );
not ( w_9795 , w_9799 );
and ( w_9798 , w_9799 , \455_b0 );
or ( \4053_b1 , \2850_b1 , w_9801 );
not ( w_9801 , w_9802 );
and ( \4053_b0 , \2850_b0 , w_9803 );
and ( w_9802 ,  , w_9803 );
buf ( w_9801 , \296_b1 );
not ( w_9801 , w_9804 );
not (  , w_9805 );
and ( w_9804 , w_9805 , \296_b0 );
or ( \4054_b1 , \4053_b1 , w_9806 );
xor ( \4054_b0 , \4053_b0 , w_9808 );
not ( w_9808 , w_9809 );
and ( w_9809 , w_9806 , w_9807 );
buf ( w_9806 , \303_b1 );
not ( w_9806 , w_9810 );
not ( w_9807 , w_9811 );
and ( w_9810 , w_9811 , \303_b0 );
or ( \4055_b1 , \4052_b1 , \4054_b1 );
not ( \4054_b1 , w_9812 );
and ( \4055_b0 , \4052_b0 , w_9813 );
and ( w_9812 , w_9813 , \4054_b0 );
or ( \4056_b1 , \4048_b1 , \4055_b1 );
not ( \4055_b1 , w_9814 );
and ( \4056_b0 , \4048_b0 , w_9815 );
and ( w_9814 , w_9815 , \4055_b0 );
or ( \4057_b1 , \2850_b1 , \298_b1 );
not ( \298_b1 , w_9816 );
and ( \4057_b0 , \2850_b0 , w_9817 );
and ( w_9816 , w_9817 , \298_b0 );
or ( \4058_b1 , \2763_b1 , \296_b1 );
not ( \296_b1 , w_9818 );
and ( \4058_b0 , \2763_b0 , w_9819 );
and ( w_9818 , w_9819 , \296_b0 );
or ( \4059_b1 , \4057_b1 , w_9821 );
not ( w_9821 , w_9822 );
and ( \4059_b0 , \4057_b0 , w_9823 );
and ( w_9822 ,  , w_9823 );
buf ( w_9821 , \4058_b1 );
not ( w_9821 , w_9824 );
not (  , w_9825 );
and ( w_9824 , w_9825 , \4058_b0 );
or ( \4060_b1 , \4059_b1 , w_9826 );
xor ( \4060_b0 , \4059_b0 , w_9828 );
not ( w_9828 , w_9829 );
and ( w_9829 , w_9826 , w_9827 );
buf ( w_9826 , \303_b1 );
not ( w_9826 , w_9830 );
not ( w_9827 , w_9831 );
and ( w_9830 , w_9831 , \303_b0 );
or ( \4061_b1 , \4055_b1 , \4060_b1 );
not ( \4060_b1 , w_9832 );
and ( \4061_b0 , \4055_b0 , w_9833 );
and ( w_9832 , w_9833 , \4060_b0 );
or ( \4062_b1 , \4048_b1 , \4060_b1 );
not ( \4060_b1 , w_9834 );
and ( \4062_b0 , \4048_b0 , w_9835 );
and ( w_9834 , w_9835 , \4060_b0 );
or ( \4064_b1 , \4032_b1 , \4063_b1 );
not ( \4063_b1 , w_9836 );
and ( \4064_b0 , \4032_b0 , w_9837 );
and ( w_9836 , w_9837 , \4063_b0 );
or ( \4065_b1 , \3864_b1 , \3868_b1 );
xor ( \4065_b0 , \3864_b0 , w_9838 );
not ( w_9838 , w_9839 );
and ( w_9839 , \3868_b1 , \3868_b0 );
or ( \4066_b1 , \4065_b1 , \3873_b1 );
xor ( \4066_b0 , \4065_b0 , w_9840 );
not ( w_9840 , w_9841 );
and ( w_9841 , \3873_b1 , \3873_b0 );
or ( \4067_b1 , \3927_b1 , \3931_b1 );
xor ( \4067_b0 , \3927_b0 , w_9842 );
not ( w_9842 , w_9843 );
and ( w_9843 , \3931_b1 , \3931_b0 );
or ( \4068_b1 , \4067_b1 , \3936_b1 );
xor ( \4068_b0 , \4067_b0 , w_9844 );
not ( w_9844 , w_9845 );
and ( w_9845 , \3936_b1 , \3936_b0 );
or ( \4069_b1 , \4066_b1 , \4068_b1 );
not ( \4068_b1 , w_9846 );
and ( \4069_b0 , \4066_b0 , w_9847 );
and ( w_9846 , w_9847 , \4068_b0 );
or ( \4070_b1 , \3897_b1 , \3901_b1 );
xor ( \4070_b0 , \3897_b0 , w_9848 );
not ( w_9848 , w_9849 );
and ( w_9849 , \3901_b1 , \3901_b0 );
or ( \4071_b1 , \4070_b1 , \3906_b1 );
xor ( \4071_b0 , \4070_b0 , w_9850 );
not ( w_9850 , w_9851 );
and ( w_9851 , \3906_b1 , \3906_b0 );
or ( \4072_b1 , \4068_b1 , \4071_b1 );
not ( \4071_b1 , w_9852 );
and ( \4072_b0 , \4068_b0 , w_9853 );
and ( w_9852 , w_9853 , \4071_b0 );
or ( \4073_b1 , \4066_b1 , \4071_b1 );
not ( \4071_b1 , w_9854 );
and ( \4073_b0 , \4066_b0 , w_9855 );
and ( w_9854 , w_9855 , \4071_b0 );
or ( \4075_b1 , \4063_b1 , \4074_b1 );
not ( \4074_b1 , w_9856 );
and ( \4075_b0 , \4063_b0 , w_9857 );
and ( w_9856 , w_9857 , \4074_b0 );
or ( \4076_b1 , \4032_b1 , \4074_b1 );
not ( \4074_b1 , w_9858 );
and ( \4076_b0 , \4032_b0 , w_9859 );
and ( w_9858 , w_9859 , \4074_b0 );
or ( \4078_b1 , \3876_b1 , \3892_b1 );
xor ( \4078_b0 , \3876_b0 , w_9860 );
not ( w_9860 , w_9861 );
and ( w_9861 , \3892_b1 , \3892_b0 );
or ( \4079_b1 , \4078_b1 , \3909_b1 );
xor ( \4079_b0 , \4078_b0 , w_9862 );
not ( w_9862 , w_9863 );
and ( w_9863 , \3909_b1 , \3909_b0 );
or ( \4080_b1 , \3914_b1 , \3916_b1 );
xor ( \4080_b0 , \3914_b0 , w_9864 );
not ( w_9864 , w_9865 );
and ( w_9865 , \3916_b1 , \3916_b0 );
or ( \4081_b1 , \4080_b1 , \3919_b1 );
xor ( \4081_b0 , \4080_b0 , w_9866 );
not ( w_9866 , w_9867 );
and ( w_9867 , \3919_b1 , \3919_b0 );
or ( \4082_b1 , \4079_b1 , \4081_b1 );
not ( \4081_b1 , w_9868 );
and ( \4082_b0 , \4079_b0 , w_9869 );
and ( w_9868 , w_9869 , \4081_b0 );
or ( \4083_b1 , \3939_b1 , \3941_b1 );
xor ( \4083_b0 , \3939_b0 , w_9870 );
not ( w_9870 , w_9871 );
and ( w_9871 , \3941_b1 , \3941_b0 );
or ( \4084_b1 , \4083_b1 , \3944_b1 );
xor ( \4084_b0 , \4083_b0 , w_9872 );
not ( w_9872 , w_9873 );
and ( w_9873 , \3944_b1 , \3944_b0 );
or ( \4085_b1 , \4081_b1 , \4084_b1 );
not ( \4084_b1 , w_9874 );
and ( \4085_b0 , \4081_b0 , w_9875 );
and ( w_9874 , w_9875 , \4084_b0 );
or ( \4086_b1 , \4079_b1 , \4084_b1 );
not ( \4084_b1 , w_9876 );
and ( \4086_b0 , \4079_b0 , w_9877 );
and ( w_9876 , w_9877 , \4084_b0 );
or ( \4088_b1 , \4077_b1 , \4087_b1 );
not ( \4087_b1 , w_9878 );
and ( \4088_b0 , \4077_b0 , w_9879 );
and ( w_9878 , w_9879 , \4087_b0 );
or ( \4089_b1 , \3732_b1 , \3746_b1 );
xor ( \4089_b0 , \3732_b0 , w_9880 );
not ( w_9880 , w_9881 );
and ( w_9881 , \3746_b1 , \3746_b0 );
or ( \4090_b1 , \4089_b1 , \3751_b1 );
xor ( \4090_b0 , \4089_b0 , w_9882 );
not ( w_9882 , w_9883 );
and ( w_9883 , \3751_b1 , \3751_b0 );
or ( \4091_b1 , \4087_b1 , \4090_b1 );
not ( \4090_b1 , w_9884 );
and ( \4091_b0 , \4087_b0 , w_9885 );
and ( w_9884 , w_9885 , \4090_b0 );
or ( \4092_b1 , \4077_b1 , \4090_b1 );
not ( \4090_b1 , w_9886 );
and ( \4092_b0 , \4077_b0 , w_9887 );
and ( w_9886 , w_9887 , \4090_b0 );
or ( \4094_b1 , \3770_b1 , \3782_b1 );
xor ( \4094_b0 , \3770_b0 , w_9888 );
not ( w_9888 , w_9889 );
and ( w_9889 , \3782_b1 , \3782_b0 );
or ( \4095_b1 , \4094_b1 , \3799_b1 );
xor ( \4095_b0 , \4094_b0 , w_9890 );
not ( w_9890 , w_9891 );
and ( w_9891 , \3799_b1 , \3799_b0 );
or ( \4096_b1 , \3912_b1 , \3922_b1 );
xor ( \4096_b0 , \3912_b0 , w_9892 );
not ( w_9892 , w_9893 );
and ( w_9893 , \3922_b1 , \3922_b0 );
or ( \4097_b1 , \4096_b1 , \3947_b1 );
xor ( \4097_b0 , \4096_b0 , w_9894 );
not ( w_9894 , w_9895 );
and ( w_9895 , \3947_b1 , \3947_b0 );
or ( \4098_b1 , \4095_b1 , \4097_b1 );
not ( \4097_b1 , w_9896 );
and ( \4098_b0 , \4095_b0 , w_9897 );
and ( w_9896 , w_9897 , \4097_b0 );
or ( \4099_b1 , \3952_b1 , \3954_b1 );
xor ( \4099_b0 , \3952_b0 , w_9898 );
not ( w_9898 , w_9899 );
and ( w_9899 , \3954_b1 , \3954_b0 );
or ( \4100_b1 , \4099_b1 , \3957_b1 );
xor ( \4100_b0 , \4099_b0 , w_9900 );
not ( w_9900 , w_9901 );
and ( w_9901 , \3957_b1 , \3957_b0 );
or ( \4101_b1 , \4097_b1 , \4100_b1 );
not ( \4100_b1 , w_9902 );
and ( \4101_b0 , \4097_b0 , w_9903 );
and ( w_9902 , w_9903 , \4100_b0 );
or ( \4102_b1 , \4095_b1 , \4100_b1 );
not ( \4100_b1 , w_9904 );
and ( \4102_b0 , \4095_b0 , w_9905 );
and ( w_9904 , w_9905 , \4100_b0 );
or ( \4104_b1 , \4093_b1 , \4103_b1 );
not ( \4103_b1 , w_9906 );
and ( \4104_b0 , \4093_b0 , w_9907 );
and ( w_9906 , w_9907 , \4103_b0 );
or ( \4105_b1 , \3820_b1 , \3822_b1 );
xor ( \4105_b0 , \3820_b0 , w_9908 );
not ( w_9908 , w_9909 );
and ( w_9909 , \3822_b1 , \3822_b0 );
or ( \4106_b1 , \4105_b1 , \3825_b1 );
xor ( \4106_b0 , \4105_b0 , w_9910 );
not ( w_9910 , w_9911 );
and ( w_9911 , \3825_b1 , \3825_b0 );
or ( \4107_b1 , \4103_b1 , \4106_b1 );
not ( \4106_b1 , w_9912 );
and ( \4107_b0 , \4103_b0 , w_9913 );
and ( w_9912 , w_9913 , \4106_b0 );
or ( \4108_b1 , \4093_b1 , \4106_b1 );
not ( \4106_b1 , w_9914 );
and ( \4108_b0 , \4093_b0 , w_9915 );
and ( w_9914 , w_9915 , \4106_b0 );
or ( \4110_b1 , \3754_b1 , \3802_b1 );
xor ( \4110_b0 , \3754_b0 , w_9916 );
not ( w_9916 , w_9917 );
and ( w_9917 , \3802_b1 , \3802_b0 );
or ( \4111_b1 , \4110_b1 , \3815_b1 );
xor ( \4111_b0 , \4110_b0 , w_9918 );
not ( w_9918 , w_9919 );
and ( w_9919 , \3815_b1 , \3815_b0 );
or ( \4112_b1 , \3950_b1 , \3960_b1 );
xor ( \4112_b0 , \3950_b0 , w_9920 );
not ( w_9920 , w_9921 );
and ( w_9921 , \3960_b1 , \3960_b0 );
or ( \4113_b1 , \4112_b1 , \3963_b1 );
xor ( \4113_b0 , \4112_b0 , w_9922 );
not ( w_9922 , w_9923 );
and ( w_9923 , \3963_b1 , \3963_b0 );
or ( \4114_b1 , \4111_b1 , \4113_b1 );
not ( \4113_b1 , w_9924 );
and ( \4114_b0 , \4111_b0 , w_9925 );
and ( w_9924 , w_9925 , \4113_b0 );
or ( \4115_b1 , \4109_b1 , \4114_b1 );
not ( \4114_b1 , w_9926 );
and ( \4115_b0 , \4109_b0 , w_9927 );
and ( w_9926 , w_9927 , \4114_b0 );
or ( \4116_b1 , \3966_b1 , \3968_b1 );
xor ( \4116_b0 , \3966_b0 , w_9928 );
not ( w_9928 , w_9929 );
and ( w_9929 , \3968_b1 , \3968_b0 );
or ( \4117_b1 , \4116_b1 , \3970_b1 );
xor ( \4117_b0 , \4116_b0 , w_9930 );
not ( w_9930 , w_9931 );
and ( w_9931 , \3970_b1 , \3970_b0 );
or ( \4118_b1 , \4114_b1 , \4117_b1 );
not ( \4117_b1 , w_9932 );
and ( \4118_b0 , \4114_b0 , w_9933 );
and ( w_9932 , w_9933 , \4117_b0 );
or ( \4119_b1 , \4109_b1 , \4117_b1 );
not ( \4117_b1 , w_9934 );
and ( \4119_b0 , \4109_b0 , w_9935 );
and ( w_9934 , w_9935 , \4117_b0 );
or ( \4121_b1 , \3984_b1 , \4120_b1 );
not ( \4120_b1 , w_9936 );
and ( \4121_b0 , \3984_b0 , w_9937 );
and ( w_9936 , w_9937 , \4120_b0 );
or ( \4122_b1 , \3984_b1 , \4120_b1 );
xor ( \4122_b0 , \3984_b0 , w_9938 );
not ( w_9938 , w_9939 );
and ( w_9939 , \4120_b1 , \4120_b0 );
or ( \4123_b1 , \4109_b1 , \4114_b1 );
xor ( \4123_b0 , \4109_b0 , w_9940 );
not ( w_9940 , w_9941 );
and ( w_9941 , \4114_b1 , \4114_b0 );
or ( \4124_b1 , \4123_b1 , \4117_b1 );
xor ( \4124_b0 , \4123_b0 , w_9942 );
not ( w_9942 , w_9943 );
and ( w_9943 , \4117_b1 , \4117_b0 );
or ( \4125_b1 , \904_b1 , \1955_b1 );
not ( \1955_b1 , w_9944 );
and ( \4125_b0 , \904_b0 , w_9945 );
and ( w_9944 , w_9945 , \1955_b0 );
or ( \4126_b1 , \841_b1 , \1953_b1 );
not ( \1953_b1 , w_9946 );
and ( \4126_b0 , \841_b0 , w_9947 );
and ( w_9946 , w_9947 , \1953_b0 );
or ( \4127_b1 , \4125_b1 , w_9949 );
not ( w_9949 , w_9950 );
and ( \4127_b0 , \4125_b0 , w_9951 );
and ( w_9950 ,  , w_9951 );
buf ( w_9949 , \4126_b1 );
not ( w_9949 , w_9952 );
not (  , w_9953 );
and ( w_9952 , w_9953 , \4126_b0 );
or ( \4128_b1 , \4127_b1 , w_9954 );
xor ( \4128_b0 , \4127_b0 , w_9956 );
not ( w_9956 , w_9957 );
and ( w_9957 , w_9954 , w_9955 );
buf ( w_9954 , \1835_b1 );
not ( w_9954 , w_9958 );
not ( w_9955 , w_9959 );
and ( w_9958 , w_9959 , \1835_b0 );
or ( \4129_b1 , \1194_b1 , \1742_b1 );
not ( \1742_b1 , w_9960 );
and ( \4129_b0 , \1194_b0 , w_9961 );
and ( w_9960 , w_9961 , \1742_b0 );
or ( \4130_b1 , \1104_b1 , \1740_b1 );
not ( \1740_b1 , w_9962 );
and ( \4130_b0 , \1104_b0 , w_9963 );
and ( w_9962 , w_9963 , \1740_b0 );
or ( \4131_b1 , \4129_b1 , w_9965 );
not ( w_9965 , w_9966 );
and ( \4131_b0 , \4129_b0 , w_9967 );
and ( w_9966 ,  , w_9967 );
buf ( w_9965 , \4130_b1 );
not ( w_9965 , w_9968 );
not (  , w_9969 );
and ( w_9968 , w_9969 , \4130_b0 );
or ( \4132_b1 , \4131_b1 , w_9970 );
xor ( \4132_b0 , \4131_b0 , w_9972 );
not ( w_9972 , w_9973 );
and ( w_9973 , w_9970 , w_9971 );
buf ( w_9970 , \1610_b1 );
not ( w_9970 , w_9974 );
not ( w_9971 , w_9975 );
and ( w_9974 , w_9975 , \1610_b0 );
or ( \4133_b1 , \4128_b1 , \4132_b1 );
not ( \4132_b1 , w_9976 );
and ( \4133_b0 , \4128_b0 , w_9977 );
and ( w_9976 , w_9977 , \4132_b0 );
or ( \4134_b1 , \1304_b1 , \1476_b1 );
not ( \1476_b1 , w_9978 );
and ( \4134_b0 , \1304_b0 , w_9979 );
and ( w_9978 , w_9979 , \1476_b0 );
or ( \4135_b1 , \1299_b1 , \1474_b1 );
not ( \1474_b1 , w_9980 );
and ( \4135_b0 , \1299_b0 , w_9981 );
and ( w_9980 , w_9981 , \1474_b0 );
or ( \4136_b1 , \4134_b1 , w_9983 );
not ( w_9983 , w_9984 );
and ( \4136_b0 , \4134_b0 , w_9985 );
and ( w_9984 ,  , w_9985 );
buf ( w_9983 , \4135_b1 );
not ( w_9983 , w_9986 );
not (  , w_9987 );
and ( w_9986 , w_9987 , \4135_b0 );
or ( \4137_b1 , \4136_b1 , w_9988 );
xor ( \4137_b0 , \4136_b0 , w_9990 );
not ( w_9990 , w_9991 );
and ( w_9991 , w_9988 , w_9989 );
buf ( w_9988 , \1363_b1 );
not ( w_9988 , w_9992 );
not ( w_9989 , w_9993 );
and ( w_9992 , w_9993 , \1363_b0 );
or ( \4138_b1 , \4132_b1 , \4137_b1 );
not ( \4137_b1 , w_9994 );
and ( \4138_b0 , \4132_b0 , w_9995 );
and ( w_9994 , w_9995 , \4137_b0 );
or ( \4139_b1 , \4128_b1 , \4137_b1 );
not ( \4137_b1 , w_9996 );
and ( \4139_b0 , \4128_b0 , w_9997 );
and ( w_9996 , w_9997 , \4137_b0 );
or ( \4141_b1 , \1537_b1 , \1280_b1 );
not ( \1280_b1 , w_9998 );
and ( \4141_b0 , \1537_b0 , w_9999 );
and ( w_9998 , w_9999 , \1280_b0 );
or ( \4142_b1 , \1422_b1 , \1278_b1 );
not ( \1278_b1 , w_10000 );
and ( \4142_b0 , \1422_b0 , w_10001 );
and ( w_10000 , w_10001 , \1278_b0 );
or ( \4143_b1 , \4141_b1 , w_10003 );
not ( w_10003 , w_10004 );
and ( \4143_b0 , \4141_b0 , w_10005 );
and ( w_10004 ,  , w_10005 );
buf ( w_10003 , \4142_b1 );
not ( w_10003 , w_10006 );
not (  , w_10007 );
and ( w_10006 , w_10007 , \4142_b0 );
or ( \4144_b1 , \4143_b1 , w_10008 );
xor ( \4144_b0 , \4143_b0 , w_10010 );
not ( w_10010 , w_10011 );
and ( w_10011 , w_10008 , w_10009 );
buf ( w_10008 , \1177_b1 );
not ( w_10008 , w_10012 );
not ( w_10009 , w_10013 );
and ( w_10012 , w_10013 , \1177_b0 );
or ( \4145_b1 , \1778_b1 , \1062_b1 );
not ( \1062_b1 , w_10014 );
and ( \4145_b0 , \1778_b0 , w_10015 );
and ( w_10014 , w_10015 , \1062_b0 );
or ( \4146_b1 , \1770_b1 , \1060_b1 );
not ( \1060_b1 , w_10016 );
and ( \4146_b0 , \1770_b0 , w_10017 );
and ( w_10016 , w_10017 , \1060_b0 );
or ( \4147_b1 , \4145_b1 , w_10019 );
not ( w_10019 , w_10020 );
and ( \4147_b0 , \4145_b0 , w_10021 );
and ( w_10020 ,  , w_10021 );
buf ( w_10019 , \4146_b1 );
not ( w_10019 , w_10022 );
not (  , w_10023 );
and ( w_10022 , w_10023 , \4146_b0 );
or ( \4148_b1 , \4147_b1 , w_10024 );
xor ( \4148_b0 , \4147_b0 , w_10026 );
not ( w_10026 , w_10027 );
and ( w_10027 , w_10024 , w_10025 );
buf ( w_10024 , \984_b1 );
not ( w_10024 , w_10028 );
not ( w_10025 , w_10029 );
and ( w_10028 , w_10029 , \984_b0 );
or ( \4149_b1 , \4144_b1 , \4148_b1 );
not ( \4148_b1 , w_10030 );
and ( \4149_b0 , \4144_b0 , w_10031 );
and ( w_10030 , w_10031 , \4148_b0 );
or ( \4150_b1 , \2028_b1 , \912_b1 );
not ( \912_b1 , w_10032 );
and ( \4150_b0 , \2028_b0 , w_10033 );
and ( w_10032 , w_10033 , \912_b0 );
or ( \4151_b1 , \2023_b1 , \910_b1 );
not ( \910_b1 , w_10034 );
and ( \4151_b0 , \2023_b0 , w_10035 );
and ( w_10034 , w_10035 , \910_b0 );
or ( \4152_b1 , \4150_b1 , w_10037 );
not ( w_10037 , w_10038 );
and ( \4152_b0 , \4150_b0 , w_10039 );
and ( w_10038 ,  , w_10039 );
buf ( w_10037 , \4151_b1 );
not ( w_10037 , w_10040 );
not (  , w_10041 );
and ( w_10040 , w_10041 , \4151_b0 );
or ( \4153_b1 , \4152_b1 , w_10042 );
xor ( \4153_b0 , \4152_b0 , w_10044 );
not ( w_10044 , w_10045 );
and ( w_10045 , w_10042 , w_10043 );
buf ( w_10042 , \818_b1 );
not ( w_10042 , w_10046 );
not ( w_10043 , w_10047 );
and ( w_10046 , w_10047 , \818_b0 );
or ( \4154_b1 , \4148_b1 , \4153_b1 );
not ( \4153_b1 , w_10048 );
and ( \4154_b0 , \4148_b0 , w_10049 );
and ( w_10048 , w_10049 , \4153_b0 );
or ( \4155_b1 , \4144_b1 , \4153_b1 );
not ( \4153_b1 , w_10050 );
and ( \4155_b0 , \4144_b0 , w_10051 );
and ( w_10050 , w_10051 , \4153_b0 );
or ( \4157_b1 , \4140_b1 , \4156_b1 );
not ( \4156_b1 , w_10052 );
and ( \4157_b0 , \4140_b0 , w_10053 );
and ( w_10052 , w_10053 , \4156_b0 );
or ( \4158_b1 , \495_b1 , \2913_b1 );
not ( \2913_b1 , w_10054 );
and ( \4158_b0 , \495_b0 , w_10055 );
and ( w_10054 , w_10055 , \2913_b0 );
or ( \4159_b1 , \444_b1 , \2910_b1 );
not ( \2910_b1 , w_10056 );
and ( \4159_b0 , \444_b0 , w_10057 );
and ( w_10056 , w_10057 , \2910_b0 );
or ( \4160_b1 , \4158_b1 , w_10059 );
not ( w_10059 , w_10060 );
and ( \4160_b0 , \4158_b0 , w_10061 );
and ( w_10060 ,  , w_10061 );
buf ( w_10059 , \4159_b1 );
not ( w_10059 , w_10062 );
not (  , w_10063 );
and ( w_10062 , w_10063 , \4159_b0 );
or ( \4161_b1 , \4160_b1 , w_10064 );
xor ( \4161_b0 , \4160_b0 , w_10066 );
not ( w_10066 , w_10067 );
and ( w_10067 , w_10064 , w_10065 );
buf ( w_10064 , \2371_b1 );
not ( w_10064 , w_10068 );
not ( w_10065 , w_10069 );
and ( w_10068 , w_10069 , \2371_b0 );
or ( \4162_b1 , \621_b1 , \2550_b1 );
not ( \2550_b1 , w_10070 );
and ( \4162_b0 , \621_b0 , w_10071 );
and ( w_10070 , w_10071 , \2550_b0 );
or ( \4163_b1 , \593_b1 , \2548_b1 );
not ( \2548_b1 , w_10072 );
and ( \4163_b0 , \593_b0 , w_10073 );
and ( w_10072 , w_10073 , \2548_b0 );
or ( \4164_b1 , \4162_b1 , w_10075 );
not ( w_10075 , w_10076 );
and ( \4164_b0 , \4162_b0 , w_10077 );
and ( w_10076 ,  , w_10077 );
buf ( w_10075 , \4163_b1 );
not ( w_10075 , w_10078 );
not (  , w_10079 );
and ( w_10078 , w_10079 , \4163_b0 );
or ( \4165_b1 , \4164_b1 , w_10080 );
xor ( \4165_b0 , \4164_b0 , w_10082 );
not ( w_10082 , w_10083 );
and ( w_10083 , w_10080 , w_10081 );
buf ( w_10080 , \2374_b1 );
not ( w_10080 , w_10084 );
not ( w_10081 , w_10085 );
and ( w_10084 , w_10085 , \2374_b0 );
or ( \4166_b1 , \4161_b1 , \4165_b1 );
not ( \4165_b1 , w_10086 );
and ( \4166_b0 , \4161_b0 , w_10087 );
and ( w_10086 , w_10087 , \4165_b0 );
or ( \4167_b1 , \777_b1 , \2261_b1 );
not ( \2261_b1 , w_10088 );
and ( \4167_b0 , \777_b0 , w_10089 );
and ( w_10088 , w_10089 , \2261_b0 );
or ( \4168_b1 , \703_b1 , \2259_b1 );
not ( \2259_b1 , w_10090 );
and ( \4168_b0 , \703_b0 , w_10091 );
and ( w_10090 , w_10091 , \2259_b0 );
or ( \4169_b1 , \4167_b1 , w_10093 );
not ( w_10093 , w_10094 );
and ( \4169_b0 , \4167_b0 , w_10095 );
and ( w_10094 ,  , w_10095 );
buf ( w_10093 , \4168_b1 );
not ( w_10093 , w_10096 );
not (  , w_10097 );
and ( w_10096 , w_10097 , \4168_b0 );
or ( \4170_b1 , \4169_b1 , w_10098 );
xor ( \4170_b0 , \4169_b0 , w_10100 );
not ( w_10100 , w_10101 );
and ( w_10101 , w_10098 , w_10099 );
buf ( w_10098 , \2124_b1 );
not ( w_10098 , w_10102 );
not ( w_10099 , w_10103 );
and ( w_10102 , w_10103 , \2124_b0 );
or ( \4171_b1 , \4165_b1 , \4170_b1 );
not ( \4170_b1 , w_10104 );
and ( \4171_b0 , \4165_b0 , w_10105 );
and ( w_10104 , w_10105 , \4170_b0 );
or ( \4172_b1 , \4161_b1 , \4170_b1 );
not ( \4170_b1 , w_10106 );
and ( \4172_b0 , \4161_b0 , w_10107 );
and ( w_10106 , w_10107 , \4170_b0 );
or ( \4174_b1 , \4156_b1 , \4173_b1 );
not ( \4173_b1 , w_10108 );
and ( \4174_b0 , \4156_b0 , w_10109 );
and ( w_10108 , w_10109 , \4173_b0 );
or ( \4175_b1 , \4140_b1 , \4173_b1 );
not ( \4173_b1 , w_10110 );
and ( \4175_b0 , \4140_b0 , w_10111 );
and ( w_10110 , w_10111 , \4173_b0 );
or ( \4177_b1 , \3988_b1 , \3992_b1 );
xor ( \4177_b0 , \3988_b0 , w_10112 );
not ( w_10112 , w_10113 );
and ( w_10113 , \3992_b1 , \3992_b0 );
or ( \4178_b1 , \4177_b1 , \3997_b1 );
xor ( \4178_b0 , \4177_b0 , w_10114 );
not ( w_10114 , w_10115 );
and ( w_10115 , \3997_b1 , \3997_b0 );
or ( \4179_b1 , \4004_b1 , \4008_b1 );
xor ( \4179_b0 , \4004_b0 , w_10116 );
not ( w_10116 , w_10117 );
and ( w_10117 , \4008_b1 , \4008_b0 );
or ( \4180_b1 , \4179_b1 , \303_b1 );
xor ( \4180_b0 , \4179_b0 , w_10118 );
not ( w_10118 , w_10119 );
and ( w_10119 , \303_b1 , \303_b0 );
or ( \4181_b1 , \4178_b1 , \4180_b1 );
not ( \4180_b1 , w_10120 );
and ( \4181_b0 , \4178_b0 , w_10121 );
and ( w_10120 , w_10121 , \4180_b0 );
or ( \4182_b1 , \4017_b1 , \4021_b1 );
xor ( \4182_b0 , \4017_b0 , w_10122 );
not ( w_10122 , w_10123 );
and ( w_10123 , \4021_b1 , \4021_b0 );
or ( \4183_b1 , \4182_b1 , \4026_b1 );
xor ( \4183_b0 , \4182_b0 , w_10124 );
not ( w_10124 , w_10125 );
and ( w_10125 , \4026_b1 , \4026_b0 );
or ( \4184_b1 , \4180_b1 , \4183_b1 );
not ( \4183_b1 , w_10126 );
and ( \4184_b0 , \4180_b0 , w_10127 );
and ( w_10126 , w_10127 , \4183_b0 );
or ( \4185_b1 , \4178_b1 , \4183_b1 );
not ( \4183_b1 , w_10128 );
and ( \4185_b0 , \4178_b0 , w_10129 );
and ( w_10128 , w_10129 , \4183_b0 );
or ( \4187_b1 , \4176_b1 , \4186_b1 );
not ( \4186_b1 , w_10130 );
and ( \4187_b0 , \4176_b0 , w_10131 );
and ( w_10130 , w_10131 , \4186_b0 );
or ( \4188_b1 , \2305_b1 , \740_b1 );
not ( \740_b1 , w_10132 );
and ( \4188_b0 , \2305_b0 , w_10133 );
and ( w_10132 , w_10133 , \740_b0 );
or ( \4189_b1 , \2161_b1 , \738_b1 );
not ( \738_b1 , w_10134 );
and ( \4189_b0 , \2161_b0 , w_10135 );
and ( w_10134 , w_10135 , \738_b0 );
or ( \4190_b1 , \4188_b1 , w_10137 );
not ( w_10137 , w_10138 );
and ( \4190_b0 , \4188_b0 , w_10139 );
and ( w_10138 ,  , w_10139 );
buf ( w_10137 , \4189_b1 );
not ( w_10137 , w_10140 );
not (  , w_10141 );
and ( w_10140 , w_10141 , \4189_b0 );
or ( \4191_b1 , \4190_b1 , w_10142 );
xor ( \4191_b0 , \4190_b0 , w_10144 );
not ( w_10144 , w_10145 );
and ( w_10145 , w_10142 , w_10143 );
buf ( w_10142 , \668_b1 );
not ( w_10142 , w_10146 );
not ( w_10143 , w_10147 );
and ( w_10146 , w_10147 , \668_b0 );
or ( \4192_b1 , \2541_b1 , \604_b1 );
not ( \604_b1 , w_10148 );
and ( \4192_b0 , \2541_b0 , w_10149 );
and ( w_10148 , w_10149 , \604_b0 );
or ( \4193_b1 , \2532_b1 , \602_b1 );
not ( \602_b1 , w_10150 );
and ( \4193_b0 , \2532_b0 , w_10151 );
and ( w_10150 , w_10151 , \602_b0 );
or ( \4194_b1 , \4192_b1 , w_10153 );
not ( w_10153 , w_10154 );
and ( \4194_b0 , \4192_b0 , w_10155 );
and ( w_10154 ,  , w_10155 );
buf ( w_10153 , \4193_b1 );
not ( w_10153 , w_10156 );
not (  , w_10157 );
and ( w_10156 , w_10157 , \4193_b0 );
or ( \4195_b1 , \4194_b1 , w_10158 );
xor ( \4195_b0 , \4194_b0 , w_10160 );
not ( w_10160 , w_10161 );
and ( w_10161 , w_10158 , w_10159 );
buf ( w_10158 , \561_b1 );
not ( w_10158 , w_10162 );
not ( w_10159 , w_10163 );
and ( w_10162 , w_10163 , \561_b0 );
or ( \4196_b1 , \4191_b1 , \4195_b1 );
not ( \4195_b1 , w_10164 );
and ( \4196_b0 , \4191_b0 , w_10165 );
and ( w_10164 , w_10165 , \4195_b0 );
or ( \4197_b1 , \2850_b1 , \503_b1 );
not ( \503_b1 , w_10166 );
and ( \4197_b0 , \2850_b0 , w_10167 );
and ( w_10166 , w_10167 , \503_b0 );
or ( \4198_b1 , \2763_b1 , \501_b1 );
not ( \501_b1 , w_10168 );
and ( \4198_b0 , \2763_b0 , w_10169 );
and ( w_10168 , w_10169 , \501_b0 );
or ( \4199_b1 , \4197_b1 , w_10171 );
not ( w_10171 , w_10172 );
and ( \4199_b0 , \4197_b0 , w_10173 );
and ( w_10172 ,  , w_10173 );
buf ( w_10171 , \4198_b1 );
not ( w_10171 , w_10174 );
not (  , w_10175 );
and ( w_10174 , w_10175 , \4198_b0 );
or ( \4200_b1 , \4199_b1 , w_10176 );
xor ( \4200_b0 , \4199_b0 , w_10178 );
not ( w_10178 , w_10179 );
and ( w_10179 , w_10176 , w_10177 );
buf ( w_10176 , \455_b1 );
not ( w_10176 , w_10180 );
not ( w_10177 , w_10181 );
and ( w_10180 , w_10181 , \455_b0 );
or ( \4201_b1 , \4195_b1 , \4200_b1 );
not ( \4200_b1 , w_10182 );
and ( \4201_b0 , \4195_b0 , w_10183 );
and ( w_10182 , w_10183 , \4200_b0 );
or ( \4202_b1 , \4191_b1 , \4200_b1 );
not ( \4200_b1 , w_10184 );
and ( \4202_b0 , \4191_b0 , w_10185 );
and ( w_10184 , w_10185 , \4200_b0 );
or ( \4204_b1 , \4036_b1 , \4040_b1 );
xor ( \4204_b0 , \4036_b0 , w_10186 );
not ( w_10186 , w_10187 );
and ( w_10187 , \4040_b1 , \4040_b0 );
or ( \4205_b1 , \4204_b1 , \4045_b1 );
xor ( \4205_b0 , \4204_b0 , w_10188 );
not ( w_10188 , w_10189 );
and ( w_10189 , \4045_b1 , \4045_b0 );
or ( \4206_b1 , \4203_b1 , \4205_b1 );
not ( \4205_b1 , w_10190 );
and ( \4206_b0 , \4203_b0 , w_10191 );
and ( w_10190 , w_10191 , \4205_b0 );
or ( \4207_b1 , \4052_b1 , \4054_b1 );
xor ( \4207_b0 , \4052_b0 , w_10192 );
not ( w_10192 , w_10193 );
and ( w_10193 , \4054_b1 , \4054_b0 );
or ( \4208_b1 , \4205_b1 , \4207_b1 );
not ( \4207_b1 , w_10194 );
and ( \4208_b0 , \4205_b0 , w_10195 );
and ( w_10194 , w_10195 , \4207_b0 );
or ( \4209_b1 , \4203_b1 , \4207_b1 );
not ( \4207_b1 , w_10196 );
and ( \4209_b0 , \4203_b0 , w_10197 );
and ( w_10196 , w_10197 , \4207_b0 );
or ( \4211_b1 , \4186_b1 , \4210_b1 );
not ( \4210_b1 , w_10198 );
and ( \4211_b0 , \4186_b0 , w_10199 );
and ( w_10198 , w_10199 , \4210_b0 );
or ( \4212_b1 , \4176_b1 , \4210_b1 );
not ( \4210_b1 , w_10200 );
and ( \4212_b0 , \4176_b0 , w_10201 );
and ( w_10200 , w_10201 , \4210_b0 );
or ( \4214_b1 , \3880_b1 , \3884_b1 );
xor ( \4214_b0 , \3880_b0 , w_10202 );
not ( w_10202 , w_10203 );
and ( w_10203 , \3884_b1 , \3884_b0 );
or ( \4215_b1 , \4214_b1 , \3889_b1 );
xor ( \4215_b0 , \4214_b0 , w_10204 );
not ( w_10204 , w_10205 );
and ( w_10205 , \3889_b1 , \3889_b0 );
or ( \4216_b1 , \4048_b1 , \4055_b1 );
xor ( \4216_b0 , \4048_b0 , w_10206 );
not ( w_10206 , w_10207 );
and ( w_10207 , \4055_b1 , \4055_b0 );
or ( \4217_b1 , \4216_b1 , \4060_b1 );
xor ( \4217_b0 , \4216_b0 , w_10208 );
not ( w_10208 , w_10209 );
and ( w_10209 , \4060_b1 , \4060_b0 );
or ( \4218_b1 , \4215_b1 , \4217_b1 );
not ( \4217_b1 , w_10210 );
and ( \4218_b0 , \4215_b0 , w_10211 );
and ( w_10210 , w_10211 , \4217_b0 );
or ( \4219_b1 , \4066_b1 , \4068_b1 );
xor ( \4219_b0 , \4066_b0 , w_10212 );
not ( w_10212 , w_10213 );
and ( w_10213 , \4068_b1 , \4068_b0 );
or ( \4220_b1 , \4219_b1 , \4071_b1 );
xor ( \4220_b0 , \4219_b0 , w_10214 );
not ( w_10214 , w_10215 );
and ( w_10215 , \4071_b1 , \4071_b0 );
or ( \4221_b1 , \4217_b1 , \4220_b1 );
not ( \4220_b1 , w_10216 );
and ( \4221_b0 , \4217_b0 , w_10217 );
and ( w_10216 , w_10217 , \4220_b0 );
or ( \4222_b1 , \4215_b1 , \4220_b1 );
not ( \4220_b1 , w_10218 );
and ( \4222_b0 , \4215_b0 , w_10219 );
and ( w_10218 , w_10219 , \4220_b0 );
or ( \4224_b1 , \4213_b1 , \4223_b1 );
not ( \4223_b1 , w_10220 );
and ( \4224_b0 , \4213_b0 , w_10221 );
and ( w_10220 , w_10221 , \4223_b0 );
or ( \4225_b1 , \4079_b1 , \4081_b1 );
xor ( \4225_b0 , \4079_b0 , w_10222 );
not ( w_10222 , w_10223 );
and ( w_10223 , \4081_b1 , \4081_b0 );
or ( \4226_b1 , \4225_b1 , \4084_b1 );
xor ( \4226_b0 , \4225_b0 , w_10224 );
not ( w_10224 , w_10225 );
and ( w_10225 , \4084_b1 , \4084_b0 );
or ( \4227_b1 , \4223_b1 , \4226_b1 );
not ( \4226_b1 , w_10226 );
and ( \4227_b0 , \4223_b0 , w_10227 );
and ( w_10226 , w_10227 , \4226_b0 );
or ( \4228_b1 , \4213_b1 , \4226_b1 );
not ( \4226_b1 , w_10228 );
and ( \4228_b0 , \4213_b0 , w_10229 );
and ( w_10228 , w_10229 , \4226_b0 );
or ( \4230_b1 , \4077_b1 , \4087_b1 );
xor ( \4230_b0 , \4077_b0 , w_10230 );
not ( w_10230 , w_10231 );
and ( w_10231 , \4087_b1 , \4087_b0 );
or ( \4231_b1 , \4230_b1 , \4090_b1 );
xor ( \4231_b0 , \4230_b0 , w_10232 );
not ( w_10232 , w_10233 );
and ( w_10233 , \4090_b1 , \4090_b0 );
or ( \4232_b1 , \4229_b1 , \4231_b1 );
not ( \4231_b1 , w_10234 );
and ( \4232_b0 , \4229_b0 , w_10235 );
and ( w_10234 , w_10235 , \4231_b0 );
or ( \4233_b1 , \4095_b1 , \4097_b1 );
xor ( \4233_b0 , \4095_b0 , w_10236 );
not ( w_10236 , w_10237 );
and ( w_10237 , \4097_b1 , \4097_b0 );
or ( \4234_b1 , \4233_b1 , \4100_b1 );
xor ( \4234_b0 , \4233_b0 , w_10238 );
not ( w_10238 , w_10239 );
and ( w_10239 , \4100_b1 , \4100_b0 );
or ( \4235_b1 , \4231_b1 , \4234_b1 );
not ( \4234_b1 , w_10240 );
and ( \4235_b0 , \4231_b0 , w_10241 );
and ( w_10240 , w_10241 , \4234_b0 );
or ( \4236_b1 , \4229_b1 , \4234_b1 );
not ( \4234_b1 , w_10242 );
and ( \4236_b0 , \4229_b0 , w_10243 );
and ( w_10242 , w_10243 , \4234_b0 );
or ( \4238_b1 , \4093_b1 , \4103_b1 );
xor ( \4238_b0 , \4093_b0 , w_10244 );
not ( w_10244 , w_10245 );
and ( w_10245 , \4103_b1 , \4103_b0 );
or ( \4239_b1 , \4238_b1 , \4106_b1 );
xor ( \4239_b0 , \4238_b0 , w_10246 );
not ( w_10246 , w_10247 );
and ( w_10247 , \4106_b1 , \4106_b0 );
or ( \4240_b1 , \4237_b1 , \4239_b1 );
not ( \4239_b1 , w_10248 );
and ( \4240_b0 , \4237_b0 , w_10249 );
and ( w_10248 , w_10249 , \4239_b0 );
or ( \4241_b1 , \4111_b1 , \4113_b1 );
xor ( \4241_b0 , \4111_b0 , w_10250 );
not ( w_10250 , w_10251 );
and ( w_10251 , \4113_b1 , \4113_b0 );
or ( \4242_b1 , \4239_b1 , \4241_b1 );
not ( \4241_b1 , w_10252 );
and ( \4242_b0 , \4239_b0 , w_10253 );
and ( w_10252 , w_10253 , \4241_b0 );
or ( \4243_b1 , \4237_b1 , \4241_b1 );
not ( \4241_b1 , w_10254 );
and ( \4243_b0 , \4237_b0 , w_10255 );
and ( w_10254 , w_10255 , \4241_b0 );
or ( \4245_b1 , \4124_b1 , \4244_b1 );
not ( \4244_b1 , w_10256 );
and ( \4245_b0 , \4124_b0 , w_10257 );
and ( w_10256 , w_10257 , \4244_b0 );
or ( \4246_b1 , \4124_b1 , \4244_b1 );
xor ( \4246_b0 , \4124_b0 , w_10258 );
not ( w_10258 , w_10259 );
and ( w_10259 , \4244_b1 , \4244_b0 );
or ( \4247_b1 , \4237_b1 , \4239_b1 );
xor ( \4247_b0 , \4237_b0 , w_10260 );
not ( w_10260 , w_10261 );
and ( w_10261 , \4239_b1 , \4239_b0 );
or ( \4248_b1 , \4247_b1 , \4241_b1 );
xor ( \4248_b0 , \4247_b0 , w_10262 );
not ( w_10262 , w_10263 );
and ( w_10263 , \4241_b1 , \4241_b0 );
or ( \4249_b1 , \841_b1 , \2261_b1 );
not ( \2261_b1 , w_10264 );
and ( \4249_b0 , \841_b0 , w_10265 );
and ( w_10264 , w_10265 , \2261_b0 );
or ( \4250_b1 , \777_b1 , \2259_b1 );
not ( \2259_b1 , w_10266 );
and ( \4250_b0 , \777_b0 , w_10267 );
and ( w_10266 , w_10267 , \2259_b0 );
or ( \4251_b1 , \4249_b1 , w_10269 );
not ( w_10269 , w_10270 );
and ( \4251_b0 , \4249_b0 , w_10271 );
and ( w_10270 ,  , w_10271 );
buf ( w_10269 , \4250_b1 );
not ( w_10269 , w_10272 );
not (  , w_10273 );
and ( w_10272 , w_10273 , \4250_b0 );
or ( \4252_b1 , \4251_b1 , w_10274 );
xor ( \4252_b0 , \4251_b0 , w_10276 );
not ( w_10276 , w_10277 );
and ( w_10277 , w_10274 , w_10275 );
buf ( w_10274 , \2124_b1 );
not ( w_10274 , w_10278 );
not ( w_10275 , w_10279 );
and ( w_10278 , w_10279 , \2124_b0 );
or ( \4253_b1 , \1104_b1 , \1955_b1 );
not ( \1955_b1 , w_10280 );
and ( \4253_b0 , \1104_b0 , w_10281 );
and ( w_10280 , w_10281 , \1955_b0 );
or ( \4254_b1 , \904_b1 , \1953_b1 );
not ( \1953_b1 , w_10282 );
and ( \4254_b0 , \904_b0 , w_10283 );
and ( w_10282 , w_10283 , \1953_b0 );
or ( \4255_b1 , \4253_b1 , w_10285 );
not ( w_10285 , w_10286 );
and ( \4255_b0 , \4253_b0 , w_10287 );
and ( w_10286 ,  , w_10287 );
buf ( w_10285 , \4254_b1 );
not ( w_10285 , w_10288 );
not (  , w_10289 );
and ( w_10288 , w_10289 , \4254_b0 );
or ( \4256_b1 , \4255_b1 , w_10290 );
xor ( \4256_b0 , \4255_b0 , w_10292 );
not ( w_10292 , w_10293 );
and ( w_10293 , w_10290 , w_10291 );
buf ( w_10290 , \1835_b1 );
not ( w_10290 , w_10294 );
not ( w_10291 , w_10295 );
and ( w_10294 , w_10295 , \1835_b0 );
or ( \4257_b1 , \4252_b1 , \4256_b1 );
not ( \4256_b1 , w_10296 );
and ( \4257_b0 , \4252_b0 , w_10297 );
and ( w_10296 , w_10297 , \4256_b0 );
or ( \4258_b1 , \1299_b1 , \1742_b1 );
not ( \1742_b1 , w_10298 );
and ( \4258_b0 , \1299_b0 , w_10299 );
and ( w_10298 , w_10299 , \1742_b0 );
or ( \4259_b1 , \1194_b1 , \1740_b1 );
not ( \1740_b1 , w_10300 );
and ( \4259_b0 , \1194_b0 , w_10301 );
and ( w_10300 , w_10301 , \1740_b0 );
or ( \4260_b1 , \4258_b1 , w_10303 );
not ( w_10303 , w_10304 );
and ( \4260_b0 , \4258_b0 , w_10305 );
and ( w_10304 ,  , w_10305 );
buf ( w_10303 , \4259_b1 );
not ( w_10303 , w_10306 );
not (  , w_10307 );
and ( w_10306 , w_10307 , \4259_b0 );
or ( \4261_b1 , \4260_b1 , w_10308 );
xor ( \4261_b0 , \4260_b0 , w_10310 );
not ( w_10310 , w_10311 );
and ( w_10311 , w_10308 , w_10309 );
buf ( w_10308 , \1610_b1 );
not ( w_10308 , w_10312 );
not ( w_10309 , w_10313 );
and ( w_10312 , w_10313 , \1610_b0 );
or ( \4262_b1 , \4256_b1 , \4261_b1 );
not ( \4261_b1 , w_10314 );
and ( \4262_b0 , \4256_b0 , w_10315 );
and ( w_10314 , w_10315 , \4261_b0 );
or ( \4263_b1 , \4252_b1 , \4261_b1 );
not ( \4261_b1 , w_10316 );
and ( \4263_b0 , \4252_b0 , w_10317 );
and ( w_10316 , w_10317 , \4261_b0 );
or ( \4265_b1 , \1422_b1 , \1476_b1 );
not ( \1476_b1 , w_10318 );
and ( \4265_b0 , \1422_b0 , w_10319 );
and ( w_10318 , w_10319 , \1476_b0 );
or ( \4266_b1 , \1304_b1 , \1474_b1 );
not ( \1474_b1 , w_10320 );
and ( \4266_b0 , \1304_b0 , w_10321 );
and ( w_10320 , w_10321 , \1474_b0 );
or ( \4267_b1 , \4265_b1 , w_10323 );
not ( w_10323 , w_10324 );
and ( \4267_b0 , \4265_b0 , w_10325 );
and ( w_10324 ,  , w_10325 );
buf ( w_10323 , \4266_b1 );
not ( w_10323 , w_10326 );
not (  , w_10327 );
and ( w_10326 , w_10327 , \4266_b0 );
or ( \4268_b1 , \4267_b1 , w_10328 );
xor ( \4268_b0 , \4267_b0 , w_10330 );
not ( w_10330 , w_10331 );
and ( w_10331 , w_10328 , w_10329 );
buf ( w_10328 , \1363_b1 );
not ( w_10328 , w_10332 );
not ( w_10329 , w_10333 );
and ( w_10332 , w_10333 , \1363_b0 );
or ( \4269_b1 , \1770_b1 , \1280_b1 );
not ( \1280_b1 , w_10334 );
and ( \4269_b0 , \1770_b0 , w_10335 );
and ( w_10334 , w_10335 , \1280_b0 );
or ( \4270_b1 , \1537_b1 , \1278_b1 );
not ( \1278_b1 , w_10336 );
and ( \4270_b0 , \1537_b0 , w_10337 );
and ( w_10336 , w_10337 , \1278_b0 );
or ( \4271_b1 , \4269_b1 , w_10339 );
not ( w_10339 , w_10340 );
and ( \4271_b0 , \4269_b0 , w_10341 );
and ( w_10340 ,  , w_10341 );
buf ( w_10339 , \4270_b1 );
not ( w_10339 , w_10342 );
not (  , w_10343 );
and ( w_10342 , w_10343 , \4270_b0 );
or ( \4272_b1 , \4271_b1 , w_10344 );
xor ( \4272_b0 , \4271_b0 , w_10346 );
not ( w_10346 , w_10347 );
and ( w_10347 , w_10344 , w_10345 );
buf ( w_10344 , \1177_b1 );
not ( w_10344 , w_10348 );
not ( w_10345 , w_10349 );
and ( w_10348 , w_10349 , \1177_b0 );
or ( \4273_b1 , \4268_b1 , \4272_b1 );
not ( \4272_b1 , w_10350 );
and ( \4273_b0 , \4268_b0 , w_10351 );
and ( w_10350 , w_10351 , \4272_b0 );
or ( \4274_b1 , \2023_b1 , \1062_b1 );
not ( \1062_b1 , w_10352 );
and ( \4274_b0 , \2023_b0 , w_10353 );
and ( w_10352 , w_10353 , \1062_b0 );
or ( \4275_b1 , \1778_b1 , \1060_b1 );
not ( \1060_b1 , w_10354 );
and ( \4275_b0 , \1778_b0 , w_10355 );
and ( w_10354 , w_10355 , \1060_b0 );
or ( \4276_b1 , \4274_b1 , w_10357 );
not ( w_10357 , w_10358 );
and ( \4276_b0 , \4274_b0 , w_10359 );
and ( w_10358 ,  , w_10359 );
buf ( w_10357 , \4275_b1 );
not ( w_10357 , w_10360 );
not (  , w_10361 );
and ( w_10360 , w_10361 , \4275_b0 );
or ( \4277_b1 , \4276_b1 , w_10362 );
xor ( \4277_b0 , \4276_b0 , w_10364 );
not ( w_10364 , w_10365 );
and ( w_10365 , w_10362 , w_10363 );
buf ( w_10362 , \984_b1 );
not ( w_10362 , w_10366 );
not ( w_10363 , w_10367 );
and ( w_10366 , w_10367 , \984_b0 );
or ( \4278_b1 , \4272_b1 , \4277_b1 );
not ( \4277_b1 , w_10368 );
and ( \4278_b0 , \4272_b0 , w_10369 );
and ( w_10368 , w_10369 , \4277_b0 );
or ( \4279_b1 , \4268_b1 , \4277_b1 );
not ( \4277_b1 , w_10370 );
and ( \4279_b0 , \4268_b0 , w_10371 );
and ( w_10370 , w_10371 , \4277_b0 );
or ( \4281_b1 , \4264_b1 , \4280_b1 );
not ( \4280_b1 , w_10372 );
and ( \4281_b0 , \4264_b0 , w_10373 );
and ( w_10372 , w_10373 , \4280_b0 );
or ( \4282_b1 , \593_b1 , \2913_b1 );
not ( \2913_b1 , w_10374 );
and ( \4282_b0 , \593_b0 , w_10375 );
and ( w_10374 , w_10375 , \2913_b0 );
or ( \4283_b1 , \495_b1 , \2910_b1 );
not ( \2910_b1 , w_10376 );
and ( \4283_b0 , \495_b0 , w_10377 );
and ( w_10376 , w_10377 , \2910_b0 );
or ( \4284_b1 , \4282_b1 , w_10379 );
not ( w_10379 , w_10380 );
and ( \4284_b0 , \4282_b0 , w_10381 );
and ( w_10380 ,  , w_10381 );
buf ( w_10379 , \4283_b1 );
not ( w_10379 , w_10382 );
not (  , w_10383 );
and ( w_10382 , w_10383 , \4283_b0 );
or ( \4285_b1 , \4284_b1 , w_10384 );
xor ( \4285_b0 , \4284_b0 , w_10386 );
not ( w_10386 , w_10387 );
and ( w_10387 , w_10384 , w_10385 );
buf ( w_10384 , \2371_b1 );
not ( w_10384 , w_10388 );
not ( w_10385 , w_10389 );
and ( w_10388 , w_10389 , \2371_b0 );
or ( \4286_b1 , \703_b1 , \2550_b1 );
not ( \2550_b1 , w_10390 );
and ( \4286_b0 , \703_b0 , w_10391 );
and ( w_10390 , w_10391 , \2550_b0 );
or ( \4287_b1 , \621_b1 , \2548_b1 );
not ( \2548_b1 , w_10392 );
and ( \4287_b0 , \621_b0 , w_10393 );
and ( w_10392 , w_10393 , \2548_b0 );
or ( \4288_b1 , \4286_b1 , w_10395 );
not ( w_10395 , w_10396 );
and ( \4288_b0 , \4286_b0 , w_10397 );
and ( w_10396 ,  , w_10397 );
buf ( w_10395 , \4287_b1 );
not ( w_10395 , w_10398 );
not (  , w_10399 );
and ( w_10398 , w_10399 , \4287_b0 );
or ( \4289_b1 , \4288_b1 , w_10400 );
xor ( \4289_b0 , \4288_b0 , w_10402 );
not ( w_10402 , w_10403 );
and ( w_10403 , w_10400 , w_10401 );
buf ( w_10400 , \2374_b1 );
not ( w_10400 , w_10404 );
not ( w_10401 , w_10405 );
and ( w_10404 , w_10405 , \2374_b0 );
or ( \4290_b1 , \4285_b1 , \4289_b1 );
not ( \4289_b1 , w_10406 );
and ( \4290_b0 , \4285_b0 , w_10407 );
and ( w_10406 , w_10407 , \4289_b0 );
or ( \4291_b1 , \4289_b1 , \455_b1 );
not ( \455_b1 , w_10408 );
and ( \4291_b0 , \4289_b0 , w_10409 );
and ( w_10408 , w_10409 , \455_b0 );
or ( \4292_b1 , \4285_b1 , \455_b1 );
not ( \455_b1 , w_10410 );
and ( \4292_b0 , \4285_b0 , w_10411 );
and ( w_10410 , w_10411 , \455_b0 );
or ( \4294_b1 , \4280_b1 , \4293_b1 );
not ( \4293_b1 , w_10412 );
and ( \4294_b0 , \4280_b0 , w_10413 );
and ( w_10412 , w_10413 , \4293_b0 );
or ( \4295_b1 , \4264_b1 , \4293_b1 );
not ( \4293_b1 , w_10414 );
and ( \4295_b0 , \4264_b0 , w_10415 );
and ( w_10414 , w_10415 , \4293_b0 );
or ( \4297_b1 , \2161_b1 , \912_b1 );
not ( \912_b1 , w_10416 );
and ( \4297_b0 , \2161_b0 , w_10417 );
and ( w_10416 , w_10417 , \912_b0 );
or ( \4298_b1 , \2028_b1 , \910_b1 );
not ( \910_b1 , w_10418 );
and ( \4298_b0 , \2028_b0 , w_10419 );
and ( w_10418 , w_10419 , \910_b0 );
or ( \4299_b1 , \4297_b1 , w_10421 );
not ( w_10421 , w_10422 );
and ( \4299_b0 , \4297_b0 , w_10423 );
and ( w_10422 ,  , w_10423 );
buf ( w_10421 , \4298_b1 );
not ( w_10421 , w_10424 );
not (  , w_10425 );
and ( w_10424 , w_10425 , \4298_b0 );
or ( \4300_b1 , \4299_b1 , w_10426 );
xor ( \4300_b0 , \4299_b0 , w_10428 );
not ( w_10428 , w_10429 );
and ( w_10429 , w_10426 , w_10427 );
buf ( w_10426 , \818_b1 );
not ( w_10426 , w_10430 );
not ( w_10427 , w_10431 );
and ( w_10430 , w_10431 , \818_b0 );
or ( \4301_b1 , \2532_b1 , \740_b1 );
not ( \740_b1 , w_10432 );
and ( \4301_b0 , \2532_b0 , w_10433 );
and ( w_10432 , w_10433 , \740_b0 );
or ( \4302_b1 , \2305_b1 , \738_b1 );
not ( \738_b1 , w_10434 );
and ( \4302_b0 , \2305_b0 , w_10435 );
and ( w_10434 , w_10435 , \738_b0 );
or ( \4303_b1 , \4301_b1 , w_10437 );
not ( w_10437 , w_10438 );
and ( \4303_b0 , \4301_b0 , w_10439 );
and ( w_10438 ,  , w_10439 );
buf ( w_10437 , \4302_b1 );
not ( w_10437 , w_10440 );
not (  , w_10441 );
and ( w_10440 , w_10441 , \4302_b0 );
or ( \4304_b1 , \4303_b1 , w_10442 );
xor ( \4304_b0 , \4303_b0 , w_10444 );
not ( w_10444 , w_10445 );
and ( w_10445 , w_10442 , w_10443 );
buf ( w_10442 , \668_b1 );
not ( w_10442 , w_10446 );
not ( w_10443 , w_10447 );
and ( w_10446 , w_10447 , \668_b0 );
or ( \4305_b1 , \4300_b1 , \4304_b1 );
not ( \4304_b1 , w_10448 );
and ( \4305_b0 , \4300_b0 , w_10449 );
and ( w_10448 , w_10449 , \4304_b0 );
or ( \4306_b1 , \2763_b1 , \604_b1 );
not ( \604_b1 , w_10450 );
and ( \4306_b0 , \2763_b0 , w_10451 );
and ( w_10450 , w_10451 , \604_b0 );
or ( \4307_b1 , \2541_b1 , \602_b1 );
not ( \602_b1 , w_10452 );
and ( \4307_b0 , \2541_b0 , w_10453 );
and ( w_10452 , w_10453 , \602_b0 );
or ( \4308_b1 , \4306_b1 , w_10455 );
not ( w_10455 , w_10456 );
and ( \4308_b0 , \4306_b0 , w_10457 );
and ( w_10456 ,  , w_10457 );
buf ( w_10455 , \4307_b1 );
not ( w_10455 , w_10458 );
not (  , w_10459 );
and ( w_10458 , w_10459 , \4307_b0 );
or ( \4309_b1 , \4308_b1 , w_10460 );
xor ( \4309_b0 , \4308_b0 , w_10462 );
not ( w_10462 , w_10463 );
and ( w_10463 , w_10460 , w_10461 );
buf ( w_10460 , \561_b1 );
not ( w_10460 , w_10464 );
not ( w_10461 , w_10465 );
and ( w_10464 , w_10465 , \561_b0 );
or ( \4310_b1 , \4304_b1 , \4309_b1 );
not ( \4309_b1 , w_10466 );
and ( \4310_b0 , \4304_b0 , w_10467 );
and ( w_10466 , w_10467 , \4309_b0 );
or ( \4311_b1 , \4300_b1 , \4309_b1 );
not ( \4309_b1 , w_10468 );
and ( \4311_b0 , \4300_b0 , w_10469 );
and ( w_10468 , w_10469 , \4309_b0 );
or ( \4313_b1 , \4144_b1 , \4148_b1 );
xor ( \4313_b0 , \4144_b0 , w_10470 );
not ( w_10470 , w_10471 );
and ( w_10471 , \4148_b1 , \4148_b0 );
or ( \4314_b1 , \4313_b1 , \4153_b1 );
xor ( \4314_b0 , \4313_b0 , w_10472 );
not ( w_10472 , w_10473 );
and ( w_10473 , \4153_b1 , \4153_b0 );
or ( \4315_b1 , \4312_b1 , \4314_b1 );
not ( \4314_b1 , w_10474 );
and ( \4315_b0 , \4312_b0 , w_10475 );
and ( w_10474 , w_10475 , \4314_b0 );
or ( \4316_b1 , \4191_b1 , \4195_b1 );
xor ( \4316_b0 , \4191_b0 , w_10476 );
not ( w_10476 , w_10477 );
and ( w_10477 , \4195_b1 , \4195_b0 );
or ( \4317_b1 , \4316_b1 , \4200_b1 );
xor ( \4317_b0 , \4316_b0 , w_10478 );
not ( w_10478 , w_10479 );
and ( w_10479 , \4200_b1 , \4200_b0 );
or ( \4318_b1 , \4314_b1 , \4317_b1 );
not ( \4317_b1 , w_10480 );
and ( \4318_b0 , \4314_b0 , w_10481 );
and ( w_10480 , w_10481 , \4317_b0 );
or ( \4319_b1 , \4312_b1 , \4317_b1 );
not ( \4317_b1 , w_10482 );
and ( \4319_b0 , \4312_b0 , w_10483 );
and ( w_10482 , w_10483 , \4317_b0 );
or ( \4321_b1 , \4296_b1 , \4320_b1 );
not ( \4320_b1 , w_10484 );
and ( \4321_b0 , \4296_b0 , w_10485 );
and ( w_10484 , w_10485 , \4320_b0 );
or ( \4322_b1 , \4128_b1 , \4132_b1 );
xor ( \4322_b0 , \4128_b0 , w_10486 );
not ( w_10486 , w_10487 );
and ( w_10487 , \4132_b1 , \4132_b0 );
or ( \4323_b1 , \4322_b1 , \4137_b1 );
xor ( \4323_b0 , \4322_b0 , w_10488 );
not ( w_10488 , w_10489 );
and ( w_10489 , \4137_b1 , \4137_b0 );
or ( \4324_b1 , \4161_b1 , \4165_b1 );
xor ( \4324_b0 , \4161_b0 , w_10490 );
not ( w_10490 , w_10491 );
and ( w_10491 , \4165_b1 , \4165_b0 );
or ( \4325_b1 , \4324_b1 , \4170_b1 );
xor ( \4325_b0 , \4324_b0 , w_10492 );
not ( w_10492 , w_10493 );
and ( w_10493 , \4170_b1 , \4170_b0 );
or ( \4326_b1 , \4323_b1 , \4325_b1 );
not ( \4325_b1 , w_10494 );
and ( \4326_b0 , \4323_b0 , w_10495 );
and ( w_10494 , w_10495 , \4325_b0 );
or ( \4327_b1 , \4320_b1 , \4326_b1 );
not ( \4326_b1 , w_10496 );
and ( \4327_b0 , \4320_b0 , w_10497 );
and ( w_10496 , w_10497 , \4326_b0 );
or ( \4328_b1 , \4296_b1 , \4326_b1 );
not ( \4326_b1 , w_10498 );
and ( \4328_b0 , \4296_b0 , w_10499 );
and ( w_10498 , w_10499 , \4326_b0 );
or ( \4330_b1 , \4140_b1 , \4156_b1 );
xor ( \4330_b0 , \4140_b0 , w_10500 );
not ( w_10500 , w_10501 );
and ( w_10501 , \4156_b1 , \4156_b0 );
or ( \4331_b1 , \4330_b1 , \4173_b1 );
xor ( \4331_b0 , \4330_b0 , w_10502 );
not ( w_10502 , w_10503 );
and ( w_10503 , \4173_b1 , \4173_b0 );
or ( \4332_b1 , \4178_b1 , \4180_b1 );
xor ( \4332_b0 , \4178_b0 , w_10504 );
not ( w_10504 , w_10505 );
and ( w_10505 , \4180_b1 , \4180_b0 );
or ( \4333_b1 , \4332_b1 , \4183_b1 );
xor ( \4333_b0 , \4332_b0 , w_10506 );
not ( w_10506 , w_10507 );
and ( w_10507 , \4183_b1 , \4183_b0 );
or ( \4334_b1 , \4331_b1 , \4333_b1 );
not ( \4333_b1 , w_10508 );
and ( \4334_b0 , \4331_b0 , w_10509 );
and ( w_10508 , w_10509 , \4333_b0 );
or ( \4335_b1 , \4203_b1 , \4205_b1 );
xor ( \4335_b0 , \4203_b0 , w_10510 );
not ( w_10510 , w_10511 );
and ( w_10511 , \4205_b1 , \4205_b0 );
or ( \4336_b1 , \4335_b1 , \4207_b1 );
xor ( \4336_b0 , \4335_b0 , w_10512 );
not ( w_10512 , w_10513 );
and ( w_10513 , \4207_b1 , \4207_b0 );
or ( \4337_b1 , \4333_b1 , \4336_b1 );
not ( \4336_b1 , w_10514 );
and ( \4337_b0 , \4333_b0 , w_10515 );
and ( w_10514 , w_10515 , \4336_b0 );
or ( \4338_b1 , \4331_b1 , \4336_b1 );
not ( \4336_b1 , w_10516 );
and ( \4338_b0 , \4331_b0 , w_10517 );
and ( w_10516 , w_10517 , \4336_b0 );
or ( \4340_b1 , \4329_b1 , \4339_b1 );
not ( \4339_b1 , w_10518 );
and ( \4340_b0 , \4329_b0 , w_10519 );
and ( w_10518 , w_10519 , \4339_b0 );
or ( \4341_b1 , \4000_b1 , \4012_b1 );
xor ( \4341_b0 , \4000_b0 , w_10520 );
not ( w_10520 , w_10521 );
and ( w_10521 , \4012_b1 , \4012_b0 );
or ( \4342_b1 , \4341_b1 , \4029_b1 );
xor ( \4342_b0 , \4341_b0 , w_10522 );
not ( w_10522 , w_10523 );
and ( w_10523 , \4029_b1 , \4029_b0 );
or ( \4343_b1 , \4339_b1 , \4342_b1 );
not ( \4342_b1 , w_10524 );
and ( \4343_b0 , \4339_b0 , w_10525 );
and ( w_10524 , w_10525 , \4342_b0 );
or ( \4344_b1 , \4329_b1 , \4342_b1 );
not ( \4342_b1 , w_10526 );
and ( \4344_b0 , \4329_b0 , w_10527 );
and ( w_10526 , w_10527 , \4342_b0 );
or ( \4346_b1 , \4176_b1 , \4186_b1 );
xor ( \4346_b0 , \4176_b0 , w_10528 );
not ( w_10528 , w_10529 );
and ( w_10529 , \4186_b1 , \4186_b0 );
or ( \4347_b1 , \4346_b1 , \4210_b1 );
xor ( \4347_b0 , \4346_b0 , w_10530 );
not ( w_10530 , w_10531 );
and ( w_10531 , \4210_b1 , \4210_b0 );
or ( \4348_b1 , \4215_b1 , \4217_b1 );
xor ( \4348_b0 , \4215_b0 , w_10532 );
not ( w_10532 , w_10533 );
and ( w_10533 , \4217_b1 , \4217_b0 );
or ( \4349_b1 , \4348_b1 , \4220_b1 );
xor ( \4349_b0 , \4348_b0 , w_10534 );
not ( w_10534 , w_10535 );
and ( w_10535 , \4220_b1 , \4220_b0 );
or ( \4350_b1 , \4347_b1 , \4349_b1 );
not ( \4349_b1 , w_10536 );
and ( \4350_b0 , \4347_b0 , w_10537 );
and ( w_10536 , w_10537 , \4349_b0 );
or ( \4351_b1 , \4345_b1 , \4350_b1 );
not ( \4350_b1 , w_10538 );
and ( \4351_b0 , \4345_b0 , w_10539 );
and ( w_10538 , w_10539 , \4350_b0 );
or ( \4352_b1 , \4032_b1 , \4063_b1 );
xor ( \4352_b0 , \4032_b0 , w_10540 );
not ( w_10540 , w_10541 );
and ( w_10541 , \4063_b1 , \4063_b0 );
or ( \4353_b1 , \4352_b1 , \4074_b1 );
xor ( \4353_b0 , \4352_b0 , w_10542 );
not ( w_10542 , w_10543 );
and ( w_10543 , \4074_b1 , \4074_b0 );
or ( \4354_b1 , \4350_b1 , \4353_b1 );
not ( \4353_b1 , w_10544 );
and ( \4354_b0 , \4350_b0 , w_10545 );
and ( w_10544 , w_10545 , \4353_b0 );
or ( \4355_b1 , \4345_b1 , \4353_b1 );
not ( \4353_b1 , w_10546 );
and ( \4355_b0 , \4345_b0 , w_10547 );
and ( w_10546 , w_10547 , \4353_b0 );
or ( \4357_b1 , \4229_b1 , \4231_b1 );
xor ( \4357_b0 , \4229_b0 , w_10548 );
not ( w_10548 , w_10549 );
and ( w_10549 , \4231_b1 , \4231_b0 );
or ( \4358_b1 , \4357_b1 , \4234_b1 );
xor ( \4358_b0 , \4357_b0 , w_10550 );
not ( w_10550 , w_10551 );
and ( w_10551 , \4234_b1 , \4234_b0 );
or ( \4359_b1 , \4356_b1 , \4358_b1 );
not ( \4358_b1 , w_10552 );
and ( \4359_b0 , \4356_b0 , w_10553 );
and ( w_10552 , w_10553 , \4358_b0 );
or ( \4360_b1 , \4248_b1 , \4359_b1 );
not ( \4359_b1 , w_10554 );
and ( \4360_b0 , \4248_b0 , w_10555 );
and ( w_10554 , w_10555 , \4359_b0 );
or ( \4361_b1 , \4248_b1 , \4359_b1 );
xor ( \4361_b0 , \4248_b0 , w_10556 );
not ( w_10556 , w_10557 );
and ( w_10557 , \4359_b1 , \4359_b0 );
or ( \4362_b1 , \4356_b1 , \4358_b1 );
xor ( \4362_b0 , \4356_b0 , w_10558 );
not ( w_10558 , w_10559 );
and ( w_10559 , \4358_b1 , \4358_b0 );
or ( \4363_b1 , \4345_b1 , \4350_b1 );
xor ( \4363_b0 , \4345_b0 , w_10560 );
not ( w_10560 , w_10561 );
and ( w_10561 , \4350_b1 , \4350_b0 );
or ( \4364_b1 , \4363_b1 , \4353_b1 );
xor ( \4364_b0 , \4363_b0 , w_10562 );
not ( w_10562 , w_10563 );
and ( w_10563 , \4353_b1 , \4353_b0 );
or ( \4365_b1 , \4213_b1 , \4223_b1 );
xor ( \4365_b0 , \4213_b0 , w_10564 );
not ( w_10564 , w_10565 );
and ( w_10565 , \4223_b1 , \4223_b0 );
or ( \4366_b1 , \4365_b1 , \4226_b1 );
xor ( \4366_b0 , \4365_b0 , w_10566 );
not ( w_10566 , w_10567 );
and ( w_10567 , \4226_b1 , \4226_b0 );
or ( \4367_b1 , \4364_b1 , \4366_b1 );
not ( \4366_b1 , w_10568 );
and ( \4367_b0 , \4364_b0 , w_10569 );
and ( w_10568 , w_10569 , \4366_b0 );
or ( \4368_b1 , \4362_b1 , \4367_b1 );
not ( \4367_b1 , w_10570 );
and ( \4368_b0 , \4362_b0 , w_10571 );
and ( w_10570 , w_10571 , \4367_b0 );
or ( \4369_b1 , \4362_b1 , \4367_b1 );
xor ( \4369_b0 , \4362_b0 , w_10572 );
not ( w_10572 , w_10573 );
and ( w_10573 , \4367_b1 , \4367_b0 );
or ( \4370_b1 , \4364_b1 , \4366_b1 );
xor ( \4370_b0 , \4364_b0 , w_10574 );
not ( w_10574 , w_10575 );
and ( w_10575 , \4366_b1 , \4366_b0 );
or ( \4371_b1 , \621_b1 , \2913_b1 );
not ( \2913_b1 , w_10576 );
and ( \4371_b0 , \621_b0 , w_10577 );
and ( w_10576 , w_10577 , \2913_b0 );
or ( \4372_b1 , \593_b1 , \2910_b1 );
not ( \2910_b1 , w_10578 );
and ( \4372_b0 , \593_b0 , w_10579 );
and ( w_10578 , w_10579 , \2910_b0 );
or ( \4373_b1 , \4371_b1 , w_10581 );
not ( w_10581 , w_10582 );
and ( \4373_b0 , \4371_b0 , w_10583 );
and ( w_10582 ,  , w_10583 );
buf ( w_10581 , \4372_b1 );
not ( w_10581 , w_10584 );
not (  , w_10585 );
and ( w_10584 , w_10585 , \4372_b0 );
or ( \4374_b1 , \4373_b1 , w_10586 );
xor ( \4374_b0 , \4373_b0 , w_10588 );
not ( w_10588 , w_10589 );
and ( w_10589 , w_10586 , w_10587 );
buf ( w_10586 , \2371_b1 );
not ( w_10586 , w_10590 );
not ( w_10587 , w_10591 );
and ( w_10590 , w_10591 , \2371_b0 );
or ( \4375_b1 , \777_b1 , \2550_b1 );
not ( \2550_b1 , w_10592 );
and ( \4375_b0 , \777_b0 , w_10593 );
and ( w_10592 , w_10593 , \2550_b0 );
or ( \4376_b1 , \703_b1 , \2548_b1 );
not ( \2548_b1 , w_10594 );
and ( \4376_b0 , \703_b0 , w_10595 );
and ( w_10594 , w_10595 , \2548_b0 );
or ( \4377_b1 , \4375_b1 , w_10597 );
not ( w_10597 , w_10598 );
and ( \4377_b0 , \4375_b0 , w_10599 );
and ( w_10598 ,  , w_10599 );
buf ( w_10597 , \4376_b1 );
not ( w_10597 , w_10600 );
not (  , w_10601 );
and ( w_10600 , w_10601 , \4376_b0 );
or ( \4378_b1 , \4377_b1 , w_10602 );
xor ( \4378_b0 , \4377_b0 , w_10604 );
not ( w_10604 , w_10605 );
and ( w_10605 , w_10602 , w_10603 );
buf ( w_10602 , \2374_b1 );
not ( w_10602 , w_10606 );
not ( w_10603 , w_10607 );
and ( w_10606 , w_10607 , \2374_b0 );
or ( \4379_b1 , \4374_b1 , \4378_b1 );
not ( \4378_b1 , w_10608 );
and ( \4379_b0 , \4374_b0 , w_10609 );
and ( w_10608 , w_10609 , \4378_b0 );
or ( \4380_b1 , \904_b1 , \2261_b1 );
not ( \2261_b1 , w_10610 );
and ( \4380_b0 , \904_b0 , w_10611 );
and ( w_10610 , w_10611 , \2261_b0 );
or ( \4381_b1 , \841_b1 , \2259_b1 );
not ( \2259_b1 , w_10612 );
and ( \4381_b0 , \841_b0 , w_10613 );
and ( w_10612 , w_10613 , \2259_b0 );
or ( \4382_b1 , \4380_b1 , w_10615 );
not ( w_10615 , w_10616 );
and ( \4382_b0 , \4380_b0 , w_10617 );
and ( w_10616 ,  , w_10617 );
buf ( w_10615 , \4381_b1 );
not ( w_10615 , w_10618 );
not (  , w_10619 );
and ( w_10618 , w_10619 , \4381_b0 );
or ( \4383_b1 , \4382_b1 , w_10620 );
xor ( \4383_b0 , \4382_b0 , w_10622 );
not ( w_10622 , w_10623 );
and ( w_10623 , w_10620 , w_10621 );
buf ( w_10620 , \2124_b1 );
not ( w_10620 , w_10624 );
not ( w_10621 , w_10625 );
and ( w_10624 , w_10625 , \2124_b0 );
or ( \4384_b1 , \4378_b1 , \4383_b1 );
not ( \4383_b1 , w_10626 );
and ( \4384_b0 , \4378_b0 , w_10627 );
and ( w_10626 , w_10627 , \4383_b0 );
or ( \4385_b1 , \4374_b1 , \4383_b1 );
not ( \4383_b1 , w_10628 );
and ( \4385_b0 , \4374_b0 , w_10629 );
and ( w_10628 , w_10629 , \4383_b0 );
or ( \4387_b1 , \1778_b1 , \1280_b1 );
not ( \1280_b1 , w_10630 );
and ( \4387_b0 , \1778_b0 , w_10631 );
and ( w_10630 , w_10631 , \1280_b0 );
or ( \4388_b1 , \1770_b1 , \1278_b1 );
not ( \1278_b1 , w_10632 );
and ( \4388_b0 , \1770_b0 , w_10633 );
and ( w_10632 , w_10633 , \1278_b0 );
or ( \4389_b1 , \4387_b1 , w_10635 );
not ( w_10635 , w_10636 );
and ( \4389_b0 , \4387_b0 , w_10637 );
and ( w_10636 ,  , w_10637 );
buf ( w_10635 , \4388_b1 );
not ( w_10635 , w_10638 );
not (  , w_10639 );
and ( w_10638 , w_10639 , \4388_b0 );
or ( \4390_b1 , \4389_b1 , w_10640 );
xor ( \4390_b0 , \4389_b0 , w_10642 );
not ( w_10642 , w_10643 );
and ( w_10643 , w_10640 , w_10641 );
buf ( w_10640 , \1177_b1 );
not ( w_10640 , w_10644 );
not ( w_10641 , w_10645 );
and ( w_10644 , w_10645 , \1177_b0 );
or ( \4391_b1 , \2028_b1 , \1062_b1 );
not ( \1062_b1 , w_10646 );
and ( \4391_b0 , \2028_b0 , w_10647 );
and ( w_10646 , w_10647 , \1062_b0 );
or ( \4392_b1 , \2023_b1 , \1060_b1 );
not ( \1060_b1 , w_10648 );
and ( \4392_b0 , \2023_b0 , w_10649 );
and ( w_10648 , w_10649 , \1060_b0 );
or ( \4393_b1 , \4391_b1 , w_10651 );
not ( w_10651 , w_10652 );
and ( \4393_b0 , \4391_b0 , w_10653 );
and ( w_10652 ,  , w_10653 );
buf ( w_10651 , \4392_b1 );
not ( w_10651 , w_10654 );
not (  , w_10655 );
and ( w_10654 , w_10655 , \4392_b0 );
or ( \4394_b1 , \4393_b1 , w_10656 );
xor ( \4394_b0 , \4393_b0 , w_10658 );
not ( w_10658 , w_10659 );
and ( w_10659 , w_10656 , w_10657 );
buf ( w_10656 , \984_b1 );
not ( w_10656 , w_10660 );
not ( w_10657 , w_10661 );
and ( w_10660 , w_10661 , \984_b0 );
or ( \4395_b1 , \4390_b1 , \4394_b1 );
not ( \4394_b1 , w_10662 );
and ( \4395_b0 , \4390_b0 , w_10663 );
and ( w_10662 , w_10663 , \4394_b0 );
or ( \4396_b1 , \2305_b1 , \912_b1 );
not ( \912_b1 , w_10664 );
and ( \4396_b0 , \2305_b0 , w_10665 );
and ( w_10664 , w_10665 , \912_b0 );
or ( \4397_b1 , \2161_b1 , \910_b1 );
not ( \910_b1 , w_10666 );
and ( \4397_b0 , \2161_b0 , w_10667 );
and ( w_10666 , w_10667 , \910_b0 );
or ( \4398_b1 , \4396_b1 , w_10669 );
not ( w_10669 , w_10670 );
and ( \4398_b0 , \4396_b0 , w_10671 );
and ( w_10670 ,  , w_10671 );
buf ( w_10669 , \4397_b1 );
not ( w_10669 , w_10672 );
not (  , w_10673 );
and ( w_10672 , w_10673 , \4397_b0 );
or ( \4399_b1 , \4398_b1 , w_10674 );
xor ( \4399_b0 , \4398_b0 , w_10676 );
not ( w_10676 , w_10677 );
and ( w_10677 , w_10674 , w_10675 );
buf ( w_10674 , \818_b1 );
not ( w_10674 , w_10678 );
not ( w_10675 , w_10679 );
and ( w_10678 , w_10679 , \818_b0 );
or ( \4400_b1 , \4394_b1 , \4399_b1 );
not ( \4399_b1 , w_10680 );
and ( \4400_b0 , \4394_b0 , w_10681 );
and ( w_10680 , w_10681 , \4399_b0 );
or ( \4401_b1 , \4390_b1 , \4399_b1 );
not ( \4399_b1 , w_10682 );
and ( \4401_b0 , \4390_b0 , w_10683 );
and ( w_10682 , w_10683 , \4399_b0 );
or ( \4403_b1 , \4386_b1 , \4402_b1 );
not ( \4402_b1 , w_10684 );
and ( \4403_b0 , \4386_b0 , w_10685 );
and ( w_10684 , w_10685 , \4402_b0 );
or ( \4404_b1 , \1194_b1 , \1955_b1 );
not ( \1955_b1 , w_10686 );
and ( \4404_b0 , \1194_b0 , w_10687 );
and ( w_10686 , w_10687 , \1955_b0 );
or ( \4405_b1 , \1104_b1 , \1953_b1 );
not ( \1953_b1 , w_10688 );
and ( \4405_b0 , \1104_b0 , w_10689 );
and ( w_10688 , w_10689 , \1953_b0 );
or ( \4406_b1 , \4404_b1 , w_10691 );
not ( w_10691 , w_10692 );
and ( \4406_b0 , \4404_b0 , w_10693 );
and ( w_10692 ,  , w_10693 );
buf ( w_10691 , \4405_b1 );
not ( w_10691 , w_10694 );
not (  , w_10695 );
and ( w_10694 , w_10695 , \4405_b0 );
or ( \4407_b1 , \4406_b1 , w_10696 );
xor ( \4407_b0 , \4406_b0 , w_10698 );
not ( w_10698 , w_10699 );
and ( w_10699 , w_10696 , w_10697 );
buf ( w_10696 , \1835_b1 );
not ( w_10696 , w_10700 );
not ( w_10697 , w_10701 );
and ( w_10700 , w_10701 , \1835_b0 );
or ( \4408_b1 , \1304_b1 , \1742_b1 );
not ( \1742_b1 , w_10702 );
and ( \4408_b0 , \1304_b0 , w_10703 );
and ( w_10702 , w_10703 , \1742_b0 );
or ( \4409_b1 , \1299_b1 , \1740_b1 );
not ( \1740_b1 , w_10704 );
and ( \4409_b0 , \1299_b0 , w_10705 );
and ( w_10704 , w_10705 , \1740_b0 );
or ( \4410_b1 , \4408_b1 , w_10707 );
not ( w_10707 , w_10708 );
and ( \4410_b0 , \4408_b0 , w_10709 );
and ( w_10708 ,  , w_10709 );
buf ( w_10707 , \4409_b1 );
not ( w_10707 , w_10710 );
not (  , w_10711 );
and ( w_10710 , w_10711 , \4409_b0 );
or ( \4411_b1 , \4410_b1 , w_10712 );
xor ( \4411_b0 , \4410_b0 , w_10714 );
not ( w_10714 , w_10715 );
and ( w_10715 , w_10712 , w_10713 );
buf ( w_10712 , \1610_b1 );
not ( w_10712 , w_10716 );
not ( w_10713 , w_10717 );
and ( w_10716 , w_10717 , \1610_b0 );
or ( \4412_b1 , \4407_b1 , \4411_b1 );
not ( \4411_b1 , w_10718 );
and ( \4412_b0 , \4407_b0 , w_10719 );
and ( w_10718 , w_10719 , \4411_b0 );
or ( \4413_b1 , \1537_b1 , \1476_b1 );
not ( \1476_b1 , w_10720 );
and ( \4413_b0 , \1537_b0 , w_10721 );
and ( w_10720 , w_10721 , \1476_b0 );
or ( \4414_b1 , \1422_b1 , \1474_b1 );
not ( \1474_b1 , w_10722 );
and ( \4414_b0 , \1422_b0 , w_10723 );
and ( w_10722 , w_10723 , \1474_b0 );
or ( \4415_b1 , \4413_b1 , w_10725 );
not ( w_10725 , w_10726 );
and ( \4415_b0 , \4413_b0 , w_10727 );
and ( w_10726 ,  , w_10727 );
buf ( w_10725 , \4414_b1 );
not ( w_10725 , w_10728 );
not (  , w_10729 );
and ( w_10728 , w_10729 , \4414_b0 );
or ( \4416_b1 , \4415_b1 , w_10730 );
xor ( \4416_b0 , \4415_b0 , w_10732 );
not ( w_10732 , w_10733 );
and ( w_10733 , w_10730 , w_10731 );
buf ( w_10730 , \1363_b1 );
not ( w_10730 , w_10734 );
not ( w_10731 , w_10735 );
and ( w_10734 , w_10735 , \1363_b0 );
or ( \4417_b1 , \4411_b1 , \4416_b1 );
not ( \4416_b1 , w_10736 );
and ( \4417_b0 , \4411_b0 , w_10737 );
and ( w_10736 , w_10737 , \4416_b0 );
or ( \4418_b1 , \4407_b1 , \4416_b1 );
not ( \4416_b1 , w_10738 );
and ( \4418_b0 , \4407_b0 , w_10739 );
and ( w_10738 , w_10739 , \4416_b0 );
or ( \4420_b1 , \4402_b1 , \4419_b1 );
not ( \4419_b1 , w_10740 );
and ( \4420_b0 , \4402_b0 , w_10741 );
and ( w_10740 , w_10741 , \4419_b0 );
or ( \4421_b1 , \4386_b1 , \4419_b1 );
not ( \4419_b1 , w_10742 );
and ( \4421_b0 , \4386_b0 , w_10743 );
and ( w_10742 , w_10743 , \4419_b0 );
or ( \4423_b1 , \2850_b1 , w_10745 );
not ( w_10745 , w_10746 );
and ( \4423_b0 , \2850_b0 , w_10747 );
and ( w_10746 ,  , w_10747 );
buf ( w_10745 , \501_b1 );
not ( w_10745 , w_10748 );
not (  , w_10749 );
and ( w_10748 , w_10749 , \501_b0 );
or ( \4424_b1 , \4423_b1 , w_10750 );
xor ( \4424_b0 , \4423_b0 , w_10752 );
not ( w_10752 , w_10753 );
and ( w_10753 , w_10750 , w_10751 );
buf ( w_10750 , \455_b1 );
not ( w_10750 , w_10754 );
not ( w_10751 , w_10755 );
and ( w_10754 , w_10755 , \455_b0 );
or ( \4425_b1 , \4268_b1 , \4272_b1 );
xor ( \4425_b0 , \4268_b0 , w_10756 );
not ( w_10756 , w_10757 );
and ( w_10757 , \4272_b1 , \4272_b0 );
or ( \4426_b1 , \4425_b1 , \4277_b1 );
xor ( \4426_b0 , \4425_b0 , w_10758 );
not ( w_10758 , w_10759 );
and ( w_10759 , \4277_b1 , \4277_b0 );
or ( \4427_b1 , \4424_b1 , \4426_b1 );
not ( \4426_b1 , w_10760 );
and ( \4427_b0 , \4424_b0 , w_10761 );
and ( w_10760 , w_10761 , \4426_b0 );
or ( \4428_b1 , \4300_b1 , \4304_b1 );
xor ( \4428_b0 , \4300_b0 , w_10762 );
not ( w_10762 , w_10763 );
and ( w_10763 , \4304_b1 , \4304_b0 );
or ( \4429_b1 , \4428_b1 , \4309_b1 );
xor ( \4429_b0 , \4428_b0 , w_10764 );
not ( w_10764 , w_10765 );
and ( w_10765 , \4309_b1 , \4309_b0 );
or ( \4430_b1 , \4426_b1 , \4429_b1 );
not ( \4429_b1 , w_10766 );
and ( \4430_b0 , \4426_b0 , w_10767 );
and ( w_10766 , w_10767 , \4429_b0 );
or ( \4431_b1 , \4424_b1 , \4429_b1 );
not ( \4429_b1 , w_10768 );
and ( \4431_b0 , \4424_b0 , w_10769 );
and ( w_10768 , w_10769 , \4429_b0 );
or ( \4433_b1 , \4422_b1 , \4432_b1 );
not ( \4432_b1 , w_10770 );
and ( \4433_b0 , \4422_b0 , w_10771 );
and ( w_10770 , w_10771 , \4432_b0 );
or ( \4434_b1 , \4252_b1 , \4256_b1 );
xor ( \4434_b0 , \4252_b0 , w_10772 );
not ( w_10772 , w_10773 );
and ( w_10773 , \4256_b1 , \4256_b0 );
or ( \4435_b1 , \4434_b1 , \4261_b1 );
xor ( \4435_b0 , \4434_b0 , w_10774 );
not ( w_10774 , w_10775 );
and ( w_10775 , \4261_b1 , \4261_b0 );
or ( \4436_b1 , \4285_b1 , \4289_b1 );
xor ( \4436_b0 , \4285_b0 , w_10776 );
not ( w_10776 , w_10777 );
and ( w_10777 , \4289_b1 , \4289_b0 );
or ( \4437_b1 , \4436_b1 , \455_b1 );
xor ( \4437_b0 , \4436_b0 , w_10778 );
not ( w_10778 , w_10779 );
and ( w_10779 , \455_b1 , \455_b0 );
or ( \4438_b1 , \4435_b1 , \4437_b1 );
not ( \4437_b1 , w_10780 );
and ( \4438_b0 , \4435_b0 , w_10781 );
and ( w_10780 , w_10781 , \4437_b0 );
or ( \4439_b1 , \4432_b1 , \4438_b1 );
not ( \4438_b1 , w_10782 );
and ( \4439_b0 , \4432_b0 , w_10783 );
and ( w_10782 , w_10783 , \4438_b0 );
or ( \4440_b1 , \4422_b1 , \4438_b1 );
not ( \4438_b1 , w_10784 );
and ( \4440_b0 , \4422_b0 , w_10785 );
and ( w_10784 , w_10785 , \4438_b0 );
or ( \4442_b1 , \4264_b1 , \4280_b1 );
xor ( \4442_b0 , \4264_b0 , w_10786 );
not ( w_10786 , w_10787 );
and ( w_10787 , \4280_b1 , \4280_b0 );
or ( \4443_b1 , \4442_b1 , \4293_b1 );
xor ( \4443_b0 , \4442_b0 , w_10788 );
not ( w_10788 , w_10789 );
and ( w_10789 , \4293_b1 , \4293_b0 );
or ( \4444_b1 , \4312_b1 , \4314_b1 );
xor ( \4444_b0 , \4312_b0 , w_10790 );
not ( w_10790 , w_10791 );
and ( w_10791 , \4314_b1 , \4314_b0 );
or ( \4445_b1 , \4444_b1 , \4317_b1 );
xor ( \4445_b0 , \4444_b0 , w_10792 );
not ( w_10792 , w_10793 );
and ( w_10793 , \4317_b1 , \4317_b0 );
or ( \4446_b1 , \4443_b1 , \4445_b1 );
not ( \4445_b1 , w_10794 );
and ( \4446_b0 , \4443_b0 , w_10795 );
and ( w_10794 , w_10795 , \4445_b0 );
or ( \4447_b1 , \4323_b1 , \4325_b1 );
xor ( \4447_b0 , \4323_b0 , w_10796 );
not ( w_10796 , w_10797 );
and ( w_10797 , \4325_b1 , \4325_b0 );
or ( \4448_b1 , \4445_b1 , \4447_b1 );
not ( \4447_b1 , w_10798 );
and ( \4448_b0 , \4445_b0 , w_10799 );
and ( w_10798 , w_10799 , \4447_b0 );
or ( \4449_b1 , \4443_b1 , \4447_b1 );
not ( \4447_b1 , w_10800 );
and ( \4449_b0 , \4443_b0 , w_10801 );
and ( w_10800 , w_10801 , \4447_b0 );
or ( \4451_b1 , \4441_b1 , \4450_b1 );
not ( \4450_b1 , w_10802 );
and ( \4451_b0 , \4441_b0 , w_10803 );
and ( w_10802 , w_10803 , \4450_b0 );
or ( \4452_b1 , \4331_b1 , \4333_b1 );
xor ( \4452_b0 , \4331_b0 , w_10804 );
not ( w_10804 , w_10805 );
and ( w_10805 , \4333_b1 , \4333_b0 );
or ( \4453_b1 , \4452_b1 , \4336_b1 );
xor ( \4453_b0 , \4452_b0 , w_10806 );
not ( w_10806 , w_10807 );
and ( w_10807 , \4336_b1 , \4336_b0 );
or ( \4454_b1 , \4450_b1 , \4453_b1 );
not ( \4453_b1 , w_10808 );
and ( \4454_b0 , \4450_b0 , w_10809 );
and ( w_10808 , w_10809 , \4453_b0 );
or ( \4455_b1 , \4441_b1 , \4453_b1 );
not ( \4453_b1 , w_10810 );
and ( \4455_b0 , \4441_b0 , w_10811 );
and ( w_10810 , w_10811 , \4453_b0 );
or ( \4457_b1 , \4329_b1 , \4339_b1 );
xor ( \4457_b0 , \4329_b0 , w_10812 );
not ( w_10812 , w_10813 );
and ( w_10813 , \4339_b1 , \4339_b0 );
or ( \4458_b1 , \4457_b1 , \4342_b1 );
xor ( \4458_b0 , \4457_b0 , w_10814 );
not ( w_10814 , w_10815 );
and ( w_10815 , \4342_b1 , \4342_b0 );
or ( \4459_b1 , \4456_b1 , \4458_b1 );
not ( \4458_b1 , w_10816 );
and ( \4459_b0 , \4456_b0 , w_10817 );
and ( w_10816 , w_10817 , \4458_b0 );
or ( \4460_b1 , \4347_b1 , \4349_b1 );
xor ( \4460_b0 , \4347_b0 , w_10818 );
not ( w_10818 , w_10819 );
and ( w_10819 , \4349_b1 , \4349_b0 );
or ( \4461_b1 , \4458_b1 , \4460_b1 );
not ( \4460_b1 , w_10820 );
and ( \4461_b0 , \4458_b0 , w_10821 );
and ( w_10820 , w_10821 , \4460_b0 );
or ( \4462_b1 , \4456_b1 , \4460_b1 );
not ( \4460_b1 , w_10822 );
and ( \4462_b0 , \4456_b0 , w_10823 );
and ( w_10822 , w_10823 , \4460_b0 );
or ( \4464_b1 , \4370_b1 , \4463_b1 );
not ( \4463_b1 , w_10824 );
and ( \4464_b0 , \4370_b0 , w_10825 );
and ( w_10824 , w_10825 , \4463_b0 );
or ( \4465_b1 , \4370_b1 , \4463_b1 );
xor ( \4465_b0 , \4370_b0 , w_10826 );
not ( w_10826 , w_10827 );
and ( w_10827 , \4463_b1 , \4463_b0 );
or ( \4466_b1 , \4456_b1 , \4458_b1 );
xor ( \4466_b0 , \4456_b0 , w_10828 );
not ( w_10828 , w_10829 );
and ( w_10829 , \4458_b1 , \4458_b0 );
or ( \4467_b1 , \4466_b1 , \4460_b1 );
xor ( \4467_b0 , \4466_b0 , w_10830 );
not ( w_10830 , w_10831 );
and ( w_10831 , \4460_b1 , \4460_b0 );
or ( \4468_b1 , \2532_b1 , \912_b1 );
not ( \912_b1 , w_10832 );
and ( \4468_b0 , \2532_b0 , w_10833 );
and ( w_10832 , w_10833 , \912_b0 );
or ( \4469_b1 , \2305_b1 , \910_b1 );
not ( \910_b1 , w_10834 );
and ( \4469_b0 , \2305_b0 , w_10835 );
and ( w_10834 , w_10835 , \910_b0 );
or ( \4470_b1 , \4468_b1 , w_10837 );
not ( w_10837 , w_10838 );
and ( \4470_b0 , \4468_b0 , w_10839 );
and ( w_10838 ,  , w_10839 );
buf ( w_10837 , \4469_b1 );
not ( w_10837 , w_10840 );
not (  , w_10841 );
and ( w_10840 , w_10841 , \4469_b0 );
or ( \4471_b1 , \4470_b1 , w_10842 );
xor ( \4471_b0 , \4470_b0 , w_10844 );
not ( w_10844 , w_10845 );
and ( w_10845 , w_10842 , w_10843 );
buf ( w_10842 , \818_b1 );
not ( w_10842 , w_10846 );
not ( w_10843 , w_10847 );
and ( w_10846 , w_10847 , \818_b0 );
or ( \4472_b1 , \2763_b1 , \740_b1 );
not ( \740_b1 , w_10848 );
and ( \4472_b0 , \2763_b0 , w_10849 );
and ( w_10848 , w_10849 , \740_b0 );
or ( \4473_b1 , \2541_b1 , \738_b1 );
not ( \738_b1 , w_10850 );
and ( \4473_b0 , \2541_b0 , w_10851 );
and ( w_10850 , w_10851 , \738_b0 );
or ( \4474_b1 , \4472_b1 , w_10853 );
not ( w_10853 , w_10854 );
and ( \4474_b0 , \4472_b0 , w_10855 );
and ( w_10854 ,  , w_10855 );
buf ( w_10853 , \4473_b1 );
not ( w_10853 , w_10856 );
not (  , w_10857 );
and ( w_10856 , w_10857 , \4473_b0 );
or ( \4475_b1 , \4474_b1 , w_10858 );
xor ( \4475_b0 , \4474_b0 , w_10860 );
not ( w_10860 , w_10861 );
and ( w_10861 , w_10858 , w_10859 );
buf ( w_10858 , \668_b1 );
not ( w_10858 , w_10862 );
not ( w_10859 , w_10863 );
and ( w_10862 , w_10863 , \668_b0 );
or ( \4476_b1 , \4471_b1 , \4475_b1 );
not ( \4475_b1 , w_10864 );
and ( \4476_b0 , \4471_b0 , w_10865 );
and ( w_10864 , w_10865 , \4475_b0 );
or ( \4477_b1 , \2850_b1 , w_10867 );
not ( w_10867 , w_10868 );
and ( \4477_b0 , \2850_b0 , w_10869 );
and ( w_10868 ,  , w_10869 );
buf ( w_10867 , \602_b1 );
not ( w_10867 , w_10870 );
not (  , w_10871 );
and ( w_10870 , w_10871 , \602_b0 );
or ( \4478_b1 , \4477_b1 , w_10872 );
xor ( \4478_b0 , \4477_b0 , w_10874 );
not ( w_10874 , w_10875 );
and ( w_10875 , w_10872 , w_10873 );
buf ( w_10872 , \561_b1 );
not ( w_10872 , w_10876 );
not ( w_10873 , w_10877 );
and ( w_10876 , w_10877 , \561_b0 );
or ( \4479_b1 , \4475_b1 , \4478_b1 );
not ( \4478_b1 , w_10878 );
and ( \4479_b0 , \4475_b0 , w_10879 );
and ( w_10878 , w_10879 , \4478_b0 );
or ( \4480_b1 , \4471_b1 , \4478_b1 );
not ( \4478_b1 , w_10880 );
and ( \4480_b0 , \4471_b0 , w_10881 );
and ( w_10880 , w_10881 , \4478_b0 );
or ( \4482_b1 , \2541_b1 , \740_b1 );
not ( \740_b1 , w_10882 );
and ( \4482_b0 , \2541_b0 , w_10883 );
and ( w_10882 , w_10883 , \740_b0 );
or ( \4483_b1 , \2532_b1 , \738_b1 );
not ( \738_b1 , w_10884 );
and ( \4483_b0 , \2532_b0 , w_10885 );
and ( w_10884 , w_10885 , \738_b0 );
or ( \4484_b1 , \4482_b1 , w_10887 );
not ( w_10887 , w_10888 );
and ( \4484_b0 , \4482_b0 , w_10889 );
and ( w_10888 ,  , w_10889 );
buf ( w_10887 , \4483_b1 );
not ( w_10887 , w_10890 );
not (  , w_10891 );
and ( w_10890 , w_10891 , \4483_b0 );
or ( \4485_b1 , \4484_b1 , w_10892 );
xor ( \4485_b0 , \4484_b0 , w_10894 );
not ( w_10894 , w_10895 );
and ( w_10895 , w_10892 , w_10893 );
buf ( w_10892 , \668_b1 );
not ( w_10892 , w_10896 );
not ( w_10893 , w_10897 );
and ( w_10896 , w_10897 , \668_b0 );
or ( \4486_b1 , \4481_b1 , \4485_b1 );
not ( \4485_b1 , w_10898 );
and ( \4486_b0 , \4481_b0 , w_10899 );
and ( w_10898 , w_10899 , \4485_b0 );
or ( \4487_b1 , \2850_b1 , \604_b1 );
not ( \604_b1 , w_10900 );
and ( \4487_b0 , \2850_b0 , w_10901 );
and ( w_10900 , w_10901 , \604_b0 );
or ( \4488_b1 , \2763_b1 , \602_b1 );
not ( \602_b1 , w_10902 );
and ( \4488_b0 , \2763_b0 , w_10903 );
and ( w_10902 , w_10903 , \602_b0 );
or ( \4489_b1 , \4487_b1 , w_10905 );
not ( w_10905 , w_10906 );
and ( \4489_b0 , \4487_b0 , w_10907 );
and ( w_10906 ,  , w_10907 );
buf ( w_10905 , \4488_b1 );
not ( w_10905 , w_10908 );
not (  , w_10909 );
and ( w_10908 , w_10909 , \4488_b0 );
or ( \4490_b1 , \4489_b1 , w_10910 );
xor ( \4490_b0 , \4489_b0 , w_10912 );
not ( w_10912 , w_10913 );
and ( w_10913 , w_10910 , w_10911 );
buf ( w_10910 , \561_b1 );
not ( w_10910 , w_10914 );
not ( w_10911 , w_10915 );
and ( w_10914 , w_10915 , \561_b0 );
or ( \4491_b1 , \4485_b1 , \4490_b1 );
not ( \4490_b1 , w_10916 );
and ( \4491_b0 , \4485_b0 , w_10917 );
and ( w_10916 , w_10917 , \4490_b0 );
or ( \4492_b1 , \4481_b1 , \4490_b1 );
not ( \4490_b1 , w_10918 );
and ( \4492_b0 , \4481_b0 , w_10919 );
and ( w_10918 , w_10919 , \4490_b0 );
or ( \4494_b1 , \703_b1 , \2913_b1 );
not ( \2913_b1 , w_10920 );
and ( \4494_b0 , \703_b0 , w_10921 );
and ( w_10920 , w_10921 , \2913_b0 );
or ( \4495_b1 , \621_b1 , \2910_b1 );
not ( \2910_b1 , w_10922 );
and ( \4495_b0 , \621_b0 , w_10923 );
and ( w_10922 , w_10923 , \2910_b0 );
or ( \4496_b1 , \4494_b1 , w_10925 );
not ( w_10925 , w_10926 );
and ( \4496_b0 , \4494_b0 , w_10927 );
and ( w_10926 ,  , w_10927 );
buf ( w_10925 , \4495_b1 );
not ( w_10925 , w_10928 );
not (  , w_10929 );
and ( w_10928 , w_10929 , \4495_b0 );
or ( \4497_b1 , \4496_b1 , w_10930 );
xor ( \4497_b0 , \4496_b0 , w_10932 );
not ( w_10932 , w_10933 );
and ( w_10933 , w_10930 , w_10931 );
buf ( w_10930 , \2371_b1 );
not ( w_10930 , w_10934 );
not ( w_10931 , w_10935 );
and ( w_10934 , w_10935 , \2371_b0 );
or ( \4498_b1 , \841_b1 , \2550_b1 );
not ( \2550_b1 , w_10936 );
and ( \4498_b0 , \841_b0 , w_10937 );
and ( w_10936 , w_10937 , \2550_b0 );
or ( \4499_b1 , \777_b1 , \2548_b1 );
not ( \2548_b1 , w_10938 );
and ( \4499_b0 , \777_b0 , w_10939 );
and ( w_10938 , w_10939 , \2548_b0 );
or ( \4500_b1 , \4498_b1 , w_10941 );
not ( w_10941 , w_10942 );
and ( \4500_b0 , \4498_b0 , w_10943 );
and ( w_10942 ,  , w_10943 );
buf ( w_10941 , \4499_b1 );
not ( w_10941 , w_10944 );
not (  , w_10945 );
and ( w_10944 , w_10945 , \4499_b0 );
or ( \4501_b1 , \4500_b1 , w_10946 );
xor ( \4501_b0 , \4500_b0 , w_10948 );
not ( w_10948 , w_10949 );
and ( w_10949 , w_10946 , w_10947 );
buf ( w_10946 , \2374_b1 );
not ( w_10946 , w_10950 );
not ( w_10947 , w_10951 );
and ( w_10950 , w_10951 , \2374_b0 );
or ( \4502_b1 , \4497_b1 , \4501_b1 );
not ( \4501_b1 , w_10952 );
and ( \4502_b0 , \4497_b0 , w_10953 );
and ( w_10952 , w_10953 , \4501_b0 );
or ( \4503_b1 , \4501_b1 , \561_b1 );
not ( \561_b1 , w_10954 );
and ( \4503_b0 , \4501_b0 , w_10955 );
and ( w_10954 , w_10955 , \561_b0 );
or ( \4504_b1 , \4497_b1 , \561_b1 );
not ( \561_b1 , w_10956 );
and ( \4504_b0 , \4497_b0 , w_10957 );
and ( w_10956 , w_10957 , \561_b0 );
or ( \4506_b1 , \1104_b1 , \2261_b1 );
not ( \2261_b1 , w_10958 );
and ( \4506_b0 , \1104_b0 , w_10959 );
and ( w_10958 , w_10959 , \2261_b0 );
or ( \4507_b1 , \904_b1 , \2259_b1 );
not ( \2259_b1 , w_10960 );
and ( \4507_b0 , \904_b0 , w_10961 );
and ( w_10960 , w_10961 , \2259_b0 );
or ( \4508_b1 , \4506_b1 , w_10963 );
not ( w_10963 , w_10964 );
and ( \4508_b0 , \4506_b0 , w_10965 );
and ( w_10964 ,  , w_10965 );
buf ( w_10963 , \4507_b1 );
not ( w_10963 , w_10966 );
not (  , w_10967 );
and ( w_10966 , w_10967 , \4507_b0 );
or ( \4509_b1 , \4508_b1 , w_10968 );
xor ( \4509_b0 , \4508_b0 , w_10970 );
not ( w_10970 , w_10971 );
and ( w_10971 , w_10968 , w_10969 );
buf ( w_10968 , \2124_b1 );
not ( w_10968 , w_10972 );
not ( w_10969 , w_10973 );
and ( w_10972 , w_10973 , \2124_b0 );
or ( \4510_b1 , \1299_b1 , \1955_b1 );
not ( \1955_b1 , w_10974 );
and ( \4510_b0 , \1299_b0 , w_10975 );
and ( w_10974 , w_10975 , \1955_b0 );
or ( \4511_b1 , \1194_b1 , \1953_b1 );
not ( \1953_b1 , w_10976 );
and ( \4511_b0 , \1194_b0 , w_10977 );
and ( w_10976 , w_10977 , \1953_b0 );
or ( \4512_b1 , \4510_b1 , w_10979 );
not ( w_10979 , w_10980 );
and ( \4512_b0 , \4510_b0 , w_10981 );
and ( w_10980 ,  , w_10981 );
buf ( w_10979 , \4511_b1 );
not ( w_10979 , w_10982 );
not (  , w_10983 );
and ( w_10982 , w_10983 , \4511_b0 );
or ( \4513_b1 , \4512_b1 , w_10984 );
xor ( \4513_b0 , \4512_b0 , w_10986 );
not ( w_10986 , w_10987 );
and ( w_10987 , w_10984 , w_10985 );
buf ( w_10984 , \1835_b1 );
not ( w_10984 , w_10988 );
not ( w_10985 , w_10989 );
and ( w_10988 , w_10989 , \1835_b0 );
or ( \4514_b1 , \4509_b1 , \4513_b1 );
not ( \4513_b1 , w_10990 );
and ( \4514_b0 , \4509_b0 , w_10991 );
and ( w_10990 , w_10991 , \4513_b0 );
or ( \4515_b1 , \1422_b1 , \1742_b1 );
not ( \1742_b1 , w_10992 );
and ( \4515_b0 , \1422_b0 , w_10993 );
and ( w_10992 , w_10993 , \1742_b0 );
or ( \4516_b1 , \1304_b1 , \1740_b1 );
not ( \1740_b1 , w_10994 );
and ( \4516_b0 , \1304_b0 , w_10995 );
and ( w_10994 , w_10995 , \1740_b0 );
or ( \4517_b1 , \4515_b1 , w_10997 );
not ( w_10997 , w_10998 );
and ( \4517_b0 , \4515_b0 , w_10999 );
and ( w_10998 ,  , w_10999 );
buf ( w_10997 , \4516_b1 );
not ( w_10997 , w_11000 );
not (  , w_11001 );
and ( w_11000 , w_11001 , \4516_b0 );
or ( \4518_b1 , \4517_b1 , w_11002 );
xor ( \4518_b0 , \4517_b0 , w_11004 );
not ( w_11004 , w_11005 );
and ( w_11005 , w_11002 , w_11003 );
buf ( w_11002 , \1610_b1 );
not ( w_11002 , w_11006 );
not ( w_11003 , w_11007 );
and ( w_11006 , w_11007 , \1610_b0 );
or ( \4519_b1 , \4513_b1 , \4518_b1 );
not ( \4518_b1 , w_11008 );
and ( \4519_b0 , \4513_b0 , w_11009 );
and ( w_11008 , w_11009 , \4518_b0 );
or ( \4520_b1 , \4509_b1 , \4518_b1 );
not ( \4518_b1 , w_11010 );
and ( \4520_b0 , \4509_b0 , w_11011 );
and ( w_11010 , w_11011 , \4518_b0 );
or ( \4522_b1 , \4505_b1 , \4521_b1 );
not ( \4521_b1 , w_11012 );
and ( \4522_b0 , \4505_b0 , w_11013 );
and ( w_11012 , w_11013 , \4521_b0 );
or ( \4523_b1 , \1770_b1 , \1476_b1 );
not ( \1476_b1 , w_11014 );
and ( \4523_b0 , \1770_b0 , w_11015 );
and ( w_11014 , w_11015 , \1476_b0 );
or ( \4524_b1 , \1537_b1 , \1474_b1 );
not ( \1474_b1 , w_11016 );
and ( \4524_b0 , \1537_b0 , w_11017 );
and ( w_11016 , w_11017 , \1474_b0 );
or ( \4525_b1 , \4523_b1 , w_11019 );
not ( w_11019 , w_11020 );
and ( \4525_b0 , \4523_b0 , w_11021 );
and ( w_11020 ,  , w_11021 );
buf ( w_11019 , \4524_b1 );
not ( w_11019 , w_11022 );
not (  , w_11023 );
and ( w_11022 , w_11023 , \4524_b0 );
or ( \4526_b1 , \4525_b1 , w_11024 );
xor ( \4526_b0 , \4525_b0 , w_11026 );
not ( w_11026 , w_11027 );
and ( w_11027 , w_11024 , w_11025 );
buf ( w_11024 , \1363_b1 );
not ( w_11024 , w_11028 );
not ( w_11025 , w_11029 );
and ( w_11028 , w_11029 , \1363_b0 );
or ( \4527_b1 , \2023_b1 , \1280_b1 );
not ( \1280_b1 , w_11030 );
and ( \4527_b0 , \2023_b0 , w_11031 );
and ( w_11030 , w_11031 , \1280_b0 );
or ( \4528_b1 , \1778_b1 , \1278_b1 );
not ( \1278_b1 , w_11032 );
and ( \4528_b0 , \1778_b0 , w_11033 );
and ( w_11032 , w_11033 , \1278_b0 );
or ( \4529_b1 , \4527_b1 , w_11035 );
not ( w_11035 , w_11036 );
and ( \4529_b0 , \4527_b0 , w_11037 );
and ( w_11036 ,  , w_11037 );
buf ( w_11035 , \4528_b1 );
not ( w_11035 , w_11038 );
not (  , w_11039 );
and ( w_11038 , w_11039 , \4528_b0 );
or ( \4530_b1 , \4529_b1 , w_11040 );
xor ( \4530_b0 , \4529_b0 , w_11042 );
not ( w_11042 , w_11043 );
and ( w_11043 , w_11040 , w_11041 );
buf ( w_11040 , \1177_b1 );
not ( w_11040 , w_11044 );
not ( w_11041 , w_11045 );
and ( w_11044 , w_11045 , \1177_b0 );
or ( \4531_b1 , \4526_b1 , \4530_b1 );
not ( \4530_b1 , w_11046 );
and ( \4531_b0 , \4526_b0 , w_11047 );
and ( w_11046 , w_11047 , \4530_b0 );
or ( \4532_b1 , \2161_b1 , \1062_b1 );
not ( \1062_b1 , w_11048 );
and ( \4532_b0 , \2161_b0 , w_11049 );
and ( w_11048 , w_11049 , \1062_b0 );
or ( \4533_b1 , \2028_b1 , \1060_b1 );
not ( \1060_b1 , w_11050 );
and ( \4533_b0 , \2028_b0 , w_11051 );
and ( w_11050 , w_11051 , \1060_b0 );
or ( \4534_b1 , \4532_b1 , w_11053 );
not ( w_11053 , w_11054 );
and ( \4534_b0 , \4532_b0 , w_11055 );
and ( w_11054 ,  , w_11055 );
buf ( w_11053 , \4533_b1 );
not ( w_11053 , w_11056 );
not (  , w_11057 );
and ( w_11056 , w_11057 , \4533_b0 );
or ( \4535_b1 , \4534_b1 , w_11058 );
xor ( \4535_b0 , \4534_b0 , w_11060 );
not ( w_11060 , w_11061 );
and ( w_11061 , w_11058 , w_11059 );
buf ( w_11058 , \984_b1 );
not ( w_11058 , w_11062 );
not ( w_11059 , w_11063 );
and ( w_11062 , w_11063 , \984_b0 );
or ( \4536_b1 , \4530_b1 , \4535_b1 );
not ( \4535_b1 , w_11064 );
and ( \4536_b0 , \4530_b0 , w_11065 );
and ( w_11064 , w_11065 , \4535_b0 );
or ( \4537_b1 , \4526_b1 , \4535_b1 );
not ( \4535_b1 , w_11066 );
and ( \4537_b0 , \4526_b0 , w_11067 );
and ( w_11066 , w_11067 , \4535_b0 );
or ( \4539_b1 , \4521_b1 , \4538_b1 );
not ( \4538_b1 , w_11068 );
and ( \4539_b0 , \4521_b0 , w_11069 );
and ( w_11068 , w_11069 , \4538_b0 );
or ( \4540_b1 , \4505_b1 , \4538_b1 );
not ( \4538_b1 , w_11070 );
and ( \4540_b0 , \4505_b0 , w_11071 );
and ( w_11070 , w_11071 , \4538_b0 );
or ( \4542_b1 , \4493_b1 , \4541_b1 );
not ( \4541_b1 , w_11072 );
and ( \4542_b0 , \4493_b0 , w_11073 );
and ( w_11072 , w_11073 , \4541_b0 );
or ( \4543_b1 , \4374_b1 , \4378_b1 );
xor ( \4543_b0 , \4374_b0 , w_11074 );
not ( w_11074 , w_11075 );
and ( w_11075 , \4378_b1 , \4378_b0 );
or ( \4544_b1 , \4543_b1 , \4383_b1 );
xor ( \4544_b0 , \4543_b0 , w_11076 );
not ( w_11076 , w_11077 );
and ( w_11077 , \4383_b1 , \4383_b0 );
or ( \4545_b1 , \4390_b1 , \4394_b1 );
xor ( \4545_b0 , \4390_b0 , w_11078 );
not ( w_11078 , w_11079 );
and ( w_11079 , \4394_b1 , \4394_b0 );
or ( \4546_b1 , \4545_b1 , \4399_b1 );
xor ( \4546_b0 , \4545_b0 , w_11080 );
not ( w_11080 , w_11081 );
and ( w_11081 , \4399_b1 , \4399_b0 );
or ( \4547_b1 , \4544_b1 , \4546_b1 );
not ( \4546_b1 , w_11082 );
and ( \4547_b0 , \4544_b0 , w_11083 );
and ( w_11082 , w_11083 , \4546_b0 );
or ( \4548_b1 , \4407_b1 , \4411_b1 );
xor ( \4548_b0 , \4407_b0 , w_11084 );
not ( w_11084 , w_11085 );
and ( w_11085 , \4411_b1 , \4411_b0 );
or ( \4549_b1 , \4548_b1 , \4416_b1 );
xor ( \4549_b0 , \4548_b0 , w_11086 );
not ( w_11086 , w_11087 );
and ( w_11087 , \4416_b1 , \4416_b0 );
or ( \4550_b1 , \4546_b1 , \4549_b1 );
not ( \4549_b1 , w_11088 );
and ( \4550_b0 , \4546_b0 , w_11089 );
and ( w_11088 , w_11089 , \4549_b0 );
or ( \4551_b1 , \4544_b1 , \4549_b1 );
not ( \4549_b1 , w_11090 );
and ( \4551_b0 , \4544_b0 , w_11091 );
and ( w_11090 , w_11091 , \4549_b0 );
or ( \4553_b1 , \4541_b1 , \4552_b1 );
not ( \4552_b1 , w_11092 );
and ( \4553_b0 , \4541_b0 , w_11093 );
and ( w_11092 , w_11093 , \4552_b0 );
or ( \4554_b1 , \4493_b1 , \4552_b1 );
not ( \4552_b1 , w_11094 );
and ( \4554_b0 , \4493_b0 , w_11095 );
and ( w_11094 , w_11095 , \4552_b0 );
or ( \4556_b1 , \4386_b1 , \4402_b1 );
xor ( \4556_b0 , \4386_b0 , w_11096 );
not ( w_11096 , w_11097 );
and ( w_11097 , \4402_b1 , \4402_b0 );
or ( \4557_b1 , \4556_b1 , \4419_b1 );
xor ( \4557_b0 , \4556_b0 , w_11098 );
not ( w_11098 , w_11099 );
and ( w_11099 , \4419_b1 , \4419_b0 );
or ( \4558_b1 , \4424_b1 , \4426_b1 );
xor ( \4558_b0 , \4424_b0 , w_11100 );
not ( w_11100 , w_11101 );
and ( w_11101 , \4426_b1 , \4426_b0 );
or ( \4559_b1 , \4558_b1 , \4429_b1 );
xor ( \4559_b0 , \4558_b0 , w_11102 );
not ( w_11102 , w_11103 );
and ( w_11103 , \4429_b1 , \4429_b0 );
or ( \4560_b1 , \4557_b1 , \4559_b1 );
not ( \4559_b1 , w_11104 );
and ( \4560_b0 , \4557_b0 , w_11105 );
and ( w_11104 , w_11105 , \4559_b0 );
or ( \4561_b1 , \4435_b1 , \4437_b1 );
xor ( \4561_b0 , \4435_b0 , w_11106 );
not ( w_11106 , w_11107 );
and ( w_11107 , \4437_b1 , \4437_b0 );
or ( \4562_b1 , \4559_b1 , \4561_b1 );
not ( \4561_b1 , w_11108 );
and ( \4562_b0 , \4559_b0 , w_11109 );
and ( w_11108 , w_11109 , \4561_b0 );
or ( \4563_b1 , \4557_b1 , \4561_b1 );
not ( \4561_b1 , w_11110 );
and ( \4563_b0 , \4557_b0 , w_11111 );
and ( w_11110 , w_11111 , \4561_b0 );
or ( \4565_b1 , \4555_b1 , \4564_b1 );
not ( \4564_b1 , w_11112 );
and ( \4565_b0 , \4555_b0 , w_11113 );
and ( w_11112 , w_11113 , \4564_b0 );
or ( \4566_b1 , \4443_b1 , \4445_b1 );
xor ( \4566_b0 , \4443_b0 , w_11114 );
not ( w_11114 , w_11115 );
and ( w_11115 , \4445_b1 , \4445_b0 );
or ( \4567_b1 , \4566_b1 , \4447_b1 );
xor ( \4567_b0 , \4566_b0 , w_11116 );
not ( w_11116 , w_11117 );
and ( w_11117 , \4447_b1 , \4447_b0 );
or ( \4568_b1 , \4564_b1 , \4567_b1 );
not ( \4567_b1 , w_11118 );
and ( \4568_b0 , \4564_b0 , w_11119 );
and ( w_11118 , w_11119 , \4567_b0 );
or ( \4569_b1 , \4555_b1 , \4567_b1 );
not ( \4567_b1 , w_11120 );
and ( \4569_b0 , \4555_b0 , w_11121 );
and ( w_11120 , w_11121 , \4567_b0 );
or ( \4571_b1 , \4296_b1 , \4320_b1 );
xor ( \4571_b0 , \4296_b0 , w_11122 );
not ( w_11122 , w_11123 );
and ( w_11123 , \4320_b1 , \4320_b0 );
or ( \4572_b1 , \4571_b1 , \4326_b1 );
xor ( \4572_b0 , \4571_b0 , w_11124 );
not ( w_11124 , w_11125 );
and ( w_11125 , \4326_b1 , \4326_b0 );
or ( \4573_b1 , \4570_b1 , \4572_b1 );
not ( \4572_b1 , w_11126 );
and ( \4573_b0 , \4570_b0 , w_11127 );
and ( w_11126 , w_11127 , \4572_b0 );
or ( \4574_b1 , \4441_b1 , \4450_b1 );
xor ( \4574_b0 , \4441_b0 , w_11128 );
not ( w_11128 , w_11129 );
and ( w_11129 , \4450_b1 , \4450_b0 );
or ( \4575_b1 , \4574_b1 , \4453_b1 );
xor ( \4575_b0 , \4574_b0 , w_11130 );
not ( w_11130 , w_11131 );
and ( w_11131 , \4453_b1 , \4453_b0 );
or ( \4576_b1 , \4572_b1 , \4575_b1 );
not ( \4575_b1 , w_11132 );
and ( \4576_b0 , \4572_b0 , w_11133 );
and ( w_11132 , w_11133 , \4575_b0 );
or ( \4577_b1 , \4570_b1 , \4575_b1 );
not ( \4575_b1 , w_11134 );
and ( \4577_b0 , \4570_b0 , w_11135 );
and ( w_11134 , w_11135 , \4575_b0 );
or ( \4579_b1 , \4467_b1 , \4578_b1 );
not ( \4578_b1 , w_11136 );
and ( \4579_b0 , \4467_b0 , w_11137 );
and ( w_11136 , w_11137 , \4578_b0 );
or ( \4580_b1 , \4467_b1 , \4578_b1 );
xor ( \4580_b0 , \4467_b0 , w_11138 );
not ( w_11138 , w_11139 );
and ( w_11139 , \4578_b1 , \4578_b0 );
or ( \4581_b1 , \4570_b1 , \4572_b1 );
xor ( \4581_b0 , \4570_b0 , w_11140 );
not ( w_11140 , w_11141 );
and ( w_11141 , \4572_b1 , \4572_b0 );
or ( \4582_b1 , \4581_b1 , \4575_b1 );
xor ( \4582_b0 , \4581_b0 , w_11142 );
not ( w_11142 , w_11143 );
and ( w_11143 , \4575_b1 , \4575_b0 );
or ( \4583_b1 , \2028_b1 , \1280_b1 );
not ( \1280_b1 , w_11144 );
and ( \4583_b0 , \2028_b0 , w_11145 );
and ( w_11144 , w_11145 , \1280_b0 );
or ( \4584_b1 , \2023_b1 , \1278_b1 );
not ( \1278_b1 , w_11146 );
and ( \4584_b0 , \2023_b0 , w_11147 );
and ( w_11146 , w_11147 , \1278_b0 );
or ( \4585_b1 , \4583_b1 , w_11149 );
not ( w_11149 , w_11150 );
and ( \4585_b0 , \4583_b0 , w_11151 );
and ( w_11150 ,  , w_11151 );
buf ( w_11149 , \4584_b1 );
not ( w_11149 , w_11152 );
not (  , w_11153 );
and ( w_11152 , w_11153 , \4584_b0 );
or ( \4586_b1 , \4585_b1 , w_11154 );
xor ( \4586_b0 , \4585_b0 , w_11156 );
not ( w_11156 , w_11157 );
and ( w_11157 , w_11154 , w_11155 );
buf ( w_11154 , \1177_b1 );
not ( w_11154 , w_11158 );
not ( w_11155 , w_11159 );
and ( w_11158 , w_11159 , \1177_b0 );
or ( \4587_b1 , \2305_b1 , \1062_b1 );
not ( \1062_b1 , w_11160 );
and ( \4587_b0 , \2305_b0 , w_11161 );
and ( w_11160 , w_11161 , \1062_b0 );
or ( \4588_b1 , \2161_b1 , \1060_b1 );
not ( \1060_b1 , w_11162 );
and ( \4588_b0 , \2161_b0 , w_11163 );
and ( w_11162 , w_11163 , \1060_b0 );
or ( \4589_b1 , \4587_b1 , w_11165 );
not ( w_11165 , w_11166 );
and ( \4589_b0 , \4587_b0 , w_11167 );
and ( w_11166 ,  , w_11167 );
buf ( w_11165 , \4588_b1 );
not ( w_11165 , w_11168 );
not (  , w_11169 );
and ( w_11168 , w_11169 , \4588_b0 );
or ( \4590_b1 , \4589_b1 , w_11170 );
xor ( \4590_b0 , \4589_b0 , w_11172 );
not ( w_11172 , w_11173 );
and ( w_11173 , w_11170 , w_11171 );
buf ( w_11170 , \984_b1 );
not ( w_11170 , w_11174 );
not ( w_11171 , w_11175 );
and ( w_11174 , w_11175 , \984_b0 );
or ( \4591_b1 , \4586_b1 , \4590_b1 );
not ( \4590_b1 , w_11176 );
and ( \4591_b0 , \4586_b0 , w_11177 );
and ( w_11176 , w_11177 , \4590_b0 );
or ( \4592_b1 , \2541_b1 , \912_b1 );
not ( \912_b1 , w_11178 );
and ( \4592_b0 , \2541_b0 , w_11179 );
and ( w_11178 , w_11179 , \912_b0 );
or ( \4593_b1 , \2532_b1 , \910_b1 );
not ( \910_b1 , w_11180 );
and ( \4593_b0 , \2532_b0 , w_11181 );
and ( w_11180 , w_11181 , \910_b0 );
or ( \4594_b1 , \4592_b1 , w_11183 );
not ( w_11183 , w_11184 );
and ( \4594_b0 , \4592_b0 , w_11185 );
and ( w_11184 ,  , w_11185 );
buf ( w_11183 , \4593_b1 );
not ( w_11183 , w_11186 );
not (  , w_11187 );
and ( w_11186 , w_11187 , \4593_b0 );
or ( \4595_b1 , \4594_b1 , w_11188 );
xor ( \4595_b0 , \4594_b0 , w_11190 );
not ( w_11190 , w_11191 );
and ( w_11191 , w_11188 , w_11189 );
buf ( w_11188 , \818_b1 );
not ( w_11188 , w_11192 );
not ( w_11189 , w_11193 );
and ( w_11192 , w_11193 , \818_b0 );
or ( \4596_b1 , \4590_b1 , \4595_b1 );
not ( \4595_b1 , w_11194 );
and ( \4596_b0 , \4590_b0 , w_11195 );
and ( w_11194 , w_11195 , \4595_b0 );
or ( \4597_b1 , \4586_b1 , \4595_b1 );
not ( \4595_b1 , w_11196 );
and ( \4597_b0 , \4586_b0 , w_11197 );
and ( w_11196 , w_11197 , \4595_b0 );
or ( \4599_b1 , \777_b1 , \2913_b1 );
not ( \2913_b1 , w_11198 );
and ( \4599_b0 , \777_b0 , w_11199 );
and ( w_11198 , w_11199 , \2913_b0 );
or ( \4600_b1 , \703_b1 , \2910_b1 );
not ( \2910_b1 , w_11200 );
and ( \4600_b0 , \703_b0 , w_11201 );
and ( w_11200 , w_11201 , \2910_b0 );
or ( \4601_b1 , \4599_b1 , w_11203 );
not ( w_11203 , w_11204 );
and ( \4601_b0 , \4599_b0 , w_11205 );
and ( w_11204 ,  , w_11205 );
buf ( w_11203 , \4600_b1 );
not ( w_11203 , w_11206 );
not (  , w_11207 );
and ( w_11206 , w_11207 , \4600_b0 );
or ( \4602_b1 , \4601_b1 , w_11208 );
xor ( \4602_b0 , \4601_b0 , w_11210 );
not ( w_11210 , w_11211 );
and ( w_11211 , w_11208 , w_11209 );
buf ( w_11208 , \2371_b1 );
not ( w_11208 , w_11212 );
not ( w_11209 , w_11213 );
and ( w_11212 , w_11213 , \2371_b0 );
or ( \4603_b1 , \904_b1 , \2550_b1 );
not ( \2550_b1 , w_11214 );
and ( \4603_b0 , \904_b0 , w_11215 );
and ( w_11214 , w_11215 , \2550_b0 );
or ( \4604_b1 , \841_b1 , \2548_b1 );
not ( \2548_b1 , w_11216 );
and ( \4604_b0 , \841_b0 , w_11217 );
and ( w_11216 , w_11217 , \2548_b0 );
or ( \4605_b1 , \4603_b1 , w_11219 );
not ( w_11219 , w_11220 );
and ( \4605_b0 , \4603_b0 , w_11221 );
and ( w_11220 ,  , w_11221 );
buf ( w_11219 , \4604_b1 );
not ( w_11219 , w_11222 );
not (  , w_11223 );
and ( w_11222 , w_11223 , \4604_b0 );
or ( \4606_b1 , \4605_b1 , w_11224 );
xor ( \4606_b0 , \4605_b0 , w_11226 );
not ( w_11226 , w_11227 );
and ( w_11227 , w_11224 , w_11225 );
buf ( w_11224 , \2374_b1 );
not ( w_11224 , w_11228 );
not ( w_11225 , w_11229 );
and ( w_11228 , w_11229 , \2374_b0 );
or ( \4607_b1 , \4602_b1 , \4606_b1 );
not ( \4606_b1 , w_11230 );
and ( \4607_b0 , \4602_b0 , w_11231 );
and ( w_11230 , w_11231 , \4606_b0 );
or ( \4608_b1 , \1194_b1 , \2261_b1 );
not ( \2261_b1 , w_11232 );
and ( \4608_b0 , \1194_b0 , w_11233 );
and ( w_11232 , w_11233 , \2261_b0 );
or ( \4609_b1 , \1104_b1 , \2259_b1 );
not ( \2259_b1 , w_11234 );
and ( \4609_b0 , \1104_b0 , w_11235 );
and ( w_11234 , w_11235 , \2259_b0 );
or ( \4610_b1 , \4608_b1 , w_11237 );
not ( w_11237 , w_11238 );
and ( \4610_b0 , \4608_b0 , w_11239 );
and ( w_11238 ,  , w_11239 );
buf ( w_11237 , \4609_b1 );
not ( w_11237 , w_11240 );
not (  , w_11241 );
and ( w_11240 , w_11241 , \4609_b0 );
or ( \4611_b1 , \4610_b1 , w_11242 );
xor ( \4611_b0 , \4610_b0 , w_11244 );
not ( w_11244 , w_11245 );
and ( w_11245 , w_11242 , w_11243 );
buf ( w_11242 , \2124_b1 );
not ( w_11242 , w_11246 );
not ( w_11243 , w_11247 );
and ( w_11246 , w_11247 , \2124_b0 );
or ( \4612_b1 , \4606_b1 , \4611_b1 );
not ( \4611_b1 , w_11248 );
and ( \4612_b0 , \4606_b0 , w_11249 );
and ( w_11248 , w_11249 , \4611_b0 );
or ( \4613_b1 , \4602_b1 , \4611_b1 );
not ( \4611_b1 , w_11250 );
and ( \4613_b0 , \4602_b0 , w_11251 );
and ( w_11250 , w_11251 , \4611_b0 );
or ( \4615_b1 , \4598_b1 , \4614_b1 );
not ( \4614_b1 , w_11252 );
and ( \4615_b0 , \4598_b0 , w_11253 );
and ( w_11252 , w_11253 , \4614_b0 );
or ( \4616_b1 , \1304_b1 , \1955_b1 );
not ( \1955_b1 , w_11254 );
and ( \4616_b0 , \1304_b0 , w_11255 );
and ( w_11254 , w_11255 , \1955_b0 );
or ( \4617_b1 , \1299_b1 , \1953_b1 );
not ( \1953_b1 , w_11256 );
and ( \4617_b0 , \1299_b0 , w_11257 );
and ( w_11256 , w_11257 , \1953_b0 );
or ( \4618_b1 , \4616_b1 , w_11259 );
not ( w_11259 , w_11260 );
and ( \4618_b0 , \4616_b0 , w_11261 );
and ( w_11260 ,  , w_11261 );
buf ( w_11259 , \4617_b1 );
not ( w_11259 , w_11262 );
not (  , w_11263 );
and ( w_11262 , w_11263 , \4617_b0 );
or ( \4619_b1 , \4618_b1 , w_11264 );
xor ( \4619_b0 , \4618_b0 , w_11266 );
not ( w_11266 , w_11267 );
and ( w_11267 , w_11264 , w_11265 );
buf ( w_11264 , \1835_b1 );
not ( w_11264 , w_11268 );
not ( w_11265 , w_11269 );
and ( w_11268 , w_11269 , \1835_b0 );
or ( \4620_b1 , \1537_b1 , \1742_b1 );
not ( \1742_b1 , w_11270 );
and ( \4620_b0 , \1537_b0 , w_11271 );
and ( w_11270 , w_11271 , \1742_b0 );
or ( \4621_b1 , \1422_b1 , \1740_b1 );
not ( \1740_b1 , w_11272 );
and ( \4621_b0 , \1422_b0 , w_11273 );
and ( w_11272 , w_11273 , \1740_b0 );
or ( \4622_b1 , \4620_b1 , w_11275 );
not ( w_11275 , w_11276 );
and ( \4622_b0 , \4620_b0 , w_11277 );
and ( w_11276 ,  , w_11277 );
buf ( w_11275 , \4621_b1 );
not ( w_11275 , w_11278 );
not (  , w_11279 );
and ( w_11278 , w_11279 , \4621_b0 );
or ( \4623_b1 , \4622_b1 , w_11280 );
xor ( \4623_b0 , \4622_b0 , w_11282 );
not ( w_11282 , w_11283 );
and ( w_11283 , w_11280 , w_11281 );
buf ( w_11280 , \1610_b1 );
not ( w_11280 , w_11284 );
not ( w_11281 , w_11285 );
and ( w_11284 , w_11285 , \1610_b0 );
or ( \4624_b1 , \4619_b1 , \4623_b1 );
not ( \4623_b1 , w_11286 );
and ( \4624_b0 , \4619_b0 , w_11287 );
and ( w_11286 , w_11287 , \4623_b0 );
or ( \4625_b1 , \1778_b1 , \1476_b1 );
not ( \1476_b1 , w_11288 );
and ( \4625_b0 , \1778_b0 , w_11289 );
and ( w_11288 , w_11289 , \1476_b0 );
or ( \4626_b1 , \1770_b1 , \1474_b1 );
not ( \1474_b1 , w_11290 );
and ( \4626_b0 , \1770_b0 , w_11291 );
and ( w_11290 , w_11291 , \1474_b0 );
or ( \4627_b1 , \4625_b1 , w_11293 );
not ( w_11293 , w_11294 );
and ( \4627_b0 , \4625_b0 , w_11295 );
and ( w_11294 ,  , w_11295 );
buf ( w_11293 , \4626_b1 );
not ( w_11293 , w_11296 );
not (  , w_11297 );
and ( w_11296 , w_11297 , \4626_b0 );
or ( \4628_b1 , \4627_b1 , w_11298 );
xor ( \4628_b0 , \4627_b0 , w_11300 );
not ( w_11300 , w_11301 );
and ( w_11301 , w_11298 , w_11299 );
buf ( w_11298 , \1363_b1 );
not ( w_11298 , w_11302 );
not ( w_11299 , w_11303 );
and ( w_11302 , w_11303 , \1363_b0 );
or ( \4629_b1 , \4623_b1 , \4628_b1 );
not ( \4628_b1 , w_11304 );
and ( \4629_b0 , \4623_b0 , w_11305 );
and ( w_11304 , w_11305 , \4628_b0 );
or ( \4630_b1 , \4619_b1 , \4628_b1 );
not ( \4628_b1 , w_11306 );
and ( \4630_b0 , \4619_b0 , w_11307 );
and ( w_11306 , w_11307 , \4628_b0 );
or ( \4632_b1 , \4614_b1 , \4631_b1 );
not ( \4631_b1 , w_11308 );
and ( \4632_b0 , \4614_b0 , w_11309 );
and ( w_11308 , w_11309 , \4631_b0 );
or ( \4633_b1 , \4598_b1 , \4631_b1 );
not ( \4631_b1 , w_11310 );
and ( \4633_b0 , \4598_b0 , w_11311 );
and ( w_11310 , w_11311 , \4631_b0 );
or ( \4635_b1 , \4509_b1 , \4513_b1 );
xor ( \4635_b0 , \4509_b0 , w_11312 );
not ( w_11312 , w_11313 );
and ( w_11313 , \4513_b1 , \4513_b0 );
or ( \4636_b1 , \4635_b1 , \4518_b1 );
xor ( \4636_b0 , \4635_b0 , w_11314 );
not ( w_11314 , w_11315 );
and ( w_11315 , \4518_b1 , \4518_b0 );
or ( \4637_b1 , \4471_b1 , \4475_b1 );
xor ( \4637_b0 , \4471_b0 , w_11316 );
not ( w_11316 , w_11317 );
and ( w_11317 , \4475_b1 , \4475_b0 );
or ( \4638_b1 , \4637_b1 , \4478_b1 );
xor ( \4638_b0 , \4637_b0 , w_11318 );
not ( w_11318 , w_11319 );
and ( w_11319 , \4478_b1 , \4478_b0 );
or ( \4639_b1 , \4636_b1 , \4638_b1 );
not ( \4638_b1 , w_11320 );
and ( \4639_b0 , \4636_b0 , w_11321 );
and ( w_11320 , w_11321 , \4638_b0 );
or ( \4640_b1 , \4526_b1 , \4530_b1 );
xor ( \4640_b0 , \4526_b0 , w_11322 );
not ( w_11322 , w_11323 );
and ( w_11323 , \4530_b1 , \4530_b0 );
or ( \4641_b1 , \4640_b1 , \4535_b1 );
xor ( \4641_b0 , \4640_b0 , w_11324 );
not ( w_11324 , w_11325 );
and ( w_11325 , \4535_b1 , \4535_b0 );
or ( \4642_b1 , \4638_b1 , \4641_b1 );
not ( \4641_b1 , w_11326 );
and ( \4642_b0 , \4638_b0 , w_11327 );
and ( w_11326 , w_11327 , \4641_b0 );
or ( \4643_b1 , \4636_b1 , \4641_b1 );
not ( \4641_b1 , w_11328 );
and ( \4643_b0 , \4636_b0 , w_11329 );
and ( w_11328 , w_11329 , \4641_b0 );
or ( \4645_b1 , \4634_b1 , \4644_b1 );
not ( \4644_b1 , w_11330 );
and ( \4645_b0 , \4634_b0 , w_11331 );
and ( w_11330 , w_11331 , \4644_b0 );
or ( \4646_b1 , \4544_b1 , \4546_b1 );
xor ( \4646_b0 , \4544_b0 , w_11332 );
not ( w_11332 , w_11333 );
and ( w_11333 , \4546_b1 , \4546_b0 );
or ( \4647_b1 , \4646_b1 , \4549_b1 );
xor ( \4647_b0 , \4646_b0 , w_11334 );
not ( w_11334 , w_11335 );
and ( w_11335 , \4549_b1 , \4549_b0 );
or ( \4648_b1 , \4644_b1 , \4647_b1 );
not ( \4647_b1 , w_11336 );
and ( \4648_b0 , \4644_b0 , w_11337 );
and ( w_11336 , w_11337 , \4647_b0 );
or ( \4649_b1 , \4634_b1 , \4647_b1 );
not ( \4647_b1 , w_11338 );
and ( \4649_b0 , \4634_b0 , w_11339 );
and ( w_11338 , w_11339 , \4647_b0 );
or ( \4651_b1 , \4493_b1 , \4541_b1 );
xor ( \4651_b0 , \4493_b0 , w_11340 );
not ( w_11340 , w_11341 );
and ( w_11341 , \4541_b1 , \4541_b0 );
or ( \4652_b1 , \4651_b1 , \4552_b1 );
xor ( \4652_b0 , \4651_b0 , w_11342 );
not ( w_11342 , w_11343 );
and ( w_11343 , \4552_b1 , \4552_b0 );
or ( \4653_b1 , \4650_b1 , \4652_b1 );
not ( \4652_b1 , w_11344 );
and ( \4653_b0 , \4650_b0 , w_11345 );
and ( w_11344 , w_11345 , \4652_b0 );
or ( \4654_b1 , \4557_b1 , \4559_b1 );
xor ( \4654_b0 , \4557_b0 , w_11346 );
not ( w_11346 , w_11347 );
and ( w_11347 , \4559_b1 , \4559_b0 );
or ( \4655_b1 , \4654_b1 , \4561_b1 );
xor ( \4655_b0 , \4654_b0 , w_11348 );
not ( w_11348 , w_11349 );
and ( w_11349 , \4561_b1 , \4561_b0 );
or ( \4656_b1 , \4652_b1 , \4655_b1 );
not ( \4655_b1 , w_11350 );
and ( \4656_b0 , \4652_b0 , w_11351 );
and ( w_11350 , w_11351 , \4655_b0 );
or ( \4657_b1 , \4650_b1 , \4655_b1 );
not ( \4655_b1 , w_11352 );
and ( \4657_b0 , \4650_b0 , w_11353 );
and ( w_11352 , w_11353 , \4655_b0 );
or ( \4659_b1 , \4422_b1 , \4432_b1 );
xor ( \4659_b0 , \4422_b0 , w_11354 );
not ( w_11354 , w_11355 );
and ( w_11355 , \4432_b1 , \4432_b0 );
or ( \4660_b1 , \4659_b1 , \4438_b1 );
xor ( \4660_b0 , \4659_b0 , w_11356 );
not ( w_11356 , w_11357 );
and ( w_11357 , \4438_b1 , \4438_b0 );
or ( \4661_b1 , \4658_b1 , \4660_b1 );
not ( \4660_b1 , w_11358 );
and ( \4661_b0 , \4658_b0 , w_11359 );
and ( w_11358 , w_11359 , \4660_b0 );
or ( \4662_b1 , \4555_b1 , \4564_b1 );
xor ( \4662_b0 , \4555_b0 , w_11360 );
not ( w_11360 , w_11361 );
and ( w_11361 , \4564_b1 , \4564_b0 );
or ( \4663_b1 , \4662_b1 , \4567_b1 );
xor ( \4663_b0 , \4662_b0 , w_11362 );
not ( w_11362 , w_11363 );
and ( w_11363 , \4567_b1 , \4567_b0 );
or ( \4664_b1 , \4660_b1 , \4663_b1 );
not ( \4663_b1 , w_11364 );
and ( \4664_b0 , \4660_b0 , w_11365 );
and ( w_11364 , w_11365 , \4663_b0 );
or ( \4665_b1 , \4658_b1 , \4663_b1 );
not ( \4663_b1 , w_11366 );
and ( \4665_b0 , \4658_b0 , w_11367 );
and ( w_11366 , w_11367 , \4663_b0 );
or ( \4667_b1 , \4582_b1 , \4666_b1 );
not ( \4666_b1 , w_11368 );
and ( \4667_b0 , \4582_b0 , w_11369 );
and ( w_11368 , w_11369 , \4666_b0 );
or ( \4668_b1 , \4582_b1 , \4666_b1 );
xor ( \4668_b0 , \4582_b0 , w_11370 );
not ( w_11370 , w_11371 );
and ( w_11371 , \4666_b1 , \4666_b0 );
or ( \4669_b1 , \4658_b1 , \4660_b1 );
xor ( \4669_b0 , \4658_b0 , w_11372 );
not ( w_11372 , w_11373 );
and ( w_11373 , \4660_b1 , \4660_b0 );
or ( \4670_b1 , \4669_b1 , \4663_b1 );
xor ( \4670_b0 , \4669_b0 , w_11374 );
not ( w_11374 , w_11375 );
and ( w_11375 , \4663_b1 , \4663_b0 );
or ( \4671_b1 , \841_b1 , \2913_b1 );
not ( \2913_b1 , w_11376 );
and ( \4671_b0 , \841_b0 , w_11377 );
and ( w_11376 , w_11377 , \2913_b0 );
or ( \4672_b1 , \777_b1 , \2910_b1 );
not ( \2910_b1 , w_11378 );
and ( \4672_b0 , \777_b0 , w_11379 );
and ( w_11378 , w_11379 , \2910_b0 );
or ( \4673_b1 , \4671_b1 , w_11381 );
not ( w_11381 , w_11382 );
and ( \4673_b0 , \4671_b0 , w_11383 );
and ( w_11382 ,  , w_11383 );
buf ( w_11381 , \4672_b1 );
not ( w_11381 , w_11384 );
not (  , w_11385 );
and ( w_11384 , w_11385 , \4672_b0 );
or ( \4674_b1 , \4673_b1 , w_11386 );
xor ( \4674_b0 , \4673_b0 , w_11388 );
not ( w_11388 , w_11389 );
and ( w_11389 , w_11386 , w_11387 );
buf ( w_11386 , \2371_b1 );
not ( w_11386 , w_11390 );
not ( w_11387 , w_11391 );
and ( w_11390 , w_11391 , \2371_b0 );
or ( \4675_b1 , \1104_b1 , \2550_b1 );
not ( \2550_b1 , w_11392 );
and ( \4675_b0 , \1104_b0 , w_11393 );
and ( w_11392 , w_11393 , \2550_b0 );
or ( \4676_b1 , \904_b1 , \2548_b1 );
not ( \2548_b1 , w_11394 );
and ( \4676_b0 , \904_b0 , w_11395 );
and ( w_11394 , w_11395 , \2548_b0 );
or ( \4677_b1 , \4675_b1 , w_11397 );
not ( w_11397 , w_11398 );
and ( \4677_b0 , \4675_b0 , w_11399 );
and ( w_11398 ,  , w_11399 );
buf ( w_11397 , \4676_b1 );
not ( w_11397 , w_11400 );
not (  , w_11401 );
and ( w_11400 , w_11401 , \4676_b0 );
or ( \4678_b1 , \4677_b1 , w_11402 );
xor ( \4678_b0 , \4677_b0 , w_11404 );
not ( w_11404 , w_11405 );
and ( w_11405 , w_11402 , w_11403 );
buf ( w_11402 , \2374_b1 );
not ( w_11402 , w_11406 );
not ( w_11403 , w_11407 );
and ( w_11406 , w_11407 , \2374_b0 );
or ( \4679_b1 , \4674_b1 , \4678_b1 );
not ( \4678_b1 , w_11408 );
and ( \4679_b0 , \4674_b0 , w_11409 );
and ( w_11408 , w_11409 , \4678_b0 );
or ( \4680_b1 , \4678_b1 , \668_b1 );
not ( \668_b1 , w_11410 );
and ( \4680_b0 , \4678_b0 , w_11411 );
and ( w_11410 , w_11411 , \668_b0 );
or ( \4681_b1 , \4674_b1 , \668_b1 );
not ( \668_b1 , w_11412 );
and ( \4681_b0 , \4674_b0 , w_11413 );
and ( w_11412 , w_11413 , \668_b0 );
or ( \4683_b1 , \2023_b1 , \1476_b1 );
not ( \1476_b1 , w_11414 );
and ( \4683_b0 , \2023_b0 , w_11415 );
and ( w_11414 , w_11415 , \1476_b0 );
or ( \4684_b1 , \1778_b1 , \1474_b1 );
not ( \1474_b1 , w_11416 );
and ( \4684_b0 , \1778_b0 , w_11417 );
and ( w_11416 , w_11417 , \1474_b0 );
or ( \4685_b1 , \4683_b1 , w_11419 );
not ( w_11419 , w_11420 );
and ( \4685_b0 , \4683_b0 , w_11421 );
and ( w_11420 ,  , w_11421 );
buf ( w_11419 , \4684_b1 );
not ( w_11419 , w_11422 );
not (  , w_11423 );
and ( w_11422 , w_11423 , \4684_b0 );
or ( \4686_b1 , \4685_b1 , w_11424 );
xor ( \4686_b0 , \4685_b0 , w_11426 );
not ( w_11426 , w_11427 );
and ( w_11427 , w_11424 , w_11425 );
buf ( w_11424 , \1363_b1 );
not ( w_11424 , w_11428 );
not ( w_11425 , w_11429 );
and ( w_11428 , w_11429 , \1363_b0 );
or ( \4687_b1 , \2161_b1 , \1280_b1 );
not ( \1280_b1 , w_11430 );
and ( \4687_b0 , \2161_b0 , w_11431 );
and ( w_11430 , w_11431 , \1280_b0 );
or ( \4688_b1 , \2028_b1 , \1278_b1 );
not ( \1278_b1 , w_11432 );
and ( \4688_b0 , \2028_b0 , w_11433 );
and ( w_11432 , w_11433 , \1278_b0 );
or ( \4689_b1 , \4687_b1 , w_11435 );
not ( w_11435 , w_11436 );
and ( \4689_b0 , \4687_b0 , w_11437 );
and ( w_11436 ,  , w_11437 );
buf ( w_11435 , \4688_b1 );
not ( w_11435 , w_11438 );
not (  , w_11439 );
and ( w_11438 , w_11439 , \4688_b0 );
or ( \4690_b1 , \4689_b1 , w_11440 );
xor ( \4690_b0 , \4689_b0 , w_11442 );
not ( w_11442 , w_11443 );
and ( w_11443 , w_11440 , w_11441 );
buf ( w_11440 , \1177_b1 );
not ( w_11440 , w_11444 );
not ( w_11441 , w_11445 );
and ( w_11444 , w_11445 , \1177_b0 );
or ( \4691_b1 , \4686_b1 , \4690_b1 );
not ( \4690_b1 , w_11446 );
and ( \4691_b0 , \4686_b0 , w_11447 );
and ( w_11446 , w_11447 , \4690_b0 );
or ( \4692_b1 , \2532_b1 , \1062_b1 );
not ( \1062_b1 , w_11448 );
and ( \4692_b0 , \2532_b0 , w_11449 );
and ( w_11448 , w_11449 , \1062_b0 );
or ( \4693_b1 , \2305_b1 , \1060_b1 );
not ( \1060_b1 , w_11450 );
and ( \4693_b0 , \2305_b0 , w_11451 );
and ( w_11450 , w_11451 , \1060_b0 );
or ( \4694_b1 , \4692_b1 , w_11453 );
not ( w_11453 , w_11454 );
and ( \4694_b0 , \4692_b0 , w_11455 );
and ( w_11454 ,  , w_11455 );
buf ( w_11453 , \4693_b1 );
not ( w_11453 , w_11456 );
not (  , w_11457 );
and ( w_11456 , w_11457 , \4693_b0 );
or ( \4695_b1 , \4694_b1 , w_11458 );
xor ( \4695_b0 , \4694_b0 , w_11460 );
not ( w_11460 , w_11461 );
and ( w_11461 , w_11458 , w_11459 );
buf ( w_11458 , \984_b1 );
not ( w_11458 , w_11462 );
not ( w_11459 , w_11463 );
and ( w_11462 , w_11463 , \984_b0 );
or ( \4696_b1 , \4690_b1 , \4695_b1 );
not ( \4695_b1 , w_11464 );
and ( \4696_b0 , \4690_b0 , w_11465 );
and ( w_11464 , w_11465 , \4695_b0 );
or ( \4697_b1 , \4686_b1 , \4695_b1 );
not ( \4695_b1 , w_11466 );
and ( \4697_b0 , \4686_b0 , w_11467 );
and ( w_11466 , w_11467 , \4695_b0 );
or ( \4699_b1 , \4682_b1 , \4698_b1 );
not ( \4698_b1 , w_11468 );
and ( \4699_b0 , \4682_b0 , w_11469 );
and ( w_11468 , w_11469 , \4698_b0 );
or ( \4700_b1 , \1299_b1 , \2261_b1 );
not ( \2261_b1 , w_11470 );
and ( \4700_b0 , \1299_b0 , w_11471 );
and ( w_11470 , w_11471 , \2261_b0 );
or ( \4701_b1 , \1194_b1 , \2259_b1 );
not ( \2259_b1 , w_11472 );
and ( \4701_b0 , \1194_b0 , w_11473 );
and ( w_11472 , w_11473 , \2259_b0 );
or ( \4702_b1 , \4700_b1 , w_11475 );
not ( w_11475 , w_11476 );
and ( \4702_b0 , \4700_b0 , w_11477 );
and ( w_11476 ,  , w_11477 );
buf ( w_11475 , \4701_b1 );
not ( w_11475 , w_11478 );
not (  , w_11479 );
and ( w_11478 , w_11479 , \4701_b0 );
or ( \4703_b1 , \4702_b1 , w_11480 );
xor ( \4703_b0 , \4702_b0 , w_11482 );
not ( w_11482 , w_11483 );
and ( w_11483 , w_11480 , w_11481 );
buf ( w_11480 , \2124_b1 );
not ( w_11480 , w_11484 );
not ( w_11481 , w_11485 );
and ( w_11484 , w_11485 , \2124_b0 );
or ( \4704_b1 , \1422_b1 , \1955_b1 );
not ( \1955_b1 , w_11486 );
and ( \4704_b0 , \1422_b0 , w_11487 );
and ( w_11486 , w_11487 , \1955_b0 );
or ( \4705_b1 , \1304_b1 , \1953_b1 );
not ( \1953_b1 , w_11488 );
and ( \4705_b0 , \1304_b0 , w_11489 );
and ( w_11488 , w_11489 , \1953_b0 );
or ( \4706_b1 , \4704_b1 , w_11491 );
not ( w_11491 , w_11492 );
and ( \4706_b0 , \4704_b0 , w_11493 );
and ( w_11492 ,  , w_11493 );
buf ( w_11491 , \4705_b1 );
not ( w_11491 , w_11494 );
not (  , w_11495 );
and ( w_11494 , w_11495 , \4705_b0 );
or ( \4707_b1 , \4706_b1 , w_11496 );
xor ( \4707_b0 , \4706_b0 , w_11498 );
not ( w_11498 , w_11499 );
and ( w_11499 , w_11496 , w_11497 );
buf ( w_11496 , \1835_b1 );
not ( w_11496 , w_11500 );
not ( w_11497 , w_11501 );
and ( w_11500 , w_11501 , \1835_b0 );
or ( \4708_b1 , \4703_b1 , \4707_b1 );
not ( \4707_b1 , w_11502 );
and ( \4708_b0 , \4703_b0 , w_11503 );
and ( w_11502 , w_11503 , \4707_b0 );
or ( \4709_b1 , \1770_b1 , \1742_b1 );
not ( \1742_b1 , w_11504 );
and ( \4709_b0 , \1770_b0 , w_11505 );
and ( w_11504 , w_11505 , \1742_b0 );
or ( \4710_b1 , \1537_b1 , \1740_b1 );
not ( \1740_b1 , w_11506 );
and ( \4710_b0 , \1537_b0 , w_11507 );
and ( w_11506 , w_11507 , \1740_b0 );
or ( \4711_b1 , \4709_b1 , w_11509 );
not ( w_11509 , w_11510 );
and ( \4711_b0 , \4709_b0 , w_11511 );
and ( w_11510 ,  , w_11511 );
buf ( w_11509 , \4710_b1 );
not ( w_11509 , w_11512 );
not (  , w_11513 );
and ( w_11512 , w_11513 , \4710_b0 );
or ( \4712_b1 , \4711_b1 , w_11514 );
xor ( \4712_b0 , \4711_b0 , w_11516 );
not ( w_11516 , w_11517 );
and ( w_11517 , w_11514 , w_11515 );
buf ( w_11514 , \1610_b1 );
not ( w_11514 , w_11518 );
not ( w_11515 , w_11519 );
and ( w_11518 , w_11519 , \1610_b0 );
or ( \4713_b1 , \4707_b1 , \4712_b1 );
not ( \4712_b1 , w_11520 );
and ( \4713_b0 , \4707_b0 , w_11521 );
and ( w_11520 , w_11521 , \4712_b0 );
or ( \4714_b1 , \4703_b1 , \4712_b1 );
not ( \4712_b1 , w_11522 );
and ( \4714_b0 , \4703_b0 , w_11523 );
and ( w_11522 , w_11523 , \4712_b0 );
or ( \4716_b1 , \4698_b1 , \4715_b1 );
not ( \4715_b1 , w_11524 );
and ( \4716_b0 , \4698_b0 , w_11525 );
and ( w_11524 , w_11525 , \4715_b0 );
or ( \4717_b1 , \4682_b1 , \4715_b1 );
not ( \4715_b1 , w_11526 );
and ( \4717_b0 , \4682_b0 , w_11527 );
and ( w_11526 , w_11527 , \4715_b0 );
or ( \4719_b1 , \2850_b1 , \740_b1 );
not ( \740_b1 , w_11528 );
and ( \4719_b0 , \2850_b0 , w_11529 );
and ( w_11528 , w_11529 , \740_b0 );
or ( \4720_b1 , \2763_b1 , \738_b1 );
not ( \738_b1 , w_11530 );
and ( \4720_b0 , \2763_b0 , w_11531 );
and ( w_11530 , w_11531 , \738_b0 );
or ( \4721_b1 , \4719_b1 , w_11533 );
not ( w_11533 , w_11534 );
and ( \4721_b0 , \4719_b0 , w_11535 );
and ( w_11534 ,  , w_11535 );
buf ( w_11533 , \4720_b1 );
not ( w_11533 , w_11536 );
not (  , w_11537 );
and ( w_11536 , w_11537 , \4720_b0 );
or ( \4722_b1 , \4721_b1 , w_11538 );
xor ( \4722_b0 , \4721_b0 , w_11540 );
not ( w_11540 , w_11541 );
and ( w_11541 , w_11538 , w_11539 );
buf ( w_11538 , \668_b1 );
not ( w_11538 , w_11542 );
not ( w_11539 , w_11543 );
and ( w_11542 , w_11543 , \668_b0 );
or ( \4723_b1 , \4586_b1 , \4590_b1 );
xor ( \4723_b0 , \4586_b0 , w_11544 );
not ( w_11544 , w_11545 );
and ( w_11545 , \4590_b1 , \4590_b0 );
or ( \4724_b1 , \4723_b1 , \4595_b1 );
xor ( \4724_b0 , \4723_b0 , w_11546 );
not ( w_11546 , w_11547 );
and ( w_11547 , \4595_b1 , \4595_b0 );
or ( \4725_b1 , \4722_b1 , \4724_b1 );
not ( \4724_b1 , w_11548 );
and ( \4725_b0 , \4722_b0 , w_11549 );
and ( w_11548 , w_11549 , \4724_b0 );
or ( \4726_b1 , \4619_b1 , \4623_b1 );
xor ( \4726_b0 , \4619_b0 , w_11550 );
not ( w_11550 , w_11551 );
and ( w_11551 , \4623_b1 , \4623_b0 );
or ( \4727_b1 , \4726_b1 , \4628_b1 );
xor ( \4727_b0 , \4726_b0 , w_11552 );
not ( w_11552 , w_11553 );
and ( w_11553 , \4628_b1 , \4628_b0 );
or ( \4728_b1 , \4724_b1 , \4727_b1 );
not ( \4727_b1 , w_11554 );
and ( \4728_b0 , \4724_b0 , w_11555 );
and ( w_11554 , w_11555 , \4727_b0 );
or ( \4729_b1 , \4722_b1 , \4727_b1 );
not ( \4727_b1 , w_11556 );
and ( \4729_b0 , \4722_b0 , w_11557 );
and ( w_11556 , w_11557 , \4727_b0 );
or ( \4731_b1 , \4718_b1 , \4730_b1 );
not ( \4730_b1 , w_11558 );
and ( \4731_b0 , \4718_b0 , w_11559 );
and ( w_11558 , w_11559 , \4730_b0 );
or ( \4732_b1 , \4497_b1 , \4501_b1 );
xor ( \4732_b0 , \4497_b0 , w_11560 );
not ( w_11560 , w_11561 );
and ( w_11561 , \4501_b1 , \4501_b0 );
or ( \4733_b1 , \4732_b1 , \561_b1 );
xor ( \4733_b0 , \4732_b0 , w_11562 );
not ( w_11562 , w_11563 );
and ( w_11563 , \561_b1 , \561_b0 );
or ( \4734_b1 , \4730_b1 , \4733_b1 );
not ( \4733_b1 , w_11564 );
and ( \4734_b0 , \4730_b0 , w_11565 );
and ( w_11564 , w_11565 , \4733_b0 );
or ( \4735_b1 , \4718_b1 , \4733_b1 );
not ( \4733_b1 , w_11566 );
and ( \4735_b0 , \4718_b0 , w_11567 );
and ( w_11566 , w_11567 , \4733_b0 );
or ( \4737_b1 , \4598_b1 , \4614_b1 );
xor ( \4737_b0 , \4598_b0 , w_11568 );
not ( w_11568 , w_11569 );
and ( w_11569 , \4614_b1 , \4614_b0 );
or ( \4738_b1 , \4737_b1 , \4631_b1 );
xor ( \4738_b0 , \4737_b0 , w_11570 );
not ( w_11570 , w_11571 );
and ( w_11571 , \4631_b1 , \4631_b0 );
or ( \4739_b1 , \4636_b1 , \4638_b1 );
xor ( \4739_b0 , \4636_b0 , w_11572 );
not ( w_11572 , w_11573 );
and ( w_11573 , \4638_b1 , \4638_b0 );
or ( \4740_b1 , \4739_b1 , \4641_b1 );
xor ( \4740_b0 , \4739_b0 , w_11574 );
not ( w_11574 , w_11575 );
and ( w_11575 , \4641_b1 , \4641_b0 );
or ( \4741_b1 , \4738_b1 , \4740_b1 );
not ( \4740_b1 , w_11576 );
and ( \4741_b0 , \4738_b0 , w_11577 );
and ( w_11576 , w_11577 , \4740_b0 );
or ( \4742_b1 , \4736_b1 , \4741_b1 );
not ( \4741_b1 , w_11578 );
and ( \4742_b0 , \4736_b0 , w_11579 );
and ( w_11578 , w_11579 , \4741_b0 );
or ( \4743_b1 , \4481_b1 , \4485_b1 );
xor ( \4743_b0 , \4481_b0 , w_11580 );
not ( w_11580 , w_11581 );
and ( w_11581 , \4485_b1 , \4485_b0 );
or ( \4744_b1 , \4743_b1 , \4490_b1 );
xor ( \4744_b0 , \4743_b0 , w_11582 );
not ( w_11582 , w_11583 );
and ( w_11583 , \4490_b1 , \4490_b0 );
or ( \4745_b1 , \4741_b1 , \4744_b1 );
not ( \4744_b1 , w_11584 );
and ( \4745_b0 , \4741_b0 , w_11585 );
and ( w_11584 , w_11585 , \4744_b0 );
or ( \4746_b1 , \4736_b1 , \4744_b1 );
not ( \4744_b1 , w_11586 );
and ( \4746_b0 , \4736_b0 , w_11587 );
and ( w_11586 , w_11587 , \4744_b0 );
or ( \4748_b1 , \4505_b1 , \4521_b1 );
xor ( \4748_b0 , \4505_b0 , w_11588 );
not ( w_11588 , w_11589 );
and ( w_11589 , \4521_b1 , \4521_b0 );
or ( \4749_b1 , \4748_b1 , \4538_b1 );
xor ( \4749_b0 , \4748_b0 , w_11590 );
not ( w_11590 , w_11591 );
and ( w_11591 , \4538_b1 , \4538_b0 );
or ( \4750_b1 , \4634_b1 , \4644_b1 );
xor ( \4750_b0 , \4634_b0 , w_11592 );
not ( w_11592 , w_11593 );
and ( w_11593 , \4644_b1 , \4644_b0 );
or ( \4751_b1 , \4750_b1 , \4647_b1 );
xor ( \4751_b0 , \4750_b0 , w_11594 );
not ( w_11594 , w_11595 );
and ( w_11595 , \4647_b1 , \4647_b0 );
or ( \4752_b1 , \4749_b1 , \4751_b1 );
not ( \4751_b1 , w_11596 );
and ( \4752_b0 , \4749_b0 , w_11597 );
and ( w_11596 , w_11597 , \4751_b0 );
or ( \4753_b1 , \4747_b1 , \4752_b1 );
not ( \4752_b1 , w_11598 );
and ( \4753_b0 , \4747_b0 , w_11599 );
and ( w_11598 , w_11599 , \4752_b0 );
or ( \4754_b1 , \4650_b1 , \4652_b1 );
xor ( \4754_b0 , \4650_b0 , w_11600 );
not ( w_11600 , w_11601 );
and ( w_11601 , \4652_b1 , \4652_b0 );
or ( \4755_b1 , \4754_b1 , \4655_b1 );
xor ( \4755_b0 , \4754_b0 , w_11602 );
not ( w_11602 , w_11603 );
and ( w_11603 , \4655_b1 , \4655_b0 );
or ( \4756_b1 , \4752_b1 , \4755_b1 );
not ( \4755_b1 , w_11604 );
and ( \4756_b0 , \4752_b0 , w_11605 );
and ( w_11604 , w_11605 , \4755_b0 );
or ( \4757_b1 , \4747_b1 , \4755_b1 );
not ( \4755_b1 , w_11606 );
and ( \4757_b0 , \4747_b0 , w_11607 );
and ( w_11606 , w_11607 , \4755_b0 );
or ( \4759_b1 , \4670_b1 , \4758_b1 );
not ( \4758_b1 , w_11608 );
and ( \4759_b0 , \4670_b0 , w_11609 );
and ( w_11608 , w_11609 , \4758_b0 );
or ( \4760_b1 , \4670_b1 , \4758_b1 );
xor ( \4760_b0 , \4670_b0 , w_11610 );
not ( w_11610 , w_11611 );
and ( w_11611 , \4758_b1 , \4758_b0 );
or ( \4761_b1 , \4747_b1 , \4752_b1 );
xor ( \4761_b0 , \4747_b0 , w_11612 );
not ( w_11612 , w_11613 );
and ( w_11613 , \4752_b1 , \4752_b0 );
or ( \4762_b1 , \4761_b1 , \4755_b1 );
xor ( \4762_b0 , \4761_b0 , w_11614 );
not ( w_11614 , w_11615 );
and ( w_11615 , \4755_b1 , \4755_b0 );
or ( \4763_b1 , \1537_b1 , \1955_b1 );
not ( \1955_b1 , w_11616 );
and ( \4763_b0 , \1537_b0 , w_11617 );
and ( w_11616 , w_11617 , \1955_b0 );
or ( \4764_b1 , \1422_b1 , \1953_b1 );
not ( \1953_b1 , w_11618 );
and ( \4764_b0 , \1422_b0 , w_11619 );
and ( w_11618 , w_11619 , \1953_b0 );
or ( \4765_b1 , \4763_b1 , w_11621 );
not ( w_11621 , w_11622 );
and ( \4765_b0 , \4763_b0 , w_11623 );
and ( w_11622 ,  , w_11623 );
buf ( w_11621 , \4764_b1 );
not ( w_11621 , w_11624 );
not (  , w_11625 );
and ( w_11624 , w_11625 , \4764_b0 );
or ( \4766_b1 , \4765_b1 , w_11626 );
xor ( \4766_b0 , \4765_b0 , w_11628 );
not ( w_11628 , w_11629 );
and ( w_11629 , w_11626 , w_11627 );
buf ( w_11626 , \1835_b1 );
not ( w_11626 , w_11630 );
not ( w_11627 , w_11631 );
and ( w_11630 , w_11631 , \1835_b0 );
or ( \4767_b1 , \1778_b1 , \1742_b1 );
not ( \1742_b1 , w_11632 );
and ( \4767_b0 , \1778_b0 , w_11633 );
and ( w_11632 , w_11633 , \1742_b0 );
or ( \4768_b1 , \1770_b1 , \1740_b1 );
not ( \1740_b1 , w_11634 );
and ( \4768_b0 , \1770_b0 , w_11635 );
and ( w_11634 , w_11635 , \1740_b0 );
or ( \4769_b1 , \4767_b1 , w_11637 );
not ( w_11637 , w_11638 );
and ( \4769_b0 , \4767_b0 , w_11639 );
and ( w_11638 ,  , w_11639 );
buf ( w_11637 , \4768_b1 );
not ( w_11637 , w_11640 );
not (  , w_11641 );
and ( w_11640 , w_11641 , \4768_b0 );
or ( \4770_b1 , \4769_b1 , w_11642 );
xor ( \4770_b0 , \4769_b0 , w_11644 );
not ( w_11644 , w_11645 );
and ( w_11645 , w_11642 , w_11643 );
buf ( w_11642 , \1610_b1 );
not ( w_11642 , w_11646 );
not ( w_11643 , w_11647 );
and ( w_11646 , w_11647 , \1610_b0 );
or ( \4771_b1 , \4766_b1 , \4770_b1 );
not ( \4770_b1 , w_11648 );
and ( \4771_b0 , \4766_b0 , w_11649 );
and ( w_11648 , w_11649 , \4770_b0 );
or ( \4772_b1 , \2028_b1 , \1476_b1 );
not ( \1476_b1 , w_11650 );
and ( \4772_b0 , \2028_b0 , w_11651 );
and ( w_11650 , w_11651 , \1476_b0 );
or ( \4773_b1 , \2023_b1 , \1474_b1 );
not ( \1474_b1 , w_11652 );
and ( \4773_b0 , \2023_b0 , w_11653 );
and ( w_11652 , w_11653 , \1474_b0 );
or ( \4774_b1 , \4772_b1 , w_11655 );
not ( w_11655 , w_11656 );
and ( \4774_b0 , \4772_b0 , w_11657 );
and ( w_11656 ,  , w_11657 );
buf ( w_11655 , \4773_b1 );
not ( w_11655 , w_11658 );
not (  , w_11659 );
and ( w_11658 , w_11659 , \4773_b0 );
or ( \4775_b1 , \4774_b1 , w_11660 );
xor ( \4775_b0 , \4774_b0 , w_11662 );
not ( w_11662 , w_11663 );
and ( w_11663 , w_11660 , w_11661 );
buf ( w_11660 , \1363_b1 );
not ( w_11660 , w_11664 );
not ( w_11661 , w_11665 );
and ( w_11664 , w_11665 , \1363_b0 );
or ( \4776_b1 , \4770_b1 , \4775_b1 );
not ( \4775_b1 , w_11666 );
and ( \4776_b0 , \4770_b0 , w_11667 );
and ( w_11666 , w_11667 , \4775_b0 );
or ( \4777_b1 , \4766_b1 , \4775_b1 );
not ( \4775_b1 , w_11668 );
and ( \4777_b0 , \4766_b0 , w_11669 );
and ( w_11668 , w_11669 , \4775_b0 );
or ( \4779_b1 , \904_b1 , \2913_b1 );
not ( \2913_b1 , w_11670 );
and ( \4779_b0 , \904_b0 , w_11671 );
and ( w_11670 , w_11671 , \2913_b0 );
or ( \4780_b1 , \841_b1 , \2910_b1 );
not ( \2910_b1 , w_11672 );
and ( \4780_b0 , \841_b0 , w_11673 );
and ( w_11672 , w_11673 , \2910_b0 );
or ( \4781_b1 , \4779_b1 , w_11675 );
not ( w_11675 , w_11676 );
and ( \4781_b0 , \4779_b0 , w_11677 );
and ( w_11676 ,  , w_11677 );
buf ( w_11675 , \4780_b1 );
not ( w_11675 , w_11678 );
not (  , w_11679 );
and ( w_11678 , w_11679 , \4780_b0 );
or ( \4782_b1 , \4781_b1 , w_11680 );
xor ( \4782_b0 , \4781_b0 , w_11682 );
not ( w_11682 , w_11683 );
and ( w_11683 , w_11680 , w_11681 );
buf ( w_11680 , \2371_b1 );
not ( w_11680 , w_11684 );
not ( w_11681 , w_11685 );
and ( w_11684 , w_11685 , \2371_b0 );
or ( \4783_b1 , \1194_b1 , \2550_b1 );
not ( \2550_b1 , w_11686 );
and ( \4783_b0 , \1194_b0 , w_11687 );
and ( w_11686 , w_11687 , \2550_b0 );
or ( \4784_b1 , \1104_b1 , \2548_b1 );
not ( \2548_b1 , w_11688 );
and ( \4784_b0 , \1104_b0 , w_11689 );
and ( w_11688 , w_11689 , \2548_b0 );
or ( \4785_b1 , \4783_b1 , w_11691 );
not ( w_11691 , w_11692 );
and ( \4785_b0 , \4783_b0 , w_11693 );
and ( w_11692 ,  , w_11693 );
buf ( w_11691 , \4784_b1 );
not ( w_11691 , w_11694 );
not (  , w_11695 );
and ( w_11694 , w_11695 , \4784_b0 );
or ( \4786_b1 , \4785_b1 , w_11696 );
xor ( \4786_b0 , \4785_b0 , w_11698 );
not ( w_11698 , w_11699 );
and ( w_11699 , w_11696 , w_11697 );
buf ( w_11696 , \2374_b1 );
not ( w_11696 , w_11700 );
not ( w_11697 , w_11701 );
and ( w_11700 , w_11701 , \2374_b0 );
or ( \4787_b1 , \4782_b1 , \4786_b1 );
not ( \4786_b1 , w_11702 );
and ( \4787_b0 , \4782_b0 , w_11703 );
and ( w_11702 , w_11703 , \4786_b0 );
or ( \4788_b1 , \1304_b1 , \2261_b1 );
not ( \2261_b1 , w_11704 );
and ( \4788_b0 , \1304_b0 , w_11705 );
and ( w_11704 , w_11705 , \2261_b0 );
or ( \4789_b1 , \1299_b1 , \2259_b1 );
not ( \2259_b1 , w_11706 );
and ( \4789_b0 , \1299_b0 , w_11707 );
and ( w_11706 , w_11707 , \2259_b0 );
or ( \4790_b1 , \4788_b1 , w_11709 );
not ( w_11709 , w_11710 );
and ( \4790_b0 , \4788_b0 , w_11711 );
and ( w_11710 ,  , w_11711 );
buf ( w_11709 , \4789_b1 );
not ( w_11709 , w_11712 );
not (  , w_11713 );
and ( w_11712 , w_11713 , \4789_b0 );
or ( \4791_b1 , \4790_b1 , w_11714 );
xor ( \4791_b0 , \4790_b0 , w_11716 );
not ( w_11716 , w_11717 );
and ( w_11717 , w_11714 , w_11715 );
buf ( w_11714 , \2124_b1 );
not ( w_11714 , w_11718 );
not ( w_11715 , w_11719 );
and ( w_11718 , w_11719 , \2124_b0 );
or ( \4792_b1 , \4786_b1 , \4791_b1 );
not ( \4791_b1 , w_11720 );
and ( \4792_b0 , \4786_b0 , w_11721 );
and ( w_11720 , w_11721 , \4791_b0 );
or ( \4793_b1 , \4782_b1 , \4791_b1 );
not ( \4791_b1 , w_11722 );
and ( \4793_b0 , \4782_b0 , w_11723 );
and ( w_11722 , w_11723 , \4791_b0 );
or ( \4795_b1 , \4778_b1 , \4794_b1 );
not ( \4794_b1 , w_11724 );
and ( \4795_b0 , \4778_b0 , w_11725 );
and ( w_11724 , w_11725 , \4794_b0 );
or ( \4796_b1 , \2305_b1 , \1280_b1 );
not ( \1280_b1 , w_11726 );
and ( \4796_b0 , \2305_b0 , w_11727 );
and ( w_11726 , w_11727 , \1280_b0 );
or ( \4797_b1 , \2161_b1 , \1278_b1 );
not ( \1278_b1 , w_11728 );
and ( \4797_b0 , \2161_b0 , w_11729 );
and ( w_11728 , w_11729 , \1278_b0 );
or ( \4798_b1 , \4796_b1 , w_11731 );
not ( w_11731 , w_11732 );
and ( \4798_b0 , \4796_b0 , w_11733 );
and ( w_11732 ,  , w_11733 );
buf ( w_11731 , \4797_b1 );
not ( w_11731 , w_11734 );
not (  , w_11735 );
and ( w_11734 , w_11735 , \4797_b0 );
or ( \4799_b1 , \4798_b1 , w_11736 );
xor ( \4799_b0 , \4798_b0 , w_11738 );
not ( w_11738 , w_11739 );
and ( w_11739 , w_11736 , w_11737 );
buf ( w_11736 , \1177_b1 );
not ( w_11736 , w_11740 );
not ( w_11737 , w_11741 );
and ( w_11740 , w_11741 , \1177_b0 );
or ( \4800_b1 , \2541_b1 , \1062_b1 );
not ( \1062_b1 , w_11742 );
and ( \4800_b0 , \2541_b0 , w_11743 );
and ( w_11742 , w_11743 , \1062_b0 );
or ( \4801_b1 , \2532_b1 , \1060_b1 );
not ( \1060_b1 , w_11744 );
and ( \4801_b0 , \2532_b0 , w_11745 );
and ( w_11744 , w_11745 , \1060_b0 );
or ( \4802_b1 , \4800_b1 , w_11747 );
not ( w_11747 , w_11748 );
and ( \4802_b0 , \4800_b0 , w_11749 );
and ( w_11748 ,  , w_11749 );
buf ( w_11747 , \4801_b1 );
not ( w_11747 , w_11750 );
not (  , w_11751 );
and ( w_11750 , w_11751 , \4801_b0 );
or ( \4803_b1 , \4802_b1 , w_11752 );
xor ( \4803_b0 , \4802_b0 , w_11754 );
not ( w_11754 , w_11755 );
and ( w_11755 , w_11752 , w_11753 );
buf ( w_11752 , \984_b1 );
not ( w_11752 , w_11756 );
not ( w_11753 , w_11757 );
and ( w_11756 , w_11757 , \984_b0 );
or ( \4804_b1 , \4799_b1 , \4803_b1 );
not ( \4803_b1 , w_11758 );
and ( \4804_b0 , \4799_b0 , w_11759 );
and ( w_11758 , w_11759 , \4803_b0 );
or ( \4805_b1 , \2850_b1 , \912_b1 );
not ( \912_b1 , w_11760 );
and ( \4805_b0 , \2850_b0 , w_11761 );
and ( w_11760 , w_11761 , \912_b0 );
or ( \4806_b1 , \2763_b1 , \910_b1 );
not ( \910_b1 , w_11762 );
and ( \4806_b0 , \2763_b0 , w_11763 );
and ( w_11762 , w_11763 , \910_b0 );
or ( \4807_b1 , \4805_b1 , w_11765 );
not ( w_11765 , w_11766 );
and ( \4807_b0 , \4805_b0 , w_11767 );
and ( w_11766 ,  , w_11767 );
buf ( w_11765 , \4806_b1 );
not ( w_11765 , w_11768 );
not (  , w_11769 );
and ( w_11768 , w_11769 , \4806_b0 );
or ( \4808_b1 , \4807_b1 , w_11770 );
xor ( \4808_b0 , \4807_b0 , w_11772 );
not ( w_11772 , w_11773 );
and ( w_11773 , w_11770 , w_11771 );
buf ( w_11770 , \818_b1 );
not ( w_11770 , w_11774 );
not ( w_11771 , w_11775 );
and ( w_11774 , w_11775 , \818_b0 );
or ( \4809_b1 , \4803_b1 , \4808_b1 );
not ( \4808_b1 , w_11776 );
and ( \4809_b0 , \4803_b0 , w_11777 );
and ( w_11776 , w_11777 , \4808_b0 );
or ( \4810_b1 , \4799_b1 , \4808_b1 );
not ( \4808_b1 , w_11778 );
and ( \4810_b0 , \4799_b0 , w_11779 );
and ( w_11778 , w_11779 , \4808_b0 );
or ( \4812_b1 , \4794_b1 , \4811_b1 );
not ( \4811_b1 , w_11780 );
and ( \4812_b0 , \4794_b0 , w_11781 );
and ( w_11780 , w_11781 , \4811_b0 );
or ( \4813_b1 , \4778_b1 , \4811_b1 );
not ( \4811_b1 , w_11782 );
and ( \4813_b0 , \4778_b0 , w_11783 );
and ( w_11782 , w_11783 , \4811_b0 );
or ( \4815_b1 , \2763_b1 , \912_b1 );
not ( \912_b1 , w_11784 );
and ( \4815_b0 , \2763_b0 , w_11785 );
and ( w_11784 , w_11785 , \912_b0 );
or ( \4816_b1 , \2541_b1 , \910_b1 );
not ( \910_b1 , w_11786 );
and ( \4816_b0 , \2541_b0 , w_11787 );
and ( w_11786 , w_11787 , \910_b0 );
or ( \4817_b1 , \4815_b1 , w_11789 );
not ( w_11789 , w_11790 );
and ( \4817_b0 , \4815_b0 , w_11791 );
and ( w_11790 ,  , w_11791 );
buf ( w_11789 , \4816_b1 );
not ( w_11789 , w_11792 );
not (  , w_11793 );
and ( w_11792 , w_11793 , \4816_b0 );
or ( \4818_b1 , \4817_b1 , w_11794 );
xor ( \4818_b0 , \4817_b0 , w_11796 );
not ( w_11796 , w_11797 );
and ( w_11797 , w_11794 , w_11795 );
buf ( w_11794 , \818_b1 );
not ( w_11794 , w_11798 );
not ( w_11795 , w_11799 );
and ( w_11798 , w_11799 , \818_b0 );
or ( \4819_b1 , \2850_b1 , w_11801 );
not ( w_11801 , w_11802 );
and ( \4819_b0 , \2850_b0 , w_11803 );
and ( w_11802 ,  , w_11803 );
buf ( w_11801 , \738_b1 );
not ( w_11801 , w_11804 );
not (  , w_11805 );
and ( w_11804 , w_11805 , \738_b0 );
or ( \4820_b1 , \4819_b1 , w_11806 );
xor ( \4820_b0 , \4819_b0 , w_11808 );
not ( w_11808 , w_11809 );
and ( w_11809 , w_11806 , w_11807 );
buf ( w_11806 , \668_b1 );
not ( w_11806 , w_11810 );
not ( w_11807 , w_11811 );
and ( w_11810 , w_11811 , \668_b0 );
or ( \4821_b1 , \4818_b1 , \4820_b1 );
not ( \4820_b1 , w_11812 );
and ( \4821_b0 , \4818_b0 , w_11813 );
and ( w_11812 , w_11813 , \4820_b0 );
or ( \4822_b1 , \4686_b1 , \4690_b1 );
xor ( \4822_b0 , \4686_b0 , w_11814 );
not ( w_11814 , w_11815 );
and ( w_11815 , \4690_b1 , \4690_b0 );
or ( \4823_b1 , \4822_b1 , \4695_b1 );
xor ( \4823_b0 , \4822_b0 , w_11816 );
not ( w_11816 , w_11817 );
and ( w_11817 , \4695_b1 , \4695_b0 );
or ( \4824_b1 , \4820_b1 , \4823_b1 );
not ( \4823_b1 , w_11818 );
and ( \4824_b0 , \4820_b0 , w_11819 );
and ( w_11818 , w_11819 , \4823_b0 );
or ( \4825_b1 , \4818_b1 , \4823_b1 );
not ( \4823_b1 , w_11820 );
and ( \4825_b0 , \4818_b0 , w_11821 );
and ( w_11820 , w_11821 , \4823_b0 );
or ( \4827_b1 , \4814_b1 , \4826_b1 );
not ( \4826_b1 , w_11822 );
and ( \4827_b0 , \4814_b0 , w_11823 );
and ( w_11822 , w_11823 , \4826_b0 );
or ( \4828_b1 , \4602_b1 , \4606_b1 );
xor ( \4828_b0 , \4602_b0 , w_11824 );
not ( w_11824 , w_11825 );
and ( w_11825 , \4606_b1 , \4606_b0 );
or ( \4829_b1 , \4828_b1 , \4611_b1 );
xor ( \4829_b0 , \4828_b0 , w_11826 );
not ( w_11826 , w_11827 );
and ( w_11827 , \4611_b1 , \4611_b0 );
or ( \4830_b1 , \4826_b1 , \4829_b1 );
not ( \4829_b1 , w_11828 );
and ( \4830_b0 , \4826_b0 , w_11829 );
and ( w_11828 , w_11829 , \4829_b0 );
or ( \4831_b1 , \4814_b1 , \4829_b1 );
not ( \4829_b1 , w_11830 );
and ( \4831_b0 , \4814_b0 , w_11831 );
and ( w_11830 , w_11831 , \4829_b0 );
or ( \4833_b1 , \4718_b1 , \4730_b1 );
xor ( \4833_b0 , \4718_b0 , w_11832 );
not ( w_11832 , w_11833 );
and ( w_11833 , \4730_b1 , \4730_b0 );
or ( \4834_b1 , \4833_b1 , \4733_b1 );
xor ( \4834_b0 , \4833_b0 , w_11834 );
not ( w_11834 , w_11835 );
and ( w_11835 , \4733_b1 , \4733_b0 );
or ( \4835_b1 , \4832_b1 , \4834_b1 );
not ( \4834_b1 , w_11836 );
and ( \4835_b0 , \4832_b0 , w_11837 );
and ( w_11836 , w_11837 , \4834_b0 );
or ( \4836_b1 , \4738_b1 , \4740_b1 );
xor ( \4836_b0 , \4738_b0 , w_11838 );
not ( w_11838 , w_11839 );
and ( w_11839 , \4740_b1 , \4740_b0 );
or ( \4837_b1 , \4834_b1 , \4836_b1 );
not ( \4836_b1 , w_11840 );
and ( \4837_b0 , \4834_b0 , w_11841 );
and ( w_11840 , w_11841 , \4836_b0 );
or ( \4838_b1 , \4832_b1 , \4836_b1 );
not ( \4836_b1 , w_11842 );
and ( \4838_b0 , \4832_b0 , w_11843 );
and ( w_11842 , w_11843 , \4836_b0 );
or ( \4840_b1 , \4736_b1 , \4741_b1 );
xor ( \4840_b0 , \4736_b0 , w_11844 );
not ( w_11844 , w_11845 );
and ( w_11845 , \4741_b1 , \4741_b0 );
or ( \4841_b1 , \4840_b1 , \4744_b1 );
xor ( \4841_b0 , \4840_b0 , w_11846 );
not ( w_11846 , w_11847 );
and ( w_11847 , \4744_b1 , \4744_b0 );
or ( \4842_b1 , \4839_b1 , \4841_b1 );
not ( \4841_b1 , w_11848 );
and ( \4842_b0 , \4839_b0 , w_11849 );
and ( w_11848 , w_11849 , \4841_b0 );
or ( \4843_b1 , \4749_b1 , \4751_b1 );
xor ( \4843_b0 , \4749_b0 , w_11850 );
not ( w_11850 , w_11851 );
and ( w_11851 , \4751_b1 , \4751_b0 );
or ( \4844_b1 , \4841_b1 , \4843_b1 );
not ( \4843_b1 , w_11852 );
and ( \4844_b0 , \4841_b0 , w_11853 );
and ( w_11852 , w_11853 , \4843_b0 );
or ( \4845_b1 , \4839_b1 , \4843_b1 );
not ( \4843_b1 , w_11854 );
and ( \4845_b0 , \4839_b0 , w_11855 );
and ( w_11854 , w_11855 , \4843_b0 );
or ( \4847_b1 , \4762_b1 , \4846_b1 );
not ( \4846_b1 , w_11856 );
and ( \4847_b0 , \4762_b0 , w_11857 );
and ( w_11856 , w_11857 , \4846_b0 );
or ( \4848_b1 , \4762_b1 , \4846_b1 );
xor ( \4848_b0 , \4762_b0 , w_11858 );
not ( w_11858 , w_11859 );
and ( w_11859 , \4846_b1 , \4846_b0 );
or ( \4849_b1 , \4839_b1 , \4841_b1 );
xor ( \4849_b0 , \4839_b0 , w_11860 );
not ( w_11860 , w_11861 );
and ( w_11861 , \4841_b1 , \4841_b0 );
or ( \4850_b1 , \4849_b1 , \4843_b1 );
xor ( \4850_b0 , \4849_b0 , w_11862 );
not ( w_11862 , w_11863 );
and ( w_11863 , \4843_b1 , \4843_b0 );
or ( \4851_b1 , \1422_b1 , \2261_b1 );
not ( \2261_b1 , w_11864 );
and ( \4851_b0 , \1422_b0 , w_11865 );
and ( w_11864 , w_11865 , \2261_b0 );
or ( \4852_b1 , \1304_b1 , \2259_b1 );
not ( \2259_b1 , w_11866 );
and ( \4852_b0 , \1304_b0 , w_11867 );
and ( w_11866 , w_11867 , \2259_b0 );
or ( \4853_b1 , \4851_b1 , w_11869 );
not ( w_11869 , w_11870 );
and ( \4853_b0 , \4851_b0 , w_11871 );
and ( w_11870 ,  , w_11871 );
buf ( w_11869 , \4852_b1 );
not ( w_11869 , w_11872 );
not (  , w_11873 );
and ( w_11872 , w_11873 , \4852_b0 );
or ( \4854_b1 , \4853_b1 , w_11874 );
xor ( \4854_b0 , \4853_b0 , w_11876 );
not ( w_11876 , w_11877 );
and ( w_11877 , w_11874 , w_11875 );
buf ( w_11874 , \2124_b1 );
not ( w_11874 , w_11878 );
not ( w_11875 , w_11879 );
and ( w_11878 , w_11879 , \2124_b0 );
or ( \4855_b1 , \1770_b1 , \1955_b1 );
not ( \1955_b1 , w_11880 );
and ( \4855_b0 , \1770_b0 , w_11881 );
and ( w_11880 , w_11881 , \1955_b0 );
or ( \4856_b1 , \1537_b1 , \1953_b1 );
not ( \1953_b1 , w_11882 );
and ( \4856_b0 , \1537_b0 , w_11883 );
and ( w_11882 , w_11883 , \1953_b0 );
or ( \4857_b1 , \4855_b1 , w_11885 );
not ( w_11885 , w_11886 );
and ( \4857_b0 , \4855_b0 , w_11887 );
and ( w_11886 ,  , w_11887 );
buf ( w_11885 , \4856_b1 );
not ( w_11885 , w_11888 );
not (  , w_11889 );
and ( w_11888 , w_11889 , \4856_b0 );
or ( \4858_b1 , \4857_b1 , w_11890 );
xor ( \4858_b0 , \4857_b0 , w_11892 );
not ( w_11892 , w_11893 );
and ( w_11893 , w_11890 , w_11891 );
buf ( w_11890 , \1835_b1 );
not ( w_11890 , w_11894 );
not ( w_11891 , w_11895 );
and ( w_11894 , w_11895 , \1835_b0 );
or ( \4859_b1 , \4854_b1 , \4858_b1 );
not ( \4858_b1 , w_11896 );
and ( \4859_b0 , \4854_b0 , w_11897 );
and ( w_11896 , w_11897 , \4858_b0 );
or ( \4860_b1 , \2023_b1 , \1742_b1 );
not ( \1742_b1 , w_11898 );
and ( \4860_b0 , \2023_b0 , w_11899 );
and ( w_11898 , w_11899 , \1742_b0 );
or ( \4861_b1 , \1778_b1 , \1740_b1 );
not ( \1740_b1 , w_11900 );
and ( \4861_b0 , \1778_b0 , w_11901 );
and ( w_11900 , w_11901 , \1740_b0 );
or ( \4862_b1 , \4860_b1 , w_11903 );
not ( w_11903 , w_11904 );
and ( \4862_b0 , \4860_b0 , w_11905 );
and ( w_11904 ,  , w_11905 );
buf ( w_11903 , \4861_b1 );
not ( w_11903 , w_11906 );
not (  , w_11907 );
and ( w_11906 , w_11907 , \4861_b0 );
or ( \4863_b1 , \4862_b1 , w_11908 );
xor ( \4863_b0 , \4862_b0 , w_11910 );
not ( w_11910 , w_11911 );
and ( w_11911 , w_11908 , w_11909 );
buf ( w_11908 , \1610_b1 );
not ( w_11908 , w_11912 );
not ( w_11909 , w_11913 );
and ( w_11912 , w_11913 , \1610_b0 );
or ( \4864_b1 , \4858_b1 , \4863_b1 );
not ( \4863_b1 , w_11914 );
and ( \4864_b0 , \4858_b0 , w_11915 );
and ( w_11914 , w_11915 , \4863_b0 );
or ( \4865_b1 , \4854_b1 , \4863_b1 );
not ( \4863_b1 , w_11916 );
and ( \4865_b0 , \4854_b0 , w_11917 );
and ( w_11916 , w_11917 , \4863_b0 );
or ( \4867_b1 , \1104_b1 , \2913_b1 );
not ( \2913_b1 , w_11918 );
and ( \4867_b0 , \1104_b0 , w_11919 );
and ( w_11918 , w_11919 , \2913_b0 );
or ( \4868_b1 , \904_b1 , \2910_b1 );
not ( \2910_b1 , w_11920 );
and ( \4868_b0 , \904_b0 , w_11921 );
and ( w_11920 , w_11921 , \2910_b0 );
or ( \4869_b1 , \4867_b1 , w_11923 );
not ( w_11923 , w_11924 );
and ( \4869_b0 , \4867_b0 , w_11925 );
and ( w_11924 ,  , w_11925 );
buf ( w_11923 , \4868_b1 );
not ( w_11923 , w_11926 );
not (  , w_11927 );
and ( w_11926 , w_11927 , \4868_b0 );
or ( \4870_b1 , \4869_b1 , w_11928 );
xor ( \4870_b0 , \4869_b0 , w_11930 );
not ( w_11930 , w_11931 );
and ( w_11931 , w_11928 , w_11929 );
buf ( w_11928 , \2371_b1 );
not ( w_11928 , w_11932 );
not ( w_11929 , w_11933 );
and ( w_11932 , w_11933 , \2371_b0 );
or ( \4871_b1 , \1299_b1 , \2550_b1 );
not ( \2550_b1 , w_11934 );
and ( \4871_b0 , \1299_b0 , w_11935 );
and ( w_11934 , w_11935 , \2550_b0 );
or ( \4872_b1 , \1194_b1 , \2548_b1 );
not ( \2548_b1 , w_11936 );
and ( \4872_b0 , \1194_b0 , w_11937 );
and ( w_11936 , w_11937 , \2548_b0 );
or ( \4873_b1 , \4871_b1 , w_11939 );
not ( w_11939 , w_11940 );
and ( \4873_b0 , \4871_b0 , w_11941 );
and ( w_11940 ,  , w_11941 );
buf ( w_11939 , \4872_b1 );
not ( w_11939 , w_11942 );
not (  , w_11943 );
and ( w_11942 , w_11943 , \4872_b0 );
or ( \4874_b1 , \4873_b1 , w_11944 );
xor ( \4874_b0 , \4873_b0 , w_11946 );
not ( w_11946 , w_11947 );
and ( w_11947 , w_11944 , w_11945 );
buf ( w_11944 , \2374_b1 );
not ( w_11944 , w_11948 );
not ( w_11945 , w_11949 );
and ( w_11948 , w_11949 , \2374_b0 );
or ( \4875_b1 , \4870_b1 , \4874_b1 );
not ( \4874_b1 , w_11950 );
and ( \4875_b0 , \4870_b0 , w_11951 );
and ( w_11950 , w_11951 , \4874_b0 );
or ( \4876_b1 , \4874_b1 , \818_b1 );
not ( \818_b1 , w_11952 );
and ( \4876_b0 , \4874_b0 , w_11953 );
and ( w_11952 , w_11953 , \818_b0 );
or ( \4877_b1 , \4870_b1 , \818_b1 );
not ( \818_b1 , w_11954 );
and ( \4877_b0 , \4870_b0 , w_11955 );
and ( w_11954 , w_11955 , \818_b0 );
or ( \4879_b1 , \4866_b1 , \4878_b1 );
not ( \4878_b1 , w_11956 );
and ( \4879_b0 , \4866_b0 , w_11957 );
and ( w_11956 , w_11957 , \4878_b0 );
or ( \4880_b1 , \2161_b1 , \1476_b1 );
not ( \1476_b1 , w_11958 );
and ( \4880_b0 , \2161_b0 , w_11959 );
and ( w_11958 , w_11959 , \1476_b0 );
or ( \4881_b1 , \2028_b1 , \1474_b1 );
not ( \1474_b1 , w_11960 );
and ( \4881_b0 , \2028_b0 , w_11961 );
and ( w_11960 , w_11961 , \1474_b0 );
or ( \4882_b1 , \4880_b1 , w_11963 );
not ( w_11963 , w_11964 );
and ( \4882_b0 , \4880_b0 , w_11965 );
and ( w_11964 ,  , w_11965 );
buf ( w_11963 , \4881_b1 );
not ( w_11963 , w_11966 );
not (  , w_11967 );
and ( w_11966 , w_11967 , \4881_b0 );
or ( \4883_b1 , \4882_b1 , w_11968 );
xor ( \4883_b0 , \4882_b0 , w_11970 );
not ( w_11970 , w_11971 );
and ( w_11971 , w_11968 , w_11969 );
buf ( w_11968 , \1363_b1 );
not ( w_11968 , w_11972 );
not ( w_11969 , w_11973 );
and ( w_11972 , w_11973 , \1363_b0 );
or ( \4884_b1 , \2532_b1 , \1280_b1 );
not ( \1280_b1 , w_11974 );
and ( \4884_b0 , \2532_b0 , w_11975 );
and ( w_11974 , w_11975 , \1280_b0 );
or ( \4885_b1 , \2305_b1 , \1278_b1 );
not ( \1278_b1 , w_11976 );
and ( \4885_b0 , \2305_b0 , w_11977 );
and ( w_11976 , w_11977 , \1278_b0 );
or ( \4886_b1 , \4884_b1 , w_11979 );
not ( w_11979 , w_11980 );
and ( \4886_b0 , \4884_b0 , w_11981 );
and ( w_11980 ,  , w_11981 );
buf ( w_11979 , \4885_b1 );
not ( w_11979 , w_11982 );
not (  , w_11983 );
and ( w_11982 , w_11983 , \4885_b0 );
or ( \4887_b1 , \4886_b1 , w_11984 );
xor ( \4887_b0 , \4886_b0 , w_11986 );
not ( w_11986 , w_11987 );
and ( w_11987 , w_11984 , w_11985 );
buf ( w_11984 , \1177_b1 );
not ( w_11984 , w_11988 );
not ( w_11985 , w_11989 );
and ( w_11988 , w_11989 , \1177_b0 );
or ( \4888_b1 , \4883_b1 , \4887_b1 );
not ( \4887_b1 , w_11990 );
and ( \4888_b0 , \4883_b0 , w_11991 );
and ( w_11990 , w_11991 , \4887_b0 );
or ( \4889_b1 , \2763_b1 , \1062_b1 );
not ( \1062_b1 , w_11992 );
and ( \4889_b0 , \2763_b0 , w_11993 );
and ( w_11992 , w_11993 , \1062_b0 );
or ( \4890_b1 , \2541_b1 , \1060_b1 );
not ( \1060_b1 , w_11994 );
and ( \4890_b0 , \2541_b0 , w_11995 );
and ( w_11994 , w_11995 , \1060_b0 );
or ( \4891_b1 , \4889_b1 , w_11997 );
not ( w_11997 , w_11998 );
and ( \4891_b0 , \4889_b0 , w_11999 );
and ( w_11998 ,  , w_11999 );
buf ( w_11997 , \4890_b1 );
not ( w_11997 , w_12000 );
not (  , w_12001 );
and ( w_12000 , w_12001 , \4890_b0 );
or ( \4892_b1 , \4891_b1 , w_12002 );
xor ( \4892_b0 , \4891_b0 , w_12004 );
not ( w_12004 , w_12005 );
and ( w_12005 , w_12002 , w_12003 );
buf ( w_12002 , \984_b1 );
not ( w_12002 , w_12006 );
not ( w_12003 , w_12007 );
and ( w_12006 , w_12007 , \984_b0 );
or ( \4893_b1 , \4887_b1 , \4892_b1 );
not ( \4892_b1 , w_12008 );
and ( \4893_b0 , \4887_b0 , w_12009 );
and ( w_12008 , w_12009 , \4892_b0 );
or ( \4894_b1 , \4883_b1 , \4892_b1 );
not ( \4892_b1 , w_12010 );
and ( \4894_b0 , \4883_b0 , w_12011 );
and ( w_12010 , w_12011 , \4892_b0 );
or ( \4896_b1 , \4878_b1 , \4895_b1 );
not ( \4895_b1 , w_12012 );
and ( \4896_b0 , \4878_b0 , w_12013 );
and ( w_12012 , w_12013 , \4895_b0 );
or ( \4897_b1 , \4866_b1 , \4895_b1 );
not ( \4895_b1 , w_12014 );
and ( \4897_b0 , \4866_b0 , w_12015 );
and ( w_12014 , w_12015 , \4895_b0 );
or ( \4899_b1 , \4766_b1 , \4770_b1 );
xor ( \4899_b0 , \4766_b0 , w_12016 );
not ( w_12016 , w_12017 );
and ( w_12017 , \4770_b1 , \4770_b0 );
or ( \4900_b1 , \4899_b1 , \4775_b1 );
xor ( \4900_b0 , \4899_b0 , w_12018 );
not ( w_12018 , w_12019 );
and ( w_12019 , \4775_b1 , \4775_b0 );
or ( \4901_b1 , \4782_b1 , \4786_b1 );
xor ( \4901_b0 , \4782_b0 , w_12020 );
not ( w_12020 , w_12021 );
and ( w_12021 , \4786_b1 , \4786_b0 );
or ( \4902_b1 , \4901_b1 , \4791_b1 );
xor ( \4902_b0 , \4901_b0 , w_12022 );
not ( w_12022 , w_12023 );
and ( w_12023 , \4791_b1 , \4791_b0 );
or ( \4903_b1 , \4900_b1 , \4902_b1 );
not ( \4902_b1 , w_12024 );
and ( \4903_b0 , \4900_b0 , w_12025 );
and ( w_12024 , w_12025 , \4902_b0 );
or ( \4904_b1 , \4799_b1 , \4803_b1 );
xor ( \4904_b0 , \4799_b0 , w_12026 );
not ( w_12026 , w_12027 );
and ( w_12027 , \4803_b1 , \4803_b0 );
or ( \4905_b1 , \4904_b1 , \4808_b1 );
xor ( \4905_b0 , \4904_b0 , w_12028 );
not ( w_12028 , w_12029 );
and ( w_12029 , \4808_b1 , \4808_b0 );
or ( \4906_b1 , \4902_b1 , \4905_b1 );
not ( \4905_b1 , w_12030 );
and ( \4906_b0 , \4902_b0 , w_12031 );
and ( w_12030 , w_12031 , \4905_b0 );
or ( \4907_b1 , \4900_b1 , \4905_b1 );
not ( \4905_b1 , w_12032 );
and ( \4907_b0 , \4900_b0 , w_12033 );
and ( w_12032 , w_12033 , \4905_b0 );
or ( \4909_b1 , \4898_b1 , \4908_b1 );
not ( \4908_b1 , w_12034 );
and ( \4909_b0 , \4898_b0 , w_12035 );
and ( w_12034 , w_12035 , \4908_b0 );
or ( \4910_b1 , \4703_b1 , \4707_b1 );
xor ( \4910_b0 , \4703_b0 , w_12036 );
not ( w_12036 , w_12037 );
and ( w_12037 , \4707_b1 , \4707_b0 );
or ( \4911_b1 , \4910_b1 , \4712_b1 );
xor ( \4911_b0 , \4910_b0 , w_12038 );
not ( w_12038 , w_12039 );
and ( w_12039 , \4712_b1 , \4712_b0 );
or ( \4912_b1 , \4908_b1 , \4911_b1 );
not ( \4911_b1 , w_12040 );
and ( \4912_b0 , \4908_b0 , w_12041 );
and ( w_12040 , w_12041 , \4911_b0 );
or ( \4913_b1 , \4898_b1 , \4911_b1 );
not ( \4911_b1 , w_12042 );
and ( \4913_b0 , \4898_b0 , w_12043 );
and ( w_12042 , w_12043 , \4911_b0 );
or ( \4915_b1 , \4674_b1 , \4678_b1 );
xor ( \4915_b0 , \4674_b0 , w_12044 );
not ( w_12044 , w_12045 );
and ( w_12045 , \4678_b1 , \4678_b0 );
or ( \4916_b1 , \4915_b1 , \668_b1 );
xor ( \4916_b0 , \4915_b0 , w_12046 );
not ( w_12046 , w_12047 );
and ( w_12047 , \668_b1 , \668_b0 );
or ( \4917_b1 , \4778_b1 , \4794_b1 );
xor ( \4917_b0 , \4778_b0 , w_12048 );
not ( w_12048 , w_12049 );
and ( w_12049 , \4794_b1 , \4794_b0 );
or ( \4918_b1 , \4917_b1 , \4811_b1 );
xor ( \4918_b0 , \4917_b0 , w_12050 );
not ( w_12050 , w_12051 );
and ( w_12051 , \4811_b1 , \4811_b0 );
or ( \4919_b1 , \4916_b1 , \4918_b1 );
not ( \4918_b1 , w_12052 );
and ( \4919_b0 , \4916_b0 , w_12053 );
and ( w_12052 , w_12053 , \4918_b0 );
or ( \4920_b1 , \4818_b1 , \4820_b1 );
xor ( \4920_b0 , \4818_b0 , w_12054 );
not ( w_12054 , w_12055 );
and ( w_12055 , \4820_b1 , \4820_b0 );
or ( \4921_b1 , \4920_b1 , \4823_b1 );
xor ( \4921_b0 , \4920_b0 , w_12056 );
not ( w_12056 , w_12057 );
and ( w_12057 , \4823_b1 , \4823_b0 );
or ( \4922_b1 , \4918_b1 , \4921_b1 );
not ( \4921_b1 , w_12058 );
and ( \4922_b0 , \4918_b0 , w_12059 );
and ( w_12058 , w_12059 , \4921_b0 );
or ( \4923_b1 , \4916_b1 , \4921_b1 );
not ( \4921_b1 , w_12060 );
and ( \4923_b0 , \4916_b0 , w_12061 );
and ( w_12060 , w_12061 , \4921_b0 );
or ( \4925_b1 , \4914_b1 , \4924_b1 );
not ( \4924_b1 , w_12062 );
and ( \4925_b0 , \4914_b0 , w_12063 );
and ( w_12062 , w_12063 , \4924_b0 );
or ( \4926_b1 , \4722_b1 , \4724_b1 );
xor ( \4926_b0 , \4722_b0 , w_12064 );
not ( w_12064 , w_12065 );
and ( w_12065 , \4724_b1 , \4724_b0 );
or ( \4927_b1 , \4926_b1 , \4727_b1 );
xor ( \4927_b0 , \4926_b0 , w_12066 );
not ( w_12066 , w_12067 );
and ( w_12067 , \4727_b1 , \4727_b0 );
or ( \4928_b1 , \4924_b1 , \4927_b1 );
not ( \4927_b1 , w_12068 );
and ( \4928_b0 , \4924_b0 , w_12069 );
and ( w_12068 , w_12069 , \4927_b0 );
or ( \4929_b1 , \4914_b1 , \4927_b1 );
not ( \4927_b1 , w_12070 );
and ( \4929_b0 , \4914_b0 , w_12071 );
and ( w_12070 , w_12071 , \4927_b0 );
or ( \4931_b1 , \4682_b1 , \4698_b1 );
xor ( \4931_b0 , \4682_b0 , w_12072 );
not ( w_12072 , w_12073 );
and ( w_12073 , \4698_b1 , \4698_b0 );
or ( \4932_b1 , \4931_b1 , \4715_b1 );
xor ( \4932_b0 , \4931_b0 , w_12074 );
not ( w_12074 , w_12075 );
and ( w_12075 , \4715_b1 , \4715_b0 );
or ( \4933_b1 , \4814_b1 , \4826_b1 );
xor ( \4933_b0 , \4814_b0 , w_12076 );
not ( w_12076 , w_12077 );
and ( w_12077 , \4826_b1 , \4826_b0 );
or ( \4934_b1 , \4933_b1 , \4829_b1 );
xor ( \4934_b0 , \4933_b0 , w_12078 );
not ( w_12078 , w_12079 );
and ( w_12079 , \4829_b1 , \4829_b0 );
or ( \4935_b1 , \4932_b1 , \4934_b1 );
not ( \4934_b1 , w_12080 );
and ( \4935_b0 , \4932_b0 , w_12081 );
and ( w_12080 , w_12081 , \4934_b0 );
or ( \4936_b1 , \4930_b1 , \4935_b1 );
not ( \4935_b1 , w_12082 );
and ( \4936_b0 , \4930_b0 , w_12083 );
and ( w_12082 , w_12083 , \4935_b0 );
or ( \4937_b1 , \4832_b1 , \4834_b1 );
xor ( \4937_b0 , \4832_b0 , w_12084 );
not ( w_12084 , w_12085 );
and ( w_12085 , \4834_b1 , \4834_b0 );
or ( \4938_b1 , \4937_b1 , \4836_b1 );
xor ( \4938_b0 , \4937_b0 , w_12086 );
not ( w_12086 , w_12087 );
and ( w_12087 , \4836_b1 , \4836_b0 );
or ( \4939_b1 , \4935_b1 , \4938_b1 );
not ( \4938_b1 , w_12088 );
and ( \4939_b0 , \4935_b0 , w_12089 );
and ( w_12088 , w_12089 , \4938_b0 );
or ( \4940_b1 , \4930_b1 , \4938_b1 );
not ( \4938_b1 , w_12090 );
and ( \4940_b0 , \4930_b0 , w_12091 );
and ( w_12090 , w_12091 , \4938_b0 );
or ( \4942_b1 , \4850_b1 , \4941_b1 );
not ( \4941_b1 , w_12092 );
and ( \4942_b0 , \4850_b0 , w_12093 );
and ( w_12092 , w_12093 , \4941_b0 );
or ( \4943_b1 , \4850_b1 , \4941_b1 );
xor ( \4943_b0 , \4850_b0 , w_12094 );
not ( w_12094 , w_12095 );
and ( w_12095 , \4941_b1 , \4941_b0 );
or ( \4944_b1 , \4930_b1 , \4935_b1 );
xor ( \4944_b0 , \4930_b0 , w_12096 );
not ( w_12096 , w_12097 );
and ( w_12097 , \4935_b1 , \4935_b0 );
or ( \4945_b1 , \4944_b1 , \4938_b1 );
xor ( \4945_b0 , \4944_b0 , w_12098 );
not ( w_12098 , w_12099 );
and ( w_12099 , \4938_b1 , \4938_b0 );
or ( \4946_b1 , \1194_b1 , \2913_b1 );
not ( \2913_b1 , w_12100 );
and ( \4946_b0 , \1194_b0 , w_12101 );
and ( w_12100 , w_12101 , \2913_b0 );
or ( \4947_b1 , \1104_b1 , \2910_b1 );
not ( \2910_b1 , w_12102 );
and ( \4947_b0 , \1104_b0 , w_12103 );
and ( w_12102 , w_12103 , \2910_b0 );
or ( \4948_b1 , \4946_b1 , w_12105 );
not ( w_12105 , w_12106 );
and ( \4948_b0 , \4946_b0 , w_12107 );
and ( w_12106 ,  , w_12107 );
buf ( w_12105 , \4947_b1 );
not ( w_12105 , w_12108 );
not (  , w_12109 );
and ( w_12108 , w_12109 , \4947_b0 );
or ( \4949_b1 , \4948_b1 , w_12110 );
xor ( \4949_b0 , \4948_b0 , w_12112 );
not ( w_12112 , w_12113 );
and ( w_12113 , w_12110 , w_12111 );
buf ( w_12110 , \2371_b1 );
not ( w_12110 , w_12114 );
not ( w_12111 , w_12115 );
and ( w_12114 , w_12115 , \2371_b0 );
or ( \4950_b1 , \1304_b1 , \2550_b1 );
not ( \2550_b1 , w_12116 );
and ( \4950_b0 , \1304_b0 , w_12117 );
and ( w_12116 , w_12117 , \2550_b0 );
or ( \4951_b1 , \1299_b1 , \2548_b1 );
not ( \2548_b1 , w_12118 );
and ( \4951_b0 , \1299_b0 , w_12119 );
and ( w_12118 , w_12119 , \2548_b0 );
or ( \4952_b1 , \4950_b1 , w_12121 );
not ( w_12121 , w_12122 );
and ( \4952_b0 , \4950_b0 , w_12123 );
and ( w_12122 ,  , w_12123 );
buf ( w_12121 , \4951_b1 );
not ( w_12121 , w_12124 );
not (  , w_12125 );
and ( w_12124 , w_12125 , \4951_b0 );
or ( \4953_b1 , \4952_b1 , w_12126 );
xor ( \4953_b0 , \4952_b0 , w_12128 );
not ( w_12128 , w_12129 );
and ( w_12129 , w_12126 , w_12127 );
buf ( w_12126 , \2374_b1 );
not ( w_12126 , w_12130 );
not ( w_12127 , w_12131 );
and ( w_12130 , w_12131 , \2374_b0 );
or ( \4954_b1 , \4949_b1 , \4953_b1 );
not ( \4953_b1 , w_12132 );
and ( \4954_b0 , \4949_b0 , w_12133 );
and ( w_12132 , w_12133 , \4953_b0 );
or ( \4955_b1 , \1537_b1 , \2261_b1 );
not ( \2261_b1 , w_12134 );
and ( \4955_b0 , \1537_b0 , w_12135 );
and ( w_12134 , w_12135 , \2261_b0 );
or ( \4956_b1 , \1422_b1 , \2259_b1 );
not ( \2259_b1 , w_12136 );
and ( \4956_b0 , \1422_b0 , w_12137 );
and ( w_12136 , w_12137 , \2259_b0 );
or ( \4957_b1 , \4955_b1 , w_12139 );
not ( w_12139 , w_12140 );
and ( \4957_b0 , \4955_b0 , w_12141 );
and ( w_12140 ,  , w_12141 );
buf ( w_12139 , \4956_b1 );
not ( w_12139 , w_12142 );
not (  , w_12143 );
and ( w_12142 , w_12143 , \4956_b0 );
or ( \4958_b1 , \4957_b1 , w_12144 );
xor ( \4958_b0 , \4957_b0 , w_12146 );
not ( w_12146 , w_12147 );
and ( w_12147 , w_12144 , w_12145 );
buf ( w_12144 , \2124_b1 );
not ( w_12144 , w_12148 );
not ( w_12145 , w_12149 );
and ( w_12148 , w_12149 , \2124_b0 );
or ( \4959_b1 , \4953_b1 , \4958_b1 );
not ( \4958_b1 , w_12150 );
and ( \4959_b0 , \4953_b0 , w_12151 );
and ( w_12150 , w_12151 , \4958_b0 );
or ( \4960_b1 , \4949_b1 , \4958_b1 );
not ( \4958_b1 , w_12152 );
and ( \4960_b0 , \4949_b0 , w_12153 );
and ( w_12152 , w_12153 , \4958_b0 );
or ( \4962_b1 , \1778_b1 , \1955_b1 );
not ( \1955_b1 , w_12154 );
and ( \4962_b0 , \1778_b0 , w_12155 );
and ( w_12154 , w_12155 , \1955_b0 );
or ( \4963_b1 , \1770_b1 , \1953_b1 );
not ( \1953_b1 , w_12156 );
and ( \4963_b0 , \1770_b0 , w_12157 );
and ( w_12156 , w_12157 , \1953_b0 );
or ( \4964_b1 , \4962_b1 , w_12159 );
not ( w_12159 , w_12160 );
and ( \4964_b0 , \4962_b0 , w_12161 );
and ( w_12160 ,  , w_12161 );
buf ( w_12159 , \4963_b1 );
not ( w_12159 , w_12162 );
not (  , w_12163 );
and ( w_12162 , w_12163 , \4963_b0 );
or ( \4965_b1 , \4964_b1 , w_12164 );
xor ( \4965_b0 , \4964_b0 , w_12166 );
not ( w_12166 , w_12167 );
and ( w_12167 , w_12164 , w_12165 );
buf ( w_12164 , \1835_b1 );
not ( w_12164 , w_12168 );
not ( w_12165 , w_12169 );
and ( w_12168 , w_12169 , \1835_b0 );
or ( \4966_b1 , \2028_b1 , \1742_b1 );
not ( \1742_b1 , w_12170 );
and ( \4966_b0 , \2028_b0 , w_12171 );
and ( w_12170 , w_12171 , \1742_b0 );
or ( \4967_b1 , \2023_b1 , \1740_b1 );
not ( \1740_b1 , w_12172 );
and ( \4967_b0 , \2023_b0 , w_12173 );
and ( w_12172 , w_12173 , \1740_b0 );
or ( \4968_b1 , \4966_b1 , w_12175 );
not ( w_12175 , w_12176 );
and ( \4968_b0 , \4966_b0 , w_12177 );
and ( w_12176 ,  , w_12177 );
buf ( w_12175 , \4967_b1 );
not ( w_12175 , w_12178 );
not (  , w_12179 );
and ( w_12178 , w_12179 , \4967_b0 );
or ( \4969_b1 , \4968_b1 , w_12180 );
xor ( \4969_b0 , \4968_b0 , w_12182 );
not ( w_12182 , w_12183 );
and ( w_12183 , w_12180 , w_12181 );
buf ( w_12180 , \1610_b1 );
not ( w_12180 , w_12184 );
not ( w_12181 , w_12185 );
and ( w_12184 , w_12185 , \1610_b0 );
or ( \4970_b1 , \4965_b1 , \4969_b1 );
not ( \4969_b1 , w_12186 );
and ( \4970_b0 , \4965_b0 , w_12187 );
and ( w_12186 , w_12187 , \4969_b0 );
or ( \4971_b1 , \2305_b1 , \1476_b1 );
not ( \1476_b1 , w_12188 );
and ( \4971_b0 , \2305_b0 , w_12189 );
and ( w_12188 , w_12189 , \1476_b0 );
or ( \4972_b1 , \2161_b1 , \1474_b1 );
not ( \1474_b1 , w_12190 );
and ( \4972_b0 , \2161_b0 , w_12191 );
and ( w_12190 , w_12191 , \1474_b0 );
or ( \4973_b1 , \4971_b1 , w_12193 );
not ( w_12193 , w_12194 );
and ( \4973_b0 , \4971_b0 , w_12195 );
and ( w_12194 ,  , w_12195 );
buf ( w_12193 , \4972_b1 );
not ( w_12193 , w_12196 );
not (  , w_12197 );
and ( w_12196 , w_12197 , \4972_b0 );
or ( \4974_b1 , \4973_b1 , w_12198 );
xor ( \4974_b0 , \4973_b0 , w_12200 );
not ( w_12200 , w_12201 );
and ( w_12201 , w_12198 , w_12199 );
buf ( w_12198 , \1363_b1 );
not ( w_12198 , w_12202 );
not ( w_12199 , w_12203 );
and ( w_12202 , w_12203 , \1363_b0 );
or ( \4975_b1 , \4969_b1 , \4974_b1 );
not ( \4974_b1 , w_12204 );
and ( \4975_b0 , \4969_b0 , w_12205 );
and ( w_12204 , w_12205 , \4974_b0 );
or ( \4976_b1 , \4965_b1 , \4974_b1 );
not ( \4974_b1 , w_12206 );
and ( \4976_b0 , \4965_b0 , w_12207 );
and ( w_12206 , w_12207 , \4974_b0 );
or ( \4978_b1 , \4961_b1 , \4977_b1 );
not ( \4977_b1 , w_12208 );
and ( \4978_b0 , \4961_b0 , w_12209 );
and ( w_12208 , w_12209 , \4977_b0 );
or ( \4979_b1 , \2541_b1 , \1280_b1 );
not ( \1280_b1 , w_12210 );
and ( \4979_b0 , \2541_b0 , w_12211 );
and ( w_12210 , w_12211 , \1280_b0 );
or ( \4980_b1 , \2532_b1 , \1278_b1 );
not ( \1278_b1 , w_12212 );
and ( \4980_b0 , \2532_b0 , w_12213 );
and ( w_12212 , w_12213 , \1278_b0 );
or ( \4981_b1 , \4979_b1 , w_12215 );
not ( w_12215 , w_12216 );
and ( \4981_b0 , \4979_b0 , w_12217 );
and ( w_12216 ,  , w_12217 );
buf ( w_12215 , \4980_b1 );
not ( w_12215 , w_12218 );
not (  , w_12219 );
and ( w_12218 , w_12219 , \4980_b0 );
or ( \4982_b1 , \4981_b1 , w_12220 );
xor ( \4982_b0 , \4981_b0 , w_12222 );
not ( w_12222 , w_12223 );
and ( w_12223 , w_12220 , w_12221 );
buf ( w_12220 , \1177_b1 );
not ( w_12220 , w_12224 );
not ( w_12221 , w_12225 );
and ( w_12224 , w_12225 , \1177_b0 );
or ( \4983_b1 , \2850_b1 , \1062_b1 );
not ( \1062_b1 , w_12226 );
and ( \4983_b0 , \2850_b0 , w_12227 );
and ( w_12226 , w_12227 , \1062_b0 );
or ( \4984_b1 , \2763_b1 , \1060_b1 );
not ( \1060_b1 , w_12228 );
and ( \4984_b0 , \2763_b0 , w_12229 );
and ( w_12228 , w_12229 , \1060_b0 );
or ( \4985_b1 , \4983_b1 , w_12231 );
not ( w_12231 , w_12232 );
and ( \4985_b0 , \4983_b0 , w_12233 );
and ( w_12232 ,  , w_12233 );
buf ( w_12231 , \4984_b1 );
not ( w_12231 , w_12234 );
not (  , w_12235 );
and ( w_12234 , w_12235 , \4984_b0 );
or ( \4986_b1 , \4985_b1 , w_12236 );
xor ( \4986_b0 , \4985_b0 , w_12238 );
not ( w_12238 , w_12239 );
and ( w_12239 , w_12236 , w_12237 );
buf ( w_12236 , \984_b1 );
not ( w_12236 , w_12240 );
not ( w_12237 , w_12241 );
and ( w_12240 , w_12241 , \984_b0 );
or ( \4987_b1 , \4982_b1 , \4986_b1 );
not ( \4986_b1 , w_12242 );
and ( \4987_b0 , \4982_b0 , w_12243 );
and ( w_12242 , w_12243 , \4986_b0 );
or ( \4988_b1 , \4977_b1 , \4987_b1 );
not ( \4987_b1 , w_12244 );
and ( \4988_b0 , \4977_b0 , w_12245 );
and ( w_12244 , w_12245 , \4987_b0 );
or ( \4989_b1 , \4961_b1 , \4987_b1 );
not ( \4987_b1 , w_12246 );
and ( \4989_b0 , \4961_b0 , w_12247 );
and ( w_12246 , w_12247 , \4987_b0 );
or ( \4991_b1 , \2850_b1 , w_12249 );
not ( w_12249 , w_12250 );
and ( \4991_b0 , \2850_b0 , w_12251 );
and ( w_12250 ,  , w_12251 );
buf ( w_12249 , \910_b1 );
not ( w_12249 , w_12252 );
not (  , w_12253 );
and ( w_12252 , w_12253 , \910_b0 );
or ( \4992_b1 , \4991_b1 , w_12254 );
xor ( \4992_b0 , \4991_b0 , w_12256 );
not ( w_12256 , w_12257 );
and ( w_12257 , w_12254 , w_12255 );
buf ( w_12254 , \818_b1 );
not ( w_12254 , w_12258 );
not ( w_12255 , w_12259 );
and ( w_12258 , w_12259 , \818_b0 );
or ( \4993_b1 , \4854_b1 , \4858_b1 );
xor ( \4993_b0 , \4854_b0 , w_12260 );
not ( w_12260 , w_12261 );
and ( w_12261 , \4858_b1 , \4858_b0 );
or ( \4994_b1 , \4993_b1 , \4863_b1 );
xor ( \4994_b0 , \4993_b0 , w_12262 );
not ( w_12262 , w_12263 );
and ( w_12263 , \4863_b1 , \4863_b0 );
or ( \4995_b1 , \4992_b1 , \4994_b1 );
not ( \4994_b1 , w_12264 );
and ( \4995_b0 , \4992_b0 , w_12265 );
and ( w_12264 , w_12265 , \4994_b0 );
or ( \4996_b1 , \4883_b1 , \4887_b1 );
xor ( \4996_b0 , \4883_b0 , w_12266 );
not ( w_12266 , w_12267 );
and ( w_12267 , \4887_b1 , \4887_b0 );
or ( \4997_b1 , \4996_b1 , \4892_b1 );
xor ( \4997_b0 , \4996_b0 , w_12268 );
not ( w_12268 , w_12269 );
and ( w_12269 , \4892_b1 , \4892_b0 );
or ( \4998_b1 , \4994_b1 , \4997_b1 );
not ( \4997_b1 , w_12270 );
and ( \4998_b0 , \4994_b0 , w_12271 );
and ( w_12270 , w_12271 , \4997_b0 );
or ( \4999_b1 , \4992_b1 , \4997_b1 );
not ( \4997_b1 , w_12272 );
and ( \4999_b0 , \4992_b0 , w_12273 );
and ( w_12272 , w_12273 , \4997_b0 );
or ( \5001_b1 , \4990_b1 , \5000_b1 );
not ( \5000_b1 , w_12274 );
and ( \5001_b0 , \4990_b0 , w_12275 );
and ( w_12274 , w_12275 , \5000_b0 );
or ( \5002_b1 , \4900_b1 , \4902_b1 );
xor ( \5002_b0 , \4900_b0 , w_12276 );
not ( w_12276 , w_12277 );
and ( w_12277 , \4902_b1 , \4902_b0 );
or ( \5003_b1 , \5002_b1 , \4905_b1 );
xor ( \5003_b0 , \5002_b0 , w_12278 );
not ( w_12278 , w_12279 );
and ( w_12279 , \4905_b1 , \4905_b0 );
or ( \5004_b1 , \5000_b1 , \5003_b1 );
not ( \5003_b1 , w_12280 );
and ( \5004_b0 , \5000_b0 , w_12281 );
and ( w_12280 , w_12281 , \5003_b0 );
or ( \5005_b1 , \4990_b1 , \5003_b1 );
not ( \5003_b1 , w_12282 );
and ( \5005_b0 , \4990_b0 , w_12283 );
and ( w_12282 , w_12283 , \5003_b0 );
or ( \5007_b1 , \4898_b1 , \4908_b1 );
xor ( \5007_b0 , \4898_b0 , w_12284 );
not ( w_12284 , w_12285 );
and ( w_12285 , \4908_b1 , \4908_b0 );
or ( \5008_b1 , \5007_b1 , \4911_b1 );
xor ( \5008_b0 , \5007_b0 , w_12286 );
not ( w_12286 , w_12287 );
and ( w_12287 , \4911_b1 , \4911_b0 );
or ( \5009_b1 , \5006_b1 , \5008_b1 );
not ( \5008_b1 , w_12288 );
and ( \5009_b0 , \5006_b0 , w_12289 );
and ( w_12288 , w_12289 , \5008_b0 );
or ( \5010_b1 , \4916_b1 , \4918_b1 );
xor ( \5010_b0 , \4916_b0 , w_12290 );
not ( w_12290 , w_12291 );
and ( w_12291 , \4918_b1 , \4918_b0 );
or ( \5011_b1 , \5010_b1 , \4921_b1 );
xor ( \5011_b0 , \5010_b0 , w_12292 );
not ( w_12292 , w_12293 );
and ( w_12293 , \4921_b1 , \4921_b0 );
or ( \5012_b1 , \5008_b1 , \5011_b1 );
not ( \5011_b1 , w_12294 );
and ( \5012_b0 , \5008_b0 , w_12295 );
and ( w_12294 , w_12295 , \5011_b0 );
or ( \5013_b1 , \5006_b1 , \5011_b1 );
not ( \5011_b1 , w_12296 );
and ( \5013_b0 , \5006_b0 , w_12297 );
and ( w_12296 , w_12297 , \5011_b0 );
or ( \5015_b1 , \4914_b1 , \4924_b1 );
xor ( \5015_b0 , \4914_b0 , w_12298 );
not ( w_12298 , w_12299 );
and ( w_12299 , \4924_b1 , \4924_b0 );
or ( \5016_b1 , \5015_b1 , \4927_b1 );
xor ( \5016_b0 , \5015_b0 , w_12300 );
not ( w_12300 , w_12301 );
and ( w_12301 , \4927_b1 , \4927_b0 );
or ( \5017_b1 , \5014_b1 , \5016_b1 );
not ( \5016_b1 , w_12302 );
and ( \5017_b0 , \5014_b0 , w_12303 );
and ( w_12302 , w_12303 , \5016_b0 );
or ( \5018_b1 , \4932_b1 , \4934_b1 );
xor ( \5018_b0 , \4932_b0 , w_12304 );
not ( w_12304 , w_12305 );
and ( w_12305 , \4934_b1 , \4934_b0 );
or ( \5019_b1 , \5016_b1 , \5018_b1 );
not ( \5018_b1 , w_12306 );
and ( \5019_b0 , \5016_b0 , w_12307 );
and ( w_12306 , w_12307 , \5018_b0 );
or ( \5020_b1 , \5014_b1 , \5018_b1 );
not ( \5018_b1 , w_12308 );
and ( \5020_b0 , \5014_b0 , w_12309 );
and ( w_12308 , w_12309 , \5018_b0 );
or ( \5022_b1 , \4945_b1 , \5021_b1 );
not ( \5021_b1 , w_12310 );
and ( \5022_b0 , \4945_b0 , w_12311 );
and ( w_12310 , w_12311 , \5021_b0 );
or ( \5023_b1 , \4945_b1 , \5021_b1 );
xor ( \5023_b0 , \4945_b0 , w_12312 );
not ( w_12312 , w_12313 );
and ( w_12313 , \5021_b1 , \5021_b0 );
or ( \5024_b1 , \5014_b1 , \5016_b1 );
xor ( \5024_b0 , \5014_b0 , w_12314 );
not ( w_12314 , w_12315 );
and ( w_12315 , \5016_b1 , \5016_b0 );
or ( \5025_b1 , \5024_b1 , \5018_b1 );
xor ( \5025_b0 , \5024_b0 , w_12316 );
not ( w_12316 , w_12317 );
and ( w_12317 , \5018_b1 , \5018_b0 );
or ( \5026_b1 , \2532_b1 , \1476_b1 );
not ( \1476_b1 , w_12318 );
and ( \5026_b0 , \2532_b0 , w_12319 );
and ( w_12318 , w_12319 , \1476_b0 );
or ( \5027_b1 , \2305_b1 , \1474_b1 );
not ( \1474_b1 , w_12320 );
and ( \5027_b0 , \2305_b0 , w_12321 );
and ( w_12320 , w_12321 , \1474_b0 );
or ( \5028_b1 , \5026_b1 , w_12323 );
not ( w_12323 , w_12324 );
and ( \5028_b0 , \5026_b0 , w_12325 );
and ( w_12324 ,  , w_12325 );
buf ( w_12323 , \5027_b1 );
not ( w_12323 , w_12326 );
not (  , w_12327 );
and ( w_12326 , w_12327 , \5027_b0 );
or ( \5029_b1 , \5028_b1 , w_12328 );
xor ( \5029_b0 , \5028_b0 , w_12330 );
not ( w_12330 , w_12331 );
and ( w_12331 , w_12328 , w_12329 );
buf ( w_12328 , \1363_b1 );
not ( w_12328 , w_12332 );
not ( w_12329 , w_12333 );
and ( w_12332 , w_12333 , \1363_b0 );
or ( \5030_b1 , \2763_b1 , \1280_b1 );
not ( \1280_b1 , w_12334 );
and ( \5030_b0 , \2763_b0 , w_12335 );
and ( w_12334 , w_12335 , \1280_b0 );
or ( \5031_b1 , \2541_b1 , \1278_b1 );
not ( \1278_b1 , w_12336 );
and ( \5031_b0 , \2541_b0 , w_12337 );
and ( w_12336 , w_12337 , \1278_b0 );
or ( \5032_b1 , \5030_b1 , w_12339 );
not ( w_12339 , w_12340 );
and ( \5032_b0 , \5030_b0 , w_12341 );
and ( w_12340 ,  , w_12341 );
buf ( w_12339 , \5031_b1 );
not ( w_12339 , w_12342 );
not (  , w_12343 );
and ( w_12342 , w_12343 , \5031_b0 );
or ( \5033_b1 , \5032_b1 , w_12344 );
xor ( \5033_b0 , \5032_b0 , w_12346 );
not ( w_12346 , w_12347 );
and ( w_12347 , w_12344 , w_12345 );
buf ( w_12344 , \1177_b1 );
not ( w_12344 , w_12348 );
not ( w_12345 , w_12349 );
and ( w_12348 , w_12349 , \1177_b0 );
or ( \5034_b1 , \5029_b1 , \5033_b1 );
not ( \5033_b1 , w_12350 );
and ( \5034_b0 , \5029_b0 , w_12351 );
and ( w_12350 , w_12351 , \5033_b0 );
or ( \5035_b1 , \2850_b1 , w_12353 );
not ( w_12353 , w_12354 );
and ( \5035_b0 , \2850_b0 , w_12355 );
and ( w_12354 ,  , w_12355 );
buf ( w_12353 , \1060_b1 );
not ( w_12353 , w_12356 );
not (  , w_12357 );
and ( w_12356 , w_12357 , \1060_b0 );
or ( \5036_b1 , \5035_b1 , w_12358 );
xor ( \5036_b0 , \5035_b0 , w_12360 );
not ( w_12360 , w_12361 );
and ( w_12361 , w_12358 , w_12359 );
buf ( w_12358 , \984_b1 );
not ( w_12358 , w_12362 );
not ( w_12359 , w_12363 );
and ( w_12362 , w_12363 , \984_b0 );
or ( \5037_b1 , \5033_b1 , \5036_b1 );
not ( \5036_b1 , w_12364 );
and ( \5037_b0 , \5033_b0 , w_12365 );
and ( w_12364 , w_12365 , \5036_b0 );
or ( \5038_b1 , \5029_b1 , \5036_b1 );
not ( \5036_b1 , w_12366 );
and ( \5038_b0 , \5029_b0 , w_12367 );
and ( w_12366 , w_12367 , \5036_b0 );
or ( \5040_b1 , \1299_b1 , \2913_b1 );
not ( \2913_b1 , w_12368 );
and ( \5040_b0 , \1299_b0 , w_12369 );
and ( w_12368 , w_12369 , \2913_b0 );
or ( \5041_b1 , \1194_b1 , \2910_b1 );
not ( \2910_b1 , w_12370 );
and ( \5041_b0 , \1194_b0 , w_12371 );
and ( w_12370 , w_12371 , \2910_b0 );
or ( \5042_b1 , \5040_b1 , w_12373 );
not ( w_12373 , w_12374 );
and ( \5042_b0 , \5040_b0 , w_12375 );
and ( w_12374 ,  , w_12375 );
buf ( w_12373 , \5041_b1 );
not ( w_12373 , w_12376 );
not (  , w_12377 );
and ( w_12376 , w_12377 , \5041_b0 );
or ( \5043_b1 , \5042_b1 , w_12378 );
xor ( \5043_b0 , \5042_b0 , w_12380 );
not ( w_12380 , w_12381 );
and ( w_12381 , w_12378 , w_12379 );
buf ( w_12378 , \2371_b1 );
not ( w_12378 , w_12382 );
not ( w_12379 , w_12383 );
and ( w_12382 , w_12383 , \2371_b0 );
or ( \5044_b1 , \1422_b1 , \2550_b1 );
not ( \2550_b1 , w_12384 );
and ( \5044_b0 , \1422_b0 , w_12385 );
and ( w_12384 , w_12385 , \2550_b0 );
or ( \5045_b1 , \1304_b1 , \2548_b1 );
not ( \2548_b1 , w_12386 );
and ( \5045_b0 , \1304_b0 , w_12387 );
and ( w_12386 , w_12387 , \2548_b0 );
or ( \5046_b1 , \5044_b1 , w_12389 );
not ( w_12389 , w_12390 );
and ( \5046_b0 , \5044_b0 , w_12391 );
and ( w_12390 ,  , w_12391 );
buf ( w_12389 , \5045_b1 );
not ( w_12389 , w_12392 );
not (  , w_12393 );
and ( w_12392 , w_12393 , \5045_b0 );
or ( \5047_b1 , \5046_b1 , w_12394 );
xor ( \5047_b0 , \5046_b0 , w_12396 );
not ( w_12396 , w_12397 );
and ( w_12397 , w_12394 , w_12395 );
buf ( w_12394 , \2374_b1 );
not ( w_12394 , w_12398 );
not ( w_12395 , w_12399 );
and ( w_12398 , w_12399 , \2374_b0 );
or ( \5048_b1 , \5043_b1 , \5047_b1 );
not ( \5047_b1 , w_12400 );
and ( \5048_b0 , \5043_b0 , w_12401 );
and ( w_12400 , w_12401 , \5047_b0 );
or ( \5049_b1 , \5047_b1 , \984_b1 );
not ( \984_b1 , w_12402 );
and ( \5049_b0 , \5047_b0 , w_12403 );
and ( w_12402 , w_12403 , \984_b0 );
or ( \5050_b1 , \5043_b1 , \984_b1 );
not ( \984_b1 , w_12404 );
and ( \5050_b0 , \5043_b0 , w_12405 );
and ( w_12404 , w_12405 , \984_b0 );
or ( \5052_b1 , \5039_b1 , \5051_b1 );
not ( \5051_b1 , w_12406 );
and ( \5052_b0 , \5039_b0 , w_12407 );
and ( w_12406 , w_12407 , \5051_b0 );
or ( \5053_b1 , \1770_b1 , \2261_b1 );
not ( \2261_b1 , w_12408 );
and ( \5053_b0 , \1770_b0 , w_12409 );
and ( w_12408 , w_12409 , \2261_b0 );
or ( \5054_b1 , \1537_b1 , \2259_b1 );
not ( \2259_b1 , w_12410 );
and ( \5054_b0 , \1537_b0 , w_12411 );
and ( w_12410 , w_12411 , \2259_b0 );
or ( \5055_b1 , \5053_b1 , w_12413 );
not ( w_12413 , w_12414 );
and ( \5055_b0 , \5053_b0 , w_12415 );
and ( w_12414 ,  , w_12415 );
buf ( w_12413 , \5054_b1 );
not ( w_12413 , w_12416 );
not (  , w_12417 );
and ( w_12416 , w_12417 , \5054_b0 );
or ( \5056_b1 , \5055_b1 , w_12418 );
xor ( \5056_b0 , \5055_b0 , w_12420 );
not ( w_12420 , w_12421 );
and ( w_12421 , w_12418 , w_12419 );
buf ( w_12418 , \2124_b1 );
not ( w_12418 , w_12422 );
not ( w_12419 , w_12423 );
and ( w_12422 , w_12423 , \2124_b0 );
or ( \5057_b1 , \2023_b1 , \1955_b1 );
not ( \1955_b1 , w_12424 );
and ( \5057_b0 , \2023_b0 , w_12425 );
and ( w_12424 , w_12425 , \1955_b0 );
or ( \5058_b1 , \1778_b1 , \1953_b1 );
not ( \1953_b1 , w_12426 );
and ( \5058_b0 , \1778_b0 , w_12427 );
and ( w_12426 , w_12427 , \1953_b0 );
or ( \5059_b1 , \5057_b1 , w_12429 );
not ( w_12429 , w_12430 );
and ( \5059_b0 , \5057_b0 , w_12431 );
and ( w_12430 ,  , w_12431 );
buf ( w_12429 , \5058_b1 );
not ( w_12429 , w_12432 );
not (  , w_12433 );
and ( w_12432 , w_12433 , \5058_b0 );
or ( \5060_b1 , \5059_b1 , w_12434 );
xor ( \5060_b0 , \5059_b0 , w_12436 );
not ( w_12436 , w_12437 );
and ( w_12437 , w_12434 , w_12435 );
buf ( w_12434 , \1835_b1 );
not ( w_12434 , w_12438 );
not ( w_12435 , w_12439 );
and ( w_12438 , w_12439 , \1835_b0 );
or ( \5061_b1 , \5056_b1 , \5060_b1 );
not ( \5060_b1 , w_12440 );
and ( \5061_b0 , \5056_b0 , w_12441 );
and ( w_12440 , w_12441 , \5060_b0 );
or ( \5062_b1 , \2161_b1 , \1742_b1 );
not ( \1742_b1 , w_12442 );
and ( \5062_b0 , \2161_b0 , w_12443 );
and ( w_12442 , w_12443 , \1742_b0 );
or ( \5063_b1 , \2028_b1 , \1740_b1 );
not ( \1740_b1 , w_12444 );
and ( \5063_b0 , \2028_b0 , w_12445 );
and ( w_12444 , w_12445 , \1740_b0 );
or ( \5064_b1 , \5062_b1 , w_12447 );
not ( w_12447 , w_12448 );
and ( \5064_b0 , \5062_b0 , w_12449 );
and ( w_12448 ,  , w_12449 );
buf ( w_12447 , \5063_b1 );
not ( w_12447 , w_12450 );
not (  , w_12451 );
and ( w_12450 , w_12451 , \5063_b0 );
or ( \5065_b1 , \5064_b1 , w_12452 );
xor ( \5065_b0 , \5064_b0 , w_12454 );
not ( w_12454 , w_12455 );
and ( w_12455 , w_12452 , w_12453 );
buf ( w_12452 , \1610_b1 );
not ( w_12452 , w_12456 );
not ( w_12453 , w_12457 );
and ( w_12456 , w_12457 , \1610_b0 );
or ( \5066_b1 , \5060_b1 , \5065_b1 );
not ( \5065_b1 , w_12458 );
and ( \5066_b0 , \5060_b0 , w_12459 );
and ( w_12458 , w_12459 , \5065_b0 );
or ( \5067_b1 , \5056_b1 , \5065_b1 );
not ( \5065_b1 , w_12460 );
and ( \5067_b0 , \5056_b0 , w_12461 );
and ( w_12460 , w_12461 , \5065_b0 );
or ( \5069_b1 , \5051_b1 , \5068_b1 );
not ( \5068_b1 , w_12462 );
and ( \5069_b0 , \5051_b0 , w_12463 );
and ( w_12462 , w_12463 , \5068_b0 );
or ( \5070_b1 , \5039_b1 , \5068_b1 );
not ( \5068_b1 , w_12464 );
and ( \5070_b0 , \5039_b0 , w_12465 );
and ( w_12464 , w_12465 , \5068_b0 );
or ( \5072_b1 , \4949_b1 , \4953_b1 );
xor ( \5072_b0 , \4949_b0 , w_12466 );
not ( w_12466 , w_12467 );
and ( w_12467 , \4953_b1 , \4953_b0 );
or ( \5073_b1 , \5072_b1 , \4958_b1 );
xor ( \5073_b0 , \5072_b0 , w_12468 );
not ( w_12468 , w_12469 );
and ( w_12469 , \4958_b1 , \4958_b0 );
or ( \5074_b1 , \4965_b1 , \4969_b1 );
xor ( \5074_b0 , \4965_b0 , w_12470 );
not ( w_12470 , w_12471 );
and ( w_12471 , \4969_b1 , \4969_b0 );
or ( \5075_b1 , \5074_b1 , \4974_b1 );
xor ( \5075_b0 , \5074_b0 , w_12472 );
not ( w_12472 , w_12473 );
and ( w_12473 , \4974_b1 , \4974_b0 );
or ( \5076_b1 , \5073_b1 , \5075_b1 );
not ( \5075_b1 , w_12474 );
and ( \5076_b0 , \5073_b0 , w_12475 );
and ( w_12474 , w_12475 , \5075_b0 );
or ( \5077_b1 , \4982_b1 , \4986_b1 );
xor ( \5077_b0 , \4982_b0 , w_12476 );
not ( w_12476 , w_12477 );
and ( w_12477 , \4986_b1 , \4986_b0 );
or ( \5078_b1 , \5075_b1 , \5077_b1 );
not ( \5077_b1 , w_12478 );
and ( \5078_b0 , \5075_b0 , w_12479 );
and ( w_12478 , w_12479 , \5077_b0 );
or ( \5079_b1 , \5073_b1 , \5077_b1 );
not ( \5077_b1 , w_12480 );
and ( \5079_b0 , \5073_b0 , w_12481 );
and ( w_12480 , w_12481 , \5077_b0 );
or ( \5081_b1 , \5071_b1 , \5080_b1 );
not ( \5080_b1 , w_12482 );
and ( \5081_b0 , \5071_b0 , w_12483 );
and ( w_12482 , w_12483 , \5080_b0 );
or ( \5082_b1 , \4870_b1 , \4874_b1 );
xor ( \5082_b0 , \4870_b0 , w_12484 );
not ( w_12484 , w_12485 );
and ( w_12485 , \4874_b1 , \4874_b0 );
or ( \5083_b1 , \5082_b1 , \818_b1 );
xor ( \5083_b0 , \5082_b0 , w_12486 );
not ( w_12486 , w_12487 );
and ( w_12487 , \818_b1 , \818_b0 );
or ( \5084_b1 , \5080_b1 , \5083_b1 );
not ( \5083_b1 , w_12488 );
and ( \5084_b0 , \5080_b0 , w_12489 );
and ( w_12488 , w_12489 , \5083_b0 );
or ( \5085_b1 , \5071_b1 , \5083_b1 );
not ( \5083_b1 , w_12490 );
and ( \5085_b0 , \5071_b0 , w_12491 );
and ( w_12490 , w_12491 , \5083_b0 );
or ( \5087_b1 , \4961_b1 , \4977_b1 );
xor ( \5087_b0 , \4961_b0 , w_12492 );
not ( w_12492 , w_12493 );
and ( w_12493 , \4977_b1 , \4977_b0 );
or ( \5088_b1 , \5087_b1 , \4987_b1 );
xor ( \5088_b0 , \5087_b0 , w_12494 );
not ( w_12494 , w_12495 );
and ( w_12495 , \4987_b1 , \4987_b0 );
or ( \5089_b1 , \4992_b1 , \4994_b1 );
xor ( \5089_b0 , \4992_b0 , w_12496 );
not ( w_12496 , w_12497 );
and ( w_12497 , \4994_b1 , \4994_b0 );
or ( \5090_b1 , \5089_b1 , \4997_b1 );
xor ( \5090_b0 , \5089_b0 , w_12498 );
not ( w_12498 , w_12499 );
and ( w_12499 , \4997_b1 , \4997_b0 );
or ( \5091_b1 , \5088_b1 , \5090_b1 );
not ( \5090_b1 , w_12500 );
and ( \5091_b0 , \5088_b0 , w_12501 );
and ( w_12500 , w_12501 , \5090_b0 );
or ( \5092_b1 , \5086_b1 , \5091_b1 );
not ( \5091_b1 , w_12502 );
and ( \5092_b0 , \5086_b0 , w_12503 );
and ( w_12502 , w_12503 , \5091_b0 );
or ( \5093_b1 , \4866_b1 , \4878_b1 );
xor ( \5093_b0 , \4866_b0 , w_12504 );
not ( w_12504 , w_12505 );
and ( w_12505 , \4878_b1 , \4878_b0 );
or ( \5094_b1 , \5093_b1 , \4895_b1 );
xor ( \5094_b0 , \5093_b0 , w_12506 );
not ( w_12506 , w_12507 );
and ( w_12507 , \4895_b1 , \4895_b0 );
or ( \5095_b1 , \5091_b1 , \5094_b1 );
not ( \5094_b1 , w_12508 );
and ( \5095_b0 , \5091_b0 , w_12509 );
and ( w_12508 , w_12509 , \5094_b0 );
or ( \5096_b1 , \5086_b1 , \5094_b1 );
not ( \5094_b1 , w_12510 );
and ( \5096_b0 , \5086_b0 , w_12511 );
and ( w_12510 , w_12511 , \5094_b0 );
or ( \5098_b1 , \5006_b1 , \5008_b1 );
xor ( \5098_b0 , \5006_b0 , w_12512 );
not ( w_12512 , w_12513 );
and ( w_12513 , \5008_b1 , \5008_b0 );
or ( \5099_b1 , \5098_b1 , \5011_b1 );
xor ( \5099_b0 , \5098_b0 , w_12514 );
not ( w_12514 , w_12515 );
and ( w_12515 , \5011_b1 , \5011_b0 );
or ( \5100_b1 , \5097_b1 , \5099_b1 );
not ( \5099_b1 , w_12516 );
and ( \5100_b0 , \5097_b0 , w_12517 );
and ( w_12516 , w_12517 , \5099_b0 );
or ( \5101_b1 , \5025_b1 , \5100_b1 );
not ( \5100_b1 , w_12518 );
and ( \5101_b0 , \5025_b0 , w_12519 );
and ( w_12518 , w_12519 , \5100_b0 );
or ( \5102_b1 , \5025_b1 , \5100_b1 );
xor ( \5102_b0 , \5025_b0 , w_12520 );
not ( w_12520 , w_12521 );
and ( w_12521 , \5100_b1 , \5100_b0 );
or ( \5103_b1 , \5097_b1 , \5099_b1 );
xor ( \5103_b0 , \5097_b0 , w_12522 );
not ( w_12522 , w_12523 );
and ( w_12523 , \5099_b1 , \5099_b0 );
or ( \5104_b1 , \5086_b1 , \5091_b1 );
xor ( \5104_b0 , \5086_b0 , w_12524 );
not ( w_12524 , w_12525 );
and ( w_12525 , \5091_b1 , \5091_b0 );
or ( \5105_b1 , \5104_b1 , \5094_b1 );
xor ( \5105_b0 , \5104_b0 , w_12526 );
not ( w_12526 , w_12527 );
and ( w_12527 , \5094_b1 , \5094_b0 );
or ( \5106_b1 , \4990_b1 , \5000_b1 );
xor ( \5106_b0 , \4990_b0 , w_12528 );
not ( w_12528 , w_12529 );
and ( w_12529 , \5000_b1 , \5000_b0 );
or ( \5107_b1 , \5106_b1 , \5003_b1 );
xor ( \5107_b0 , \5106_b0 , w_12530 );
not ( w_12530 , w_12531 );
and ( w_12531 , \5003_b1 , \5003_b0 );
or ( \5108_b1 , \5105_b1 , \5107_b1 );
not ( \5107_b1 , w_12532 );
and ( \5108_b0 , \5105_b0 , w_12533 );
and ( w_12532 , w_12533 , \5107_b0 );
or ( \5109_b1 , \5103_b1 , \5108_b1 );
not ( \5108_b1 , w_12534 );
and ( \5109_b0 , \5103_b0 , w_12535 );
and ( w_12534 , w_12535 , \5108_b0 );
or ( \5110_b1 , \5103_b1 , \5108_b1 );
xor ( \5110_b0 , \5103_b0 , w_12536 );
not ( w_12536 , w_12537 );
and ( w_12537 , \5108_b1 , \5108_b0 );
or ( \5111_b1 , \5105_b1 , \5107_b1 );
xor ( \5111_b0 , \5105_b0 , w_12538 );
not ( w_12538 , w_12539 );
and ( w_12539 , \5107_b1 , \5107_b0 );
or ( \5112_b1 , \1304_b1 , \2913_b1 );
not ( \2913_b1 , w_12540 );
and ( \5112_b0 , \1304_b0 , w_12541 );
and ( w_12540 , w_12541 , \2913_b0 );
or ( \5113_b1 , \1299_b1 , \2910_b1 );
not ( \2910_b1 , w_12542 );
and ( \5113_b0 , \1299_b0 , w_12543 );
and ( w_12542 , w_12543 , \2910_b0 );
or ( \5114_b1 , \5112_b1 , w_12545 );
not ( w_12545 , w_12546 );
and ( \5114_b0 , \5112_b0 , w_12547 );
and ( w_12546 ,  , w_12547 );
buf ( w_12545 , \5113_b1 );
not ( w_12545 , w_12548 );
not (  , w_12549 );
and ( w_12548 , w_12549 , \5113_b0 );
or ( \5115_b1 , \5114_b1 , w_12550 );
xor ( \5115_b0 , \5114_b0 , w_12552 );
not ( w_12552 , w_12553 );
and ( w_12553 , w_12550 , w_12551 );
buf ( w_12550 , \2371_b1 );
not ( w_12550 , w_12554 );
not ( w_12551 , w_12555 );
and ( w_12554 , w_12555 , \2371_b0 );
or ( \5116_b1 , \1537_b1 , \2550_b1 );
not ( \2550_b1 , w_12556 );
and ( \5116_b0 , \1537_b0 , w_12557 );
and ( w_12556 , w_12557 , \2550_b0 );
or ( \5117_b1 , \1422_b1 , \2548_b1 );
not ( \2548_b1 , w_12558 );
and ( \5117_b0 , \1422_b0 , w_12559 );
and ( w_12558 , w_12559 , \2548_b0 );
or ( \5118_b1 , \5116_b1 , w_12561 );
not ( w_12561 , w_12562 );
and ( \5118_b0 , \5116_b0 , w_12563 );
and ( w_12562 ,  , w_12563 );
buf ( w_12561 , \5117_b1 );
not ( w_12561 , w_12564 );
not (  , w_12565 );
and ( w_12564 , w_12565 , \5117_b0 );
or ( \5119_b1 , \5118_b1 , w_12566 );
xor ( \5119_b0 , \5118_b0 , w_12568 );
not ( w_12568 , w_12569 );
and ( w_12569 , w_12566 , w_12567 );
buf ( w_12566 , \2374_b1 );
not ( w_12566 , w_12570 );
not ( w_12567 , w_12571 );
and ( w_12570 , w_12571 , \2374_b0 );
or ( \5120_b1 , \5115_b1 , \5119_b1 );
not ( \5119_b1 , w_12572 );
and ( \5120_b0 , \5115_b0 , w_12573 );
and ( w_12572 , w_12573 , \5119_b0 );
or ( \5121_b1 , \1778_b1 , \2261_b1 );
not ( \2261_b1 , w_12574 );
and ( \5121_b0 , \1778_b0 , w_12575 );
and ( w_12574 , w_12575 , \2261_b0 );
or ( \5122_b1 , \1770_b1 , \2259_b1 );
not ( \2259_b1 , w_12576 );
and ( \5122_b0 , \1770_b0 , w_12577 );
and ( w_12576 , w_12577 , \2259_b0 );
or ( \5123_b1 , \5121_b1 , w_12579 );
not ( w_12579 , w_12580 );
and ( \5123_b0 , \5121_b0 , w_12581 );
and ( w_12580 ,  , w_12581 );
buf ( w_12579 , \5122_b1 );
not ( w_12579 , w_12582 );
not (  , w_12583 );
and ( w_12582 , w_12583 , \5122_b0 );
or ( \5124_b1 , \5123_b1 , w_12584 );
xor ( \5124_b0 , \5123_b0 , w_12586 );
not ( w_12586 , w_12587 );
and ( w_12587 , w_12584 , w_12585 );
buf ( w_12584 , \2124_b1 );
not ( w_12584 , w_12588 );
not ( w_12585 , w_12589 );
and ( w_12588 , w_12589 , \2124_b0 );
or ( \5125_b1 , \5119_b1 , \5124_b1 );
not ( \5124_b1 , w_12590 );
and ( \5125_b0 , \5119_b0 , w_12591 );
and ( w_12590 , w_12591 , \5124_b0 );
or ( \5126_b1 , \5115_b1 , \5124_b1 );
not ( \5124_b1 , w_12592 );
and ( \5126_b0 , \5115_b0 , w_12593 );
and ( w_12592 , w_12593 , \5124_b0 );
or ( \5128_b1 , \2028_b1 , \1955_b1 );
not ( \1955_b1 , w_12594 );
and ( \5128_b0 , \2028_b0 , w_12595 );
and ( w_12594 , w_12595 , \1955_b0 );
or ( \5129_b1 , \2023_b1 , \1953_b1 );
not ( \1953_b1 , w_12596 );
and ( \5129_b0 , \2023_b0 , w_12597 );
and ( w_12596 , w_12597 , \1953_b0 );
or ( \5130_b1 , \5128_b1 , w_12599 );
not ( w_12599 , w_12600 );
and ( \5130_b0 , \5128_b0 , w_12601 );
and ( w_12600 ,  , w_12601 );
buf ( w_12599 , \5129_b1 );
not ( w_12599 , w_12602 );
not (  , w_12603 );
and ( w_12602 , w_12603 , \5129_b0 );
or ( \5131_b1 , \5130_b1 , w_12604 );
xor ( \5131_b0 , \5130_b0 , w_12606 );
not ( w_12606 , w_12607 );
and ( w_12607 , w_12604 , w_12605 );
buf ( w_12604 , \1835_b1 );
not ( w_12604 , w_12608 );
not ( w_12605 , w_12609 );
and ( w_12608 , w_12609 , \1835_b0 );
or ( \5132_b1 , \2305_b1 , \1742_b1 );
not ( \1742_b1 , w_12610 );
and ( \5132_b0 , \2305_b0 , w_12611 );
and ( w_12610 , w_12611 , \1742_b0 );
or ( \5133_b1 , \2161_b1 , \1740_b1 );
not ( \1740_b1 , w_12612 );
and ( \5133_b0 , \2161_b0 , w_12613 );
and ( w_12612 , w_12613 , \1740_b0 );
or ( \5134_b1 , \5132_b1 , w_12615 );
not ( w_12615 , w_12616 );
and ( \5134_b0 , \5132_b0 , w_12617 );
and ( w_12616 ,  , w_12617 );
buf ( w_12615 , \5133_b1 );
not ( w_12615 , w_12618 );
not (  , w_12619 );
and ( w_12618 , w_12619 , \5133_b0 );
or ( \5135_b1 , \5134_b1 , w_12620 );
xor ( \5135_b0 , \5134_b0 , w_12622 );
not ( w_12622 , w_12623 );
and ( w_12623 , w_12620 , w_12621 );
buf ( w_12620 , \1610_b1 );
not ( w_12620 , w_12624 );
not ( w_12621 , w_12625 );
and ( w_12624 , w_12625 , \1610_b0 );
or ( \5136_b1 , \5131_b1 , \5135_b1 );
not ( \5135_b1 , w_12626 );
and ( \5136_b0 , \5131_b0 , w_12627 );
and ( w_12626 , w_12627 , \5135_b0 );
or ( \5137_b1 , \2541_b1 , \1476_b1 );
not ( \1476_b1 , w_12628 );
and ( \5137_b0 , \2541_b0 , w_12629 );
and ( w_12628 , w_12629 , \1476_b0 );
or ( \5138_b1 , \2532_b1 , \1474_b1 );
not ( \1474_b1 , w_12630 );
and ( \5138_b0 , \2532_b0 , w_12631 );
and ( w_12630 , w_12631 , \1474_b0 );
or ( \5139_b1 , \5137_b1 , w_12633 );
not ( w_12633 , w_12634 );
and ( \5139_b0 , \5137_b0 , w_12635 );
and ( w_12634 ,  , w_12635 );
buf ( w_12633 , \5138_b1 );
not ( w_12633 , w_12636 );
not (  , w_12637 );
and ( w_12636 , w_12637 , \5138_b0 );
or ( \5140_b1 , \5139_b1 , w_12638 );
xor ( \5140_b0 , \5139_b0 , w_12640 );
not ( w_12640 , w_12641 );
and ( w_12641 , w_12638 , w_12639 );
buf ( w_12638 , \1363_b1 );
not ( w_12638 , w_12642 );
not ( w_12639 , w_12643 );
and ( w_12642 , w_12643 , \1363_b0 );
or ( \5141_b1 , \5135_b1 , \5140_b1 );
not ( \5140_b1 , w_12644 );
and ( \5141_b0 , \5135_b0 , w_12645 );
and ( w_12644 , w_12645 , \5140_b0 );
or ( \5142_b1 , \5131_b1 , \5140_b1 );
not ( \5140_b1 , w_12646 );
and ( \5142_b0 , \5131_b0 , w_12647 );
and ( w_12646 , w_12647 , \5140_b0 );
or ( \5144_b1 , \5127_b1 , \5143_b1 );
not ( \5143_b1 , w_12648 );
and ( \5144_b0 , \5127_b0 , w_12649 );
and ( w_12648 , w_12649 , \5143_b0 );
or ( \5145_b1 , \5029_b1 , \5033_b1 );
xor ( \5145_b0 , \5029_b0 , w_12650 );
not ( w_12650 , w_12651 );
and ( w_12651 , \5033_b1 , \5033_b0 );
or ( \5146_b1 , \5145_b1 , \5036_b1 );
xor ( \5146_b0 , \5145_b0 , w_12652 );
not ( w_12652 , w_12653 );
and ( w_12653 , \5036_b1 , \5036_b0 );
or ( \5147_b1 , \5143_b1 , \5146_b1 );
not ( \5146_b1 , w_12654 );
and ( \5147_b0 , \5143_b0 , w_12655 );
and ( w_12654 , w_12655 , \5146_b0 );
or ( \5148_b1 , \5127_b1 , \5146_b1 );
not ( \5146_b1 , w_12656 );
and ( \5148_b0 , \5127_b0 , w_12657 );
and ( w_12656 , w_12657 , \5146_b0 );
or ( \5150_b1 , \5043_b1 , \5047_b1 );
xor ( \5150_b0 , \5043_b0 , w_12658 );
not ( w_12658 , w_12659 );
and ( w_12659 , \5047_b1 , \5047_b0 );
or ( \5151_b1 , \5150_b1 , \984_b1 );
xor ( \5151_b0 , \5150_b0 , w_12660 );
not ( w_12660 , w_12661 );
and ( w_12661 , \984_b1 , \984_b0 );
or ( \5152_b1 , \5056_b1 , \5060_b1 );
xor ( \5152_b0 , \5056_b0 , w_12662 );
not ( w_12662 , w_12663 );
and ( w_12663 , \5060_b1 , \5060_b0 );
or ( \5153_b1 , \5152_b1 , \5065_b1 );
xor ( \5153_b0 , \5152_b0 , w_12664 );
not ( w_12664 , w_12665 );
and ( w_12665 , \5065_b1 , \5065_b0 );
or ( \5154_b1 , \5151_b1 , \5153_b1 );
not ( \5153_b1 , w_12666 );
and ( \5154_b0 , \5151_b0 , w_12667 );
and ( w_12666 , w_12667 , \5153_b0 );
or ( \5155_b1 , \5149_b1 , \5154_b1 );
not ( \5154_b1 , w_12668 );
and ( \5155_b0 , \5149_b0 , w_12669 );
and ( w_12668 , w_12669 , \5154_b0 );
or ( \5156_b1 , \5073_b1 , \5075_b1 );
xor ( \5156_b0 , \5073_b0 , w_12670 );
not ( w_12670 , w_12671 );
and ( w_12671 , \5075_b1 , \5075_b0 );
or ( \5157_b1 , \5156_b1 , \5077_b1 );
xor ( \5157_b0 , \5156_b0 , w_12672 );
not ( w_12672 , w_12673 );
and ( w_12673 , \5077_b1 , \5077_b0 );
or ( \5158_b1 , \5154_b1 , \5157_b1 );
not ( \5157_b1 , w_12674 );
and ( \5158_b0 , \5154_b0 , w_12675 );
and ( w_12674 , w_12675 , \5157_b0 );
or ( \5159_b1 , \5149_b1 , \5157_b1 );
not ( \5157_b1 , w_12676 );
and ( \5159_b0 , \5149_b0 , w_12677 );
and ( w_12676 , w_12677 , \5157_b0 );
or ( \5161_b1 , \5071_b1 , \5080_b1 );
xor ( \5161_b0 , \5071_b0 , w_12678 );
not ( w_12678 , w_12679 );
and ( w_12679 , \5080_b1 , \5080_b0 );
or ( \5162_b1 , \5161_b1 , \5083_b1 );
xor ( \5162_b0 , \5161_b0 , w_12680 );
not ( w_12680 , w_12681 );
and ( w_12681 , \5083_b1 , \5083_b0 );
or ( \5163_b1 , \5160_b1 , \5162_b1 );
not ( \5162_b1 , w_12682 );
and ( \5163_b0 , \5160_b0 , w_12683 );
and ( w_12682 , w_12683 , \5162_b0 );
or ( \5164_b1 , \5088_b1 , \5090_b1 );
xor ( \5164_b0 , \5088_b0 , w_12684 );
not ( w_12684 , w_12685 );
and ( w_12685 , \5090_b1 , \5090_b0 );
or ( \5165_b1 , \5162_b1 , \5164_b1 );
not ( \5164_b1 , w_12686 );
and ( \5165_b0 , \5162_b0 , w_12687 );
and ( w_12686 , w_12687 , \5164_b0 );
or ( \5166_b1 , \5160_b1 , \5164_b1 );
not ( \5164_b1 , w_12688 );
and ( \5166_b0 , \5160_b0 , w_12689 );
and ( w_12688 , w_12689 , \5164_b0 );
or ( \5168_b1 , \5111_b1 , \5167_b1 );
not ( \5167_b1 , w_12690 );
and ( \5168_b0 , \5111_b0 , w_12691 );
and ( w_12690 , w_12691 , \5167_b0 );
or ( \5169_b1 , \5111_b1 , \5167_b1 );
xor ( \5169_b0 , \5111_b0 , w_12692 );
not ( w_12692 , w_12693 );
and ( w_12693 , \5167_b1 , \5167_b0 );
or ( \5170_b1 , \5160_b1 , \5162_b1 );
xor ( \5170_b0 , \5160_b0 , w_12694 );
not ( w_12694 , w_12695 );
and ( w_12695 , \5162_b1 , \5162_b0 );
or ( \5171_b1 , \5170_b1 , \5164_b1 );
xor ( \5171_b0 , \5170_b0 , w_12696 );
not ( w_12696 , w_12697 );
and ( w_12697 , \5164_b1 , \5164_b0 );
or ( \5172_b1 , \1422_b1 , \2913_b1 );
not ( \2913_b1 , w_12698 );
and ( \5172_b0 , \1422_b0 , w_12699 );
and ( w_12698 , w_12699 , \2913_b0 );
or ( \5173_b1 , \1304_b1 , \2910_b1 );
not ( \2910_b1 , w_12700 );
and ( \5173_b0 , \1304_b0 , w_12701 );
and ( w_12700 , w_12701 , \2910_b0 );
or ( \5174_b1 , \5172_b1 , w_12703 );
not ( w_12703 , w_12704 );
and ( \5174_b0 , \5172_b0 , w_12705 );
and ( w_12704 ,  , w_12705 );
buf ( w_12703 , \5173_b1 );
not ( w_12703 , w_12706 );
not (  , w_12707 );
and ( w_12706 , w_12707 , \5173_b0 );
or ( \5175_b1 , \5174_b1 , w_12708 );
xor ( \5175_b0 , \5174_b0 , w_12710 );
not ( w_12710 , w_12711 );
and ( w_12711 , w_12708 , w_12709 );
buf ( w_12708 , \2371_b1 );
not ( w_12708 , w_12712 );
not ( w_12709 , w_12713 );
and ( w_12712 , w_12713 , \2371_b0 );
or ( \5176_b1 , \1770_b1 , \2550_b1 );
not ( \2550_b1 , w_12714 );
and ( \5176_b0 , \1770_b0 , w_12715 );
and ( w_12714 , w_12715 , \2550_b0 );
or ( \5177_b1 , \1537_b1 , \2548_b1 );
not ( \2548_b1 , w_12716 );
and ( \5177_b0 , \1537_b0 , w_12717 );
and ( w_12716 , w_12717 , \2548_b0 );
or ( \5178_b1 , \5176_b1 , w_12719 );
not ( w_12719 , w_12720 );
and ( \5178_b0 , \5176_b0 , w_12721 );
and ( w_12720 ,  , w_12721 );
buf ( w_12719 , \5177_b1 );
not ( w_12719 , w_12722 );
not (  , w_12723 );
and ( w_12722 , w_12723 , \5177_b0 );
or ( \5179_b1 , \5178_b1 , w_12724 );
xor ( \5179_b0 , \5178_b0 , w_12726 );
not ( w_12726 , w_12727 );
and ( w_12727 , w_12724 , w_12725 );
buf ( w_12724 , \2374_b1 );
not ( w_12724 , w_12728 );
not ( w_12725 , w_12729 );
and ( w_12728 , w_12729 , \2374_b0 );
or ( \5180_b1 , \5175_b1 , \5179_b1 );
not ( \5179_b1 , w_12730 );
and ( \5180_b0 , \5175_b0 , w_12731 );
and ( w_12730 , w_12731 , \5179_b0 );
or ( \5181_b1 , \5179_b1 , \1177_b1 );
not ( \1177_b1 , w_12732 );
and ( \5181_b0 , \5179_b0 , w_12733 );
and ( w_12732 , w_12733 , \1177_b0 );
or ( \5182_b1 , \5175_b1 , \1177_b1 );
not ( \1177_b1 , w_12734 );
and ( \5182_b0 , \5175_b0 , w_12735 );
and ( w_12734 , w_12735 , \1177_b0 );
or ( \5184_b1 , \2023_b1 , \2261_b1 );
not ( \2261_b1 , w_12736 );
and ( \5184_b0 , \2023_b0 , w_12737 );
and ( w_12736 , w_12737 , \2261_b0 );
or ( \5185_b1 , \1778_b1 , \2259_b1 );
not ( \2259_b1 , w_12738 );
and ( \5185_b0 , \1778_b0 , w_12739 );
and ( w_12738 , w_12739 , \2259_b0 );
or ( \5186_b1 , \5184_b1 , w_12741 );
not ( w_12741 , w_12742 );
and ( \5186_b0 , \5184_b0 , w_12743 );
and ( w_12742 ,  , w_12743 );
buf ( w_12741 , \5185_b1 );
not ( w_12741 , w_12744 );
not (  , w_12745 );
and ( w_12744 , w_12745 , \5185_b0 );
or ( \5187_b1 , \5186_b1 , w_12746 );
xor ( \5187_b0 , \5186_b0 , w_12748 );
not ( w_12748 , w_12749 );
and ( w_12749 , w_12746 , w_12747 );
buf ( w_12746 , \2124_b1 );
not ( w_12746 , w_12750 );
not ( w_12747 , w_12751 );
and ( w_12750 , w_12751 , \2124_b0 );
or ( \5188_b1 , \2161_b1 , \1955_b1 );
not ( \1955_b1 , w_12752 );
and ( \5188_b0 , \2161_b0 , w_12753 );
and ( w_12752 , w_12753 , \1955_b0 );
or ( \5189_b1 , \2028_b1 , \1953_b1 );
not ( \1953_b1 , w_12754 );
and ( \5189_b0 , \2028_b0 , w_12755 );
and ( w_12754 , w_12755 , \1953_b0 );
or ( \5190_b1 , \5188_b1 , w_12757 );
not ( w_12757 , w_12758 );
and ( \5190_b0 , \5188_b0 , w_12759 );
and ( w_12758 ,  , w_12759 );
buf ( w_12757 , \5189_b1 );
not ( w_12757 , w_12760 );
not (  , w_12761 );
and ( w_12760 , w_12761 , \5189_b0 );
or ( \5191_b1 , \5190_b1 , w_12762 );
xor ( \5191_b0 , \5190_b0 , w_12764 );
not ( w_12764 , w_12765 );
and ( w_12765 , w_12762 , w_12763 );
buf ( w_12762 , \1835_b1 );
not ( w_12762 , w_12766 );
not ( w_12763 , w_12767 );
and ( w_12766 , w_12767 , \1835_b0 );
or ( \5192_b1 , \5187_b1 , \5191_b1 );
not ( \5191_b1 , w_12768 );
and ( \5192_b0 , \5187_b0 , w_12769 );
and ( w_12768 , w_12769 , \5191_b0 );
or ( \5193_b1 , \2532_b1 , \1742_b1 );
not ( \1742_b1 , w_12770 );
and ( \5193_b0 , \2532_b0 , w_12771 );
and ( w_12770 , w_12771 , \1742_b0 );
or ( \5194_b1 , \2305_b1 , \1740_b1 );
not ( \1740_b1 , w_12772 );
and ( \5194_b0 , \2305_b0 , w_12773 );
and ( w_12772 , w_12773 , \1740_b0 );
or ( \5195_b1 , \5193_b1 , w_12775 );
not ( w_12775 , w_12776 );
and ( \5195_b0 , \5193_b0 , w_12777 );
and ( w_12776 ,  , w_12777 );
buf ( w_12775 , \5194_b1 );
not ( w_12775 , w_12778 );
not (  , w_12779 );
and ( w_12778 , w_12779 , \5194_b0 );
or ( \5196_b1 , \5195_b1 , w_12780 );
xor ( \5196_b0 , \5195_b0 , w_12782 );
not ( w_12782 , w_12783 );
and ( w_12783 , w_12780 , w_12781 );
buf ( w_12780 , \1610_b1 );
not ( w_12780 , w_12784 );
not ( w_12781 , w_12785 );
and ( w_12784 , w_12785 , \1610_b0 );
or ( \5197_b1 , \5191_b1 , \5196_b1 );
not ( \5196_b1 , w_12786 );
and ( \5197_b0 , \5191_b0 , w_12787 );
and ( w_12786 , w_12787 , \5196_b0 );
or ( \5198_b1 , \5187_b1 , \5196_b1 );
not ( \5196_b1 , w_12788 );
and ( \5198_b0 , \5187_b0 , w_12789 );
and ( w_12788 , w_12789 , \5196_b0 );
or ( \5200_b1 , \5183_b1 , \5199_b1 );
not ( \5199_b1 , w_12790 );
and ( \5200_b0 , \5183_b0 , w_12791 );
and ( w_12790 , w_12791 , \5199_b0 );
or ( \5201_b1 , \2850_b1 , \1280_b1 );
not ( \1280_b1 , w_12792 );
and ( \5201_b0 , \2850_b0 , w_12793 );
and ( w_12792 , w_12793 , \1280_b0 );
or ( \5202_b1 , \2763_b1 , \1278_b1 );
not ( \1278_b1 , w_12794 );
and ( \5202_b0 , \2763_b0 , w_12795 );
and ( w_12794 , w_12795 , \1278_b0 );
or ( \5203_b1 , \5201_b1 , w_12797 );
not ( w_12797 , w_12798 );
and ( \5203_b0 , \5201_b0 , w_12799 );
and ( w_12798 ,  , w_12799 );
buf ( w_12797 , \5202_b1 );
not ( w_12797 , w_12800 );
not (  , w_12801 );
and ( w_12800 , w_12801 , \5202_b0 );
or ( \5204_b1 , \5203_b1 , w_12802 );
xor ( \5204_b0 , \5203_b0 , w_12804 );
not ( w_12804 , w_12805 );
and ( w_12805 , w_12802 , w_12803 );
buf ( w_12802 , \1177_b1 );
not ( w_12802 , w_12806 );
not ( w_12803 , w_12807 );
and ( w_12806 , w_12807 , \1177_b0 );
or ( \5205_b1 , \5199_b1 , \5204_b1 );
not ( \5204_b1 , w_12808 );
and ( \5205_b0 , \5199_b0 , w_12809 );
and ( w_12808 , w_12809 , \5204_b0 );
or ( \5206_b1 , \5183_b1 , \5204_b1 );
not ( \5204_b1 , w_12810 );
and ( \5206_b0 , \5183_b0 , w_12811 );
and ( w_12810 , w_12811 , \5204_b0 );
or ( \5208_b1 , \5127_b1 , \5143_b1 );
xor ( \5208_b0 , \5127_b0 , w_12812 );
not ( w_12812 , w_12813 );
and ( w_12813 , \5143_b1 , \5143_b0 );
or ( \5209_b1 , \5208_b1 , \5146_b1 );
xor ( \5209_b0 , \5208_b0 , w_12814 );
not ( w_12814 , w_12815 );
and ( w_12815 , \5146_b1 , \5146_b0 );
or ( \5210_b1 , \5207_b1 , \5209_b1 );
not ( \5209_b1 , w_12816 );
and ( \5210_b0 , \5207_b0 , w_12817 );
and ( w_12816 , w_12817 , \5209_b0 );
or ( \5211_b1 , \5151_b1 , \5153_b1 );
xor ( \5211_b0 , \5151_b0 , w_12818 );
not ( w_12818 , w_12819 );
and ( w_12819 , \5153_b1 , \5153_b0 );
or ( \5212_b1 , \5209_b1 , \5211_b1 );
not ( \5211_b1 , w_12820 );
and ( \5212_b0 , \5209_b0 , w_12821 );
and ( w_12820 , w_12821 , \5211_b0 );
or ( \5213_b1 , \5207_b1 , \5211_b1 );
not ( \5211_b1 , w_12822 );
and ( \5213_b0 , \5207_b0 , w_12823 );
and ( w_12822 , w_12823 , \5211_b0 );
or ( \5215_b1 , \5039_b1 , \5051_b1 );
xor ( \5215_b0 , \5039_b0 , w_12824 );
not ( w_12824 , w_12825 );
and ( w_12825 , \5051_b1 , \5051_b0 );
or ( \5216_b1 , \5215_b1 , \5068_b1 );
xor ( \5216_b0 , \5215_b0 , w_12826 );
not ( w_12826 , w_12827 );
and ( w_12827 , \5068_b1 , \5068_b0 );
or ( \5217_b1 , \5214_b1 , \5216_b1 );
not ( \5216_b1 , w_12828 );
and ( \5217_b0 , \5214_b0 , w_12829 );
and ( w_12828 , w_12829 , \5216_b0 );
or ( \5218_b1 , \5149_b1 , \5154_b1 );
xor ( \5218_b0 , \5149_b0 , w_12830 );
not ( w_12830 , w_12831 );
and ( w_12831 , \5154_b1 , \5154_b0 );
or ( \5219_b1 , \5218_b1 , \5157_b1 );
xor ( \5219_b0 , \5218_b0 , w_12832 );
not ( w_12832 , w_12833 );
and ( w_12833 , \5157_b1 , \5157_b0 );
or ( \5220_b1 , \5216_b1 , \5219_b1 );
not ( \5219_b1 , w_12834 );
and ( \5220_b0 , \5216_b0 , w_12835 );
and ( w_12834 , w_12835 , \5219_b0 );
or ( \5221_b1 , \5214_b1 , \5219_b1 );
not ( \5219_b1 , w_12836 );
and ( \5221_b0 , \5214_b0 , w_12837 );
and ( w_12836 , w_12837 , \5219_b0 );
or ( \5223_b1 , \5171_b1 , \5222_b1 );
not ( \5222_b1 , w_12838 );
and ( \5223_b0 , \5171_b0 , w_12839 );
and ( w_12838 , w_12839 , \5222_b0 );
or ( \5224_b1 , \5171_b1 , \5222_b1 );
xor ( \5224_b0 , \5171_b0 , w_12840 );
not ( w_12840 , w_12841 );
and ( w_12841 , \5222_b1 , \5222_b0 );
or ( \5225_b1 , \5214_b1 , \5216_b1 );
xor ( \5225_b0 , \5214_b0 , w_12842 );
not ( w_12842 , w_12843 );
and ( w_12843 , \5216_b1 , \5216_b0 );
or ( \5226_b1 , \5225_b1 , \5219_b1 );
xor ( \5226_b0 , \5225_b0 , w_12844 );
not ( w_12844 , w_12845 );
and ( w_12845 , \5219_b1 , \5219_b0 );
or ( \5227_b1 , \2305_b1 , \1955_b1 );
not ( \1955_b1 , w_12846 );
and ( \5227_b0 , \2305_b0 , w_12847 );
and ( w_12846 , w_12847 , \1955_b0 );
or ( \5228_b1 , \2161_b1 , \1953_b1 );
not ( \1953_b1 , w_12848 );
and ( \5228_b0 , \2161_b0 , w_12849 );
and ( w_12848 , w_12849 , \1953_b0 );
or ( \5229_b1 , \5227_b1 , w_12851 );
not ( w_12851 , w_12852 );
and ( \5229_b0 , \5227_b0 , w_12853 );
and ( w_12852 ,  , w_12853 );
buf ( w_12851 , \5228_b1 );
not ( w_12851 , w_12854 );
not (  , w_12855 );
and ( w_12854 , w_12855 , \5228_b0 );
or ( \5230_b1 , \5229_b1 , w_12856 );
xor ( \5230_b0 , \5229_b0 , w_12858 );
not ( w_12858 , w_12859 );
and ( w_12859 , w_12856 , w_12857 );
buf ( w_12856 , \1835_b1 );
not ( w_12856 , w_12860 );
not ( w_12857 , w_12861 );
and ( w_12860 , w_12861 , \1835_b0 );
or ( \5231_b1 , \2541_b1 , \1742_b1 );
not ( \1742_b1 , w_12862 );
and ( \5231_b0 , \2541_b0 , w_12863 );
and ( w_12862 , w_12863 , \1742_b0 );
or ( \5232_b1 , \2532_b1 , \1740_b1 );
not ( \1740_b1 , w_12864 );
and ( \5232_b0 , \2532_b0 , w_12865 );
and ( w_12864 , w_12865 , \1740_b0 );
or ( \5233_b1 , \5231_b1 , w_12867 );
not ( w_12867 , w_12868 );
and ( \5233_b0 , \5231_b0 , w_12869 );
and ( w_12868 ,  , w_12869 );
buf ( w_12867 , \5232_b1 );
not ( w_12867 , w_12870 );
not (  , w_12871 );
and ( w_12870 , w_12871 , \5232_b0 );
or ( \5234_b1 , \5233_b1 , w_12872 );
xor ( \5234_b0 , \5233_b0 , w_12874 );
not ( w_12874 , w_12875 );
and ( w_12875 , w_12872 , w_12873 );
buf ( w_12872 , \1610_b1 );
not ( w_12872 , w_12876 );
not ( w_12873 , w_12877 );
and ( w_12876 , w_12877 , \1610_b0 );
or ( \5235_b1 , \5230_b1 , \5234_b1 );
not ( \5234_b1 , w_12878 );
and ( \5235_b0 , \5230_b0 , w_12879 );
and ( w_12878 , w_12879 , \5234_b0 );
or ( \5236_b1 , \2850_b1 , \1476_b1 );
not ( \1476_b1 , w_12880 );
and ( \5236_b0 , \2850_b0 , w_12881 );
and ( w_12880 , w_12881 , \1476_b0 );
or ( \5237_b1 , \2763_b1 , \1474_b1 );
not ( \1474_b1 , w_12882 );
and ( \5237_b0 , \2763_b0 , w_12883 );
and ( w_12882 , w_12883 , \1474_b0 );
or ( \5238_b1 , \5236_b1 , w_12885 );
not ( w_12885 , w_12886 );
and ( \5238_b0 , \5236_b0 , w_12887 );
and ( w_12886 ,  , w_12887 );
buf ( w_12885 , \5237_b1 );
not ( w_12885 , w_12888 );
not (  , w_12889 );
and ( w_12888 , w_12889 , \5237_b0 );
or ( \5239_b1 , \5238_b1 , w_12890 );
xor ( \5239_b0 , \5238_b0 , w_12892 );
not ( w_12892 , w_12893 );
and ( w_12893 , w_12890 , w_12891 );
buf ( w_12890 , \1363_b1 );
not ( w_12890 , w_12894 );
not ( w_12891 , w_12895 );
and ( w_12894 , w_12895 , \1363_b0 );
or ( \5240_b1 , \5234_b1 , \5239_b1 );
not ( \5239_b1 , w_12896 );
and ( \5240_b0 , \5234_b0 , w_12897 );
and ( w_12896 , w_12897 , \5239_b0 );
or ( \5241_b1 , \5230_b1 , \5239_b1 );
not ( \5239_b1 , w_12898 );
and ( \5241_b0 , \5230_b0 , w_12899 );
and ( w_12898 , w_12899 , \5239_b0 );
or ( \5243_b1 , \1537_b1 , \2913_b1 );
not ( \2913_b1 , w_12900 );
and ( \5243_b0 , \1537_b0 , w_12901 );
and ( w_12900 , w_12901 , \2913_b0 );
or ( \5244_b1 , \1422_b1 , \2910_b1 );
not ( \2910_b1 , w_12902 );
and ( \5244_b0 , \1422_b0 , w_12903 );
and ( w_12902 , w_12903 , \2910_b0 );
or ( \5245_b1 , \5243_b1 , w_12905 );
not ( w_12905 , w_12906 );
and ( \5245_b0 , \5243_b0 , w_12907 );
and ( w_12906 ,  , w_12907 );
buf ( w_12905 , \5244_b1 );
not ( w_12905 , w_12908 );
not (  , w_12909 );
and ( w_12908 , w_12909 , \5244_b0 );
or ( \5246_b1 , \5245_b1 , w_12910 );
xor ( \5246_b0 , \5245_b0 , w_12912 );
not ( w_12912 , w_12913 );
and ( w_12913 , w_12910 , w_12911 );
buf ( w_12910 , \2371_b1 );
not ( w_12910 , w_12914 );
not ( w_12911 , w_12915 );
and ( w_12914 , w_12915 , \2371_b0 );
or ( \5247_b1 , \1778_b1 , \2550_b1 );
not ( \2550_b1 , w_12916 );
and ( \5247_b0 , \1778_b0 , w_12917 );
and ( w_12916 , w_12917 , \2550_b0 );
or ( \5248_b1 , \1770_b1 , \2548_b1 );
not ( \2548_b1 , w_12918 );
and ( \5248_b0 , \1770_b0 , w_12919 );
and ( w_12918 , w_12919 , \2548_b0 );
or ( \5249_b1 , \5247_b1 , w_12921 );
not ( w_12921 , w_12922 );
and ( \5249_b0 , \5247_b0 , w_12923 );
and ( w_12922 ,  , w_12923 );
buf ( w_12921 , \5248_b1 );
not ( w_12921 , w_12924 );
not (  , w_12925 );
and ( w_12924 , w_12925 , \5248_b0 );
or ( \5250_b1 , \5249_b1 , w_12926 );
xor ( \5250_b0 , \5249_b0 , w_12928 );
not ( w_12928 , w_12929 );
and ( w_12929 , w_12926 , w_12927 );
buf ( w_12926 , \2374_b1 );
not ( w_12926 , w_12930 );
not ( w_12927 , w_12931 );
and ( w_12930 , w_12931 , \2374_b0 );
or ( \5251_b1 , \5246_b1 , \5250_b1 );
not ( \5250_b1 , w_12932 );
and ( \5251_b0 , \5246_b0 , w_12933 );
and ( w_12932 , w_12933 , \5250_b0 );
or ( \5252_b1 , \2028_b1 , \2261_b1 );
not ( \2261_b1 , w_12934 );
and ( \5252_b0 , \2028_b0 , w_12935 );
and ( w_12934 , w_12935 , \2261_b0 );
or ( \5253_b1 , \2023_b1 , \2259_b1 );
not ( \2259_b1 , w_12936 );
and ( \5253_b0 , \2023_b0 , w_12937 );
and ( w_12936 , w_12937 , \2259_b0 );
or ( \5254_b1 , \5252_b1 , w_12939 );
not ( w_12939 , w_12940 );
and ( \5254_b0 , \5252_b0 , w_12941 );
and ( w_12940 ,  , w_12941 );
buf ( w_12939 , \5253_b1 );
not ( w_12939 , w_12942 );
not (  , w_12943 );
and ( w_12942 , w_12943 , \5253_b0 );
or ( \5255_b1 , \5254_b1 , w_12944 );
xor ( \5255_b0 , \5254_b0 , w_12946 );
not ( w_12946 , w_12947 );
and ( w_12947 , w_12944 , w_12945 );
buf ( w_12944 , \2124_b1 );
not ( w_12944 , w_12948 );
not ( w_12945 , w_12949 );
and ( w_12948 , w_12949 , \2124_b0 );
or ( \5256_b1 , \5250_b1 , \5255_b1 );
not ( \5255_b1 , w_12950 );
and ( \5256_b0 , \5250_b0 , w_12951 );
and ( w_12950 , w_12951 , \5255_b0 );
or ( \5257_b1 , \5246_b1 , \5255_b1 );
not ( \5255_b1 , w_12952 );
and ( \5257_b0 , \5246_b0 , w_12953 );
and ( w_12952 , w_12953 , \5255_b0 );
or ( \5259_b1 , \5242_b1 , \5258_b1 );
not ( \5258_b1 , w_12954 );
and ( \5259_b0 , \5242_b0 , w_12955 );
and ( w_12954 , w_12955 , \5258_b0 );
or ( \5260_b1 , \2763_b1 , \1476_b1 );
not ( \1476_b1 , w_12956 );
and ( \5260_b0 , \2763_b0 , w_12957 );
and ( w_12956 , w_12957 , \1476_b0 );
or ( \5261_b1 , \2541_b1 , \1474_b1 );
not ( \1474_b1 , w_12958 );
and ( \5261_b0 , \2541_b0 , w_12959 );
and ( w_12958 , w_12959 , \1474_b0 );
or ( \5262_b1 , \5260_b1 , w_12961 );
not ( w_12961 , w_12962 );
and ( \5262_b0 , \5260_b0 , w_12963 );
and ( w_12962 ,  , w_12963 );
buf ( w_12961 , \5261_b1 );
not ( w_12961 , w_12964 );
not (  , w_12965 );
and ( w_12964 , w_12965 , \5261_b0 );
or ( \5263_b1 , \5262_b1 , w_12966 );
xor ( \5263_b0 , \5262_b0 , w_12968 );
not ( w_12968 , w_12969 );
and ( w_12969 , w_12966 , w_12967 );
buf ( w_12966 , \1363_b1 );
not ( w_12966 , w_12970 );
not ( w_12967 , w_12971 );
and ( w_12970 , w_12971 , \1363_b0 );
or ( \5264_b1 , \5258_b1 , \5263_b1 );
not ( \5263_b1 , w_12972 );
and ( \5264_b0 , \5258_b0 , w_12973 );
and ( w_12972 , w_12973 , \5263_b0 );
or ( \5265_b1 , \5242_b1 , \5263_b1 );
not ( \5263_b1 , w_12974 );
and ( \5265_b0 , \5242_b0 , w_12975 );
and ( w_12974 , w_12975 , \5263_b0 );
or ( \5267_b1 , \2850_b1 , w_12977 );
not ( w_12977 , w_12978 );
and ( \5267_b0 , \2850_b0 , w_12979 );
and ( w_12978 ,  , w_12979 );
buf ( w_12977 , \1278_b1 );
not ( w_12977 , w_12980 );
not (  , w_12981 );
and ( w_12980 , w_12981 , \1278_b0 );
or ( \5268_b1 , \5267_b1 , w_12982 );
xor ( \5268_b0 , \5267_b0 , w_12984 );
not ( w_12984 , w_12985 );
and ( w_12985 , w_12982 , w_12983 );
buf ( w_12982 , \1177_b1 );
not ( w_12982 , w_12986 );
not ( w_12983 , w_12987 );
and ( w_12986 , w_12987 , \1177_b0 );
or ( \5269_b1 , \5175_b1 , \5179_b1 );
xor ( \5269_b0 , \5175_b0 , w_12988 );
not ( w_12988 , w_12989 );
and ( w_12989 , \5179_b1 , \5179_b0 );
or ( \5270_b1 , \5269_b1 , \1177_b1 );
xor ( \5270_b0 , \5269_b0 , w_12990 );
not ( w_12990 , w_12991 );
and ( w_12991 , \1177_b1 , \1177_b0 );
or ( \5271_b1 , \5268_b1 , \5270_b1 );
not ( \5270_b1 , w_12992 );
and ( \5271_b0 , \5268_b0 , w_12993 );
and ( w_12992 , w_12993 , \5270_b0 );
or ( \5272_b1 , \5187_b1 , \5191_b1 );
xor ( \5272_b0 , \5187_b0 , w_12994 );
not ( w_12994 , w_12995 );
and ( w_12995 , \5191_b1 , \5191_b0 );
or ( \5273_b1 , \5272_b1 , \5196_b1 );
xor ( \5273_b0 , \5272_b0 , w_12996 );
not ( w_12996 , w_12997 );
and ( w_12997 , \5196_b1 , \5196_b0 );
or ( \5274_b1 , \5270_b1 , \5273_b1 );
not ( \5273_b1 , w_12998 );
and ( \5274_b0 , \5270_b0 , w_12999 );
and ( w_12998 , w_12999 , \5273_b0 );
or ( \5275_b1 , \5268_b1 , \5273_b1 );
not ( \5273_b1 , w_13000 );
and ( \5275_b0 , \5268_b0 , w_13001 );
and ( w_13000 , w_13001 , \5273_b0 );
or ( \5277_b1 , \5266_b1 , \5276_b1 );
not ( \5276_b1 , w_13002 );
and ( \5277_b0 , \5266_b0 , w_13003 );
and ( w_13002 , w_13003 , \5276_b0 );
or ( \5278_b1 , \5131_b1 , \5135_b1 );
xor ( \5278_b0 , \5131_b0 , w_13004 );
not ( w_13004 , w_13005 );
and ( w_13005 , \5135_b1 , \5135_b0 );
or ( \5279_b1 , \5278_b1 , \5140_b1 );
xor ( \5279_b0 , \5278_b0 , w_13006 );
not ( w_13006 , w_13007 );
and ( w_13007 , \5140_b1 , \5140_b0 );
or ( \5280_b1 , \5276_b1 , \5279_b1 );
not ( \5279_b1 , w_13008 );
and ( \5280_b0 , \5276_b0 , w_13009 );
and ( w_13008 , w_13009 , \5279_b0 );
or ( \5281_b1 , \5266_b1 , \5279_b1 );
not ( \5279_b1 , w_13010 );
and ( \5281_b0 , \5266_b0 , w_13011 );
and ( w_13010 , w_13011 , \5279_b0 );
or ( \5283_b1 , \5115_b1 , \5119_b1 );
xor ( \5283_b0 , \5115_b0 , w_13012 );
not ( w_13012 , w_13013 );
and ( w_13013 , \5119_b1 , \5119_b0 );
or ( \5284_b1 , \5283_b1 , \5124_b1 );
xor ( \5284_b0 , \5283_b0 , w_13014 );
not ( w_13014 , w_13015 );
and ( w_13015 , \5124_b1 , \5124_b0 );
or ( \5285_b1 , \5183_b1 , \5199_b1 );
xor ( \5285_b0 , \5183_b0 , w_13016 );
not ( w_13016 , w_13017 );
and ( w_13017 , \5199_b1 , \5199_b0 );
or ( \5286_b1 , \5285_b1 , \5204_b1 );
xor ( \5286_b0 , \5285_b0 , w_13018 );
not ( w_13018 , w_13019 );
and ( w_13019 , \5204_b1 , \5204_b0 );
or ( \5287_b1 , \5284_b1 , \5286_b1 );
not ( \5286_b1 , w_13020 );
and ( \5287_b0 , \5284_b0 , w_13021 );
and ( w_13020 , w_13021 , \5286_b0 );
or ( \5288_b1 , \5282_b1 , \5287_b1 );
not ( \5287_b1 , w_13022 );
and ( \5288_b0 , \5282_b0 , w_13023 );
and ( w_13022 , w_13023 , \5287_b0 );
or ( \5289_b1 , \5207_b1 , \5209_b1 );
xor ( \5289_b0 , \5207_b0 , w_13024 );
not ( w_13024 , w_13025 );
and ( w_13025 , \5209_b1 , \5209_b0 );
or ( \5290_b1 , \5289_b1 , \5211_b1 );
xor ( \5290_b0 , \5289_b0 , w_13026 );
not ( w_13026 , w_13027 );
and ( w_13027 , \5211_b1 , \5211_b0 );
or ( \5291_b1 , \5287_b1 , \5290_b1 );
not ( \5290_b1 , w_13028 );
and ( \5291_b0 , \5287_b0 , w_13029 );
and ( w_13028 , w_13029 , \5290_b0 );
or ( \5292_b1 , \5282_b1 , \5290_b1 );
not ( \5290_b1 , w_13030 );
and ( \5292_b0 , \5282_b0 , w_13031 );
and ( w_13030 , w_13031 , \5290_b0 );
or ( \5294_b1 , \5226_b1 , \5293_b1 );
not ( \5293_b1 , w_13032 );
and ( \5294_b0 , \5226_b0 , w_13033 );
and ( w_13032 , w_13033 , \5293_b0 );
or ( \5295_b1 , \5226_b1 , \5293_b1 );
xor ( \5295_b0 , \5226_b0 , w_13034 );
not ( w_13034 , w_13035 );
and ( w_13035 , \5293_b1 , \5293_b0 );
or ( \5296_b1 , \5282_b1 , \5287_b1 );
xor ( \5296_b0 , \5282_b0 , w_13036 );
not ( w_13036 , w_13037 );
and ( w_13037 , \5287_b1 , \5287_b0 );
or ( \5297_b1 , \5296_b1 , \5290_b1 );
xor ( \5297_b0 , \5296_b0 , w_13038 );
not ( w_13038 , w_13039 );
and ( w_13039 , \5290_b1 , \5290_b0 );
or ( \5298_b1 , \2161_b1 , \2261_b1 );
not ( \2261_b1 , w_13040 );
and ( \5298_b0 , \2161_b0 , w_13041 );
and ( w_13040 , w_13041 , \2261_b0 );
or ( \5299_b1 , \2028_b1 , \2259_b1 );
not ( \2259_b1 , w_13042 );
and ( \5299_b0 , \2028_b0 , w_13043 );
and ( w_13042 , w_13043 , \2259_b0 );
or ( \5300_b1 , \5298_b1 , w_13045 );
not ( w_13045 , w_13046 );
and ( \5300_b0 , \5298_b0 , w_13047 );
and ( w_13046 ,  , w_13047 );
buf ( w_13045 , \5299_b1 );
not ( w_13045 , w_13048 );
not (  , w_13049 );
and ( w_13048 , w_13049 , \5299_b0 );
or ( \5301_b1 , \5300_b1 , w_13050 );
xor ( \5301_b0 , \5300_b0 , w_13052 );
not ( w_13052 , w_13053 );
and ( w_13053 , w_13050 , w_13051 );
buf ( w_13050 , \2124_b1 );
not ( w_13050 , w_13054 );
not ( w_13051 , w_13055 );
and ( w_13054 , w_13055 , \2124_b0 );
or ( \5302_b1 , \2532_b1 , \1955_b1 );
not ( \1955_b1 , w_13056 );
and ( \5302_b0 , \2532_b0 , w_13057 );
and ( w_13056 , w_13057 , \1955_b0 );
or ( \5303_b1 , \2305_b1 , \1953_b1 );
not ( \1953_b1 , w_13058 );
and ( \5303_b0 , \2305_b0 , w_13059 );
and ( w_13058 , w_13059 , \1953_b0 );
or ( \5304_b1 , \5302_b1 , w_13061 );
not ( w_13061 , w_13062 );
and ( \5304_b0 , \5302_b0 , w_13063 );
and ( w_13062 ,  , w_13063 );
buf ( w_13061 , \5303_b1 );
not ( w_13061 , w_13064 );
not (  , w_13065 );
and ( w_13064 , w_13065 , \5303_b0 );
or ( \5305_b1 , \5304_b1 , w_13066 );
xor ( \5305_b0 , \5304_b0 , w_13068 );
not ( w_13068 , w_13069 );
and ( w_13069 , w_13066 , w_13067 );
buf ( w_13066 , \1835_b1 );
not ( w_13066 , w_13070 );
not ( w_13067 , w_13071 );
and ( w_13070 , w_13071 , \1835_b0 );
or ( \5306_b1 , \5301_b1 , \5305_b1 );
not ( \5305_b1 , w_13072 );
and ( \5306_b0 , \5301_b0 , w_13073 );
and ( w_13072 , w_13073 , \5305_b0 );
or ( \5307_b1 , \2763_b1 , \1742_b1 );
not ( \1742_b1 , w_13074 );
and ( \5307_b0 , \2763_b0 , w_13075 );
and ( w_13074 , w_13075 , \1742_b0 );
or ( \5308_b1 , \2541_b1 , \1740_b1 );
not ( \1740_b1 , w_13076 );
and ( \5308_b0 , \2541_b0 , w_13077 );
and ( w_13076 , w_13077 , \1740_b0 );
or ( \5309_b1 , \5307_b1 , w_13079 );
not ( w_13079 , w_13080 );
and ( \5309_b0 , \5307_b0 , w_13081 );
and ( w_13080 ,  , w_13081 );
buf ( w_13079 , \5308_b1 );
not ( w_13079 , w_13082 );
not (  , w_13083 );
and ( w_13082 , w_13083 , \5308_b0 );
or ( \5310_b1 , \5309_b1 , w_13084 );
xor ( \5310_b0 , \5309_b0 , w_13086 );
not ( w_13086 , w_13087 );
and ( w_13087 , w_13084 , w_13085 );
buf ( w_13084 , \1610_b1 );
not ( w_13084 , w_13088 );
not ( w_13085 , w_13089 );
and ( w_13088 , w_13089 , \1610_b0 );
or ( \5311_b1 , \5305_b1 , \5310_b1 );
not ( \5310_b1 , w_13090 );
and ( \5311_b0 , \5305_b0 , w_13091 );
and ( w_13090 , w_13091 , \5310_b0 );
or ( \5312_b1 , \5301_b1 , \5310_b1 );
not ( \5310_b1 , w_13092 );
and ( \5312_b0 , \5301_b0 , w_13093 );
and ( w_13092 , w_13093 , \5310_b0 );
or ( \5314_b1 , \1770_b1 , \2913_b1 );
not ( \2913_b1 , w_13094 );
and ( \5314_b0 , \1770_b0 , w_13095 );
and ( w_13094 , w_13095 , \2913_b0 );
or ( \5315_b1 , \1537_b1 , \2910_b1 );
not ( \2910_b1 , w_13096 );
and ( \5315_b0 , \1537_b0 , w_13097 );
and ( w_13096 , w_13097 , \2910_b0 );
or ( \5316_b1 , \5314_b1 , w_13099 );
not ( w_13099 , w_13100 );
and ( \5316_b0 , \5314_b0 , w_13101 );
and ( w_13100 ,  , w_13101 );
buf ( w_13099 , \5315_b1 );
not ( w_13099 , w_13102 );
not (  , w_13103 );
and ( w_13102 , w_13103 , \5315_b0 );
or ( \5317_b1 , \5316_b1 , w_13104 );
xor ( \5317_b0 , \5316_b0 , w_13106 );
not ( w_13106 , w_13107 );
and ( w_13107 , w_13104 , w_13105 );
buf ( w_13104 , \2371_b1 );
not ( w_13104 , w_13108 );
not ( w_13105 , w_13109 );
and ( w_13108 , w_13109 , \2371_b0 );
or ( \5318_b1 , \2023_b1 , \2550_b1 );
not ( \2550_b1 , w_13110 );
and ( \5318_b0 , \2023_b0 , w_13111 );
and ( w_13110 , w_13111 , \2550_b0 );
or ( \5319_b1 , \1778_b1 , \2548_b1 );
not ( \2548_b1 , w_13112 );
and ( \5319_b0 , \1778_b0 , w_13113 );
and ( w_13112 , w_13113 , \2548_b0 );
or ( \5320_b1 , \5318_b1 , w_13115 );
not ( w_13115 , w_13116 );
and ( \5320_b0 , \5318_b0 , w_13117 );
and ( w_13116 ,  , w_13117 );
buf ( w_13115 , \5319_b1 );
not ( w_13115 , w_13118 );
not (  , w_13119 );
and ( w_13118 , w_13119 , \5319_b0 );
or ( \5321_b1 , \5320_b1 , w_13120 );
xor ( \5321_b0 , \5320_b0 , w_13122 );
not ( w_13122 , w_13123 );
and ( w_13123 , w_13120 , w_13121 );
buf ( w_13120 , \2374_b1 );
not ( w_13120 , w_13124 );
not ( w_13121 , w_13125 );
and ( w_13124 , w_13125 , \2374_b0 );
or ( \5322_b1 , \5317_b1 , \5321_b1 );
not ( \5321_b1 , w_13126 );
and ( \5322_b0 , \5317_b0 , w_13127 );
and ( w_13126 , w_13127 , \5321_b0 );
or ( \5323_b1 , \5321_b1 , \1363_b1 );
not ( \1363_b1 , w_13128 );
and ( \5323_b0 , \5321_b0 , w_13129 );
and ( w_13128 , w_13129 , \1363_b0 );
or ( \5324_b1 , \5317_b1 , \1363_b1 );
not ( \1363_b1 , w_13130 );
and ( \5324_b0 , \5317_b0 , w_13131 );
and ( w_13130 , w_13131 , \1363_b0 );
or ( \5326_b1 , \5313_b1 , \5325_b1 );
not ( \5325_b1 , w_13132 );
and ( \5326_b0 , \5313_b0 , w_13133 );
and ( w_13132 , w_13133 , \5325_b0 );
or ( \5327_b1 , \5230_b1 , \5234_b1 );
xor ( \5327_b0 , \5230_b0 , w_13134 );
not ( w_13134 , w_13135 );
and ( w_13135 , \5234_b1 , \5234_b0 );
or ( \5328_b1 , \5327_b1 , \5239_b1 );
xor ( \5328_b0 , \5327_b0 , w_13136 );
not ( w_13136 , w_13137 );
and ( w_13137 , \5239_b1 , \5239_b0 );
or ( \5329_b1 , \5325_b1 , \5328_b1 );
not ( \5328_b1 , w_13138 );
and ( \5329_b0 , \5325_b0 , w_13139 );
and ( w_13138 , w_13139 , \5328_b0 );
or ( \5330_b1 , \5313_b1 , \5328_b1 );
not ( \5328_b1 , w_13140 );
and ( \5330_b0 , \5313_b0 , w_13141 );
and ( w_13140 , w_13141 , \5328_b0 );
or ( \5332_b1 , \5242_b1 , \5258_b1 );
xor ( \5332_b0 , \5242_b0 , w_13142 );
not ( w_13142 , w_13143 );
and ( w_13143 , \5258_b1 , \5258_b0 );
or ( \5333_b1 , \5332_b1 , \5263_b1 );
xor ( \5333_b0 , \5332_b0 , w_13144 );
not ( w_13144 , w_13145 );
and ( w_13145 , \5263_b1 , \5263_b0 );
or ( \5334_b1 , \5331_b1 , \5333_b1 );
not ( \5333_b1 , w_13146 );
and ( \5334_b0 , \5331_b0 , w_13147 );
and ( w_13146 , w_13147 , \5333_b0 );
or ( \5335_b1 , \5268_b1 , \5270_b1 );
xor ( \5335_b0 , \5268_b0 , w_13148 );
not ( w_13148 , w_13149 );
and ( w_13149 , \5270_b1 , \5270_b0 );
or ( \5336_b1 , \5335_b1 , \5273_b1 );
xor ( \5336_b0 , \5335_b0 , w_13150 );
not ( w_13150 , w_13151 );
and ( w_13151 , \5273_b1 , \5273_b0 );
or ( \5337_b1 , \5333_b1 , \5336_b1 );
not ( \5336_b1 , w_13152 );
and ( \5337_b0 , \5333_b0 , w_13153 );
and ( w_13152 , w_13153 , \5336_b0 );
or ( \5338_b1 , \5331_b1 , \5336_b1 );
not ( \5336_b1 , w_13154 );
and ( \5338_b0 , \5331_b0 , w_13155 );
and ( w_13154 , w_13155 , \5336_b0 );
or ( \5340_b1 , \5266_b1 , \5276_b1 );
xor ( \5340_b0 , \5266_b0 , w_13156 );
not ( w_13156 , w_13157 );
and ( w_13157 , \5276_b1 , \5276_b0 );
or ( \5341_b1 , \5340_b1 , \5279_b1 );
xor ( \5341_b0 , \5340_b0 , w_13158 );
not ( w_13158 , w_13159 );
and ( w_13159 , \5279_b1 , \5279_b0 );
or ( \5342_b1 , \5339_b1 , \5341_b1 );
not ( \5341_b1 , w_13160 );
and ( \5342_b0 , \5339_b0 , w_13161 );
and ( w_13160 , w_13161 , \5341_b0 );
or ( \5343_b1 , \5284_b1 , \5286_b1 );
xor ( \5343_b0 , \5284_b0 , w_13162 );
not ( w_13162 , w_13163 );
and ( w_13163 , \5286_b1 , \5286_b0 );
or ( \5344_b1 , \5341_b1 , \5343_b1 );
not ( \5343_b1 , w_13164 );
and ( \5344_b0 , \5341_b0 , w_13165 );
and ( w_13164 , w_13165 , \5343_b0 );
or ( \5345_b1 , \5339_b1 , \5343_b1 );
not ( \5343_b1 , w_13166 );
and ( \5345_b0 , \5339_b0 , w_13167 );
and ( w_13166 , w_13167 , \5343_b0 );
or ( \5347_b1 , \5297_b1 , \5346_b1 );
not ( \5346_b1 , w_13168 );
and ( \5347_b0 , \5297_b0 , w_13169 );
and ( w_13168 , w_13169 , \5346_b0 );
or ( \5348_b1 , \5297_b1 , \5346_b1 );
xor ( \5348_b0 , \5297_b0 , w_13170 );
not ( w_13170 , w_13171 );
and ( w_13171 , \5346_b1 , \5346_b0 );
or ( \5349_b1 , \5339_b1 , \5341_b1 );
xor ( \5349_b0 , \5339_b0 , w_13172 );
not ( w_13172 , w_13173 );
and ( w_13173 , \5341_b1 , \5341_b0 );
or ( \5350_b1 , \5349_b1 , \5343_b1 );
xor ( \5350_b0 , \5349_b0 , w_13174 );
not ( w_13174 , w_13175 );
and ( w_13175 , \5343_b1 , \5343_b0 );
or ( \5351_b1 , \1778_b1 , \2913_b1 );
not ( \2913_b1 , w_13176 );
and ( \5351_b0 , \1778_b0 , w_13177 );
and ( w_13176 , w_13177 , \2913_b0 );
or ( \5352_b1 , \1770_b1 , \2910_b1 );
not ( \2910_b1 , w_13178 );
and ( \5352_b0 , \1770_b0 , w_13179 );
and ( w_13178 , w_13179 , \2910_b0 );
or ( \5353_b1 , \5351_b1 , w_13181 );
not ( w_13181 , w_13182 );
and ( \5353_b0 , \5351_b0 , w_13183 );
and ( w_13182 ,  , w_13183 );
buf ( w_13181 , \5352_b1 );
not ( w_13181 , w_13184 );
not (  , w_13185 );
and ( w_13184 , w_13185 , \5352_b0 );
or ( \5354_b1 , \5353_b1 , w_13186 );
xor ( \5354_b0 , \5353_b0 , w_13188 );
not ( w_13188 , w_13189 );
and ( w_13189 , w_13186 , w_13187 );
buf ( w_13186 , \2371_b1 );
not ( w_13186 , w_13190 );
not ( w_13187 , w_13191 );
and ( w_13190 , w_13191 , \2371_b0 );
or ( \5355_b1 , \2028_b1 , \2550_b1 );
not ( \2550_b1 , w_13192 );
and ( \5355_b0 , \2028_b0 , w_13193 );
and ( w_13192 , w_13193 , \2550_b0 );
or ( \5356_b1 , \2023_b1 , \2548_b1 );
not ( \2548_b1 , w_13194 );
and ( \5356_b0 , \2023_b0 , w_13195 );
and ( w_13194 , w_13195 , \2548_b0 );
or ( \5357_b1 , \5355_b1 , w_13197 );
not ( w_13197 , w_13198 );
and ( \5357_b0 , \5355_b0 , w_13199 );
and ( w_13198 ,  , w_13199 );
buf ( w_13197 , \5356_b1 );
not ( w_13197 , w_13200 );
not (  , w_13201 );
and ( w_13200 , w_13201 , \5356_b0 );
or ( \5358_b1 , \5357_b1 , w_13202 );
xor ( \5358_b0 , \5357_b0 , w_13204 );
not ( w_13204 , w_13205 );
and ( w_13205 , w_13202 , w_13203 );
buf ( w_13202 , \2374_b1 );
not ( w_13202 , w_13206 );
not ( w_13203 , w_13207 );
and ( w_13206 , w_13207 , \2374_b0 );
or ( \5359_b1 , \5354_b1 , \5358_b1 );
not ( \5358_b1 , w_13208 );
and ( \5359_b0 , \5354_b0 , w_13209 );
and ( w_13208 , w_13209 , \5358_b0 );
or ( \5360_b1 , \2305_b1 , \2261_b1 );
not ( \2261_b1 , w_13210 );
and ( \5360_b0 , \2305_b0 , w_13211 );
and ( w_13210 , w_13211 , \2261_b0 );
or ( \5361_b1 , \2161_b1 , \2259_b1 );
not ( \2259_b1 , w_13212 );
and ( \5361_b0 , \2161_b0 , w_13213 );
and ( w_13212 , w_13213 , \2259_b0 );
or ( \5362_b1 , \5360_b1 , w_13215 );
not ( w_13215 , w_13216 );
and ( \5362_b0 , \5360_b0 , w_13217 );
and ( w_13216 ,  , w_13217 );
buf ( w_13215 , \5361_b1 );
not ( w_13215 , w_13218 );
not (  , w_13219 );
and ( w_13218 , w_13219 , \5361_b0 );
or ( \5363_b1 , \5362_b1 , w_13220 );
xor ( \5363_b0 , \5362_b0 , w_13222 );
not ( w_13222 , w_13223 );
and ( w_13223 , w_13220 , w_13221 );
buf ( w_13220 , \2124_b1 );
not ( w_13220 , w_13224 );
not ( w_13221 , w_13225 );
and ( w_13224 , w_13225 , \2124_b0 );
or ( \5364_b1 , \5358_b1 , \5363_b1 );
not ( \5363_b1 , w_13226 );
and ( \5364_b0 , \5358_b0 , w_13227 );
and ( w_13226 , w_13227 , \5363_b0 );
or ( \5365_b1 , \5354_b1 , \5363_b1 );
not ( \5363_b1 , w_13228 );
and ( \5365_b0 , \5354_b0 , w_13229 );
and ( w_13228 , w_13229 , \5363_b0 );
or ( \5367_b1 , \2850_b1 , w_13231 );
not ( w_13231 , w_13232 );
and ( \5367_b0 , \2850_b0 , w_13233 );
and ( w_13232 ,  , w_13233 );
buf ( w_13231 , \1474_b1 );
not ( w_13231 , w_13234 );
not (  , w_13235 );
and ( w_13234 , w_13235 , \1474_b0 );
or ( \5368_b1 , \5367_b1 , w_13236 );
xor ( \5368_b0 , \5367_b0 , w_13238 );
not ( w_13238 , w_13239 );
and ( w_13239 , w_13236 , w_13237 );
buf ( w_13236 , \1363_b1 );
not ( w_13236 , w_13240 );
not ( w_13237 , w_13241 );
and ( w_13240 , w_13241 , \1363_b0 );
or ( \5369_b1 , \5366_b1 , \5368_b1 );
not ( \5368_b1 , w_13242 );
and ( \5369_b0 , \5366_b0 , w_13243 );
and ( w_13242 , w_13243 , \5368_b0 );
or ( \5370_b1 , \5301_b1 , \5305_b1 );
xor ( \5370_b0 , \5301_b0 , w_13244 );
not ( w_13244 , w_13245 );
and ( w_13245 , \5305_b1 , \5305_b0 );
or ( \5371_b1 , \5370_b1 , \5310_b1 );
xor ( \5371_b0 , \5370_b0 , w_13246 );
not ( w_13246 , w_13247 );
and ( w_13247 , \5310_b1 , \5310_b0 );
or ( \5372_b1 , \5368_b1 , \5371_b1 );
not ( \5371_b1 , w_13248 );
and ( \5372_b0 , \5368_b0 , w_13249 );
and ( w_13248 , w_13249 , \5371_b0 );
or ( \5373_b1 , \5366_b1 , \5371_b1 );
not ( \5371_b1 , w_13250 );
and ( \5373_b0 , \5366_b0 , w_13251 );
and ( w_13250 , w_13251 , \5371_b0 );
or ( \5375_b1 , \5246_b1 , \5250_b1 );
xor ( \5375_b0 , \5246_b0 , w_13252 );
not ( w_13252 , w_13253 );
and ( w_13253 , \5250_b1 , \5250_b0 );
or ( \5376_b1 , \5375_b1 , \5255_b1 );
xor ( \5376_b0 , \5375_b0 , w_13254 );
not ( w_13254 , w_13255 );
and ( w_13255 , \5255_b1 , \5255_b0 );
or ( \5377_b1 , \5374_b1 , \5376_b1 );
not ( \5376_b1 , w_13256 );
and ( \5377_b0 , \5374_b0 , w_13257 );
and ( w_13256 , w_13257 , \5376_b0 );
or ( \5378_b1 , \5313_b1 , \5325_b1 );
xor ( \5378_b0 , \5313_b0 , w_13258 );
not ( w_13258 , w_13259 );
and ( w_13259 , \5325_b1 , \5325_b0 );
or ( \5379_b1 , \5378_b1 , \5328_b1 );
xor ( \5379_b0 , \5378_b0 , w_13260 );
not ( w_13260 , w_13261 );
and ( w_13261 , \5328_b1 , \5328_b0 );
or ( \5380_b1 , \5376_b1 , \5379_b1 );
not ( \5379_b1 , w_13262 );
and ( \5380_b0 , \5376_b0 , w_13263 );
and ( w_13262 , w_13263 , \5379_b0 );
or ( \5381_b1 , \5374_b1 , \5379_b1 );
not ( \5379_b1 , w_13264 );
and ( \5381_b0 , \5374_b0 , w_13265 );
and ( w_13264 , w_13265 , \5379_b0 );
or ( \5383_b1 , \5331_b1 , \5333_b1 );
xor ( \5383_b0 , \5331_b0 , w_13266 );
not ( w_13266 , w_13267 );
and ( w_13267 , \5333_b1 , \5333_b0 );
or ( \5384_b1 , \5383_b1 , \5336_b1 );
xor ( \5384_b0 , \5383_b0 , w_13268 );
not ( w_13268 , w_13269 );
and ( w_13269 , \5336_b1 , \5336_b0 );
or ( \5385_b1 , \5382_b1 , \5384_b1 );
not ( \5384_b1 , w_13270 );
and ( \5385_b0 , \5382_b0 , w_13271 );
and ( w_13270 , w_13271 , \5384_b0 );
or ( \5386_b1 , \5350_b1 , \5385_b1 );
not ( \5385_b1 , w_13272 );
and ( \5386_b0 , \5350_b0 , w_13273 );
and ( w_13272 , w_13273 , \5385_b0 );
or ( \5387_b1 , \5350_b1 , \5385_b1 );
xor ( \5387_b0 , \5350_b0 , w_13274 );
not ( w_13274 , w_13275 );
and ( w_13275 , \5385_b1 , \5385_b0 );
or ( \5388_b1 , \5382_b1 , \5384_b1 );
xor ( \5388_b0 , \5382_b0 , w_13276 );
not ( w_13276 , w_13277 );
and ( w_13277 , \5384_b1 , \5384_b0 );
or ( \5389_b1 , \2532_b1 , \2261_b1 );
not ( \2261_b1 , w_13278 );
and ( \5389_b0 , \2532_b0 , w_13279 );
and ( w_13278 , w_13279 , \2261_b0 );
or ( \5390_b1 , \2305_b1 , \2259_b1 );
not ( \2259_b1 , w_13280 );
and ( \5390_b0 , \2305_b0 , w_13281 );
and ( w_13280 , w_13281 , \2259_b0 );
or ( \5391_b1 , \5389_b1 , w_13283 );
not ( w_13283 , w_13284 );
and ( \5391_b0 , \5389_b0 , w_13285 );
and ( w_13284 ,  , w_13285 );
buf ( w_13283 , \5390_b1 );
not ( w_13283 , w_13286 );
not (  , w_13287 );
and ( w_13286 , w_13287 , \5390_b0 );
or ( \5392_b1 , \5391_b1 , w_13288 );
xor ( \5392_b0 , \5391_b0 , w_13290 );
not ( w_13290 , w_13291 );
and ( w_13291 , w_13288 , w_13289 );
buf ( w_13288 , \2124_b1 );
not ( w_13288 , w_13292 );
not ( w_13289 , w_13293 );
and ( w_13292 , w_13293 , \2124_b0 );
or ( \5393_b1 , \2763_b1 , \1955_b1 );
not ( \1955_b1 , w_13294 );
and ( \5393_b0 , \2763_b0 , w_13295 );
and ( w_13294 , w_13295 , \1955_b0 );
or ( \5394_b1 , \2541_b1 , \1953_b1 );
not ( \1953_b1 , w_13296 );
and ( \5394_b0 , \2541_b0 , w_13297 );
and ( w_13296 , w_13297 , \1953_b0 );
or ( \5395_b1 , \5393_b1 , w_13299 );
not ( w_13299 , w_13300 );
and ( \5395_b0 , \5393_b0 , w_13301 );
and ( w_13300 ,  , w_13301 );
buf ( w_13299 , \5394_b1 );
not ( w_13299 , w_13302 );
not (  , w_13303 );
and ( w_13302 , w_13303 , \5394_b0 );
or ( \5396_b1 , \5395_b1 , w_13304 );
xor ( \5396_b0 , \5395_b0 , w_13306 );
not ( w_13306 , w_13307 );
and ( w_13307 , w_13304 , w_13305 );
buf ( w_13304 , \1835_b1 );
not ( w_13304 , w_13308 );
not ( w_13305 , w_13309 );
and ( w_13308 , w_13309 , \1835_b0 );
or ( \5397_b1 , \5392_b1 , \5396_b1 );
not ( \5396_b1 , w_13310 );
and ( \5397_b0 , \5392_b0 , w_13311 );
and ( w_13310 , w_13311 , \5396_b0 );
or ( \5398_b1 , \2850_b1 , w_13313 );
not ( w_13313 , w_13314 );
and ( \5398_b0 , \2850_b0 , w_13315 );
and ( w_13314 ,  , w_13315 );
buf ( w_13313 , \1740_b1 );
not ( w_13313 , w_13316 );
not (  , w_13317 );
and ( w_13316 , w_13317 , \1740_b0 );
or ( \5399_b1 , \5398_b1 , w_13318 );
xor ( \5399_b0 , \5398_b0 , w_13320 );
not ( w_13320 , w_13321 );
and ( w_13321 , w_13318 , w_13319 );
buf ( w_13318 , \1610_b1 );
not ( w_13318 , w_13322 );
not ( w_13319 , w_13323 );
and ( w_13322 , w_13323 , \1610_b0 );
or ( \5400_b1 , \5396_b1 , \5399_b1 );
not ( \5399_b1 , w_13324 );
and ( \5400_b0 , \5396_b0 , w_13325 );
and ( w_13324 , w_13325 , \5399_b0 );
or ( \5401_b1 , \5392_b1 , \5399_b1 );
not ( \5399_b1 , w_13326 );
and ( \5401_b0 , \5392_b0 , w_13327 );
and ( w_13326 , w_13327 , \5399_b0 );
or ( \5403_b1 , \2023_b1 , \2913_b1 );
not ( \2913_b1 , w_13328 );
and ( \5403_b0 , \2023_b0 , w_13329 );
and ( w_13328 , w_13329 , \2913_b0 );
or ( \5404_b1 , \1778_b1 , \2910_b1 );
not ( \2910_b1 , w_13330 );
and ( \5404_b0 , \1778_b0 , w_13331 );
and ( w_13330 , w_13331 , \2910_b0 );
or ( \5405_b1 , \5403_b1 , w_13333 );
not ( w_13333 , w_13334 );
and ( \5405_b0 , \5403_b0 , w_13335 );
and ( w_13334 ,  , w_13335 );
buf ( w_13333 , \5404_b1 );
not ( w_13333 , w_13336 );
not (  , w_13337 );
and ( w_13336 , w_13337 , \5404_b0 );
or ( \5406_b1 , \5405_b1 , w_13338 );
xor ( \5406_b0 , \5405_b0 , w_13340 );
not ( w_13340 , w_13341 );
and ( w_13341 , w_13338 , w_13339 );
buf ( w_13338 , \2371_b1 );
not ( w_13338 , w_13342 );
not ( w_13339 , w_13343 );
and ( w_13342 , w_13343 , \2371_b0 );
or ( \5407_b1 , \2161_b1 , \2550_b1 );
not ( \2550_b1 , w_13344 );
and ( \5407_b0 , \2161_b0 , w_13345 );
and ( w_13344 , w_13345 , \2550_b0 );
or ( \5408_b1 , \2028_b1 , \2548_b1 );
not ( \2548_b1 , w_13346 );
and ( \5408_b0 , \2028_b0 , w_13347 );
and ( w_13346 , w_13347 , \2548_b0 );
or ( \5409_b1 , \5407_b1 , w_13349 );
not ( w_13349 , w_13350 );
and ( \5409_b0 , \5407_b0 , w_13351 );
and ( w_13350 ,  , w_13351 );
buf ( w_13349 , \5408_b1 );
not ( w_13349 , w_13352 );
not (  , w_13353 );
and ( w_13352 , w_13353 , \5408_b0 );
or ( \5410_b1 , \5409_b1 , w_13354 );
xor ( \5410_b0 , \5409_b0 , w_13356 );
not ( w_13356 , w_13357 );
and ( w_13357 , w_13354 , w_13355 );
buf ( w_13354 , \2374_b1 );
not ( w_13354 , w_13358 );
not ( w_13355 , w_13359 );
and ( w_13358 , w_13359 , \2374_b0 );
or ( \5411_b1 , \5406_b1 , \5410_b1 );
not ( \5410_b1 , w_13360 );
and ( \5411_b0 , \5406_b0 , w_13361 );
and ( w_13360 , w_13361 , \5410_b0 );
or ( \5412_b1 , \5410_b1 , \1610_b1 );
not ( \1610_b1 , w_13362 );
and ( \5412_b0 , \5410_b0 , w_13363 );
and ( w_13362 , w_13363 , \1610_b0 );
or ( \5413_b1 , \5406_b1 , \1610_b1 );
not ( \1610_b1 , w_13364 );
and ( \5413_b0 , \5406_b0 , w_13365 );
and ( w_13364 , w_13365 , \1610_b0 );
or ( \5415_b1 , \5402_b1 , \5414_b1 );
not ( \5414_b1 , w_13366 );
and ( \5415_b0 , \5402_b0 , w_13367 );
and ( w_13366 , w_13367 , \5414_b0 );
or ( \5416_b1 , \2541_b1 , \1955_b1 );
not ( \1955_b1 , w_13368 );
and ( \5416_b0 , \2541_b0 , w_13369 );
and ( w_13368 , w_13369 , \1955_b0 );
or ( \5417_b1 , \2532_b1 , \1953_b1 );
not ( \1953_b1 , w_13370 );
and ( \5417_b0 , \2532_b0 , w_13371 );
and ( w_13370 , w_13371 , \1953_b0 );
or ( \5418_b1 , \5416_b1 , w_13373 );
not ( w_13373 , w_13374 );
and ( \5418_b0 , \5416_b0 , w_13375 );
and ( w_13374 ,  , w_13375 );
buf ( w_13373 , \5417_b1 );
not ( w_13373 , w_13376 );
not (  , w_13377 );
and ( w_13376 , w_13377 , \5417_b0 );
or ( \5419_b1 , \5418_b1 , w_13378 );
xor ( \5419_b0 , \5418_b0 , w_13380 );
not ( w_13380 , w_13381 );
and ( w_13381 , w_13378 , w_13379 );
buf ( w_13378 , \1835_b1 );
not ( w_13378 , w_13382 );
not ( w_13379 , w_13383 );
and ( w_13382 , w_13383 , \1835_b0 );
or ( \5420_b1 , \5414_b1 , \5419_b1 );
not ( \5419_b1 , w_13384 );
and ( \5420_b0 , \5414_b0 , w_13385 );
and ( w_13384 , w_13385 , \5419_b0 );
or ( \5421_b1 , \5402_b1 , \5419_b1 );
not ( \5419_b1 , w_13386 );
and ( \5421_b0 , \5402_b0 , w_13387 );
and ( w_13386 , w_13387 , \5419_b0 );
or ( \5423_b1 , \2850_b1 , \1742_b1 );
not ( \1742_b1 , w_13388 );
and ( \5423_b0 , \2850_b0 , w_13389 );
and ( w_13388 , w_13389 , \1742_b0 );
or ( \5424_b1 , \2763_b1 , \1740_b1 );
not ( \1740_b1 , w_13390 );
and ( \5424_b0 , \2763_b0 , w_13391 );
and ( w_13390 , w_13391 , \1740_b0 );
or ( \5425_b1 , \5423_b1 , w_13393 );
not ( w_13393 , w_13394 );
and ( \5425_b0 , \5423_b0 , w_13395 );
and ( w_13394 ,  , w_13395 );
buf ( w_13393 , \5424_b1 );
not ( w_13393 , w_13396 );
not (  , w_13397 );
and ( w_13396 , w_13397 , \5424_b0 );
or ( \5426_b1 , \5425_b1 , w_13398 );
xor ( \5426_b0 , \5425_b0 , w_13400 );
not ( w_13400 , w_13401 );
and ( w_13401 , w_13398 , w_13399 );
buf ( w_13398 , \1610_b1 );
not ( w_13398 , w_13402 );
not ( w_13399 , w_13403 );
and ( w_13402 , w_13403 , \1610_b0 );
or ( \5427_b1 , \5354_b1 , \5358_b1 );
xor ( \5427_b0 , \5354_b0 , w_13404 );
not ( w_13404 , w_13405 );
and ( w_13405 , \5358_b1 , \5358_b0 );
or ( \5428_b1 , \5427_b1 , \5363_b1 );
xor ( \5428_b0 , \5427_b0 , w_13406 );
not ( w_13406 , w_13407 );
and ( w_13407 , \5363_b1 , \5363_b0 );
or ( \5429_b1 , \5426_b1 , \5428_b1 );
not ( \5428_b1 , w_13408 );
and ( \5429_b0 , \5426_b0 , w_13409 );
and ( w_13408 , w_13409 , \5428_b0 );
or ( \5430_b1 , \5422_b1 , \5429_b1 );
not ( \5429_b1 , w_13410 );
and ( \5430_b0 , \5422_b0 , w_13411 );
and ( w_13410 , w_13411 , \5429_b0 );
or ( \5431_b1 , \5317_b1 , \5321_b1 );
xor ( \5431_b0 , \5317_b0 , w_13412 );
not ( w_13412 , w_13413 );
and ( w_13413 , \5321_b1 , \5321_b0 );
or ( \5432_b1 , \5431_b1 , \1363_b1 );
xor ( \5432_b0 , \5431_b0 , w_13414 );
not ( w_13414 , w_13415 );
and ( w_13415 , \1363_b1 , \1363_b0 );
or ( \5433_b1 , \5429_b1 , \5432_b1 );
not ( \5432_b1 , w_13416 );
and ( \5433_b0 , \5429_b0 , w_13417 );
and ( w_13416 , w_13417 , \5432_b0 );
or ( \5434_b1 , \5422_b1 , \5432_b1 );
not ( \5432_b1 , w_13418 );
and ( \5434_b0 , \5422_b0 , w_13419 );
and ( w_13418 , w_13419 , \5432_b0 );
or ( \5436_b1 , \5374_b1 , \5376_b1 );
xor ( \5436_b0 , \5374_b0 , w_13420 );
not ( w_13420 , w_13421 );
and ( w_13421 , \5376_b1 , \5376_b0 );
or ( \5437_b1 , \5436_b1 , \5379_b1 );
xor ( \5437_b0 , \5436_b0 , w_13422 );
not ( w_13422 , w_13423 );
and ( w_13423 , \5379_b1 , \5379_b0 );
or ( \5438_b1 , \5435_b1 , \5437_b1 );
not ( \5437_b1 , w_13424 );
and ( \5438_b0 , \5435_b0 , w_13425 );
and ( w_13424 , w_13425 , \5437_b0 );
or ( \5439_b1 , \5388_b1 , \5438_b1 );
not ( \5438_b1 , w_13426 );
and ( \5439_b0 , \5388_b0 , w_13427 );
and ( w_13426 , w_13427 , \5438_b0 );
or ( \5440_b1 , \5388_b1 , \5438_b1 );
xor ( \5440_b0 , \5388_b0 , w_13428 );
not ( w_13428 , w_13429 );
and ( w_13429 , \5438_b1 , \5438_b0 );
or ( \5441_b1 , \5435_b1 , \5437_b1 );
xor ( \5441_b0 , \5435_b0 , w_13430 );
not ( w_13430 , w_13431 );
and ( w_13431 , \5437_b1 , \5437_b0 );
or ( \5442_b1 , \5366_b1 , \5368_b1 );
xor ( \5442_b0 , \5366_b0 , w_13432 );
not ( w_13432 , w_13433 );
and ( w_13433 , \5368_b1 , \5368_b0 );
or ( \5443_b1 , \5442_b1 , \5371_b1 );
xor ( \5443_b0 , \5442_b0 , w_13434 );
not ( w_13434 , w_13435 );
and ( w_13435 , \5371_b1 , \5371_b0 );
or ( \5444_b1 , \5422_b1 , \5429_b1 );
xor ( \5444_b0 , \5422_b0 , w_13436 );
not ( w_13436 , w_13437 );
and ( w_13437 , \5429_b1 , \5429_b0 );
or ( \5445_b1 , \5444_b1 , \5432_b1 );
xor ( \5445_b0 , \5444_b0 , w_13438 );
not ( w_13438 , w_13439 );
and ( w_13439 , \5432_b1 , \5432_b0 );
or ( \5446_b1 , \5443_b1 , \5445_b1 );
not ( \5445_b1 , w_13440 );
and ( \5446_b0 , \5443_b0 , w_13441 );
and ( w_13440 , w_13441 , \5445_b0 );
or ( \5447_b1 , \5441_b1 , \5446_b1 );
not ( \5446_b1 , w_13442 );
and ( \5447_b0 , \5441_b0 , w_13443 );
and ( w_13442 , w_13443 , \5446_b0 );
or ( \5448_b1 , \5441_b1 , \5446_b1 );
xor ( \5448_b0 , \5441_b0 , w_13444 );
not ( w_13444 , w_13445 );
and ( w_13445 , \5446_b1 , \5446_b0 );
or ( \5449_b1 , \5443_b1 , \5445_b1 );
xor ( \5449_b0 , \5443_b0 , w_13446 );
not ( w_13446 , w_13447 );
and ( w_13447 , \5445_b1 , \5445_b0 );
or ( \5450_b1 , \2028_b1 , \2913_b1 );
not ( \2913_b1 , w_13448 );
and ( \5450_b0 , \2028_b0 , w_13449 );
and ( w_13448 , w_13449 , \2913_b0 );
or ( \5451_b1 , \2023_b1 , \2910_b1 );
not ( \2910_b1 , w_13450 );
and ( \5451_b0 , \2023_b0 , w_13451 );
and ( w_13450 , w_13451 , \2910_b0 );
or ( \5452_b1 , \5450_b1 , w_13453 );
not ( w_13453 , w_13454 );
and ( \5452_b0 , \5450_b0 , w_13455 );
and ( w_13454 ,  , w_13455 );
buf ( w_13453 , \5451_b1 );
not ( w_13453 , w_13456 );
not (  , w_13457 );
and ( w_13456 , w_13457 , \5451_b0 );
or ( \5453_b1 , \5452_b1 , w_13458 );
xor ( \5453_b0 , \5452_b0 , w_13460 );
not ( w_13460 , w_13461 );
and ( w_13461 , w_13458 , w_13459 );
buf ( w_13458 , \2371_b1 );
not ( w_13458 , w_13462 );
not ( w_13459 , w_13463 );
and ( w_13462 , w_13463 , \2371_b0 );
or ( \5454_b1 , \2305_b1 , \2550_b1 );
not ( \2550_b1 , w_13464 );
and ( \5454_b0 , \2305_b0 , w_13465 );
and ( w_13464 , w_13465 , \2550_b0 );
or ( \5455_b1 , \2161_b1 , \2548_b1 );
not ( \2548_b1 , w_13466 );
and ( \5455_b0 , \2161_b0 , w_13467 );
and ( w_13466 , w_13467 , \2548_b0 );
or ( \5456_b1 , \5454_b1 , w_13469 );
not ( w_13469 , w_13470 );
and ( \5456_b0 , \5454_b0 , w_13471 );
and ( w_13470 ,  , w_13471 );
buf ( w_13469 , \5455_b1 );
not ( w_13469 , w_13472 );
not (  , w_13473 );
and ( w_13472 , w_13473 , \5455_b0 );
or ( \5457_b1 , \5456_b1 , w_13474 );
xor ( \5457_b0 , \5456_b0 , w_13476 );
not ( w_13476 , w_13477 );
and ( w_13477 , w_13474 , w_13475 );
buf ( w_13474 , \2374_b1 );
not ( w_13474 , w_13478 );
not ( w_13475 , w_13479 );
and ( w_13478 , w_13479 , \2374_b0 );
or ( \5458_b1 , \5453_b1 , \5457_b1 );
not ( \5457_b1 , w_13480 );
and ( \5458_b0 , \5453_b0 , w_13481 );
and ( w_13480 , w_13481 , \5457_b0 );
or ( \5459_b1 , \2541_b1 , \2261_b1 );
not ( \2261_b1 , w_13482 );
and ( \5459_b0 , \2541_b0 , w_13483 );
and ( w_13482 , w_13483 , \2261_b0 );
or ( \5460_b1 , \2532_b1 , \2259_b1 );
not ( \2259_b1 , w_13484 );
and ( \5460_b0 , \2532_b0 , w_13485 );
and ( w_13484 , w_13485 , \2259_b0 );
or ( \5461_b1 , \5459_b1 , w_13487 );
not ( w_13487 , w_13488 );
and ( \5461_b0 , \5459_b0 , w_13489 );
and ( w_13488 ,  , w_13489 );
buf ( w_13487 , \5460_b1 );
not ( w_13487 , w_13490 );
not (  , w_13491 );
and ( w_13490 , w_13491 , \5460_b0 );
or ( \5462_b1 , \5461_b1 , w_13492 );
xor ( \5462_b0 , \5461_b0 , w_13494 );
not ( w_13494 , w_13495 );
and ( w_13495 , w_13492 , w_13493 );
buf ( w_13492 , \2124_b1 );
not ( w_13492 , w_13496 );
not ( w_13493 , w_13497 );
and ( w_13496 , w_13497 , \2124_b0 );
or ( \5463_b1 , \5457_b1 , \5462_b1 );
not ( \5462_b1 , w_13498 );
and ( \5463_b0 , \5457_b0 , w_13499 );
and ( w_13498 , w_13499 , \5462_b0 );
or ( \5464_b1 , \5453_b1 , \5462_b1 );
not ( \5462_b1 , w_13500 );
and ( \5464_b0 , \5453_b0 , w_13501 );
and ( w_13500 , w_13501 , \5462_b0 );
or ( \5466_b1 , \5392_b1 , \5396_b1 );
xor ( \5466_b0 , \5392_b0 , w_13502 );
not ( w_13502 , w_13503 );
and ( w_13503 , \5396_b1 , \5396_b0 );
or ( \5467_b1 , \5466_b1 , \5399_b1 );
xor ( \5467_b0 , \5466_b0 , w_13504 );
not ( w_13504 , w_13505 );
and ( w_13505 , \5399_b1 , \5399_b0 );
or ( \5468_b1 , \5465_b1 , \5467_b1 );
not ( \5467_b1 , w_13506 );
and ( \5468_b0 , \5465_b0 , w_13507 );
and ( w_13506 , w_13507 , \5467_b0 );
or ( \5469_b1 , \5406_b1 , \5410_b1 );
xor ( \5469_b0 , \5406_b0 , w_13508 );
not ( w_13508 , w_13509 );
and ( w_13509 , \5410_b1 , \5410_b0 );
or ( \5470_b1 , \5469_b1 , \1610_b1 );
xor ( \5470_b0 , \5469_b0 , w_13510 );
not ( w_13510 , w_13511 );
and ( w_13511 , \1610_b1 , \1610_b0 );
or ( \5471_b1 , \5467_b1 , \5470_b1 );
not ( \5470_b1 , w_13512 );
and ( \5471_b0 , \5467_b0 , w_13513 );
and ( w_13512 , w_13513 , \5470_b0 );
or ( \5472_b1 , \5465_b1 , \5470_b1 );
not ( \5470_b1 , w_13514 );
and ( \5472_b0 , \5465_b0 , w_13515 );
and ( w_13514 , w_13515 , \5470_b0 );
or ( \5474_b1 , \5402_b1 , \5414_b1 );
xor ( \5474_b0 , \5402_b0 , w_13516 );
not ( w_13516 , w_13517 );
and ( w_13517 , \5414_b1 , \5414_b0 );
or ( \5475_b1 , \5474_b1 , \5419_b1 );
xor ( \5475_b0 , \5474_b0 , w_13518 );
not ( w_13518 , w_13519 );
and ( w_13519 , \5419_b1 , \5419_b0 );
or ( \5476_b1 , \5473_b1 , \5475_b1 );
not ( \5475_b1 , w_13520 );
and ( \5476_b0 , \5473_b0 , w_13521 );
and ( w_13520 , w_13521 , \5475_b0 );
or ( \5477_b1 , \5426_b1 , \5428_b1 );
xor ( \5477_b0 , \5426_b0 , w_13522 );
not ( w_13522 , w_13523 );
and ( w_13523 , \5428_b1 , \5428_b0 );
or ( \5478_b1 , \5475_b1 , \5477_b1 );
not ( \5477_b1 , w_13524 );
and ( \5478_b0 , \5475_b0 , w_13525 );
and ( w_13524 , w_13525 , \5477_b0 );
or ( \5479_b1 , \5473_b1 , \5477_b1 );
not ( \5477_b1 , w_13526 );
and ( \5479_b0 , \5473_b0 , w_13527 );
and ( w_13526 , w_13527 , \5477_b0 );
or ( \5481_b1 , \5449_b1 , \5480_b1 );
not ( \5480_b1 , w_13528 );
and ( \5481_b0 , \5449_b0 , w_13529 );
and ( w_13528 , w_13529 , \5480_b0 );
or ( \5482_b1 , \5449_b1 , \5480_b1 );
xor ( \5482_b0 , \5449_b0 , w_13530 );
not ( w_13530 , w_13531 );
and ( w_13531 , \5480_b1 , \5480_b0 );
or ( \5483_b1 , \5473_b1 , \5475_b1 );
xor ( \5483_b0 , \5473_b0 , w_13532 );
not ( w_13532 , w_13533 );
and ( w_13533 , \5475_b1 , \5475_b0 );
or ( \5484_b1 , \5483_b1 , \5477_b1 );
xor ( \5484_b0 , \5483_b0 , w_13534 );
not ( w_13534 , w_13535 );
and ( w_13535 , \5477_b1 , \5477_b0 );
or ( \5485_b1 , \2161_b1 , \2913_b1 );
not ( \2913_b1 , w_13536 );
and ( \5485_b0 , \2161_b0 , w_13537 );
and ( w_13536 , w_13537 , \2913_b0 );
or ( \5486_b1 , \2028_b1 , \2910_b1 );
not ( \2910_b1 , w_13538 );
and ( \5486_b0 , \2028_b0 , w_13539 );
and ( w_13538 , w_13539 , \2910_b0 );
or ( \5487_b1 , \5485_b1 , w_13541 );
not ( w_13541 , w_13542 );
and ( \5487_b0 , \5485_b0 , w_13543 );
and ( w_13542 ,  , w_13543 );
buf ( w_13541 , \5486_b1 );
not ( w_13541 , w_13544 );
not (  , w_13545 );
and ( w_13544 , w_13545 , \5486_b0 );
or ( \5488_b1 , \5487_b1 , w_13546 );
xor ( \5488_b0 , \5487_b0 , w_13548 );
not ( w_13548 , w_13549 );
and ( w_13549 , w_13546 , w_13547 );
buf ( w_13546 , \2371_b1 );
not ( w_13546 , w_13550 );
not ( w_13547 , w_13551 );
and ( w_13550 , w_13551 , \2371_b0 );
or ( \5489_b1 , \2532_b1 , \2550_b1 );
not ( \2550_b1 , w_13552 );
and ( \5489_b0 , \2532_b0 , w_13553 );
and ( w_13552 , w_13553 , \2550_b0 );
or ( \5490_b1 , \2305_b1 , \2548_b1 );
not ( \2548_b1 , w_13554 );
and ( \5490_b0 , \2305_b0 , w_13555 );
and ( w_13554 , w_13555 , \2548_b0 );
or ( \5491_b1 , \5489_b1 , w_13557 );
not ( w_13557 , w_13558 );
and ( \5491_b0 , \5489_b0 , w_13559 );
and ( w_13558 ,  , w_13559 );
buf ( w_13557 , \5490_b1 );
not ( w_13557 , w_13560 );
not (  , w_13561 );
and ( w_13560 , w_13561 , \5490_b0 );
or ( \5492_b1 , \5491_b1 , w_13562 );
xor ( \5492_b0 , \5491_b0 , w_13564 );
not ( w_13564 , w_13565 );
and ( w_13565 , w_13562 , w_13563 );
buf ( w_13562 , \2374_b1 );
not ( w_13562 , w_13566 );
not ( w_13563 , w_13567 );
and ( w_13566 , w_13567 , \2374_b0 );
or ( \5493_b1 , \5488_b1 , \5492_b1 );
not ( \5492_b1 , w_13568 );
and ( \5493_b0 , \5488_b0 , w_13569 );
and ( w_13568 , w_13569 , \5492_b0 );
or ( \5494_b1 , \5492_b1 , \1835_b1 );
not ( \1835_b1 , w_13570 );
and ( \5494_b0 , \5492_b0 , w_13571 );
and ( w_13570 , w_13571 , \1835_b0 );
or ( \5495_b1 , \5488_b1 , \1835_b1 );
not ( \1835_b1 , w_13572 );
and ( \5495_b0 , \5488_b0 , w_13573 );
and ( w_13572 , w_13573 , \1835_b0 );
or ( \5497_b1 , \2763_b1 , \2261_b1 );
not ( \2261_b1 , w_13574 );
and ( \5497_b0 , \2763_b0 , w_13575 );
and ( w_13574 , w_13575 , \2261_b0 );
or ( \5498_b1 , \2541_b1 , \2259_b1 );
not ( \2259_b1 , w_13576 );
and ( \5498_b0 , \2541_b0 , w_13577 );
and ( w_13576 , w_13577 , \2259_b0 );
or ( \5499_b1 , \5497_b1 , w_13579 );
not ( w_13579 , w_13580 );
and ( \5499_b0 , \5497_b0 , w_13581 );
and ( w_13580 ,  , w_13581 );
buf ( w_13579 , \5498_b1 );
not ( w_13579 , w_13582 );
not (  , w_13583 );
and ( w_13582 , w_13583 , \5498_b0 );
or ( \5500_b1 , \5499_b1 , w_13584 );
xor ( \5500_b0 , \5499_b0 , w_13586 );
not ( w_13586 , w_13587 );
and ( w_13587 , w_13584 , w_13585 );
buf ( w_13584 , \2124_b1 );
not ( w_13584 , w_13588 );
not ( w_13585 , w_13589 );
and ( w_13588 , w_13589 , \2124_b0 );
or ( \5501_b1 , \2850_b1 , w_13591 );
not ( w_13591 , w_13592 );
and ( \5501_b0 , \2850_b0 , w_13593 );
and ( w_13592 ,  , w_13593 );
buf ( w_13591 , \1953_b1 );
not ( w_13591 , w_13594 );
not (  , w_13595 );
and ( w_13594 , w_13595 , \1953_b0 );
or ( \5502_b1 , \5501_b1 , w_13596 );
xor ( \5502_b0 , \5501_b0 , w_13598 );
not ( w_13598 , w_13599 );
and ( w_13599 , w_13596 , w_13597 );
buf ( w_13596 , \1835_b1 );
not ( w_13596 , w_13600 );
not ( w_13597 , w_13601 );
and ( w_13600 , w_13601 , \1835_b0 );
or ( \5503_b1 , \5500_b1 , \5502_b1 );
not ( \5502_b1 , w_13602 );
and ( \5503_b0 , \5500_b0 , w_13603 );
and ( w_13602 , w_13603 , \5502_b0 );
or ( \5504_b1 , \5496_b1 , \5503_b1 );
not ( \5503_b1 , w_13604 );
and ( \5504_b0 , \5496_b0 , w_13605 );
and ( w_13604 , w_13605 , \5503_b0 );
or ( \5505_b1 , \2850_b1 , \1955_b1 );
not ( \1955_b1 , w_13606 );
and ( \5505_b0 , \2850_b0 , w_13607 );
and ( w_13606 , w_13607 , \1955_b0 );
or ( \5506_b1 , \2763_b1 , \1953_b1 );
not ( \1953_b1 , w_13608 );
and ( \5506_b0 , \2763_b0 , w_13609 );
and ( w_13608 , w_13609 , \1953_b0 );
or ( \5507_b1 , \5505_b1 , w_13611 );
not ( w_13611 , w_13612 );
and ( \5507_b0 , \5505_b0 , w_13613 );
and ( w_13612 ,  , w_13613 );
buf ( w_13611 , \5506_b1 );
not ( w_13611 , w_13614 );
not (  , w_13615 );
and ( w_13614 , w_13615 , \5506_b0 );
or ( \5508_b1 , \5507_b1 , w_13616 );
xor ( \5508_b0 , \5507_b0 , w_13618 );
not ( w_13618 , w_13619 );
and ( w_13619 , w_13616 , w_13617 );
buf ( w_13616 , \1835_b1 );
not ( w_13616 , w_13620 );
not ( w_13617 , w_13621 );
and ( w_13620 , w_13621 , \1835_b0 );
or ( \5509_b1 , \5503_b1 , \5508_b1 );
not ( \5508_b1 , w_13622 );
and ( \5509_b0 , \5503_b0 , w_13623 );
and ( w_13622 , w_13623 , \5508_b0 );
or ( \5510_b1 , \5496_b1 , \5508_b1 );
not ( \5508_b1 , w_13624 );
and ( \5510_b0 , \5496_b0 , w_13625 );
and ( w_13624 , w_13625 , \5508_b0 );
or ( \5512_b1 , \5465_b1 , \5467_b1 );
xor ( \5512_b0 , \5465_b0 , w_13626 );
not ( w_13626 , w_13627 );
and ( w_13627 , \5467_b1 , \5467_b0 );
or ( \5513_b1 , \5512_b1 , \5470_b1 );
xor ( \5513_b0 , \5512_b0 , w_13628 );
not ( w_13628 , w_13629 );
and ( w_13629 , \5470_b1 , \5470_b0 );
or ( \5514_b1 , \5511_b1 , \5513_b1 );
not ( \5513_b1 , w_13630 );
and ( \5514_b0 , \5511_b0 , w_13631 );
and ( w_13630 , w_13631 , \5513_b0 );
or ( \5515_b1 , \5484_b1 , \5514_b1 );
not ( \5514_b1 , w_13632 );
and ( \5515_b0 , \5484_b0 , w_13633 );
and ( w_13632 , w_13633 , \5514_b0 );
or ( \5516_b1 , \5484_b1 , \5514_b1 );
xor ( \5516_b0 , \5484_b0 , w_13634 );
not ( w_13634 , w_13635 );
and ( w_13635 , \5514_b1 , \5514_b0 );
or ( \5517_b1 , \5511_b1 , \5513_b1 );
xor ( \5517_b0 , \5511_b0 , w_13636 );
not ( w_13636 , w_13637 );
and ( w_13637 , \5513_b1 , \5513_b0 );
or ( \5518_b1 , \5453_b1 , \5457_b1 );
xor ( \5518_b0 , \5453_b0 , w_13638 );
not ( w_13638 , w_13639 );
and ( w_13639 , \5457_b1 , \5457_b0 );
or ( \5519_b1 , \5518_b1 , \5462_b1 );
xor ( \5519_b0 , \5518_b0 , w_13640 );
not ( w_13640 , w_13641 );
and ( w_13641 , \5462_b1 , \5462_b0 );
or ( \5520_b1 , \5496_b1 , \5503_b1 );
xor ( \5520_b0 , \5496_b0 , w_13642 );
not ( w_13642 , w_13643 );
and ( w_13643 , \5503_b1 , \5503_b0 );
or ( \5521_b1 , \5520_b1 , \5508_b1 );
xor ( \5521_b0 , \5520_b0 , w_13644 );
not ( w_13644 , w_13645 );
and ( w_13645 , \5508_b1 , \5508_b0 );
or ( \5522_b1 , \5519_b1 , \5521_b1 );
not ( \5521_b1 , w_13646 );
and ( \5522_b0 , \5519_b0 , w_13647 );
and ( w_13646 , w_13647 , \5521_b0 );
or ( \5523_b1 , \5517_b1 , \5522_b1 );
not ( \5522_b1 , w_13648 );
and ( \5523_b0 , \5517_b0 , w_13649 );
and ( w_13648 , w_13649 , \5522_b0 );
or ( \5524_b1 , \5517_b1 , \5522_b1 );
xor ( \5524_b0 , \5517_b0 , w_13650 );
not ( w_13650 , w_13651 );
and ( w_13651 , \5522_b1 , \5522_b0 );
or ( \5525_b1 , \5519_b1 , \5521_b1 );
xor ( \5525_b0 , \5519_b0 , w_13652 );
not ( w_13652 , w_13653 );
and ( w_13653 , \5521_b1 , \5521_b0 );
or ( \5526_b1 , \2305_b1 , \2913_b1 );
not ( \2913_b1 , w_13654 );
and ( \5526_b0 , \2305_b0 , w_13655 );
and ( w_13654 , w_13655 , \2913_b0 );
or ( \5527_b1 , \2161_b1 , \2910_b1 );
not ( \2910_b1 , w_13656 );
and ( \5527_b0 , \2161_b0 , w_13657 );
and ( w_13656 , w_13657 , \2910_b0 );
or ( \5528_b1 , \5526_b1 , w_13659 );
not ( w_13659 , w_13660 );
and ( \5528_b0 , \5526_b0 , w_13661 );
and ( w_13660 ,  , w_13661 );
buf ( w_13659 , \5527_b1 );
not ( w_13659 , w_13662 );
not (  , w_13663 );
and ( w_13662 , w_13663 , \5527_b0 );
or ( \5529_b1 , \5528_b1 , w_13664 );
xor ( \5529_b0 , \5528_b0 , w_13666 );
not ( w_13666 , w_13667 );
and ( w_13667 , w_13664 , w_13665 );
buf ( w_13664 , \2371_b1 );
not ( w_13664 , w_13668 );
not ( w_13665 , w_13669 );
and ( w_13668 , w_13669 , \2371_b0 );
or ( \5530_b1 , \2541_b1 , \2550_b1 );
not ( \2550_b1 , w_13670 );
and ( \5530_b0 , \2541_b0 , w_13671 );
and ( w_13670 , w_13671 , \2550_b0 );
or ( \5531_b1 , \2532_b1 , \2548_b1 );
not ( \2548_b1 , w_13672 );
and ( \5531_b0 , \2532_b0 , w_13673 );
and ( w_13672 , w_13673 , \2548_b0 );
or ( \5532_b1 , \5530_b1 , w_13675 );
not ( w_13675 , w_13676 );
and ( \5532_b0 , \5530_b0 , w_13677 );
and ( w_13676 ,  , w_13677 );
buf ( w_13675 , \5531_b1 );
not ( w_13675 , w_13678 );
not (  , w_13679 );
and ( w_13678 , w_13679 , \5531_b0 );
or ( \5533_b1 , \5532_b1 , w_13680 );
xor ( \5533_b0 , \5532_b0 , w_13682 );
not ( w_13682 , w_13683 );
and ( w_13683 , w_13680 , w_13681 );
buf ( w_13680 , \2374_b1 );
not ( w_13680 , w_13684 );
not ( w_13681 , w_13685 );
and ( w_13684 , w_13685 , \2374_b0 );
or ( \5534_b1 , \5529_b1 , \5533_b1 );
not ( \5533_b1 , w_13686 );
and ( \5534_b0 , \5529_b0 , w_13687 );
and ( w_13686 , w_13687 , \5533_b0 );
or ( \5535_b1 , \2850_b1 , \2261_b1 );
not ( \2261_b1 , w_13688 );
and ( \5535_b0 , \2850_b0 , w_13689 );
and ( w_13688 , w_13689 , \2261_b0 );
or ( \5536_b1 , \2763_b1 , \2259_b1 );
not ( \2259_b1 , w_13690 );
and ( \5536_b0 , \2763_b0 , w_13691 );
and ( w_13690 , w_13691 , \2259_b0 );
or ( \5537_b1 , \5535_b1 , w_13693 );
not ( w_13693 , w_13694 );
and ( \5537_b0 , \5535_b0 , w_13695 );
and ( w_13694 ,  , w_13695 );
buf ( w_13693 , \5536_b1 );
not ( w_13693 , w_13696 );
not (  , w_13697 );
and ( w_13696 , w_13697 , \5536_b0 );
or ( \5538_b1 , \5537_b1 , w_13698 );
xor ( \5538_b0 , \5537_b0 , w_13700 );
not ( w_13700 , w_13701 );
and ( w_13701 , w_13698 , w_13699 );
buf ( w_13698 , \2124_b1 );
not ( w_13698 , w_13702 );
not ( w_13699 , w_13703 );
and ( w_13702 , w_13703 , \2124_b0 );
or ( \5539_b1 , \5533_b1 , \5538_b1 );
not ( \5538_b1 , w_13704 );
and ( \5539_b0 , \5533_b0 , w_13705 );
and ( w_13704 , w_13705 , \5538_b0 );
or ( \5540_b1 , \5529_b1 , \5538_b1 );
not ( \5538_b1 , w_13706 );
and ( \5540_b0 , \5529_b0 , w_13707 );
and ( w_13706 , w_13707 , \5538_b0 );
or ( \5542_b1 , \5488_b1 , \5492_b1 );
xor ( \5542_b0 , \5488_b0 , w_13708 );
not ( w_13708 , w_13709 );
and ( w_13709 , \5492_b1 , \5492_b0 );
or ( \5543_b1 , \5542_b1 , \1835_b1 );
xor ( \5543_b0 , \5542_b0 , w_13710 );
not ( w_13710 , w_13711 );
and ( w_13711 , \1835_b1 , \1835_b0 );
or ( \5544_b1 , \5541_b1 , \5543_b1 );
not ( \5543_b1 , w_13712 );
and ( \5544_b0 , \5541_b0 , w_13713 );
and ( w_13712 , w_13713 , \5543_b0 );
or ( \5545_b1 , \5500_b1 , \5502_b1 );
xor ( \5545_b0 , \5500_b0 , w_13714 );
not ( w_13714 , w_13715 );
and ( w_13715 , \5502_b1 , \5502_b0 );
or ( \5546_b1 , \5543_b1 , \5545_b1 );
not ( \5545_b1 , w_13716 );
and ( \5546_b0 , \5543_b0 , w_13717 );
and ( w_13716 , w_13717 , \5545_b0 );
or ( \5547_b1 , \5541_b1 , \5545_b1 );
not ( \5545_b1 , w_13718 );
and ( \5547_b0 , \5541_b0 , w_13719 );
and ( w_13718 , w_13719 , \5545_b0 );
or ( \5549_b1 , \5525_b1 , \5548_b1 );
not ( \5548_b1 , w_13720 );
and ( \5549_b0 , \5525_b0 , w_13721 );
and ( w_13720 , w_13721 , \5548_b0 );
or ( \5550_b1 , \5525_b1 , \5548_b1 );
xor ( \5550_b0 , \5525_b0 , w_13722 );
not ( w_13722 , w_13723 );
and ( w_13723 , \5548_b1 , \5548_b0 );
or ( \5551_b1 , \5541_b1 , \5543_b1 );
xor ( \5551_b0 , \5541_b0 , w_13724 );
not ( w_13724 , w_13725 );
and ( w_13725 , \5543_b1 , \5543_b0 );
or ( \5552_b1 , \5551_b1 , \5545_b1 );
xor ( \5552_b0 , \5551_b0 , w_13726 );
not ( w_13726 , w_13727 );
and ( w_13727 , \5545_b1 , \5545_b0 );
or ( \5553_b1 , \2532_b1 , \2913_b1 );
not ( \2913_b1 , w_13728 );
and ( \5553_b0 , \2532_b0 , w_13729 );
and ( w_13728 , w_13729 , \2913_b0 );
or ( \5554_b1 , \2305_b1 , \2910_b1 );
not ( \2910_b1 , w_13730 );
and ( \5554_b0 , \2305_b0 , w_13731 );
and ( w_13730 , w_13731 , \2910_b0 );
or ( \5555_b1 , \5553_b1 , w_13733 );
not ( w_13733 , w_13734 );
and ( \5555_b0 , \5553_b0 , w_13735 );
and ( w_13734 ,  , w_13735 );
buf ( w_13733 , \5554_b1 );
not ( w_13733 , w_13736 );
not (  , w_13737 );
and ( w_13736 , w_13737 , \5554_b0 );
or ( \5556_b1 , \5555_b1 , w_13738 );
xor ( \5556_b0 , \5555_b0 , w_13740 );
not ( w_13740 , w_13741 );
and ( w_13741 , w_13738 , w_13739 );
buf ( w_13738 , \2371_b1 );
not ( w_13738 , w_13742 );
not ( w_13739 , w_13743 );
and ( w_13742 , w_13743 , \2371_b0 );
or ( \5557_b1 , \2763_b1 , \2550_b1 );
not ( \2550_b1 , w_13744 );
and ( \5557_b0 , \2763_b0 , w_13745 );
and ( w_13744 , w_13745 , \2550_b0 );
or ( \5558_b1 , \2541_b1 , \2548_b1 );
not ( \2548_b1 , w_13746 );
and ( \5558_b0 , \2541_b0 , w_13747 );
and ( w_13746 , w_13747 , \2548_b0 );
or ( \5559_b1 , \5557_b1 , w_13749 );
not ( w_13749 , w_13750 );
and ( \5559_b0 , \5557_b0 , w_13751 );
and ( w_13750 ,  , w_13751 );
buf ( w_13749 , \5558_b1 );
not ( w_13749 , w_13752 );
not (  , w_13753 );
and ( w_13752 , w_13753 , \5558_b0 );
or ( \5560_b1 , \5559_b1 , w_13754 );
xor ( \5560_b0 , \5559_b0 , w_13756 );
not ( w_13756 , w_13757 );
and ( w_13757 , w_13754 , w_13755 );
buf ( w_13754 , \2374_b1 );
not ( w_13754 , w_13758 );
not ( w_13755 , w_13759 );
and ( w_13758 , w_13759 , \2374_b0 );
or ( \5561_b1 , \5556_b1 , \5560_b1 );
not ( \5560_b1 , w_13760 );
and ( \5561_b0 , \5556_b0 , w_13761 );
and ( w_13760 , w_13761 , \5560_b0 );
or ( \5562_b1 , \5560_b1 , \2124_b1 );
not ( \2124_b1 , w_13762 );
and ( \5562_b0 , \5560_b0 , w_13763 );
and ( w_13762 , w_13763 , \2124_b0 );
or ( \5563_b1 , \5556_b1 , \2124_b1 );
not ( \2124_b1 , w_13764 );
and ( \5563_b0 , \5556_b0 , w_13765 );
and ( w_13764 , w_13765 , \2124_b0 );
or ( \5565_b1 , \5529_b1 , \5533_b1 );
xor ( \5565_b0 , \5529_b0 , w_13766 );
not ( w_13766 , w_13767 );
and ( w_13767 , \5533_b1 , \5533_b0 );
or ( \5566_b1 , \5565_b1 , \5538_b1 );
xor ( \5566_b0 , \5565_b0 , w_13768 );
not ( w_13768 , w_13769 );
and ( w_13769 , \5538_b1 , \5538_b0 );
or ( \5567_b1 , \5564_b1 , \5566_b1 );
not ( \5566_b1 , w_13770 );
and ( \5567_b0 , \5564_b0 , w_13771 );
and ( w_13770 , w_13771 , \5566_b0 );
or ( \5568_b1 , \5552_b1 , \5567_b1 );
not ( \5567_b1 , w_13772 );
and ( \5568_b0 , \5552_b0 , w_13773 );
and ( w_13772 , w_13773 , \5567_b0 );
or ( \5569_b1 , \5552_b1 , \5567_b1 );
xor ( \5569_b0 , \5552_b0 , w_13774 );
not ( w_13774 , w_13775 );
and ( w_13775 , \5567_b1 , \5567_b0 );
or ( \5570_b1 , \5564_b1 , \5566_b1 );
xor ( \5570_b0 , \5564_b0 , w_13776 );
not ( w_13776 , w_13777 );
and ( w_13777 , \5566_b1 , \5566_b0 );
or ( \5571_b1 , \2850_b1 , w_13779 );
not ( w_13779 , w_13780 );
and ( \5571_b0 , \2850_b0 , w_13781 );
and ( w_13780 ,  , w_13781 );
buf ( w_13779 , \2259_b1 );
not ( w_13779 , w_13782 );
not (  , w_13783 );
and ( w_13782 , w_13783 , \2259_b0 );
or ( \5572_b1 , \5571_b1 , w_13784 );
xor ( \5572_b0 , \5571_b0 , w_13786 );
not ( w_13786 , w_13787 );
and ( w_13787 , w_13784 , w_13785 );
buf ( w_13784 , \2124_b1 );
not ( w_13784 , w_13788 );
not ( w_13785 , w_13789 );
and ( w_13788 , w_13789 , \2124_b0 );
or ( \5573_b1 , \5556_b1 , \5560_b1 );
xor ( \5573_b0 , \5556_b0 , w_13790 );
not ( w_13790 , w_13791 );
and ( w_13791 , \5560_b1 , \5560_b0 );
or ( \5574_b1 , \5573_b1 , \2124_b1 );
xor ( \5574_b0 , \5573_b0 , w_13792 );
not ( w_13792 , w_13793 );
and ( w_13793 , \2124_b1 , \2124_b0 );
or ( \5575_b1 , \5572_b1 , \5574_b1 );
not ( \5574_b1 , w_13794 );
and ( \5575_b0 , \5572_b0 , w_13795 );
and ( w_13794 , w_13795 , \5574_b0 );
or ( \5576_b1 , \5570_b1 , \5575_b1 );
not ( \5575_b1 , w_13796 );
and ( \5576_b0 , \5570_b0 , w_13797 );
and ( w_13796 , w_13797 , \5575_b0 );
or ( \5577_b1 , \5570_b1 , \5575_b1 );
xor ( \5577_b0 , \5570_b0 , w_13798 );
not ( w_13798 , w_13799 );
and ( w_13799 , \5575_b1 , \5575_b0 );
or ( \5578_b1 , \5572_b1 , \5574_b1 );
xor ( \5578_b0 , \5572_b0 , w_13800 );
not ( w_13800 , w_13801 );
and ( w_13801 , \5574_b1 , \5574_b0 );
or ( \5579_b1 , \2541_b1 , \2913_b1 );
not ( \2913_b1 , w_13802 );
and ( \5579_b0 , \2541_b0 , w_13803 );
and ( w_13802 , w_13803 , \2913_b0 );
or ( \5580_b1 , \2532_b1 , \2910_b1 );
not ( \2910_b1 , w_13804 );
and ( \5580_b0 , \2532_b0 , w_13805 );
and ( w_13804 , w_13805 , \2910_b0 );
or ( \5581_b1 , \5579_b1 , w_13807 );
not ( w_13807 , w_13808 );
and ( \5581_b0 , \5579_b0 , w_13809 );
and ( w_13808 ,  , w_13809 );
buf ( w_13807 , \5580_b1 );
not ( w_13807 , w_13810 );
not (  , w_13811 );
and ( w_13810 , w_13811 , \5580_b0 );
or ( \5582_b1 , \5581_b1 , w_13812 );
xor ( \5582_b0 , \5581_b0 , w_13814 );
not ( w_13814 , w_13815 );
and ( w_13815 , w_13812 , w_13813 );
buf ( w_13812 , \2371_b1 );
not ( w_13812 , w_13816 );
not ( w_13813 , w_13817 );
and ( w_13816 , w_13817 , \2371_b0 );
or ( \5583_b1 , \2850_b1 , \2550_b1 );
not ( \2550_b1 , w_13818 );
and ( \5583_b0 , \2850_b0 , w_13819 );
and ( w_13818 , w_13819 , \2550_b0 );
or ( \5584_b1 , \2763_b1 , \2548_b1 );
not ( \2548_b1 , w_13820 );
and ( \5584_b0 , \2763_b0 , w_13821 );
and ( w_13820 , w_13821 , \2548_b0 );
or ( \5585_b1 , \5583_b1 , w_13823 );
not ( w_13823 , w_13824 );
and ( \5585_b0 , \5583_b0 , w_13825 );
and ( w_13824 ,  , w_13825 );
buf ( w_13823 , \5584_b1 );
not ( w_13823 , w_13826 );
not (  , w_13827 );
and ( w_13826 , w_13827 , \5584_b0 );
or ( \5586_b1 , \5585_b1 , w_13828 );
xor ( \5586_b0 , \5585_b0 , w_13830 );
not ( w_13830 , w_13831 );
and ( w_13831 , w_13828 , w_13829 );
buf ( w_13828 , \2374_b1 );
not ( w_13828 , w_13832 );
not ( w_13829 , w_13833 );
and ( w_13832 , w_13833 , \2374_b0 );
or ( \5587_b1 , \5582_b1 , \5586_b1 );
not ( \5586_b1 , w_13834 );
and ( \5587_b0 , \5582_b0 , w_13835 );
and ( w_13834 , w_13835 , \5586_b0 );
or ( \5588_b1 , \5578_b1 , \5587_b1 );
not ( \5587_b1 , w_13836 );
and ( \5588_b0 , \5578_b0 , w_13837 );
and ( w_13836 , w_13837 , \5587_b0 );
or ( \5589_b1 , \5578_b1 , \5587_b1 );
xor ( \5589_b0 , \5578_b0 , w_13838 );
not ( w_13838 , w_13839 );
and ( w_13839 , \5587_b1 , \5587_b0 );
or ( \5590_b1 , \5582_b1 , \5586_b1 );
xor ( \5590_b0 , \5582_b0 , w_13840 );
not ( w_13840 , w_13841 );
and ( w_13841 , \5586_b1 , \5586_b0 );
or ( \5591_b1 , \2763_b1 , \2913_b1 );
not ( \2913_b1 , w_13842 );
and ( \5591_b0 , \2763_b0 , w_13843 );
and ( w_13842 , w_13843 , \2913_b0 );
or ( \5592_b1 , \2541_b1 , \2910_b1 );
not ( \2910_b1 , w_13844 );
and ( \5592_b0 , \2541_b0 , w_13845 );
and ( w_13844 , w_13845 , \2910_b0 );
or ( \5593_b1 , \5591_b1 , w_13847 );
not ( w_13847 , w_13848 );
and ( \5593_b0 , \5591_b0 , w_13849 );
and ( w_13848 ,  , w_13849 );
buf ( w_13847 , \5592_b1 );
not ( w_13847 , w_13850 );
not (  , w_13851 );
and ( w_13850 , w_13851 , \5592_b0 );
or ( \5594_b1 , \5593_b1 , w_13852 );
xor ( \5594_b0 , \5593_b0 , w_13854 );
not ( w_13854 , w_13855 );
and ( w_13855 , w_13852 , w_13853 );
buf ( w_13852 , \2371_b1 );
not ( w_13852 , w_13856 );
not ( w_13853 , w_13857 );
and ( w_13856 , w_13857 , \2371_b0 );
or ( \5595_b1 , \5594_b1 , \2374_b1 );
not ( \2374_b1 , w_13858 );
and ( \5595_b0 , \5594_b0 , w_13859 );
and ( w_13858 , w_13859 , \2374_b0 );
or ( \5596_b1 , \5590_b1 , \5595_b1 );
not ( \5595_b1 , w_13860 );
and ( \5596_b0 , \5590_b0 , w_13861 );
and ( w_13860 , w_13861 , \5595_b0 );
or ( \5597_b1 , \5590_b1 , \5595_b1 );
xor ( \5597_b0 , \5590_b0 , w_13862 );
not ( w_13862 , w_13863 );
and ( w_13863 , \5595_b1 , \5595_b0 );
or ( \5598_b1 , \2850_b1 , w_13865 );
not ( w_13865 , w_13866 );
and ( \5598_b0 , \2850_b0 , w_13867 );
and ( w_13866 ,  , w_13867 );
buf ( w_13865 , \2548_b1 );
not ( w_13865 , w_13868 );
not (  , w_13869 );
and ( w_13868 , w_13869 , \2548_b0 );
or ( \5599_b1 , \5598_b1 , w_13870 );
xor ( \5599_b0 , \5598_b0 , w_13872 );
not ( w_13872 , w_13873 );
and ( w_13873 , w_13870 , w_13871 );
buf ( w_13870 , \2374_b1 );
not ( w_13870 , w_13874 );
not ( w_13871 , w_13875 );
and ( w_13874 , w_13875 , \2374_b0 );
or ( \5600_b1 , \5594_b1 , \2374_b1 );
xor ( \5600_b0 , \5594_b0 , w_13876 );
not ( w_13876 , w_13877 );
and ( w_13877 , \2374_b1 , \2374_b0 );
or ( \5601_b1 , \5599_b1 , \5600_b1 );
not ( \5600_b1 , w_13878 );
and ( \5601_b0 , \5599_b0 , w_13879 );
and ( w_13878 , w_13879 , \5600_b0 );
or ( \5602_b1 , \5599_b1 , \5600_b1 );
xor ( \5602_b0 , \5599_b0 , w_13880 );
not ( w_13880 , w_13881 );
and ( w_13881 , \5600_b1 , \5600_b0 );
or ( \5603_b1 , \2850_b1 , \2913_b1 );
not ( \2913_b1 , w_13882 );
and ( \5603_b0 , \2850_b0 , w_13883 );
and ( w_13882 , w_13883 , \2913_b0 );
or ( \5604_b1 , \2763_b1 , \2910_b1 );
not ( \2910_b1 , w_13884 );
and ( \5604_b0 , \2763_b0 , w_13885 );
and ( w_13884 , w_13885 , \2910_b0 );
or ( \5605_b1 , \5603_b1 , w_13887 );
not ( w_13887 , w_13888 );
and ( \5605_b0 , \5603_b0 , w_13889 );
and ( w_13888 ,  , w_13889 );
buf ( w_13887 , \5604_b1 );
not ( w_13887 , w_13890 );
not (  , w_13891 );
and ( w_13890 , w_13891 , \5604_b0 );
or ( \5606_b1 , \5605_b1 , w_13892 );
xor ( \5606_b0 , \5605_b0 , w_13894 );
not ( w_13894 , w_13895 );
and ( w_13895 , w_13892 , w_13893 );
buf ( w_13892 , \2371_b1 );
not ( w_13892 , w_13896 );
not ( w_13893 , w_13897 );
and ( w_13896 , w_13897 , \2371_b0 );
or ( \5607_b1 , \2850_b1 , w_13899 );
not ( w_13899 , w_13900 );
and ( \5607_b0 , \2850_b0 , w_13901 );
and ( w_13900 ,  , w_13901 );
buf ( w_13899 , \2910_b1 );
not ( w_13899 , w_13902 );
not (  , w_13903 );
and ( w_13902 , w_13903 , \2910_b0 );
or ( \5608_b1 , \5607_b1 , w_13904 );
xor ( \5608_b0 , \5607_b0 , w_13906 );
not ( w_13906 , w_13907 );
and ( w_13907 , w_13904 , w_13905 );
buf ( w_13904 , \2371_b1 );
not ( w_13904 , w_13908 );
not ( w_13905 , w_13909 );
and ( w_13908 , w_13909 , \2371_b0 );
or ( \5609_b1 , \5608_b1 , \2371_b1 );
not ( \2371_b1 , w_13910 );
and ( \5609_b0 , \5608_b0 , w_13911 );
and ( w_13910 , w_13911 , \2371_b0 );
or ( \5610_b1 , \5606_b1 , \5609_b1 );
not ( \5609_b1 , w_13912 );
and ( \5610_b0 , \5606_b0 , w_13913 );
and ( w_13912 , w_13913 , \5609_b0 );
or ( \5611_b1 , \5602_b1 , \5610_b1 );
not ( \5610_b1 , w_13914 );
and ( \5611_b0 , \5602_b0 , w_13915 );
and ( w_13914 , w_13915 , \5610_b0 );
or ( \5612_b1 , \5601_b1 , w_13916 );
or ( \5612_b0 , \5601_b0 , \5611_b0 );
not ( \5611_b0 , w_13917 );
and ( w_13917 , w_13916 , \5611_b1 );
or ( \5613_b1 , \5597_b1 , \5612_b1 );
not ( \5612_b1 , w_13918 );
and ( \5613_b0 , \5597_b0 , w_13919 );
and ( w_13918 , w_13919 , \5612_b0 );
or ( \5614_b1 , \5596_b1 , w_13920 );
or ( \5614_b0 , \5596_b0 , \5613_b0 );
not ( \5613_b0 , w_13921 );
and ( w_13921 , w_13920 , \5613_b1 );
or ( \5615_b1 , \5589_b1 , \5614_b1 );
not ( \5614_b1 , w_13922 );
and ( \5615_b0 , \5589_b0 , w_13923 );
and ( w_13922 , w_13923 , \5614_b0 );
or ( \5616_b1 , \5588_b1 , w_13924 );
or ( \5616_b0 , \5588_b0 , \5615_b0 );
not ( \5615_b0 , w_13925 );
and ( w_13925 , w_13924 , \5615_b1 );
or ( \5617_b1 , \5577_b1 , \5616_b1 );
not ( \5616_b1 , w_13926 );
and ( \5617_b0 , \5577_b0 , w_13927 );
and ( w_13926 , w_13927 , \5616_b0 );
or ( \5618_b1 , \5576_b1 , w_13928 );
or ( \5618_b0 , \5576_b0 , \5617_b0 );
not ( \5617_b0 , w_13929 );
and ( w_13929 , w_13928 , \5617_b1 );
or ( \5619_b1 , \5569_b1 , \5618_b1 );
not ( \5618_b1 , w_13930 );
and ( \5619_b0 , \5569_b0 , w_13931 );
and ( w_13930 , w_13931 , \5618_b0 );
or ( \5620_b1 , \5568_b1 , w_13932 );
or ( \5620_b0 , \5568_b0 , \5619_b0 );
not ( \5619_b0 , w_13933 );
and ( w_13933 , w_13932 , \5619_b1 );
or ( \5621_b1 , \5550_b1 , \5620_b1 );
not ( \5620_b1 , w_13934 );
and ( \5621_b0 , \5550_b0 , w_13935 );
and ( w_13934 , w_13935 , \5620_b0 );
or ( \5622_b1 , \5549_b1 , w_13936 );
or ( \5622_b0 , \5549_b0 , \5621_b0 );
not ( \5621_b0 , w_13937 );
and ( w_13937 , w_13936 , \5621_b1 );
or ( \5623_b1 , \5524_b1 , \5622_b1 );
not ( \5622_b1 , w_13938 );
and ( \5623_b0 , \5524_b0 , w_13939 );
and ( w_13938 , w_13939 , \5622_b0 );
or ( \5624_b1 , \5523_b1 , w_13940 );
or ( \5624_b0 , \5523_b0 , \5623_b0 );
not ( \5623_b0 , w_13941 );
and ( w_13941 , w_13940 , \5623_b1 );
or ( \5625_b1 , \5516_b1 , \5624_b1 );
not ( \5624_b1 , w_13942 );
and ( \5625_b0 , \5516_b0 , w_13943 );
and ( w_13942 , w_13943 , \5624_b0 );
or ( \5626_b1 , \5515_b1 , w_13944 );
or ( \5626_b0 , \5515_b0 , \5625_b0 );
not ( \5625_b0 , w_13945 );
and ( w_13945 , w_13944 , \5625_b1 );
or ( \5627_b1 , \5482_b1 , \5626_b1 );
not ( \5626_b1 , w_13946 );
and ( \5627_b0 , \5482_b0 , w_13947 );
and ( w_13946 , w_13947 , \5626_b0 );
or ( \5628_b1 , \5481_b1 , w_13948 );
or ( \5628_b0 , \5481_b0 , \5627_b0 );
not ( \5627_b0 , w_13949 );
and ( w_13949 , w_13948 , \5627_b1 );
or ( \5629_b1 , \5448_b1 , \5628_b1 );
not ( \5628_b1 , w_13950 );
and ( \5629_b0 , \5448_b0 , w_13951 );
and ( w_13950 , w_13951 , \5628_b0 );
or ( \5630_b1 , \5447_b1 , w_13952 );
or ( \5630_b0 , \5447_b0 , \5629_b0 );
not ( \5629_b0 , w_13953 );
and ( w_13953 , w_13952 , \5629_b1 );
or ( \5631_b1 , \5440_b1 , \5630_b1 );
not ( \5630_b1 , w_13954 );
and ( \5631_b0 , \5440_b0 , w_13955 );
and ( w_13954 , w_13955 , \5630_b0 );
or ( \5632_b1 , \5439_b1 , w_13956 );
or ( \5632_b0 , \5439_b0 , \5631_b0 );
not ( \5631_b0 , w_13957 );
and ( w_13957 , w_13956 , \5631_b1 );
or ( \5633_b1 , \5387_b1 , \5632_b1 );
not ( \5632_b1 , w_13958 );
and ( \5633_b0 , \5387_b0 , w_13959 );
and ( w_13958 , w_13959 , \5632_b0 );
or ( \5634_b1 , \5386_b1 , w_13960 );
or ( \5634_b0 , \5386_b0 , \5633_b0 );
not ( \5633_b0 , w_13961 );
and ( w_13961 , w_13960 , \5633_b1 );
or ( \5635_b1 , \5348_b1 , \5634_b1 );
not ( \5634_b1 , w_13962 );
and ( \5635_b0 , \5348_b0 , w_13963 );
and ( w_13962 , w_13963 , \5634_b0 );
or ( \5636_b1 , \5347_b1 , w_13964 );
or ( \5636_b0 , \5347_b0 , \5635_b0 );
not ( \5635_b0 , w_13965 );
and ( w_13965 , w_13964 , \5635_b1 );
or ( \5637_b1 , \5295_b1 , \5636_b1 );
not ( \5636_b1 , w_13966 );
and ( \5637_b0 , \5295_b0 , w_13967 );
and ( w_13966 , w_13967 , \5636_b0 );
or ( \5638_b1 , \5294_b1 , w_13968 );
or ( \5638_b0 , \5294_b0 , \5637_b0 );
not ( \5637_b0 , w_13969 );
and ( w_13969 , w_13968 , \5637_b1 );
or ( \5639_b1 , \5224_b1 , \5638_b1 );
not ( \5638_b1 , w_13970 );
and ( \5639_b0 , \5224_b0 , w_13971 );
and ( w_13970 , w_13971 , \5638_b0 );
or ( \5640_b1 , \5223_b1 , w_13972 );
or ( \5640_b0 , \5223_b0 , \5639_b0 );
not ( \5639_b0 , w_13973 );
and ( w_13973 , w_13972 , \5639_b1 );
or ( \5641_b1 , \5169_b1 , \5640_b1 );
not ( \5640_b1 , w_13974 );
and ( \5641_b0 , \5169_b0 , w_13975 );
and ( w_13974 , w_13975 , \5640_b0 );
or ( \5642_b1 , \5168_b1 , w_13976 );
or ( \5642_b0 , \5168_b0 , \5641_b0 );
not ( \5641_b0 , w_13977 );
and ( w_13977 , w_13976 , \5641_b1 );
or ( \5643_b1 , \5110_b1 , \5642_b1 );
not ( \5642_b1 , w_13978 );
and ( \5643_b0 , \5110_b0 , w_13979 );
and ( w_13978 , w_13979 , \5642_b0 );
or ( \5644_b1 , \5109_b1 , w_13980 );
or ( \5644_b0 , \5109_b0 , \5643_b0 );
not ( \5643_b0 , w_13981 );
and ( w_13981 , w_13980 , \5643_b1 );
or ( \5645_b1 , \5102_b1 , \5644_b1 );
not ( \5644_b1 , w_13982 );
and ( \5645_b0 , \5102_b0 , w_13983 );
and ( w_13982 , w_13983 , \5644_b0 );
or ( \5646_b1 , \5101_b1 , w_13984 );
or ( \5646_b0 , \5101_b0 , \5645_b0 );
not ( \5645_b0 , w_13985 );
and ( w_13985 , w_13984 , \5645_b1 );
or ( \5647_b1 , \5023_b1 , \5646_b1 );
not ( \5646_b1 , w_13986 );
and ( \5647_b0 , \5023_b0 , w_13987 );
and ( w_13986 , w_13987 , \5646_b0 );
or ( \5648_b1 , \5022_b1 , w_13988 );
or ( \5648_b0 , \5022_b0 , \5647_b0 );
not ( \5647_b0 , w_13989 );
and ( w_13989 , w_13988 , \5647_b1 );
or ( \5649_b1 , \4943_b1 , \5648_b1 );
not ( \5648_b1 , w_13990 );
and ( \5649_b0 , \4943_b0 , w_13991 );
and ( w_13990 , w_13991 , \5648_b0 );
or ( \5650_b1 , \4942_b1 , w_13992 );
or ( \5650_b0 , \4942_b0 , \5649_b0 );
not ( \5649_b0 , w_13993 );
and ( w_13993 , w_13992 , \5649_b1 );
or ( \5651_b1 , \4848_b1 , \5650_b1 );
not ( \5650_b1 , w_13994 );
and ( \5651_b0 , \4848_b0 , w_13995 );
and ( w_13994 , w_13995 , \5650_b0 );
or ( \5652_b1 , \4847_b1 , w_13996 );
or ( \5652_b0 , \4847_b0 , \5651_b0 );
not ( \5651_b0 , w_13997 );
and ( w_13997 , w_13996 , \5651_b1 );
or ( \5653_b1 , \4760_b1 , \5652_b1 );
not ( \5652_b1 , w_13998 );
and ( \5653_b0 , \4760_b0 , w_13999 );
and ( w_13998 , w_13999 , \5652_b0 );
or ( \5654_b1 , \4759_b1 , w_14000 );
or ( \5654_b0 , \4759_b0 , \5653_b0 );
not ( \5653_b0 , w_14001 );
and ( w_14001 , w_14000 , \5653_b1 );
or ( \5655_b1 , \4668_b1 , \5654_b1 );
not ( \5654_b1 , w_14002 );
and ( \5655_b0 , \4668_b0 , w_14003 );
and ( w_14002 , w_14003 , \5654_b0 );
or ( \5656_b1 , \4667_b1 , w_14004 );
or ( \5656_b0 , \4667_b0 , \5655_b0 );
not ( \5655_b0 , w_14005 );
and ( w_14005 , w_14004 , \5655_b1 );
or ( \5657_b1 , \4580_b1 , \5656_b1 );
not ( \5656_b1 , w_14006 );
and ( \5657_b0 , \4580_b0 , w_14007 );
and ( w_14006 , w_14007 , \5656_b0 );
or ( \5658_b1 , \4579_b1 , w_14008 );
or ( \5658_b0 , \4579_b0 , \5657_b0 );
not ( \5657_b0 , w_14009 );
and ( w_14009 , w_14008 , \5657_b1 );
or ( \5659_b1 , \4465_b1 , \5658_b1 );
not ( \5658_b1 , w_14010 );
and ( \5659_b0 , \4465_b0 , w_14011 );
and ( w_14010 , w_14011 , \5658_b0 );
or ( \5660_b1 , \4464_b1 , w_14012 );
or ( \5660_b0 , \4464_b0 , \5659_b0 );
not ( \5659_b0 , w_14013 );
and ( w_14013 , w_14012 , \5659_b1 );
or ( \5661_b1 , \4369_b1 , \5660_b1 );
not ( \5660_b1 , w_14014 );
and ( \5661_b0 , \4369_b0 , w_14015 );
and ( w_14014 , w_14015 , \5660_b0 );
or ( \5662_b1 , \4368_b1 , w_14016 );
or ( \5662_b0 , \4368_b0 , \5661_b0 );
not ( \5661_b0 , w_14017 );
and ( w_14017 , w_14016 , \5661_b1 );
or ( \5663_b1 , \4361_b1 , \5662_b1 );
not ( \5662_b1 , w_14018 );
and ( \5663_b0 , \4361_b0 , w_14019 );
and ( w_14018 , w_14019 , \5662_b0 );
or ( \5664_b1 , \4360_b1 , w_14020 );
or ( \5664_b0 , \4360_b0 , \5663_b0 );
not ( \5663_b0 , w_14021 );
and ( w_14021 , w_14020 , \5663_b1 );
or ( \5665_b1 , \4246_b1 , \5664_b1 );
not ( \5664_b1 , w_14022 );
and ( \5665_b0 , \4246_b0 , w_14023 );
and ( w_14022 , w_14023 , \5664_b0 );
or ( \5666_b1 , \4245_b1 , w_14024 );
or ( \5666_b0 , \4245_b0 , \5665_b0 );
not ( \5665_b0 , w_14025 );
and ( w_14025 , w_14024 , \5665_b1 );
or ( \5667_b1 , \4122_b1 , \5666_b1 );
not ( \5666_b1 , w_14026 );
and ( \5667_b0 , \4122_b0 , w_14027 );
and ( w_14026 , w_14027 , \5666_b0 );
or ( \5668_b1 , \4121_b1 , w_14028 );
or ( \5668_b0 , \4121_b0 , \5667_b0 );
not ( \5667_b0 , w_14029 );
and ( w_14029 , w_14028 , \5667_b1 );
or ( \5669_b1 , \3982_b1 , \5668_b1 );
not ( \5668_b1 , w_14030 );
and ( \5669_b0 , \3982_b0 , w_14031 );
and ( w_14030 , w_14031 , \5668_b0 );
or ( \5670_b1 , \3981_b1 , w_14032 );
or ( \5670_b0 , \3981_b0 , \5669_b0 );
not ( \5669_b0 , w_14033 );
and ( w_14033 , w_14032 , \5669_b1 );
or ( \5671_b1 , \3858_b1 , \5670_b1 );
not ( \5670_b1 , w_14034 );
and ( \5671_b0 , \3858_b0 , w_14035 );
and ( w_14034 , w_14035 , \5670_b0 );
or ( \5672_b1 , \3857_b1 , w_14036 );
or ( \5672_b0 , \3857_b0 , \5671_b0 );
not ( \5671_b0 , w_14037 );
and ( w_14037 , w_14036 , \5671_b1 );
or ( \5673_b1 , \3714_b1 , \5672_b1 );
not ( \5672_b1 , w_14038 );
and ( \5673_b0 , \3714_b0 , w_14039 );
and ( w_14038 , w_14039 , \5672_b0 );
or ( \5674_b1 , \3713_b1 , w_14040 );
or ( \5674_b0 , \3713_b0 , \5673_b0 );
not ( \5673_b0 , w_14041 );
and ( w_14041 , w_14040 , \5673_b1 );
or ( \5675_b1 , \3589_b1 , \5674_b1 );
not ( \5674_b1 , w_14042 );
and ( \5675_b0 , \3589_b0 , w_14043 );
and ( w_14042 , w_14043 , \5674_b0 );
or ( \5676_b1 , \3588_b1 , w_14044 );
or ( \5676_b0 , \3588_b0 , \5675_b0 );
not ( \5675_b0 , w_14045 );
and ( w_14045 , w_14044 , \5675_b1 );
or ( \5677_b1 , \3450_b1 , \5676_b1 );
not ( \5676_b1 , w_14046 );
and ( \5677_b0 , \3450_b0 , w_14047 );
and ( w_14046 , w_14047 , \5676_b0 );
or ( \5678_b1 , \3449_b1 , w_14048 );
or ( \5678_b0 , \3449_b0 , \5677_b0 );
not ( \5677_b0 , w_14049 );
and ( w_14049 , w_14048 , \5677_b1 );
or ( \5679_b1 , \3285_b1 , \5678_b1 );
not ( \5678_b1 , w_14050 );
and ( \5679_b0 , \3285_b0 , w_14051 );
and ( w_14050 , w_14051 , \5678_b0 );
or ( \5680_b1 , \3284_b1 , w_14052 );
or ( \5680_b0 , \3284_b0 , \5679_b0 );
not ( \5679_b0 , w_14053 );
and ( w_14053 , w_14052 , \5679_b1 );
or ( \5681_b1 , \3137_b1 , \5680_b1 );
not ( \5680_b1 , w_14054 );
and ( \5681_b0 , \3137_b0 , w_14055 );
and ( w_14054 , w_14055 , \5680_b0 );
or ( \5682_b1 , \3136_b1 , w_14056 );
or ( \5682_b0 , \3136_b0 , \5681_b0 );
not ( \5681_b0 , w_14057 );
and ( w_14057 , w_14056 , \5681_b1 );
or ( \5683_b1 , \2990_b1 , \5682_b1 );
not ( \5682_b1 , w_14058 );
and ( \5683_b0 , \2990_b0 , w_14059 );
and ( w_14058 , w_14059 , \5682_b0 );
or ( \5684_b1 , \2989_b1 , w_14060 );
or ( \5684_b0 , \2989_b0 , \5683_b0 );
not ( \5683_b0 , w_14061 );
and ( w_14061 , w_14060 , \5683_b1 );
or ( \5685_b1 , \2822_b1 , \5684_b1 );
not ( \5684_b1 , w_14062 );
and ( \5685_b0 , \2822_b0 , w_14063 );
and ( w_14062 , w_14063 , \5684_b0 );
or ( \5686_b1 , \2821_b1 , w_14064 );
or ( \5686_b0 , \2821_b0 , \5685_b0 );
not ( \5685_b0 , w_14065 );
and ( w_14065 , w_14064 , \5685_b1 );
or ( \5687_b1 , \2674_b1 , \5686_b1 );
not ( \5686_b1 , w_14066 );
and ( \5687_b0 , \2674_b0 , w_14067 );
and ( w_14066 , w_14067 , \5686_b0 );
or ( \5688_b1 , \2673_b1 , w_14068 );
or ( \5688_b0 , \2673_b0 , \5687_b0 );
not ( \5687_b0 , w_14069 );
and ( w_14069 , w_14068 , \5687_b1 );
or ( \5689_b1 , \2504_b1 , \5688_b1 );
not ( \5688_b1 , w_14070 );
and ( \5689_b0 , \2504_b0 , w_14071 );
and ( w_14070 , w_14071 , \5688_b0 );
or ( \5690_b1 , \2503_b1 , w_14072 );
or ( \5690_b0 , \2503_b0 , \5689_b0 );
not ( \5689_b0 , w_14073 );
and ( w_14073 , w_14072 , \5689_b1 );
or ( \5691_b1 , \2366_b1 , \5690_b1 );
not ( \5690_b1 , w_14074 );
and ( \5691_b0 , \2366_b0 , w_14075 );
and ( w_14074 , w_14075 , \5690_b0 );
or ( \5692_b1 , \2365_b1 , w_14076 );
or ( \5692_b0 , \2365_b0 , \5691_b0 );
not ( \5691_b0 , w_14077 );
and ( w_14077 , w_14076 , \5691_b1 );
or ( \5693_b1 , \2222_b1 , \5692_b1 );
not ( \5692_b1 , w_14078 );
and ( \5693_b0 , \2222_b0 , w_14079 );
and ( w_14078 , w_14079 , \5692_b0 );
or ( \5694_b1 , \2221_b1 , w_14080 );
or ( \5694_b0 , \2221_b0 , \5693_b0 );
not ( \5693_b0 , w_14081 );
and ( w_14081 , w_14080 , \5693_b1 );
or ( \5695_b1 , \2083_b1 , \5694_b1 );
not ( \5694_b1 , w_14082 );
and ( \5695_b0 , \2083_b0 , w_14083 );
and ( w_14082 , w_14083 , \5694_b0 );
or ( \5696_b1 , \2082_b1 , w_14084 );
or ( \5696_b0 , \2082_b0 , \5695_b0 );
not ( \5695_b0 , w_14085 );
and ( w_14085 , w_14084 , \5695_b1 );
or ( \5697_b1 , \1950_b1 , \5696_b1 );
not ( \5696_b1 , w_14086 );
and ( \5697_b0 , \1950_b0 , w_14087 );
and ( w_14086 , w_14087 , \5696_b0 );
or ( \5698_b1 , \1949_b1 , w_14088 );
or ( \5698_b0 , \1949_b0 , \5697_b0 );
not ( \5697_b0 , w_14089 );
and ( w_14089 , w_14088 , \5697_b1 );
or ( \5699_b1 , \1827_b1 , \5698_b1 );
not ( \5698_b1 , w_14090 );
and ( \5699_b0 , \1827_b0 , w_14091 );
and ( w_14090 , w_14091 , \5698_b0 );
or ( \5700_b1 , \1826_b1 , w_14092 );
or ( \5700_b0 , \1826_b0 , \5699_b0 );
not ( \5699_b0 , w_14093 );
and ( w_14093 , w_14092 , \5699_b1 );
or ( \5701_b1 , \1704_b1 , \5700_b1 );
not ( \5700_b1 , w_14094 );
and ( \5701_b0 , \1704_b0 , w_14095 );
and ( w_14094 , w_14095 , \5700_b0 );
or ( \5702_b1 , \1703_b1 , w_14096 );
or ( \5702_b0 , \1703_b0 , \5701_b0 );
not ( \5701_b0 , w_14097 );
and ( w_14097 , w_14096 , \5701_b1 );
or ( \5703_b1 , \1586_b1 , \5702_b1 );
not ( \5702_b1 , w_14098 );
and ( \5703_b0 , \1586_b0 , w_14099 );
and ( w_14098 , w_14099 , \5702_b0 );
or ( \5704_b1 , \1585_b1 , w_14100 );
or ( \5704_b0 , \1585_b0 , \5703_b0 );
not ( \5703_b0 , w_14101 );
and ( w_14101 , w_14100 , \5703_b1 );
or ( \5705_b1 , \1471_b1 , \5704_b1 );
not ( \5704_b1 , w_14102 );
and ( \5705_b0 , \1471_b0 , w_14103 );
and ( w_14102 , w_14103 , \5704_b0 );
or ( \5706_b1 , \1470_b1 , w_14104 );
or ( \5706_b0 , \1470_b0 , \5705_b0 );
not ( \5705_b0 , w_14105 );
and ( w_14105 , w_14104 , \5705_b1 );
or ( \5707_b1 , \1355_b1 , \5706_b1 );
not ( \5706_b1 , w_14106 );
and ( \5707_b0 , \1355_b0 , w_14107 );
and ( w_14106 , w_14107 , \5706_b0 );
or ( \5708_b1 , \1354_b1 , w_14108 );
or ( \5708_b0 , \1354_b0 , \5707_b0 );
not ( \5707_b0 , w_14109 );
and ( w_14109 , w_14108 , \5707_b1 );
or ( \5709_b1 , \1241_b1 , \5708_b1 );
not ( \5708_b1 , w_14110 );
and ( \5709_b0 , \1241_b0 , w_14111 );
and ( w_14110 , w_14111 , \5708_b0 );
or ( \5710_b1 , \1240_b1 , w_14112 );
or ( \5710_b0 , \1240_b0 , \5709_b0 );
not ( \5709_b0 , w_14113 );
and ( w_14113 , w_14112 , \5709_b1 );
or ( \5711_b1 , \1057_b1 , \5710_b1 );
not ( \5710_b1 , w_14114 );
and ( \5711_b0 , \1057_b0 , w_14115 );
and ( w_14114 , w_14115 , \5710_b0 );
or ( \5712_b1 , \1056_b1 , w_14116 );
or ( \5712_b0 , \1056_b0 , \5711_b0 );
not ( \5711_b0 , w_14117 );
and ( w_14117 , w_14116 , \5711_b1 );
or ( \5713_b1 , \976_b1 , \5712_b1 );
not ( \5712_b1 , w_14118 );
and ( \5713_b0 , \976_b0 , w_14119 );
and ( w_14118 , w_14119 , \5712_b0 );
or ( \5714_b1 , \975_b1 , w_14120 );
or ( \5714_b0 , \975_b0 , \5713_b0 );
not ( \5713_b0 , w_14121 );
and ( w_14121 , w_14120 , \5713_b1 );
or ( \5715_b1 , \893_b1 , \5714_b1 );
not ( \5714_b1 , w_14122 );
and ( \5715_b0 , \893_b0 , w_14123 );
and ( w_14122 , w_14123 , \5714_b0 );
or ( \5716_b1 , \892_b1 , w_14124 );
or ( \5716_b0 , \892_b0 , \5715_b0 );
not ( \5715_b0 , w_14125 );
and ( w_14125 , w_14124 , \5715_b1 );
or ( \5717_b1 , \810_b1 , \5716_b1 );
not ( \5716_b1 , w_14126 );
and ( \5717_b0 , \810_b0 , w_14127 );
and ( w_14126 , w_14127 , \5716_b0 );
or ( \5718_b1 , \809_b1 , w_14128 );
or ( \5718_b0 , \809_b0 , \5717_b0 );
not ( \5717_b0 , w_14129 );
and ( w_14129 , w_14128 , \5717_b1 );
or ( \5719_b1 , \735_b1 , \5718_b1 );
not ( \5718_b1 , w_14130 );
and ( \5719_b0 , \735_b0 , w_14131 );
and ( w_14130 , w_14131 , \5718_b0 );
or ( \5720_b1 , \734_b1 , w_14132 );
or ( \5720_b0 , \734_b0 , \5719_b0 );
not ( \5719_b0 , w_14133 );
and ( w_14133 , w_14132 , \5719_b1 );
or ( \5721_b1 , \659_b1 , \5720_b1 );
not ( \5720_b1 , w_14134 );
and ( \5721_b0 , \659_b0 , w_14135 );
and ( w_14134 , w_14135 , \5720_b0 );
or ( \5722_b1 , \658_b1 , w_14136 );
or ( \5722_b0 , \658_b0 , \5721_b0 );
not ( \5721_b0 , w_14137 );
and ( w_14137 , w_14136 , \5721_b1 );
or ( \5723_b1 , \537_b1 , \5722_b1 );
not ( \5722_b1 , w_14138 );
and ( \5723_b0 , \537_b0 , w_14139 );
and ( w_14138 , w_14139 , \5722_b0 );
or ( \5724_b1 , \536_b1 , w_14140 );
or ( \5724_b0 , \536_b0 , \5723_b0 );
not ( \5723_b0 , w_14141 );
and ( w_14141 , w_14140 , \5723_b1 );
or ( \5725_b1 , \484_b1 , \5724_b1 );
xor ( \5725_b0 , \484_b0 , w_14142 );
not ( w_14142 , w_14143 );
and ( w_14143 , \5724_b1 , \5724_b0 );
buf ( \5726_b1 , \5725_b1 );
buf ( \5726_b0 , \5725_b0 );
buf ( \5727_b1 , \5726_b1 );
buf ( \5727_b0 , \5726_b0 );
or ( \5728_b1 , \537_b1 , \5722_b1 );
xor ( \5728_b0 , \537_b0 , w_14144 );
not ( w_14144 , w_14145 );
and ( w_14145 , \5722_b1 , \5722_b0 );
buf ( \5729_b1 , \5728_b1 );
buf ( \5729_b0 , \5728_b0 );
buf ( \5730_b1 , \5729_b1 );
buf ( \5730_b0 , \5729_b0 );
or ( \5731_b1 , \659_b1 , \5720_b1 );
xor ( \5731_b0 , \659_b0 , w_14146 );
not ( w_14146 , w_14147 );
and ( w_14147 , \5720_b1 , \5720_b0 );
buf ( \5732_b1 , \5731_b1 );
buf ( \5732_b0 , \5731_b0 );
buf ( \5733_b1 , \5732_b1 );
buf ( \5733_b0 , \5732_b0 );
or ( \5734_b1 , \5730_b1 , \5733_b1 );
not ( \5733_b1 , w_14148 );
and ( \5734_b0 , \5730_b0 , w_14149 );
and ( w_14148 , w_14149 , \5733_b0 );
buf ( \5735_b1 , \5734_b1 );
not ( \5735_b1 , w_14150 );
not ( \5735_b0 , w_14151 );
and ( w_14150 , w_14151 , \5734_b0 );
or ( \5736_b1 , \5727_b1 , \5735_b1 );
not ( \5735_b1 , w_14152 );
and ( \5736_b0 , \5727_b0 , w_14153 );
and ( w_14152 , w_14153 , \5735_b0 );
buf ( \5737_b1 , RIa167a08_1_b1 );
buf ( \5737_b0 , RIa167a08_1_b0 );
or ( \5738_b1 , \4369_b1 , \5660_b1 );
xor ( \5738_b0 , \4369_b0 , w_14154 );
not ( w_14154 , w_14155 );
and ( w_14155 , \5660_b1 , \5660_b0 );
buf ( \5739_b1 , \5738_b1 );
buf ( \5739_b0 , \5738_b0 );
buf ( \5740_b1 , \5739_b1 );
buf ( \5740_b0 , \5739_b0 );
or ( \5741_b1 , \4465_b1 , \5658_b1 );
xor ( \5741_b0 , \4465_b0 , w_14156 );
not ( w_14156 , w_14157 );
and ( w_14157 , \5658_b1 , \5658_b0 );
buf ( \5742_b1 , \5741_b1 );
buf ( \5742_b0 , \5741_b0 );
buf ( \5743_b1 , \5742_b1 );
buf ( \5743_b0 , \5742_b0 );
or ( \5744_b1 , \5740_b1 , \5743_b1 );
xor ( \5744_b0 , \5740_b0 , w_14158 );
not ( w_14158 , w_14159 );
and ( w_14159 , \5743_b1 , \5743_b0 );
or ( \5745_b1 , \4580_b1 , \5656_b1 );
xor ( \5745_b0 , \4580_b0 , w_14160 );
not ( w_14160 , w_14161 );
and ( w_14161 , \5656_b1 , \5656_b0 );
buf ( \5746_b1 , \5745_b1 );
buf ( \5746_b0 , \5745_b0 );
buf ( \5747_b1 , \5746_b1 );
buf ( \5747_b0 , \5746_b0 );
or ( \5748_b1 , \5743_b1 , \5747_b1 );
xor ( \5748_b0 , \5743_b0 , w_14162 );
not ( w_14162 , w_14163 );
and ( w_14163 , \5747_b1 , \5747_b0 );
buf ( \5749_b1 , \5748_b1 );
not ( \5749_b1 , w_14164 );
not ( \5749_b0 , w_14165 );
and ( w_14164 , w_14165 , \5748_b0 );
or ( \5750_b1 , \5744_b1 , \5749_b1 );
not ( \5749_b1 , w_14166 );
and ( \5750_b0 , \5744_b0 , w_14167 );
and ( w_14166 , w_14167 , \5749_b0 );
or ( \5751_b1 , \5737_b1 , \5750_b1 );
not ( \5750_b1 , w_14168 );
and ( \5751_b0 , \5737_b0 , w_14169 );
and ( w_14168 , w_14169 , \5750_b0 );
buf ( \5752_b1 , \5751_b1 );
not ( \5752_b1 , w_14170 );
not ( \5752_b0 , w_14171 );
and ( w_14170 , w_14171 , \5751_b0 );
or ( \5753_b1 , \5743_b1 , \5747_b1 );
not ( \5747_b1 , w_14172 );
and ( \5753_b0 , \5743_b0 , w_14173 );
and ( w_14172 , w_14173 , \5747_b0 );
buf ( \5754_b1 , \5753_b1 );
not ( \5754_b1 , w_14174 );
not ( \5754_b0 , w_14175 );
and ( w_14174 , w_14175 , \5753_b0 );
or ( \5755_b1 , \5740_b1 , \5754_b1 );
not ( \5754_b1 , w_14176 );
and ( \5755_b0 , \5740_b0 , w_14177 );
and ( w_14176 , w_14177 , \5754_b0 );
or ( \5756_b1 , \5752_b1 , w_14178 );
xor ( \5756_b0 , \5752_b0 , w_14180 );
not ( w_14180 , w_14181 );
and ( w_14181 , w_14178 , w_14179 );
buf ( w_14178 , \5755_b1 );
not ( w_14178 , w_14182 );
not ( w_14179 , w_14183 );
and ( w_14182 , w_14183 , \5755_b0 );
or ( \5757_b1 , \5736_b1 , \5756_b1 );
not ( \5756_b1 , w_14184 );
and ( \5757_b0 , \5736_b0 , w_14185 );
and ( w_14184 , w_14185 , \5756_b0 );
buf ( \5758_b1 , RIa167918_3_b1 );
buf ( \5758_b0 , RIa167918_3_b0 );
or ( \5759_b1 , \4246_b1 , \5664_b1 );
xor ( \5759_b0 , \4246_b0 , w_14186 );
not ( w_14186 , w_14187 );
and ( w_14187 , \5664_b1 , \5664_b0 );
buf ( \5760_b1 , \5759_b1 );
buf ( \5760_b0 , \5759_b0 );
buf ( \5761_b1 , \5760_b1 );
buf ( \5761_b0 , \5760_b0 );
or ( \5762_b1 , \4361_b1 , \5662_b1 );
xor ( \5762_b0 , \4361_b0 , w_14188 );
not ( w_14188 , w_14189 );
and ( w_14189 , \5662_b1 , \5662_b0 );
buf ( \5763_b1 , \5762_b1 );
buf ( \5763_b0 , \5762_b0 );
buf ( \5764_b1 , \5763_b1 );
buf ( \5764_b0 , \5763_b0 );
or ( \5765_b1 , \5761_b1 , \5764_b1 );
xor ( \5765_b0 , \5761_b0 , w_14190 );
not ( w_14190 , w_14191 );
and ( w_14191 , \5764_b1 , \5764_b0 );
or ( \5766_b1 , \5764_b1 , \5740_b1 );
xor ( \5766_b0 , \5764_b0 , w_14192 );
not ( w_14192 , w_14193 );
and ( w_14193 , \5740_b1 , \5740_b0 );
buf ( \5767_b1 , \5766_b1 );
not ( \5767_b1 , w_14194 );
not ( \5767_b0 , w_14195 );
and ( w_14194 , w_14195 , \5766_b0 );
or ( \5768_b1 , \5765_b1 , \5767_b1 );
not ( \5767_b1 , w_14196 );
and ( \5768_b0 , \5765_b0 , w_14197 );
and ( w_14196 , w_14197 , \5767_b0 );
or ( \5769_b1 , \5758_b1 , \5768_b1 );
not ( \5768_b1 , w_14198 );
and ( \5769_b0 , \5758_b0 , w_14199 );
and ( w_14198 , w_14199 , \5768_b0 );
buf ( \5770_b1 , RIa167990_2_b1 );
buf ( \5770_b0 , RIa167990_2_b0 );
or ( \5771_b1 , \5770_b1 , \5766_b1 );
not ( \5766_b1 , w_14200 );
and ( \5771_b0 , \5770_b0 , w_14201 );
and ( w_14200 , w_14201 , \5766_b0 );
or ( \5772_b1 , \5769_b1 , w_14203 );
not ( w_14203 , w_14204 );
and ( \5772_b0 , \5769_b0 , w_14205 );
and ( w_14204 ,  , w_14205 );
buf ( w_14203 , \5771_b1 );
not ( w_14203 , w_14206 );
not (  , w_14207 );
and ( w_14206 , w_14207 , \5771_b0 );
or ( \5773_b1 , \5764_b1 , \5740_b1 );
not ( \5740_b1 , w_14208 );
and ( \5773_b0 , \5764_b0 , w_14209 );
and ( w_14208 , w_14209 , \5740_b0 );
buf ( \5774_b1 , \5773_b1 );
not ( \5774_b1 , w_14210 );
not ( \5774_b0 , w_14211 );
and ( w_14210 , w_14211 , \5773_b0 );
or ( \5775_b1 , \5761_b1 , \5774_b1 );
not ( \5774_b1 , w_14212 );
and ( \5775_b0 , \5761_b0 , w_14213 );
and ( w_14212 , w_14213 , \5774_b0 );
or ( \5776_b1 , \5772_b1 , w_14214 );
xor ( \5776_b0 , \5772_b0 , w_14216 );
not ( w_14216 , w_14217 );
and ( w_14217 , w_14214 , w_14215 );
buf ( w_14214 , \5775_b1 );
not ( w_14214 , w_14218 );
not ( w_14215 , w_14219 );
and ( w_14218 , w_14219 , \5775_b0 );
or ( \5777_b1 , \5756_b1 , \5776_b1 );
not ( \5776_b1 , w_14220 );
and ( \5777_b0 , \5756_b0 , w_14221 );
and ( w_14220 , w_14221 , \5776_b0 );
or ( \5778_b1 , \5736_b1 , \5776_b1 );
not ( \5776_b1 , w_14222 );
and ( \5778_b0 , \5736_b0 , w_14223 );
and ( w_14222 , w_14223 , \5776_b0 );
buf ( \5780_b1 , RIa167828_5_b1 );
buf ( \5780_b0 , RIa167828_5_b0 );
or ( \5781_b1 , \3982_b1 , \5668_b1 );
xor ( \5781_b0 , \3982_b0 , w_14224 );
not ( w_14224 , w_14225 );
and ( w_14225 , \5668_b1 , \5668_b0 );
buf ( \5782_b1 , \5781_b1 );
buf ( \5782_b0 , \5781_b0 );
buf ( \5783_b1 , \5782_b1 );
buf ( \5783_b0 , \5782_b0 );
or ( \5784_b1 , \4122_b1 , \5666_b1 );
xor ( \5784_b0 , \4122_b0 , w_14226 );
not ( w_14226 , w_14227 );
and ( w_14227 , \5666_b1 , \5666_b0 );
buf ( \5785_b1 , \5784_b1 );
buf ( \5785_b0 , \5784_b0 );
buf ( \5786_b1 , \5785_b1 );
buf ( \5786_b0 , \5785_b0 );
or ( \5787_b1 , \5783_b1 , \5786_b1 );
xor ( \5787_b0 , \5783_b0 , w_14228 );
not ( w_14228 , w_14229 );
and ( w_14229 , \5786_b1 , \5786_b0 );
or ( \5788_b1 , \5786_b1 , \5761_b1 );
xor ( \5788_b0 , \5786_b0 , w_14230 );
not ( w_14230 , w_14231 );
and ( w_14231 , \5761_b1 , \5761_b0 );
buf ( \5789_b1 , \5788_b1 );
not ( \5789_b1 , w_14232 );
not ( \5789_b0 , w_14233 );
and ( w_14232 , w_14233 , \5788_b0 );
or ( \5790_b1 , \5787_b1 , \5789_b1 );
not ( \5789_b1 , w_14234 );
and ( \5790_b0 , \5787_b0 , w_14235 );
and ( w_14234 , w_14235 , \5789_b0 );
or ( \5791_b1 , \5780_b1 , \5790_b1 );
not ( \5790_b1 , w_14236 );
and ( \5791_b0 , \5780_b0 , w_14237 );
and ( w_14236 , w_14237 , \5790_b0 );
buf ( \5792_b1 , RIa1678a0_4_b1 );
buf ( \5792_b0 , RIa1678a0_4_b0 );
or ( \5793_b1 , \5792_b1 , \5788_b1 );
not ( \5788_b1 , w_14238 );
and ( \5793_b0 , \5792_b0 , w_14239 );
and ( w_14238 , w_14239 , \5788_b0 );
or ( \5794_b1 , \5791_b1 , w_14241 );
not ( w_14241 , w_14242 );
and ( \5794_b0 , \5791_b0 , w_14243 );
and ( w_14242 ,  , w_14243 );
buf ( w_14241 , \5793_b1 );
not ( w_14241 , w_14244 );
not (  , w_14245 );
and ( w_14244 , w_14245 , \5793_b0 );
or ( \5795_b1 , \5786_b1 , \5761_b1 );
not ( \5761_b1 , w_14246 );
and ( \5795_b0 , \5786_b0 , w_14247 );
and ( w_14246 , w_14247 , \5761_b0 );
buf ( \5796_b1 , \5795_b1 );
not ( \5796_b1 , w_14248 );
not ( \5796_b0 , w_14249 );
and ( w_14248 , w_14249 , \5795_b0 );
or ( \5797_b1 , \5783_b1 , \5796_b1 );
not ( \5796_b1 , w_14250 );
and ( \5797_b0 , \5783_b0 , w_14251 );
and ( w_14250 , w_14251 , \5796_b0 );
or ( \5798_b1 , \5794_b1 , w_14252 );
xor ( \5798_b0 , \5794_b0 , w_14254 );
not ( w_14254 , w_14255 );
and ( w_14255 , w_14252 , w_14253 );
buf ( w_14252 , \5797_b1 );
not ( w_14252 , w_14256 );
not ( w_14253 , w_14257 );
and ( w_14256 , w_14257 , \5797_b0 );
buf ( \5799_b1 , RIa167738_7_b1 );
buf ( \5799_b0 , RIa167738_7_b0 );
or ( \5800_b1 , \3714_b1 , \5672_b1 );
xor ( \5800_b0 , \3714_b0 , w_14258 );
not ( w_14258 , w_14259 );
and ( w_14259 , \5672_b1 , \5672_b0 );
buf ( \5801_b1 , \5800_b1 );
buf ( \5801_b0 , \5800_b0 );
buf ( \5802_b1 , \5801_b1 );
buf ( \5802_b0 , \5801_b0 );
or ( \5803_b1 , \3858_b1 , \5670_b1 );
xor ( \5803_b0 , \3858_b0 , w_14260 );
not ( w_14260 , w_14261 );
and ( w_14261 , \5670_b1 , \5670_b0 );
buf ( \5804_b1 , \5803_b1 );
buf ( \5804_b0 , \5803_b0 );
buf ( \5805_b1 , \5804_b1 );
buf ( \5805_b0 , \5804_b0 );
or ( \5806_b1 , \5802_b1 , \5805_b1 );
xor ( \5806_b0 , \5802_b0 , w_14262 );
not ( w_14262 , w_14263 );
and ( w_14263 , \5805_b1 , \5805_b0 );
or ( \5807_b1 , \5805_b1 , \5783_b1 );
xor ( \5807_b0 , \5805_b0 , w_14264 );
not ( w_14264 , w_14265 );
and ( w_14265 , \5783_b1 , \5783_b0 );
buf ( \5808_b1 , \5807_b1 );
not ( \5808_b1 , w_14266 );
not ( \5808_b0 , w_14267 );
and ( w_14266 , w_14267 , \5807_b0 );
or ( \5809_b1 , \5806_b1 , \5808_b1 );
not ( \5808_b1 , w_14268 );
and ( \5809_b0 , \5806_b0 , w_14269 );
and ( w_14268 , w_14269 , \5808_b0 );
or ( \5810_b1 , \5799_b1 , \5809_b1 );
not ( \5809_b1 , w_14270 );
and ( \5810_b0 , \5799_b0 , w_14271 );
and ( w_14270 , w_14271 , \5809_b0 );
buf ( \5811_b1 , RIa1677b0_6_b1 );
buf ( \5811_b0 , RIa1677b0_6_b0 );
or ( \5812_b1 , \5811_b1 , \5807_b1 );
not ( \5807_b1 , w_14272 );
and ( \5812_b0 , \5811_b0 , w_14273 );
and ( w_14272 , w_14273 , \5807_b0 );
or ( \5813_b1 , \5810_b1 , w_14275 );
not ( w_14275 , w_14276 );
and ( \5813_b0 , \5810_b0 , w_14277 );
and ( w_14276 ,  , w_14277 );
buf ( w_14275 , \5812_b1 );
not ( w_14275 , w_14278 );
not (  , w_14279 );
and ( w_14278 , w_14279 , \5812_b0 );
or ( \5814_b1 , \5805_b1 , \5783_b1 );
not ( \5783_b1 , w_14280 );
and ( \5814_b0 , \5805_b0 , w_14281 );
and ( w_14280 , w_14281 , \5783_b0 );
buf ( \5815_b1 , \5814_b1 );
not ( \5815_b1 , w_14282 );
not ( \5815_b0 , w_14283 );
and ( w_14282 , w_14283 , \5814_b0 );
or ( \5816_b1 , \5802_b1 , \5815_b1 );
not ( \5815_b1 , w_14284 );
and ( \5816_b0 , \5802_b0 , w_14285 );
and ( w_14284 , w_14285 , \5815_b0 );
or ( \5817_b1 , \5813_b1 , w_14286 );
xor ( \5817_b0 , \5813_b0 , w_14288 );
not ( w_14288 , w_14289 );
and ( w_14289 , w_14286 , w_14287 );
buf ( w_14286 , \5816_b1 );
not ( w_14286 , w_14290 );
not ( w_14287 , w_14291 );
and ( w_14290 , w_14291 , \5816_b0 );
or ( \5818_b1 , \5798_b1 , \5817_b1 );
not ( \5817_b1 , w_14292 );
and ( \5818_b0 , \5798_b0 , w_14293 );
and ( w_14292 , w_14293 , \5817_b0 );
buf ( \5819_b1 , RIa167648_9_b1 );
buf ( \5819_b0 , RIa167648_9_b0 );
or ( \5820_b1 , \3450_b1 , \5676_b1 );
xor ( \5820_b0 , \3450_b0 , w_14294 );
not ( w_14294 , w_14295 );
and ( w_14295 , \5676_b1 , \5676_b0 );
buf ( \5821_b1 , \5820_b1 );
buf ( \5821_b0 , \5820_b0 );
buf ( \5822_b1 , \5821_b1 );
buf ( \5822_b0 , \5821_b0 );
or ( \5823_b1 , \3589_b1 , \5674_b1 );
xor ( \5823_b0 , \3589_b0 , w_14296 );
not ( w_14296 , w_14297 );
and ( w_14297 , \5674_b1 , \5674_b0 );
buf ( \5824_b1 , \5823_b1 );
buf ( \5824_b0 , \5823_b0 );
buf ( \5825_b1 , \5824_b1 );
buf ( \5825_b0 , \5824_b0 );
or ( \5826_b1 , \5822_b1 , \5825_b1 );
xor ( \5826_b0 , \5822_b0 , w_14298 );
not ( w_14298 , w_14299 );
and ( w_14299 , \5825_b1 , \5825_b0 );
or ( \5827_b1 , \5825_b1 , \5802_b1 );
xor ( \5827_b0 , \5825_b0 , w_14300 );
not ( w_14300 , w_14301 );
and ( w_14301 , \5802_b1 , \5802_b0 );
buf ( \5828_b1 , \5827_b1 );
not ( \5828_b1 , w_14302 );
not ( \5828_b0 , w_14303 );
and ( w_14302 , w_14303 , \5827_b0 );
or ( \5829_b1 , \5826_b1 , \5828_b1 );
not ( \5828_b1 , w_14304 );
and ( \5829_b0 , \5826_b0 , w_14305 );
and ( w_14304 , w_14305 , \5828_b0 );
or ( \5830_b1 , \5819_b1 , \5829_b1 );
not ( \5829_b1 , w_14306 );
and ( \5830_b0 , \5819_b0 , w_14307 );
and ( w_14306 , w_14307 , \5829_b0 );
buf ( \5831_b1 , RIa1676c0_8_b1 );
buf ( \5831_b0 , RIa1676c0_8_b0 );
or ( \5832_b1 , \5831_b1 , \5827_b1 );
not ( \5827_b1 , w_14308 );
and ( \5832_b0 , \5831_b0 , w_14309 );
and ( w_14308 , w_14309 , \5827_b0 );
or ( \5833_b1 , \5830_b1 , w_14311 );
not ( w_14311 , w_14312 );
and ( \5833_b0 , \5830_b0 , w_14313 );
and ( w_14312 ,  , w_14313 );
buf ( w_14311 , \5832_b1 );
not ( w_14311 , w_14314 );
not (  , w_14315 );
and ( w_14314 , w_14315 , \5832_b0 );
or ( \5834_b1 , \5825_b1 , \5802_b1 );
not ( \5802_b1 , w_14316 );
and ( \5834_b0 , \5825_b0 , w_14317 );
and ( w_14316 , w_14317 , \5802_b0 );
buf ( \5835_b1 , \5834_b1 );
not ( \5835_b1 , w_14318 );
not ( \5835_b0 , w_14319 );
and ( w_14318 , w_14319 , \5834_b0 );
or ( \5836_b1 , \5822_b1 , \5835_b1 );
not ( \5835_b1 , w_14320 );
and ( \5836_b0 , \5822_b0 , w_14321 );
and ( w_14320 , w_14321 , \5835_b0 );
or ( \5837_b1 , \5833_b1 , w_14322 );
xor ( \5837_b0 , \5833_b0 , w_14324 );
not ( w_14324 , w_14325 );
and ( w_14325 , w_14322 , w_14323 );
buf ( w_14322 , \5836_b1 );
not ( w_14322 , w_14326 );
not ( w_14323 , w_14327 );
and ( w_14326 , w_14327 , \5836_b0 );
or ( \5838_b1 , \5817_b1 , \5837_b1 );
not ( \5837_b1 , w_14328 );
and ( \5838_b0 , \5817_b0 , w_14329 );
and ( w_14328 , w_14329 , \5837_b0 );
or ( \5839_b1 , \5798_b1 , \5837_b1 );
not ( \5837_b1 , w_14330 );
and ( \5839_b0 , \5798_b0 , w_14331 );
and ( w_14330 , w_14331 , \5837_b0 );
or ( \5841_b1 , \5779_b1 , \5840_b1 );
not ( \5840_b1 , w_14332 );
and ( \5841_b0 , \5779_b0 , w_14333 );
and ( w_14332 , w_14333 , \5840_b0 );
buf ( \5842_b1 , RIa167558_11_b1 );
buf ( \5842_b0 , RIa167558_11_b0 );
or ( \5843_b1 , \3137_b1 , \5680_b1 );
xor ( \5843_b0 , \3137_b0 , w_14334 );
not ( w_14334 , w_14335 );
and ( w_14335 , \5680_b1 , \5680_b0 );
buf ( \5844_b1 , \5843_b1 );
buf ( \5844_b0 , \5843_b0 );
buf ( \5845_b1 , \5844_b1 );
buf ( \5845_b0 , \5844_b0 );
or ( \5846_b1 , \3285_b1 , \5678_b1 );
xor ( \5846_b0 , \3285_b0 , w_14336 );
not ( w_14336 , w_14337 );
and ( w_14337 , \5678_b1 , \5678_b0 );
buf ( \5847_b1 , \5846_b1 );
buf ( \5847_b0 , \5846_b0 );
buf ( \5848_b1 , \5847_b1 );
buf ( \5848_b0 , \5847_b0 );
or ( \5849_b1 , \5845_b1 , \5848_b1 );
xor ( \5849_b0 , \5845_b0 , w_14338 );
not ( w_14338 , w_14339 );
and ( w_14339 , \5848_b1 , \5848_b0 );
or ( \5850_b1 , \5848_b1 , \5822_b1 );
xor ( \5850_b0 , \5848_b0 , w_14340 );
not ( w_14340 , w_14341 );
and ( w_14341 , \5822_b1 , \5822_b0 );
buf ( \5851_b1 , \5850_b1 );
not ( \5851_b1 , w_14342 );
not ( \5851_b0 , w_14343 );
and ( w_14342 , w_14343 , \5850_b0 );
or ( \5852_b1 , \5849_b1 , \5851_b1 );
not ( \5851_b1 , w_14344 );
and ( \5852_b0 , \5849_b0 , w_14345 );
and ( w_14344 , w_14345 , \5851_b0 );
or ( \5853_b1 , \5842_b1 , \5852_b1 );
not ( \5852_b1 , w_14346 );
and ( \5853_b0 , \5842_b0 , w_14347 );
and ( w_14346 , w_14347 , \5852_b0 );
buf ( \5854_b1 , RIa1675d0_10_b1 );
buf ( \5854_b0 , RIa1675d0_10_b0 );
or ( \5855_b1 , \5854_b1 , \5850_b1 );
not ( \5850_b1 , w_14348 );
and ( \5855_b0 , \5854_b0 , w_14349 );
and ( w_14348 , w_14349 , \5850_b0 );
or ( \5856_b1 , \5853_b1 , w_14351 );
not ( w_14351 , w_14352 );
and ( \5856_b0 , \5853_b0 , w_14353 );
and ( w_14352 ,  , w_14353 );
buf ( w_14351 , \5855_b1 );
not ( w_14351 , w_14354 );
not (  , w_14355 );
and ( w_14354 , w_14355 , \5855_b0 );
or ( \5857_b1 , \5848_b1 , \5822_b1 );
not ( \5822_b1 , w_14356 );
and ( \5857_b0 , \5848_b0 , w_14357 );
and ( w_14356 , w_14357 , \5822_b0 );
buf ( \5858_b1 , \5857_b1 );
not ( \5858_b1 , w_14358 );
not ( \5858_b0 , w_14359 );
and ( w_14358 , w_14359 , \5857_b0 );
or ( \5859_b1 , \5845_b1 , \5858_b1 );
not ( \5858_b1 , w_14360 );
and ( \5859_b0 , \5845_b0 , w_14361 );
and ( w_14360 , w_14361 , \5858_b0 );
or ( \5860_b1 , \5856_b1 , w_14362 );
xor ( \5860_b0 , \5856_b0 , w_14364 );
not ( w_14364 , w_14365 );
and ( w_14365 , w_14362 , w_14363 );
buf ( w_14362 , \5859_b1 );
not ( w_14362 , w_14366 );
not ( w_14363 , w_14367 );
and ( w_14366 , w_14367 , \5859_b0 );
buf ( \5861_b1 , RIa167468_13_b1 );
buf ( \5861_b0 , RIa167468_13_b0 );
or ( \5862_b1 , \2822_b1 , \5684_b1 );
xor ( \5862_b0 , \2822_b0 , w_14368 );
not ( w_14368 , w_14369 );
and ( w_14369 , \5684_b1 , \5684_b0 );
buf ( \5863_b1 , \5862_b1 );
buf ( \5863_b0 , \5862_b0 );
buf ( \5864_b1 , \5863_b1 );
buf ( \5864_b0 , \5863_b0 );
or ( \5865_b1 , \2990_b1 , \5682_b1 );
xor ( \5865_b0 , \2990_b0 , w_14370 );
not ( w_14370 , w_14371 );
and ( w_14371 , \5682_b1 , \5682_b0 );
buf ( \5866_b1 , \5865_b1 );
buf ( \5866_b0 , \5865_b0 );
buf ( \5867_b1 , \5866_b1 );
buf ( \5867_b0 , \5866_b0 );
or ( \5868_b1 , \5864_b1 , \5867_b1 );
xor ( \5868_b0 , \5864_b0 , w_14372 );
not ( w_14372 , w_14373 );
and ( w_14373 , \5867_b1 , \5867_b0 );
or ( \5869_b1 , \5867_b1 , \5845_b1 );
xor ( \5869_b0 , \5867_b0 , w_14374 );
not ( w_14374 , w_14375 );
and ( w_14375 , \5845_b1 , \5845_b0 );
buf ( \5870_b1 , \5869_b1 );
not ( \5870_b1 , w_14376 );
not ( \5870_b0 , w_14377 );
and ( w_14376 , w_14377 , \5869_b0 );
or ( \5871_b1 , \5868_b1 , \5870_b1 );
not ( \5870_b1 , w_14378 );
and ( \5871_b0 , \5868_b0 , w_14379 );
and ( w_14378 , w_14379 , \5870_b0 );
or ( \5872_b1 , \5861_b1 , \5871_b1 );
not ( \5871_b1 , w_14380 );
and ( \5872_b0 , \5861_b0 , w_14381 );
and ( w_14380 , w_14381 , \5871_b0 );
buf ( \5873_b1 , RIa1674e0_12_b1 );
buf ( \5873_b0 , RIa1674e0_12_b0 );
or ( \5874_b1 , \5873_b1 , \5869_b1 );
not ( \5869_b1 , w_14382 );
and ( \5874_b0 , \5873_b0 , w_14383 );
and ( w_14382 , w_14383 , \5869_b0 );
or ( \5875_b1 , \5872_b1 , w_14385 );
not ( w_14385 , w_14386 );
and ( \5875_b0 , \5872_b0 , w_14387 );
and ( w_14386 ,  , w_14387 );
buf ( w_14385 , \5874_b1 );
not ( w_14385 , w_14388 );
not (  , w_14389 );
and ( w_14388 , w_14389 , \5874_b0 );
or ( \5876_b1 , \5867_b1 , \5845_b1 );
not ( \5845_b1 , w_14390 );
and ( \5876_b0 , \5867_b0 , w_14391 );
and ( w_14390 , w_14391 , \5845_b0 );
buf ( \5877_b1 , \5876_b1 );
not ( \5877_b1 , w_14392 );
not ( \5877_b0 , w_14393 );
and ( w_14392 , w_14393 , \5876_b0 );
or ( \5878_b1 , \5864_b1 , \5877_b1 );
not ( \5877_b1 , w_14394 );
and ( \5878_b0 , \5864_b0 , w_14395 );
and ( w_14394 , w_14395 , \5877_b0 );
or ( \5879_b1 , \5875_b1 , w_14396 );
xor ( \5879_b0 , \5875_b0 , w_14398 );
not ( w_14398 , w_14399 );
and ( w_14399 , w_14396 , w_14397 );
buf ( w_14396 , \5878_b1 );
not ( w_14396 , w_14400 );
not ( w_14397 , w_14401 );
and ( w_14400 , w_14401 , \5878_b0 );
or ( \5880_b1 , \5860_b1 , \5879_b1 );
not ( \5879_b1 , w_14402 );
and ( \5880_b0 , \5860_b0 , w_14403 );
and ( w_14402 , w_14403 , \5879_b0 );
buf ( \5881_b1 , RIa167378_15_b1 );
buf ( \5881_b0 , RIa167378_15_b0 );
or ( \5882_b1 , \2504_b1 , \5688_b1 );
xor ( \5882_b0 , \2504_b0 , w_14404 );
not ( w_14404 , w_14405 );
and ( w_14405 , \5688_b1 , \5688_b0 );
buf ( \5883_b1 , \5882_b1 );
buf ( \5883_b0 , \5882_b0 );
buf ( \5884_b1 , \5883_b1 );
buf ( \5884_b0 , \5883_b0 );
or ( \5885_b1 , \2674_b1 , \5686_b1 );
xor ( \5885_b0 , \2674_b0 , w_14406 );
not ( w_14406 , w_14407 );
and ( w_14407 , \5686_b1 , \5686_b0 );
buf ( \5886_b1 , \5885_b1 );
buf ( \5886_b0 , \5885_b0 );
buf ( \5887_b1 , \5886_b1 );
buf ( \5887_b0 , \5886_b0 );
or ( \5888_b1 , \5884_b1 , \5887_b1 );
xor ( \5888_b0 , \5884_b0 , w_14408 );
not ( w_14408 , w_14409 );
and ( w_14409 , \5887_b1 , \5887_b0 );
or ( \5889_b1 , \5887_b1 , \5864_b1 );
xor ( \5889_b0 , \5887_b0 , w_14410 );
not ( w_14410 , w_14411 );
and ( w_14411 , \5864_b1 , \5864_b0 );
buf ( \5890_b1 , \5889_b1 );
not ( \5890_b1 , w_14412 );
not ( \5890_b0 , w_14413 );
and ( w_14412 , w_14413 , \5889_b0 );
or ( \5891_b1 , \5888_b1 , \5890_b1 );
not ( \5890_b1 , w_14414 );
and ( \5891_b0 , \5888_b0 , w_14415 );
and ( w_14414 , w_14415 , \5890_b0 );
or ( \5892_b1 , \5881_b1 , \5891_b1 );
not ( \5891_b1 , w_14416 );
and ( \5892_b0 , \5881_b0 , w_14417 );
and ( w_14416 , w_14417 , \5891_b0 );
buf ( \5893_b1 , RIa1673f0_14_b1 );
buf ( \5893_b0 , RIa1673f0_14_b0 );
or ( \5894_b1 , \5893_b1 , \5889_b1 );
not ( \5889_b1 , w_14418 );
and ( \5894_b0 , \5893_b0 , w_14419 );
and ( w_14418 , w_14419 , \5889_b0 );
or ( \5895_b1 , \5892_b1 , w_14421 );
not ( w_14421 , w_14422 );
and ( \5895_b0 , \5892_b0 , w_14423 );
and ( w_14422 ,  , w_14423 );
buf ( w_14421 , \5894_b1 );
not ( w_14421 , w_14424 );
not (  , w_14425 );
and ( w_14424 , w_14425 , \5894_b0 );
or ( \5896_b1 , \5887_b1 , \5864_b1 );
not ( \5864_b1 , w_14426 );
and ( \5896_b0 , \5887_b0 , w_14427 );
and ( w_14426 , w_14427 , \5864_b0 );
buf ( \5897_b1 , \5896_b1 );
not ( \5897_b1 , w_14428 );
not ( \5897_b0 , w_14429 );
and ( w_14428 , w_14429 , \5896_b0 );
or ( \5898_b1 , \5884_b1 , \5897_b1 );
not ( \5897_b1 , w_14430 );
and ( \5898_b0 , \5884_b0 , w_14431 );
and ( w_14430 , w_14431 , \5897_b0 );
or ( \5899_b1 , \5895_b1 , w_14432 );
xor ( \5899_b0 , \5895_b0 , w_14434 );
not ( w_14434 , w_14435 );
and ( w_14435 , w_14432 , w_14433 );
buf ( w_14432 , \5898_b1 );
not ( w_14432 , w_14436 );
not ( w_14433 , w_14437 );
and ( w_14436 , w_14437 , \5898_b0 );
or ( \5900_b1 , \5879_b1 , \5899_b1 );
not ( \5899_b1 , w_14438 );
and ( \5900_b0 , \5879_b0 , w_14439 );
and ( w_14438 , w_14439 , \5899_b0 );
or ( \5901_b1 , \5860_b1 , \5899_b1 );
not ( \5899_b1 , w_14440 );
and ( \5901_b0 , \5860_b0 , w_14441 );
and ( w_14440 , w_14441 , \5899_b0 );
or ( \5903_b1 , \5840_b1 , \5902_b1 );
not ( \5902_b1 , w_14442 );
and ( \5903_b0 , \5840_b0 , w_14443 );
and ( w_14442 , w_14443 , \5902_b0 );
or ( \5904_b1 , \5779_b1 , \5902_b1 );
not ( \5902_b1 , w_14444 );
and ( \5904_b0 , \5779_b0 , w_14445 );
and ( w_14444 , w_14445 , \5902_b0 );
buf ( \5906_b1 , RIa167288_17_b1 );
buf ( \5906_b0 , RIa167288_17_b0 );
or ( \5907_b1 , \2222_b1 , \5692_b1 );
xor ( \5907_b0 , \2222_b0 , w_14446 );
not ( w_14446 , w_14447 );
and ( w_14447 , \5692_b1 , \5692_b0 );
buf ( \5908_b1 , \5907_b1 );
buf ( \5908_b0 , \5907_b0 );
buf ( \5909_b1 , \5908_b1 );
buf ( \5909_b0 , \5908_b0 );
or ( \5910_b1 , \2366_b1 , \5690_b1 );
xor ( \5910_b0 , \2366_b0 , w_14448 );
not ( w_14448 , w_14449 );
and ( w_14449 , \5690_b1 , \5690_b0 );
buf ( \5911_b1 , \5910_b1 );
buf ( \5911_b0 , \5910_b0 );
buf ( \5912_b1 , \5911_b1 );
buf ( \5912_b0 , \5911_b0 );
or ( \5913_b1 , \5909_b1 , \5912_b1 );
xor ( \5913_b0 , \5909_b0 , w_14450 );
not ( w_14450 , w_14451 );
and ( w_14451 , \5912_b1 , \5912_b0 );
or ( \5914_b1 , \5912_b1 , \5884_b1 );
xor ( \5914_b0 , \5912_b0 , w_14452 );
not ( w_14452 , w_14453 );
and ( w_14453 , \5884_b1 , \5884_b0 );
buf ( \5915_b1 , \5914_b1 );
not ( \5915_b1 , w_14454 );
not ( \5915_b0 , w_14455 );
and ( w_14454 , w_14455 , \5914_b0 );
or ( \5916_b1 , \5913_b1 , \5915_b1 );
not ( \5915_b1 , w_14456 );
and ( \5916_b0 , \5913_b0 , w_14457 );
and ( w_14456 , w_14457 , \5915_b0 );
or ( \5917_b1 , \5906_b1 , \5916_b1 );
not ( \5916_b1 , w_14458 );
and ( \5917_b0 , \5906_b0 , w_14459 );
and ( w_14458 , w_14459 , \5916_b0 );
buf ( \5918_b1 , RIa167300_16_b1 );
buf ( \5918_b0 , RIa167300_16_b0 );
or ( \5919_b1 , \5918_b1 , \5914_b1 );
not ( \5914_b1 , w_14460 );
and ( \5919_b0 , \5918_b0 , w_14461 );
and ( w_14460 , w_14461 , \5914_b0 );
or ( \5920_b1 , \5917_b1 , w_14463 );
not ( w_14463 , w_14464 );
and ( \5920_b0 , \5917_b0 , w_14465 );
and ( w_14464 ,  , w_14465 );
buf ( w_14463 , \5919_b1 );
not ( w_14463 , w_14466 );
not (  , w_14467 );
and ( w_14466 , w_14467 , \5919_b0 );
or ( \5921_b1 , \5912_b1 , \5884_b1 );
not ( \5884_b1 , w_14468 );
and ( \5921_b0 , \5912_b0 , w_14469 );
and ( w_14468 , w_14469 , \5884_b0 );
buf ( \5922_b1 , \5921_b1 );
not ( \5922_b1 , w_14470 );
not ( \5922_b0 , w_14471 );
and ( w_14470 , w_14471 , \5921_b0 );
or ( \5923_b1 , \5909_b1 , \5922_b1 );
not ( \5922_b1 , w_14472 );
and ( \5923_b0 , \5909_b0 , w_14473 );
and ( w_14472 , w_14473 , \5922_b0 );
or ( \5924_b1 , \5920_b1 , w_14474 );
xor ( \5924_b0 , \5920_b0 , w_14476 );
not ( w_14476 , w_14477 );
and ( w_14477 , w_14474 , w_14475 );
buf ( w_14474 , \5923_b1 );
not ( w_14474 , w_14478 );
not ( w_14475 , w_14479 );
and ( w_14478 , w_14479 , \5923_b0 );
buf ( \5925_b1 , RIa167198_19_b1 );
buf ( \5925_b0 , RIa167198_19_b0 );
or ( \5926_b1 , \1950_b1 , \5696_b1 );
xor ( \5926_b0 , \1950_b0 , w_14480 );
not ( w_14480 , w_14481 );
and ( w_14481 , \5696_b1 , \5696_b0 );
buf ( \5927_b1 , \5926_b1 );
buf ( \5927_b0 , \5926_b0 );
buf ( \5928_b1 , \5927_b1 );
buf ( \5928_b0 , \5927_b0 );
or ( \5929_b1 , \2083_b1 , \5694_b1 );
xor ( \5929_b0 , \2083_b0 , w_14482 );
not ( w_14482 , w_14483 );
and ( w_14483 , \5694_b1 , \5694_b0 );
buf ( \5930_b1 , \5929_b1 );
buf ( \5930_b0 , \5929_b0 );
buf ( \5931_b1 , \5930_b1 );
buf ( \5931_b0 , \5930_b0 );
or ( \5932_b1 , \5928_b1 , \5931_b1 );
xor ( \5932_b0 , \5928_b0 , w_14484 );
not ( w_14484 , w_14485 );
and ( w_14485 , \5931_b1 , \5931_b0 );
or ( \5933_b1 , \5931_b1 , \5909_b1 );
xor ( \5933_b0 , \5931_b0 , w_14486 );
not ( w_14486 , w_14487 );
and ( w_14487 , \5909_b1 , \5909_b0 );
buf ( \5934_b1 , \5933_b1 );
not ( \5934_b1 , w_14488 );
not ( \5934_b0 , w_14489 );
and ( w_14488 , w_14489 , \5933_b0 );
or ( \5935_b1 , \5932_b1 , \5934_b1 );
not ( \5934_b1 , w_14490 );
and ( \5935_b0 , \5932_b0 , w_14491 );
and ( w_14490 , w_14491 , \5934_b0 );
or ( \5936_b1 , \5925_b1 , \5935_b1 );
not ( \5935_b1 , w_14492 );
and ( \5936_b0 , \5925_b0 , w_14493 );
and ( w_14492 , w_14493 , \5935_b0 );
buf ( \5937_b1 , RIa167210_18_b1 );
buf ( \5937_b0 , RIa167210_18_b0 );
or ( \5938_b1 , \5937_b1 , \5933_b1 );
not ( \5933_b1 , w_14494 );
and ( \5938_b0 , \5937_b0 , w_14495 );
and ( w_14494 , w_14495 , \5933_b0 );
or ( \5939_b1 , \5936_b1 , w_14497 );
not ( w_14497 , w_14498 );
and ( \5939_b0 , \5936_b0 , w_14499 );
and ( w_14498 ,  , w_14499 );
buf ( w_14497 , \5938_b1 );
not ( w_14497 , w_14500 );
not (  , w_14501 );
and ( w_14500 , w_14501 , \5938_b0 );
or ( \5940_b1 , \5931_b1 , \5909_b1 );
not ( \5909_b1 , w_14502 );
and ( \5940_b0 , \5931_b0 , w_14503 );
and ( w_14502 , w_14503 , \5909_b0 );
buf ( \5941_b1 , \5940_b1 );
not ( \5941_b1 , w_14504 );
not ( \5941_b0 , w_14505 );
and ( w_14504 , w_14505 , \5940_b0 );
or ( \5942_b1 , \5928_b1 , \5941_b1 );
not ( \5941_b1 , w_14506 );
and ( \5942_b0 , \5928_b0 , w_14507 );
and ( w_14506 , w_14507 , \5941_b0 );
or ( \5943_b1 , \5939_b1 , w_14508 );
xor ( \5943_b0 , \5939_b0 , w_14510 );
not ( w_14510 , w_14511 );
and ( w_14511 , w_14508 , w_14509 );
buf ( w_14508 , \5942_b1 );
not ( w_14508 , w_14512 );
not ( w_14509 , w_14513 );
and ( w_14512 , w_14513 , \5942_b0 );
or ( \5944_b1 , \5924_b1 , \5943_b1 );
not ( \5943_b1 , w_14514 );
and ( \5944_b0 , \5924_b0 , w_14515 );
and ( w_14514 , w_14515 , \5943_b0 );
buf ( \5945_b1 , RIa1670a8_21_b1 );
buf ( \5945_b0 , RIa1670a8_21_b0 );
or ( \5946_b1 , \1704_b1 , \5700_b1 );
xor ( \5946_b0 , \1704_b0 , w_14516 );
not ( w_14516 , w_14517 );
and ( w_14517 , \5700_b1 , \5700_b0 );
buf ( \5947_b1 , \5946_b1 );
buf ( \5947_b0 , \5946_b0 );
buf ( \5948_b1 , \5947_b1 );
buf ( \5948_b0 , \5947_b0 );
or ( \5949_b1 , \1827_b1 , \5698_b1 );
xor ( \5949_b0 , \1827_b0 , w_14518 );
not ( w_14518 , w_14519 );
and ( w_14519 , \5698_b1 , \5698_b0 );
buf ( \5950_b1 , \5949_b1 );
buf ( \5950_b0 , \5949_b0 );
buf ( \5951_b1 , \5950_b1 );
buf ( \5951_b0 , \5950_b0 );
or ( \5952_b1 , \5948_b1 , \5951_b1 );
xor ( \5952_b0 , \5948_b0 , w_14520 );
not ( w_14520 , w_14521 );
and ( w_14521 , \5951_b1 , \5951_b0 );
or ( \5953_b1 , \5951_b1 , \5928_b1 );
xor ( \5953_b0 , \5951_b0 , w_14522 );
not ( w_14522 , w_14523 );
and ( w_14523 , \5928_b1 , \5928_b0 );
buf ( \5954_b1 , \5953_b1 );
not ( \5954_b1 , w_14524 );
not ( \5954_b0 , w_14525 );
and ( w_14524 , w_14525 , \5953_b0 );
or ( \5955_b1 , \5952_b1 , \5954_b1 );
not ( \5954_b1 , w_14526 );
and ( \5955_b0 , \5952_b0 , w_14527 );
and ( w_14526 , w_14527 , \5954_b0 );
or ( \5956_b1 , \5945_b1 , \5955_b1 );
not ( \5955_b1 , w_14528 );
and ( \5956_b0 , \5945_b0 , w_14529 );
and ( w_14528 , w_14529 , \5955_b0 );
buf ( \5957_b1 , RIa167120_20_b1 );
buf ( \5957_b0 , RIa167120_20_b0 );
or ( \5958_b1 , \5957_b1 , \5953_b1 );
not ( \5953_b1 , w_14530 );
and ( \5958_b0 , \5957_b0 , w_14531 );
and ( w_14530 , w_14531 , \5953_b0 );
or ( \5959_b1 , \5956_b1 , w_14533 );
not ( w_14533 , w_14534 );
and ( \5959_b0 , \5956_b0 , w_14535 );
and ( w_14534 ,  , w_14535 );
buf ( w_14533 , \5958_b1 );
not ( w_14533 , w_14536 );
not (  , w_14537 );
and ( w_14536 , w_14537 , \5958_b0 );
or ( \5960_b1 , \5951_b1 , \5928_b1 );
not ( \5928_b1 , w_14538 );
and ( \5960_b0 , \5951_b0 , w_14539 );
and ( w_14538 , w_14539 , \5928_b0 );
buf ( \5961_b1 , \5960_b1 );
not ( \5961_b1 , w_14540 );
not ( \5961_b0 , w_14541 );
and ( w_14540 , w_14541 , \5960_b0 );
or ( \5962_b1 , \5948_b1 , \5961_b1 );
not ( \5961_b1 , w_14542 );
and ( \5962_b0 , \5948_b0 , w_14543 );
and ( w_14542 , w_14543 , \5961_b0 );
or ( \5963_b1 , \5959_b1 , w_14544 );
xor ( \5963_b0 , \5959_b0 , w_14546 );
not ( w_14546 , w_14547 );
and ( w_14547 , w_14544 , w_14545 );
buf ( w_14544 , \5962_b1 );
not ( w_14544 , w_14548 );
not ( w_14545 , w_14549 );
and ( w_14548 , w_14549 , \5962_b0 );
or ( \5964_b1 , \5943_b1 , \5963_b1 );
not ( \5963_b1 , w_14550 );
and ( \5964_b0 , \5943_b0 , w_14551 );
and ( w_14550 , w_14551 , \5963_b0 );
or ( \5965_b1 , \5924_b1 , \5963_b1 );
not ( \5963_b1 , w_14552 );
and ( \5965_b0 , \5924_b0 , w_14553 );
and ( w_14552 , w_14553 , \5963_b0 );
buf ( \5967_b1 , RIa166fb8_23_b1 );
buf ( \5967_b0 , RIa166fb8_23_b0 );
or ( \5968_b1 , \1471_b1 , \5704_b1 );
xor ( \5968_b0 , \1471_b0 , w_14554 );
not ( w_14554 , w_14555 );
and ( w_14555 , \5704_b1 , \5704_b0 );
buf ( \5969_b1 , \5968_b1 );
buf ( \5969_b0 , \5968_b0 );
buf ( \5970_b1 , \5969_b1 );
buf ( \5970_b0 , \5969_b0 );
or ( \5971_b1 , \1586_b1 , \5702_b1 );
xor ( \5971_b0 , \1586_b0 , w_14556 );
not ( w_14556 , w_14557 );
and ( w_14557 , \5702_b1 , \5702_b0 );
buf ( \5972_b1 , \5971_b1 );
buf ( \5972_b0 , \5971_b0 );
buf ( \5973_b1 , \5972_b1 );
buf ( \5973_b0 , \5972_b0 );
or ( \5974_b1 , \5970_b1 , \5973_b1 );
xor ( \5974_b0 , \5970_b0 , w_14558 );
not ( w_14558 , w_14559 );
and ( w_14559 , \5973_b1 , \5973_b0 );
or ( \5975_b1 , \5973_b1 , \5948_b1 );
xor ( \5975_b0 , \5973_b0 , w_14560 );
not ( w_14560 , w_14561 );
and ( w_14561 , \5948_b1 , \5948_b0 );
buf ( \5976_b1 , \5975_b1 );
not ( \5976_b1 , w_14562 );
not ( \5976_b0 , w_14563 );
and ( w_14562 , w_14563 , \5975_b0 );
or ( \5977_b1 , \5974_b1 , \5976_b1 );
not ( \5976_b1 , w_14564 );
and ( \5977_b0 , \5974_b0 , w_14565 );
and ( w_14564 , w_14565 , \5976_b0 );
or ( \5978_b1 , \5967_b1 , \5977_b1 );
not ( \5977_b1 , w_14566 );
and ( \5978_b0 , \5967_b0 , w_14567 );
and ( w_14566 , w_14567 , \5977_b0 );
buf ( \5979_b1 , RIa167030_22_b1 );
buf ( \5979_b0 , RIa167030_22_b0 );
or ( \5980_b1 , \5979_b1 , \5975_b1 );
not ( \5975_b1 , w_14568 );
and ( \5980_b0 , \5979_b0 , w_14569 );
and ( w_14568 , w_14569 , \5975_b0 );
or ( \5981_b1 , \5978_b1 , w_14571 );
not ( w_14571 , w_14572 );
and ( \5981_b0 , \5978_b0 , w_14573 );
and ( w_14572 ,  , w_14573 );
buf ( w_14571 , \5980_b1 );
not ( w_14571 , w_14574 );
not (  , w_14575 );
and ( w_14574 , w_14575 , \5980_b0 );
or ( \5982_b1 , \5973_b1 , \5948_b1 );
not ( \5948_b1 , w_14576 );
and ( \5982_b0 , \5973_b0 , w_14577 );
and ( w_14576 , w_14577 , \5948_b0 );
buf ( \5983_b1 , \5982_b1 );
not ( \5983_b1 , w_14578 );
not ( \5983_b0 , w_14579 );
and ( w_14578 , w_14579 , \5982_b0 );
or ( \5984_b1 , \5970_b1 , \5983_b1 );
not ( \5983_b1 , w_14580 );
and ( \5984_b0 , \5970_b0 , w_14581 );
and ( w_14580 , w_14581 , \5983_b0 );
or ( \5985_b1 , \5981_b1 , w_14582 );
xor ( \5985_b0 , \5981_b0 , w_14584 );
not ( w_14584 , w_14585 );
and ( w_14585 , w_14582 , w_14583 );
buf ( w_14582 , \5984_b1 );
not ( w_14582 , w_14586 );
not ( w_14583 , w_14587 );
and ( w_14586 , w_14587 , \5984_b0 );
buf ( \5986_b1 , RIa166ec8_25_b1 );
buf ( \5986_b0 , RIa166ec8_25_b0 );
or ( \5987_b1 , \1241_b1 , \5708_b1 );
xor ( \5987_b0 , \1241_b0 , w_14588 );
not ( w_14588 , w_14589 );
and ( w_14589 , \5708_b1 , \5708_b0 );
buf ( \5988_b1 , \5987_b1 );
buf ( \5988_b0 , \5987_b0 );
buf ( \5989_b1 , \5988_b1 );
buf ( \5989_b0 , \5988_b0 );
or ( \5990_b1 , \1355_b1 , \5706_b1 );
xor ( \5990_b0 , \1355_b0 , w_14590 );
not ( w_14590 , w_14591 );
and ( w_14591 , \5706_b1 , \5706_b0 );
buf ( \5991_b1 , \5990_b1 );
buf ( \5991_b0 , \5990_b0 );
buf ( \5992_b1 , \5991_b1 );
buf ( \5992_b0 , \5991_b0 );
or ( \5993_b1 , \5989_b1 , \5992_b1 );
xor ( \5993_b0 , \5989_b0 , w_14592 );
not ( w_14592 , w_14593 );
and ( w_14593 , \5992_b1 , \5992_b0 );
or ( \5994_b1 , \5992_b1 , \5970_b1 );
xor ( \5994_b0 , \5992_b0 , w_14594 );
not ( w_14594 , w_14595 );
and ( w_14595 , \5970_b1 , \5970_b0 );
buf ( \5995_b1 , \5994_b1 );
not ( \5995_b1 , w_14596 );
not ( \5995_b0 , w_14597 );
and ( w_14596 , w_14597 , \5994_b0 );
or ( \5996_b1 , \5993_b1 , \5995_b1 );
not ( \5995_b1 , w_14598 );
and ( \5996_b0 , \5993_b0 , w_14599 );
and ( w_14598 , w_14599 , \5995_b0 );
or ( \5997_b1 , \5986_b1 , \5996_b1 );
not ( \5996_b1 , w_14600 );
and ( \5997_b0 , \5986_b0 , w_14601 );
and ( w_14600 , w_14601 , \5996_b0 );
buf ( \5998_b1 , RIa166f40_24_b1 );
buf ( \5998_b0 , RIa166f40_24_b0 );
or ( \5999_b1 , \5998_b1 , \5994_b1 );
not ( \5994_b1 , w_14602 );
and ( \5999_b0 , \5998_b0 , w_14603 );
and ( w_14602 , w_14603 , \5994_b0 );
or ( \6000_b1 , \5997_b1 , w_14605 );
not ( w_14605 , w_14606 );
and ( \6000_b0 , \5997_b0 , w_14607 );
and ( w_14606 ,  , w_14607 );
buf ( w_14605 , \5999_b1 );
not ( w_14605 , w_14608 );
not (  , w_14609 );
and ( w_14608 , w_14609 , \5999_b0 );
or ( \6001_b1 , \5992_b1 , \5970_b1 );
not ( \5970_b1 , w_14610 );
and ( \6001_b0 , \5992_b0 , w_14611 );
and ( w_14610 , w_14611 , \5970_b0 );
buf ( \6002_b1 , \6001_b1 );
not ( \6002_b1 , w_14612 );
not ( \6002_b0 , w_14613 );
and ( w_14612 , w_14613 , \6001_b0 );
or ( \6003_b1 , \5989_b1 , \6002_b1 );
not ( \6002_b1 , w_14614 );
and ( \6003_b0 , \5989_b0 , w_14615 );
and ( w_14614 , w_14615 , \6002_b0 );
or ( \6004_b1 , \6000_b1 , w_14616 );
xor ( \6004_b0 , \6000_b0 , w_14618 );
not ( w_14618 , w_14619 );
and ( w_14619 , w_14616 , w_14617 );
buf ( w_14616 , \6003_b1 );
not ( w_14616 , w_14620 );
not ( w_14617 , w_14621 );
and ( w_14620 , w_14621 , \6003_b0 );
or ( \6005_b1 , \5985_b1 , \6004_b1 );
not ( \6004_b1 , w_14622 );
and ( \6005_b0 , \5985_b0 , w_14623 );
and ( w_14622 , w_14623 , \6004_b0 );
buf ( \6006_b1 , RIa166dd8_27_b1 );
buf ( \6006_b0 , RIa166dd8_27_b0 );
or ( \6007_b1 , \976_b1 , \5712_b1 );
xor ( \6007_b0 , \976_b0 , w_14624 );
not ( w_14624 , w_14625 );
and ( w_14625 , \5712_b1 , \5712_b0 );
buf ( \6008_b1 , \6007_b1 );
buf ( \6008_b0 , \6007_b0 );
buf ( \6009_b1 , \6008_b1 );
buf ( \6009_b0 , \6008_b0 );
or ( \6010_b1 , \1057_b1 , \5710_b1 );
xor ( \6010_b0 , \1057_b0 , w_14626 );
not ( w_14626 , w_14627 );
and ( w_14627 , \5710_b1 , \5710_b0 );
buf ( \6011_b1 , \6010_b1 );
buf ( \6011_b0 , \6010_b0 );
buf ( \6012_b1 , \6011_b1 );
buf ( \6012_b0 , \6011_b0 );
or ( \6013_b1 , \6009_b1 , \6012_b1 );
xor ( \6013_b0 , \6009_b0 , w_14628 );
not ( w_14628 , w_14629 );
and ( w_14629 , \6012_b1 , \6012_b0 );
or ( \6014_b1 , \6012_b1 , \5989_b1 );
xor ( \6014_b0 , \6012_b0 , w_14630 );
not ( w_14630 , w_14631 );
and ( w_14631 , \5989_b1 , \5989_b0 );
buf ( \6015_b1 , \6014_b1 );
not ( \6015_b1 , w_14632 );
not ( \6015_b0 , w_14633 );
and ( w_14632 , w_14633 , \6014_b0 );
or ( \6016_b1 , \6013_b1 , \6015_b1 );
not ( \6015_b1 , w_14634 );
and ( \6016_b0 , \6013_b0 , w_14635 );
and ( w_14634 , w_14635 , \6015_b0 );
or ( \6017_b1 , \6006_b1 , \6016_b1 );
not ( \6016_b1 , w_14636 );
and ( \6017_b0 , \6006_b0 , w_14637 );
and ( w_14636 , w_14637 , \6016_b0 );
buf ( \6018_b1 , RIa166e50_26_b1 );
buf ( \6018_b0 , RIa166e50_26_b0 );
or ( \6019_b1 , \6018_b1 , \6014_b1 );
not ( \6014_b1 , w_14638 );
and ( \6019_b0 , \6018_b0 , w_14639 );
and ( w_14638 , w_14639 , \6014_b0 );
or ( \6020_b1 , \6017_b1 , w_14641 );
not ( w_14641 , w_14642 );
and ( \6020_b0 , \6017_b0 , w_14643 );
and ( w_14642 ,  , w_14643 );
buf ( w_14641 , \6019_b1 );
not ( w_14641 , w_14644 );
not (  , w_14645 );
and ( w_14644 , w_14645 , \6019_b0 );
or ( \6021_b1 , \6012_b1 , \5989_b1 );
not ( \5989_b1 , w_14646 );
and ( \6021_b0 , \6012_b0 , w_14647 );
and ( w_14646 , w_14647 , \5989_b0 );
buf ( \6022_b1 , \6021_b1 );
not ( \6022_b1 , w_14648 );
not ( \6022_b0 , w_14649 );
and ( w_14648 , w_14649 , \6021_b0 );
or ( \6023_b1 , \6009_b1 , \6022_b1 );
not ( \6022_b1 , w_14650 );
and ( \6023_b0 , \6009_b0 , w_14651 );
and ( w_14650 , w_14651 , \6022_b0 );
or ( \6024_b1 , \6020_b1 , w_14652 );
xor ( \6024_b0 , \6020_b0 , w_14654 );
not ( w_14654 , w_14655 );
and ( w_14655 , w_14652 , w_14653 );
buf ( w_14652 , \6023_b1 );
not ( w_14652 , w_14656 );
not ( w_14653 , w_14657 );
and ( w_14656 , w_14657 , \6023_b0 );
or ( \6025_b1 , \6004_b1 , \6024_b1 );
not ( \6024_b1 , w_14658 );
and ( \6025_b0 , \6004_b0 , w_14659 );
and ( w_14658 , w_14659 , \6024_b0 );
or ( \6026_b1 , \5985_b1 , \6024_b1 );
not ( \6024_b1 , w_14660 );
and ( \6026_b0 , \5985_b0 , w_14661 );
and ( w_14660 , w_14661 , \6024_b0 );
or ( \6028_b1 , \5966_b1 , \6027_b1 );
not ( \6027_b1 , w_14662 );
and ( \6028_b0 , \5966_b0 , w_14663 );
and ( w_14662 , w_14663 , \6027_b0 );
buf ( \6029_b1 , RIa166ce8_29_b1 );
buf ( \6029_b0 , RIa166ce8_29_b0 );
or ( \6030_b1 , \810_b1 , \5716_b1 );
xor ( \6030_b0 , \810_b0 , w_14664 );
not ( w_14664 , w_14665 );
and ( w_14665 , \5716_b1 , \5716_b0 );
buf ( \6031_b1 , \6030_b1 );
buf ( \6031_b0 , \6030_b0 );
buf ( \6032_b1 , \6031_b1 );
buf ( \6032_b0 , \6031_b0 );
or ( \6033_b1 , \893_b1 , \5714_b1 );
xor ( \6033_b0 , \893_b0 , w_14666 );
not ( w_14666 , w_14667 );
and ( w_14667 , \5714_b1 , \5714_b0 );
buf ( \6034_b1 , \6033_b1 );
buf ( \6034_b0 , \6033_b0 );
buf ( \6035_b1 , \6034_b1 );
buf ( \6035_b0 , \6034_b0 );
or ( \6036_b1 , \6032_b1 , \6035_b1 );
xor ( \6036_b0 , \6032_b0 , w_14668 );
not ( w_14668 , w_14669 );
and ( w_14669 , \6035_b1 , \6035_b0 );
or ( \6037_b1 , \6035_b1 , \6009_b1 );
xor ( \6037_b0 , \6035_b0 , w_14670 );
not ( w_14670 , w_14671 );
and ( w_14671 , \6009_b1 , \6009_b0 );
buf ( \6038_b1 , \6037_b1 );
not ( \6038_b1 , w_14672 );
not ( \6038_b0 , w_14673 );
and ( w_14672 , w_14673 , \6037_b0 );
or ( \6039_b1 , \6036_b1 , \6038_b1 );
not ( \6038_b1 , w_14674 );
and ( \6039_b0 , \6036_b0 , w_14675 );
and ( w_14674 , w_14675 , \6038_b0 );
or ( \6040_b1 , \6029_b1 , \6039_b1 );
not ( \6039_b1 , w_14676 );
and ( \6040_b0 , \6029_b0 , w_14677 );
and ( w_14676 , w_14677 , \6039_b0 );
buf ( \6041_b1 , RIa166d60_28_b1 );
buf ( \6041_b0 , RIa166d60_28_b0 );
or ( \6042_b1 , \6041_b1 , \6037_b1 );
not ( \6037_b1 , w_14678 );
and ( \6042_b0 , \6041_b0 , w_14679 );
and ( w_14678 , w_14679 , \6037_b0 );
or ( \6043_b1 , \6040_b1 , w_14681 );
not ( w_14681 , w_14682 );
and ( \6043_b0 , \6040_b0 , w_14683 );
and ( w_14682 ,  , w_14683 );
buf ( w_14681 , \6042_b1 );
not ( w_14681 , w_14684 );
not (  , w_14685 );
and ( w_14684 , w_14685 , \6042_b0 );
or ( \6044_b1 , \6035_b1 , \6009_b1 );
not ( \6009_b1 , w_14686 );
and ( \6044_b0 , \6035_b0 , w_14687 );
and ( w_14686 , w_14687 , \6009_b0 );
buf ( \6045_b1 , \6044_b1 );
not ( \6045_b1 , w_14688 );
not ( \6045_b0 , w_14689 );
and ( w_14688 , w_14689 , \6044_b0 );
or ( \6046_b1 , \6032_b1 , \6045_b1 );
not ( \6045_b1 , w_14690 );
and ( \6046_b0 , \6032_b0 , w_14691 );
and ( w_14690 , w_14691 , \6045_b0 );
or ( \6047_b1 , \6043_b1 , w_14692 );
xor ( \6047_b0 , \6043_b0 , w_14694 );
not ( w_14694 , w_14695 );
and ( w_14695 , w_14692 , w_14693 );
buf ( w_14692 , \6046_b1 );
not ( w_14692 , w_14696 );
not ( w_14693 , w_14697 );
and ( w_14696 , w_14697 , \6046_b0 );
buf ( \6048_b1 , RIb4ca4d8_31_b1 );
buf ( \6048_b0 , RIb4ca4d8_31_b0 );
or ( \6049_b1 , \735_b1 , \5718_b1 );
xor ( \6049_b0 , \735_b0 , w_14698 );
not ( w_14698 , w_14699 );
and ( w_14699 , \5718_b1 , \5718_b0 );
buf ( \6050_b1 , \6049_b1 );
buf ( \6050_b0 , \6049_b0 );
buf ( \6051_b1 , \6050_b1 );
buf ( \6051_b0 , \6050_b0 );
or ( \6052_b1 , \5733_b1 , \6051_b1 );
xor ( \6052_b0 , \5733_b0 , w_14700 );
not ( w_14700 , w_14701 );
and ( w_14701 , \6051_b1 , \6051_b0 );
or ( \6053_b1 , \6051_b1 , \6032_b1 );
xor ( \6053_b0 , \6051_b0 , w_14702 );
not ( w_14702 , w_14703 );
and ( w_14703 , \6032_b1 , \6032_b0 );
buf ( \6054_b1 , \6053_b1 );
not ( \6054_b1 , w_14704 );
not ( \6054_b0 , w_14705 );
and ( w_14704 , w_14705 , \6053_b0 );
or ( \6055_b1 , \6052_b1 , \6054_b1 );
not ( \6054_b1 , w_14706 );
and ( \6055_b0 , \6052_b0 , w_14707 );
and ( w_14706 , w_14707 , \6054_b0 );
or ( \6056_b1 , \6048_b1 , \6055_b1 );
not ( \6055_b1 , w_14708 );
and ( \6056_b0 , \6048_b0 , w_14709 );
and ( w_14708 , w_14709 , \6055_b0 );
buf ( \6057_b1 , RIa166c70_30_b1 );
buf ( \6057_b0 , RIa166c70_30_b0 );
or ( \6058_b1 , \6057_b1 , \6053_b1 );
not ( \6053_b1 , w_14710 );
and ( \6058_b0 , \6057_b0 , w_14711 );
and ( w_14710 , w_14711 , \6053_b0 );
or ( \6059_b1 , \6056_b1 , w_14713 );
not ( w_14713 , w_14714 );
and ( \6059_b0 , \6056_b0 , w_14715 );
and ( w_14714 ,  , w_14715 );
buf ( w_14713 , \6058_b1 );
not ( w_14713 , w_14716 );
not (  , w_14717 );
and ( w_14716 , w_14717 , \6058_b0 );
or ( \6060_b1 , \6051_b1 , \6032_b1 );
not ( \6032_b1 , w_14718 );
and ( \6060_b0 , \6051_b0 , w_14719 );
and ( w_14718 , w_14719 , \6032_b0 );
buf ( \6061_b1 , \6060_b1 );
not ( \6061_b1 , w_14720 );
not ( \6061_b0 , w_14721 );
and ( w_14720 , w_14721 , \6060_b0 );
or ( \6062_b1 , \5733_b1 , \6061_b1 );
not ( \6061_b1 , w_14722 );
and ( \6062_b0 , \5733_b0 , w_14723 );
and ( w_14722 , w_14723 , \6061_b0 );
or ( \6063_b1 , \6059_b1 , w_14724 );
xor ( \6063_b0 , \6059_b0 , w_14726 );
not ( w_14726 , w_14727 );
and ( w_14727 , w_14724 , w_14725 );
buf ( w_14724 , \6062_b1 );
not ( w_14724 , w_14728 );
not ( w_14725 , w_14729 );
and ( w_14728 , w_14729 , \6062_b0 );
or ( \6064_b1 , \6047_b1 , \6063_b1 );
not ( \6063_b1 , w_14730 );
and ( \6064_b0 , \6047_b0 , w_14731 );
and ( w_14730 , w_14731 , \6063_b0 );
buf ( \6065_b1 , RIb4ca460_32_b1 );
buf ( \6065_b0 , RIb4ca460_32_b0 );
or ( \6066_b1 , \5730_b1 , \5733_b1 );
xor ( \6066_b0 , \5730_b0 , w_14732 );
not ( w_14732 , w_14733 );
and ( w_14733 , \5733_b1 , \5733_b0 );
or ( \6067_b1 , \6065_b1 , w_14735 );
not ( w_14735 , w_14736 );
and ( \6067_b0 , \6065_b0 , w_14737 );
and ( w_14736 ,  , w_14737 );
buf ( w_14735 , \6066_b1 );
not ( w_14735 , w_14738 );
not (  , w_14739 );
and ( w_14738 , w_14739 , \6066_b0 );
or ( \6068_b1 , \6067_b1 , w_14740 );
xor ( \6068_b0 , \6067_b0 , w_14742 );
not ( w_14742 , w_14743 );
and ( w_14743 , w_14740 , w_14741 );
buf ( w_14740 , \5736_b1 );
not ( w_14740 , w_14744 );
not ( w_14741 , w_14745 );
and ( w_14744 , w_14745 , \5736_b0 );
or ( \6069_b1 , \6063_b1 , \6068_b1 );
not ( \6068_b1 , w_14746 );
and ( \6069_b0 , \6063_b0 , w_14747 );
and ( w_14746 , w_14747 , \6068_b0 );
or ( \6070_b1 , \6047_b1 , \6068_b1 );
not ( \6068_b1 , w_14748 );
and ( \6070_b0 , \6047_b0 , w_14749 );
and ( w_14748 , w_14749 , \6068_b0 );
or ( \6072_b1 , \6027_b1 , \6071_b1 );
not ( \6071_b1 , w_14750 );
and ( \6072_b0 , \6027_b0 , w_14751 );
and ( w_14750 , w_14751 , \6071_b0 );
or ( \6073_b1 , \5966_b1 , \6071_b1 );
not ( \6071_b1 , w_14752 );
and ( \6073_b0 , \5966_b0 , w_14753 );
and ( w_14752 , w_14753 , \6071_b0 );
or ( \6075_b1 , \5905_b1 , \6074_b1 );
not ( \6074_b1 , w_14754 );
and ( \6075_b0 , \5905_b0 , w_14755 );
and ( w_14754 , w_14755 , \6074_b0 );
or ( \6076_b1 , \6057_b1 , \6055_b1 );
not ( \6055_b1 , w_14756 );
and ( \6076_b0 , \6057_b0 , w_14757 );
and ( w_14756 , w_14757 , \6055_b0 );
or ( \6077_b1 , \6029_b1 , \6053_b1 );
not ( \6053_b1 , w_14758 );
and ( \6077_b0 , \6029_b0 , w_14759 );
and ( w_14758 , w_14759 , \6053_b0 );
or ( \6078_b1 , \6076_b1 , w_14761 );
not ( w_14761 , w_14762 );
and ( \6078_b0 , \6076_b0 , w_14763 );
and ( w_14762 ,  , w_14763 );
buf ( w_14761 , \6077_b1 );
not ( w_14761 , w_14764 );
not (  , w_14765 );
and ( w_14764 , w_14765 , \6077_b0 );
or ( \6079_b1 , \6078_b1 , w_14766 );
xor ( \6079_b0 , \6078_b0 , w_14768 );
not ( w_14768 , w_14769 );
and ( w_14769 , w_14766 , w_14767 );
buf ( w_14766 , \6062_b1 );
not ( w_14766 , w_14770 );
not ( w_14767 , w_14771 );
and ( w_14770 , w_14771 , \6062_b0 );
or ( \6080_b1 , \5727_b1 , \5730_b1 );
xor ( \6080_b0 , \5727_b0 , w_14772 );
not ( w_14772 , w_14773 );
and ( w_14773 , \5730_b1 , \5730_b0 );
buf ( \6081_b1 , \6066_b1 );
not ( \6081_b1 , w_14774 );
not ( \6081_b0 , w_14775 );
and ( w_14774 , w_14775 , \6066_b0 );
or ( \6082_b1 , \6080_b1 , \6081_b1 );
not ( \6081_b1 , w_14776 );
and ( \6082_b0 , \6080_b0 , w_14777 );
and ( w_14776 , w_14777 , \6081_b0 );
or ( \6083_b1 , \6065_b1 , \6082_b1 );
not ( \6082_b1 , w_14778 );
and ( \6083_b0 , \6065_b0 , w_14779 );
and ( w_14778 , w_14779 , \6082_b0 );
or ( \6084_b1 , \6048_b1 , \6066_b1 );
not ( \6066_b1 , w_14780 );
and ( \6084_b0 , \6048_b0 , w_14781 );
and ( w_14780 , w_14781 , \6066_b0 );
or ( \6085_b1 , \6083_b1 , w_14783 );
not ( w_14783 , w_14784 );
and ( \6085_b0 , \6083_b0 , w_14785 );
and ( w_14784 ,  , w_14785 );
buf ( w_14783 , \6084_b1 );
not ( w_14783 , w_14786 );
not (  , w_14787 );
and ( w_14786 , w_14787 , \6084_b0 );
or ( \6086_b1 , \6085_b1 , w_14788 );
xor ( \6086_b0 , \6085_b0 , w_14790 );
not ( w_14790 , w_14791 );
and ( w_14791 , w_14788 , w_14789 );
buf ( w_14788 , \5736_b1 );
not ( w_14788 , w_14792 );
not ( w_14789 , w_14793 );
and ( w_14792 , w_14793 , \5736_b0 );
or ( \6087_b1 , \6079_b1 , \6086_b1 );
xor ( \6087_b0 , \6079_b0 , w_14794 );
not ( w_14794 , w_14795 );
and ( w_14795 , \6086_b1 , \6086_b0 );
or ( \6088_b1 , \5998_b1 , \5996_b1 );
not ( \5996_b1 , w_14796 );
and ( \6088_b0 , \5998_b0 , w_14797 );
and ( w_14796 , w_14797 , \5996_b0 );
or ( \6089_b1 , \5967_b1 , \5994_b1 );
not ( \5994_b1 , w_14798 );
and ( \6089_b0 , \5967_b0 , w_14799 );
and ( w_14798 , w_14799 , \5994_b0 );
or ( \6090_b1 , \6088_b1 , w_14801 );
not ( w_14801 , w_14802 );
and ( \6090_b0 , \6088_b0 , w_14803 );
and ( w_14802 ,  , w_14803 );
buf ( w_14801 , \6089_b1 );
not ( w_14801 , w_14804 );
not (  , w_14805 );
and ( w_14804 , w_14805 , \6089_b0 );
or ( \6091_b1 , \6090_b1 , w_14806 );
xor ( \6091_b0 , \6090_b0 , w_14808 );
not ( w_14808 , w_14809 );
and ( w_14809 , w_14806 , w_14807 );
buf ( w_14806 , \6003_b1 );
not ( w_14806 , w_14810 );
not ( w_14807 , w_14811 );
and ( w_14810 , w_14811 , \6003_b0 );
or ( \6092_b1 , \6018_b1 , \6016_b1 );
not ( \6016_b1 , w_14812 );
and ( \6092_b0 , \6018_b0 , w_14813 );
and ( w_14812 , w_14813 , \6016_b0 );
or ( \6093_b1 , \5986_b1 , \6014_b1 );
not ( \6014_b1 , w_14814 );
and ( \6093_b0 , \5986_b0 , w_14815 );
and ( w_14814 , w_14815 , \6014_b0 );
or ( \6094_b1 , \6092_b1 , w_14817 );
not ( w_14817 , w_14818 );
and ( \6094_b0 , \6092_b0 , w_14819 );
and ( w_14818 ,  , w_14819 );
buf ( w_14817 , \6093_b1 );
not ( w_14817 , w_14820 );
not (  , w_14821 );
and ( w_14820 , w_14821 , \6093_b0 );
or ( \6095_b1 , \6094_b1 , w_14822 );
xor ( \6095_b0 , \6094_b0 , w_14824 );
not ( w_14824 , w_14825 );
and ( w_14825 , w_14822 , w_14823 );
buf ( w_14822 , \6023_b1 );
not ( w_14822 , w_14826 );
not ( w_14823 , w_14827 );
and ( w_14826 , w_14827 , \6023_b0 );
or ( \6096_b1 , \6091_b1 , \6095_b1 );
xor ( \6096_b0 , \6091_b0 , w_14828 );
not ( w_14828 , w_14829 );
and ( w_14829 , \6095_b1 , \6095_b0 );
or ( \6097_b1 , \6041_b1 , \6039_b1 );
not ( \6039_b1 , w_14830 );
and ( \6097_b0 , \6041_b0 , w_14831 );
and ( w_14830 , w_14831 , \6039_b0 );
or ( \6098_b1 , \6006_b1 , \6037_b1 );
not ( \6037_b1 , w_14832 );
and ( \6098_b0 , \6006_b0 , w_14833 );
and ( w_14832 , w_14833 , \6037_b0 );
or ( \6099_b1 , \6097_b1 , w_14835 );
not ( w_14835 , w_14836 );
and ( \6099_b0 , \6097_b0 , w_14837 );
and ( w_14836 ,  , w_14837 );
buf ( w_14835 , \6098_b1 );
not ( w_14835 , w_14838 );
not (  , w_14839 );
and ( w_14838 , w_14839 , \6098_b0 );
or ( \6100_b1 , \6099_b1 , w_14840 );
xor ( \6100_b0 , \6099_b0 , w_14842 );
not ( w_14842 , w_14843 );
and ( w_14843 , w_14840 , w_14841 );
buf ( w_14840 , \6046_b1 );
not ( w_14840 , w_14844 );
not ( w_14841 , w_14845 );
and ( w_14844 , w_14845 , \6046_b0 );
or ( \6101_b1 , \6096_b1 , \6100_b1 );
xor ( \6101_b0 , \6096_b0 , w_14846 );
not ( w_14846 , w_14847 );
and ( w_14847 , \6100_b1 , \6100_b0 );
or ( \6102_b1 , \6087_b1 , \6101_b1 );
not ( \6101_b1 , w_14848 );
and ( \6102_b0 , \6087_b0 , w_14849 );
and ( w_14848 , w_14849 , \6101_b0 );
or ( \6103_b1 , \5937_b1 , \5935_b1 );
not ( \5935_b1 , w_14850 );
and ( \6103_b0 , \5937_b0 , w_14851 );
and ( w_14850 , w_14851 , \5935_b0 );
or ( \6104_b1 , \5906_b1 , \5933_b1 );
not ( \5933_b1 , w_14852 );
and ( \6104_b0 , \5906_b0 , w_14853 );
and ( w_14852 , w_14853 , \5933_b0 );
or ( \6105_b1 , \6103_b1 , w_14855 );
not ( w_14855 , w_14856 );
and ( \6105_b0 , \6103_b0 , w_14857 );
and ( w_14856 ,  , w_14857 );
buf ( w_14855 , \6104_b1 );
not ( w_14855 , w_14858 );
not (  , w_14859 );
and ( w_14858 , w_14859 , \6104_b0 );
or ( \6106_b1 , \6105_b1 , w_14860 );
xor ( \6106_b0 , \6105_b0 , w_14862 );
not ( w_14862 , w_14863 );
and ( w_14863 , w_14860 , w_14861 );
buf ( w_14860 , \5942_b1 );
not ( w_14860 , w_14864 );
not ( w_14861 , w_14865 );
and ( w_14864 , w_14865 , \5942_b0 );
or ( \6107_b1 , \5957_b1 , \5955_b1 );
not ( \5955_b1 , w_14866 );
and ( \6107_b0 , \5957_b0 , w_14867 );
and ( w_14866 , w_14867 , \5955_b0 );
or ( \6108_b1 , \5925_b1 , \5953_b1 );
not ( \5953_b1 , w_14868 );
and ( \6108_b0 , \5925_b0 , w_14869 );
and ( w_14868 , w_14869 , \5953_b0 );
or ( \6109_b1 , \6107_b1 , w_14871 );
not ( w_14871 , w_14872 );
and ( \6109_b0 , \6107_b0 , w_14873 );
and ( w_14872 ,  , w_14873 );
buf ( w_14871 , \6108_b1 );
not ( w_14871 , w_14874 );
not (  , w_14875 );
and ( w_14874 , w_14875 , \6108_b0 );
or ( \6110_b1 , \6109_b1 , w_14876 );
xor ( \6110_b0 , \6109_b0 , w_14878 );
not ( w_14878 , w_14879 );
and ( w_14879 , w_14876 , w_14877 );
buf ( w_14876 , \5962_b1 );
not ( w_14876 , w_14880 );
not ( w_14877 , w_14881 );
and ( w_14880 , w_14881 , \5962_b0 );
or ( \6111_b1 , \6106_b1 , \6110_b1 );
xor ( \6111_b0 , \6106_b0 , w_14882 );
not ( w_14882 , w_14883 );
and ( w_14883 , \6110_b1 , \6110_b0 );
or ( \6112_b1 , \5979_b1 , \5977_b1 );
not ( \5977_b1 , w_14884 );
and ( \6112_b0 , \5979_b0 , w_14885 );
and ( w_14884 , w_14885 , \5977_b0 );
or ( \6113_b1 , \5945_b1 , \5975_b1 );
not ( \5975_b1 , w_14886 );
and ( \6113_b0 , \5945_b0 , w_14887 );
and ( w_14886 , w_14887 , \5975_b0 );
or ( \6114_b1 , \6112_b1 , w_14889 );
not ( w_14889 , w_14890 );
and ( \6114_b0 , \6112_b0 , w_14891 );
and ( w_14890 ,  , w_14891 );
buf ( w_14889 , \6113_b1 );
not ( w_14889 , w_14892 );
not (  , w_14893 );
and ( w_14892 , w_14893 , \6113_b0 );
or ( \6115_b1 , \6114_b1 , w_14894 );
xor ( \6115_b0 , \6114_b0 , w_14896 );
not ( w_14896 , w_14897 );
and ( w_14897 , w_14894 , w_14895 );
buf ( w_14894 , \5984_b1 );
not ( w_14894 , w_14898 );
not ( w_14895 , w_14899 );
and ( w_14898 , w_14899 , \5984_b0 );
or ( \6116_b1 , \6111_b1 , \6115_b1 );
xor ( \6116_b0 , \6111_b0 , w_14900 );
not ( w_14900 , w_14901 );
and ( w_14901 , \6115_b1 , \6115_b0 );
or ( \6117_b1 , \6101_b1 , \6116_b1 );
not ( \6116_b1 , w_14902 );
and ( \6117_b0 , \6101_b0 , w_14903 );
and ( w_14902 , w_14903 , \6116_b0 );
or ( \6118_b1 , \6087_b1 , \6116_b1 );
not ( \6116_b1 , w_14904 );
and ( \6118_b0 , \6087_b0 , w_14905 );
and ( w_14904 , w_14905 , \6116_b0 );
or ( \6120_b1 , \6074_b1 , \6119_b1 );
not ( \6119_b1 , w_14906 );
and ( \6120_b0 , \6074_b0 , w_14907 );
and ( w_14906 , w_14907 , \6119_b0 );
or ( \6121_b1 , \5905_b1 , \6119_b1 );
not ( \6119_b1 , w_14908 );
and ( \6121_b0 , \5905_b0 , w_14909 );
and ( w_14908 , w_14909 , \6119_b0 );
or ( \6123_b1 , \5873_b1 , \5871_b1 );
not ( \5871_b1 , w_14910 );
and ( \6123_b0 , \5873_b0 , w_14911 );
and ( w_14910 , w_14911 , \5871_b0 );
or ( \6124_b1 , \5842_b1 , \5869_b1 );
not ( \5869_b1 , w_14912 );
and ( \6124_b0 , \5842_b0 , w_14913 );
and ( w_14912 , w_14913 , \5869_b0 );
or ( \6125_b1 , \6123_b1 , w_14915 );
not ( w_14915 , w_14916 );
and ( \6125_b0 , \6123_b0 , w_14917 );
and ( w_14916 ,  , w_14917 );
buf ( w_14915 , \6124_b1 );
not ( w_14915 , w_14918 );
not (  , w_14919 );
and ( w_14918 , w_14919 , \6124_b0 );
or ( \6126_b1 , \6125_b1 , w_14920 );
xor ( \6126_b0 , \6125_b0 , w_14922 );
not ( w_14922 , w_14923 );
and ( w_14923 , w_14920 , w_14921 );
buf ( w_14920 , \5878_b1 );
not ( w_14920 , w_14924 );
not ( w_14921 , w_14925 );
and ( w_14924 , w_14925 , \5878_b0 );
or ( \6127_b1 , \5893_b1 , \5891_b1 );
not ( \5891_b1 , w_14926 );
and ( \6127_b0 , \5893_b0 , w_14927 );
and ( w_14926 , w_14927 , \5891_b0 );
or ( \6128_b1 , \5861_b1 , \5889_b1 );
not ( \5889_b1 , w_14928 );
and ( \6128_b0 , \5861_b0 , w_14929 );
and ( w_14928 , w_14929 , \5889_b0 );
or ( \6129_b1 , \6127_b1 , w_14931 );
not ( w_14931 , w_14932 );
and ( \6129_b0 , \6127_b0 , w_14933 );
and ( w_14932 ,  , w_14933 );
buf ( w_14931 , \6128_b1 );
not ( w_14931 , w_14934 );
not (  , w_14935 );
and ( w_14934 , w_14935 , \6128_b0 );
or ( \6130_b1 , \6129_b1 , w_14936 );
xor ( \6130_b0 , \6129_b0 , w_14938 );
not ( w_14938 , w_14939 );
and ( w_14939 , w_14936 , w_14937 );
buf ( w_14936 , \5898_b1 );
not ( w_14936 , w_14940 );
not ( w_14937 , w_14941 );
and ( w_14940 , w_14941 , \5898_b0 );
or ( \6131_b1 , \6126_b1 , \6130_b1 );
xor ( \6131_b0 , \6126_b0 , w_14942 );
not ( w_14942 , w_14943 );
and ( w_14943 , \6130_b1 , \6130_b0 );
or ( \6132_b1 , \5918_b1 , \5916_b1 );
not ( \5916_b1 , w_14944 );
and ( \6132_b0 , \5918_b0 , w_14945 );
and ( w_14944 , w_14945 , \5916_b0 );
or ( \6133_b1 , \5881_b1 , \5914_b1 );
not ( \5914_b1 , w_14946 );
and ( \6133_b0 , \5881_b0 , w_14947 );
and ( w_14946 , w_14947 , \5914_b0 );
or ( \6134_b1 , \6132_b1 , w_14949 );
not ( w_14949 , w_14950 );
and ( \6134_b0 , \6132_b0 , w_14951 );
and ( w_14950 ,  , w_14951 );
buf ( w_14949 , \6133_b1 );
not ( w_14949 , w_14952 );
not (  , w_14953 );
and ( w_14952 , w_14953 , \6133_b0 );
or ( \6135_b1 , \6134_b1 , w_14954 );
xor ( \6135_b0 , \6134_b0 , w_14956 );
not ( w_14956 , w_14957 );
and ( w_14957 , w_14954 , w_14955 );
buf ( w_14954 , \5923_b1 );
not ( w_14954 , w_14958 );
not ( w_14955 , w_14959 );
and ( w_14958 , w_14959 , \5923_b0 );
or ( \6136_b1 , \6131_b1 , \6135_b1 );
xor ( \6136_b0 , \6131_b0 , w_14960 );
not ( w_14960 , w_14961 );
and ( w_14961 , \6135_b1 , \6135_b0 );
or ( \6137_b1 , \5811_b1 , \5809_b1 );
not ( \5809_b1 , w_14962 );
and ( \6137_b0 , \5811_b0 , w_14963 );
and ( w_14962 , w_14963 , \5809_b0 );
or ( \6138_b1 , \5780_b1 , \5807_b1 );
not ( \5807_b1 , w_14964 );
and ( \6138_b0 , \5780_b0 , w_14965 );
and ( w_14964 , w_14965 , \5807_b0 );
or ( \6139_b1 , \6137_b1 , w_14967 );
not ( w_14967 , w_14968 );
and ( \6139_b0 , \6137_b0 , w_14969 );
and ( w_14968 ,  , w_14969 );
buf ( w_14967 , \6138_b1 );
not ( w_14967 , w_14970 );
not (  , w_14971 );
and ( w_14970 , w_14971 , \6138_b0 );
or ( \6140_b1 , \6139_b1 , w_14972 );
xor ( \6140_b0 , \6139_b0 , w_14974 );
not ( w_14974 , w_14975 );
and ( w_14975 , w_14972 , w_14973 );
buf ( w_14972 , \5816_b1 );
not ( w_14972 , w_14976 );
not ( w_14973 , w_14977 );
and ( w_14976 , w_14977 , \5816_b0 );
or ( \6141_b1 , \5831_b1 , \5829_b1 );
not ( \5829_b1 , w_14978 );
and ( \6141_b0 , \5831_b0 , w_14979 );
and ( w_14978 , w_14979 , \5829_b0 );
or ( \6142_b1 , \5799_b1 , \5827_b1 );
not ( \5827_b1 , w_14980 );
and ( \6142_b0 , \5799_b0 , w_14981 );
and ( w_14980 , w_14981 , \5827_b0 );
or ( \6143_b1 , \6141_b1 , w_14983 );
not ( w_14983 , w_14984 );
and ( \6143_b0 , \6141_b0 , w_14985 );
and ( w_14984 ,  , w_14985 );
buf ( w_14983 , \6142_b1 );
not ( w_14983 , w_14986 );
not (  , w_14987 );
and ( w_14986 , w_14987 , \6142_b0 );
or ( \6144_b1 , \6143_b1 , w_14988 );
xor ( \6144_b0 , \6143_b0 , w_14990 );
not ( w_14990 , w_14991 );
and ( w_14991 , w_14988 , w_14989 );
buf ( w_14988 , \5836_b1 );
not ( w_14988 , w_14992 );
not ( w_14989 , w_14993 );
and ( w_14992 , w_14993 , \5836_b0 );
or ( \6145_b1 , \6140_b1 , \6144_b1 );
xor ( \6145_b0 , \6140_b0 , w_14994 );
not ( w_14994 , w_14995 );
and ( w_14995 , \6144_b1 , \6144_b0 );
or ( \6146_b1 , \5854_b1 , \5852_b1 );
not ( \5852_b1 , w_14996 );
and ( \6146_b0 , \5854_b0 , w_14997 );
and ( w_14996 , w_14997 , \5852_b0 );
or ( \6147_b1 , \5819_b1 , \5850_b1 );
not ( \5850_b1 , w_14998 );
and ( \6147_b0 , \5819_b0 , w_14999 );
and ( w_14998 , w_14999 , \5850_b0 );
or ( \6148_b1 , \6146_b1 , w_15001 );
not ( w_15001 , w_15002 );
and ( \6148_b0 , \6146_b0 , w_15003 );
and ( w_15002 ,  , w_15003 );
buf ( w_15001 , \6147_b1 );
not ( w_15001 , w_15004 );
not (  , w_15005 );
and ( w_15004 , w_15005 , \6147_b0 );
or ( \6149_b1 , \6148_b1 , w_15006 );
xor ( \6149_b0 , \6148_b0 , w_15008 );
not ( w_15008 , w_15009 );
and ( w_15009 , w_15006 , w_15007 );
buf ( w_15006 , \5859_b1 );
not ( w_15006 , w_15010 );
not ( w_15007 , w_15011 );
and ( w_15010 , w_15011 , \5859_b0 );
or ( \6150_b1 , \6145_b1 , \6149_b1 );
xor ( \6150_b0 , \6145_b0 , w_15012 );
not ( w_15012 , w_15013 );
and ( w_15013 , \6149_b1 , \6149_b0 );
or ( \6151_b1 , \6136_b1 , \6150_b1 );
not ( \6150_b1 , w_15014 );
and ( \6151_b0 , \6136_b0 , w_15015 );
and ( w_15014 , w_15015 , \6150_b0 );
buf ( \6152_b1 , \5755_b1 );
not ( \6152_b1 , w_15016 );
not ( \6152_b0 , w_15017 );
and ( w_15016 , w_15017 , \5755_b0 );
or ( \6153_b1 , \5770_b1 , \5768_b1 );
not ( \5768_b1 , w_15018 );
and ( \6153_b0 , \5770_b0 , w_15019 );
and ( w_15018 , w_15019 , \5768_b0 );
or ( \6154_b1 , \5737_b1 , \5766_b1 );
not ( \5766_b1 , w_15020 );
and ( \6154_b0 , \5737_b0 , w_15021 );
and ( w_15020 , w_15021 , \5766_b0 );
or ( \6155_b1 , \6153_b1 , w_15023 );
not ( w_15023 , w_15024 );
and ( \6155_b0 , \6153_b0 , w_15025 );
and ( w_15024 ,  , w_15025 );
buf ( w_15023 , \6154_b1 );
not ( w_15023 , w_15026 );
not (  , w_15027 );
and ( w_15026 , w_15027 , \6154_b0 );
or ( \6156_b1 , \6155_b1 , w_15028 );
xor ( \6156_b0 , \6155_b0 , w_15030 );
not ( w_15030 , w_15031 );
and ( w_15031 , w_15028 , w_15029 );
buf ( w_15028 , \5775_b1 );
not ( w_15028 , w_15032 );
not ( w_15029 , w_15033 );
and ( w_15032 , w_15033 , \5775_b0 );
or ( \6157_b1 , \6152_b1 , \6156_b1 );
xor ( \6157_b0 , \6152_b0 , w_15034 );
not ( w_15034 , w_15035 );
and ( w_15035 , \6156_b1 , \6156_b0 );
or ( \6158_b1 , \5792_b1 , \5790_b1 );
not ( \5790_b1 , w_15036 );
and ( \6158_b0 , \5792_b0 , w_15037 );
and ( w_15036 , w_15037 , \5790_b0 );
or ( \6159_b1 , \5758_b1 , \5788_b1 );
not ( \5788_b1 , w_15038 );
and ( \6159_b0 , \5758_b0 , w_15039 );
and ( w_15038 , w_15039 , \5788_b0 );
or ( \6160_b1 , \6158_b1 , w_15041 );
not ( w_15041 , w_15042 );
and ( \6160_b0 , \6158_b0 , w_15043 );
and ( w_15042 ,  , w_15043 );
buf ( w_15041 , \6159_b1 );
not ( w_15041 , w_15044 );
not (  , w_15045 );
and ( w_15044 , w_15045 , \6159_b0 );
or ( \6161_b1 , \6160_b1 , w_15046 );
xor ( \6161_b0 , \6160_b0 , w_15048 );
not ( w_15048 , w_15049 );
and ( w_15049 , w_15046 , w_15047 );
buf ( w_15046 , \5797_b1 );
not ( w_15046 , w_15050 );
not ( w_15047 , w_15051 );
and ( w_15050 , w_15051 , \5797_b0 );
or ( \6162_b1 , \6157_b1 , \6161_b1 );
xor ( \6162_b0 , \6157_b0 , w_15052 );
not ( w_15052 , w_15053 );
and ( w_15053 , \6161_b1 , \6161_b0 );
or ( \6163_b1 , \6150_b1 , \6162_b1 );
not ( \6162_b1 , w_15054 );
and ( \6163_b0 , \6150_b0 , w_15055 );
and ( w_15054 , w_15055 , \6162_b0 );
or ( \6164_b1 , \6136_b1 , \6162_b1 );
not ( \6162_b1 , w_15056 );
and ( \6164_b0 , \6136_b0 , w_15057 );
and ( w_15056 , w_15057 , \6162_b0 );
or ( \6166_b1 , \159_b1 , \331_b1 );
not ( \331_b1 , w_15058 );
and ( \6166_b0 , \159_b0 , w_15059 );
and ( w_15058 , w_15059 , \331_b0 );
buf ( \6167_b1 , \6166_b1 );
not ( \6167_b1 , w_15060 );
not ( \6167_b0 , w_15061 );
and ( w_15060 , w_15061 , \6166_b0 );
or ( \6168_b1 , \6167_b1 , w_15062 );
xor ( \6168_b0 , \6167_b0 , w_15064 );
not ( w_15064 , w_15065 );
and ( w_15065 , w_15062 , w_15063 );
buf ( w_15062 , \338_b1 );
not ( w_15062 , w_15066 );
not ( w_15063 , w_15067 );
and ( w_15066 , w_15067 , \338_b0 );
or ( \6169_b1 , \305_b1 , \351_b1 );
not ( \351_b1 , w_15068 );
and ( \6169_b0 , \305_b0 , w_15069 );
and ( w_15068 , w_15069 , \351_b0 );
or ( \6170_b1 , \315_b1 , \349_b1 );
not ( \349_b1 , w_15070 );
and ( \6170_b0 , \315_b0 , w_15071 );
and ( w_15070 , w_15071 , \349_b0 );
or ( \6171_b1 , \6169_b1 , w_15073 );
not ( w_15073 , w_15074 );
and ( \6171_b0 , \6169_b0 , w_15075 );
and ( w_15074 ,  , w_15075 );
buf ( w_15073 , \6170_b1 );
not ( w_15073 , w_15076 );
not (  , w_15077 );
and ( w_15076 , w_15077 , \6170_b0 );
or ( \6172_b1 , \6171_b1 , w_15078 );
xor ( \6172_b0 , \6171_b0 , w_15080 );
not ( w_15080 , w_15081 );
and ( w_15081 , w_15078 , w_15079 );
buf ( w_15078 , \358_b1 );
not ( w_15078 , w_15082 );
not ( w_15079 , w_15083 );
and ( w_15082 , w_15083 , \358_b0 );
or ( \6173_b1 , \6168_b1 , \6172_b1 );
not ( \6172_b1 , w_15084 );
and ( \6173_b0 , \6168_b0 , w_15085 );
and ( w_15084 , w_15085 , \6172_b0 );
or ( \6174_b1 , \333_b1 , \345_b1 );
not ( \345_b1 , w_15086 );
and ( \6174_b0 , \333_b0 , w_15087 );
and ( w_15086 , w_15087 , \345_b0 );
or ( \6175_b1 , \6172_b1 , \6174_b1 );
not ( \6174_b1 , w_15088 );
and ( \6175_b0 , \6172_b0 , w_15089 );
and ( w_15088 , w_15089 , \6174_b0 );
or ( \6176_b1 , \6168_b1 , \6174_b1 );
not ( \6174_b1 , w_15090 );
and ( \6176_b0 , \6168_b0 , w_15091 );
and ( w_15090 , w_15091 , \6174_b0 );
or ( \6178_b1 , \413_b1 , \417_b1 );
not ( \417_b1 , w_15092 );
and ( \6178_b0 , \413_b0 , w_15093 );
and ( w_15092 , w_15093 , \417_b0 );
or ( \6179_b1 , \417_b1 , \422_b1 );
not ( \422_b1 , w_15094 );
and ( \6179_b0 , \417_b0 , w_15095 );
and ( w_15094 , w_15095 , \422_b0 );
or ( \6180_b1 , \413_b1 , \422_b1 );
not ( \422_b1 , w_15096 );
and ( \6180_b0 , \413_b0 , w_15097 );
and ( w_15096 , w_15097 , \422_b0 );
or ( \6182_b1 , \6168_b1 , \6172_b1 );
xor ( \6182_b0 , \6168_b0 , w_15098 );
not ( w_15098 , w_15099 );
and ( w_15099 , \6172_b1 , \6172_b0 );
or ( \6183_b1 , \6182_b1 , \6174_b1 );
xor ( \6183_b0 , \6182_b0 , w_15100 );
not ( w_15100 , w_15101 );
and ( w_15101 , \6174_b1 , \6174_b0 );
or ( \6184_b1 , \6181_b1 , w_15102 );
or ( \6184_b0 , \6181_b0 , \6183_b0 );
not ( \6183_b0 , w_15103 );
and ( w_15103 , w_15102 , \6183_b1 );
or ( \6185_b1 , \6177_b1 , \6184_b1 );
xor ( \6185_b0 , \6177_b0 , w_15104 );
not ( w_15104 , w_15105 );
and ( w_15105 , \6184_b1 , \6184_b0 );
buf ( \6186_b1 , \338_b1 );
not ( \6186_b1 , w_15106 );
not ( \6186_b0 , w_15107 );
and ( w_15106 , w_15107 , \338_b0 );
or ( \6187_b1 , \315_b1 , \351_b1 );
not ( \351_b1 , w_15108 );
and ( \6187_b0 , \315_b0 , w_15109 );
and ( w_15108 , w_15109 , \351_b0 );
or ( \6188_b1 , \159_b1 , \349_b1 );
not ( \349_b1 , w_15110 );
and ( \6188_b0 , \159_b0 , w_15111 );
and ( w_15110 , w_15111 , \349_b0 );
or ( \6189_b1 , \6187_b1 , w_15113 );
not ( w_15113 , w_15114 );
and ( \6189_b0 , \6187_b0 , w_15115 );
and ( w_15114 ,  , w_15115 );
buf ( w_15113 , \6188_b1 );
not ( w_15113 , w_15116 );
not (  , w_15117 );
and ( w_15116 , w_15117 , \6188_b0 );
or ( \6190_b1 , \6189_b1 , w_15118 );
xor ( \6190_b0 , \6189_b0 , w_15120 );
not ( w_15120 , w_15121 );
and ( w_15121 , w_15118 , w_15119 );
buf ( w_15118 , \358_b1 );
not ( w_15118 , w_15122 );
not ( w_15119 , w_15123 );
and ( w_15122 , w_15123 , \358_b0 );
or ( \6191_b1 , \6186_b1 , \6190_b1 );
xor ( \6191_b0 , \6186_b0 , w_15124 );
not ( w_15124 , w_15125 );
and ( w_15125 , \6190_b1 , \6190_b0 );
or ( \6192_b1 , \305_b1 , \345_b1 );
not ( \345_b1 , w_15126 );
and ( \6192_b0 , \305_b0 , w_15127 );
and ( w_15126 , w_15127 , \345_b0 );
or ( \6193_b1 , \6191_b1 , \6192_b1 );
xor ( \6193_b0 , \6191_b0 , w_15128 );
not ( w_15128 , w_15129 );
and ( w_15129 , \6192_b1 , \6192_b0 );
or ( \6194_b1 , \6185_b1 , \6193_b1 );
xor ( \6194_b0 , \6185_b0 , w_15130 );
not ( w_15130 , w_15131 );
and ( w_15131 , \6193_b1 , \6193_b0 );
or ( \6195_b1 , \428_b1 , \429_b1 );
not ( \429_b1 , w_15132 );
and ( \6195_b0 , \428_b0 , w_15133 );
and ( w_15132 , w_15133 , \429_b0 );
or ( \6196_b1 , \429_b1 , \431_b1 );
not ( \431_b1 , w_15134 );
and ( \6196_b0 , \429_b0 , w_15135 );
and ( w_15134 , w_15135 , \431_b0 );
or ( \6197_b1 , \428_b1 , \431_b1 );
not ( \431_b1 , w_15136 );
and ( \6197_b0 , \428_b0 , w_15137 );
and ( w_15136 , w_15137 , \431_b0 );
or ( \6199_b1 , \412_b1 , \423_b1 );
not ( \423_b1 , w_15138 );
and ( \6199_b0 , \412_b0 , w_15139 );
and ( w_15138 , w_15139 , \423_b0 );
or ( \6200_b1 , \423_b1 , \432_b1 );
not ( \432_b1 , w_15140 );
and ( \6200_b0 , \423_b0 , w_15141 );
and ( w_15140 , w_15141 , \432_b0 );
or ( \6201_b1 , \412_b1 , \432_b1 );
not ( \432_b1 , w_15142 );
and ( \6201_b0 , \412_b0 , w_15143 );
and ( w_15142 , w_15143 , \432_b0 );
or ( \6203_b1 , \6198_b1 , \6202_b1 );
not ( \6202_b1 , w_15144 );
and ( \6203_b0 , \6198_b0 , w_15145 );
and ( w_15144 , w_15145 , \6202_b0 );
or ( \6204_b1 , \6181_b1 , w_15146 );
xor ( \6204_b0 , \6181_b0 , w_15148 );
not ( w_15148 , w_15149 );
and ( w_15149 , w_15146 , w_15147 );
buf ( w_15146 , \6183_b1 );
not ( w_15146 , w_15150 );
not ( w_15147 , w_15151 );
and ( w_15150 , w_15151 , \6183_b0 );
or ( \6205_b1 , \6202_b1 , \6204_b1 );
not ( \6204_b1 , w_15152 );
and ( \6205_b0 , \6202_b0 , w_15153 );
and ( w_15152 , w_15153 , \6204_b0 );
or ( \6206_b1 , \6198_b1 , \6204_b1 );
not ( \6204_b1 , w_15154 );
and ( \6206_b0 , \6198_b0 , w_15155 );
and ( w_15154 , w_15155 , \6204_b0 );
or ( \6208_b1 , \6194_b1 , \6207_b1 );
xor ( \6208_b0 , \6194_b0 , w_15156 );
not ( w_15156 , w_15157 );
and ( w_15157 , \6207_b1 , \6207_b0 );
or ( \6209_b1 , \6198_b1 , \6202_b1 );
xor ( \6209_b0 , \6198_b0 , w_15158 );
not ( w_15158 , w_15159 );
and ( w_15159 , \6202_b1 , \6202_b0 );
or ( \6210_b1 , \6209_b1 , \6204_b1 );
xor ( \6210_b0 , \6209_b0 , w_15160 );
not ( w_15160 , w_15161 );
and ( w_15161 , \6204_b1 , \6204_b0 );
or ( \6211_b1 , \408_b1 , \433_b1 );
not ( \433_b1 , w_15162 );
and ( \6211_b0 , \408_b0 , w_15163 );
and ( w_15162 , w_15163 , \433_b0 );
or ( \6212_b1 , \6210_b1 , \6211_b1 );
not ( \6211_b1 , w_15164 );
and ( \6212_b0 , \6210_b0 , w_15165 );
and ( w_15164 , w_15165 , \6211_b0 );
or ( \6213_b1 , \6210_b1 , \6211_b1 );
xor ( \6213_b0 , \6210_b0 , w_15166 );
not ( w_15166 , w_15167 );
and ( w_15167 , \6211_b1 , \6211_b0 );
or ( \6214_b1 , \434_b1 , \483_b1 );
not ( \483_b1 , w_15168 );
and ( \6214_b0 , \434_b0 , w_15169 );
and ( w_15168 , w_15169 , \483_b0 );
or ( \6215_b1 , \484_b1 , \5724_b1 );
not ( \5724_b1 , w_15170 );
and ( \6215_b0 , \484_b0 , w_15171 );
and ( w_15170 , w_15171 , \5724_b0 );
or ( \6216_b1 , \6214_b1 , w_15172 );
or ( \6216_b0 , \6214_b0 , \6215_b0 );
not ( \6215_b0 , w_15173 );
and ( w_15173 , w_15172 , \6215_b1 );
or ( \6217_b1 , \6213_b1 , \6216_b1 );
not ( \6216_b1 , w_15174 );
and ( \6217_b0 , \6213_b0 , w_15175 );
and ( w_15174 , w_15175 , \6216_b0 );
or ( \6218_b1 , \6212_b1 , w_15176 );
or ( \6218_b0 , \6212_b0 , \6217_b0 );
not ( \6217_b0 , w_15177 );
and ( w_15177 , w_15176 , \6217_b1 );
or ( \6219_b1 , \6208_b1 , \6218_b1 );
xor ( \6219_b0 , \6208_b0 , w_15178 );
not ( w_15178 , w_15179 );
and ( w_15179 , \6218_b1 , \6218_b0 );
buf ( \6220_b1 , \6219_b1 );
buf ( \6220_b0 , \6219_b0 );
buf ( \6221_b1 , \6220_b1 );
buf ( \6221_b0 , \6220_b0 );
or ( \6222_b1 , \6213_b1 , \6216_b1 );
xor ( \6222_b0 , \6213_b0 , w_15180 );
not ( w_15180 , w_15181 );
and ( w_15181 , \6216_b1 , \6216_b0 );
buf ( \6223_b1 , \6222_b1 );
buf ( \6223_b0 , \6222_b0 );
buf ( \6224_b1 , \6223_b1 );
buf ( \6224_b0 , \6223_b0 );
or ( \6225_b1 , \6224_b1 , \5727_b1 );
not ( \5727_b1 , w_15182 );
and ( \6225_b0 , \6224_b0 , w_15183 );
and ( w_15182 , w_15183 , \5727_b0 );
buf ( \6226_b1 , \6225_b1 );
not ( \6226_b1 , w_15184 );
not ( \6226_b0 , w_15185 );
and ( w_15184 , w_15185 , \6225_b0 );
or ( \6227_b1 , \6221_b1 , \6226_b1 );
not ( \6226_b1 , w_15186 );
and ( \6227_b0 , \6221_b0 , w_15187 );
and ( w_15186 , w_15187 , \6226_b0 );
or ( \6228_b1 , \5737_b1 , \5768_b1 );
not ( \5768_b1 , w_15188 );
and ( \6228_b0 , \5737_b0 , w_15189 );
and ( w_15188 , w_15189 , \5768_b0 );
buf ( \6229_b1 , \6228_b1 );
not ( \6229_b1 , w_15190 );
not ( \6229_b0 , w_15191 );
and ( w_15190 , w_15191 , \6228_b0 );
or ( \6230_b1 , \6229_b1 , w_15192 );
xor ( \6230_b0 , \6229_b0 , w_15194 );
not ( w_15194 , w_15195 );
and ( w_15195 , w_15192 , w_15193 );
buf ( w_15192 , \5775_b1 );
not ( w_15192 , w_15196 );
not ( w_15193 , w_15197 );
and ( w_15196 , w_15197 , \5775_b0 );
or ( \6231_b1 , \6227_b1 , \6230_b1 );
xor ( \6231_b0 , \6227_b0 , w_15198 );
not ( w_15198 , w_15199 );
and ( w_15199 , \6230_b1 , \6230_b0 );
or ( \6232_b1 , \5758_b1 , \5790_b1 );
not ( \5790_b1 , w_15200 );
and ( \6232_b0 , \5758_b0 , w_15201 );
and ( w_15200 , w_15201 , \5790_b0 );
or ( \6233_b1 , \5770_b1 , \5788_b1 );
not ( \5788_b1 , w_15202 );
and ( \6233_b0 , \5770_b0 , w_15203 );
and ( w_15202 , w_15203 , \5788_b0 );
or ( \6234_b1 , \6232_b1 , w_15205 );
not ( w_15205 , w_15206 );
and ( \6234_b0 , \6232_b0 , w_15207 );
and ( w_15206 ,  , w_15207 );
buf ( w_15205 , \6233_b1 );
not ( w_15205 , w_15208 );
not (  , w_15209 );
and ( w_15208 , w_15209 , \6233_b0 );
or ( \6235_b1 , \6234_b1 , w_15210 );
xor ( \6235_b0 , \6234_b0 , w_15212 );
not ( w_15212 , w_15213 );
and ( w_15213 , w_15210 , w_15211 );
buf ( w_15210 , \5797_b1 );
not ( w_15210 , w_15214 );
not ( w_15211 , w_15215 );
and ( w_15214 , w_15215 , \5797_b0 );
or ( \6236_b1 , \6231_b1 , \6235_b1 );
xor ( \6236_b0 , \6231_b0 , w_15216 );
not ( w_15216 , w_15217 );
and ( w_15217 , \6235_b1 , \6235_b0 );
or ( \6237_b1 , \6165_b1 , \6236_b1 );
not ( \6236_b1 , w_15218 );
and ( \6237_b0 , \6165_b0 , w_15219 );
and ( w_15218 , w_15219 , \6236_b0 );
or ( \6238_b1 , \5906_b1 , \5935_b1 );
not ( \5935_b1 , w_15220 );
and ( \6238_b0 , \5906_b0 , w_15221 );
and ( w_15220 , w_15221 , \5935_b0 );
or ( \6239_b1 , \5918_b1 , \5933_b1 );
not ( \5933_b1 , w_15222 );
and ( \6239_b0 , \5918_b0 , w_15223 );
and ( w_15222 , w_15223 , \5933_b0 );
or ( \6240_b1 , \6238_b1 , w_15225 );
not ( w_15225 , w_15226 );
and ( \6240_b0 , \6238_b0 , w_15227 );
and ( w_15226 ,  , w_15227 );
buf ( w_15225 , \6239_b1 );
not ( w_15225 , w_15228 );
not (  , w_15229 );
and ( w_15228 , w_15229 , \6239_b0 );
or ( \6241_b1 , \6240_b1 , w_15230 );
xor ( \6241_b0 , \6240_b0 , w_15232 );
not ( w_15232 , w_15233 );
and ( w_15233 , w_15230 , w_15231 );
buf ( w_15230 , \5942_b1 );
not ( w_15230 , w_15234 );
not ( w_15231 , w_15235 );
and ( w_15234 , w_15235 , \5942_b0 );
or ( \6242_b1 , \5925_b1 , \5955_b1 );
not ( \5955_b1 , w_15236 );
and ( \6242_b0 , \5925_b0 , w_15237 );
and ( w_15236 , w_15237 , \5955_b0 );
or ( \6243_b1 , \5937_b1 , \5953_b1 );
not ( \5953_b1 , w_15238 );
and ( \6243_b0 , \5937_b0 , w_15239 );
and ( w_15238 , w_15239 , \5953_b0 );
or ( \6244_b1 , \6242_b1 , w_15241 );
not ( w_15241 , w_15242 );
and ( \6244_b0 , \6242_b0 , w_15243 );
and ( w_15242 ,  , w_15243 );
buf ( w_15241 , \6243_b1 );
not ( w_15241 , w_15244 );
not (  , w_15245 );
and ( w_15244 , w_15245 , \6243_b0 );
or ( \6245_b1 , \6244_b1 , w_15246 );
xor ( \6245_b0 , \6244_b0 , w_15248 );
not ( w_15248 , w_15249 );
and ( w_15249 , w_15246 , w_15247 );
buf ( w_15246 , \5962_b1 );
not ( w_15246 , w_15250 );
not ( w_15247 , w_15251 );
and ( w_15250 , w_15251 , \5962_b0 );
or ( \6246_b1 , \6241_b1 , \6245_b1 );
xor ( \6246_b0 , \6241_b0 , w_15252 );
not ( w_15252 , w_15253 );
and ( w_15253 , \6245_b1 , \6245_b0 );
or ( \6247_b1 , \5945_b1 , \5977_b1 );
not ( \5977_b1 , w_15254 );
and ( \6247_b0 , \5945_b0 , w_15255 );
and ( w_15254 , w_15255 , \5977_b0 );
or ( \6248_b1 , \5957_b1 , \5975_b1 );
not ( \5975_b1 , w_15256 );
and ( \6248_b0 , \5957_b0 , w_15257 );
and ( w_15256 , w_15257 , \5975_b0 );
or ( \6249_b1 , \6247_b1 , w_15259 );
not ( w_15259 , w_15260 );
and ( \6249_b0 , \6247_b0 , w_15261 );
and ( w_15260 ,  , w_15261 );
buf ( w_15259 , \6248_b1 );
not ( w_15259 , w_15262 );
not (  , w_15263 );
and ( w_15262 , w_15263 , \6248_b0 );
or ( \6250_b1 , \6249_b1 , w_15264 );
xor ( \6250_b0 , \6249_b0 , w_15266 );
not ( w_15266 , w_15267 );
and ( w_15267 , w_15264 , w_15265 );
buf ( w_15264 , \5984_b1 );
not ( w_15264 , w_15268 );
not ( w_15265 , w_15269 );
and ( w_15268 , w_15269 , \5984_b0 );
or ( \6251_b1 , \6246_b1 , \6250_b1 );
xor ( \6251_b0 , \6246_b0 , w_15270 );
not ( w_15270 , w_15271 );
and ( w_15271 , \6250_b1 , \6250_b0 );
or ( \6252_b1 , \5842_b1 , \5871_b1 );
not ( \5871_b1 , w_15272 );
and ( \6252_b0 , \5842_b0 , w_15273 );
and ( w_15272 , w_15273 , \5871_b0 );
or ( \6253_b1 , \5854_b1 , \5869_b1 );
not ( \5869_b1 , w_15274 );
and ( \6253_b0 , \5854_b0 , w_15275 );
and ( w_15274 , w_15275 , \5869_b0 );
or ( \6254_b1 , \6252_b1 , w_15277 );
not ( w_15277 , w_15278 );
and ( \6254_b0 , \6252_b0 , w_15279 );
and ( w_15278 ,  , w_15279 );
buf ( w_15277 , \6253_b1 );
not ( w_15277 , w_15280 );
not (  , w_15281 );
and ( w_15280 , w_15281 , \6253_b0 );
or ( \6255_b1 , \6254_b1 , w_15282 );
xor ( \6255_b0 , \6254_b0 , w_15284 );
not ( w_15284 , w_15285 );
and ( w_15285 , w_15282 , w_15283 );
buf ( w_15282 , \5878_b1 );
not ( w_15282 , w_15286 );
not ( w_15283 , w_15287 );
and ( w_15286 , w_15287 , \5878_b0 );
or ( \6256_b1 , \5861_b1 , \5891_b1 );
not ( \5891_b1 , w_15288 );
and ( \6256_b0 , \5861_b0 , w_15289 );
and ( w_15288 , w_15289 , \5891_b0 );
or ( \6257_b1 , \5873_b1 , \5889_b1 );
not ( \5889_b1 , w_15290 );
and ( \6257_b0 , \5873_b0 , w_15291 );
and ( w_15290 , w_15291 , \5889_b0 );
or ( \6258_b1 , \6256_b1 , w_15293 );
not ( w_15293 , w_15294 );
and ( \6258_b0 , \6256_b0 , w_15295 );
and ( w_15294 ,  , w_15295 );
buf ( w_15293 , \6257_b1 );
not ( w_15293 , w_15296 );
not (  , w_15297 );
and ( w_15296 , w_15297 , \6257_b0 );
or ( \6259_b1 , \6258_b1 , w_15298 );
xor ( \6259_b0 , \6258_b0 , w_15300 );
not ( w_15300 , w_15301 );
and ( w_15301 , w_15298 , w_15299 );
buf ( w_15298 , \5898_b1 );
not ( w_15298 , w_15302 );
not ( w_15299 , w_15303 );
and ( w_15302 , w_15303 , \5898_b0 );
or ( \6260_b1 , \6255_b1 , \6259_b1 );
xor ( \6260_b0 , \6255_b0 , w_15304 );
not ( w_15304 , w_15305 );
and ( w_15305 , \6259_b1 , \6259_b0 );
or ( \6261_b1 , \5881_b1 , \5916_b1 );
not ( \5916_b1 , w_15306 );
and ( \6261_b0 , \5881_b0 , w_15307 );
and ( w_15306 , w_15307 , \5916_b0 );
or ( \6262_b1 , \5893_b1 , \5914_b1 );
not ( \5914_b1 , w_15308 );
and ( \6262_b0 , \5893_b0 , w_15309 );
and ( w_15308 , w_15309 , \5914_b0 );
or ( \6263_b1 , \6261_b1 , w_15311 );
not ( w_15311 , w_15312 );
and ( \6263_b0 , \6261_b0 , w_15313 );
and ( w_15312 ,  , w_15313 );
buf ( w_15311 , \6262_b1 );
not ( w_15311 , w_15314 );
not (  , w_15315 );
and ( w_15314 , w_15315 , \6262_b0 );
or ( \6264_b1 , \6263_b1 , w_15316 );
xor ( \6264_b0 , \6263_b0 , w_15318 );
not ( w_15318 , w_15319 );
and ( w_15319 , w_15316 , w_15317 );
buf ( w_15316 , \5923_b1 );
not ( w_15316 , w_15320 );
not ( w_15317 , w_15321 );
and ( w_15320 , w_15321 , \5923_b0 );
or ( \6265_b1 , \6260_b1 , \6264_b1 );
xor ( \6265_b0 , \6260_b0 , w_15322 );
not ( w_15322 , w_15323 );
and ( w_15323 , \6264_b1 , \6264_b0 );
or ( \6266_b1 , \6251_b1 , \6265_b1 );
xor ( \6266_b0 , \6251_b0 , w_15324 );
not ( w_15324 , w_15325 );
and ( w_15325 , \6265_b1 , \6265_b0 );
or ( \6267_b1 , \5780_b1 , \5809_b1 );
not ( \5809_b1 , w_15326 );
and ( \6267_b0 , \5780_b0 , w_15327 );
and ( w_15326 , w_15327 , \5809_b0 );
or ( \6268_b1 , \5792_b1 , \5807_b1 );
not ( \5807_b1 , w_15328 );
and ( \6268_b0 , \5792_b0 , w_15329 );
and ( w_15328 , w_15329 , \5807_b0 );
or ( \6269_b1 , \6267_b1 , w_15331 );
not ( w_15331 , w_15332 );
and ( \6269_b0 , \6267_b0 , w_15333 );
and ( w_15332 ,  , w_15333 );
buf ( w_15331 , \6268_b1 );
not ( w_15331 , w_15334 );
not (  , w_15335 );
and ( w_15334 , w_15335 , \6268_b0 );
or ( \6270_b1 , \6269_b1 , w_15336 );
xor ( \6270_b0 , \6269_b0 , w_15338 );
not ( w_15338 , w_15339 );
and ( w_15339 , w_15336 , w_15337 );
buf ( w_15336 , \5816_b1 );
not ( w_15336 , w_15340 );
not ( w_15337 , w_15341 );
and ( w_15340 , w_15341 , \5816_b0 );
or ( \6271_b1 , \5799_b1 , \5829_b1 );
not ( \5829_b1 , w_15342 );
and ( \6271_b0 , \5799_b0 , w_15343 );
and ( w_15342 , w_15343 , \5829_b0 );
or ( \6272_b1 , \5811_b1 , \5827_b1 );
not ( \5827_b1 , w_15344 );
and ( \6272_b0 , \5811_b0 , w_15345 );
and ( w_15344 , w_15345 , \5827_b0 );
or ( \6273_b1 , \6271_b1 , w_15347 );
not ( w_15347 , w_15348 );
and ( \6273_b0 , \6271_b0 , w_15349 );
and ( w_15348 ,  , w_15349 );
buf ( w_15347 , \6272_b1 );
not ( w_15347 , w_15350 );
not (  , w_15351 );
and ( w_15350 , w_15351 , \6272_b0 );
or ( \6274_b1 , \6273_b1 , w_15352 );
xor ( \6274_b0 , \6273_b0 , w_15354 );
not ( w_15354 , w_15355 );
and ( w_15355 , w_15352 , w_15353 );
buf ( w_15352 , \5836_b1 );
not ( w_15352 , w_15356 );
not ( w_15353 , w_15357 );
and ( w_15356 , w_15357 , \5836_b0 );
or ( \6275_b1 , \6270_b1 , \6274_b1 );
xor ( \6275_b0 , \6270_b0 , w_15358 );
not ( w_15358 , w_15359 );
and ( w_15359 , \6274_b1 , \6274_b0 );
or ( \6276_b1 , \5819_b1 , \5852_b1 );
not ( \5852_b1 , w_15360 );
and ( \6276_b0 , \5819_b0 , w_15361 );
and ( w_15360 , w_15361 , \5852_b0 );
or ( \6277_b1 , \5831_b1 , \5850_b1 );
not ( \5850_b1 , w_15362 );
and ( \6277_b0 , \5831_b0 , w_15363 );
and ( w_15362 , w_15363 , \5850_b0 );
or ( \6278_b1 , \6276_b1 , w_15365 );
not ( w_15365 , w_15366 );
and ( \6278_b0 , \6276_b0 , w_15367 );
and ( w_15366 ,  , w_15367 );
buf ( w_15365 , \6277_b1 );
not ( w_15365 , w_15368 );
not (  , w_15369 );
and ( w_15368 , w_15369 , \6277_b0 );
or ( \6279_b1 , \6278_b1 , w_15370 );
xor ( \6279_b0 , \6278_b0 , w_15372 );
not ( w_15372 , w_15373 );
and ( w_15373 , w_15370 , w_15371 );
buf ( w_15370 , \5859_b1 );
not ( w_15370 , w_15374 );
not ( w_15371 , w_15375 );
and ( w_15374 , w_15375 , \5859_b0 );
or ( \6280_b1 , \6275_b1 , \6279_b1 );
xor ( \6280_b0 , \6275_b0 , w_15376 );
not ( w_15376 , w_15377 );
and ( w_15377 , \6279_b1 , \6279_b0 );
or ( \6281_b1 , \6266_b1 , \6280_b1 );
xor ( \6281_b0 , \6266_b0 , w_15378 );
not ( w_15378 , w_15379 );
and ( w_15379 , \6280_b1 , \6280_b0 );
or ( \6282_b1 , \6236_b1 , \6281_b1 );
not ( \6281_b1 , w_15380 );
and ( \6282_b0 , \6236_b0 , w_15381 );
and ( w_15380 , w_15381 , \6281_b0 );
or ( \6283_b1 , \6165_b1 , \6281_b1 );
not ( \6281_b1 , w_15382 );
and ( \6283_b0 , \6165_b0 , w_15383 );
and ( w_15382 , w_15383 , \6281_b0 );
or ( \6285_b1 , \6122_b1 , \6284_b1 );
not ( \6284_b1 , w_15384 );
and ( \6285_b0 , \6122_b0 , w_15385 );
and ( w_15384 , w_15385 , \6284_b0 );
or ( \6286_b1 , \6029_b1 , \6055_b1 );
not ( \6055_b1 , w_15386 );
and ( \6286_b0 , \6029_b0 , w_15387 );
and ( w_15386 , w_15387 , \6055_b0 );
or ( \6287_b1 , \6041_b1 , \6053_b1 );
not ( \6053_b1 , w_15388 );
and ( \6287_b0 , \6041_b0 , w_15389 );
and ( w_15388 , w_15389 , \6053_b0 );
or ( \6288_b1 , \6286_b1 , w_15391 );
not ( w_15391 , w_15392 );
and ( \6288_b0 , \6286_b0 , w_15393 );
and ( w_15392 ,  , w_15393 );
buf ( w_15391 , \6287_b1 );
not ( w_15391 , w_15394 );
not (  , w_15395 );
and ( w_15394 , w_15395 , \6287_b0 );
or ( \6289_b1 , \6288_b1 , w_15396 );
xor ( \6289_b0 , \6288_b0 , w_15398 );
not ( w_15398 , w_15399 );
and ( w_15399 , w_15396 , w_15397 );
buf ( w_15396 , \6062_b1 );
not ( w_15396 , w_15400 );
not ( w_15397 , w_15401 );
and ( w_15400 , w_15401 , \6062_b0 );
or ( \6290_b1 , \6048_b1 , \6082_b1 );
not ( \6082_b1 , w_15402 );
and ( \6290_b0 , \6048_b0 , w_15403 );
and ( w_15402 , w_15403 , \6082_b0 );
or ( \6291_b1 , \6057_b1 , \6066_b1 );
not ( \6066_b1 , w_15404 );
and ( \6291_b0 , \6057_b0 , w_15405 );
and ( w_15404 , w_15405 , \6066_b0 );
or ( \6292_b1 , \6290_b1 , w_15407 );
not ( w_15407 , w_15408 );
and ( \6292_b0 , \6290_b0 , w_15409 );
and ( w_15408 ,  , w_15409 );
buf ( w_15407 , \6291_b1 );
not ( w_15407 , w_15410 );
not (  , w_15411 );
and ( w_15410 , w_15411 , \6291_b0 );
or ( \6293_b1 , \6292_b1 , w_15412 );
xor ( \6293_b0 , \6292_b0 , w_15414 );
not ( w_15414 , w_15415 );
and ( w_15415 , w_15412 , w_15413 );
buf ( w_15412 , \5736_b1 );
not ( w_15412 , w_15416 );
not ( w_15413 , w_15417 );
and ( w_15416 , w_15417 , \5736_b0 );
or ( \6294_b1 , \6289_b1 , \6293_b1 );
xor ( \6294_b0 , \6289_b0 , w_15418 );
not ( w_15418 , w_15419 );
and ( w_15419 , \6293_b1 , \6293_b0 );
or ( \6295_b1 , \6224_b1 , \5727_b1 );
xor ( \6295_b0 , \6224_b0 , w_15420 );
not ( w_15420 , w_15421 );
and ( w_15421 , \5727_b1 , \5727_b0 );
or ( \6296_b1 , \6065_b1 , w_15423 );
not ( w_15423 , w_15424 );
and ( \6296_b0 , \6065_b0 , w_15425 );
and ( w_15424 ,  , w_15425 );
buf ( w_15423 , \6295_b1 );
not ( w_15423 , w_15426 );
not (  , w_15427 );
and ( w_15426 , w_15427 , \6295_b0 );
or ( \6297_b1 , \6296_b1 , w_15428 );
xor ( \6297_b0 , \6296_b0 , w_15430 );
not ( w_15430 , w_15431 );
and ( w_15431 , w_15428 , w_15429 );
buf ( w_15428 , \6227_b1 );
not ( w_15428 , w_15432 );
not ( w_15429 , w_15433 );
and ( w_15432 , w_15433 , \6227_b0 );
or ( \6298_b1 , \6294_b1 , \6297_b1 );
xor ( \6298_b0 , \6294_b0 , w_15434 );
not ( w_15434 , w_15435 );
and ( w_15435 , \6297_b1 , \6297_b0 );
or ( \6299_b1 , \5967_b1 , \5996_b1 );
not ( \5996_b1 , w_15436 );
and ( \6299_b0 , \5967_b0 , w_15437 );
and ( w_15436 , w_15437 , \5996_b0 );
or ( \6300_b1 , \5979_b1 , \5994_b1 );
not ( \5994_b1 , w_15438 );
and ( \6300_b0 , \5979_b0 , w_15439 );
and ( w_15438 , w_15439 , \5994_b0 );
or ( \6301_b1 , \6299_b1 , w_15441 );
not ( w_15441 , w_15442 );
and ( \6301_b0 , \6299_b0 , w_15443 );
and ( w_15442 ,  , w_15443 );
buf ( w_15441 , \6300_b1 );
not ( w_15441 , w_15444 );
not (  , w_15445 );
and ( w_15444 , w_15445 , \6300_b0 );
or ( \6302_b1 , \6301_b1 , w_15446 );
xor ( \6302_b0 , \6301_b0 , w_15448 );
not ( w_15448 , w_15449 );
and ( w_15449 , w_15446 , w_15447 );
buf ( w_15446 , \6003_b1 );
not ( w_15446 , w_15450 );
not ( w_15447 , w_15451 );
and ( w_15450 , w_15451 , \6003_b0 );
or ( \6303_b1 , \5986_b1 , \6016_b1 );
not ( \6016_b1 , w_15452 );
and ( \6303_b0 , \5986_b0 , w_15453 );
and ( w_15452 , w_15453 , \6016_b0 );
or ( \6304_b1 , \5998_b1 , \6014_b1 );
not ( \6014_b1 , w_15454 );
and ( \6304_b0 , \5998_b0 , w_15455 );
and ( w_15454 , w_15455 , \6014_b0 );
or ( \6305_b1 , \6303_b1 , w_15457 );
not ( w_15457 , w_15458 );
and ( \6305_b0 , \6303_b0 , w_15459 );
and ( w_15458 ,  , w_15459 );
buf ( w_15457 , \6304_b1 );
not ( w_15457 , w_15460 );
not (  , w_15461 );
and ( w_15460 , w_15461 , \6304_b0 );
or ( \6306_b1 , \6305_b1 , w_15462 );
xor ( \6306_b0 , \6305_b0 , w_15464 );
not ( w_15464 , w_15465 );
and ( w_15465 , w_15462 , w_15463 );
buf ( w_15462 , \6023_b1 );
not ( w_15462 , w_15466 );
not ( w_15463 , w_15467 );
and ( w_15466 , w_15467 , \6023_b0 );
or ( \6307_b1 , \6302_b1 , \6306_b1 );
xor ( \6307_b0 , \6302_b0 , w_15468 );
not ( w_15468 , w_15469 );
and ( w_15469 , \6306_b1 , \6306_b0 );
or ( \6308_b1 , \6006_b1 , \6039_b1 );
not ( \6039_b1 , w_15470 );
and ( \6308_b0 , \6006_b0 , w_15471 );
and ( w_15470 , w_15471 , \6039_b0 );
or ( \6309_b1 , \6018_b1 , \6037_b1 );
not ( \6037_b1 , w_15472 );
and ( \6309_b0 , \6018_b0 , w_15473 );
and ( w_15472 , w_15473 , \6037_b0 );
or ( \6310_b1 , \6308_b1 , w_15475 );
not ( w_15475 , w_15476 );
and ( \6310_b0 , \6308_b0 , w_15477 );
and ( w_15476 ,  , w_15477 );
buf ( w_15475 , \6309_b1 );
not ( w_15475 , w_15478 );
not (  , w_15479 );
and ( w_15478 , w_15479 , \6309_b0 );
or ( \6311_b1 , \6310_b1 , w_15480 );
xor ( \6311_b0 , \6310_b0 , w_15482 );
not ( w_15482 , w_15483 );
and ( w_15483 , w_15480 , w_15481 );
buf ( w_15480 , \6046_b1 );
not ( w_15480 , w_15484 );
not ( w_15481 , w_15485 );
and ( w_15484 , w_15485 , \6046_b0 );
or ( \6312_b1 , \6307_b1 , \6311_b1 );
xor ( \6312_b0 , \6307_b0 , w_15486 );
not ( w_15486 , w_15487 );
and ( w_15487 , \6311_b1 , \6311_b0 );
or ( \6313_b1 , \6298_b1 , w_15488 );
xor ( \6313_b0 , \6298_b0 , w_15490 );
not ( w_15490 , w_15491 );
and ( w_15491 , w_15488 , w_15489 );
buf ( w_15488 , \6312_b1 );
not ( w_15488 , w_15492 );
not ( w_15489 , w_15493 );
and ( w_15492 , w_15493 , \6312_b0 );
or ( \6314_b1 , \6106_b1 , \6110_b1 );
not ( \6110_b1 , w_15494 );
and ( \6314_b0 , \6106_b0 , w_15495 );
and ( w_15494 , w_15495 , \6110_b0 );
or ( \6315_b1 , \6110_b1 , \6115_b1 );
not ( \6115_b1 , w_15496 );
and ( \6315_b0 , \6110_b0 , w_15497 );
and ( w_15496 , w_15497 , \6115_b0 );
or ( \6316_b1 , \6106_b1 , \6115_b1 );
not ( \6115_b1 , w_15498 );
and ( \6316_b0 , \6106_b0 , w_15499 );
and ( w_15498 , w_15499 , \6115_b0 );
or ( \6318_b1 , \6091_b1 , \6095_b1 );
not ( \6095_b1 , w_15500 );
and ( \6318_b0 , \6091_b0 , w_15501 );
and ( w_15500 , w_15501 , \6095_b0 );
or ( \6319_b1 , \6095_b1 , \6100_b1 );
not ( \6100_b1 , w_15502 );
and ( \6319_b0 , \6095_b0 , w_15503 );
and ( w_15502 , w_15503 , \6100_b0 );
or ( \6320_b1 , \6091_b1 , \6100_b1 );
not ( \6100_b1 , w_15504 );
and ( \6320_b0 , \6091_b0 , w_15505 );
and ( w_15504 , w_15505 , \6100_b0 );
or ( \6322_b1 , \6317_b1 , \6321_b1 );
xor ( \6322_b0 , \6317_b0 , w_15506 );
not ( w_15506 , w_15507 );
and ( w_15507 , \6321_b1 , \6321_b0 );
or ( \6323_b1 , \6079_b1 , \6086_b1 );
not ( \6086_b1 , w_15508 );
and ( \6323_b0 , \6079_b0 , w_15509 );
and ( w_15508 , w_15509 , \6086_b0 );
or ( \6324_b1 , \6322_b1 , \6323_b1 );
xor ( \6324_b0 , \6322_b0 , w_15510 );
not ( w_15510 , w_15511 );
and ( w_15511 , \6323_b1 , \6323_b0 );
or ( \6325_b1 , \6313_b1 , \6324_b1 );
not ( \6324_b1 , w_15512 );
and ( \6325_b0 , \6313_b0 , w_15513 );
and ( w_15512 , w_15513 , \6324_b0 );
or ( \6326_b1 , \6152_b1 , \6156_b1 );
not ( \6156_b1 , w_15514 );
and ( \6326_b0 , \6152_b0 , w_15515 );
and ( w_15514 , w_15515 , \6156_b0 );
or ( \6327_b1 , \6156_b1 , \6161_b1 );
not ( \6161_b1 , w_15516 );
and ( \6327_b0 , \6156_b0 , w_15517 );
and ( w_15516 , w_15517 , \6161_b0 );
or ( \6328_b1 , \6152_b1 , \6161_b1 );
not ( \6161_b1 , w_15518 );
and ( \6328_b0 , \6152_b0 , w_15519 );
and ( w_15518 , w_15519 , \6161_b0 );
or ( \6330_b1 , \6140_b1 , \6144_b1 );
not ( \6144_b1 , w_15520 );
and ( \6330_b0 , \6140_b0 , w_15521 );
and ( w_15520 , w_15521 , \6144_b0 );
or ( \6331_b1 , \6144_b1 , \6149_b1 );
not ( \6149_b1 , w_15522 );
and ( \6331_b0 , \6144_b0 , w_15523 );
and ( w_15522 , w_15523 , \6149_b0 );
or ( \6332_b1 , \6140_b1 , \6149_b1 );
not ( \6149_b1 , w_15524 );
and ( \6332_b0 , \6140_b0 , w_15525 );
and ( w_15524 , w_15525 , \6149_b0 );
or ( \6334_b1 , \6329_b1 , \6333_b1 );
xor ( \6334_b0 , \6329_b0 , w_15526 );
not ( w_15526 , w_15527 );
and ( w_15527 , \6333_b1 , \6333_b0 );
or ( \6335_b1 , \6126_b1 , \6130_b1 );
not ( \6130_b1 , w_15528 );
and ( \6335_b0 , \6126_b0 , w_15529 );
and ( w_15528 , w_15529 , \6130_b0 );
or ( \6336_b1 , \6130_b1 , \6135_b1 );
not ( \6135_b1 , w_15530 );
and ( \6336_b0 , \6130_b0 , w_15531 );
and ( w_15530 , w_15531 , \6135_b0 );
or ( \6337_b1 , \6126_b1 , \6135_b1 );
not ( \6135_b1 , w_15532 );
and ( \6337_b0 , \6126_b0 , w_15533 );
and ( w_15532 , w_15533 , \6135_b0 );
or ( \6339_b1 , \6334_b1 , \6338_b1 );
xor ( \6339_b0 , \6334_b0 , w_15534 );
not ( w_15534 , w_15535 );
and ( w_15535 , \6338_b1 , \6338_b0 );
or ( \6340_b1 , \6324_b1 , \6339_b1 );
not ( \6339_b1 , w_15536 );
and ( \6340_b0 , \6324_b0 , w_15537 );
and ( w_15536 , w_15537 , \6339_b0 );
or ( \6341_b1 , \6313_b1 , \6339_b1 );
not ( \6339_b1 , w_15538 );
and ( \6341_b0 , \6313_b0 , w_15539 );
and ( w_15538 , w_15539 , \6339_b0 );
or ( \6343_b1 , \6284_b1 , \6342_b1 );
not ( \6342_b1 , w_15540 );
and ( \6343_b0 , \6284_b0 , w_15541 );
and ( w_15540 , w_15541 , \6342_b0 );
or ( \6344_b1 , \6122_b1 , \6342_b1 );
not ( \6342_b1 , w_15542 );
and ( \6344_b0 , \6122_b0 , w_15543 );
and ( w_15542 , w_15543 , \6342_b0 );
or ( \6346_b1 , \6241_b1 , \6245_b1 );
not ( \6245_b1 , w_15544 );
and ( \6346_b0 , \6241_b0 , w_15545 );
and ( w_15544 , w_15545 , \6245_b0 );
or ( \6347_b1 , \6245_b1 , \6250_b1 );
not ( \6250_b1 , w_15546 );
and ( \6347_b0 , \6245_b0 , w_15547 );
and ( w_15546 , w_15547 , \6250_b0 );
or ( \6348_b1 , \6241_b1 , \6250_b1 );
not ( \6250_b1 , w_15548 );
and ( \6348_b0 , \6241_b0 , w_15549 );
and ( w_15548 , w_15549 , \6250_b0 );
or ( \6350_b1 , \6302_b1 , \6306_b1 );
not ( \6306_b1 , w_15550 );
and ( \6350_b0 , \6302_b0 , w_15551 );
and ( w_15550 , w_15551 , \6306_b0 );
or ( \6351_b1 , \6306_b1 , \6311_b1 );
not ( \6311_b1 , w_15552 );
and ( \6351_b0 , \6306_b0 , w_15553 );
and ( w_15552 , w_15553 , \6311_b0 );
or ( \6352_b1 , \6302_b1 , \6311_b1 );
not ( \6311_b1 , w_15554 );
and ( \6352_b0 , \6302_b0 , w_15555 );
and ( w_15554 , w_15555 , \6311_b0 );
or ( \6354_b1 , \6349_b1 , \6353_b1 );
xor ( \6354_b0 , \6349_b0 , w_15556 );
not ( w_15556 , w_15557 );
and ( w_15557 , \6353_b1 , \6353_b0 );
or ( \6355_b1 , \6289_b1 , \6293_b1 );
not ( \6293_b1 , w_15558 );
and ( \6355_b0 , \6289_b0 , w_15559 );
and ( w_15558 , w_15559 , \6293_b0 );
or ( \6356_b1 , \6293_b1 , \6297_b1 );
not ( \6297_b1 , w_15560 );
and ( \6356_b0 , \6293_b0 , w_15561 );
and ( w_15560 , w_15561 , \6297_b0 );
or ( \6357_b1 , \6289_b1 , \6297_b1 );
not ( \6297_b1 , w_15562 );
and ( \6357_b0 , \6289_b0 , w_15563 );
and ( w_15562 , w_15563 , \6297_b0 );
or ( \6359_b1 , \6354_b1 , \6358_b1 );
xor ( \6359_b0 , \6354_b0 , w_15564 );
not ( w_15564 , w_15565 );
and ( w_15565 , \6358_b1 , \6358_b0 );
or ( \6360_b1 , \6227_b1 , \6230_b1 );
not ( \6230_b1 , w_15566 );
and ( \6360_b0 , \6227_b0 , w_15567 );
and ( w_15566 , w_15567 , \6230_b0 );
or ( \6361_b1 , \6230_b1 , \6235_b1 );
not ( \6235_b1 , w_15568 );
and ( \6361_b0 , \6230_b0 , w_15569 );
and ( w_15568 , w_15569 , \6235_b0 );
or ( \6362_b1 , \6227_b1 , \6235_b1 );
not ( \6235_b1 , w_15570 );
and ( \6362_b0 , \6227_b0 , w_15571 );
and ( w_15570 , w_15571 , \6235_b0 );
or ( \6364_b1 , \6270_b1 , \6274_b1 );
not ( \6274_b1 , w_15572 );
and ( \6364_b0 , \6270_b0 , w_15573 );
and ( w_15572 , w_15573 , \6274_b0 );
or ( \6365_b1 , \6274_b1 , \6279_b1 );
not ( \6279_b1 , w_15574 );
and ( \6365_b0 , \6274_b0 , w_15575 );
and ( w_15574 , w_15575 , \6279_b0 );
or ( \6366_b1 , \6270_b1 , \6279_b1 );
not ( \6279_b1 , w_15576 );
and ( \6366_b0 , \6270_b0 , w_15577 );
and ( w_15576 , w_15577 , \6279_b0 );
or ( \6368_b1 , \6363_b1 , \6367_b1 );
xor ( \6368_b0 , \6363_b0 , w_15578 );
not ( w_15578 , w_15579 );
and ( w_15579 , \6367_b1 , \6367_b0 );
or ( \6369_b1 , \6255_b1 , \6259_b1 );
not ( \6259_b1 , w_15580 );
and ( \6369_b0 , \6255_b0 , w_15581 );
and ( w_15580 , w_15581 , \6259_b0 );
or ( \6370_b1 , \6259_b1 , \6264_b1 );
not ( \6264_b1 , w_15582 );
and ( \6370_b0 , \6259_b0 , w_15583 );
and ( w_15582 , w_15583 , \6264_b0 );
or ( \6371_b1 , \6255_b1 , \6264_b1 );
not ( \6264_b1 , w_15584 );
and ( \6371_b0 , \6255_b0 , w_15585 );
and ( w_15584 , w_15585 , \6264_b0 );
or ( \6373_b1 , \6368_b1 , \6372_b1 );
xor ( \6373_b0 , \6368_b0 , w_15586 );
not ( w_15586 , w_15587 );
and ( w_15587 , \6372_b1 , \6372_b0 );
or ( \6374_b1 , \6359_b1 , \6373_b1 );
xor ( \6374_b0 , \6359_b0 , w_15588 );
not ( w_15588 , w_15589 );
and ( w_15589 , \6373_b1 , \6373_b0 );
or ( \6375_b1 , \6251_b1 , \6265_b1 );
not ( \6265_b1 , w_15590 );
and ( \6375_b0 , \6251_b0 , w_15591 );
and ( w_15590 , w_15591 , \6265_b0 );
or ( \6376_b1 , \6265_b1 , \6280_b1 );
not ( \6280_b1 , w_15592 );
and ( \6376_b0 , \6265_b0 , w_15593 );
and ( w_15592 , w_15593 , \6280_b0 );
or ( \6377_b1 , \6251_b1 , \6280_b1 );
not ( \6280_b1 , w_15594 );
and ( \6377_b0 , \6251_b0 , w_15595 );
and ( w_15594 , w_15595 , \6280_b0 );
or ( \6379_b1 , \5873_b1 , \5891_b1 );
not ( \5891_b1 , w_15596 );
and ( \6379_b0 , \5873_b0 , w_15597 );
and ( w_15596 , w_15597 , \5891_b0 );
or ( \6380_b1 , \5842_b1 , \5889_b1 );
not ( \5889_b1 , w_15598 );
and ( \6380_b0 , \5842_b0 , w_15599 );
and ( w_15598 , w_15599 , \5889_b0 );
or ( \6381_b1 , \6379_b1 , w_15601 );
not ( w_15601 , w_15602 );
and ( \6381_b0 , \6379_b0 , w_15603 );
and ( w_15602 ,  , w_15603 );
buf ( w_15601 , \6380_b1 );
not ( w_15601 , w_15604 );
not (  , w_15605 );
and ( w_15604 , w_15605 , \6380_b0 );
or ( \6382_b1 , \6381_b1 , w_15606 );
xor ( \6382_b0 , \6381_b0 , w_15608 );
not ( w_15608 , w_15609 );
and ( w_15609 , w_15606 , w_15607 );
buf ( w_15606 , \5898_b1 );
not ( w_15606 , w_15610 );
not ( w_15607 , w_15611 );
and ( w_15610 , w_15611 , \5898_b0 );
or ( \6383_b1 , \5893_b1 , \5916_b1 );
not ( \5916_b1 , w_15612 );
and ( \6383_b0 , \5893_b0 , w_15613 );
and ( w_15612 , w_15613 , \5916_b0 );
or ( \6384_b1 , \5861_b1 , \5914_b1 );
not ( \5914_b1 , w_15614 );
and ( \6384_b0 , \5861_b0 , w_15615 );
and ( w_15614 , w_15615 , \5914_b0 );
or ( \6385_b1 , \6383_b1 , w_15617 );
not ( w_15617 , w_15618 );
and ( \6385_b0 , \6383_b0 , w_15619 );
and ( w_15618 ,  , w_15619 );
buf ( w_15617 , \6384_b1 );
not ( w_15617 , w_15620 );
not (  , w_15621 );
and ( w_15620 , w_15621 , \6384_b0 );
or ( \6386_b1 , \6385_b1 , w_15622 );
xor ( \6386_b0 , \6385_b0 , w_15624 );
not ( w_15624 , w_15625 );
and ( w_15625 , w_15622 , w_15623 );
buf ( w_15622 , \5923_b1 );
not ( w_15622 , w_15626 );
not ( w_15623 , w_15627 );
and ( w_15626 , w_15627 , \5923_b0 );
or ( \6387_b1 , \6382_b1 , \6386_b1 );
xor ( \6387_b0 , \6382_b0 , w_15628 );
not ( w_15628 , w_15629 );
and ( w_15629 , \6386_b1 , \6386_b0 );
or ( \6388_b1 , \5918_b1 , \5935_b1 );
not ( \5935_b1 , w_15630 );
and ( \6388_b0 , \5918_b0 , w_15631 );
and ( w_15630 , w_15631 , \5935_b0 );
or ( \6389_b1 , \5881_b1 , \5933_b1 );
not ( \5933_b1 , w_15632 );
and ( \6389_b0 , \5881_b0 , w_15633 );
and ( w_15632 , w_15633 , \5933_b0 );
or ( \6390_b1 , \6388_b1 , w_15635 );
not ( w_15635 , w_15636 );
and ( \6390_b0 , \6388_b0 , w_15637 );
and ( w_15636 ,  , w_15637 );
buf ( w_15635 , \6389_b1 );
not ( w_15635 , w_15638 );
not (  , w_15639 );
and ( w_15638 , w_15639 , \6389_b0 );
or ( \6391_b1 , \6390_b1 , w_15640 );
xor ( \6391_b0 , \6390_b0 , w_15642 );
not ( w_15642 , w_15643 );
and ( w_15643 , w_15640 , w_15641 );
buf ( w_15640 , \5942_b1 );
not ( w_15640 , w_15644 );
not ( w_15641 , w_15645 );
and ( w_15644 , w_15645 , \5942_b0 );
or ( \6392_b1 , \6387_b1 , \6391_b1 );
xor ( \6392_b0 , \6387_b0 , w_15646 );
not ( w_15646 , w_15647 );
and ( w_15647 , \6391_b1 , \6391_b0 );
or ( \6393_b1 , \5811_b1 , \5829_b1 );
not ( \5829_b1 , w_15648 );
and ( \6393_b0 , \5811_b0 , w_15649 );
and ( w_15648 , w_15649 , \5829_b0 );
or ( \6394_b1 , \5780_b1 , \5827_b1 );
not ( \5827_b1 , w_15650 );
and ( \6394_b0 , \5780_b0 , w_15651 );
and ( w_15650 , w_15651 , \5827_b0 );
or ( \6395_b1 , \6393_b1 , w_15653 );
not ( w_15653 , w_15654 );
and ( \6395_b0 , \6393_b0 , w_15655 );
and ( w_15654 ,  , w_15655 );
buf ( w_15653 , \6394_b1 );
not ( w_15653 , w_15656 );
not (  , w_15657 );
and ( w_15656 , w_15657 , \6394_b0 );
or ( \6396_b1 , \6395_b1 , w_15658 );
xor ( \6396_b0 , \6395_b0 , w_15660 );
not ( w_15660 , w_15661 );
and ( w_15661 , w_15658 , w_15659 );
buf ( w_15658 , \5836_b1 );
not ( w_15658 , w_15662 );
not ( w_15659 , w_15663 );
and ( w_15662 , w_15663 , \5836_b0 );
or ( \6397_b1 , \5831_b1 , \5852_b1 );
not ( \5852_b1 , w_15664 );
and ( \6397_b0 , \5831_b0 , w_15665 );
and ( w_15664 , w_15665 , \5852_b0 );
or ( \6398_b1 , \5799_b1 , \5850_b1 );
not ( \5850_b1 , w_15666 );
and ( \6398_b0 , \5799_b0 , w_15667 );
and ( w_15666 , w_15667 , \5850_b0 );
or ( \6399_b1 , \6397_b1 , w_15669 );
not ( w_15669 , w_15670 );
and ( \6399_b0 , \6397_b0 , w_15671 );
and ( w_15670 ,  , w_15671 );
buf ( w_15669 , \6398_b1 );
not ( w_15669 , w_15672 );
not (  , w_15673 );
and ( w_15672 , w_15673 , \6398_b0 );
or ( \6400_b1 , \6399_b1 , w_15674 );
xor ( \6400_b0 , \6399_b0 , w_15676 );
not ( w_15676 , w_15677 );
and ( w_15677 , w_15674 , w_15675 );
buf ( w_15674 , \5859_b1 );
not ( w_15674 , w_15678 );
not ( w_15675 , w_15679 );
and ( w_15678 , w_15679 , \5859_b0 );
or ( \6401_b1 , \6396_b1 , \6400_b1 );
xor ( \6401_b0 , \6396_b0 , w_15680 );
not ( w_15680 , w_15681 );
and ( w_15681 , \6400_b1 , \6400_b0 );
or ( \6402_b1 , \5854_b1 , \5871_b1 );
not ( \5871_b1 , w_15682 );
and ( \6402_b0 , \5854_b0 , w_15683 );
and ( w_15682 , w_15683 , \5871_b0 );
or ( \6403_b1 , \5819_b1 , \5869_b1 );
not ( \5869_b1 , w_15684 );
and ( \6403_b0 , \5819_b0 , w_15685 );
and ( w_15684 , w_15685 , \5869_b0 );
or ( \6404_b1 , \6402_b1 , w_15687 );
not ( w_15687 , w_15688 );
and ( \6404_b0 , \6402_b0 , w_15689 );
and ( w_15688 ,  , w_15689 );
buf ( w_15687 , \6403_b1 );
not ( w_15687 , w_15690 );
not (  , w_15691 );
and ( w_15690 , w_15691 , \6403_b0 );
or ( \6405_b1 , \6404_b1 , w_15692 );
xor ( \6405_b0 , \6404_b0 , w_15694 );
not ( w_15694 , w_15695 );
and ( w_15695 , w_15692 , w_15693 );
buf ( w_15692 , \5878_b1 );
not ( w_15692 , w_15696 );
not ( w_15693 , w_15697 );
and ( w_15696 , w_15697 , \5878_b0 );
or ( \6406_b1 , \6401_b1 , \6405_b1 );
xor ( \6406_b0 , \6401_b0 , w_15698 );
not ( w_15698 , w_15699 );
and ( w_15699 , \6405_b1 , \6405_b0 );
or ( \6407_b1 , \6392_b1 , \6406_b1 );
xor ( \6407_b0 , \6392_b0 , w_15700 );
not ( w_15700 , w_15701 );
and ( w_15701 , \6406_b1 , \6406_b0 );
buf ( \6408_b1 , \5775_b1 );
not ( \6408_b1 , w_15702 );
not ( \6408_b0 , w_15703 );
and ( w_15702 , w_15703 , \5775_b0 );
or ( \6409_b1 , \5770_b1 , \5790_b1 );
not ( \5790_b1 , w_15704 );
and ( \6409_b0 , \5770_b0 , w_15705 );
and ( w_15704 , w_15705 , \5790_b0 );
or ( \6410_b1 , \5737_b1 , \5788_b1 );
not ( \5788_b1 , w_15706 );
and ( \6410_b0 , \5737_b0 , w_15707 );
and ( w_15706 , w_15707 , \5788_b0 );
or ( \6411_b1 , \6409_b1 , w_15709 );
not ( w_15709 , w_15710 );
and ( \6411_b0 , \6409_b0 , w_15711 );
and ( w_15710 ,  , w_15711 );
buf ( w_15709 , \6410_b1 );
not ( w_15709 , w_15712 );
not (  , w_15713 );
and ( w_15712 , w_15713 , \6410_b0 );
or ( \6412_b1 , \6411_b1 , w_15714 );
xor ( \6412_b0 , \6411_b0 , w_15716 );
not ( w_15716 , w_15717 );
and ( w_15717 , w_15714 , w_15715 );
buf ( w_15714 , \5797_b1 );
not ( w_15714 , w_15718 );
not ( w_15715 , w_15719 );
and ( w_15718 , w_15719 , \5797_b0 );
or ( \6413_b1 , \6408_b1 , \6412_b1 );
xor ( \6413_b0 , \6408_b0 , w_15720 );
not ( w_15720 , w_15721 );
and ( w_15721 , \6412_b1 , \6412_b0 );
or ( \6414_b1 , \5792_b1 , \5809_b1 );
not ( \5809_b1 , w_15722 );
and ( \6414_b0 , \5792_b0 , w_15723 );
and ( w_15722 , w_15723 , \5809_b0 );
or ( \6415_b1 , \5758_b1 , \5807_b1 );
not ( \5807_b1 , w_15724 );
and ( \6415_b0 , \5758_b0 , w_15725 );
and ( w_15724 , w_15725 , \5807_b0 );
or ( \6416_b1 , \6414_b1 , w_15727 );
not ( w_15727 , w_15728 );
and ( \6416_b0 , \6414_b0 , w_15729 );
and ( w_15728 ,  , w_15729 );
buf ( w_15727 , \6415_b1 );
not ( w_15727 , w_15730 );
not (  , w_15731 );
and ( w_15730 , w_15731 , \6415_b0 );
or ( \6417_b1 , \6416_b1 , w_15732 );
xor ( \6417_b0 , \6416_b0 , w_15734 );
not ( w_15734 , w_15735 );
and ( w_15735 , w_15732 , w_15733 );
buf ( w_15732 , \5816_b1 );
not ( w_15732 , w_15736 );
not ( w_15733 , w_15737 );
and ( w_15736 , w_15737 , \5816_b0 );
or ( \6418_b1 , \6413_b1 , \6417_b1 );
xor ( \6418_b0 , \6413_b0 , w_15738 );
not ( w_15738 , w_15739 );
and ( w_15739 , \6417_b1 , \6417_b0 );
or ( \6419_b1 , \6407_b1 , \6418_b1 );
xor ( \6419_b0 , \6407_b0 , w_15740 );
not ( w_15740 , w_15741 );
and ( w_15741 , \6418_b1 , \6418_b0 );
or ( \6420_b1 , \6378_b1 , \6419_b1 );
xor ( \6420_b0 , \6378_b0 , w_15742 );
not ( w_15742 , w_15743 );
and ( w_15743 , \6419_b1 , \6419_b0 );
or ( \6421_b1 , \6057_b1 , \6082_b1 );
not ( \6082_b1 , w_15744 );
and ( \6421_b0 , \6057_b0 , w_15745 );
and ( w_15744 , w_15745 , \6082_b0 );
or ( \6422_b1 , \6029_b1 , \6066_b1 );
not ( \6066_b1 , w_15746 );
and ( \6422_b0 , \6029_b0 , w_15747 );
and ( w_15746 , w_15747 , \6066_b0 );
or ( \6423_b1 , \6421_b1 , w_15749 );
not ( w_15749 , w_15750 );
and ( \6423_b0 , \6421_b0 , w_15751 );
and ( w_15750 ,  , w_15751 );
buf ( w_15749 , \6422_b1 );
not ( w_15749 , w_15752 );
not (  , w_15753 );
and ( w_15752 , w_15753 , \6422_b0 );
or ( \6424_b1 , \6423_b1 , w_15754 );
xor ( \6424_b0 , \6423_b0 , w_15756 );
not ( w_15756 , w_15757 );
and ( w_15757 , w_15754 , w_15755 );
buf ( w_15754 , \5736_b1 );
not ( w_15754 , w_15758 );
not ( w_15755 , w_15759 );
and ( w_15758 , w_15759 , \5736_b0 );
or ( \6425_b1 , \6221_b1 , \6224_b1 );
xor ( \6425_b0 , \6221_b0 , w_15760 );
not ( w_15760 , w_15761 );
and ( w_15761 , \6224_b1 , \6224_b0 );
buf ( \6426_b1 , \6295_b1 );
not ( \6426_b1 , w_15762 );
not ( \6426_b0 , w_15763 );
and ( w_15762 , w_15763 , \6295_b0 );
or ( \6427_b1 , \6425_b1 , \6426_b1 );
not ( \6426_b1 , w_15764 );
and ( \6427_b0 , \6425_b0 , w_15765 );
and ( w_15764 , w_15765 , \6426_b0 );
or ( \6428_b1 , \6065_b1 , \6427_b1 );
not ( \6427_b1 , w_15766 );
and ( \6428_b0 , \6065_b0 , w_15767 );
and ( w_15766 , w_15767 , \6427_b0 );
or ( \6429_b1 , \6048_b1 , \6295_b1 );
not ( \6295_b1 , w_15768 );
and ( \6429_b0 , \6048_b0 , w_15769 );
and ( w_15768 , w_15769 , \6295_b0 );
or ( \6430_b1 , \6428_b1 , w_15771 );
not ( w_15771 , w_15772 );
and ( \6430_b0 , \6428_b0 , w_15773 );
and ( w_15772 ,  , w_15773 );
buf ( w_15771 , \6429_b1 );
not ( w_15771 , w_15774 );
not (  , w_15775 );
and ( w_15774 , w_15775 , \6429_b0 );
or ( \6431_b1 , \6430_b1 , w_15776 );
xor ( \6431_b0 , \6430_b0 , w_15778 );
not ( w_15778 , w_15779 );
and ( w_15779 , w_15776 , w_15777 );
buf ( w_15776 , \6227_b1 );
not ( w_15776 , w_15780 );
not ( w_15777 , w_15781 );
and ( w_15780 , w_15781 , \6227_b0 );
or ( \6432_b1 , \6424_b1 , \6431_b1 );
xor ( \6432_b0 , \6424_b0 , w_15782 );
not ( w_15782 , w_15783 );
and ( w_15783 , \6431_b1 , \6431_b0 );
or ( \6433_b1 , \5998_b1 , \6016_b1 );
not ( \6016_b1 , w_15784 );
and ( \6433_b0 , \5998_b0 , w_15785 );
and ( w_15784 , w_15785 , \6016_b0 );
or ( \6434_b1 , \5967_b1 , \6014_b1 );
not ( \6014_b1 , w_15786 );
and ( \6434_b0 , \5967_b0 , w_15787 );
and ( w_15786 , w_15787 , \6014_b0 );
or ( \6435_b1 , \6433_b1 , w_15789 );
not ( w_15789 , w_15790 );
and ( \6435_b0 , \6433_b0 , w_15791 );
and ( w_15790 ,  , w_15791 );
buf ( w_15789 , \6434_b1 );
not ( w_15789 , w_15792 );
not (  , w_15793 );
and ( w_15792 , w_15793 , \6434_b0 );
or ( \6436_b1 , \6435_b1 , w_15794 );
xor ( \6436_b0 , \6435_b0 , w_15796 );
not ( w_15796 , w_15797 );
and ( w_15797 , w_15794 , w_15795 );
buf ( w_15794 , \6023_b1 );
not ( w_15794 , w_15798 );
not ( w_15795 , w_15799 );
and ( w_15798 , w_15799 , \6023_b0 );
or ( \6437_b1 , \6018_b1 , \6039_b1 );
not ( \6039_b1 , w_15800 );
and ( \6437_b0 , \6018_b0 , w_15801 );
and ( w_15800 , w_15801 , \6039_b0 );
or ( \6438_b1 , \5986_b1 , \6037_b1 );
not ( \6037_b1 , w_15802 );
and ( \6438_b0 , \5986_b0 , w_15803 );
and ( w_15802 , w_15803 , \6037_b0 );
or ( \6439_b1 , \6437_b1 , w_15805 );
not ( w_15805 , w_15806 );
and ( \6439_b0 , \6437_b0 , w_15807 );
and ( w_15806 ,  , w_15807 );
buf ( w_15805 , \6438_b1 );
not ( w_15805 , w_15808 );
not (  , w_15809 );
and ( w_15808 , w_15809 , \6438_b0 );
or ( \6440_b1 , \6439_b1 , w_15810 );
xor ( \6440_b0 , \6439_b0 , w_15812 );
not ( w_15812 , w_15813 );
and ( w_15813 , w_15810 , w_15811 );
buf ( w_15810 , \6046_b1 );
not ( w_15810 , w_15814 );
not ( w_15811 , w_15815 );
and ( w_15814 , w_15815 , \6046_b0 );
or ( \6441_b1 , \6436_b1 , \6440_b1 );
xor ( \6441_b0 , \6436_b0 , w_15816 );
not ( w_15816 , w_15817 );
and ( w_15817 , \6440_b1 , \6440_b0 );
or ( \6442_b1 , \6041_b1 , \6055_b1 );
not ( \6055_b1 , w_15818 );
and ( \6442_b0 , \6041_b0 , w_15819 );
and ( w_15818 , w_15819 , \6055_b0 );
or ( \6443_b1 , \6006_b1 , \6053_b1 );
not ( \6053_b1 , w_15820 );
and ( \6443_b0 , \6006_b0 , w_15821 );
and ( w_15820 , w_15821 , \6053_b0 );
or ( \6444_b1 , \6442_b1 , w_15823 );
not ( w_15823 , w_15824 );
and ( \6444_b0 , \6442_b0 , w_15825 );
and ( w_15824 ,  , w_15825 );
buf ( w_15823 , \6443_b1 );
not ( w_15823 , w_15826 );
not (  , w_15827 );
and ( w_15826 , w_15827 , \6443_b0 );
or ( \6445_b1 , \6444_b1 , w_15828 );
xor ( \6445_b0 , \6444_b0 , w_15830 );
not ( w_15830 , w_15831 );
and ( w_15831 , w_15828 , w_15829 );
buf ( w_15828 , \6062_b1 );
not ( w_15828 , w_15832 );
not ( w_15829 , w_15833 );
and ( w_15832 , w_15833 , \6062_b0 );
or ( \6446_b1 , \6441_b1 , \6445_b1 );
xor ( \6446_b0 , \6441_b0 , w_15834 );
not ( w_15834 , w_15835 );
and ( w_15835 , \6445_b1 , \6445_b0 );
or ( \6447_b1 , \6432_b1 , \6446_b1 );
xor ( \6447_b0 , \6432_b0 , w_15836 );
not ( w_15836 , w_15837 );
and ( w_15837 , \6446_b1 , \6446_b0 );
or ( \6448_b1 , \5937_b1 , \5955_b1 );
not ( \5955_b1 , w_15838 );
and ( \6448_b0 , \5937_b0 , w_15839 );
and ( w_15838 , w_15839 , \5955_b0 );
or ( \6449_b1 , \5906_b1 , \5953_b1 );
not ( \5953_b1 , w_15840 );
and ( \6449_b0 , \5906_b0 , w_15841 );
and ( w_15840 , w_15841 , \5953_b0 );
or ( \6450_b1 , \6448_b1 , w_15843 );
not ( w_15843 , w_15844 );
and ( \6450_b0 , \6448_b0 , w_15845 );
and ( w_15844 ,  , w_15845 );
buf ( w_15843 , \6449_b1 );
not ( w_15843 , w_15846 );
not (  , w_15847 );
and ( w_15846 , w_15847 , \6449_b0 );
or ( \6451_b1 , \6450_b1 , w_15848 );
xor ( \6451_b0 , \6450_b0 , w_15850 );
not ( w_15850 , w_15851 );
and ( w_15851 , w_15848 , w_15849 );
buf ( w_15848 , \5962_b1 );
not ( w_15848 , w_15852 );
not ( w_15849 , w_15853 );
and ( w_15852 , w_15853 , \5962_b0 );
or ( \6452_b1 , \5957_b1 , \5977_b1 );
not ( \5977_b1 , w_15854 );
and ( \6452_b0 , \5957_b0 , w_15855 );
and ( w_15854 , w_15855 , \5977_b0 );
or ( \6453_b1 , \5925_b1 , \5975_b1 );
not ( \5975_b1 , w_15856 );
and ( \6453_b0 , \5925_b0 , w_15857 );
and ( w_15856 , w_15857 , \5975_b0 );
or ( \6454_b1 , \6452_b1 , w_15859 );
not ( w_15859 , w_15860 );
and ( \6454_b0 , \6452_b0 , w_15861 );
and ( w_15860 ,  , w_15861 );
buf ( w_15859 , \6453_b1 );
not ( w_15859 , w_15862 );
not (  , w_15863 );
and ( w_15862 , w_15863 , \6453_b0 );
or ( \6455_b1 , \6454_b1 , w_15864 );
xor ( \6455_b0 , \6454_b0 , w_15866 );
not ( w_15866 , w_15867 );
and ( w_15867 , w_15864 , w_15865 );
buf ( w_15864 , \5984_b1 );
not ( w_15864 , w_15868 );
not ( w_15865 , w_15869 );
and ( w_15868 , w_15869 , \5984_b0 );
or ( \6456_b1 , \6451_b1 , \6455_b1 );
xor ( \6456_b0 , \6451_b0 , w_15870 );
not ( w_15870 , w_15871 );
and ( w_15871 , \6455_b1 , \6455_b0 );
or ( \6457_b1 , \5979_b1 , \5996_b1 );
not ( \5996_b1 , w_15872 );
and ( \6457_b0 , \5979_b0 , w_15873 );
and ( w_15872 , w_15873 , \5996_b0 );
or ( \6458_b1 , \5945_b1 , \5994_b1 );
not ( \5994_b1 , w_15874 );
and ( \6458_b0 , \5945_b0 , w_15875 );
and ( w_15874 , w_15875 , \5994_b0 );
or ( \6459_b1 , \6457_b1 , w_15877 );
not ( w_15877 , w_15878 );
and ( \6459_b0 , \6457_b0 , w_15879 );
and ( w_15878 ,  , w_15879 );
buf ( w_15877 , \6458_b1 );
not ( w_15877 , w_15880 );
not (  , w_15881 );
and ( w_15880 , w_15881 , \6458_b0 );
or ( \6460_b1 , \6459_b1 , w_15882 );
xor ( \6460_b0 , \6459_b0 , w_15884 );
not ( w_15884 , w_15885 );
and ( w_15885 , w_15882 , w_15883 );
buf ( w_15882 , \6003_b1 );
not ( w_15882 , w_15886 );
not ( w_15883 , w_15887 );
and ( w_15886 , w_15887 , \6003_b0 );
or ( \6461_b1 , \6456_b1 , \6460_b1 );
xor ( \6461_b0 , \6456_b0 , w_15888 );
not ( w_15888 , w_15889 );
and ( w_15889 , \6460_b1 , \6460_b0 );
or ( \6462_b1 , \6447_b1 , \6461_b1 );
xor ( \6462_b0 , \6447_b0 , w_15890 );
not ( w_15890 , w_15891 );
and ( w_15891 , \6461_b1 , \6461_b0 );
or ( \6463_b1 , \6420_b1 , \6462_b1 );
xor ( \6463_b0 , \6420_b0 , w_15892 );
not ( w_15892 , w_15893 );
and ( w_15893 , \6462_b1 , \6462_b0 );
or ( \6464_b1 , \6374_b1 , \6463_b1 );
not ( \6463_b1 , w_15894 );
and ( \6464_b0 , \6374_b0 , w_15895 );
and ( w_15894 , w_15895 , \6463_b0 );
or ( \6465_b1 , \6329_b1 , \6333_b1 );
not ( \6333_b1 , w_15896 );
and ( \6465_b0 , \6329_b0 , w_15897 );
and ( w_15896 , w_15897 , \6333_b0 );
or ( \6466_b1 , \6333_b1 , \6338_b1 );
not ( \6338_b1 , w_15898 );
and ( \6466_b0 , \6333_b0 , w_15899 );
and ( w_15898 , w_15899 , \6338_b0 );
or ( \6467_b1 , \6329_b1 , \6338_b1 );
not ( \6338_b1 , w_15900 );
and ( \6467_b0 , \6329_b0 , w_15901 );
and ( w_15900 , w_15901 , \6338_b0 );
or ( \6469_b1 , \6317_b1 , \6321_b1 );
not ( \6321_b1 , w_15902 );
and ( \6469_b0 , \6317_b0 , w_15903 );
and ( w_15902 , w_15903 , \6321_b0 );
or ( \6470_b1 , \6321_b1 , \6323_b1 );
not ( \6323_b1 , w_15904 );
and ( \6470_b0 , \6321_b0 , w_15905 );
and ( w_15904 , w_15905 , \6323_b0 );
or ( \6471_b1 , \6317_b1 , \6323_b1 );
not ( \6323_b1 , w_15906 );
and ( \6471_b0 , \6317_b0 , w_15907 );
and ( w_15906 , w_15907 , \6323_b0 );
or ( \6473_b1 , \6468_b1 , \6472_b1 );
xor ( \6473_b0 , \6468_b0 , w_15908 );
not ( w_15908 , w_15909 );
and ( w_15909 , \6472_b1 , \6472_b0 );
or ( \6474_b1 , \6298_b1 , w_15910 );
or ( \6474_b0 , \6298_b0 , \6312_b0 );
not ( \6312_b0 , w_15911 );
and ( w_15911 , w_15910 , \6312_b1 );
or ( \6475_b1 , \6473_b1 , \6474_b1 );
xor ( \6475_b0 , \6473_b0 , w_15912 );
not ( w_15912 , w_15913 );
and ( w_15913 , \6474_b1 , \6474_b0 );
or ( \6476_b1 , \6463_b1 , \6475_b1 );
not ( \6475_b1 , w_15914 );
and ( \6476_b0 , \6463_b0 , w_15915 );
and ( w_15914 , w_15915 , \6475_b0 );
or ( \6477_b1 , \6374_b1 , \6475_b1 );
not ( \6475_b1 , w_15916 );
and ( \6477_b0 , \6374_b0 , w_15917 );
and ( w_15916 , w_15917 , \6475_b0 );
or ( \6479_b1 , \6345_b1 , \6478_b1 );
not ( \6478_b1 , w_15918 );
and ( \6479_b0 , \6345_b0 , w_15919 );
and ( w_15918 , w_15919 , \6478_b0 );
or ( \6480_b1 , \6029_b1 , \6082_b1 );
not ( \6082_b1 , w_15920 );
and ( \6480_b0 , \6029_b0 , w_15921 );
and ( w_15920 , w_15921 , \6082_b0 );
or ( \6481_b1 , \6041_b1 , \6066_b1 );
not ( \6066_b1 , w_15922 );
and ( \6481_b0 , \6041_b0 , w_15923 );
and ( w_15922 , w_15923 , \6066_b0 );
or ( \6482_b1 , \6480_b1 , w_15925 );
not ( w_15925 , w_15926 );
and ( \6482_b0 , \6480_b0 , w_15927 );
and ( w_15926 ,  , w_15927 );
buf ( w_15925 , \6481_b1 );
not ( w_15925 , w_15928 );
not (  , w_15929 );
and ( w_15928 , w_15929 , \6481_b0 );
or ( \6483_b1 , \6482_b1 , w_15930 );
xor ( \6483_b0 , \6482_b0 , w_15932 );
not ( w_15932 , w_15933 );
and ( w_15933 , w_15930 , w_15931 );
buf ( w_15930 , \5736_b1 );
not ( w_15930 , w_15934 );
not ( w_15931 , w_15935 );
and ( w_15934 , w_15935 , \5736_b0 );
or ( \6484_b1 , \6048_b1 , \6427_b1 );
not ( \6427_b1 , w_15936 );
and ( \6484_b0 , \6048_b0 , w_15937 );
and ( w_15936 , w_15937 , \6427_b0 );
or ( \6485_b1 , \6057_b1 , \6295_b1 );
not ( \6295_b1 , w_15938 );
and ( \6485_b0 , \6057_b0 , w_15939 );
and ( w_15938 , w_15939 , \6295_b0 );
or ( \6486_b1 , \6484_b1 , w_15941 );
not ( w_15941 , w_15942 );
and ( \6486_b0 , \6484_b0 , w_15943 );
and ( w_15942 ,  , w_15943 );
buf ( w_15941 , \6485_b1 );
not ( w_15941 , w_15944 );
not (  , w_15945 );
and ( w_15944 , w_15945 , \6485_b0 );
or ( \6487_b1 , \6486_b1 , w_15946 );
xor ( \6487_b0 , \6486_b0 , w_15948 );
not ( w_15948 , w_15949 );
and ( w_15949 , w_15946 , w_15947 );
buf ( w_15946 , \6227_b1 );
not ( w_15946 , w_15950 );
not ( w_15947 , w_15951 );
and ( w_15950 , w_15951 , \6227_b0 );
or ( \6488_b1 , \6483_b1 , \6487_b1 );
xor ( \6488_b0 , \6483_b0 , w_15952 );
not ( w_15952 , w_15953 );
and ( w_15953 , \6487_b1 , \6487_b0 );
or ( \6489_b1 , \6186_b1 , \6190_b1 );
not ( \6190_b1 , w_15954 );
and ( \6489_b0 , \6186_b0 , w_15955 );
and ( w_15954 , w_15955 , \6190_b0 );
or ( \6490_b1 , \6190_b1 , \6192_b1 );
not ( \6192_b1 , w_15956 );
and ( \6490_b0 , \6190_b0 , w_15957 );
and ( w_15956 , w_15957 , \6192_b0 );
or ( \6491_b1 , \6186_b1 , \6192_b1 );
not ( \6192_b1 , w_15958 );
and ( \6491_b0 , \6186_b0 , w_15959 );
and ( w_15958 , w_15959 , \6192_b0 );
or ( \6493_b1 , \159_b1 , \351_b1 );
not ( \351_b1 , w_15960 );
and ( \6493_b0 , \159_b0 , w_15961 );
and ( w_15960 , w_15961 , \351_b0 );
buf ( \6494_b1 , \6493_b1 );
not ( \6494_b1 , w_15962 );
not ( \6494_b0 , w_15963 );
and ( w_15962 , w_15963 , \6493_b0 );
or ( \6495_b1 , \6494_b1 , w_15964 );
xor ( \6495_b0 , \6494_b0 , w_15966 );
not ( w_15966 , w_15967 );
and ( w_15967 , w_15964 , w_15965 );
buf ( w_15964 , \358_b1 );
not ( w_15964 , w_15968 );
not ( w_15965 , w_15969 );
and ( w_15968 , w_15969 , \358_b0 );
or ( \6496_b1 , \315_b1 , \345_b1 );
not ( \345_b1 , w_15970 );
and ( \6496_b0 , \315_b0 , w_15971 );
and ( w_15970 , w_15971 , \345_b0 );
or ( \6497_b1 , \6495_b1 , w_15972 );
xor ( \6497_b0 , \6495_b0 , w_15974 );
not ( w_15974 , w_15975 );
and ( w_15975 , w_15972 , w_15973 );
buf ( w_15972 , \6496_b1 );
not ( w_15972 , w_15976 );
not ( w_15973 , w_15977 );
and ( w_15976 , w_15977 , \6496_b0 );
or ( \6498_b1 , \6492_b1 , \6497_b1 );
xor ( \6498_b0 , \6492_b0 , w_15978 );
not ( w_15978 , w_15979 );
and ( w_15979 , \6497_b1 , \6497_b0 );
or ( \6499_b1 , \6177_b1 , \6184_b1 );
not ( \6184_b1 , w_15980 );
and ( \6499_b0 , \6177_b0 , w_15981 );
and ( w_15980 , w_15981 , \6184_b0 );
or ( \6500_b1 , \6184_b1 , \6193_b1 );
not ( \6193_b1 , w_15982 );
and ( \6500_b0 , \6184_b0 , w_15983 );
and ( w_15982 , w_15983 , \6193_b0 );
or ( \6501_b1 , \6177_b1 , \6193_b1 );
not ( \6193_b1 , w_15984 );
and ( \6501_b0 , \6177_b0 , w_15985 );
and ( w_15984 , w_15985 , \6193_b0 );
or ( \6503_b1 , \6498_b1 , \6502_b1 );
xor ( \6503_b0 , \6498_b0 , w_15986 );
not ( w_15986 , w_15987 );
and ( w_15987 , \6502_b1 , \6502_b0 );
or ( \6504_b1 , \6194_b1 , \6207_b1 );
not ( \6207_b1 , w_15988 );
and ( \6504_b0 , \6194_b0 , w_15989 );
and ( w_15988 , w_15989 , \6207_b0 );
or ( \6505_b1 , \6208_b1 , \6218_b1 );
not ( \6218_b1 , w_15990 );
and ( \6505_b0 , \6208_b0 , w_15991 );
and ( w_15990 , w_15991 , \6218_b0 );
or ( \6506_b1 , \6504_b1 , w_15992 );
or ( \6506_b0 , \6504_b0 , \6505_b0 );
not ( \6505_b0 , w_15993 );
and ( w_15993 , w_15992 , \6505_b1 );
or ( \6507_b1 , \6503_b1 , \6506_b1 );
xor ( \6507_b0 , \6503_b0 , w_15994 );
not ( w_15994 , w_15995 );
and ( w_15995 , \6506_b1 , \6506_b0 );
buf ( \6508_b1 , \6507_b1 );
buf ( \6508_b0 , \6507_b0 );
buf ( \6509_b1 , \6508_b1 );
buf ( \6509_b0 , \6508_b0 );
or ( \6510_b1 , \6509_b1 , \6221_b1 );
xor ( \6510_b0 , \6509_b0 , w_15996 );
not ( w_15996 , w_15997 );
and ( w_15997 , \6221_b1 , \6221_b0 );
or ( \6511_b1 , \6065_b1 , w_15999 );
not ( w_15999 , w_16000 );
and ( \6511_b0 , \6065_b0 , w_16001 );
and ( w_16000 ,  , w_16001 );
buf ( w_15999 , \6510_b1 );
not ( w_15999 , w_16002 );
not (  , w_16003 );
and ( w_16002 , w_16003 , \6510_b0 );
or ( \6512_b1 , \6495_b1 , w_16004 );
or ( \6512_b0 , \6495_b0 , \6496_b0 );
not ( \6496_b0 , w_16005 );
and ( w_16005 , w_16004 , \6496_b1 );
buf ( \6513_b1 , \358_b1 );
not ( \6513_b1 , w_16006 );
not ( \6513_b0 , w_16007 );
and ( w_16006 , w_16007 , \358_b0 );
or ( \6514_b1 , \6512_b1 , \6513_b1 );
xor ( \6514_b0 , \6512_b0 , w_16008 );
not ( w_16008 , w_16009 );
and ( w_16009 , \6513_b1 , \6513_b0 );
or ( \6515_b1 , \159_b1 , \345_b1 );
not ( \345_b1 , w_16010 );
and ( \6515_b0 , \159_b0 , w_16011 );
and ( w_16010 , w_16011 , \345_b0 );
or ( \6516_b1 , \6514_b1 , \6515_b1 );
xor ( \6516_b0 , \6514_b0 , w_16012 );
not ( w_16012 , w_16013 );
and ( w_16013 , \6515_b1 , \6515_b0 );
or ( \6517_b1 , \6492_b1 , \6497_b1 );
not ( \6497_b1 , w_16014 );
and ( \6517_b0 , \6492_b0 , w_16015 );
and ( w_16014 , w_16015 , \6497_b0 );
or ( \6518_b1 , \6516_b1 , \6517_b1 );
xor ( \6518_b0 , \6516_b0 , w_16016 );
not ( w_16016 , w_16017 );
and ( w_16017 , \6517_b1 , \6517_b0 );
or ( \6519_b1 , \6498_b1 , \6502_b1 );
not ( \6502_b1 , w_16018 );
and ( \6519_b0 , \6498_b0 , w_16019 );
and ( w_16018 , w_16019 , \6502_b0 );
or ( \6520_b1 , \6503_b1 , \6506_b1 );
not ( \6506_b1 , w_16020 );
and ( \6520_b0 , \6503_b0 , w_16021 );
and ( w_16020 , w_16021 , \6506_b0 );
or ( \6521_b1 , \6519_b1 , w_16022 );
or ( \6521_b0 , \6519_b0 , \6520_b0 );
not ( \6520_b0 , w_16023 );
and ( w_16023 , w_16022 , \6520_b1 );
or ( \6522_b1 , \6518_b1 , \6521_b1 );
xor ( \6522_b0 , \6518_b0 , w_16024 );
not ( w_16024 , w_16025 );
and ( w_16025 , \6521_b1 , \6521_b0 );
buf ( \6523_b1 , \6522_b1 );
buf ( \6523_b0 , \6522_b0 );
buf ( \6524_b1 , \6523_b1 );
buf ( \6524_b0 , \6523_b0 );
or ( \6525_b1 , \6509_b1 , \6221_b1 );
not ( \6221_b1 , w_16026 );
and ( \6525_b0 , \6509_b0 , w_16027 );
and ( w_16026 , w_16027 , \6221_b0 );
buf ( \6526_b1 , \6525_b1 );
not ( \6526_b1 , w_16028 );
not ( \6526_b0 , w_16029 );
and ( w_16028 , w_16029 , \6525_b0 );
or ( \6527_b1 , \6524_b1 , \6526_b1 );
not ( \6526_b1 , w_16030 );
and ( \6527_b0 , \6524_b0 , w_16031 );
and ( w_16030 , w_16031 , \6526_b0 );
or ( \6528_b1 , \6511_b1 , w_16032 );
xor ( \6528_b0 , \6511_b0 , w_16034 );
not ( w_16034 , w_16035 );
and ( w_16035 , w_16032 , w_16033 );
buf ( w_16032 , \6527_b1 );
not ( w_16032 , w_16036 );
not ( w_16033 , w_16037 );
and ( w_16036 , w_16037 , \6527_b0 );
or ( \6529_b1 , \6488_b1 , \6528_b1 );
xor ( \6529_b0 , \6488_b0 , w_16038 );
not ( w_16038 , w_16039 );
and ( w_16039 , \6528_b1 , \6528_b0 );
or ( \6530_b1 , \5967_b1 , \6016_b1 );
not ( \6016_b1 , w_16040 );
and ( \6530_b0 , \5967_b0 , w_16041 );
and ( w_16040 , w_16041 , \6016_b0 );
or ( \6531_b1 , \5979_b1 , \6014_b1 );
not ( \6014_b1 , w_16042 );
and ( \6531_b0 , \5979_b0 , w_16043 );
and ( w_16042 , w_16043 , \6014_b0 );
or ( \6532_b1 , \6530_b1 , w_16045 );
not ( w_16045 , w_16046 );
and ( \6532_b0 , \6530_b0 , w_16047 );
and ( w_16046 ,  , w_16047 );
buf ( w_16045 , \6531_b1 );
not ( w_16045 , w_16048 );
not (  , w_16049 );
and ( w_16048 , w_16049 , \6531_b0 );
or ( \6533_b1 , \6532_b1 , w_16050 );
xor ( \6533_b0 , \6532_b0 , w_16052 );
not ( w_16052 , w_16053 );
and ( w_16053 , w_16050 , w_16051 );
buf ( w_16050 , \6023_b1 );
not ( w_16050 , w_16054 );
not ( w_16051 , w_16055 );
and ( w_16054 , w_16055 , \6023_b0 );
or ( \6534_b1 , \5986_b1 , \6039_b1 );
not ( \6039_b1 , w_16056 );
and ( \6534_b0 , \5986_b0 , w_16057 );
and ( w_16056 , w_16057 , \6039_b0 );
or ( \6535_b1 , \5998_b1 , \6037_b1 );
not ( \6037_b1 , w_16058 );
and ( \6535_b0 , \5998_b0 , w_16059 );
and ( w_16058 , w_16059 , \6037_b0 );
or ( \6536_b1 , \6534_b1 , w_16061 );
not ( w_16061 , w_16062 );
and ( \6536_b0 , \6534_b0 , w_16063 );
and ( w_16062 ,  , w_16063 );
buf ( w_16061 , \6535_b1 );
not ( w_16061 , w_16064 );
not (  , w_16065 );
and ( w_16064 , w_16065 , \6535_b0 );
or ( \6537_b1 , \6536_b1 , w_16066 );
xor ( \6537_b0 , \6536_b0 , w_16068 );
not ( w_16068 , w_16069 );
and ( w_16069 , w_16066 , w_16067 );
buf ( w_16066 , \6046_b1 );
not ( w_16066 , w_16070 );
not ( w_16067 , w_16071 );
and ( w_16070 , w_16071 , \6046_b0 );
or ( \6538_b1 , \6533_b1 , \6537_b1 );
xor ( \6538_b0 , \6533_b0 , w_16072 );
not ( w_16072 , w_16073 );
and ( w_16073 , \6537_b1 , \6537_b0 );
or ( \6539_b1 , \6006_b1 , \6055_b1 );
not ( \6055_b1 , w_16074 );
and ( \6539_b0 , \6006_b0 , w_16075 );
and ( w_16074 , w_16075 , \6055_b0 );
or ( \6540_b1 , \6018_b1 , \6053_b1 );
not ( \6053_b1 , w_16076 );
and ( \6540_b0 , \6018_b0 , w_16077 );
and ( w_16076 , w_16077 , \6053_b0 );
or ( \6541_b1 , \6539_b1 , w_16079 );
not ( w_16079 , w_16080 );
and ( \6541_b0 , \6539_b0 , w_16081 );
and ( w_16080 ,  , w_16081 );
buf ( w_16079 , \6540_b1 );
not ( w_16079 , w_16082 );
not (  , w_16083 );
and ( w_16082 , w_16083 , \6540_b0 );
or ( \6542_b1 , \6541_b1 , w_16084 );
xor ( \6542_b0 , \6541_b0 , w_16086 );
not ( w_16086 , w_16087 );
and ( w_16087 , w_16084 , w_16085 );
buf ( w_16084 , \6062_b1 );
not ( w_16084 , w_16088 );
not ( w_16085 , w_16089 );
and ( w_16088 , w_16089 , \6062_b0 );
or ( \6543_b1 , \6538_b1 , \6542_b1 );
xor ( \6543_b0 , \6538_b0 , w_16090 );
not ( w_16090 , w_16091 );
and ( w_16091 , \6542_b1 , \6542_b0 );
or ( \6544_b1 , \6529_b1 , w_16092 );
xor ( \6544_b0 , \6529_b0 , w_16094 );
not ( w_16094 , w_16095 );
and ( w_16095 , w_16092 , w_16093 );
buf ( w_16092 , \6543_b1 );
not ( w_16092 , w_16096 );
not ( w_16093 , w_16097 );
and ( w_16096 , w_16097 , \6543_b0 );
or ( \6545_b1 , \6451_b1 , \6455_b1 );
not ( \6455_b1 , w_16098 );
and ( \6545_b0 , \6451_b0 , w_16099 );
and ( w_16098 , w_16099 , \6455_b0 );
or ( \6546_b1 , \6455_b1 , \6460_b1 );
not ( \6460_b1 , w_16100 );
and ( \6546_b0 , \6455_b0 , w_16101 );
and ( w_16100 , w_16101 , \6460_b0 );
or ( \6547_b1 , \6451_b1 , \6460_b1 );
not ( \6460_b1 , w_16102 );
and ( \6547_b0 , \6451_b0 , w_16103 );
and ( w_16102 , w_16103 , \6460_b0 );
or ( \6549_b1 , \6436_b1 , \6440_b1 );
not ( \6440_b1 , w_16104 );
and ( \6549_b0 , \6436_b0 , w_16105 );
and ( w_16104 , w_16105 , \6440_b0 );
or ( \6550_b1 , \6440_b1 , \6445_b1 );
not ( \6445_b1 , w_16106 );
and ( \6550_b0 , \6440_b0 , w_16107 );
and ( w_16106 , w_16107 , \6445_b0 );
or ( \6551_b1 , \6436_b1 , \6445_b1 );
not ( \6445_b1 , w_16108 );
and ( \6551_b0 , \6436_b0 , w_16109 );
and ( w_16108 , w_16109 , \6445_b0 );
or ( \6553_b1 , \6548_b1 , \6552_b1 );
xor ( \6553_b0 , \6548_b0 , w_16110 );
not ( w_16110 , w_16111 );
and ( w_16111 , \6552_b1 , \6552_b0 );
or ( \6554_b1 , \6424_b1 , \6431_b1 );
not ( \6431_b1 , w_16112 );
and ( \6554_b0 , \6424_b0 , w_16113 );
and ( w_16112 , w_16113 , \6431_b0 );
or ( \6555_b1 , \6553_b1 , \6554_b1 );
xor ( \6555_b0 , \6553_b0 , w_16114 );
not ( w_16114 , w_16115 );
and ( w_16115 , \6554_b1 , \6554_b0 );
or ( \6556_b1 , \6544_b1 , \6555_b1 );
xor ( \6556_b0 , \6544_b0 , w_16116 );
not ( w_16116 , w_16117 );
and ( w_16117 , \6555_b1 , \6555_b0 );
or ( \6557_b1 , \6408_b1 , \6412_b1 );
not ( \6412_b1 , w_16118 );
and ( \6557_b0 , \6408_b0 , w_16119 );
and ( w_16118 , w_16119 , \6412_b0 );
or ( \6558_b1 , \6412_b1 , \6417_b1 );
not ( \6417_b1 , w_16120 );
and ( \6558_b0 , \6412_b0 , w_16121 );
and ( w_16120 , w_16121 , \6417_b0 );
or ( \6559_b1 , \6408_b1 , \6417_b1 );
not ( \6417_b1 , w_16122 );
and ( \6559_b0 , \6408_b0 , w_16123 );
and ( w_16122 , w_16123 , \6417_b0 );
or ( \6561_b1 , \6396_b1 , \6400_b1 );
not ( \6400_b1 , w_16124 );
and ( \6561_b0 , \6396_b0 , w_16125 );
and ( w_16124 , w_16125 , \6400_b0 );
or ( \6562_b1 , \6400_b1 , \6405_b1 );
not ( \6405_b1 , w_16126 );
and ( \6562_b0 , \6400_b0 , w_16127 );
and ( w_16126 , w_16127 , \6405_b0 );
or ( \6563_b1 , \6396_b1 , \6405_b1 );
not ( \6405_b1 , w_16128 );
and ( \6563_b0 , \6396_b0 , w_16129 );
and ( w_16128 , w_16129 , \6405_b0 );
or ( \6565_b1 , \6560_b1 , \6564_b1 );
xor ( \6565_b0 , \6560_b0 , w_16130 );
not ( w_16130 , w_16131 );
and ( w_16131 , \6564_b1 , \6564_b0 );
or ( \6566_b1 , \6382_b1 , \6386_b1 );
not ( \6386_b1 , w_16132 );
and ( \6566_b0 , \6382_b0 , w_16133 );
and ( w_16132 , w_16133 , \6386_b0 );
or ( \6567_b1 , \6386_b1 , \6391_b1 );
not ( \6391_b1 , w_16134 );
and ( \6567_b0 , \6386_b0 , w_16135 );
and ( w_16134 , w_16135 , \6391_b0 );
or ( \6568_b1 , \6382_b1 , \6391_b1 );
not ( \6391_b1 , w_16136 );
and ( \6568_b0 , \6382_b0 , w_16137 );
and ( w_16136 , w_16137 , \6391_b0 );
or ( \6570_b1 , \6565_b1 , \6569_b1 );
xor ( \6570_b0 , \6565_b0 , w_16138 );
not ( w_16138 , w_16139 );
and ( w_16139 , \6569_b1 , \6569_b0 );
or ( \6571_b1 , \6556_b1 , \6570_b1 );
xor ( \6571_b0 , \6556_b0 , w_16140 );
not ( w_16140 , w_16141 );
and ( w_16141 , \6570_b1 , \6570_b0 );
or ( \6572_b1 , \6392_b1 , \6406_b1 );
not ( \6406_b1 , w_16142 );
and ( \6572_b0 , \6392_b0 , w_16143 );
and ( w_16142 , w_16143 , \6406_b0 );
or ( \6573_b1 , \6406_b1 , \6418_b1 );
not ( \6418_b1 , w_16144 );
and ( \6573_b0 , \6406_b0 , w_16145 );
and ( w_16144 , w_16145 , \6418_b0 );
or ( \6574_b1 , \6392_b1 , \6418_b1 );
not ( \6418_b1 , w_16146 );
and ( \6574_b0 , \6392_b0 , w_16147 );
and ( w_16146 , w_16147 , \6418_b0 );
or ( \6576_b1 , \5737_b1 , \5790_b1 );
not ( \5790_b1 , w_16148 );
and ( \6576_b0 , \5737_b0 , w_16149 );
and ( w_16148 , w_16149 , \5790_b0 );
buf ( \6577_b1 , \6576_b1 );
not ( \6577_b1 , w_16150 );
not ( \6577_b0 , w_16151 );
and ( w_16150 , w_16151 , \6576_b0 );
or ( \6578_b1 , \6577_b1 , w_16152 );
xor ( \6578_b0 , \6577_b0 , w_16154 );
not ( w_16154 , w_16155 );
and ( w_16155 , w_16152 , w_16153 );
buf ( w_16152 , \5797_b1 );
not ( w_16152 , w_16156 );
not ( w_16153 , w_16157 );
and ( w_16156 , w_16157 , \5797_b0 );
or ( \6579_b1 , \6527_b1 , \6578_b1 );
xor ( \6579_b0 , \6527_b0 , w_16158 );
not ( w_16158 , w_16159 );
and ( w_16159 , \6578_b1 , \6578_b0 );
or ( \6580_b1 , \5758_b1 , \5809_b1 );
not ( \5809_b1 , w_16160 );
and ( \6580_b0 , \5758_b0 , w_16161 );
and ( w_16160 , w_16161 , \5809_b0 );
or ( \6581_b1 , \5770_b1 , \5807_b1 );
not ( \5807_b1 , w_16162 );
and ( \6581_b0 , \5770_b0 , w_16163 );
and ( w_16162 , w_16163 , \5807_b0 );
or ( \6582_b1 , \6580_b1 , w_16165 );
not ( w_16165 , w_16166 );
and ( \6582_b0 , \6580_b0 , w_16167 );
and ( w_16166 ,  , w_16167 );
buf ( w_16165 , \6581_b1 );
not ( w_16165 , w_16168 );
not (  , w_16169 );
and ( w_16168 , w_16169 , \6581_b0 );
or ( \6583_b1 , \6582_b1 , w_16170 );
xor ( \6583_b0 , \6582_b0 , w_16172 );
not ( w_16172 , w_16173 );
and ( w_16173 , w_16170 , w_16171 );
buf ( w_16170 , \5816_b1 );
not ( w_16170 , w_16174 );
not ( w_16171 , w_16175 );
and ( w_16174 , w_16175 , \5816_b0 );
or ( \6584_b1 , \6579_b1 , \6583_b1 );
xor ( \6584_b0 , \6579_b0 , w_16176 );
not ( w_16176 , w_16177 );
and ( w_16177 , \6583_b1 , \6583_b0 );
or ( \6585_b1 , \6575_b1 , \6584_b1 );
xor ( \6585_b0 , \6575_b0 , w_16178 );
not ( w_16178 , w_16179 );
and ( w_16179 , \6584_b1 , \6584_b0 );
or ( \6586_b1 , \5906_b1 , \5955_b1 );
not ( \5955_b1 , w_16180 );
and ( \6586_b0 , \5906_b0 , w_16181 );
and ( w_16180 , w_16181 , \5955_b0 );
or ( \6587_b1 , \5918_b1 , \5953_b1 );
not ( \5953_b1 , w_16182 );
and ( \6587_b0 , \5918_b0 , w_16183 );
and ( w_16182 , w_16183 , \5953_b0 );
or ( \6588_b1 , \6586_b1 , w_16185 );
not ( w_16185 , w_16186 );
and ( \6588_b0 , \6586_b0 , w_16187 );
and ( w_16186 ,  , w_16187 );
buf ( w_16185 , \6587_b1 );
not ( w_16185 , w_16188 );
not (  , w_16189 );
and ( w_16188 , w_16189 , \6587_b0 );
or ( \6589_b1 , \6588_b1 , w_16190 );
xor ( \6589_b0 , \6588_b0 , w_16192 );
not ( w_16192 , w_16193 );
and ( w_16193 , w_16190 , w_16191 );
buf ( w_16190 , \5962_b1 );
not ( w_16190 , w_16194 );
not ( w_16191 , w_16195 );
and ( w_16194 , w_16195 , \5962_b0 );
or ( \6590_b1 , \5925_b1 , \5977_b1 );
not ( \5977_b1 , w_16196 );
and ( \6590_b0 , \5925_b0 , w_16197 );
and ( w_16196 , w_16197 , \5977_b0 );
or ( \6591_b1 , \5937_b1 , \5975_b1 );
not ( \5975_b1 , w_16198 );
and ( \6591_b0 , \5937_b0 , w_16199 );
and ( w_16198 , w_16199 , \5975_b0 );
or ( \6592_b1 , \6590_b1 , w_16201 );
not ( w_16201 , w_16202 );
and ( \6592_b0 , \6590_b0 , w_16203 );
and ( w_16202 ,  , w_16203 );
buf ( w_16201 , \6591_b1 );
not ( w_16201 , w_16204 );
not (  , w_16205 );
and ( w_16204 , w_16205 , \6591_b0 );
or ( \6593_b1 , \6592_b1 , w_16206 );
xor ( \6593_b0 , \6592_b0 , w_16208 );
not ( w_16208 , w_16209 );
and ( w_16209 , w_16206 , w_16207 );
buf ( w_16206 , \5984_b1 );
not ( w_16206 , w_16210 );
not ( w_16207 , w_16211 );
and ( w_16210 , w_16211 , \5984_b0 );
or ( \6594_b1 , \6589_b1 , \6593_b1 );
xor ( \6594_b0 , \6589_b0 , w_16212 );
not ( w_16212 , w_16213 );
and ( w_16213 , \6593_b1 , \6593_b0 );
or ( \6595_b1 , \5945_b1 , \5996_b1 );
not ( \5996_b1 , w_16214 );
and ( \6595_b0 , \5945_b0 , w_16215 );
and ( w_16214 , w_16215 , \5996_b0 );
or ( \6596_b1 , \5957_b1 , \5994_b1 );
not ( \5994_b1 , w_16216 );
and ( \6596_b0 , \5957_b0 , w_16217 );
and ( w_16216 , w_16217 , \5994_b0 );
or ( \6597_b1 , \6595_b1 , w_16219 );
not ( w_16219 , w_16220 );
and ( \6597_b0 , \6595_b0 , w_16221 );
and ( w_16220 ,  , w_16221 );
buf ( w_16219 , \6596_b1 );
not ( w_16219 , w_16222 );
not (  , w_16223 );
and ( w_16222 , w_16223 , \6596_b0 );
or ( \6598_b1 , \6597_b1 , w_16224 );
xor ( \6598_b0 , \6597_b0 , w_16226 );
not ( w_16226 , w_16227 );
and ( w_16227 , w_16224 , w_16225 );
buf ( w_16224 , \6003_b1 );
not ( w_16224 , w_16228 );
not ( w_16225 , w_16229 );
and ( w_16228 , w_16229 , \6003_b0 );
or ( \6599_b1 , \6594_b1 , \6598_b1 );
xor ( \6599_b0 , \6594_b0 , w_16230 );
not ( w_16230 , w_16231 );
and ( w_16231 , \6598_b1 , \6598_b0 );
or ( \6600_b1 , \5842_b1 , \5891_b1 );
not ( \5891_b1 , w_16232 );
and ( \6600_b0 , \5842_b0 , w_16233 );
and ( w_16232 , w_16233 , \5891_b0 );
or ( \6601_b1 , \5854_b1 , \5889_b1 );
not ( \5889_b1 , w_16234 );
and ( \6601_b0 , \5854_b0 , w_16235 );
and ( w_16234 , w_16235 , \5889_b0 );
or ( \6602_b1 , \6600_b1 , w_16237 );
not ( w_16237 , w_16238 );
and ( \6602_b0 , \6600_b0 , w_16239 );
and ( w_16238 ,  , w_16239 );
buf ( w_16237 , \6601_b1 );
not ( w_16237 , w_16240 );
not (  , w_16241 );
and ( w_16240 , w_16241 , \6601_b0 );
or ( \6603_b1 , \6602_b1 , w_16242 );
xor ( \6603_b0 , \6602_b0 , w_16244 );
not ( w_16244 , w_16245 );
and ( w_16245 , w_16242 , w_16243 );
buf ( w_16242 , \5898_b1 );
not ( w_16242 , w_16246 );
not ( w_16243 , w_16247 );
and ( w_16246 , w_16247 , \5898_b0 );
or ( \6604_b1 , \5861_b1 , \5916_b1 );
not ( \5916_b1 , w_16248 );
and ( \6604_b0 , \5861_b0 , w_16249 );
and ( w_16248 , w_16249 , \5916_b0 );
or ( \6605_b1 , \5873_b1 , \5914_b1 );
not ( \5914_b1 , w_16250 );
and ( \6605_b0 , \5873_b0 , w_16251 );
and ( w_16250 , w_16251 , \5914_b0 );
or ( \6606_b1 , \6604_b1 , w_16253 );
not ( w_16253 , w_16254 );
and ( \6606_b0 , \6604_b0 , w_16255 );
and ( w_16254 ,  , w_16255 );
buf ( w_16253 , \6605_b1 );
not ( w_16253 , w_16256 );
not (  , w_16257 );
and ( w_16256 , w_16257 , \6605_b0 );
or ( \6607_b1 , \6606_b1 , w_16258 );
xor ( \6607_b0 , \6606_b0 , w_16260 );
not ( w_16260 , w_16261 );
and ( w_16261 , w_16258 , w_16259 );
buf ( w_16258 , \5923_b1 );
not ( w_16258 , w_16262 );
not ( w_16259 , w_16263 );
and ( w_16262 , w_16263 , \5923_b0 );
or ( \6608_b1 , \6603_b1 , \6607_b1 );
xor ( \6608_b0 , \6603_b0 , w_16264 );
not ( w_16264 , w_16265 );
and ( w_16265 , \6607_b1 , \6607_b0 );
or ( \6609_b1 , \5881_b1 , \5935_b1 );
not ( \5935_b1 , w_16266 );
and ( \6609_b0 , \5881_b0 , w_16267 );
and ( w_16266 , w_16267 , \5935_b0 );
or ( \6610_b1 , \5893_b1 , \5933_b1 );
not ( \5933_b1 , w_16268 );
and ( \6610_b0 , \5893_b0 , w_16269 );
and ( w_16268 , w_16269 , \5933_b0 );
or ( \6611_b1 , \6609_b1 , w_16271 );
not ( w_16271 , w_16272 );
and ( \6611_b0 , \6609_b0 , w_16273 );
and ( w_16272 ,  , w_16273 );
buf ( w_16271 , \6610_b1 );
not ( w_16271 , w_16274 );
not (  , w_16275 );
and ( w_16274 , w_16275 , \6610_b0 );
or ( \6612_b1 , \6611_b1 , w_16276 );
xor ( \6612_b0 , \6611_b0 , w_16278 );
not ( w_16278 , w_16279 );
and ( w_16279 , w_16276 , w_16277 );
buf ( w_16276 , \5942_b1 );
not ( w_16276 , w_16280 );
not ( w_16277 , w_16281 );
and ( w_16280 , w_16281 , \5942_b0 );
or ( \6613_b1 , \6608_b1 , \6612_b1 );
xor ( \6613_b0 , \6608_b0 , w_16282 );
not ( w_16282 , w_16283 );
and ( w_16283 , \6612_b1 , \6612_b0 );
or ( \6614_b1 , \6599_b1 , \6613_b1 );
xor ( \6614_b0 , \6599_b0 , w_16284 );
not ( w_16284 , w_16285 );
and ( w_16285 , \6613_b1 , \6613_b0 );
or ( \6615_b1 , \5780_b1 , \5829_b1 );
not ( \5829_b1 , w_16286 );
and ( \6615_b0 , \5780_b0 , w_16287 );
and ( w_16286 , w_16287 , \5829_b0 );
or ( \6616_b1 , \5792_b1 , \5827_b1 );
not ( \5827_b1 , w_16288 );
and ( \6616_b0 , \5792_b0 , w_16289 );
and ( w_16288 , w_16289 , \5827_b0 );
or ( \6617_b1 , \6615_b1 , w_16291 );
not ( w_16291 , w_16292 );
and ( \6617_b0 , \6615_b0 , w_16293 );
and ( w_16292 ,  , w_16293 );
buf ( w_16291 , \6616_b1 );
not ( w_16291 , w_16294 );
not (  , w_16295 );
and ( w_16294 , w_16295 , \6616_b0 );
or ( \6618_b1 , \6617_b1 , w_16296 );
xor ( \6618_b0 , \6617_b0 , w_16298 );
not ( w_16298 , w_16299 );
and ( w_16299 , w_16296 , w_16297 );
buf ( w_16296 , \5836_b1 );
not ( w_16296 , w_16300 );
not ( w_16297 , w_16301 );
and ( w_16300 , w_16301 , \5836_b0 );
or ( \6619_b1 , \5799_b1 , \5852_b1 );
not ( \5852_b1 , w_16302 );
and ( \6619_b0 , \5799_b0 , w_16303 );
and ( w_16302 , w_16303 , \5852_b0 );
or ( \6620_b1 , \5811_b1 , \5850_b1 );
not ( \5850_b1 , w_16304 );
and ( \6620_b0 , \5811_b0 , w_16305 );
and ( w_16304 , w_16305 , \5850_b0 );
or ( \6621_b1 , \6619_b1 , w_16307 );
not ( w_16307 , w_16308 );
and ( \6621_b0 , \6619_b0 , w_16309 );
and ( w_16308 ,  , w_16309 );
buf ( w_16307 , \6620_b1 );
not ( w_16307 , w_16310 );
not (  , w_16311 );
and ( w_16310 , w_16311 , \6620_b0 );
or ( \6622_b1 , \6621_b1 , w_16312 );
xor ( \6622_b0 , \6621_b0 , w_16314 );
not ( w_16314 , w_16315 );
and ( w_16315 , w_16312 , w_16313 );
buf ( w_16312 , \5859_b1 );
not ( w_16312 , w_16316 );
not ( w_16313 , w_16317 );
and ( w_16316 , w_16317 , \5859_b0 );
or ( \6623_b1 , \6618_b1 , \6622_b1 );
xor ( \6623_b0 , \6618_b0 , w_16318 );
not ( w_16318 , w_16319 );
and ( w_16319 , \6622_b1 , \6622_b0 );
or ( \6624_b1 , \5819_b1 , \5871_b1 );
not ( \5871_b1 , w_16320 );
and ( \6624_b0 , \5819_b0 , w_16321 );
and ( w_16320 , w_16321 , \5871_b0 );
or ( \6625_b1 , \5831_b1 , \5869_b1 );
not ( \5869_b1 , w_16322 );
and ( \6625_b0 , \5831_b0 , w_16323 );
and ( w_16322 , w_16323 , \5869_b0 );
or ( \6626_b1 , \6624_b1 , w_16325 );
not ( w_16325 , w_16326 );
and ( \6626_b0 , \6624_b0 , w_16327 );
and ( w_16326 ,  , w_16327 );
buf ( w_16325 , \6625_b1 );
not ( w_16325 , w_16328 );
not (  , w_16329 );
and ( w_16328 , w_16329 , \6625_b0 );
or ( \6627_b1 , \6626_b1 , w_16330 );
xor ( \6627_b0 , \6626_b0 , w_16332 );
not ( w_16332 , w_16333 );
and ( w_16333 , w_16330 , w_16331 );
buf ( w_16330 , \5878_b1 );
not ( w_16330 , w_16334 );
not ( w_16331 , w_16335 );
and ( w_16334 , w_16335 , \5878_b0 );
or ( \6628_b1 , \6623_b1 , \6627_b1 );
xor ( \6628_b0 , \6623_b0 , w_16336 );
not ( w_16336 , w_16337 );
and ( w_16337 , \6627_b1 , \6627_b0 );
or ( \6629_b1 , \6614_b1 , \6628_b1 );
xor ( \6629_b0 , \6614_b0 , w_16338 );
not ( w_16338 , w_16339 );
and ( w_16339 , \6628_b1 , \6628_b0 );
or ( \6630_b1 , \6585_b1 , \6629_b1 );
xor ( \6630_b0 , \6585_b0 , w_16340 );
not ( w_16340 , w_16341 );
and ( w_16341 , \6629_b1 , \6629_b0 );
or ( \6631_b1 , \6571_b1 , \6630_b1 );
xor ( \6631_b0 , \6571_b0 , w_16342 );
not ( w_16342 , w_16343 );
and ( w_16343 , \6630_b1 , \6630_b0 );
or ( \6632_b1 , \6363_b1 , \6367_b1 );
not ( \6367_b1 , w_16344 );
and ( \6632_b0 , \6363_b0 , w_16345 );
and ( w_16344 , w_16345 , \6367_b0 );
or ( \6633_b1 , \6367_b1 , \6372_b1 );
not ( \6372_b1 , w_16346 );
and ( \6633_b0 , \6367_b0 , w_16347 );
and ( w_16346 , w_16347 , \6372_b0 );
or ( \6634_b1 , \6363_b1 , \6372_b1 );
not ( \6372_b1 , w_16348 );
and ( \6634_b0 , \6363_b0 , w_16349 );
and ( w_16348 , w_16349 , \6372_b0 );
or ( \6636_b1 , \6349_b1 , \6353_b1 );
not ( \6353_b1 , w_16350 );
and ( \6636_b0 , \6349_b0 , w_16351 );
and ( w_16350 , w_16351 , \6353_b0 );
or ( \6637_b1 , \6353_b1 , \6358_b1 );
not ( \6358_b1 , w_16352 );
and ( \6637_b0 , \6353_b0 , w_16353 );
and ( w_16352 , w_16353 , \6358_b0 );
or ( \6638_b1 , \6349_b1 , \6358_b1 );
not ( \6358_b1 , w_16354 );
and ( \6638_b0 , \6349_b0 , w_16355 );
and ( w_16354 , w_16355 , \6358_b0 );
or ( \6640_b1 , \6635_b1 , \6639_b1 );
xor ( \6640_b0 , \6635_b0 , w_16356 );
not ( w_16356 , w_16357 );
and ( w_16357 , \6639_b1 , \6639_b0 );
or ( \6641_b1 , \6432_b1 , \6446_b1 );
not ( \6446_b1 , w_16358 );
and ( \6641_b0 , \6432_b0 , w_16359 );
and ( w_16358 , w_16359 , \6446_b0 );
or ( \6642_b1 , \6446_b1 , \6461_b1 );
not ( \6461_b1 , w_16360 );
and ( \6642_b0 , \6446_b0 , w_16361 );
and ( w_16360 , w_16361 , \6461_b0 );
or ( \6643_b1 , \6432_b1 , \6461_b1 );
not ( \6461_b1 , w_16362 );
and ( \6643_b0 , \6432_b0 , w_16363 );
and ( w_16362 , w_16363 , \6461_b0 );
or ( \6645_b1 , \6640_b1 , \6644_b1 );
xor ( \6645_b0 , \6640_b0 , w_16364 );
not ( w_16364 , w_16365 );
and ( w_16365 , \6644_b1 , \6644_b0 );
or ( \6646_b1 , \6631_b1 , \6645_b1 );
xor ( \6646_b0 , \6631_b0 , w_16366 );
not ( w_16366 , w_16367 );
and ( w_16367 , \6645_b1 , \6645_b0 );
or ( \6647_b1 , \6478_b1 , \6646_b1 );
not ( \6646_b1 , w_16368 );
and ( \6647_b0 , \6478_b0 , w_16369 );
and ( w_16368 , w_16369 , \6646_b0 );
or ( \6648_b1 , \6345_b1 , \6646_b1 );
not ( \6646_b1 , w_16370 );
and ( \6648_b0 , \6345_b0 , w_16371 );
and ( w_16370 , w_16371 , \6646_b0 );
or ( \6650_b1 , \6635_b1 , \6639_b1 );
not ( \6639_b1 , w_16372 );
and ( \6650_b0 , \6635_b0 , w_16373 );
and ( w_16372 , w_16373 , \6639_b0 );
or ( \6651_b1 , \6639_b1 , \6644_b1 );
not ( \6644_b1 , w_16374 );
and ( \6651_b0 , \6639_b0 , w_16375 );
and ( w_16374 , w_16375 , \6644_b0 );
or ( \6652_b1 , \6635_b1 , \6644_b1 );
not ( \6644_b1 , w_16376 );
and ( \6652_b0 , \6635_b0 , w_16377 );
and ( w_16376 , w_16377 , \6644_b0 );
or ( \6654_b1 , \6575_b1 , \6584_b1 );
not ( \6584_b1 , w_16378 );
and ( \6654_b0 , \6575_b0 , w_16379 );
and ( w_16378 , w_16379 , \6584_b0 );
or ( \6655_b1 , \6584_b1 , \6629_b1 );
not ( \6629_b1 , w_16380 );
and ( \6655_b0 , \6584_b0 , w_16381 );
and ( w_16380 , w_16381 , \6629_b0 );
or ( \6656_b1 , \6575_b1 , \6629_b1 );
not ( \6629_b1 , w_16382 );
and ( \6656_b0 , \6575_b0 , w_16383 );
and ( w_16382 , w_16383 , \6629_b0 );
or ( \6658_b1 , \6653_b1 , \6657_b1 );
xor ( \6658_b0 , \6653_b0 , w_16384 );
not ( w_16384 , w_16385 );
and ( w_16385 , \6657_b1 , \6657_b0 );
or ( \6659_b1 , \6544_b1 , \6555_b1 );
not ( \6555_b1 , w_16386 );
and ( \6659_b0 , \6544_b0 , w_16387 );
and ( w_16386 , w_16387 , \6555_b0 );
or ( \6660_b1 , \6555_b1 , \6570_b1 );
not ( \6570_b1 , w_16388 );
and ( \6660_b0 , \6555_b0 , w_16389 );
and ( w_16388 , w_16389 , \6570_b0 );
or ( \6661_b1 , \6544_b1 , \6570_b1 );
not ( \6570_b1 , w_16390 );
and ( \6661_b0 , \6544_b0 , w_16391 );
and ( w_16390 , w_16391 , \6570_b0 );
or ( \6663_b1 , \6658_b1 , \6662_b1 );
xor ( \6663_b0 , \6658_b0 , w_16392 );
not ( w_16392 , w_16393 );
and ( w_16393 , \6662_b1 , \6662_b0 );
or ( \6664_b1 , \6649_b1 , \6663_b1 );
xor ( \6664_b0 , \6649_b0 , w_16394 );
not ( w_16394 , w_16395 );
and ( w_16395 , \6663_b1 , \6663_b0 );
or ( \6665_b1 , \6468_b1 , \6472_b1 );
not ( \6472_b1 , w_16396 );
and ( \6665_b0 , \6468_b0 , w_16397 );
and ( w_16396 , w_16397 , \6472_b0 );
or ( \6666_b1 , \6472_b1 , \6474_b1 );
not ( \6474_b1 , w_16398 );
and ( \6666_b0 , \6472_b0 , w_16399 );
and ( w_16398 , w_16399 , \6474_b0 );
or ( \6667_b1 , \6468_b1 , \6474_b1 );
not ( \6474_b1 , w_16400 );
and ( \6667_b0 , \6468_b0 , w_16401 );
and ( w_16400 , w_16401 , \6474_b0 );
or ( \6669_b1 , \6378_b1 , \6419_b1 );
not ( \6419_b1 , w_16402 );
and ( \6669_b0 , \6378_b0 , w_16403 );
and ( w_16402 , w_16403 , \6419_b0 );
or ( \6670_b1 , \6419_b1 , \6462_b1 );
not ( \6462_b1 , w_16404 );
and ( \6670_b0 , \6419_b0 , w_16405 );
and ( w_16404 , w_16405 , \6462_b0 );
or ( \6671_b1 , \6378_b1 , \6462_b1 );
not ( \6462_b1 , w_16406 );
and ( \6671_b0 , \6378_b0 , w_16407 );
and ( w_16406 , w_16407 , \6462_b0 );
or ( \6673_b1 , \6668_b1 , \6672_b1 );
not ( \6672_b1 , w_16408 );
and ( \6673_b0 , \6668_b0 , w_16409 );
and ( w_16408 , w_16409 , \6672_b0 );
or ( \6674_b1 , \6359_b1 , \6373_b1 );
not ( \6373_b1 , w_16410 );
and ( \6674_b0 , \6359_b0 , w_16411 );
and ( w_16410 , w_16411 , \6373_b0 );
or ( \6675_b1 , \6672_b1 , \6674_b1 );
not ( \6674_b1 , w_16412 );
and ( \6675_b0 , \6672_b0 , w_16413 );
and ( w_16412 , w_16413 , \6674_b0 );
or ( \6676_b1 , \6668_b1 , \6674_b1 );
not ( \6674_b1 , w_16414 );
and ( \6676_b0 , \6668_b0 , w_16415 );
and ( w_16414 , w_16415 , \6674_b0 );
or ( \6678_b1 , \6571_b1 , \6630_b1 );
not ( \6630_b1 , w_16416 );
and ( \6678_b0 , \6571_b0 , w_16417 );
and ( w_16416 , w_16417 , \6630_b0 );
or ( \6679_b1 , \6630_b1 , \6645_b1 );
not ( \6645_b1 , w_16418 );
and ( \6679_b0 , \6630_b0 , w_16419 );
and ( w_16418 , w_16419 , \6645_b0 );
or ( \6680_b1 , \6571_b1 , \6645_b1 );
not ( \6645_b1 , w_16420 );
and ( \6680_b0 , \6571_b0 , w_16421 );
and ( w_16420 , w_16421 , \6645_b0 );
or ( \6682_b1 , \6677_b1 , \6681_b1 );
xor ( \6682_b0 , \6677_b0 , w_16422 );
not ( w_16422 , w_16423 );
and ( w_16423 , \6681_b1 , \6681_b0 );
or ( \6683_b1 , \6589_b1 , \6593_b1 );
not ( \6593_b1 , w_16424 );
and ( \6683_b0 , \6589_b0 , w_16425 );
and ( w_16424 , w_16425 , \6593_b0 );
or ( \6684_b1 , \6593_b1 , \6598_b1 );
not ( \6598_b1 , w_16426 );
and ( \6684_b0 , \6593_b0 , w_16427 );
and ( w_16426 , w_16427 , \6598_b0 );
or ( \6685_b1 , \6589_b1 , \6598_b1 );
not ( \6598_b1 , w_16428 );
and ( \6685_b0 , \6589_b0 , w_16429 );
and ( w_16428 , w_16429 , \6598_b0 );
or ( \6687_b1 , \6533_b1 , \6537_b1 );
not ( \6537_b1 , w_16430 );
and ( \6687_b0 , \6533_b0 , w_16431 );
and ( w_16430 , w_16431 , \6537_b0 );
or ( \6688_b1 , \6537_b1 , \6542_b1 );
not ( \6542_b1 , w_16432 );
and ( \6688_b0 , \6537_b0 , w_16433 );
and ( w_16432 , w_16433 , \6542_b0 );
or ( \6689_b1 , \6533_b1 , \6542_b1 );
not ( \6542_b1 , w_16434 );
and ( \6689_b0 , \6533_b0 , w_16435 );
and ( w_16434 , w_16435 , \6542_b0 );
or ( \6691_b1 , \6686_b1 , \6690_b1 );
xor ( \6691_b0 , \6686_b0 , w_16436 );
not ( w_16436 , w_16437 );
and ( w_16437 , \6690_b1 , \6690_b0 );
or ( \6692_b1 , \6483_b1 , \6487_b1 );
not ( \6487_b1 , w_16438 );
and ( \6692_b0 , \6483_b0 , w_16439 );
and ( w_16438 , w_16439 , \6487_b0 );
or ( \6693_b1 , \6487_b1 , \6528_b1 );
not ( \6528_b1 , w_16440 );
and ( \6693_b0 , \6487_b0 , w_16441 );
and ( w_16440 , w_16441 , \6528_b0 );
or ( \6694_b1 , \6483_b1 , \6528_b1 );
not ( \6528_b1 , w_16442 );
and ( \6694_b0 , \6483_b0 , w_16443 );
and ( w_16442 , w_16443 , \6528_b0 );
or ( \6696_b1 , \6691_b1 , \6695_b1 );
xor ( \6696_b0 , \6691_b0 , w_16444 );
not ( w_16444 , w_16445 );
and ( w_16445 , \6695_b1 , \6695_b0 );
or ( \6697_b1 , \6527_b1 , \6578_b1 );
not ( \6578_b1 , w_16446 );
and ( \6697_b0 , \6527_b0 , w_16447 );
and ( w_16446 , w_16447 , \6578_b0 );
or ( \6698_b1 , \6578_b1 , \6583_b1 );
not ( \6583_b1 , w_16448 );
and ( \6698_b0 , \6578_b0 , w_16449 );
and ( w_16448 , w_16449 , \6583_b0 );
or ( \6699_b1 , \6527_b1 , \6583_b1 );
not ( \6583_b1 , w_16450 );
and ( \6699_b0 , \6527_b0 , w_16451 );
and ( w_16450 , w_16451 , \6583_b0 );
or ( \6701_b1 , \6618_b1 , \6622_b1 );
not ( \6622_b1 , w_16452 );
and ( \6701_b0 , \6618_b0 , w_16453 );
and ( w_16452 , w_16453 , \6622_b0 );
or ( \6702_b1 , \6622_b1 , \6627_b1 );
not ( \6627_b1 , w_16454 );
and ( \6702_b0 , \6622_b0 , w_16455 );
and ( w_16454 , w_16455 , \6627_b0 );
or ( \6703_b1 , \6618_b1 , \6627_b1 );
not ( \6627_b1 , w_16456 );
and ( \6703_b0 , \6618_b0 , w_16457 );
and ( w_16456 , w_16457 , \6627_b0 );
or ( \6705_b1 , \6700_b1 , \6704_b1 );
xor ( \6705_b0 , \6700_b0 , w_16458 );
not ( w_16458 , w_16459 );
and ( w_16459 , \6704_b1 , \6704_b0 );
or ( \6706_b1 , \6603_b1 , \6607_b1 );
not ( \6607_b1 , w_16460 );
and ( \6706_b0 , \6603_b0 , w_16461 );
and ( w_16460 , w_16461 , \6607_b0 );
or ( \6707_b1 , \6607_b1 , \6612_b1 );
not ( \6612_b1 , w_16462 );
and ( \6707_b0 , \6607_b0 , w_16463 );
and ( w_16462 , w_16463 , \6612_b0 );
or ( \6708_b1 , \6603_b1 , \6612_b1 );
not ( \6612_b1 , w_16464 );
and ( \6708_b0 , \6603_b0 , w_16465 );
and ( w_16464 , w_16465 , \6612_b0 );
or ( \6710_b1 , \6705_b1 , \6709_b1 );
xor ( \6710_b0 , \6705_b0 , w_16466 );
not ( w_16466 , w_16467 );
and ( w_16467 , \6709_b1 , \6709_b0 );
or ( \6711_b1 , \6696_b1 , \6710_b1 );
xor ( \6711_b0 , \6696_b0 , w_16468 );
not ( w_16468 , w_16469 );
and ( w_16469 , \6710_b1 , \6710_b0 );
or ( \6712_b1 , \6599_b1 , \6613_b1 );
not ( \6613_b1 , w_16470 );
and ( \6712_b0 , \6599_b0 , w_16471 );
and ( w_16470 , w_16471 , \6613_b0 );
or ( \6713_b1 , \6613_b1 , \6628_b1 );
not ( \6628_b1 , w_16472 );
and ( \6713_b0 , \6613_b0 , w_16473 );
and ( w_16472 , w_16473 , \6628_b0 );
or ( \6714_b1 , \6599_b1 , \6628_b1 );
not ( \6628_b1 , w_16474 );
and ( \6714_b0 , \6599_b0 , w_16475 );
and ( w_16474 , w_16475 , \6628_b0 );
or ( \6716_b1 , \5873_b1 , \5916_b1 );
not ( \5916_b1 , w_16476 );
and ( \6716_b0 , \5873_b0 , w_16477 );
and ( w_16476 , w_16477 , \5916_b0 );
or ( \6717_b1 , \5842_b1 , \5914_b1 );
not ( \5914_b1 , w_16478 );
and ( \6717_b0 , \5842_b0 , w_16479 );
and ( w_16478 , w_16479 , \5914_b0 );
or ( \6718_b1 , \6716_b1 , w_16481 );
not ( w_16481 , w_16482 );
and ( \6718_b0 , \6716_b0 , w_16483 );
and ( w_16482 ,  , w_16483 );
buf ( w_16481 , \6717_b1 );
not ( w_16481 , w_16484 );
not (  , w_16485 );
and ( w_16484 , w_16485 , \6717_b0 );
or ( \6719_b1 , \6718_b1 , w_16486 );
xor ( \6719_b0 , \6718_b0 , w_16488 );
not ( w_16488 , w_16489 );
and ( w_16489 , w_16486 , w_16487 );
buf ( w_16486 , \5923_b1 );
not ( w_16486 , w_16490 );
not ( w_16487 , w_16491 );
and ( w_16490 , w_16491 , \5923_b0 );
or ( \6720_b1 , \5893_b1 , \5935_b1 );
not ( \5935_b1 , w_16492 );
and ( \6720_b0 , \5893_b0 , w_16493 );
and ( w_16492 , w_16493 , \5935_b0 );
or ( \6721_b1 , \5861_b1 , \5933_b1 );
not ( \5933_b1 , w_16494 );
and ( \6721_b0 , \5861_b0 , w_16495 );
and ( w_16494 , w_16495 , \5933_b0 );
or ( \6722_b1 , \6720_b1 , w_16497 );
not ( w_16497 , w_16498 );
and ( \6722_b0 , \6720_b0 , w_16499 );
and ( w_16498 ,  , w_16499 );
buf ( w_16497 , \6721_b1 );
not ( w_16497 , w_16500 );
not (  , w_16501 );
and ( w_16500 , w_16501 , \6721_b0 );
or ( \6723_b1 , \6722_b1 , w_16502 );
xor ( \6723_b0 , \6722_b0 , w_16504 );
not ( w_16504 , w_16505 );
and ( w_16505 , w_16502 , w_16503 );
buf ( w_16502 , \5942_b1 );
not ( w_16502 , w_16506 );
not ( w_16503 , w_16507 );
and ( w_16506 , w_16507 , \5942_b0 );
or ( \6724_b1 , \6719_b1 , \6723_b1 );
xor ( \6724_b0 , \6719_b0 , w_16508 );
not ( w_16508 , w_16509 );
and ( w_16509 , \6723_b1 , \6723_b0 );
or ( \6725_b1 , \5918_b1 , \5955_b1 );
not ( \5955_b1 , w_16510 );
and ( \6725_b0 , \5918_b0 , w_16511 );
and ( w_16510 , w_16511 , \5955_b0 );
or ( \6726_b1 , \5881_b1 , \5953_b1 );
not ( \5953_b1 , w_16512 );
and ( \6726_b0 , \5881_b0 , w_16513 );
and ( w_16512 , w_16513 , \5953_b0 );
or ( \6727_b1 , \6725_b1 , w_16515 );
not ( w_16515 , w_16516 );
and ( \6727_b0 , \6725_b0 , w_16517 );
and ( w_16516 ,  , w_16517 );
buf ( w_16515 , \6726_b1 );
not ( w_16515 , w_16518 );
not (  , w_16519 );
and ( w_16518 , w_16519 , \6726_b0 );
or ( \6728_b1 , \6727_b1 , w_16520 );
xor ( \6728_b0 , \6727_b0 , w_16522 );
not ( w_16522 , w_16523 );
and ( w_16523 , w_16520 , w_16521 );
buf ( w_16520 , \5962_b1 );
not ( w_16520 , w_16524 );
not ( w_16521 , w_16525 );
and ( w_16524 , w_16525 , \5962_b0 );
or ( \6729_b1 , \6724_b1 , \6728_b1 );
xor ( \6729_b0 , \6724_b0 , w_16526 );
not ( w_16526 , w_16527 );
and ( w_16527 , \6728_b1 , \6728_b0 );
or ( \6730_b1 , \5811_b1 , \5852_b1 );
not ( \5852_b1 , w_16528 );
and ( \6730_b0 , \5811_b0 , w_16529 );
and ( w_16528 , w_16529 , \5852_b0 );
or ( \6731_b1 , \5780_b1 , \5850_b1 );
not ( \5850_b1 , w_16530 );
and ( \6731_b0 , \5780_b0 , w_16531 );
and ( w_16530 , w_16531 , \5850_b0 );
or ( \6732_b1 , \6730_b1 , w_16533 );
not ( w_16533 , w_16534 );
and ( \6732_b0 , \6730_b0 , w_16535 );
and ( w_16534 ,  , w_16535 );
buf ( w_16533 , \6731_b1 );
not ( w_16533 , w_16536 );
not (  , w_16537 );
and ( w_16536 , w_16537 , \6731_b0 );
or ( \6733_b1 , \6732_b1 , w_16538 );
xor ( \6733_b0 , \6732_b0 , w_16540 );
not ( w_16540 , w_16541 );
and ( w_16541 , w_16538 , w_16539 );
buf ( w_16538 , \5859_b1 );
not ( w_16538 , w_16542 );
not ( w_16539 , w_16543 );
and ( w_16542 , w_16543 , \5859_b0 );
or ( \6734_b1 , \5831_b1 , \5871_b1 );
not ( \5871_b1 , w_16544 );
and ( \6734_b0 , \5831_b0 , w_16545 );
and ( w_16544 , w_16545 , \5871_b0 );
or ( \6735_b1 , \5799_b1 , \5869_b1 );
not ( \5869_b1 , w_16546 );
and ( \6735_b0 , \5799_b0 , w_16547 );
and ( w_16546 , w_16547 , \5869_b0 );
or ( \6736_b1 , \6734_b1 , w_16549 );
not ( w_16549 , w_16550 );
and ( \6736_b0 , \6734_b0 , w_16551 );
and ( w_16550 ,  , w_16551 );
buf ( w_16549 , \6735_b1 );
not ( w_16549 , w_16552 );
not (  , w_16553 );
and ( w_16552 , w_16553 , \6735_b0 );
or ( \6737_b1 , \6736_b1 , w_16554 );
xor ( \6737_b0 , \6736_b0 , w_16556 );
not ( w_16556 , w_16557 );
and ( w_16557 , w_16554 , w_16555 );
buf ( w_16554 , \5878_b1 );
not ( w_16554 , w_16558 );
not ( w_16555 , w_16559 );
and ( w_16558 , w_16559 , \5878_b0 );
or ( \6738_b1 , \6733_b1 , \6737_b1 );
xor ( \6738_b0 , \6733_b0 , w_16560 );
not ( w_16560 , w_16561 );
and ( w_16561 , \6737_b1 , \6737_b0 );
or ( \6739_b1 , \5854_b1 , \5891_b1 );
not ( \5891_b1 , w_16562 );
and ( \6739_b0 , \5854_b0 , w_16563 );
and ( w_16562 , w_16563 , \5891_b0 );
or ( \6740_b1 , \5819_b1 , \5889_b1 );
not ( \5889_b1 , w_16564 );
and ( \6740_b0 , \5819_b0 , w_16565 );
and ( w_16564 , w_16565 , \5889_b0 );
or ( \6741_b1 , \6739_b1 , w_16567 );
not ( w_16567 , w_16568 );
and ( \6741_b0 , \6739_b0 , w_16569 );
and ( w_16568 ,  , w_16569 );
buf ( w_16567 , \6740_b1 );
not ( w_16567 , w_16570 );
not (  , w_16571 );
and ( w_16570 , w_16571 , \6740_b0 );
or ( \6742_b1 , \6741_b1 , w_16572 );
xor ( \6742_b0 , \6741_b0 , w_16574 );
not ( w_16574 , w_16575 );
and ( w_16575 , w_16572 , w_16573 );
buf ( w_16572 , \5898_b1 );
not ( w_16572 , w_16576 );
not ( w_16573 , w_16577 );
and ( w_16576 , w_16577 , \5898_b0 );
or ( \6743_b1 , \6738_b1 , \6742_b1 );
xor ( \6743_b0 , \6738_b0 , w_16578 );
not ( w_16578 , w_16579 );
and ( w_16579 , \6742_b1 , \6742_b0 );
or ( \6744_b1 , \6729_b1 , \6743_b1 );
xor ( \6744_b0 , \6729_b0 , w_16580 );
not ( w_16580 , w_16581 );
and ( w_16581 , \6743_b1 , \6743_b0 );
buf ( \6745_b1 , \5797_b1 );
not ( \6745_b1 , w_16582 );
not ( \6745_b0 , w_16583 );
and ( w_16582 , w_16583 , \5797_b0 );
or ( \6746_b1 , \5770_b1 , \5809_b1 );
not ( \5809_b1 , w_16584 );
and ( \6746_b0 , \5770_b0 , w_16585 );
and ( w_16584 , w_16585 , \5809_b0 );
or ( \6747_b1 , \5737_b1 , \5807_b1 );
not ( \5807_b1 , w_16586 );
and ( \6747_b0 , \5737_b0 , w_16587 );
and ( w_16586 , w_16587 , \5807_b0 );
or ( \6748_b1 , \6746_b1 , w_16589 );
not ( w_16589 , w_16590 );
and ( \6748_b0 , \6746_b0 , w_16591 );
and ( w_16590 ,  , w_16591 );
buf ( w_16589 , \6747_b1 );
not ( w_16589 , w_16592 );
not (  , w_16593 );
and ( w_16592 , w_16593 , \6747_b0 );
or ( \6749_b1 , \6748_b1 , w_16594 );
xor ( \6749_b0 , \6748_b0 , w_16596 );
not ( w_16596 , w_16597 );
and ( w_16597 , w_16594 , w_16595 );
buf ( w_16594 , \5816_b1 );
not ( w_16594 , w_16598 );
not ( w_16595 , w_16599 );
and ( w_16598 , w_16599 , \5816_b0 );
or ( \6750_b1 , \6745_b1 , \6749_b1 );
xor ( \6750_b0 , \6745_b0 , w_16600 );
not ( w_16600 , w_16601 );
and ( w_16601 , \6749_b1 , \6749_b0 );
or ( \6751_b1 , \5792_b1 , \5829_b1 );
not ( \5829_b1 , w_16602 );
and ( \6751_b0 , \5792_b0 , w_16603 );
and ( w_16602 , w_16603 , \5829_b0 );
or ( \6752_b1 , \5758_b1 , \5827_b1 );
not ( \5827_b1 , w_16604 );
and ( \6752_b0 , \5758_b0 , w_16605 );
and ( w_16604 , w_16605 , \5827_b0 );
or ( \6753_b1 , \6751_b1 , w_16607 );
not ( w_16607 , w_16608 );
and ( \6753_b0 , \6751_b0 , w_16609 );
and ( w_16608 ,  , w_16609 );
buf ( w_16607 , \6752_b1 );
not ( w_16607 , w_16610 );
not (  , w_16611 );
and ( w_16610 , w_16611 , \6752_b0 );
or ( \6754_b1 , \6753_b1 , w_16612 );
xor ( \6754_b0 , \6753_b0 , w_16614 );
not ( w_16614 , w_16615 );
and ( w_16615 , w_16612 , w_16613 );
buf ( w_16612 , \5836_b1 );
not ( w_16612 , w_16616 );
not ( w_16613 , w_16617 );
and ( w_16616 , w_16617 , \5836_b0 );
or ( \6755_b1 , \6750_b1 , \6754_b1 );
xor ( \6755_b0 , \6750_b0 , w_16618 );
not ( w_16618 , w_16619 );
and ( w_16619 , \6754_b1 , \6754_b0 );
or ( \6756_b1 , \6744_b1 , \6755_b1 );
xor ( \6756_b0 , \6744_b0 , w_16620 );
not ( w_16620 , w_16621 );
and ( w_16621 , \6755_b1 , \6755_b0 );
or ( \6757_b1 , \6715_b1 , \6756_b1 );
xor ( \6757_b0 , \6715_b0 , w_16622 );
not ( w_16622 , w_16623 );
and ( w_16623 , \6756_b1 , \6756_b0 );
or ( \6758_b1 , \6057_b1 , \6427_b1 );
not ( \6427_b1 , w_16624 );
and ( \6758_b0 , \6057_b0 , w_16625 );
and ( w_16624 , w_16625 , \6427_b0 );
or ( \6759_b1 , \6029_b1 , \6295_b1 );
not ( \6295_b1 , w_16626 );
and ( \6759_b0 , \6029_b0 , w_16627 );
and ( w_16626 , w_16627 , \6295_b0 );
or ( \6760_b1 , \6758_b1 , w_16629 );
not ( w_16629 , w_16630 );
and ( \6760_b0 , \6758_b0 , w_16631 );
and ( w_16630 ,  , w_16631 );
buf ( w_16629 , \6759_b1 );
not ( w_16629 , w_16632 );
not (  , w_16633 );
and ( w_16632 , w_16633 , \6759_b0 );
or ( \6761_b1 , \6760_b1 , w_16634 );
xor ( \6761_b0 , \6760_b0 , w_16636 );
not ( w_16636 , w_16637 );
and ( w_16637 , w_16634 , w_16635 );
buf ( w_16634 , \6227_b1 );
not ( w_16634 , w_16638 );
not ( w_16635 , w_16639 );
and ( w_16638 , w_16639 , \6227_b0 );
or ( \6762_b1 , \6524_b1 , \6509_b1 );
xor ( \6762_b0 , \6524_b0 , w_16640 );
not ( w_16640 , w_16641 );
and ( w_16641 , \6509_b1 , \6509_b0 );
buf ( \6763_b1 , \6510_b1 );
not ( \6763_b1 , w_16642 );
not ( \6763_b0 , w_16643 );
and ( w_16642 , w_16643 , \6510_b0 );
or ( \6764_b1 , \6762_b1 , \6763_b1 );
not ( \6763_b1 , w_16644 );
and ( \6764_b0 , \6762_b0 , w_16645 );
and ( w_16644 , w_16645 , \6763_b0 );
or ( \6765_b1 , \6065_b1 , \6764_b1 );
not ( \6764_b1 , w_16646 );
and ( \6765_b0 , \6065_b0 , w_16647 );
and ( w_16646 , w_16647 , \6764_b0 );
or ( \6766_b1 , \6048_b1 , \6510_b1 );
not ( \6510_b1 , w_16648 );
and ( \6766_b0 , \6048_b0 , w_16649 );
and ( w_16648 , w_16649 , \6510_b0 );
or ( \6767_b1 , \6765_b1 , w_16651 );
not ( w_16651 , w_16652 );
and ( \6767_b0 , \6765_b0 , w_16653 );
and ( w_16652 ,  , w_16653 );
buf ( w_16651 , \6766_b1 );
not ( w_16651 , w_16654 );
not (  , w_16655 );
and ( w_16654 , w_16655 , \6766_b0 );
or ( \6768_b1 , \6767_b1 , w_16656 );
xor ( \6768_b0 , \6767_b0 , w_16658 );
not ( w_16658 , w_16659 );
and ( w_16659 , w_16656 , w_16657 );
buf ( w_16656 , \6527_b1 );
not ( w_16656 , w_16660 );
not ( w_16657 , w_16661 );
and ( w_16660 , w_16661 , \6527_b0 );
or ( \6769_b1 , \6761_b1 , \6768_b1 );
xor ( \6769_b0 , \6761_b0 , w_16662 );
not ( w_16662 , w_16663 );
and ( w_16663 , \6768_b1 , \6768_b0 );
or ( \6770_b1 , \5998_b1 , \6039_b1 );
not ( \6039_b1 , w_16664 );
and ( \6770_b0 , \5998_b0 , w_16665 );
and ( w_16664 , w_16665 , \6039_b0 );
or ( \6771_b1 , \5967_b1 , \6037_b1 );
not ( \6037_b1 , w_16666 );
and ( \6771_b0 , \5967_b0 , w_16667 );
and ( w_16666 , w_16667 , \6037_b0 );
or ( \6772_b1 , \6770_b1 , w_16669 );
not ( w_16669 , w_16670 );
and ( \6772_b0 , \6770_b0 , w_16671 );
and ( w_16670 ,  , w_16671 );
buf ( w_16669 , \6771_b1 );
not ( w_16669 , w_16672 );
not (  , w_16673 );
and ( w_16672 , w_16673 , \6771_b0 );
or ( \6773_b1 , \6772_b1 , w_16674 );
xor ( \6773_b0 , \6772_b0 , w_16676 );
not ( w_16676 , w_16677 );
and ( w_16677 , w_16674 , w_16675 );
buf ( w_16674 , \6046_b1 );
not ( w_16674 , w_16678 );
not ( w_16675 , w_16679 );
and ( w_16678 , w_16679 , \6046_b0 );
or ( \6774_b1 , \6018_b1 , \6055_b1 );
not ( \6055_b1 , w_16680 );
and ( \6774_b0 , \6018_b0 , w_16681 );
and ( w_16680 , w_16681 , \6055_b0 );
or ( \6775_b1 , \5986_b1 , \6053_b1 );
not ( \6053_b1 , w_16682 );
and ( \6775_b0 , \5986_b0 , w_16683 );
and ( w_16682 , w_16683 , \6053_b0 );
or ( \6776_b1 , \6774_b1 , w_16685 );
not ( w_16685 , w_16686 );
and ( \6776_b0 , \6774_b0 , w_16687 );
and ( w_16686 ,  , w_16687 );
buf ( w_16685 , \6775_b1 );
not ( w_16685 , w_16688 );
not (  , w_16689 );
and ( w_16688 , w_16689 , \6775_b0 );
or ( \6777_b1 , \6776_b1 , w_16690 );
xor ( \6777_b0 , \6776_b0 , w_16692 );
not ( w_16692 , w_16693 );
and ( w_16693 , w_16690 , w_16691 );
buf ( w_16690 , \6062_b1 );
not ( w_16690 , w_16694 );
not ( w_16691 , w_16695 );
and ( w_16694 , w_16695 , \6062_b0 );
or ( \6778_b1 , \6773_b1 , \6777_b1 );
xor ( \6778_b0 , \6773_b0 , w_16696 );
not ( w_16696 , w_16697 );
and ( w_16697 , \6777_b1 , \6777_b0 );
or ( \6779_b1 , \6041_b1 , \6082_b1 );
not ( \6082_b1 , w_16698 );
and ( \6779_b0 , \6041_b0 , w_16699 );
and ( w_16698 , w_16699 , \6082_b0 );
or ( \6780_b1 , \6006_b1 , \6066_b1 );
not ( \6066_b1 , w_16700 );
and ( \6780_b0 , \6006_b0 , w_16701 );
and ( w_16700 , w_16701 , \6066_b0 );
or ( \6781_b1 , \6779_b1 , w_16703 );
not ( w_16703 , w_16704 );
and ( \6781_b0 , \6779_b0 , w_16705 );
and ( w_16704 ,  , w_16705 );
buf ( w_16703 , \6780_b1 );
not ( w_16703 , w_16706 );
not (  , w_16707 );
and ( w_16706 , w_16707 , \6780_b0 );
or ( \6782_b1 , \6781_b1 , w_16708 );
xor ( \6782_b0 , \6781_b0 , w_16710 );
not ( w_16710 , w_16711 );
and ( w_16711 , w_16708 , w_16709 );
buf ( w_16708 , \5736_b1 );
not ( w_16708 , w_16712 );
not ( w_16709 , w_16713 );
and ( w_16712 , w_16713 , \5736_b0 );
or ( \6783_b1 , \6778_b1 , \6782_b1 );
xor ( \6783_b0 , \6778_b0 , w_16714 );
not ( w_16714 , w_16715 );
and ( w_16715 , \6782_b1 , \6782_b0 );
or ( \6784_b1 , \6769_b1 , \6783_b1 );
xor ( \6784_b0 , \6769_b0 , w_16716 );
not ( w_16716 , w_16717 );
and ( w_16717 , \6783_b1 , \6783_b0 );
or ( \6785_b1 , \5937_b1 , \5977_b1 );
not ( \5977_b1 , w_16718 );
and ( \6785_b0 , \5937_b0 , w_16719 );
and ( w_16718 , w_16719 , \5977_b0 );
or ( \6786_b1 , \5906_b1 , \5975_b1 );
not ( \5975_b1 , w_16720 );
and ( \6786_b0 , \5906_b0 , w_16721 );
and ( w_16720 , w_16721 , \5975_b0 );
or ( \6787_b1 , \6785_b1 , w_16723 );
not ( w_16723 , w_16724 );
and ( \6787_b0 , \6785_b0 , w_16725 );
and ( w_16724 ,  , w_16725 );
buf ( w_16723 , \6786_b1 );
not ( w_16723 , w_16726 );
not (  , w_16727 );
and ( w_16726 , w_16727 , \6786_b0 );
or ( \6788_b1 , \6787_b1 , w_16728 );
xor ( \6788_b0 , \6787_b0 , w_16730 );
not ( w_16730 , w_16731 );
and ( w_16731 , w_16728 , w_16729 );
buf ( w_16728 , \5984_b1 );
not ( w_16728 , w_16732 );
not ( w_16729 , w_16733 );
and ( w_16732 , w_16733 , \5984_b0 );
or ( \6789_b1 , \5957_b1 , \5996_b1 );
not ( \5996_b1 , w_16734 );
and ( \6789_b0 , \5957_b0 , w_16735 );
and ( w_16734 , w_16735 , \5996_b0 );
or ( \6790_b1 , \5925_b1 , \5994_b1 );
not ( \5994_b1 , w_16736 );
and ( \6790_b0 , \5925_b0 , w_16737 );
and ( w_16736 , w_16737 , \5994_b0 );
or ( \6791_b1 , \6789_b1 , w_16739 );
not ( w_16739 , w_16740 );
and ( \6791_b0 , \6789_b0 , w_16741 );
and ( w_16740 ,  , w_16741 );
buf ( w_16739 , \6790_b1 );
not ( w_16739 , w_16742 );
not (  , w_16743 );
and ( w_16742 , w_16743 , \6790_b0 );
or ( \6792_b1 , \6791_b1 , w_16744 );
xor ( \6792_b0 , \6791_b0 , w_16746 );
not ( w_16746 , w_16747 );
and ( w_16747 , w_16744 , w_16745 );
buf ( w_16744 , \6003_b1 );
not ( w_16744 , w_16748 );
not ( w_16745 , w_16749 );
and ( w_16748 , w_16749 , \6003_b0 );
or ( \6793_b1 , \6788_b1 , \6792_b1 );
xor ( \6793_b0 , \6788_b0 , w_16750 );
not ( w_16750 , w_16751 );
and ( w_16751 , \6792_b1 , \6792_b0 );
or ( \6794_b1 , \5979_b1 , \6016_b1 );
not ( \6016_b1 , w_16752 );
and ( \6794_b0 , \5979_b0 , w_16753 );
and ( w_16752 , w_16753 , \6016_b0 );
or ( \6795_b1 , \5945_b1 , \6014_b1 );
not ( \6014_b1 , w_16754 );
and ( \6795_b0 , \5945_b0 , w_16755 );
and ( w_16754 , w_16755 , \6014_b0 );
or ( \6796_b1 , \6794_b1 , w_16757 );
not ( w_16757 , w_16758 );
and ( \6796_b0 , \6794_b0 , w_16759 );
and ( w_16758 ,  , w_16759 );
buf ( w_16757 , \6795_b1 );
not ( w_16757 , w_16760 );
not (  , w_16761 );
and ( w_16760 , w_16761 , \6795_b0 );
or ( \6797_b1 , \6796_b1 , w_16762 );
xor ( \6797_b0 , \6796_b0 , w_16764 );
not ( w_16764 , w_16765 );
and ( w_16765 , w_16762 , w_16763 );
buf ( w_16762 , \6023_b1 );
not ( w_16762 , w_16766 );
not ( w_16763 , w_16767 );
and ( w_16766 , w_16767 , \6023_b0 );
or ( \6798_b1 , \6793_b1 , \6797_b1 );
xor ( \6798_b0 , \6793_b0 , w_16768 );
not ( w_16768 , w_16769 );
and ( w_16769 , \6797_b1 , \6797_b0 );
or ( \6799_b1 , \6784_b1 , \6798_b1 );
xor ( \6799_b0 , \6784_b0 , w_16770 );
not ( w_16770 , w_16771 );
and ( w_16771 , \6798_b1 , \6798_b0 );
or ( \6800_b1 , \6757_b1 , \6799_b1 );
xor ( \6800_b0 , \6757_b0 , w_16772 );
not ( w_16772 , w_16773 );
and ( w_16773 , \6799_b1 , \6799_b0 );
or ( \6801_b1 , \6711_b1 , \6800_b1 );
xor ( \6801_b0 , \6711_b0 , w_16774 );
not ( w_16774 , w_16775 );
and ( w_16775 , \6800_b1 , \6800_b0 );
or ( \6802_b1 , \6560_b1 , \6564_b1 );
not ( \6564_b1 , w_16776 );
and ( \6802_b0 , \6560_b0 , w_16777 );
and ( w_16776 , w_16777 , \6564_b0 );
or ( \6803_b1 , \6564_b1 , \6569_b1 );
not ( \6569_b1 , w_16778 );
and ( \6803_b0 , \6564_b0 , w_16779 );
and ( w_16778 , w_16779 , \6569_b0 );
or ( \6804_b1 , \6560_b1 , \6569_b1 );
not ( \6569_b1 , w_16780 );
and ( \6804_b0 , \6560_b0 , w_16781 );
and ( w_16780 , w_16781 , \6569_b0 );
or ( \6806_b1 , \6548_b1 , \6552_b1 );
not ( \6552_b1 , w_16782 );
and ( \6806_b0 , \6548_b0 , w_16783 );
and ( w_16782 , w_16783 , \6552_b0 );
or ( \6807_b1 , \6552_b1 , \6554_b1 );
not ( \6554_b1 , w_16784 );
and ( \6807_b0 , \6552_b0 , w_16785 );
and ( w_16784 , w_16785 , \6554_b0 );
or ( \6808_b1 , \6548_b1 , \6554_b1 );
not ( \6554_b1 , w_16786 );
and ( \6808_b0 , \6548_b0 , w_16787 );
and ( w_16786 , w_16787 , \6554_b0 );
or ( \6810_b1 , \6805_b1 , \6809_b1 );
xor ( \6810_b0 , \6805_b0 , w_16788 );
not ( w_16788 , w_16789 );
and ( w_16789 , \6809_b1 , \6809_b0 );
or ( \6811_b1 , \6529_b1 , w_16790 );
or ( \6811_b0 , \6529_b0 , \6543_b0 );
not ( \6543_b0 , w_16791 );
and ( w_16791 , w_16790 , \6543_b1 );
or ( \6812_b1 , \6810_b1 , \6811_b1 );
xor ( \6812_b0 , \6810_b0 , w_16792 );
not ( w_16792 , w_16793 );
and ( w_16793 , \6811_b1 , \6811_b0 );
or ( \6813_b1 , \6801_b1 , \6812_b1 );
xor ( \6813_b0 , \6801_b0 , w_16794 );
not ( w_16794 , w_16795 );
and ( w_16795 , \6812_b1 , \6812_b0 );
or ( \6814_b1 , \6682_b1 , \6813_b1 );
xor ( \6814_b0 , \6682_b0 , w_16796 );
not ( w_16796 , w_16797 );
and ( w_16797 , \6813_b1 , \6813_b0 );
or ( \6815_b1 , \6664_b1 , \6814_b1 );
xor ( \6815_b0 , \6664_b0 , w_16798 );
not ( w_16798 , w_16799 );
and ( w_16799 , \6814_b1 , \6814_b0 );
or ( \6816_b1 , \4668_b1 , \5654_b1 );
xor ( \6816_b0 , \4668_b0 , w_16800 );
not ( w_16800 , w_16801 );
and ( w_16801 , \5654_b1 , \5654_b0 );
buf ( \6817_b1 , \6816_b1 );
buf ( \6817_b0 , \6816_b0 );
buf ( \6818_b1 , \6817_b1 );
buf ( \6818_b0 , \6817_b0 );
or ( \6819_b1 , \4760_b1 , \5652_b1 );
xor ( \6819_b0 , \4760_b0 , w_16802 );
not ( w_16802 , w_16803 );
and ( w_16803 , \5652_b1 , \5652_b0 );
buf ( \6820_b1 , \6819_b1 );
buf ( \6820_b0 , \6819_b0 );
buf ( \6821_b1 , \6820_b1 );
buf ( \6821_b0 , \6820_b0 );
or ( \6822_b1 , \6818_b1 , \6821_b1 );
not ( \6821_b1 , w_16804 );
and ( \6822_b0 , \6818_b0 , w_16805 );
and ( w_16804 , w_16805 , \6821_b0 );
buf ( \6823_b1 , \6822_b1 );
not ( \6823_b1 , w_16806 );
not ( \6823_b0 , w_16807 );
and ( w_16806 , w_16807 , \6822_b0 );
or ( \6824_b1 , \5747_b1 , \6823_b1 );
not ( \6823_b1 , w_16808 );
and ( \6824_b0 , \5747_b0 , w_16809 );
and ( w_16808 , w_16809 , \6823_b0 );
buf ( \6825_b1 , \6824_b1 );
not ( \6825_b1 , w_16810 );
not ( \6825_b0 , w_16811 );
and ( w_16810 , w_16811 , \6824_b0 );
or ( \6826_b1 , \5770_b1 , \5750_b1 );
not ( \5750_b1 , w_16812 );
and ( \6826_b0 , \5770_b0 , w_16813 );
and ( w_16812 , w_16813 , \5750_b0 );
or ( \6827_b1 , \5737_b1 , \5748_b1 );
not ( \5748_b1 , w_16814 );
and ( \6827_b0 , \5737_b0 , w_16815 );
and ( w_16814 , w_16815 , \5748_b0 );
or ( \6828_b1 , \6826_b1 , w_16817 );
not ( w_16817 , w_16818 );
and ( \6828_b0 , \6826_b0 , w_16819 );
and ( w_16818 ,  , w_16819 );
buf ( w_16817 , \6827_b1 );
not ( w_16817 , w_16820 );
not (  , w_16821 );
and ( w_16820 , w_16821 , \6827_b0 );
or ( \6829_b1 , \6828_b1 , w_16822 );
xor ( \6829_b0 , \6828_b0 , w_16824 );
not ( w_16824 , w_16825 );
and ( w_16825 , w_16822 , w_16823 );
buf ( w_16822 , \5755_b1 );
not ( w_16822 , w_16826 );
not ( w_16823 , w_16827 );
and ( w_16826 , w_16827 , \5755_b0 );
or ( \6830_b1 , \6825_b1 , \6829_b1 );
not ( \6829_b1 , w_16828 );
and ( \6830_b0 , \6825_b0 , w_16829 );
and ( w_16828 , w_16829 , \6829_b0 );
or ( \6831_b1 , \5792_b1 , \5768_b1 );
not ( \5768_b1 , w_16830 );
and ( \6831_b0 , \5792_b0 , w_16831 );
and ( w_16830 , w_16831 , \5768_b0 );
or ( \6832_b1 , \5758_b1 , \5766_b1 );
not ( \5766_b1 , w_16832 );
and ( \6832_b0 , \5758_b0 , w_16833 );
and ( w_16832 , w_16833 , \5766_b0 );
or ( \6833_b1 , \6831_b1 , w_16835 );
not ( w_16835 , w_16836 );
and ( \6833_b0 , \6831_b0 , w_16837 );
and ( w_16836 ,  , w_16837 );
buf ( w_16835 , \6832_b1 );
not ( w_16835 , w_16838 );
not (  , w_16839 );
and ( w_16838 , w_16839 , \6832_b0 );
or ( \6834_b1 , \6833_b1 , w_16840 );
xor ( \6834_b0 , \6833_b0 , w_16842 );
not ( w_16842 , w_16843 );
and ( w_16843 , w_16840 , w_16841 );
buf ( w_16840 , \5775_b1 );
not ( w_16840 , w_16844 );
not ( w_16841 , w_16845 );
and ( w_16844 , w_16845 , \5775_b0 );
or ( \6835_b1 , \6829_b1 , \6834_b1 );
not ( \6834_b1 , w_16846 );
and ( \6835_b0 , \6829_b0 , w_16847 );
and ( w_16846 , w_16847 , \6834_b0 );
or ( \6836_b1 , \6825_b1 , \6834_b1 );
not ( \6834_b1 , w_16848 );
and ( \6836_b0 , \6825_b0 , w_16849 );
and ( w_16848 , w_16849 , \6834_b0 );
or ( \6838_b1 , \5811_b1 , \5790_b1 );
not ( \5790_b1 , w_16850 );
and ( \6838_b0 , \5811_b0 , w_16851 );
and ( w_16850 , w_16851 , \5790_b0 );
or ( \6839_b1 , \5780_b1 , \5788_b1 );
not ( \5788_b1 , w_16852 );
and ( \6839_b0 , \5780_b0 , w_16853 );
and ( w_16852 , w_16853 , \5788_b0 );
or ( \6840_b1 , \6838_b1 , w_16855 );
not ( w_16855 , w_16856 );
and ( \6840_b0 , \6838_b0 , w_16857 );
and ( w_16856 ,  , w_16857 );
buf ( w_16855 , \6839_b1 );
not ( w_16855 , w_16858 );
not (  , w_16859 );
and ( w_16858 , w_16859 , \6839_b0 );
or ( \6841_b1 , \6840_b1 , w_16860 );
xor ( \6841_b0 , \6840_b0 , w_16862 );
not ( w_16862 , w_16863 );
and ( w_16863 , w_16860 , w_16861 );
buf ( w_16860 , \5797_b1 );
not ( w_16860 , w_16864 );
not ( w_16861 , w_16865 );
and ( w_16864 , w_16865 , \5797_b0 );
or ( \6842_b1 , \5831_b1 , \5809_b1 );
not ( \5809_b1 , w_16866 );
and ( \6842_b0 , \5831_b0 , w_16867 );
and ( w_16866 , w_16867 , \5809_b0 );
or ( \6843_b1 , \5799_b1 , \5807_b1 );
not ( \5807_b1 , w_16868 );
and ( \6843_b0 , \5799_b0 , w_16869 );
and ( w_16868 , w_16869 , \5807_b0 );
or ( \6844_b1 , \6842_b1 , w_16871 );
not ( w_16871 , w_16872 );
and ( \6844_b0 , \6842_b0 , w_16873 );
and ( w_16872 ,  , w_16873 );
buf ( w_16871 , \6843_b1 );
not ( w_16871 , w_16874 );
not (  , w_16875 );
and ( w_16874 , w_16875 , \6843_b0 );
or ( \6845_b1 , \6844_b1 , w_16876 );
xor ( \6845_b0 , \6844_b0 , w_16878 );
not ( w_16878 , w_16879 );
and ( w_16879 , w_16876 , w_16877 );
buf ( w_16876 , \5816_b1 );
not ( w_16876 , w_16880 );
not ( w_16877 , w_16881 );
and ( w_16880 , w_16881 , \5816_b0 );
or ( \6846_b1 , \6841_b1 , \6845_b1 );
not ( \6845_b1 , w_16882 );
and ( \6846_b0 , \6841_b0 , w_16883 );
and ( w_16882 , w_16883 , \6845_b0 );
or ( \6847_b1 , \5854_b1 , \5829_b1 );
not ( \5829_b1 , w_16884 );
and ( \6847_b0 , \5854_b0 , w_16885 );
and ( w_16884 , w_16885 , \5829_b0 );
or ( \6848_b1 , \5819_b1 , \5827_b1 );
not ( \5827_b1 , w_16886 );
and ( \6848_b0 , \5819_b0 , w_16887 );
and ( w_16886 , w_16887 , \5827_b0 );
or ( \6849_b1 , \6847_b1 , w_16889 );
not ( w_16889 , w_16890 );
and ( \6849_b0 , \6847_b0 , w_16891 );
and ( w_16890 ,  , w_16891 );
buf ( w_16889 , \6848_b1 );
not ( w_16889 , w_16892 );
not (  , w_16893 );
and ( w_16892 , w_16893 , \6848_b0 );
or ( \6850_b1 , \6849_b1 , w_16894 );
xor ( \6850_b0 , \6849_b0 , w_16896 );
not ( w_16896 , w_16897 );
and ( w_16897 , w_16894 , w_16895 );
buf ( w_16894 , \5836_b1 );
not ( w_16894 , w_16898 );
not ( w_16895 , w_16899 );
and ( w_16898 , w_16899 , \5836_b0 );
or ( \6851_b1 , \6845_b1 , \6850_b1 );
not ( \6850_b1 , w_16900 );
and ( \6851_b0 , \6845_b0 , w_16901 );
and ( w_16900 , w_16901 , \6850_b0 );
or ( \6852_b1 , \6841_b1 , \6850_b1 );
not ( \6850_b1 , w_16902 );
and ( \6852_b0 , \6841_b0 , w_16903 );
and ( w_16902 , w_16903 , \6850_b0 );
or ( \6854_b1 , \6837_b1 , \6853_b1 );
not ( \6853_b1 , w_16904 );
and ( \6854_b0 , \6837_b0 , w_16905 );
and ( w_16904 , w_16905 , \6853_b0 );
or ( \6855_b1 , \5873_b1 , \5852_b1 );
not ( \5852_b1 , w_16906 );
and ( \6855_b0 , \5873_b0 , w_16907 );
and ( w_16906 , w_16907 , \5852_b0 );
or ( \6856_b1 , \5842_b1 , \5850_b1 );
not ( \5850_b1 , w_16908 );
and ( \6856_b0 , \5842_b0 , w_16909 );
and ( w_16908 , w_16909 , \5850_b0 );
or ( \6857_b1 , \6855_b1 , w_16911 );
not ( w_16911 , w_16912 );
and ( \6857_b0 , \6855_b0 , w_16913 );
and ( w_16912 ,  , w_16913 );
buf ( w_16911 , \6856_b1 );
not ( w_16911 , w_16914 );
not (  , w_16915 );
and ( w_16914 , w_16915 , \6856_b0 );
or ( \6858_b1 , \6857_b1 , w_16916 );
xor ( \6858_b0 , \6857_b0 , w_16918 );
not ( w_16918 , w_16919 );
and ( w_16919 , w_16916 , w_16917 );
buf ( w_16916 , \5859_b1 );
not ( w_16916 , w_16920 );
not ( w_16917 , w_16921 );
and ( w_16920 , w_16921 , \5859_b0 );
or ( \6859_b1 , \5893_b1 , \5871_b1 );
not ( \5871_b1 , w_16922 );
and ( \6859_b0 , \5893_b0 , w_16923 );
and ( w_16922 , w_16923 , \5871_b0 );
or ( \6860_b1 , \5861_b1 , \5869_b1 );
not ( \5869_b1 , w_16924 );
and ( \6860_b0 , \5861_b0 , w_16925 );
and ( w_16924 , w_16925 , \5869_b0 );
or ( \6861_b1 , \6859_b1 , w_16927 );
not ( w_16927 , w_16928 );
and ( \6861_b0 , \6859_b0 , w_16929 );
and ( w_16928 ,  , w_16929 );
buf ( w_16927 , \6860_b1 );
not ( w_16927 , w_16930 );
not (  , w_16931 );
and ( w_16930 , w_16931 , \6860_b0 );
or ( \6862_b1 , \6861_b1 , w_16932 );
xor ( \6862_b0 , \6861_b0 , w_16934 );
not ( w_16934 , w_16935 );
and ( w_16935 , w_16932 , w_16933 );
buf ( w_16932 , \5878_b1 );
not ( w_16932 , w_16936 );
not ( w_16933 , w_16937 );
and ( w_16936 , w_16937 , \5878_b0 );
or ( \6863_b1 , \6858_b1 , \6862_b1 );
not ( \6862_b1 , w_16938 );
and ( \6863_b0 , \6858_b0 , w_16939 );
and ( w_16938 , w_16939 , \6862_b0 );
or ( \6864_b1 , \5918_b1 , \5891_b1 );
not ( \5891_b1 , w_16940 );
and ( \6864_b0 , \5918_b0 , w_16941 );
and ( w_16940 , w_16941 , \5891_b0 );
or ( \6865_b1 , \5881_b1 , \5889_b1 );
not ( \5889_b1 , w_16942 );
and ( \6865_b0 , \5881_b0 , w_16943 );
and ( w_16942 , w_16943 , \5889_b0 );
or ( \6866_b1 , \6864_b1 , w_16945 );
not ( w_16945 , w_16946 );
and ( \6866_b0 , \6864_b0 , w_16947 );
and ( w_16946 ,  , w_16947 );
buf ( w_16945 , \6865_b1 );
not ( w_16945 , w_16948 );
not (  , w_16949 );
and ( w_16948 , w_16949 , \6865_b0 );
or ( \6867_b1 , \6866_b1 , w_16950 );
xor ( \6867_b0 , \6866_b0 , w_16952 );
not ( w_16952 , w_16953 );
and ( w_16953 , w_16950 , w_16951 );
buf ( w_16950 , \5898_b1 );
not ( w_16950 , w_16954 );
not ( w_16951 , w_16955 );
and ( w_16954 , w_16955 , \5898_b0 );
or ( \6868_b1 , \6862_b1 , \6867_b1 );
not ( \6867_b1 , w_16956 );
and ( \6868_b0 , \6862_b0 , w_16957 );
and ( w_16956 , w_16957 , \6867_b0 );
or ( \6869_b1 , \6858_b1 , \6867_b1 );
not ( \6867_b1 , w_16958 );
and ( \6869_b0 , \6858_b0 , w_16959 );
and ( w_16958 , w_16959 , \6867_b0 );
or ( \6871_b1 , \6853_b1 , \6870_b1 );
not ( \6870_b1 , w_16960 );
and ( \6871_b0 , \6853_b0 , w_16961 );
and ( w_16960 , w_16961 , \6870_b0 );
or ( \6872_b1 , \6837_b1 , \6870_b1 );
not ( \6870_b1 , w_16962 );
and ( \6872_b0 , \6837_b0 , w_16963 );
and ( w_16962 , w_16963 , \6870_b0 );
or ( \6874_b1 , \5937_b1 , \5916_b1 );
not ( \5916_b1 , w_16964 );
and ( \6874_b0 , \5937_b0 , w_16965 );
and ( w_16964 , w_16965 , \5916_b0 );
or ( \6875_b1 , \5906_b1 , \5914_b1 );
not ( \5914_b1 , w_16966 );
and ( \6875_b0 , \5906_b0 , w_16967 );
and ( w_16966 , w_16967 , \5914_b0 );
or ( \6876_b1 , \6874_b1 , w_16969 );
not ( w_16969 , w_16970 );
and ( \6876_b0 , \6874_b0 , w_16971 );
and ( w_16970 ,  , w_16971 );
buf ( w_16969 , \6875_b1 );
not ( w_16969 , w_16972 );
not (  , w_16973 );
and ( w_16972 , w_16973 , \6875_b0 );
or ( \6877_b1 , \6876_b1 , w_16974 );
xor ( \6877_b0 , \6876_b0 , w_16976 );
not ( w_16976 , w_16977 );
and ( w_16977 , w_16974 , w_16975 );
buf ( w_16974 , \5923_b1 );
not ( w_16974 , w_16978 );
not ( w_16975 , w_16979 );
and ( w_16978 , w_16979 , \5923_b0 );
or ( \6878_b1 , \5957_b1 , \5935_b1 );
not ( \5935_b1 , w_16980 );
and ( \6878_b0 , \5957_b0 , w_16981 );
and ( w_16980 , w_16981 , \5935_b0 );
or ( \6879_b1 , \5925_b1 , \5933_b1 );
not ( \5933_b1 , w_16982 );
and ( \6879_b0 , \5925_b0 , w_16983 );
and ( w_16982 , w_16983 , \5933_b0 );
or ( \6880_b1 , \6878_b1 , w_16985 );
not ( w_16985 , w_16986 );
and ( \6880_b0 , \6878_b0 , w_16987 );
and ( w_16986 ,  , w_16987 );
buf ( w_16985 , \6879_b1 );
not ( w_16985 , w_16988 );
not (  , w_16989 );
and ( w_16988 , w_16989 , \6879_b0 );
or ( \6881_b1 , \6880_b1 , w_16990 );
xor ( \6881_b0 , \6880_b0 , w_16992 );
not ( w_16992 , w_16993 );
and ( w_16993 , w_16990 , w_16991 );
buf ( w_16990 , \5942_b1 );
not ( w_16990 , w_16994 );
not ( w_16991 , w_16995 );
and ( w_16994 , w_16995 , \5942_b0 );
or ( \6882_b1 , \6877_b1 , \6881_b1 );
not ( \6881_b1 , w_16996 );
and ( \6882_b0 , \6877_b0 , w_16997 );
and ( w_16996 , w_16997 , \6881_b0 );
or ( \6883_b1 , \5979_b1 , \5955_b1 );
not ( \5955_b1 , w_16998 );
and ( \6883_b0 , \5979_b0 , w_16999 );
and ( w_16998 , w_16999 , \5955_b0 );
or ( \6884_b1 , \5945_b1 , \5953_b1 );
not ( \5953_b1 , w_17000 );
and ( \6884_b0 , \5945_b0 , w_17001 );
and ( w_17000 , w_17001 , \5953_b0 );
or ( \6885_b1 , \6883_b1 , w_17003 );
not ( w_17003 , w_17004 );
and ( \6885_b0 , \6883_b0 , w_17005 );
and ( w_17004 ,  , w_17005 );
buf ( w_17003 , \6884_b1 );
not ( w_17003 , w_17006 );
not (  , w_17007 );
and ( w_17006 , w_17007 , \6884_b0 );
or ( \6886_b1 , \6885_b1 , w_17008 );
xor ( \6886_b0 , \6885_b0 , w_17010 );
not ( w_17010 , w_17011 );
and ( w_17011 , w_17008 , w_17009 );
buf ( w_17008 , \5962_b1 );
not ( w_17008 , w_17012 );
not ( w_17009 , w_17013 );
and ( w_17012 , w_17013 , \5962_b0 );
or ( \6887_b1 , \6881_b1 , \6886_b1 );
not ( \6886_b1 , w_17014 );
and ( \6887_b0 , \6881_b0 , w_17015 );
and ( w_17014 , w_17015 , \6886_b0 );
or ( \6888_b1 , \6877_b1 , \6886_b1 );
not ( \6886_b1 , w_17016 );
and ( \6888_b0 , \6877_b0 , w_17017 );
and ( w_17016 , w_17017 , \6886_b0 );
or ( \6890_b1 , \5998_b1 , \5977_b1 );
not ( \5977_b1 , w_17018 );
and ( \6890_b0 , \5998_b0 , w_17019 );
and ( w_17018 , w_17019 , \5977_b0 );
or ( \6891_b1 , \5967_b1 , \5975_b1 );
not ( \5975_b1 , w_17020 );
and ( \6891_b0 , \5967_b0 , w_17021 );
and ( w_17020 , w_17021 , \5975_b0 );
or ( \6892_b1 , \6890_b1 , w_17023 );
not ( w_17023 , w_17024 );
and ( \6892_b0 , \6890_b0 , w_17025 );
and ( w_17024 ,  , w_17025 );
buf ( w_17023 , \6891_b1 );
not ( w_17023 , w_17026 );
not (  , w_17027 );
and ( w_17026 , w_17027 , \6891_b0 );
or ( \6893_b1 , \6892_b1 , w_17028 );
xor ( \6893_b0 , \6892_b0 , w_17030 );
not ( w_17030 , w_17031 );
and ( w_17031 , w_17028 , w_17029 );
buf ( w_17028 , \5984_b1 );
not ( w_17028 , w_17032 );
not ( w_17029 , w_17033 );
and ( w_17032 , w_17033 , \5984_b0 );
or ( \6894_b1 , \6018_b1 , \5996_b1 );
not ( \5996_b1 , w_17034 );
and ( \6894_b0 , \6018_b0 , w_17035 );
and ( w_17034 , w_17035 , \5996_b0 );
or ( \6895_b1 , \5986_b1 , \5994_b1 );
not ( \5994_b1 , w_17036 );
and ( \6895_b0 , \5986_b0 , w_17037 );
and ( w_17036 , w_17037 , \5994_b0 );
or ( \6896_b1 , \6894_b1 , w_17039 );
not ( w_17039 , w_17040 );
and ( \6896_b0 , \6894_b0 , w_17041 );
and ( w_17040 ,  , w_17041 );
buf ( w_17039 , \6895_b1 );
not ( w_17039 , w_17042 );
not (  , w_17043 );
and ( w_17042 , w_17043 , \6895_b0 );
or ( \6897_b1 , \6896_b1 , w_17044 );
xor ( \6897_b0 , \6896_b0 , w_17046 );
not ( w_17046 , w_17047 );
and ( w_17047 , w_17044 , w_17045 );
buf ( w_17044 , \6003_b1 );
not ( w_17044 , w_17048 );
not ( w_17045 , w_17049 );
and ( w_17048 , w_17049 , \6003_b0 );
or ( \6898_b1 , \6893_b1 , \6897_b1 );
not ( \6897_b1 , w_17050 );
and ( \6898_b0 , \6893_b0 , w_17051 );
and ( w_17050 , w_17051 , \6897_b0 );
or ( \6899_b1 , \6041_b1 , \6016_b1 );
not ( \6016_b1 , w_17052 );
and ( \6899_b0 , \6041_b0 , w_17053 );
and ( w_17052 , w_17053 , \6016_b0 );
or ( \6900_b1 , \6006_b1 , \6014_b1 );
not ( \6014_b1 , w_17054 );
and ( \6900_b0 , \6006_b0 , w_17055 );
and ( w_17054 , w_17055 , \6014_b0 );
or ( \6901_b1 , \6899_b1 , w_17057 );
not ( w_17057 , w_17058 );
and ( \6901_b0 , \6899_b0 , w_17059 );
and ( w_17058 ,  , w_17059 );
buf ( w_17057 , \6900_b1 );
not ( w_17057 , w_17060 );
not (  , w_17061 );
and ( w_17060 , w_17061 , \6900_b0 );
or ( \6902_b1 , \6901_b1 , w_17062 );
xor ( \6902_b0 , \6901_b0 , w_17064 );
not ( w_17064 , w_17065 );
and ( w_17065 , w_17062 , w_17063 );
buf ( w_17062 , \6023_b1 );
not ( w_17062 , w_17066 );
not ( w_17063 , w_17067 );
and ( w_17066 , w_17067 , \6023_b0 );
or ( \6903_b1 , \6897_b1 , \6902_b1 );
not ( \6902_b1 , w_17068 );
and ( \6903_b0 , \6897_b0 , w_17069 );
and ( w_17068 , w_17069 , \6902_b0 );
or ( \6904_b1 , \6893_b1 , \6902_b1 );
not ( \6902_b1 , w_17070 );
and ( \6904_b0 , \6893_b0 , w_17071 );
and ( w_17070 , w_17071 , \6902_b0 );
or ( \6906_b1 , \6889_b1 , \6905_b1 );
not ( \6905_b1 , w_17072 );
and ( \6906_b0 , \6889_b0 , w_17073 );
and ( w_17072 , w_17073 , \6905_b0 );
or ( \6907_b1 , \6057_b1 , \6039_b1 );
not ( \6039_b1 , w_17074 );
and ( \6907_b0 , \6057_b0 , w_17075 );
and ( w_17074 , w_17075 , \6039_b0 );
or ( \6908_b1 , \6029_b1 , \6037_b1 );
not ( \6037_b1 , w_17076 );
and ( \6908_b0 , \6029_b0 , w_17077 );
and ( w_17076 , w_17077 , \6037_b0 );
or ( \6909_b1 , \6907_b1 , w_17079 );
not ( w_17079 , w_17080 );
and ( \6909_b0 , \6907_b0 , w_17081 );
and ( w_17080 ,  , w_17081 );
buf ( w_17079 , \6908_b1 );
not ( w_17079 , w_17082 );
not (  , w_17083 );
and ( w_17082 , w_17083 , \6908_b0 );
or ( \6910_b1 , \6909_b1 , w_17084 );
xor ( \6910_b0 , \6909_b0 , w_17086 );
not ( w_17086 , w_17087 );
and ( w_17087 , w_17084 , w_17085 );
buf ( w_17084 , \6046_b1 );
not ( w_17084 , w_17088 );
not ( w_17085 , w_17089 );
and ( w_17088 , w_17089 , \6046_b0 );
or ( \6911_b1 , \6065_b1 , \6055_b1 );
not ( \6055_b1 , w_17090 );
and ( \6911_b0 , \6065_b0 , w_17091 );
and ( w_17090 , w_17091 , \6055_b0 );
or ( \6912_b1 , \6048_b1 , \6053_b1 );
not ( \6053_b1 , w_17092 );
and ( \6912_b0 , \6048_b0 , w_17093 );
and ( w_17092 , w_17093 , \6053_b0 );
or ( \6913_b1 , \6911_b1 , w_17095 );
not ( w_17095 , w_17096 );
and ( \6913_b0 , \6911_b0 , w_17097 );
and ( w_17096 ,  , w_17097 );
buf ( w_17095 , \6912_b1 );
not ( w_17095 , w_17098 );
not (  , w_17099 );
and ( w_17098 , w_17099 , \6912_b0 );
or ( \6914_b1 , \6913_b1 , w_17100 );
xor ( \6914_b0 , \6913_b0 , w_17102 );
not ( w_17102 , w_17103 );
and ( w_17103 , w_17100 , w_17101 );
buf ( w_17100 , \6062_b1 );
not ( w_17100 , w_17104 );
not ( w_17101 , w_17105 );
and ( w_17104 , w_17105 , \6062_b0 );
or ( \6915_b1 , \6910_b1 , \6914_b1 );
not ( \6914_b1 , w_17106 );
and ( \6915_b0 , \6910_b0 , w_17107 );
and ( w_17106 , w_17107 , \6914_b0 );
or ( \6916_b1 , \6905_b1 , \6915_b1 );
not ( \6915_b1 , w_17108 );
and ( \6916_b0 , \6905_b0 , w_17109 );
and ( w_17108 , w_17109 , \6915_b0 );
or ( \6917_b1 , \6889_b1 , \6915_b1 );
not ( \6915_b1 , w_17110 );
and ( \6917_b0 , \6889_b0 , w_17111 );
and ( w_17110 , w_17111 , \6915_b0 );
or ( \6919_b1 , \6873_b1 , \6918_b1 );
not ( \6918_b1 , w_17112 );
and ( \6919_b0 , \6873_b0 , w_17113 );
and ( w_17112 , w_17113 , \6918_b0 );
or ( \6920_b1 , \6047_b1 , \6063_b1 );
xor ( \6920_b0 , \6047_b0 , w_17114 );
not ( w_17114 , w_17115 );
and ( w_17115 , \6063_b1 , \6063_b0 );
or ( \6921_b1 , \6920_b1 , \6068_b1 );
xor ( \6921_b0 , \6920_b0 , w_17116 );
not ( w_17116 , w_17117 );
and ( w_17117 , \6068_b1 , \6068_b0 );
or ( \6922_b1 , \5985_b1 , \6004_b1 );
xor ( \6922_b0 , \5985_b0 , w_17118 );
not ( w_17118 , w_17119 );
and ( w_17119 , \6004_b1 , \6004_b0 );
or ( \6923_b1 , \6922_b1 , \6024_b1 );
xor ( \6923_b0 , \6922_b0 , w_17120 );
not ( w_17120 , w_17121 );
and ( w_17121 , \6024_b1 , \6024_b0 );
or ( \6924_b1 , \6921_b1 , w_17122 );
or ( \6924_b0 , \6921_b0 , \6923_b0 );
not ( \6923_b0 , w_17123 );
and ( w_17123 , w_17122 , \6923_b1 );
or ( \6925_b1 , \6918_b1 , \6924_b1 );
not ( \6924_b1 , w_17124 );
and ( \6925_b0 , \6918_b0 , w_17125 );
and ( w_17124 , w_17125 , \6924_b0 );
or ( \6926_b1 , \6873_b1 , \6924_b1 );
not ( \6924_b1 , w_17126 );
and ( \6926_b0 , \6873_b0 , w_17127 );
and ( w_17126 , w_17127 , \6924_b0 );
or ( \6928_b1 , \5924_b1 , \5943_b1 );
xor ( \6928_b0 , \5924_b0 , w_17128 );
not ( w_17128 , w_17129 );
and ( w_17129 , \5943_b1 , \5943_b0 );
or ( \6929_b1 , \6928_b1 , \5963_b1 );
xor ( \6929_b0 , \6928_b0 , w_17130 );
not ( w_17130 , w_17131 );
and ( w_17131 , \5963_b1 , \5963_b0 );
or ( \6930_b1 , \5860_b1 , \5879_b1 );
xor ( \6930_b0 , \5860_b0 , w_17132 );
not ( w_17132 , w_17133 );
and ( w_17133 , \5879_b1 , \5879_b0 );
or ( \6931_b1 , \6930_b1 , \5899_b1 );
xor ( \6931_b0 , \6930_b0 , w_17134 );
not ( w_17134 , w_17135 );
and ( w_17135 , \5899_b1 , \5899_b0 );
or ( \6932_b1 , \6929_b1 , \6931_b1 );
not ( \6931_b1 , w_17136 );
and ( \6932_b0 , \6929_b0 , w_17137 );
and ( w_17136 , w_17137 , \6931_b0 );
or ( \6933_b1 , \5798_b1 , \5817_b1 );
xor ( \6933_b0 , \5798_b0 , w_17138 );
not ( w_17138 , w_17139 );
and ( w_17139 , \5817_b1 , \5817_b0 );
or ( \6934_b1 , \6933_b1 , \5837_b1 );
xor ( \6934_b0 , \6933_b0 , w_17140 );
not ( w_17140 , w_17141 );
and ( w_17141 , \5837_b1 , \5837_b0 );
or ( \6935_b1 , \6931_b1 , \6934_b1 );
not ( \6934_b1 , w_17142 );
and ( \6935_b0 , \6931_b0 , w_17143 );
and ( w_17142 , w_17143 , \6934_b0 );
or ( \6936_b1 , \6929_b1 , \6934_b1 );
not ( \6934_b1 , w_17144 );
and ( \6936_b0 , \6929_b0 , w_17145 );
and ( w_17144 , w_17145 , \6934_b0 );
or ( \6938_b1 , \6136_b1 , \6150_b1 );
xor ( \6938_b0 , \6136_b0 , w_17146 );
not ( w_17146 , w_17147 );
and ( w_17147 , \6150_b1 , \6150_b0 );
or ( \6939_b1 , \6938_b1 , \6162_b1 );
xor ( \6939_b0 , \6938_b0 , w_17148 );
not ( w_17148 , w_17149 );
and ( w_17149 , \6162_b1 , \6162_b0 );
or ( \6940_b1 , \6937_b1 , \6939_b1 );
not ( \6939_b1 , w_17150 );
and ( \6940_b0 , \6937_b0 , w_17151 );
and ( w_17150 , w_17151 , \6939_b0 );
or ( \6941_b1 , \6087_b1 , \6101_b1 );
xor ( \6941_b0 , \6087_b0 , w_17152 );
not ( w_17152 , w_17153 );
and ( w_17153 , \6101_b1 , \6101_b0 );
or ( \6942_b1 , \6941_b1 , \6116_b1 );
xor ( \6942_b0 , \6941_b0 , w_17154 );
not ( w_17154 , w_17155 );
and ( w_17155 , \6116_b1 , \6116_b0 );
or ( \6943_b1 , \6939_b1 , \6942_b1 );
not ( \6942_b1 , w_17156 );
and ( \6943_b0 , \6939_b0 , w_17157 );
and ( w_17156 , w_17157 , \6942_b0 );
or ( \6944_b1 , \6937_b1 , \6942_b1 );
not ( \6942_b1 , w_17158 );
and ( \6944_b0 , \6937_b0 , w_17159 );
and ( w_17158 , w_17159 , \6942_b0 );
or ( \6946_b1 , \6927_b1 , \6945_b1 );
not ( \6945_b1 , w_17160 );
and ( \6946_b0 , \6927_b0 , w_17161 );
and ( w_17160 , w_17161 , \6945_b0 );
or ( \6947_b1 , \5966_b1 , \6027_b1 );
xor ( \6947_b0 , \5966_b0 , w_17162 );
not ( w_17162 , w_17163 );
and ( w_17163 , \6027_b1 , \6027_b0 );
or ( \6948_b1 , \6947_b1 , \6071_b1 );
xor ( \6948_b0 , \6947_b0 , w_17164 );
not ( w_17164 , w_17165 );
and ( w_17165 , \6071_b1 , \6071_b0 );
or ( \6949_b1 , \5779_b1 , \5840_b1 );
xor ( \6949_b0 , \5779_b0 , w_17166 );
not ( w_17166 , w_17167 );
and ( w_17167 , \5840_b1 , \5840_b0 );
or ( \6950_b1 , \6949_b1 , \5902_b1 );
xor ( \6950_b0 , \6949_b0 , w_17168 );
not ( w_17168 , w_17169 );
and ( w_17169 , \5902_b1 , \5902_b0 );
or ( \6951_b1 , \6948_b1 , \6950_b1 );
not ( \6950_b1 , w_17170 );
and ( \6951_b0 , \6948_b0 , w_17171 );
and ( w_17170 , w_17171 , \6950_b0 );
or ( \6952_b1 , \6945_b1 , \6951_b1 );
not ( \6951_b1 , w_17172 );
and ( \6952_b0 , \6945_b0 , w_17173 );
and ( w_17172 , w_17173 , \6951_b0 );
or ( \6953_b1 , \6927_b1 , \6951_b1 );
not ( \6951_b1 , w_17174 );
and ( \6953_b0 , \6927_b0 , w_17175 );
and ( w_17174 , w_17175 , \6951_b0 );
or ( \6955_b1 , \6313_b1 , \6324_b1 );
xor ( \6955_b0 , \6313_b0 , w_17176 );
not ( w_17176 , w_17177 );
and ( w_17177 , \6324_b1 , \6324_b0 );
or ( \6956_b1 , \6955_b1 , \6339_b1 );
xor ( \6956_b0 , \6955_b0 , w_17178 );
not ( w_17178 , w_17179 );
and ( w_17179 , \6339_b1 , \6339_b0 );
or ( \6957_b1 , \6165_b1 , \6236_b1 );
xor ( \6957_b0 , \6165_b0 , w_17180 );
not ( w_17180 , w_17181 );
and ( w_17181 , \6236_b1 , \6236_b0 );
or ( \6958_b1 , \6957_b1 , \6281_b1 );
xor ( \6958_b0 , \6957_b0 , w_17182 );
not ( w_17182 , w_17183 );
and ( w_17183 , \6281_b1 , \6281_b0 );
or ( \6959_b1 , \6956_b1 , \6958_b1 );
not ( \6958_b1 , w_17184 );
and ( \6959_b0 , \6956_b0 , w_17185 );
and ( w_17184 , w_17185 , \6958_b0 );
or ( \6960_b1 , \5905_b1 , \6074_b1 );
xor ( \6960_b0 , \5905_b0 , w_17186 );
not ( w_17186 , w_17187 );
and ( w_17187 , \6074_b1 , \6074_b0 );
or ( \6961_b1 , \6960_b1 , \6119_b1 );
xor ( \6961_b0 , \6960_b0 , w_17188 );
not ( w_17188 , w_17189 );
and ( w_17189 , \6119_b1 , \6119_b0 );
or ( \6962_b1 , \6958_b1 , \6961_b1 );
not ( \6961_b1 , w_17190 );
and ( \6962_b0 , \6958_b0 , w_17191 );
and ( w_17190 , w_17191 , \6961_b0 );
or ( \6963_b1 , \6956_b1 , \6961_b1 );
not ( \6961_b1 , w_17192 );
and ( \6963_b0 , \6956_b0 , w_17193 );
and ( w_17192 , w_17193 , \6961_b0 );
or ( \6965_b1 , \6954_b1 , \6964_b1 );
not ( \6964_b1 , w_17194 );
and ( \6965_b0 , \6954_b0 , w_17195 );
and ( w_17194 , w_17195 , \6964_b0 );
or ( \6966_b1 , \6374_b1 , \6463_b1 );
xor ( \6966_b0 , \6374_b0 , w_17196 );
not ( w_17196 , w_17197 );
and ( w_17197 , \6463_b1 , \6463_b0 );
or ( \6967_b1 , \6966_b1 , \6475_b1 );
xor ( \6967_b0 , \6966_b0 , w_17198 );
not ( w_17198 , w_17199 );
and ( w_17199 , \6475_b1 , \6475_b0 );
or ( \6968_b1 , \6964_b1 , \6967_b1 );
not ( \6967_b1 , w_17200 );
and ( \6968_b0 , \6964_b0 , w_17201 );
and ( w_17200 , w_17201 , \6967_b0 );
or ( \6969_b1 , \6954_b1 , \6967_b1 );
not ( \6967_b1 , w_17202 );
and ( \6969_b0 , \6954_b0 , w_17203 );
and ( w_17202 , w_17203 , \6967_b0 );
or ( \6971_b1 , \6668_b1 , \6672_b1 );
xor ( \6971_b0 , \6668_b0 , w_17204 );
not ( w_17204 , w_17205 );
and ( w_17205 , \6672_b1 , \6672_b0 );
or ( \6972_b1 , \6971_b1 , \6674_b1 );
xor ( \6972_b0 , \6971_b0 , w_17206 );
not ( w_17206 , w_17207 );
and ( w_17207 , \6674_b1 , \6674_b0 );
or ( \6973_b1 , \6970_b1 , \6972_b1 );
not ( \6972_b1 , w_17208 );
and ( \6973_b0 , \6970_b0 , w_17209 );
and ( w_17208 , w_17209 , \6972_b0 );
or ( \6974_b1 , \6345_b1 , \6478_b1 );
xor ( \6974_b0 , \6345_b0 , w_17210 );
not ( w_17210 , w_17211 );
and ( w_17211 , \6478_b1 , \6478_b0 );
or ( \6975_b1 , \6974_b1 , \6646_b1 );
xor ( \6975_b0 , \6974_b0 , w_17212 );
not ( w_17212 , w_17213 );
and ( w_17213 , \6646_b1 , \6646_b0 );
or ( \6976_b1 , \6972_b1 , \6975_b1 );
not ( \6975_b1 , w_17214 );
and ( \6976_b0 , \6972_b0 , w_17215 );
and ( w_17214 , w_17215 , \6975_b0 );
or ( \6977_b1 , \6970_b1 , \6975_b1 );
not ( \6975_b1 , w_17216 );
and ( \6977_b0 , \6970_b0 , w_17217 );
and ( w_17216 , w_17217 , \6975_b0 );
or ( \6979_b1 , \6815_b1 , w_17219 );
not ( w_17219 , w_17220 );
and ( \6979_b0 , \6815_b0 , w_17221 );
and ( w_17220 ,  , w_17221 );
buf ( w_17219 , \6978_b1 );
not ( w_17219 , w_17222 );
not (  , w_17223 );
and ( w_17222 , w_17223 , \6978_b0 );
or ( \6980_b1 , \6815_b1 , w_17225 );
not ( w_17225 , w_17226 );
and ( \6980_b0 , \6815_b0 , w_17227 );
and ( w_17226 ,  , w_17227 );
buf ( w_17225 , \6978_b1 );
not ( w_17225 , w_17228 );
not (  , w_17229 );
and ( w_17228 , w_17229 , \6978_b0 );
buf ( \6981_b1 , \6980_b1 );
not ( \6981_b1 , w_17230 );
not ( \6981_b0 , w_17231 );
and ( w_17230 , w_17231 , \6980_b0 );
or ( \6982_b1 , \6979_b1 , w_17233 );
not ( w_17233 , w_17234 );
and ( \6982_b0 , \6979_b0 , w_17235 );
and ( w_17234 ,  , w_17235 );
buf ( w_17233 , \6981_b1 );
not ( w_17233 , w_17236 );
not (  , w_17237 );
and ( w_17236 , w_17237 , \6981_b0 );
or ( \6983_b1 , \5606_b1 , \5609_b1 );
xor ( \6983_b0 , \5606_b0 , w_17238 );
not ( w_17238 , w_17239 );
and ( w_17239 , \5609_b1 , \5609_b0 );
buf ( \6984_b1 , \6983_b1 );
buf ( \6984_b0 , \6983_b0 );
buf ( \6985_b1 , \6984_b1 );
buf ( \6985_b0 , \6984_b0 );
or ( \6986_b1 , \5608_b1 , \2371_b1 );
xor ( \6986_b0 , \5608_b0 , w_17240 );
not ( w_17240 , w_17241 );
and ( w_17241 , \2371_b1 , \2371_b0 );
buf ( \6987_b1 , \6986_b1 );
buf ( \6987_b0 , \6986_b0 );
buf ( \6988_b1 , \6987_b1 );
buf ( \6988_b0 , \6987_b0 );
or ( \6989_b1 , \6985_b1 , \6988_b1 );
xor ( \6989_b0 , \6985_b0 , w_17242 );
not ( w_17242 , w_17243 );
and ( w_17243 , \6988_b1 , \6988_b0 );
buf ( \6990_b1 , \6988_b1 );
not ( \6990_b1 , w_17244 );
not ( \6990_b0 , w_17245 );
and ( w_17244 , w_17245 , \6988_b0 );
or ( \6991_b1 , \6989_b1 , \6990_b1 );
not ( \6990_b1 , w_17246 );
and ( \6991_b0 , \6989_b0 , w_17247 );
and ( w_17246 , w_17247 , \6990_b0 );
or ( \6992_b1 , \5799_b1 , \6991_b1 );
not ( \6991_b1 , w_17248 );
and ( \6992_b0 , \5799_b0 , w_17249 );
and ( w_17248 , w_17249 , \6991_b0 );
or ( \6993_b1 , \5811_b1 , \6988_b1 );
not ( \6988_b1 , w_17250 );
and ( \6993_b0 , \5811_b0 , w_17251 );
and ( w_17250 , w_17251 , \6988_b0 );
or ( \6994_b1 , \6992_b1 , w_17253 );
not ( w_17253 , w_17254 );
and ( \6994_b0 , \6992_b0 , w_17255 );
and ( w_17254 ,  , w_17255 );
buf ( w_17253 , \6993_b1 );
not ( w_17253 , w_17256 );
not (  , w_17257 );
and ( w_17256 , w_17257 , \6993_b0 );
or ( \6995_b1 , \6994_b1 , w_17258 );
xor ( \6995_b0 , \6994_b0 , w_17260 );
not ( w_17260 , w_17261 );
and ( w_17261 , w_17258 , w_17259 );
buf ( w_17258 , \6985_b1 );
not ( w_17258 , w_17262 );
not ( w_17259 , w_17263 );
and ( w_17262 , w_17263 , \6985_b0 );
or ( \6996_b1 , \5755_b1 , \6995_b1 );
not ( \6995_b1 , w_17264 );
and ( \6996_b0 , \5755_b0 , w_17265 );
and ( w_17264 , w_17265 , \6995_b0 );
or ( \6997_b1 , \5597_b1 , \5612_b1 );
xor ( \6997_b0 , \5597_b0 , w_17266 );
not ( w_17266 , w_17267 );
and ( w_17267 , \5612_b1 , \5612_b0 );
buf ( \6998_b1 , \6997_b1 );
buf ( \6998_b0 , \6997_b0 );
buf ( \6999_b1 , \6998_b1 );
buf ( \6999_b0 , \6998_b0 );
or ( \7000_b1 , \5602_b1 , \5610_b1 );
xor ( \7000_b0 , \5602_b0 , w_17268 );
not ( w_17268 , w_17269 );
and ( w_17269 , \5610_b1 , \5610_b0 );
buf ( \7001_b1 , \7000_b1 );
buf ( \7001_b0 , \7000_b0 );
buf ( \7002_b1 , \7001_b1 );
buf ( \7002_b0 , \7001_b0 );
or ( \7003_b1 , \6999_b1 , \7002_b1 );
xor ( \7003_b0 , \6999_b0 , w_17270 );
not ( w_17270 , w_17271 );
and ( w_17271 , \7002_b1 , \7002_b0 );
or ( \7004_b1 , \7002_b1 , \6985_b1 );
xor ( \7004_b0 , \7002_b0 , w_17272 );
not ( w_17272 , w_17273 );
and ( w_17273 , \6985_b1 , \6985_b0 );
buf ( \7005_b1 , \7004_b1 );
not ( \7005_b1 , w_17274 );
not ( \7005_b0 , w_17275 );
and ( w_17274 , w_17275 , \7004_b0 );
or ( \7006_b1 , \7003_b1 , \7005_b1 );
not ( \7005_b1 , w_17276 );
and ( \7006_b0 , \7003_b0 , w_17277 );
and ( w_17276 , w_17277 , \7005_b0 );
or ( \7007_b1 , \5819_b1 , \7006_b1 );
not ( \7006_b1 , w_17278 );
and ( \7007_b0 , \5819_b0 , w_17279 );
and ( w_17278 , w_17279 , \7006_b0 );
or ( \7008_b1 , \5831_b1 , \7004_b1 );
not ( \7004_b1 , w_17280 );
and ( \7008_b0 , \5831_b0 , w_17281 );
and ( w_17280 , w_17281 , \7004_b0 );
or ( \7009_b1 , \7007_b1 , w_17283 );
not ( w_17283 , w_17284 );
and ( \7009_b0 , \7007_b0 , w_17285 );
and ( w_17284 ,  , w_17285 );
buf ( w_17283 , \7008_b1 );
not ( w_17283 , w_17286 );
not (  , w_17287 );
and ( w_17286 , w_17287 , \7008_b0 );
or ( \7010_b1 , \7002_b1 , \6985_b1 );
not ( \6985_b1 , w_17288 );
and ( \7010_b0 , \7002_b0 , w_17289 );
and ( w_17288 , w_17289 , \6985_b0 );
buf ( \7011_b1 , \7010_b1 );
not ( \7011_b1 , w_17290 );
not ( \7011_b0 , w_17291 );
and ( w_17290 , w_17291 , \7010_b0 );
or ( \7012_b1 , \6999_b1 , \7011_b1 );
not ( \7011_b1 , w_17292 );
and ( \7012_b0 , \6999_b0 , w_17293 );
and ( w_17292 , w_17293 , \7011_b0 );
or ( \7013_b1 , \7009_b1 , w_17294 );
xor ( \7013_b0 , \7009_b0 , w_17296 );
not ( w_17296 , w_17297 );
and ( w_17297 , w_17294 , w_17295 );
buf ( w_17294 , \7012_b1 );
not ( w_17294 , w_17298 );
not ( w_17295 , w_17299 );
and ( w_17298 , w_17299 , \7012_b0 );
or ( \7014_b1 , \6995_b1 , \7013_b1 );
not ( \7013_b1 , w_17300 );
and ( \7014_b0 , \6995_b0 , w_17301 );
and ( w_17300 , w_17301 , \7013_b0 );
or ( \7015_b1 , \5755_b1 , \7013_b1 );
not ( \7013_b1 , w_17302 );
and ( \7015_b0 , \5755_b0 , w_17303 );
and ( w_17302 , w_17303 , \7013_b0 );
or ( \7017_b1 , \5577_b1 , \5616_b1 );
xor ( \7017_b0 , \5577_b0 , w_17304 );
not ( w_17304 , w_17305 );
and ( w_17305 , \5616_b1 , \5616_b0 );
buf ( \7018_b1 , \7017_b1 );
buf ( \7018_b0 , \7017_b0 );
buf ( \7019_b1 , \7018_b1 );
buf ( \7019_b0 , \7018_b0 );
or ( \7020_b1 , \5589_b1 , \5614_b1 );
xor ( \7020_b0 , \5589_b0 , w_17306 );
not ( w_17306 , w_17307 );
and ( w_17307 , \5614_b1 , \5614_b0 );
buf ( \7021_b1 , \7020_b1 );
buf ( \7021_b0 , \7020_b0 );
buf ( \7022_b1 , \7021_b1 );
buf ( \7022_b0 , \7021_b0 );
or ( \7023_b1 , \7019_b1 , \7022_b1 );
xor ( \7023_b0 , \7019_b0 , w_17308 );
not ( w_17308 , w_17309 );
and ( w_17309 , \7022_b1 , \7022_b0 );
or ( \7024_b1 , \7022_b1 , \6999_b1 );
xor ( \7024_b0 , \7022_b0 , w_17310 );
not ( w_17310 , w_17311 );
and ( w_17311 , \6999_b1 , \6999_b0 );
buf ( \7025_b1 , \7024_b1 );
not ( \7025_b1 , w_17312 );
not ( \7025_b0 , w_17313 );
and ( w_17312 , w_17313 , \7024_b0 );
or ( \7026_b1 , \7023_b1 , \7025_b1 );
not ( \7025_b1 , w_17314 );
and ( \7026_b0 , \7023_b0 , w_17315 );
and ( w_17314 , w_17315 , \7025_b0 );
or ( \7027_b1 , \5842_b1 , \7026_b1 );
not ( \7026_b1 , w_17316 );
and ( \7027_b0 , \5842_b0 , w_17317 );
and ( w_17316 , w_17317 , \7026_b0 );
or ( \7028_b1 , \5854_b1 , \7024_b1 );
not ( \7024_b1 , w_17318 );
and ( \7028_b0 , \5854_b0 , w_17319 );
and ( w_17318 , w_17319 , \7024_b0 );
or ( \7029_b1 , \7027_b1 , w_17321 );
not ( w_17321 , w_17322 );
and ( \7029_b0 , \7027_b0 , w_17323 );
and ( w_17322 ,  , w_17323 );
buf ( w_17321 , \7028_b1 );
not ( w_17321 , w_17324 );
not (  , w_17325 );
and ( w_17324 , w_17325 , \7028_b0 );
or ( \7030_b1 , \7022_b1 , \6999_b1 );
not ( \6999_b1 , w_17326 );
and ( \7030_b0 , \7022_b0 , w_17327 );
and ( w_17326 , w_17327 , \6999_b0 );
buf ( \7031_b1 , \7030_b1 );
not ( \7031_b1 , w_17328 );
not ( \7031_b0 , w_17329 );
and ( w_17328 , w_17329 , \7030_b0 );
or ( \7032_b1 , \7019_b1 , \7031_b1 );
not ( \7031_b1 , w_17330 );
and ( \7032_b0 , \7019_b0 , w_17331 );
and ( w_17330 , w_17331 , \7031_b0 );
or ( \7033_b1 , \7029_b1 , w_17332 );
xor ( \7033_b0 , \7029_b0 , w_17334 );
not ( w_17334 , w_17335 );
and ( w_17335 , w_17332 , w_17333 );
buf ( w_17332 , \7032_b1 );
not ( w_17332 , w_17336 );
not ( w_17333 , w_17337 );
and ( w_17336 , w_17337 , \7032_b0 );
or ( \7034_b1 , \5550_b1 , \5620_b1 );
xor ( \7034_b0 , \5550_b0 , w_17338 );
not ( w_17338 , w_17339 );
and ( w_17339 , \5620_b1 , \5620_b0 );
buf ( \7035_b1 , \7034_b1 );
buf ( \7035_b0 , \7034_b0 );
buf ( \7036_b1 , \7035_b1 );
buf ( \7036_b0 , \7035_b0 );
or ( \7037_b1 , \5569_b1 , \5618_b1 );
xor ( \7037_b0 , \5569_b0 , w_17340 );
not ( w_17340 , w_17341 );
and ( w_17341 , \5618_b1 , \5618_b0 );
buf ( \7038_b1 , \7037_b1 );
buf ( \7038_b0 , \7037_b0 );
buf ( \7039_b1 , \7038_b1 );
buf ( \7039_b0 , \7038_b0 );
or ( \7040_b1 , \7036_b1 , \7039_b1 );
xor ( \7040_b0 , \7036_b0 , w_17342 );
not ( w_17342 , w_17343 );
and ( w_17343 , \7039_b1 , \7039_b0 );
or ( \7041_b1 , \7039_b1 , \7019_b1 );
xor ( \7041_b0 , \7039_b0 , w_17344 );
not ( w_17344 , w_17345 );
and ( w_17345 , \7019_b1 , \7019_b0 );
buf ( \7042_b1 , \7041_b1 );
not ( \7042_b1 , w_17346 );
not ( \7042_b0 , w_17347 );
and ( w_17346 , w_17347 , \7041_b0 );
or ( \7043_b1 , \7040_b1 , \7042_b1 );
not ( \7042_b1 , w_17348 );
and ( \7043_b0 , \7040_b0 , w_17349 );
and ( w_17348 , w_17349 , \7042_b0 );
or ( \7044_b1 , \5861_b1 , \7043_b1 );
not ( \7043_b1 , w_17350 );
and ( \7044_b0 , \5861_b0 , w_17351 );
and ( w_17350 , w_17351 , \7043_b0 );
or ( \7045_b1 , \5873_b1 , \7041_b1 );
not ( \7041_b1 , w_17352 );
and ( \7045_b0 , \5873_b0 , w_17353 );
and ( w_17352 , w_17353 , \7041_b0 );
or ( \7046_b1 , \7044_b1 , w_17355 );
not ( w_17355 , w_17356 );
and ( \7046_b0 , \7044_b0 , w_17357 );
and ( w_17356 ,  , w_17357 );
buf ( w_17355 , \7045_b1 );
not ( w_17355 , w_17358 );
not (  , w_17359 );
and ( w_17358 , w_17359 , \7045_b0 );
or ( \7047_b1 , \7039_b1 , \7019_b1 );
not ( \7019_b1 , w_17360 );
and ( \7047_b0 , \7039_b0 , w_17361 );
and ( w_17360 , w_17361 , \7019_b0 );
buf ( \7048_b1 , \7047_b1 );
not ( \7048_b1 , w_17362 );
not ( \7048_b0 , w_17363 );
and ( w_17362 , w_17363 , \7047_b0 );
or ( \7049_b1 , \7036_b1 , \7048_b1 );
not ( \7048_b1 , w_17364 );
and ( \7049_b0 , \7036_b0 , w_17365 );
and ( w_17364 , w_17365 , \7048_b0 );
or ( \7050_b1 , \7046_b1 , w_17366 );
xor ( \7050_b0 , \7046_b0 , w_17368 );
not ( w_17368 , w_17369 );
and ( w_17369 , w_17366 , w_17367 );
buf ( w_17366 , \7049_b1 );
not ( w_17366 , w_17370 );
not ( w_17367 , w_17371 );
and ( w_17370 , w_17371 , \7049_b0 );
or ( \7051_b1 , \7033_b1 , \7050_b1 );
not ( \7050_b1 , w_17372 );
and ( \7051_b0 , \7033_b0 , w_17373 );
and ( w_17372 , w_17373 , \7050_b0 );
or ( \7052_b1 , \5516_b1 , \5624_b1 );
xor ( \7052_b0 , \5516_b0 , w_17374 );
not ( w_17374 , w_17375 );
and ( w_17375 , \5624_b1 , \5624_b0 );
buf ( \7053_b1 , \7052_b1 );
buf ( \7053_b0 , \7052_b0 );
buf ( \7054_b1 , \7053_b1 );
buf ( \7054_b0 , \7053_b0 );
or ( \7055_b1 , \5524_b1 , \5622_b1 );
xor ( \7055_b0 , \5524_b0 , w_17376 );
not ( w_17376 , w_17377 );
and ( w_17377 , \5622_b1 , \5622_b0 );
buf ( \7056_b1 , \7055_b1 );
buf ( \7056_b0 , \7055_b0 );
buf ( \7057_b1 , \7056_b1 );
buf ( \7057_b0 , \7056_b0 );
or ( \7058_b1 , \7054_b1 , \7057_b1 );
xor ( \7058_b0 , \7054_b0 , w_17378 );
not ( w_17378 , w_17379 );
and ( w_17379 , \7057_b1 , \7057_b0 );
or ( \7059_b1 , \7057_b1 , \7036_b1 );
xor ( \7059_b0 , \7057_b0 , w_17380 );
not ( w_17380 , w_17381 );
and ( w_17381 , \7036_b1 , \7036_b0 );
buf ( \7060_b1 , \7059_b1 );
not ( \7060_b1 , w_17382 );
not ( \7060_b0 , w_17383 );
and ( w_17382 , w_17383 , \7059_b0 );
or ( \7061_b1 , \7058_b1 , \7060_b1 );
not ( \7060_b1 , w_17384 );
and ( \7061_b0 , \7058_b0 , w_17385 );
and ( w_17384 , w_17385 , \7060_b0 );
or ( \7062_b1 , \5881_b1 , \7061_b1 );
not ( \7061_b1 , w_17386 );
and ( \7062_b0 , \5881_b0 , w_17387 );
and ( w_17386 , w_17387 , \7061_b0 );
or ( \7063_b1 , \5893_b1 , \7059_b1 );
not ( \7059_b1 , w_17388 );
and ( \7063_b0 , \5893_b0 , w_17389 );
and ( w_17388 , w_17389 , \7059_b0 );
or ( \7064_b1 , \7062_b1 , w_17391 );
not ( w_17391 , w_17392 );
and ( \7064_b0 , \7062_b0 , w_17393 );
and ( w_17392 ,  , w_17393 );
buf ( w_17391 , \7063_b1 );
not ( w_17391 , w_17394 );
not (  , w_17395 );
and ( w_17394 , w_17395 , \7063_b0 );
or ( \7065_b1 , \7057_b1 , \7036_b1 );
not ( \7036_b1 , w_17396 );
and ( \7065_b0 , \7057_b0 , w_17397 );
and ( w_17396 , w_17397 , \7036_b0 );
buf ( \7066_b1 , \7065_b1 );
not ( \7066_b1 , w_17398 );
not ( \7066_b0 , w_17399 );
and ( w_17398 , w_17399 , \7065_b0 );
or ( \7067_b1 , \7054_b1 , \7066_b1 );
not ( \7066_b1 , w_17400 );
and ( \7067_b0 , \7054_b0 , w_17401 );
and ( w_17400 , w_17401 , \7066_b0 );
or ( \7068_b1 , \7064_b1 , w_17402 );
xor ( \7068_b0 , \7064_b0 , w_17404 );
not ( w_17404 , w_17405 );
and ( w_17405 , w_17402 , w_17403 );
buf ( w_17402 , \7067_b1 );
not ( w_17402 , w_17406 );
not ( w_17403 , w_17407 );
and ( w_17406 , w_17407 , \7067_b0 );
or ( \7069_b1 , \7050_b1 , \7068_b1 );
not ( \7068_b1 , w_17408 );
and ( \7069_b0 , \7050_b0 , w_17409 );
and ( w_17408 , w_17409 , \7068_b0 );
or ( \7070_b1 , \7033_b1 , \7068_b1 );
not ( \7068_b1 , w_17410 );
and ( \7070_b0 , \7033_b0 , w_17411 );
and ( w_17410 , w_17411 , \7068_b0 );
or ( \7072_b1 , \7016_b1 , \7071_b1 );
not ( \7071_b1 , w_17412 );
and ( \7072_b0 , \7016_b0 , w_17413 );
and ( w_17412 , w_17413 , \7071_b0 );
or ( \7073_b1 , \5448_b1 , \5628_b1 );
xor ( \7073_b0 , \5448_b0 , w_17414 );
not ( w_17414 , w_17415 );
and ( w_17415 , \5628_b1 , \5628_b0 );
buf ( \7074_b1 , \7073_b1 );
buf ( \7074_b0 , \7073_b0 );
buf ( \7075_b1 , \7074_b1 );
buf ( \7075_b0 , \7074_b0 );
or ( \7076_b1 , \5482_b1 , \5626_b1 );
xor ( \7076_b0 , \5482_b0 , w_17416 );
not ( w_17416 , w_17417 );
and ( w_17417 , \5626_b1 , \5626_b0 );
buf ( \7077_b1 , \7076_b1 );
buf ( \7077_b0 , \7076_b0 );
buf ( \7078_b1 , \7077_b1 );
buf ( \7078_b0 , \7077_b0 );
or ( \7079_b1 , \7075_b1 , \7078_b1 );
xor ( \7079_b0 , \7075_b0 , w_17418 );
not ( w_17418 , w_17419 );
and ( w_17419 , \7078_b1 , \7078_b0 );
or ( \7080_b1 , \7078_b1 , \7054_b1 );
xor ( \7080_b0 , \7078_b0 , w_17420 );
not ( w_17420 , w_17421 );
and ( w_17421 , \7054_b1 , \7054_b0 );
buf ( \7081_b1 , \7080_b1 );
not ( \7081_b1 , w_17422 );
not ( \7081_b0 , w_17423 );
and ( w_17422 , w_17423 , \7080_b0 );
or ( \7082_b1 , \7079_b1 , \7081_b1 );
not ( \7081_b1 , w_17424 );
and ( \7082_b0 , \7079_b0 , w_17425 );
and ( w_17424 , w_17425 , \7081_b0 );
or ( \7083_b1 , \5906_b1 , \7082_b1 );
not ( \7082_b1 , w_17426 );
and ( \7083_b0 , \5906_b0 , w_17427 );
and ( w_17426 , w_17427 , \7082_b0 );
or ( \7084_b1 , \5918_b1 , \7080_b1 );
not ( \7080_b1 , w_17428 );
and ( \7084_b0 , \5918_b0 , w_17429 );
and ( w_17428 , w_17429 , \7080_b0 );
or ( \7085_b1 , \7083_b1 , w_17431 );
not ( w_17431 , w_17432 );
and ( \7085_b0 , \7083_b0 , w_17433 );
and ( w_17432 ,  , w_17433 );
buf ( w_17431 , \7084_b1 );
not ( w_17431 , w_17434 );
not (  , w_17435 );
and ( w_17434 , w_17435 , \7084_b0 );
or ( \7086_b1 , \7078_b1 , \7054_b1 );
not ( \7054_b1 , w_17436 );
and ( \7086_b0 , \7078_b0 , w_17437 );
and ( w_17436 , w_17437 , \7054_b0 );
buf ( \7087_b1 , \7086_b1 );
not ( \7087_b1 , w_17438 );
not ( \7087_b0 , w_17439 );
and ( w_17438 , w_17439 , \7086_b0 );
or ( \7088_b1 , \7075_b1 , \7087_b1 );
not ( \7087_b1 , w_17440 );
and ( \7088_b0 , \7075_b0 , w_17441 );
and ( w_17440 , w_17441 , \7087_b0 );
or ( \7089_b1 , \7085_b1 , w_17442 );
xor ( \7089_b0 , \7085_b0 , w_17444 );
not ( w_17444 , w_17445 );
and ( w_17445 , w_17442 , w_17443 );
buf ( w_17442 , \7088_b1 );
not ( w_17442 , w_17446 );
not ( w_17443 , w_17447 );
and ( w_17446 , w_17447 , \7088_b0 );
or ( \7090_b1 , \5387_b1 , \5632_b1 );
xor ( \7090_b0 , \5387_b0 , w_17448 );
not ( w_17448 , w_17449 );
and ( w_17449 , \5632_b1 , \5632_b0 );
buf ( \7091_b1 , \7090_b1 );
buf ( \7091_b0 , \7090_b0 );
buf ( \7092_b1 , \7091_b1 );
buf ( \7092_b0 , \7091_b0 );
or ( \7093_b1 , \5440_b1 , \5630_b1 );
xor ( \7093_b0 , \5440_b0 , w_17450 );
not ( w_17450 , w_17451 );
and ( w_17451 , \5630_b1 , \5630_b0 );
buf ( \7094_b1 , \7093_b1 );
buf ( \7094_b0 , \7093_b0 );
buf ( \7095_b1 , \7094_b1 );
buf ( \7095_b0 , \7094_b0 );
or ( \7096_b1 , \7092_b1 , \7095_b1 );
xor ( \7096_b0 , \7092_b0 , w_17452 );
not ( w_17452 , w_17453 );
and ( w_17453 , \7095_b1 , \7095_b0 );
or ( \7097_b1 , \7095_b1 , \7075_b1 );
xor ( \7097_b0 , \7095_b0 , w_17454 );
not ( w_17454 , w_17455 );
and ( w_17455 , \7075_b1 , \7075_b0 );
buf ( \7098_b1 , \7097_b1 );
not ( \7098_b1 , w_17456 );
not ( \7098_b0 , w_17457 );
and ( w_17456 , w_17457 , \7097_b0 );
or ( \7099_b1 , \7096_b1 , \7098_b1 );
not ( \7098_b1 , w_17458 );
and ( \7099_b0 , \7096_b0 , w_17459 );
and ( w_17458 , w_17459 , \7098_b0 );
or ( \7100_b1 , \5925_b1 , \7099_b1 );
not ( \7099_b1 , w_17460 );
and ( \7100_b0 , \5925_b0 , w_17461 );
and ( w_17460 , w_17461 , \7099_b0 );
or ( \7101_b1 , \5937_b1 , \7097_b1 );
not ( \7097_b1 , w_17462 );
and ( \7101_b0 , \5937_b0 , w_17463 );
and ( w_17462 , w_17463 , \7097_b0 );
or ( \7102_b1 , \7100_b1 , w_17465 );
not ( w_17465 , w_17466 );
and ( \7102_b0 , \7100_b0 , w_17467 );
and ( w_17466 ,  , w_17467 );
buf ( w_17465 , \7101_b1 );
not ( w_17465 , w_17468 );
not (  , w_17469 );
and ( w_17468 , w_17469 , \7101_b0 );
or ( \7103_b1 , \7095_b1 , \7075_b1 );
not ( \7075_b1 , w_17470 );
and ( \7103_b0 , \7095_b0 , w_17471 );
and ( w_17470 , w_17471 , \7075_b0 );
buf ( \7104_b1 , \7103_b1 );
not ( \7104_b1 , w_17472 );
not ( \7104_b0 , w_17473 );
and ( w_17472 , w_17473 , \7103_b0 );
or ( \7105_b1 , \7092_b1 , \7104_b1 );
not ( \7104_b1 , w_17474 );
and ( \7105_b0 , \7092_b0 , w_17475 );
and ( w_17474 , w_17475 , \7104_b0 );
or ( \7106_b1 , \7102_b1 , w_17476 );
xor ( \7106_b0 , \7102_b0 , w_17478 );
not ( w_17478 , w_17479 );
and ( w_17479 , w_17476 , w_17477 );
buf ( w_17476 , \7105_b1 );
not ( w_17476 , w_17480 );
not ( w_17477 , w_17481 );
and ( w_17480 , w_17481 , \7105_b0 );
or ( \7107_b1 , \7089_b1 , \7106_b1 );
not ( \7106_b1 , w_17482 );
and ( \7107_b0 , \7089_b0 , w_17483 );
and ( w_17482 , w_17483 , \7106_b0 );
or ( \7108_b1 , \5295_b1 , \5636_b1 );
xor ( \7108_b0 , \5295_b0 , w_17484 );
not ( w_17484 , w_17485 );
and ( w_17485 , \5636_b1 , \5636_b0 );
buf ( \7109_b1 , \7108_b1 );
buf ( \7109_b0 , \7108_b0 );
buf ( \7110_b1 , \7109_b1 );
buf ( \7110_b0 , \7109_b0 );
or ( \7111_b1 , \5348_b1 , \5634_b1 );
xor ( \7111_b0 , \5348_b0 , w_17486 );
not ( w_17486 , w_17487 );
and ( w_17487 , \5634_b1 , \5634_b0 );
buf ( \7112_b1 , \7111_b1 );
buf ( \7112_b0 , \7111_b0 );
buf ( \7113_b1 , \7112_b1 );
buf ( \7113_b0 , \7112_b0 );
or ( \7114_b1 , \7110_b1 , \7113_b1 );
xor ( \7114_b0 , \7110_b0 , w_17488 );
not ( w_17488 , w_17489 );
and ( w_17489 , \7113_b1 , \7113_b0 );
or ( \7115_b1 , \7113_b1 , \7092_b1 );
xor ( \7115_b0 , \7113_b0 , w_17490 );
not ( w_17490 , w_17491 );
and ( w_17491 , \7092_b1 , \7092_b0 );
buf ( \7116_b1 , \7115_b1 );
not ( \7116_b1 , w_17492 );
not ( \7116_b0 , w_17493 );
and ( w_17492 , w_17493 , \7115_b0 );
or ( \7117_b1 , \7114_b1 , \7116_b1 );
not ( \7116_b1 , w_17494 );
and ( \7117_b0 , \7114_b0 , w_17495 );
and ( w_17494 , w_17495 , \7116_b0 );
or ( \7118_b1 , \5945_b1 , \7117_b1 );
not ( \7117_b1 , w_17496 );
and ( \7118_b0 , \5945_b0 , w_17497 );
and ( w_17496 , w_17497 , \7117_b0 );
or ( \7119_b1 , \5957_b1 , \7115_b1 );
not ( \7115_b1 , w_17498 );
and ( \7119_b0 , \5957_b0 , w_17499 );
and ( w_17498 , w_17499 , \7115_b0 );
or ( \7120_b1 , \7118_b1 , w_17501 );
not ( w_17501 , w_17502 );
and ( \7120_b0 , \7118_b0 , w_17503 );
and ( w_17502 ,  , w_17503 );
buf ( w_17501 , \7119_b1 );
not ( w_17501 , w_17504 );
not (  , w_17505 );
and ( w_17504 , w_17505 , \7119_b0 );
or ( \7121_b1 , \7113_b1 , \7092_b1 );
not ( \7092_b1 , w_17506 );
and ( \7121_b0 , \7113_b0 , w_17507 );
and ( w_17506 , w_17507 , \7092_b0 );
buf ( \7122_b1 , \7121_b1 );
not ( \7122_b1 , w_17508 );
not ( \7122_b0 , w_17509 );
and ( w_17508 , w_17509 , \7121_b0 );
or ( \7123_b1 , \7110_b1 , \7122_b1 );
not ( \7122_b1 , w_17510 );
and ( \7123_b0 , \7110_b0 , w_17511 );
and ( w_17510 , w_17511 , \7122_b0 );
or ( \7124_b1 , \7120_b1 , w_17512 );
xor ( \7124_b0 , \7120_b0 , w_17514 );
not ( w_17514 , w_17515 );
and ( w_17515 , w_17512 , w_17513 );
buf ( w_17512 , \7123_b1 );
not ( w_17512 , w_17516 );
not ( w_17513 , w_17517 );
and ( w_17516 , w_17517 , \7123_b0 );
or ( \7125_b1 , \7106_b1 , \7124_b1 );
not ( \7124_b1 , w_17518 );
and ( \7125_b0 , \7106_b0 , w_17519 );
and ( w_17518 , w_17519 , \7124_b0 );
or ( \7126_b1 , \7089_b1 , \7124_b1 );
not ( \7124_b1 , w_17520 );
and ( \7126_b0 , \7089_b0 , w_17521 );
and ( w_17520 , w_17521 , \7124_b0 );
or ( \7128_b1 , \7071_b1 , \7127_b1 );
not ( \7127_b1 , w_17522 );
and ( \7128_b0 , \7071_b0 , w_17523 );
and ( w_17522 , w_17523 , \7127_b0 );
or ( \7129_b1 , \7016_b1 , \7127_b1 );
not ( \7127_b1 , w_17524 );
and ( \7129_b0 , \7016_b0 , w_17525 );
and ( w_17524 , w_17525 , \7127_b0 );
or ( \7131_b1 , \5169_b1 , \5640_b1 );
xor ( \7131_b0 , \5169_b0 , w_17526 );
not ( w_17526 , w_17527 );
and ( w_17527 , \5640_b1 , \5640_b0 );
buf ( \7132_b1 , \7131_b1 );
buf ( \7132_b0 , \7131_b0 );
buf ( \7133_b1 , \7132_b1 );
buf ( \7133_b0 , \7132_b0 );
or ( \7134_b1 , \5224_b1 , \5638_b1 );
xor ( \7134_b0 , \5224_b0 , w_17528 );
not ( w_17528 , w_17529 );
and ( w_17529 , \5638_b1 , \5638_b0 );
buf ( \7135_b1 , \7134_b1 );
buf ( \7135_b0 , \7134_b0 );
buf ( \7136_b1 , \7135_b1 );
buf ( \7136_b0 , \7135_b0 );
or ( \7137_b1 , \7133_b1 , \7136_b1 );
xor ( \7137_b0 , \7133_b0 , w_17530 );
not ( w_17530 , w_17531 );
and ( w_17531 , \7136_b1 , \7136_b0 );
or ( \7138_b1 , \7136_b1 , \7110_b1 );
xor ( \7138_b0 , \7136_b0 , w_17532 );
not ( w_17532 , w_17533 );
and ( w_17533 , \7110_b1 , \7110_b0 );
buf ( \7139_b1 , \7138_b1 );
not ( \7139_b1 , w_17534 );
not ( \7139_b0 , w_17535 );
and ( w_17534 , w_17535 , \7138_b0 );
or ( \7140_b1 , \7137_b1 , \7139_b1 );
not ( \7139_b1 , w_17536 );
and ( \7140_b0 , \7137_b0 , w_17537 );
and ( w_17536 , w_17537 , \7139_b0 );
or ( \7141_b1 , \5967_b1 , \7140_b1 );
not ( \7140_b1 , w_17538 );
and ( \7141_b0 , \5967_b0 , w_17539 );
and ( w_17538 , w_17539 , \7140_b0 );
or ( \7142_b1 , \5979_b1 , \7138_b1 );
not ( \7138_b1 , w_17540 );
and ( \7142_b0 , \5979_b0 , w_17541 );
and ( w_17540 , w_17541 , \7138_b0 );
or ( \7143_b1 , \7141_b1 , w_17543 );
not ( w_17543 , w_17544 );
and ( \7143_b0 , \7141_b0 , w_17545 );
and ( w_17544 ,  , w_17545 );
buf ( w_17543 , \7142_b1 );
not ( w_17543 , w_17546 );
not (  , w_17547 );
and ( w_17546 , w_17547 , \7142_b0 );
or ( \7144_b1 , \7136_b1 , \7110_b1 );
not ( \7110_b1 , w_17548 );
and ( \7144_b0 , \7136_b0 , w_17549 );
and ( w_17548 , w_17549 , \7110_b0 );
buf ( \7145_b1 , \7144_b1 );
not ( \7145_b1 , w_17550 );
not ( \7145_b0 , w_17551 );
and ( w_17550 , w_17551 , \7144_b0 );
or ( \7146_b1 , \7133_b1 , \7145_b1 );
not ( \7145_b1 , w_17552 );
and ( \7146_b0 , \7133_b0 , w_17553 );
and ( w_17552 , w_17553 , \7145_b0 );
or ( \7147_b1 , \7143_b1 , w_17554 );
xor ( \7147_b0 , \7143_b0 , w_17556 );
not ( w_17556 , w_17557 );
and ( w_17557 , w_17554 , w_17555 );
buf ( w_17554 , \7146_b1 );
not ( w_17554 , w_17558 );
not ( w_17555 , w_17559 );
and ( w_17558 , w_17559 , \7146_b0 );
or ( \7148_b1 , \5102_b1 , \5644_b1 );
xor ( \7148_b0 , \5102_b0 , w_17560 );
not ( w_17560 , w_17561 );
and ( w_17561 , \5644_b1 , \5644_b0 );
buf ( \7149_b1 , \7148_b1 );
buf ( \7149_b0 , \7148_b0 );
buf ( \7150_b1 , \7149_b1 );
buf ( \7150_b0 , \7149_b0 );
or ( \7151_b1 , \5110_b1 , \5642_b1 );
xor ( \7151_b0 , \5110_b0 , w_17562 );
not ( w_17562 , w_17563 );
and ( w_17563 , \5642_b1 , \5642_b0 );
buf ( \7152_b1 , \7151_b1 );
buf ( \7152_b0 , \7151_b0 );
buf ( \7153_b1 , \7152_b1 );
buf ( \7153_b0 , \7152_b0 );
or ( \7154_b1 , \7150_b1 , \7153_b1 );
xor ( \7154_b0 , \7150_b0 , w_17564 );
not ( w_17564 , w_17565 );
and ( w_17565 , \7153_b1 , \7153_b0 );
or ( \7155_b1 , \7153_b1 , \7133_b1 );
xor ( \7155_b0 , \7153_b0 , w_17566 );
not ( w_17566 , w_17567 );
and ( w_17567 , \7133_b1 , \7133_b0 );
buf ( \7156_b1 , \7155_b1 );
not ( \7156_b1 , w_17568 );
not ( \7156_b0 , w_17569 );
and ( w_17568 , w_17569 , \7155_b0 );
or ( \7157_b1 , \7154_b1 , \7156_b1 );
not ( \7156_b1 , w_17570 );
and ( \7157_b0 , \7154_b0 , w_17571 );
and ( w_17570 , w_17571 , \7156_b0 );
or ( \7158_b1 , \5986_b1 , \7157_b1 );
not ( \7157_b1 , w_17572 );
and ( \7158_b0 , \5986_b0 , w_17573 );
and ( w_17572 , w_17573 , \7157_b0 );
or ( \7159_b1 , \5998_b1 , \7155_b1 );
not ( \7155_b1 , w_17574 );
and ( \7159_b0 , \5998_b0 , w_17575 );
and ( w_17574 , w_17575 , \7155_b0 );
or ( \7160_b1 , \7158_b1 , w_17577 );
not ( w_17577 , w_17578 );
and ( \7160_b0 , \7158_b0 , w_17579 );
and ( w_17578 ,  , w_17579 );
buf ( w_17577 , \7159_b1 );
not ( w_17577 , w_17580 );
not (  , w_17581 );
and ( w_17580 , w_17581 , \7159_b0 );
or ( \7161_b1 , \7153_b1 , \7133_b1 );
not ( \7133_b1 , w_17582 );
and ( \7161_b0 , \7153_b0 , w_17583 );
and ( w_17582 , w_17583 , \7133_b0 );
buf ( \7162_b1 , \7161_b1 );
not ( \7162_b1 , w_17584 );
not ( \7162_b0 , w_17585 );
and ( w_17584 , w_17585 , \7161_b0 );
or ( \7163_b1 , \7150_b1 , \7162_b1 );
not ( \7162_b1 , w_17586 );
and ( \7163_b0 , \7150_b0 , w_17587 );
and ( w_17586 , w_17587 , \7162_b0 );
or ( \7164_b1 , \7160_b1 , w_17588 );
xor ( \7164_b0 , \7160_b0 , w_17590 );
not ( w_17590 , w_17591 );
and ( w_17591 , w_17588 , w_17589 );
buf ( w_17588 , \7163_b1 );
not ( w_17588 , w_17592 );
not ( w_17589 , w_17593 );
and ( w_17592 , w_17593 , \7163_b0 );
or ( \7165_b1 , \7147_b1 , \7164_b1 );
not ( \7164_b1 , w_17594 );
and ( \7165_b0 , \7147_b0 , w_17595 );
and ( w_17594 , w_17595 , \7164_b0 );
or ( \7166_b1 , \4943_b1 , \5648_b1 );
xor ( \7166_b0 , \4943_b0 , w_17596 );
not ( w_17596 , w_17597 );
and ( w_17597 , \5648_b1 , \5648_b0 );
buf ( \7167_b1 , \7166_b1 );
buf ( \7167_b0 , \7166_b0 );
buf ( \7168_b1 , \7167_b1 );
buf ( \7168_b0 , \7167_b0 );
or ( \7169_b1 , \5023_b1 , \5646_b1 );
xor ( \7169_b0 , \5023_b0 , w_17598 );
not ( w_17598 , w_17599 );
and ( w_17599 , \5646_b1 , \5646_b0 );
buf ( \7170_b1 , \7169_b1 );
buf ( \7170_b0 , \7169_b0 );
buf ( \7171_b1 , \7170_b1 );
buf ( \7171_b0 , \7170_b0 );
or ( \7172_b1 , \7168_b1 , \7171_b1 );
xor ( \7172_b0 , \7168_b0 , w_17600 );
not ( w_17600 , w_17601 );
and ( w_17601 , \7171_b1 , \7171_b0 );
or ( \7173_b1 , \7171_b1 , \7150_b1 );
xor ( \7173_b0 , \7171_b0 , w_17602 );
not ( w_17602 , w_17603 );
and ( w_17603 , \7150_b1 , \7150_b0 );
buf ( \7174_b1 , \7173_b1 );
not ( \7174_b1 , w_17604 );
not ( \7174_b0 , w_17605 );
and ( w_17604 , w_17605 , \7173_b0 );
or ( \7175_b1 , \7172_b1 , \7174_b1 );
not ( \7174_b1 , w_17606 );
and ( \7175_b0 , \7172_b0 , w_17607 );
and ( w_17606 , w_17607 , \7174_b0 );
or ( \7176_b1 , \6006_b1 , \7175_b1 );
not ( \7175_b1 , w_17608 );
and ( \7176_b0 , \6006_b0 , w_17609 );
and ( w_17608 , w_17609 , \7175_b0 );
or ( \7177_b1 , \6018_b1 , \7173_b1 );
not ( \7173_b1 , w_17610 );
and ( \7177_b0 , \6018_b0 , w_17611 );
and ( w_17610 , w_17611 , \7173_b0 );
or ( \7178_b1 , \7176_b1 , w_17613 );
not ( w_17613 , w_17614 );
and ( \7178_b0 , \7176_b0 , w_17615 );
and ( w_17614 ,  , w_17615 );
buf ( w_17613 , \7177_b1 );
not ( w_17613 , w_17616 );
not (  , w_17617 );
and ( w_17616 , w_17617 , \7177_b0 );
or ( \7179_b1 , \7171_b1 , \7150_b1 );
not ( \7150_b1 , w_17618 );
and ( \7179_b0 , \7171_b0 , w_17619 );
and ( w_17618 , w_17619 , \7150_b0 );
buf ( \7180_b1 , \7179_b1 );
not ( \7180_b1 , w_17620 );
not ( \7180_b0 , w_17621 );
and ( w_17620 , w_17621 , \7179_b0 );
or ( \7181_b1 , \7168_b1 , \7180_b1 );
not ( \7180_b1 , w_17622 );
and ( \7181_b0 , \7168_b0 , w_17623 );
and ( w_17622 , w_17623 , \7180_b0 );
or ( \7182_b1 , \7178_b1 , w_17624 );
xor ( \7182_b0 , \7178_b0 , w_17626 );
not ( w_17626 , w_17627 );
and ( w_17627 , w_17624 , w_17625 );
buf ( w_17624 , \7181_b1 );
not ( w_17624 , w_17628 );
not ( w_17625 , w_17629 );
and ( w_17628 , w_17629 , \7181_b0 );
or ( \7183_b1 , \7164_b1 , \7182_b1 );
not ( \7182_b1 , w_17630 );
and ( \7183_b0 , \7164_b0 , w_17631 );
and ( w_17630 , w_17631 , \7182_b0 );
or ( \7184_b1 , \7147_b1 , \7182_b1 );
not ( \7182_b1 , w_17632 );
and ( \7184_b0 , \7147_b0 , w_17633 );
and ( w_17632 , w_17633 , \7182_b0 );
or ( \7186_b1 , \4848_b1 , \5650_b1 );
xor ( \7186_b0 , \4848_b0 , w_17634 );
not ( w_17634 , w_17635 );
and ( w_17635 , \5650_b1 , \5650_b0 );
buf ( \7187_b1 , \7186_b1 );
buf ( \7187_b0 , \7186_b0 );
buf ( \7188_b1 , \7187_b1 );
buf ( \7188_b0 , \7187_b0 );
or ( \7189_b1 , \6821_b1 , \7188_b1 );
xor ( \7189_b0 , \6821_b0 , w_17636 );
not ( w_17636 , w_17637 );
and ( w_17637 , \7188_b1 , \7188_b0 );
or ( \7190_b1 , \7188_b1 , \7168_b1 );
xor ( \7190_b0 , \7188_b0 , w_17638 );
not ( w_17638 , w_17639 );
and ( w_17639 , \7168_b1 , \7168_b0 );
buf ( \7191_b1 , \7190_b1 );
not ( \7191_b1 , w_17640 );
not ( \7191_b0 , w_17641 );
and ( w_17640 , w_17641 , \7190_b0 );
or ( \7192_b1 , \7189_b1 , \7191_b1 );
not ( \7191_b1 , w_17642 );
and ( \7192_b0 , \7189_b0 , w_17643 );
and ( w_17642 , w_17643 , \7191_b0 );
or ( \7193_b1 , \6029_b1 , \7192_b1 );
not ( \7192_b1 , w_17644 );
and ( \7193_b0 , \6029_b0 , w_17645 );
and ( w_17644 , w_17645 , \7192_b0 );
or ( \7194_b1 , \6041_b1 , \7190_b1 );
not ( \7190_b1 , w_17646 );
and ( \7194_b0 , \6041_b0 , w_17647 );
and ( w_17646 , w_17647 , \7190_b0 );
or ( \7195_b1 , \7193_b1 , w_17649 );
not ( w_17649 , w_17650 );
and ( \7195_b0 , \7193_b0 , w_17651 );
and ( w_17650 ,  , w_17651 );
buf ( w_17649 , \7194_b1 );
not ( w_17649 , w_17652 );
not (  , w_17653 );
and ( w_17652 , w_17653 , \7194_b0 );
or ( \7196_b1 , \7188_b1 , \7168_b1 );
not ( \7168_b1 , w_17654 );
and ( \7196_b0 , \7188_b0 , w_17655 );
and ( w_17654 , w_17655 , \7168_b0 );
buf ( \7197_b1 , \7196_b1 );
not ( \7197_b1 , w_17656 );
not ( \7197_b0 , w_17657 );
and ( w_17656 , w_17657 , \7196_b0 );
or ( \7198_b1 , \6821_b1 , \7197_b1 );
not ( \7197_b1 , w_17658 );
and ( \7198_b0 , \6821_b0 , w_17659 );
and ( w_17658 , w_17659 , \7197_b0 );
or ( \7199_b1 , \7195_b1 , w_17660 );
xor ( \7199_b0 , \7195_b0 , w_17662 );
not ( w_17662 , w_17663 );
and ( w_17663 , w_17660 , w_17661 );
buf ( w_17660 , \7198_b1 );
not ( w_17660 , w_17664 );
not ( w_17661 , w_17665 );
and ( w_17664 , w_17665 , \7198_b0 );
or ( \7200_b1 , \5747_b1 , \6818_b1 );
xor ( \7200_b0 , \5747_b0 , w_17666 );
not ( w_17666 , w_17667 );
and ( w_17667 , \6818_b1 , \6818_b0 );
or ( \7201_b1 , \6818_b1 , \6821_b1 );
xor ( \7201_b0 , \6818_b0 , w_17668 );
not ( w_17668 , w_17669 );
and ( w_17669 , \6821_b1 , \6821_b0 );
buf ( \7202_b1 , \7201_b1 );
not ( \7202_b1 , w_17670 );
not ( \7202_b0 , w_17671 );
and ( w_17670 , w_17671 , \7201_b0 );
or ( \7203_b1 , \7200_b1 , \7202_b1 );
not ( \7202_b1 , w_17672 );
and ( \7203_b0 , \7200_b0 , w_17673 );
and ( w_17672 , w_17673 , \7202_b0 );
or ( \7204_b1 , \6048_b1 , \7203_b1 );
not ( \7203_b1 , w_17674 );
and ( \7204_b0 , \6048_b0 , w_17675 );
and ( w_17674 , w_17675 , \7203_b0 );
or ( \7205_b1 , \6057_b1 , \7201_b1 );
not ( \7201_b1 , w_17676 );
and ( \7205_b0 , \6057_b0 , w_17677 );
and ( w_17676 , w_17677 , \7201_b0 );
or ( \7206_b1 , \7204_b1 , w_17679 );
not ( w_17679 , w_17680 );
and ( \7206_b0 , \7204_b0 , w_17681 );
and ( w_17680 ,  , w_17681 );
buf ( w_17679 , \7205_b1 );
not ( w_17679 , w_17682 );
not (  , w_17683 );
and ( w_17682 , w_17683 , \7205_b0 );
or ( \7207_b1 , \7206_b1 , w_17684 );
xor ( \7207_b0 , \7206_b0 , w_17686 );
not ( w_17686 , w_17687 );
and ( w_17687 , w_17684 , w_17685 );
buf ( w_17684 , \6824_b1 );
not ( w_17684 , w_17688 );
not ( w_17685 , w_17689 );
and ( w_17688 , w_17689 , \6824_b0 );
or ( \7208_b1 , \7199_b1 , \7207_b1 );
not ( \7207_b1 , w_17690 );
and ( \7208_b0 , \7199_b0 , w_17691 );
and ( w_17690 , w_17691 , \7207_b0 );
or ( \7209_b1 , \6065_b1 , w_17693 );
not ( w_17693 , w_17694 );
and ( \7209_b0 , \6065_b0 , w_17695 );
and ( w_17694 ,  , w_17695 );
buf ( w_17693 , \5748_b1 );
not ( w_17693 , w_17696 );
not (  , w_17697 );
and ( w_17696 , w_17697 , \5748_b0 );
or ( \7210_b1 , \7209_b1 , w_17698 );
xor ( \7210_b0 , \7209_b0 , w_17700 );
not ( w_17700 , w_17701 );
and ( w_17701 , w_17698 , w_17699 );
buf ( w_17698 , \5755_b1 );
not ( w_17698 , w_17702 );
not ( w_17699 , w_17703 );
and ( w_17702 , w_17703 , \5755_b0 );
or ( \7211_b1 , \7207_b1 , \7210_b1 );
not ( \7210_b1 , w_17704 );
and ( \7211_b0 , \7207_b0 , w_17705 );
and ( w_17704 , w_17705 , \7210_b0 );
or ( \7212_b1 , \7199_b1 , \7210_b1 );
not ( \7210_b1 , w_17706 );
and ( \7212_b0 , \7199_b0 , w_17707 );
and ( w_17706 , w_17707 , \7210_b0 );
or ( \7214_b1 , \7185_b1 , \7213_b1 );
not ( \7213_b1 , w_17708 );
and ( \7214_b0 , \7185_b0 , w_17709 );
and ( w_17708 , w_17709 , \7213_b0 );
or ( \7215_b1 , \6057_b1 , \7203_b1 );
not ( \7203_b1 , w_17710 );
and ( \7215_b0 , \6057_b0 , w_17711 );
and ( w_17710 , w_17711 , \7203_b0 );
or ( \7216_b1 , \6029_b1 , \7201_b1 );
not ( \7201_b1 , w_17712 );
and ( \7216_b0 , \6029_b0 , w_17713 );
and ( w_17712 , w_17713 , \7201_b0 );
or ( \7217_b1 , \7215_b1 , w_17715 );
not ( w_17715 , w_17716 );
and ( \7217_b0 , \7215_b0 , w_17717 );
and ( w_17716 ,  , w_17717 );
buf ( w_17715 , \7216_b1 );
not ( w_17715 , w_17718 );
not (  , w_17719 );
and ( w_17718 , w_17719 , \7216_b0 );
or ( \7218_b1 , \7217_b1 , w_17720 );
xor ( \7218_b0 , \7217_b0 , w_17722 );
not ( w_17722 , w_17723 );
and ( w_17723 , w_17720 , w_17721 );
buf ( w_17720 , \6824_b1 );
not ( w_17720 , w_17724 );
not ( w_17721 , w_17725 );
and ( w_17724 , w_17725 , \6824_b0 );
or ( \7219_b1 , \7213_b1 , \7218_b1 );
not ( \7218_b1 , w_17726 );
and ( \7219_b0 , \7213_b0 , w_17727 );
and ( w_17726 , w_17727 , \7218_b0 );
or ( \7220_b1 , \7185_b1 , \7218_b1 );
not ( \7218_b1 , w_17728 );
and ( \7220_b0 , \7185_b0 , w_17729 );
and ( w_17728 , w_17729 , \7218_b0 );
or ( \7222_b1 , \7130_b1 , \7221_b1 );
not ( \7221_b1 , w_17730 );
and ( \7222_b0 , \7130_b0 , w_17731 );
and ( w_17730 , w_17731 , \7221_b0 );
or ( \7223_b1 , \6065_b1 , \5750_b1 );
not ( \5750_b1 , w_17732 );
and ( \7223_b0 , \6065_b0 , w_17733 );
and ( w_17732 , w_17733 , \5750_b0 );
or ( \7224_b1 , \6048_b1 , \5748_b1 );
not ( \5748_b1 , w_17734 );
and ( \7224_b0 , \6048_b0 , w_17735 );
and ( w_17734 , w_17735 , \5748_b0 );
or ( \7225_b1 , \7223_b1 , w_17737 );
not ( w_17737 , w_17738 );
and ( \7225_b0 , \7223_b0 , w_17739 );
and ( w_17738 ,  , w_17739 );
buf ( w_17737 , \7224_b1 );
not ( w_17737 , w_17740 );
not (  , w_17741 );
and ( w_17740 , w_17741 , \7224_b0 );
or ( \7226_b1 , \7225_b1 , w_17742 );
xor ( \7226_b0 , \7225_b0 , w_17744 );
not ( w_17744 , w_17745 );
and ( w_17745 , w_17742 , w_17743 );
buf ( w_17742 , \5755_b1 );
not ( w_17742 , w_17746 );
not ( w_17743 , w_17747 );
and ( w_17746 , w_17747 , \5755_b0 );
or ( \7227_b1 , \5998_b1 , \7157_b1 );
not ( \7157_b1 , w_17748 );
and ( \7227_b0 , \5998_b0 , w_17749 );
and ( w_17748 , w_17749 , \7157_b0 );
or ( \7228_b1 , \5967_b1 , \7155_b1 );
not ( \7155_b1 , w_17750 );
and ( \7228_b0 , \5967_b0 , w_17751 );
and ( w_17750 , w_17751 , \7155_b0 );
or ( \7229_b1 , \7227_b1 , w_17753 );
not ( w_17753 , w_17754 );
and ( \7229_b0 , \7227_b0 , w_17755 );
and ( w_17754 ,  , w_17755 );
buf ( w_17753 , \7228_b1 );
not ( w_17753 , w_17756 );
not (  , w_17757 );
and ( w_17756 , w_17757 , \7228_b0 );
or ( \7230_b1 , \7229_b1 , w_17758 );
xor ( \7230_b0 , \7229_b0 , w_17760 );
not ( w_17760 , w_17761 );
and ( w_17761 , w_17758 , w_17759 );
buf ( w_17758 , \7163_b1 );
not ( w_17758 , w_17762 );
not ( w_17759 , w_17763 );
and ( w_17762 , w_17763 , \7163_b0 );
or ( \7231_b1 , \6018_b1 , \7175_b1 );
not ( \7175_b1 , w_17764 );
and ( \7231_b0 , \6018_b0 , w_17765 );
and ( w_17764 , w_17765 , \7175_b0 );
or ( \7232_b1 , \5986_b1 , \7173_b1 );
not ( \7173_b1 , w_17766 );
and ( \7232_b0 , \5986_b0 , w_17767 );
and ( w_17766 , w_17767 , \7173_b0 );
or ( \7233_b1 , \7231_b1 , w_17769 );
not ( w_17769 , w_17770 );
and ( \7233_b0 , \7231_b0 , w_17771 );
and ( w_17770 ,  , w_17771 );
buf ( w_17769 , \7232_b1 );
not ( w_17769 , w_17772 );
not (  , w_17773 );
and ( w_17772 , w_17773 , \7232_b0 );
or ( \7234_b1 , \7233_b1 , w_17774 );
xor ( \7234_b0 , \7233_b0 , w_17776 );
not ( w_17776 , w_17777 );
and ( w_17777 , w_17774 , w_17775 );
buf ( w_17774 , \7181_b1 );
not ( w_17774 , w_17778 );
not ( w_17775 , w_17779 );
and ( w_17778 , w_17779 , \7181_b0 );
or ( \7235_b1 , \7230_b1 , \7234_b1 );
xor ( \7235_b0 , \7230_b0 , w_17780 );
not ( w_17780 , w_17781 );
and ( w_17781 , \7234_b1 , \7234_b0 );
or ( \7236_b1 , \6041_b1 , \7192_b1 );
not ( \7192_b1 , w_17782 );
and ( \7236_b0 , \6041_b0 , w_17783 );
and ( w_17782 , w_17783 , \7192_b0 );
or ( \7237_b1 , \6006_b1 , \7190_b1 );
not ( \7190_b1 , w_17784 );
and ( \7237_b0 , \6006_b0 , w_17785 );
and ( w_17784 , w_17785 , \7190_b0 );
or ( \7238_b1 , \7236_b1 , w_17787 );
not ( w_17787 , w_17788 );
and ( \7238_b0 , \7236_b0 , w_17789 );
and ( w_17788 ,  , w_17789 );
buf ( w_17787 , \7237_b1 );
not ( w_17787 , w_17790 );
not (  , w_17791 );
and ( w_17790 , w_17791 , \7237_b0 );
or ( \7239_b1 , \7238_b1 , w_17792 );
xor ( \7239_b0 , \7238_b0 , w_17794 );
not ( w_17794 , w_17795 );
and ( w_17795 , w_17792 , w_17793 );
buf ( w_17792 , \7198_b1 );
not ( w_17792 , w_17796 );
not ( w_17793 , w_17797 );
and ( w_17796 , w_17797 , \7198_b0 );
or ( \7240_b1 , \7235_b1 , \7239_b1 );
xor ( \7240_b0 , \7235_b0 , w_17798 );
not ( w_17798 , w_17799 );
and ( w_17799 , \7239_b1 , \7239_b0 );
or ( \7241_b1 , \7226_b1 , \7240_b1 );
not ( \7240_b1 , w_17800 );
and ( \7241_b0 , \7226_b0 , w_17801 );
and ( w_17800 , w_17801 , \7240_b0 );
or ( \7242_b1 , \5937_b1 , \7099_b1 );
not ( \7099_b1 , w_17802 );
and ( \7242_b0 , \5937_b0 , w_17803 );
and ( w_17802 , w_17803 , \7099_b0 );
or ( \7243_b1 , \5906_b1 , \7097_b1 );
not ( \7097_b1 , w_17804 );
and ( \7243_b0 , \5906_b0 , w_17805 );
and ( w_17804 , w_17805 , \7097_b0 );
or ( \7244_b1 , \7242_b1 , w_17807 );
not ( w_17807 , w_17808 );
and ( \7244_b0 , \7242_b0 , w_17809 );
and ( w_17808 ,  , w_17809 );
buf ( w_17807 , \7243_b1 );
not ( w_17807 , w_17810 );
not (  , w_17811 );
and ( w_17810 , w_17811 , \7243_b0 );
or ( \7245_b1 , \7244_b1 , w_17812 );
xor ( \7245_b0 , \7244_b0 , w_17814 );
not ( w_17814 , w_17815 );
and ( w_17815 , w_17812 , w_17813 );
buf ( w_17812 , \7105_b1 );
not ( w_17812 , w_17816 );
not ( w_17813 , w_17817 );
and ( w_17816 , w_17817 , \7105_b0 );
or ( \7246_b1 , \5957_b1 , \7117_b1 );
not ( \7117_b1 , w_17818 );
and ( \7246_b0 , \5957_b0 , w_17819 );
and ( w_17818 , w_17819 , \7117_b0 );
or ( \7247_b1 , \5925_b1 , \7115_b1 );
not ( \7115_b1 , w_17820 );
and ( \7247_b0 , \5925_b0 , w_17821 );
and ( w_17820 , w_17821 , \7115_b0 );
or ( \7248_b1 , \7246_b1 , w_17823 );
not ( w_17823 , w_17824 );
and ( \7248_b0 , \7246_b0 , w_17825 );
and ( w_17824 ,  , w_17825 );
buf ( w_17823 , \7247_b1 );
not ( w_17823 , w_17826 );
not (  , w_17827 );
and ( w_17826 , w_17827 , \7247_b0 );
or ( \7249_b1 , \7248_b1 , w_17828 );
xor ( \7249_b0 , \7248_b0 , w_17830 );
not ( w_17830 , w_17831 );
and ( w_17831 , w_17828 , w_17829 );
buf ( w_17828 , \7123_b1 );
not ( w_17828 , w_17832 );
not ( w_17829 , w_17833 );
and ( w_17832 , w_17833 , \7123_b0 );
or ( \7250_b1 , \7245_b1 , \7249_b1 );
xor ( \7250_b0 , \7245_b0 , w_17834 );
not ( w_17834 , w_17835 );
and ( w_17835 , \7249_b1 , \7249_b0 );
or ( \7251_b1 , \5979_b1 , \7140_b1 );
not ( \7140_b1 , w_17836 );
and ( \7251_b0 , \5979_b0 , w_17837 );
and ( w_17836 , w_17837 , \7140_b0 );
or ( \7252_b1 , \5945_b1 , \7138_b1 );
not ( \7138_b1 , w_17838 );
and ( \7252_b0 , \5945_b0 , w_17839 );
and ( w_17838 , w_17839 , \7138_b0 );
or ( \7253_b1 , \7251_b1 , w_17841 );
not ( w_17841 , w_17842 );
and ( \7253_b0 , \7251_b0 , w_17843 );
and ( w_17842 ,  , w_17843 );
buf ( w_17841 , \7252_b1 );
not ( w_17841 , w_17844 );
not (  , w_17845 );
and ( w_17844 , w_17845 , \7252_b0 );
or ( \7254_b1 , \7253_b1 , w_17846 );
xor ( \7254_b0 , \7253_b0 , w_17848 );
not ( w_17848 , w_17849 );
and ( w_17849 , w_17846 , w_17847 );
buf ( w_17846 , \7146_b1 );
not ( w_17846 , w_17850 );
not ( w_17847 , w_17851 );
and ( w_17850 , w_17851 , \7146_b0 );
or ( \7255_b1 , \7250_b1 , \7254_b1 );
xor ( \7255_b0 , \7250_b0 , w_17852 );
not ( w_17852 , w_17853 );
and ( w_17853 , \7254_b1 , \7254_b0 );
or ( \7256_b1 , \7240_b1 , \7255_b1 );
not ( \7255_b1 , w_17854 );
and ( \7256_b0 , \7240_b0 , w_17855 );
and ( w_17854 , w_17855 , \7255_b0 );
or ( \7257_b1 , \7226_b1 , \7255_b1 );
not ( \7255_b1 , w_17856 );
and ( \7257_b0 , \7226_b0 , w_17857 );
and ( w_17856 , w_17857 , \7255_b0 );
or ( \7259_b1 , \7221_b1 , \7258_b1 );
not ( \7258_b1 , w_17858 );
and ( \7259_b0 , \7221_b0 , w_17859 );
and ( w_17858 , w_17859 , \7258_b0 );
or ( \7260_b1 , \7130_b1 , \7258_b1 );
not ( \7258_b1 , w_17860 );
and ( \7260_b0 , \7130_b0 , w_17861 );
and ( w_17860 , w_17861 , \7258_b0 );
or ( \7262_b1 , \5780_b1 , \6991_b1 );
not ( \6991_b1 , w_17862 );
and ( \7262_b0 , \5780_b0 , w_17863 );
and ( w_17862 , w_17863 , \6991_b0 );
or ( \7263_b1 , \5792_b1 , \6988_b1 );
not ( \6988_b1 , w_17864 );
and ( \7263_b0 , \5792_b0 , w_17865 );
and ( w_17864 , w_17865 , \6988_b0 );
or ( \7264_b1 , \7262_b1 , w_17867 );
not ( w_17867 , w_17868 );
and ( \7264_b0 , \7262_b0 , w_17869 );
and ( w_17868 ,  , w_17869 );
buf ( w_17867 , \7263_b1 );
not ( w_17867 , w_17870 );
not (  , w_17871 );
and ( w_17870 , w_17871 , \7263_b0 );
or ( \7265_b1 , \7264_b1 , w_17872 );
xor ( \7265_b0 , \7264_b0 , w_17874 );
not ( w_17874 , w_17875 );
and ( w_17875 , w_17872 , w_17873 );
buf ( w_17872 , \6985_b1 );
not ( w_17872 , w_17876 );
not ( w_17873 , w_17877 );
and ( w_17876 , w_17877 , \6985_b0 );
or ( \7266_b1 , \5775_b1 , \7265_b1 );
xor ( \7266_b0 , \5775_b0 , w_17878 );
not ( w_17878 , w_17879 );
and ( w_17879 , \7265_b1 , \7265_b0 );
or ( \7267_b1 , \5799_b1 , \7006_b1 );
not ( \7006_b1 , w_17880 );
and ( \7267_b0 , \5799_b0 , w_17881 );
and ( w_17880 , w_17881 , \7006_b0 );
or ( \7268_b1 , \5811_b1 , \7004_b1 );
not ( \7004_b1 , w_17882 );
and ( \7268_b0 , \5811_b0 , w_17883 );
and ( w_17882 , w_17883 , \7004_b0 );
or ( \7269_b1 , \7267_b1 , w_17885 );
not ( w_17885 , w_17886 );
and ( \7269_b0 , \7267_b0 , w_17887 );
and ( w_17886 ,  , w_17887 );
buf ( w_17885 , \7268_b1 );
not ( w_17885 , w_17888 );
not (  , w_17889 );
and ( w_17888 , w_17889 , \7268_b0 );
or ( \7270_b1 , \7269_b1 , w_17890 );
xor ( \7270_b0 , \7269_b0 , w_17892 );
not ( w_17892 , w_17893 );
and ( w_17893 , w_17890 , w_17891 );
buf ( w_17890 , \7012_b1 );
not ( w_17890 , w_17894 );
not ( w_17891 , w_17895 );
and ( w_17894 , w_17895 , \7012_b0 );
or ( \7271_b1 , \7266_b1 , \7270_b1 );
xor ( \7271_b0 , \7266_b0 , w_17896 );
not ( w_17896 , w_17897 );
and ( w_17897 , \7270_b1 , \7270_b0 );
or ( \7272_b1 , \5945_b1 , \7140_b1 );
not ( \7140_b1 , w_17898 );
and ( \7272_b0 , \5945_b0 , w_17899 );
and ( w_17898 , w_17899 , \7140_b0 );
or ( \7273_b1 , \5957_b1 , \7138_b1 );
not ( \7138_b1 , w_17900 );
and ( \7273_b0 , \5957_b0 , w_17901 );
and ( w_17900 , w_17901 , \7138_b0 );
or ( \7274_b1 , \7272_b1 , w_17903 );
not ( w_17903 , w_17904 );
and ( \7274_b0 , \7272_b0 , w_17905 );
and ( w_17904 ,  , w_17905 );
buf ( w_17903 , \7273_b1 );
not ( w_17903 , w_17906 );
not (  , w_17907 );
and ( w_17906 , w_17907 , \7273_b0 );
or ( \7275_b1 , \7274_b1 , w_17908 );
xor ( \7275_b0 , \7274_b0 , w_17910 );
not ( w_17910 , w_17911 );
and ( w_17911 , w_17908 , w_17909 );
buf ( w_17908 , \7146_b1 );
not ( w_17908 , w_17912 );
not ( w_17909 , w_17913 );
and ( w_17912 , w_17913 , \7146_b0 );
or ( \7276_b1 , \5967_b1 , \7157_b1 );
not ( \7157_b1 , w_17914 );
and ( \7276_b0 , \5967_b0 , w_17915 );
and ( w_17914 , w_17915 , \7157_b0 );
or ( \7277_b1 , \5979_b1 , \7155_b1 );
not ( \7155_b1 , w_17916 );
and ( \7277_b0 , \5979_b0 , w_17917 );
and ( w_17916 , w_17917 , \7155_b0 );
or ( \7278_b1 , \7276_b1 , w_17919 );
not ( w_17919 , w_17920 );
and ( \7278_b0 , \7276_b0 , w_17921 );
and ( w_17920 ,  , w_17921 );
buf ( w_17919 , \7277_b1 );
not ( w_17919 , w_17922 );
not (  , w_17923 );
and ( w_17922 , w_17923 , \7277_b0 );
or ( \7279_b1 , \7278_b1 , w_17924 );
xor ( \7279_b0 , \7278_b0 , w_17926 );
not ( w_17926 , w_17927 );
and ( w_17927 , w_17924 , w_17925 );
buf ( w_17924 , \7163_b1 );
not ( w_17924 , w_17928 );
not ( w_17925 , w_17929 );
and ( w_17928 , w_17929 , \7163_b0 );
or ( \7280_b1 , \7275_b1 , \7279_b1 );
xor ( \7280_b0 , \7275_b0 , w_17930 );
not ( w_17930 , w_17931 );
and ( w_17931 , \7279_b1 , \7279_b0 );
or ( \7281_b1 , \5986_b1 , \7175_b1 );
not ( \7175_b1 , w_17932 );
and ( \7281_b0 , \5986_b0 , w_17933 );
and ( w_17932 , w_17933 , \7175_b0 );
or ( \7282_b1 , \5998_b1 , \7173_b1 );
not ( \7173_b1 , w_17934 );
and ( \7282_b0 , \5998_b0 , w_17935 );
and ( w_17934 , w_17935 , \7173_b0 );
or ( \7283_b1 , \7281_b1 , w_17937 );
not ( w_17937 , w_17938 );
and ( \7283_b0 , \7281_b0 , w_17939 );
and ( w_17938 ,  , w_17939 );
buf ( w_17937 , \7282_b1 );
not ( w_17937 , w_17940 );
not (  , w_17941 );
and ( w_17940 , w_17941 , \7282_b0 );
or ( \7284_b1 , \7283_b1 , w_17942 );
xor ( \7284_b0 , \7283_b0 , w_17944 );
not ( w_17944 , w_17945 );
and ( w_17945 , w_17942 , w_17943 );
buf ( w_17942 , \7181_b1 );
not ( w_17942 , w_17946 );
not ( w_17943 , w_17947 );
and ( w_17946 , w_17947 , \7181_b0 );
or ( \7285_b1 , \7280_b1 , \7284_b1 );
xor ( \7285_b0 , \7280_b0 , w_17948 );
not ( w_17948 , w_17949 );
and ( w_17949 , \7284_b1 , \7284_b0 );
or ( \7286_b1 , \5881_b1 , \7082_b1 );
not ( \7082_b1 , w_17950 );
and ( \7286_b0 , \5881_b0 , w_17951 );
and ( w_17950 , w_17951 , \7082_b0 );
or ( \7287_b1 , \5893_b1 , \7080_b1 );
not ( \7080_b1 , w_17952 );
and ( \7287_b0 , \5893_b0 , w_17953 );
and ( w_17952 , w_17953 , \7080_b0 );
or ( \7288_b1 , \7286_b1 , w_17955 );
not ( w_17955 , w_17956 );
and ( \7288_b0 , \7286_b0 , w_17957 );
and ( w_17956 ,  , w_17957 );
buf ( w_17955 , \7287_b1 );
not ( w_17955 , w_17958 );
not (  , w_17959 );
and ( w_17958 , w_17959 , \7287_b0 );
or ( \7289_b1 , \7288_b1 , w_17960 );
xor ( \7289_b0 , \7288_b0 , w_17962 );
not ( w_17962 , w_17963 );
and ( w_17963 , w_17960 , w_17961 );
buf ( w_17960 , \7088_b1 );
not ( w_17960 , w_17964 );
not ( w_17961 , w_17965 );
and ( w_17964 , w_17965 , \7088_b0 );
or ( \7290_b1 , \5906_b1 , \7099_b1 );
not ( \7099_b1 , w_17966 );
and ( \7290_b0 , \5906_b0 , w_17967 );
and ( w_17966 , w_17967 , \7099_b0 );
or ( \7291_b1 , \5918_b1 , \7097_b1 );
not ( \7097_b1 , w_17968 );
and ( \7291_b0 , \5918_b0 , w_17969 );
and ( w_17968 , w_17969 , \7097_b0 );
or ( \7292_b1 , \7290_b1 , w_17971 );
not ( w_17971 , w_17972 );
and ( \7292_b0 , \7290_b0 , w_17973 );
and ( w_17972 ,  , w_17973 );
buf ( w_17971 , \7291_b1 );
not ( w_17971 , w_17974 );
not (  , w_17975 );
and ( w_17974 , w_17975 , \7291_b0 );
or ( \7293_b1 , \7292_b1 , w_17976 );
xor ( \7293_b0 , \7292_b0 , w_17978 );
not ( w_17978 , w_17979 );
and ( w_17979 , w_17976 , w_17977 );
buf ( w_17976 , \7105_b1 );
not ( w_17976 , w_17980 );
not ( w_17977 , w_17981 );
and ( w_17980 , w_17981 , \7105_b0 );
or ( \7294_b1 , \7289_b1 , \7293_b1 );
xor ( \7294_b0 , \7289_b0 , w_17982 );
not ( w_17982 , w_17983 );
and ( w_17983 , \7293_b1 , \7293_b0 );
or ( \7295_b1 , \5925_b1 , \7117_b1 );
not ( \7117_b1 , w_17984 );
and ( \7295_b0 , \5925_b0 , w_17985 );
and ( w_17984 , w_17985 , \7117_b0 );
or ( \7296_b1 , \5937_b1 , \7115_b1 );
not ( \7115_b1 , w_17986 );
and ( \7296_b0 , \5937_b0 , w_17987 );
and ( w_17986 , w_17987 , \7115_b0 );
or ( \7297_b1 , \7295_b1 , w_17989 );
not ( w_17989 , w_17990 );
and ( \7297_b0 , \7295_b0 , w_17991 );
and ( w_17990 ,  , w_17991 );
buf ( w_17989 , \7296_b1 );
not ( w_17989 , w_17992 );
not (  , w_17993 );
and ( w_17992 , w_17993 , \7296_b0 );
or ( \7298_b1 , \7297_b1 , w_17994 );
xor ( \7298_b0 , \7297_b0 , w_17996 );
not ( w_17996 , w_17997 );
and ( w_17997 , w_17994 , w_17995 );
buf ( w_17994 , \7123_b1 );
not ( w_17994 , w_17998 );
not ( w_17995 , w_17999 );
and ( w_17998 , w_17999 , \7123_b0 );
or ( \7299_b1 , \7294_b1 , \7298_b1 );
xor ( \7299_b0 , \7294_b0 , w_18000 );
not ( w_18000 , w_18001 );
and ( w_18001 , \7298_b1 , \7298_b0 );
or ( \7300_b1 , \7285_b1 , \7299_b1 );
xor ( \7300_b0 , \7285_b0 , w_18002 );
not ( w_18002 , w_18003 );
and ( w_18003 , \7299_b1 , \7299_b0 );
or ( \7301_b1 , \5819_b1 , \7026_b1 );
not ( \7026_b1 , w_18004 );
and ( \7301_b0 , \5819_b0 , w_18005 );
and ( w_18004 , w_18005 , \7026_b0 );
or ( \7302_b1 , \5831_b1 , \7024_b1 );
not ( \7024_b1 , w_18006 );
and ( \7302_b0 , \5831_b0 , w_18007 );
and ( w_18006 , w_18007 , \7024_b0 );
or ( \7303_b1 , \7301_b1 , w_18009 );
not ( w_18009 , w_18010 );
and ( \7303_b0 , \7301_b0 , w_18011 );
and ( w_18010 ,  , w_18011 );
buf ( w_18009 , \7302_b1 );
not ( w_18009 , w_18012 );
not (  , w_18013 );
and ( w_18012 , w_18013 , \7302_b0 );
or ( \7304_b1 , \7303_b1 , w_18014 );
xor ( \7304_b0 , \7303_b0 , w_18016 );
not ( w_18016 , w_18017 );
and ( w_18017 , w_18014 , w_18015 );
buf ( w_18014 , \7032_b1 );
not ( w_18014 , w_18018 );
not ( w_18015 , w_18019 );
and ( w_18018 , w_18019 , \7032_b0 );
or ( \7305_b1 , \5842_b1 , \7043_b1 );
not ( \7043_b1 , w_18020 );
and ( \7305_b0 , \5842_b0 , w_18021 );
and ( w_18020 , w_18021 , \7043_b0 );
or ( \7306_b1 , \5854_b1 , \7041_b1 );
not ( \7041_b1 , w_18022 );
and ( \7306_b0 , \5854_b0 , w_18023 );
and ( w_18022 , w_18023 , \7041_b0 );
or ( \7307_b1 , \7305_b1 , w_18025 );
not ( w_18025 , w_18026 );
and ( \7307_b0 , \7305_b0 , w_18027 );
and ( w_18026 ,  , w_18027 );
buf ( w_18025 , \7306_b1 );
not ( w_18025 , w_18028 );
not (  , w_18029 );
and ( w_18028 , w_18029 , \7306_b0 );
or ( \7308_b1 , \7307_b1 , w_18030 );
xor ( \7308_b0 , \7307_b0 , w_18032 );
not ( w_18032 , w_18033 );
and ( w_18033 , w_18030 , w_18031 );
buf ( w_18030 , \7049_b1 );
not ( w_18030 , w_18034 );
not ( w_18031 , w_18035 );
and ( w_18034 , w_18035 , \7049_b0 );
or ( \7309_b1 , \7304_b1 , \7308_b1 );
xor ( \7309_b0 , \7304_b0 , w_18036 );
not ( w_18036 , w_18037 );
and ( w_18037 , \7308_b1 , \7308_b0 );
or ( \7310_b1 , \5861_b1 , \7061_b1 );
not ( \7061_b1 , w_18038 );
and ( \7310_b0 , \5861_b0 , w_18039 );
and ( w_18038 , w_18039 , \7061_b0 );
or ( \7311_b1 , \5873_b1 , \7059_b1 );
not ( \7059_b1 , w_18040 );
and ( \7311_b0 , \5873_b0 , w_18041 );
and ( w_18040 , w_18041 , \7059_b0 );
or ( \7312_b1 , \7310_b1 , w_18043 );
not ( w_18043 , w_18044 );
and ( \7312_b0 , \7310_b0 , w_18045 );
and ( w_18044 ,  , w_18045 );
buf ( w_18043 , \7311_b1 );
not ( w_18043 , w_18046 );
not (  , w_18047 );
and ( w_18046 , w_18047 , \7311_b0 );
or ( \7313_b1 , \7312_b1 , w_18048 );
xor ( \7313_b0 , \7312_b0 , w_18050 );
not ( w_18050 , w_18051 );
and ( w_18051 , w_18048 , w_18049 );
buf ( w_18048 , \7067_b1 );
not ( w_18048 , w_18052 );
not ( w_18049 , w_18053 );
and ( w_18052 , w_18053 , \7067_b0 );
or ( \7314_b1 , \7309_b1 , \7313_b1 );
xor ( \7314_b0 , \7309_b0 , w_18054 );
not ( w_18054 , w_18055 );
and ( w_18055 , \7313_b1 , \7313_b0 );
or ( \7315_b1 , \7300_b1 , \7314_b1 );
xor ( \7315_b0 , \7300_b0 , w_18056 );
not ( w_18056 , w_18057 );
and ( w_18057 , \7314_b1 , \7314_b0 );
or ( \7316_b1 , \7271_b1 , \7315_b1 );
not ( \7315_b1 , w_18058 );
and ( \7316_b0 , \7271_b0 , w_18059 );
and ( w_18058 , w_18059 , \7315_b0 );
or ( \7317_b1 , \7230_b1 , \7234_b1 );
not ( \7234_b1 , w_18060 );
and ( \7317_b0 , \7230_b0 , w_18061 );
and ( w_18060 , w_18061 , \7234_b0 );
or ( \7318_b1 , \7234_b1 , \7239_b1 );
not ( \7239_b1 , w_18062 );
and ( \7318_b0 , \7234_b0 , w_18063 );
and ( w_18062 , w_18063 , \7239_b0 );
or ( \7319_b1 , \7230_b1 , \7239_b1 );
not ( \7239_b1 , w_18064 );
and ( \7319_b0 , \7230_b0 , w_18065 );
and ( w_18064 , w_18065 , \7239_b0 );
or ( \7321_b1 , \6065_b1 , w_18067 );
not ( w_18067 , w_18068 );
and ( \7321_b0 , \6065_b0 , w_18069 );
and ( w_18068 ,  , w_18069 );
buf ( w_18067 , \5766_b1 );
not ( w_18067 , w_18070 );
not (  , w_18071 );
and ( w_18070 , w_18071 , \5766_b0 );
or ( \7322_b1 , \7321_b1 , w_18072 );
xor ( \7322_b0 , \7321_b0 , w_18074 );
not ( w_18074 , w_18075 );
and ( w_18075 , w_18072 , w_18073 );
buf ( w_18072 , \5775_b1 );
not ( w_18072 , w_18076 );
not ( w_18073 , w_18077 );
and ( w_18076 , w_18077 , \5775_b0 );
or ( \7323_b1 , \7320_b1 , \7322_b1 );
xor ( \7323_b0 , \7320_b0 , w_18078 );
not ( w_18078 , w_18079 );
and ( w_18079 , \7322_b1 , \7322_b0 );
or ( \7324_b1 , \6006_b1 , \7192_b1 );
not ( \7192_b1 , w_18080 );
and ( \7324_b0 , \6006_b0 , w_18081 );
and ( w_18080 , w_18081 , \7192_b0 );
or ( \7325_b1 , \6018_b1 , \7190_b1 );
not ( \7190_b1 , w_18082 );
and ( \7325_b0 , \6018_b0 , w_18083 );
and ( w_18082 , w_18083 , \7190_b0 );
or ( \7326_b1 , \7324_b1 , w_18085 );
not ( w_18085 , w_18086 );
and ( \7326_b0 , \7324_b0 , w_18087 );
and ( w_18086 ,  , w_18087 );
buf ( w_18085 , \7325_b1 );
not ( w_18085 , w_18088 );
not (  , w_18089 );
and ( w_18088 , w_18089 , \7325_b0 );
or ( \7327_b1 , \7326_b1 , w_18090 );
xor ( \7327_b0 , \7326_b0 , w_18092 );
not ( w_18092 , w_18093 );
and ( w_18093 , w_18090 , w_18091 );
buf ( w_18090 , \7198_b1 );
not ( w_18090 , w_18094 );
not ( w_18091 , w_18095 );
and ( w_18094 , w_18095 , \7198_b0 );
or ( \7328_b1 , \6029_b1 , \7203_b1 );
not ( \7203_b1 , w_18096 );
and ( \7328_b0 , \6029_b0 , w_18097 );
and ( w_18096 , w_18097 , \7203_b0 );
or ( \7329_b1 , \6041_b1 , \7201_b1 );
not ( \7201_b1 , w_18098 );
and ( \7329_b0 , \6041_b0 , w_18099 );
and ( w_18098 , w_18099 , \7201_b0 );
or ( \7330_b1 , \7328_b1 , w_18101 );
not ( w_18101 , w_18102 );
and ( \7330_b0 , \7328_b0 , w_18103 );
and ( w_18102 ,  , w_18103 );
buf ( w_18101 , \7329_b1 );
not ( w_18101 , w_18104 );
not (  , w_18105 );
and ( w_18104 , w_18105 , \7329_b0 );
or ( \7331_b1 , \7330_b1 , w_18106 );
xor ( \7331_b0 , \7330_b0 , w_18108 );
not ( w_18108 , w_18109 );
and ( w_18109 , w_18106 , w_18107 );
buf ( w_18106 , \6824_b1 );
not ( w_18106 , w_18110 );
not ( w_18107 , w_18111 );
and ( w_18110 , w_18111 , \6824_b0 );
or ( \7332_b1 , \7327_b1 , \7331_b1 );
xor ( \7332_b0 , \7327_b0 , w_18112 );
not ( w_18112 , w_18113 );
and ( w_18113 , \7331_b1 , \7331_b0 );
or ( \7333_b1 , \6048_b1 , \5750_b1 );
not ( \5750_b1 , w_18114 );
and ( \7333_b0 , \6048_b0 , w_18115 );
and ( w_18114 , w_18115 , \5750_b0 );
or ( \7334_b1 , \6057_b1 , \5748_b1 );
not ( \5748_b1 , w_18116 );
and ( \7334_b0 , \6057_b0 , w_18117 );
and ( w_18116 , w_18117 , \5748_b0 );
or ( \7335_b1 , \7333_b1 , w_18119 );
not ( w_18119 , w_18120 );
and ( \7335_b0 , \7333_b0 , w_18121 );
and ( w_18120 ,  , w_18121 );
buf ( w_18119 , \7334_b1 );
not ( w_18119 , w_18122 );
not (  , w_18123 );
and ( w_18122 , w_18123 , \7334_b0 );
or ( \7336_b1 , \7335_b1 , w_18124 );
xor ( \7336_b0 , \7335_b0 , w_18126 );
not ( w_18126 , w_18127 );
and ( w_18127 , w_18124 , w_18125 );
buf ( w_18124 , \5755_b1 );
not ( w_18124 , w_18128 );
not ( w_18125 , w_18129 );
and ( w_18128 , w_18129 , \5755_b0 );
or ( \7337_b1 , \7332_b1 , \7336_b1 );
xor ( \7337_b0 , \7332_b0 , w_18130 );
not ( w_18130 , w_18131 );
and ( w_18131 , \7336_b1 , \7336_b0 );
or ( \7338_b1 , \7323_b1 , \7337_b1 );
xor ( \7338_b0 , \7323_b0 , w_18132 );
not ( w_18132 , w_18133 );
and ( w_18133 , \7337_b1 , \7337_b0 );
or ( \7339_b1 , \7315_b1 , \7338_b1 );
not ( \7338_b1 , w_18134 );
and ( \7339_b0 , \7315_b0 , w_18135 );
and ( w_18134 , w_18135 , \7338_b0 );
or ( \7340_b1 , \7271_b1 , \7338_b1 );
not ( \7338_b1 , w_18136 );
and ( \7340_b0 , \7271_b0 , w_18137 );
and ( w_18136 , w_18137 , \7338_b0 );
or ( \7342_b1 , \7261_b1 , \7341_b1 );
not ( \7341_b1 , w_18138 );
and ( \7342_b0 , \7261_b0 , w_18139 );
and ( w_18138 , w_18139 , \7341_b0 );
or ( \7343_b1 , \5775_b1 , \7265_b1 );
not ( \7265_b1 , w_18140 );
and ( \7343_b0 , \5775_b0 , w_18141 );
and ( w_18140 , w_18141 , \7265_b0 );
or ( \7344_b1 , \7265_b1 , \7270_b1 );
not ( \7270_b1 , w_18142 );
and ( \7344_b0 , \7265_b0 , w_18143 );
and ( w_18142 , w_18143 , \7270_b0 );
or ( \7345_b1 , \5775_b1 , \7270_b1 );
not ( \7270_b1 , w_18144 );
and ( \7345_b0 , \5775_b0 , w_18145 );
and ( w_18144 , w_18145 , \7270_b0 );
or ( \7347_b1 , \7304_b1 , \7308_b1 );
not ( \7308_b1 , w_18146 );
and ( \7347_b0 , \7304_b0 , w_18147 );
and ( w_18146 , w_18147 , \7308_b0 );
or ( \7348_b1 , \7308_b1 , \7313_b1 );
not ( \7313_b1 , w_18148 );
and ( \7348_b0 , \7308_b0 , w_18149 );
and ( w_18148 , w_18149 , \7313_b0 );
or ( \7349_b1 , \7304_b1 , \7313_b1 );
not ( \7313_b1 , w_18150 );
and ( \7349_b0 , \7304_b0 , w_18151 );
and ( w_18150 , w_18151 , \7313_b0 );
or ( \7351_b1 , \7346_b1 , \7350_b1 );
xor ( \7351_b0 , \7346_b0 , w_18152 );
not ( w_18152 , w_18153 );
and ( w_18153 , \7350_b1 , \7350_b0 );
or ( \7352_b1 , \7289_b1 , \7293_b1 );
not ( \7293_b1 , w_18154 );
and ( \7352_b0 , \7289_b0 , w_18155 );
and ( w_18154 , w_18155 , \7293_b0 );
or ( \7353_b1 , \7293_b1 , \7298_b1 );
not ( \7298_b1 , w_18156 );
and ( \7353_b0 , \7293_b0 , w_18157 );
and ( w_18156 , w_18157 , \7298_b0 );
or ( \7354_b1 , \7289_b1 , \7298_b1 );
not ( \7298_b1 , w_18158 );
and ( \7354_b0 , \7289_b0 , w_18159 );
and ( w_18158 , w_18159 , \7298_b0 );
or ( \7356_b1 , \7351_b1 , \7355_b1 );
xor ( \7356_b0 , \7351_b0 , w_18160 );
not ( w_18160 , w_18161 );
and ( w_18161 , \7355_b1 , \7355_b0 );
or ( \7357_b1 , \7341_b1 , \7356_b1 );
not ( \7356_b1 , w_18162 );
and ( \7357_b0 , \7341_b0 , w_18163 );
and ( w_18162 , w_18163 , \7356_b0 );
or ( \7358_b1 , \7261_b1 , \7356_b1 );
not ( \7356_b1 , w_18164 );
and ( \7358_b0 , \7261_b0 , w_18165 );
and ( w_18164 , w_18165 , \7356_b0 );
or ( \7360_b1 , \5792_b1 , \6991_b1 );
not ( \6991_b1 , w_18166 );
and ( \7360_b0 , \5792_b0 , w_18167 );
and ( w_18166 , w_18167 , \6991_b0 );
or ( \7361_b1 , \5758_b1 , \6988_b1 );
not ( \6988_b1 , w_18168 );
and ( \7361_b0 , \5758_b0 , w_18169 );
and ( w_18168 , w_18169 , \6988_b0 );
or ( \7362_b1 , \7360_b1 , w_18171 );
not ( w_18171 , w_18172 );
and ( \7362_b0 , \7360_b0 , w_18173 );
and ( w_18172 ,  , w_18173 );
buf ( w_18171 , \7361_b1 );
not ( w_18171 , w_18174 );
not (  , w_18175 );
and ( w_18174 , w_18175 , \7361_b0 );
or ( \7363_b1 , \7362_b1 , w_18176 );
xor ( \7363_b0 , \7362_b0 , w_18178 );
not ( w_18178 , w_18179 );
and ( w_18179 , w_18176 , w_18177 );
buf ( w_18176 , \6985_b1 );
not ( w_18176 , w_18180 );
not ( w_18177 , w_18181 );
and ( w_18180 , w_18181 , \6985_b0 );
or ( \7364_b1 , \5811_b1 , \7006_b1 );
not ( \7006_b1 , w_18182 );
and ( \7364_b0 , \5811_b0 , w_18183 );
and ( w_18182 , w_18183 , \7006_b0 );
or ( \7365_b1 , \5780_b1 , \7004_b1 );
not ( \7004_b1 , w_18184 );
and ( \7365_b0 , \5780_b0 , w_18185 );
and ( w_18184 , w_18185 , \7004_b0 );
or ( \7366_b1 , \7364_b1 , w_18187 );
not ( w_18187 , w_18188 );
and ( \7366_b0 , \7364_b0 , w_18189 );
and ( w_18188 ,  , w_18189 );
buf ( w_18187 , \7365_b1 );
not ( w_18187 , w_18190 );
not (  , w_18191 );
and ( w_18190 , w_18191 , \7365_b0 );
or ( \7367_b1 , \7366_b1 , w_18192 );
xor ( \7367_b0 , \7366_b0 , w_18194 );
not ( w_18194 , w_18195 );
and ( w_18195 , w_18192 , w_18193 );
buf ( w_18192 , \7012_b1 );
not ( w_18192 , w_18196 );
not ( w_18193 , w_18197 );
and ( w_18196 , w_18197 , \7012_b0 );
or ( \7368_b1 , \7363_b1 , \7367_b1 );
xor ( \7368_b0 , \7363_b0 , w_18198 );
not ( w_18198 , w_18199 );
and ( w_18199 , \7367_b1 , \7367_b0 );
or ( \7369_b1 , \5831_b1 , \7026_b1 );
not ( \7026_b1 , w_18200 );
and ( \7369_b0 , \5831_b0 , w_18201 );
and ( w_18200 , w_18201 , \7026_b0 );
or ( \7370_b1 , \5799_b1 , \7024_b1 );
not ( \7024_b1 , w_18202 );
and ( \7370_b0 , \5799_b0 , w_18203 );
and ( w_18202 , w_18203 , \7024_b0 );
or ( \7371_b1 , \7369_b1 , w_18205 );
not ( w_18205 , w_18206 );
and ( \7371_b0 , \7369_b0 , w_18207 );
and ( w_18206 ,  , w_18207 );
buf ( w_18205 , \7370_b1 );
not ( w_18205 , w_18208 );
not (  , w_18209 );
and ( w_18208 , w_18209 , \7370_b0 );
or ( \7372_b1 , \7371_b1 , w_18210 );
xor ( \7372_b0 , \7371_b0 , w_18212 );
not ( w_18212 , w_18213 );
and ( w_18213 , w_18210 , w_18211 );
buf ( w_18210 , \7032_b1 );
not ( w_18210 , w_18214 );
not ( w_18211 , w_18215 );
and ( w_18214 , w_18215 , \7032_b0 );
or ( \7373_b1 , \7368_b1 , \7372_b1 );
xor ( \7373_b0 , \7368_b0 , w_18216 );
not ( w_18216 , w_18217 );
and ( w_18217 , \7372_b1 , \7372_b0 );
or ( \7374_b1 , \5979_b1 , \7157_b1 );
not ( \7157_b1 , w_18218 );
and ( \7374_b0 , \5979_b0 , w_18219 );
and ( w_18218 , w_18219 , \7157_b0 );
or ( \7375_b1 , \5945_b1 , \7155_b1 );
not ( \7155_b1 , w_18220 );
and ( \7375_b0 , \5945_b0 , w_18221 );
and ( w_18220 , w_18221 , \7155_b0 );
or ( \7376_b1 , \7374_b1 , w_18223 );
not ( w_18223 , w_18224 );
and ( \7376_b0 , \7374_b0 , w_18225 );
and ( w_18224 ,  , w_18225 );
buf ( w_18223 , \7375_b1 );
not ( w_18223 , w_18226 );
not (  , w_18227 );
and ( w_18226 , w_18227 , \7375_b0 );
or ( \7377_b1 , \7376_b1 , w_18228 );
xor ( \7377_b0 , \7376_b0 , w_18230 );
not ( w_18230 , w_18231 );
and ( w_18231 , w_18228 , w_18229 );
buf ( w_18228 , \7163_b1 );
not ( w_18228 , w_18232 );
not ( w_18229 , w_18233 );
and ( w_18232 , w_18233 , \7163_b0 );
or ( \7378_b1 , \5998_b1 , \7175_b1 );
not ( \7175_b1 , w_18234 );
and ( \7378_b0 , \5998_b0 , w_18235 );
and ( w_18234 , w_18235 , \7175_b0 );
or ( \7379_b1 , \5967_b1 , \7173_b1 );
not ( \7173_b1 , w_18236 );
and ( \7379_b0 , \5967_b0 , w_18237 );
and ( w_18236 , w_18237 , \7173_b0 );
or ( \7380_b1 , \7378_b1 , w_18239 );
not ( w_18239 , w_18240 );
and ( \7380_b0 , \7378_b0 , w_18241 );
and ( w_18240 ,  , w_18241 );
buf ( w_18239 , \7379_b1 );
not ( w_18239 , w_18242 );
not (  , w_18243 );
and ( w_18242 , w_18243 , \7379_b0 );
or ( \7381_b1 , \7380_b1 , w_18244 );
xor ( \7381_b0 , \7380_b0 , w_18246 );
not ( w_18246 , w_18247 );
and ( w_18247 , w_18244 , w_18245 );
buf ( w_18244 , \7181_b1 );
not ( w_18244 , w_18248 );
not ( w_18245 , w_18249 );
and ( w_18248 , w_18249 , \7181_b0 );
or ( \7382_b1 , \7377_b1 , \7381_b1 );
xor ( \7382_b0 , \7377_b0 , w_18250 );
not ( w_18250 , w_18251 );
and ( w_18251 , \7381_b1 , \7381_b0 );
or ( \7383_b1 , \6018_b1 , \7192_b1 );
not ( \7192_b1 , w_18252 );
and ( \7383_b0 , \6018_b0 , w_18253 );
and ( w_18252 , w_18253 , \7192_b0 );
or ( \7384_b1 , \5986_b1 , \7190_b1 );
not ( \7190_b1 , w_18254 );
and ( \7384_b0 , \5986_b0 , w_18255 );
and ( w_18254 , w_18255 , \7190_b0 );
or ( \7385_b1 , \7383_b1 , w_18257 );
not ( w_18257 , w_18258 );
and ( \7385_b0 , \7383_b0 , w_18259 );
and ( w_18258 ,  , w_18259 );
buf ( w_18257 , \7384_b1 );
not ( w_18257 , w_18260 );
not (  , w_18261 );
and ( w_18260 , w_18261 , \7384_b0 );
or ( \7386_b1 , \7385_b1 , w_18262 );
xor ( \7386_b0 , \7385_b0 , w_18264 );
not ( w_18264 , w_18265 );
and ( w_18265 , w_18262 , w_18263 );
buf ( w_18262 , \7198_b1 );
not ( w_18262 , w_18266 );
not ( w_18263 , w_18267 );
and ( w_18266 , w_18267 , \7198_b0 );
or ( \7387_b1 , \7382_b1 , \7386_b1 );
xor ( \7387_b0 , \7382_b0 , w_18268 );
not ( w_18268 , w_18269 );
and ( w_18269 , \7386_b1 , \7386_b0 );
or ( \7388_b1 , \5918_b1 , \7099_b1 );
not ( \7099_b1 , w_18270 );
and ( \7388_b0 , \5918_b0 , w_18271 );
and ( w_18270 , w_18271 , \7099_b0 );
or ( \7389_b1 , \5881_b1 , \7097_b1 );
not ( \7097_b1 , w_18272 );
and ( \7389_b0 , \5881_b0 , w_18273 );
and ( w_18272 , w_18273 , \7097_b0 );
or ( \7390_b1 , \7388_b1 , w_18275 );
not ( w_18275 , w_18276 );
and ( \7390_b0 , \7388_b0 , w_18277 );
and ( w_18276 ,  , w_18277 );
buf ( w_18275 , \7389_b1 );
not ( w_18275 , w_18278 );
not (  , w_18279 );
and ( w_18278 , w_18279 , \7389_b0 );
or ( \7391_b1 , \7390_b1 , w_18280 );
xor ( \7391_b0 , \7390_b0 , w_18282 );
not ( w_18282 , w_18283 );
and ( w_18283 , w_18280 , w_18281 );
buf ( w_18280 , \7105_b1 );
not ( w_18280 , w_18284 );
not ( w_18281 , w_18285 );
and ( w_18284 , w_18285 , \7105_b0 );
or ( \7392_b1 , \5937_b1 , \7117_b1 );
not ( \7117_b1 , w_18286 );
and ( \7392_b0 , \5937_b0 , w_18287 );
and ( w_18286 , w_18287 , \7117_b0 );
or ( \7393_b1 , \5906_b1 , \7115_b1 );
not ( \7115_b1 , w_18288 );
and ( \7393_b0 , \5906_b0 , w_18289 );
and ( w_18288 , w_18289 , \7115_b0 );
or ( \7394_b1 , \7392_b1 , w_18291 );
not ( w_18291 , w_18292 );
and ( \7394_b0 , \7392_b0 , w_18293 );
and ( w_18292 ,  , w_18293 );
buf ( w_18291 , \7393_b1 );
not ( w_18291 , w_18294 );
not (  , w_18295 );
and ( w_18294 , w_18295 , \7393_b0 );
or ( \7395_b1 , \7394_b1 , w_18296 );
xor ( \7395_b0 , \7394_b0 , w_18298 );
not ( w_18298 , w_18299 );
and ( w_18299 , w_18296 , w_18297 );
buf ( w_18296 , \7123_b1 );
not ( w_18296 , w_18300 );
not ( w_18297 , w_18301 );
and ( w_18300 , w_18301 , \7123_b0 );
or ( \7396_b1 , \7391_b1 , \7395_b1 );
xor ( \7396_b0 , \7391_b0 , w_18302 );
not ( w_18302 , w_18303 );
and ( w_18303 , \7395_b1 , \7395_b0 );
or ( \7397_b1 , \5957_b1 , \7140_b1 );
not ( \7140_b1 , w_18304 );
and ( \7397_b0 , \5957_b0 , w_18305 );
and ( w_18304 , w_18305 , \7140_b0 );
or ( \7398_b1 , \5925_b1 , \7138_b1 );
not ( \7138_b1 , w_18306 );
and ( \7398_b0 , \5925_b0 , w_18307 );
and ( w_18306 , w_18307 , \7138_b0 );
or ( \7399_b1 , \7397_b1 , w_18309 );
not ( w_18309 , w_18310 );
and ( \7399_b0 , \7397_b0 , w_18311 );
and ( w_18310 ,  , w_18311 );
buf ( w_18309 , \7398_b1 );
not ( w_18309 , w_18312 );
not (  , w_18313 );
and ( w_18312 , w_18313 , \7398_b0 );
or ( \7400_b1 , \7399_b1 , w_18314 );
xor ( \7400_b0 , \7399_b0 , w_18316 );
not ( w_18316 , w_18317 );
and ( w_18317 , w_18314 , w_18315 );
buf ( w_18314 , \7146_b1 );
not ( w_18314 , w_18318 );
not ( w_18315 , w_18319 );
and ( w_18318 , w_18319 , \7146_b0 );
or ( \7401_b1 , \7396_b1 , \7400_b1 );
xor ( \7401_b0 , \7396_b0 , w_18320 );
not ( w_18320 , w_18321 );
and ( w_18321 , \7400_b1 , \7400_b0 );
or ( \7402_b1 , \7387_b1 , \7401_b1 );
xor ( \7402_b0 , \7387_b0 , w_18322 );
not ( w_18322 , w_18323 );
and ( w_18323 , \7401_b1 , \7401_b0 );
or ( \7403_b1 , \5854_b1 , \7043_b1 );
not ( \7043_b1 , w_18324 );
and ( \7403_b0 , \5854_b0 , w_18325 );
and ( w_18324 , w_18325 , \7043_b0 );
or ( \7404_b1 , \5819_b1 , \7041_b1 );
not ( \7041_b1 , w_18326 );
and ( \7404_b0 , \5819_b0 , w_18327 );
and ( w_18326 , w_18327 , \7041_b0 );
or ( \7405_b1 , \7403_b1 , w_18329 );
not ( w_18329 , w_18330 );
and ( \7405_b0 , \7403_b0 , w_18331 );
and ( w_18330 ,  , w_18331 );
buf ( w_18329 , \7404_b1 );
not ( w_18329 , w_18332 );
not (  , w_18333 );
and ( w_18332 , w_18333 , \7404_b0 );
or ( \7406_b1 , \7405_b1 , w_18334 );
xor ( \7406_b0 , \7405_b0 , w_18336 );
not ( w_18336 , w_18337 );
and ( w_18337 , w_18334 , w_18335 );
buf ( w_18334 , \7049_b1 );
not ( w_18334 , w_18338 );
not ( w_18335 , w_18339 );
and ( w_18338 , w_18339 , \7049_b0 );
or ( \7407_b1 , \5873_b1 , \7061_b1 );
not ( \7061_b1 , w_18340 );
and ( \7407_b0 , \5873_b0 , w_18341 );
and ( w_18340 , w_18341 , \7061_b0 );
or ( \7408_b1 , \5842_b1 , \7059_b1 );
not ( \7059_b1 , w_18342 );
and ( \7408_b0 , \5842_b0 , w_18343 );
and ( w_18342 , w_18343 , \7059_b0 );
or ( \7409_b1 , \7407_b1 , w_18345 );
not ( w_18345 , w_18346 );
and ( \7409_b0 , \7407_b0 , w_18347 );
and ( w_18346 ,  , w_18347 );
buf ( w_18345 , \7408_b1 );
not ( w_18345 , w_18348 );
not (  , w_18349 );
and ( w_18348 , w_18349 , \7408_b0 );
or ( \7410_b1 , \7409_b1 , w_18350 );
xor ( \7410_b0 , \7409_b0 , w_18352 );
not ( w_18352 , w_18353 );
and ( w_18353 , w_18350 , w_18351 );
buf ( w_18350 , \7067_b1 );
not ( w_18350 , w_18354 );
not ( w_18351 , w_18355 );
and ( w_18354 , w_18355 , \7067_b0 );
or ( \7411_b1 , \7406_b1 , \7410_b1 );
xor ( \7411_b0 , \7406_b0 , w_18356 );
not ( w_18356 , w_18357 );
and ( w_18357 , \7410_b1 , \7410_b0 );
or ( \7412_b1 , \5893_b1 , \7082_b1 );
not ( \7082_b1 , w_18358 );
and ( \7412_b0 , \5893_b0 , w_18359 );
and ( w_18358 , w_18359 , \7082_b0 );
or ( \7413_b1 , \5861_b1 , \7080_b1 );
not ( \7080_b1 , w_18360 );
and ( \7413_b0 , \5861_b0 , w_18361 );
and ( w_18360 , w_18361 , \7080_b0 );
or ( \7414_b1 , \7412_b1 , w_18363 );
not ( w_18363 , w_18364 );
and ( \7414_b0 , \7412_b0 , w_18365 );
and ( w_18364 ,  , w_18365 );
buf ( w_18363 , \7413_b1 );
not ( w_18363 , w_18366 );
not (  , w_18367 );
and ( w_18366 , w_18367 , \7413_b0 );
or ( \7415_b1 , \7414_b1 , w_18368 );
xor ( \7415_b0 , \7414_b0 , w_18370 );
not ( w_18370 , w_18371 );
and ( w_18371 , w_18368 , w_18369 );
buf ( w_18368 , \7088_b1 );
not ( w_18368 , w_18372 );
not ( w_18369 , w_18373 );
and ( w_18372 , w_18373 , \7088_b0 );
or ( \7416_b1 , \7411_b1 , \7415_b1 );
xor ( \7416_b0 , \7411_b0 , w_18374 );
not ( w_18374 , w_18375 );
and ( w_18375 , \7415_b1 , \7415_b0 );
or ( \7417_b1 , \7402_b1 , \7416_b1 );
xor ( \7417_b0 , \7402_b0 , w_18376 );
not ( w_18376 , w_18377 );
and ( w_18377 , \7416_b1 , \7416_b0 );
or ( \7418_b1 , \7373_b1 , \7417_b1 );
xor ( \7418_b0 , \7373_b0 , w_18378 );
not ( w_18378 , w_18379 );
and ( w_18379 , \7417_b1 , \7417_b0 );
or ( \7419_b1 , \7275_b1 , \7279_b1 );
not ( \7279_b1 , w_18380 );
and ( \7419_b0 , \7275_b0 , w_18381 );
and ( w_18380 , w_18381 , \7279_b0 );
or ( \7420_b1 , \7279_b1 , \7284_b1 );
not ( \7284_b1 , w_18382 );
and ( \7420_b0 , \7279_b0 , w_18383 );
and ( w_18382 , w_18383 , \7284_b0 );
or ( \7421_b1 , \7275_b1 , \7284_b1 );
not ( \7284_b1 , w_18384 );
and ( \7421_b0 , \7275_b0 , w_18385 );
and ( w_18384 , w_18385 , \7284_b0 );
or ( \7423_b1 , \7327_b1 , \7331_b1 );
not ( \7331_b1 , w_18386 );
and ( \7423_b0 , \7327_b0 , w_18387 );
and ( w_18386 , w_18387 , \7331_b0 );
or ( \7424_b1 , \7331_b1 , \7336_b1 );
not ( \7336_b1 , w_18388 );
and ( \7424_b0 , \7331_b0 , w_18389 );
and ( w_18388 , w_18389 , \7336_b0 );
or ( \7425_b1 , \7327_b1 , \7336_b1 );
not ( \7336_b1 , w_18390 );
and ( \7425_b0 , \7327_b0 , w_18391 );
and ( w_18390 , w_18391 , \7336_b0 );
or ( \7427_b1 , \7422_b1 , \7426_b1 );
xor ( \7427_b0 , \7422_b0 , w_18392 );
not ( w_18392 , w_18393 );
and ( w_18393 , \7426_b1 , \7426_b0 );
or ( \7428_b1 , \6041_b1 , \7203_b1 );
not ( \7203_b1 , w_18394 );
and ( \7428_b0 , \6041_b0 , w_18395 );
and ( w_18394 , w_18395 , \7203_b0 );
or ( \7429_b1 , \6006_b1 , \7201_b1 );
not ( \7201_b1 , w_18396 );
and ( \7429_b0 , \6006_b0 , w_18397 );
and ( w_18396 , w_18397 , \7201_b0 );
or ( \7430_b1 , \7428_b1 , w_18399 );
not ( w_18399 , w_18400 );
and ( \7430_b0 , \7428_b0 , w_18401 );
and ( w_18400 ,  , w_18401 );
buf ( w_18399 , \7429_b1 );
not ( w_18399 , w_18402 );
not (  , w_18403 );
and ( w_18402 , w_18403 , \7429_b0 );
or ( \7431_b1 , \7430_b1 , w_18404 );
xor ( \7431_b0 , \7430_b0 , w_18406 );
not ( w_18406 , w_18407 );
and ( w_18407 , w_18404 , w_18405 );
buf ( w_18404 , \6824_b1 );
not ( w_18404 , w_18408 );
not ( w_18405 , w_18409 );
and ( w_18408 , w_18409 , \6824_b0 );
or ( \7432_b1 , \6057_b1 , \5750_b1 );
not ( \5750_b1 , w_18410 );
and ( \7432_b0 , \6057_b0 , w_18411 );
and ( w_18410 , w_18411 , \5750_b0 );
or ( \7433_b1 , \6029_b1 , \5748_b1 );
not ( \5748_b1 , w_18412 );
and ( \7433_b0 , \6029_b0 , w_18413 );
and ( w_18412 , w_18413 , \5748_b0 );
or ( \7434_b1 , \7432_b1 , w_18415 );
not ( w_18415 , w_18416 );
and ( \7434_b0 , \7432_b0 , w_18417 );
and ( w_18416 ,  , w_18417 );
buf ( w_18415 , \7433_b1 );
not ( w_18415 , w_18418 );
not (  , w_18419 );
and ( w_18418 , w_18419 , \7433_b0 );
or ( \7435_b1 , \7434_b1 , w_18420 );
xor ( \7435_b0 , \7434_b0 , w_18422 );
not ( w_18422 , w_18423 );
and ( w_18423 , w_18420 , w_18421 );
buf ( w_18420 , \5755_b1 );
not ( w_18420 , w_18424 );
not ( w_18421 , w_18425 );
and ( w_18424 , w_18425 , \5755_b0 );
or ( \7436_b1 , \7431_b1 , \7435_b1 );
xor ( \7436_b0 , \7431_b0 , w_18426 );
not ( w_18426 , w_18427 );
and ( w_18427 , \7435_b1 , \7435_b0 );
or ( \7437_b1 , \6065_b1 , \5768_b1 );
not ( \5768_b1 , w_18428 );
and ( \7437_b0 , \6065_b0 , w_18429 );
and ( w_18428 , w_18429 , \5768_b0 );
or ( \7438_b1 , \6048_b1 , \5766_b1 );
not ( \5766_b1 , w_18430 );
and ( \7438_b0 , \6048_b0 , w_18431 );
and ( w_18430 , w_18431 , \5766_b0 );
or ( \7439_b1 , \7437_b1 , w_18433 );
not ( w_18433 , w_18434 );
and ( \7439_b0 , \7437_b0 , w_18435 );
and ( w_18434 ,  , w_18435 );
buf ( w_18433 , \7438_b1 );
not ( w_18433 , w_18436 );
not (  , w_18437 );
and ( w_18436 , w_18437 , \7438_b0 );
or ( \7440_b1 , \7439_b1 , w_18438 );
xor ( \7440_b0 , \7439_b0 , w_18440 );
not ( w_18440 , w_18441 );
and ( w_18441 , w_18438 , w_18439 );
buf ( w_18438 , \5775_b1 );
not ( w_18438 , w_18442 );
not ( w_18439 , w_18443 );
and ( w_18442 , w_18443 , \5775_b0 );
or ( \7441_b1 , \7436_b1 , \7440_b1 );
xor ( \7441_b0 , \7436_b0 , w_18444 );
not ( w_18444 , w_18445 );
and ( w_18445 , \7440_b1 , \7440_b0 );
or ( \7442_b1 , \7427_b1 , \7441_b1 );
xor ( \7442_b0 , \7427_b0 , w_18446 );
not ( w_18446 , w_18447 );
and ( w_18447 , \7441_b1 , \7441_b0 );
or ( \7443_b1 , \7418_b1 , \7442_b1 );
xor ( \7443_b0 , \7418_b0 , w_18448 );
not ( w_18448 , w_18449 );
and ( w_18449 , \7442_b1 , \7442_b0 );
or ( \7444_b1 , \5811_b1 , \6991_b1 );
not ( \6991_b1 , w_18450 );
and ( \7444_b0 , \5811_b0 , w_18451 );
and ( w_18450 , w_18451 , \6991_b0 );
or ( \7445_b1 , \5780_b1 , \6988_b1 );
not ( \6988_b1 , w_18452 );
and ( \7445_b0 , \5780_b0 , w_18453 );
and ( w_18452 , w_18453 , \6988_b0 );
or ( \7446_b1 , \7444_b1 , w_18455 );
not ( w_18455 , w_18456 );
and ( \7446_b0 , \7444_b0 , w_18457 );
and ( w_18456 ,  , w_18457 );
buf ( w_18455 , \7445_b1 );
not ( w_18455 , w_18458 );
not (  , w_18459 );
and ( w_18458 , w_18459 , \7445_b0 );
or ( \7447_b1 , \7446_b1 , w_18460 );
xor ( \7447_b0 , \7446_b0 , w_18462 );
not ( w_18462 , w_18463 );
and ( w_18463 , w_18460 , w_18461 );
buf ( w_18460 , \6985_b1 );
not ( w_18460 , w_18464 );
not ( w_18461 , w_18465 );
and ( w_18464 , w_18465 , \6985_b0 );
or ( \7448_b1 , \5831_b1 , \7006_b1 );
not ( \7006_b1 , w_18466 );
and ( \7448_b0 , \5831_b0 , w_18467 );
and ( w_18466 , w_18467 , \7006_b0 );
or ( \7449_b1 , \5799_b1 , \7004_b1 );
not ( \7004_b1 , w_18468 );
and ( \7449_b0 , \5799_b0 , w_18469 );
and ( w_18468 , w_18469 , \7004_b0 );
or ( \7450_b1 , \7448_b1 , w_18471 );
not ( w_18471 , w_18472 );
and ( \7450_b0 , \7448_b0 , w_18473 );
and ( w_18472 ,  , w_18473 );
buf ( w_18471 , \7449_b1 );
not ( w_18471 , w_18474 );
not (  , w_18475 );
and ( w_18474 , w_18475 , \7449_b0 );
or ( \7451_b1 , \7450_b1 , w_18476 );
xor ( \7451_b0 , \7450_b0 , w_18478 );
not ( w_18478 , w_18479 );
and ( w_18479 , w_18476 , w_18477 );
buf ( w_18476 , \7012_b1 );
not ( w_18476 , w_18480 );
not ( w_18477 , w_18481 );
and ( w_18480 , w_18481 , \7012_b0 );
or ( \7452_b1 , \7447_b1 , \7451_b1 );
not ( \7451_b1 , w_18482 );
and ( \7452_b0 , \7447_b0 , w_18483 );
and ( w_18482 , w_18483 , \7451_b0 );
or ( \7453_b1 , \5854_b1 , \7026_b1 );
not ( \7026_b1 , w_18484 );
and ( \7453_b0 , \5854_b0 , w_18485 );
and ( w_18484 , w_18485 , \7026_b0 );
or ( \7454_b1 , \5819_b1 , \7024_b1 );
not ( \7024_b1 , w_18486 );
and ( \7454_b0 , \5819_b0 , w_18487 );
and ( w_18486 , w_18487 , \7024_b0 );
or ( \7455_b1 , \7453_b1 , w_18489 );
not ( w_18489 , w_18490 );
and ( \7455_b0 , \7453_b0 , w_18491 );
and ( w_18490 ,  , w_18491 );
buf ( w_18489 , \7454_b1 );
not ( w_18489 , w_18492 );
not (  , w_18493 );
and ( w_18492 , w_18493 , \7454_b0 );
or ( \7456_b1 , \7455_b1 , w_18494 );
xor ( \7456_b0 , \7455_b0 , w_18496 );
not ( w_18496 , w_18497 );
and ( w_18497 , w_18494 , w_18495 );
buf ( w_18494 , \7032_b1 );
not ( w_18494 , w_18498 );
not ( w_18495 , w_18499 );
and ( w_18498 , w_18499 , \7032_b0 );
or ( \7457_b1 , \7451_b1 , \7456_b1 );
not ( \7456_b1 , w_18500 );
and ( \7457_b0 , \7451_b0 , w_18501 );
and ( w_18500 , w_18501 , \7456_b0 );
or ( \7458_b1 , \7447_b1 , \7456_b1 );
not ( \7456_b1 , w_18502 );
and ( \7458_b0 , \7447_b0 , w_18503 );
and ( w_18502 , w_18503 , \7456_b0 );
or ( \7460_b1 , \5873_b1 , \7043_b1 );
not ( \7043_b1 , w_18504 );
and ( \7460_b0 , \5873_b0 , w_18505 );
and ( w_18504 , w_18505 , \7043_b0 );
or ( \7461_b1 , \5842_b1 , \7041_b1 );
not ( \7041_b1 , w_18506 );
and ( \7461_b0 , \5842_b0 , w_18507 );
and ( w_18506 , w_18507 , \7041_b0 );
or ( \7462_b1 , \7460_b1 , w_18509 );
not ( w_18509 , w_18510 );
and ( \7462_b0 , \7460_b0 , w_18511 );
and ( w_18510 ,  , w_18511 );
buf ( w_18509 , \7461_b1 );
not ( w_18509 , w_18512 );
not (  , w_18513 );
and ( w_18512 , w_18513 , \7461_b0 );
or ( \7463_b1 , \7462_b1 , w_18514 );
xor ( \7463_b0 , \7462_b0 , w_18516 );
not ( w_18516 , w_18517 );
and ( w_18517 , w_18514 , w_18515 );
buf ( w_18514 , \7049_b1 );
not ( w_18514 , w_18518 );
not ( w_18515 , w_18519 );
and ( w_18518 , w_18519 , \7049_b0 );
or ( \7464_b1 , \5893_b1 , \7061_b1 );
not ( \7061_b1 , w_18520 );
and ( \7464_b0 , \5893_b0 , w_18521 );
and ( w_18520 , w_18521 , \7061_b0 );
or ( \7465_b1 , \5861_b1 , \7059_b1 );
not ( \7059_b1 , w_18522 );
and ( \7465_b0 , \5861_b0 , w_18523 );
and ( w_18522 , w_18523 , \7059_b0 );
or ( \7466_b1 , \7464_b1 , w_18525 );
not ( w_18525 , w_18526 );
and ( \7466_b0 , \7464_b0 , w_18527 );
and ( w_18526 ,  , w_18527 );
buf ( w_18525 , \7465_b1 );
not ( w_18525 , w_18528 );
not (  , w_18529 );
and ( w_18528 , w_18529 , \7465_b0 );
or ( \7467_b1 , \7466_b1 , w_18530 );
xor ( \7467_b0 , \7466_b0 , w_18532 );
not ( w_18532 , w_18533 );
and ( w_18533 , w_18530 , w_18531 );
buf ( w_18530 , \7067_b1 );
not ( w_18530 , w_18534 );
not ( w_18531 , w_18535 );
and ( w_18534 , w_18535 , \7067_b0 );
or ( \7468_b1 , \7463_b1 , \7467_b1 );
not ( \7467_b1 , w_18536 );
and ( \7468_b0 , \7463_b0 , w_18537 );
and ( w_18536 , w_18537 , \7467_b0 );
or ( \7469_b1 , \5918_b1 , \7082_b1 );
not ( \7082_b1 , w_18538 );
and ( \7469_b0 , \5918_b0 , w_18539 );
and ( w_18538 , w_18539 , \7082_b0 );
or ( \7470_b1 , \5881_b1 , \7080_b1 );
not ( \7080_b1 , w_18540 );
and ( \7470_b0 , \5881_b0 , w_18541 );
and ( w_18540 , w_18541 , \7080_b0 );
or ( \7471_b1 , \7469_b1 , w_18543 );
not ( w_18543 , w_18544 );
and ( \7471_b0 , \7469_b0 , w_18545 );
and ( w_18544 ,  , w_18545 );
buf ( w_18543 , \7470_b1 );
not ( w_18543 , w_18546 );
not (  , w_18547 );
and ( w_18546 , w_18547 , \7470_b0 );
or ( \7472_b1 , \7471_b1 , w_18548 );
xor ( \7472_b0 , \7471_b0 , w_18550 );
not ( w_18550 , w_18551 );
and ( w_18551 , w_18548 , w_18549 );
buf ( w_18548 , \7088_b1 );
not ( w_18548 , w_18552 );
not ( w_18549 , w_18553 );
and ( w_18552 , w_18553 , \7088_b0 );
or ( \7473_b1 , \7467_b1 , \7472_b1 );
not ( \7472_b1 , w_18554 );
and ( \7473_b0 , \7467_b0 , w_18555 );
and ( w_18554 , w_18555 , \7472_b0 );
or ( \7474_b1 , \7463_b1 , \7472_b1 );
not ( \7472_b1 , w_18556 );
and ( \7474_b0 , \7463_b0 , w_18557 );
and ( w_18556 , w_18557 , \7472_b0 );
or ( \7476_b1 , \7459_b1 , \7475_b1 );
not ( \7475_b1 , w_18558 );
and ( \7476_b0 , \7459_b0 , w_18559 );
and ( w_18558 , w_18559 , \7475_b0 );
or ( \7477_b1 , \7245_b1 , \7249_b1 );
not ( \7249_b1 , w_18560 );
and ( \7477_b0 , \7245_b0 , w_18561 );
and ( w_18560 , w_18561 , \7249_b0 );
or ( \7478_b1 , \7249_b1 , \7254_b1 );
not ( \7254_b1 , w_18562 );
and ( \7478_b0 , \7249_b0 , w_18563 );
and ( w_18562 , w_18563 , \7254_b0 );
or ( \7479_b1 , \7245_b1 , \7254_b1 );
not ( \7254_b1 , w_18564 );
and ( \7479_b0 , \7245_b0 , w_18565 );
and ( w_18564 , w_18565 , \7254_b0 );
or ( \7481_b1 , \7475_b1 , \7480_b1 );
not ( \7480_b1 , w_18566 );
and ( \7481_b0 , \7475_b0 , w_18567 );
and ( w_18566 , w_18567 , \7480_b0 );
or ( \7482_b1 , \7459_b1 , \7480_b1 );
not ( \7480_b1 , w_18568 );
and ( \7482_b0 , \7459_b0 , w_18569 );
and ( w_18568 , w_18569 , \7480_b0 );
or ( \7484_b1 , \7320_b1 , \7322_b1 );
not ( \7322_b1 , w_18570 );
and ( \7484_b0 , \7320_b0 , w_18571 );
and ( w_18570 , w_18571 , \7322_b0 );
or ( \7485_b1 , \7322_b1 , \7337_b1 );
not ( \7337_b1 , w_18572 );
and ( \7485_b0 , \7322_b0 , w_18573 );
and ( w_18572 , w_18573 , \7337_b0 );
or ( \7486_b1 , \7320_b1 , \7337_b1 );
not ( \7337_b1 , w_18574 );
and ( \7486_b0 , \7320_b0 , w_18575 );
and ( w_18574 , w_18575 , \7337_b0 );
or ( \7488_b1 , \7483_b1 , \7487_b1 );
xor ( \7488_b0 , \7483_b0 , w_18576 );
not ( w_18576 , w_18577 );
and ( w_18577 , \7487_b1 , \7487_b0 );
or ( \7489_b1 , \7285_b1 , \7299_b1 );
not ( \7299_b1 , w_18578 );
and ( \7489_b0 , \7285_b0 , w_18579 );
and ( w_18578 , w_18579 , \7299_b0 );
or ( \7490_b1 , \7299_b1 , \7314_b1 );
not ( \7314_b1 , w_18580 );
and ( \7490_b0 , \7299_b0 , w_18581 );
and ( w_18580 , w_18581 , \7314_b0 );
or ( \7491_b1 , \7285_b1 , \7314_b1 );
not ( \7314_b1 , w_18582 );
and ( \7491_b0 , \7285_b0 , w_18583 );
and ( w_18582 , w_18583 , \7314_b0 );
or ( \7493_b1 , \7488_b1 , \7492_b1 );
xor ( \7493_b0 , \7488_b0 , w_18584 );
not ( w_18584 , w_18585 );
and ( w_18585 , \7492_b1 , \7492_b0 );
or ( \7494_b1 , \7443_b1 , \7493_b1 );
not ( \7493_b1 , w_18586 );
and ( \7494_b0 , \7443_b0 , w_18587 );
and ( w_18586 , w_18587 , \7493_b0 );
or ( \7495_b1 , \7359_b1 , \7494_b1 );
not ( \7494_b1 , w_18588 );
and ( \7495_b0 , \7359_b0 , w_18589 );
and ( w_18588 , w_18589 , \7494_b0 );
or ( \7496_b1 , \5861_b1 , \7082_b1 );
not ( \7082_b1 , w_18590 );
and ( \7496_b0 , \5861_b0 , w_18591 );
and ( w_18590 , w_18591 , \7082_b0 );
or ( \7497_b1 , \5873_b1 , \7080_b1 );
not ( \7080_b1 , w_18592 );
and ( \7497_b0 , \5873_b0 , w_18593 );
and ( w_18592 , w_18593 , \7080_b0 );
or ( \7498_b1 , \7496_b1 , w_18595 );
not ( w_18595 , w_18596 );
and ( \7498_b0 , \7496_b0 , w_18597 );
and ( w_18596 ,  , w_18597 );
buf ( w_18595 , \7497_b1 );
not ( w_18595 , w_18598 );
not (  , w_18599 );
and ( w_18598 , w_18599 , \7497_b0 );
or ( \7499_b1 , \7498_b1 , w_18600 );
xor ( \7499_b0 , \7498_b0 , w_18602 );
not ( w_18602 , w_18603 );
and ( w_18603 , w_18600 , w_18601 );
buf ( w_18600 , \7088_b1 );
not ( w_18600 , w_18604 );
not ( w_18601 , w_18605 );
and ( w_18604 , w_18605 , \7088_b0 );
or ( \7500_b1 , \5881_b1 , \7099_b1 );
not ( \7099_b1 , w_18606 );
and ( \7500_b0 , \5881_b0 , w_18607 );
and ( w_18606 , w_18607 , \7099_b0 );
or ( \7501_b1 , \5893_b1 , \7097_b1 );
not ( \7097_b1 , w_18608 );
and ( \7501_b0 , \5893_b0 , w_18609 );
and ( w_18608 , w_18609 , \7097_b0 );
or ( \7502_b1 , \7500_b1 , w_18611 );
not ( w_18611 , w_18612 );
and ( \7502_b0 , \7500_b0 , w_18613 );
and ( w_18612 ,  , w_18613 );
buf ( w_18611 , \7501_b1 );
not ( w_18611 , w_18614 );
not (  , w_18615 );
and ( w_18614 , w_18615 , \7501_b0 );
or ( \7503_b1 , \7502_b1 , w_18616 );
xor ( \7503_b0 , \7502_b0 , w_18618 );
not ( w_18618 , w_18619 );
and ( w_18619 , w_18616 , w_18617 );
buf ( w_18616 , \7105_b1 );
not ( w_18616 , w_18620 );
not ( w_18617 , w_18621 );
and ( w_18620 , w_18621 , \7105_b0 );
or ( \7504_b1 , \7499_b1 , \7503_b1 );
xor ( \7504_b0 , \7499_b0 , w_18622 );
not ( w_18622 , w_18623 );
and ( w_18623 , \7503_b1 , \7503_b0 );
or ( \7505_b1 , \5906_b1 , \7117_b1 );
not ( \7117_b1 , w_18624 );
and ( \7505_b0 , \5906_b0 , w_18625 );
and ( w_18624 , w_18625 , \7117_b0 );
or ( \7506_b1 , \5918_b1 , \7115_b1 );
not ( \7115_b1 , w_18626 );
and ( \7506_b0 , \5918_b0 , w_18627 );
and ( w_18626 , w_18627 , \7115_b0 );
or ( \7507_b1 , \7505_b1 , w_18629 );
not ( w_18629 , w_18630 );
and ( \7507_b0 , \7505_b0 , w_18631 );
and ( w_18630 ,  , w_18631 );
buf ( w_18629 , \7506_b1 );
not ( w_18629 , w_18632 );
not (  , w_18633 );
and ( w_18632 , w_18633 , \7506_b0 );
or ( \7508_b1 , \7507_b1 , w_18634 );
xor ( \7508_b0 , \7507_b0 , w_18636 );
not ( w_18636 , w_18637 );
and ( w_18637 , w_18634 , w_18635 );
buf ( w_18634 , \7123_b1 );
not ( w_18634 , w_18638 );
not ( w_18635 , w_18639 );
and ( w_18638 , w_18639 , \7123_b0 );
or ( \7509_b1 , \7504_b1 , \7508_b1 );
xor ( \7509_b0 , \7504_b0 , w_18640 );
not ( w_18640 , w_18641 );
and ( w_18641 , \7508_b1 , \7508_b0 );
or ( \7510_b1 , \5799_b1 , \7026_b1 );
not ( \7026_b1 , w_18642 );
and ( \7510_b0 , \5799_b0 , w_18643 );
and ( w_18642 , w_18643 , \7026_b0 );
or ( \7511_b1 , \5811_b1 , \7024_b1 );
not ( \7024_b1 , w_18644 );
and ( \7511_b0 , \5811_b0 , w_18645 );
and ( w_18644 , w_18645 , \7024_b0 );
or ( \7512_b1 , \7510_b1 , w_18647 );
not ( w_18647 , w_18648 );
and ( \7512_b0 , \7510_b0 , w_18649 );
and ( w_18648 ,  , w_18649 );
buf ( w_18647 , \7511_b1 );
not ( w_18647 , w_18650 );
not (  , w_18651 );
and ( w_18650 , w_18651 , \7511_b0 );
or ( \7513_b1 , \7512_b1 , w_18652 );
xor ( \7513_b0 , \7512_b0 , w_18654 );
not ( w_18654 , w_18655 );
and ( w_18655 , w_18652 , w_18653 );
buf ( w_18652 , \7032_b1 );
not ( w_18652 , w_18656 );
not ( w_18653 , w_18657 );
and ( w_18656 , w_18657 , \7032_b0 );
or ( \7514_b1 , \5819_b1 , \7043_b1 );
not ( \7043_b1 , w_18658 );
and ( \7514_b0 , \5819_b0 , w_18659 );
and ( w_18658 , w_18659 , \7043_b0 );
or ( \7515_b1 , \5831_b1 , \7041_b1 );
not ( \7041_b1 , w_18660 );
and ( \7515_b0 , \5831_b0 , w_18661 );
and ( w_18660 , w_18661 , \7041_b0 );
or ( \7516_b1 , \7514_b1 , w_18663 );
not ( w_18663 , w_18664 );
and ( \7516_b0 , \7514_b0 , w_18665 );
and ( w_18664 ,  , w_18665 );
buf ( w_18663 , \7515_b1 );
not ( w_18663 , w_18666 );
not (  , w_18667 );
and ( w_18666 , w_18667 , \7515_b0 );
or ( \7517_b1 , \7516_b1 , w_18668 );
xor ( \7517_b0 , \7516_b0 , w_18670 );
not ( w_18670 , w_18671 );
and ( w_18671 , w_18668 , w_18669 );
buf ( w_18668 , \7049_b1 );
not ( w_18668 , w_18672 );
not ( w_18669 , w_18673 );
and ( w_18672 , w_18673 , \7049_b0 );
or ( \7518_b1 , \7513_b1 , \7517_b1 );
xor ( \7518_b0 , \7513_b0 , w_18674 );
not ( w_18674 , w_18675 );
and ( w_18675 , \7517_b1 , \7517_b0 );
or ( \7519_b1 , \5842_b1 , \7061_b1 );
not ( \7061_b1 , w_18676 );
and ( \7519_b0 , \5842_b0 , w_18677 );
and ( w_18676 , w_18677 , \7061_b0 );
or ( \7520_b1 , \5854_b1 , \7059_b1 );
not ( \7059_b1 , w_18678 );
and ( \7520_b0 , \5854_b0 , w_18679 );
and ( w_18678 , w_18679 , \7059_b0 );
or ( \7521_b1 , \7519_b1 , w_18681 );
not ( w_18681 , w_18682 );
and ( \7521_b0 , \7519_b0 , w_18683 );
and ( w_18682 ,  , w_18683 );
buf ( w_18681 , \7520_b1 );
not ( w_18681 , w_18684 );
not (  , w_18685 );
and ( w_18684 , w_18685 , \7520_b0 );
or ( \7522_b1 , \7521_b1 , w_18686 );
xor ( \7522_b0 , \7521_b0 , w_18688 );
not ( w_18688 , w_18689 );
and ( w_18689 , w_18686 , w_18687 );
buf ( w_18686 , \7067_b1 );
not ( w_18686 , w_18690 );
not ( w_18687 , w_18691 );
and ( w_18690 , w_18691 , \7067_b0 );
or ( \7523_b1 , \7518_b1 , \7522_b1 );
xor ( \7523_b0 , \7518_b0 , w_18692 );
not ( w_18692 , w_18693 );
and ( w_18693 , \7522_b1 , \7522_b0 );
or ( \7524_b1 , \7509_b1 , \7523_b1 );
xor ( \7524_b0 , \7509_b0 , w_18694 );
not ( w_18694 , w_18695 );
and ( w_18695 , \7523_b1 , \7523_b0 );
or ( \7525_b1 , \5758_b1 , \6991_b1 );
not ( \6991_b1 , w_18696 );
and ( \7525_b0 , \5758_b0 , w_18697 );
and ( w_18696 , w_18697 , \6991_b0 );
or ( \7526_b1 , \5770_b1 , \6988_b1 );
not ( \6988_b1 , w_18698 );
and ( \7526_b0 , \5770_b0 , w_18699 );
and ( w_18698 , w_18699 , \6988_b0 );
or ( \7527_b1 , \7525_b1 , w_18701 );
not ( w_18701 , w_18702 );
and ( \7527_b0 , \7525_b0 , w_18703 );
and ( w_18702 ,  , w_18703 );
buf ( w_18701 , \7526_b1 );
not ( w_18701 , w_18704 );
not (  , w_18705 );
and ( w_18704 , w_18705 , \7526_b0 );
or ( \7528_b1 , \7527_b1 , w_18706 );
xor ( \7528_b0 , \7527_b0 , w_18708 );
not ( w_18708 , w_18709 );
and ( w_18709 , w_18706 , w_18707 );
buf ( w_18706 , \6985_b1 );
not ( w_18706 , w_18710 );
not ( w_18707 , w_18711 );
and ( w_18710 , w_18711 , \6985_b0 );
or ( \7529_b1 , \5797_b1 , \7528_b1 );
xor ( \7529_b0 , \5797_b0 , w_18712 );
not ( w_18712 , w_18713 );
and ( w_18713 , \7528_b1 , \7528_b0 );
or ( \7530_b1 , \5780_b1 , \7006_b1 );
not ( \7006_b1 , w_18714 );
and ( \7530_b0 , \5780_b0 , w_18715 );
and ( w_18714 , w_18715 , \7006_b0 );
or ( \7531_b1 , \5792_b1 , \7004_b1 );
not ( \7004_b1 , w_18716 );
and ( \7531_b0 , \5792_b0 , w_18717 );
and ( w_18716 , w_18717 , \7004_b0 );
or ( \7532_b1 , \7530_b1 , w_18719 );
not ( w_18719 , w_18720 );
and ( \7532_b0 , \7530_b0 , w_18721 );
and ( w_18720 ,  , w_18721 );
buf ( w_18719 , \7531_b1 );
not ( w_18719 , w_18722 );
not (  , w_18723 );
and ( w_18722 , w_18723 , \7531_b0 );
or ( \7533_b1 , \7532_b1 , w_18724 );
xor ( \7533_b0 , \7532_b0 , w_18726 );
not ( w_18726 , w_18727 );
and ( w_18727 , w_18724 , w_18725 );
buf ( w_18724 , \7012_b1 );
not ( w_18724 , w_18728 );
not ( w_18725 , w_18729 );
and ( w_18728 , w_18729 , \7012_b0 );
or ( \7534_b1 , \7529_b1 , \7533_b1 );
xor ( \7534_b0 , \7529_b0 , w_18730 );
not ( w_18730 , w_18731 );
and ( w_18731 , \7533_b1 , \7533_b0 );
or ( \7535_b1 , \7524_b1 , \7534_b1 );
xor ( \7535_b0 , \7524_b0 , w_18732 );
not ( w_18732 , w_18733 );
and ( w_18733 , \7534_b1 , \7534_b0 );
or ( \7536_b1 , \6065_b1 , w_18735 );
not ( w_18735 , w_18736 );
and ( \7536_b0 , \6065_b0 , w_18737 );
and ( w_18736 ,  , w_18737 );
buf ( w_18735 , \5788_b1 );
not ( w_18735 , w_18738 );
not (  , w_18739 );
and ( w_18738 , w_18739 , \5788_b0 );
or ( \7537_b1 , \7536_b1 , w_18740 );
xor ( \7537_b0 , \7536_b0 , w_18742 );
not ( w_18742 , w_18743 );
and ( w_18743 , w_18740 , w_18741 );
buf ( w_18740 , \5797_b1 );
not ( w_18740 , w_18744 );
not ( w_18741 , w_18745 );
and ( w_18744 , w_18745 , \5797_b0 );
or ( \7538_b1 , \5986_b1 , \7192_b1 );
not ( \7192_b1 , w_18746 );
and ( \7538_b0 , \5986_b0 , w_18747 );
and ( w_18746 , w_18747 , \7192_b0 );
or ( \7539_b1 , \5998_b1 , \7190_b1 );
not ( \7190_b1 , w_18748 );
and ( \7539_b0 , \5998_b0 , w_18749 );
and ( w_18748 , w_18749 , \7190_b0 );
or ( \7540_b1 , \7538_b1 , w_18751 );
not ( w_18751 , w_18752 );
and ( \7540_b0 , \7538_b0 , w_18753 );
and ( w_18752 ,  , w_18753 );
buf ( w_18751 , \7539_b1 );
not ( w_18751 , w_18754 );
not (  , w_18755 );
and ( w_18754 , w_18755 , \7539_b0 );
or ( \7541_b1 , \7540_b1 , w_18756 );
xor ( \7541_b0 , \7540_b0 , w_18758 );
not ( w_18758 , w_18759 );
and ( w_18759 , w_18756 , w_18757 );
buf ( w_18756 , \7198_b1 );
not ( w_18756 , w_18760 );
not ( w_18757 , w_18761 );
and ( w_18760 , w_18761 , \7198_b0 );
or ( \7542_b1 , \6006_b1 , \7203_b1 );
not ( \7203_b1 , w_18762 );
and ( \7542_b0 , \6006_b0 , w_18763 );
and ( w_18762 , w_18763 , \7203_b0 );
or ( \7543_b1 , \6018_b1 , \7201_b1 );
not ( \7201_b1 , w_18764 );
and ( \7543_b0 , \6018_b0 , w_18765 );
and ( w_18764 , w_18765 , \7201_b0 );
or ( \7544_b1 , \7542_b1 , w_18767 );
not ( w_18767 , w_18768 );
and ( \7544_b0 , \7542_b0 , w_18769 );
and ( w_18768 ,  , w_18769 );
buf ( w_18767 , \7543_b1 );
not ( w_18767 , w_18770 );
not (  , w_18771 );
and ( w_18770 , w_18771 , \7543_b0 );
or ( \7545_b1 , \7544_b1 , w_18772 );
xor ( \7545_b0 , \7544_b0 , w_18774 );
not ( w_18774 , w_18775 );
and ( w_18775 , w_18772 , w_18773 );
buf ( w_18772 , \6824_b1 );
not ( w_18772 , w_18776 );
not ( w_18773 , w_18777 );
and ( w_18776 , w_18777 , \6824_b0 );
or ( \7546_b1 , \7541_b1 , \7545_b1 );
xor ( \7546_b0 , \7541_b0 , w_18778 );
not ( w_18778 , w_18779 );
and ( w_18779 , \7545_b1 , \7545_b0 );
or ( \7547_b1 , \6029_b1 , \5750_b1 );
not ( \5750_b1 , w_18780 );
and ( \7547_b0 , \6029_b0 , w_18781 );
and ( w_18780 , w_18781 , \5750_b0 );
or ( \7548_b1 , \6041_b1 , \5748_b1 );
not ( \5748_b1 , w_18782 );
and ( \7548_b0 , \6041_b0 , w_18783 );
and ( w_18782 , w_18783 , \5748_b0 );
or ( \7549_b1 , \7547_b1 , w_18785 );
not ( w_18785 , w_18786 );
and ( \7549_b0 , \7547_b0 , w_18787 );
and ( w_18786 ,  , w_18787 );
buf ( w_18785 , \7548_b1 );
not ( w_18785 , w_18788 );
not (  , w_18789 );
and ( w_18788 , w_18789 , \7548_b0 );
or ( \7550_b1 , \7549_b1 , w_18790 );
xor ( \7550_b0 , \7549_b0 , w_18792 );
not ( w_18792 , w_18793 );
and ( w_18793 , w_18790 , w_18791 );
buf ( w_18790 , \5755_b1 );
not ( w_18790 , w_18794 );
not ( w_18791 , w_18795 );
and ( w_18794 , w_18795 , \5755_b0 );
or ( \7551_b1 , \7546_b1 , \7550_b1 );
xor ( \7551_b0 , \7546_b0 , w_18796 );
not ( w_18796 , w_18797 );
and ( w_18797 , \7550_b1 , \7550_b0 );
or ( \7552_b1 , \7537_b1 , \7551_b1 );
xor ( \7552_b0 , \7537_b0 , w_18798 );
not ( w_18798 , w_18799 );
and ( w_18799 , \7551_b1 , \7551_b0 );
or ( \7553_b1 , \5925_b1 , \7140_b1 );
not ( \7140_b1 , w_18800 );
and ( \7553_b0 , \5925_b0 , w_18801 );
and ( w_18800 , w_18801 , \7140_b0 );
or ( \7554_b1 , \5937_b1 , \7138_b1 );
not ( \7138_b1 , w_18802 );
and ( \7554_b0 , \5937_b0 , w_18803 );
and ( w_18802 , w_18803 , \7138_b0 );
or ( \7555_b1 , \7553_b1 , w_18805 );
not ( w_18805 , w_18806 );
and ( \7555_b0 , \7553_b0 , w_18807 );
and ( w_18806 ,  , w_18807 );
buf ( w_18805 , \7554_b1 );
not ( w_18805 , w_18808 );
not (  , w_18809 );
and ( w_18808 , w_18809 , \7554_b0 );
or ( \7556_b1 , \7555_b1 , w_18810 );
xor ( \7556_b0 , \7555_b0 , w_18812 );
not ( w_18812 , w_18813 );
and ( w_18813 , w_18810 , w_18811 );
buf ( w_18810 , \7146_b1 );
not ( w_18810 , w_18814 );
not ( w_18811 , w_18815 );
and ( w_18814 , w_18815 , \7146_b0 );
or ( \7557_b1 , \5945_b1 , \7157_b1 );
not ( \7157_b1 , w_18816 );
and ( \7557_b0 , \5945_b0 , w_18817 );
and ( w_18816 , w_18817 , \7157_b0 );
or ( \7558_b1 , \5957_b1 , \7155_b1 );
not ( \7155_b1 , w_18818 );
and ( \7558_b0 , \5957_b0 , w_18819 );
and ( w_18818 , w_18819 , \7155_b0 );
or ( \7559_b1 , \7557_b1 , w_18821 );
not ( w_18821 , w_18822 );
and ( \7559_b0 , \7557_b0 , w_18823 );
and ( w_18822 ,  , w_18823 );
buf ( w_18821 , \7558_b1 );
not ( w_18821 , w_18824 );
not (  , w_18825 );
and ( w_18824 , w_18825 , \7558_b0 );
or ( \7560_b1 , \7559_b1 , w_18826 );
xor ( \7560_b0 , \7559_b0 , w_18828 );
not ( w_18828 , w_18829 );
and ( w_18829 , w_18826 , w_18827 );
buf ( w_18826 , \7163_b1 );
not ( w_18826 , w_18830 );
not ( w_18827 , w_18831 );
and ( w_18830 , w_18831 , \7163_b0 );
or ( \7561_b1 , \7556_b1 , \7560_b1 );
xor ( \7561_b0 , \7556_b0 , w_18832 );
not ( w_18832 , w_18833 );
and ( w_18833 , \7560_b1 , \7560_b0 );
or ( \7562_b1 , \5967_b1 , \7175_b1 );
not ( \7175_b1 , w_18834 );
and ( \7562_b0 , \5967_b0 , w_18835 );
and ( w_18834 , w_18835 , \7175_b0 );
or ( \7563_b1 , \5979_b1 , \7173_b1 );
not ( \7173_b1 , w_18836 );
and ( \7563_b0 , \5979_b0 , w_18837 );
and ( w_18836 , w_18837 , \7173_b0 );
or ( \7564_b1 , \7562_b1 , w_18839 );
not ( w_18839 , w_18840 );
and ( \7564_b0 , \7562_b0 , w_18841 );
and ( w_18840 ,  , w_18841 );
buf ( w_18839 , \7563_b1 );
not ( w_18839 , w_18842 );
not (  , w_18843 );
and ( w_18842 , w_18843 , \7563_b0 );
or ( \7565_b1 , \7564_b1 , w_18844 );
xor ( \7565_b0 , \7564_b0 , w_18846 );
not ( w_18846 , w_18847 );
and ( w_18847 , w_18844 , w_18845 );
buf ( w_18844 , \7181_b1 );
not ( w_18844 , w_18848 );
not ( w_18845 , w_18849 );
and ( w_18848 , w_18849 , \7181_b0 );
or ( \7566_b1 , \7561_b1 , \7565_b1 );
xor ( \7566_b0 , \7561_b0 , w_18850 );
not ( w_18850 , w_18851 );
and ( w_18851 , \7565_b1 , \7565_b0 );
or ( \7567_b1 , \7552_b1 , \7566_b1 );
xor ( \7567_b0 , \7552_b0 , w_18852 );
not ( w_18852 , w_18853 );
and ( w_18853 , \7566_b1 , \7566_b0 );
or ( \7568_b1 , \7535_b1 , \7567_b1 );
xor ( \7568_b0 , \7535_b0 , w_18854 );
not ( w_18854 , w_18855 );
and ( w_18855 , \7567_b1 , \7567_b0 );
or ( \7569_b1 , \7377_b1 , \7381_b1 );
not ( \7381_b1 , w_18856 );
and ( \7569_b0 , \7377_b0 , w_18857 );
and ( w_18856 , w_18857 , \7381_b0 );
or ( \7570_b1 , \7381_b1 , \7386_b1 );
not ( \7386_b1 , w_18858 );
and ( \7570_b0 , \7381_b0 , w_18859 );
and ( w_18858 , w_18859 , \7386_b0 );
or ( \7571_b1 , \7377_b1 , \7386_b1 );
not ( \7386_b1 , w_18860 );
and ( \7571_b0 , \7377_b0 , w_18861 );
and ( w_18860 , w_18861 , \7386_b0 );
or ( \7573_b1 , \7431_b1 , \7435_b1 );
not ( \7435_b1 , w_18862 );
and ( \7573_b0 , \7431_b0 , w_18863 );
and ( w_18862 , w_18863 , \7435_b0 );
or ( \7574_b1 , \7435_b1 , \7440_b1 );
not ( \7440_b1 , w_18864 );
and ( \7574_b0 , \7435_b0 , w_18865 );
and ( w_18864 , w_18865 , \7440_b0 );
or ( \7575_b1 , \7431_b1 , \7440_b1 );
not ( \7440_b1 , w_18866 );
and ( \7575_b0 , \7431_b0 , w_18867 );
and ( w_18866 , w_18867 , \7440_b0 );
or ( \7577_b1 , \7572_b1 , \7576_b1 );
xor ( \7577_b0 , \7572_b0 , w_18868 );
not ( w_18868 , w_18869 );
and ( w_18869 , \7576_b1 , \7576_b0 );
or ( \7578_b1 , \6048_b1 , \5768_b1 );
not ( \5768_b1 , w_18870 );
and ( \7578_b0 , \6048_b0 , w_18871 );
and ( w_18870 , w_18871 , \5768_b0 );
or ( \7579_b1 , \6057_b1 , \5766_b1 );
not ( \5766_b1 , w_18872 );
and ( \7579_b0 , \6057_b0 , w_18873 );
and ( w_18872 , w_18873 , \5766_b0 );
or ( \7580_b1 , \7578_b1 , w_18875 );
not ( w_18875 , w_18876 );
and ( \7580_b0 , \7578_b0 , w_18877 );
and ( w_18876 ,  , w_18877 );
buf ( w_18875 , \7579_b1 );
not ( w_18875 , w_18878 );
not (  , w_18879 );
and ( w_18878 , w_18879 , \7579_b0 );
or ( \7581_b1 , \7580_b1 , w_18880 );
xor ( \7581_b0 , \7580_b0 , w_18882 );
not ( w_18882 , w_18883 );
and ( w_18883 , w_18880 , w_18881 );
buf ( w_18880 , \5775_b1 );
not ( w_18880 , w_18884 );
not ( w_18881 , w_18885 );
and ( w_18884 , w_18885 , \5775_b0 );
or ( \7582_b1 , \7577_b1 , \7581_b1 );
xor ( \7582_b0 , \7577_b0 , w_18886 );
not ( w_18886 , w_18887 );
and ( w_18887 , \7581_b1 , \7581_b0 );
or ( \7583_b1 , \7568_b1 , \7582_b1 );
xor ( \7583_b0 , \7568_b0 , w_18888 );
not ( w_18888 , w_18889 );
and ( w_18889 , \7582_b1 , \7582_b0 );
or ( \7584_b1 , \7494_b1 , \7583_b1 );
not ( \7583_b1 , w_18890 );
and ( \7584_b0 , \7494_b0 , w_18891 );
and ( w_18890 , w_18891 , \7583_b0 );
or ( \7585_b1 , \7359_b1 , \7583_b1 );
not ( \7583_b1 , w_18892 );
and ( \7585_b0 , \7359_b0 , w_18893 );
and ( w_18892 , w_18893 , \7583_b0 );
or ( \7587_b1 , \7346_b1 , \7350_b1 );
not ( \7350_b1 , w_18894 );
and ( \7587_b0 , \7346_b0 , w_18895 );
and ( w_18894 , w_18895 , \7350_b0 );
or ( \7588_b1 , \7350_b1 , \7355_b1 );
not ( \7355_b1 , w_18896 );
and ( \7588_b0 , \7350_b0 , w_18897 );
and ( w_18896 , w_18897 , \7355_b0 );
or ( \7589_b1 , \7346_b1 , \7355_b1 );
not ( \7355_b1 , w_18898 );
and ( \7589_b0 , \7346_b0 , w_18899 );
and ( w_18898 , w_18899 , \7355_b0 );
or ( \7591_b1 , \7422_b1 , \7426_b1 );
not ( \7426_b1 , w_18900 );
and ( \7591_b0 , \7422_b0 , w_18901 );
and ( w_18900 , w_18901 , \7426_b0 );
or ( \7592_b1 , \7426_b1 , \7441_b1 );
not ( \7441_b1 , w_18902 );
and ( \7592_b0 , \7426_b0 , w_18903 );
and ( w_18902 , w_18903 , \7441_b0 );
or ( \7593_b1 , \7422_b1 , \7441_b1 );
not ( \7441_b1 , w_18904 );
and ( \7593_b0 , \7422_b0 , w_18905 );
and ( w_18904 , w_18905 , \7441_b0 );
or ( \7595_b1 , \7590_b1 , \7594_b1 );
xor ( \7595_b0 , \7590_b0 , w_18906 );
not ( w_18906 , w_18907 );
and ( w_18907 , \7594_b1 , \7594_b0 );
or ( \7596_b1 , \7387_b1 , \7401_b1 );
not ( \7401_b1 , w_18908 );
and ( \7596_b0 , \7387_b0 , w_18909 );
and ( w_18908 , w_18909 , \7401_b0 );
or ( \7597_b1 , \7401_b1 , \7416_b1 );
not ( \7416_b1 , w_18910 );
and ( \7597_b0 , \7401_b0 , w_18911 );
and ( w_18910 , w_18911 , \7416_b0 );
or ( \7598_b1 , \7387_b1 , \7416_b1 );
not ( \7416_b1 , w_18912 );
and ( \7598_b0 , \7387_b0 , w_18913 );
and ( w_18912 , w_18913 , \7416_b0 );
or ( \7600_b1 , \7595_b1 , \7599_b1 );
xor ( \7600_b0 , \7595_b0 , w_18914 );
not ( w_18914 , w_18915 );
and ( w_18915 , \7599_b1 , \7599_b0 );
or ( \7601_b1 , \7483_b1 , \7487_b1 );
not ( \7487_b1 , w_18916 );
and ( \7601_b0 , \7483_b0 , w_18917 );
and ( w_18916 , w_18917 , \7487_b0 );
or ( \7602_b1 , \7487_b1 , \7492_b1 );
not ( \7492_b1 , w_18918 );
and ( \7602_b0 , \7487_b0 , w_18919 );
and ( w_18918 , w_18919 , \7492_b0 );
or ( \7603_b1 , \7483_b1 , \7492_b1 );
not ( \7492_b1 , w_18920 );
and ( \7603_b0 , \7483_b0 , w_18921 );
and ( w_18920 , w_18921 , \7492_b0 );
or ( \7605_b1 , \7373_b1 , \7417_b1 );
not ( \7417_b1 , w_18922 );
and ( \7605_b0 , \7373_b0 , w_18923 );
and ( w_18922 , w_18923 , \7417_b0 );
or ( \7606_b1 , \7417_b1 , \7442_b1 );
not ( \7442_b1 , w_18924 );
and ( \7606_b0 , \7417_b0 , w_18925 );
and ( w_18924 , w_18925 , \7442_b0 );
or ( \7607_b1 , \7373_b1 , \7442_b1 );
not ( \7442_b1 , w_18926 );
and ( \7607_b0 , \7373_b0 , w_18927 );
and ( w_18926 , w_18927 , \7442_b0 );
or ( \7609_b1 , \7604_b1 , \7608_b1 );
xor ( \7609_b0 , \7604_b0 , w_18928 );
not ( w_18928 , w_18929 );
and ( w_18929 , \7608_b1 , \7608_b0 );
or ( \7610_b1 , \7363_b1 , \7367_b1 );
not ( \7367_b1 , w_18930 );
and ( \7610_b0 , \7363_b0 , w_18931 );
and ( w_18930 , w_18931 , \7367_b0 );
or ( \7611_b1 , \7367_b1 , \7372_b1 );
not ( \7372_b1 , w_18932 );
and ( \7611_b0 , \7367_b0 , w_18933 );
and ( w_18932 , w_18933 , \7372_b0 );
or ( \7612_b1 , \7363_b1 , \7372_b1 );
not ( \7372_b1 , w_18934 );
and ( \7612_b0 , \7363_b0 , w_18935 );
and ( w_18934 , w_18935 , \7372_b0 );
or ( \7614_b1 , \7406_b1 , \7410_b1 );
not ( \7410_b1 , w_18936 );
and ( \7614_b0 , \7406_b0 , w_18937 );
and ( w_18936 , w_18937 , \7410_b0 );
or ( \7615_b1 , \7410_b1 , \7415_b1 );
not ( \7415_b1 , w_18938 );
and ( \7615_b0 , \7410_b0 , w_18939 );
and ( w_18938 , w_18939 , \7415_b0 );
or ( \7616_b1 , \7406_b1 , \7415_b1 );
not ( \7415_b1 , w_18940 );
and ( \7616_b0 , \7406_b0 , w_18941 );
and ( w_18940 , w_18941 , \7415_b0 );
or ( \7618_b1 , \7613_b1 , \7617_b1 );
xor ( \7618_b0 , \7613_b0 , w_18942 );
not ( w_18942 , w_18943 );
and ( w_18943 , \7617_b1 , \7617_b0 );
or ( \7619_b1 , \7391_b1 , \7395_b1 );
not ( \7395_b1 , w_18944 );
and ( \7619_b0 , \7391_b0 , w_18945 );
and ( w_18944 , w_18945 , \7395_b0 );
or ( \7620_b1 , \7395_b1 , \7400_b1 );
not ( \7400_b1 , w_18946 );
and ( \7620_b0 , \7395_b0 , w_18947 );
and ( w_18946 , w_18947 , \7400_b0 );
or ( \7621_b1 , \7391_b1 , \7400_b1 );
not ( \7400_b1 , w_18948 );
and ( \7621_b0 , \7391_b0 , w_18949 );
and ( w_18948 , w_18949 , \7400_b0 );
or ( \7623_b1 , \7618_b1 , \7622_b1 );
xor ( \7623_b0 , \7618_b0 , w_18950 );
not ( w_18950 , w_18951 );
and ( w_18951 , \7622_b1 , \7622_b0 );
or ( \7624_b1 , \7609_b1 , \7623_b1 );
xor ( \7624_b0 , \7609_b0 , w_18952 );
not ( w_18952 , w_18953 );
and ( w_18953 , \7623_b1 , \7623_b0 );
or ( \7625_b1 , \7600_b1 , \7624_b1 );
not ( \7624_b1 , w_18954 );
and ( \7625_b0 , \7600_b0 , w_18955 );
and ( w_18954 , w_18955 , \7624_b0 );
or ( \7626_b1 , \7586_b1 , \7625_b1 );
xor ( \7626_b0 , \7586_b0 , w_18956 );
not ( w_18956 , w_18957 );
and ( w_18957 , \7625_b1 , \7625_b0 );
or ( \7627_b1 , \7604_b1 , \7608_b1 );
not ( \7608_b1 , w_18958 );
and ( \7627_b0 , \7604_b0 , w_18959 );
and ( w_18958 , w_18959 , \7608_b0 );
or ( \7628_b1 , \7608_b1 , \7623_b1 );
not ( \7623_b1 , w_18960 );
and ( \7628_b0 , \7608_b0 , w_18961 );
and ( w_18960 , w_18961 , \7623_b0 );
or ( \7629_b1 , \7604_b1 , \7623_b1 );
not ( \7623_b1 , w_18962 );
and ( \7629_b0 , \7604_b0 , w_18963 );
and ( w_18962 , w_18963 , \7623_b0 );
or ( \7631_b1 , \7509_b1 , \7523_b1 );
not ( \7523_b1 , w_18964 );
and ( \7631_b0 , \7509_b0 , w_18965 );
and ( w_18964 , w_18965 , \7523_b0 );
or ( \7632_b1 , \7523_b1 , \7534_b1 );
not ( \7534_b1 , w_18966 );
and ( \7632_b0 , \7523_b0 , w_18967 );
and ( w_18966 , w_18967 , \7534_b0 );
or ( \7633_b1 , \7509_b1 , \7534_b1 );
not ( \7534_b1 , w_18968 );
and ( \7633_b0 , \7509_b0 , w_18969 );
and ( w_18968 , w_18969 , \7534_b0 );
or ( \7635_b1 , \5831_b1 , \7043_b1 );
not ( \7043_b1 , w_18970 );
and ( \7635_b0 , \5831_b0 , w_18971 );
and ( w_18970 , w_18971 , \7043_b0 );
or ( \7636_b1 , \5799_b1 , \7041_b1 );
not ( \7041_b1 , w_18972 );
and ( \7636_b0 , \5799_b0 , w_18973 );
and ( w_18972 , w_18973 , \7041_b0 );
or ( \7637_b1 , \7635_b1 , w_18975 );
not ( w_18975 , w_18976 );
and ( \7637_b0 , \7635_b0 , w_18977 );
and ( w_18976 ,  , w_18977 );
buf ( w_18975 , \7636_b1 );
not ( w_18975 , w_18978 );
not (  , w_18979 );
and ( w_18978 , w_18979 , \7636_b0 );
or ( \7638_b1 , \7637_b1 , w_18980 );
xor ( \7638_b0 , \7637_b0 , w_18982 );
not ( w_18982 , w_18983 );
and ( w_18983 , w_18980 , w_18981 );
buf ( w_18980 , \7049_b1 );
not ( w_18980 , w_18984 );
not ( w_18981 , w_18985 );
and ( w_18984 , w_18985 , \7049_b0 );
or ( \7639_b1 , \5854_b1 , \7061_b1 );
not ( \7061_b1 , w_18986 );
and ( \7639_b0 , \5854_b0 , w_18987 );
and ( w_18986 , w_18987 , \7061_b0 );
or ( \7640_b1 , \5819_b1 , \7059_b1 );
not ( \7059_b1 , w_18988 );
and ( \7640_b0 , \5819_b0 , w_18989 );
and ( w_18988 , w_18989 , \7059_b0 );
or ( \7641_b1 , \7639_b1 , w_18991 );
not ( w_18991 , w_18992 );
and ( \7641_b0 , \7639_b0 , w_18993 );
and ( w_18992 ,  , w_18993 );
buf ( w_18991 , \7640_b1 );
not ( w_18991 , w_18994 );
not (  , w_18995 );
and ( w_18994 , w_18995 , \7640_b0 );
or ( \7642_b1 , \7641_b1 , w_18996 );
xor ( \7642_b0 , \7641_b0 , w_18998 );
not ( w_18998 , w_18999 );
and ( w_18999 , w_18996 , w_18997 );
buf ( w_18996 , \7067_b1 );
not ( w_18996 , w_19000 );
not ( w_18997 , w_19001 );
and ( w_19000 , w_19001 , \7067_b0 );
or ( \7643_b1 , \7638_b1 , \7642_b1 );
xor ( \7643_b0 , \7638_b0 , w_19002 );
not ( w_19002 , w_19003 );
and ( w_19003 , \7642_b1 , \7642_b0 );
or ( \7644_b1 , \5873_b1 , \7082_b1 );
not ( \7082_b1 , w_19004 );
and ( \7644_b0 , \5873_b0 , w_19005 );
and ( w_19004 , w_19005 , \7082_b0 );
or ( \7645_b1 , \5842_b1 , \7080_b1 );
not ( \7080_b1 , w_19006 );
and ( \7645_b0 , \5842_b0 , w_19007 );
and ( w_19006 , w_19007 , \7080_b0 );
or ( \7646_b1 , \7644_b1 , w_19009 );
not ( w_19009 , w_19010 );
and ( \7646_b0 , \7644_b0 , w_19011 );
and ( w_19010 ,  , w_19011 );
buf ( w_19009 , \7645_b1 );
not ( w_19009 , w_19012 );
not (  , w_19013 );
and ( w_19012 , w_19013 , \7645_b0 );
or ( \7647_b1 , \7646_b1 , w_19014 );
xor ( \7647_b0 , \7646_b0 , w_19016 );
not ( w_19016 , w_19017 );
and ( w_19017 , w_19014 , w_19015 );
buf ( w_19014 , \7088_b1 );
not ( w_19014 , w_19018 );
not ( w_19015 , w_19019 );
and ( w_19018 , w_19019 , \7088_b0 );
or ( \7648_b1 , \7643_b1 , \7647_b1 );
xor ( \7648_b0 , \7643_b0 , w_19020 );
not ( w_19020 , w_19021 );
and ( w_19021 , \7647_b1 , \7647_b0 );
or ( \7649_b1 , \7634_b1 , \7648_b1 );
xor ( \7649_b0 , \7634_b0 , w_19022 );
not ( w_19022 , w_19023 );
and ( w_19023 , \7648_b1 , \7648_b0 );
or ( \7650_b1 , \5770_b1 , \6991_b1 );
not ( \6991_b1 , w_19024 );
and ( \7650_b0 , \5770_b0 , w_19025 );
and ( w_19024 , w_19025 , \6991_b0 );
or ( \7651_b1 , \5737_b1 , \6988_b1 );
not ( \6988_b1 , w_19026 );
and ( \7651_b0 , \5737_b0 , w_19027 );
and ( w_19026 , w_19027 , \6988_b0 );
or ( \7652_b1 , \7650_b1 , w_19029 );
not ( w_19029 , w_19030 );
and ( \7652_b0 , \7650_b0 , w_19031 );
and ( w_19030 ,  , w_19031 );
buf ( w_19029 , \7651_b1 );
not ( w_19029 , w_19032 );
not (  , w_19033 );
and ( w_19032 , w_19033 , \7651_b0 );
or ( \7653_b1 , \7652_b1 , w_19034 );
xor ( \7653_b0 , \7652_b0 , w_19036 );
not ( w_19036 , w_19037 );
and ( w_19037 , w_19034 , w_19035 );
buf ( w_19034 , \6985_b1 );
not ( w_19034 , w_19038 );
not ( w_19035 , w_19039 );
and ( w_19038 , w_19039 , \6985_b0 );
or ( \7654_b1 , \5792_b1 , \7006_b1 );
not ( \7006_b1 , w_19040 );
and ( \7654_b0 , \5792_b0 , w_19041 );
and ( w_19040 , w_19041 , \7006_b0 );
or ( \7655_b1 , \5758_b1 , \7004_b1 );
not ( \7004_b1 , w_19042 );
and ( \7655_b0 , \5758_b0 , w_19043 );
and ( w_19042 , w_19043 , \7004_b0 );
or ( \7656_b1 , \7654_b1 , w_19045 );
not ( w_19045 , w_19046 );
and ( \7656_b0 , \7654_b0 , w_19047 );
and ( w_19046 ,  , w_19047 );
buf ( w_19045 , \7655_b1 );
not ( w_19045 , w_19048 );
not (  , w_19049 );
and ( w_19048 , w_19049 , \7655_b0 );
or ( \7657_b1 , \7656_b1 , w_19050 );
xor ( \7657_b0 , \7656_b0 , w_19052 );
not ( w_19052 , w_19053 );
and ( w_19053 , w_19050 , w_19051 );
buf ( w_19050 , \7012_b1 );
not ( w_19050 , w_19054 );
not ( w_19051 , w_19055 );
and ( w_19054 , w_19055 , \7012_b0 );
or ( \7658_b1 , \7653_b1 , \7657_b1 );
xor ( \7658_b0 , \7653_b0 , w_19056 );
not ( w_19056 , w_19057 );
and ( w_19057 , \7657_b1 , \7657_b0 );
or ( \7659_b1 , \5811_b1 , \7026_b1 );
not ( \7026_b1 , w_19058 );
and ( \7659_b0 , \5811_b0 , w_19059 );
and ( w_19058 , w_19059 , \7026_b0 );
or ( \7660_b1 , \5780_b1 , \7024_b1 );
not ( \7024_b1 , w_19060 );
and ( \7660_b0 , \5780_b0 , w_19061 );
and ( w_19060 , w_19061 , \7024_b0 );
or ( \7661_b1 , \7659_b1 , w_19063 );
not ( w_19063 , w_19064 );
and ( \7661_b0 , \7659_b0 , w_19065 );
and ( w_19064 ,  , w_19065 );
buf ( w_19063 , \7660_b1 );
not ( w_19063 , w_19066 );
not (  , w_19067 );
and ( w_19066 , w_19067 , \7660_b0 );
or ( \7662_b1 , \7661_b1 , w_19068 );
xor ( \7662_b0 , \7661_b0 , w_19070 );
not ( w_19070 , w_19071 );
and ( w_19071 , w_19068 , w_19069 );
buf ( w_19068 , \7032_b1 );
not ( w_19068 , w_19072 );
not ( w_19069 , w_19073 );
and ( w_19072 , w_19073 , \7032_b0 );
or ( \7663_b1 , \7658_b1 , \7662_b1 );
xor ( \7663_b0 , \7658_b0 , w_19074 );
not ( w_19074 , w_19075 );
and ( w_19075 , \7662_b1 , \7662_b0 );
or ( \7664_b1 , \7649_b1 , \7663_b1 );
xor ( \7664_b0 , \7649_b0 , w_19076 );
not ( w_19076 , w_19077 );
and ( w_19077 , \7663_b1 , \7663_b0 );
or ( \7665_b1 , \7613_b1 , \7617_b1 );
not ( \7617_b1 , w_19078 );
and ( \7665_b0 , \7613_b0 , w_19079 );
and ( w_19078 , w_19079 , \7617_b0 );
or ( \7666_b1 , \7617_b1 , \7622_b1 );
not ( \7622_b1 , w_19080 );
and ( \7666_b0 , \7617_b0 , w_19081 );
and ( w_19080 , w_19081 , \7622_b0 );
or ( \7667_b1 , \7613_b1 , \7622_b1 );
not ( \7622_b1 , w_19082 );
and ( \7667_b0 , \7613_b0 , w_19083 );
and ( w_19082 , w_19083 , \7622_b0 );
or ( \7669_b1 , \7572_b1 , \7576_b1 );
not ( \7576_b1 , w_19084 );
and ( \7669_b0 , \7572_b0 , w_19085 );
and ( w_19084 , w_19085 , \7576_b0 );
or ( \7670_b1 , \7576_b1 , \7581_b1 );
not ( \7581_b1 , w_19086 );
and ( \7670_b0 , \7576_b0 , w_19087 );
and ( w_19086 , w_19087 , \7581_b0 );
or ( \7671_b1 , \7572_b1 , \7581_b1 );
not ( \7581_b1 , w_19088 );
and ( \7671_b0 , \7572_b0 , w_19089 );
and ( w_19088 , w_19089 , \7581_b0 );
or ( \7673_b1 , \7668_b1 , \7672_b1 );
xor ( \7673_b0 , \7668_b0 , w_19090 );
not ( w_19090 , w_19091 );
and ( w_19091 , \7672_b1 , \7672_b0 );
or ( \7674_b1 , \7537_b1 , \7551_b1 );
not ( \7551_b1 , w_19092 );
and ( \7674_b0 , \7537_b0 , w_19093 );
and ( w_19092 , w_19093 , \7551_b0 );
or ( \7675_b1 , \7551_b1 , \7566_b1 );
not ( \7566_b1 , w_19094 );
and ( \7675_b0 , \7551_b0 , w_19095 );
and ( w_19094 , w_19095 , \7566_b0 );
or ( \7676_b1 , \7537_b1 , \7566_b1 );
not ( \7566_b1 , w_19096 );
and ( \7676_b0 , \7537_b0 , w_19097 );
and ( w_19096 , w_19097 , \7566_b0 );
or ( \7678_b1 , \7673_b1 , \7677_b1 );
xor ( \7678_b0 , \7673_b0 , w_19098 );
not ( w_19098 , w_19099 );
and ( w_19099 , \7677_b1 , \7677_b0 );
or ( \7679_b1 , \7664_b1 , \7678_b1 );
xor ( \7679_b0 , \7664_b0 , w_19100 );
not ( w_19100 , w_19101 );
and ( w_19101 , \7678_b1 , \7678_b0 );
or ( \7680_b1 , \7630_b1 , \7679_b1 );
xor ( \7680_b0 , \7630_b0 , w_19102 );
not ( w_19102 , w_19103 );
and ( w_19103 , \7679_b1 , \7679_b0 );
or ( \7681_b1 , \7590_b1 , \7594_b1 );
not ( \7594_b1 , w_19104 );
and ( \7681_b0 , \7590_b0 , w_19105 );
and ( w_19104 , w_19105 , \7594_b0 );
or ( \7682_b1 , \7594_b1 , \7599_b1 );
not ( \7599_b1 , w_19106 );
and ( \7682_b0 , \7594_b0 , w_19107 );
and ( w_19106 , w_19107 , \7599_b0 );
or ( \7683_b1 , \7590_b1 , \7599_b1 );
not ( \7599_b1 , w_19108 );
and ( \7683_b0 , \7590_b0 , w_19109 );
and ( w_19108 , w_19109 , \7599_b0 );
or ( \7685_b1 , \7535_b1 , \7567_b1 );
not ( \7567_b1 , w_19110 );
and ( \7685_b0 , \7535_b0 , w_19111 );
and ( w_19110 , w_19111 , \7567_b0 );
or ( \7686_b1 , \7567_b1 , \7582_b1 );
not ( \7582_b1 , w_19112 );
and ( \7686_b0 , \7567_b0 , w_19113 );
and ( w_19112 , w_19113 , \7582_b0 );
or ( \7687_b1 , \7535_b1 , \7582_b1 );
not ( \7582_b1 , w_19114 );
and ( \7687_b0 , \7535_b0 , w_19115 );
and ( w_19114 , w_19115 , \7582_b0 );
or ( \7689_b1 , \7684_b1 , \7688_b1 );
xor ( \7689_b0 , \7684_b0 , w_19116 );
not ( w_19116 , w_19117 );
and ( w_19117 , \7688_b1 , \7688_b0 );
or ( \7690_b1 , \6018_b1 , \7203_b1 );
not ( \7203_b1 , w_19118 );
and ( \7690_b0 , \6018_b0 , w_19119 );
and ( w_19118 , w_19119 , \7203_b0 );
or ( \7691_b1 , \5986_b1 , \7201_b1 );
not ( \7201_b1 , w_19120 );
and ( \7691_b0 , \5986_b0 , w_19121 );
and ( w_19120 , w_19121 , \7201_b0 );
or ( \7692_b1 , \7690_b1 , w_19123 );
not ( w_19123 , w_19124 );
and ( \7692_b0 , \7690_b0 , w_19125 );
and ( w_19124 ,  , w_19125 );
buf ( w_19123 , \7691_b1 );
not ( w_19123 , w_19126 );
not (  , w_19127 );
and ( w_19126 , w_19127 , \7691_b0 );
or ( \7693_b1 , \7692_b1 , w_19128 );
xor ( \7693_b0 , \7692_b0 , w_19130 );
not ( w_19130 , w_19131 );
and ( w_19131 , w_19128 , w_19129 );
buf ( w_19128 , \6824_b1 );
not ( w_19128 , w_19132 );
not ( w_19129 , w_19133 );
and ( w_19132 , w_19133 , \6824_b0 );
or ( \7694_b1 , \6041_b1 , \5750_b1 );
not ( \5750_b1 , w_19134 );
and ( \7694_b0 , \6041_b0 , w_19135 );
and ( w_19134 , w_19135 , \5750_b0 );
or ( \7695_b1 , \6006_b1 , \5748_b1 );
not ( \5748_b1 , w_19136 );
and ( \7695_b0 , \6006_b0 , w_19137 );
and ( w_19136 , w_19137 , \5748_b0 );
or ( \7696_b1 , \7694_b1 , w_19139 );
not ( w_19139 , w_19140 );
and ( \7696_b0 , \7694_b0 , w_19141 );
and ( w_19140 ,  , w_19141 );
buf ( w_19139 , \7695_b1 );
not ( w_19139 , w_19142 );
not (  , w_19143 );
and ( w_19142 , w_19143 , \7695_b0 );
or ( \7697_b1 , \7696_b1 , w_19144 );
xor ( \7697_b0 , \7696_b0 , w_19146 );
not ( w_19146 , w_19147 );
and ( w_19147 , w_19144 , w_19145 );
buf ( w_19144 , \5755_b1 );
not ( w_19144 , w_19148 );
not ( w_19145 , w_19149 );
and ( w_19148 , w_19149 , \5755_b0 );
or ( \7698_b1 , \7693_b1 , \7697_b1 );
xor ( \7698_b0 , \7693_b0 , w_19150 );
not ( w_19150 , w_19151 );
and ( w_19151 , \7697_b1 , \7697_b0 );
or ( \7699_b1 , \6057_b1 , \5768_b1 );
not ( \5768_b1 , w_19152 );
and ( \7699_b0 , \6057_b0 , w_19153 );
and ( w_19152 , w_19153 , \5768_b0 );
or ( \7700_b1 , \6029_b1 , \5766_b1 );
not ( \5766_b1 , w_19154 );
and ( \7700_b0 , \6029_b0 , w_19155 );
and ( w_19154 , w_19155 , \5766_b0 );
or ( \7701_b1 , \7699_b1 , w_19157 );
not ( w_19157 , w_19158 );
and ( \7701_b0 , \7699_b0 , w_19159 );
and ( w_19158 ,  , w_19159 );
buf ( w_19157 , \7700_b1 );
not ( w_19157 , w_19160 );
not (  , w_19161 );
and ( w_19160 , w_19161 , \7700_b0 );
or ( \7702_b1 , \7701_b1 , w_19162 );
xor ( \7702_b0 , \7701_b0 , w_19164 );
not ( w_19164 , w_19165 );
and ( w_19165 , w_19162 , w_19163 );
buf ( w_19162 , \5775_b1 );
not ( w_19162 , w_19166 );
not ( w_19163 , w_19167 );
and ( w_19166 , w_19167 , \5775_b0 );
or ( \7703_b1 , \7698_b1 , \7702_b1 );
xor ( \7703_b0 , \7698_b0 , w_19168 );
not ( w_19168 , w_19169 );
and ( w_19169 , \7702_b1 , \7702_b0 );
or ( \7704_b1 , \5957_b1 , \7157_b1 );
not ( \7157_b1 , w_19170 );
and ( \7704_b0 , \5957_b0 , w_19171 );
and ( w_19170 , w_19171 , \7157_b0 );
or ( \7705_b1 , \5925_b1 , \7155_b1 );
not ( \7155_b1 , w_19172 );
and ( \7705_b0 , \5925_b0 , w_19173 );
and ( w_19172 , w_19173 , \7155_b0 );
or ( \7706_b1 , \7704_b1 , w_19175 );
not ( w_19175 , w_19176 );
and ( \7706_b0 , \7704_b0 , w_19177 );
and ( w_19176 ,  , w_19177 );
buf ( w_19175 , \7705_b1 );
not ( w_19175 , w_19178 );
not (  , w_19179 );
and ( w_19178 , w_19179 , \7705_b0 );
or ( \7707_b1 , \7706_b1 , w_19180 );
xor ( \7707_b0 , \7706_b0 , w_19182 );
not ( w_19182 , w_19183 );
and ( w_19183 , w_19180 , w_19181 );
buf ( w_19180 , \7163_b1 );
not ( w_19180 , w_19184 );
not ( w_19181 , w_19185 );
and ( w_19184 , w_19185 , \7163_b0 );
or ( \7708_b1 , \5979_b1 , \7175_b1 );
not ( \7175_b1 , w_19186 );
and ( \7708_b0 , \5979_b0 , w_19187 );
and ( w_19186 , w_19187 , \7175_b0 );
or ( \7709_b1 , \5945_b1 , \7173_b1 );
not ( \7173_b1 , w_19188 );
and ( \7709_b0 , \5945_b0 , w_19189 );
and ( w_19188 , w_19189 , \7173_b0 );
or ( \7710_b1 , \7708_b1 , w_19191 );
not ( w_19191 , w_19192 );
and ( \7710_b0 , \7708_b0 , w_19193 );
and ( w_19192 ,  , w_19193 );
buf ( w_19191 , \7709_b1 );
not ( w_19191 , w_19194 );
not (  , w_19195 );
and ( w_19194 , w_19195 , \7709_b0 );
or ( \7711_b1 , \7710_b1 , w_19196 );
xor ( \7711_b0 , \7710_b0 , w_19198 );
not ( w_19198 , w_19199 );
and ( w_19199 , w_19196 , w_19197 );
buf ( w_19196 , \7181_b1 );
not ( w_19196 , w_19200 );
not ( w_19197 , w_19201 );
and ( w_19200 , w_19201 , \7181_b0 );
or ( \7712_b1 , \7707_b1 , \7711_b1 );
xor ( \7712_b0 , \7707_b0 , w_19202 );
not ( w_19202 , w_19203 );
and ( w_19203 , \7711_b1 , \7711_b0 );
or ( \7713_b1 , \5998_b1 , \7192_b1 );
not ( \7192_b1 , w_19204 );
and ( \7713_b0 , \5998_b0 , w_19205 );
and ( w_19204 , w_19205 , \7192_b0 );
or ( \7714_b1 , \5967_b1 , \7190_b1 );
not ( \7190_b1 , w_19206 );
and ( \7714_b0 , \5967_b0 , w_19207 );
and ( w_19206 , w_19207 , \7190_b0 );
or ( \7715_b1 , \7713_b1 , w_19209 );
not ( w_19209 , w_19210 );
and ( \7715_b0 , \7713_b0 , w_19211 );
and ( w_19210 ,  , w_19211 );
buf ( w_19209 , \7714_b1 );
not ( w_19209 , w_19212 );
not (  , w_19213 );
and ( w_19212 , w_19213 , \7714_b0 );
or ( \7716_b1 , \7715_b1 , w_19214 );
xor ( \7716_b0 , \7715_b0 , w_19216 );
not ( w_19216 , w_19217 );
and ( w_19217 , w_19214 , w_19215 );
buf ( w_19214 , \7198_b1 );
not ( w_19214 , w_19218 );
not ( w_19215 , w_19219 );
and ( w_19218 , w_19219 , \7198_b0 );
or ( \7717_b1 , \7712_b1 , \7716_b1 );
xor ( \7717_b0 , \7712_b0 , w_19220 );
not ( w_19220 , w_19221 );
and ( w_19221 , \7716_b1 , \7716_b0 );
or ( \7718_b1 , \7703_b1 , \7717_b1 );
xor ( \7718_b0 , \7703_b0 , w_19222 );
not ( w_19222 , w_19223 );
and ( w_19223 , \7717_b1 , \7717_b0 );
or ( \7719_b1 , \5893_b1 , \7099_b1 );
not ( \7099_b1 , w_19224 );
and ( \7719_b0 , \5893_b0 , w_19225 );
and ( w_19224 , w_19225 , \7099_b0 );
or ( \7720_b1 , \5861_b1 , \7097_b1 );
not ( \7097_b1 , w_19226 );
and ( \7720_b0 , \5861_b0 , w_19227 );
and ( w_19226 , w_19227 , \7097_b0 );
or ( \7721_b1 , \7719_b1 , w_19229 );
not ( w_19229 , w_19230 );
and ( \7721_b0 , \7719_b0 , w_19231 );
and ( w_19230 ,  , w_19231 );
buf ( w_19229 , \7720_b1 );
not ( w_19229 , w_19232 );
not (  , w_19233 );
and ( w_19232 , w_19233 , \7720_b0 );
or ( \7722_b1 , \7721_b1 , w_19234 );
xor ( \7722_b0 , \7721_b0 , w_19236 );
not ( w_19236 , w_19237 );
and ( w_19237 , w_19234 , w_19235 );
buf ( w_19234 , \7105_b1 );
not ( w_19234 , w_19238 );
not ( w_19235 , w_19239 );
and ( w_19238 , w_19239 , \7105_b0 );
or ( \7723_b1 , \5918_b1 , \7117_b1 );
not ( \7117_b1 , w_19240 );
and ( \7723_b0 , \5918_b0 , w_19241 );
and ( w_19240 , w_19241 , \7117_b0 );
or ( \7724_b1 , \5881_b1 , \7115_b1 );
not ( \7115_b1 , w_19242 );
and ( \7724_b0 , \5881_b0 , w_19243 );
and ( w_19242 , w_19243 , \7115_b0 );
or ( \7725_b1 , \7723_b1 , w_19245 );
not ( w_19245 , w_19246 );
and ( \7725_b0 , \7723_b0 , w_19247 );
and ( w_19246 ,  , w_19247 );
buf ( w_19245 , \7724_b1 );
not ( w_19245 , w_19248 );
not (  , w_19249 );
and ( w_19248 , w_19249 , \7724_b0 );
or ( \7726_b1 , \7725_b1 , w_19250 );
xor ( \7726_b0 , \7725_b0 , w_19252 );
not ( w_19252 , w_19253 );
and ( w_19253 , w_19250 , w_19251 );
buf ( w_19250 , \7123_b1 );
not ( w_19250 , w_19254 );
not ( w_19251 , w_19255 );
and ( w_19254 , w_19255 , \7123_b0 );
or ( \7727_b1 , \7722_b1 , \7726_b1 );
xor ( \7727_b0 , \7722_b0 , w_19256 );
not ( w_19256 , w_19257 );
and ( w_19257 , \7726_b1 , \7726_b0 );
or ( \7728_b1 , \5937_b1 , \7140_b1 );
not ( \7140_b1 , w_19258 );
and ( \7728_b0 , \5937_b0 , w_19259 );
and ( w_19258 , w_19259 , \7140_b0 );
or ( \7729_b1 , \5906_b1 , \7138_b1 );
not ( \7138_b1 , w_19260 );
and ( \7729_b0 , \5906_b0 , w_19261 );
and ( w_19260 , w_19261 , \7138_b0 );
or ( \7730_b1 , \7728_b1 , w_19263 );
not ( w_19263 , w_19264 );
and ( \7730_b0 , \7728_b0 , w_19265 );
and ( w_19264 ,  , w_19265 );
buf ( w_19263 , \7729_b1 );
not ( w_19263 , w_19266 );
not (  , w_19267 );
and ( w_19266 , w_19267 , \7729_b0 );
or ( \7731_b1 , \7730_b1 , w_19268 );
xor ( \7731_b0 , \7730_b0 , w_19270 );
not ( w_19270 , w_19271 );
and ( w_19271 , w_19268 , w_19269 );
buf ( w_19268 , \7146_b1 );
not ( w_19268 , w_19272 );
not ( w_19269 , w_19273 );
and ( w_19272 , w_19273 , \7146_b0 );
or ( \7732_b1 , \7727_b1 , \7731_b1 );
xor ( \7732_b0 , \7727_b0 , w_19274 );
not ( w_19274 , w_19275 );
and ( w_19275 , \7731_b1 , \7731_b0 );
or ( \7733_b1 , \7718_b1 , \7732_b1 );
xor ( \7733_b0 , \7718_b0 , w_19276 );
not ( w_19276 , w_19277 );
and ( w_19277 , \7732_b1 , \7732_b0 );
or ( \7734_b1 , \7556_b1 , \7560_b1 );
not ( \7560_b1 , w_19278 );
and ( \7734_b0 , \7556_b0 , w_19279 );
and ( w_19278 , w_19279 , \7560_b0 );
or ( \7735_b1 , \7560_b1 , \7565_b1 );
not ( \7565_b1 , w_19280 );
and ( \7735_b0 , \7560_b0 , w_19281 );
and ( w_19280 , w_19281 , \7565_b0 );
or ( \7736_b1 , \7556_b1 , \7565_b1 );
not ( \7565_b1 , w_19282 );
and ( \7736_b0 , \7556_b0 , w_19283 );
and ( w_19282 , w_19283 , \7565_b0 );
or ( \7738_b1 , \7541_b1 , \7545_b1 );
not ( \7545_b1 , w_19284 );
and ( \7738_b0 , \7541_b0 , w_19285 );
and ( w_19284 , w_19285 , \7545_b0 );
or ( \7739_b1 , \7545_b1 , \7550_b1 );
not ( \7550_b1 , w_19286 );
and ( \7739_b0 , \7545_b0 , w_19287 );
and ( w_19286 , w_19287 , \7550_b0 );
or ( \7740_b1 , \7541_b1 , \7550_b1 );
not ( \7550_b1 , w_19288 );
and ( \7740_b0 , \7541_b0 , w_19289 );
and ( w_19288 , w_19289 , \7550_b0 );
or ( \7742_b1 , \7737_b1 , \7741_b1 );
xor ( \7742_b0 , \7737_b0 , w_19290 );
not ( w_19290 , w_19291 );
and ( w_19291 , \7741_b1 , \7741_b0 );
or ( \7743_b1 , \6065_b1 , \5790_b1 );
not ( \5790_b1 , w_19292 );
and ( \7743_b0 , \6065_b0 , w_19293 );
and ( w_19292 , w_19293 , \5790_b0 );
or ( \7744_b1 , \6048_b1 , \5788_b1 );
not ( \5788_b1 , w_19294 );
and ( \7744_b0 , \6048_b0 , w_19295 );
and ( w_19294 , w_19295 , \5788_b0 );
or ( \7745_b1 , \7743_b1 , w_19297 );
not ( w_19297 , w_19298 );
and ( \7745_b0 , \7743_b0 , w_19299 );
and ( w_19298 ,  , w_19299 );
buf ( w_19297 , \7744_b1 );
not ( w_19297 , w_19300 );
not (  , w_19301 );
and ( w_19300 , w_19301 , \7744_b0 );
or ( \7746_b1 , \7745_b1 , w_19302 );
xor ( \7746_b0 , \7745_b0 , w_19304 );
not ( w_19304 , w_19305 );
and ( w_19305 , w_19302 , w_19303 );
buf ( w_19302 , \5797_b1 );
not ( w_19302 , w_19306 );
not ( w_19303 , w_19307 );
and ( w_19306 , w_19307 , \5797_b0 );
or ( \7747_b1 , \7742_b1 , \7746_b1 );
xor ( \7747_b0 , \7742_b0 , w_19308 );
not ( w_19308 , w_19309 );
and ( w_19309 , \7746_b1 , \7746_b0 );
or ( \7748_b1 , \7733_b1 , \7747_b1 );
xor ( \7748_b0 , \7733_b0 , w_19310 );
not ( w_19310 , w_19311 );
and ( w_19311 , \7747_b1 , \7747_b0 );
or ( \7749_b1 , \5797_b1 , \7528_b1 );
not ( \7528_b1 , w_19312 );
and ( \7749_b0 , \5797_b0 , w_19313 );
and ( w_19312 , w_19313 , \7528_b0 );
or ( \7750_b1 , \7528_b1 , \7533_b1 );
not ( \7533_b1 , w_19314 );
and ( \7750_b0 , \7528_b0 , w_19315 );
and ( w_19314 , w_19315 , \7533_b0 );
or ( \7751_b1 , \5797_b1 , \7533_b1 );
not ( \7533_b1 , w_19316 );
and ( \7751_b0 , \5797_b0 , w_19317 );
and ( w_19316 , w_19317 , \7533_b0 );
or ( \7753_b1 , \7513_b1 , \7517_b1 );
not ( \7517_b1 , w_19318 );
and ( \7753_b0 , \7513_b0 , w_19319 );
and ( w_19318 , w_19319 , \7517_b0 );
or ( \7754_b1 , \7517_b1 , \7522_b1 );
not ( \7522_b1 , w_19320 );
and ( \7754_b0 , \7517_b0 , w_19321 );
and ( w_19320 , w_19321 , \7522_b0 );
or ( \7755_b1 , \7513_b1 , \7522_b1 );
not ( \7522_b1 , w_19322 );
and ( \7755_b0 , \7513_b0 , w_19323 );
and ( w_19322 , w_19323 , \7522_b0 );
or ( \7757_b1 , \7752_b1 , \7756_b1 );
xor ( \7757_b0 , \7752_b0 , w_19324 );
not ( w_19324 , w_19325 );
and ( w_19325 , \7756_b1 , \7756_b0 );
or ( \7758_b1 , \7499_b1 , \7503_b1 );
not ( \7503_b1 , w_19326 );
and ( \7758_b0 , \7499_b0 , w_19327 );
and ( w_19326 , w_19327 , \7503_b0 );
or ( \7759_b1 , \7503_b1 , \7508_b1 );
not ( \7508_b1 , w_19328 );
and ( \7759_b0 , \7503_b0 , w_19329 );
and ( w_19328 , w_19329 , \7508_b0 );
or ( \7760_b1 , \7499_b1 , \7508_b1 );
not ( \7508_b1 , w_19330 );
and ( \7760_b0 , \7499_b0 , w_19331 );
and ( w_19330 , w_19331 , \7508_b0 );
or ( \7762_b1 , \7757_b1 , \7761_b1 );
xor ( \7762_b0 , \7757_b0 , w_19332 );
not ( w_19332 , w_19333 );
and ( w_19333 , \7761_b1 , \7761_b0 );
or ( \7763_b1 , \7748_b1 , \7762_b1 );
xor ( \7763_b0 , \7748_b0 , w_19334 );
not ( w_19334 , w_19335 );
and ( w_19335 , \7762_b1 , \7762_b0 );
or ( \7764_b1 , \7689_b1 , \7763_b1 );
xor ( \7764_b0 , \7689_b0 , w_19336 );
not ( w_19336 , w_19337 );
and ( w_19337 , \7763_b1 , \7763_b0 );
or ( \7765_b1 , \7680_b1 , \7764_b1 );
xor ( \7765_b0 , \7680_b0 , w_19338 );
not ( w_19338 , w_19339 );
and ( w_19339 , \7764_b1 , \7764_b0 );
or ( \7766_b1 , \7626_b1 , \7765_b1 );
xor ( \7766_b0 , \7626_b0 , w_19340 );
not ( w_19340 , w_19341 );
and ( w_19341 , \7765_b1 , \7765_b0 );
or ( \7767_b1 , \5831_b1 , \6991_b1 );
not ( \6991_b1 , w_19342 );
and ( \7767_b0 , \5831_b0 , w_19343 );
and ( w_19342 , w_19343 , \6991_b0 );
or ( \7768_b1 , \5799_b1 , \6988_b1 );
not ( \6988_b1 , w_19344 );
and ( \7768_b0 , \5799_b0 , w_19345 );
and ( w_19344 , w_19345 , \6988_b0 );
or ( \7769_b1 , \7767_b1 , w_19347 );
not ( w_19347 , w_19348 );
and ( \7769_b0 , \7767_b0 , w_19349 );
and ( w_19348 ,  , w_19349 );
buf ( w_19347 , \7768_b1 );
not ( w_19347 , w_19350 );
not (  , w_19351 );
and ( w_19350 , w_19351 , \7768_b0 );
or ( \7770_b1 , \7769_b1 , w_19352 );
xor ( \7770_b0 , \7769_b0 , w_19354 );
not ( w_19354 , w_19355 );
and ( w_19355 , w_19352 , w_19353 );
buf ( w_19352 , \6985_b1 );
not ( w_19352 , w_19356 );
not ( w_19353 , w_19357 );
and ( w_19356 , w_19357 , \6985_b0 );
or ( \7771_b1 , \5854_b1 , \7006_b1 );
not ( \7006_b1 , w_19358 );
and ( \7771_b0 , \5854_b0 , w_19359 );
and ( w_19358 , w_19359 , \7006_b0 );
or ( \7772_b1 , \5819_b1 , \7004_b1 );
not ( \7004_b1 , w_19360 );
and ( \7772_b0 , \5819_b0 , w_19361 );
and ( w_19360 , w_19361 , \7004_b0 );
or ( \7773_b1 , \7771_b1 , w_19363 );
not ( w_19363 , w_19364 );
and ( \7773_b0 , \7771_b0 , w_19365 );
and ( w_19364 ,  , w_19365 );
buf ( w_19363 , \7772_b1 );
not ( w_19363 , w_19366 );
not (  , w_19367 );
and ( w_19366 , w_19367 , \7772_b0 );
or ( \7774_b1 , \7773_b1 , w_19368 );
xor ( \7774_b0 , \7773_b0 , w_19370 );
not ( w_19370 , w_19371 );
and ( w_19371 , w_19368 , w_19369 );
buf ( w_19368 , \7012_b1 );
not ( w_19368 , w_19372 );
not ( w_19369 , w_19373 );
and ( w_19372 , w_19373 , \7012_b0 );
or ( \7775_b1 , \7770_b1 , \7774_b1 );
not ( \7774_b1 , w_19374 );
and ( \7775_b0 , \7770_b0 , w_19375 );
and ( w_19374 , w_19375 , \7774_b0 );
or ( \7776_b1 , \5873_b1 , \7026_b1 );
not ( \7026_b1 , w_19376 );
and ( \7776_b0 , \5873_b0 , w_19377 );
and ( w_19376 , w_19377 , \7026_b0 );
or ( \7777_b1 , \5842_b1 , \7024_b1 );
not ( \7024_b1 , w_19378 );
and ( \7777_b0 , \5842_b0 , w_19379 );
and ( w_19378 , w_19379 , \7024_b0 );
or ( \7778_b1 , \7776_b1 , w_19381 );
not ( w_19381 , w_19382 );
and ( \7778_b0 , \7776_b0 , w_19383 );
and ( w_19382 ,  , w_19383 );
buf ( w_19381 , \7777_b1 );
not ( w_19381 , w_19384 );
not (  , w_19385 );
and ( w_19384 , w_19385 , \7777_b0 );
or ( \7779_b1 , \7778_b1 , w_19386 );
xor ( \7779_b0 , \7778_b0 , w_19388 );
not ( w_19388 , w_19389 );
and ( w_19389 , w_19386 , w_19387 );
buf ( w_19386 , \7032_b1 );
not ( w_19386 , w_19390 );
not ( w_19387 , w_19391 );
and ( w_19390 , w_19391 , \7032_b0 );
or ( \7780_b1 , \7774_b1 , \7779_b1 );
not ( \7779_b1 , w_19392 );
and ( \7780_b0 , \7774_b0 , w_19393 );
and ( w_19392 , w_19393 , \7779_b0 );
or ( \7781_b1 , \7770_b1 , \7779_b1 );
not ( \7779_b1 , w_19394 );
and ( \7781_b0 , \7770_b0 , w_19395 );
and ( w_19394 , w_19395 , \7779_b0 );
or ( \7783_b1 , \5893_b1 , \7043_b1 );
not ( \7043_b1 , w_19396 );
and ( \7783_b0 , \5893_b0 , w_19397 );
and ( w_19396 , w_19397 , \7043_b0 );
or ( \7784_b1 , \5861_b1 , \7041_b1 );
not ( \7041_b1 , w_19398 );
and ( \7784_b0 , \5861_b0 , w_19399 );
and ( w_19398 , w_19399 , \7041_b0 );
or ( \7785_b1 , \7783_b1 , w_19401 );
not ( w_19401 , w_19402 );
and ( \7785_b0 , \7783_b0 , w_19403 );
and ( w_19402 ,  , w_19403 );
buf ( w_19401 , \7784_b1 );
not ( w_19401 , w_19404 );
not (  , w_19405 );
and ( w_19404 , w_19405 , \7784_b0 );
or ( \7786_b1 , \7785_b1 , w_19406 );
xor ( \7786_b0 , \7785_b0 , w_19408 );
not ( w_19408 , w_19409 );
and ( w_19409 , w_19406 , w_19407 );
buf ( w_19406 , \7049_b1 );
not ( w_19406 , w_19410 );
not ( w_19407 , w_19411 );
and ( w_19410 , w_19411 , \7049_b0 );
or ( \7787_b1 , \5918_b1 , \7061_b1 );
not ( \7061_b1 , w_19412 );
and ( \7787_b0 , \5918_b0 , w_19413 );
and ( w_19412 , w_19413 , \7061_b0 );
or ( \7788_b1 , \5881_b1 , \7059_b1 );
not ( \7059_b1 , w_19414 );
and ( \7788_b0 , \5881_b0 , w_19415 );
and ( w_19414 , w_19415 , \7059_b0 );
or ( \7789_b1 , \7787_b1 , w_19417 );
not ( w_19417 , w_19418 );
and ( \7789_b0 , \7787_b0 , w_19419 );
and ( w_19418 ,  , w_19419 );
buf ( w_19417 , \7788_b1 );
not ( w_19417 , w_19420 );
not (  , w_19421 );
and ( w_19420 , w_19421 , \7788_b0 );
or ( \7790_b1 , \7789_b1 , w_19422 );
xor ( \7790_b0 , \7789_b0 , w_19424 );
not ( w_19424 , w_19425 );
and ( w_19425 , w_19422 , w_19423 );
buf ( w_19422 , \7067_b1 );
not ( w_19422 , w_19426 );
not ( w_19423 , w_19427 );
and ( w_19426 , w_19427 , \7067_b0 );
or ( \7791_b1 , \7786_b1 , \7790_b1 );
not ( \7790_b1 , w_19428 );
and ( \7791_b0 , \7786_b0 , w_19429 );
and ( w_19428 , w_19429 , \7790_b0 );
or ( \7792_b1 , \5937_b1 , \7082_b1 );
not ( \7082_b1 , w_19430 );
and ( \7792_b0 , \5937_b0 , w_19431 );
and ( w_19430 , w_19431 , \7082_b0 );
or ( \7793_b1 , \5906_b1 , \7080_b1 );
not ( \7080_b1 , w_19432 );
and ( \7793_b0 , \5906_b0 , w_19433 );
and ( w_19432 , w_19433 , \7080_b0 );
or ( \7794_b1 , \7792_b1 , w_19435 );
not ( w_19435 , w_19436 );
and ( \7794_b0 , \7792_b0 , w_19437 );
and ( w_19436 ,  , w_19437 );
buf ( w_19435 , \7793_b1 );
not ( w_19435 , w_19438 );
not (  , w_19439 );
and ( w_19438 , w_19439 , \7793_b0 );
or ( \7795_b1 , \7794_b1 , w_19440 );
xor ( \7795_b0 , \7794_b0 , w_19442 );
not ( w_19442 , w_19443 );
and ( w_19443 , w_19440 , w_19441 );
buf ( w_19440 , \7088_b1 );
not ( w_19440 , w_19444 );
not ( w_19441 , w_19445 );
and ( w_19444 , w_19445 , \7088_b0 );
or ( \7796_b1 , \7790_b1 , \7795_b1 );
not ( \7795_b1 , w_19446 );
and ( \7796_b0 , \7790_b0 , w_19447 );
and ( w_19446 , w_19447 , \7795_b0 );
or ( \7797_b1 , \7786_b1 , \7795_b1 );
not ( \7795_b1 , w_19448 );
and ( \7797_b0 , \7786_b0 , w_19449 );
and ( w_19448 , w_19449 , \7795_b0 );
or ( \7799_b1 , \7782_b1 , \7798_b1 );
not ( \7798_b1 , w_19450 );
and ( \7799_b0 , \7782_b0 , w_19451 );
and ( w_19450 , w_19451 , \7798_b0 );
or ( \7800_b1 , \5957_b1 , \7099_b1 );
not ( \7099_b1 , w_19452 );
and ( \7800_b0 , \5957_b0 , w_19453 );
and ( w_19452 , w_19453 , \7099_b0 );
or ( \7801_b1 , \5925_b1 , \7097_b1 );
not ( \7097_b1 , w_19454 );
and ( \7801_b0 , \5925_b0 , w_19455 );
and ( w_19454 , w_19455 , \7097_b0 );
or ( \7802_b1 , \7800_b1 , w_19457 );
not ( w_19457 , w_19458 );
and ( \7802_b0 , \7800_b0 , w_19459 );
and ( w_19458 ,  , w_19459 );
buf ( w_19457 , \7801_b1 );
not ( w_19457 , w_19460 );
not (  , w_19461 );
and ( w_19460 , w_19461 , \7801_b0 );
or ( \7803_b1 , \7802_b1 , w_19462 );
xor ( \7803_b0 , \7802_b0 , w_19464 );
not ( w_19464 , w_19465 );
and ( w_19465 , w_19462 , w_19463 );
buf ( w_19462 , \7105_b1 );
not ( w_19462 , w_19466 );
not ( w_19463 , w_19467 );
and ( w_19466 , w_19467 , \7105_b0 );
or ( \7804_b1 , \5979_b1 , \7117_b1 );
not ( \7117_b1 , w_19468 );
and ( \7804_b0 , \5979_b0 , w_19469 );
and ( w_19468 , w_19469 , \7117_b0 );
or ( \7805_b1 , \5945_b1 , \7115_b1 );
not ( \7115_b1 , w_19470 );
and ( \7805_b0 , \5945_b0 , w_19471 );
and ( w_19470 , w_19471 , \7115_b0 );
or ( \7806_b1 , \7804_b1 , w_19473 );
not ( w_19473 , w_19474 );
and ( \7806_b0 , \7804_b0 , w_19475 );
and ( w_19474 ,  , w_19475 );
buf ( w_19473 , \7805_b1 );
not ( w_19473 , w_19476 );
not (  , w_19477 );
and ( w_19476 , w_19477 , \7805_b0 );
or ( \7807_b1 , \7806_b1 , w_19478 );
xor ( \7807_b0 , \7806_b0 , w_19480 );
not ( w_19480 , w_19481 );
and ( w_19481 , w_19478 , w_19479 );
buf ( w_19478 , \7123_b1 );
not ( w_19478 , w_19482 );
not ( w_19479 , w_19483 );
and ( w_19482 , w_19483 , \7123_b0 );
or ( \7808_b1 , \7803_b1 , \7807_b1 );
not ( \7807_b1 , w_19484 );
and ( \7808_b0 , \7803_b0 , w_19485 );
and ( w_19484 , w_19485 , \7807_b0 );
or ( \7809_b1 , \5998_b1 , \7140_b1 );
not ( \7140_b1 , w_19486 );
and ( \7809_b0 , \5998_b0 , w_19487 );
and ( w_19486 , w_19487 , \7140_b0 );
or ( \7810_b1 , \5967_b1 , \7138_b1 );
not ( \7138_b1 , w_19488 );
and ( \7810_b0 , \5967_b0 , w_19489 );
and ( w_19488 , w_19489 , \7138_b0 );
or ( \7811_b1 , \7809_b1 , w_19491 );
not ( w_19491 , w_19492 );
and ( \7811_b0 , \7809_b0 , w_19493 );
and ( w_19492 ,  , w_19493 );
buf ( w_19491 , \7810_b1 );
not ( w_19491 , w_19494 );
not (  , w_19495 );
and ( w_19494 , w_19495 , \7810_b0 );
or ( \7812_b1 , \7811_b1 , w_19496 );
xor ( \7812_b0 , \7811_b0 , w_19498 );
not ( w_19498 , w_19499 );
and ( w_19499 , w_19496 , w_19497 );
buf ( w_19496 , \7146_b1 );
not ( w_19496 , w_19500 );
not ( w_19497 , w_19501 );
and ( w_19500 , w_19501 , \7146_b0 );
or ( \7813_b1 , \7807_b1 , \7812_b1 );
not ( \7812_b1 , w_19502 );
and ( \7813_b0 , \7807_b0 , w_19503 );
and ( w_19502 , w_19503 , \7812_b0 );
or ( \7814_b1 , \7803_b1 , \7812_b1 );
not ( \7812_b1 , w_19504 );
and ( \7814_b0 , \7803_b0 , w_19505 );
and ( w_19504 , w_19505 , \7812_b0 );
or ( \7816_b1 , \7798_b1 , \7815_b1 );
not ( \7815_b1 , w_19506 );
and ( \7816_b0 , \7798_b0 , w_19507 );
and ( w_19506 , w_19507 , \7815_b0 );
or ( \7817_b1 , \7782_b1 , \7815_b1 );
not ( \7815_b1 , w_19508 );
and ( \7817_b0 , \7782_b0 , w_19509 );
and ( w_19508 , w_19509 , \7815_b0 );
or ( \7819_b1 , \6018_b1 , \7157_b1 );
not ( \7157_b1 , w_19510 );
and ( \7819_b0 , \6018_b0 , w_19511 );
and ( w_19510 , w_19511 , \7157_b0 );
or ( \7820_b1 , \5986_b1 , \7155_b1 );
not ( \7155_b1 , w_19512 );
and ( \7820_b0 , \5986_b0 , w_19513 );
and ( w_19512 , w_19513 , \7155_b0 );
or ( \7821_b1 , \7819_b1 , w_19515 );
not ( w_19515 , w_19516 );
and ( \7821_b0 , \7819_b0 , w_19517 );
and ( w_19516 ,  , w_19517 );
buf ( w_19515 , \7820_b1 );
not ( w_19515 , w_19518 );
not (  , w_19519 );
and ( w_19518 , w_19519 , \7820_b0 );
or ( \7822_b1 , \7821_b1 , w_19520 );
xor ( \7822_b0 , \7821_b0 , w_19522 );
not ( w_19522 , w_19523 );
and ( w_19523 , w_19520 , w_19521 );
buf ( w_19520 , \7163_b1 );
not ( w_19520 , w_19524 );
not ( w_19521 , w_19525 );
and ( w_19524 , w_19525 , \7163_b0 );
or ( \7823_b1 , \6041_b1 , \7175_b1 );
not ( \7175_b1 , w_19526 );
and ( \7823_b0 , \6041_b0 , w_19527 );
and ( w_19526 , w_19527 , \7175_b0 );
or ( \7824_b1 , \6006_b1 , \7173_b1 );
not ( \7173_b1 , w_19528 );
and ( \7824_b0 , \6006_b0 , w_19529 );
and ( w_19528 , w_19529 , \7173_b0 );
or ( \7825_b1 , \7823_b1 , w_19531 );
not ( w_19531 , w_19532 );
and ( \7825_b0 , \7823_b0 , w_19533 );
and ( w_19532 ,  , w_19533 );
buf ( w_19531 , \7824_b1 );
not ( w_19531 , w_19534 );
not (  , w_19535 );
and ( w_19534 , w_19535 , \7824_b0 );
or ( \7826_b1 , \7825_b1 , w_19536 );
xor ( \7826_b0 , \7825_b0 , w_19538 );
not ( w_19538 , w_19539 );
and ( w_19539 , w_19536 , w_19537 );
buf ( w_19536 , \7181_b1 );
not ( w_19536 , w_19540 );
not ( w_19537 , w_19541 );
and ( w_19540 , w_19541 , \7181_b0 );
or ( \7827_b1 , \7822_b1 , \7826_b1 );
not ( \7826_b1 , w_19542 );
and ( \7827_b0 , \7822_b0 , w_19543 );
and ( w_19542 , w_19543 , \7826_b0 );
or ( \7828_b1 , \6057_b1 , \7192_b1 );
not ( \7192_b1 , w_19544 );
and ( \7828_b0 , \6057_b0 , w_19545 );
and ( w_19544 , w_19545 , \7192_b0 );
or ( \7829_b1 , \6029_b1 , \7190_b1 );
not ( \7190_b1 , w_19546 );
and ( \7829_b0 , \6029_b0 , w_19547 );
and ( w_19546 , w_19547 , \7190_b0 );
or ( \7830_b1 , \7828_b1 , w_19549 );
not ( w_19549 , w_19550 );
and ( \7830_b0 , \7828_b0 , w_19551 );
and ( w_19550 ,  , w_19551 );
buf ( w_19549 , \7829_b1 );
not ( w_19549 , w_19552 );
not (  , w_19553 );
and ( w_19552 , w_19553 , \7829_b0 );
or ( \7831_b1 , \7830_b1 , w_19554 );
xor ( \7831_b0 , \7830_b0 , w_19556 );
not ( w_19556 , w_19557 );
and ( w_19557 , w_19554 , w_19555 );
buf ( w_19554 , \7198_b1 );
not ( w_19554 , w_19558 );
not ( w_19555 , w_19559 );
and ( w_19558 , w_19559 , \7198_b0 );
or ( \7832_b1 , \7826_b1 , \7831_b1 );
not ( \7831_b1 , w_19560 );
and ( \7832_b0 , \7826_b0 , w_19561 );
and ( w_19560 , w_19561 , \7831_b0 );
or ( \7833_b1 , \7822_b1 , \7831_b1 );
not ( \7831_b1 , w_19562 );
and ( \7833_b0 , \7822_b0 , w_19563 );
and ( w_19562 , w_19563 , \7831_b0 );
or ( \7835_b1 , \7199_b1 , \7207_b1 );
xor ( \7835_b0 , \7199_b0 , w_19564 );
not ( w_19564 , w_19565 );
and ( w_19565 , \7207_b1 , \7207_b0 );
or ( \7836_b1 , \7835_b1 , \7210_b1 );
xor ( \7836_b0 , \7835_b0 , w_19566 );
not ( w_19566 , w_19567 );
and ( w_19567 , \7210_b1 , \7210_b0 );
or ( \7837_b1 , \7834_b1 , \7836_b1 );
not ( \7836_b1 , w_19568 );
and ( \7837_b0 , \7834_b0 , w_19569 );
and ( w_19568 , w_19569 , \7836_b0 );
or ( \7838_b1 , \7147_b1 , \7164_b1 );
xor ( \7838_b0 , \7147_b0 , w_19570 );
not ( w_19570 , w_19571 );
and ( w_19571 , \7164_b1 , \7164_b0 );
or ( \7839_b1 , \7838_b1 , \7182_b1 );
xor ( \7839_b0 , \7838_b0 , w_19572 );
not ( w_19572 , w_19573 );
and ( w_19573 , \7182_b1 , \7182_b0 );
or ( \7840_b1 , \7836_b1 , \7839_b1 );
not ( \7839_b1 , w_19574 );
and ( \7840_b0 , \7836_b0 , w_19575 );
and ( w_19574 , w_19575 , \7839_b0 );
or ( \7841_b1 , \7834_b1 , \7839_b1 );
not ( \7839_b1 , w_19576 );
and ( \7841_b0 , \7834_b0 , w_19577 );
and ( w_19576 , w_19577 , \7839_b0 );
or ( \7843_b1 , \7818_b1 , \7842_b1 );
not ( \7842_b1 , w_19578 );
and ( \7843_b0 , \7818_b0 , w_19579 );
and ( w_19578 , w_19579 , \7842_b0 );
or ( \7844_b1 , \7089_b1 , \7106_b1 );
xor ( \7844_b0 , \7089_b0 , w_19580 );
not ( w_19580 , w_19581 );
and ( w_19581 , \7106_b1 , \7106_b0 );
or ( \7845_b1 , \7844_b1 , \7124_b1 );
xor ( \7845_b0 , \7844_b0 , w_19582 );
not ( w_19582 , w_19583 );
and ( w_19583 , \7124_b1 , \7124_b0 );
or ( \7846_b1 , \7033_b1 , \7050_b1 );
xor ( \7846_b0 , \7033_b0 , w_19584 );
not ( w_19584 , w_19585 );
and ( w_19585 , \7050_b1 , \7050_b0 );
or ( \7847_b1 , \7846_b1 , \7068_b1 );
xor ( \7847_b0 , \7846_b0 , w_19586 );
not ( w_19586 , w_19587 );
and ( w_19587 , \7068_b1 , \7068_b0 );
or ( \7848_b1 , \7845_b1 , \7847_b1 );
not ( \7847_b1 , w_19588 );
and ( \7848_b0 , \7845_b0 , w_19589 );
and ( w_19588 , w_19589 , \7847_b0 );
or ( \7849_b1 , \5755_b1 , \6995_b1 );
xor ( \7849_b0 , \5755_b0 , w_19590 );
not ( w_19590 , w_19591 );
and ( w_19591 , \6995_b1 , \6995_b0 );
or ( \7850_b1 , \7849_b1 , \7013_b1 );
xor ( \7850_b0 , \7849_b0 , w_19592 );
not ( w_19592 , w_19593 );
and ( w_19593 , \7013_b1 , \7013_b0 );
or ( \7851_b1 , \7847_b1 , \7850_b1 );
not ( \7850_b1 , w_19594 );
and ( \7851_b0 , \7847_b0 , w_19595 );
and ( w_19594 , w_19595 , \7850_b0 );
or ( \7852_b1 , \7845_b1 , \7850_b1 );
not ( \7850_b1 , w_19596 );
and ( \7852_b0 , \7845_b0 , w_19597 );
and ( w_19596 , w_19597 , \7850_b0 );
or ( \7854_b1 , \7842_b1 , \7853_b1 );
not ( \7853_b1 , w_19598 );
and ( \7854_b0 , \7842_b0 , w_19599 );
and ( w_19598 , w_19599 , \7853_b0 );
or ( \7855_b1 , \7818_b1 , \7853_b1 );
not ( \7853_b1 , w_19600 );
and ( \7855_b0 , \7818_b0 , w_19601 );
and ( w_19600 , w_19601 , \7853_b0 );
or ( \7857_b1 , \7463_b1 , \7467_b1 );
xor ( \7857_b0 , \7463_b0 , w_19602 );
not ( w_19602 , w_19603 );
and ( w_19603 , \7467_b1 , \7467_b0 );
or ( \7858_b1 , \7857_b1 , \7472_b1 );
xor ( \7858_b0 , \7857_b0 , w_19604 );
not ( w_19604 , w_19605 );
and ( w_19605 , \7472_b1 , \7472_b0 );
or ( \7859_b1 , \7447_b1 , \7451_b1 );
xor ( \7859_b0 , \7447_b0 , w_19606 );
not ( w_19606 , w_19607 );
and ( w_19607 , \7451_b1 , \7451_b0 );
or ( \7860_b1 , \7859_b1 , \7456_b1 );
xor ( \7860_b0 , \7859_b0 , w_19608 );
not ( w_19608 , w_19609 );
and ( w_19609 , \7456_b1 , \7456_b0 );
or ( \7861_b1 , \7858_b1 , \7860_b1 );
not ( \7860_b1 , w_19610 );
and ( \7861_b0 , \7858_b0 , w_19611 );
and ( w_19610 , w_19611 , \7860_b0 );
or ( \7862_b1 , \7226_b1 , \7240_b1 );
xor ( \7862_b0 , \7226_b0 , w_19612 );
not ( w_19612 , w_19613 );
and ( w_19613 , \7240_b1 , \7240_b0 );
or ( \7863_b1 , \7862_b1 , \7255_b1 );
xor ( \7863_b0 , \7862_b0 , w_19614 );
not ( w_19614 , w_19615 );
and ( w_19615 , \7255_b1 , \7255_b0 );
or ( \7864_b1 , \7860_b1 , \7863_b1 );
not ( \7863_b1 , w_19616 );
and ( \7864_b0 , \7860_b0 , w_19617 );
and ( w_19616 , w_19617 , \7863_b0 );
or ( \7865_b1 , \7858_b1 , \7863_b1 );
not ( \7863_b1 , w_19618 );
and ( \7865_b0 , \7858_b0 , w_19619 );
and ( w_19618 , w_19619 , \7863_b0 );
or ( \7867_b1 , \7856_b1 , \7866_b1 );
not ( \7866_b1 , w_19620 );
and ( \7867_b0 , \7856_b0 , w_19621 );
and ( w_19620 , w_19621 , \7866_b0 );
or ( \7868_b1 , \7459_b1 , \7475_b1 );
xor ( \7868_b0 , \7459_b0 , w_19622 );
not ( w_19622 , w_19623 );
and ( w_19623 , \7475_b1 , \7475_b0 );
or ( \7869_b1 , \7868_b1 , \7480_b1 );
xor ( \7869_b0 , \7868_b0 , w_19624 );
not ( w_19624 , w_19625 );
and ( w_19625 , \7480_b1 , \7480_b0 );
or ( \7870_b1 , \7866_b1 , \7869_b1 );
not ( \7869_b1 , w_19626 );
and ( \7870_b0 , \7866_b0 , w_19627 );
and ( w_19626 , w_19627 , \7869_b0 );
or ( \7871_b1 , \7856_b1 , \7869_b1 );
not ( \7869_b1 , w_19628 );
and ( \7871_b0 , \7856_b0 , w_19629 );
and ( w_19628 , w_19629 , \7869_b0 );
or ( \7873_b1 , \7443_b1 , \7493_b1 );
xor ( \7873_b0 , \7443_b0 , w_19630 );
not ( w_19630 , w_19631 );
and ( w_19631 , \7493_b1 , \7493_b0 );
or ( \7874_b1 , \7872_b1 , \7873_b1 );
not ( \7873_b1 , w_19632 );
and ( \7874_b0 , \7872_b0 , w_19633 );
and ( w_19632 , w_19633 , \7873_b0 );
or ( \7875_b1 , \7261_b1 , \7341_b1 );
xor ( \7875_b0 , \7261_b0 , w_19634 );
not ( w_19634 , w_19635 );
and ( w_19635 , \7341_b1 , \7341_b0 );
or ( \7876_b1 , \7875_b1 , \7356_b1 );
xor ( \7876_b0 , \7875_b0 , w_19636 );
not ( w_19636 , w_19637 );
and ( w_19637 , \7356_b1 , \7356_b0 );
or ( \7877_b1 , \7873_b1 , \7876_b1 );
not ( \7876_b1 , w_19638 );
and ( \7877_b0 , \7873_b0 , w_19639 );
and ( w_19638 , w_19639 , \7876_b0 );
or ( \7878_b1 , \7872_b1 , \7876_b1 );
not ( \7876_b1 , w_19640 );
and ( \7878_b0 , \7872_b0 , w_19641 );
and ( w_19640 , w_19641 , \7876_b0 );
or ( \7880_b1 , \7600_b1 , \7624_b1 );
xor ( \7880_b0 , \7600_b0 , w_19642 );
not ( w_19642 , w_19643 );
and ( w_19643 , \7624_b1 , \7624_b0 );
or ( \7881_b1 , \7879_b1 , \7880_b1 );
not ( \7880_b1 , w_19644 );
and ( \7881_b0 , \7879_b0 , w_19645 );
and ( w_19644 , w_19645 , \7880_b0 );
or ( \7882_b1 , \7359_b1 , \7494_b1 );
xor ( \7882_b0 , \7359_b0 , w_19646 );
not ( w_19646 , w_19647 );
and ( w_19647 , \7494_b1 , \7494_b0 );
or ( \7883_b1 , \7882_b1 , \7583_b1 );
xor ( \7883_b0 , \7882_b0 , w_19648 );
not ( w_19648 , w_19649 );
and ( w_19649 , \7583_b1 , \7583_b0 );
or ( \7884_b1 , \7880_b1 , \7883_b1 );
not ( \7883_b1 , w_19650 );
and ( \7884_b0 , \7880_b0 , w_19651 );
and ( w_19650 , w_19651 , \7883_b0 );
or ( \7885_b1 , \7879_b1 , \7883_b1 );
not ( \7883_b1 , w_19652 );
and ( \7885_b0 , \7879_b0 , w_19653 );
and ( w_19652 , w_19653 , \7883_b0 );
or ( \7887_b1 , \7766_b1 , w_19655 );
not ( w_19655 , w_19656 );
and ( \7887_b0 , \7766_b0 , w_19657 );
and ( w_19656 ,  , w_19657 );
buf ( w_19655 , \7886_b1 );
not ( w_19655 , w_19658 );
not (  , w_19659 );
and ( w_19658 , w_19659 , \7886_b0 );
or ( \7888_b1 , \7630_b1 , \7679_b1 );
not ( \7679_b1 , w_19660 );
and ( \7888_b0 , \7630_b0 , w_19661 );
and ( w_19660 , w_19661 , \7679_b0 );
or ( \7889_b1 , \7679_b1 , \7764_b1 );
not ( \7764_b1 , w_19662 );
and ( \7889_b0 , \7679_b0 , w_19663 );
and ( w_19662 , w_19663 , \7764_b0 );
or ( \7890_b1 , \7630_b1 , \7764_b1 );
not ( \7764_b1 , w_19664 );
and ( \7890_b0 , \7630_b0 , w_19665 );
and ( w_19664 , w_19665 , \7764_b0 );
or ( \7892_b1 , \7668_b1 , \7672_b1 );
not ( \7672_b1 , w_19666 );
and ( \7892_b0 , \7668_b0 , w_19667 );
and ( w_19666 , w_19667 , \7672_b0 );
or ( \7893_b1 , \7672_b1 , \7677_b1 );
not ( \7677_b1 , w_19668 );
and ( \7893_b0 , \7672_b0 , w_19669 );
and ( w_19668 , w_19669 , \7677_b0 );
or ( \7894_b1 , \7668_b1 , \7677_b1 );
not ( \7677_b1 , w_19670 );
and ( \7894_b0 , \7668_b0 , w_19671 );
and ( w_19670 , w_19671 , \7677_b0 );
or ( \7896_b1 , \7634_b1 , \7648_b1 );
not ( \7648_b1 , w_19672 );
and ( \7896_b0 , \7634_b0 , w_19673 );
and ( w_19672 , w_19673 , \7648_b0 );
or ( \7897_b1 , \7648_b1 , \7663_b1 );
not ( \7663_b1 , w_19674 );
and ( \7897_b0 , \7648_b0 , w_19675 );
and ( w_19674 , w_19675 , \7663_b0 );
or ( \7898_b1 , \7634_b1 , \7663_b1 );
not ( \7663_b1 , w_19676 );
and ( \7898_b0 , \7634_b0 , w_19677 );
and ( w_19676 , w_19677 , \7663_b0 );
or ( \7900_b1 , \7895_b1 , \7899_b1 );
xor ( \7900_b0 , \7895_b0 , w_19678 );
not ( w_19678 , w_19679 );
and ( w_19679 , \7899_b1 , \7899_b0 );
or ( \7901_b1 , \7733_b1 , \7747_b1 );
not ( \7747_b1 , w_19680 );
and ( \7901_b0 , \7733_b0 , w_19681 );
and ( w_19680 , w_19681 , \7747_b0 );
or ( \7902_b1 , \7747_b1 , \7762_b1 );
not ( \7762_b1 , w_19682 );
and ( \7902_b0 , \7747_b0 , w_19683 );
and ( w_19682 , w_19683 , \7762_b0 );
or ( \7903_b1 , \7733_b1 , \7762_b1 );
not ( \7762_b1 , w_19684 );
and ( \7903_b0 , \7733_b0 , w_19685 );
and ( w_19684 , w_19685 , \7762_b0 );
or ( \7905_b1 , \7900_b1 , \7904_b1 );
xor ( \7905_b0 , \7900_b0 , w_19686 );
not ( w_19686 , w_19687 );
and ( w_19687 , \7904_b1 , \7904_b0 );
or ( \7906_b1 , \7891_b1 , \7905_b1 );
xor ( \7906_b0 , \7891_b0 , w_19688 );
not ( w_19688 , w_19689 );
and ( w_19689 , \7905_b1 , \7905_b0 );
or ( \7907_b1 , \7684_b1 , \7688_b1 );
not ( \7688_b1 , w_19690 );
and ( \7907_b0 , \7684_b0 , w_19691 );
and ( w_19690 , w_19691 , \7688_b0 );
or ( \7908_b1 , \7688_b1 , \7763_b1 );
not ( \7763_b1 , w_19692 );
and ( \7908_b0 , \7688_b0 , w_19693 );
and ( w_19692 , w_19693 , \7763_b0 );
or ( \7909_b1 , \7684_b1 , \7763_b1 );
not ( \7763_b1 , w_19694 );
and ( \7909_b0 , \7684_b0 , w_19695 );
and ( w_19694 , w_19695 , \7763_b0 );
or ( \7911_b1 , \7664_b1 , \7678_b1 );
not ( \7678_b1 , w_19696 );
and ( \7911_b0 , \7664_b0 , w_19697 );
and ( w_19696 , w_19697 , \7678_b0 );
or ( \7912_b1 , \7910_b1 , \7911_b1 );
xor ( \7912_b0 , \7910_b0 , w_19698 );
not ( w_19698 , w_19699 );
and ( w_19699 , \7911_b1 , \7911_b0 );
or ( \7913_b1 , \7707_b1 , \7711_b1 );
not ( \7711_b1 , w_19700 );
and ( \7913_b0 , \7707_b0 , w_19701 );
and ( w_19700 , w_19701 , \7711_b0 );
or ( \7914_b1 , \7711_b1 , \7716_b1 );
not ( \7716_b1 , w_19702 );
and ( \7914_b0 , \7711_b0 , w_19703 );
and ( w_19702 , w_19703 , \7716_b0 );
or ( \7915_b1 , \7707_b1 , \7716_b1 );
not ( \7716_b1 , w_19704 );
and ( \7915_b0 , \7707_b0 , w_19705 );
and ( w_19704 , w_19705 , \7716_b0 );
or ( \7917_b1 , \7693_b1 , \7697_b1 );
not ( \7697_b1 , w_19706 );
and ( \7917_b0 , \7693_b0 , w_19707 );
and ( w_19706 , w_19707 , \7697_b0 );
or ( \7918_b1 , \7697_b1 , \7702_b1 );
not ( \7702_b1 , w_19708 );
and ( \7918_b0 , \7697_b0 , w_19709 );
and ( w_19708 , w_19709 , \7702_b0 );
or ( \7919_b1 , \7693_b1 , \7702_b1 );
not ( \7702_b1 , w_19710 );
and ( \7919_b0 , \7693_b0 , w_19711 );
and ( w_19710 , w_19711 , \7702_b0 );
or ( \7921_b1 , \7916_b1 , \7920_b1 );
xor ( \7921_b0 , \7916_b0 , w_19712 );
not ( w_19712 , w_19713 );
and ( w_19713 , \7920_b1 , \7920_b0 );
or ( \7922_b1 , \6029_b1 , \5768_b1 );
not ( \5768_b1 , w_19714 );
and ( \7922_b0 , \6029_b0 , w_19715 );
and ( w_19714 , w_19715 , \5768_b0 );
or ( \7923_b1 , \6041_b1 , \5766_b1 );
not ( \5766_b1 , w_19716 );
and ( \7923_b0 , \6041_b0 , w_19717 );
and ( w_19716 , w_19717 , \5766_b0 );
or ( \7924_b1 , \7922_b1 , w_19719 );
not ( w_19719 , w_19720 );
and ( \7924_b0 , \7922_b0 , w_19721 );
and ( w_19720 ,  , w_19721 );
buf ( w_19719 , \7923_b1 );
not ( w_19719 , w_19722 );
not (  , w_19723 );
and ( w_19722 , w_19723 , \7923_b0 );
or ( \7925_b1 , \7924_b1 , w_19724 );
xor ( \7925_b0 , \7924_b0 , w_19726 );
not ( w_19726 , w_19727 );
and ( w_19727 , w_19724 , w_19725 );
buf ( w_19724 , \5775_b1 );
not ( w_19724 , w_19728 );
not ( w_19725 , w_19729 );
and ( w_19728 , w_19729 , \5775_b0 );
or ( \7926_b1 , \6048_b1 , \5790_b1 );
not ( \5790_b1 , w_19730 );
and ( \7926_b0 , \6048_b0 , w_19731 );
and ( w_19730 , w_19731 , \5790_b0 );
or ( \7927_b1 , \6057_b1 , \5788_b1 );
not ( \5788_b1 , w_19732 );
and ( \7927_b0 , \6057_b0 , w_19733 );
and ( w_19732 , w_19733 , \5788_b0 );
or ( \7928_b1 , \7926_b1 , w_19735 );
not ( w_19735 , w_19736 );
and ( \7928_b0 , \7926_b0 , w_19737 );
and ( w_19736 ,  , w_19737 );
buf ( w_19735 , \7927_b1 );
not ( w_19735 , w_19738 );
not (  , w_19739 );
and ( w_19738 , w_19739 , \7927_b0 );
or ( \7929_b1 , \7928_b1 , w_19740 );
xor ( \7929_b0 , \7928_b0 , w_19742 );
not ( w_19742 , w_19743 );
and ( w_19743 , w_19740 , w_19741 );
buf ( w_19740 , \5797_b1 );
not ( w_19740 , w_19744 );
not ( w_19741 , w_19745 );
and ( w_19744 , w_19745 , \5797_b0 );
or ( \7930_b1 , \7925_b1 , \7929_b1 );
xor ( \7930_b0 , \7925_b0 , w_19746 );
not ( w_19746 , w_19747 );
and ( w_19747 , \7929_b1 , \7929_b0 );
or ( \7931_b1 , \6065_b1 , w_19749 );
not ( w_19749 , w_19750 );
and ( \7931_b0 , \6065_b0 , w_19751 );
and ( w_19750 ,  , w_19751 );
buf ( w_19749 , \5807_b1 );
not ( w_19749 , w_19752 );
not (  , w_19753 );
and ( w_19752 , w_19753 , \5807_b0 );
or ( \7932_b1 , \7931_b1 , w_19754 );
xor ( \7932_b0 , \7931_b0 , w_19756 );
not ( w_19756 , w_19757 );
and ( w_19757 , w_19754 , w_19755 );
buf ( w_19754 , \5816_b1 );
not ( w_19754 , w_19758 );
not ( w_19755 , w_19759 );
and ( w_19758 , w_19759 , \5816_b0 );
or ( \7933_b1 , \7930_b1 , \7932_b1 );
xor ( \7933_b0 , \7930_b0 , w_19760 );
not ( w_19760 , w_19761 );
and ( w_19761 , \7932_b1 , \7932_b0 );
or ( \7934_b1 , \7921_b1 , \7933_b1 );
xor ( \7934_b0 , \7921_b0 , w_19762 );
not ( w_19762 , w_19763 );
and ( w_19763 , \7933_b1 , \7933_b0 );
or ( \7935_b1 , \7653_b1 , \7657_b1 );
not ( \7657_b1 , w_19764 );
and ( \7935_b0 , \7653_b0 , w_19765 );
and ( w_19764 , w_19765 , \7657_b0 );
or ( \7936_b1 , \7657_b1 , \7662_b1 );
not ( \7662_b1 , w_19766 );
and ( \7936_b0 , \7657_b0 , w_19767 );
and ( w_19766 , w_19767 , \7662_b0 );
or ( \7937_b1 , \7653_b1 , \7662_b1 );
not ( \7662_b1 , w_19768 );
and ( \7937_b0 , \7653_b0 , w_19769 );
and ( w_19768 , w_19769 , \7662_b0 );
or ( \7939_b1 , \7638_b1 , \7642_b1 );
not ( \7642_b1 , w_19770 );
and ( \7939_b0 , \7638_b0 , w_19771 );
and ( w_19770 , w_19771 , \7642_b0 );
or ( \7940_b1 , \7642_b1 , \7647_b1 );
not ( \7647_b1 , w_19772 );
and ( \7940_b0 , \7642_b0 , w_19773 );
and ( w_19772 , w_19773 , \7647_b0 );
or ( \7941_b1 , \7638_b1 , \7647_b1 );
not ( \7647_b1 , w_19774 );
and ( \7941_b0 , \7638_b0 , w_19775 );
and ( w_19774 , w_19775 , \7647_b0 );
or ( \7943_b1 , \7938_b1 , \7942_b1 );
xor ( \7943_b0 , \7938_b0 , w_19776 );
not ( w_19776 , w_19777 );
and ( w_19777 , \7942_b1 , \7942_b0 );
or ( \7944_b1 , \7722_b1 , \7726_b1 );
not ( \7726_b1 , w_19778 );
and ( \7944_b0 , \7722_b0 , w_19779 );
and ( w_19778 , w_19779 , \7726_b0 );
or ( \7945_b1 , \7726_b1 , \7731_b1 );
not ( \7731_b1 , w_19780 );
and ( \7945_b0 , \7726_b0 , w_19781 );
and ( w_19780 , w_19781 , \7731_b0 );
or ( \7946_b1 , \7722_b1 , \7731_b1 );
not ( \7731_b1 , w_19782 );
and ( \7946_b0 , \7722_b0 , w_19783 );
and ( w_19782 , w_19783 , \7731_b0 );
or ( \7948_b1 , \7943_b1 , \7947_b1 );
xor ( \7948_b0 , \7943_b0 , w_19784 );
not ( w_19784 , w_19785 );
and ( w_19785 , \7947_b1 , \7947_b0 );
or ( \7949_b1 , \7934_b1 , \7948_b1 );
xor ( \7949_b0 , \7934_b0 , w_19786 );
not ( w_19786 , w_19787 );
and ( w_19787 , \7948_b1 , \7948_b0 );
or ( \7950_b1 , \5780_b1 , \7026_b1 );
not ( \7026_b1 , w_19788 );
and ( \7950_b0 , \5780_b0 , w_19789 );
and ( w_19788 , w_19789 , \7026_b0 );
or ( \7951_b1 , \5792_b1 , \7024_b1 );
not ( \7024_b1 , w_19790 );
and ( \7951_b0 , \5792_b0 , w_19791 );
and ( w_19790 , w_19791 , \7024_b0 );
or ( \7952_b1 , \7950_b1 , w_19793 );
not ( w_19793 , w_19794 );
and ( \7952_b0 , \7950_b0 , w_19795 );
and ( w_19794 ,  , w_19795 );
buf ( w_19793 , \7951_b1 );
not ( w_19793 , w_19796 );
not (  , w_19797 );
and ( w_19796 , w_19797 , \7951_b0 );
or ( \7953_b1 , \7952_b1 , w_19798 );
xor ( \7953_b0 , \7952_b0 , w_19800 );
not ( w_19800 , w_19801 );
and ( w_19801 , w_19798 , w_19799 );
buf ( w_19798 , \7032_b1 );
not ( w_19798 , w_19802 );
not ( w_19799 , w_19803 );
and ( w_19802 , w_19803 , \7032_b0 );
or ( \7954_b1 , \5799_b1 , \7043_b1 );
not ( \7043_b1 , w_19804 );
and ( \7954_b0 , \5799_b0 , w_19805 );
and ( w_19804 , w_19805 , \7043_b0 );
or ( \7955_b1 , \5811_b1 , \7041_b1 );
not ( \7041_b1 , w_19806 );
and ( \7955_b0 , \5811_b0 , w_19807 );
and ( w_19806 , w_19807 , \7041_b0 );
or ( \7956_b1 , \7954_b1 , w_19809 );
not ( w_19809 , w_19810 );
and ( \7956_b0 , \7954_b0 , w_19811 );
and ( w_19810 ,  , w_19811 );
buf ( w_19809 , \7955_b1 );
not ( w_19809 , w_19812 );
not (  , w_19813 );
and ( w_19812 , w_19813 , \7955_b0 );
or ( \7957_b1 , \7956_b1 , w_19814 );
xor ( \7957_b0 , \7956_b0 , w_19816 );
not ( w_19816 , w_19817 );
and ( w_19817 , w_19814 , w_19815 );
buf ( w_19814 , \7049_b1 );
not ( w_19814 , w_19818 );
not ( w_19815 , w_19819 );
and ( w_19818 , w_19819 , \7049_b0 );
or ( \7958_b1 , \7953_b1 , \7957_b1 );
xor ( \7958_b0 , \7953_b0 , w_19820 );
not ( w_19820 , w_19821 );
and ( w_19821 , \7957_b1 , \7957_b0 );
or ( \7959_b1 , \5819_b1 , \7061_b1 );
not ( \7061_b1 , w_19822 );
and ( \7959_b0 , \5819_b0 , w_19823 );
and ( w_19822 , w_19823 , \7061_b0 );
or ( \7960_b1 , \5831_b1 , \7059_b1 );
not ( \7059_b1 , w_19824 );
and ( \7960_b0 , \5831_b0 , w_19825 );
and ( w_19824 , w_19825 , \7059_b0 );
or ( \7961_b1 , \7959_b1 , w_19827 );
not ( w_19827 , w_19828 );
and ( \7961_b0 , \7959_b0 , w_19829 );
and ( w_19828 ,  , w_19829 );
buf ( w_19827 , \7960_b1 );
not ( w_19827 , w_19830 );
not (  , w_19831 );
and ( w_19830 , w_19831 , \7960_b0 );
or ( \7962_b1 , \7961_b1 , w_19832 );
xor ( \7962_b0 , \7961_b0 , w_19834 );
not ( w_19834 , w_19835 );
and ( w_19835 , w_19832 , w_19833 );
buf ( w_19832 , \7067_b1 );
not ( w_19832 , w_19836 );
not ( w_19833 , w_19837 );
and ( w_19836 , w_19837 , \7067_b0 );
or ( \7963_b1 , \7958_b1 , \7962_b1 );
xor ( \7963_b0 , \7958_b0 , w_19838 );
not ( w_19838 , w_19839 );
and ( w_19839 , \7962_b1 , \7962_b0 );
or ( \7964_b1 , \5737_b1 , \6991_b1 );
not ( \6991_b1 , w_19840 );
and ( \7964_b0 , \5737_b0 , w_19841 );
and ( w_19840 , w_19841 , \6991_b0 );
buf ( \7965_b1 , \7964_b1 );
not ( \7965_b1 , w_19842 );
not ( \7965_b0 , w_19843 );
and ( w_19842 , w_19843 , \7964_b0 );
or ( \7966_b1 , \7965_b1 , w_19844 );
xor ( \7966_b0 , \7965_b0 , w_19846 );
not ( w_19846 , w_19847 );
and ( w_19847 , w_19844 , w_19845 );
buf ( w_19844 , \6985_b1 );
not ( w_19844 , w_19848 );
not ( w_19845 , w_19849 );
and ( w_19848 , w_19849 , \6985_b0 );
or ( \7967_b1 , \5816_b1 , \7966_b1 );
xor ( \7967_b0 , \5816_b0 , w_19850 );
not ( w_19850 , w_19851 );
and ( w_19851 , \7966_b1 , \7966_b0 );
or ( \7968_b1 , \5758_b1 , \7006_b1 );
not ( \7006_b1 , w_19852 );
and ( \7968_b0 , \5758_b0 , w_19853 );
and ( w_19852 , w_19853 , \7006_b0 );
or ( \7969_b1 , \5770_b1 , \7004_b1 );
not ( \7004_b1 , w_19854 );
and ( \7969_b0 , \5770_b0 , w_19855 );
and ( w_19854 , w_19855 , \7004_b0 );
or ( \7970_b1 , \7968_b1 , w_19857 );
not ( w_19857 , w_19858 );
and ( \7970_b0 , \7968_b0 , w_19859 );
and ( w_19858 ,  , w_19859 );
buf ( w_19857 , \7969_b1 );
not ( w_19857 , w_19860 );
not (  , w_19861 );
and ( w_19860 , w_19861 , \7969_b0 );
or ( \7971_b1 , \7970_b1 , w_19862 );
xor ( \7971_b0 , \7970_b0 , w_19864 );
not ( w_19864 , w_19865 );
and ( w_19865 , w_19862 , w_19863 );
buf ( w_19862 , \7012_b1 );
not ( w_19862 , w_19866 );
not ( w_19863 , w_19867 );
and ( w_19866 , w_19867 , \7012_b0 );
or ( \7972_b1 , \7967_b1 , \7971_b1 );
xor ( \7972_b0 , \7967_b0 , w_19868 );
not ( w_19868 , w_19869 );
and ( w_19869 , \7971_b1 , \7971_b0 );
or ( \7973_b1 , \7963_b1 , \7972_b1 );
xor ( \7973_b0 , \7963_b0 , w_19870 );
not ( w_19870 , w_19871 );
and ( w_19871 , \7972_b1 , \7972_b0 );
or ( \7974_b1 , \5967_b1 , \7192_b1 );
not ( \7192_b1 , w_19872 );
and ( \7974_b0 , \5967_b0 , w_19873 );
and ( w_19872 , w_19873 , \7192_b0 );
or ( \7975_b1 , \5979_b1 , \7190_b1 );
not ( \7190_b1 , w_19874 );
and ( \7975_b0 , \5979_b0 , w_19875 );
and ( w_19874 , w_19875 , \7190_b0 );
or ( \7976_b1 , \7974_b1 , w_19877 );
not ( w_19877 , w_19878 );
and ( \7976_b0 , \7974_b0 , w_19879 );
and ( w_19878 ,  , w_19879 );
buf ( w_19877 , \7975_b1 );
not ( w_19877 , w_19880 );
not (  , w_19881 );
and ( w_19880 , w_19881 , \7975_b0 );
or ( \7977_b1 , \7976_b1 , w_19882 );
xor ( \7977_b0 , \7976_b0 , w_19884 );
not ( w_19884 , w_19885 );
and ( w_19885 , w_19882 , w_19883 );
buf ( w_19882 , \7198_b1 );
not ( w_19882 , w_19886 );
not ( w_19883 , w_19887 );
and ( w_19886 , w_19887 , \7198_b0 );
or ( \7978_b1 , \5986_b1 , \7203_b1 );
not ( \7203_b1 , w_19888 );
and ( \7978_b0 , \5986_b0 , w_19889 );
and ( w_19888 , w_19889 , \7203_b0 );
or ( \7979_b1 , \5998_b1 , \7201_b1 );
not ( \7201_b1 , w_19890 );
and ( \7979_b0 , \5998_b0 , w_19891 );
and ( w_19890 , w_19891 , \7201_b0 );
or ( \7980_b1 , \7978_b1 , w_19893 );
not ( w_19893 , w_19894 );
and ( \7980_b0 , \7978_b0 , w_19895 );
and ( w_19894 ,  , w_19895 );
buf ( w_19893 , \7979_b1 );
not ( w_19893 , w_19896 );
not (  , w_19897 );
and ( w_19896 , w_19897 , \7979_b0 );
or ( \7981_b1 , \7980_b1 , w_19898 );
xor ( \7981_b0 , \7980_b0 , w_19900 );
not ( w_19900 , w_19901 );
and ( w_19901 , w_19898 , w_19899 );
buf ( w_19898 , \6824_b1 );
not ( w_19898 , w_19902 );
not ( w_19899 , w_19903 );
and ( w_19902 , w_19903 , \6824_b0 );
or ( \7982_b1 , \7977_b1 , \7981_b1 );
xor ( \7982_b0 , \7977_b0 , w_19904 );
not ( w_19904 , w_19905 );
and ( w_19905 , \7981_b1 , \7981_b0 );
or ( \7983_b1 , \6006_b1 , \5750_b1 );
not ( \5750_b1 , w_19906 );
and ( \7983_b0 , \6006_b0 , w_19907 );
and ( w_19906 , w_19907 , \5750_b0 );
or ( \7984_b1 , \6018_b1 , \5748_b1 );
not ( \5748_b1 , w_19908 );
and ( \7984_b0 , \6018_b0 , w_19909 );
and ( w_19908 , w_19909 , \5748_b0 );
or ( \7985_b1 , \7983_b1 , w_19911 );
not ( w_19911 , w_19912 );
and ( \7985_b0 , \7983_b0 , w_19913 );
and ( w_19912 ,  , w_19913 );
buf ( w_19911 , \7984_b1 );
not ( w_19911 , w_19914 );
not (  , w_19915 );
and ( w_19914 , w_19915 , \7984_b0 );
or ( \7986_b1 , \7985_b1 , w_19916 );
xor ( \7986_b0 , \7985_b0 , w_19918 );
not ( w_19918 , w_19919 );
and ( w_19919 , w_19916 , w_19917 );
buf ( w_19916 , \5755_b1 );
not ( w_19916 , w_19920 );
not ( w_19917 , w_19921 );
and ( w_19920 , w_19921 , \5755_b0 );
or ( \7987_b1 , \7982_b1 , \7986_b1 );
xor ( \7987_b0 , \7982_b0 , w_19922 );
not ( w_19922 , w_19923 );
and ( w_19923 , \7986_b1 , \7986_b0 );
or ( \7988_b1 , \5906_b1 , \7140_b1 );
not ( \7140_b1 , w_19924 );
and ( \7988_b0 , \5906_b0 , w_19925 );
and ( w_19924 , w_19925 , \7140_b0 );
or ( \7989_b1 , \5918_b1 , \7138_b1 );
not ( \7138_b1 , w_19926 );
and ( \7989_b0 , \5918_b0 , w_19927 );
and ( w_19926 , w_19927 , \7138_b0 );
or ( \7990_b1 , \7988_b1 , w_19929 );
not ( w_19929 , w_19930 );
and ( \7990_b0 , \7988_b0 , w_19931 );
and ( w_19930 ,  , w_19931 );
buf ( w_19929 , \7989_b1 );
not ( w_19929 , w_19932 );
not (  , w_19933 );
and ( w_19932 , w_19933 , \7989_b0 );
or ( \7991_b1 , \7990_b1 , w_19934 );
xor ( \7991_b0 , \7990_b0 , w_19936 );
not ( w_19936 , w_19937 );
and ( w_19937 , w_19934 , w_19935 );
buf ( w_19934 , \7146_b1 );
not ( w_19934 , w_19938 );
not ( w_19935 , w_19939 );
and ( w_19938 , w_19939 , \7146_b0 );
or ( \7992_b1 , \5925_b1 , \7157_b1 );
not ( \7157_b1 , w_19940 );
and ( \7992_b0 , \5925_b0 , w_19941 );
and ( w_19940 , w_19941 , \7157_b0 );
or ( \7993_b1 , \5937_b1 , \7155_b1 );
not ( \7155_b1 , w_19942 );
and ( \7993_b0 , \5937_b0 , w_19943 );
and ( w_19942 , w_19943 , \7155_b0 );
or ( \7994_b1 , \7992_b1 , w_19945 );
not ( w_19945 , w_19946 );
and ( \7994_b0 , \7992_b0 , w_19947 );
and ( w_19946 ,  , w_19947 );
buf ( w_19945 , \7993_b1 );
not ( w_19945 , w_19948 );
not (  , w_19949 );
and ( w_19948 , w_19949 , \7993_b0 );
or ( \7995_b1 , \7994_b1 , w_19950 );
xor ( \7995_b0 , \7994_b0 , w_19952 );
not ( w_19952 , w_19953 );
and ( w_19953 , w_19950 , w_19951 );
buf ( w_19950 , \7163_b1 );
not ( w_19950 , w_19954 );
not ( w_19951 , w_19955 );
and ( w_19954 , w_19955 , \7163_b0 );
or ( \7996_b1 , \7991_b1 , \7995_b1 );
xor ( \7996_b0 , \7991_b0 , w_19956 );
not ( w_19956 , w_19957 );
and ( w_19957 , \7995_b1 , \7995_b0 );
or ( \7997_b1 , \5945_b1 , \7175_b1 );
not ( \7175_b1 , w_19958 );
and ( \7997_b0 , \5945_b0 , w_19959 );
and ( w_19958 , w_19959 , \7175_b0 );
or ( \7998_b1 , \5957_b1 , \7173_b1 );
not ( \7173_b1 , w_19960 );
and ( \7998_b0 , \5957_b0 , w_19961 );
and ( w_19960 , w_19961 , \7173_b0 );
or ( \7999_b1 , \7997_b1 , w_19963 );
not ( w_19963 , w_19964 );
and ( \7999_b0 , \7997_b0 , w_19965 );
and ( w_19964 ,  , w_19965 );
buf ( w_19963 , \7998_b1 );
not ( w_19963 , w_19966 );
not (  , w_19967 );
and ( w_19966 , w_19967 , \7998_b0 );
or ( \8000_b1 , \7999_b1 , w_19968 );
xor ( \8000_b0 , \7999_b0 , w_19970 );
not ( w_19970 , w_19971 );
and ( w_19971 , w_19968 , w_19969 );
buf ( w_19968 , \7181_b1 );
not ( w_19968 , w_19972 );
not ( w_19969 , w_19973 );
and ( w_19972 , w_19973 , \7181_b0 );
or ( \8001_b1 , \7996_b1 , \8000_b1 );
xor ( \8001_b0 , \7996_b0 , w_19974 );
not ( w_19974 , w_19975 );
and ( w_19975 , \8000_b1 , \8000_b0 );
or ( \8002_b1 , \7987_b1 , \8001_b1 );
xor ( \8002_b0 , \7987_b0 , w_19976 );
not ( w_19976 , w_19977 );
and ( w_19977 , \8001_b1 , \8001_b0 );
or ( \8003_b1 , \5842_b1 , \7082_b1 );
not ( \7082_b1 , w_19978 );
and ( \8003_b0 , \5842_b0 , w_19979 );
and ( w_19978 , w_19979 , \7082_b0 );
or ( \8004_b1 , \5854_b1 , \7080_b1 );
not ( \7080_b1 , w_19980 );
and ( \8004_b0 , \5854_b0 , w_19981 );
and ( w_19980 , w_19981 , \7080_b0 );
or ( \8005_b1 , \8003_b1 , w_19983 );
not ( w_19983 , w_19984 );
and ( \8005_b0 , \8003_b0 , w_19985 );
and ( w_19984 ,  , w_19985 );
buf ( w_19983 , \8004_b1 );
not ( w_19983 , w_19986 );
not (  , w_19987 );
and ( w_19986 , w_19987 , \8004_b0 );
or ( \8006_b1 , \8005_b1 , w_19988 );
xor ( \8006_b0 , \8005_b0 , w_19990 );
not ( w_19990 , w_19991 );
and ( w_19991 , w_19988 , w_19989 );
buf ( w_19988 , \7088_b1 );
not ( w_19988 , w_19992 );
not ( w_19989 , w_19993 );
and ( w_19992 , w_19993 , \7088_b0 );
or ( \8007_b1 , \5861_b1 , \7099_b1 );
not ( \7099_b1 , w_19994 );
and ( \8007_b0 , \5861_b0 , w_19995 );
and ( w_19994 , w_19995 , \7099_b0 );
or ( \8008_b1 , \5873_b1 , \7097_b1 );
not ( \7097_b1 , w_19996 );
and ( \8008_b0 , \5873_b0 , w_19997 );
and ( w_19996 , w_19997 , \7097_b0 );
or ( \8009_b1 , \8007_b1 , w_19999 );
not ( w_19999 , w_20000 );
and ( \8009_b0 , \8007_b0 , w_20001 );
and ( w_20000 ,  , w_20001 );
buf ( w_19999 , \8008_b1 );
not ( w_19999 , w_20002 );
not (  , w_20003 );
and ( w_20002 , w_20003 , \8008_b0 );
or ( \8010_b1 , \8009_b1 , w_20004 );
xor ( \8010_b0 , \8009_b0 , w_20006 );
not ( w_20006 , w_20007 );
and ( w_20007 , w_20004 , w_20005 );
buf ( w_20004 , \7105_b1 );
not ( w_20004 , w_20008 );
not ( w_20005 , w_20009 );
and ( w_20008 , w_20009 , \7105_b0 );
or ( \8011_b1 , \8006_b1 , \8010_b1 );
xor ( \8011_b0 , \8006_b0 , w_20010 );
not ( w_20010 , w_20011 );
and ( w_20011 , \8010_b1 , \8010_b0 );
or ( \8012_b1 , \5881_b1 , \7117_b1 );
not ( \7117_b1 , w_20012 );
and ( \8012_b0 , \5881_b0 , w_20013 );
and ( w_20012 , w_20013 , \7117_b0 );
or ( \8013_b1 , \5893_b1 , \7115_b1 );
not ( \7115_b1 , w_20014 );
and ( \8013_b0 , \5893_b0 , w_20015 );
and ( w_20014 , w_20015 , \7115_b0 );
or ( \8014_b1 , \8012_b1 , w_20017 );
not ( w_20017 , w_20018 );
and ( \8014_b0 , \8012_b0 , w_20019 );
and ( w_20018 ,  , w_20019 );
buf ( w_20017 , \8013_b1 );
not ( w_20017 , w_20020 );
not (  , w_20021 );
and ( w_20020 , w_20021 , \8013_b0 );
or ( \8015_b1 , \8014_b1 , w_20022 );
xor ( \8015_b0 , \8014_b0 , w_20024 );
not ( w_20024 , w_20025 );
and ( w_20025 , w_20022 , w_20023 );
buf ( w_20022 , \7123_b1 );
not ( w_20022 , w_20026 );
not ( w_20023 , w_20027 );
and ( w_20026 , w_20027 , \7123_b0 );
or ( \8016_b1 , \8011_b1 , \8015_b1 );
xor ( \8016_b0 , \8011_b0 , w_20028 );
not ( w_20028 , w_20029 );
and ( w_20029 , \8015_b1 , \8015_b0 );
or ( \8017_b1 , \8002_b1 , \8016_b1 );
xor ( \8017_b0 , \8002_b0 , w_20030 );
not ( w_20030 , w_20031 );
and ( w_20031 , \8016_b1 , \8016_b0 );
or ( \8018_b1 , \7973_b1 , \8017_b1 );
xor ( \8018_b0 , \7973_b0 , w_20032 );
not ( w_20032 , w_20033 );
and ( w_20033 , \8017_b1 , \8017_b0 );
or ( \8019_b1 , \7949_b1 , \8018_b1 );
xor ( \8019_b0 , \7949_b0 , w_20034 );
not ( w_20034 , w_20035 );
and ( w_20035 , \8018_b1 , \8018_b0 );
or ( \8020_b1 , \7752_b1 , \7756_b1 );
not ( \7756_b1 , w_20036 );
and ( \8020_b0 , \7752_b0 , w_20037 );
and ( w_20036 , w_20037 , \7756_b0 );
or ( \8021_b1 , \7756_b1 , \7761_b1 );
not ( \7761_b1 , w_20038 );
and ( \8021_b0 , \7756_b0 , w_20039 );
and ( w_20038 , w_20039 , \7761_b0 );
or ( \8022_b1 , \7752_b1 , \7761_b1 );
not ( \7761_b1 , w_20040 );
and ( \8022_b0 , \7752_b0 , w_20041 );
and ( w_20040 , w_20041 , \7761_b0 );
or ( \8024_b1 , \7737_b1 , \7741_b1 );
not ( \7741_b1 , w_20042 );
and ( \8024_b0 , \7737_b0 , w_20043 );
and ( w_20042 , w_20043 , \7741_b0 );
or ( \8025_b1 , \7741_b1 , \7746_b1 );
not ( \7746_b1 , w_20044 );
and ( \8025_b0 , \7741_b0 , w_20045 );
and ( w_20044 , w_20045 , \7746_b0 );
or ( \8026_b1 , \7737_b1 , \7746_b1 );
not ( \7746_b1 , w_20046 );
and ( \8026_b0 , \7737_b0 , w_20047 );
and ( w_20046 , w_20047 , \7746_b0 );
or ( \8028_b1 , \8023_b1 , \8027_b1 );
xor ( \8028_b0 , \8023_b0 , w_20048 );
not ( w_20048 , w_20049 );
and ( w_20049 , \8027_b1 , \8027_b0 );
or ( \8029_b1 , \7703_b1 , \7717_b1 );
not ( \7717_b1 , w_20050 );
and ( \8029_b0 , \7703_b0 , w_20051 );
and ( w_20050 , w_20051 , \7717_b0 );
or ( \8030_b1 , \7717_b1 , \7732_b1 );
not ( \7732_b1 , w_20052 );
and ( \8030_b0 , \7717_b0 , w_20053 );
and ( w_20052 , w_20053 , \7732_b0 );
or ( \8031_b1 , \7703_b1 , \7732_b1 );
not ( \7732_b1 , w_20054 );
and ( \8031_b0 , \7703_b0 , w_20055 );
and ( w_20054 , w_20055 , \7732_b0 );
or ( \8033_b1 , \8028_b1 , \8032_b1 );
xor ( \8033_b0 , \8028_b0 , w_20056 );
not ( w_20056 , w_20057 );
and ( w_20057 , \8032_b1 , \8032_b0 );
or ( \8034_b1 , \8019_b1 , \8033_b1 );
xor ( \8034_b0 , \8019_b0 , w_20058 );
not ( w_20058 , w_20059 );
and ( w_20059 , \8033_b1 , \8033_b0 );
or ( \8035_b1 , \7912_b1 , \8034_b1 );
xor ( \8035_b0 , \7912_b0 , w_20060 );
not ( w_20060 , w_20061 );
and ( w_20061 , \8034_b1 , \8034_b0 );
or ( \8036_b1 , \7906_b1 , \8035_b1 );
xor ( \8036_b0 , \7906_b0 , w_20062 );
not ( w_20062 , w_20063 );
and ( w_20063 , \8035_b1 , \8035_b0 );
or ( \8037_b1 , \7586_b1 , \7625_b1 );
not ( \7625_b1 , w_20064 );
and ( \8037_b0 , \7586_b0 , w_20065 );
and ( w_20064 , w_20065 , \7625_b0 );
or ( \8038_b1 , \7625_b1 , \7765_b1 );
not ( \7765_b1 , w_20066 );
and ( \8038_b0 , \7625_b0 , w_20067 );
and ( w_20066 , w_20067 , \7765_b0 );
or ( \8039_b1 , \7586_b1 , \7765_b1 );
not ( \7765_b1 , w_20068 );
and ( \8039_b0 , \7586_b0 , w_20069 );
and ( w_20068 , w_20069 , \7765_b0 );
or ( \8041_b1 , \8036_b1 , w_20071 );
not ( w_20071 , w_20072 );
and ( \8041_b0 , \8036_b0 , w_20073 );
and ( w_20072 ,  , w_20073 );
buf ( w_20071 , \8040_b1 );
not ( w_20071 , w_20074 );
not (  , w_20075 );
and ( w_20074 , w_20075 , \8040_b0 );
or ( \8042_b1 , \7887_b1 , w_20077 );
not ( w_20077 , w_20078 );
and ( \8042_b0 , \7887_b0 , w_20079 );
and ( w_20078 ,  , w_20079 );
buf ( w_20077 , \8041_b1 );
not ( w_20077 , w_20080 );
not (  , w_20081 );
and ( w_20080 , w_20081 , \8041_b0 );
or ( \8043_b1 , \7910_b1 , \7911_b1 );
not ( \7911_b1 , w_20082 );
and ( \8043_b0 , \7910_b0 , w_20083 );
and ( w_20082 , w_20083 , \7911_b0 );
or ( \8044_b1 , \7911_b1 , \8034_b1 );
not ( \8034_b1 , w_20084 );
and ( \8044_b0 , \7911_b0 , w_20085 );
and ( w_20084 , w_20085 , \8034_b0 );
or ( \8045_b1 , \7910_b1 , \8034_b1 );
not ( \8034_b1 , w_20086 );
and ( \8045_b0 , \7910_b0 , w_20087 );
and ( w_20086 , w_20087 , \8034_b0 );
or ( \8047_b1 , \8023_b1 , \8027_b1 );
not ( \8027_b1 , w_20088 );
and ( \8047_b0 , \8023_b0 , w_20089 );
and ( w_20088 , w_20089 , \8027_b0 );
or ( \8048_b1 , \8027_b1 , \8032_b1 );
not ( \8032_b1 , w_20090 );
and ( \8048_b0 , \8027_b0 , w_20091 );
and ( w_20090 , w_20091 , \8032_b0 );
or ( \8049_b1 , \8023_b1 , \8032_b1 );
not ( \8032_b1 , w_20092 );
and ( \8049_b0 , \8023_b0 , w_20093 );
and ( w_20092 , w_20093 , \8032_b0 );
or ( \8051_b1 , \7963_b1 , \7972_b1 );
not ( \7972_b1 , w_20094 );
and ( \8051_b0 , \7963_b0 , w_20095 );
and ( w_20094 , w_20095 , \7972_b0 );
or ( \8052_b1 , \7972_b1 , \8017_b1 );
not ( \8017_b1 , w_20096 );
and ( \8052_b0 , \7972_b0 , w_20097 );
and ( w_20096 , w_20097 , \8017_b0 );
or ( \8053_b1 , \7963_b1 , \8017_b1 );
not ( \8017_b1 , w_20098 );
and ( \8053_b0 , \7963_b0 , w_20099 );
and ( w_20098 , w_20099 , \8017_b0 );
or ( \8055_b1 , \8050_b1 , \8054_b1 );
xor ( \8055_b0 , \8050_b0 , w_20100 );
not ( w_20100 , w_20101 );
and ( w_20101 , \8054_b1 , \8054_b0 );
or ( \8056_b1 , \7934_b1 , \7948_b1 );
not ( \7948_b1 , w_20102 );
and ( \8056_b0 , \7934_b0 , w_20103 );
and ( w_20102 , w_20103 , \7948_b0 );
or ( \8057_b1 , \8055_b1 , \8056_b1 );
xor ( \8057_b0 , \8055_b0 , w_20104 );
not ( w_20104 , w_20105 );
and ( w_20105 , \8056_b1 , \8056_b0 );
or ( \8058_b1 , \8046_b1 , \8057_b1 );
xor ( \8058_b0 , \8046_b0 , w_20106 );
not ( w_20106 , w_20107 );
and ( w_20107 , \8057_b1 , \8057_b0 );
or ( \8059_b1 , \7895_b1 , \7899_b1 );
not ( \7899_b1 , w_20108 );
and ( \8059_b0 , \7895_b0 , w_20109 );
and ( w_20108 , w_20109 , \7899_b0 );
or ( \8060_b1 , \7899_b1 , \7904_b1 );
not ( \7904_b1 , w_20110 );
and ( \8060_b0 , \7899_b0 , w_20111 );
and ( w_20110 , w_20111 , \7904_b0 );
or ( \8061_b1 , \7895_b1 , \7904_b1 );
not ( \7904_b1 , w_20112 );
and ( \8061_b0 , \7895_b0 , w_20113 );
and ( w_20112 , w_20113 , \7904_b0 );
or ( \8063_b1 , \7949_b1 , \8018_b1 );
not ( \8018_b1 , w_20114 );
and ( \8063_b0 , \7949_b0 , w_20115 );
and ( w_20114 , w_20115 , \8018_b0 );
or ( \8064_b1 , \8018_b1 , \8033_b1 );
not ( \8033_b1 , w_20116 );
and ( \8064_b0 , \8018_b0 , w_20117 );
and ( w_20116 , w_20117 , \8033_b0 );
or ( \8065_b1 , \7949_b1 , \8033_b1 );
not ( \8033_b1 , w_20118 );
and ( \8065_b0 , \7949_b0 , w_20119 );
and ( w_20118 , w_20119 , \8033_b0 );
or ( \8067_b1 , \8062_b1 , \8066_b1 );
xor ( \8067_b0 , \8062_b0 , w_20120 );
not ( w_20120 , w_20121 );
and ( w_20121 , \8066_b1 , \8066_b0 );
or ( \8068_b1 , \5816_b1 , \7966_b1 );
not ( \7966_b1 , w_20122 );
and ( \8068_b0 , \5816_b0 , w_20123 );
and ( w_20122 , w_20123 , \7966_b0 );
or ( \8069_b1 , \7966_b1 , \7971_b1 );
not ( \7971_b1 , w_20124 );
and ( \8069_b0 , \7966_b0 , w_20125 );
and ( w_20124 , w_20125 , \7971_b0 );
or ( \8070_b1 , \5816_b1 , \7971_b1 );
not ( \7971_b1 , w_20126 );
and ( \8070_b0 , \5816_b0 , w_20127 );
and ( w_20126 , w_20127 , \7971_b0 );
or ( \8072_b1 , \7953_b1 , \7957_b1 );
not ( \7957_b1 , w_20128 );
and ( \8072_b0 , \7953_b0 , w_20129 );
and ( w_20128 , w_20129 , \7957_b0 );
or ( \8073_b1 , \7957_b1 , \7962_b1 );
not ( \7962_b1 , w_20130 );
and ( \8073_b0 , \7957_b0 , w_20131 );
and ( w_20130 , w_20131 , \7962_b0 );
or ( \8074_b1 , \7953_b1 , \7962_b1 );
not ( \7962_b1 , w_20132 );
and ( \8074_b0 , \7953_b0 , w_20133 );
and ( w_20132 , w_20133 , \7962_b0 );
or ( \8076_b1 , \8071_b1 , \8075_b1 );
xor ( \8076_b0 , \8071_b0 , w_20134 );
not ( w_20134 , w_20135 );
and ( w_20135 , \8075_b1 , \8075_b0 );
or ( \8077_b1 , \8006_b1 , \8010_b1 );
not ( \8010_b1 , w_20136 );
and ( \8077_b0 , \8006_b0 , w_20137 );
and ( w_20136 , w_20137 , \8010_b0 );
or ( \8078_b1 , \8010_b1 , \8015_b1 );
not ( \8015_b1 , w_20138 );
and ( \8078_b0 , \8010_b0 , w_20139 );
and ( w_20138 , w_20139 , \8015_b0 );
or ( \8079_b1 , \8006_b1 , \8015_b1 );
not ( \8015_b1 , w_20140 );
and ( \8079_b0 , \8006_b0 , w_20141 );
and ( w_20140 , w_20141 , \8015_b0 );
or ( \8081_b1 , \8076_b1 , \8080_b1 );
xor ( \8081_b0 , \8076_b0 , w_20142 );
not ( w_20142 , w_20143 );
and ( w_20143 , \8080_b1 , \8080_b0 );
or ( \8082_b1 , \5873_b1 , \7099_b1 );
not ( \7099_b1 , w_20144 );
and ( \8082_b0 , \5873_b0 , w_20145 );
and ( w_20144 , w_20145 , \7099_b0 );
or ( \8083_b1 , \5842_b1 , \7097_b1 );
not ( \7097_b1 , w_20146 );
and ( \8083_b0 , \5842_b0 , w_20147 );
and ( w_20146 , w_20147 , \7097_b0 );
or ( \8084_b1 , \8082_b1 , w_20149 );
not ( w_20149 , w_20150 );
and ( \8084_b0 , \8082_b0 , w_20151 );
and ( w_20150 ,  , w_20151 );
buf ( w_20149 , \8083_b1 );
not ( w_20149 , w_20152 );
not (  , w_20153 );
and ( w_20152 , w_20153 , \8083_b0 );
or ( \8085_b1 , \8084_b1 , w_20154 );
xor ( \8085_b0 , \8084_b0 , w_20156 );
not ( w_20156 , w_20157 );
and ( w_20157 , w_20154 , w_20155 );
buf ( w_20154 , \7105_b1 );
not ( w_20154 , w_20158 );
not ( w_20155 , w_20159 );
and ( w_20158 , w_20159 , \7105_b0 );
or ( \8086_b1 , \5893_b1 , \7117_b1 );
not ( \7117_b1 , w_20160 );
and ( \8086_b0 , \5893_b0 , w_20161 );
and ( w_20160 , w_20161 , \7117_b0 );
or ( \8087_b1 , \5861_b1 , \7115_b1 );
not ( \7115_b1 , w_20162 );
and ( \8087_b0 , \5861_b0 , w_20163 );
and ( w_20162 , w_20163 , \7115_b0 );
or ( \8088_b1 , \8086_b1 , w_20165 );
not ( w_20165 , w_20166 );
and ( \8088_b0 , \8086_b0 , w_20167 );
and ( w_20166 ,  , w_20167 );
buf ( w_20165 , \8087_b1 );
not ( w_20165 , w_20168 );
not (  , w_20169 );
and ( w_20168 , w_20169 , \8087_b0 );
or ( \8089_b1 , \8088_b1 , w_20170 );
xor ( \8089_b0 , \8088_b0 , w_20172 );
not ( w_20172 , w_20173 );
and ( w_20173 , w_20170 , w_20171 );
buf ( w_20170 , \7123_b1 );
not ( w_20170 , w_20174 );
not ( w_20171 , w_20175 );
and ( w_20174 , w_20175 , \7123_b0 );
or ( \8090_b1 , \8085_b1 , \8089_b1 );
xor ( \8090_b0 , \8085_b0 , w_20176 );
not ( w_20176 , w_20177 );
and ( w_20177 , \8089_b1 , \8089_b0 );
or ( \8091_b1 , \5918_b1 , \7140_b1 );
not ( \7140_b1 , w_20178 );
and ( \8091_b0 , \5918_b0 , w_20179 );
and ( w_20178 , w_20179 , \7140_b0 );
or ( \8092_b1 , \5881_b1 , \7138_b1 );
not ( \7138_b1 , w_20180 );
and ( \8092_b0 , \5881_b0 , w_20181 );
and ( w_20180 , w_20181 , \7138_b0 );
or ( \8093_b1 , \8091_b1 , w_20183 );
not ( w_20183 , w_20184 );
and ( \8093_b0 , \8091_b0 , w_20185 );
and ( w_20184 ,  , w_20185 );
buf ( w_20183 , \8092_b1 );
not ( w_20183 , w_20186 );
not (  , w_20187 );
and ( w_20186 , w_20187 , \8092_b0 );
or ( \8094_b1 , \8093_b1 , w_20188 );
xor ( \8094_b0 , \8093_b0 , w_20190 );
not ( w_20190 , w_20191 );
and ( w_20191 , w_20188 , w_20189 );
buf ( w_20188 , \7146_b1 );
not ( w_20188 , w_20192 );
not ( w_20189 , w_20193 );
and ( w_20192 , w_20193 , \7146_b0 );
or ( \8095_b1 , \8090_b1 , \8094_b1 );
xor ( \8095_b0 , \8090_b0 , w_20194 );
not ( w_20194 , w_20195 );
and ( w_20195 , \8094_b1 , \8094_b0 );
or ( \8096_b1 , \5811_b1 , \7043_b1 );
not ( \7043_b1 , w_20196 );
and ( \8096_b0 , \5811_b0 , w_20197 );
and ( w_20196 , w_20197 , \7043_b0 );
or ( \8097_b1 , \5780_b1 , \7041_b1 );
not ( \7041_b1 , w_20198 );
and ( \8097_b0 , \5780_b0 , w_20199 );
and ( w_20198 , w_20199 , \7041_b0 );
or ( \8098_b1 , \8096_b1 , w_20201 );
not ( w_20201 , w_20202 );
and ( \8098_b0 , \8096_b0 , w_20203 );
and ( w_20202 ,  , w_20203 );
buf ( w_20201 , \8097_b1 );
not ( w_20201 , w_20204 );
not (  , w_20205 );
and ( w_20204 , w_20205 , \8097_b0 );
or ( \8099_b1 , \8098_b1 , w_20206 );
xor ( \8099_b0 , \8098_b0 , w_20208 );
not ( w_20208 , w_20209 );
and ( w_20209 , w_20206 , w_20207 );
buf ( w_20206 , \7049_b1 );
not ( w_20206 , w_20210 );
not ( w_20207 , w_20211 );
and ( w_20210 , w_20211 , \7049_b0 );
or ( \8100_b1 , \5831_b1 , \7061_b1 );
not ( \7061_b1 , w_20212 );
and ( \8100_b0 , \5831_b0 , w_20213 );
and ( w_20212 , w_20213 , \7061_b0 );
or ( \8101_b1 , \5799_b1 , \7059_b1 );
not ( \7059_b1 , w_20214 );
and ( \8101_b0 , \5799_b0 , w_20215 );
and ( w_20214 , w_20215 , \7059_b0 );
or ( \8102_b1 , \8100_b1 , w_20217 );
not ( w_20217 , w_20218 );
and ( \8102_b0 , \8100_b0 , w_20219 );
and ( w_20218 ,  , w_20219 );
buf ( w_20217 , \8101_b1 );
not ( w_20217 , w_20220 );
not (  , w_20221 );
and ( w_20220 , w_20221 , \8101_b0 );
or ( \8103_b1 , \8102_b1 , w_20222 );
xor ( \8103_b0 , \8102_b0 , w_20224 );
not ( w_20224 , w_20225 );
and ( w_20225 , w_20222 , w_20223 );
buf ( w_20222 , \7067_b1 );
not ( w_20222 , w_20226 );
not ( w_20223 , w_20227 );
and ( w_20226 , w_20227 , \7067_b0 );
or ( \8104_b1 , \8099_b1 , \8103_b1 );
xor ( \8104_b0 , \8099_b0 , w_20228 );
not ( w_20228 , w_20229 );
and ( w_20229 , \8103_b1 , \8103_b0 );
or ( \8105_b1 , \5854_b1 , \7082_b1 );
not ( \7082_b1 , w_20230 );
and ( \8105_b0 , \5854_b0 , w_20231 );
and ( w_20230 , w_20231 , \7082_b0 );
or ( \8106_b1 , \5819_b1 , \7080_b1 );
not ( \7080_b1 , w_20232 );
and ( \8106_b0 , \5819_b0 , w_20233 );
and ( w_20232 , w_20233 , \7080_b0 );
or ( \8107_b1 , \8105_b1 , w_20235 );
not ( w_20235 , w_20236 );
and ( \8107_b0 , \8105_b0 , w_20237 );
and ( w_20236 ,  , w_20237 );
buf ( w_20235 , \8106_b1 );
not ( w_20235 , w_20238 );
not (  , w_20239 );
and ( w_20238 , w_20239 , \8106_b0 );
or ( \8108_b1 , \8107_b1 , w_20240 );
xor ( \8108_b0 , \8107_b0 , w_20242 );
not ( w_20242 , w_20243 );
and ( w_20243 , w_20240 , w_20241 );
buf ( w_20240 , \7088_b1 );
not ( w_20240 , w_20244 );
not ( w_20241 , w_20245 );
and ( w_20244 , w_20245 , \7088_b0 );
or ( \8109_b1 , \8104_b1 , \8108_b1 );
xor ( \8109_b0 , \8104_b0 , w_20246 );
not ( w_20246 , w_20247 );
and ( w_20247 , \8108_b1 , \8108_b0 );
or ( \8110_b1 , \8095_b1 , \8109_b1 );
xor ( \8110_b0 , \8095_b0 , w_20248 );
not ( w_20248 , w_20249 );
and ( w_20249 , \8109_b1 , \8109_b0 );
buf ( \8111_b1 , \6985_b1 );
not ( \8111_b1 , w_20250 );
not ( \8111_b0 , w_20251 );
and ( w_20250 , w_20251 , \6985_b0 );
or ( \8112_b1 , \5770_b1 , \7006_b1 );
not ( \7006_b1 , w_20252 );
and ( \8112_b0 , \5770_b0 , w_20253 );
and ( w_20252 , w_20253 , \7006_b0 );
or ( \8113_b1 , \5737_b1 , \7004_b1 );
not ( \7004_b1 , w_20254 );
and ( \8113_b0 , \5737_b0 , w_20255 );
and ( w_20254 , w_20255 , \7004_b0 );
or ( \8114_b1 , \8112_b1 , w_20257 );
not ( w_20257 , w_20258 );
and ( \8114_b0 , \8112_b0 , w_20259 );
and ( w_20258 ,  , w_20259 );
buf ( w_20257 , \8113_b1 );
not ( w_20257 , w_20260 );
not (  , w_20261 );
and ( w_20260 , w_20261 , \8113_b0 );
or ( \8115_b1 , \8114_b1 , w_20262 );
xor ( \8115_b0 , \8114_b0 , w_20264 );
not ( w_20264 , w_20265 );
and ( w_20265 , w_20262 , w_20263 );
buf ( w_20262 , \7012_b1 );
not ( w_20262 , w_20266 );
not ( w_20263 , w_20267 );
and ( w_20266 , w_20267 , \7012_b0 );
or ( \8116_b1 , \8111_b1 , \8115_b1 );
xor ( \8116_b0 , \8111_b0 , w_20268 );
not ( w_20268 , w_20269 );
and ( w_20269 , \8115_b1 , \8115_b0 );
or ( \8117_b1 , \5792_b1 , \7026_b1 );
not ( \7026_b1 , w_20270 );
and ( \8117_b0 , \5792_b0 , w_20271 );
and ( w_20270 , w_20271 , \7026_b0 );
or ( \8118_b1 , \5758_b1 , \7024_b1 );
not ( \7024_b1 , w_20272 );
and ( \8118_b0 , \5758_b0 , w_20273 );
and ( w_20272 , w_20273 , \7024_b0 );
or ( \8119_b1 , \8117_b1 , w_20275 );
not ( w_20275 , w_20276 );
and ( \8119_b0 , \8117_b0 , w_20277 );
and ( w_20276 ,  , w_20277 );
buf ( w_20275 , \8118_b1 );
not ( w_20275 , w_20278 );
not (  , w_20279 );
and ( w_20278 , w_20279 , \8118_b0 );
or ( \8120_b1 , \8119_b1 , w_20280 );
xor ( \8120_b0 , \8119_b0 , w_20282 );
not ( w_20282 , w_20283 );
and ( w_20283 , w_20280 , w_20281 );
buf ( w_20280 , \7032_b1 );
not ( w_20280 , w_20284 );
not ( w_20281 , w_20285 );
and ( w_20284 , w_20285 , \7032_b0 );
or ( \8121_b1 , \8116_b1 , \8120_b1 );
xor ( \8121_b0 , \8116_b0 , w_20286 );
not ( w_20286 , w_20287 );
and ( w_20287 , \8120_b1 , \8120_b0 );
or ( \8122_b1 , \8110_b1 , \8121_b1 );
xor ( \8122_b0 , \8110_b0 , w_20288 );
not ( w_20288 , w_20289 );
and ( w_20289 , \8121_b1 , \8121_b0 );
or ( \8123_b1 , \6057_b1 , \5790_b1 );
not ( \5790_b1 , w_20290 );
and ( \8123_b0 , \6057_b0 , w_20291 );
and ( w_20290 , w_20291 , \5790_b0 );
or ( \8124_b1 , \6029_b1 , \5788_b1 );
not ( \5788_b1 , w_20292 );
and ( \8124_b0 , \6029_b0 , w_20293 );
and ( w_20292 , w_20293 , \5788_b0 );
or ( \8125_b1 , \8123_b1 , w_20295 );
not ( w_20295 , w_20296 );
and ( \8125_b0 , \8123_b0 , w_20297 );
and ( w_20296 ,  , w_20297 );
buf ( w_20295 , \8124_b1 );
not ( w_20295 , w_20298 );
not (  , w_20299 );
and ( w_20298 , w_20299 , \8124_b0 );
or ( \8126_b1 , \8125_b1 , w_20300 );
xor ( \8126_b0 , \8125_b0 , w_20302 );
not ( w_20302 , w_20303 );
and ( w_20303 , w_20300 , w_20301 );
buf ( w_20300 , \5797_b1 );
not ( w_20300 , w_20304 );
not ( w_20301 , w_20305 );
and ( w_20304 , w_20305 , \5797_b0 );
or ( \8127_b1 , \6065_b1 , \5809_b1 );
not ( \5809_b1 , w_20306 );
and ( \8127_b0 , \6065_b0 , w_20307 );
and ( w_20306 , w_20307 , \5809_b0 );
or ( \8128_b1 , \6048_b1 , \5807_b1 );
not ( \5807_b1 , w_20308 );
and ( \8128_b0 , \6048_b0 , w_20309 );
and ( w_20308 , w_20309 , \5807_b0 );
or ( \8129_b1 , \8127_b1 , w_20311 );
not ( w_20311 , w_20312 );
and ( \8129_b0 , \8127_b0 , w_20313 );
and ( w_20312 ,  , w_20313 );
buf ( w_20311 , \8128_b1 );
not ( w_20311 , w_20314 );
not (  , w_20315 );
and ( w_20314 , w_20315 , \8128_b0 );
or ( \8130_b1 , \8129_b1 , w_20316 );
xor ( \8130_b0 , \8129_b0 , w_20318 );
not ( w_20318 , w_20319 );
and ( w_20319 , w_20316 , w_20317 );
buf ( w_20316 , \5816_b1 );
not ( w_20316 , w_20320 );
not ( w_20317 , w_20321 );
and ( w_20320 , w_20321 , \5816_b0 );
or ( \8131_b1 , \8126_b1 , w_20322 );
xor ( \8131_b0 , \8126_b0 , w_20324 );
not ( w_20324 , w_20325 );
and ( w_20325 , w_20322 , w_20323 );
buf ( w_20322 , \8130_b1 );
not ( w_20322 , w_20326 );
not ( w_20323 , w_20327 );
and ( w_20326 , w_20327 , \8130_b0 );
or ( \8132_b1 , \5998_b1 , \7203_b1 );
not ( \7203_b1 , w_20328 );
and ( \8132_b0 , \5998_b0 , w_20329 );
and ( w_20328 , w_20329 , \7203_b0 );
or ( \8133_b1 , \5967_b1 , \7201_b1 );
not ( \7201_b1 , w_20330 );
and ( \8133_b0 , \5967_b0 , w_20331 );
and ( w_20330 , w_20331 , \7201_b0 );
or ( \8134_b1 , \8132_b1 , w_20333 );
not ( w_20333 , w_20334 );
and ( \8134_b0 , \8132_b0 , w_20335 );
and ( w_20334 ,  , w_20335 );
buf ( w_20333 , \8133_b1 );
not ( w_20333 , w_20336 );
not (  , w_20337 );
and ( w_20336 , w_20337 , \8133_b0 );
or ( \8135_b1 , \8134_b1 , w_20338 );
xor ( \8135_b0 , \8134_b0 , w_20340 );
not ( w_20340 , w_20341 );
and ( w_20341 , w_20338 , w_20339 );
buf ( w_20338 , \6824_b1 );
not ( w_20338 , w_20342 );
not ( w_20339 , w_20343 );
and ( w_20342 , w_20343 , \6824_b0 );
or ( \8136_b1 , \6018_b1 , \5750_b1 );
not ( \5750_b1 , w_20344 );
and ( \8136_b0 , \6018_b0 , w_20345 );
and ( w_20344 , w_20345 , \5750_b0 );
or ( \8137_b1 , \5986_b1 , \5748_b1 );
not ( \5748_b1 , w_20346 );
and ( \8137_b0 , \5986_b0 , w_20347 );
and ( w_20346 , w_20347 , \5748_b0 );
or ( \8138_b1 , \8136_b1 , w_20349 );
not ( w_20349 , w_20350 );
and ( \8138_b0 , \8136_b0 , w_20351 );
and ( w_20350 ,  , w_20351 );
buf ( w_20349 , \8137_b1 );
not ( w_20349 , w_20352 );
not (  , w_20353 );
and ( w_20352 , w_20353 , \8137_b0 );
or ( \8139_b1 , \8138_b1 , w_20354 );
xor ( \8139_b0 , \8138_b0 , w_20356 );
not ( w_20356 , w_20357 );
and ( w_20357 , w_20354 , w_20355 );
buf ( w_20354 , \5755_b1 );
not ( w_20354 , w_20358 );
not ( w_20355 , w_20359 );
and ( w_20358 , w_20359 , \5755_b0 );
or ( \8140_b1 , \8135_b1 , \8139_b1 );
xor ( \8140_b0 , \8135_b0 , w_20360 );
not ( w_20360 , w_20361 );
and ( w_20361 , \8139_b1 , \8139_b0 );
or ( \8141_b1 , \6041_b1 , \5768_b1 );
not ( \5768_b1 , w_20362 );
and ( \8141_b0 , \6041_b0 , w_20363 );
and ( w_20362 , w_20363 , \5768_b0 );
or ( \8142_b1 , \6006_b1 , \5766_b1 );
not ( \5766_b1 , w_20364 );
and ( \8142_b0 , \6006_b0 , w_20365 );
and ( w_20364 , w_20365 , \5766_b0 );
or ( \8143_b1 , \8141_b1 , w_20367 );
not ( w_20367 , w_20368 );
and ( \8143_b0 , \8141_b0 , w_20369 );
and ( w_20368 ,  , w_20369 );
buf ( w_20367 , \8142_b1 );
not ( w_20367 , w_20370 );
not (  , w_20371 );
and ( w_20370 , w_20371 , \8142_b0 );
or ( \8144_b1 , \8143_b1 , w_20372 );
xor ( \8144_b0 , \8143_b0 , w_20374 );
not ( w_20374 , w_20375 );
and ( w_20375 , w_20372 , w_20373 );
buf ( w_20372 , \5775_b1 );
not ( w_20372 , w_20376 );
not ( w_20373 , w_20377 );
and ( w_20376 , w_20377 , \5775_b0 );
or ( \8145_b1 , \8140_b1 , \8144_b1 );
xor ( \8145_b0 , \8140_b0 , w_20378 );
not ( w_20378 , w_20379 );
and ( w_20379 , \8144_b1 , \8144_b0 );
or ( \8146_b1 , \8131_b1 , \8145_b1 );
xor ( \8146_b0 , \8131_b0 , w_20380 );
not ( w_20380 , w_20381 );
and ( w_20381 , \8145_b1 , \8145_b0 );
or ( \8147_b1 , \5937_b1 , \7157_b1 );
not ( \7157_b1 , w_20382 );
and ( \8147_b0 , \5937_b0 , w_20383 );
and ( w_20382 , w_20383 , \7157_b0 );
or ( \8148_b1 , \5906_b1 , \7155_b1 );
not ( \7155_b1 , w_20384 );
and ( \8148_b0 , \5906_b0 , w_20385 );
and ( w_20384 , w_20385 , \7155_b0 );
or ( \8149_b1 , \8147_b1 , w_20387 );
not ( w_20387 , w_20388 );
and ( \8149_b0 , \8147_b0 , w_20389 );
and ( w_20388 ,  , w_20389 );
buf ( w_20387 , \8148_b1 );
not ( w_20387 , w_20390 );
not (  , w_20391 );
and ( w_20390 , w_20391 , \8148_b0 );
or ( \8150_b1 , \8149_b1 , w_20392 );
xor ( \8150_b0 , \8149_b0 , w_20394 );
not ( w_20394 , w_20395 );
and ( w_20395 , w_20392 , w_20393 );
buf ( w_20392 , \7163_b1 );
not ( w_20392 , w_20396 );
not ( w_20393 , w_20397 );
and ( w_20396 , w_20397 , \7163_b0 );
or ( \8151_b1 , \5957_b1 , \7175_b1 );
not ( \7175_b1 , w_20398 );
and ( \8151_b0 , \5957_b0 , w_20399 );
and ( w_20398 , w_20399 , \7175_b0 );
or ( \8152_b1 , \5925_b1 , \7173_b1 );
not ( \7173_b1 , w_20400 );
and ( \8152_b0 , \5925_b0 , w_20401 );
and ( w_20400 , w_20401 , \7173_b0 );
or ( \8153_b1 , \8151_b1 , w_20403 );
not ( w_20403 , w_20404 );
and ( \8153_b0 , \8151_b0 , w_20405 );
and ( w_20404 ,  , w_20405 );
buf ( w_20403 , \8152_b1 );
not ( w_20403 , w_20406 );
not (  , w_20407 );
and ( w_20406 , w_20407 , \8152_b0 );
or ( \8154_b1 , \8153_b1 , w_20408 );
xor ( \8154_b0 , \8153_b0 , w_20410 );
not ( w_20410 , w_20411 );
and ( w_20411 , w_20408 , w_20409 );
buf ( w_20408 , \7181_b1 );
not ( w_20408 , w_20412 );
not ( w_20409 , w_20413 );
and ( w_20412 , w_20413 , \7181_b0 );
or ( \8155_b1 , \8150_b1 , \8154_b1 );
xor ( \8155_b0 , \8150_b0 , w_20414 );
not ( w_20414 , w_20415 );
and ( w_20415 , \8154_b1 , \8154_b0 );
or ( \8156_b1 , \5979_b1 , \7192_b1 );
not ( \7192_b1 , w_20416 );
and ( \8156_b0 , \5979_b0 , w_20417 );
and ( w_20416 , w_20417 , \7192_b0 );
or ( \8157_b1 , \5945_b1 , \7190_b1 );
not ( \7190_b1 , w_20418 );
and ( \8157_b0 , \5945_b0 , w_20419 );
and ( w_20418 , w_20419 , \7190_b0 );
or ( \8158_b1 , \8156_b1 , w_20421 );
not ( w_20421 , w_20422 );
and ( \8158_b0 , \8156_b0 , w_20423 );
and ( w_20422 ,  , w_20423 );
buf ( w_20421 , \8157_b1 );
not ( w_20421 , w_20424 );
not (  , w_20425 );
and ( w_20424 , w_20425 , \8157_b0 );
or ( \8159_b1 , \8158_b1 , w_20426 );
xor ( \8159_b0 , \8158_b0 , w_20428 );
not ( w_20428 , w_20429 );
and ( w_20429 , w_20426 , w_20427 );
buf ( w_20426 , \7198_b1 );
not ( w_20426 , w_20430 );
not ( w_20427 , w_20431 );
and ( w_20430 , w_20431 , \7198_b0 );
or ( \8160_b1 , \8155_b1 , \8159_b1 );
xor ( \8160_b0 , \8155_b0 , w_20432 );
not ( w_20432 , w_20433 );
and ( w_20433 , \8159_b1 , \8159_b0 );
or ( \8161_b1 , \8146_b1 , \8160_b1 );
xor ( \8161_b0 , \8146_b0 , w_20434 );
not ( w_20434 , w_20435 );
and ( w_20435 , \8160_b1 , \8160_b0 );
or ( \8162_b1 , \8122_b1 , \8161_b1 );
xor ( \8162_b0 , \8122_b0 , w_20436 );
not ( w_20436 , w_20437 );
and ( w_20437 , \8161_b1 , \8161_b0 );
or ( \8163_b1 , \7991_b1 , \7995_b1 );
not ( \7995_b1 , w_20438 );
and ( \8163_b0 , \7991_b0 , w_20439 );
and ( w_20438 , w_20439 , \7995_b0 );
or ( \8164_b1 , \7995_b1 , \8000_b1 );
not ( \8000_b1 , w_20440 );
and ( \8164_b0 , \7995_b0 , w_20441 );
and ( w_20440 , w_20441 , \8000_b0 );
or ( \8165_b1 , \7991_b1 , \8000_b1 );
not ( \8000_b1 , w_20442 );
and ( \8165_b0 , \7991_b0 , w_20443 );
and ( w_20442 , w_20443 , \8000_b0 );
or ( \8167_b1 , \7977_b1 , \7981_b1 );
not ( \7981_b1 , w_20444 );
and ( \8167_b0 , \7977_b0 , w_20445 );
and ( w_20444 , w_20445 , \7981_b0 );
or ( \8168_b1 , \7981_b1 , \7986_b1 );
not ( \7986_b1 , w_20446 );
and ( \8168_b0 , \7981_b0 , w_20447 );
and ( w_20446 , w_20447 , \7986_b0 );
or ( \8169_b1 , \7977_b1 , \7986_b1 );
not ( \7986_b1 , w_20448 );
and ( \8169_b0 , \7977_b0 , w_20449 );
and ( w_20448 , w_20449 , \7986_b0 );
or ( \8171_b1 , \8166_b1 , \8170_b1 );
xor ( \8171_b0 , \8166_b0 , w_20450 );
not ( w_20450 , w_20451 );
and ( w_20451 , \8170_b1 , \8170_b0 );
or ( \8172_b1 , \7925_b1 , \7929_b1 );
not ( \7929_b1 , w_20452 );
and ( \8172_b0 , \7925_b0 , w_20453 );
and ( w_20452 , w_20453 , \7929_b0 );
or ( \8173_b1 , \7929_b1 , \7932_b1 );
not ( \7932_b1 , w_20454 );
and ( \8173_b0 , \7929_b0 , w_20455 );
and ( w_20454 , w_20455 , \7932_b0 );
or ( \8174_b1 , \7925_b1 , \7932_b1 );
not ( \7932_b1 , w_20456 );
and ( \8174_b0 , \7925_b0 , w_20457 );
and ( w_20456 , w_20457 , \7932_b0 );
or ( \8176_b1 , \8171_b1 , \8175_b1 );
xor ( \8176_b0 , \8171_b0 , w_20458 );
not ( w_20458 , w_20459 );
and ( w_20459 , \8175_b1 , \8175_b0 );
or ( \8177_b1 , \8162_b1 , \8176_b1 );
xor ( \8177_b0 , \8162_b0 , w_20460 );
not ( w_20460 , w_20461 );
and ( w_20461 , \8176_b1 , \8176_b0 );
or ( \8178_b1 , \8081_b1 , \8177_b1 );
xor ( \8178_b0 , \8081_b0 , w_20462 );
not ( w_20462 , w_20463 );
and ( w_20463 , \8177_b1 , \8177_b0 );
or ( \8179_b1 , \7938_b1 , \7942_b1 );
not ( \7942_b1 , w_20464 );
and ( \8179_b0 , \7938_b0 , w_20465 );
and ( w_20464 , w_20465 , \7942_b0 );
or ( \8180_b1 , \7942_b1 , \7947_b1 );
not ( \7947_b1 , w_20466 );
and ( \8180_b0 , \7942_b0 , w_20467 );
and ( w_20466 , w_20467 , \7947_b0 );
or ( \8181_b1 , \7938_b1 , \7947_b1 );
not ( \7947_b1 , w_20468 );
and ( \8181_b0 , \7938_b0 , w_20469 );
and ( w_20468 , w_20469 , \7947_b0 );
or ( \8183_b1 , \7916_b1 , \7920_b1 );
not ( \7920_b1 , w_20470 );
and ( \8183_b0 , \7916_b0 , w_20471 );
and ( w_20470 , w_20471 , \7920_b0 );
or ( \8184_b1 , \7920_b1 , \7933_b1 );
not ( \7933_b1 , w_20472 );
and ( \8184_b0 , \7920_b0 , w_20473 );
and ( w_20472 , w_20473 , \7933_b0 );
or ( \8185_b1 , \7916_b1 , \7933_b1 );
not ( \7933_b1 , w_20474 );
and ( \8185_b0 , \7916_b0 , w_20475 );
and ( w_20474 , w_20475 , \7933_b0 );
or ( \8187_b1 , \8182_b1 , \8186_b1 );
xor ( \8187_b0 , \8182_b0 , w_20476 );
not ( w_20476 , w_20477 );
and ( w_20477 , \8186_b1 , \8186_b0 );
or ( \8188_b1 , \7987_b1 , \8001_b1 );
not ( \8001_b1 , w_20478 );
and ( \8188_b0 , \7987_b0 , w_20479 );
and ( w_20478 , w_20479 , \8001_b0 );
or ( \8189_b1 , \8001_b1 , \8016_b1 );
not ( \8016_b1 , w_20480 );
and ( \8189_b0 , \8001_b0 , w_20481 );
and ( w_20480 , w_20481 , \8016_b0 );
or ( \8190_b1 , \7987_b1 , \8016_b1 );
not ( \8016_b1 , w_20482 );
and ( \8190_b0 , \7987_b0 , w_20483 );
and ( w_20482 , w_20483 , \8016_b0 );
or ( \8192_b1 , \8187_b1 , \8191_b1 );
xor ( \8192_b0 , \8187_b0 , w_20484 );
not ( w_20484 , w_20485 );
and ( w_20485 , \8191_b1 , \8191_b0 );
or ( \8193_b1 , \8178_b1 , \8192_b1 );
xor ( \8193_b0 , \8178_b0 , w_20486 );
not ( w_20486 , w_20487 );
and ( w_20487 , \8192_b1 , \8192_b0 );
or ( \8194_b1 , \8067_b1 , \8193_b1 );
xor ( \8194_b0 , \8067_b0 , w_20488 );
not ( w_20488 , w_20489 );
and ( w_20489 , \8193_b1 , \8193_b0 );
or ( \8195_b1 , \8058_b1 , \8194_b1 );
xor ( \8195_b0 , \8058_b0 , w_20490 );
not ( w_20490 , w_20491 );
and ( w_20491 , \8194_b1 , \8194_b0 );
or ( \8196_b1 , \7891_b1 , \7905_b1 );
not ( \7905_b1 , w_20492 );
and ( \8196_b0 , \7891_b0 , w_20493 );
and ( w_20492 , w_20493 , \7905_b0 );
or ( \8197_b1 , \7905_b1 , \8035_b1 );
not ( \8035_b1 , w_20494 );
and ( \8197_b0 , \7905_b0 , w_20495 );
and ( w_20494 , w_20495 , \8035_b0 );
or ( \8198_b1 , \7891_b1 , \8035_b1 );
not ( \8035_b1 , w_20496 );
and ( \8198_b0 , \7891_b0 , w_20497 );
and ( w_20496 , w_20497 , \8035_b0 );
or ( \8200_b1 , \8195_b1 , w_20499 );
not ( w_20499 , w_20500 );
and ( \8200_b0 , \8195_b0 , w_20501 );
and ( w_20500 ,  , w_20501 );
buf ( w_20499 , \8199_b1 );
not ( w_20499 , w_20502 );
not (  , w_20503 );
and ( w_20502 , w_20503 , \8199_b0 );
or ( \8201_b1 , \8062_b1 , \8066_b1 );
not ( \8066_b1 , w_20504 );
and ( \8201_b0 , \8062_b0 , w_20505 );
and ( w_20504 , w_20505 , \8066_b0 );
or ( \8202_b1 , \8066_b1 , \8193_b1 );
not ( \8193_b1 , w_20506 );
and ( \8202_b0 , \8066_b0 , w_20507 );
and ( w_20506 , w_20507 , \8193_b0 );
or ( \8203_b1 , \8062_b1 , \8193_b1 );
not ( \8193_b1 , w_20508 );
and ( \8203_b0 , \8062_b0 , w_20509 );
and ( w_20508 , w_20509 , \8193_b0 );
or ( \8205_b1 , \8071_b1 , \8075_b1 );
not ( \8075_b1 , w_20510 );
and ( \8205_b0 , \8071_b0 , w_20511 );
and ( w_20510 , w_20511 , \8075_b0 );
or ( \8206_b1 , \8075_b1 , \8080_b1 );
not ( \8080_b1 , w_20512 );
and ( \8206_b0 , \8075_b0 , w_20513 );
and ( w_20512 , w_20513 , \8080_b0 );
or ( \8207_b1 , \8071_b1 , \8080_b1 );
not ( \8080_b1 , w_20514 );
and ( \8207_b0 , \8071_b0 , w_20515 );
and ( w_20514 , w_20515 , \8080_b0 );
or ( \8209_b1 , \8166_b1 , \8170_b1 );
not ( \8170_b1 , w_20516 );
and ( \8209_b0 , \8166_b0 , w_20517 );
and ( w_20516 , w_20517 , \8170_b0 );
or ( \8210_b1 , \8170_b1 , \8175_b1 );
not ( \8175_b1 , w_20518 );
and ( \8210_b0 , \8170_b0 , w_20519 );
and ( w_20518 , w_20519 , \8175_b0 );
or ( \8211_b1 , \8166_b1 , \8175_b1 );
not ( \8175_b1 , w_20520 );
and ( \8211_b0 , \8166_b0 , w_20521 );
and ( w_20520 , w_20521 , \8175_b0 );
or ( \8213_b1 , \8208_b1 , \8212_b1 );
xor ( \8213_b0 , \8208_b0 , w_20522 );
not ( w_20522 , w_20523 );
and ( w_20523 , \8212_b1 , \8212_b0 );
or ( \8214_b1 , \8131_b1 , \8145_b1 );
not ( \8145_b1 , w_20524 );
and ( \8214_b0 , \8131_b0 , w_20525 );
and ( w_20524 , w_20525 , \8145_b0 );
or ( \8215_b1 , \8145_b1 , \8160_b1 );
not ( \8160_b1 , w_20526 );
and ( \8215_b0 , \8145_b0 , w_20527 );
and ( w_20526 , w_20527 , \8160_b0 );
or ( \8216_b1 , \8131_b1 , \8160_b1 );
not ( \8160_b1 , w_20528 );
and ( \8216_b0 , \8131_b0 , w_20529 );
and ( w_20528 , w_20529 , \8160_b0 );
or ( \8218_b1 , \8213_b1 , \8217_b1 );
xor ( \8218_b0 , \8213_b0 , w_20530 );
not ( w_20530 , w_20531 );
and ( w_20531 , \8217_b1 , \8217_b0 );
or ( \8219_b1 , \8182_b1 , \8186_b1 );
not ( \8186_b1 , w_20532 );
and ( \8219_b0 , \8182_b0 , w_20533 );
and ( w_20532 , w_20533 , \8186_b0 );
or ( \8220_b1 , \8186_b1 , \8191_b1 );
not ( \8191_b1 , w_20534 );
and ( \8220_b0 , \8186_b0 , w_20535 );
and ( w_20534 , w_20535 , \8191_b0 );
or ( \8221_b1 , \8182_b1 , \8191_b1 );
not ( \8191_b1 , w_20536 );
and ( \8221_b0 , \8182_b0 , w_20537 );
and ( w_20536 , w_20537 , \8191_b0 );
or ( \8223_b1 , \8122_b1 , \8161_b1 );
not ( \8161_b1 , w_20538 );
and ( \8223_b0 , \8122_b0 , w_20539 );
and ( w_20538 , w_20539 , \8161_b0 );
or ( \8224_b1 , \8161_b1 , \8176_b1 );
not ( \8176_b1 , w_20540 );
and ( \8224_b0 , \8161_b0 , w_20541 );
and ( w_20540 , w_20541 , \8176_b0 );
or ( \8225_b1 , \8122_b1 , \8176_b1 );
not ( \8176_b1 , w_20542 );
and ( \8225_b0 , \8122_b0 , w_20543 );
and ( w_20542 , w_20543 , \8176_b0 );
or ( \8227_b1 , \8222_b1 , \8226_b1 );
xor ( \8227_b0 , \8222_b0 , w_20544 );
not ( w_20544 , w_20545 );
and ( w_20545 , \8226_b1 , \8226_b0 );
or ( \8228_b1 , \6029_b1 , \5790_b1 );
not ( \5790_b1 , w_20546 );
and ( \8228_b0 , \6029_b0 , w_20547 );
and ( w_20546 , w_20547 , \5790_b0 );
or ( \8229_b1 , \6041_b1 , \5788_b1 );
not ( \5788_b1 , w_20548 );
and ( \8229_b0 , \6041_b0 , w_20549 );
and ( w_20548 , w_20549 , \5788_b0 );
or ( \8230_b1 , \8228_b1 , w_20551 );
not ( w_20551 , w_20552 );
and ( \8230_b0 , \8228_b0 , w_20553 );
and ( w_20552 ,  , w_20553 );
buf ( w_20551 , \8229_b1 );
not ( w_20551 , w_20554 );
not (  , w_20555 );
and ( w_20554 , w_20555 , \8229_b0 );
or ( \8231_b1 , \8230_b1 , w_20556 );
xor ( \8231_b0 , \8230_b0 , w_20558 );
not ( w_20558 , w_20559 );
and ( w_20559 , w_20556 , w_20557 );
buf ( w_20556 , \5797_b1 );
not ( w_20556 , w_20560 );
not ( w_20557 , w_20561 );
and ( w_20560 , w_20561 , \5797_b0 );
or ( \8232_b1 , \6048_b1 , \5809_b1 );
not ( \5809_b1 , w_20562 );
and ( \8232_b0 , \6048_b0 , w_20563 );
and ( w_20562 , w_20563 , \5809_b0 );
or ( \8233_b1 , \6057_b1 , \5807_b1 );
not ( \5807_b1 , w_20564 );
and ( \8233_b0 , \6057_b0 , w_20565 );
and ( w_20564 , w_20565 , \5807_b0 );
or ( \8234_b1 , \8232_b1 , w_20567 );
not ( w_20567 , w_20568 );
and ( \8234_b0 , \8232_b0 , w_20569 );
and ( w_20568 ,  , w_20569 );
buf ( w_20567 , \8233_b1 );
not ( w_20567 , w_20570 );
not (  , w_20571 );
and ( w_20570 , w_20571 , \8233_b0 );
or ( \8235_b1 , \8234_b1 , w_20572 );
xor ( \8235_b0 , \8234_b0 , w_20574 );
not ( w_20574 , w_20575 );
and ( w_20575 , w_20572 , w_20573 );
buf ( w_20572 , \5816_b1 );
not ( w_20572 , w_20576 );
not ( w_20573 , w_20577 );
and ( w_20576 , w_20577 , \5816_b0 );
or ( \8236_b1 , \8231_b1 , \8235_b1 );
xor ( \8236_b0 , \8231_b0 , w_20578 );
not ( w_20578 , w_20579 );
and ( w_20579 , \8235_b1 , \8235_b0 );
or ( \8237_b1 , \6065_b1 , w_20581 );
not ( w_20581 , w_20582 );
and ( \8237_b0 , \6065_b0 , w_20583 );
and ( w_20582 ,  , w_20583 );
buf ( w_20581 , \5827_b1 );
not ( w_20581 , w_20584 );
not (  , w_20585 );
and ( w_20584 , w_20585 , \5827_b0 );
or ( \8238_b1 , \8237_b1 , w_20586 );
xor ( \8238_b0 , \8237_b0 , w_20588 );
not ( w_20588 , w_20589 );
and ( w_20589 , w_20586 , w_20587 );
buf ( w_20586 , \5836_b1 );
not ( w_20586 , w_20590 );
not ( w_20587 , w_20591 );
and ( w_20590 , w_20591 , \5836_b0 );
or ( \8239_b1 , \8236_b1 , \8238_b1 );
xor ( \8239_b0 , \8236_b0 , w_20592 );
not ( w_20592 , w_20593 );
and ( w_20593 , \8238_b1 , \8238_b0 );
or ( \8240_b1 , \5967_b1 , \7203_b1 );
not ( \7203_b1 , w_20594 );
and ( \8240_b0 , \5967_b0 , w_20595 );
and ( w_20594 , w_20595 , \7203_b0 );
or ( \8241_b1 , \5979_b1 , \7201_b1 );
not ( \7201_b1 , w_20596 );
and ( \8241_b0 , \5979_b0 , w_20597 );
and ( w_20596 , w_20597 , \7201_b0 );
or ( \8242_b1 , \8240_b1 , w_20599 );
not ( w_20599 , w_20600 );
and ( \8242_b0 , \8240_b0 , w_20601 );
and ( w_20600 ,  , w_20601 );
buf ( w_20599 , \8241_b1 );
not ( w_20599 , w_20602 );
not (  , w_20603 );
and ( w_20602 , w_20603 , \8241_b0 );
or ( \8243_b1 , \8242_b1 , w_20604 );
xor ( \8243_b0 , \8242_b0 , w_20606 );
not ( w_20606 , w_20607 );
and ( w_20607 , w_20604 , w_20605 );
buf ( w_20604 , \6824_b1 );
not ( w_20604 , w_20608 );
not ( w_20605 , w_20609 );
and ( w_20608 , w_20609 , \6824_b0 );
or ( \8244_b1 , \5986_b1 , \5750_b1 );
not ( \5750_b1 , w_20610 );
and ( \8244_b0 , \5986_b0 , w_20611 );
and ( w_20610 , w_20611 , \5750_b0 );
or ( \8245_b1 , \5998_b1 , \5748_b1 );
not ( \5748_b1 , w_20612 );
and ( \8245_b0 , \5998_b0 , w_20613 );
and ( w_20612 , w_20613 , \5748_b0 );
or ( \8246_b1 , \8244_b1 , w_20615 );
not ( w_20615 , w_20616 );
and ( \8246_b0 , \8244_b0 , w_20617 );
and ( w_20616 ,  , w_20617 );
buf ( w_20615 , \8245_b1 );
not ( w_20615 , w_20618 );
not (  , w_20619 );
and ( w_20618 , w_20619 , \8245_b0 );
or ( \8247_b1 , \8246_b1 , w_20620 );
xor ( \8247_b0 , \8246_b0 , w_20622 );
not ( w_20622 , w_20623 );
and ( w_20623 , w_20620 , w_20621 );
buf ( w_20620 , \5755_b1 );
not ( w_20620 , w_20624 );
not ( w_20621 , w_20625 );
and ( w_20624 , w_20625 , \5755_b0 );
or ( \8248_b1 , \8243_b1 , \8247_b1 );
xor ( \8248_b0 , \8243_b0 , w_20626 );
not ( w_20626 , w_20627 );
and ( w_20627 , \8247_b1 , \8247_b0 );
or ( \8249_b1 , \6006_b1 , \5768_b1 );
not ( \5768_b1 , w_20628 );
and ( \8249_b0 , \6006_b0 , w_20629 );
and ( w_20628 , w_20629 , \5768_b0 );
or ( \8250_b1 , \6018_b1 , \5766_b1 );
not ( \5766_b1 , w_20630 );
and ( \8250_b0 , \6018_b0 , w_20631 );
and ( w_20630 , w_20631 , \5766_b0 );
or ( \8251_b1 , \8249_b1 , w_20633 );
not ( w_20633 , w_20634 );
and ( \8251_b0 , \8249_b0 , w_20635 );
and ( w_20634 ,  , w_20635 );
buf ( w_20633 , \8250_b1 );
not ( w_20633 , w_20636 );
not (  , w_20637 );
and ( w_20636 , w_20637 , \8250_b0 );
or ( \8252_b1 , \8251_b1 , w_20638 );
xor ( \8252_b0 , \8251_b0 , w_20640 );
not ( w_20640 , w_20641 );
and ( w_20641 , w_20638 , w_20639 );
buf ( w_20638 , \5775_b1 );
not ( w_20638 , w_20642 );
not ( w_20639 , w_20643 );
and ( w_20642 , w_20643 , \5775_b0 );
or ( \8253_b1 , \8248_b1 , \8252_b1 );
xor ( \8253_b0 , \8248_b0 , w_20644 );
not ( w_20644 , w_20645 );
and ( w_20645 , \8252_b1 , \8252_b0 );
or ( \8254_b1 , \8239_b1 , w_20646 );
xor ( \8254_b0 , \8239_b0 , w_20648 );
not ( w_20648 , w_20649 );
and ( w_20649 , w_20646 , w_20647 );
buf ( w_20646 , \8253_b1 );
not ( w_20646 , w_20650 );
not ( w_20647 , w_20651 );
and ( w_20650 , w_20651 , \8253_b0 );
or ( \8255_b1 , \8150_b1 , \8154_b1 );
not ( \8154_b1 , w_20652 );
and ( \8255_b0 , \8150_b0 , w_20653 );
and ( w_20652 , w_20653 , \8154_b0 );
or ( \8256_b1 , \8154_b1 , \8159_b1 );
not ( \8159_b1 , w_20654 );
and ( \8256_b0 , \8154_b0 , w_20655 );
and ( w_20654 , w_20655 , \8159_b0 );
or ( \8257_b1 , \8150_b1 , \8159_b1 );
not ( \8159_b1 , w_20656 );
and ( \8257_b0 , \8150_b0 , w_20657 );
and ( w_20656 , w_20657 , \8159_b0 );
or ( \8259_b1 , \8135_b1 , \8139_b1 );
not ( \8139_b1 , w_20658 );
and ( \8259_b0 , \8135_b0 , w_20659 );
and ( w_20658 , w_20659 , \8139_b0 );
or ( \8260_b1 , \8139_b1 , \8144_b1 );
not ( \8144_b1 , w_20660 );
and ( \8260_b0 , \8139_b0 , w_20661 );
and ( w_20660 , w_20661 , \8144_b0 );
or ( \8261_b1 , \8135_b1 , \8144_b1 );
not ( \8144_b1 , w_20662 );
and ( \8261_b0 , \8135_b0 , w_20663 );
and ( w_20662 , w_20663 , \8144_b0 );
or ( \8263_b1 , \8258_b1 , \8262_b1 );
xor ( \8263_b0 , \8258_b0 , w_20664 );
not ( w_20664 , w_20665 );
and ( w_20665 , \8262_b1 , \8262_b0 );
or ( \8264_b1 , \8126_b1 , w_20666 );
or ( \8264_b0 , \8126_b0 , \8130_b0 );
not ( \8130_b0 , w_20667 );
and ( w_20667 , w_20666 , \8130_b1 );
or ( \8265_b1 , \8263_b1 , \8264_b1 );
xor ( \8265_b0 , \8263_b0 , w_20668 );
not ( w_20668 , w_20669 );
and ( w_20669 , \8264_b1 , \8264_b0 );
or ( \8266_b1 , \8254_b1 , \8265_b1 );
xor ( \8266_b0 , \8254_b0 , w_20670 );
not ( w_20670 , w_20671 );
and ( w_20671 , \8265_b1 , \8265_b0 );
or ( \8267_b1 , \8111_b1 , \8115_b1 );
not ( \8115_b1 , w_20672 );
and ( \8267_b0 , \8111_b0 , w_20673 );
and ( w_20672 , w_20673 , \8115_b0 );
or ( \8268_b1 , \8115_b1 , \8120_b1 );
not ( \8120_b1 , w_20674 );
and ( \8268_b0 , \8115_b0 , w_20675 );
and ( w_20674 , w_20675 , \8120_b0 );
or ( \8269_b1 , \8111_b1 , \8120_b1 );
not ( \8120_b1 , w_20676 );
and ( \8269_b0 , \8111_b0 , w_20677 );
and ( w_20676 , w_20677 , \8120_b0 );
or ( \8271_b1 , \8099_b1 , \8103_b1 );
not ( \8103_b1 , w_20678 );
and ( \8271_b0 , \8099_b0 , w_20679 );
and ( w_20678 , w_20679 , \8103_b0 );
or ( \8272_b1 , \8103_b1 , \8108_b1 );
not ( \8108_b1 , w_20680 );
and ( \8272_b0 , \8103_b0 , w_20681 );
and ( w_20680 , w_20681 , \8108_b0 );
or ( \8273_b1 , \8099_b1 , \8108_b1 );
not ( \8108_b1 , w_20682 );
and ( \8273_b0 , \8099_b0 , w_20683 );
and ( w_20682 , w_20683 , \8108_b0 );
or ( \8275_b1 , \8270_b1 , \8274_b1 );
xor ( \8275_b0 , \8270_b0 , w_20684 );
not ( w_20684 , w_20685 );
and ( w_20685 , \8274_b1 , \8274_b0 );
or ( \8276_b1 , \8085_b1 , \8089_b1 );
not ( \8089_b1 , w_20686 );
and ( \8276_b0 , \8085_b0 , w_20687 );
and ( w_20686 , w_20687 , \8089_b0 );
or ( \8277_b1 , \8089_b1 , \8094_b1 );
not ( \8094_b1 , w_20688 );
and ( \8277_b0 , \8089_b0 , w_20689 );
and ( w_20688 , w_20689 , \8094_b0 );
or ( \8278_b1 , \8085_b1 , \8094_b1 );
not ( \8094_b1 , w_20690 );
and ( \8278_b0 , \8085_b0 , w_20691 );
and ( w_20690 , w_20691 , \8094_b0 );
or ( \8280_b1 , \8275_b1 , \8279_b1 );
xor ( \8280_b0 , \8275_b0 , w_20692 );
not ( w_20692 , w_20693 );
and ( w_20693 , \8279_b1 , \8279_b0 );
or ( \8281_b1 , \8266_b1 , \8280_b1 );
xor ( \8281_b0 , \8266_b0 , w_20694 );
not ( w_20694 , w_20695 );
and ( w_20695 , \8280_b1 , \8280_b0 );
or ( \8282_b1 , \8227_b1 , \8281_b1 );
xor ( \8282_b0 , \8227_b0 , w_20696 );
not ( w_20696 , w_20697 );
and ( w_20697 , \8281_b1 , \8281_b0 );
or ( \8283_b1 , \8218_b1 , \8282_b1 );
xor ( \8283_b0 , \8218_b0 , w_20698 );
not ( w_20698 , w_20699 );
and ( w_20699 , \8282_b1 , \8282_b0 );
or ( \8284_b1 , \8204_b1 , \8283_b1 );
xor ( \8284_b0 , \8204_b0 , w_20700 );
not ( w_20700 , w_20701 );
and ( w_20701 , \8283_b1 , \8283_b0 );
or ( \8285_b1 , \8050_b1 , \8054_b1 );
not ( \8054_b1 , w_20702 );
and ( \8285_b0 , \8050_b0 , w_20703 );
and ( w_20702 , w_20703 , \8054_b0 );
or ( \8286_b1 , \8054_b1 , \8056_b1 );
not ( \8056_b1 , w_20704 );
and ( \8286_b0 , \8054_b0 , w_20705 );
and ( w_20704 , w_20705 , \8056_b0 );
or ( \8287_b1 , \8050_b1 , \8056_b1 );
not ( \8056_b1 , w_20706 );
and ( \8287_b0 , \8050_b0 , w_20707 );
and ( w_20706 , w_20707 , \8056_b0 );
or ( \8289_b1 , \8081_b1 , \8177_b1 );
not ( \8177_b1 , w_20708 );
and ( \8289_b0 , \8081_b0 , w_20709 );
and ( w_20708 , w_20709 , \8177_b0 );
or ( \8290_b1 , \8177_b1 , \8192_b1 );
not ( \8192_b1 , w_20710 );
and ( \8290_b0 , \8177_b0 , w_20711 );
and ( w_20710 , w_20711 , \8192_b0 );
or ( \8291_b1 , \8081_b1 , \8192_b1 );
not ( \8192_b1 , w_20712 );
and ( \8291_b0 , \8081_b0 , w_20713 );
and ( w_20712 , w_20713 , \8192_b0 );
or ( \8293_b1 , \8288_b1 , \8292_b1 );
xor ( \8293_b0 , \8288_b0 , w_20714 );
not ( w_20714 , w_20715 );
and ( w_20715 , \8292_b1 , \8292_b0 );
or ( \8294_b1 , \8095_b1 , \8109_b1 );
not ( \8109_b1 , w_20716 );
and ( \8294_b0 , \8095_b0 , w_20717 );
and ( w_20716 , w_20717 , \8109_b0 );
or ( \8295_b1 , \8109_b1 , \8121_b1 );
not ( \8121_b1 , w_20718 );
and ( \8295_b0 , \8109_b0 , w_20719 );
and ( w_20718 , w_20719 , \8121_b0 );
or ( \8296_b1 , \8095_b1 , \8121_b1 );
not ( \8121_b1 , w_20720 );
and ( \8296_b0 , \8095_b0 , w_20721 );
and ( w_20720 , w_20721 , \8121_b0 );
or ( \8298_b1 , \5737_b1 , \7006_b1 );
not ( \7006_b1 , w_20722 );
and ( \8298_b0 , \5737_b0 , w_20723 );
and ( w_20722 , w_20723 , \7006_b0 );
buf ( \8299_b1 , \8298_b1 );
not ( \8299_b1 , w_20724 );
not ( \8299_b0 , w_20725 );
and ( w_20724 , w_20725 , \8298_b0 );
or ( \8300_b1 , \8299_b1 , w_20726 );
xor ( \8300_b0 , \8299_b0 , w_20728 );
not ( w_20728 , w_20729 );
and ( w_20729 , w_20726 , w_20727 );
buf ( w_20726 , \7012_b1 );
not ( w_20726 , w_20730 );
not ( w_20727 , w_20731 );
and ( w_20730 , w_20731 , \7012_b0 );
or ( \8301_b1 , \5836_b1 , \8300_b1 );
xor ( \8301_b0 , \5836_b0 , w_20732 );
not ( w_20732 , w_20733 );
and ( w_20733 , \8300_b1 , \8300_b0 );
or ( \8302_b1 , \5758_b1 , \7026_b1 );
not ( \7026_b1 , w_20734 );
and ( \8302_b0 , \5758_b0 , w_20735 );
and ( w_20734 , w_20735 , \7026_b0 );
or ( \8303_b1 , \5770_b1 , \7024_b1 );
not ( \7024_b1 , w_20736 );
and ( \8303_b0 , \5770_b0 , w_20737 );
and ( w_20736 , w_20737 , \7024_b0 );
or ( \8304_b1 , \8302_b1 , w_20739 );
not ( w_20739 , w_20740 );
and ( \8304_b0 , \8302_b0 , w_20741 );
and ( w_20740 ,  , w_20741 );
buf ( w_20739 , \8303_b1 );
not ( w_20739 , w_20742 );
not (  , w_20743 );
and ( w_20742 , w_20743 , \8303_b0 );
or ( \8305_b1 , \8304_b1 , w_20744 );
xor ( \8305_b0 , \8304_b0 , w_20746 );
not ( w_20746 , w_20747 );
and ( w_20747 , w_20744 , w_20745 );
buf ( w_20744 , \7032_b1 );
not ( w_20744 , w_20748 );
not ( w_20745 , w_20749 );
and ( w_20748 , w_20749 , \7032_b0 );
or ( \8306_b1 , \8301_b1 , \8305_b1 );
xor ( \8306_b0 , \8301_b0 , w_20750 );
not ( w_20750 , w_20751 );
and ( w_20751 , \8305_b1 , \8305_b0 );
or ( \8307_b1 , \8297_b1 , \8306_b1 );
xor ( \8307_b0 , \8297_b0 , w_20752 );
not ( w_20752 , w_20753 );
and ( w_20753 , \8306_b1 , \8306_b0 );
or ( \8308_b1 , \5906_b1 , \7157_b1 );
not ( \7157_b1 , w_20754 );
and ( \8308_b0 , \5906_b0 , w_20755 );
and ( w_20754 , w_20755 , \7157_b0 );
or ( \8309_b1 , \5918_b1 , \7155_b1 );
not ( \7155_b1 , w_20756 );
and ( \8309_b0 , \5918_b0 , w_20757 );
and ( w_20756 , w_20757 , \7155_b0 );
or ( \8310_b1 , \8308_b1 , w_20759 );
not ( w_20759 , w_20760 );
and ( \8310_b0 , \8308_b0 , w_20761 );
and ( w_20760 ,  , w_20761 );
buf ( w_20759 , \8309_b1 );
not ( w_20759 , w_20762 );
not (  , w_20763 );
and ( w_20762 , w_20763 , \8309_b0 );
or ( \8311_b1 , \8310_b1 , w_20764 );
xor ( \8311_b0 , \8310_b0 , w_20766 );
not ( w_20766 , w_20767 );
and ( w_20767 , w_20764 , w_20765 );
buf ( w_20764 , \7163_b1 );
not ( w_20764 , w_20768 );
not ( w_20765 , w_20769 );
and ( w_20768 , w_20769 , \7163_b0 );
or ( \8312_b1 , \5925_b1 , \7175_b1 );
not ( \7175_b1 , w_20770 );
and ( \8312_b0 , \5925_b0 , w_20771 );
and ( w_20770 , w_20771 , \7175_b0 );
or ( \8313_b1 , \5937_b1 , \7173_b1 );
not ( \7173_b1 , w_20772 );
and ( \8313_b0 , \5937_b0 , w_20773 );
and ( w_20772 , w_20773 , \7173_b0 );
or ( \8314_b1 , \8312_b1 , w_20775 );
not ( w_20775 , w_20776 );
and ( \8314_b0 , \8312_b0 , w_20777 );
and ( w_20776 ,  , w_20777 );
buf ( w_20775 , \8313_b1 );
not ( w_20775 , w_20778 );
not (  , w_20779 );
and ( w_20778 , w_20779 , \8313_b0 );
or ( \8315_b1 , \8314_b1 , w_20780 );
xor ( \8315_b0 , \8314_b0 , w_20782 );
not ( w_20782 , w_20783 );
and ( w_20783 , w_20780 , w_20781 );
buf ( w_20780 , \7181_b1 );
not ( w_20780 , w_20784 );
not ( w_20781 , w_20785 );
and ( w_20784 , w_20785 , \7181_b0 );
or ( \8316_b1 , \8311_b1 , \8315_b1 );
xor ( \8316_b0 , \8311_b0 , w_20786 );
not ( w_20786 , w_20787 );
and ( w_20787 , \8315_b1 , \8315_b0 );
or ( \8317_b1 , \5945_b1 , \7192_b1 );
not ( \7192_b1 , w_20788 );
and ( \8317_b0 , \5945_b0 , w_20789 );
and ( w_20788 , w_20789 , \7192_b0 );
or ( \8318_b1 , \5957_b1 , \7190_b1 );
not ( \7190_b1 , w_20790 );
and ( \8318_b0 , \5957_b0 , w_20791 );
and ( w_20790 , w_20791 , \7190_b0 );
or ( \8319_b1 , \8317_b1 , w_20793 );
not ( w_20793 , w_20794 );
and ( \8319_b0 , \8317_b0 , w_20795 );
and ( w_20794 ,  , w_20795 );
buf ( w_20793 , \8318_b1 );
not ( w_20793 , w_20796 );
not (  , w_20797 );
and ( w_20796 , w_20797 , \8318_b0 );
or ( \8320_b1 , \8319_b1 , w_20798 );
xor ( \8320_b0 , \8319_b0 , w_20800 );
not ( w_20800 , w_20801 );
and ( w_20801 , w_20798 , w_20799 );
buf ( w_20798 , \7198_b1 );
not ( w_20798 , w_20802 );
not ( w_20799 , w_20803 );
and ( w_20802 , w_20803 , \7198_b0 );
or ( \8321_b1 , \8316_b1 , \8320_b1 );
xor ( \8321_b0 , \8316_b0 , w_20804 );
not ( w_20804 , w_20805 );
and ( w_20805 , \8320_b1 , \8320_b0 );
or ( \8322_b1 , \5842_b1 , \7099_b1 );
not ( \7099_b1 , w_20806 );
and ( \8322_b0 , \5842_b0 , w_20807 );
and ( w_20806 , w_20807 , \7099_b0 );
or ( \8323_b1 , \5854_b1 , \7097_b1 );
not ( \7097_b1 , w_20808 );
and ( \8323_b0 , \5854_b0 , w_20809 );
and ( w_20808 , w_20809 , \7097_b0 );
or ( \8324_b1 , \8322_b1 , w_20811 );
not ( w_20811 , w_20812 );
and ( \8324_b0 , \8322_b0 , w_20813 );
and ( w_20812 ,  , w_20813 );
buf ( w_20811 , \8323_b1 );
not ( w_20811 , w_20814 );
not (  , w_20815 );
and ( w_20814 , w_20815 , \8323_b0 );
or ( \8325_b1 , \8324_b1 , w_20816 );
xor ( \8325_b0 , \8324_b0 , w_20818 );
not ( w_20818 , w_20819 );
and ( w_20819 , w_20816 , w_20817 );
buf ( w_20816 , \7105_b1 );
not ( w_20816 , w_20820 );
not ( w_20817 , w_20821 );
and ( w_20820 , w_20821 , \7105_b0 );
or ( \8326_b1 , \5861_b1 , \7117_b1 );
not ( \7117_b1 , w_20822 );
and ( \8326_b0 , \5861_b0 , w_20823 );
and ( w_20822 , w_20823 , \7117_b0 );
or ( \8327_b1 , \5873_b1 , \7115_b1 );
not ( \7115_b1 , w_20824 );
and ( \8327_b0 , \5873_b0 , w_20825 );
and ( w_20824 , w_20825 , \7115_b0 );
or ( \8328_b1 , \8326_b1 , w_20827 );
not ( w_20827 , w_20828 );
and ( \8328_b0 , \8326_b0 , w_20829 );
and ( w_20828 ,  , w_20829 );
buf ( w_20827 , \8327_b1 );
not ( w_20827 , w_20830 );
not (  , w_20831 );
and ( w_20830 , w_20831 , \8327_b0 );
or ( \8329_b1 , \8328_b1 , w_20832 );
xor ( \8329_b0 , \8328_b0 , w_20834 );
not ( w_20834 , w_20835 );
and ( w_20835 , w_20832 , w_20833 );
buf ( w_20832 , \7123_b1 );
not ( w_20832 , w_20836 );
not ( w_20833 , w_20837 );
and ( w_20836 , w_20837 , \7123_b0 );
or ( \8330_b1 , \8325_b1 , \8329_b1 );
xor ( \8330_b0 , \8325_b0 , w_20838 );
not ( w_20838 , w_20839 );
and ( w_20839 , \8329_b1 , \8329_b0 );
or ( \8331_b1 , \5881_b1 , \7140_b1 );
not ( \7140_b1 , w_20840 );
and ( \8331_b0 , \5881_b0 , w_20841 );
and ( w_20840 , w_20841 , \7140_b0 );
or ( \8332_b1 , \5893_b1 , \7138_b1 );
not ( \7138_b1 , w_20842 );
and ( \8332_b0 , \5893_b0 , w_20843 );
and ( w_20842 , w_20843 , \7138_b0 );
or ( \8333_b1 , \8331_b1 , w_20845 );
not ( w_20845 , w_20846 );
and ( \8333_b0 , \8331_b0 , w_20847 );
and ( w_20846 ,  , w_20847 );
buf ( w_20845 , \8332_b1 );
not ( w_20845 , w_20848 );
not (  , w_20849 );
and ( w_20848 , w_20849 , \8332_b0 );
or ( \8334_b1 , \8333_b1 , w_20850 );
xor ( \8334_b0 , \8333_b0 , w_20852 );
not ( w_20852 , w_20853 );
and ( w_20853 , w_20850 , w_20851 );
buf ( w_20850 , \7146_b1 );
not ( w_20850 , w_20854 );
not ( w_20851 , w_20855 );
and ( w_20854 , w_20855 , \7146_b0 );
or ( \8335_b1 , \8330_b1 , \8334_b1 );
xor ( \8335_b0 , \8330_b0 , w_20856 );
not ( w_20856 , w_20857 );
and ( w_20857 , \8334_b1 , \8334_b0 );
or ( \8336_b1 , \8321_b1 , \8335_b1 );
xor ( \8336_b0 , \8321_b0 , w_20858 );
not ( w_20858 , w_20859 );
and ( w_20859 , \8335_b1 , \8335_b0 );
or ( \8337_b1 , \5780_b1 , \7043_b1 );
not ( \7043_b1 , w_20860 );
and ( \8337_b0 , \5780_b0 , w_20861 );
and ( w_20860 , w_20861 , \7043_b0 );
or ( \8338_b1 , \5792_b1 , \7041_b1 );
not ( \7041_b1 , w_20862 );
and ( \8338_b0 , \5792_b0 , w_20863 );
and ( w_20862 , w_20863 , \7041_b0 );
or ( \8339_b1 , \8337_b1 , w_20865 );
not ( w_20865 , w_20866 );
and ( \8339_b0 , \8337_b0 , w_20867 );
and ( w_20866 ,  , w_20867 );
buf ( w_20865 , \8338_b1 );
not ( w_20865 , w_20868 );
not (  , w_20869 );
and ( w_20868 , w_20869 , \8338_b0 );
or ( \8340_b1 , \8339_b1 , w_20870 );
xor ( \8340_b0 , \8339_b0 , w_20872 );
not ( w_20872 , w_20873 );
and ( w_20873 , w_20870 , w_20871 );
buf ( w_20870 , \7049_b1 );
not ( w_20870 , w_20874 );
not ( w_20871 , w_20875 );
and ( w_20874 , w_20875 , \7049_b0 );
or ( \8341_b1 , \5799_b1 , \7061_b1 );
not ( \7061_b1 , w_20876 );
and ( \8341_b0 , \5799_b0 , w_20877 );
and ( w_20876 , w_20877 , \7061_b0 );
or ( \8342_b1 , \5811_b1 , \7059_b1 );
not ( \7059_b1 , w_20878 );
and ( \8342_b0 , \5811_b0 , w_20879 );
and ( w_20878 , w_20879 , \7059_b0 );
or ( \8343_b1 , \8341_b1 , w_20881 );
not ( w_20881 , w_20882 );
and ( \8343_b0 , \8341_b0 , w_20883 );
and ( w_20882 ,  , w_20883 );
buf ( w_20881 , \8342_b1 );
not ( w_20881 , w_20884 );
not (  , w_20885 );
and ( w_20884 , w_20885 , \8342_b0 );
or ( \8344_b1 , \8343_b1 , w_20886 );
xor ( \8344_b0 , \8343_b0 , w_20888 );
not ( w_20888 , w_20889 );
and ( w_20889 , w_20886 , w_20887 );
buf ( w_20886 , \7067_b1 );
not ( w_20886 , w_20890 );
not ( w_20887 , w_20891 );
and ( w_20890 , w_20891 , \7067_b0 );
or ( \8345_b1 , \8340_b1 , \8344_b1 );
xor ( \8345_b0 , \8340_b0 , w_20892 );
not ( w_20892 , w_20893 );
and ( w_20893 , \8344_b1 , \8344_b0 );
or ( \8346_b1 , \5819_b1 , \7082_b1 );
not ( \7082_b1 , w_20894 );
and ( \8346_b0 , \5819_b0 , w_20895 );
and ( w_20894 , w_20895 , \7082_b0 );
or ( \8347_b1 , \5831_b1 , \7080_b1 );
not ( \7080_b1 , w_20896 );
and ( \8347_b0 , \5831_b0 , w_20897 );
and ( w_20896 , w_20897 , \7080_b0 );
or ( \8348_b1 , \8346_b1 , w_20899 );
not ( w_20899 , w_20900 );
and ( \8348_b0 , \8346_b0 , w_20901 );
and ( w_20900 ,  , w_20901 );
buf ( w_20899 , \8347_b1 );
not ( w_20899 , w_20902 );
not (  , w_20903 );
and ( w_20902 , w_20903 , \8347_b0 );
or ( \8349_b1 , \8348_b1 , w_20904 );
xor ( \8349_b0 , \8348_b0 , w_20906 );
not ( w_20906 , w_20907 );
and ( w_20907 , w_20904 , w_20905 );
buf ( w_20904 , \7088_b1 );
not ( w_20904 , w_20908 );
not ( w_20905 , w_20909 );
and ( w_20908 , w_20909 , \7088_b0 );
or ( \8350_b1 , \8345_b1 , \8349_b1 );
xor ( \8350_b0 , \8345_b0 , w_20910 );
not ( w_20910 , w_20911 );
and ( w_20911 , \8349_b1 , \8349_b0 );
or ( \8351_b1 , \8336_b1 , \8350_b1 );
xor ( \8351_b0 , \8336_b0 , w_20912 );
not ( w_20912 , w_20913 );
and ( w_20913 , \8350_b1 , \8350_b0 );
or ( \8352_b1 , \8307_b1 , \8351_b1 );
xor ( \8352_b0 , \8307_b0 , w_20914 );
not ( w_20914 , w_20915 );
and ( w_20915 , \8351_b1 , \8351_b0 );
or ( \8353_b1 , \8293_b1 , \8352_b1 );
xor ( \8353_b0 , \8293_b0 , w_20916 );
not ( w_20916 , w_20917 );
and ( w_20917 , \8352_b1 , \8352_b0 );
or ( \8354_b1 , \8284_b1 , \8353_b1 );
xor ( \8354_b0 , \8284_b0 , w_20918 );
not ( w_20918 , w_20919 );
and ( w_20919 , \8353_b1 , \8353_b0 );
or ( \8355_b1 , \8046_b1 , \8057_b1 );
not ( \8057_b1 , w_20920 );
and ( \8355_b0 , \8046_b0 , w_20921 );
and ( w_20920 , w_20921 , \8057_b0 );
or ( \8356_b1 , \8057_b1 , \8194_b1 );
not ( \8194_b1 , w_20922 );
and ( \8356_b0 , \8057_b0 , w_20923 );
and ( w_20922 , w_20923 , \8194_b0 );
or ( \8357_b1 , \8046_b1 , \8194_b1 );
not ( \8194_b1 , w_20924 );
and ( \8357_b0 , \8046_b0 , w_20925 );
and ( w_20924 , w_20925 , \8194_b0 );
or ( \8359_b1 , \8354_b1 , w_20927 );
not ( w_20927 , w_20928 );
and ( \8359_b0 , \8354_b0 , w_20929 );
and ( w_20928 ,  , w_20929 );
buf ( w_20927 , \8358_b1 );
not ( w_20927 , w_20930 );
not (  , w_20931 );
and ( w_20930 , w_20931 , \8358_b0 );
or ( \8360_b1 , \8200_b1 , w_20933 );
not ( w_20933 , w_20934 );
and ( \8360_b0 , \8200_b0 , w_20935 );
and ( w_20934 ,  , w_20935 );
buf ( w_20933 , \8359_b1 );
not ( w_20933 , w_20936 );
not (  , w_20937 );
and ( w_20936 , w_20937 , \8359_b0 );
or ( \8361_b1 , \8042_b1 , w_20939 );
not ( w_20939 , w_20940 );
and ( \8361_b0 , \8042_b0 , w_20941 );
and ( w_20940 ,  , w_20941 );
buf ( w_20939 , \8360_b1 );
not ( w_20939 , w_20942 );
not (  , w_20943 );
and ( w_20942 , w_20943 , \8360_b0 );
or ( \8362_b1 , \8288_b1 , \8292_b1 );
not ( \8292_b1 , w_20944 );
and ( \8362_b0 , \8288_b0 , w_20945 );
and ( w_20944 , w_20945 , \8292_b0 );
or ( \8363_b1 , \8292_b1 , \8352_b1 );
not ( \8352_b1 , w_20946 );
and ( \8363_b0 , \8292_b0 , w_20947 );
and ( w_20946 , w_20947 , \8352_b0 );
or ( \8364_b1 , \8288_b1 , \8352_b1 );
not ( \8352_b1 , w_20948 );
and ( \8364_b0 , \8288_b0 , w_20949 );
and ( w_20948 , w_20949 , \8352_b0 );
or ( \8366_b1 , \8218_b1 , \8282_b1 );
not ( \8282_b1 , w_20950 );
and ( \8366_b0 , \8218_b0 , w_20951 );
and ( w_20950 , w_20951 , \8282_b0 );
or ( \8367_b1 , \8365_b1 , \8366_b1 );
xor ( \8367_b0 , \8365_b0 , w_20952 );
not ( w_20952 , w_20953 );
and ( w_20953 , \8366_b1 , \8366_b0 );
or ( \8368_b1 , \8222_b1 , \8226_b1 );
not ( \8226_b1 , w_20954 );
and ( \8368_b0 , \8222_b0 , w_20955 );
and ( w_20954 , w_20955 , \8226_b0 );
or ( \8369_b1 , \8226_b1 , \8281_b1 );
not ( \8281_b1 , w_20956 );
and ( \8369_b0 , \8226_b0 , w_20957 );
and ( w_20956 , w_20957 , \8281_b0 );
or ( \8370_b1 , \8222_b1 , \8281_b1 );
not ( \8281_b1 , w_20958 );
and ( \8370_b0 , \8222_b0 , w_20959 );
and ( w_20958 , w_20959 , \8281_b0 );
or ( \8372_b1 , \8311_b1 , \8315_b1 );
not ( \8315_b1 , w_20960 );
and ( \8372_b0 , \8311_b0 , w_20961 );
and ( w_20960 , w_20961 , \8315_b0 );
or ( \8373_b1 , \8315_b1 , \8320_b1 );
not ( \8320_b1 , w_20962 );
and ( \8373_b0 , \8315_b0 , w_20963 );
and ( w_20962 , w_20963 , \8320_b0 );
or ( \8374_b1 , \8311_b1 , \8320_b1 );
not ( \8320_b1 , w_20964 );
and ( \8374_b0 , \8311_b0 , w_20965 );
and ( w_20964 , w_20965 , \8320_b0 );
or ( \8376_b1 , \8243_b1 , \8247_b1 );
not ( \8247_b1 , w_20966 );
and ( \8376_b0 , \8243_b0 , w_20967 );
and ( w_20966 , w_20967 , \8247_b0 );
or ( \8377_b1 , \8247_b1 , \8252_b1 );
not ( \8252_b1 , w_20968 );
and ( \8377_b0 , \8247_b0 , w_20969 );
and ( w_20968 , w_20969 , \8252_b0 );
or ( \8378_b1 , \8243_b1 , \8252_b1 );
not ( \8252_b1 , w_20970 );
and ( \8378_b0 , \8243_b0 , w_20971 );
and ( w_20970 , w_20971 , \8252_b0 );
or ( \8380_b1 , \8375_b1 , \8379_b1 );
xor ( \8380_b0 , \8375_b0 , w_20972 );
not ( w_20972 , w_20973 );
and ( w_20973 , \8379_b1 , \8379_b0 );
or ( \8381_b1 , \8231_b1 , \8235_b1 );
not ( \8235_b1 , w_20974 );
and ( \8381_b0 , \8231_b0 , w_20975 );
and ( w_20974 , w_20975 , \8235_b0 );
or ( \8382_b1 , \8235_b1 , \8238_b1 );
not ( \8238_b1 , w_20976 );
and ( \8382_b0 , \8235_b0 , w_20977 );
and ( w_20976 , w_20977 , \8238_b0 );
or ( \8383_b1 , \8231_b1 , \8238_b1 );
not ( \8238_b1 , w_20978 );
and ( \8383_b0 , \8231_b0 , w_20979 );
and ( w_20978 , w_20979 , \8238_b0 );
or ( \8385_b1 , \8380_b1 , \8384_b1 );
xor ( \8385_b0 , \8380_b0 , w_20980 );
not ( w_20980 , w_20981 );
and ( w_20981 , \8384_b1 , \8384_b0 );
or ( \8386_b1 , \5836_b1 , \8300_b1 );
not ( \8300_b1 , w_20982 );
and ( \8386_b0 , \5836_b0 , w_20983 );
and ( w_20982 , w_20983 , \8300_b0 );
or ( \8387_b1 , \8300_b1 , \8305_b1 );
not ( \8305_b1 , w_20984 );
and ( \8387_b0 , \8300_b0 , w_20985 );
and ( w_20984 , w_20985 , \8305_b0 );
or ( \8388_b1 , \5836_b1 , \8305_b1 );
not ( \8305_b1 , w_20986 );
and ( \8388_b0 , \5836_b0 , w_20987 );
and ( w_20986 , w_20987 , \8305_b0 );
or ( \8390_b1 , \8340_b1 , \8344_b1 );
not ( \8344_b1 , w_20988 );
and ( \8390_b0 , \8340_b0 , w_20989 );
and ( w_20988 , w_20989 , \8344_b0 );
or ( \8391_b1 , \8344_b1 , \8349_b1 );
not ( \8349_b1 , w_20990 );
and ( \8391_b0 , \8344_b0 , w_20991 );
and ( w_20990 , w_20991 , \8349_b0 );
or ( \8392_b1 , \8340_b1 , \8349_b1 );
not ( \8349_b1 , w_20992 );
and ( \8392_b0 , \8340_b0 , w_20993 );
and ( w_20992 , w_20993 , \8349_b0 );
or ( \8394_b1 , \8389_b1 , \8393_b1 );
xor ( \8394_b0 , \8389_b0 , w_20994 );
not ( w_20994 , w_20995 );
and ( w_20995 , \8393_b1 , \8393_b0 );
or ( \8395_b1 , \8325_b1 , \8329_b1 );
not ( \8329_b1 , w_20996 );
and ( \8395_b0 , \8325_b0 , w_20997 );
and ( w_20996 , w_20997 , \8329_b0 );
or ( \8396_b1 , \8329_b1 , \8334_b1 );
not ( \8334_b1 , w_20998 );
and ( \8396_b0 , \8329_b0 , w_20999 );
and ( w_20998 , w_20999 , \8334_b0 );
or ( \8397_b1 , \8325_b1 , \8334_b1 );
not ( \8334_b1 , w_21000 );
and ( \8397_b0 , \8325_b0 , w_21001 );
and ( w_21000 , w_21001 , \8334_b0 );
or ( \8399_b1 , \8394_b1 , \8398_b1 );
xor ( \8399_b0 , \8394_b0 , w_21002 );
not ( w_21002 , w_21003 );
and ( w_21003 , \8398_b1 , \8398_b0 );
or ( \8400_b1 , \8385_b1 , \8399_b1 );
xor ( \8400_b0 , \8385_b0 , w_21004 );
not ( w_21004 , w_21005 );
and ( w_21005 , \8399_b1 , \8399_b0 );
or ( \8401_b1 , \8321_b1 , \8335_b1 );
not ( \8335_b1 , w_21006 );
and ( \8401_b0 , \8321_b0 , w_21007 );
and ( w_21006 , w_21007 , \8335_b0 );
or ( \8402_b1 , \8335_b1 , \8350_b1 );
not ( \8350_b1 , w_21008 );
and ( \8402_b0 , \8335_b0 , w_21009 );
and ( w_21008 , w_21009 , \8350_b0 );
or ( \8403_b1 , \8321_b1 , \8350_b1 );
not ( \8350_b1 , w_21010 );
and ( \8403_b0 , \8321_b0 , w_21011 );
and ( w_21010 , w_21011 , \8350_b0 );
or ( \8405_b1 , \5873_b1 , \7117_b1 );
not ( \7117_b1 , w_21012 );
and ( \8405_b0 , \5873_b0 , w_21013 );
and ( w_21012 , w_21013 , \7117_b0 );
or ( \8406_b1 , \5842_b1 , \7115_b1 );
not ( \7115_b1 , w_21014 );
and ( \8406_b0 , \5842_b0 , w_21015 );
and ( w_21014 , w_21015 , \7115_b0 );
or ( \8407_b1 , \8405_b1 , w_21017 );
not ( w_21017 , w_21018 );
and ( \8407_b0 , \8405_b0 , w_21019 );
and ( w_21018 ,  , w_21019 );
buf ( w_21017 , \8406_b1 );
not ( w_21017 , w_21020 );
not (  , w_21021 );
and ( w_21020 , w_21021 , \8406_b0 );
or ( \8408_b1 , \8407_b1 , w_21022 );
xor ( \8408_b0 , \8407_b0 , w_21024 );
not ( w_21024 , w_21025 );
and ( w_21025 , w_21022 , w_21023 );
buf ( w_21022 , \7123_b1 );
not ( w_21022 , w_21026 );
not ( w_21023 , w_21027 );
and ( w_21026 , w_21027 , \7123_b0 );
or ( \8409_b1 , \5893_b1 , \7140_b1 );
not ( \7140_b1 , w_21028 );
and ( \8409_b0 , \5893_b0 , w_21029 );
and ( w_21028 , w_21029 , \7140_b0 );
or ( \8410_b1 , \5861_b1 , \7138_b1 );
not ( \7138_b1 , w_21030 );
and ( \8410_b0 , \5861_b0 , w_21031 );
and ( w_21030 , w_21031 , \7138_b0 );
or ( \8411_b1 , \8409_b1 , w_21033 );
not ( w_21033 , w_21034 );
and ( \8411_b0 , \8409_b0 , w_21035 );
and ( w_21034 ,  , w_21035 );
buf ( w_21033 , \8410_b1 );
not ( w_21033 , w_21036 );
not (  , w_21037 );
and ( w_21036 , w_21037 , \8410_b0 );
or ( \8412_b1 , \8411_b1 , w_21038 );
xor ( \8412_b0 , \8411_b0 , w_21040 );
not ( w_21040 , w_21041 );
and ( w_21041 , w_21038 , w_21039 );
buf ( w_21038 , \7146_b1 );
not ( w_21038 , w_21042 );
not ( w_21039 , w_21043 );
and ( w_21042 , w_21043 , \7146_b0 );
or ( \8413_b1 , \8408_b1 , \8412_b1 );
xor ( \8413_b0 , \8408_b0 , w_21044 );
not ( w_21044 , w_21045 );
and ( w_21045 , \8412_b1 , \8412_b0 );
or ( \8414_b1 , \5918_b1 , \7157_b1 );
not ( \7157_b1 , w_21046 );
and ( \8414_b0 , \5918_b0 , w_21047 );
and ( w_21046 , w_21047 , \7157_b0 );
or ( \8415_b1 , \5881_b1 , \7155_b1 );
not ( \7155_b1 , w_21048 );
and ( \8415_b0 , \5881_b0 , w_21049 );
and ( w_21048 , w_21049 , \7155_b0 );
or ( \8416_b1 , \8414_b1 , w_21051 );
not ( w_21051 , w_21052 );
and ( \8416_b0 , \8414_b0 , w_21053 );
and ( w_21052 ,  , w_21053 );
buf ( w_21051 , \8415_b1 );
not ( w_21051 , w_21054 );
not (  , w_21055 );
and ( w_21054 , w_21055 , \8415_b0 );
or ( \8417_b1 , \8416_b1 , w_21056 );
xor ( \8417_b0 , \8416_b0 , w_21058 );
not ( w_21058 , w_21059 );
and ( w_21059 , w_21056 , w_21057 );
buf ( w_21056 , \7163_b1 );
not ( w_21056 , w_21060 );
not ( w_21057 , w_21061 );
and ( w_21060 , w_21061 , \7163_b0 );
or ( \8418_b1 , \8413_b1 , \8417_b1 );
xor ( \8418_b0 , \8413_b0 , w_21062 );
not ( w_21062 , w_21063 );
and ( w_21063 , \8417_b1 , \8417_b0 );
or ( \8419_b1 , \5811_b1 , \7061_b1 );
not ( \7061_b1 , w_21064 );
and ( \8419_b0 , \5811_b0 , w_21065 );
and ( w_21064 , w_21065 , \7061_b0 );
or ( \8420_b1 , \5780_b1 , \7059_b1 );
not ( \7059_b1 , w_21066 );
and ( \8420_b0 , \5780_b0 , w_21067 );
and ( w_21066 , w_21067 , \7059_b0 );
or ( \8421_b1 , \8419_b1 , w_21069 );
not ( w_21069 , w_21070 );
and ( \8421_b0 , \8419_b0 , w_21071 );
and ( w_21070 ,  , w_21071 );
buf ( w_21069 , \8420_b1 );
not ( w_21069 , w_21072 );
not (  , w_21073 );
and ( w_21072 , w_21073 , \8420_b0 );
or ( \8422_b1 , \8421_b1 , w_21074 );
xor ( \8422_b0 , \8421_b0 , w_21076 );
not ( w_21076 , w_21077 );
and ( w_21077 , w_21074 , w_21075 );
buf ( w_21074 , \7067_b1 );
not ( w_21074 , w_21078 );
not ( w_21075 , w_21079 );
and ( w_21078 , w_21079 , \7067_b0 );
or ( \8423_b1 , \5831_b1 , \7082_b1 );
not ( \7082_b1 , w_21080 );
and ( \8423_b0 , \5831_b0 , w_21081 );
and ( w_21080 , w_21081 , \7082_b0 );
or ( \8424_b1 , \5799_b1 , \7080_b1 );
not ( \7080_b1 , w_21082 );
and ( \8424_b0 , \5799_b0 , w_21083 );
and ( w_21082 , w_21083 , \7080_b0 );
or ( \8425_b1 , \8423_b1 , w_21085 );
not ( w_21085 , w_21086 );
and ( \8425_b0 , \8423_b0 , w_21087 );
and ( w_21086 ,  , w_21087 );
buf ( w_21085 , \8424_b1 );
not ( w_21085 , w_21088 );
not (  , w_21089 );
and ( w_21088 , w_21089 , \8424_b0 );
or ( \8426_b1 , \8425_b1 , w_21090 );
xor ( \8426_b0 , \8425_b0 , w_21092 );
not ( w_21092 , w_21093 );
and ( w_21093 , w_21090 , w_21091 );
buf ( w_21090 , \7088_b1 );
not ( w_21090 , w_21094 );
not ( w_21091 , w_21095 );
and ( w_21094 , w_21095 , \7088_b0 );
or ( \8427_b1 , \8422_b1 , \8426_b1 );
xor ( \8427_b0 , \8422_b0 , w_21096 );
not ( w_21096 , w_21097 );
and ( w_21097 , \8426_b1 , \8426_b0 );
or ( \8428_b1 , \5854_b1 , \7099_b1 );
not ( \7099_b1 , w_21098 );
and ( \8428_b0 , \5854_b0 , w_21099 );
and ( w_21098 , w_21099 , \7099_b0 );
or ( \8429_b1 , \5819_b1 , \7097_b1 );
not ( \7097_b1 , w_21100 );
and ( \8429_b0 , \5819_b0 , w_21101 );
and ( w_21100 , w_21101 , \7097_b0 );
or ( \8430_b1 , \8428_b1 , w_21103 );
not ( w_21103 , w_21104 );
and ( \8430_b0 , \8428_b0 , w_21105 );
and ( w_21104 ,  , w_21105 );
buf ( w_21103 , \8429_b1 );
not ( w_21103 , w_21106 );
not (  , w_21107 );
and ( w_21106 , w_21107 , \8429_b0 );
or ( \8431_b1 , \8430_b1 , w_21108 );
xor ( \8431_b0 , \8430_b0 , w_21110 );
not ( w_21110 , w_21111 );
and ( w_21111 , w_21108 , w_21109 );
buf ( w_21108 , \7105_b1 );
not ( w_21108 , w_21112 );
not ( w_21109 , w_21113 );
and ( w_21112 , w_21113 , \7105_b0 );
or ( \8432_b1 , \8427_b1 , \8431_b1 );
xor ( \8432_b0 , \8427_b0 , w_21114 );
not ( w_21114 , w_21115 );
and ( w_21115 , \8431_b1 , \8431_b0 );
or ( \8433_b1 , \8418_b1 , \8432_b1 );
xor ( \8433_b0 , \8418_b0 , w_21116 );
not ( w_21116 , w_21117 );
and ( w_21117 , \8432_b1 , \8432_b0 );
buf ( \8434_b1 , \7012_b1 );
not ( \8434_b1 , w_21118 );
not ( \8434_b0 , w_21119 );
and ( w_21118 , w_21119 , \7012_b0 );
or ( \8435_b1 , \5770_b1 , \7026_b1 );
not ( \7026_b1 , w_21120 );
and ( \8435_b0 , \5770_b0 , w_21121 );
and ( w_21120 , w_21121 , \7026_b0 );
or ( \8436_b1 , \5737_b1 , \7024_b1 );
not ( \7024_b1 , w_21122 );
and ( \8436_b0 , \5737_b0 , w_21123 );
and ( w_21122 , w_21123 , \7024_b0 );
or ( \8437_b1 , \8435_b1 , w_21125 );
not ( w_21125 , w_21126 );
and ( \8437_b0 , \8435_b0 , w_21127 );
and ( w_21126 ,  , w_21127 );
buf ( w_21125 , \8436_b1 );
not ( w_21125 , w_21128 );
not (  , w_21129 );
and ( w_21128 , w_21129 , \8436_b0 );
or ( \8438_b1 , \8437_b1 , w_21130 );
xor ( \8438_b0 , \8437_b0 , w_21132 );
not ( w_21132 , w_21133 );
and ( w_21133 , w_21130 , w_21131 );
buf ( w_21130 , \7032_b1 );
not ( w_21130 , w_21134 );
not ( w_21131 , w_21135 );
and ( w_21134 , w_21135 , \7032_b0 );
or ( \8439_b1 , \8434_b1 , \8438_b1 );
xor ( \8439_b0 , \8434_b0 , w_21136 );
not ( w_21136 , w_21137 );
and ( w_21137 , \8438_b1 , \8438_b0 );
or ( \8440_b1 , \5792_b1 , \7043_b1 );
not ( \7043_b1 , w_21138 );
and ( \8440_b0 , \5792_b0 , w_21139 );
and ( w_21138 , w_21139 , \7043_b0 );
or ( \8441_b1 , \5758_b1 , \7041_b1 );
not ( \7041_b1 , w_21140 );
and ( \8441_b0 , \5758_b0 , w_21141 );
and ( w_21140 , w_21141 , \7041_b0 );
or ( \8442_b1 , \8440_b1 , w_21143 );
not ( w_21143 , w_21144 );
and ( \8442_b0 , \8440_b0 , w_21145 );
and ( w_21144 ,  , w_21145 );
buf ( w_21143 , \8441_b1 );
not ( w_21143 , w_21146 );
not (  , w_21147 );
and ( w_21146 , w_21147 , \8441_b0 );
or ( \8443_b1 , \8442_b1 , w_21148 );
xor ( \8443_b0 , \8442_b0 , w_21150 );
not ( w_21150 , w_21151 );
and ( w_21151 , w_21148 , w_21149 );
buf ( w_21148 , \7049_b1 );
not ( w_21148 , w_21152 );
not ( w_21149 , w_21153 );
and ( w_21152 , w_21153 , \7049_b0 );
or ( \8444_b1 , \8439_b1 , \8443_b1 );
xor ( \8444_b0 , \8439_b0 , w_21154 );
not ( w_21154 , w_21155 );
and ( w_21155 , \8443_b1 , \8443_b0 );
or ( \8445_b1 , \8433_b1 , \8444_b1 );
xor ( \8445_b0 , \8433_b0 , w_21156 );
not ( w_21156 , w_21157 );
and ( w_21157 , \8444_b1 , \8444_b0 );
or ( \8446_b1 , \8404_b1 , \8445_b1 );
xor ( \8446_b0 , \8404_b0 , w_21158 );
not ( w_21158 , w_21159 );
and ( w_21159 , \8445_b1 , \8445_b0 );
or ( \8447_b1 , \6057_b1 , \5809_b1 );
not ( \5809_b1 , w_21160 );
and ( \8447_b0 , \6057_b0 , w_21161 );
and ( w_21160 , w_21161 , \5809_b0 );
or ( \8448_b1 , \6029_b1 , \5807_b1 );
not ( \5807_b1 , w_21162 );
and ( \8448_b0 , \6029_b0 , w_21163 );
and ( w_21162 , w_21163 , \5807_b0 );
or ( \8449_b1 , \8447_b1 , w_21165 );
not ( w_21165 , w_21166 );
and ( \8449_b0 , \8447_b0 , w_21167 );
and ( w_21166 ,  , w_21167 );
buf ( w_21165 , \8448_b1 );
not ( w_21165 , w_21168 );
not (  , w_21169 );
and ( w_21168 , w_21169 , \8448_b0 );
or ( \8450_b1 , \8449_b1 , w_21170 );
xor ( \8450_b0 , \8449_b0 , w_21172 );
not ( w_21172 , w_21173 );
and ( w_21173 , w_21170 , w_21171 );
buf ( w_21170 , \5816_b1 );
not ( w_21170 , w_21174 );
not ( w_21171 , w_21175 );
and ( w_21174 , w_21175 , \5816_b0 );
or ( \8451_b1 , \6065_b1 , \5829_b1 );
not ( \5829_b1 , w_21176 );
and ( \8451_b0 , \6065_b0 , w_21177 );
and ( w_21176 , w_21177 , \5829_b0 );
or ( \8452_b1 , \6048_b1 , \5827_b1 );
not ( \5827_b1 , w_21178 );
and ( \8452_b0 , \6048_b0 , w_21179 );
and ( w_21178 , w_21179 , \5827_b0 );
or ( \8453_b1 , \8451_b1 , w_21181 );
not ( w_21181 , w_21182 );
and ( \8453_b0 , \8451_b0 , w_21183 );
and ( w_21182 ,  , w_21183 );
buf ( w_21181 , \8452_b1 );
not ( w_21181 , w_21184 );
not (  , w_21185 );
and ( w_21184 , w_21185 , \8452_b0 );
or ( \8454_b1 , \8453_b1 , w_21186 );
xor ( \8454_b0 , \8453_b0 , w_21188 );
not ( w_21188 , w_21189 );
and ( w_21189 , w_21186 , w_21187 );
buf ( w_21186 , \5836_b1 );
not ( w_21186 , w_21190 );
not ( w_21187 , w_21191 );
and ( w_21190 , w_21191 , \5836_b0 );
or ( \8455_b1 , \8450_b1 , \8454_b1 );
xor ( \8455_b0 , \8450_b0 , w_21192 );
not ( w_21192 , w_21193 );
and ( w_21193 , \8454_b1 , \8454_b0 );
or ( \8456_b1 , \5998_b1 , \5750_b1 );
not ( \5750_b1 , w_21194 );
and ( \8456_b0 , \5998_b0 , w_21195 );
and ( w_21194 , w_21195 , \5750_b0 );
or ( \8457_b1 , \5967_b1 , \5748_b1 );
not ( \5748_b1 , w_21196 );
and ( \8457_b0 , \5967_b0 , w_21197 );
and ( w_21196 , w_21197 , \5748_b0 );
or ( \8458_b1 , \8456_b1 , w_21199 );
not ( w_21199 , w_21200 );
and ( \8458_b0 , \8456_b0 , w_21201 );
and ( w_21200 ,  , w_21201 );
buf ( w_21199 , \8457_b1 );
not ( w_21199 , w_21202 );
not (  , w_21203 );
and ( w_21202 , w_21203 , \8457_b0 );
or ( \8459_b1 , \8458_b1 , w_21204 );
xor ( \8459_b0 , \8458_b0 , w_21206 );
not ( w_21206 , w_21207 );
and ( w_21207 , w_21204 , w_21205 );
buf ( w_21204 , \5755_b1 );
not ( w_21204 , w_21208 );
not ( w_21205 , w_21209 );
and ( w_21208 , w_21209 , \5755_b0 );
or ( \8460_b1 , \6018_b1 , \5768_b1 );
not ( \5768_b1 , w_21210 );
and ( \8460_b0 , \6018_b0 , w_21211 );
and ( w_21210 , w_21211 , \5768_b0 );
or ( \8461_b1 , \5986_b1 , \5766_b1 );
not ( \5766_b1 , w_21212 );
and ( \8461_b0 , \5986_b0 , w_21213 );
and ( w_21212 , w_21213 , \5766_b0 );
or ( \8462_b1 , \8460_b1 , w_21215 );
not ( w_21215 , w_21216 );
and ( \8462_b0 , \8460_b0 , w_21217 );
and ( w_21216 ,  , w_21217 );
buf ( w_21215 , \8461_b1 );
not ( w_21215 , w_21218 );
not (  , w_21219 );
and ( w_21218 , w_21219 , \8461_b0 );
or ( \8463_b1 , \8462_b1 , w_21220 );
xor ( \8463_b0 , \8462_b0 , w_21222 );
not ( w_21222 , w_21223 );
and ( w_21223 , w_21220 , w_21221 );
buf ( w_21220 , \5775_b1 );
not ( w_21220 , w_21224 );
not ( w_21221 , w_21225 );
and ( w_21224 , w_21225 , \5775_b0 );
or ( \8464_b1 , \8459_b1 , \8463_b1 );
xor ( \8464_b0 , \8459_b0 , w_21226 );
not ( w_21226 , w_21227 );
and ( w_21227 , \8463_b1 , \8463_b0 );
or ( \8465_b1 , \6041_b1 , \5790_b1 );
not ( \5790_b1 , w_21228 );
and ( \8465_b0 , \6041_b0 , w_21229 );
and ( w_21228 , w_21229 , \5790_b0 );
or ( \8466_b1 , \6006_b1 , \5788_b1 );
not ( \5788_b1 , w_21230 );
and ( \8466_b0 , \6006_b0 , w_21231 );
and ( w_21230 , w_21231 , \5788_b0 );
or ( \8467_b1 , \8465_b1 , w_21233 );
not ( w_21233 , w_21234 );
and ( \8467_b0 , \8465_b0 , w_21235 );
and ( w_21234 ,  , w_21235 );
buf ( w_21233 , \8466_b1 );
not ( w_21233 , w_21236 );
not (  , w_21237 );
and ( w_21236 , w_21237 , \8466_b0 );
or ( \8468_b1 , \8467_b1 , w_21238 );
xor ( \8468_b0 , \8467_b0 , w_21240 );
not ( w_21240 , w_21241 );
and ( w_21241 , w_21238 , w_21239 );
buf ( w_21238 , \5797_b1 );
not ( w_21238 , w_21242 );
not ( w_21239 , w_21243 );
and ( w_21242 , w_21243 , \5797_b0 );
or ( \8469_b1 , \8464_b1 , \8468_b1 );
xor ( \8469_b0 , \8464_b0 , w_21244 );
not ( w_21244 , w_21245 );
and ( w_21245 , \8468_b1 , \8468_b0 );
or ( \8470_b1 , \8455_b1 , \8469_b1 );
xor ( \8470_b0 , \8455_b0 , w_21246 );
not ( w_21246 , w_21247 );
and ( w_21247 , \8469_b1 , \8469_b0 );
or ( \8471_b1 , \5937_b1 , \7175_b1 );
not ( \7175_b1 , w_21248 );
and ( \8471_b0 , \5937_b0 , w_21249 );
and ( w_21248 , w_21249 , \7175_b0 );
or ( \8472_b1 , \5906_b1 , \7173_b1 );
not ( \7173_b1 , w_21250 );
and ( \8472_b0 , \5906_b0 , w_21251 );
and ( w_21250 , w_21251 , \7173_b0 );
or ( \8473_b1 , \8471_b1 , w_21253 );
not ( w_21253 , w_21254 );
and ( \8473_b0 , \8471_b0 , w_21255 );
and ( w_21254 ,  , w_21255 );
buf ( w_21253 , \8472_b1 );
not ( w_21253 , w_21256 );
not (  , w_21257 );
and ( w_21256 , w_21257 , \8472_b0 );
or ( \8474_b1 , \8473_b1 , w_21258 );
xor ( \8474_b0 , \8473_b0 , w_21260 );
not ( w_21260 , w_21261 );
and ( w_21261 , w_21258 , w_21259 );
buf ( w_21258 , \7181_b1 );
not ( w_21258 , w_21262 );
not ( w_21259 , w_21263 );
and ( w_21262 , w_21263 , \7181_b0 );
or ( \8475_b1 , \5957_b1 , \7192_b1 );
not ( \7192_b1 , w_21264 );
and ( \8475_b0 , \5957_b0 , w_21265 );
and ( w_21264 , w_21265 , \7192_b0 );
or ( \8476_b1 , \5925_b1 , \7190_b1 );
not ( \7190_b1 , w_21266 );
and ( \8476_b0 , \5925_b0 , w_21267 );
and ( w_21266 , w_21267 , \7190_b0 );
or ( \8477_b1 , \8475_b1 , w_21269 );
not ( w_21269 , w_21270 );
and ( \8477_b0 , \8475_b0 , w_21271 );
and ( w_21270 ,  , w_21271 );
buf ( w_21269 , \8476_b1 );
not ( w_21269 , w_21272 );
not (  , w_21273 );
and ( w_21272 , w_21273 , \8476_b0 );
or ( \8478_b1 , \8477_b1 , w_21274 );
xor ( \8478_b0 , \8477_b0 , w_21276 );
not ( w_21276 , w_21277 );
and ( w_21277 , w_21274 , w_21275 );
buf ( w_21274 , \7198_b1 );
not ( w_21274 , w_21278 );
not ( w_21275 , w_21279 );
and ( w_21278 , w_21279 , \7198_b0 );
or ( \8479_b1 , \8474_b1 , \8478_b1 );
xor ( \8479_b0 , \8474_b0 , w_21280 );
not ( w_21280 , w_21281 );
and ( w_21281 , \8478_b1 , \8478_b0 );
or ( \8480_b1 , \5979_b1 , \7203_b1 );
not ( \7203_b1 , w_21282 );
and ( \8480_b0 , \5979_b0 , w_21283 );
and ( w_21282 , w_21283 , \7203_b0 );
or ( \8481_b1 , \5945_b1 , \7201_b1 );
not ( \7201_b1 , w_21284 );
and ( \8481_b0 , \5945_b0 , w_21285 );
and ( w_21284 , w_21285 , \7201_b0 );
or ( \8482_b1 , \8480_b1 , w_21287 );
not ( w_21287 , w_21288 );
and ( \8482_b0 , \8480_b0 , w_21289 );
and ( w_21288 ,  , w_21289 );
buf ( w_21287 , \8481_b1 );
not ( w_21287 , w_21290 );
not (  , w_21291 );
and ( w_21290 , w_21291 , \8481_b0 );
or ( \8483_b1 , \8482_b1 , w_21292 );
xor ( \8483_b0 , \8482_b0 , w_21294 );
not ( w_21294 , w_21295 );
and ( w_21295 , w_21292 , w_21293 );
buf ( w_21292 , \6824_b1 );
not ( w_21292 , w_21296 );
not ( w_21293 , w_21297 );
and ( w_21296 , w_21297 , \6824_b0 );
or ( \8484_b1 , \8479_b1 , \8483_b1 );
xor ( \8484_b0 , \8479_b0 , w_21298 );
not ( w_21298 , w_21299 );
and ( w_21299 , \8483_b1 , \8483_b0 );
or ( \8485_b1 , \8470_b1 , \8484_b1 );
xor ( \8485_b0 , \8470_b0 , w_21300 );
not ( w_21300 , w_21301 );
and ( w_21301 , \8484_b1 , \8484_b0 );
or ( \8486_b1 , \8446_b1 , \8485_b1 );
xor ( \8486_b0 , \8446_b0 , w_21302 );
not ( w_21302 , w_21303 );
and ( w_21303 , \8485_b1 , \8485_b0 );
or ( \8487_b1 , \8400_b1 , \8486_b1 );
xor ( \8487_b0 , \8400_b0 , w_21304 );
not ( w_21304 , w_21305 );
and ( w_21305 , \8486_b1 , \8486_b0 );
or ( \8488_b1 , \8270_b1 , \8274_b1 );
not ( \8274_b1 , w_21306 );
and ( \8488_b0 , \8270_b0 , w_21307 );
and ( w_21306 , w_21307 , \8274_b0 );
or ( \8489_b1 , \8274_b1 , \8279_b1 );
not ( \8279_b1 , w_21308 );
and ( \8489_b0 , \8274_b0 , w_21309 );
and ( w_21308 , w_21309 , \8279_b0 );
or ( \8490_b1 , \8270_b1 , \8279_b1 );
not ( \8279_b1 , w_21310 );
and ( \8490_b0 , \8270_b0 , w_21311 );
and ( w_21310 , w_21311 , \8279_b0 );
or ( \8492_b1 , \8258_b1 , \8262_b1 );
not ( \8262_b1 , w_21312 );
and ( \8492_b0 , \8258_b0 , w_21313 );
and ( w_21312 , w_21313 , \8262_b0 );
or ( \8493_b1 , \8262_b1 , \8264_b1 );
not ( \8264_b1 , w_21314 );
and ( \8493_b0 , \8262_b0 , w_21315 );
and ( w_21314 , w_21315 , \8264_b0 );
or ( \8494_b1 , \8258_b1 , \8264_b1 );
not ( \8264_b1 , w_21316 );
and ( \8494_b0 , \8258_b0 , w_21317 );
and ( w_21316 , w_21317 , \8264_b0 );
or ( \8496_b1 , \8491_b1 , \8495_b1 );
xor ( \8496_b0 , \8491_b0 , w_21318 );
not ( w_21318 , w_21319 );
and ( w_21319 , \8495_b1 , \8495_b0 );
or ( \8497_b1 , \8239_b1 , w_21320 );
or ( \8497_b0 , \8239_b0 , \8253_b0 );
not ( \8253_b0 , w_21321 );
and ( w_21321 , w_21320 , \8253_b1 );
or ( \8498_b1 , \8496_b1 , \8497_b1 );
xor ( \8498_b0 , \8496_b0 , w_21322 );
not ( w_21322 , w_21323 );
and ( w_21323 , \8497_b1 , \8497_b0 );
or ( \8499_b1 , \8487_b1 , \8498_b1 );
xor ( \8499_b0 , \8487_b0 , w_21324 );
not ( w_21324 , w_21325 );
and ( w_21325 , \8498_b1 , \8498_b0 );
or ( \8500_b1 , \8371_b1 , \8499_b1 );
xor ( \8500_b0 , \8371_b0 , w_21326 );
not ( w_21326 , w_21327 );
and ( w_21327 , \8499_b1 , \8499_b0 );
or ( \8501_b1 , \8208_b1 , \8212_b1 );
not ( \8212_b1 , w_21328 );
and ( \8501_b0 , \8208_b0 , w_21329 );
and ( w_21328 , w_21329 , \8212_b0 );
or ( \8502_b1 , \8212_b1 , \8217_b1 );
not ( \8217_b1 , w_21330 );
and ( \8502_b0 , \8212_b0 , w_21331 );
and ( w_21330 , w_21331 , \8217_b0 );
or ( \8503_b1 , \8208_b1 , \8217_b1 );
not ( \8217_b1 , w_21332 );
and ( \8503_b0 , \8208_b0 , w_21333 );
and ( w_21332 , w_21333 , \8217_b0 );
or ( \8505_b1 , \8297_b1 , \8306_b1 );
not ( \8306_b1 , w_21334 );
and ( \8505_b0 , \8297_b0 , w_21335 );
and ( w_21334 , w_21335 , \8306_b0 );
or ( \8506_b1 , \8306_b1 , \8351_b1 );
not ( \8351_b1 , w_21336 );
and ( \8506_b0 , \8306_b0 , w_21337 );
and ( w_21336 , w_21337 , \8351_b0 );
or ( \8507_b1 , \8297_b1 , \8351_b1 );
not ( \8351_b1 , w_21338 );
and ( \8507_b0 , \8297_b0 , w_21339 );
and ( w_21338 , w_21339 , \8351_b0 );
or ( \8509_b1 , \8504_b1 , \8508_b1 );
xor ( \8509_b0 , \8504_b0 , w_21340 );
not ( w_21340 , w_21341 );
and ( w_21341 , \8508_b1 , \8508_b0 );
or ( \8510_b1 , \8254_b1 , \8265_b1 );
not ( \8265_b1 , w_21342 );
and ( \8510_b0 , \8254_b0 , w_21343 );
and ( w_21342 , w_21343 , \8265_b0 );
or ( \8511_b1 , \8265_b1 , \8280_b1 );
not ( \8280_b1 , w_21344 );
and ( \8511_b0 , \8265_b0 , w_21345 );
and ( w_21344 , w_21345 , \8280_b0 );
or ( \8512_b1 , \8254_b1 , \8280_b1 );
not ( \8280_b1 , w_21346 );
and ( \8512_b0 , \8254_b0 , w_21347 );
and ( w_21346 , w_21347 , \8280_b0 );
or ( \8514_b1 , \8509_b1 , \8513_b1 );
xor ( \8514_b0 , \8509_b0 , w_21348 );
not ( w_21348 , w_21349 );
and ( w_21349 , \8513_b1 , \8513_b0 );
or ( \8515_b1 , \8500_b1 , \8514_b1 );
xor ( \8515_b0 , \8500_b0 , w_21350 );
not ( w_21350 , w_21351 );
and ( w_21351 , \8514_b1 , \8514_b0 );
or ( \8516_b1 , \8367_b1 , \8515_b1 );
xor ( \8516_b0 , \8367_b0 , w_21352 );
not ( w_21352 , w_21353 );
and ( w_21353 , \8515_b1 , \8515_b0 );
or ( \8517_b1 , \8204_b1 , \8283_b1 );
not ( \8283_b1 , w_21354 );
and ( \8517_b0 , \8204_b0 , w_21355 );
and ( w_21354 , w_21355 , \8283_b0 );
or ( \8518_b1 , \8283_b1 , \8353_b1 );
not ( \8353_b1 , w_21356 );
and ( \8518_b0 , \8283_b0 , w_21357 );
and ( w_21356 , w_21357 , \8353_b0 );
or ( \8519_b1 , \8204_b1 , \8353_b1 );
not ( \8353_b1 , w_21358 );
and ( \8519_b0 , \8204_b0 , w_21359 );
and ( w_21358 , w_21359 , \8353_b0 );
or ( \8521_b1 , \8516_b1 , w_21361 );
not ( w_21361 , w_21362 );
and ( \8521_b0 , \8516_b0 , w_21363 );
and ( w_21362 ,  , w_21363 );
buf ( w_21361 , \8520_b1 );
not ( w_21361 , w_21364 );
not (  , w_21365 );
and ( w_21364 , w_21365 , \8520_b0 );
or ( \8522_b1 , \8371_b1 , \8499_b1 );
not ( \8499_b1 , w_21366 );
and ( \8522_b0 , \8371_b0 , w_21367 );
and ( w_21366 , w_21367 , \8499_b0 );
or ( \8523_b1 , \8499_b1 , \8514_b1 );
not ( \8514_b1 , w_21368 );
and ( \8523_b0 , \8499_b0 , w_21369 );
and ( w_21368 , w_21369 , \8514_b0 );
or ( \8524_b1 , \8371_b1 , \8514_b1 );
not ( \8514_b1 , w_21370 );
and ( \8524_b0 , \8371_b0 , w_21371 );
and ( w_21370 , w_21371 , \8514_b0 );
or ( \8526_b1 , \8491_b1 , \8495_b1 );
not ( \8495_b1 , w_21372 );
and ( \8526_b0 , \8491_b0 , w_21373 );
and ( w_21372 , w_21373 , \8495_b0 );
or ( \8527_b1 , \8495_b1 , \8497_b1 );
not ( \8497_b1 , w_21374 );
and ( \8527_b0 , \8495_b0 , w_21375 );
and ( w_21374 , w_21375 , \8497_b0 );
or ( \8528_b1 , \8491_b1 , \8497_b1 );
not ( \8497_b1 , w_21376 );
and ( \8528_b0 , \8491_b0 , w_21377 );
and ( w_21376 , w_21377 , \8497_b0 );
or ( \8530_b1 , \8404_b1 , \8445_b1 );
not ( \8445_b1 , w_21378 );
and ( \8530_b0 , \8404_b0 , w_21379 );
and ( w_21378 , w_21379 , \8445_b0 );
or ( \8531_b1 , \8445_b1 , \8485_b1 );
not ( \8485_b1 , w_21380 );
and ( \8531_b0 , \8445_b0 , w_21381 );
and ( w_21380 , w_21381 , \8485_b0 );
or ( \8532_b1 , \8404_b1 , \8485_b1 );
not ( \8485_b1 , w_21382 );
and ( \8532_b0 , \8404_b0 , w_21383 );
and ( w_21382 , w_21383 , \8485_b0 );
or ( \8534_b1 , \8529_b1 , \8533_b1 );
xor ( \8534_b0 , \8529_b0 , w_21384 );
not ( w_21384 , w_21385 );
and ( w_21385 , \8533_b1 , \8533_b0 );
or ( \8535_b1 , \8385_b1 , \8399_b1 );
not ( \8399_b1 , w_21386 );
and ( \8535_b0 , \8385_b0 , w_21387 );
and ( w_21386 , w_21387 , \8399_b0 );
or ( \8536_b1 , \8534_b1 , \8535_b1 );
xor ( \8536_b0 , \8534_b0 , w_21388 );
not ( w_21388 , w_21389 );
and ( w_21389 , \8535_b1 , \8535_b0 );
or ( \8537_b1 , \8525_b1 , \8536_b1 );
xor ( \8537_b0 , \8525_b0 , w_21390 );
not ( w_21390 , w_21391 );
and ( w_21391 , \8536_b1 , \8536_b0 );
or ( \8538_b1 , \8504_b1 , \8508_b1 );
not ( \8508_b1 , w_21392 );
and ( \8538_b0 , \8504_b0 , w_21393 );
and ( w_21392 , w_21393 , \8508_b0 );
or ( \8539_b1 , \8508_b1 , \8513_b1 );
not ( \8513_b1 , w_21394 );
and ( \8539_b0 , \8508_b0 , w_21395 );
and ( w_21394 , w_21395 , \8513_b0 );
or ( \8540_b1 , \8504_b1 , \8513_b1 );
not ( \8513_b1 , w_21396 );
and ( \8540_b0 , \8504_b0 , w_21397 );
and ( w_21396 , w_21397 , \8513_b0 );
or ( \8542_b1 , \8400_b1 , \8486_b1 );
not ( \8486_b1 , w_21398 );
and ( \8542_b0 , \8400_b0 , w_21399 );
and ( w_21398 , w_21399 , \8486_b0 );
or ( \8543_b1 , \8486_b1 , \8498_b1 );
not ( \8498_b1 , w_21400 );
and ( \8543_b0 , \8486_b0 , w_21401 );
and ( w_21400 , w_21401 , \8498_b0 );
or ( \8544_b1 , \8400_b1 , \8498_b1 );
not ( \8498_b1 , w_21402 );
and ( \8544_b0 , \8400_b0 , w_21403 );
and ( w_21402 , w_21403 , \8498_b0 );
or ( \8546_b1 , \8541_b1 , \8545_b1 );
xor ( \8546_b0 , \8541_b0 , w_21404 );
not ( w_21404 , w_21405 );
and ( w_21405 , \8545_b1 , \8545_b0 );
or ( \8547_b1 , \6029_b1 , \5809_b1 );
not ( \5809_b1 , w_21406 );
and ( \8547_b0 , \6029_b0 , w_21407 );
and ( w_21406 , w_21407 , \5809_b0 );
or ( \8548_b1 , \6041_b1 , \5807_b1 );
not ( \5807_b1 , w_21408 );
and ( \8548_b0 , \6041_b0 , w_21409 );
and ( w_21408 , w_21409 , \5807_b0 );
or ( \8549_b1 , \8547_b1 , w_21411 );
not ( w_21411 , w_21412 );
and ( \8549_b0 , \8547_b0 , w_21413 );
and ( w_21412 ,  , w_21413 );
buf ( w_21411 , \8548_b1 );
not ( w_21411 , w_21414 );
not (  , w_21415 );
and ( w_21414 , w_21415 , \8548_b0 );
or ( \8550_b1 , \8549_b1 , w_21416 );
xor ( \8550_b0 , \8549_b0 , w_21418 );
not ( w_21418 , w_21419 );
and ( w_21419 , w_21416 , w_21417 );
buf ( w_21416 , \5816_b1 );
not ( w_21416 , w_21420 );
not ( w_21417 , w_21421 );
and ( w_21420 , w_21421 , \5816_b0 );
or ( \8551_b1 , \6048_b1 , \5829_b1 );
not ( \5829_b1 , w_21422 );
and ( \8551_b0 , \6048_b0 , w_21423 );
and ( w_21422 , w_21423 , \5829_b0 );
or ( \8552_b1 , \6057_b1 , \5827_b1 );
not ( \5827_b1 , w_21424 );
and ( \8552_b0 , \6057_b0 , w_21425 );
and ( w_21424 , w_21425 , \5827_b0 );
or ( \8553_b1 , \8551_b1 , w_21427 );
not ( w_21427 , w_21428 );
and ( \8553_b0 , \8551_b0 , w_21429 );
and ( w_21428 ,  , w_21429 );
buf ( w_21427 , \8552_b1 );
not ( w_21427 , w_21430 );
not (  , w_21431 );
and ( w_21430 , w_21431 , \8552_b0 );
or ( \8554_b1 , \8553_b1 , w_21432 );
xor ( \8554_b0 , \8553_b0 , w_21434 );
not ( w_21434 , w_21435 );
and ( w_21435 , w_21432 , w_21433 );
buf ( w_21432 , \5836_b1 );
not ( w_21432 , w_21436 );
not ( w_21433 , w_21437 );
and ( w_21436 , w_21437 , \5836_b0 );
or ( \8555_b1 , \8550_b1 , \8554_b1 );
xor ( \8555_b0 , \8550_b0 , w_21438 );
not ( w_21438 , w_21439 );
and ( w_21439 , \8554_b1 , \8554_b0 );
or ( \8556_b1 , \6065_b1 , w_21441 );
not ( w_21441 , w_21442 );
and ( \8556_b0 , \6065_b0 , w_21443 );
and ( w_21442 ,  , w_21443 );
buf ( w_21441 , \5850_b1 );
not ( w_21441 , w_21444 );
not (  , w_21445 );
and ( w_21444 , w_21445 , \5850_b0 );
or ( \8557_b1 , \8556_b1 , w_21446 );
xor ( \8557_b0 , \8556_b0 , w_21448 );
not ( w_21448 , w_21449 );
and ( w_21449 , w_21446 , w_21447 );
buf ( w_21446 , \5859_b1 );
not ( w_21446 , w_21450 );
not ( w_21447 , w_21451 );
and ( w_21450 , w_21451 , \5859_b0 );
or ( \8558_b1 , \8555_b1 , \8557_b1 );
xor ( \8558_b0 , \8555_b0 , w_21452 );
not ( w_21452 , w_21453 );
and ( w_21453 , \8557_b1 , \8557_b0 );
or ( \8559_b1 , \5967_b1 , \5750_b1 );
not ( \5750_b1 , w_21454 );
and ( \8559_b0 , \5967_b0 , w_21455 );
and ( w_21454 , w_21455 , \5750_b0 );
or ( \8560_b1 , \5979_b1 , \5748_b1 );
not ( \5748_b1 , w_21456 );
and ( \8560_b0 , \5979_b0 , w_21457 );
and ( w_21456 , w_21457 , \5748_b0 );
or ( \8561_b1 , \8559_b1 , w_21459 );
not ( w_21459 , w_21460 );
and ( \8561_b0 , \8559_b0 , w_21461 );
and ( w_21460 ,  , w_21461 );
buf ( w_21459 , \8560_b1 );
not ( w_21459 , w_21462 );
not (  , w_21463 );
and ( w_21462 , w_21463 , \8560_b0 );
or ( \8562_b1 , \8561_b1 , w_21464 );
xor ( \8562_b0 , \8561_b0 , w_21466 );
not ( w_21466 , w_21467 );
and ( w_21467 , w_21464 , w_21465 );
buf ( w_21464 , \5755_b1 );
not ( w_21464 , w_21468 );
not ( w_21465 , w_21469 );
and ( w_21468 , w_21469 , \5755_b0 );
or ( \8563_b1 , \5986_b1 , \5768_b1 );
not ( \5768_b1 , w_21470 );
and ( \8563_b0 , \5986_b0 , w_21471 );
and ( w_21470 , w_21471 , \5768_b0 );
or ( \8564_b1 , \5998_b1 , \5766_b1 );
not ( \5766_b1 , w_21472 );
and ( \8564_b0 , \5998_b0 , w_21473 );
and ( w_21472 , w_21473 , \5766_b0 );
or ( \8565_b1 , \8563_b1 , w_21475 );
not ( w_21475 , w_21476 );
and ( \8565_b0 , \8563_b0 , w_21477 );
and ( w_21476 ,  , w_21477 );
buf ( w_21475 , \8564_b1 );
not ( w_21475 , w_21478 );
not (  , w_21479 );
and ( w_21478 , w_21479 , \8564_b0 );
or ( \8566_b1 , \8565_b1 , w_21480 );
xor ( \8566_b0 , \8565_b0 , w_21482 );
not ( w_21482 , w_21483 );
and ( w_21483 , w_21480 , w_21481 );
buf ( w_21480 , \5775_b1 );
not ( w_21480 , w_21484 );
not ( w_21481 , w_21485 );
and ( w_21484 , w_21485 , \5775_b0 );
or ( \8567_b1 , \8562_b1 , \8566_b1 );
xor ( \8567_b0 , \8562_b0 , w_21486 );
not ( w_21486 , w_21487 );
and ( w_21487 , \8566_b1 , \8566_b0 );
or ( \8568_b1 , \6006_b1 , \5790_b1 );
not ( \5790_b1 , w_21488 );
and ( \8568_b0 , \6006_b0 , w_21489 );
and ( w_21488 , w_21489 , \5790_b0 );
or ( \8569_b1 , \6018_b1 , \5788_b1 );
not ( \5788_b1 , w_21490 );
and ( \8569_b0 , \6018_b0 , w_21491 );
and ( w_21490 , w_21491 , \5788_b0 );
or ( \8570_b1 , \8568_b1 , w_21493 );
not ( w_21493 , w_21494 );
and ( \8570_b0 , \8568_b0 , w_21495 );
and ( w_21494 ,  , w_21495 );
buf ( w_21493 , \8569_b1 );
not ( w_21493 , w_21496 );
not (  , w_21497 );
and ( w_21496 , w_21497 , \8569_b0 );
or ( \8571_b1 , \8570_b1 , w_21498 );
xor ( \8571_b0 , \8570_b0 , w_21500 );
not ( w_21500 , w_21501 );
and ( w_21501 , w_21498 , w_21499 );
buf ( w_21498 , \5797_b1 );
not ( w_21498 , w_21502 );
not ( w_21499 , w_21503 );
and ( w_21502 , w_21503 , \5797_b0 );
or ( \8572_b1 , \8567_b1 , \8571_b1 );
xor ( \8572_b0 , \8567_b0 , w_21504 );
not ( w_21504 , w_21505 );
and ( w_21505 , \8571_b1 , \8571_b0 );
or ( \8573_b1 , \8558_b1 , w_21506 );
xor ( \8573_b0 , \8558_b0 , w_21508 );
not ( w_21508 , w_21509 );
and ( w_21509 , w_21506 , w_21507 );
buf ( w_21506 , \8572_b1 );
not ( w_21506 , w_21510 );
not ( w_21507 , w_21511 );
and ( w_21510 , w_21511 , \8572_b0 );
or ( \8574_b1 , \8474_b1 , \8478_b1 );
not ( \8478_b1 , w_21512 );
and ( \8574_b0 , \8474_b0 , w_21513 );
and ( w_21512 , w_21513 , \8478_b0 );
or ( \8575_b1 , \8478_b1 , \8483_b1 );
not ( \8483_b1 , w_21514 );
and ( \8575_b0 , \8478_b0 , w_21515 );
and ( w_21514 , w_21515 , \8483_b0 );
or ( \8576_b1 , \8474_b1 , \8483_b1 );
not ( \8483_b1 , w_21516 );
and ( \8576_b0 , \8474_b0 , w_21517 );
and ( w_21516 , w_21517 , \8483_b0 );
or ( \8578_b1 , \8459_b1 , \8463_b1 );
not ( \8463_b1 , w_21518 );
and ( \8578_b0 , \8459_b0 , w_21519 );
and ( w_21518 , w_21519 , \8463_b0 );
or ( \8579_b1 , \8463_b1 , \8468_b1 );
not ( \8468_b1 , w_21520 );
and ( \8579_b0 , \8463_b0 , w_21521 );
and ( w_21520 , w_21521 , \8468_b0 );
or ( \8580_b1 , \8459_b1 , \8468_b1 );
not ( \8468_b1 , w_21522 );
and ( \8580_b0 , \8459_b0 , w_21523 );
and ( w_21522 , w_21523 , \8468_b0 );
or ( \8582_b1 , \8577_b1 , \8581_b1 );
xor ( \8582_b0 , \8577_b0 , w_21524 );
not ( w_21524 , w_21525 );
and ( w_21525 , \8581_b1 , \8581_b0 );
or ( \8583_b1 , \8450_b1 , \8454_b1 );
not ( \8454_b1 , w_21526 );
and ( \8583_b0 , \8450_b0 , w_21527 );
and ( w_21526 , w_21527 , \8454_b0 );
or ( \8584_b1 , \8582_b1 , \8583_b1 );
xor ( \8584_b0 , \8582_b0 , w_21528 );
not ( w_21528 , w_21529 );
and ( w_21529 , \8583_b1 , \8583_b0 );
or ( \8585_b1 , \8573_b1 , \8584_b1 );
xor ( \8585_b0 , \8573_b0 , w_21530 );
not ( w_21530 , w_21531 );
and ( w_21531 , \8584_b1 , \8584_b0 );
or ( \8586_b1 , \8434_b1 , \8438_b1 );
not ( \8438_b1 , w_21532 );
and ( \8586_b0 , \8434_b0 , w_21533 );
and ( w_21532 , w_21533 , \8438_b0 );
or ( \8587_b1 , \8438_b1 , \8443_b1 );
not ( \8443_b1 , w_21534 );
and ( \8587_b0 , \8438_b0 , w_21535 );
and ( w_21534 , w_21535 , \8443_b0 );
or ( \8588_b1 , \8434_b1 , \8443_b1 );
not ( \8443_b1 , w_21536 );
and ( \8588_b0 , \8434_b0 , w_21537 );
and ( w_21536 , w_21537 , \8443_b0 );
or ( \8590_b1 , \8422_b1 , \8426_b1 );
not ( \8426_b1 , w_21538 );
and ( \8590_b0 , \8422_b0 , w_21539 );
and ( w_21538 , w_21539 , \8426_b0 );
or ( \8591_b1 , \8426_b1 , \8431_b1 );
not ( \8431_b1 , w_21540 );
and ( \8591_b0 , \8426_b0 , w_21541 );
and ( w_21540 , w_21541 , \8431_b0 );
or ( \8592_b1 , \8422_b1 , \8431_b1 );
not ( \8431_b1 , w_21542 );
and ( \8592_b0 , \8422_b0 , w_21543 );
and ( w_21542 , w_21543 , \8431_b0 );
or ( \8594_b1 , \8589_b1 , \8593_b1 );
xor ( \8594_b0 , \8589_b0 , w_21544 );
not ( w_21544 , w_21545 );
and ( w_21545 , \8593_b1 , \8593_b0 );
or ( \8595_b1 , \8408_b1 , \8412_b1 );
not ( \8412_b1 , w_21546 );
and ( \8595_b0 , \8408_b0 , w_21547 );
and ( w_21546 , w_21547 , \8412_b0 );
or ( \8596_b1 , \8412_b1 , \8417_b1 );
not ( \8417_b1 , w_21548 );
and ( \8596_b0 , \8412_b0 , w_21549 );
and ( w_21548 , w_21549 , \8417_b0 );
or ( \8597_b1 , \8408_b1 , \8417_b1 );
not ( \8417_b1 , w_21550 );
and ( \8597_b0 , \8408_b0 , w_21551 );
and ( w_21550 , w_21551 , \8417_b0 );
or ( \8599_b1 , \8594_b1 , \8598_b1 );
xor ( \8599_b0 , \8594_b0 , w_21552 );
not ( w_21552 , w_21553 );
and ( w_21553 , \8598_b1 , \8598_b0 );
or ( \8600_b1 , \8585_b1 , \8599_b1 );
xor ( \8600_b0 , \8585_b0 , w_21554 );
not ( w_21554 , w_21555 );
and ( w_21555 , \8599_b1 , \8599_b0 );
or ( \8601_b1 , \8418_b1 , \8432_b1 );
not ( \8432_b1 , w_21556 );
and ( \8601_b0 , \8418_b0 , w_21557 );
and ( w_21556 , w_21557 , \8432_b0 );
or ( \8602_b1 , \8432_b1 , \8444_b1 );
not ( \8444_b1 , w_21558 );
and ( \8602_b0 , \8432_b0 , w_21559 );
and ( w_21558 , w_21559 , \8444_b0 );
or ( \8603_b1 , \8418_b1 , \8444_b1 );
not ( \8444_b1 , w_21560 );
and ( \8603_b0 , \8418_b0 , w_21561 );
and ( w_21560 , w_21561 , \8444_b0 );
or ( \8605_b1 , \5737_b1 , \7026_b1 );
not ( \7026_b1 , w_21562 );
and ( \8605_b0 , \5737_b0 , w_21563 );
and ( w_21562 , w_21563 , \7026_b0 );
buf ( \8606_b1 , \8605_b1 );
not ( \8606_b1 , w_21564 );
not ( \8606_b0 , w_21565 );
and ( w_21564 , w_21565 , \8605_b0 );
or ( \8607_b1 , \8606_b1 , w_21566 );
xor ( \8607_b0 , \8606_b0 , w_21568 );
not ( w_21568 , w_21569 );
and ( w_21569 , w_21566 , w_21567 );
buf ( w_21566 , \7032_b1 );
not ( w_21566 , w_21570 );
not ( w_21567 , w_21571 );
and ( w_21570 , w_21571 , \7032_b0 );
or ( \8608_b1 , \5859_b1 , \8607_b1 );
xor ( \8608_b0 , \5859_b0 , w_21572 );
not ( w_21572 , w_21573 );
and ( w_21573 , \8607_b1 , \8607_b0 );
or ( \8609_b1 , \5758_b1 , \7043_b1 );
not ( \7043_b1 , w_21574 );
and ( \8609_b0 , \5758_b0 , w_21575 );
and ( w_21574 , w_21575 , \7043_b0 );
or ( \8610_b1 , \5770_b1 , \7041_b1 );
not ( \7041_b1 , w_21576 );
and ( \8610_b0 , \5770_b0 , w_21577 );
and ( w_21576 , w_21577 , \7041_b0 );
or ( \8611_b1 , \8609_b1 , w_21579 );
not ( w_21579 , w_21580 );
and ( \8611_b0 , \8609_b0 , w_21581 );
and ( w_21580 ,  , w_21581 );
buf ( w_21579 , \8610_b1 );
not ( w_21579 , w_21582 );
not (  , w_21583 );
and ( w_21582 , w_21583 , \8610_b0 );
or ( \8612_b1 , \8611_b1 , w_21584 );
xor ( \8612_b0 , \8611_b0 , w_21586 );
not ( w_21586 , w_21587 );
and ( w_21587 , w_21584 , w_21585 );
buf ( w_21584 , \7049_b1 );
not ( w_21584 , w_21588 );
not ( w_21585 , w_21589 );
and ( w_21588 , w_21589 , \7049_b0 );
or ( \8613_b1 , \8608_b1 , \8612_b1 );
xor ( \8613_b0 , \8608_b0 , w_21590 );
not ( w_21590 , w_21591 );
and ( w_21591 , \8612_b1 , \8612_b0 );
or ( \8614_b1 , \8604_b1 , \8613_b1 );
xor ( \8614_b0 , \8604_b0 , w_21592 );
not ( w_21592 , w_21593 );
and ( w_21593 , \8613_b1 , \8613_b0 );
or ( \8615_b1 , \5906_b1 , \7175_b1 );
not ( \7175_b1 , w_21594 );
and ( \8615_b0 , \5906_b0 , w_21595 );
and ( w_21594 , w_21595 , \7175_b0 );
or ( \8616_b1 , \5918_b1 , \7173_b1 );
not ( \7173_b1 , w_21596 );
and ( \8616_b0 , \5918_b0 , w_21597 );
and ( w_21596 , w_21597 , \7173_b0 );
or ( \8617_b1 , \8615_b1 , w_21599 );
not ( w_21599 , w_21600 );
and ( \8617_b0 , \8615_b0 , w_21601 );
and ( w_21600 ,  , w_21601 );
buf ( w_21599 , \8616_b1 );
not ( w_21599 , w_21602 );
not (  , w_21603 );
and ( w_21602 , w_21603 , \8616_b0 );
or ( \8618_b1 , \8617_b1 , w_21604 );
xor ( \8618_b0 , \8617_b0 , w_21606 );
not ( w_21606 , w_21607 );
and ( w_21607 , w_21604 , w_21605 );
buf ( w_21604 , \7181_b1 );
not ( w_21604 , w_21608 );
not ( w_21605 , w_21609 );
and ( w_21608 , w_21609 , \7181_b0 );
or ( \8619_b1 , \5925_b1 , \7192_b1 );
not ( \7192_b1 , w_21610 );
and ( \8619_b0 , \5925_b0 , w_21611 );
and ( w_21610 , w_21611 , \7192_b0 );
or ( \8620_b1 , \5937_b1 , \7190_b1 );
not ( \7190_b1 , w_21612 );
and ( \8620_b0 , \5937_b0 , w_21613 );
and ( w_21612 , w_21613 , \7190_b0 );
or ( \8621_b1 , \8619_b1 , w_21615 );
not ( w_21615 , w_21616 );
and ( \8621_b0 , \8619_b0 , w_21617 );
and ( w_21616 ,  , w_21617 );
buf ( w_21615 , \8620_b1 );
not ( w_21615 , w_21618 );
not (  , w_21619 );
and ( w_21618 , w_21619 , \8620_b0 );
or ( \8622_b1 , \8621_b1 , w_21620 );
xor ( \8622_b0 , \8621_b0 , w_21622 );
not ( w_21622 , w_21623 );
and ( w_21623 , w_21620 , w_21621 );
buf ( w_21620 , \7198_b1 );
not ( w_21620 , w_21624 );
not ( w_21621 , w_21625 );
and ( w_21624 , w_21625 , \7198_b0 );
or ( \8623_b1 , \8618_b1 , \8622_b1 );
xor ( \8623_b0 , \8618_b0 , w_21626 );
not ( w_21626 , w_21627 );
and ( w_21627 , \8622_b1 , \8622_b0 );
or ( \8624_b1 , \5945_b1 , \7203_b1 );
not ( \7203_b1 , w_21628 );
and ( \8624_b0 , \5945_b0 , w_21629 );
and ( w_21628 , w_21629 , \7203_b0 );
or ( \8625_b1 , \5957_b1 , \7201_b1 );
not ( \7201_b1 , w_21630 );
and ( \8625_b0 , \5957_b0 , w_21631 );
and ( w_21630 , w_21631 , \7201_b0 );
or ( \8626_b1 , \8624_b1 , w_21633 );
not ( w_21633 , w_21634 );
and ( \8626_b0 , \8624_b0 , w_21635 );
and ( w_21634 ,  , w_21635 );
buf ( w_21633 , \8625_b1 );
not ( w_21633 , w_21636 );
not (  , w_21637 );
and ( w_21636 , w_21637 , \8625_b0 );
or ( \8627_b1 , \8626_b1 , w_21638 );
xor ( \8627_b0 , \8626_b0 , w_21640 );
not ( w_21640 , w_21641 );
and ( w_21641 , w_21638 , w_21639 );
buf ( w_21638 , \6824_b1 );
not ( w_21638 , w_21642 );
not ( w_21639 , w_21643 );
and ( w_21642 , w_21643 , \6824_b0 );
or ( \8628_b1 , \8623_b1 , \8627_b1 );
xor ( \8628_b0 , \8623_b0 , w_21644 );
not ( w_21644 , w_21645 );
and ( w_21645 , \8627_b1 , \8627_b0 );
or ( \8629_b1 , \5842_b1 , \7117_b1 );
not ( \7117_b1 , w_21646 );
and ( \8629_b0 , \5842_b0 , w_21647 );
and ( w_21646 , w_21647 , \7117_b0 );
or ( \8630_b1 , \5854_b1 , \7115_b1 );
not ( \7115_b1 , w_21648 );
and ( \8630_b0 , \5854_b0 , w_21649 );
and ( w_21648 , w_21649 , \7115_b0 );
or ( \8631_b1 , \8629_b1 , w_21651 );
not ( w_21651 , w_21652 );
and ( \8631_b0 , \8629_b0 , w_21653 );
and ( w_21652 ,  , w_21653 );
buf ( w_21651 , \8630_b1 );
not ( w_21651 , w_21654 );
not (  , w_21655 );
and ( w_21654 , w_21655 , \8630_b0 );
or ( \8632_b1 , \8631_b1 , w_21656 );
xor ( \8632_b0 , \8631_b0 , w_21658 );
not ( w_21658 , w_21659 );
and ( w_21659 , w_21656 , w_21657 );
buf ( w_21656 , \7123_b1 );
not ( w_21656 , w_21660 );
not ( w_21657 , w_21661 );
and ( w_21660 , w_21661 , \7123_b0 );
or ( \8633_b1 , \5861_b1 , \7140_b1 );
not ( \7140_b1 , w_21662 );
and ( \8633_b0 , \5861_b0 , w_21663 );
and ( w_21662 , w_21663 , \7140_b0 );
or ( \8634_b1 , \5873_b1 , \7138_b1 );
not ( \7138_b1 , w_21664 );
and ( \8634_b0 , \5873_b0 , w_21665 );
and ( w_21664 , w_21665 , \7138_b0 );
or ( \8635_b1 , \8633_b1 , w_21667 );
not ( w_21667 , w_21668 );
and ( \8635_b0 , \8633_b0 , w_21669 );
and ( w_21668 ,  , w_21669 );
buf ( w_21667 , \8634_b1 );
not ( w_21667 , w_21670 );
not (  , w_21671 );
and ( w_21670 , w_21671 , \8634_b0 );
or ( \8636_b1 , \8635_b1 , w_21672 );
xor ( \8636_b0 , \8635_b0 , w_21674 );
not ( w_21674 , w_21675 );
and ( w_21675 , w_21672 , w_21673 );
buf ( w_21672 , \7146_b1 );
not ( w_21672 , w_21676 );
not ( w_21673 , w_21677 );
and ( w_21676 , w_21677 , \7146_b0 );
or ( \8637_b1 , \8632_b1 , \8636_b1 );
xor ( \8637_b0 , \8632_b0 , w_21678 );
not ( w_21678 , w_21679 );
and ( w_21679 , \8636_b1 , \8636_b0 );
or ( \8638_b1 , \5881_b1 , \7157_b1 );
not ( \7157_b1 , w_21680 );
and ( \8638_b0 , \5881_b0 , w_21681 );
and ( w_21680 , w_21681 , \7157_b0 );
or ( \8639_b1 , \5893_b1 , \7155_b1 );
not ( \7155_b1 , w_21682 );
and ( \8639_b0 , \5893_b0 , w_21683 );
and ( w_21682 , w_21683 , \7155_b0 );
or ( \8640_b1 , \8638_b1 , w_21685 );
not ( w_21685 , w_21686 );
and ( \8640_b0 , \8638_b0 , w_21687 );
and ( w_21686 ,  , w_21687 );
buf ( w_21685 , \8639_b1 );
not ( w_21685 , w_21688 );
not (  , w_21689 );
and ( w_21688 , w_21689 , \8639_b0 );
or ( \8641_b1 , \8640_b1 , w_21690 );
xor ( \8641_b0 , \8640_b0 , w_21692 );
not ( w_21692 , w_21693 );
and ( w_21693 , w_21690 , w_21691 );
buf ( w_21690 , \7163_b1 );
not ( w_21690 , w_21694 );
not ( w_21691 , w_21695 );
and ( w_21694 , w_21695 , \7163_b0 );
or ( \8642_b1 , \8637_b1 , \8641_b1 );
xor ( \8642_b0 , \8637_b0 , w_21696 );
not ( w_21696 , w_21697 );
and ( w_21697 , \8641_b1 , \8641_b0 );
or ( \8643_b1 , \8628_b1 , \8642_b1 );
xor ( \8643_b0 , \8628_b0 , w_21698 );
not ( w_21698 , w_21699 );
and ( w_21699 , \8642_b1 , \8642_b0 );
or ( \8644_b1 , \5780_b1 , \7061_b1 );
not ( \7061_b1 , w_21700 );
and ( \8644_b0 , \5780_b0 , w_21701 );
and ( w_21700 , w_21701 , \7061_b0 );
or ( \8645_b1 , \5792_b1 , \7059_b1 );
not ( \7059_b1 , w_21702 );
and ( \8645_b0 , \5792_b0 , w_21703 );
and ( w_21702 , w_21703 , \7059_b0 );
or ( \8646_b1 , \8644_b1 , w_21705 );
not ( w_21705 , w_21706 );
and ( \8646_b0 , \8644_b0 , w_21707 );
and ( w_21706 ,  , w_21707 );
buf ( w_21705 , \8645_b1 );
not ( w_21705 , w_21708 );
not (  , w_21709 );
and ( w_21708 , w_21709 , \8645_b0 );
or ( \8647_b1 , \8646_b1 , w_21710 );
xor ( \8647_b0 , \8646_b0 , w_21712 );
not ( w_21712 , w_21713 );
and ( w_21713 , w_21710 , w_21711 );
buf ( w_21710 , \7067_b1 );
not ( w_21710 , w_21714 );
not ( w_21711 , w_21715 );
and ( w_21714 , w_21715 , \7067_b0 );
or ( \8648_b1 , \5799_b1 , \7082_b1 );
not ( \7082_b1 , w_21716 );
and ( \8648_b0 , \5799_b0 , w_21717 );
and ( w_21716 , w_21717 , \7082_b0 );
or ( \8649_b1 , \5811_b1 , \7080_b1 );
not ( \7080_b1 , w_21718 );
and ( \8649_b0 , \5811_b0 , w_21719 );
and ( w_21718 , w_21719 , \7080_b0 );
or ( \8650_b1 , \8648_b1 , w_21721 );
not ( w_21721 , w_21722 );
and ( \8650_b0 , \8648_b0 , w_21723 );
and ( w_21722 ,  , w_21723 );
buf ( w_21721 , \8649_b1 );
not ( w_21721 , w_21724 );
not (  , w_21725 );
and ( w_21724 , w_21725 , \8649_b0 );
or ( \8651_b1 , \8650_b1 , w_21726 );
xor ( \8651_b0 , \8650_b0 , w_21728 );
not ( w_21728 , w_21729 );
and ( w_21729 , w_21726 , w_21727 );
buf ( w_21726 , \7088_b1 );
not ( w_21726 , w_21730 );
not ( w_21727 , w_21731 );
and ( w_21730 , w_21731 , \7088_b0 );
or ( \8652_b1 , \8647_b1 , \8651_b1 );
xor ( \8652_b0 , \8647_b0 , w_21732 );
not ( w_21732 , w_21733 );
and ( w_21733 , \8651_b1 , \8651_b0 );
or ( \8653_b1 , \5819_b1 , \7099_b1 );
not ( \7099_b1 , w_21734 );
and ( \8653_b0 , \5819_b0 , w_21735 );
and ( w_21734 , w_21735 , \7099_b0 );
or ( \8654_b1 , \5831_b1 , \7097_b1 );
not ( \7097_b1 , w_21736 );
and ( \8654_b0 , \5831_b0 , w_21737 );
and ( w_21736 , w_21737 , \7097_b0 );
or ( \8655_b1 , \8653_b1 , w_21739 );
not ( w_21739 , w_21740 );
and ( \8655_b0 , \8653_b0 , w_21741 );
and ( w_21740 ,  , w_21741 );
buf ( w_21739 , \8654_b1 );
not ( w_21739 , w_21742 );
not (  , w_21743 );
and ( w_21742 , w_21743 , \8654_b0 );
or ( \8656_b1 , \8655_b1 , w_21744 );
xor ( \8656_b0 , \8655_b0 , w_21746 );
not ( w_21746 , w_21747 );
and ( w_21747 , w_21744 , w_21745 );
buf ( w_21744 , \7105_b1 );
not ( w_21744 , w_21748 );
not ( w_21745 , w_21749 );
and ( w_21748 , w_21749 , \7105_b0 );
or ( \8657_b1 , \8652_b1 , \8656_b1 );
xor ( \8657_b0 , \8652_b0 , w_21750 );
not ( w_21750 , w_21751 );
and ( w_21751 , \8656_b1 , \8656_b0 );
or ( \8658_b1 , \8643_b1 , \8657_b1 );
xor ( \8658_b0 , \8643_b0 , w_21752 );
not ( w_21752 , w_21753 );
and ( w_21753 , \8657_b1 , \8657_b0 );
or ( \8659_b1 , \8614_b1 , \8658_b1 );
xor ( \8659_b0 , \8614_b0 , w_21754 );
not ( w_21754 , w_21755 );
and ( w_21755 , \8658_b1 , \8658_b0 );
or ( \8660_b1 , \8600_b1 , \8659_b1 );
xor ( \8660_b0 , \8600_b0 , w_21756 );
not ( w_21756 , w_21757 );
and ( w_21757 , \8659_b1 , \8659_b0 );
or ( \8661_b1 , \8389_b1 , \8393_b1 );
not ( \8393_b1 , w_21758 );
and ( \8661_b0 , \8389_b0 , w_21759 );
and ( w_21758 , w_21759 , \8393_b0 );
or ( \8662_b1 , \8393_b1 , \8398_b1 );
not ( \8398_b1 , w_21760 );
and ( \8662_b0 , \8393_b0 , w_21761 );
and ( w_21760 , w_21761 , \8398_b0 );
or ( \8663_b1 , \8389_b1 , \8398_b1 );
not ( \8398_b1 , w_21762 );
and ( \8663_b0 , \8389_b0 , w_21763 );
and ( w_21762 , w_21763 , \8398_b0 );
or ( \8665_b1 , \8375_b1 , \8379_b1 );
not ( \8379_b1 , w_21764 );
and ( \8665_b0 , \8375_b0 , w_21765 );
and ( w_21764 , w_21765 , \8379_b0 );
or ( \8666_b1 , \8379_b1 , \8384_b1 );
not ( \8384_b1 , w_21766 );
and ( \8666_b0 , \8379_b0 , w_21767 );
and ( w_21766 , w_21767 , \8384_b0 );
or ( \8667_b1 , \8375_b1 , \8384_b1 );
not ( \8384_b1 , w_21768 );
and ( \8667_b0 , \8375_b0 , w_21769 );
and ( w_21768 , w_21769 , \8384_b0 );
or ( \8669_b1 , \8664_b1 , \8668_b1 );
xor ( \8669_b0 , \8664_b0 , w_21770 );
not ( w_21770 , w_21771 );
and ( w_21771 , \8668_b1 , \8668_b0 );
or ( \8670_b1 , \8455_b1 , \8469_b1 );
not ( \8469_b1 , w_21772 );
and ( \8670_b0 , \8455_b0 , w_21773 );
and ( w_21772 , w_21773 , \8469_b0 );
or ( \8671_b1 , \8469_b1 , \8484_b1 );
not ( \8484_b1 , w_21774 );
and ( \8671_b0 , \8469_b0 , w_21775 );
and ( w_21774 , w_21775 , \8484_b0 );
or ( \8672_b1 , \8455_b1 , \8484_b1 );
not ( \8484_b1 , w_21776 );
and ( \8672_b0 , \8455_b0 , w_21777 );
and ( w_21776 , w_21777 , \8484_b0 );
or ( \8674_b1 , \8669_b1 , \8673_b1 );
xor ( \8674_b0 , \8669_b0 , w_21778 );
not ( w_21778 , w_21779 );
and ( w_21779 , \8673_b1 , \8673_b0 );
or ( \8675_b1 , \8660_b1 , \8674_b1 );
xor ( \8675_b0 , \8660_b0 , w_21780 );
not ( w_21780 , w_21781 );
and ( w_21781 , \8674_b1 , \8674_b0 );
or ( \8676_b1 , \8546_b1 , \8675_b1 );
xor ( \8676_b0 , \8546_b0 , w_21782 );
not ( w_21782 , w_21783 );
and ( w_21783 , \8675_b1 , \8675_b0 );
or ( \8677_b1 , \8537_b1 , \8676_b1 );
xor ( \8677_b0 , \8537_b0 , w_21784 );
not ( w_21784 , w_21785 );
and ( w_21785 , \8676_b1 , \8676_b0 );
or ( \8678_b1 , \8365_b1 , \8366_b1 );
not ( \8366_b1 , w_21786 );
and ( \8678_b0 , \8365_b0 , w_21787 );
and ( w_21786 , w_21787 , \8366_b0 );
or ( \8679_b1 , \8366_b1 , \8515_b1 );
not ( \8515_b1 , w_21788 );
and ( \8679_b0 , \8366_b0 , w_21789 );
and ( w_21788 , w_21789 , \8515_b0 );
or ( \8680_b1 , \8365_b1 , \8515_b1 );
not ( \8515_b1 , w_21790 );
and ( \8680_b0 , \8365_b0 , w_21791 );
and ( w_21790 , w_21791 , \8515_b0 );
or ( \8682_b1 , \8677_b1 , w_21793 );
not ( w_21793 , w_21794 );
and ( \8682_b0 , \8677_b0 , w_21795 );
and ( w_21794 ,  , w_21795 );
buf ( w_21793 , \8681_b1 );
not ( w_21793 , w_21796 );
not (  , w_21797 );
and ( w_21796 , w_21797 , \8681_b0 );
or ( \8683_b1 , \8521_b1 , w_21799 );
not ( w_21799 , w_21800 );
and ( \8683_b0 , \8521_b0 , w_21801 );
and ( w_21800 ,  , w_21801 );
buf ( w_21799 , \8682_b1 );
not ( w_21799 , w_21802 );
not (  , w_21803 );
and ( w_21802 , w_21803 , \8682_b0 );
or ( \8684_b1 , \8541_b1 , \8545_b1 );
not ( \8545_b1 , w_21804 );
and ( \8684_b0 , \8541_b0 , w_21805 );
and ( w_21804 , w_21805 , \8545_b0 );
or ( \8685_b1 , \8545_b1 , \8675_b1 );
not ( \8675_b1 , w_21806 );
and ( \8685_b0 , \8545_b0 , w_21807 );
and ( w_21806 , w_21807 , \8675_b0 );
or ( \8686_b1 , \8541_b1 , \8675_b1 );
not ( \8675_b1 , w_21808 );
and ( \8686_b0 , \8541_b0 , w_21809 );
and ( w_21808 , w_21809 , \8675_b0 );
or ( \8688_b1 , \8664_b1 , \8668_b1 );
not ( \8668_b1 , w_21810 );
and ( \8688_b0 , \8664_b0 , w_21811 );
and ( w_21810 , w_21811 , \8668_b0 );
or ( \8689_b1 , \8668_b1 , \8673_b1 );
not ( \8673_b1 , w_21812 );
and ( \8689_b0 , \8668_b0 , w_21813 );
and ( w_21812 , w_21813 , \8673_b0 );
or ( \8690_b1 , \8664_b1 , \8673_b1 );
not ( \8673_b1 , w_21814 );
and ( \8690_b0 , \8664_b0 , w_21815 );
and ( w_21814 , w_21815 , \8673_b0 );
or ( \8692_b1 , \8604_b1 , \8613_b1 );
not ( \8613_b1 , w_21816 );
and ( \8692_b0 , \8604_b0 , w_21817 );
and ( w_21816 , w_21817 , \8613_b0 );
or ( \8693_b1 , \8613_b1 , \8658_b1 );
not ( \8658_b1 , w_21818 );
and ( \8693_b0 , \8613_b0 , w_21819 );
and ( w_21818 , w_21819 , \8658_b0 );
or ( \8694_b1 , \8604_b1 , \8658_b1 );
not ( \8658_b1 , w_21820 );
and ( \8694_b0 , \8604_b0 , w_21821 );
and ( w_21820 , w_21821 , \8658_b0 );
or ( \8696_b1 , \8691_b1 , \8695_b1 );
xor ( \8696_b0 , \8691_b0 , w_21822 );
not ( w_21822 , w_21823 );
and ( w_21823 , \8695_b1 , \8695_b0 );
or ( \8697_b1 , \8573_b1 , \8584_b1 );
not ( \8584_b1 , w_21824 );
and ( \8697_b0 , \8573_b0 , w_21825 );
and ( w_21824 , w_21825 , \8584_b0 );
or ( \8698_b1 , \8584_b1 , \8599_b1 );
not ( \8599_b1 , w_21826 );
and ( \8698_b0 , \8584_b0 , w_21827 );
and ( w_21826 , w_21827 , \8599_b0 );
or ( \8699_b1 , \8573_b1 , \8599_b1 );
not ( \8599_b1 , w_21828 );
and ( \8699_b0 , \8573_b0 , w_21829 );
and ( w_21828 , w_21829 , \8599_b0 );
or ( \8701_b1 , \8696_b1 , \8700_b1 );
xor ( \8701_b0 , \8696_b0 , w_21830 );
not ( w_21830 , w_21831 );
and ( w_21831 , \8700_b1 , \8700_b0 );
or ( \8702_b1 , \8687_b1 , \8701_b1 );
xor ( \8702_b0 , \8687_b0 , w_21832 );
not ( w_21832 , w_21833 );
and ( w_21833 , \8701_b1 , \8701_b0 );
or ( \8703_b1 , \8529_b1 , \8533_b1 );
not ( \8533_b1 , w_21834 );
and ( \8703_b0 , \8529_b0 , w_21835 );
and ( w_21834 , w_21835 , \8533_b0 );
or ( \8704_b1 , \8533_b1 , \8535_b1 );
not ( \8535_b1 , w_21836 );
and ( \8704_b0 , \8533_b0 , w_21837 );
and ( w_21836 , w_21837 , \8535_b0 );
or ( \8705_b1 , \8529_b1 , \8535_b1 );
not ( \8535_b1 , w_21838 );
and ( \8705_b0 , \8529_b0 , w_21839 );
and ( w_21838 , w_21839 , \8535_b0 );
or ( \8707_b1 , \8600_b1 , \8659_b1 );
not ( \8659_b1 , w_21840 );
and ( \8707_b0 , \8600_b0 , w_21841 );
and ( w_21840 , w_21841 , \8659_b0 );
or ( \8708_b1 , \8659_b1 , \8674_b1 );
not ( \8674_b1 , w_21842 );
and ( \8708_b0 , \8659_b0 , w_21843 );
and ( w_21842 , w_21843 , \8674_b0 );
or ( \8709_b1 , \8600_b1 , \8674_b1 );
not ( \8674_b1 , w_21844 );
and ( \8709_b0 , \8600_b0 , w_21845 );
and ( w_21844 , w_21845 , \8674_b0 );
or ( \8711_b1 , \8706_b1 , \8710_b1 );
xor ( \8711_b0 , \8706_b0 , w_21846 );
not ( w_21846 , w_21847 );
and ( w_21847 , \8710_b1 , \8710_b0 );
or ( \8712_b1 , \8618_b1 , \8622_b1 );
not ( \8622_b1 , w_21848 );
and ( \8712_b0 , \8618_b0 , w_21849 );
and ( w_21848 , w_21849 , \8622_b0 );
or ( \8713_b1 , \8622_b1 , \8627_b1 );
not ( \8627_b1 , w_21850 );
and ( \8713_b0 , \8622_b0 , w_21851 );
and ( w_21850 , w_21851 , \8627_b0 );
or ( \8714_b1 , \8618_b1 , \8627_b1 );
not ( \8627_b1 , w_21852 );
and ( \8714_b0 , \8618_b0 , w_21853 );
and ( w_21852 , w_21853 , \8627_b0 );
or ( \8716_b1 , \8562_b1 , \8566_b1 );
not ( \8566_b1 , w_21854 );
and ( \8716_b0 , \8562_b0 , w_21855 );
and ( w_21854 , w_21855 , \8566_b0 );
or ( \8717_b1 , \8566_b1 , \8571_b1 );
not ( \8571_b1 , w_21856 );
and ( \8717_b0 , \8566_b0 , w_21857 );
and ( w_21856 , w_21857 , \8571_b0 );
or ( \8718_b1 , \8562_b1 , \8571_b1 );
not ( \8571_b1 , w_21858 );
and ( \8718_b0 , \8562_b0 , w_21859 );
and ( w_21858 , w_21859 , \8571_b0 );
or ( \8720_b1 , \8715_b1 , \8719_b1 );
xor ( \8720_b0 , \8715_b0 , w_21860 );
not ( w_21860 , w_21861 );
and ( w_21861 , \8719_b1 , \8719_b0 );
or ( \8721_b1 , \8550_b1 , \8554_b1 );
not ( \8554_b1 , w_21862 );
and ( \8721_b0 , \8550_b0 , w_21863 );
and ( w_21862 , w_21863 , \8554_b0 );
or ( \8722_b1 , \8554_b1 , \8557_b1 );
not ( \8557_b1 , w_21864 );
and ( \8722_b0 , \8554_b0 , w_21865 );
and ( w_21864 , w_21865 , \8557_b0 );
or ( \8723_b1 , \8550_b1 , \8557_b1 );
not ( \8557_b1 , w_21866 );
and ( \8723_b0 , \8550_b0 , w_21867 );
and ( w_21866 , w_21867 , \8557_b0 );
or ( \8725_b1 , \8720_b1 , \8724_b1 );
xor ( \8725_b0 , \8720_b0 , w_21868 );
not ( w_21868 , w_21869 );
and ( w_21869 , \8724_b1 , \8724_b0 );
or ( \8726_b1 , \5859_b1 , \8607_b1 );
not ( \8607_b1 , w_21870 );
and ( \8726_b0 , \5859_b0 , w_21871 );
and ( w_21870 , w_21871 , \8607_b0 );
or ( \8727_b1 , \8607_b1 , \8612_b1 );
not ( \8612_b1 , w_21872 );
and ( \8727_b0 , \8607_b0 , w_21873 );
and ( w_21872 , w_21873 , \8612_b0 );
or ( \8728_b1 , \5859_b1 , \8612_b1 );
not ( \8612_b1 , w_21874 );
and ( \8728_b0 , \5859_b0 , w_21875 );
and ( w_21874 , w_21875 , \8612_b0 );
or ( \8730_b1 , \8647_b1 , \8651_b1 );
not ( \8651_b1 , w_21876 );
and ( \8730_b0 , \8647_b0 , w_21877 );
and ( w_21876 , w_21877 , \8651_b0 );
or ( \8731_b1 , \8651_b1 , \8656_b1 );
not ( \8656_b1 , w_21878 );
and ( \8731_b0 , \8651_b0 , w_21879 );
and ( w_21878 , w_21879 , \8656_b0 );
or ( \8732_b1 , \8647_b1 , \8656_b1 );
not ( \8656_b1 , w_21880 );
and ( \8732_b0 , \8647_b0 , w_21881 );
and ( w_21880 , w_21881 , \8656_b0 );
or ( \8734_b1 , \8729_b1 , \8733_b1 );
xor ( \8734_b0 , \8729_b0 , w_21882 );
not ( w_21882 , w_21883 );
and ( w_21883 , \8733_b1 , \8733_b0 );
or ( \8735_b1 , \8632_b1 , \8636_b1 );
not ( \8636_b1 , w_21884 );
and ( \8735_b0 , \8632_b0 , w_21885 );
and ( w_21884 , w_21885 , \8636_b0 );
or ( \8736_b1 , \8636_b1 , \8641_b1 );
not ( \8641_b1 , w_21886 );
and ( \8736_b0 , \8636_b0 , w_21887 );
and ( w_21886 , w_21887 , \8641_b0 );
or ( \8737_b1 , \8632_b1 , \8641_b1 );
not ( \8641_b1 , w_21888 );
and ( \8737_b0 , \8632_b0 , w_21889 );
and ( w_21888 , w_21889 , \8641_b0 );
or ( \8739_b1 , \8734_b1 , \8738_b1 );
xor ( \8739_b0 , \8734_b0 , w_21890 );
not ( w_21890 , w_21891 );
and ( w_21891 , \8738_b1 , \8738_b0 );
or ( \8740_b1 , \8725_b1 , \8739_b1 );
xor ( \8740_b0 , \8725_b0 , w_21892 );
not ( w_21892 , w_21893 );
and ( w_21893 , \8739_b1 , \8739_b0 );
or ( \8741_b1 , \8628_b1 , \8642_b1 );
not ( \8642_b1 , w_21894 );
and ( \8741_b0 , \8628_b0 , w_21895 );
and ( w_21894 , w_21895 , \8642_b0 );
or ( \8742_b1 , \8642_b1 , \8657_b1 );
not ( \8657_b1 , w_21896 );
and ( \8742_b0 , \8642_b0 , w_21897 );
and ( w_21896 , w_21897 , \8657_b0 );
or ( \8743_b1 , \8628_b1 , \8657_b1 );
not ( \8657_b1 , w_21898 );
and ( \8743_b0 , \8628_b0 , w_21899 );
and ( w_21898 , w_21899 , \8657_b0 );
or ( \8745_b1 , \5873_b1 , \7140_b1 );
not ( \7140_b1 , w_21900 );
and ( \8745_b0 , \5873_b0 , w_21901 );
and ( w_21900 , w_21901 , \7140_b0 );
or ( \8746_b1 , \5842_b1 , \7138_b1 );
not ( \7138_b1 , w_21902 );
and ( \8746_b0 , \5842_b0 , w_21903 );
and ( w_21902 , w_21903 , \7138_b0 );
or ( \8747_b1 , \8745_b1 , w_21905 );
not ( w_21905 , w_21906 );
and ( \8747_b0 , \8745_b0 , w_21907 );
and ( w_21906 ,  , w_21907 );
buf ( w_21905 , \8746_b1 );
not ( w_21905 , w_21908 );
not (  , w_21909 );
and ( w_21908 , w_21909 , \8746_b0 );
or ( \8748_b1 , \8747_b1 , w_21910 );
xor ( \8748_b0 , \8747_b0 , w_21912 );
not ( w_21912 , w_21913 );
and ( w_21913 , w_21910 , w_21911 );
buf ( w_21910 , \7146_b1 );
not ( w_21910 , w_21914 );
not ( w_21911 , w_21915 );
and ( w_21914 , w_21915 , \7146_b0 );
or ( \8749_b1 , \5893_b1 , \7157_b1 );
not ( \7157_b1 , w_21916 );
and ( \8749_b0 , \5893_b0 , w_21917 );
and ( w_21916 , w_21917 , \7157_b0 );
or ( \8750_b1 , \5861_b1 , \7155_b1 );
not ( \7155_b1 , w_21918 );
and ( \8750_b0 , \5861_b0 , w_21919 );
and ( w_21918 , w_21919 , \7155_b0 );
or ( \8751_b1 , \8749_b1 , w_21921 );
not ( w_21921 , w_21922 );
and ( \8751_b0 , \8749_b0 , w_21923 );
and ( w_21922 ,  , w_21923 );
buf ( w_21921 , \8750_b1 );
not ( w_21921 , w_21924 );
not (  , w_21925 );
and ( w_21924 , w_21925 , \8750_b0 );
or ( \8752_b1 , \8751_b1 , w_21926 );
xor ( \8752_b0 , \8751_b0 , w_21928 );
not ( w_21928 , w_21929 );
and ( w_21929 , w_21926 , w_21927 );
buf ( w_21926 , \7163_b1 );
not ( w_21926 , w_21930 );
not ( w_21927 , w_21931 );
and ( w_21930 , w_21931 , \7163_b0 );
or ( \8753_b1 , \8748_b1 , \8752_b1 );
xor ( \8753_b0 , \8748_b0 , w_21932 );
not ( w_21932 , w_21933 );
and ( w_21933 , \8752_b1 , \8752_b0 );
or ( \8754_b1 , \5918_b1 , \7175_b1 );
not ( \7175_b1 , w_21934 );
and ( \8754_b0 , \5918_b0 , w_21935 );
and ( w_21934 , w_21935 , \7175_b0 );
or ( \8755_b1 , \5881_b1 , \7173_b1 );
not ( \7173_b1 , w_21936 );
and ( \8755_b0 , \5881_b0 , w_21937 );
and ( w_21936 , w_21937 , \7173_b0 );
or ( \8756_b1 , \8754_b1 , w_21939 );
not ( w_21939 , w_21940 );
and ( \8756_b0 , \8754_b0 , w_21941 );
and ( w_21940 ,  , w_21941 );
buf ( w_21939 , \8755_b1 );
not ( w_21939 , w_21942 );
not (  , w_21943 );
and ( w_21942 , w_21943 , \8755_b0 );
or ( \8757_b1 , \8756_b1 , w_21944 );
xor ( \8757_b0 , \8756_b0 , w_21946 );
not ( w_21946 , w_21947 );
and ( w_21947 , w_21944 , w_21945 );
buf ( w_21944 , \7181_b1 );
not ( w_21944 , w_21948 );
not ( w_21945 , w_21949 );
and ( w_21948 , w_21949 , \7181_b0 );
or ( \8758_b1 , \8753_b1 , \8757_b1 );
xor ( \8758_b0 , \8753_b0 , w_21950 );
not ( w_21950 , w_21951 );
and ( w_21951 , \8757_b1 , \8757_b0 );
or ( \8759_b1 , \5811_b1 , \7082_b1 );
not ( \7082_b1 , w_21952 );
and ( \8759_b0 , \5811_b0 , w_21953 );
and ( w_21952 , w_21953 , \7082_b0 );
or ( \8760_b1 , \5780_b1 , \7080_b1 );
not ( \7080_b1 , w_21954 );
and ( \8760_b0 , \5780_b0 , w_21955 );
and ( w_21954 , w_21955 , \7080_b0 );
or ( \8761_b1 , \8759_b1 , w_21957 );
not ( w_21957 , w_21958 );
and ( \8761_b0 , \8759_b0 , w_21959 );
and ( w_21958 ,  , w_21959 );
buf ( w_21957 , \8760_b1 );
not ( w_21957 , w_21960 );
not (  , w_21961 );
and ( w_21960 , w_21961 , \8760_b0 );
or ( \8762_b1 , \8761_b1 , w_21962 );
xor ( \8762_b0 , \8761_b0 , w_21964 );
not ( w_21964 , w_21965 );
and ( w_21965 , w_21962 , w_21963 );
buf ( w_21962 , \7088_b1 );
not ( w_21962 , w_21966 );
not ( w_21963 , w_21967 );
and ( w_21966 , w_21967 , \7088_b0 );
or ( \8763_b1 , \5831_b1 , \7099_b1 );
not ( \7099_b1 , w_21968 );
and ( \8763_b0 , \5831_b0 , w_21969 );
and ( w_21968 , w_21969 , \7099_b0 );
or ( \8764_b1 , \5799_b1 , \7097_b1 );
not ( \7097_b1 , w_21970 );
and ( \8764_b0 , \5799_b0 , w_21971 );
and ( w_21970 , w_21971 , \7097_b0 );
or ( \8765_b1 , \8763_b1 , w_21973 );
not ( w_21973 , w_21974 );
and ( \8765_b0 , \8763_b0 , w_21975 );
and ( w_21974 ,  , w_21975 );
buf ( w_21973 , \8764_b1 );
not ( w_21973 , w_21976 );
not (  , w_21977 );
and ( w_21976 , w_21977 , \8764_b0 );
or ( \8766_b1 , \8765_b1 , w_21978 );
xor ( \8766_b0 , \8765_b0 , w_21980 );
not ( w_21980 , w_21981 );
and ( w_21981 , w_21978 , w_21979 );
buf ( w_21978 , \7105_b1 );
not ( w_21978 , w_21982 );
not ( w_21979 , w_21983 );
and ( w_21982 , w_21983 , \7105_b0 );
or ( \8767_b1 , \8762_b1 , \8766_b1 );
xor ( \8767_b0 , \8762_b0 , w_21984 );
not ( w_21984 , w_21985 );
and ( w_21985 , \8766_b1 , \8766_b0 );
or ( \8768_b1 , \5854_b1 , \7117_b1 );
not ( \7117_b1 , w_21986 );
and ( \8768_b0 , \5854_b0 , w_21987 );
and ( w_21986 , w_21987 , \7117_b0 );
or ( \8769_b1 , \5819_b1 , \7115_b1 );
not ( \7115_b1 , w_21988 );
and ( \8769_b0 , \5819_b0 , w_21989 );
and ( w_21988 , w_21989 , \7115_b0 );
or ( \8770_b1 , \8768_b1 , w_21991 );
not ( w_21991 , w_21992 );
and ( \8770_b0 , \8768_b0 , w_21993 );
and ( w_21992 ,  , w_21993 );
buf ( w_21991 , \8769_b1 );
not ( w_21991 , w_21994 );
not (  , w_21995 );
and ( w_21994 , w_21995 , \8769_b0 );
or ( \8771_b1 , \8770_b1 , w_21996 );
xor ( \8771_b0 , \8770_b0 , w_21998 );
not ( w_21998 , w_21999 );
and ( w_21999 , w_21996 , w_21997 );
buf ( w_21996 , \7123_b1 );
not ( w_21996 , w_22000 );
not ( w_21997 , w_22001 );
and ( w_22000 , w_22001 , \7123_b0 );
or ( \8772_b1 , \8767_b1 , \8771_b1 );
xor ( \8772_b0 , \8767_b0 , w_22002 );
not ( w_22002 , w_22003 );
and ( w_22003 , \8771_b1 , \8771_b0 );
or ( \8773_b1 , \8758_b1 , \8772_b1 );
xor ( \8773_b0 , \8758_b0 , w_22004 );
not ( w_22004 , w_22005 );
and ( w_22005 , \8772_b1 , \8772_b0 );
buf ( \8774_b1 , \7032_b1 );
not ( \8774_b1 , w_22006 );
not ( \8774_b0 , w_22007 );
and ( w_22006 , w_22007 , \7032_b0 );
or ( \8775_b1 , \5770_b1 , \7043_b1 );
not ( \7043_b1 , w_22008 );
and ( \8775_b0 , \5770_b0 , w_22009 );
and ( w_22008 , w_22009 , \7043_b0 );
or ( \8776_b1 , \5737_b1 , \7041_b1 );
not ( \7041_b1 , w_22010 );
and ( \8776_b0 , \5737_b0 , w_22011 );
and ( w_22010 , w_22011 , \7041_b0 );
or ( \8777_b1 , \8775_b1 , w_22013 );
not ( w_22013 , w_22014 );
and ( \8777_b0 , \8775_b0 , w_22015 );
and ( w_22014 ,  , w_22015 );
buf ( w_22013 , \8776_b1 );
not ( w_22013 , w_22016 );
not (  , w_22017 );
and ( w_22016 , w_22017 , \8776_b0 );
or ( \8778_b1 , \8777_b1 , w_22018 );
xor ( \8778_b0 , \8777_b0 , w_22020 );
not ( w_22020 , w_22021 );
and ( w_22021 , w_22018 , w_22019 );
buf ( w_22018 , \7049_b1 );
not ( w_22018 , w_22022 );
not ( w_22019 , w_22023 );
and ( w_22022 , w_22023 , \7049_b0 );
or ( \8779_b1 , \8774_b1 , \8778_b1 );
xor ( \8779_b0 , \8774_b0 , w_22024 );
not ( w_22024 , w_22025 );
and ( w_22025 , \8778_b1 , \8778_b0 );
or ( \8780_b1 , \5792_b1 , \7061_b1 );
not ( \7061_b1 , w_22026 );
and ( \8780_b0 , \5792_b0 , w_22027 );
and ( w_22026 , w_22027 , \7061_b0 );
or ( \8781_b1 , \5758_b1 , \7059_b1 );
not ( \7059_b1 , w_22028 );
and ( \8781_b0 , \5758_b0 , w_22029 );
and ( w_22028 , w_22029 , \7059_b0 );
or ( \8782_b1 , \8780_b1 , w_22031 );
not ( w_22031 , w_22032 );
and ( \8782_b0 , \8780_b0 , w_22033 );
and ( w_22032 ,  , w_22033 );
buf ( w_22031 , \8781_b1 );
not ( w_22031 , w_22034 );
not (  , w_22035 );
and ( w_22034 , w_22035 , \8781_b0 );
or ( \8783_b1 , \8782_b1 , w_22036 );
xor ( \8783_b0 , \8782_b0 , w_22038 );
not ( w_22038 , w_22039 );
and ( w_22039 , w_22036 , w_22037 );
buf ( w_22036 , \7067_b1 );
not ( w_22036 , w_22040 );
not ( w_22037 , w_22041 );
and ( w_22040 , w_22041 , \7067_b0 );
or ( \8784_b1 , \8779_b1 , \8783_b1 );
xor ( \8784_b0 , \8779_b0 , w_22042 );
not ( w_22042 , w_22043 );
and ( w_22043 , \8783_b1 , \8783_b0 );
or ( \8785_b1 , \8773_b1 , \8784_b1 );
xor ( \8785_b0 , \8773_b0 , w_22044 );
not ( w_22044 , w_22045 );
and ( w_22045 , \8784_b1 , \8784_b0 );
or ( \8786_b1 , \8744_b1 , \8785_b1 );
xor ( \8786_b0 , \8744_b0 , w_22046 );
not ( w_22046 , w_22047 );
and ( w_22047 , \8785_b1 , \8785_b0 );
or ( \8787_b1 , \6057_b1 , \5829_b1 );
not ( \5829_b1 , w_22048 );
and ( \8787_b0 , \6057_b0 , w_22049 );
and ( w_22048 , w_22049 , \5829_b0 );
or ( \8788_b1 , \6029_b1 , \5827_b1 );
not ( \5827_b1 , w_22050 );
and ( \8788_b0 , \6029_b0 , w_22051 );
and ( w_22050 , w_22051 , \5827_b0 );
or ( \8789_b1 , \8787_b1 , w_22053 );
not ( w_22053 , w_22054 );
and ( \8789_b0 , \8787_b0 , w_22055 );
and ( w_22054 ,  , w_22055 );
buf ( w_22053 , \8788_b1 );
not ( w_22053 , w_22056 );
not (  , w_22057 );
and ( w_22056 , w_22057 , \8788_b0 );
or ( \8790_b1 , \8789_b1 , w_22058 );
xor ( \8790_b0 , \8789_b0 , w_22060 );
not ( w_22060 , w_22061 );
and ( w_22061 , w_22058 , w_22059 );
buf ( w_22058 , \5836_b1 );
not ( w_22058 , w_22062 );
not ( w_22059 , w_22063 );
and ( w_22062 , w_22063 , \5836_b0 );
or ( \8791_b1 , \6065_b1 , \5852_b1 );
not ( \5852_b1 , w_22064 );
and ( \8791_b0 , \6065_b0 , w_22065 );
and ( w_22064 , w_22065 , \5852_b0 );
or ( \8792_b1 , \6048_b1 , \5850_b1 );
not ( \5850_b1 , w_22066 );
and ( \8792_b0 , \6048_b0 , w_22067 );
and ( w_22066 , w_22067 , \5850_b0 );
or ( \8793_b1 , \8791_b1 , w_22069 );
not ( w_22069 , w_22070 );
and ( \8793_b0 , \8791_b0 , w_22071 );
and ( w_22070 ,  , w_22071 );
buf ( w_22069 , \8792_b1 );
not ( w_22069 , w_22072 );
not (  , w_22073 );
and ( w_22072 , w_22073 , \8792_b0 );
or ( \8794_b1 , \8793_b1 , w_22074 );
xor ( \8794_b0 , \8793_b0 , w_22076 );
not ( w_22076 , w_22077 );
and ( w_22077 , w_22074 , w_22075 );
buf ( w_22074 , \5859_b1 );
not ( w_22074 , w_22078 );
not ( w_22075 , w_22079 );
and ( w_22078 , w_22079 , \5859_b0 );
or ( \8795_b1 , \8790_b1 , \8794_b1 );
xor ( \8795_b0 , \8790_b0 , w_22080 );
not ( w_22080 , w_22081 );
and ( w_22081 , \8794_b1 , \8794_b0 );
or ( \8796_b1 , \5998_b1 , \5768_b1 );
not ( \5768_b1 , w_22082 );
and ( \8796_b0 , \5998_b0 , w_22083 );
and ( w_22082 , w_22083 , \5768_b0 );
or ( \8797_b1 , \5967_b1 , \5766_b1 );
not ( \5766_b1 , w_22084 );
and ( \8797_b0 , \5967_b0 , w_22085 );
and ( w_22084 , w_22085 , \5766_b0 );
or ( \8798_b1 , \8796_b1 , w_22087 );
not ( w_22087 , w_22088 );
and ( \8798_b0 , \8796_b0 , w_22089 );
and ( w_22088 ,  , w_22089 );
buf ( w_22087 , \8797_b1 );
not ( w_22087 , w_22090 );
not (  , w_22091 );
and ( w_22090 , w_22091 , \8797_b0 );
or ( \8799_b1 , \8798_b1 , w_22092 );
xor ( \8799_b0 , \8798_b0 , w_22094 );
not ( w_22094 , w_22095 );
and ( w_22095 , w_22092 , w_22093 );
buf ( w_22092 , \5775_b1 );
not ( w_22092 , w_22096 );
not ( w_22093 , w_22097 );
and ( w_22096 , w_22097 , \5775_b0 );
or ( \8800_b1 , \6018_b1 , \5790_b1 );
not ( \5790_b1 , w_22098 );
and ( \8800_b0 , \6018_b0 , w_22099 );
and ( w_22098 , w_22099 , \5790_b0 );
or ( \8801_b1 , \5986_b1 , \5788_b1 );
not ( \5788_b1 , w_22100 );
and ( \8801_b0 , \5986_b0 , w_22101 );
and ( w_22100 , w_22101 , \5788_b0 );
or ( \8802_b1 , \8800_b1 , w_22103 );
not ( w_22103 , w_22104 );
and ( \8802_b0 , \8800_b0 , w_22105 );
and ( w_22104 ,  , w_22105 );
buf ( w_22103 , \8801_b1 );
not ( w_22103 , w_22106 );
not (  , w_22107 );
and ( w_22106 , w_22107 , \8801_b0 );
or ( \8803_b1 , \8802_b1 , w_22108 );
xor ( \8803_b0 , \8802_b0 , w_22110 );
not ( w_22110 , w_22111 );
and ( w_22111 , w_22108 , w_22109 );
buf ( w_22108 , \5797_b1 );
not ( w_22108 , w_22112 );
not ( w_22109 , w_22113 );
and ( w_22112 , w_22113 , \5797_b0 );
or ( \8804_b1 , \8799_b1 , \8803_b1 );
xor ( \8804_b0 , \8799_b0 , w_22114 );
not ( w_22114 , w_22115 );
and ( w_22115 , \8803_b1 , \8803_b0 );
or ( \8805_b1 , \6041_b1 , \5809_b1 );
not ( \5809_b1 , w_22116 );
and ( \8805_b0 , \6041_b0 , w_22117 );
and ( w_22116 , w_22117 , \5809_b0 );
or ( \8806_b1 , \6006_b1 , \5807_b1 );
not ( \5807_b1 , w_22118 );
and ( \8806_b0 , \6006_b0 , w_22119 );
and ( w_22118 , w_22119 , \5807_b0 );
or ( \8807_b1 , \8805_b1 , w_22121 );
not ( w_22121 , w_22122 );
and ( \8807_b0 , \8805_b0 , w_22123 );
and ( w_22122 ,  , w_22123 );
buf ( w_22121 , \8806_b1 );
not ( w_22121 , w_22124 );
not (  , w_22125 );
and ( w_22124 , w_22125 , \8806_b0 );
or ( \8808_b1 , \8807_b1 , w_22126 );
xor ( \8808_b0 , \8807_b0 , w_22128 );
not ( w_22128 , w_22129 );
and ( w_22129 , w_22126 , w_22127 );
buf ( w_22126 , \5816_b1 );
not ( w_22126 , w_22130 );
not ( w_22127 , w_22131 );
and ( w_22130 , w_22131 , \5816_b0 );
or ( \8809_b1 , \8804_b1 , \8808_b1 );
xor ( \8809_b0 , \8804_b0 , w_22132 );
not ( w_22132 , w_22133 );
and ( w_22133 , \8808_b1 , \8808_b0 );
or ( \8810_b1 , \8795_b1 , \8809_b1 );
xor ( \8810_b0 , \8795_b0 , w_22134 );
not ( w_22134 , w_22135 );
and ( w_22135 , \8809_b1 , \8809_b0 );
or ( \8811_b1 , \5937_b1 , \7192_b1 );
not ( \7192_b1 , w_22136 );
and ( \8811_b0 , \5937_b0 , w_22137 );
and ( w_22136 , w_22137 , \7192_b0 );
or ( \8812_b1 , \5906_b1 , \7190_b1 );
not ( \7190_b1 , w_22138 );
and ( \8812_b0 , \5906_b0 , w_22139 );
and ( w_22138 , w_22139 , \7190_b0 );
or ( \8813_b1 , \8811_b1 , w_22141 );
not ( w_22141 , w_22142 );
and ( \8813_b0 , \8811_b0 , w_22143 );
and ( w_22142 ,  , w_22143 );
buf ( w_22141 , \8812_b1 );
not ( w_22141 , w_22144 );
not (  , w_22145 );
and ( w_22144 , w_22145 , \8812_b0 );
or ( \8814_b1 , \8813_b1 , w_22146 );
xor ( \8814_b0 , \8813_b0 , w_22148 );
not ( w_22148 , w_22149 );
and ( w_22149 , w_22146 , w_22147 );
buf ( w_22146 , \7198_b1 );
not ( w_22146 , w_22150 );
not ( w_22147 , w_22151 );
and ( w_22150 , w_22151 , \7198_b0 );
or ( \8815_b1 , \5957_b1 , \7203_b1 );
not ( \7203_b1 , w_22152 );
and ( \8815_b0 , \5957_b0 , w_22153 );
and ( w_22152 , w_22153 , \7203_b0 );
or ( \8816_b1 , \5925_b1 , \7201_b1 );
not ( \7201_b1 , w_22154 );
and ( \8816_b0 , \5925_b0 , w_22155 );
and ( w_22154 , w_22155 , \7201_b0 );
or ( \8817_b1 , \8815_b1 , w_22157 );
not ( w_22157 , w_22158 );
and ( \8817_b0 , \8815_b0 , w_22159 );
and ( w_22158 ,  , w_22159 );
buf ( w_22157 , \8816_b1 );
not ( w_22157 , w_22160 );
not (  , w_22161 );
and ( w_22160 , w_22161 , \8816_b0 );
or ( \8818_b1 , \8817_b1 , w_22162 );
xor ( \8818_b0 , \8817_b0 , w_22164 );
not ( w_22164 , w_22165 );
and ( w_22165 , w_22162 , w_22163 );
buf ( w_22162 , \6824_b1 );
not ( w_22162 , w_22166 );
not ( w_22163 , w_22167 );
and ( w_22166 , w_22167 , \6824_b0 );
or ( \8819_b1 , \8814_b1 , \8818_b1 );
xor ( \8819_b0 , \8814_b0 , w_22168 );
not ( w_22168 , w_22169 );
and ( w_22169 , \8818_b1 , \8818_b0 );
or ( \8820_b1 , \5979_b1 , \5750_b1 );
not ( \5750_b1 , w_22170 );
and ( \8820_b0 , \5979_b0 , w_22171 );
and ( w_22170 , w_22171 , \5750_b0 );
or ( \8821_b1 , \5945_b1 , \5748_b1 );
not ( \5748_b1 , w_22172 );
and ( \8821_b0 , \5945_b0 , w_22173 );
and ( w_22172 , w_22173 , \5748_b0 );
or ( \8822_b1 , \8820_b1 , w_22175 );
not ( w_22175 , w_22176 );
and ( \8822_b0 , \8820_b0 , w_22177 );
and ( w_22176 ,  , w_22177 );
buf ( w_22175 , \8821_b1 );
not ( w_22175 , w_22178 );
not (  , w_22179 );
and ( w_22178 , w_22179 , \8821_b0 );
or ( \8823_b1 , \8822_b1 , w_22180 );
xor ( \8823_b0 , \8822_b0 , w_22182 );
not ( w_22182 , w_22183 );
and ( w_22183 , w_22180 , w_22181 );
buf ( w_22180 , \5755_b1 );
not ( w_22180 , w_22184 );
not ( w_22181 , w_22185 );
and ( w_22184 , w_22185 , \5755_b0 );
or ( \8824_b1 , \8819_b1 , \8823_b1 );
xor ( \8824_b0 , \8819_b0 , w_22186 );
not ( w_22186 , w_22187 );
and ( w_22187 , \8823_b1 , \8823_b0 );
or ( \8825_b1 , \8810_b1 , \8824_b1 );
xor ( \8825_b0 , \8810_b0 , w_22188 );
not ( w_22188 , w_22189 );
and ( w_22189 , \8824_b1 , \8824_b0 );
or ( \8826_b1 , \8786_b1 , \8825_b1 );
xor ( \8826_b0 , \8786_b0 , w_22190 );
not ( w_22190 , w_22191 );
and ( w_22191 , \8825_b1 , \8825_b0 );
or ( \8827_b1 , \8740_b1 , \8826_b1 );
xor ( \8827_b0 , \8740_b0 , w_22192 );
not ( w_22192 , w_22193 );
and ( w_22193 , \8826_b1 , \8826_b0 );
or ( \8828_b1 , \8589_b1 , \8593_b1 );
not ( \8593_b1 , w_22194 );
and ( \8828_b0 , \8589_b0 , w_22195 );
and ( w_22194 , w_22195 , \8593_b0 );
or ( \8829_b1 , \8593_b1 , \8598_b1 );
not ( \8598_b1 , w_22196 );
and ( \8829_b0 , \8593_b0 , w_22197 );
and ( w_22196 , w_22197 , \8598_b0 );
or ( \8830_b1 , \8589_b1 , \8598_b1 );
not ( \8598_b1 , w_22198 );
and ( \8830_b0 , \8589_b0 , w_22199 );
and ( w_22198 , w_22199 , \8598_b0 );
or ( \8832_b1 , \8577_b1 , \8581_b1 );
not ( \8581_b1 , w_22200 );
and ( \8832_b0 , \8577_b0 , w_22201 );
and ( w_22200 , w_22201 , \8581_b0 );
or ( \8833_b1 , \8581_b1 , \8583_b1 );
not ( \8583_b1 , w_22202 );
and ( \8833_b0 , \8581_b0 , w_22203 );
and ( w_22202 , w_22203 , \8583_b0 );
or ( \8834_b1 , \8577_b1 , \8583_b1 );
not ( \8583_b1 , w_22204 );
and ( \8834_b0 , \8577_b0 , w_22205 );
and ( w_22204 , w_22205 , \8583_b0 );
or ( \8836_b1 , \8831_b1 , \8835_b1 );
xor ( \8836_b0 , \8831_b0 , w_22206 );
not ( w_22206 , w_22207 );
and ( w_22207 , \8835_b1 , \8835_b0 );
or ( \8837_b1 , \8558_b1 , w_22208 );
or ( \8837_b0 , \8558_b0 , \8572_b0 );
not ( \8572_b0 , w_22209 );
and ( w_22209 , w_22208 , \8572_b1 );
or ( \8838_b1 , \8836_b1 , \8837_b1 );
xor ( \8838_b0 , \8836_b0 , w_22210 );
not ( w_22210 , w_22211 );
and ( w_22211 , \8837_b1 , \8837_b0 );
or ( \8839_b1 , \8827_b1 , \8838_b1 );
xor ( \8839_b0 , \8827_b0 , w_22212 );
not ( w_22212 , w_22213 );
and ( w_22213 , \8838_b1 , \8838_b0 );
or ( \8840_b1 , \8711_b1 , \8839_b1 );
xor ( \8840_b0 , \8711_b0 , w_22214 );
not ( w_22214 , w_22215 );
and ( w_22215 , \8839_b1 , \8839_b0 );
or ( \8841_b1 , \8702_b1 , \8840_b1 );
xor ( \8841_b0 , \8702_b0 , w_22216 );
not ( w_22216 , w_22217 );
and ( w_22217 , \8840_b1 , \8840_b0 );
or ( \8842_b1 , \8525_b1 , \8536_b1 );
not ( \8536_b1 , w_22218 );
and ( \8842_b0 , \8525_b0 , w_22219 );
and ( w_22218 , w_22219 , \8536_b0 );
or ( \8843_b1 , \8536_b1 , \8676_b1 );
not ( \8676_b1 , w_22220 );
and ( \8843_b0 , \8536_b0 , w_22221 );
and ( w_22220 , w_22221 , \8676_b0 );
or ( \8844_b1 , \8525_b1 , \8676_b1 );
not ( \8676_b1 , w_22222 );
and ( \8844_b0 , \8525_b0 , w_22223 );
and ( w_22222 , w_22223 , \8676_b0 );
or ( \8846_b1 , \8841_b1 , w_22225 );
not ( w_22225 , w_22226 );
and ( \8846_b0 , \8841_b0 , w_22227 );
and ( w_22226 ,  , w_22227 );
buf ( w_22225 , \8845_b1 );
not ( w_22225 , w_22228 );
not (  , w_22229 );
and ( w_22228 , w_22229 , \8845_b0 );
or ( \8847_b1 , \8706_b1 , \8710_b1 );
not ( \8710_b1 , w_22230 );
and ( \8847_b0 , \8706_b0 , w_22231 );
and ( w_22230 , w_22231 , \8710_b0 );
or ( \8848_b1 , \8710_b1 , \8839_b1 );
not ( \8839_b1 , w_22232 );
and ( \8848_b0 , \8710_b0 , w_22233 );
and ( w_22232 , w_22233 , \8839_b0 );
or ( \8849_b1 , \8706_b1 , \8839_b1 );
not ( \8839_b1 , w_22234 );
and ( \8849_b0 , \8706_b0 , w_22235 );
and ( w_22234 , w_22235 , \8839_b0 );
or ( \8851_b1 , \8831_b1 , \8835_b1 );
not ( \8835_b1 , w_22236 );
and ( \8851_b0 , \8831_b0 , w_22237 );
and ( w_22236 , w_22237 , \8835_b0 );
or ( \8852_b1 , \8835_b1 , \8837_b1 );
not ( \8837_b1 , w_22238 );
and ( \8852_b0 , \8835_b0 , w_22239 );
and ( w_22238 , w_22239 , \8837_b0 );
or ( \8853_b1 , \8831_b1 , \8837_b1 );
not ( \8837_b1 , w_22240 );
and ( \8853_b0 , \8831_b0 , w_22241 );
and ( w_22240 , w_22241 , \8837_b0 );
or ( \8855_b1 , \8744_b1 , \8785_b1 );
not ( \8785_b1 , w_22242 );
and ( \8855_b0 , \8744_b0 , w_22243 );
and ( w_22242 , w_22243 , \8785_b0 );
or ( \8856_b1 , \8785_b1 , \8825_b1 );
not ( \8825_b1 , w_22244 );
and ( \8856_b0 , \8785_b0 , w_22245 );
and ( w_22244 , w_22245 , \8825_b0 );
or ( \8857_b1 , \8744_b1 , \8825_b1 );
not ( \8825_b1 , w_22246 );
and ( \8857_b0 , \8744_b0 , w_22247 );
and ( w_22246 , w_22247 , \8825_b0 );
or ( \8859_b1 , \8854_b1 , \8858_b1 );
xor ( \8859_b0 , \8854_b0 , w_22248 );
not ( w_22248 , w_22249 );
and ( w_22249 , \8858_b1 , \8858_b0 );
or ( \8860_b1 , \8725_b1 , \8739_b1 );
not ( \8739_b1 , w_22250 );
and ( \8860_b0 , \8725_b0 , w_22251 );
and ( w_22250 , w_22251 , \8739_b0 );
or ( \8861_b1 , \8859_b1 , \8860_b1 );
xor ( \8861_b0 , \8859_b0 , w_22252 );
not ( w_22252 , w_22253 );
and ( w_22253 , \8860_b1 , \8860_b0 );
or ( \8862_b1 , \8850_b1 , \8861_b1 );
xor ( \8862_b0 , \8850_b0 , w_22254 );
not ( w_22254 , w_22255 );
and ( w_22255 , \8861_b1 , \8861_b0 );
or ( \8863_b1 , \8691_b1 , \8695_b1 );
not ( \8695_b1 , w_22256 );
and ( \8863_b0 , \8691_b0 , w_22257 );
and ( w_22256 , w_22257 , \8695_b0 );
or ( \8864_b1 , \8695_b1 , \8700_b1 );
not ( \8700_b1 , w_22258 );
and ( \8864_b0 , \8695_b0 , w_22259 );
and ( w_22258 , w_22259 , \8700_b0 );
or ( \8865_b1 , \8691_b1 , \8700_b1 );
not ( \8700_b1 , w_22260 );
and ( \8865_b0 , \8691_b0 , w_22261 );
and ( w_22260 , w_22261 , \8700_b0 );
or ( \8867_b1 , \8740_b1 , \8826_b1 );
not ( \8826_b1 , w_22262 );
and ( \8867_b0 , \8740_b0 , w_22263 );
and ( w_22262 , w_22263 , \8826_b0 );
or ( \8868_b1 , \8826_b1 , \8838_b1 );
not ( \8838_b1 , w_22264 );
and ( \8868_b0 , \8826_b0 , w_22265 );
and ( w_22264 , w_22265 , \8838_b0 );
or ( \8869_b1 , \8740_b1 , \8838_b1 );
not ( \8838_b1 , w_22266 );
and ( \8869_b0 , \8740_b0 , w_22267 );
and ( w_22266 , w_22267 , \8838_b0 );
or ( \8871_b1 , \8866_b1 , \8870_b1 );
xor ( \8871_b0 , \8866_b0 , w_22268 );
not ( w_22268 , w_22269 );
and ( w_22269 , \8870_b1 , \8870_b0 );
or ( \8872_b1 , \6029_b1 , \5829_b1 );
not ( \5829_b1 , w_22270 );
and ( \8872_b0 , \6029_b0 , w_22271 );
and ( w_22270 , w_22271 , \5829_b0 );
or ( \8873_b1 , \6041_b1 , \5827_b1 );
not ( \5827_b1 , w_22272 );
and ( \8873_b0 , \6041_b0 , w_22273 );
and ( w_22272 , w_22273 , \5827_b0 );
or ( \8874_b1 , \8872_b1 , w_22275 );
not ( w_22275 , w_22276 );
and ( \8874_b0 , \8872_b0 , w_22277 );
and ( w_22276 ,  , w_22277 );
buf ( w_22275 , \8873_b1 );
not ( w_22275 , w_22278 );
not (  , w_22279 );
and ( w_22278 , w_22279 , \8873_b0 );
or ( \8875_b1 , \8874_b1 , w_22280 );
xor ( \8875_b0 , \8874_b0 , w_22282 );
not ( w_22282 , w_22283 );
and ( w_22283 , w_22280 , w_22281 );
buf ( w_22280 , \5836_b1 );
not ( w_22280 , w_22284 );
not ( w_22281 , w_22285 );
and ( w_22284 , w_22285 , \5836_b0 );
or ( \8876_b1 , \6048_b1 , \5852_b1 );
not ( \5852_b1 , w_22286 );
and ( \8876_b0 , \6048_b0 , w_22287 );
and ( w_22286 , w_22287 , \5852_b0 );
or ( \8877_b1 , \6057_b1 , \5850_b1 );
not ( \5850_b1 , w_22288 );
and ( \8877_b0 , \6057_b0 , w_22289 );
and ( w_22288 , w_22289 , \5850_b0 );
or ( \8878_b1 , \8876_b1 , w_22291 );
not ( w_22291 , w_22292 );
and ( \8878_b0 , \8876_b0 , w_22293 );
and ( w_22292 ,  , w_22293 );
buf ( w_22291 , \8877_b1 );
not ( w_22291 , w_22294 );
not (  , w_22295 );
and ( w_22294 , w_22295 , \8877_b0 );
or ( \8879_b1 , \8878_b1 , w_22296 );
xor ( \8879_b0 , \8878_b0 , w_22298 );
not ( w_22298 , w_22299 );
and ( w_22299 , w_22296 , w_22297 );
buf ( w_22296 , \5859_b1 );
not ( w_22296 , w_22300 );
not ( w_22297 , w_22301 );
and ( w_22300 , w_22301 , \5859_b0 );
or ( \8880_b1 , \8875_b1 , \8879_b1 );
xor ( \8880_b0 , \8875_b0 , w_22302 );
not ( w_22302 , w_22303 );
and ( w_22303 , \8879_b1 , \8879_b0 );
or ( \8881_b1 , \6065_b1 , w_22305 );
not ( w_22305 , w_22306 );
and ( \8881_b0 , \6065_b0 , w_22307 );
and ( w_22306 ,  , w_22307 );
buf ( w_22305 , \5869_b1 );
not ( w_22305 , w_22308 );
not (  , w_22309 );
and ( w_22308 , w_22309 , \5869_b0 );
or ( \8882_b1 , \8881_b1 , w_22310 );
xor ( \8882_b0 , \8881_b0 , w_22312 );
not ( w_22312 , w_22313 );
and ( w_22313 , w_22310 , w_22311 );
buf ( w_22310 , \5878_b1 );
not ( w_22310 , w_22314 );
not ( w_22311 , w_22315 );
and ( w_22314 , w_22315 , \5878_b0 );
or ( \8883_b1 , \8880_b1 , \8882_b1 );
xor ( \8883_b0 , \8880_b0 , w_22316 );
not ( w_22316 , w_22317 );
and ( w_22317 , \8882_b1 , \8882_b0 );
or ( \8884_b1 , \5967_b1 , \5768_b1 );
not ( \5768_b1 , w_22318 );
and ( \8884_b0 , \5967_b0 , w_22319 );
and ( w_22318 , w_22319 , \5768_b0 );
or ( \8885_b1 , \5979_b1 , \5766_b1 );
not ( \5766_b1 , w_22320 );
and ( \8885_b0 , \5979_b0 , w_22321 );
and ( w_22320 , w_22321 , \5766_b0 );
or ( \8886_b1 , \8884_b1 , w_22323 );
not ( w_22323 , w_22324 );
and ( \8886_b0 , \8884_b0 , w_22325 );
and ( w_22324 ,  , w_22325 );
buf ( w_22323 , \8885_b1 );
not ( w_22323 , w_22326 );
not (  , w_22327 );
and ( w_22326 , w_22327 , \8885_b0 );
or ( \8887_b1 , \8886_b1 , w_22328 );
xor ( \8887_b0 , \8886_b0 , w_22330 );
not ( w_22330 , w_22331 );
and ( w_22331 , w_22328 , w_22329 );
buf ( w_22328 , \5775_b1 );
not ( w_22328 , w_22332 );
not ( w_22329 , w_22333 );
and ( w_22332 , w_22333 , \5775_b0 );
or ( \8888_b1 , \5986_b1 , \5790_b1 );
not ( \5790_b1 , w_22334 );
and ( \8888_b0 , \5986_b0 , w_22335 );
and ( w_22334 , w_22335 , \5790_b0 );
or ( \8889_b1 , \5998_b1 , \5788_b1 );
not ( \5788_b1 , w_22336 );
and ( \8889_b0 , \5998_b0 , w_22337 );
and ( w_22336 , w_22337 , \5788_b0 );
or ( \8890_b1 , \8888_b1 , w_22339 );
not ( w_22339 , w_22340 );
and ( \8890_b0 , \8888_b0 , w_22341 );
and ( w_22340 ,  , w_22341 );
buf ( w_22339 , \8889_b1 );
not ( w_22339 , w_22342 );
not (  , w_22343 );
and ( w_22342 , w_22343 , \8889_b0 );
or ( \8891_b1 , \8890_b1 , w_22344 );
xor ( \8891_b0 , \8890_b0 , w_22346 );
not ( w_22346 , w_22347 );
and ( w_22347 , w_22344 , w_22345 );
buf ( w_22344 , \5797_b1 );
not ( w_22344 , w_22348 );
not ( w_22345 , w_22349 );
and ( w_22348 , w_22349 , \5797_b0 );
or ( \8892_b1 , \8887_b1 , \8891_b1 );
xor ( \8892_b0 , \8887_b0 , w_22350 );
not ( w_22350 , w_22351 );
and ( w_22351 , \8891_b1 , \8891_b0 );
or ( \8893_b1 , \6006_b1 , \5809_b1 );
not ( \5809_b1 , w_22352 );
and ( \8893_b0 , \6006_b0 , w_22353 );
and ( w_22352 , w_22353 , \5809_b0 );
or ( \8894_b1 , \6018_b1 , \5807_b1 );
not ( \5807_b1 , w_22354 );
and ( \8894_b0 , \6018_b0 , w_22355 );
and ( w_22354 , w_22355 , \5807_b0 );
or ( \8895_b1 , \8893_b1 , w_22357 );
not ( w_22357 , w_22358 );
and ( \8895_b0 , \8893_b0 , w_22359 );
and ( w_22358 ,  , w_22359 );
buf ( w_22357 , \8894_b1 );
not ( w_22357 , w_22360 );
not (  , w_22361 );
and ( w_22360 , w_22361 , \8894_b0 );
or ( \8896_b1 , \8895_b1 , w_22362 );
xor ( \8896_b0 , \8895_b0 , w_22364 );
not ( w_22364 , w_22365 );
and ( w_22365 , w_22362 , w_22363 );
buf ( w_22362 , \5816_b1 );
not ( w_22362 , w_22366 );
not ( w_22363 , w_22367 );
and ( w_22366 , w_22367 , \5816_b0 );
or ( \8897_b1 , \8892_b1 , \8896_b1 );
xor ( \8897_b0 , \8892_b0 , w_22368 );
not ( w_22368 , w_22369 );
and ( w_22369 , \8896_b1 , \8896_b0 );
or ( \8898_b1 , \8883_b1 , w_22370 );
xor ( \8898_b0 , \8883_b0 , w_22372 );
not ( w_22372 , w_22373 );
and ( w_22373 , w_22370 , w_22371 );
buf ( w_22370 , \8897_b1 );
not ( w_22370 , w_22374 );
not ( w_22371 , w_22375 );
and ( w_22374 , w_22375 , \8897_b0 );
or ( \8899_b1 , \8814_b1 , \8818_b1 );
not ( \8818_b1 , w_22376 );
and ( \8899_b0 , \8814_b0 , w_22377 );
and ( w_22376 , w_22377 , \8818_b0 );
or ( \8900_b1 , \8818_b1 , \8823_b1 );
not ( \8823_b1 , w_22378 );
and ( \8900_b0 , \8818_b0 , w_22379 );
and ( w_22378 , w_22379 , \8823_b0 );
or ( \8901_b1 , \8814_b1 , \8823_b1 );
not ( \8823_b1 , w_22380 );
and ( \8901_b0 , \8814_b0 , w_22381 );
and ( w_22380 , w_22381 , \8823_b0 );
or ( \8903_b1 , \8799_b1 , \8803_b1 );
not ( \8803_b1 , w_22382 );
and ( \8903_b0 , \8799_b0 , w_22383 );
and ( w_22382 , w_22383 , \8803_b0 );
or ( \8904_b1 , \8803_b1 , \8808_b1 );
not ( \8808_b1 , w_22384 );
and ( \8904_b0 , \8803_b0 , w_22385 );
and ( w_22384 , w_22385 , \8808_b0 );
or ( \8905_b1 , \8799_b1 , \8808_b1 );
not ( \8808_b1 , w_22386 );
and ( \8905_b0 , \8799_b0 , w_22387 );
and ( w_22386 , w_22387 , \8808_b0 );
or ( \8907_b1 , \8902_b1 , \8906_b1 );
xor ( \8907_b0 , \8902_b0 , w_22388 );
not ( w_22388 , w_22389 );
and ( w_22389 , \8906_b1 , \8906_b0 );
or ( \8908_b1 , \8790_b1 , \8794_b1 );
not ( \8794_b1 , w_22390 );
and ( \8908_b0 , \8790_b0 , w_22391 );
and ( w_22390 , w_22391 , \8794_b0 );
or ( \8909_b1 , \8907_b1 , \8908_b1 );
xor ( \8909_b0 , \8907_b0 , w_22392 );
not ( w_22392 , w_22393 );
and ( w_22393 , \8908_b1 , \8908_b0 );
or ( \8910_b1 , \8898_b1 , \8909_b1 );
xor ( \8910_b0 , \8898_b0 , w_22394 );
not ( w_22394 , w_22395 );
and ( w_22395 , \8909_b1 , \8909_b0 );
or ( \8911_b1 , \8774_b1 , \8778_b1 );
not ( \8778_b1 , w_22396 );
and ( \8911_b0 , \8774_b0 , w_22397 );
and ( w_22396 , w_22397 , \8778_b0 );
or ( \8912_b1 , \8778_b1 , \8783_b1 );
not ( \8783_b1 , w_22398 );
and ( \8912_b0 , \8778_b0 , w_22399 );
and ( w_22398 , w_22399 , \8783_b0 );
or ( \8913_b1 , \8774_b1 , \8783_b1 );
not ( \8783_b1 , w_22400 );
and ( \8913_b0 , \8774_b0 , w_22401 );
and ( w_22400 , w_22401 , \8783_b0 );
or ( \8915_b1 , \8762_b1 , \8766_b1 );
not ( \8766_b1 , w_22402 );
and ( \8915_b0 , \8762_b0 , w_22403 );
and ( w_22402 , w_22403 , \8766_b0 );
or ( \8916_b1 , \8766_b1 , \8771_b1 );
not ( \8771_b1 , w_22404 );
and ( \8916_b0 , \8766_b0 , w_22405 );
and ( w_22404 , w_22405 , \8771_b0 );
or ( \8917_b1 , \8762_b1 , \8771_b1 );
not ( \8771_b1 , w_22406 );
and ( \8917_b0 , \8762_b0 , w_22407 );
and ( w_22406 , w_22407 , \8771_b0 );
or ( \8919_b1 , \8914_b1 , \8918_b1 );
xor ( \8919_b0 , \8914_b0 , w_22408 );
not ( w_22408 , w_22409 );
and ( w_22409 , \8918_b1 , \8918_b0 );
or ( \8920_b1 , \8748_b1 , \8752_b1 );
not ( \8752_b1 , w_22410 );
and ( \8920_b0 , \8748_b0 , w_22411 );
and ( w_22410 , w_22411 , \8752_b0 );
or ( \8921_b1 , \8752_b1 , \8757_b1 );
not ( \8757_b1 , w_22412 );
and ( \8921_b0 , \8752_b0 , w_22413 );
and ( w_22412 , w_22413 , \8757_b0 );
or ( \8922_b1 , \8748_b1 , \8757_b1 );
not ( \8757_b1 , w_22414 );
and ( \8922_b0 , \8748_b0 , w_22415 );
and ( w_22414 , w_22415 , \8757_b0 );
or ( \8924_b1 , \8919_b1 , \8923_b1 );
xor ( \8924_b0 , \8919_b0 , w_22416 );
not ( w_22416 , w_22417 );
and ( w_22417 , \8923_b1 , \8923_b0 );
or ( \8925_b1 , \8910_b1 , \8924_b1 );
xor ( \8925_b0 , \8910_b0 , w_22418 );
not ( w_22418 , w_22419 );
and ( w_22419 , \8924_b1 , \8924_b0 );
or ( \8926_b1 , \8758_b1 , \8772_b1 );
not ( \8772_b1 , w_22420 );
and ( \8926_b0 , \8758_b0 , w_22421 );
and ( w_22420 , w_22421 , \8772_b0 );
or ( \8927_b1 , \8772_b1 , \8784_b1 );
not ( \8784_b1 , w_22422 );
and ( \8927_b0 , \8772_b0 , w_22423 );
and ( w_22422 , w_22423 , \8784_b0 );
or ( \8928_b1 , \8758_b1 , \8784_b1 );
not ( \8784_b1 , w_22424 );
and ( \8928_b0 , \8758_b0 , w_22425 );
and ( w_22424 , w_22425 , \8784_b0 );
or ( \8930_b1 , \5737_b1 , \7043_b1 );
not ( \7043_b1 , w_22426 );
and ( \8930_b0 , \5737_b0 , w_22427 );
and ( w_22426 , w_22427 , \7043_b0 );
buf ( \8931_b1 , \8930_b1 );
not ( \8931_b1 , w_22428 );
not ( \8931_b0 , w_22429 );
and ( w_22428 , w_22429 , \8930_b0 );
or ( \8932_b1 , \8931_b1 , w_22430 );
xor ( \8932_b0 , \8931_b0 , w_22432 );
not ( w_22432 , w_22433 );
and ( w_22433 , w_22430 , w_22431 );
buf ( w_22430 , \7049_b1 );
not ( w_22430 , w_22434 );
not ( w_22431 , w_22435 );
and ( w_22434 , w_22435 , \7049_b0 );
or ( \8933_b1 , \5878_b1 , \8932_b1 );
xor ( \8933_b0 , \5878_b0 , w_22436 );
not ( w_22436 , w_22437 );
and ( w_22437 , \8932_b1 , \8932_b0 );
or ( \8934_b1 , \5758_b1 , \7061_b1 );
not ( \7061_b1 , w_22438 );
and ( \8934_b0 , \5758_b0 , w_22439 );
and ( w_22438 , w_22439 , \7061_b0 );
or ( \8935_b1 , \5770_b1 , \7059_b1 );
not ( \7059_b1 , w_22440 );
and ( \8935_b0 , \5770_b0 , w_22441 );
and ( w_22440 , w_22441 , \7059_b0 );
or ( \8936_b1 , \8934_b1 , w_22443 );
not ( w_22443 , w_22444 );
and ( \8936_b0 , \8934_b0 , w_22445 );
and ( w_22444 ,  , w_22445 );
buf ( w_22443 , \8935_b1 );
not ( w_22443 , w_22446 );
not (  , w_22447 );
and ( w_22446 , w_22447 , \8935_b0 );
or ( \8937_b1 , \8936_b1 , w_22448 );
xor ( \8937_b0 , \8936_b0 , w_22450 );
not ( w_22450 , w_22451 );
and ( w_22451 , w_22448 , w_22449 );
buf ( w_22448 , \7067_b1 );
not ( w_22448 , w_22452 );
not ( w_22449 , w_22453 );
and ( w_22452 , w_22453 , \7067_b0 );
or ( \8938_b1 , \8933_b1 , \8937_b1 );
xor ( \8938_b0 , \8933_b0 , w_22454 );
not ( w_22454 , w_22455 );
and ( w_22455 , \8937_b1 , \8937_b0 );
or ( \8939_b1 , \8929_b1 , \8938_b1 );
xor ( \8939_b0 , \8929_b0 , w_22456 );
not ( w_22456 , w_22457 );
and ( w_22457 , \8938_b1 , \8938_b0 );
or ( \8940_b1 , \5906_b1 , \7192_b1 );
not ( \7192_b1 , w_22458 );
and ( \8940_b0 , \5906_b0 , w_22459 );
and ( w_22458 , w_22459 , \7192_b0 );
or ( \8941_b1 , \5918_b1 , \7190_b1 );
not ( \7190_b1 , w_22460 );
and ( \8941_b0 , \5918_b0 , w_22461 );
and ( w_22460 , w_22461 , \7190_b0 );
or ( \8942_b1 , \8940_b1 , w_22463 );
not ( w_22463 , w_22464 );
and ( \8942_b0 , \8940_b0 , w_22465 );
and ( w_22464 ,  , w_22465 );
buf ( w_22463 , \8941_b1 );
not ( w_22463 , w_22466 );
not (  , w_22467 );
and ( w_22466 , w_22467 , \8941_b0 );
or ( \8943_b1 , \8942_b1 , w_22468 );
xor ( \8943_b0 , \8942_b0 , w_22470 );
not ( w_22470 , w_22471 );
and ( w_22471 , w_22468 , w_22469 );
buf ( w_22468 , \7198_b1 );
not ( w_22468 , w_22472 );
not ( w_22469 , w_22473 );
and ( w_22472 , w_22473 , \7198_b0 );
or ( \8944_b1 , \5925_b1 , \7203_b1 );
not ( \7203_b1 , w_22474 );
and ( \8944_b0 , \5925_b0 , w_22475 );
and ( w_22474 , w_22475 , \7203_b0 );
or ( \8945_b1 , \5937_b1 , \7201_b1 );
not ( \7201_b1 , w_22476 );
and ( \8945_b0 , \5937_b0 , w_22477 );
and ( w_22476 , w_22477 , \7201_b0 );
or ( \8946_b1 , \8944_b1 , w_22479 );
not ( w_22479 , w_22480 );
and ( \8946_b0 , \8944_b0 , w_22481 );
and ( w_22480 ,  , w_22481 );
buf ( w_22479 , \8945_b1 );
not ( w_22479 , w_22482 );
not (  , w_22483 );
and ( w_22482 , w_22483 , \8945_b0 );
or ( \8947_b1 , \8946_b1 , w_22484 );
xor ( \8947_b0 , \8946_b0 , w_22486 );
not ( w_22486 , w_22487 );
and ( w_22487 , w_22484 , w_22485 );
buf ( w_22484 , \6824_b1 );
not ( w_22484 , w_22488 );
not ( w_22485 , w_22489 );
and ( w_22488 , w_22489 , \6824_b0 );
or ( \8948_b1 , \8943_b1 , \8947_b1 );
xor ( \8948_b0 , \8943_b0 , w_22490 );
not ( w_22490 , w_22491 );
and ( w_22491 , \8947_b1 , \8947_b0 );
or ( \8949_b1 , \5945_b1 , \5750_b1 );
not ( \5750_b1 , w_22492 );
and ( \8949_b0 , \5945_b0 , w_22493 );
and ( w_22492 , w_22493 , \5750_b0 );
or ( \8950_b1 , \5957_b1 , \5748_b1 );
not ( \5748_b1 , w_22494 );
and ( \8950_b0 , \5957_b0 , w_22495 );
and ( w_22494 , w_22495 , \5748_b0 );
or ( \8951_b1 , \8949_b1 , w_22497 );
not ( w_22497 , w_22498 );
and ( \8951_b0 , \8949_b0 , w_22499 );
and ( w_22498 ,  , w_22499 );
buf ( w_22497 , \8950_b1 );
not ( w_22497 , w_22500 );
not (  , w_22501 );
and ( w_22500 , w_22501 , \8950_b0 );
or ( \8952_b1 , \8951_b1 , w_22502 );
xor ( \8952_b0 , \8951_b0 , w_22504 );
not ( w_22504 , w_22505 );
and ( w_22505 , w_22502 , w_22503 );
buf ( w_22502 , \5755_b1 );
not ( w_22502 , w_22506 );
not ( w_22503 , w_22507 );
and ( w_22506 , w_22507 , \5755_b0 );
or ( \8953_b1 , \8948_b1 , \8952_b1 );
xor ( \8953_b0 , \8948_b0 , w_22508 );
not ( w_22508 , w_22509 );
and ( w_22509 , \8952_b1 , \8952_b0 );
or ( \8954_b1 , \5842_b1 , \7140_b1 );
not ( \7140_b1 , w_22510 );
and ( \8954_b0 , \5842_b0 , w_22511 );
and ( w_22510 , w_22511 , \7140_b0 );
or ( \8955_b1 , \5854_b1 , \7138_b1 );
not ( \7138_b1 , w_22512 );
and ( \8955_b0 , \5854_b0 , w_22513 );
and ( w_22512 , w_22513 , \7138_b0 );
or ( \8956_b1 , \8954_b1 , w_22515 );
not ( w_22515 , w_22516 );
and ( \8956_b0 , \8954_b0 , w_22517 );
and ( w_22516 ,  , w_22517 );
buf ( w_22515 , \8955_b1 );
not ( w_22515 , w_22518 );
not (  , w_22519 );
and ( w_22518 , w_22519 , \8955_b0 );
or ( \8957_b1 , \8956_b1 , w_22520 );
xor ( \8957_b0 , \8956_b0 , w_22522 );
not ( w_22522 , w_22523 );
and ( w_22523 , w_22520 , w_22521 );
buf ( w_22520 , \7146_b1 );
not ( w_22520 , w_22524 );
not ( w_22521 , w_22525 );
and ( w_22524 , w_22525 , \7146_b0 );
or ( \8958_b1 , \5861_b1 , \7157_b1 );
not ( \7157_b1 , w_22526 );
and ( \8958_b0 , \5861_b0 , w_22527 );
and ( w_22526 , w_22527 , \7157_b0 );
or ( \8959_b1 , \5873_b1 , \7155_b1 );
not ( \7155_b1 , w_22528 );
and ( \8959_b0 , \5873_b0 , w_22529 );
and ( w_22528 , w_22529 , \7155_b0 );
or ( \8960_b1 , \8958_b1 , w_22531 );
not ( w_22531 , w_22532 );
and ( \8960_b0 , \8958_b0 , w_22533 );
and ( w_22532 ,  , w_22533 );
buf ( w_22531 , \8959_b1 );
not ( w_22531 , w_22534 );
not (  , w_22535 );
and ( w_22534 , w_22535 , \8959_b0 );
or ( \8961_b1 , \8960_b1 , w_22536 );
xor ( \8961_b0 , \8960_b0 , w_22538 );
not ( w_22538 , w_22539 );
and ( w_22539 , w_22536 , w_22537 );
buf ( w_22536 , \7163_b1 );
not ( w_22536 , w_22540 );
not ( w_22537 , w_22541 );
and ( w_22540 , w_22541 , \7163_b0 );
or ( \8962_b1 , \8957_b1 , \8961_b1 );
xor ( \8962_b0 , \8957_b0 , w_22542 );
not ( w_22542 , w_22543 );
and ( w_22543 , \8961_b1 , \8961_b0 );
or ( \8963_b1 , \5881_b1 , \7175_b1 );
not ( \7175_b1 , w_22544 );
and ( \8963_b0 , \5881_b0 , w_22545 );
and ( w_22544 , w_22545 , \7175_b0 );
or ( \8964_b1 , \5893_b1 , \7173_b1 );
not ( \7173_b1 , w_22546 );
and ( \8964_b0 , \5893_b0 , w_22547 );
and ( w_22546 , w_22547 , \7173_b0 );
or ( \8965_b1 , \8963_b1 , w_22549 );
not ( w_22549 , w_22550 );
and ( \8965_b0 , \8963_b0 , w_22551 );
and ( w_22550 ,  , w_22551 );
buf ( w_22549 , \8964_b1 );
not ( w_22549 , w_22552 );
not (  , w_22553 );
and ( w_22552 , w_22553 , \8964_b0 );
or ( \8966_b1 , \8965_b1 , w_22554 );
xor ( \8966_b0 , \8965_b0 , w_22556 );
not ( w_22556 , w_22557 );
and ( w_22557 , w_22554 , w_22555 );
buf ( w_22554 , \7181_b1 );
not ( w_22554 , w_22558 );
not ( w_22555 , w_22559 );
and ( w_22558 , w_22559 , \7181_b0 );
or ( \8967_b1 , \8962_b1 , \8966_b1 );
xor ( \8967_b0 , \8962_b0 , w_22560 );
not ( w_22560 , w_22561 );
and ( w_22561 , \8966_b1 , \8966_b0 );
or ( \8968_b1 , \8953_b1 , \8967_b1 );
xor ( \8968_b0 , \8953_b0 , w_22562 );
not ( w_22562 , w_22563 );
and ( w_22563 , \8967_b1 , \8967_b0 );
or ( \8969_b1 , \5780_b1 , \7082_b1 );
not ( \7082_b1 , w_22564 );
and ( \8969_b0 , \5780_b0 , w_22565 );
and ( w_22564 , w_22565 , \7082_b0 );
or ( \8970_b1 , \5792_b1 , \7080_b1 );
not ( \7080_b1 , w_22566 );
and ( \8970_b0 , \5792_b0 , w_22567 );
and ( w_22566 , w_22567 , \7080_b0 );
or ( \8971_b1 , \8969_b1 , w_22569 );
not ( w_22569 , w_22570 );
and ( \8971_b0 , \8969_b0 , w_22571 );
and ( w_22570 ,  , w_22571 );
buf ( w_22569 , \8970_b1 );
not ( w_22569 , w_22572 );
not (  , w_22573 );
and ( w_22572 , w_22573 , \8970_b0 );
or ( \8972_b1 , \8971_b1 , w_22574 );
xor ( \8972_b0 , \8971_b0 , w_22576 );
not ( w_22576 , w_22577 );
and ( w_22577 , w_22574 , w_22575 );
buf ( w_22574 , \7088_b1 );
not ( w_22574 , w_22578 );
not ( w_22575 , w_22579 );
and ( w_22578 , w_22579 , \7088_b0 );
or ( \8973_b1 , \5799_b1 , \7099_b1 );
not ( \7099_b1 , w_22580 );
and ( \8973_b0 , \5799_b0 , w_22581 );
and ( w_22580 , w_22581 , \7099_b0 );
or ( \8974_b1 , \5811_b1 , \7097_b1 );
not ( \7097_b1 , w_22582 );
and ( \8974_b0 , \5811_b0 , w_22583 );
and ( w_22582 , w_22583 , \7097_b0 );
or ( \8975_b1 , \8973_b1 , w_22585 );
not ( w_22585 , w_22586 );
and ( \8975_b0 , \8973_b0 , w_22587 );
and ( w_22586 ,  , w_22587 );
buf ( w_22585 , \8974_b1 );
not ( w_22585 , w_22588 );
not (  , w_22589 );
and ( w_22588 , w_22589 , \8974_b0 );
or ( \8976_b1 , \8975_b1 , w_22590 );
xor ( \8976_b0 , \8975_b0 , w_22592 );
not ( w_22592 , w_22593 );
and ( w_22593 , w_22590 , w_22591 );
buf ( w_22590 , \7105_b1 );
not ( w_22590 , w_22594 );
not ( w_22591 , w_22595 );
and ( w_22594 , w_22595 , \7105_b0 );
or ( \8977_b1 , \8972_b1 , \8976_b1 );
xor ( \8977_b0 , \8972_b0 , w_22596 );
not ( w_22596 , w_22597 );
and ( w_22597 , \8976_b1 , \8976_b0 );
or ( \8978_b1 , \5819_b1 , \7117_b1 );
not ( \7117_b1 , w_22598 );
and ( \8978_b0 , \5819_b0 , w_22599 );
and ( w_22598 , w_22599 , \7117_b0 );
or ( \8979_b1 , \5831_b1 , \7115_b1 );
not ( \7115_b1 , w_22600 );
and ( \8979_b0 , \5831_b0 , w_22601 );
and ( w_22600 , w_22601 , \7115_b0 );
or ( \8980_b1 , \8978_b1 , w_22603 );
not ( w_22603 , w_22604 );
and ( \8980_b0 , \8978_b0 , w_22605 );
and ( w_22604 ,  , w_22605 );
buf ( w_22603 , \8979_b1 );
not ( w_22603 , w_22606 );
not (  , w_22607 );
and ( w_22606 , w_22607 , \8979_b0 );
or ( \8981_b1 , \8980_b1 , w_22608 );
xor ( \8981_b0 , \8980_b0 , w_22610 );
not ( w_22610 , w_22611 );
and ( w_22611 , w_22608 , w_22609 );
buf ( w_22608 , \7123_b1 );
not ( w_22608 , w_22612 );
not ( w_22609 , w_22613 );
and ( w_22612 , w_22613 , \7123_b0 );
or ( \8982_b1 , \8977_b1 , \8981_b1 );
xor ( \8982_b0 , \8977_b0 , w_22614 );
not ( w_22614 , w_22615 );
and ( w_22615 , \8981_b1 , \8981_b0 );
or ( \8983_b1 , \8968_b1 , \8982_b1 );
xor ( \8983_b0 , \8968_b0 , w_22616 );
not ( w_22616 , w_22617 );
and ( w_22617 , \8982_b1 , \8982_b0 );
or ( \8984_b1 , \8939_b1 , \8983_b1 );
xor ( \8984_b0 , \8939_b0 , w_22618 );
not ( w_22618 , w_22619 );
and ( w_22619 , \8983_b1 , \8983_b0 );
or ( \8985_b1 , \8925_b1 , \8984_b1 );
xor ( \8985_b0 , \8925_b0 , w_22620 );
not ( w_22620 , w_22621 );
and ( w_22621 , \8984_b1 , \8984_b0 );
or ( \8986_b1 , \8729_b1 , \8733_b1 );
not ( \8733_b1 , w_22622 );
and ( \8986_b0 , \8729_b0 , w_22623 );
and ( w_22622 , w_22623 , \8733_b0 );
or ( \8987_b1 , \8733_b1 , \8738_b1 );
not ( \8738_b1 , w_22624 );
and ( \8987_b0 , \8733_b0 , w_22625 );
and ( w_22624 , w_22625 , \8738_b0 );
or ( \8988_b1 , \8729_b1 , \8738_b1 );
not ( \8738_b1 , w_22626 );
and ( \8988_b0 , \8729_b0 , w_22627 );
and ( w_22626 , w_22627 , \8738_b0 );
or ( \8990_b1 , \8715_b1 , \8719_b1 );
not ( \8719_b1 , w_22628 );
and ( \8990_b0 , \8715_b0 , w_22629 );
and ( w_22628 , w_22629 , \8719_b0 );
or ( \8991_b1 , \8719_b1 , \8724_b1 );
not ( \8724_b1 , w_22630 );
and ( \8991_b0 , \8719_b0 , w_22631 );
and ( w_22630 , w_22631 , \8724_b0 );
or ( \8992_b1 , \8715_b1 , \8724_b1 );
not ( \8724_b1 , w_22632 );
and ( \8992_b0 , \8715_b0 , w_22633 );
and ( w_22632 , w_22633 , \8724_b0 );
or ( \8994_b1 , \8989_b1 , \8993_b1 );
xor ( \8994_b0 , \8989_b0 , w_22634 );
not ( w_22634 , w_22635 );
and ( w_22635 , \8993_b1 , \8993_b0 );
or ( \8995_b1 , \8795_b1 , \8809_b1 );
not ( \8809_b1 , w_22636 );
and ( \8995_b0 , \8795_b0 , w_22637 );
and ( w_22636 , w_22637 , \8809_b0 );
or ( \8996_b1 , \8809_b1 , \8824_b1 );
not ( \8824_b1 , w_22638 );
and ( \8996_b0 , \8809_b0 , w_22639 );
and ( w_22638 , w_22639 , \8824_b0 );
or ( \8997_b1 , \8795_b1 , \8824_b1 );
not ( \8824_b1 , w_22640 );
and ( \8997_b0 , \8795_b0 , w_22641 );
and ( w_22640 , w_22641 , \8824_b0 );
or ( \8999_b1 , \8994_b1 , \8998_b1 );
xor ( \8999_b0 , \8994_b0 , w_22642 );
not ( w_22642 , w_22643 );
and ( w_22643 , \8998_b1 , \8998_b0 );
or ( \9000_b1 , \8985_b1 , \8999_b1 );
xor ( \9000_b0 , \8985_b0 , w_22644 );
not ( w_22644 , w_22645 );
and ( w_22645 , \8999_b1 , \8999_b0 );
or ( \9001_b1 , \8871_b1 , \9000_b1 );
xor ( \9001_b0 , \8871_b0 , w_22646 );
not ( w_22646 , w_22647 );
and ( w_22647 , \9000_b1 , \9000_b0 );
or ( \9002_b1 , \8862_b1 , \9001_b1 );
xor ( \9002_b0 , \8862_b0 , w_22648 );
not ( w_22648 , w_22649 );
and ( w_22649 , \9001_b1 , \9001_b0 );
or ( \9003_b1 , \8687_b1 , \8701_b1 );
not ( \8701_b1 , w_22650 );
and ( \9003_b0 , \8687_b0 , w_22651 );
and ( w_22650 , w_22651 , \8701_b0 );
or ( \9004_b1 , \8701_b1 , \8840_b1 );
not ( \8840_b1 , w_22652 );
and ( \9004_b0 , \8701_b0 , w_22653 );
and ( w_22652 , w_22653 , \8840_b0 );
or ( \9005_b1 , \8687_b1 , \8840_b1 );
not ( \8840_b1 , w_22654 );
and ( \9005_b0 , \8687_b0 , w_22655 );
and ( w_22654 , w_22655 , \8840_b0 );
or ( \9007_b1 , \9002_b1 , w_22657 );
not ( w_22657 , w_22658 );
and ( \9007_b0 , \9002_b0 , w_22659 );
and ( w_22658 ,  , w_22659 );
buf ( w_22657 , \9006_b1 );
not ( w_22657 , w_22660 );
not (  , w_22661 );
and ( w_22660 , w_22661 , \9006_b0 );
or ( \9008_b1 , \8846_b1 , w_22663 );
not ( w_22663 , w_22664 );
and ( \9008_b0 , \8846_b0 , w_22665 );
and ( w_22664 ,  , w_22665 );
buf ( w_22663 , \9007_b1 );
not ( w_22663 , w_22666 );
not (  , w_22667 );
and ( w_22666 , w_22667 , \9007_b0 );
or ( \9009_b1 , \8683_b1 , w_22669 );
not ( w_22669 , w_22670 );
and ( \9009_b0 , \8683_b0 , w_22671 );
and ( w_22670 ,  , w_22671 );
buf ( w_22669 , \9008_b1 );
not ( w_22669 , w_22672 );
not (  , w_22673 );
and ( w_22672 , w_22673 , \9008_b0 );
or ( \9010_b1 , \8361_b1 , w_22675 );
not ( w_22675 , w_22676 );
and ( \9010_b0 , \8361_b0 , w_22677 );
and ( w_22676 ,  , w_22677 );
buf ( w_22675 , \9009_b1 );
not ( w_22675 , w_22678 );
not (  , w_22679 );
and ( w_22678 , w_22679 , \9009_b0 );
or ( \9011_b1 , \8866_b1 , \8870_b1 );
not ( \8870_b1 , w_22680 );
and ( \9011_b0 , \8866_b0 , w_22681 );
and ( w_22680 , w_22681 , \8870_b0 );
or ( \9012_b1 , \8870_b1 , \9000_b1 );
not ( \9000_b1 , w_22682 );
and ( \9012_b0 , \8870_b0 , w_22683 );
and ( w_22682 , w_22683 , \9000_b0 );
or ( \9013_b1 , \8866_b1 , \9000_b1 );
not ( \9000_b1 , w_22684 );
and ( \9013_b0 , \8866_b0 , w_22685 );
and ( w_22684 , w_22685 , \9000_b0 );
or ( \9015_b1 , \8989_b1 , \8993_b1 );
not ( \8993_b1 , w_22686 );
and ( \9015_b0 , \8989_b0 , w_22687 );
and ( w_22686 , w_22687 , \8993_b0 );
or ( \9016_b1 , \8993_b1 , \8998_b1 );
not ( \8998_b1 , w_22688 );
and ( \9016_b0 , \8993_b0 , w_22689 );
and ( w_22688 , w_22689 , \8998_b0 );
or ( \9017_b1 , \8989_b1 , \8998_b1 );
not ( \8998_b1 , w_22690 );
and ( \9017_b0 , \8989_b0 , w_22691 );
and ( w_22690 , w_22691 , \8998_b0 );
or ( \9019_b1 , \8929_b1 , \8938_b1 );
not ( \8938_b1 , w_22692 );
and ( \9019_b0 , \8929_b0 , w_22693 );
and ( w_22692 , w_22693 , \8938_b0 );
or ( \9020_b1 , \8938_b1 , \8983_b1 );
not ( \8983_b1 , w_22694 );
and ( \9020_b0 , \8938_b0 , w_22695 );
and ( w_22694 , w_22695 , \8983_b0 );
or ( \9021_b1 , \8929_b1 , \8983_b1 );
not ( \8983_b1 , w_22696 );
and ( \9021_b0 , \8929_b0 , w_22697 );
and ( w_22696 , w_22697 , \8983_b0 );
or ( \9023_b1 , \9018_b1 , \9022_b1 );
xor ( \9023_b0 , \9018_b0 , w_22698 );
not ( w_22698 , w_22699 );
and ( w_22699 , \9022_b1 , \9022_b0 );
or ( \9024_b1 , \8898_b1 , \8909_b1 );
not ( \8909_b1 , w_22700 );
and ( \9024_b0 , \8898_b0 , w_22701 );
and ( w_22700 , w_22701 , \8909_b0 );
or ( \9025_b1 , \8909_b1 , \8924_b1 );
not ( \8924_b1 , w_22702 );
and ( \9025_b0 , \8909_b0 , w_22703 );
and ( w_22702 , w_22703 , \8924_b0 );
or ( \9026_b1 , \8898_b1 , \8924_b1 );
not ( \8924_b1 , w_22704 );
and ( \9026_b0 , \8898_b0 , w_22705 );
and ( w_22704 , w_22705 , \8924_b0 );
or ( \9028_b1 , \9023_b1 , \9027_b1 );
xor ( \9028_b0 , \9023_b0 , w_22706 );
not ( w_22706 , w_22707 );
and ( w_22707 , \9027_b1 , \9027_b0 );
or ( \9029_b1 , \9014_b1 , \9028_b1 );
xor ( \9029_b0 , \9014_b0 , w_22708 );
not ( w_22708 , w_22709 );
and ( w_22709 , \9028_b1 , \9028_b0 );
or ( \9030_b1 , \8854_b1 , \8858_b1 );
not ( \8858_b1 , w_22710 );
and ( \9030_b0 , \8854_b0 , w_22711 );
and ( w_22710 , w_22711 , \8858_b0 );
or ( \9031_b1 , \8858_b1 , \8860_b1 );
not ( \8860_b1 , w_22712 );
and ( \9031_b0 , \8858_b0 , w_22713 );
and ( w_22712 , w_22713 , \8860_b0 );
or ( \9032_b1 , \8854_b1 , \8860_b1 );
not ( \8860_b1 , w_22714 );
and ( \9032_b0 , \8854_b0 , w_22715 );
and ( w_22714 , w_22715 , \8860_b0 );
or ( \9034_b1 , \8925_b1 , \8984_b1 );
not ( \8984_b1 , w_22716 );
and ( \9034_b0 , \8925_b0 , w_22717 );
and ( w_22716 , w_22717 , \8984_b0 );
or ( \9035_b1 , \8984_b1 , \8999_b1 );
not ( \8999_b1 , w_22718 );
and ( \9035_b0 , \8984_b0 , w_22719 );
and ( w_22718 , w_22719 , \8999_b0 );
or ( \9036_b1 , \8925_b1 , \8999_b1 );
not ( \8999_b1 , w_22720 );
and ( \9036_b0 , \8925_b0 , w_22721 );
and ( w_22720 , w_22721 , \8999_b0 );
or ( \9038_b1 , \9033_b1 , \9037_b1 );
xor ( \9038_b0 , \9033_b0 , w_22722 );
not ( w_22722 , w_22723 );
and ( w_22723 , \9037_b1 , \9037_b0 );
or ( \9039_b1 , \8943_b1 , \8947_b1 );
not ( \8947_b1 , w_22724 );
and ( \9039_b0 , \8943_b0 , w_22725 );
and ( w_22724 , w_22725 , \8947_b0 );
or ( \9040_b1 , \8947_b1 , \8952_b1 );
not ( \8952_b1 , w_22726 );
and ( \9040_b0 , \8947_b0 , w_22727 );
and ( w_22726 , w_22727 , \8952_b0 );
or ( \9041_b1 , \8943_b1 , \8952_b1 );
not ( \8952_b1 , w_22728 );
and ( \9041_b0 , \8943_b0 , w_22729 );
and ( w_22728 , w_22729 , \8952_b0 );
or ( \9043_b1 , \8887_b1 , \8891_b1 );
not ( \8891_b1 , w_22730 );
and ( \9043_b0 , \8887_b0 , w_22731 );
and ( w_22730 , w_22731 , \8891_b0 );
or ( \9044_b1 , \8891_b1 , \8896_b1 );
not ( \8896_b1 , w_22732 );
and ( \9044_b0 , \8891_b0 , w_22733 );
and ( w_22732 , w_22733 , \8896_b0 );
or ( \9045_b1 , \8887_b1 , \8896_b1 );
not ( \8896_b1 , w_22734 );
and ( \9045_b0 , \8887_b0 , w_22735 );
and ( w_22734 , w_22735 , \8896_b0 );
or ( \9047_b1 , \9042_b1 , \9046_b1 );
xor ( \9047_b0 , \9042_b0 , w_22736 );
not ( w_22736 , w_22737 );
and ( w_22737 , \9046_b1 , \9046_b0 );
or ( \9048_b1 , \8875_b1 , \8879_b1 );
not ( \8879_b1 , w_22738 );
and ( \9048_b0 , \8875_b0 , w_22739 );
and ( w_22738 , w_22739 , \8879_b0 );
or ( \9049_b1 , \8879_b1 , \8882_b1 );
not ( \8882_b1 , w_22740 );
and ( \9049_b0 , \8879_b0 , w_22741 );
and ( w_22740 , w_22741 , \8882_b0 );
or ( \9050_b1 , \8875_b1 , \8882_b1 );
not ( \8882_b1 , w_22742 );
and ( \9050_b0 , \8875_b0 , w_22743 );
and ( w_22742 , w_22743 , \8882_b0 );
or ( \9052_b1 , \9047_b1 , \9051_b1 );
xor ( \9052_b0 , \9047_b0 , w_22744 );
not ( w_22744 , w_22745 );
and ( w_22745 , \9051_b1 , \9051_b0 );
or ( \9053_b1 , \5878_b1 , \8932_b1 );
not ( \8932_b1 , w_22746 );
and ( \9053_b0 , \5878_b0 , w_22747 );
and ( w_22746 , w_22747 , \8932_b0 );
or ( \9054_b1 , \8932_b1 , \8937_b1 );
not ( \8937_b1 , w_22748 );
and ( \9054_b0 , \8932_b0 , w_22749 );
and ( w_22748 , w_22749 , \8937_b0 );
or ( \9055_b1 , \5878_b1 , \8937_b1 );
not ( \8937_b1 , w_22750 );
and ( \9055_b0 , \5878_b0 , w_22751 );
and ( w_22750 , w_22751 , \8937_b0 );
or ( \9057_b1 , \8972_b1 , \8976_b1 );
not ( \8976_b1 , w_22752 );
and ( \9057_b0 , \8972_b0 , w_22753 );
and ( w_22752 , w_22753 , \8976_b0 );
or ( \9058_b1 , \8976_b1 , \8981_b1 );
not ( \8981_b1 , w_22754 );
and ( \9058_b0 , \8976_b0 , w_22755 );
and ( w_22754 , w_22755 , \8981_b0 );
or ( \9059_b1 , \8972_b1 , \8981_b1 );
not ( \8981_b1 , w_22756 );
and ( \9059_b0 , \8972_b0 , w_22757 );
and ( w_22756 , w_22757 , \8981_b0 );
or ( \9061_b1 , \9056_b1 , \9060_b1 );
xor ( \9061_b0 , \9056_b0 , w_22758 );
not ( w_22758 , w_22759 );
and ( w_22759 , \9060_b1 , \9060_b0 );
or ( \9062_b1 , \8957_b1 , \8961_b1 );
not ( \8961_b1 , w_22760 );
and ( \9062_b0 , \8957_b0 , w_22761 );
and ( w_22760 , w_22761 , \8961_b0 );
or ( \9063_b1 , \8961_b1 , \8966_b1 );
not ( \8966_b1 , w_22762 );
and ( \9063_b0 , \8961_b0 , w_22763 );
and ( w_22762 , w_22763 , \8966_b0 );
or ( \9064_b1 , \8957_b1 , \8966_b1 );
not ( \8966_b1 , w_22764 );
and ( \9064_b0 , \8957_b0 , w_22765 );
and ( w_22764 , w_22765 , \8966_b0 );
or ( \9066_b1 , \9061_b1 , \9065_b1 );
xor ( \9066_b0 , \9061_b0 , w_22766 );
not ( w_22766 , w_22767 );
and ( w_22767 , \9065_b1 , \9065_b0 );
or ( \9067_b1 , \9052_b1 , \9066_b1 );
xor ( \9067_b0 , \9052_b0 , w_22768 );
not ( w_22768 , w_22769 );
and ( w_22769 , \9066_b1 , \9066_b0 );
or ( \9068_b1 , \8953_b1 , \8967_b1 );
not ( \8967_b1 , w_22770 );
and ( \9068_b0 , \8953_b0 , w_22771 );
and ( w_22770 , w_22771 , \8967_b0 );
or ( \9069_b1 , \8967_b1 , \8982_b1 );
not ( \8982_b1 , w_22772 );
and ( \9069_b0 , \8967_b0 , w_22773 );
and ( w_22772 , w_22773 , \8982_b0 );
or ( \9070_b1 , \8953_b1 , \8982_b1 );
not ( \8982_b1 , w_22774 );
and ( \9070_b0 , \8953_b0 , w_22775 );
and ( w_22774 , w_22775 , \8982_b0 );
or ( \9072_b1 , \5873_b1 , \7157_b1 );
not ( \7157_b1 , w_22776 );
and ( \9072_b0 , \5873_b0 , w_22777 );
and ( w_22776 , w_22777 , \7157_b0 );
or ( \9073_b1 , \5842_b1 , \7155_b1 );
not ( \7155_b1 , w_22778 );
and ( \9073_b0 , \5842_b0 , w_22779 );
and ( w_22778 , w_22779 , \7155_b0 );
or ( \9074_b1 , \9072_b1 , w_22781 );
not ( w_22781 , w_22782 );
and ( \9074_b0 , \9072_b0 , w_22783 );
and ( w_22782 ,  , w_22783 );
buf ( w_22781 , \9073_b1 );
not ( w_22781 , w_22784 );
not (  , w_22785 );
and ( w_22784 , w_22785 , \9073_b0 );
or ( \9075_b1 , \9074_b1 , w_22786 );
xor ( \9075_b0 , \9074_b0 , w_22788 );
not ( w_22788 , w_22789 );
and ( w_22789 , w_22786 , w_22787 );
buf ( w_22786 , \7163_b1 );
not ( w_22786 , w_22790 );
not ( w_22787 , w_22791 );
and ( w_22790 , w_22791 , \7163_b0 );
or ( \9076_b1 , \5893_b1 , \7175_b1 );
not ( \7175_b1 , w_22792 );
and ( \9076_b0 , \5893_b0 , w_22793 );
and ( w_22792 , w_22793 , \7175_b0 );
or ( \9077_b1 , \5861_b1 , \7173_b1 );
not ( \7173_b1 , w_22794 );
and ( \9077_b0 , \5861_b0 , w_22795 );
and ( w_22794 , w_22795 , \7173_b0 );
or ( \9078_b1 , \9076_b1 , w_22797 );
not ( w_22797 , w_22798 );
and ( \9078_b0 , \9076_b0 , w_22799 );
and ( w_22798 ,  , w_22799 );
buf ( w_22797 , \9077_b1 );
not ( w_22797 , w_22800 );
not (  , w_22801 );
and ( w_22800 , w_22801 , \9077_b0 );
or ( \9079_b1 , \9078_b1 , w_22802 );
xor ( \9079_b0 , \9078_b0 , w_22804 );
not ( w_22804 , w_22805 );
and ( w_22805 , w_22802 , w_22803 );
buf ( w_22802 , \7181_b1 );
not ( w_22802 , w_22806 );
not ( w_22803 , w_22807 );
and ( w_22806 , w_22807 , \7181_b0 );
or ( \9080_b1 , \9075_b1 , \9079_b1 );
xor ( \9080_b0 , \9075_b0 , w_22808 );
not ( w_22808 , w_22809 );
and ( w_22809 , \9079_b1 , \9079_b0 );
or ( \9081_b1 , \5918_b1 , \7192_b1 );
not ( \7192_b1 , w_22810 );
and ( \9081_b0 , \5918_b0 , w_22811 );
and ( w_22810 , w_22811 , \7192_b0 );
or ( \9082_b1 , \5881_b1 , \7190_b1 );
not ( \7190_b1 , w_22812 );
and ( \9082_b0 , \5881_b0 , w_22813 );
and ( w_22812 , w_22813 , \7190_b0 );
or ( \9083_b1 , \9081_b1 , w_22815 );
not ( w_22815 , w_22816 );
and ( \9083_b0 , \9081_b0 , w_22817 );
and ( w_22816 ,  , w_22817 );
buf ( w_22815 , \9082_b1 );
not ( w_22815 , w_22818 );
not (  , w_22819 );
and ( w_22818 , w_22819 , \9082_b0 );
or ( \9084_b1 , \9083_b1 , w_22820 );
xor ( \9084_b0 , \9083_b0 , w_22822 );
not ( w_22822 , w_22823 );
and ( w_22823 , w_22820 , w_22821 );
buf ( w_22820 , \7198_b1 );
not ( w_22820 , w_22824 );
not ( w_22821 , w_22825 );
and ( w_22824 , w_22825 , \7198_b0 );
or ( \9085_b1 , \9080_b1 , \9084_b1 );
xor ( \9085_b0 , \9080_b0 , w_22826 );
not ( w_22826 , w_22827 );
and ( w_22827 , \9084_b1 , \9084_b0 );
or ( \9086_b1 , \5811_b1 , \7099_b1 );
not ( \7099_b1 , w_22828 );
and ( \9086_b0 , \5811_b0 , w_22829 );
and ( w_22828 , w_22829 , \7099_b0 );
or ( \9087_b1 , \5780_b1 , \7097_b1 );
not ( \7097_b1 , w_22830 );
and ( \9087_b0 , \5780_b0 , w_22831 );
and ( w_22830 , w_22831 , \7097_b0 );
or ( \9088_b1 , \9086_b1 , w_22833 );
not ( w_22833 , w_22834 );
and ( \9088_b0 , \9086_b0 , w_22835 );
and ( w_22834 ,  , w_22835 );
buf ( w_22833 , \9087_b1 );
not ( w_22833 , w_22836 );
not (  , w_22837 );
and ( w_22836 , w_22837 , \9087_b0 );
or ( \9089_b1 , \9088_b1 , w_22838 );
xor ( \9089_b0 , \9088_b0 , w_22840 );
not ( w_22840 , w_22841 );
and ( w_22841 , w_22838 , w_22839 );
buf ( w_22838 , \7105_b1 );
not ( w_22838 , w_22842 );
not ( w_22839 , w_22843 );
and ( w_22842 , w_22843 , \7105_b0 );
or ( \9090_b1 , \5831_b1 , \7117_b1 );
not ( \7117_b1 , w_22844 );
and ( \9090_b0 , \5831_b0 , w_22845 );
and ( w_22844 , w_22845 , \7117_b0 );
or ( \9091_b1 , \5799_b1 , \7115_b1 );
not ( \7115_b1 , w_22846 );
and ( \9091_b0 , \5799_b0 , w_22847 );
and ( w_22846 , w_22847 , \7115_b0 );
or ( \9092_b1 , \9090_b1 , w_22849 );
not ( w_22849 , w_22850 );
and ( \9092_b0 , \9090_b0 , w_22851 );
and ( w_22850 ,  , w_22851 );
buf ( w_22849 , \9091_b1 );
not ( w_22849 , w_22852 );
not (  , w_22853 );
and ( w_22852 , w_22853 , \9091_b0 );
or ( \9093_b1 , \9092_b1 , w_22854 );
xor ( \9093_b0 , \9092_b0 , w_22856 );
not ( w_22856 , w_22857 );
and ( w_22857 , w_22854 , w_22855 );
buf ( w_22854 , \7123_b1 );
not ( w_22854 , w_22858 );
not ( w_22855 , w_22859 );
and ( w_22858 , w_22859 , \7123_b0 );
or ( \9094_b1 , \9089_b1 , \9093_b1 );
xor ( \9094_b0 , \9089_b0 , w_22860 );
not ( w_22860 , w_22861 );
and ( w_22861 , \9093_b1 , \9093_b0 );
or ( \9095_b1 , \5854_b1 , \7140_b1 );
not ( \7140_b1 , w_22862 );
and ( \9095_b0 , \5854_b0 , w_22863 );
and ( w_22862 , w_22863 , \7140_b0 );
or ( \9096_b1 , \5819_b1 , \7138_b1 );
not ( \7138_b1 , w_22864 );
and ( \9096_b0 , \5819_b0 , w_22865 );
and ( w_22864 , w_22865 , \7138_b0 );
or ( \9097_b1 , \9095_b1 , w_22867 );
not ( w_22867 , w_22868 );
and ( \9097_b0 , \9095_b0 , w_22869 );
and ( w_22868 ,  , w_22869 );
buf ( w_22867 , \9096_b1 );
not ( w_22867 , w_22870 );
not (  , w_22871 );
and ( w_22870 , w_22871 , \9096_b0 );
or ( \9098_b1 , \9097_b1 , w_22872 );
xor ( \9098_b0 , \9097_b0 , w_22874 );
not ( w_22874 , w_22875 );
and ( w_22875 , w_22872 , w_22873 );
buf ( w_22872 , \7146_b1 );
not ( w_22872 , w_22876 );
not ( w_22873 , w_22877 );
and ( w_22876 , w_22877 , \7146_b0 );
or ( \9099_b1 , \9094_b1 , \9098_b1 );
xor ( \9099_b0 , \9094_b0 , w_22878 );
not ( w_22878 , w_22879 );
and ( w_22879 , \9098_b1 , \9098_b0 );
or ( \9100_b1 , \9085_b1 , \9099_b1 );
xor ( \9100_b0 , \9085_b0 , w_22880 );
not ( w_22880 , w_22881 );
and ( w_22881 , \9099_b1 , \9099_b0 );
buf ( \9101_b1 , \7049_b1 );
not ( \9101_b1 , w_22882 );
not ( \9101_b0 , w_22883 );
and ( w_22882 , w_22883 , \7049_b0 );
or ( \9102_b1 , \5770_b1 , \7061_b1 );
not ( \7061_b1 , w_22884 );
and ( \9102_b0 , \5770_b0 , w_22885 );
and ( w_22884 , w_22885 , \7061_b0 );
or ( \9103_b1 , \5737_b1 , \7059_b1 );
not ( \7059_b1 , w_22886 );
and ( \9103_b0 , \5737_b0 , w_22887 );
and ( w_22886 , w_22887 , \7059_b0 );
or ( \9104_b1 , \9102_b1 , w_22889 );
not ( w_22889 , w_22890 );
and ( \9104_b0 , \9102_b0 , w_22891 );
and ( w_22890 ,  , w_22891 );
buf ( w_22889 , \9103_b1 );
not ( w_22889 , w_22892 );
not (  , w_22893 );
and ( w_22892 , w_22893 , \9103_b0 );
or ( \9105_b1 , \9104_b1 , w_22894 );
xor ( \9105_b0 , \9104_b0 , w_22896 );
not ( w_22896 , w_22897 );
and ( w_22897 , w_22894 , w_22895 );
buf ( w_22894 , \7067_b1 );
not ( w_22894 , w_22898 );
not ( w_22895 , w_22899 );
and ( w_22898 , w_22899 , \7067_b0 );
or ( \9106_b1 , \9101_b1 , \9105_b1 );
xor ( \9106_b0 , \9101_b0 , w_22900 );
not ( w_22900 , w_22901 );
and ( w_22901 , \9105_b1 , \9105_b0 );
or ( \9107_b1 , \5792_b1 , \7082_b1 );
not ( \7082_b1 , w_22902 );
and ( \9107_b0 , \5792_b0 , w_22903 );
and ( w_22902 , w_22903 , \7082_b0 );
or ( \9108_b1 , \5758_b1 , \7080_b1 );
not ( \7080_b1 , w_22904 );
and ( \9108_b0 , \5758_b0 , w_22905 );
and ( w_22904 , w_22905 , \7080_b0 );
or ( \9109_b1 , \9107_b1 , w_22907 );
not ( w_22907 , w_22908 );
and ( \9109_b0 , \9107_b0 , w_22909 );
and ( w_22908 ,  , w_22909 );
buf ( w_22907 , \9108_b1 );
not ( w_22907 , w_22910 );
not (  , w_22911 );
and ( w_22910 , w_22911 , \9108_b0 );
or ( \9110_b1 , \9109_b1 , w_22912 );
xor ( \9110_b0 , \9109_b0 , w_22914 );
not ( w_22914 , w_22915 );
and ( w_22915 , w_22912 , w_22913 );
buf ( w_22912 , \7088_b1 );
not ( w_22912 , w_22916 );
not ( w_22913 , w_22917 );
and ( w_22916 , w_22917 , \7088_b0 );
or ( \9111_b1 , \9106_b1 , \9110_b1 );
xor ( \9111_b0 , \9106_b0 , w_22918 );
not ( w_22918 , w_22919 );
and ( w_22919 , \9110_b1 , \9110_b0 );
or ( \9112_b1 , \9100_b1 , \9111_b1 );
xor ( \9112_b0 , \9100_b0 , w_22920 );
not ( w_22920 , w_22921 );
and ( w_22921 , \9111_b1 , \9111_b0 );
or ( \9113_b1 , \9071_b1 , \9112_b1 );
xor ( \9113_b0 , \9071_b0 , w_22922 );
not ( w_22922 , w_22923 );
and ( w_22923 , \9112_b1 , \9112_b0 );
or ( \9114_b1 , \6057_b1 , \5852_b1 );
not ( \5852_b1 , w_22924 );
and ( \9114_b0 , \6057_b0 , w_22925 );
and ( w_22924 , w_22925 , \5852_b0 );
or ( \9115_b1 , \6029_b1 , \5850_b1 );
not ( \5850_b1 , w_22926 );
and ( \9115_b0 , \6029_b0 , w_22927 );
and ( w_22926 , w_22927 , \5850_b0 );
or ( \9116_b1 , \9114_b1 , w_22929 );
not ( w_22929 , w_22930 );
and ( \9116_b0 , \9114_b0 , w_22931 );
and ( w_22930 ,  , w_22931 );
buf ( w_22929 , \9115_b1 );
not ( w_22929 , w_22932 );
not (  , w_22933 );
and ( w_22932 , w_22933 , \9115_b0 );
or ( \9117_b1 , \9116_b1 , w_22934 );
xor ( \9117_b0 , \9116_b0 , w_22936 );
not ( w_22936 , w_22937 );
and ( w_22937 , w_22934 , w_22935 );
buf ( w_22934 , \5859_b1 );
not ( w_22934 , w_22938 );
not ( w_22935 , w_22939 );
and ( w_22938 , w_22939 , \5859_b0 );
or ( \9118_b1 , \6065_b1 , \5871_b1 );
not ( \5871_b1 , w_22940 );
and ( \9118_b0 , \6065_b0 , w_22941 );
and ( w_22940 , w_22941 , \5871_b0 );
or ( \9119_b1 , \6048_b1 , \5869_b1 );
not ( \5869_b1 , w_22942 );
and ( \9119_b0 , \6048_b0 , w_22943 );
and ( w_22942 , w_22943 , \5869_b0 );
or ( \9120_b1 , \9118_b1 , w_22945 );
not ( w_22945 , w_22946 );
and ( \9120_b0 , \9118_b0 , w_22947 );
and ( w_22946 ,  , w_22947 );
buf ( w_22945 , \9119_b1 );
not ( w_22945 , w_22948 );
not (  , w_22949 );
and ( w_22948 , w_22949 , \9119_b0 );
or ( \9121_b1 , \9120_b1 , w_22950 );
xor ( \9121_b0 , \9120_b0 , w_22952 );
not ( w_22952 , w_22953 );
and ( w_22953 , w_22950 , w_22951 );
buf ( w_22950 , \5878_b1 );
not ( w_22950 , w_22954 );
not ( w_22951 , w_22955 );
and ( w_22954 , w_22955 , \5878_b0 );
or ( \9122_b1 , \9117_b1 , \9121_b1 );
xor ( \9122_b0 , \9117_b0 , w_22956 );
not ( w_22956 , w_22957 );
and ( w_22957 , \9121_b1 , \9121_b0 );
or ( \9123_b1 , \5998_b1 , \5790_b1 );
not ( \5790_b1 , w_22958 );
and ( \9123_b0 , \5998_b0 , w_22959 );
and ( w_22958 , w_22959 , \5790_b0 );
or ( \9124_b1 , \5967_b1 , \5788_b1 );
not ( \5788_b1 , w_22960 );
and ( \9124_b0 , \5967_b0 , w_22961 );
and ( w_22960 , w_22961 , \5788_b0 );
or ( \9125_b1 , \9123_b1 , w_22963 );
not ( w_22963 , w_22964 );
and ( \9125_b0 , \9123_b0 , w_22965 );
and ( w_22964 ,  , w_22965 );
buf ( w_22963 , \9124_b1 );
not ( w_22963 , w_22966 );
not (  , w_22967 );
and ( w_22966 , w_22967 , \9124_b0 );
or ( \9126_b1 , \9125_b1 , w_22968 );
xor ( \9126_b0 , \9125_b0 , w_22970 );
not ( w_22970 , w_22971 );
and ( w_22971 , w_22968 , w_22969 );
buf ( w_22968 , \5797_b1 );
not ( w_22968 , w_22972 );
not ( w_22969 , w_22973 );
and ( w_22972 , w_22973 , \5797_b0 );
or ( \9127_b1 , \6018_b1 , \5809_b1 );
not ( \5809_b1 , w_22974 );
and ( \9127_b0 , \6018_b0 , w_22975 );
and ( w_22974 , w_22975 , \5809_b0 );
or ( \9128_b1 , \5986_b1 , \5807_b1 );
not ( \5807_b1 , w_22976 );
and ( \9128_b0 , \5986_b0 , w_22977 );
and ( w_22976 , w_22977 , \5807_b0 );
or ( \9129_b1 , \9127_b1 , w_22979 );
not ( w_22979 , w_22980 );
and ( \9129_b0 , \9127_b0 , w_22981 );
and ( w_22980 ,  , w_22981 );
buf ( w_22979 , \9128_b1 );
not ( w_22979 , w_22982 );
not (  , w_22983 );
and ( w_22982 , w_22983 , \9128_b0 );
or ( \9130_b1 , \9129_b1 , w_22984 );
xor ( \9130_b0 , \9129_b0 , w_22986 );
not ( w_22986 , w_22987 );
and ( w_22987 , w_22984 , w_22985 );
buf ( w_22984 , \5816_b1 );
not ( w_22984 , w_22988 );
not ( w_22985 , w_22989 );
and ( w_22988 , w_22989 , \5816_b0 );
or ( \9131_b1 , \9126_b1 , \9130_b1 );
xor ( \9131_b0 , \9126_b0 , w_22990 );
not ( w_22990 , w_22991 );
and ( w_22991 , \9130_b1 , \9130_b0 );
or ( \9132_b1 , \6041_b1 , \5829_b1 );
not ( \5829_b1 , w_22992 );
and ( \9132_b0 , \6041_b0 , w_22993 );
and ( w_22992 , w_22993 , \5829_b0 );
or ( \9133_b1 , \6006_b1 , \5827_b1 );
not ( \5827_b1 , w_22994 );
and ( \9133_b0 , \6006_b0 , w_22995 );
and ( w_22994 , w_22995 , \5827_b0 );
or ( \9134_b1 , \9132_b1 , w_22997 );
not ( w_22997 , w_22998 );
and ( \9134_b0 , \9132_b0 , w_22999 );
and ( w_22998 ,  , w_22999 );
buf ( w_22997 , \9133_b1 );
not ( w_22997 , w_23000 );
not (  , w_23001 );
and ( w_23000 , w_23001 , \9133_b0 );
or ( \9135_b1 , \9134_b1 , w_23002 );
xor ( \9135_b0 , \9134_b0 , w_23004 );
not ( w_23004 , w_23005 );
and ( w_23005 , w_23002 , w_23003 );
buf ( w_23002 , \5836_b1 );
not ( w_23002 , w_23006 );
not ( w_23003 , w_23007 );
and ( w_23006 , w_23007 , \5836_b0 );
or ( \9136_b1 , \9131_b1 , \9135_b1 );
xor ( \9136_b0 , \9131_b0 , w_23008 );
not ( w_23008 , w_23009 );
and ( w_23009 , \9135_b1 , \9135_b0 );
or ( \9137_b1 , \9122_b1 , \9136_b1 );
xor ( \9137_b0 , \9122_b0 , w_23010 );
not ( w_23010 , w_23011 );
and ( w_23011 , \9136_b1 , \9136_b0 );
or ( \9138_b1 , \5937_b1 , \7203_b1 );
not ( \7203_b1 , w_23012 );
and ( \9138_b0 , \5937_b0 , w_23013 );
and ( w_23012 , w_23013 , \7203_b0 );
or ( \9139_b1 , \5906_b1 , \7201_b1 );
not ( \7201_b1 , w_23014 );
and ( \9139_b0 , \5906_b0 , w_23015 );
and ( w_23014 , w_23015 , \7201_b0 );
or ( \9140_b1 , \9138_b1 , w_23017 );
not ( w_23017 , w_23018 );
and ( \9140_b0 , \9138_b0 , w_23019 );
and ( w_23018 ,  , w_23019 );
buf ( w_23017 , \9139_b1 );
not ( w_23017 , w_23020 );
not (  , w_23021 );
and ( w_23020 , w_23021 , \9139_b0 );
or ( \9141_b1 , \9140_b1 , w_23022 );
xor ( \9141_b0 , \9140_b0 , w_23024 );
not ( w_23024 , w_23025 );
and ( w_23025 , w_23022 , w_23023 );
buf ( w_23022 , \6824_b1 );
not ( w_23022 , w_23026 );
not ( w_23023 , w_23027 );
and ( w_23026 , w_23027 , \6824_b0 );
or ( \9142_b1 , \5957_b1 , \5750_b1 );
not ( \5750_b1 , w_23028 );
and ( \9142_b0 , \5957_b0 , w_23029 );
and ( w_23028 , w_23029 , \5750_b0 );
or ( \9143_b1 , \5925_b1 , \5748_b1 );
not ( \5748_b1 , w_23030 );
and ( \9143_b0 , \5925_b0 , w_23031 );
and ( w_23030 , w_23031 , \5748_b0 );
or ( \9144_b1 , \9142_b1 , w_23033 );
not ( w_23033 , w_23034 );
and ( \9144_b0 , \9142_b0 , w_23035 );
and ( w_23034 ,  , w_23035 );
buf ( w_23033 , \9143_b1 );
not ( w_23033 , w_23036 );
not (  , w_23037 );
and ( w_23036 , w_23037 , \9143_b0 );
or ( \9145_b1 , \9144_b1 , w_23038 );
xor ( \9145_b0 , \9144_b0 , w_23040 );
not ( w_23040 , w_23041 );
and ( w_23041 , w_23038 , w_23039 );
buf ( w_23038 , \5755_b1 );
not ( w_23038 , w_23042 );
not ( w_23039 , w_23043 );
and ( w_23042 , w_23043 , \5755_b0 );
or ( \9146_b1 , \9141_b1 , \9145_b1 );
xor ( \9146_b0 , \9141_b0 , w_23044 );
not ( w_23044 , w_23045 );
and ( w_23045 , \9145_b1 , \9145_b0 );
or ( \9147_b1 , \5979_b1 , \5768_b1 );
not ( \5768_b1 , w_23046 );
and ( \9147_b0 , \5979_b0 , w_23047 );
and ( w_23046 , w_23047 , \5768_b0 );
or ( \9148_b1 , \5945_b1 , \5766_b1 );
not ( \5766_b1 , w_23048 );
and ( \9148_b0 , \5945_b0 , w_23049 );
and ( w_23048 , w_23049 , \5766_b0 );
or ( \9149_b1 , \9147_b1 , w_23051 );
not ( w_23051 , w_23052 );
and ( \9149_b0 , \9147_b0 , w_23053 );
and ( w_23052 ,  , w_23053 );
buf ( w_23051 , \9148_b1 );
not ( w_23051 , w_23054 );
not (  , w_23055 );
and ( w_23054 , w_23055 , \9148_b0 );
or ( \9150_b1 , \9149_b1 , w_23056 );
xor ( \9150_b0 , \9149_b0 , w_23058 );
not ( w_23058 , w_23059 );
and ( w_23059 , w_23056 , w_23057 );
buf ( w_23056 , \5775_b1 );
not ( w_23056 , w_23060 );
not ( w_23057 , w_23061 );
and ( w_23060 , w_23061 , \5775_b0 );
or ( \9151_b1 , \9146_b1 , \9150_b1 );
xor ( \9151_b0 , \9146_b0 , w_23062 );
not ( w_23062 , w_23063 );
and ( w_23063 , \9150_b1 , \9150_b0 );
or ( \9152_b1 , \9137_b1 , \9151_b1 );
xor ( \9152_b0 , \9137_b0 , w_23064 );
not ( w_23064 , w_23065 );
and ( w_23065 , \9151_b1 , \9151_b0 );
or ( \9153_b1 , \9113_b1 , \9152_b1 );
xor ( \9153_b0 , \9113_b0 , w_23066 );
not ( w_23066 , w_23067 );
and ( w_23067 , \9152_b1 , \9152_b0 );
or ( \9154_b1 , \9067_b1 , \9153_b1 );
xor ( \9154_b0 , \9067_b0 , w_23068 );
not ( w_23068 , w_23069 );
and ( w_23069 , \9153_b1 , \9153_b0 );
or ( \9155_b1 , \8914_b1 , \8918_b1 );
not ( \8918_b1 , w_23070 );
and ( \9155_b0 , \8914_b0 , w_23071 );
and ( w_23070 , w_23071 , \8918_b0 );
or ( \9156_b1 , \8918_b1 , \8923_b1 );
not ( \8923_b1 , w_23072 );
and ( \9156_b0 , \8918_b0 , w_23073 );
and ( w_23072 , w_23073 , \8923_b0 );
or ( \9157_b1 , \8914_b1 , \8923_b1 );
not ( \8923_b1 , w_23074 );
and ( \9157_b0 , \8914_b0 , w_23075 );
and ( w_23074 , w_23075 , \8923_b0 );
or ( \9159_b1 , \8902_b1 , \8906_b1 );
not ( \8906_b1 , w_23076 );
and ( \9159_b0 , \8902_b0 , w_23077 );
and ( w_23076 , w_23077 , \8906_b0 );
or ( \9160_b1 , \8906_b1 , \8908_b1 );
not ( \8908_b1 , w_23078 );
and ( \9160_b0 , \8906_b0 , w_23079 );
and ( w_23078 , w_23079 , \8908_b0 );
or ( \9161_b1 , \8902_b1 , \8908_b1 );
not ( \8908_b1 , w_23080 );
and ( \9161_b0 , \8902_b0 , w_23081 );
and ( w_23080 , w_23081 , \8908_b0 );
or ( \9163_b1 , \9158_b1 , \9162_b1 );
xor ( \9163_b0 , \9158_b0 , w_23082 );
not ( w_23082 , w_23083 );
and ( w_23083 , \9162_b1 , \9162_b0 );
or ( \9164_b1 , \8883_b1 , w_23084 );
or ( \9164_b0 , \8883_b0 , \8897_b0 );
not ( \8897_b0 , w_23085 );
and ( w_23085 , w_23084 , \8897_b1 );
or ( \9165_b1 , \9163_b1 , \9164_b1 );
xor ( \9165_b0 , \9163_b0 , w_23086 );
not ( w_23086 , w_23087 );
and ( w_23087 , \9164_b1 , \9164_b0 );
or ( \9166_b1 , \9154_b1 , \9165_b1 );
xor ( \9166_b0 , \9154_b0 , w_23088 );
not ( w_23088 , w_23089 );
and ( w_23089 , \9165_b1 , \9165_b0 );
or ( \9167_b1 , \9038_b1 , \9166_b1 );
xor ( \9167_b0 , \9038_b0 , w_23090 );
not ( w_23090 , w_23091 );
and ( w_23091 , \9166_b1 , \9166_b0 );
or ( \9168_b1 , \9029_b1 , \9167_b1 );
xor ( \9168_b0 , \9029_b0 , w_23092 );
not ( w_23092 , w_23093 );
and ( w_23093 , \9167_b1 , \9167_b0 );
or ( \9169_b1 , \8850_b1 , \8861_b1 );
not ( \8861_b1 , w_23094 );
and ( \9169_b0 , \8850_b0 , w_23095 );
and ( w_23094 , w_23095 , \8861_b0 );
or ( \9170_b1 , \8861_b1 , \9001_b1 );
not ( \9001_b1 , w_23096 );
and ( \9170_b0 , \8861_b0 , w_23097 );
and ( w_23096 , w_23097 , \9001_b0 );
or ( \9171_b1 , \8850_b1 , \9001_b1 );
not ( \9001_b1 , w_23098 );
and ( \9171_b0 , \8850_b0 , w_23099 );
and ( w_23098 , w_23099 , \9001_b0 );
or ( \9173_b1 , \9168_b1 , w_23101 );
not ( w_23101 , w_23102 );
and ( \9173_b0 , \9168_b0 , w_23103 );
and ( w_23102 ,  , w_23103 );
buf ( w_23101 , \9172_b1 );
not ( w_23101 , w_23104 );
not (  , w_23105 );
and ( w_23104 , w_23105 , \9172_b0 );
or ( \9174_b1 , \9033_b1 , \9037_b1 );
not ( \9037_b1 , w_23106 );
and ( \9174_b0 , \9033_b0 , w_23107 );
and ( w_23106 , w_23107 , \9037_b0 );
or ( \9175_b1 , \9037_b1 , \9166_b1 );
not ( \9166_b1 , w_23108 );
and ( \9175_b0 , \9037_b0 , w_23109 );
and ( w_23108 , w_23109 , \9166_b0 );
or ( \9176_b1 , \9033_b1 , \9166_b1 );
not ( \9166_b1 , w_23110 );
and ( \9176_b0 , \9033_b0 , w_23111 );
and ( w_23110 , w_23111 , \9166_b0 );
or ( \9178_b1 , \9158_b1 , \9162_b1 );
not ( \9162_b1 , w_23112 );
and ( \9178_b0 , \9158_b0 , w_23113 );
and ( w_23112 , w_23113 , \9162_b0 );
or ( \9179_b1 , \9162_b1 , \9164_b1 );
not ( \9164_b1 , w_23114 );
and ( \9179_b0 , \9162_b0 , w_23115 );
and ( w_23114 , w_23115 , \9164_b0 );
or ( \9180_b1 , \9158_b1 , \9164_b1 );
not ( \9164_b1 , w_23116 );
and ( \9180_b0 , \9158_b0 , w_23117 );
and ( w_23116 , w_23117 , \9164_b0 );
or ( \9182_b1 , \9071_b1 , \9112_b1 );
not ( \9112_b1 , w_23118 );
and ( \9182_b0 , \9071_b0 , w_23119 );
and ( w_23118 , w_23119 , \9112_b0 );
or ( \9183_b1 , \9112_b1 , \9152_b1 );
not ( \9152_b1 , w_23120 );
and ( \9183_b0 , \9112_b0 , w_23121 );
and ( w_23120 , w_23121 , \9152_b0 );
or ( \9184_b1 , \9071_b1 , \9152_b1 );
not ( \9152_b1 , w_23122 );
and ( \9184_b0 , \9071_b0 , w_23123 );
and ( w_23122 , w_23123 , \9152_b0 );
or ( \9186_b1 , \9181_b1 , \9185_b1 );
xor ( \9186_b0 , \9181_b0 , w_23124 );
not ( w_23124 , w_23125 );
and ( w_23125 , \9185_b1 , \9185_b0 );
or ( \9187_b1 , \9052_b1 , \9066_b1 );
not ( \9066_b1 , w_23126 );
and ( \9187_b0 , \9052_b0 , w_23127 );
and ( w_23126 , w_23127 , \9066_b0 );
or ( \9188_b1 , \9186_b1 , \9187_b1 );
xor ( \9188_b0 , \9186_b0 , w_23128 );
not ( w_23128 , w_23129 );
and ( w_23129 , \9187_b1 , \9187_b0 );
or ( \9189_b1 , \9177_b1 , \9188_b1 );
xor ( \9189_b0 , \9177_b0 , w_23130 );
not ( w_23130 , w_23131 );
and ( w_23131 , \9188_b1 , \9188_b0 );
or ( \9190_b1 , \9018_b1 , \9022_b1 );
not ( \9022_b1 , w_23132 );
and ( \9190_b0 , \9018_b0 , w_23133 );
and ( w_23132 , w_23133 , \9022_b0 );
or ( \9191_b1 , \9022_b1 , \9027_b1 );
not ( \9027_b1 , w_23134 );
and ( \9191_b0 , \9022_b0 , w_23135 );
and ( w_23134 , w_23135 , \9027_b0 );
or ( \9192_b1 , \9018_b1 , \9027_b1 );
not ( \9027_b1 , w_23136 );
and ( \9192_b0 , \9018_b0 , w_23137 );
and ( w_23136 , w_23137 , \9027_b0 );
or ( \9194_b1 , \9067_b1 , \9153_b1 );
not ( \9153_b1 , w_23138 );
and ( \9194_b0 , \9067_b0 , w_23139 );
and ( w_23138 , w_23139 , \9153_b0 );
or ( \9195_b1 , \9153_b1 , \9165_b1 );
not ( \9165_b1 , w_23140 );
and ( \9195_b0 , \9153_b0 , w_23141 );
and ( w_23140 , w_23141 , \9165_b0 );
or ( \9196_b1 , \9067_b1 , \9165_b1 );
not ( \9165_b1 , w_23142 );
and ( \9196_b0 , \9067_b0 , w_23143 );
and ( w_23142 , w_23143 , \9165_b0 );
or ( \9198_b1 , \9193_b1 , \9197_b1 );
xor ( \9198_b0 , \9193_b0 , w_23144 );
not ( w_23144 , w_23145 );
and ( w_23145 , \9197_b1 , \9197_b0 );
or ( \9199_b1 , \6029_b1 , \5852_b1 );
not ( \5852_b1 , w_23146 );
and ( \9199_b0 , \6029_b0 , w_23147 );
and ( w_23146 , w_23147 , \5852_b0 );
or ( \9200_b1 , \6041_b1 , \5850_b1 );
not ( \5850_b1 , w_23148 );
and ( \9200_b0 , \6041_b0 , w_23149 );
and ( w_23148 , w_23149 , \5850_b0 );
or ( \9201_b1 , \9199_b1 , w_23151 );
not ( w_23151 , w_23152 );
and ( \9201_b0 , \9199_b0 , w_23153 );
and ( w_23152 ,  , w_23153 );
buf ( w_23151 , \9200_b1 );
not ( w_23151 , w_23154 );
not (  , w_23155 );
and ( w_23154 , w_23155 , \9200_b0 );
or ( \9202_b1 , \9201_b1 , w_23156 );
xor ( \9202_b0 , \9201_b0 , w_23158 );
not ( w_23158 , w_23159 );
and ( w_23159 , w_23156 , w_23157 );
buf ( w_23156 , \5859_b1 );
not ( w_23156 , w_23160 );
not ( w_23157 , w_23161 );
and ( w_23160 , w_23161 , \5859_b0 );
or ( \9203_b1 , \6048_b1 , \5871_b1 );
not ( \5871_b1 , w_23162 );
and ( \9203_b0 , \6048_b0 , w_23163 );
and ( w_23162 , w_23163 , \5871_b0 );
or ( \9204_b1 , \6057_b1 , \5869_b1 );
not ( \5869_b1 , w_23164 );
and ( \9204_b0 , \6057_b0 , w_23165 );
and ( w_23164 , w_23165 , \5869_b0 );
or ( \9205_b1 , \9203_b1 , w_23167 );
not ( w_23167 , w_23168 );
and ( \9205_b0 , \9203_b0 , w_23169 );
and ( w_23168 ,  , w_23169 );
buf ( w_23167 , \9204_b1 );
not ( w_23167 , w_23170 );
not (  , w_23171 );
and ( w_23170 , w_23171 , \9204_b0 );
or ( \9206_b1 , \9205_b1 , w_23172 );
xor ( \9206_b0 , \9205_b0 , w_23174 );
not ( w_23174 , w_23175 );
and ( w_23175 , w_23172 , w_23173 );
buf ( w_23172 , \5878_b1 );
not ( w_23172 , w_23176 );
not ( w_23173 , w_23177 );
and ( w_23176 , w_23177 , \5878_b0 );
or ( \9207_b1 , \9202_b1 , \9206_b1 );
xor ( \9207_b0 , \9202_b0 , w_23178 );
not ( w_23178 , w_23179 );
and ( w_23179 , \9206_b1 , \9206_b0 );
or ( \9208_b1 , \6065_b1 , w_23181 );
not ( w_23181 , w_23182 );
and ( \9208_b0 , \6065_b0 , w_23183 );
and ( w_23182 ,  , w_23183 );
buf ( w_23181 , \5889_b1 );
not ( w_23181 , w_23184 );
not (  , w_23185 );
and ( w_23184 , w_23185 , \5889_b0 );
or ( \9209_b1 , \9208_b1 , w_23186 );
xor ( \9209_b0 , \9208_b0 , w_23188 );
not ( w_23188 , w_23189 );
and ( w_23189 , w_23186 , w_23187 );
buf ( w_23186 , \5898_b1 );
not ( w_23186 , w_23190 );
not ( w_23187 , w_23191 );
and ( w_23190 , w_23191 , \5898_b0 );
or ( \9210_b1 , \9207_b1 , \9209_b1 );
xor ( \9210_b0 , \9207_b0 , w_23192 );
not ( w_23192 , w_23193 );
and ( w_23193 , \9209_b1 , \9209_b0 );
or ( \9211_b1 , \5967_b1 , \5790_b1 );
not ( \5790_b1 , w_23194 );
and ( \9211_b0 , \5967_b0 , w_23195 );
and ( w_23194 , w_23195 , \5790_b0 );
or ( \9212_b1 , \5979_b1 , \5788_b1 );
not ( \5788_b1 , w_23196 );
and ( \9212_b0 , \5979_b0 , w_23197 );
and ( w_23196 , w_23197 , \5788_b0 );
or ( \9213_b1 , \9211_b1 , w_23199 );
not ( w_23199 , w_23200 );
and ( \9213_b0 , \9211_b0 , w_23201 );
and ( w_23200 ,  , w_23201 );
buf ( w_23199 , \9212_b1 );
not ( w_23199 , w_23202 );
not (  , w_23203 );
and ( w_23202 , w_23203 , \9212_b0 );
or ( \9214_b1 , \9213_b1 , w_23204 );
xor ( \9214_b0 , \9213_b0 , w_23206 );
not ( w_23206 , w_23207 );
and ( w_23207 , w_23204 , w_23205 );
buf ( w_23204 , \5797_b1 );
not ( w_23204 , w_23208 );
not ( w_23205 , w_23209 );
and ( w_23208 , w_23209 , \5797_b0 );
or ( \9215_b1 , \5986_b1 , \5809_b1 );
not ( \5809_b1 , w_23210 );
and ( \9215_b0 , \5986_b0 , w_23211 );
and ( w_23210 , w_23211 , \5809_b0 );
or ( \9216_b1 , \5998_b1 , \5807_b1 );
not ( \5807_b1 , w_23212 );
and ( \9216_b0 , \5998_b0 , w_23213 );
and ( w_23212 , w_23213 , \5807_b0 );
or ( \9217_b1 , \9215_b1 , w_23215 );
not ( w_23215 , w_23216 );
and ( \9217_b0 , \9215_b0 , w_23217 );
and ( w_23216 ,  , w_23217 );
buf ( w_23215 , \9216_b1 );
not ( w_23215 , w_23218 );
not (  , w_23219 );
and ( w_23218 , w_23219 , \9216_b0 );
or ( \9218_b1 , \9217_b1 , w_23220 );
xor ( \9218_b0 , \9217_b0 , w_23222 );
not ( w_23222 , w_23223 );
and ( w_23223 , w_23220 , w_23221 );
buf ( w_23220 , \5816_b1 );
not ( w_23220 , w_23224 );
not ( w_23221 , w_23225 );
and ( w_23224 , w_23225 , \5816_b0 );
or ( \9219_b1 , \9214_b1 , \9218_b1 );
xor ( \9219_b0 , \9214_b0 , w_23226 );
not ( w_23226 , w_23227 );
and ( w_23227 , \9218_b1 , \9218_b0 );
or ( \9220_b1 , \6006_b1 , \5829_b1 );
not ( \5829_b1 , w_23228 );
and ( \9220_b0 , \6006_b0 , w_23229 );
and ( w_23228 , w_23229 , \5829_b0 );
or ( \9221_b1 , \6018_b1 , \5827_b1 );
not ( \5827_b1 , w_23230 );
and ( \9221_b0 , \6018_b0 , w_23231 );
and ( w_23230 , w_23231 , \5827_b0 );
or ( \9222_b1 , \9220_b1 , w_23233 );
not ( w_23233 , w_23234 );
and ( \9222_b0 , \9220_b0 , w_23235 );
and ( w_23234 ,  , w_23235 );
buf ( w_23233 , \9221_b1 );
not ( w_23233 , w_23236 );
not (  , w_23237 );
and ( w_23236 , w_23237 , \9221_b0 );
or ( \9223_b1 , \9222_b1 , w_23238 );
xor ( \9223_b0 , \9222_b0 , w_23240 );
not ( w_23240 , w_23241 );
and ( w_23241 , w_23238 , w_23239 );
buf ( w_23238 , \5836_b1 );
not ( w_23238 , w_23242 );
not ( w_23239 , w_23243 );
and ( w_23242 , w_23243 , \5836_b0 );
or ( \9224_b1 , \9219_b1 , \9223_b1 );
xor ( \9224_b0 , \9219_b0 , w_23244 );
not ( w_23244 , w_23245 );
and ( w_23245 , \9223_b1 , \9223_b0 );
or ( \9225_b1 , \9210_b1 , w_23246 );
xor ( \9225_b0 , \9210_b0 , w_23248 );
not ( w_23248 , w_23249 );
and ( w_23249 , w_23246 , w_23247 );
buf ( w_23246 , \9224_b1 );
not ( w_23246 , w_23250 );
not ( w_23247 , w_23251 );
and ( w_23250 , w_23251 , \9224_b0 );
or ( \9226_b1 , \9141_b1 , \9145_b1 );
not ( \9145_b1 , w_23252 );
and ( \9226_b0 , \9141_b0 , w_23253 );
and ( w_23252 , w_23253 , \9145_b0 );
or ( \9227_b1 , \9145_b1 , \9150_b1 );
not ( \9150_b1 , w_23254 );
and ( \9227_b0 , \9145_b0 , w_23255 );
and ( w_23254 , w_23255 , \9150_b0 );
or ( \9228_b1 , \9141_b1 , \9150_b1 );
not ( \9150_b1 , w_23256 );
and ( \9228_b0 , \9141_b0 , w_23257 );
and ( w_23256 , w_23257 , \9150_b0 );
or ( \9230_b1 , \9126_b1 , \9130_b1 );
not ( \9130_b1 , w_23258 );
and ( \9230_b0 , \9126_b0 , w_23259 );
and ( w_23258 , w_23259 , \9130_b0 );
or ( \9231_b1 , \9130_b1 , \9135_b1 );
not ( \9135_b1 , w_23260 );
and ( \9231_b0 , \9130_b0 , w_23261 );
and ( w_23260 , w_23261 , \9135_b0 );
or ( \9232_b1 , \9126_b1 , \9135_b1 );
not ( \9135_b1 , w_23262 );
and ( \9232_b0 , \9126_b0 , w_23263 );
and ( w_23262 , w_23263 , \9135_b0 );
or ( \9234_b1 , \9229_b1 , \9233_b1 );
xor ( \9234_b0 , \9229_b0 , w_23264 );
not ( w_23264 , w_23265 );
and ( w_23265 , \9233_b1 , \9233_b0 );
or ( \9235_b1 , \9117_b1 , \9121_b1 );
not ( \9121_b1 , w_23266 );
and ( \9235_b0 , \9117_b0 , w_23267 );
and ( w_23266 , w_23267 , \9121_b0 );
or ( \9236_b1 , \9234_b1 , \9235_b1 );
xor ( \9236_b0 , \9234_b0 , w_23268 );
not ( w_23268 , w_23269 );
and ( w_23269 , \9235_b1 , \9235_b0 );
or ( \9237_b1 , \9225_b1 , \9236_b1 );
xor ( \9237_b0 , \9225_b0 , w_23270 );
not ( w_23270 , w_23271 );
and ( w_23271 , \9236_b1 , \9236_b0 );
or ( \9238_b1 , \9101_b1 , \9105_b1 );
not ( \9105_b1 , w_23272 );
and ( \9238_b0 , \9101_b0 , w_23273 );
and ( w_23272 , w_23273 , \9105_b0 );
or ( \9239_b1 , \9105_b1 , \9110_b1 );
not ( \9110_b1 , w_23274 );
and ( \9239_b0 , \9105_b0 , w_23275 );
and ( w_23274 , w_23275 , \9110_b0 );
or ( \9240_b1 , \9101_b1 , \9110_b1 );
not ( \9110_b1 , w_23276 );
and ( \9240_b0 , \9101_b0 , w_23277 );
and ( w_23276 , w_23277 , \9110_b0 );
or ( \9242_b1 , \9089_b1 , \9093_b1 );
not ( \9093_b1 , w_23278 );
and ( \9242_b0 , \9089_b0 , w_23279 );
and ( w_23278 , w_23279 , \9093_b0 );
or ( \9243_b1 , \9093_b1 , \9098_b1 );
not ( \9098_b1 , w_23280 );
and ( \9243_b0 , \9093_b0 , w_23281 );
and ( w_23280 , w_23281 , \9098_b0 );
or ( \9244_b1 , \9089_b1 , \9098_b1 );
not ( \9098_b1 , w_23282 );
and ( \9244_b0 , \9089_b0 , w_23283 );
and ( w_23282 , w_23283 , \9098_b0 );
or ( \9246_b1 , \9241_b1 , \9245_b1 );
xor ( \9246_b0 , \9241_b0 , w_23284 );
not ( w_23284 , w_23285 );
and ( w_23285 , \9245_b1 , \9245_b0 );
or ( \9247_b1 , \9075_b1 , \9079_b1 );
not ( \9079_b1 , w_23286 );
and ( \9247_b0 , \9075_b0 , w_23287 );
and ( w_23286 , w_23287 , \9079_b0 );
or ( \9248_b1 , \9079_b1 , \9084_b1 );
not ( \9084_b1 , w_23288 );
and ( \9248_b0 , \9079_b0 , w_23289 );
and ( w_23288 , w_23289 , \9084_b0 );
or ( \9249_b1 , \9075_b1 , \9084_b1 );
not ( \9084_b1 , w_23290 );
and ( \9249_b0 , \9075_b0 , w_23291 );
and ( w_23290 , w_23291 , \9084_b0 );
or ( \9251_b1 , \9246_b1 , \9250_b1 );
xor ( \9251_b0 , \9246_b0 , w_23292 );
not ( w_23292 , w_23293 );
and ( w_23293 , \9250_b1 , \9250_b0 );
or ( \9252_b1 , \9237_b1 , \9251_b1 );
xor ( \9252_b0 , \9237_b0 , w_23294 );
not ( w_23294 , w_23295 );
and ( w_23295 , \9251_b1 , \9251_b0 );
or ( \9253_b1 , \9085_b1 , \9099_b1 );
not ( \9099_b1 , w_23296 );
and ( \9253_b0 , \9085_b0 , w_23297 );
and ( w_23296 , w_23297 , \9099_b0 );
or ( \9254_b1 , \9099_b1 , \9111_b1 );
not ( \9111_b1 , w_23298 );
and ( \9254_b0 , \9099_b0 , w_23299 );
and ( w_23298 , w_23299 , \9111_b0 );
or ( \9255_b1 , \9085_b1 , \9111_b1 );
not ( \9111_b1 , w_23300 );
and ( \9255_b0 , \9085_b0 , w_23301 );
and ( w_23300 , w_23301 , \9111_b0 );
or ( \9257_b1 , \5737_b1 , \7061_b1 );
not ( \7061_b1 , w_23302 );
and ( \9257_b0 , \5737_b0 , w_23303 );
and ( w_23302 , w_23303 , \7061_b0 );
buf ( \9258_b1 , \9257_b1 );
not ( \9258_b1 , w_23304 );
not ( \9258_b0 , w_23305 );
and ( w_23304 , w_23305 , \9257_b0 );
or ( \9259_b1 , \9258_b1 , w_23306 );
xor ( \9259_b0 , \9258_b0 , w_23308 );
not ( w_23308 , w_23309 );
and ( w_23309 , w_23306 , w_23307 );
buf ( w_23306 , \7067_b1 );
not ( w_23306 , w_23310 );
not ( w_23307 , w_23311 );
and ( w_23310 , w_23311 , \7067_b0 );
or ( \9260_b1 , \5898_b1 , \9259_b1 );
xor ( \9260_b0 , \5898_b0 , w_23312 );
not ( w_23312 , w_23313 );
and ( w_23313 , \9259_b1 , \9259_b0 );
or ( \9261_b1 , \5758_b1 , \7082_b1 );
not ( \7082_b1 , w_23314 );
and ( \9261_b0 , \5758_b0 , w_23315 );
and ( w_23314 , w_23315 , \7082_b0 );
or ( \9262_b1 , \5770_b1 , \7080_b1 );
not ( \7080_b1 , w_23316 );
and ( \9262_b0 , \5770_b0 , w_23317 );
and ( w_23316 , w_23317 , \7080_b0 );
or ( \9263_b1 , \9261_b1 , w_23319 );
not ( w_23319 , w_23320 );
and ( \9263_b0 , \9261_b0 , w_23321 );
and ( w_23320 ,  , w_23321 );
buf ( w_23319 , \9262_b1 );
not ( w_23319 , w_23322 );
not (  , w_23323 );
and ( w_23322 , w_23323 , \9262_b0 );
or ( \9264_b1 , \9263_b1 , w_23324 );
xor ( \9264_b0 , \9263_b0 , w_23326 );
not ( w_23326 , w_23327 );
and ( w_23327 , w_23324 , w_23325 );
buf ( w_23324 , \7088_b1 );
not ( w_23324 , w_23328 );
not ( w_23325 , w_23329 );
and ( w_23328 , w_23329 , \7088_b0 );
or ( \9265_b1 , \9260_b1 , \9264_b1 );
xor ( \9265_b0 , \9260_b0 , w_23330 );
not ( w_23330 , w_23331 );
and ( w_23331 , \9264_b1 , \9264_b0 );
or ( \9266_b1 , \9256_b1 , \9265_b1 );
xor ( \9266_b0 , \9256_b0 , w_23332 );
not ( w_23332 , w_23333 );
and ( w_23333 , \9265_b1 , \9265_b0 );
or ( \9267_b1 , \5906_b1 , \7203_b1 );
not ( \7203_b1 , w_23334 );
and ( \9267_b0 , \5906_b0 , w_23335 );
and ( w_23334 , w_23335 , \7203_b0 );
or ( \9268_b1 , \5918_b1 , \7201_b1 );
not ( \7201_b1 , w_23336 );
and ( \9268_b0 , \5918_b0 , w_23337 );
and ( w_23336 , w_23337 , \7201_b0 );
or ( \9269_b1 , \9267_b1 , w_23339 );
not ( w_23339 , w_23340 );
and ( \9269_b0 , \9267_b0 , w_23341 );
and ( w_23340 ,  , w_23341 );
buf ( w_23339 , \9268_b1 );
not ( w_23339 , w_23342 );
not (  , w_23343 );
and ( w_23342 , w_23343 , \9268_b0 );
or ( \9270_b1 , \9269_b1 , w_23344 );
xor ( \9270_b0 , \9269_b0 , w_23346 );
not ( w_23346 , w_23347 );
and ( w_23347 , w_23344 , w_23345 );
buf ( w_23344 , \6824_b1 );
not ( w_23344 , w_23348 );
not ( w_23345 , w_23349 );
and ( w_23348 , w_23349 , \6824_b0 );
or ( \9271_b1 , \5925_b1 , \5750_b1 );
not ( \5750_b1 , w_23350 );
and ( \9271_b0 , \5925_b0 , w_23351 );
and ( w_23350 , w_23351 , \5750_b0 );
or ( \9272_b1 , \5937_b1 , \5748_b1 );
not ( \5748_b1 , w_23352 );
and ( \9272_b0 , \5937_b0 , w_23353 );
and ( w_23352 , w_23353 , \5748_b0 );
or ( \9273_b1 , \9271_b1 , w_23355 );
not ( w_23355 , w_23356 );
and ( \9273_b0 , \9271_b0 , w_23357 );
and ( w_23356 ,  , w_23357 );
buf ( w_23355 , \9272_b1 );
not ( w_23355 , w_23358 );
not (  , w_23359 );
and ( w_23358 , w_23359 , \9272_b0 );
or ( \9274_b1 , \9273_b1 , w_23360 );
xor ( \9274_b0 , \9273_b0 , w_23362 );
not ( w_23362 , w_23363 );
and ( w_23363 , w_23360 , w_23361 );
buf ( w_23360 , \5755_b1 );
not ( w_23360 , w_23364 );
not ( w_23361 , w_23365 );
and ( w_23364 , w_23365 , \5755_b0 );
or ( \9275_b1 , \9270_b1 , \9274_b1 );
xor ( \9275_b0 , \9270_b0 , w_23366 );
not ( w_23366 , w_23367 );
and ( w_23367 , \9274_b1 , \9274_b0 );
or ( \9276_b1 , \5945_b1 , \5768_b1 );
not ( \5768_b1 , w_23368 );
and ( \9276_b0 , \5945_b0 , w_23369 );
and ( w_23368 , w_23369 , \5768_b0 );
or ( \9277_b1 , \5957_b1 , \5766_b1 );
not ( \5766_b1 , w_23370 );
and ( \9277_b0 , \5957_b0 , w_23371 );
and ( w_23370 , w_23371 , \5766_b0 );
or ( \9278_b1 , \9276_b1 , w_23373 );
not ( w_23373 , w_23374 );
and ( \9278_b0 , \9276_b0 , w_23375 );
and ( w_23374 ,  , w_23375 );
buf ( w_23373 , \9277_b1 );
not ( w_23373 , w_23376 );
not (  , w_23377 );
and ( w_23376 , w_23377 , \9277_b0 );
or ( \9279_b1 , \9278_b1 , w_23378 );
xor ( \9279_b0 , \9278_b0 , w_23380 );
not ( w_23380 , w_23381 );
and ( w_23381 , w_23378 , w_23379 );
buf ( w_23378 , \5775_b1 );
not ( w_23378 , w_23382 );
not ( w_23379 , w_23383 );
and ( w_23382 , w_23383 , \5775_b0 );
or ( \9280_b1 , \9275_b1 , \9279_b1 );
xor ( \9280_b0 , \9275_b0 , w_23384 );
not ( w_23384 , w_23385 );
and ( w_23385 , \9279_b1 , \9279_b0 );
or ( \9281_b1 , \5842_b1 , \7157_b1 );
not ( \7157_b1 , w_23386 );
and ( \9281_b0 , \5842_b0 , w_23387 );
and ( w_23386 , w_23387 , \7157_b0 );
or ( \9282_b1 , \5854_b1 , \7155_b1 );
not ( \7155_b1 , w_23388 );
and ( \9282_b0 , \5854_b0 , w_23389 );
and ( w_23388 , w_23389 , \7155_b0 );
or ( \9283_b1 , \9281_b1 , w_23391 );
not ( w_23391 , w_23392 );
and ( \9283_b0 , \9281_b0 , w_23393 );
and ( w_23392 ,  , w_23393 );
buf ( w_23391 , \9282_b1 );
not ( w_23391 , w_23394 );
not (  , w_23395 );
and ( w_23394 , w_23395 , \9282_b0 );
or ( \9284_b1 , \9283_b1 , w_23396 );
xor ( \9284_b0 , \9283_b0 , w_23398 );
not ( w_23398 , w_23399 );
and ( w_23399 , w_23396 , w_23397 );
buf ( w_23396 , \7163_b1 );
not ( w_23396 , w_23400 );
not ( w_23397 , w_23401 );
and ( w_23400 , w_23401 , \7163_b0 );
or ( \9285_b1 , \5861_b1 , \7175_b1 );
not ( \7175_b1 , w_23402 );
and ( \9285_b0 , \5861_b0 , w_23403 );
and ( w_23402 , w_23403 , \7175_b0 );
or ( \9286_b1 , \5873_b1 , \7173_b1 );
not ( \7173_b1 , w_23404 );
and ( \9286_b0 , \5873_b0 , w_23405 );
and ( w_23404 , w_23405 , \7173_b0 );
or ( \9287_b1 , \9285_b1 , w_23407 );
not ( w_23407 , w_23408 );
and ( \9287_b0 , \9285_b0 , w_23409 );
and ( w_23408 ,  , w_23409 );
buf ( w_23407 , \9286_b1 );
not ( w_23407 , w_23410 );
not (  , w_23411 );
and ( w_23410 , w_23411 , \9286_b0 );
or ( \9288_b1 , \9287_b1 , w_23412 );
xor ( \9288_b0 , \9287_b0 , w_23414 );
not ( w_23414 , w_23415 );
and ( w_23415 , w_23412 , w_23413 );
buf ( w_23412 , \7181_b1 );
not ( w_23412 , w_23416 );
not ( w_23413 , w_23417 );
and ( w_23416 , w_23417 , \7181_b0 );
or ( \9289_b1 , \9284_b1 , \9288_b1 );
xor ( \9289_b0 , \9284_b0 , w_23418 );
not ( w_23418 , w_23419 );
and ( w_23419 , \9288_b1 , \9288_b0 );
or ( \9290_b1 , \5881_b1 , \7192_b1 );
not ( \7192_b1 , w_23420 );
and ( \9290_b0 , \5881_b0 , w_23421 );
and ( w_23420 , w_23421 , \7192_b0 );
or ( \9291_b1 , \5893_b1 , \7190_b1 );
not ( \7190_b1 , w_23422 );
and ( \9291_b0 , \5893_b0 , w_23423 );
and ( w_23422 , w_23423 , \7190_b0 );
or ( \9292_b1 , \9290_b1 , w_23425 );
not ( w_23425 , w_23426 );
and ( \9292_b0 , \9290_b0 , w_23427 );
and ( w_23426 ,  , w_23427 );
buf ( w_23425 , \9291_b1 );
not ( w_23425 , w_23428 );
not (  , w_23429 );
and ( w_23428 , w_23429 , \9291_b0 );
or ( \9293_b1 , \9292_b1 , w_23430 );
xor ( \9293_b0 , \9292_b0 , w_23432 );
not ( w_23432 , w_23433 );
and ( w_23433 , w_23430 , w_23431 );
buf ( w_23430 , \7198_b1 );
not ( w_23430 , w_23434 );
not ( w_23431 , w_23435 );
and ( w_23434 , w_23435 , \7198_b0 );
or ( \9294_b1 , \9289_b1 , \9293_b1 );
xor ( \9294_b0 , \9289_b0 , w_23436 );
not ( w_23436 , w_23437 );
and ( w_23437 , \9293_b1 , \9293_b0 );
or ( \9295_b1 , \9280_b1 , \9294_b1 );
xor ( \9295_b0 , \9280_b0 , w_23438 );
not ( w_23438 , w_23439 );
and ( w_23439 , \9294_b1 , \9294_b0 );
or ( \9296_b1 , \5780_b1 , \7099_b1 );
not ( \7099_b1 , w_23440 );
and ( \9296_b0 , \5780_b0 , w_23441 );
and ( w_23440 , w_23441 , \7099_b0 );
or ( \9297_b1 , \5792_b1 , \7097_b1 );
not ( \7097_b1 , w_23442 );
and ( \9297_b0 , \5792_b0 , w_23443 );
and ( w_23442 , w_23443 , \7097_b0 );
or ( \9298_b1 , \9296_b1 , w_23445 );
not ( w_23445 , w_23446 );
and ( \9298_b0 , \9296_b0 , w_23447 );
and ( w_23446 ,  , w_23447 );
buf ( w_23445 , \9297_b1 );
not ( w_23445 , w_23448 );
not (  , w_23449 );
and ( w_23448 , w_23449 , \9297_b0 );
or ( \9299_b1 , \9298_b1 , w_23450 );
xor ( \9299_b0 , \9298_b0 , w_23452 );
not ( w_23452 , w_23453 );
and ( w_23453 , w_23450 , w_23451 );
buf ( w_23450 , \7105_b1 );
not ( w_23450 , w_23454 );
not ( w_23451 , w_23455 );
and ( w_23454 , w_23455 , \7105_b0 );
or ( \9300_b1 , \5799_b1 , \7117_b1 );
not ( \7117_b1 , w_23456 );
and ( \9300_b0 , \5799_b0 , w_23457 );
and ( w_23456 , w_23457 , \7117_b0 );
or ( \9301_b1 , \5811_b1 , \7115_b1 );
not ( \7115_b1 , w_23458 );
and ( \9301_b0 , \5811_b0 , w_23459 );
and ( w_23458 , w_23459 , \7115_b0 );
or ( \9302_b1 , \9300_b1 , w_23461 );
not ( w_23461 , w_23462 );
and ( \9302_b0 , \9300_b0 , w_23463 );
and ( w_23462 ,  , w_23463 );
buf ( w_23461 , \9301_b1 );
not ( w_23461 , w_23464 );
not (  , w_23465 );
and ( w_23464 , w_23465 , \9301_b0 );
or ( \9303_b1 , \9302_b1 , w_23466 );
xor ( \9303_b0 , \9302_b0 , w_23468 );
not ( w_23468 , w_23469 );
and ( w_23469 , w_23466 , w_23467 );
buf ( w_23466 , \7123_b1 );
not ( w_23466 , w_23470 );
not ( w_23467 , w_23471 );
and ( w_23470 , w_23471 , \7123_b0 );
or ( \9304_b1 , \9299_b1 , \9303_b1 );
xor ( \9304_b0 , \9299_b0 , w_23472 );
not ( w_23472 , w_23473 );
and ( w_23473 , \9303_b1 , \9303_b0 );
or ( \9305_b1 , \5819_b1 , \7140_b1 );
not ( \7140_b1 , w_23474 );
and ( \9305_b0 , \5819_b0 , w_23475 );
and ( w_23474 , w_23475 , \7140_b0 );
or ( \9306_b1 , \5831_b1 , \7138_b1 );
not ( \7138_b1 , w_23476 );
and ( \9306_b0 , \5831_b0 , w_23477 );
and ( w_23476 , w_23477 , \7138_b0 );
or ( \9307_b1 , \9305_b1 , w_23479 );
not ( w_23479 , w_23480 );
and ( \9307_b0 , \9305_b0 , w_23481 );
and ( w_23480 ,  , w_23481 );
buf ( w_23479 , \9306_b1 );
not ( w_23479 , w_23482 );
not (  , w_23483 );
and ( w_23482 , w_23483 , \9306_b0 );
or ( \9308_b1 , \9307_b1 , w_23484 );
xor ( \9308_b0 , \9307_b0 , w_23486 );
not ( w_23486 , w_23487 );
and ( w_23487 , w_23484 , w_23485 );
buf ( w_23484 , \7146_b1 );
not ( w_23484 , w_23488 );
not ( w_23485 , w_23489 );
and ( w_23488 , w_23489 , \7146_b0 );
or ( \9309_b1 , \9304_b1 , \9308_b1 );
xor ( \9309_b0 , \9304_b0 , w_23490 );
not ( w_23490 , w_23491 );
and ( w_23491 , \9308_b1 , \9308_b0 );
or ( \9310_b1 , \9295_b1 , \9309_b1 );
xor ( \9310_b0 , \9295_b0 , w_23492 );
not ( w_23492 , w_23493 );
and ( w_23493 , \9309_b1 , \9309_b0 );
or ( \9311_b1 , \9266_b1 , \9310_b1 );
xor ( \9311_b0 , \9266_b0 , w_23494 );
not ( w_23494 , w_23495 );
and ( w_23495 , \9310_b1 , \9310_b0 );
or ( \9312_b1 , \9252_b1 , \9311_b1 );
xor ( \9312_b0 , \9252_b0 , w_23496 );
not ( w_23496 , w_23497 );
and ( w_23497 , \9311_b1 , \9311_b0 );
or ( \9313_b1 , \9056_b1 , \9060_b1 );
not ( \9060_b1 , w_23498 );
and ( \9313_b0 , \9056_b0 , w_23499 );
and ( w_23498 , w_23499 , \9060_b0 );
or ( \9314_b1 , \9060_b1 , \9065_b1 );
not ( \9065_b1 , w_23500 );
and ( \9314_b0 , \9060_b0 , w_23501 );
and ( w_23500 , w_23501 , \9065_b0 );
or ( \9315_b1 , \9056_b1 , \9065_b1 );
not ( \9065_b1 , w_23502 );
and ( \9315_b0 , \9056_b0 , w_23503 );
and ( w_23502 , w_23503 , \9065_b0 );
or ( \9317_b1 , \9042_b1 , \9046_b1 );
not ( \9046_b1 , w_23504 );
and ( \9317_b0 , \9042_b0 , w_23505 );
and ( w_23504 , w_23505 , \9046_b0 );
or ( \9318_b1 , \9046_b1 , \9051_b1 );
not ( \9051_b1 , w_23506 );
and ( \9318_b0 , \9046_b0 , w_23507 );
and ( w_23506 , w_23507 , \9051_b0 );
or ( \9319_b1 , \9042_b1 , \9051_b1 );
not ( \9051_b1 , w_23508 );
and ( \9319_b0 , \9042_b0 , w_23509 );
and ( w_23508 , w_23509 , \9051_b0 );
or ( \9321_b1 , \9316_b1 , \9320_b1 );
xor ( \9321_b0 , \9316_b0 , w_23510 );
not ( w_23510 , w_23511 );
and ( w_23511 , \9320_b1 , \9320_b0 );
or ( \9322_b1 , \9122_b1 , \9136_b1 );
not ( \9136_b1 , w_23512 );
and ( \9322_b0 , \9122_b0 , w_23513 );
and ( w_23512 , w_23513 , \9136_b0 );
or ( \9323_b1 , \9136_b1 , \9151_b1 );
not ( \9151_b1 , w_23514 );
and ( \9323_b0 , \9136_b0 , w_23515 );
and ( w_23514 , w_23515 , \9151_b0 );
or ( \9324_b1 , \9122_b1 , \9151_b1 );
not ( \9151_b1 , w_23516 );
and ( \9324_b0 , \9122_b0 , w_23517 );
and ( w_23516 , w_23517 , \9151_b0 );
or ( \9326_b1 , \9321_b1 , \9325_b1 );
xor ( \9326_b0 , \9321_b0 , w_23518 );
not ( w_23518 , w_23519 );
and ( w_23519 , \9325_b1 , \9325_b0 );
or ( \9327_b1 , \9312_b1 , \9326_b1 );
xor ( \9327_b0 , \9312_b0 , w_23520 );
not ( w_23520 , w_23521 );
and ( w_23521 , \9326_b1 , \9326_b0 );
or ( \9328_b1 , \9198_b1 , \9327_b1 );
xor ( \9328_b0 , \9198_b0 , w_23522 );
not ( w_23522 , w_23523 );
and ( w_23523 , \9327_b1 , \9327_b0 );
or ( \9329_b1 , \9189_b1 , \9328_b1 );
xor ( \9329_b0 , \9189_b0 , w_23524 );
not ( w_23524 , w_23525 );
and ( w_23525 , \9328_b1 , \9328_b0 );
or ( \9330_b1 , \9014_b1 , \9028_b1 );
not ( \9028_b1 , w_23526 );
and ( \9330_b0 , \9014_b0 , w_23527 );
and ( w_23526 , w_23527 , \9028_b0 );
or ( \9331_b1 , \9028_b1 , \9167_b1 );
not ( \9167_b1 , w_23528 );
and ( \9331_b0 , \9028_b0 , w_23529 );
and ( w_23528 , w_23529 , \9167_b0 );
or ( \9332_b1 , \9014_b1 , \9167_b1 );
not ( \9167_b1 , w_23530 );
and ( \9332_b0 , \9014_b0 , w_23531 );
and ( w_23530 , w_23531 , \9167_b0 );
or ( \9334_b1 , \9329_b1 , w_23533 );
not ( w_23533 , w_23534 );
and ( \9334_b0 , \9329_b0 , w_23535 );
and ( w_23534 ,  , w_23535 );
buf ( w_23533 , \9333_b1 );
not ( w_23533 , w_23536 );
not (  , w_23537 );
and ( w_23536 , w_23537 , \9333_b0 );
or ( \9335_b1 , \9173_b1 , w_23539 );
not ( w_23539 , w_23540 );
and ( \9335_b0 , \9173_b0 , w_23541 );
and ( w_23540 ,  , w_23541 );
buf ( w_23539 , \9334_b1 );
not ( w_23539 , w_23542 );
not (  , w_23543 );
and ( w_23542 , w_23543 , \9334_b0 );
or ( \9336_b1 , \9193_b1 , \9197_b1 );
not ( \9197_b1 , w_23544 );
and ( \9336_b0 , \9193_b0 , w_23545 );
and ( w_23544 , w_23545 , \9197_b0 );
or ( \9337_b1 , \9197_b1 , \9327_b1 );
not ( \9327_b1 , w_23546 );
and ( \9337_b0 , \9197_b0 , w_23547 );
and ( w_23546 , w_23547 , \9327_b0 );
or ( \9338_b1 , \9193_b1 , \9327_b1 );
not ( \9327_b1 , w_23548 );
and ( \9338_b0 , \9193_b0 , w_23549 );
and ( w_23548 , w_23549 , \9327_b0 );
or ( \9340_b1 , \9316_b1 , \9320_b1 );
not ( \9320_b1 , w_23550 );
and ( \9340_b0 , \9316_b0 , w_23551 );
and ( w_23550 , w_23551 , \9320_b0 );
or ( \9341_b1 , \9320_b1 , \9325_b1 );
not ( \9325_b1 , w_23552 );
and ( \9341_b0 , \9320_b0 , w_23553 );
and ( w_23552 , w_23553 , \9325_b0 );
or ( \9342_b1 , \9316_b1 , \9325_b1 );
not ( \9325_b1 , w_23554 );
and ( \9342_b0 , \9316_b0 , w_23555 );
and ( w_23554 , w_23555 , \9325_b0 );
or ( \9344_b1 , \9256_b1 , \9265_b1 );
not ( \9265_b1 , w_23556 );
and ( \9344_b0 , \9256_b0 , w_23557 );
and ( w_23556 , w_23557 , \9265_b0 );
or ( \9345_b1 , \9265_b1 , \9310_b1 );
not ( \9310_b1 , w_23558 );
and ( \9345_b0 , \9265_b0 , w_23559 );
and ( w_23558 , w_23559 , \9310_b0 );
or ( \9346_b1 , \9256_b1 , \9310_b1 );
not ( \9310_b1 , w_23560 );
and ( \9346_b0 , \9256_b0 , w_23561 );
and ( w_23560 , w_23561 , \9310_b0 );
or ( \9348_b1 , \9343_b1 , \9347_b1 );
xor ( \9348_b0 , \9343_b0 , w_23562 );
not ( w_23562 , w_23563 );
and ( w_23563 , \9347_b1 , \9347_b0 );
or ( \9349_b1 , \9225_b1 , \9236_b1 );
not ( \9236_b1 , w_23564 );
and ( \9349_b0 , \9225_b0 , w_23565 );
and ( w_23564 , w_23565 , \9236_b0 );
or ( \9350_b1 , \9236_b1 , \9251_b1 );
not ( \9251_b1 , w_23566 );
and ( \9350_b0 , \9236_b0 , w_23567 );
and ( w_23566 , w_23567 , \9251_b0 );
or ( \9351_b1 , \9225_b1 , \9251_b1 );
not ( \9251_b1 , w_23568 );
and ( \9351_b0 , \9225_b0 , w_23569 );
and ( w_23568 , w_23569 , \9251_b0 );
or ( \9353_b1 , \9348_b1 , \9352_b1 );
xor ( \9353_b0 , \9348_b0 , w_23570 );
not ( w_23570 , w_23571 );
and ( w_23571 , \9352_b1 , \9352_b0 );
or ( \9354_b1 , \9339_b1 , \9353_b1 );
xor ( \9354_b0 , \9339_b0 , w_23572 );
not ( w_23572 , w_23573 );
and ( w_23573 , \9353_b1 , \9353_b0 );
or ( \9355_b1 , \9181_b1 , \9185_b1 );
not ( \9185_b1 , w_23574 );
and ( \9355_b0 , \9181_b0 , w_23575 );
and ( w_23574 , w_23575 , \9185_b0 );
or ( \9356_b1 , \9185_b1 , \9187_b1 );
not ( \9187_b1 , w_23576 );
and ( \9356_b0 , \9185_b0 , w_23577 );
and ( w_23576 , w_23577 , \9187_b0 );
or ( \9357_b1 , \9181_b1 , \9187_b1 );
not ( \9187_b1 , w_23578 );
and ( \9357_b0 , \9181_b0 , w_23579 );
and ( w_23578 , w_23579 , \9187_b0 );
or ( \9359_b1 , \9252_b1 , \9311_b1 );
not ( \9311_b1 , w_23580 );
and ( \9359_b0 , \9252_b0 , w_23581 );
and ( w_23580 , w_23581 , \9311_b0 );
or ( \9360_b1 , \9311_b1 , \9326_b1 );
not ( \9326_b1 , w_23582 );
and ( \9360_b0 , \9311_b0 , w_23583 );
and ( w_23582 , w_23583 , \9326_b0 );
or ( \9361_b1 , \9252_b1 , \9326_b1 );
not ( \9326_b1 , w_23584 );
and ( \9361_b0 , \9252_b0 , w_23585 );
and ( w_23584 , w_23585 , \9326_b0 );
or ( \9363_b1 , \9358_b1 , \9362_b1 );
xor ( \9363_b0 , \9358_b0 , w_23586 );
not ( w_23586 , w_23587 );
and ( w_23587 , \9362_b1 , \9362_b0 );
or ( \9364_b1 , \9270_b1 , \9274_b1 );
not ( \9274_b1 , w_23588 );
and ( \9364_b0 , \9270_b0 , w_23589 );
and ( w_23588 , w_23589 , \9274_b0 );
or ( \9365_b1 , \9274_b1 , \9279_b1 );
not ( \9279_b1 , w_23590 );
and ( \9365_b0 , \9274_b0 , w_23591 );
and ( w_23590 , w_23591 , \9279_b0 );
or ( \9366_b1 , \9270_b1 , \9279_b1 );
not ( \9279_b1 , w_23592 );
and ( \9366_b0 , \9270_b0 , w_23593 );
and ( w_23592 , w_23593 , \9279_b0 );
or ( \9368_b1 , \9214_b1 , \9218_b1 );
not ( \9218_b1 , w_23594 );
and ( \9368_b0 , \9214_b0 , w_23595 );
and ( w_23594 , w_23595 , \9218_b0 );
or ( \9369_b1 , \9218_b1 , \9223_b1 );
not ( \9223_b1 , w_23596 );
and ( \9369_b0 , \9218_b0 , w_23597 );
and ( w_23596 , w_23597 , \9223_b0 );
or ( \9370_b1 , \9214_b1 , \9223_b1 );
not ( \9223_b1 , w_23598 );
and ( \9370_b0 , \9214_b0 , w_23599 );
and ( w_23598 , w_23599 , \9223_b0 );
or ( \9372_b1 , \9367_b1 , \9371_b1 );
xor ( \9372_b0 , \9367_b0 , w_23600 );
not ( w_23600 , w_23601 );
and ( w_23601 , \9371_b1 , \9371_b0 );
or ( \9373_b1 , \9202_b1 , \9206_b1 );
not ( \9206_b1 , w_23602 );
and ( \9373_b0 , \9202_b0 , w_23603 );
and ( w_23602 , w_23603 , \9206_b0 );
or ( \9374_b1 , \9206_b1 , \9209_b1 );
not ( \9209_b1 , w_23604 );
and ( \9374_b0 , \9206_b0 , w_23605 );
and ( w_23604 , w_23605 , \9209_b0 );
or ( \9375_b1 , \9202_b1 , \9209_b1 );
not ( \9209_b1 , w_23606 );
and ( \9375_b0 , \9202_b0 , w_23607 );
and ( w_23606 , w_23607 , \9209_b0 );
or ( \9377_b1 , \9372_b1 , \9376_b1 );
xor ( \9377_b0 , \9372_b0 , w_23608 );
not ( w_23608 , w_23609 );
and ( w_23609 , \9376_b1 , \9376_b0 );
or ( \9378_b1 , \5898_b1 , \9259_b1 );
not ( \9259_b1 , w_23610 );
and ( \9378_b0 , \5898_b0 , w_23611 );
and ( w_23610 , w_23611 , \9259_b0 );
or ( \9379_b1 , \9259_b1 , \9264_b1 );
not ( \9264_b1 , w_23612 );
and ( \9379_b0 , \9259_b0 , w_23613 );
and ( w_23612 , w_23613 , \9264_b0 );
or ( \9380_b1 , \5898_b1 , \9264_b1 );
not ( \9264_b1 , w_23614 );
and ( \9380_b0 , \5898_b0 , w_23615 );
and ( w_23614 , w_23615 , \9264_b0 );
or ( \9382_b1 , \9299_b1 , \9303_b1 );
not ( \9303_b1 , w_23616 );
and ( \9382_b0 , \9299_b0 , w_23617 );
and ( w_23616 , w_23617 , \9303_b0 );
or ( \9383_b1 , \9303_b1 , \9308_b1 );
not ( \9308_b1 , w_23618 );
and ( \9383_b0 , \9303_b0 , w_23619 );
and ( w_23618 , w_23619 , \9308_b0 );
or ( \9384_b1 , \9299_b1 , \9308_b1 );
not ( \9308_b1 , w_23620 );
and ( \9384_b0 , \9299_b0 , w_23621 );
and ( w_23620 , w_23621 , \9308_b0 );
or ( \9386_b1 , \9381_b1 , \9385_b1 );
xor ( \9386_b0 , \9381_b0 , w_23622 );
not ( w_23622 , w_23623 );
and ( w_23623 , \9385_b1 , \9385_b0 );
or ( \9387_b1 , \9284_b1 , \9288_b1 );
not ( \9288_b1 , w_23624 );
and ( \9387_b0 , \9284_b0 , w_23625 );
and ( w_23624 , w_23625 , \9288_b0 );
or ( \9388_b1 , \9288_b1 , \9293_b1 );
not ( \9293_b1 , w_23626 );
and ( \9388_b0 , \9288_b0 , w_23627 );
and ( w_23626 , w_23627 , \9293_b0 );
or ( \9389_b1 , \9284_b1 , \9293_b1 );
not ( \9293_b1 , w_23628 );
and ( \9389_b0 , \9284_b0 , w_23629 );
and ( w_23628 , w_23629 , \9293_b0 );
or ( \9391_b1 , \9386_b1 , \9390_b1 );
xor ( \9391_b0 , \9386_b0 , w_23630 );
not ( w_23630 , w_23631 );
and ( w_23631 , \9390_b1 , \9390_b0 );
or ( \9392_b1 , \9377_b1 , \9391_b1 );
xor ( \9392_b0 , \9377_b0 , w_23632 );
not ( w_23632 , w_23633 );
and ( w_23633 , \9391_b1 , \9391_b0 );
or ( \9393_b1 , \9280_b1 , \9294_b1 );
not ( \9294_b1 , w_23634 );
and ( \9393_b0 , \9280_b0 , w_23635 );
and ( w_23634 , w_23635 , \9294_b0 );
or ( \9394_b1 , \9294_b1 , \9309_b1 );
not ( \9309_b1 , w_23636 );
and ( \9394_b0 , \9294_b0 , w_23637 );
and ( w_23636 , w_23637 , \9309_b0 );
or ( \9395_b1 , \9280_b1 , \9309_b1 );
not ( \9309_b1 , w_23638 );
and ( \9395_b0 , \9280_b0 , w_23639 );
and ( w_23638 , w_23639 , \9309_b0 );
or ( \9397_b1 , \5873_b1 , \7175_b1 );
not ( \7175_b1 , w_23640 );
and ( \9397_b0 , \5873_b0 , w_23641 );
and ( w_23640 , w_23641 , \7175_b0 );
or ( \9398_b1 , \5842_b1 , \7173_b1 );
not ( \7173_b1 , w_23642 );
and ( \9398_b0 , \5842_b0 , w_23643 );
and ( w_23642 , w_23643 , \7173_b0 );
or ( \9399_b1 , \9397_b1 , w_23645 );
not ( w_23645 , w_23646 );
and ( \9399_b0 , \9397_b0 , w_23647 );
and ( w_23646 ,  , w_23647 );
buf ( w_23645 , \9398_b1 );
not ( w_23645 , w_23648 );
not (  , w_23649 );
and ( w_23648 , w_23649 , \9398_b0 );
or ( \9400_b1 , \9399_b1 , w_23650 );
xor ( \9400_b0 , \9399_b0 , w_23652 );
not ( w_23652 , w_23653 );
and ( w_23653 , w_23650 , w_23651 );
buf ( w_23650 , \7181_b1 );
not ( w_23650 , w_23654 );
not ( w_23651 , w_23655 );
and ( w_23654 , w_23655 , \7181_b0 );
or ( \9401_b1 , \5893_b1 , \7192_b1 );
not ( \7192_b1 , w_23656 );
and ( \9401_b0 , \5893_b0 , w_23657 );
and ( w_23656 , w_23657 , \7192_b0 );
or ( \9402_b1 , \5861_b1 , \7190_b1 );
not ( \7190_b1 , w_23658 );
and ( \9402_b0 , \5861_b0 , w_23659 );
and ( w_23658 , w_23659 , \7190_b0 );
or ( \9403_b1 , \9401_b1 , w_23661 );
not ( w_23661 , w_23662 );
and ( \9403_b0 , \9401_b0 , w_23663 );
and ( w_23662 ,  , w_23663 );
buf ( w_23661 , \9402_b1 );
not ( w_23661 , w_23664 );
not (  , w_23665 );
and ( w_23664 , w_23665 , \9402_b0 );
or ( \9404_b1 , \9403_b1 , w_23666 );
xor ( \9404_b0 , \9403_b0 , w_23668 );
not ( w_23668 , w_23669 );
and ( w_23669 , w_23666 , w_23667 );
buf ( w_23666 , \7198_b1 );
not ( w_23666 , w_23670 );
not ( w_23667 , w_23671 );
and ( w_23670 , w_23671 , \7198_b0 );
or ( \9405_b1 , \9400_b1 , \9404_b1 );
xor ( \9405_b0 , \9400_b0 , w_23672 );
not ( w_23672 , w_23673 );
and ( w_23673 , \9404_b1 , \9404_b0 );
or ( \9406_b1 , \5918_b1 , \7203_b1 );
not ( \7203_b1 , w_23674 );
and ( \9406_b0 , \5918_b0 , w_23675 );
and ( w_23674 , w_23675 , \7203_b0 );
or ( \9407_b1 , \5881_b1 , \7201_b1 );
not ( \7201_b1 , w_23676 );
and ( \9407_b0 , \5881_b0 , w_23677 );
and ( w_23676 , w_23677 , \7201_b0 );
or ( \9408_b1 , \9406_b1 , w_23679 );
not ( w_23679 , w_23680 );
and ( \9408_b0 , \9406_b0 , w_23681 );
and ( w_23680 ,  , w_23681 );
buf ( w_23679 , \9407_b1 );
not ( w_23679 , w_23682 );
not (  , w_23683 );
and ( w_23682 , w_23683 , \9407_b0 );
or ( \9409_b1 , \9408_b1 , w_23684 );
xor ( \9409_b0 , \9408_b0 , w_23686 );
not ( w_23686 , w_23687 );
and ( w_23687 , w_23684 , w_23685 );
buf ( w_23684 , \6824_b1 );
not ( w_23684 , w_23688 );
not ( w_23685 , w_23689 );
and ( w_23688 , w_23689 , \6824_b0 );
or ( \9410_b1 , \9405_b1 , \9409_b1 );
xor ( \9410_b0 , \9405_b0 , w_23690 );
not ( w_23690 , w_23691 );
and ( w_23691 , \9409_b1 , \9409_b0 );
or ( \9411_b1 , \5811_b1 , \7117_b1 );
not ( \7117_b1 , w_23692 );
and ( \9411_b0 , \5811_b0 , w_23693 );
and ( w_23692 , w_23693 , \7117_b0 );
or ( \9412_b1 , \5780_b1 , \7115_b1 );
not ( \7115_b1 , w_23694 );
and ( \9412_b0 , \5780_b0 , w_23695 );
and ( w_23694 , w_23695 , \7115_b0 );
or ( \9413_b1 , \9411_b1 , w_23697 );
not ( w_23697 , w_23698 );
and ( \9413_b0 , \9411_b0 , w_23699 );
and ( w_23698 ,  , w_23699 );
buf ( w_23697 , \9412_b1 );
not ( w_23697 , w_23700 );
not (  , w_23701 );
and ( w_23700 , w_23701 , \9412_b0 );
or ( \9414_b1 , \9413_b1 , w_23702 );
xor ( \9414_b0 , \9413_b0 , w_23704 );
not ( w_23704 , w_23705 );
and ( w_23705 , w_23702 , w_23703 );
buf ( w_23702 , \7123_b1 );
not ( w_23702 , w_23706 );
not ( w_23703 , w_23707 );
and ( w_23706 , w_23707 , \7123_b0 );
or ( \9415_b1 , \5831_b1 , \7140_b1 );
not ( \7140_b1 , w_23708 );
and ( \9415_b0 , \5831_b0 , w_23709 );
and ( w_23708 , w_23709 , \7140_b0 );
or ( \9416_b1 , \5799_b1 , \7138_b1 );
not ( \7138_b1 , w_23710 );
and ( \9416_b0 , \5799_b0 , w_23711 );
and ( w_23710 , w_23711 , \7138_b0 );
or ( \9417_b1 , \9415_b1 , w_23713 );
not ( w_23713 , w_23714 );
and ( \9417_b0 , \9415_b0 , w_23715 );
and ( w_23714 ,  , w_23715 );
buf ( w_23713 , \9416_b1 );
not ( w_23713 , w_23716 );
not (  , w_23717 );
and ( w_23716 , w_23717 , \9416_b0 );
or ( \9418_b1 , \9417_b1 , w_23718 );
xor ( \9418_b0 , \9417_b0 , w_23720 );
not ( w_23720 , w_23721 );
and ( w_23721 , w_23718 , w_23719 );
buf ( w_23718 , \7146_b1 );
not ( w_23718 , w_23722 );
not ( w_23719 , w_23723 );
and ( w_23722 , w_23723 , \7146_b0 );
or ( \9419_b1 , \9414_b1 , \9418_b1 );
xor ( \9419_b0 , \9414_b0 , w_23724 );
not ( w_23724 , w_23725 );
and ( w_23725 , \9418_b1 , \9418_b0 );
or ( \9420_b1 , \5854_b1 , \7157_b1 );
not ( \7157_b1 , w_23726 );
and ( \9420_b0 , \5854_b0 , w_23727 );
and ( w_23726 , w_23727 , \7157_b0 );
or ( \9421_b1 , \5819_b1 , \7155_b1 );
not ( \7155_b1 , w_23728 );
and ( \9421_b0 , \5819_b0 , w_23729 );
and ( w_23728 , w_23729 , \7155_b0 );
or ( \9422_b1 , \9420_b1 , w_23731 );
not ( w_23731 , w_23732 );
and ( \9422_b0 , \9420_b0 , w_23733 );
and ( w_23732 ,  , w_23733 );
buf ( w_23731 , \9421_b1 );
not ( w_23731 , w_23734 );
not (  , w_23735 );
and ( w_23734 , w_23735 , \9421_b0 );
or ( \9423_b1 , \9422_b1 , w_23736 );
xor ( \9423_b0 , \9422_b0 , w_23738 );
not ( w_23738 , w_23739 );
and ( w_23739 , w_23736 , w_23737 );
buf ( w_23736 , \7163_b1 );
not ( w_23736 , w_23740 );
not ( w_23737 , w_23741 );
and ( w_23740 , w_23741 , \7163_b0 );
or ( \9424_b1 , \9419_b1 , \9423_b1 );
xor ( \9424_b0 , \9419_b0 , w_23742 );
not ( w_23742 , w_23743 );
and ( w_23743 , \9423_b1 , \9423_b0 );
or ( \9425_b1 , \9410_b1 , \9424_b1 );
xor ( \9425_b0 , \9410_b0 , w_23744 );
not ( w_23744 , w_23745 );
and ( w_23745 , \9424_b1 , \9424_b0 );
buf ( \9426_b1 , \7067_b1 );
not ( \9426_b1 , w_23746 );
not ( \9426_b0 , w_23747 );
and ( w_23746 , w_23747 , \7067_b0 );
or ( \9427_b1 , \5770_b1 , \7082_b1 );
not ( \7082_b1 , w_23748 );
and ( \9427_b0 , \5770_b0 , w_23749 );
and ( w_23748 , w_23749 , \7082_b0 );
or ( \9428_b1 , \5737_b1 , \7080_b1 );
not ( \7080_b1 , w_23750 );
and ( \9428_b0 , \5737_b0 , w_23751 );
and ( w_23750 , w_23751 , \7080_b0 );
or ( \9429_b1 , \9427_b1 , w_23753 );
not ( w_23753 , w_23754 );
and ( \9429_b0 , \9427_b0 , w_23755 );
and ( w_23754 ,  , w_23755 );
buf ( w_23753 , \9428_b1 );
not ( w_23753 , w_23756 );
not (  , w_23757 );
and ( w_23756 , w_23757 , \9428_b0 );
or ( \9430_b1 , \9429_b1 , w_23758 );
xor ( \9430_b0 , \9429_b0 , w_23760 );
not ( w_23760 , w_23761 );
and ( w_23761 , w_23758 , w_23759 );
buf ( w_23758 , \7088_b1 );
not ( w_23758 , w_23762 );
not ( w_23759 , w_23763 );
and ( w_23762 , w_23763 , \7088_b0 );
or ( \9431_b1 , \9426_b1 , \9430_b1 );
xor ( \9431_b0 , \9426_b0 , w_23764 );
not ( w_23764 , w_23765 );
and ( w_23765 , \9430_b1 , \9430_b0 );
or ( \9432_b1 , \5792_b1 , \7099_b1 );
not ( \7099_b1 , w_23766 );
and ( \9432_b0 , \5792_b0 , w_23767 );
and ( w_23766 , w_23767 , \7099_b0 );
or ( \9433_b1 , \5758_b1 , \7097_b1 );
not ( \7097_b1 , w_23768 );
and ( \9433_b0 , \5758_b0 , w_23769 );
and ( w_23768 , w_23769 , \7097_b0 );
or ( \9434_b1 , \9432_b1 , w_23771 );
not ( w_23771 , w_23772 );
and ( \9434_b0 , \9432_b0 , w_23773 );
and ( w_23772 ,  , w_23773 );
buf ( w_23771 , \9433_b1 );
not ( w_23771 , w_23774 );
not (  , w_23775 );
and ( w_23774 , w_23775 , \9433_b0 );
or ( \9435_b1 , \9434_b1 , w_23776 );
xor ( \9435_b0 , \9434_b0 , w_23778 );
not ( w_23778 , w_23779 );
and ( w_23779 , w_23776 , w_23777 );
buf ( w_23776 , \7105_b1 );
not ( w_23776 , w_23780 );
not ( w_23777 , w_23781 );
and ( w_23780 , w_23781 , \7105_b0 );
or ( \9436_b1 , \9431_b1 , \9435_b1 );
xor ( \9436_b0 , \9431_b0 , w_23782 );
not ( w_23782 , w_23783 );
and ( w_23783 , \9435_b1 , \9435_b0 );
or ( \9437_b1 , \9425_b1 , \9436_b1 );
xor ( \9437_b0 , \9425_b0 , w_23784 );
not ( w_23784 , w_23785 );
and ( w_23785 , \9436_b1 , \9436_b0 );
or ( \9438_b1 , \9396_b1 , \9437_b1 );
xor ( \9438_b0 , \9396_b0 , w_23786 );
not ( w_23786 , w_23787 );
and ( w_23787 , \9437_b1 , \9437_b0 );
or ( \9439_b1 , \6057_b1 , \5871_b1 );
not ( \5871_b1 , w_23788 );
and ( \9439_b0 , \6057_b0 , w_23789 );
and ( w_23788 , w_23789 , \5871_b0 );
or ( \9440_b1 , \6029_b1 , \5869_b1 );
not ( \5869_b1 , w_23790 );
and ( \9440_b0 , \6029_b0 , w_23791 );
and ( w_23790 , w_23791 , \5869_b0 );
or ( \9441_b1 , \9439_b1 , w_23793 );
not ( w_23793 , w_23794 );
and ( \9441_b0 , \9439_b0 , w_23795 );
and ( w_23794 ,  , w_23795 );
buf ( w_23793 , \9440_b1 );
not ( w_23793 , w_23796 );
not (  , w_23797 );
and ( w_23796 , w_23797 , \9440_b0 );
or ( \9442_b1 , \9441_b1 , w_23798 );
xor ( \9442_b0 , \9441_b0 , w_23800 );
not ( w_23800 , w_23801 );
and ( w_23801 , w_23798 , w_23799 );
buf ( w_23798 , \5878_b1 );
not ( w_23798 , w_23802 );
not ( w_23799 , w_23803 );
and ( w_23802 , w_23803 , \5878_b0 );
or ( \9443_b1 , \6065_b1 , \5891_b1 );
not ( \5891_b1 , w_23804 );
and ( \9443_b0 , \6065_b0 , w_23805 );
and ( w_23804 , w_23805 , \5891_b0 );
or ( \9444_b1 , \6048_b1 , \5889_b1 );
not ( \5889_b1 , w_23806 );
and ( \9444_b0 , \6048_b0 , w_23807 );
and ( w_23806 , w_23807 , \5889_b0 );
or ( \9445_b1 , \9443_b1 , w_23809 );
not ( w_23809 , w_23810 );
and ( \9445_b0 , \9443_b0 , w_23811 );
and ( w_23810 ,  , w_23811 );
buf ( w_23809 , \9444_b1 );
not ( w_23809 , w_23812 );
not (  , w_23813 );
and ( w_23812 , w_23813 , \9444_b0 );
or ( \9446_b1 , \9445_b1 , w_23814 );
xor ( \9446_b0 , \9445_b0 , w_23816 );
not ( w_23816 , w_23817 );
and ( w_23817 , w_23814 , w_23815 );
buf ( w_23814 , \5898_b1 );
not ( w_23814 , w_23818 );
not ( w_23815 , w_23819 );
and ( w_23818 , w_23819 , \5898_b0 );
or ( \9447_b1 , \9442_b1 , \9446_b1 );
xor ( \9447_b0 , \9442_b0 , w_23820 );
not ( w_23820 , w_23821 );
and ( w_23821 , \9446_b1 , \9446_b0 );
or ( \9448_b1 , \5998_b1 , \5809_b1 );
not ( \5809_b1 , w_23822 );
and ( \9448_b0 , \5998_b0 , w_23823 );
and ( w_23822 , w_23823 , \5809_b0 );
or ( \9449_b1 , \5967_b1 , \5807_b1 );
not ( \5807_b1 , w_23824 );
and ( \9449_b0 , \5967_b0 , w_23825 );
and ( w_23824 , w_23825 , \5807_b0 );
or ( \9450_b1 , \9448_b1 , w_23827 );
not ( w_23827 , w_23828 );
and ( \9450_b0 , \9448_b0 , w_23829 );
and ( w_23828 ,  , w_23829 );
buf ( w_23827 , \9449_b1 );
not ( w_23827 , w_23830 );
not (  , w_23831 );
and ( w_23830 , w_23831 , \9449_b0 );
or ( \9451_b1 , \9450_b1 , w_23832 );
xor ( \9451_b0 , \9450_b0 , w_23834 );
not ( w_23834 , w_23835 );
and ( w_23835 , w_23832 , w_23833 );
buf ( w_23832 , \5816_b1 );
not ( w_23832 , w_23836 );
not ( w_23833 , w_23837 );
and ( w_23836 , w_23837 , \5816_b0 );
or ( \9452_b1 , \6018_b1 , \5829_b1 );
not ( \5829_b1 , w_23838 );
and ( \9452_b0 , \6018_b0 , w_23839 );
and ( w_23838 , w_23839 , \5829_b0 );
or ( \9453_b1 , \5986_b1 , \5827_b1 );
not ( \5827_b1 , w_23840 );
and ( \9453_b0 , \5986_b0 , w_23841 );
and ( w_23840 , w_23841 , \5827_b0 );
or ( \9454_b1 , \9452_b1 , w_23843 );
not ( w_23843 , w_23844 );
and ( \9454_b0 , \9452_b0 , w_23845 );
and ( w_23844 ,  , w_23845 );
buf ( w_23843 , \9453_b1 );
not ( w_23843 , w_23846 );
not (  , w_23847 );
and ( w_23846 , w_23847 , \9453_b0 );
or ( \9455_b1 , \9454_b1 , w_23848 );
xor ( \9455_b0 , \9454_b0 , w_23850 );
not ( w_23850 , w_23851 );
and ( w_23851 , w_23848 , w_23849 );
buf ( w_23848 , \5836_b1 );
not ( w_23848 , w_23852 );
not ( w_23849 , w_23853 );
and ( w_23852 , w_23853 , \5836_b0 );
or ( \9456_b1 , \9451_b1 , \9455_b1 );
xor ( \9456_b0 , \9451_b0 , w_23854 );
not ( w_23854 , w_23855 );
and ( w_23855 , \9455_b1 , \9455_b0 );
or ( \9457_b1 , \6041_b1 , \5852_b1 );
not ( \5852_b1 , w_23856 );
and ( \9457_b0 , \6041_b0 , w_23857 );
and ( w_23856 , w_23857 , \5852_b0 );
or ( \9458_b1 , \6006_b1 , \5850_b1 );
not ( \5850_b1 , w_23858 );
and ( \9458_b0 , \6006_b0 , w_23859 );
and ( w_23858 , w_23859 , \5850_b0 );
or ( \9459_b1 , \9457_b1 , w_23861 );
not ( w_23861 , w_23862 );
and ( \9459_b0 , \9457_b0 , w_23863 );
and ( w_23862 ,  , w_23863 );
buf ( w_23861 , \9458_b1 );
not ( w_23861 , w_23864 );
not (  , w_23865 );
and ( w_23864 , w_23865 , \9458_b0 );
or ( \9460_b1 , \9459_b1 , w_23866 );
xor ( \9460_b0 , \9459_b0 , w_23868 );
not ( w_23868 , w_23869 );
and ( w_23869 , w_23866 , w_23867 );
buf ( w_23866 , \5859_b1 );
not ( w_23866 , w_23870 );
not ( w_23867 , w_23871 );
and ( w_23870 , w_23871 , \5859_b0 );
or ( \9461_b1 , \9456_b1 , \9460_b1 );
xor ( \9461_b0 , \9456_b0 , w_23872 );
not ( w_23872 , w_23873 );
and ( w_23873 , \9460_b1 , \9460_b0 );
or ( \9462_b1 , \9447_b1 , \9461_b1 );
xor ( \9462_b0 , \9447_b0 , w_23874 );
not ( w_23874 , w_23875 );
and ( w_23875 , \9461_b1 , \9461_b0 );
or ( \9463_b1 , \5937_b1 , \5750_b1 );
not ( \5750_b1 , w_23876 );
and ( \9463_b0 , \5937_b0 , w_23877 );
and ( w_23876 , w_23877 , \5750_b0 );
or ( \9464_b1 , \5906_b1 , \5748_b1 );
not ( \5748_b1 , w_23878 );
and ( \9464_b0 , \5906_b0 , w_23879 );
and ( w_23878 , w_23879 , \5748_b0 );
or ( \9465_b1 , \9463_b1 , w_23881 );
not ( w_23881 , w_23882 );
and ( \9465_b0 , \9463_b0 , w_23883 );
and ( w_23882 ,  , w_23883 );
buf ( w_23881 , \9464_b1 );
not ( w_23881 , w_23884 );
not (  , w_23885 );
and ( w_23884 , w_23885 , \9464_b0 );
or ( \9466_b1 , \9465_b1 , w_23886 );
xor ( \9466_b0 , \9465_b0 , w_23888 );
not ( w_23888 , w_23889 );
and ( w_23889 , w_23886 , w_23887 );
buf ( w_23886 , \5755_b1 );
not ( w_23886 , w_23890 );
not ( w_23887 , w_23891 );
and ( w_23890 , w_23891 , \5755_b0 );
or ( \9467_b1 , \5957_b1 , \5768_b1 );
not ( \5768_b1 , w_23892 );
and ( \9467_b0 , \5957_b0 , w_23893 );
and ( w_23892 , w_23893 , \5768_b0 );
or ( \9468_b1 , \5925_b1 , \5766_b1 );
not ( \5766_b1 , w_23894 );
and ( \9468_b0 , \5925_b0 , w_23895 );
and ( w_23894 , w_23895 , \5766_b0 );
or ( \9469_b1 , \9467_b1 , w_23897 );
not ( w_23897 , w_23898 );
and ( \9469_b0 , \9467_b0 , w_23899 );
and ( w_23898 ,  , w_23899 );
buf ( w_23897 , \9468_b1 );
not ( w_23897 , w_23900 );
not (  , w_23901 );
and ( w_23900 , w_23901 , \9468_b0 );
or ( \9470_b1 , \9469_b1 , w_23902 );
xor ( \9470_b0 , \9469_b0 , w_23904 );
not ( w_23904 , w_23905 );
and ( w_23905 , w_23902 , w_23903 );
buf ( w_23902 , \5775_b1 );
not ( w_23902 , w_23906 );
not ( w_23903 , w_23907 );
and ( w_23906 , w_23907 , \5775_b0 );
or ( \9471_b1 , \9466_b1 , \9470_b1 );
xor ( \9471_b0 , \9466_b0 , w_23908 );
not ( w_23908 , w_23909 );
and ( w_23909 , \9470_b1 , \9470_b0 );
or ( \9472_b1 , \5979_b1 , \5790_b1 );
not ( \5790_b1 , w_23910 );
and ( \9472_b0 , \5979_b0 , w_23911 );
and ( w_23910 , w_23911 , \5790_b0 );
or ( \9473_b1 , \5945_b1 , \5788_b1 );
not ( \5788_b1 , w_23912 );
and ( \9473_b0 , \5945_b0 , w_23913 );
and ( w_23912 , w_23913 , \5788_b0 );
or ( \9474_b1 , \9472_b1 , w_23915 );
not ( w_23915 , w_23916 );
and ( \9474_b0 , \9472_b0 , w_23917 );
and ( w_23916 ,  , w_23917 );
buf ( w_23915 , \9473_b1 );
not ( w_23915 , w_23918 );
not (  , w_23919 );
and ( w_23918 , w_23919 , \9473_b0 );
or ( \9475_b1 , \9474_b1 , w_23920 );
xor ( \9475_b0 , \9474_b0 , w_23922 );
not ( w_23922 , w_23923 );
and ( w_23923 , w_23920 , w_23921 );
buf ( w_23920 , \5797_b1 );
not ( w_23920 , w_23924 );
not ( w_23921 , w_23925 );
and ( w_23924 , w_23925 , \5797_b0 );
or ( \9476_b1 , \9471_b1 , \9475_b1 );
xor ( \9476_b0 , \9471_b0 , w_23926 );
not ( w_23926 , w_23927 );
and ( w_23927 , \9475_b1 , \9475_b0 );
or ( \9477_b1 , \9462_b1 , \9476_b1 );
xor ( \9477_b0 , \9462_b0 , w_23928 );
not ( w_23928 , w_23929 );
and ( w_23929 , \9476_b1 , \9476_b0 );
or ( \9478_b1 , \9438_b1 , \9477_b1 );
xor ( \9478_b0 , \9438_b0 , w_23930 );
not ( w_23930 , w_23931 );
and ( w_23931 , \9477_b1 , \9477_b0 );
or ( \9479_b1 , \9392_b1 , \9478_b1 );
xor ( \9479_b0 , \9392_b0 , w_23932 );
not ( w_23932 , w_23933 );
and ( w_23933 , \9478_b1 , \9478_b0 );
or ( \9480_b1 , \9241_b1 , \9245_b1 );
not ( \9245_b1 , w_23934 );
and ( \9480_b0 , \9241_b0 , w_23935 );
and ( w_23934 , w_23935 , \9245_b0 );
or ( \9481_b1 , \9245_b1 , \9250_b1 );
not ( \9250_b1 , w_23936 );
and ( \9481_b0 , \9245_b0 , w_23937 );
and ( w_23936 , w_23937 , \9250_b0 );
or ( \9482_b1 , \9241_b1 , \9250_b1 );
not ( \9250_b1 , w_23938 );
and ( \9482_b0 , \9241_b0 , w_23939 );
and ( w_23938 , w_23939 , \9250_b0 );
or ( \9484_b1 , \9229_b1 , \9233_b1 );
not ( \9233_b1 , w_23940 );
and ( \9484_b0 , \9229_b0 , w_23941 );
and ( w_23940 , w_23941 , \9233_b0 );
or ( \9485_b1 , \9233_b1 , \9235_b1 );
not ( \9235_b1 , w_23942 );
and ( \9485_b0 , \9233_b0 , w_23943 );
and ( w_23942 , w_23943 , \9235_b0 );
or ( \9486_b1 , \9229_b1 , \9235_b1 );
not ( \9235_b1 , w_23944 );
and ( \9486_b0 , \9229_b0 , w_23945 );
and ( w_23944 , w_23945 , \9235_b0 );
or ( \9488_b1 , \9483_b1 , \9487_b1 );
xor ( \9488_b0 , \9483_b0 , w_23946 );
not ( w_23946 , w_23947 );
and ( w_23947 , \9487_b1 , \9487_b0 );
or ( \9489_b1 , \9210_b1 , w_23948 );
or ( \9489_b0 , \9210_b0 , \9224_b0 );
not ( \9224_b0 , w_23949 );
and ( w_23949 , w_23948 , \9224_b1 );
or ( \9490_b1 , \9488_b1 , \9489_b1 );
xor ( \9490_b0 , \9488_b0 , w_23950 );
not ( w_23950 , w_23951 );
and ( w_23951 , \9489_b1 , \9489_b0 );
or ( \9491_b1 , \9479_b1 , \9490_b1 );
xor ( \9491_b0 , \9479_b0 , w_23952 );
not ( w_23952 , w_23953 );
and ( w_23953 , \9490_b1 , \9490_b0 );
or ( \9492_b1 , \9363_b1 , \9491_b1 );
xor ( \9492_b0 , \9363_b0 , w_23954 );
not ( w_23954 , w_23955 );
and ( w_23955 , \9491_b1 , \9491_b0 );
or ( \9493_b1 , \9354_b1 , \9492_b1 );
xor ( \9493_b0 , \9354_b0 , w_23956 );
not ( w_23956 , w_23957 );
and ( w_23957 , \9492_b1 , \9492_b0 );
or ( \9494_b1 , \9177_b1 , \9188_b1 );
not ( \9188_b1 , w_23958 );
and ( \9494_b0 , \9177_b0 , w_23959 );
and ( w_23958 , w_23959 , \9188_b0 );
or ( \9495_b1 , \9188_b1 , \9328_b1 );
not ( \9328_b1 , w_23960 );
and ( \9495_b0 , \9188_b0 , w_23961 );
and ( w_23960 , w_23961 , \9328_b0 );
or ( \9496_b1 , \9177_b1 , \9328_b1 );
not ( \9328_b1 , w_23962 );
and ( \9496_b0 , \9177_b0 , w_23963 );
and ( w_23962 , w_23963 , \9328_b0 );
or ( \9498_b1 , \9493_b1 , w_23965 );
not ( w_23965 , w_23966 );
and ( \9498_b0 , \9493_b0 , w_23967 );
and ( w_23966 ,  , w_23967 );
buf ( w_23965 , \9497_b1 );
not ( w_23965 , w_23968 );
not (  , w_23969 );
and ( w_23968 , w_23969 , \9497_b0 );
or ( \9499_b1 , \9358_b1 , \9362_b1 );
not ( \9362_b1 , w_23970 );
and ( \9499_b0 , \9358_b0 , w_23971 );
and ( w_23970 , w_23971 , \9362_b0 );
or ( \9500_b1 , \9362_b1 , \9491_b1 );
not ( \9491_b1 , w_23972 );
and ( \9500_b0 , \9362_b0 , w_23973 );
and ( w_23972 , w_23973 , \9491_b0 );
or ( \9501_b1 , \9358_b1 , \9491_b1 );
not ( \9491_b1 , w_23974 );
and ( \9501_b0 , \9358_b0 , w_23975 );
and ( w_23974 , w_23975 , \9491_b0 );
or ( \9503_b1 , \9483_b1 , \9487_b1 );
not ( \9487_b1 , w_23976 );
and ( \9503_b0 , \9483_b0 , w_23977 );
and ( w_23976 , w_23977 , \9487_b0 );
or ( \9504_b1 , \9487_b1 , \9489_b1 );
not ( \9489_b1 , w_23978 );
and ( \9504_b0 , \9487_b0 , w_23979 );
and ( w_23978 , w_23979 , \9489_b0 );
or ( \9505_b1 , \9483_b1 , \9489_b1 );
not ( \9489_b1 , w_23980 );
and ( \9505_b0 , \9483_b0 , w_23981 );
and ( w_23980 , w_23981 , \9489_b0 );
or ( \9507_b1 , \9396_b1 , \9437_b1 );
not ( \9437_b1 , w_23982 );
and ( \9507_b0 , \9396_b0 , w_23983 );
and ( w_23982 , w_23983 , \9437_b0 );
or ( \9508_b1 , \9437_b1 , \9477_b1 );
not ( \9477_b1 , w_23984 );
and ( \9508_b0 , \9437_b0 , w_23985 );
and ( w_23984 , w_23985 , \9477_b0 );
or ( \9509_b1 , \9396_b1 , \9477_b1 );
not ( \9477_b1 , w_23986 );
and ( \9509_b0 , \9396_b0 , w_23987 );
and ( w_23986 , w_23987 , \9477_b0 );
or ( \9511_b1 , \9506_b1 , \9510_b1 );
xor ( \9511_b0 , \9506_b0 , w_23988 );
not ( w_23988 , w_23989 );
and ( w_23989 , \9510_b1 , \9510_b0 );
or ( \9512_b1 , \9377_b1 , \9391_b1 );
not ( \9391_b1 , w_23990 );
and ( \9512_b0 , \9377_b0 , w_23991 );
and ( w_23990 , w_23991 , \9391_b0 );
or ( \9513_b1 , \9511_b1 , \9512_b1 );
xor ( \9513_b0 , \9511_b0 , w_23992 );
not ( w_23992 , w_23993 );
and ( w_23993 , \9512_b1 , \9512_b0 );
or ( \9514_b1 , \9502_b1 , \9513_b1 );
xor ( \9514_b0 , \9502_b0 , w_23994 );
not ( w_23994 , w_23995 );
and ( w_23995 , \9513_b1 , \9513_b0 );
or ( \9515_b1 , \9343_b1 , \9347_b1 );
not ( \9347_b1 , w_23996 );
and ( \9515_b0 , \9343_b0 , w_23997 );
and ( w_23996 , w_23997 , \9347_b0 );
or ( \9516_b1 , \9347_b1 , \9352_b1 );
not ( \9352_b1 , w_23998 );
and ( \9516_b0 , \9347_b0 , w_23999 );
and ( w_23998 , w_23999 , \9352_b0 );
or ( \9517_b1 , \9343_b1 , \9352_b1 );
not ( \9352_b1 , w_24000 );
and ( \9517_b0 , \9343_b0 , w_24001 );
and ( w_24000 , w_24001 , \9352_b0 );
or ( \9519_b1 , \9392_b1 , \9478_b1 );
not ( \9478_b1 , w_24002 );
and ( \9519_b0 , \9392_b0 , w_24003 );
and ( w_24002 , w_24003 , \9478_b0 );
or ( \9520_b1 , \9478_b1 , \9490_b1 );
not ( \9490_b1 , w_24004 );
and ( \9520_b0 , \9478_b0 , w_24005 );
and ( w_24004 , w_24005 , \9490_b0 );
or ( \9521_b1 , \9392_b1 , \9490_b1 );
not ( \9490_b1 , w_24006 );
and ( \9521_b0 , \9392_b0 , w_24007 );
and ( w_24006 , w_24007 , \9490_b0 );
or ( \9523_b1 , \9518_b1 , \9522_b1 );
xor ( \9523_b0 , \9518_b0 , w_24008 );
not ( w_24008 , w_24009 );
and ( w_24009 , \9522_b1 , \9522_b0 );
or ( \9524_b1 , \6029_b1 , \5871_b1 );
not ( \5871_b1 , w_24010 );
and ( \9524_b0 , \6029_b0 , w_24011 );
and ( w_24010 , w_24011 , \5871_b0 );
or ( \9525_b1 , \6041_b1 , \5869_b1 );
not ( \5869_b1 , w_24012 );
and ( \9525_b0 , \6041_b0 , w_24013 );
and ( w_24012 , w_24013 , \5869_b0 );
or ( \9526_b1 , \9524_b1 , w_24015 );
not ( w_24015 , w_24016 );
and ( \9526_b0 , \9524_b0 , w_24017 );
and ( w_24016 ,  , w_24017 );
buf ( w_24015 , \9525_b1 );
not ( w_24015 , w_24018 );
not (  , w_24019 );
and ( w_24018 , w_24019 , \9525_b0 );
or ( \9527_b1 , \9526_b1 , w_24020 );
xor ( \9527_b0 , \9526_b0 , w_24022 );
not ( w_24022 , w_24023 );
and ( w_24023 , w_24020 , w_24021 );
buf ( w_24020 , \5878_b1 );
not ( w_24020 , w_24024 );
not ( w_24021 , w_24025 );
and ( w_24024 , w_24025 , \5878_b0 );
or ( \9528_b1 , \6048_b1 , \5891_b1 );
not ( \5891_b1 , w_24026 );
and ( \9528_b0 , \6048_b0 , w_24027 );
and ( w_24026 , w_24027 , \5891_b0 );
or ( \9529_b1 , \6057_b1 , \5889_b1 );
not ( \5889_b1 , w_24028 );
and ( \9529_b0 , \6057_b0 , w_24029 );
and ( w_24028 , w_24029 , \5889_b0 );
or ( \9530_b1 , \9528_b1 , w_24031 );
not ( w_24031 , w_24032 );
and ( \9530_b0 , \9528_b0 , w_24033 );
and ( w_24032 ,  , w_24033 );
buf ( w_24031 , \9529_b1 );
not ( w_24031 , w_24034 );
not (  , w_24035 );
and ( w_24034 , w_24035 , \9529_b0 );
or ( \9531_b1 , \9530_b1 , w_24036 );
xor ( \9531_b0 , \9530_b0 , w_24038 );
not ( w_24038 , w_24039 );
and ( w_24039 , w_24036 , w_24037 );
buf ( w_24036 , \5898_b1 );
not ( w_24036 , w_24040 );
not ( w_24037 , w_24041 );
and ( w_24040 , w_24041 , \5898_b0 );
or ( \9532_b1 , \9527_b1 , \9531_b1 );
xor ( \9532_b0 , \9527_b0 , w_24042 );
not ( w_24042 , w_24043 );
and ( w_24043 , \9531_b1 , \9531_b0 );
or ( \9533_b1 , \6065_b1 , w_24045 );
not ( w_24045 , w_24046 );
and ( \9533_b0 , \6065_b0 , w_24047 );
and ( w_24046 ,  , w_24047 );
buf ( w_24045 , \5914_b1 );
not ( w_24045 , w_24048 );
not (  , w_24049 );
and ( w_24048 , w_24049 , \5914_b0 );
or ( \9534_b1 , \9533_b1 , w_24050 );
xor ( \9534_b0 , \9533_b0 , w_24052 );
not ( w_24052 , w_24053 );
and ( w_24053 , w_24050 , w_24051 );
buf ( w_24050 , \5923_b1 );
not ( w_24050 , w_24054 );
not ( w_24051 , w_24055 );
and ( w_24054 , w_24055 , \5923_b0 );
or ( \9535_b1 , \9532_b1 , \9534_b1 );
xor ( \9535_b0 , \9532_b0 , w_24056 );
not ( w_24056 , w_24057 );
and ( w_24057 , \9534_b1 , \9534_b0 );
or ( \9536_b1 , \5967_b1 , \5809_b1 );
not ( \5809_b1 , w_24058 );
and ( \9536_b0 , \5967_b0 , w_24059 );
and ( w_24058 , w_24059 , \5809_b0 );
or ( \9537_b1 , \5979_b1 , \5807_b1 );
not ( \5807_b1 , w_24060 );
and ( \9537_b0 , \5979_b0 , w_24061 );
and ( w_24060 , w_24061 , \5807_b0 );
or ( \9538_b1 , \9536_b1 , w_24063 );
not ( w_24063 , w_24064 );
and ( \9538_b0 , \9536_b0 , w_24065 );
and ( w_24064 ,  , w_24065 );
buf ( w_24063 , \9537_b1 );
not ( w_24063 , w_24066 );
not (  , w_24067 );
and ( w_24066 , w_24067 , \9537_b0 );
or ( \9539_b1 , \9538_b1 , w_24068 );
xor ( \9539_b0 , \9538_b0 , w_24070 );
not ( w_24070 , w_24071 );
and ( w_24071 , w_24068 , w_24069 );
buf ( w_24068 , \5816_b1 );
not ( w_24068 , w_24072 );
not ( w_24069 , w_24073 );
and ( w_24072 , w_24073 , \5816_b0 );
or ( \9540_b1 , \5986_b1 , \5829_b1 );
not ( \5829_b1 , w_24074 );
and ( \9540_b0 , \5986_b0 , w_24075 );
and ( w_24074 , w_24075 , \5829_b0 );
or ( \9541_b1 , \5998_b1 , \5827_b1 );
not ( \5827_b1 , w_24076 );
and ( \9541_b0 , \5998_b0 , w_24077 );
and ( w_24076 , w_24077 , \5827_b0 );
or ( \9542_b1 , \9540_b1 , w_24079 );
not ( w_24079 , w_24080 );
and ( \9542_b0 , \9540_b0 , w_24081 );
and ( w_24080 ,  , w_24081 );
buf ( w_24079 , \9541_b1 );
not ( w_24079 , w_24082 );
not (  , w_24083 );
and ( w_24082 , w_24083 , \9541_b0 );
or ( \9543_b1 , \9542_b1 , w_24084 );
xor ( \9543_b0 , \9542_b0 , w_24086 );
not ( w_24086 , w_24087 );
and ( w_24087 , w_24084 , w_24085 );
buf ( w_24084 , \5836_b1 );
not ( w_24084 , w_24088 );
not ( w_24085 , w_24089 );
and ( w_24088 , w_24089 , \5836_b0 );
or ( \9544_b1 , \9539_b1 , \9543_b1 );
xor ( \9544_b0 , \9539_b0 , w_24090 );
not ( w_24090 , w_24091 );
and ( w_24091 , \9543_b1 , \9543_b0 );
or ( \9545_b1 , \6006_b1 , \5852_b1 );
not ( \5852_b1 , w_24092 );
and ( \9545_b0 , \6006_b0 , w_24093 );
and ( w_24092 , w_24093 , \5852_b0 );
or ( \9546_b1 , \6018_b1 , \5850_b1 );
not ( \5850_b1 , w_24094 );
and ( \9546_b0 , \6018_b0 , w_24095 );
and ( w_24094 , w_24095 , \5850_b0 );
or ( \9547_b1 , \9545_b1 , w_24097 );
not ( w_24097 , w_24098 );
and ( \9547_b0 , \9545_b0 , w_24099 );
and ( w_24098 ,  , w_24099 );
buf ( w_24097 , \9546_b1 );
not ( w_24097 , w_24100 );
not (  , w_24101 );
and ( w_24100 , w_24101 , \9546_b0 );
or ( \9548_b1 , \9547_b1 , w_24102 );
xor ( \9548_b0 , \9547_b0 , w_24104 );
not ( w_24104 , w_24105 );
and ( w_24105 , w_24102 , w_24103 );
buf ( w_24102 , \5859_b1 );
not ( w_24102 , w_24106 );
not ( w_24103 , w_24107 );
and ( w_24106 , w_24107 , \5859_b0 );
or ( \9549_b1 , \9544_b1 , \9548_b1 );
xor ( \9549_b0 , \9544_b0 , w_24108 );
not ( w_24108 , w_24109 );
and ( w_24109 , \9548_b1 , \9548_b0 );
or ( \9550_b1 , \9535_b1 , w_24110 );
xor ( \9550_b0 , \9535_b0 , w_24112 );
not ( w_24112 , w_24113 );
and ( w_24113 , w_24110 , w_24111 );
buf ( w_24110 , \9549_b1 );
not ( w_24110 , w_24114 );
not ( w_24111 , w_24115 );
and ( w_24114 , w_24115 , \9549_b0 );
or ( \9551_b1 , \9466_b1 , \9470_b1 );
not ( \9470_b1 , w_24116 );
and ( \9551_b0 , \9466_b0 , w_24117 );
and ( w_24116 , w_24117 , \9470_b0 );
or ( \9552_b1 , \9470_b1 , \9475_b1 );
not ( \9475_b1 , w_24118 );
and ( \9552_b0 , \9470_b0 , w_24119 );
and ( w_24118 , w_24119 , \9475_b0 );
or ( \9553_b1 , \9466_b1 , \9475_b1 );
not ( \9475_b1 , w_24120 );
and ( \9553_b0 , \9466_b0 , w_24121 );
and ( w_24120 , w_24121 , \9475_b0 );
or ( \9555_b1 , \9451_b1 , \9455_b1 );
not ( \9455_b1 , w_24122 );
and ( \9555_b0 , \9451_b0 , w_24123 );
and ( w_24122 , w_24123 , \9455_b0 );
or ( \9556_b1 , \9455_b1 , \9460_b1 );
not ( \9460_b1 , w_24124 );
and ( \9556_b0 , \9455_b0 , w_24125 );
and ( w_24124 , w_24125 , \9460_b0 );
or ( \9557_b1 , \9451_b1 , \9460_b1 );
not ( \9460_b1 , w_24126 );
and ( \9557_b0 , \9451_b0 , w_24127 );
and ( w_24126 , w_24127 , \9460_b0 );
or ( \9559_b1 , \9554_b1 , \9558_b1 );
xor ( \9559_b0 , \9554_b0 , w_24128 );
not ( w_24128 , w_24129 );
and ( w_24129 , \9558_b1 , \9558_b0 );
or ( \9560_b1 , \9442_b1 , \9446_b1 );
not ( \9446_b1 , w_24130 );
and ( \9560_b0 , \9442_b0 , w_24131 );
and ( w_24130 , w_24131 , \9446_b0 );
or ( \9561_b1 , \9559_b1 , \9560_b1 );
xor ( \9561_b0 , \9559_b0 , w_24132 );
not ( w_24132 , w_24133 );
and ( w_24133 , \9560_b1 , \9560_b0 );
or ( \9562_b1 , \9550_b1 , \9561_b1 );
xor ( \9562_b0 , \9550_b0 , w_24134 );
not ( w_24134 , w_24135 );
and ( w_24135 , \9561_b1 , \9561_b0 );
or ( \9563_b1 , \9426_b1 , \9430_b1 );
not ( \9430_b1 , w_24136 );
and ( \9563_b0 , \9426_b0 , w_24137 );
and ( w_24136 , w_24137 , \9430_b0 );
or ( \9564_b1 , \9430_b1 , \9435_b1 );
not ( \9435_b1 , w_24138 );
and ( \9564_b0 , \9430_b0 , w_24139 );
and ( w_24138 , w_24139 , \9435_b0 );
or ( \9565_b1 , \9426_b1 , \9435_b1 );
not ( \9435_b1 , w_24140 );
and ( \9565_b0 , \9426_b0 , w_24141 );
and ( w_24140 , w_24141 , \9435_b0 );
or ( \9567_b1 , \9414_b1 , \9418_b1 );
not ( \9418_b1 , w_24142 );
and ( \9567_b0 , \9414_b0 , w_24143 );
and ( w_24142 , w_24143 , \9418_b0 );
or ( \9568_b1 , \9418_b1 , \9423_b1 );
not ( \9423_b1 , w_24144 );
and ( \9568_b0 , \9418_b0 , w_24145 );
and ( w_24144 , w_24145 , \9423_b0 );
or ( \9569_b1 , \9414_b1 , \9423_b1 );
not ( \9423_b1 , w_24146 );
and ( \9569_b0 , \9414_b0 , w_24147 );
and ( w_24146 , w_24147 , \9423_b0 );
or ( \9571_b1 , \9566_b1 , \9570_b1 );
xor ( \9571_b0 , \9566_b0 , w_24148 );
not ( w_24148 , w_24149 );
and ( w_24149 , \9570_b1 , \9570_b0 );
or ( \9572_b1 , \9400_b1 , \9404_b1 );
not ( \9404_b1 , w_24150 );
and ( \9572_b0 , \9400_b0 , w_24151 );
and ( w_24150 , w_24151 , \9404_b0 );
or ( \9573_b1 , \9404_b1 , \9409_b1 );
not ( \9409_b1 , w_24152 );
and ( \9573_b0 , \9404_b0 , w_24153 );
and ( w_24152 , w_24153 , \9409_b0 );
or ( \9574_b1 , \9400_b1 , \9409_b1 );
not ( \9409_b1 , w_24154 );
and ( \9574_b0 , \9400_b0 , w_24155 );
and ( w_24154 , w_24155 , \9409_b0 );
or ( \9576_b1 , \9571_b1 , \9575_b1 );
xor ( \9576_b0 , \9571_b0 , w_24156 );
not ( w_24156 , w_24157 );
and ( w_24157 , \9575_b1 , \9575_b0 );
or ( \9577_b1 , \9562_b1 , \9576_b1 );
xor ( \9577_b0 , \9562_b0 , w_24158 );
not ( w_24158 , w_24159 );
and ( w_24159 , \9576_b1 , \9576_b0 );
or ( \9578_b1 , \9410_b1 , \9424_b1 );
not ( \9424_b1 , w_24160 );
and ( \9578_b0 , \9410_b0 , w_24161 );
and ( w_24160 , w_24161 , \9424_b0 );
or ( \9579_b1 , \9424_b1 , \9436_b1 );
not ( \9436_b1 , w_24162 );
and ( \9579_b0 , \9424_b0 , w_24163 );
and ( w_24162 , w_24163 , \9436_b0 );
or ( \9580_b1 , \9410_b1 , \9436_b1 );
not ( \9436_b1 , w_24164 );
and ( \9580_b0 , \9410_b0 , w_24165 );
and ( w_24164 , w_24165 , \9436_b0 );
or ( \9582_b1 , \5737_b1 , \7082_b1 );
not ( \7082_b1 , w_24166 );
and ( \9582_b0 , \5737_b0 , w_24167 );
and ( w_24166 , w_24167 , \7082_b0 );
buf ( \9583_b1 , \9582_b1 );
not ( \9583_b1 , w_24168 );
not ( \9583_b0 , w_24169 );
and ( w_24168 , w_24169 , \9582_b0 );
or ( \9584_b1 , \9583_b1 , w_24170 );
xor ( \9584_b0 , \9583_b0 , w_24172 );
not ( w_24172 , w_24173 );
and ( w_24173 , w_24170 , w_24171 );
buf ( w_24170 , \7088_b1 );
not ( w_24170 , w_24174 );
not ( w_24171 , w_24175 );
and ( w_24174 , w_24175 , \7088_b0 );
or ( \9585_b1 , \5923_b1 , \9584_b1 );
xor ( \9585_b0 , \5923_b0 , w_24176 );
not ( w_24176 , w_24177 );
and ( w_24177 , \9584_b1 , \9584_b0 );
or ( \9586_b1 , \5758_b1 , \7099_b1 );
not ( \7099_b1 , w_24178 );
and ( \9586_b0 , \5758_b0 , w_24179 );
and ( w_24178 , w_24179 , \7099_b0 );
or ( \9587_b1 , \5770_b1 , \7097_b1 );
not ( \7097_b1 , w_24180 );
and ( \9587_b0 , \5770_b0 , w_24181 );
and ( w_24180 , w_24181 , \7097_b0 );
or ( \9588_b1 , \9586_b1 , w_24183 );
not ( w_24183 , w_24184 );
and ( \9588_b0 , \9586_b0 , w_24185 );
and ( w_24184 ,  , w_24185 );
buf ( w_24183 , \9587_b1 );
not ( w_24183 , w_24186 );
not (  , w_24187 );
and ( w_24186 , w_24187 , \9587_b0 );
or ( \9589_b1 , \9588_b1 , w_24188 );
xor ( \9589_b0 , \9588_b0 , w_24190 );
not ( w_24190 , w_24191 );
and ( w_24191 , w_24188 , w_24189 );
buf ( w_24188 , \7105_b1 );
not ( w_24188 , w_24192 );
not ( w_24189 , w_24193 );
and ( w_24192 , w_24193 , \7105_b0 );
or ( \9590_b1 , \9585_b1 , \9589_b1 );
xor ( \9590_b0 , \9585_b0 , w_24194 );
not ( w_24194 , w_24195 );
and ( w_24195 , \9589_b1 , \9589_b0 );
or ( \9591_b1 , \9581_b1 , \9590_b1 );
xor ( \9591_b0 , \9581_b0 , w_24196 );
not ( w_24196 , w_24197 );
and ( w_24197 , \9590_b1 , \9590_b0 );
or ( \9592_b1 , \5906_b1 , \5750_b1 );
not ( \5750_b1 , w_24198 );
and ( \9592_b0 , \5906_b0 , w_24199 );
and ( w_24198 , w_24199 , \5750_b0 );
or ( \9593_b1 , \5918_b1 , \5748_b1 );
not ( \5748_b1 , w_24200 );
and ( \9593_b0 , \5918_b0 , w_24201 );
and ( w_24200 , w_24201 , \5748_b0 );
or ( \9594_b1 , \9592_b1 , w_24203 );
not ( w_24203 , w_24204 );
and ( \9594_b0 , \9592_b0 , w_24205 );
and ( w_24204 ,  , w_24205 );
buf ( w_24203 , \9593_b1 );
not ( w_24203 , w_24206 );
not (  , w_24207 );
and ( w_24206 , w_24207 , \9593_b0 );
or ( \9595_b1 , \9594_b1 , w_24208 );
xor ( \9595_b0 , \9594_b0 , w_24210 );
not ( w_24210 , w_24211 );
and ( w_24211 , w_24208 , w_24209 );
buf ( w_24208 , \5755_b1 );
not ( w_24208 , w_24212 );
not ( w_24209 , w_24213 );
and ( w_24212 , w_24213 , \5755_b0 );
or ( \9596_b1 , \5925_b1 , \5768_b1 );
not ( \5768_b1 , w_24214 );
and ( \9596_b0 , \5925_b0 , w_24215 );
and ( w_24214 , w_24215 , \5768_b0 );
or ( \9597_b1 , \5937_b1 , \5766_b1 );
not ( \5766_b1 , w_24216 );
and ( \9597_b0 , \5937_b0 , w_24217 );
and ( w_24216 , w_24217 , \5766_b0 );
or ( \9598_b1 , \9596_b1 , w_24219 );
not ( w_24219 , w_24220 );
and ( \9598_b0 , \9596_b0 , w_24221 );
and ( w_24220 ,  , w_24221 );
buf ( w_24219 , \9597_b1 );
not ( w_24219 , w_24222 );
not (  , w_24223 );
and ( w_24222 , w_24223 , \9597_b0 );
or ( \9599_b1 , \9598_b1 , w_24224 );
xor ( \9599_b0 , \9598_b0 , w_24226 );
not ( w_24226 , w_24227 );
and ( w_24227 , w_24224 , w_24225 );
buf ( w_24224 , \5775_b1 );
not ( w_24224 , w_24228 );
not ( w_24225 , w_24229 );
and ( w_24228 , w_24229 , \5775_b0 );
or ( \9600_b1 , \9595_b1 , \9599_b1 );
xor ( \9600_b0 , \9595_b0 , w_24230 );
not ( w_24230 , w_24231 );
and ( w_24231 , \9599_b1 , \9599_b0 );
or ( \9601_b1 , \5945_b1 , \5790_b1 );
not ( \5790_b1 , w_24232 );
and ( \9601_b0 , \5945_b0 , w_24233 );
and ( w_24232 , w_24233 , \5790_b0 );
or ( \9602_b1 , \5957_b1 , \5788_b1 );
not ( \5788_b1 , w_24234 );
and ( \9602_b0 , \5957_b0 , w_24235 );
and ( w_24234 , w_24235 , \5788_b0 );
or ( \9603_b1 , \9601_b1 , w_24237 );
not ( w_24237 , w_24238 );
and ( \9603_b0 , \9601_b0 , w_24239 );
and ( w_24238 ,  , w_24239 );
buf ( w_24237 , \9602_b1 );
not ( w_24237 , w_24240 );
not (  , w_24241 );
and ( w_24240 , w_24241 , \9602_b0 );
or ( \9604_b1 , \9603_b1 , w_24242 );
xor ( \9604_b0 , \9603_b0 , w_24244 );
not ( w_24244 , w_24245 );
and ( w_24245 , w_24242 , w_24243 );
buf ( w_24242 , \5797_b1 );
not ( w_24242 , w_24246 );
not ( w_24243 , w_24247 );
and ( w_24246 , w_24247 , \5797_b0 );
or ( \9605_b1 , \9600_b1 , \9604_b1 );
xor ( \9605_b0 , \9600_b0 , w_24248 );
not ( w_24248 , w_24249 );
and ( w_24249 , \9604_b1 , \9604_b0 );
or ( \9606_b1 , \5842_b1 , \7175_b1 );
not ( \7175_b1 , w_24250 );
and ( \9606_b0 , \5842_b0 , w_24251 );
and ( w_24250 , w_24251 , \7175_b0 );
or ( \9607_b1 , \5854_b1 , \7173_b1 );
not ( \7173_b1 , w_24252 );
and ( \9607_b0 , \5854_b0 , w_24253 );
and ( w_24252 , w_24253 , \7173_b0 );
or ( \9608_b1 , \9606_b1 , w_24255 );
not ( w_24255 , w_24256 );
and ( \9608_b0 , \9606_b0 , w_24257 );
and ( w_24256 ,  , w_24257 );
buf ( w_24255 , \9607_b1 );
not ( w_24255 , w_24258 );
not (  , w_24259 );
and ( w_24258 , w_24259 , \9607_b0 );
or ( \9609_b1 , \9608_b1 , w_24260 );
xor ( \9609_b0 , \9608_b0 , w_24262 );
not ( w_24262 , w_24263 );
and ( w_24263 , w_24260 , w_24261 );
buf ( w_24260 , \7181_b1 );
not ( w_24260 , w_24264 );
not ( w_24261 , w_24265 );
and ( w_24264 , w_24265 , \7181_b0 );
or ( \9610_b1 , \5861_b1 , \7192_b1 );
not ( \7192_b1 , w_24266 );
and ( \9610_b0 , \5861_b0 , w_24267 );
and ( w_24266 , w_24267 , \7192_b0 );
or ( \9611_b1 , \5873_b1 , \7190_b1 );
not ( \7190_b1 , w_24268 );
and ( \9611_b0 , \5873_b0 , w_24269 );
and ( w_24268 , w_24269 , \7190_b0 );
or ( \9612_b1 , \9610_b1 , w_24271 );
not ( w_24271 , w_24272 );
and ( \9612_b0 , \9610_b0 , w_24273 );
and ( w_24272 ,  , w_24273 );
buf ( w_24271 , \9611_b1 );
not ( w_24271 , w_24274 );
not (  , w_24275 );
and ( w_24274 , w_24275 , \9611_b0 );
or ( \9613_b1 , \9612_b1 , w_24276 );
xor ( \9613_b0 , \9612_b0 , w_24278 );
not ( w_24278 , w_24279 );
and ( w_24279 , w_24276 , w_24277 );
buf ( w_24276 , \7198_b1 );
not ( w_24276 , w_24280 );
not ( w_24277 , w_24281 );
and ( w_24280 , w_24281 , \7198_b0 );
or ( \9614_b1 , \9609_b1 , \9613_b1 );
xor ( \9614_b0 , \9609_b0 , w_24282 );
not ( w_24282 , w_24283 );
and ( w_24283 , \9613_b1 , \9613_b0 );
or ( \9615_b1 , \5881_b1 , \7203_b1 );
not ( \7203_b1 , w_24284 );
and ( \9615_b0 , \5881_b0 , w_24285 );
and ( w_24284 , w_24285 , \7203_b0 );
or ( \9616_b1 , \5893_b1 , \7201_b1 );
not ( \7201_b1 , w_24286 );
and ( \9616_b0 , \5893_b0 , w_24287 );
and ( w_24286 , w_24287 , \7201_b0 );
or ( \9617_b1 , \9615_b1 , w_24289 );
not ( w_24289 , w_24290 );
and ( \9617_b0 , \9615_b0 , w_24291 );
and ( w_24290 ,  , w_24291 );
buf ( w_24289 , \9616_b1 );
not ( w_24289 , w_24292 );
not (  , w_24293 );
and ( w_24292 , w_24293 , \9616_b0 );
or ( \9618_b1 , \9617_b1 , w_24294 );
xor ( \9618_b0 , \9617_b0 , w_24296 );
not ( w_24296 , w_24297 );
and ( w_24297 , w_24294 , w_24295 );
buf ( w_24294 , \6824_b1 );
not ( w_24294 , w_24298 );
not ( w_24295 , w_24299 );
and ( w_24298 , w_24299 , \6824_b0 );
or ( \9619_b1 , \9614_b1 , \9618_b1 );
xor ( \9619_b0 , \9614_b0 , w_24300 );
not ( w_24300 , w_24301 );
and ( w_24301 , \9618_b1 , \9618_b0 );
or ( \9620_b1 , \9605_b1 , \9619_b1 );
xor ( \9620_b0 , \9605_b0 , w_24302 );
not ( w_24302 , w_24303 );
and ( w_24303 , \9619_b1 , \9619_b0 );
or ( \9621_b1 , \5780_b1 , \7117_b1 );
not ( \7117_b1 , w_24304 );
and ( \9621_b0 , \5780_b0 , w_24305 );
and ( w_24304 , w_24305 , \7117_b0 );
or ( \9622_b1 , \5792_b1 , \7115_b1 );
not ( \7115_b1 , w_24306 );
and ( \9622_b0 , \5792_b0 , w_24307 );
and ( w_24306 , w_24307 , \7115_b0 );
or ( \9623_b1 , \9621_b1 , w_24309 );
not ( w_24309 , w_24310 );
and ( \9623_b0 , \9621_b0 , w_24311 );
and ( w_24310 ,  , w_24311 );
buf ( w_24309 , \9622_b1 );
not ( w_24309 , w_24312 );
not (  , w_24313 );
and ( w_24312 , w_24313 , \9622_b0 );
or ( \9624_b1 , \9623_b1 , w_24314 );
xor ( \9624_b0 , \9623_b0 , w_24316 );
not ( w_24316 , w_24317 );
and ( w_24317 , w_24314 , w_24315 );
buf ( w_24314 , \7123_b1 );
not ( w_24314 , w_24318 );
not ( w_24315 , w_24319 );
and ( w_24318 , w_24319 , \7123_b0 );
or ( \9625_b1 , \5799_b1 , \7140_b1 );
not ( \7140_b1 , w_24320 );
and ( \9625_b0 , \5799_b0 , w_24321 );
and ( w_24320 , w_24321 , \7140_b0 );
or ( \9626_b1 , \5811_b1 , \7138_b1 );
not ( \7138_b1 , w_24322 );
and ( \9626_b0 , \5811_b0 , w_24323 );
and ( w_24322 , w_24323 , \7138_b0 );
or ( \9627_b1 , \9625_b1 , w_24325 );
not ( w_24325 , w_24326 );
and ( \9627_b0 , \9625_b0 , w_24327 );
and ( w_24326 ,  , w_24327 );
buf ( w_24325 , \9626_b1 );
not ( w_24325 , w_24328 );
not (  , w_24329 );
and ( w_24328 , w_24329 , \9626_b0 );
or ( \9628_b1 , \9627_b1 , w_24330 );
xor ( \9628_b0 , \9627_b0 , w_24332 );
not ( w_24332 , w_24333 );
and ( w_24333 , w_24330 , w_24331 );
buf ( w_24330 , \7146_b1 );
not ( w_24330 , w_24334 );
not ( w_24331 , w_24335 );
and ( w_24334 , w_24335 , \7146_b0 );
or ( \9629_b1 , \9624_b1 , \9628_b1 );
xor ( \9629_b0 , \9624_b0 , w_24336 );
not ( w_24336 , w_24337 );
and ( w_24337 , \9628_b1 , \9628_b0 );
or ( \9630_b1 , \5819_b1 , \7157_b1 );
not ( \7157_b1 , w_24338 );
and ( \9630_b0 , \5819_b0 , w_24339 );
and ( w_24338 , w_24339 , \7157_b0 );
or ( \9631_b1 , \5831_b1 , \7155_b1 );
not ( \7155_b1 , w_24340 );
and ( \9631_b0 , \5831_b0 , w_24341 );
and ( w_24340 , w_24341 , \7155_b0 );
or ( \9632_b1 , \9630_b1 , w_24343 );
not ( w_24343 , w_24344 );
and ( \9632_b0 , \9630_b0 , w_24345 );
and ( w_24344 ,  , w_24345 );
buf ( w_24343 , \9631_b1 );
not ( w_24343 , w_24346 );
not (  , w_24347 );
and ( w_24346 , w_24347 , \9631_b0 );
or ( \9633_b1 , \9632_b1 , w_24348 );
xor ( \9633_b0 , \9632_b0 , w_24350 );
not ( w_24350 , w_24351 );
and ( w_24351 , w_24348 , w_24349 );
buf ( w_24348 , \7163_b1 );
not ( w_24348 , w_24352 );
not ( w_24349 , w_24353 );
and ( w_24352 , w_24353 , \7163_b0 );
or ( \9634_b1 , \9629_b1 , \9633_b1 );
xor ( \9634_b0 , \9629_b0 , w_24354 );
not ( w_24354 , w_24355 );
and ( w_24355 , \9633_b1 , \9633_b0 );
or ( \9635_b1 , \9620_b1 , \9634_b1 );
xor ( \9635_b0 , \9620_b0 , w_24356 );
not ( w_24356 , w_24357 );
and ( w_24357 , \9634_b1 , \9634_b0 );
or ( \9636_b1 , \9591_b1 , \9635_b1 );
xor ( \9636_b0 , \9591_b0 , w_24358 );
not ( w_24358 , w_24359 );
and ( w_24359 , \9635_b1 , \9635_b0 );
or ( \9637_b1 , \9577_b1 , \9636_b1 );
xor ( \9637_b0 , \9577_b0 , w_24360 );
not ( w_24360 , w_24361 );
and ( w_24361 , \9636_b1 , \9636_b0 );
or ( \9638_b1 , \9381_b1 , \9385_b1 );
not ( \9385_b1 , w_24362 );
and ( \9638_b0 , \9381_b0 , w_24363 );
and ( w_24362 , w_24363 , \9385_b0 );
or ( \9639_b1 , \9385_b1 , \9390_b1 );
not ( \9390_b1 , w_24364 );
and ( \9639_b0 , \9385_b0 , w_24365 );
and ( w_24364 , w_24365 , \9390_b0 );
or ( \9640_b1 , \9381_b1 , \9390_b1 );
not ( \9390_b1 , w_24366 );
and ( \9640_b0 , \9381_b0 , w_24367 );
and ( w_24366 , w_24367 , \9390_b0 );
or ( \9642_b1 , \9367_b1 , \9371_b1 );
not ( \9371_b1 , w_24368 );
and ( \9642_b0 , \9367_b0 , w_24369 );
and ( w_24368 , w_24369 , \9371_b0 );
or ( \9643_b1 , \9371_b1 , \9376_b1 );
not ( \9376_b1 , w_24370 );
and ( \9643_b0 , \9371_b0 , w_24371 );
and ( w_24370 , w_24371 , \9376_b0 );
or ( \9644_b1 , \9367_b1 , \9376_b1 );
not ( \9376_b1 , w_24372 );
and ( \9644_b0 , \9367_b0 , w_24373 );
and ( w_24372 , w_24373 , \9376_b0 );
or ( \9646_b1 , \9641_b1 , \9645_b1 );
xor ( \9646_b0 , \9641_b0 , w_24374 );
not ( w_24374 , w_24375 );
and ( w_24375 , \9645_b1 , \9645_b0 );
or ( \9647_b1 , \9447_b1 , \9461_b1 );
not ( \9461_b1 , w_24376 );
and ( \9647_b0 , \9447_b0 , w_24377 );
and ( w_24376 , w_24377 , \9461_b0 );
or ( \9648_b1 , \9461_b1 , \9476_b1 );
not ( \9476_b1 , w_24378 );
and ( \9648_b0 , \9461_b0 , w_24379 );
and ( w_24378 , w_24379 , \9476_b0 );
or ( \9649_b1 , \9447_b1 , \9476_b1 );
not ( \9476_b1 , w_24380 );
and ( \9649_b0 , \9447_b0 , w_24381 );
and ( w_24380 , w_24381 , \9476_b0 );
or ( \9651_b1 , \9646_b1 , \9650_b1 );
xor ( \9651_b0 , \9646_b0 , w_24382 );
not ( w_24382 , w_24383 );
and ( w_24383 , \9650_b1 , \9650_b0 );
or ( \9652_b1 , \9637_b1 , \9651_b1 );
xor ( \9652_b0 , \9637_b0 , w_24384 );
not ( w_24384 , w_24385 );
and ( w_24385 , \9651_b1 , \9651_b0 );
or ( \9653_b1 , \9523_b1 , \9652_b1 );
xor ( \9653_b0 , \9523_b0 , w_24386 );
not ( w_24386 , w_24387 );
and ( w_24387 , \9652_b1 , \9652_b0 );
or ( \9654_b1 , \9514_b1 , \9653_b1 );
xor ( \9654_b0 , \9514_b0 , w_24388 );
not ( w_24388 , w_24389 );
and ( w_24389 , \9653_b1 , \9653_b0 );
or ( \9655_b1 , \9339_b1 , \9353_b1 );
not ( \9353_b1 , w_24390 );
and ( \9655_b0 , \9339_b0 , w_24391 );
and ( w_24390 , w_24391 , \9353_b0 );
or ( \9656_b1 , \9353_b1 , \9492_b1 );
not ( \9492_b1 , w_24392 );
and ( \9656_b0 , \9353_b0 , w_24393 );
and ( w_24392 , w_24393 , \9492_b0 );
or ( \9657_b1 , \9339_b1 , \9492_b1 );
not ( \9492_b1 , w_24394 );
and ( \9657_b0 , \9339_b0 , w_24395 );
and ( w_24394 , w_24395 , \9492_b0 );
or ( \9659_b1 , \9654_b1 , w_24397 );
not ( w_24397 , w_24398 );
and ( \9659_b0 , \9654_b0 , w_24399 );
and ( w_24398 ,  , w_24399 );
buf ( w_24397 , \9658_b1 );
not ( w_24397 , w_24400 );
not (  , w_24401 );
and ( w_24400 , w_24401 , \9658_b0 );
or ( \9660_b1 , \9498_b1 , w_24403 );
not ( w_24403 , w_24404 );
and ( \9660_b0 , \9498_b0 , w_24405 );
and ( w_24404 ,  , w_24405 );
buf ( w_24403 , \9659_b1 );
not ( w_24403 , w_24406 );
not (  , w_24407 );
and ( w_24406 , w_24407 , \9659_b0 );
or ( \9661_b1 , \9335_b1 , w_24409 );
not ( w_24409 , w_24410 );
and ( \9661_b0 , \9335_b0 , w_24411 );
and ( w_24410 ,  , w_24411 );
buf ( w_24409 , \9660_b1 );
not ( w_24409 , w_24412 );
not (  , w_24413 );
and ( w_24412 , w_24413 , \9660_b0 );
or ( \9662_b1 , \9518_b1 , \9522_b1 );
not ( \9522_b1 , w_24414 );
and ( \9662_b0 , \9518_b0 , w_24415 );
and ( w_24414 , w_24415 , \9522_b0 );
or ( \9663_b1 , \9522_b1 , \9652_b1 );
not ( \9652_b1 , w_24416 );
and ( \9663_b0 , \9522_b0 , w_24417 );
and ( w_24416 , w_24417 , \9652_b0 );
or ( \9664_b1 , \9518_b1 , \9652_b1 );
not ( \9652_b1 , w_24418 );
and ( \9664_b0 , \9518_b0 , w_24419 );
and ( w_24418 , w_24419 , \9652_b0 );
or ( \9666_b1 , \9641_b1 , \9645_b1 );
not ( \9645_b1 , w_24420 );
and ( \9666_b0 , \9641_b0 , w_24421 );
and ( w_24420 , w_24421 , \9645_b0 );
or ( \9667_b1 , \9645_b1 , \9650_b1 );
not ( \9650_b1 , w_24422 );
and ( \9667_b0 , \9645_b0 , w_24423 );
and ( w_24422 , w_24423 , \9650_b0 );
or ( \9668_b1 , \9641_b1 , \9650_b1 );
not ( \9650_b1 , w_24424 );
and ( \9668_b0 , \9641_b0 , w_24425 );
and ( w_24424 , w_24425 , \9650_b0 );
or ( \9670_b1 , \9581_b1 , \9590_b1 );
not ( \9590_b1 , w_24426 );
and ( \9670_b0 , \9581_b0 , w_24427 );
and ( w_24426 , w_24427 , \9590_b0 );
or ( \9671_b1 , \9590_b1 , \9635_b1 );
not ( \9635_b1 , w_24428 );
and ( \9671_b0 , \9590_b0 , w_24429 );
and ( w_24428 , w_24429 , \9635_b0 );
or ( \9672_b1 , \9581_b1 , \9635_b1 );
not ( \9635_b1 , w_24430 );
and ( \9672_b0 , \9581_b0 , w_24431 );
and ( w_24430 , w_24431 , \9635_b0 );
or ( \9674_b1 , \9669_b1 , \9673_b1 );
xor ( \9674_b0 , \9669_b0 , w_24432 );
not ( w_24432 , w_24433 );
and ( w_24433 , \9673_b1 , \9673_b0 );
or ( \9675_b1 , \9550_b1 , \9561_b1 );
not ( \9561_b1 , w_24434 );
and ( \9675_b0 , \9550_b0 , w_24435 );
and ( w_24434 , w_24435 , \9561_b0 );
or ( \9676_b1 , \9561_b1 , \9576_b1 );
not ( \9576_b1 , w_24436 );
and ( \9676_b0 , \9561_b0 , w_24437 );
and ( w_24436 , w_24437 , \9576_b0 );
or ( \9677_b1 , \9550_b1 , \9576_b1 );
not ( \9576_b1 , w_24438 );
and ( \9677_b0 , \9550_b0 , w_24439 );
and ( w_24438 , w_24439 , \9576_b0 );
or ( \9679_b1 , \9674_b1 , \9678_b1 );
xor ( \9679_b0 , \9674_b0 , w_24440 );
not ( w_24440 , w_24441 );
and ( w_24441 , \9678_b1 , \9678_b0 );
or ( \9680_b1 , \9665_b1 , \9679_b1 );
xor ( \9680_b0 , \9665_b0 , w_24442 );
not ( w_24442 , w_24443 );
and ( w_24443 , \9679_b1 , \9679_b0 );
or ( \9681_b1 , \9506_b1 , \9510_b1 );
not ( \9510_b1 , w_24444 );
and ( \9681_b0 , \9506_b0 , w_24445 );
and ( w_24444 , w_24445 , \9510_b0 );
or ( \9682_b1 , \9510_b1 , \9512_b1 );
not ( \9512_b1 , w_24446 );
and ( \9682_b0 , \9510_b0 , w_24447 );
and ( w_24446 , w_24447 , \9512_b0 );
or ( \9683_b1 , \9506_b1 , \9512_b1 );
not ( \9512_b1 , w_24448 );
and ( \9683_b0 , \9506_b0 , w_24449 );
and ( w_24448 , w_24449 , \9512_b0 );
or ( \9685_b1 , \9577_b1 , \9636_b1 );
not ( \9636_b1 , w_24450 );
and ( \9685_b0 , \9577_b0 , w_24451 );
and ( w_24450 , w_24451 , \9636_b0 );
or ( \9686_b1 , \9636_b1 , \9651_b1 );
not ( \9651_b1 , w_24452 );
and ( \9686_b0 , \9636_b0 , w_24453 );
and ( w_24452 , w_24453 , \9651_b0 );
or ( \9687_b1 , \9577_b1 , \9651_b1 );
not ( \9651_b1 , w_24454 );
and ( \9687_b0 , \9577_b0 , w_24455 );
and ( w_24454 , w_24455 , \9651_b0 );
or ( \9689_b1 , \9684_b1 , \9688_b1 );
xor ( \9689_b0 , \9684_b0 , w_24456 );
not ( w_24456 , w_24457 );
and ( w_24457 , \9688_b1 , \9688_b0 );
or ( \9690_b1 , \9595_b1 , \9599_b1 );
not ( \9599_b1 , w_24458 );
and ( \9690_b0 , \9595_b0 , w_24459 );
and ( w_24458 , w_24459 , \9599_b0 );
or ( \9691_b1 , \9599_b1 , \9604_b1 );
not ( \9604_b1 , w_24460 );
and ( \9691_b0 , \9599_b0 , w_24461 );
and ( w_24460 , w_24461 , \9604_b0 );
or ( \9692_b1 , \9595_b1 , \9604_b1 );
not ( \9604_b1 , w_24462 );
and ( \9692_b0 , \9595_b0 , w_24463 );
and ( w_24462 , w_24463 , \9604_b0 );
or ( \9694_b1 , \9539_b1 , \9543_b1 );
not ( \9543_b1 , w_24464 );
and ( \9694_b0 , \9539_b0 , w_24465 );
and ( w_24464 , w_24465 , \9543_b0 );
or ( \9695_b1 , \9543_b1 , \9548_b1 );
not ( \9548_b1 , w_24466 );
and ( \9695_b0 , \9543_b0 , w_24467 );
and ( w_24466 , w_24467 , \9548_b0 );
or ( \9696_b1 , \9539_b1 , \9548_b1 );
not ( \9548_b1 , w_24468 );
and ( \9696_b0 , \9539_b0 , w_24469 );
and ( w_24468 , w_24469 , \9548_b0 );
or ( \9698_b1 , \9693_b1 , \9697_b1 );
xor ( \9698_b0 , \9693_b0 , w_24470 );
not ( w_24470 , w_24471 );
and ( w_24471 , \9697_b1 , \9697_b0 );
or ( \9699_b1 , \9527_b1 , \9531_b1 );
not ( \9531_b1 , w_24472 );
and ( \9699_b0 , \9527_b0 , w_24473 );
and ( w_24472 , w_24473 , \9531_b0 );
or ( \9700_b1 , \9531_b1 , \9534_b1 );
not ( \9534_b1 , w_24474 );
and ( \9700_b0 , \9531_b0 , w_24475 );
and ( w_24474 , w_24475 , \9534_b0 );
or ( \9701_b1 , \9527_b1 , \9534_b1 );
not ( \9534_b1 , w_24476 );
and ( \9701_b0 , \9527_b0 , w_24477 );
and ( w_24476 , w_24477 , \9534_b0 );
or ( \9703_b1 , \9698_b1 , \9702_b1 );
xor ( \9703_b0 , \9698_b0 , w_24478 );
not ( w_24478 , w_24479 );
and ( w_24479 , \9702_b1 , \9702_b0 );
or ( \9704_b1 , \5923_b1 , \9584_b1 );
not ( \9584_b1 , w_24480 );
and ( \9704_b0 , \5923_b0 , w_24481 );
and ( w_24480 , w_24481 , \9584_b0 );
or ( \9705_b1 , \9584_b1 , \9589_b1 );
not ( \9589_b1 , w_24482 );
and ( \9705_b0 , \9584_b0 , w_24483 );
and ( w_24482 , w_24483 , \9589_b0 );
or ( \9706_b1 , \5923_b1 , \9589_b1 );
not ( \9589_b1 , w_24484 );
and ( \9706_b0 , \5923_b0 , w_24485 );
and ( w_24484 , w_24485 , \9589_b0 );
or ( \9708_b1 , \9624_b1 , \9628_b1 );
not ( \9628_b1 , w_24486 );
and ( \9708_b0 , \9624_b0 , w_24487 );
and ( w_24486 , w_24487 , \9628_b0 );
or ( \9709_b1 , \9628_b1 , \9633_b1 );
not ( \9633_b1 , w_24488 );
and ( \9709_b0 , \9628_b0 , w_24489 );
and ( w_24488 , w_24489 , \9633_b0 );
or ( \9710_b1 , \9624_b1 , \9633_b1 );
not ( \9633_b1 , w_24490 );
and ( \9710_b0 , \9624_b0 , w_24491 );
and ( w_24490 , w_24491 , \9633_b0 );
or ( \9712_b1 , \9707_b1 , \9711_b1 );
xor ( \9712_b0 , \9707_b0 , w_24492 );
not ( w_24492 , w_24493 );
and ( w_24493 , \9711_b1 , \9711_b0 );
or ( \9713_b1 , \9609_b1 , \9613_b1 );
not ( \9613_b1 , w_24494 );
and ( \9713_b0 , \9609_b0 , w_24495 );
and ( w_24494 , w_24495 , \9613_b0 );
or ( \9714_b1 , \9613_b1 , \9618_b1 );
not ( \9618_b1 , w_24496 );
and ( \9714_b0 , \9613_b0 , w_24497 );
and ( w_24496 , w_24497 , \9618_b0 );
or ( \9715_b1 , \9609_b1 , \9618_b1 );
not ( \9618_b1 , w_24498 );
and ( \9715_b0 , \9609_b0 , w_24499 );
and ( w_24498 , w_24499 , \9618_b0 );
or ( \9717_b1 , \9712_b1 , \9716_b1 );
xor ( \9717_b0 , \9712_b0 , w_24500 );
not ( w_24500 , w_24501 );
and ( w_24501 , \9716_b1 , \9716_b0 );
or ( \9718_b1 , \9703_b1 , \9717_b1 );
xor ( \9718_b0 , \9703_b0 , w_24502 );
not ( w_24502 , w_24503 );
and ( w_24503 , \9717_b1 , \9717_b0 );
or ( \9719_b1 , \9605_b1 , \9619_b1 );
not ( \9619_b1 , w_24504 );
and ( \9719_b0 , \9605_b0 , w_24505 );
and ( w_24504 , w_24505 , \9619_b0 );
or ( \9720_b1 , \9619_b1 , \9634_b1 );
not ( \9634_b1 , w_24506 );
and ( \9720_b0 , \9619_b0 , w_24507 );
and ( w_24506 , w_24507 , \9634_b0 );
or ( \9721_b1 , \9605_b1 , \9634_b1 );
not ( \9634_b1 , w_24508 );
and ( \9721_b0 , \9605_b0 , w_24509 );
and ( w_24508 , w_24509 , \9634_b0 );
or ( \9723_b1 , \5873_b1 , \7192_b1 );
not ( \7192_b1 , w_24510 );
and ( \9723_b0 , \5873_b0 , w_24511 );
and ( w_24510 , w_24511 , \7192_b0 );
or ( \9724_b1 , \5842_b1 , \7190_b1 );
not ( \7190_b1 , w_24512 );
and ( \9724_b0 , \5842_b0 , w_24513 );
and ( w_24512 , w_24513 , \7190_b0 );
or ( \9725_b1 , \9723_b1 , w_24515 );
not ( w_24515 , w_24516 );
and ( \9725_b0 , \9723_b0 , w_24517 );
and ( w_24516 ,  , w_24517 );
buf ( w_24515 , \9724_b1 );
not ( w_24515 , w_24518 );
not (  , w_24519 );
and ( w_24518 , w_24519 , \9724_b0 );
or ( \9726_b1 , \9725_b1 , w_24520 );
xor ( \9726_b0 , \9725_b0 , w_24522 );
not ( w_24522 , w_24523 );
and ( w_24523 , w_24520 , w_24521 );
buf ( w_24520 , \7198_b1 );
not ( w_24520 , w_24524 );
not ( w_24521 , w_24525 );
and ( w_24524 , w_24525 , \7198_b0 );
or ( \9727_b1 , \5893_b1 , \7203_b1 );
not ( \7203_b1 , w_24526 );
and ( \9727_b0 , \5893_b0 , w_24527 );
and ( w_24526 , w_24527 , \7203_b0 );
or ( \9728_b1 , \5861_b1 , \7201_b1 );
not ( \7201_b1 , w_24528 );
and ( \9728_b0 , \5861_b0 , w_24529 );
and ( w_24528 , w_24529 , \7201_b0 );
or ( \9729_b1 , \9727_b1 , w_24531 );
not ( w_24531 , w_24532 );
and ( \9729_b0 , \9727_b0 , w_24533 );
and ( w_24532 ,  , w_24533 );
buf ( w_24531 , \9728_b1 );
not ( w_24531 , w_24534 );
not (  , w_24535 );
and ( w_24534 , w_24535 , \9728_b0 );
or ( \9730_b1 , \9729_b1 , w_24536 );
xor ( \9730_b0 , \9729_b0 , w_24538 );
not ( w_24538 , w_24539 );
and ( w_24539 , w_24536 , w_24537 );
buf ( w_24536 , \6824_b1 );
not ( w_24536 , w_24540 );
not ( w_24537 , w_24541 );
and ( w_24540 , w_24541 , \6824_b0 );
or ( \9731_b1 , \9726_b1 , \9730_b1 );
xor ( \9731_b0 , \9726_b0 , w_24542 );
not ( w_24542 , w_24543 );
and ( w_24543 , \9730_b1 , \9730_b0 );
or ( \9732_b1 , \5918_b1 , \5750_b1 );
not ( \5750_b1 , w_24544 );
and ( \9732_b0 , \5918_b0 , w_24545 );
and ( w_24544 , w_24545 , \5750_b0 );
or ( \9733_b1 , \5881_b1 , \5748_b1 );
not ( \5748_b1 , w_24546 );
and ( \9733_b0 , \5881_b0 , w_24547 );
and ( w_24546 , w_24547 , \5748_b0 );
or ( \9734_b1 , \9732_b1 , w_24549 );
not ( w_24549 , w_24550 );
and ( \9734_b0 , \9732_b0 , w_24551 );
and ( w_24550 ,  , w_24551 );
buf ( w_24549 , \9733_b1 );
not ( w_24549 , w_24552 );
not (  , w_24553 );
and ( w_24552 , w_24553 , \9733_b0 );
or ( \9735_b1 , \9734_b1 , w_24554 );
xor ( \9735_b0 , \9734_b0 , w_24556 );
not ( w_24556 , w_24557 );
and ( w_24557 , w_24554 , w_24555 );
buf ( w_24554 , \5755_b1 );
not ( w_24554 , w_24558 );
not ( w_24555 , w_24559 );
and ( w_24558 , w_24559 , \5755_b0 );
or ( \9736_b1 , \9731_b1 , \9735_b1 );
xor ( \9736_b0 , \9731_b0 , w_24560 );
not ( w_24560 , w_24561 );
and ( w_24561 , \9735_b1 , \9735_b0 );
or ( \9737_b1 , \5811_b1 , \7140_b1 );
not ( \7140_b1 , w_24562 );
and ( \9737_b0 , \5811_b0 , w_24563 );
and ( w_24562 , w_24563 , \7140_b0 );
or ( \9738_b1 , \5780_b1 , \7138_b1 );
not ( \7138_b1 , w_24564 );
and ( \9738_b0 , \5780_b0 , w_24565 );
and ( w_24564 , w_24565 , \7138_b0 );
or ( \9739_b1 , \9737_b1 , w_24567 );
not ( w_24567 , w_24568 );
and ( \9739_b0 , \9737_b0 , w_24569 );
and ( w_24568 ,  , w_24569 );
buf ( w_24567 , \9738_b1 );
not ( w_24567 , w_24570 );
not (  , w_24571 );
and ( w_24570 , w_24571 , \9738_b0 );
or ( \9740_b1 , \9739_b1 , w_24572 );
xor ( \9740_b0 , \9739_b0 , w_24574 );
not ( w_24574 , w_24575 );
and ( w_24575 , w_24572 , w_24573 );
buf ( w_24572 , \7146_b1 );
not ( w_24572 , w_24576 );
not ( w_24573 , w_24577 );
and ( w_24576 , w_24577 , \7146_b0 );
or ( \9741_b1 , \5831_b1 , \7157_b1 );
not ( \7157_b1 , w_24578 );
and ( \9741_b0 , \5831_b0 , w_24579 );
and ( w_24578 , w_24579 , \7157_b0 );
or ( \9742_b1 , \5799_b1 , \7155_b1 );
not ( \7155_b1 , w_24580 );
and ( \9742_b0 , \5799_b0 , w_24581 );
and ( w_24580 , w_24581 , \7155_b0 );
or ( \9743_b1 , \9741_b1 , w_24583 );
not ( w_24583 , w_24584 );
and ( \9743_b0 , \9741_b0 , w_24585 );
and ( w_24584 ,  , w_24585 );
buf ( w_24583 , \9742_b1 );
not ( w_24583 , w_24586 );
not (  , w_24587 );
and ( w_24586 , w_24587 , \9742_b0 );
or ( \9744_b1 , \9743_b1 , w_24588 );
xor ( \9744_b0 , \9743_b0 , w_24590 );
not ( w_24590 , w_24591 );
and ( w_24591 , w_24588 , w_24589 );
buf ( w_24588 , \7163_b1 );
not ( w_24588 , w_24592 );
not ( w_24589 , w_24593 );
and ( w_24592 , w_24593 , \7163_b0 );
or ( \9745_b1 , \9740_b1 , \9744_b1 );
xor ( \9745_b0 , \9740_b0 , w_24594 );
not ( w_24594 , w_24595 );
and ( w_24595 , \9744_b1 , \9744_b0 );
or ( \9746_b1 , \5854_b1 , \7175_b1 );
not ( \7175_b1 , w_24596 );
and ( \9746_b0 , \5854_b0 , w_24597 );
and ( w_24596 , w_24597 , \7175_b0 );
or ( \9747_b1 , \5819_b1 , \7173_b1 );
not ( \7173_b1 , w_24598 );
and ( \9747_b0 , \5819_b0 , w_24599 );
and ( w_24598 , w_24599 , \7173_b0 );
or ( \9748_b1 , \9746_b1 , w_24601 );
not ( w_24601 , w_24602 );
and ( \9748_b0 , \9746_b0 , w_24603 );
and ( w_24602 ,  , w_24603 );
buf ( w_24601 , \9747_b1 );
not ( w_24601 , w_24604 );
not (  , w_24605 );
and ( w_24604 , w_24605 , \9747_b0 );
or ( \9749_b1 , \9748_b1 , w_24606 );
xor ( \9749_b0 , \9748_b0 , w_24608 );
not ( w_24608 , w_24609 );
and ( w_24609 , w_24606 , w_24607 );
buf ( w_24606 , \7181_b1 );
not ( w_24606 , w_24610 );
not ( w_24607 , w_24611 );
and ( w_24610 , w_24611 , \7181_b0 );
or ( \9750_b1 , \9745_b1 , \9749_b1 );
xor ( \9750_b0 , \9745_b0 , w_24612 );
not ( w_24612 , w_24613 );
and ( w_24613 , \9749_b1 , \9749_b0 );
or ( \9751_b1 , \9736_b1 , \9750_b1 );
xor ( \9751_b0 , \9736_b0 , w_24614 );
not ( w_24614 , w_24615 );
and ( w_24615 , \9750_b1 , \9750_b0 );
buf ( \9752_b1 , \7088_b1 );
not ( \9752_b1 , w_24616 );
not ( \9752_b0 , w_24617 );
and ( w_24616 , w_24617 , \7088_b0 );
or ( \9753_b1 , \5770_b1 , \7099_b1 );
not ( \7099_b1 , w_24618 );
and ( \9753_b0 , \5770_b0 , w_24619 );
and ( w_24618 , w_24619 , \7099_b0 );
or ( \9754_b1 , \5737_b1 , \7097_b1 );
not ( \7097_b1 , w_24620 );
and ( \9754_b0 , \5737_b0 , w_24621 );
and ( w_24620 , w_24621 , \7097_b0 );
or ( \9755_b1 , \9753_b1 , w_24623 );
not ( w_24623 , w_24624 );
and ( \9755_b0 , \9753_b0 , w_24625 );
and ( w_24624 ,  , w_24625 );
buf ( w_24623 , \9754_b1 );
not ( w_24623 , w_24626 );
not (  , w_24627 );
and ( w_24626 , w_24627 , \9754_b0 );
or ( \9756_b1 , \9755_b1 , w_24628 );
xor ( \9756_b0 , \9755_b0 , w_24630 );
not ( w_24630 , w_24631 );
and ( w_24631 , w_24628 , w_24629 );
buf ( w_24628 , \7105_b1 );
not ( w_24628 , w_24632 );
not ( w_24629 , w_24633 );
and ( w_24632 , w_24633 , \7105_b0 );
or ( \9757_b1 , \9752_b1 , \9756_b1 );
xor ( \9757_b0 , \9752_b0 , w_24634 );
not ( w_24634 , w_24635 );
and ( w_24635 , \9756_b1 , \9756_b0 );
or ( \9758_b1 , \5792_b1 , \7117_b1 );
not ( \7117_b1 , w_24636 );
and ( \9758_b0 , \5792_b0 , w_24637 );
and ( w_24636 , w_24637 , \7117_b0 );
or ( \9759_b1 , \5758_b1 , \7115_b1 );
not ( \7115_b1 , w_24638 );
and ( \9759_b0 , \5758_b0 , w_24639 );
and ( w_24638 , w_24639 , \7115_b0 );
or ( \9760_b1 , \9758_b1 , w_24641 );
not ( w_24641 , w_24642 );
and ( \9760_b0 , \9758_b0 , w_24643 );
and ( w_24642 ,  , w_24643 );
buf ( w_24641 , \9759_b1 );
not ( w_24641 , w_24644 );
not (  , w_24645 );
and ( w_24644 , w_24645 , \9759_b0 );
or ( \9761_b1 , \9760_b1 , w_24646 );
xor ( \9761_b0 , \9760_b0 , w_24648 );
not ( w_24648 , w_24649 );
and ( w_24649 , w_24646 , w_24647 );
buf ( w_24646 , \7123_b1 );
not ( w_24646 , w_24650 );
not ( w_24647 , w_24651 );
and ( w_24650 , w_24651 , \7123_b0 );
or ( \9762_b1 , \9757_b1 , \9761_b1 );
xor ( \9762_b0 , \9757_b0 , w_24652 );
not ( w_24652 , w_24653 );
and ( w_24653 , \9761_b1 , \9761_b0 );
or ( \9763_b1 , \9751_b1 , \9762_b1 );
xor ( \9763_b0 , \9751_b0 , w_24654 );
not ( w_24654 , w_24655 );
and ( w_24655 , \9762_b1 , \9762_b0 );
or ( \9764_b1 , \9722_b1 , \9763_b1 );
xor ( \9764_b0 , \9722_b0 , w_24656 );
not ( w_24656 , w_24657 );
and ( w_24657 , \9763_b1 , \9763_b0 );
or ( \9765_b1 , \6057_b1 , \5891_b1 );
not ( \5891_b1 , w_24658 );
and ( \9765_b0 , \6057_b0 , w_24659 );
and ( w_24658 , w_24659 , \5891_b0 );
or ( \9766_b1 , \6029_b1 , \5889_b1 );
not ( \5889_b1 , w_24660 );
and ( \9766_b0 , \6029_b0 , w_24661 );
and ( w_24660 , w_24661 , \5889_b0 );
or ( \9767_b1 , \9765_b1 , w_24663 );
not ( w_24663 , w_24664 );
and ( \9767_b0 , \9765_b0 , w_24665 );
and ( w_24664 ,  , w_24665 );
buf ( w_24663 , \9766_b1 );
not ( w_24663 , w_24666 );
not (  , w_24667 );
and ( w_24666 , w_24667 , \9766_b0 );
or ( \9768_b1 , \9767_b1 , w_24668 );
xor ( \9768_b0 , \9767_b0 , w_24670 );
not ( w_24670 , w_24671 );
and ( w_24671 , w_24668 , w_24669 );
buf ( w_24668 , \5898_b1 );
not ( w_24668 , w_24672 );
not ( w_24669 , w_24673 );
and ( w_24672 , w_24673 , \5898_b0 );
or ( \9769_b1 , \6065_b1 , \5916_b1 );
not ( \5916_b1 , w_24674 );
and ( \9769_b0 , \6065_b0 , w_24675 );
and ( w_24674 , w_24675 , \5916_b0 );
or ( \9770_b1 , \6048_b1 , \5914_b1 );
not ( \5914_b1 , w_24676 );
and ( \9770_b0 , \6048_b0 , w_24677 );
and ( w_24676 , w_24677 , \5914_b0 );
or ( \9771_b1 , \9769_b1 , w_24679 );
not ( w_24679 , w_24680 );
and ( \9771_b0 , \9769_b0 , w_24681 );
and ( w_24680 ,  , w_24681 );
buf ( w_24679 , \9770_b1 );
not ( w_24679 , w_24682 );
not (  , w_24683 );
and ( w_24682 , w_24683 , \9770_b0 );
or ( \9772_b1 , \9771_b1 , w_24684 );
xor ( \9772_b0 , \9771_b0 , w_24686 );
not ( w_24686 , w_24687 );
and ( w_24687 , w_24684 , w_24685 );
buf ( w_24684 , \5923_b1 );
not ( w_24684 , w_24688 );
not ( w_24685 , w_24689 );
and ( w_24688 , w_24689 , \5923_b0 );
or ( \9773_b1 , \9768_b1 , \9772_b1 );
xor ( \9773_b0 , \9768_b0 , w_24690 );
not ( w_24690 , w_24691 );
and ( w_24691 , \9772_b1 , \9772_b0 );
or ( \9774_b1 , \5998_b1 , \5829_b1 );
not ( \5829_b1 , w_24692 );
and ( \9774_b0 , \5998_b0 , w_24693 );
and ( w_24692 , w_24693 , \5829_b0 );
or ( \9775_b1 , \5967_b1 , \5827_b1 );
not ( \5827_b1 , w_24694 );
and ( \9775_b0 , \5967_b0 , w_24695 );
and ( w_24694 , w_24695 , \5827_b0 );
or ( \9776_b1 , \9774_b1 , w_24697 );
not ( w_24697 , w_24698 );
and ( \9776_b0 , \9774_b0 , w_24699 );
and ( w_24698 ,  , w_24699 );
buf ( w_24697 , \9775_b1 );
not ( w_24697 , w_24700 );
not (  , w_24701 );
and ( w_24700 , w_24701 , \9775_b0 );
or ( \9777_b1 , \9776_b1 , w_24702 );
xor ( \9777_b0 , \9776_b0 , w_24704 );
not ( w_24704 , w_24705 );
and ( w_24705 , w_24702 , w_24703 );
buf ( w_24702 , \5836_b1 );
not ( w_24702 , w_24706 );
not ( w_24703 , w_24707 );
and ( w_24706 , w_24707 , \5836_b0 );
or ( \9778_b1 , \6018_b1 , \5852_b1 );
not ( \5852_b1 , w_24708 );
and ( \9778_b0 , \6018_b0 , w_24709 );
and ( w_24708 , w_24709 , \5852_b0 );
or ( \9779_b1 , \5986_b1 , \5850_b1 );
not ( \5850_b1 , w_24710 );
and ( \9779_b0 , \5986_b0 , w_24711 );
and ( w_24710 , w_24711 , \5850_b0 );
or ( \9780_b1 , \9778_b1 , w_24713 );
not ( w_24713 , w_24714 );
and ( \9780_b0 , \9778_b0 , w_24715 );
and ( w_24714 ,  , w_24715 );
buf ( w_24713 , \9779_b1 );
not ( w_24713 , w_24716 );
not (  , w_24717 );
and ( w_24716 , w_24717 , \9779_b0 );
or ( \9781_b1 , \9780_b1 , w_24718 );
xor ( \9781_b0 , \9780_b0 , w_24720 );
not ( w_24720 , w_24721 );
and ( w_24721 , w_24718 , w_24719 );
buf ( w_24718 , \5859_b1 );
not ( w_24718 , w_24722 );
not ( w_24719 , w_24723 );
and ( w_24722 , w_24723 , \5859_b0 );
or ( \9782_b1 , \9777_b1 , \9781_b1 );
xor ( \9782_b0 , \9777_b0 , w_24724 );
not ( w_24724 , w_24725 );
and ( w_24725 , \9781_b1 , \9781_b0 );
or ( \9783_b1 , \6041_b1 , \5871_b1 );
not ( \5871_b1 , w_24726 );
and ( \9783_b0 , \6041_b0 , w_24727 );
and ( w_24726 , w_24727 , \5871_b0 );
or ( \9784_b1 , \6006_b1 , \5869_b1 );
not ( \5869_b1 , w_24728 );
and ( \9784_b0 , \6006_b0 , w_24729 );
and ( w_24728 , w_24729 , \5869_b0 );
or ( \9785_b1 , \9783_b1 , w_24731 );
not ( w_24731 , w_24732 );
and ( \9785_b0 , \9783_b0 , w_24733 );
and ( w_24732 ,  , w_24733 );
buf ( w_24731 , \9784_b1 );
not ( w_24731 , w_24734 );
not (  , w_24735 );
and ( w_24734 , w_24735 , \9784_b0 );
or ( \9786_b1 , \9785_b1 , w_24736 );
xor ( \9786_b0 , \9785_b0 , w_24738 );
not ( w_24738 , w_24739 );
and ( w_24739 , w_24736 , w_24737 );
buf ( w_24736 , \5878_b1 );
not ( w_24736 , w_24740 );
not ( w_24737 , w_24741 );
and ( w_24740 , w_24741 , \5878_b0 );
or ( \9787_b1 , \9782_b1 , \9786_b1 );
xor ( \9787_b0 , \9782_b0 , w_24742 );
not ( w_24742 , w_24743 );
and ( w_24743 , \9786_b1 , \9786_b0 );
or ( \9788_b1 , \9773_b1 , \9787_b1 );
xor ( \9788_b0 , \9773_b0 , w_24744 );
not ( w_24744 , w_24745 );
and ( w_24745 , \9787_b1 , \9787_b0 );
or ( \9789_b1 , \5937_b1 , \5768_b1 );
not ( \5768_b1 , w_24746 );
and ( \9789_b0 , \5937_b0 , w_24747 );
and ( w_24746 , w_24747 , \5768_b0 );
or ( \9790_b1 , \5906_b1 , \5766_b1 );
not ( \5766_b1 , w_24748 );
and ( \9790_b0 , \5906_b0 , w_24749 );
and ( w_24748 , w_24749 , \5766_b0 );
or ( \9791_b1 , \9789_b1 , w_24751 );
not ( w_24751 , w_24752 );
and ( \9791_b0 , \9789_b0 , w_24753 );
and ( w_24752 ,  , w_24753 );
buf ( w_24751 , \9790_b1 );
not ( w_24751 , w_24754 );
not (  , w_24755 );
and ( w_24754 , w_24755 , \9790_b0 );
or ( \9792_b1 , \9791_b1 , w_24756 );
xor ( \9792_b0 , \9791_b0 , w_24758 );
not ( w_24758 , w_24759 );
and ( w_24759 , w_24756 , w_24757 );
buf ( w_24756 , \5775_b1 );
not ( w_24756 , w_24760 );
not ( w_24757 , w_24761 );
and ( w_24760 , w_24761 , \5775_b0 );
or ( \9793_b1 , \5957_b1 , \5790_b1 );
not ( \5790_b1 , w_24762 );
and ( \9793_b0 , \5957_b0 , w_24763 );
and ( w_24762 , w_24763 , \5790_b0 );
or ( \9794_b1 , \5925_b1 , \5788_b1 );
not ( \5788_b1 , w_24764 );
and ( \9794_b0 , \5925_b0 , w_24765 );
and ( w_24764 , w_24765 , \5788_b0 );
or ( \9795_b1 , \9793_b1 , w_24767 );
not ( w_24767 , w_24768 );
and ( \9795_b0 , \9793_b0 , w_24769 );
and ( w_24768 ,  , w_24769 );
buf ( w_24767 , \9794_b1 );
not ( w_24767 , w_24770 );
not (  , w_24771 );
and ( w_24770 , w_24771 , \9794_b0 );
or ( \9796_b1 , \9795_b1 , w_24772 );
xor ( \9796_b0 , \9795_b0 , w_24774 );
not ( w_24774 , w_24775 );
and ( w_24775 , w_24772 , w_24773 );
buf ( w_24772 , \5797_b1 );
not ( w_24772 , w_24776 );
not ( w_24773 , w_24777 );
and ( w_24776 , w_24777 , \5797_b0 );
or ( \9797_b1 , \9792_b1 , \9796_b1 );
xor ( \9797_b0 , \9792_b0 , w_24778 );
not ( w_24778 , w_24779 );
and ( w_24779 , \9796_b1 , \9796_b0 );
or ( \9798_b1 , \5979_b1 , \5809_b1 );
not ( \5809_b1 , w_24780 );
and ( \9798_b0 , \5979_b0 , w_24781 );
and ( w_24780 , w_24781 , \5809_b0 );
or ( \9799_b1 , \5945_b1 , \5807_b1 );
not ( \5807_b1 , w_24782 );
and ( \9799_b0 , \5945_b0 , w_24783 );
and ( w_24782 , w_24783 , \5807_b0 );
or ( \9800_b1 , \9798_b1 , w_24785 );
not ( w_24785 , w_24786 );
and ( \9800_b0 , \9798_b0 , w_24787 );
and ( w_24786 ,  , w_24787 );
buf ( w_24785 , \9799_b1 );
not ( w_24785 , w_24788 );
not (  , w_24789 );
and ( w_24788 , w_24789 , \9799_b0 );
or ( \9801_b1 , \9800_b1 , w_24790 );
xor ( \9801_b0 , \9800_b0 , w_24792 );
not ( w_24792 , w_24793 );
and ( w_24793 , w_24790 , w_24791 );
buf ( w_24790 , \5816_b1 );
not ( w_24790 , w_24794 );
not ( w_24791 , w_24795 );
and ( w_24794 , w_24795 , \5816_b0 );
or ( \9802_b1 , \9797_b1 , \9801_b1 );
xor ( \9802_b0 , \9797_b0 , w_24796 );
not ( w_24796 , w_24797 );
and ( w_24797 , \9801_b1 , \9801_b0 );
or ( \9803_b1 , \9788_b1 , \9802_b1 );
xor ( \9803_b0 , \9788_b0 , w_24798 );
not ( w_24798 , w_24799 );
and ( w_24799 , \9802_b1 , \9802_b0 );
or ( \9804_b1 , \9764_b1 , \9803_b1 );
xor ( \9804_b0 , \9764_b0 , w_24800 );
not ( w_24800 , w_24801 );
and ( w_24801 , \9803_b1 , \9803_b0 );
or ( \9805_b1 , \9718_b1 , \9804_b1 );
xor ( \9805_b0 , \9718_b0 , w_24802 );
not ( w_24802 , w_24803 );
and ( w_24803 , \9804_b1 , \9804_b0 );
or ( \9806_b1 , \9566_b1 , \9570_b1 );
not ( \9570_b1 , w_24804 );
and ( \9806_b0 , \9566_b0 , w_24805 );
and ( w_24804 , w_24805 , \9570_b0 );
or ( \9807_b1 , \9570_b1 , \9575_b1 );
not ( \9575_b1 , w_24806 );
and ( \9807_b0 , \9570_b0 , w_24807 );
and ( w_24806 , w_24807 , \9575_b0 );
or ( \9808_b1 , \9566_b1 , \9575_b1 );
not ( \9575_b1 , w_24808 );
and ( \9808_b0 , \9566_b0 , w_24809 );
and ( w_24808 , w_24809 , \9575_b0 );
or ( \9810_b1 , \9554_b1 , \9558_b1 );
not ( \9558_b1 , w_24810 );
and ( \9810_b0 , \9554_b0 , w_24811 );
and ( w_24810 , w_24811 , \9558_b0 );
or ( \9811_b1 , \9558_b1 , \9560_b1 );
not ( \9560_b1 , w_24812 );
and ( \9811_b0 , \9558_b0 , w_24813 );
and ( w_24812 , w_24813 , \9560_b0 );
or ( \9812_b1 , \9554_b1 , \9560_b1 );
not ( \9560_b1 , w_24814 );
and ( \9812_b0 , \9554_b0 , w_24815 );
and ( w_24814 , w_24815 , \9560_b0 );
or ( \9814_b1 , \9809_b1 , \9813_b1 );
xor ( \9814_b0 , \9809_b0 , w_24816 );
not ( w_24816 , w_24817 );
and ( w_24817 , \9813_b1 , \9813_b0 );
or ( \9815_b1 , \9535_b1 , w_24818 );
or ( \9815_b0 , \9535_b0 , \9549_b0 );
not ( \9549_b0 , w_24819 );
and ( w_24819 , w_24818 , \9549_b1 );
or ( \9816_b1 , \9814_b1 , \9815_b1 );
xor ( \9816_b0 , \9814_b0 , w_24820 );
not ( w_24820 , w_24821 );
and ( w_24821 , \9815_b1 , \9815_b0 );
or ( \9817_b1 , \9805_b1 , \9816_b1 );
xor ( \9817_b0 , \9805_b0 , w_24822 );
not ( w_24822 , w_24823 );
and ( w_24823 , \9816_b1 , \9816_b0 );
or ( \9818_b1 , \9689_b1 , \9817_b1 );
xor ( \9818_b0 , \9689_b0 , w_24824 );
not ( w_24824 , w_24825 );
and ( w_24825 , \9817_b1 , \9817_b0 );
or ( \9819_b1 , \9680_b1 , \9818_b1 );
xor ( \9819_b0 , \9680_b0 , w_24826 );
not ( w_24826 , w_24827 );
and ( w_24827 , \9818_b1 , \9818_b0 );
or ( \9820_b1 , \9502_b1 , \9513_b1 );
not ( \9513_b1 , w_24828 );
and ( \9820_b0 , \9502_b0 , w_24829 );
and ( w_24828 , w_24829 , \9513_b0 );
or ( \9821_b1 , \9513_b1 , \9653_b1 );
not ( \9653_b1 , w_24830 );
and ( \9821_b0 , \9513_b0 , w_24831 );
and ( w_24830 , w_24831 , \9653_b0 );
or ( \9822_b1 , \9502_b1 , \9653_b1 );
not ( \9653_b1 , w_24832 );
and ( \9822_b0 , \9502_b0 , w_24833 );
and ( w_24832 , w_24833 , \9653_b0 );
or ( \9824_b1 , \9819_b1 , w_24835 );
not ( w_24835 , w_24836 );
and ( \9824_b0 , \9819_b0 , w_24837 );
and ( w_24836 ,  , w_24837 );
buf ( w_24835 , \9823_b1 );
not ( w_24835 , w_24838 );
not (  , w_24839 );
and ( w_24838 , w_24839 , \9823_b0 );
or ( \9825_b1 , \9684_b1 , \9688_b1 );
not ( \9688_b1 , w_24840 );
and ( \9825_b0 , \9684_b0 , w_24841 );
and ( w_24840 , w_24841 , \9688_b0 );
or ( \9826_b1 , \9688_b1 , \9817_b1 );
not ( \9817_b1 , w_24842 );
and ( \9826_b0 , \9688_b0 , w_24843 );
and ( w_24842 , w_24843 , \9817_b0 );
or ( \9827_b1 , \9684_b1 , \9817_b1 );
not ( \9817_b1 , w_24844 );
and ( \9827_b0 , \9684_b0 , w_24845 );
and ( w_24844 , w_24845 , \9817_b0 );
or ( \9829_b1 , \9809_b1 , \9813_b1 );
not ( \9813_b1 , w_24846 );
and ( \9829_b0 , \9809_b0 , w_24847 );
and ( w_24846 , w_24847 , \9813_b0 );
or ( \9830_b1 , \9813_b1 , \9815_b1 );
not ( \9815_b1 , w_24848 );
and ( \9830_b0 , \9813_b0 , w_24849 );
and ( w_24848 , w_24849 , \9815_b0 );
or ( \9831_b1 , \9809_b1 , \9815_b1 );
not ( \9815_b1 , w_24850 );
and ( \9831_b0 , \9809_b0 , w_24851 );
and ( w_24850 , w_24851 , \9815_b0 );
or ( \9833_b1 , \9722_b1 , \9763_b1 );
not ( \9763_b1 , w_24852 );
and ( \9833_b0 , \9722_b0 , w_24853 );
and ( w_24852 , w_24853 , \9763_b0 );
or ( \9834_b1 , \9763_b1 , \9803_b1 );
not ( \9803_b1 , w_24854 );
and ( \9834_b0 , \9763_b0 , w_24855 );
and ( w_24854 , w_24855 , \9803_b0 );
or ( \9835_b1 , \9722_b1 , \9803_b1 );
not ( \9803_b1 , w_24856 );
and ( \9835_b0 , \9722_b0 , w_24857 );
and ( w_24856 , w_24857 , \9803_b0 );
or ( \9837_b1 , \9832_b1 , \9836_b1 );
xor ( \9837_b0 , \9832_b0 , w_24858 );
not ( w_24858 , w_24859 );
and ( w_24859 , \9836_b1 , \9836_b0 );
or ( \9838_b1 , \9703_b1 , \9717_b1 );
not ( \9717_b1 , w_24860 );
and ( \9838_b0 , \9703_b0 , w_24861 );
and ( w_24860 , w_24861 , \9717_b0 );
or ( \9839_b1 , \9837_b1 , \9838_b1 );
xor ( \9839_b0 , \9837_b0 , w_24862 );
not ( w_24862 , w_24863 );
and ( w_24863 , \9838_b1 , \9838_b0 );
or ( \9840_b1 , \9828_b1 , \9839_b1 );
xor ( \9840_b0 , \9828_b0 , w_24864 );
not ( w_24864 , w_24865 );
and ( w_24865 , \9839_b1 , \9839_b0 );
or ( \9841_b1 , \9669_b1 , \9673_b1 );
not ( \9673_b1 , w_24866 );
and ( \9841_b0 , \9669_b0 , w_24867 );
and ( w_24866 , w_24867 , \9673_b0 );
or ( \9842_b1 , \9673_b1 , \9678_b1 );
not ( \9678_b1 , w_24868 );
and ( \9842_b0 , \9673_b0 , w_24869 );
and ( w_24868 , w_24869 , \9678_b0 );
or ( \9843_b1 , \9669_b1 , \9678_b1 );
not ( \9678_b1 , w_24870 );
and ( \9843_b0 , \9669_b0 , w_24871 );
and ( w_24870 , w_24871 , \9678_b0 );
or ( \9845_b1 , \9718_b1 , \9804_b1 );
not ( \9804_b1 , w_24872 );
and ( \9845_b0 , \9718_b0 , w_24873 );
and ( w_24872 , w_24873 , \9804_b0 );
or ( \9846_b1 , \9804_b1 , \9816_b1 );
not ( \9816_b1 , w_24874 );
and ( \9846_b0 , \9804_b0 , w_24875 );
and ( w_24874 , w_24875 , \9816_b0 );
or ( \9847_b1 , \9718_b1 , \9816_b1 );
not ( \9816_b1 , w_24876 );
and ( \9847_b0 , \9718_b0 , w_24877 );
and ( w_24876 , w_24877 , \9816_b0 );
or ( \9849_b1 , \9844_b1 , \9848_b1 );
xor ( \9849_b0 , \9844_b0 , w_24878 );
not ( w_24878 , w_24879 );
and ( w_24879 , \9848_b1 , \9848_b0 );
or ( \9850_b1 , \6029_b1 , \5891_b1 );
not ( \5891_b1 , w_24880 );
and ( \9850_b0 , \6029_b0 , w_24881 );
and ( w_24880 , w_24881 , \5891_b0 );
or ( \9851_b1 , \6041_b1 , \5889_b1 );
not ( \5889_b1 , w_24882 );
and ( \9851_b0 , \6041_b0 , w_24883 );
and ( w_24882 , w_24883 , \5889_b0 );
or ( \9852_b1 , \9850_b1 , w_24885 );
not ( w_24885 , w_24886 );
and ( \9852_b0 , \9850_b0 , w_24887 );
and ( w_24886 ,  , w_24887 );
buf ( w_24885 , \9851_b1 );
not ( w_24885 , w_24888 );
not (  , w_24889 );
and ( w_24888 , w_24889 , \9851_b0 );
or ( \9853_b1 , \9852_b1 , w_24890 );
xor ( \9853_b0 , \9852_b0 , w_24892 );
not ( w_24892 , w_24893 );
and ( w_24893 , w_24890 , w_24891 );
buf ( w_24890 , \5898_b1 );
not ( w_24890 , w_24894 );
not ( w_24891 , w_24895 );
and ( w_24894 , w_24895 , \5898_b0 );
or ( \9854_b1 , \6048_b1 , \5916_b1 );
not ( \5916_b1 , w_24896 );
and ( \9854_b0 , \6048_b0 , w_24897 );
and ( w_24896 , w_24897 , \5916_b0 );
or ( \9855_b1 , \6057_b1 , \5914_b1 );
not ( \5914_b1 , w_24898 );
and ( \9855_b0 , \6057_b0 , w_24899 );
and ( w_24898 , w_24899 , \5914_b0 );
or ( \9856_b1 , \9854_b1 , w_24901 );
not ( w_24901 , w_24902 );
and ( \9856_b0 , \9854_b0 , w_24903 );
and ( w_24902 ,  , w_24903 );
buf ( w_24901 , \9855_b1 );
not ( w_24901 , w_24904 );
not (  , w_24905 );
and ( w_24904 , w_24905 , \9855_b0 );
or ( \9857_b1 , \9856_b1 , w_24906 );
xor ( \9857_b0 , \9856_b0 , w_24908 );
not ( w_24908 , w_24909 );
and ( w_24909 , w_24906 , w_24907 );
buf ( w_24906 , \5923_b1 );
not ( w_24906 , w_24910 );
not ( w_24907 , w_24911 );
and ( w_24910 , w_24911 , \5923_b0 );
or ( \9858_b1 , \9853_b1 , \9857_b1 );
xor ( \9858_b0 , \9853_b0 , w_24912 );
not ( w_24912 , w_24913 );
and ( w_24913 , \9857_b1 , \9857_b0 );
or ( \9859_b1 , \6065_b1 , w_24915 );
not ( w_24915 , w_24916 );
and ( \9859_b0 , \6065_b0 , w_24917 );
and ( w_24916 ,  , w_24917 );
buf ( w_24915 , \5933_b1 );
not ( w_24915 , w_24918 );
not (  , w_24919 );
and ( w_24918 , w_24919 , \5933_b0 );
or ( \9860_b1 , \9859_b1 , w_24920 );
xor ( \9860_b0 , \9859_b0 , w_24922 );
not ( w_24922 , w_24923 );
and ( w_24923 , w_24920 , w_24921 );
buf ( w_24920 , \5942_b1 );
not ( w_24920 , w_24924 );
not ( w_24921 , w_24925 );
and ( w_24924 , w_24925 , \5942_b0 );
or ( \9861_b1 , \9858_b1 , \9860_b1 );
xor ( \9861_b0 , \9858_b0 , w_24926 );
not ( w_24926 , w_24927 );
and ( w_24927 , \9860_b1 , \9860_b0 );
or ( \9862_b1 , \5967_b1 , \5829_b1 );
not ( \5829_b1 , w_24928 );
and ( \9862_b0 , \5967_b0 , w_24929 );
and ( w_24928 , w_24929 , \5829_b0 );
or ( \9863_b1 , \5979_b1 , \5827_b1 );
not ( \5827_b1 , w_24930 );
and ( \9863_b0 , \5979_b0 , w_24931 );
and ( w_24930 , w_24931 , \5827_b0 );
or ( \9864_b1 , \9862_b1 , w_24933 );
not ( w_24933 , w_24934 );
and ( \9864_b0 , \9862_b0 , w_24935 );
and ( w_24934 ,  , w_24935 );
buf ( w_24933 , \9863_b1 );
not ( w_24933 , w_24936 );
not (  , w_24937 );
and ( w_24936 , w_24937 , \9863_b0 );
or ( \9865_b1 , \9864_b1 , w_24938 );
xor ( \9865_b0 , \9864_b0 , w_24940 );
not ( w_24940 , w_24941 );
and ( w_24941 , w_24938 , w_24939 );
buf ( w_24938 , \5836_b1 );
not ( w_24938 , w_24942 );
not ( w_24939 , w_24943 );
and ( w_24942 , w_24943 , \5836_b0 );
or ( \9866_b1 , \5986_b1 , \5852_b1 );
not ( \5852_b1 , w_24944 );
and ( \9866_b0 , \5986_b0 , w_24945 );
and ( w_24944 , w_24945 , \5852_b0 );
or ( \9867_b1 , \5998_b1 , \5850_b1 );
not ( \5850_b1 , w_24946 );
and ( \9867_b0 , \5998_b0 , w_24947 );
and ( w_24946 , w_24947 , \5850_b0 );
or ( \9868_b1 , \9866_b1 , w_24949 );
not ( w_24949 , w_24950 );
and ( \9868_b0 , \9866_b0 , w_24951 );
and ( w_24950 ,  , w_24951 );
buf ( w_24949 , \9867_b1 );
not ( w_24949 , w_24952 );
not (  , w_24953 );
and ( w_24952 , w_24953 , \9867_b0 );
or ( \9869_b1 , \9868_b1 , w_24954 );
xor ( \9869_b0 , \9868_b0 , w_24956 );
not ( w_24956 , w_24957 );
and ( w_24957 , w_24954 , w_24955 );
buf ( w_24954 , \5859_b1 );
not ( w_24954 , w_24958 );
not ( w_24955 , w_24959 );
and ( w_24958 , w_24959 , \5859_b0 );
or ( \9870_b1 , \9865_b1 , \9869_b1 );
xor ( \9870_b0 , \9865_b0 , w_24960 );
not ( w_24960 , w_24961 );
and ( w_24961 , \9869_b1 , \9869_b0 );
or ( \9871_b1 , \6006_b1 , \5871_b1 );
not ( \5871_b1 , w_24962 );
and ( \9871_b0 , \6006_b0 , w_24963 );
and ( w_24962 , w_24963 , \5871_b0 );
or ( \9872_b1 , \6018_b1 , \5869_b1 );
not ( \5869_b1 , w_24964 );
and ( \9872_b0 , \6018_b0 , w_24965 );
and ( w_24964 , w_24965 , \5869_b0 );
or ( \9873_b1 , \9871_b1 , w_24967 );
not ( w_24967 , w_24968 );
and ( \9873_b0 , \9871_b0 , w_24969 );
and ( w_24968 ,  , w_24969 );
buf ( w_24967 , \9872_b1 );
not ( w_24967 , w_24970 );
not (  , w_24971 );
and ( w_24970 , w_24971 , \9872_b0 );
or ( \9874_b1 , \9873_b1 , w_24972 );
xor ( \9874_b0 , \9873_b0 , w_24974 );
not ( w_24974 , w_24975 );
and ( w_24975 , w_24972 , w_24973 );
buf ( w_24972 , \5878_b1 );
not ( w_24972 , w_24976 );
not ( w_24973 , w_24977 );
and ( w_24976 , w_24977 , \5878_b0 );
or ( \9875_b1 , \9870_b1 , \9874_b1 );
xor ( \9875_b0 , \9870_b0 , w_24978 );
not ( w_24978 , w_24979 );
and ( w_24979 , \9874_b1 , \9874_b0 );
or ( \9876_b1 , \9861_b1 , w_24980 );
xor ( \9876_b0 , \9861_b0 , w_24982 );
not ( w_24982 , w_24983 );
and ( w_24983 , w_24980 , w_24981 );
buf ( w_24980 , \9875_b1 );
not ( w_24980 , w_24984 );
not ( w_24981 , w_24985 );
and ( w_24984 , w_24985 , \9875_b0 );
or ( \9877_b1 , \9792_b1 , \9796_b1 );
not ( \9796_b1 , w_24986 );
and ( \9877_b0 , \9792_b0 , w_24987 );
and ( w_24986 , w_24987 , \9796_b0 );
or ( \9878_b1 , \9796_b1 , \9801_b1 );
not ( \9801_b1 , w_24988 );
and ( \9878_b0 , \9796_b0 , w_24989 );
and ( w_24988 , w_24989 , \9801_b0 );
or ( \9879_b1 , \9792_b1 , \9801_b1 );
not ( \9801_b1 , w_24990 );
and ( \9879_b0 , \9792_b0 , w_24991 );
and ( w_24990 , w_24991 , \9801_b0 );
or ( \9881_b1 , \9777_b1 , \9781_b1 );
not ( \9781_b1 , w_24992 );
and ( \9881_b0 , \9777_b0 , w_24993 );
and ( w_24992 , w_24993 , \9781_b0 );
or ( \9882_b1 , \9781_b1 , \9786_b1 );
not ( \9786_b1 , w_24994 );
and ( \9882_b0 , \9781_b0 , w_24995 );
and ( w_24994 , w_24995 , \9786_b0 );
or ( \9883_b1 , \9777_b1 , \9786_b1 );
not ( \9786_b1 , w_24996 );
and ( \9883_b0 , \9777_b0 , w_24997 );
and ( w_24996 , w_24997 , \9786_b0 );
or ( \9885_b1 , \9880_b1 , \9884_b1 );
xor ( \9885_b0 , \9880_b0 , w_24998 );
not ( w_24998 , w_24999 );
and ( w_24999 , \9884_b1 , \9884_b0 );
or ( \9886_b1 , \9768_b1 , \9772_b1 );
not ( \9772_b1 , w_25000 );
and ( \9886_b0 , \9768_b0 , w_25001 );
and ( w_25000 , w_25001 , \9772_b0 );
or ( \9887_b1 , \9885_b1 , \9886_b1 );
xor ( \9887_b0 , \9885_b0 , w_25002 );
not ( w_25002 , w_25003 );
and ( w_25003 , \9886_b1 , \9886_b0 );
or ( \9888_b1 , \9876_b1 , \9887_b1 );
xor ( \9888_b0 , \9876_b0 , w_25004 );
not ( w_25004 , w_25005 );
and ( w_25005 , \9887_b1 , \9887_b0 );
or ( \9889_b1 , \9752_b1 , \9756_b1 );
not ( \9756_b1 , w_25006 );
and ( \9889_b0 , \9752_b0 , w_25007 );
and ( w_25006 , w_25007 , \9756_b0 );
or ( \9890_b1 , \9756_b1 , \9761_b1 );
not ( \9761_b1 , w_25008 );
and ( \9890_b0 , \9756_b0 , w_25009 );
and ( w_25008 , w_25009 , \9761_b0 );
or ( \9891_b1 , \9752_b1 , \9761_b1 );
not ( \9761_b1 , w_25010 );
and ( \9891_b0 , \9752_b0 , w_25011 );
and ( w_25010 , w_25011 , \9761_b0 );
or ( \9893_b1 , \9740_b1 , \9744_b1 );
not ( \9744_b1 , w_25012 );
and ( \9893_b0 , \9740_b0 , w_25013 );
and ( w_25012 , w_25013 , \9744_b0 );
or ( \9894_b1 , \9744_b1 , \9749_b1 );
not ( \9749_b1 , w_25014 );
and ( \9894_b0 , \9744_b0 , w_25015 );
and ( w_25014 , w_25015 , \9749_b0 );
or ( \9895_b1 , \9740_b1 , \9749_b1 );
not ( \9749_b1 , w_25016 );
and ( \9895_b0 , \9740_b0 , w_25017 );
and ( w_25016 , w_25017 , \9749_b0 );
or ( \9897_b1 , \9892_b1 , \9896_b1 );
xor ( \9897_b0 , \9892_b0 , w_25018 );
not ( w_25018 , w_25019 );
and ( w_25019 , \9896_b1 , \9896_b0 );
or ( \9898_b1 , \9726_b1 , \9730_b1 );
not ( \9730_b1 , w_25020 );
and ( \9898_b0 , \9726_b0 , w_25021 );
and ( w_25020 , w_25021 , \9730_b0 );
or ( \9899_b1 , \9730_b1 , \9735_b1 );
not ( \9735_b1 , w_25022 );
and ( \9899_b0 , \9730_b0 , w_25023 );
and ( w_25022 , w_25023 , \9735_b0 );
or ( \9900_b1 , \9726_b1 , \9735_b1 );
not ( \9735_b1 , w_25024 );
and ( \9900_b0 , \9726_b0 , w_25025 );
and ( w_25024 , w_25025 , \9735_b0 );
or ( \9902_b1 , \9897_b1 , \9901_b1 );
xor ( \9902_b0 , \9897_b0 , w_25026 );
not ( w_25026 , w_25027 );
and ( w_25027 , \9901_b1 , \9901_b0 );
or ( \9903_b1 , \9888_b1 , \9902_b1 );
xor ( \9903_b0 , \9888_b0 , w_25028 );
not ( w_25028 , w_25029 );
and ( w_25029 , \9902_b1 , \9902_b0 );
or ( \9904_b1 , \9736_b1 , \9750_b1 );
not ( \9750_b1 , w_25030 );
and ( \9904_b0 , \9736_b0 , w_25031 );
and ( w_25030 , w_25031 , \9750_b0 );
or ( \9905_b1 , \9750_b1 , \9762_b1 );
not ( \9762_b1 , w_25032 );
and ( \9905_b0 , \9750_b0 , w_25033 );
and ( w_25032 , w_25033 , \9762_b0 );
or ( \9906_b1 , \9736_b1 , \9762_b1 );
not ( \9762_b1 , w_25034 );
and ( \9906_b0 , \9736_b0 , w_25035 );
and ( w_25034 , w_25035 , \9762_b0 );
or ( \9908_b1 , \5737_b1 , \7099_b1 );
not ( \7099_b1 , w_25036 );
and ( \9908_b0 , \5737_b0 , w_25037 );
and ( w_25036 , w_25037 , \7099_b0 );
buf ( \9909_b1 , \9908_b1 );
not ( \9909_b1 , w_25038 );
not ( \9909_b0 , w_25039 );
and ( w_25038 , w_25039 , \9908_b0 );
or ( \9910_b1 , \9909_b1 , w_25040 );
xor ( \9910_b0 , \9909_b0 , w_25042 );
not ( w_25042 , w_25043 );
and ( w_25043 , w_25040 , w_25041 );
buf ( w_25040 , \7105_b1 );
not ( w_25040 , w_25044 );
not ( w_25041 , w_25045 );
and ( w_25044 , w_25045 , \7105_b0 );
or ( \9911_b1 , \5942_b1 , \9910_b1 );
xor ( \9911_b0 , \5942_b0 , w_25046 );
not ( w_25046 , w_25047 );
and ( w_25047 , \9910_b1 , \9910_b0 );
or ( \9912_b1 , \5758_b1 , \7117_b1 );
not ( \7117_b1 , w_25048 );
and ( \9912_b0 , \5758_b0 , w_25049 );
and ( w_25048 , w_25049 , \7117_b0 );
or ( \9913_b1 , \5770_b1 , \7115_b1 );
not ( \7115_b1 , w_25050 );
and ( \9913_b0 , \5770_b0 , w_25051 );
and ( w_25050 , w_25051 , \7115_b0 );
or ( \9914_b1 , \9912_b1 , w_25053 );
not ( w_25053 , w_25054 );
and ( \9914_b0 , \9912_b0 , w_25055 );
and ( w_25054 ,  , w_25055 );
buf ( w_25053 , \9913_b1 );
not ( w_25053 , w_25056 );
not (  , w_25057 );
and ( w_25056 , w_25057 , \9913_b0 );
or ( \9915_b1 , \9914_b1 , w_25058 );
xor ( \9915_b0 , \9914_b0 , w_25060 );
not ( w_25060 , w_25061 );
and ( w_25061 , w_25058 , w_25059 );
buf ( w_25058 , \7123_b1 );
not ( w_25058 , w_25062 );
not ( w_25059 , w_25063 );
and ( w_25062 , w_25063 , \7123_b0 );
or ( \9916_b1 , \9911_b1 , \9915_b1 );
xor ( \9916_b0 , \9911_b0 , w_25064 );
not ( w_25064 , w_25065 );
and ( w_25065 , \9915_b1 , \9915_b0 );
or ( \9917_b1 , \9907_b1 , \9916_b1 );
xor ( \9917_b0 , \9907_b0 , w_25066 );
not ( w_25066 , w_25067 );
and ( w_25067 , \9916_b1 , \9916_b0 );
or ( \9918_b1 , \5906_b1 , \5768_b1 );
not ( \5768_b1 , w_25068 );
and ( \9918_b0 , \5906_b0 , w_25069 );
and ( w_25068 , w_25069 , \5768_b0 );
or ( \9919_b1 , \5918_b1 , \5766_b1 );
not ( \5766_b1 , w_25070 );
and ( \9919_b0 , \5918_b0 , w_25071 );
and ( w_25070 , w_25071 , \5766_b0 );
or ( \9920_b1 , \9918_b1 , w_25073 );
not ( w_25073 , w_25074 );
and ( \9920_b0 , \9918_b0 , w_25075 );
and ( w_25074 ,  , w_25075 );
buf ( w_25073 , \9919_b1 );
not ( w_25073 , w_25076 );
not (  , w_25077 );
and ( w_25076 , w_25077 , \9919_b0 );
or ( \9921_b1 , \9920_b1 , w_25078 );
xor ( \9921_b0 , \9920_b0 , w_25080 );
not ( w_25080 , w_25081 );
and ( w_25081 , w_25078 , w_25079 );
buf ( w_25078 , \5775_b1 );
not ( w_25078 , w_25082 );
not ( w_25079 , w_25083 );
and ( w_25082 , w_25083 , \5775_b0 );
or ( \9922_b1 , \5925_b1 , \5790_b1 );
not ( \5790_b1 , w_25084 );
and ( \9922_b0 , \5925_b0 , w_25085 );
and ( w_25084 , w_25085 , \5790_b0 );
or ( \9923_b1 , \5937_b1 , \5788_b1 );
not ( \5788_b1 , w_25086 );
and ( \9923_b0 , \5937_b0 , w_25087 );
and ( w_25086 , w_25087 , \5788_b0 );
or ( \9924_b1 , \9922_b1 , w_25089 );
not ( w_25089 , w_25090 );
and ( \9924_b0 , \9922_b0 , w_25091 );
and ( w_25090 ,  , w_25091 );
buf ( w_25089 , \9923_b1 );
not ( w_25089 , w_25092 );
not (  , w_25093 );
and ( w_25092 , w_25093 , \9923_b0 );
or ( \9925_b1 , \9924_b1 , w_25094 );
xor ( \9925_b0 , \9924_b0 , w_25096 );
not ( w_25096 , w_25097 );
and ( w_25097 , w_25094 , w_25095 );
buf ( w_25094 , \5797_b1 );
not ( w_25094 , w_25098 );
not ( w_25095 , w_25099 );
and ( w_25098 , w_25099 , \5797_b0 );
or ( \9926_b1 , \9921_b1 , \9925_b1 );
xor ( \9926_b0 , \9921_b0 , w_25100 );
not ( w_25100 , w_25101 );
and ( w_25101 , \9925_b1 , \9925_b0 );
or ( \9927_b1 , \5945_b1 , \5809_b1 );
not ( \5809_b1 , w_25102 );
and ( \9927_b0 , \5945_b0 , w_25103 );
and ( w_25102 , w_25103 , \5809_b0 );
or ( \9928_b1 , \5957_b1 , \5807_b1 );
not ( \5807_b1 , w_25104 );
and ( \9928_b0 , \5957_b0 , w_25105 );
and ( w_25104 , w_25105 , \5807_b0 );
or ( \9929_b1 , \9927_b1 , w_25107 );
not ( w_25107 , w_25108 );
and ( \9929_b0 , \9927_b0 , w_25109 );
and ( w_25108 ,  , w_25109 );
buf ( w_25107 , \9928_b1 );
not ( w_25107 , w_25110 );
not (  , w_25111 );
and ( w_25110 , w_25111 , \9928_b0 );
or ( \9930_b1 , \9929_b1 , w_25112 );
xor ( \9930_b0 , \9929_b0 , w_25114 );
not ( w_25114 , w_25115 );
and ( w_25115 , w_25112 , w_25113 );
buf ( w_25112 , \5816_b1 );
not ( w_25112 , w_25116 );
not ( w_25113 , w_25117 );
and ( w_25116 , w_25117 , \5816_b0 );
or ( \9931_b1 , \9926_b1 , \9930_b1 );
xor ( \9931_b0 , \9926_b0 , w_25118 );
not ( w_25118 , w_25119 );
and ( w_25119 , \9930_b1 , \9930_b0 );
or ( \9932_b1 , \5842_b1 , \7192_b1 );
not ( \7192_b1 , w_25120 );
and ( \9932_b0 , \5842_b0 , w_25121 );
and ( w_25120 , w_25121 , \7192_b0 );
or ( \9933_b1 , \5854_b1 , \7190_b1 );
not ( \7190_b1 , w_25122 );
and ( \9933_b0 , \5854_b0 , w_25123 );
and ( w_25122 , w_25123 , \7190_b0 );
or ( \9934_b1 , \9932_b1 , w_25125 );
not ( w_25125 , w_25126 );
and ( \9934_b0 , \9932_b0 , w_25127 );
and ( w_25126 ,  , w_25127 );
buf ( w_25125 , \9933_b1 );
not ( w_25125 , w_25128 );
not (  , w_25129 );
and ( w_25128 , w_25129 , \9933_b0 );
or ( \9935_b1 , \9934_b1 , w_25130 );
xor ( \9935_b0 , \9934_b0 , w_25132 );
not ( w_25132 , w_25133 );
and ( w_25133 , w_25130 , w_25131 );
buf ( w_25130 , \7198_b1 );
not ( w_25130 , w_25134 );
not ( w_25131 , w_25135 );
and ( w_25134 , w_25135 , \7198_b0 );
or ( \9936_b1 , \5861_b1 , \7203_b1 );
not ( \7203_b1 , w_25136 );
and ( \9936_b0 , \5861_b0 , w_25137 );
and ( w_25136 , w_25137 , \7203_b0 );
or ( \9937_b1 , \5873_b1 , \7201_b1 );
not ( \7201_b1 , w_25138 );
and ( \9937_b0 , \5873_b0 , w_25139 );
and ( w_25138 , w_25139 , \7201_b0 );
or ( \9938_b1 , \9936_b1 , w_25141 );
not ( w_25141 , w_25142 );
and ( \9938_b0 , \9936_b0 , w_25143 );
and ( w_25142 ,  , w_25143 );
buf ( w_25141 , \9937_b1 );
not ( w_25141 , w_25144 );
not (  , w_25145 );
and ( w_25144 , w_25145 , \9937_b0 );
or ( \9939_b1 , \9938_b1 , w_25146 );
xor ( \9939_b0 , \9938_b0 , w_25148 );
not ( w_25148 , w_25149 );
and ( w_25149 , w_25146 , w_25147 );
buf ( w_25146 , \6824_b1 );
not ( w_25146 , w_25150 );
not ( w_25147 , w_25151 );
and ( w_25150 , w_25151 , \6824_b0 );
or ( \9940_b1 , \9935_b1 , \9939_b1 );
xor ( \9940_b0 , \9935_b0 , w_25152 );
not ( w_25152 , w_25153 );
and ( w_25153 , \9939_b1 , \9939_b0 );
or ( \9941_b1 , \5881_b1 , \5750_b1 );
not ( \5750_b1 , w_25154 );
and ( \9941_b0 , \5881_b0 , w_25155 );
and ( w_25154 , w_25155 , \5750_b0 );
or ( \9942_b1 , \5893_b1 , \5748_b1 );
not ( \5748_b1 , w_25156 );
and ( \9942_b0 , \5893_b0 , w_25157 );
and ( w_25156 , w_25157 , \5748_b0 );
or ( \9943_b1 , \9941_b1 , w_25159 );
not ( w_25159 , w_25160 );
and ( \9943_b0 , \9941_b0 , w_25161 );
and ( w_25160 ,  , w_25161 );
buf ( w_25159 , \9942_b1 );
not ( w_25159 , w_25162 );
not (  , w_25163 );
and ( w_25162 , w_25163 , \9942_b0 );
or ( \9944_b1 , \9943_b1 , w_25164 );
xor ( \9944_b0 , \9943_b0 , w_25166 );
not ( w_25166 , w_25167 );
and ( w_25167 , w_25164 , w_25165 );
buf ( w_25164 , \5755_b1 );
not ( w_25164 , w_25168 );
not ( w_25165 , w_25169 );
and ( w_25168 , w_25169 , \5755_b0 );
or ( \9945_b1 , \9940_b1 , \9944_b1 );
xor ( \9945_b0 , \9940_b0 , w_25170 );
not ( w_25170 , w_25171 );
and ( w_25171 , \9944_b1 , \9944_b0 );
or ( \9946_b1 , \9931_b1 , \9945_b1 );
xor ( \9946_b0 , \9931_b0 , w_25172 );
not ( w_25172 , w_25173 );
and ( w_25173 , \9945_b1 , \9945_b0 );
or ( \9947_b1 , \5780_b1 , \7140_b1 );
not ( \7140_b1 , w_25174 );
and ( \9947_b0 , \5780_b0 , w_25175 );
and ( w_25174 , w_25175 , \7140_b0 );
or ( \9948_b1 , \5792_b1 , \7138_b1 );
not ( \7138_b1 , w_25176 );
and ( \9948_b0 , \5792_b0 , w_25177 );
and ( w_25176 , w_25177 , \7138_b0 );
or ( \9949_b1 , \9947_b1 , w_25179 );
not ( w_25179 , w_25180 );
and ( \9949_b0 , \9947_b0 , w_25181 );
and ( w_25180 ,  , w_25181 );
buf ( w_25179 , \9948_b1 );
not ( w_25179 , w_25182 );
not (  , w_25183 );
and ( w_25182 , w_25183 , \9948_b0 );
or ( \9950_b1 , \9949_b1 , w_25184 );
xor ( \9950_b0 , \9949_b0 , w_25186 );
not ( w_25186 , w_25187 );
and ( w_25187 , w_25184 , w_25185 );
buf ( w_25184 , \7146_b1 );
not ( w_25184 , w_25188 );
not ( w_25185 , w_25189 );
and ( w_25188 , w_25189 , \7146_b0 );
or ( \9951_b1 , \5799_b1 , \7157_b1 );
not ( \7157_b1 , w_25190 );
and ( \9951_b0 , \5799_b0 , w_25191 );
and ( w_25190 , w_25191 , \7157_b0 );
or ( \9952_b1 , \5811_b1 , \7155_b1 );
not ( \7155_b1 , w_25192 );
and ( \9952_b0 , \5811_b0 , w_25193 );
and ( w_25192 , w_25193 , \7155_b0 );
or ( \9953_b1 , \9951_b1 , w_25195 );
not ( w_25195 , w_25196 );
and ( \9953_b0 , \9951_b0 , w_25197 );
and ( w_25196 ,  , w_25197 );
buf ( w_25195 , \9952_b1 );
not ( w_25195 , w_25198 );
not (  , w_25199 );
and ( w_25198 , w_25199 , \9952_b0 );
or ( \9954_b1 , \9953_b1 , w_25200 );
xor ( \9954_b0 , \9953_b0 , w_25202 );
not ( w_25202 , w_25203 );
and ( w_25203 , w_25200 , w_25201 );
buf ( w_25200 , \7163_b1 );
not ( w_25200 , w_25204 );
not ( w_25201 , w_25205 );
and ( w_25204 , w_25205 , \7163_b0 );
or ( \9955_b1 , \9950_b1 , \9954_b1 );
xor ( \9955_b0 , \9950_b0 , w_25206 );
not ( w_25206 , w_25207 );
and ( w_25207 , \9954_b1 , \9954_b0 );
or ( \9956_b1 , \5819_b1 , \7175_b1 );
not ( \7175_b1 , w_25208 );
and ( \9956_b0 , \5819_b0 , w_25209 );
and ( w_25208 , w_25209 , \7175_b0 );
or ( \9957_b1 , \5831_b1 , \7173_b1 );
not ( \7173_b1 , w_25210 );
and ( \9957_b0 , \5831_b0 , w_25211 );
and ( w_25210 , w_25211 , \7173_b0 );
or ( \9958_b1 , \9956_b1 , w_25213 );
not ( w_25213 , w_25214 );
and ( \9958_b0 , \9956_b0 , w_25215 );
and ( w_25214 ,  , w_25215 );
buf ( w_25213 , \9957_b1 );
not ( w_25213 , w_25216 );
not (  , w_25217 );
and ( w_25216 , w_25217 , \9957_b0 );
or ( \9959_b1 , \9958_b1 , w_25218 );
xor ( \9959_b0 , \9958_b0 , w_25220 );
not ( w_25220 , w_25221 );
and ( w_25221 , w_25218 , w_25219 );
buf ( w_25218 , \7181_b1 );
not ( w_25218 , w_25222 );
not ( w_25219 , w_25223 );
and ( w_25222 , w_25223 , \7181_b0 );
or ( \9960_b1 , \9955_b1 , \9959_b1 );
xor ( \9960_b0 , \9955_b0 , w_25224 );
not ( w_25224 , w_25225 );
and ( w_25225 , \9959_b1 , \9959_b0 );
or ( \9961_b1 , \9946_b1 , \9960_b1 );
xor ( \9961_b0 , \9946_b0 , w_25226 );
not ( w_25226 , w_25227 );
and ( w_25227 , \9960_b1 , \9960_b0 );
or ( \9962_b1 , \9917_b1 , \9961_b1 );
xor ( \9962_b0 , \9917_b0 , w_25228 );
not ( w_25228 , w_25229 );
and ( w_25229 , \9961_b1 , \9961_b0 );
or ( \9963_b1 , \9903_b1 , \9962_b1 );
xor ( \9963_b0 , \9903_b0 , w_25230 );
not ( w_25230 , w_25231 );
and ( w_25231 , \9962_b1 , \9962_b0 );
or ( \9964_b1 , \9707_b1 , \9711_b1 );
not ( \9711_b1 , w_25232 );
and ( \9964_b0 , \9707_b0 , w_25233 );
and ( w_25232 , w_25233 , \9711_b0 );
or ( \9965_b1 , \9711_b1 , \9716_b1 );
not ( \9716_b1 , w_25234 );
and ( \9965_b0 , \9711_b0 , w_25235 );
and ( w_25234 , w_25235 , \9716_b0 );
or ( \9966_b1 , \9707_b1 , \9716_b1 );
not ( \9716_b1 , w_25236 );
and ( \9966_b0 , \9707_b0 , w_25237 );
and ( w_25236 , w_25237 , \9716_b0 );
or ( \9968_b1 , \9693_b1 , \9697_b1 );
not ( \9697_b1 , w_25238 );
and ( \9968_b0 , \9693_b0 , w_25239 );
and ( w_25238 , w_25239 , \9697_b0 );
or ( \9969_b1 , \9697_b1 , \9702_b1 );
not ( \9702_b1 , w_25240 );
and ( \9969_b0 , \9697_b0 , w_25241 );
and ( w_25240 , w_25241 , \9702_b0 );
or ( \9970_b1 , \9693_b1 , \9702_b1 );
not ( \9702_b1 , w_25242 );
and ( \9970_b0 , \9693_b0 , w_25243 );
and ( w_25242 , w_25243 , \9702_b0 );
or ( \9972_b1 , \9967_b1 , \9971_b1 );
xor ( \9972_b0 , \9967_b0 , w_25244 );
not ( w_25244 , w_25245 );
and ( w_25245 , \9971_b1 , \9971_b0 );
or ( \9973_b1 , \9773_b1 , \9787_b1 );
not ( \9787_b1 , w_25246 );
and ( \9973_b0 , \9773_b0 , w_25247 );
and ( w_25246 , w_25247 , \9787_b0 );
or ( \9974_b1 , \9787_b1 , \9802_b1 );
not ( \9802_b1 , w_25248 );
and ( \9974_b0 , \9787_b0 , w_25249 );
and ( w_25248 , w_25249 , \9802_b0 );
or ( \9975_b1 , \9773_b1 , \9802_b1 );
not ( \9802_b1 , w_25250 );
and ( \9975_b0 , \9773_b0 , w_25251 );
and ( w_25250 , w_25251 , \9802_b0 );
or ( \9977_b1 , \9972_b1 , \9976_b1 );
xor ( \9977_b0 , \9972_b0 , w_25252 );
not ( w_25252 , w_25253 );
and ( w_25253 , \9976_b1 , \9976_b0 );
or ( \9978_b1 , \9963_b1 , \9977_b1 );
xor ( \9978_b0 , \9963_b0 , w_25254 );
not ( w_25254 , w_25255 );
and ( w_25255 , \9977_b1 , \9977_b0 );
or ( \9979_b1 , \9849_b1 , \9978_b1 );
xor ( \9979_b0 , \9849_b0 , w_25256 );
not ( w_25256 , w_25257 );
and ( w_25257 , \9978_b1 , \9978_b0 );
or ( \9980_b1 , \9840_b1 , \9979_b1 );
xor ( \9980_b0 , \9840_b0 , w_25258 );
not ( w_25258 , w_25259 );
and ( w_25259 , \9979_b1 , \9979_b0 );
or ( \9981_b1 , \9665_b1 , \9679_b1 );
not ( \9679_b1 , w_25260 );
and ( \9981_b0 , \9665_b0 , w_25261 );
and ( w_25260 , w_25261 , \9679_b0 );
or ( \9982_b1 , \9679_b1 , \9818_b1 );
not ( \9818_b1 , w_25262 );
and ( \9982_b0 , \9679_b0 , w_25263 );
and ( w_25262 , w_25263 , \9818_b0 );
or ( \9983_b1 , \9665_b1 , \9818_b1 );
not ( \9818_b1 , w_25264 );
and ( \9983_b0 , \9665_b0 , w_25265 );
and ( w_25264 , w_25265 , \9818_b0 );
or ( \9985_b1 , \9980_b1 , w_25267 );
not ( w_25267 , w_25268 );
and ( \9985_b0 , \9980_b0 , w_25269 );
and ( w_25268 ,  , w_25269 );
buf ( w_25267 , \9984_b1 );
not ( w_25267 , w_25270 );
not (  , w_25271 );
and ( w_25270 , w_25271 , \9984_b0 );
or ( \9986_b1 , \9824_b1 , w_25273 );
not ( w_25273 , w_25274 );
and ( \9986_b0 , \9824_b0 , w_25275 );
and ( w_25274 ,  , w_25275 );
buf ( w_25273 , \9985_b1 );
not ( w_25273 , w_25276 );
not (  , w_25277 );
and ( w_25276 , w_25277 , \9985_b0 );
or ( \9987_b1 , \9844_b1 , \9848_b1 );
not ( \9848_b1 , w_25278 );
and ( \9987_b0 , \9844_b0 , w_25279 );
and ( w_25278 , w_25279 , \9848_b0 );
or ( \9988_b1 , \9848_b1 , \9978_b1 );
not ( \9978_b1 , w_25280 );
and ( \9988_b0 , \9848_b0 , w_25281 );
and ( w_25280 , w_25281 , \9978_b0 );
or ( \9989_b1 , \9844_b1 , \9978_b1 );
not ( \9978_b1 , w_25282 );
and ( \9989_b0 , \9844_b0 , w_25283 );
and ( w_25282 , w_25283 , \9978_b0 );
or ( \9991_b1 , \9967_b1 , \9971_b1 );
not ( \9971_b1 , w_25284 );
and ( \9991_b0 , \9967_b0 , w_25285 );
and ( w_25284 , w_25285 , \9971_b0 );
or ( \9992_b1 , \9971_b1 , \9976_b1 );
not ( \9976_b1 , w_25286 );
and ( \9992_b0 , \9971_b0 , w_25287 );
and ( w_25286 , w_25287 , \9976_b0 );
or ( \9993_b1 , \9967_b1 , \9976_b1 );
not ( \9976_b1 , w_25288 );
and ( \9993_b0 , \9967_b0 , w_25289 );
and ( w_25288 , w_25289 , \9976_b0 );
or ( \9995_b1 , \9907_b1 , \9916_b1 );
not ( \9916_b1 , w_25290 );
and ( \9995_b0 , \9907_b0 , w_25291 );
and ( w_25290 , w_25291 , \9916_b0 );
or ( \9996_b1 , \9916_b1 , \9961_b1 );
not ( \9961_b1 , w_25292 );
and ( \9996_b0 , \9916_b0 , w_25293 );
and ( w_25292 , w_25293 , \9961_b0 );
or ( \9997_b1 , \9907_b1 , \9961_b1 );
not ( \9961_b1 , w_25294 );
and ( \9997_b0 , \9907_b0 , w_25295 );
and ( w_25294 , w_25295 , \9961_b0 );
or ( \9999_b1 , \9994_b1 , \9998_b1 );
xor ( \9999_b0 , \9994_b0 , w_25296 );
not ( w_25296 , w_25297 );
and ( w_25297 , \9998_b1 , \9998_b0 );
or ( \10000_b1 , \9876_b1 , \9887_b1 );
not ( \9887_b1 , w_25298 );
and ( \10000_b0 , \9876_b0 , w_25299 );
and ( w_25298 , w_25299 , \9887_b0 );
or ( \10001_b1 , \9887_b1 , \9902_b1 );
not ( \9902_b1 , w_25300 );
and ( \10001_b0 , \9887_b0 , w_25301 );
and ( w_25300 , w_25301 , \9902_b0 );
or ( \10002_b1 , \9876_b1 , \9902_b1 );
not ( \9902_b1 , w_25302 );
and ( \10002_b0 , \9876_b0 , w_25303 );
and ( w_25302 , w_25303 , \9902_b0 );
or ( \10004_b1 , \9999_b1 , \10003_b1 );
xor ( \10004_b0 , \9999_b0 , w_25304 );
not ( w_25304 , w_25305 );
and ( w_25305 , \10003_b1 , \10003_b0 );
or ( \10005_b1 , \9990_b1 , \10004_b1 );
xor ( \10005_b0 , \9990_b0 , w_25306 );
not ( w_25306 , w_25307 );
and ( w_25307 , \10004_b1 , \10004_b0 );
or ( \10006_b1 , \9832_b1 , \9836_b1 );
not ( \9836_b1 , w_25308 );
and ( \10006_b0 , \9832_b0 , w_25309 );
and ( w_25308 , w_25309 , \9836_b0 );
or ( \10007_b1 , \9836_b1 , \9838_b1 );
not ( \9838_b1 , w_25310 );
and ( \10007_b0 , \9836_b0 , w_25311 );
and ( w_25310 , w_25311 , \9838_b0 );
or ( \10008_b1 , \9832_b1 , \9838_b1 );
not ( \9838_b1 , w_25312 );
and ( \10008_b0 , \9832_b0 , w_25313 );
and ( w_25312 , w_25313 , \9838_b0 );
or ( \10010_b1 , \9903_b1 , \9962_b1 );
not ( \9962_b1 , w_25314 );
and ( \10010_b0 , \9903_b0 , w_25315 );
and ( w_25314 , w_25315 , \9962_b0 );
or ( \10011_b1 , \9962_b1 , \9977_b1 );
not ( \9977_b1 , w_25316 );
and ( \10011_b0 , \9962_b0 , w_25317 );
and ( w_25316 , w_25317 , \9977_b0 );
or ( \10012_b1 , \9903_b1 , \9977_b1 );
not ( \9977_b1 , w_25318 );
and ( \10012_b0 , \9903_b0 , w_25319 );
and ( w_25318 , w_25319 , \9977_b0 );
or ( \10014_b1 , \10009_b1 , \10013_b1 );
xor ( \10014_b0 , \10009_b0 , w_25320 );
not ( w_25320 , w_25321 );
and ( w_25321 , \10013_b1 , \10013_b0 );
or ( \10015_b1 , \9921_b1 , \9925_b1 );
not ( \9925_b1 , w_25322 );
and ( \10015_b0 , \9921_b0 , w_25323 );
and ( w_25322 , w_25323 , \9925_b0 );
or ( \10016_b1 , \9925_b1 , \9930_b1 );
not ( \9930_b1 , w_25324 );
and ( \10016_b0 , \9925_b0 , w_25325 );
and ( w_25324 , w_25325 , \9930_b0 );
or ( \10017_b1 , \9921_b1 , \9930_b1 );
not ( \9930_b1 , w_25326 );
and ( \10017_b0 , \9921_b0 , w_25327 );
and ( w_25326 , w_25327 , \9930_b0 );
or ( \10019_b1 , \9865_b1 , \9869_b1 );
not ( \9869_b1 , w_25328 );
and ( \10019_b0 , \9865_b0 , w_25329 );
and ( w_25328 , w_25329 , \9869_b0 );
or ( \10020_b1 , \9869_b1 , \9874_b1 );
not ( \9874_b1 , w_25330 );
and ( \10020_b0 , \9869_b0 , w_25331 );
and ( w_25330 , w_25331 , \9874_b0 );
or ( \10021_b1 , \9865_b1 , \9874_b1 );
not ( \9874_b1 , w_25332 );
and ( \10021_b0 , \9865_b0 , w_25333 );
and ( w_25332 , w_25333 , \9874_b0 );
or ( \10023_b1 , \10018_b1 , \10022_b1 );
xor ( \10023_b0 , \10018_b0 , w_25334 );
not ( w_25334 , w_25335 );
and ( w_25335 , \10022_b1 , \10022_b0 );
or ( \10024_b1 , \9853_b1 , \9857_b1 );
not ( \9857_b1 , w_25336 );
and ( \10024_b0 , \9853_b0 , w_25337 );
and ( w_25336 , w_25337 , \9857_b0 );
or ( \10025_b1 , \9857_b1 , \9860_b1 );
not ( \9860_b1 , w_25338 );
and ( \10025_b0 , \9857_b0 , w_25339 );
and ( w_25338 , w_25339 , \9860_b0 );
or ( \10026_b1 , \9853_b1 , \9860_b1 );
not ( \9860_b1 , w_25340 );
and ( \10026_b0 , \9853_b0 , w_25341 );
and ( w_25340 , w_25341 , \9860_b0 );
or ( \10028_b1 , \10023_b1 , \10027_b1 );
xor ( \10028_b0 , \10023_b0 , w_25342 );
not ( w_25342 , w_25343 );
and ( w_25343 , \10027_b1 , \10027_b0 );
or ( \10029_b1 , \5942_b1 , \9910_b1 );
not ( \9910_b1 , w_25344 );
and ( \10029_b0 , \5942_b0 , w_25345 );
and ( w_25344 , w_25345 , \9910_b0 );
or ( \10030_b1 , \9910_b1 , \9915_b1 );
not ( \9915_b1 , w_25346 );
and ( \10030_b0 , \9910_b0 , w_25347 );
and ( w_25346 , w_25347 , \9915_b0 );
or ( \10031_b1 , \5942_b1 , \9915_b1 );
not ( \9915_b1 , w_25348 );
and ( \10031_b0 , \5942_b0 , w_25349 );
and ( w_25348 , w_25349 , \9915_b0 );
or ( \10033_b1 , \9950_b1 , \9954_b1 );
not ( \9954_b1 , w_25350 );
and ( \10033_b0 , \9950_b0 , w_25351 );
and ( w_25350 , w_25351 , \9954_b0 );
or ( \10034_b1 , \9954_b1 , \9959_b1 );
not ( \9959_b1 , w_25352 );
and ( \10034_b0 , \9954_b0 , w_25353 );
and ( w_25352 , w_25353 , \9959_b0 );
or ( \10035_b1 , \9950_b1 , \9959_b1 );
not ( \9959_b1 , w_25354 );
and ( \10035_b0 , \9950_b0 , w_25355 );
and ( w_25354 , w_25355 , \9959_b0 );
or ( \10037_b1 , \10032_b1 , \10036_b1 );
xor ( \10037_b0 , \10032_b0 , w_25356 );
not ( w_25356 , w_25357 );
and ( w_25357 , \10036_b1 , \10036_b0 );
or ( \10038_b1 , \9935_b1 , \9939_b1 );
not ( \9939_b1 , w_25358 );
and ( \10038_b0 , \9935_b0 , w_25359 );
and ( w_25358 , w_25359 , \9939_b0 );
or ( \10039_b1 , \9939_b1 , \9944_b1 );
not ( \9944_b1 , w_25360 );
and ( \10039_b0 , \9939_b0 , w_25361 );
and ( w_25360 , w_25361 , \9944_b0 );
or ( \10040_b1 , \9935_b1 , \9944_b1 );
not ( \9944_b1 , w_25362 );
and ( \10040_b0 , \9935_b0 , w_25363 );
and ( w_25362 , w_25363 , \9944_b0 );
or ( \10042_b1 , \10037_b1 , \10041_b1 );
xor ( \10042_b0 , \10037_b0 , w_25364 );
not ( w_25364 , w_25365 );
and ( w_25365 , \10041_b1 , \10041_b0 );
or ( \10043_b1 , \10028_b1 , \10042_b1 );
xor ( \10043_b0 , \10028_b0 , w_25366 );
not ( w_25366 , w_25367 );
and ( w_25367 , \10042_b1 , \10042_b0 );
or ( \10044_b1 , \9931_b1 , \9945_b1 );
not ( \9945_b1 , w_25368 );
and ( \10044_b0 , \9931_b0 , w_25369 );
and ( w_25368 , w_25369 , \9945_b0 );
or ( \10045_b1 , \9945_b1 , \9960_b1 );
not ( \9960_b1 , w_25370 );
and ( \10045_b0 , \9945_b0 , w_25371 );
and ( w_25370 , w_25371 , \9960_b0 );
or ( \10046_b1 , \9931_b1 , \9960_b1 );
not ( \9960_b1 , w_25372 );
and ( \10046_b0 , \9931_b0 , w_25373 );
and ( w_25372 , w_25373 , \9960_b0 );
or ( \10048_b1 , \5873_b1 , \7203_b1 );
not ( \7203_b1 , w_25374 );
and ( \10048_b0 , \5873_b0 , w_25375 );
and ( w_25374 , w_25375 , \7203_b0 );
or ( \10049_b1 , \5842_b1 , \7201_b1 );
not ( \7201_b1 , w_25376 );
and ( \10049_b0 , \5842_b0 , w_25377 );
and ( w_25376 , w_25377 , \7201_b0 );
or ( \10050_b1 , \10048_b1 , w_25379 );
not ( w_25379 , w_25380 );
and ( \10050_b0 , \10048_b0 , w_25381 );
and ( w_25380 ,  , w_25381 );
buf ( w_25379 , \10049_b1 );
not ( w_25379 , w_25382 );
not (  , w_25383 );
and ( w_25382 , w_25383 , \10049_b0 );
or ( \10051_b1 , \10050_b1 , w_25384 );
xor ( \10051_b0 , \10050_b0 , w_25386 );
not ( w_25386 , w_25387 );
and ( w_25387 , w_25384 , w_25385 );
buf ( w_25384 , \6824_b1 );
not ( w_25384 , w_25388 );
not ( w_25385 , w_25389 );
and ( w_25388 , w_25389 , \6824_b0 );
or ( \10052_b1 , \5893_b1 , \5750_b1 );
not ( \5750_b1 , w_25390 );
and ( \10052_b0 , \5893_b0 , w_25391 );
and ( w_25390 , w_25391 , \5750_b0 );
or ( \10053_b1 , \5861_b1 , \5748_b1 );
not ( \5748_b1 , w_25392 );
and ( \10053_b0 , \5861_b0 , w_25393 );
and ( w_25392 , w_25393 , \5748_b0 );
or ( \10054_b1 , \10052_b1 , w_25395 );
not ( w_25395 , w_25396 );
and ( \10054_b0 , \10052_b0 , w_25397 );
and ( w_25396 ,  , w_25397 );
buf ( w_25395 , \10053_b1 );
not ( w_25395 , w_25398 );
not (  , w_25399 );
and ( w_25398 , w_25399 , \10053_b0 );
or ( \10055_b1 , \10054_b1 , w_25400 );
xor ( \10055_b0 , \10054_b0 , w_25402 );
not ( w_25402 , w_25403 );
and ( w_25403 , w_25400 , w_25401 );
buf ( w_25400 , \5755_b1 );
not ( w_25400 , w_25404 );
not ( w_25401 , w_25405 );
and ( w_25404 , w_25405 , \5755_b0 );
or ( \10056_b1 , \10051_b1 , \10055_b1 );
xor ( \10056_b0 , \10051_b0 , w_25406 );
not ( w_25406 , w_25407 );
and ( w_25407 , \10055_b1 , \10055_b0 );
or ( \10057_b1 , \5918_b1 , \5768_b1 );
not ( \5768_b1 , w_25408 );
and ( \10057_b0 , \5918_b0 , w_25409 );
and ( w_25408 , w_25409 , \5768_b0 );
or ( \10058_b1 , \5881_b1 , \5766_b1 );
not ( \5766_b1 , w_25410 );
and ( \10058_b0 , \5881_b0 , w_25411 );
and ( w_25410 , w_25411 , \5766_b0 );
or ( \10059_b1 , \10057_b1 , w_25413 );
not ( w_25413 , w_25414 );
and ( \10059_b0 , \10057_b0 , w_25415 );
and ( w_25414 ,  , w_25415 );
buf ( w_25413 , \10058_b1 );
not ( w_25413 , w_25416 );
not (  , w_25417 );
and ( w_25416 , w_25417 , \10058_b0 );
or ( \10060_b1 , \10059_b1 , w_25418 );
xor ( \10060_b0 , \10059_b0 , w_25420 );
not ( w_25420 , w_25421 );
and ( w_25421 , w_25418 , w_25419 );
buf ( w_25418 , \5775_b1 );
not ( w_25418 , w_25422 );
not ( w_25419 , w_25423 );
and ( w_25422 , w_25423 , \5775_b0 );
or ( \10061_b1 , \10056_b1 , \10060_b1 );
xor ( \10061_b0 , \10056_b0 , w_25424 );
not ( w_25424 , w_25425 );
and ( w_25425 , \10060_b1 , \10060_b0 );
or ( \10062_b1 , \5811_b1 , \7157_b1 );
not ( \7157_b1 , w_25426 );
and ( \10062_b0 , \5811_b0 , w_25427 );
and ( w_25426 , w_25427 , \7157_b0 );
or ( \10063_b1 , \5780_b1 , \7155_b1 );
not ( \7155_b1 , w_25428 );
and ( \10063_b0 , \5780_b0 , w_25429 );
and ( w_25428 , w_25429 , \7155_b0 );
or ( \10064_b1 , \10062_b1 , w_25431 );
not ( w_25431 , w_25432 );
and ( \10064_b0 , \10062_b0 , w_25433 );
and ( w_25432 ,  , w_25433 );
buf ( w_25431 , \10063_b1 );
not ( w_25431 , w_25434 );
not (  , w_25435 );
and ( w_25434 , w_25435 , \10063_b0 );
or ( \10065_b1 , \10064_b1 , w_25436 );
xor ( \10065_b0 , \10064_b0 , w_25438 );
not ( w_25438 , w_25439 );
and ( w_25439 , w_25436 , w_25437 );
buf ( w_25436 , \7163_b1 );
not ( w_25436 , w_25440 );
not ( w_25437 , w_25441 );
and ( w_25440 , w_25441 , \7163_b0 );
or ( \10066_b1 , \5831_b1 , \7175_b1 );
not ( \7175_b1 , w_25442 );
and ( \10066_b0 , \5831_b0 , w_25443 );
and ( w_25442 , w_25443 , \7175_b0 );
or ( \10067_b1 , \5799_b1 , \7173_b1 );
not ( \7173_b1 , w_25444 );
and ( \10067_b0 , \5799_b0 , w_25445 );
and ( w_25444 , w_25445 , \7173_b0 );
or ( \10068_b1 , \10066_b1 , w_25447 );
not ( w_25447 , w_25448 );
and ( \10068_b0 , \10066_b0 , w_25449 );
and ( w_25448 ,  , w_25449 );
buf ( w_25447 , \10067_b1 );
not ( w_25447 , w_25450 );
not (  , w_25451 );
and ( w_25450 , w_25451 , \10067_b0 );
or ( \10069_b1 , \10068_b1 , w_25452 );
xor ( \10069_b0 , \10068_b0 , w_25454 );
not ( w_25454 , w_25455 );
and ( w_25455 , w_25452 , w_25453 );
buf ( w_25452 , \7181_b1 );
not ( w_25452 , w_25456 );
not ( w_25453 , w_25457 );
and ( w_25456 , w_25457 , \7181_b0 );
or ( \10070_b1 , \10065_b1 , \10069_b1 );
xor ( \10070_b0 , \10065_b0 , w_25458 );
not ( w_25458 , w_25459 );
and ( w_25459 , \10069_b1 , \10069_b0 );
or ( \10071_b1 , \5854_b1 , \7192_b1 );
not ( \7192_b1 , w_25460 );
and ( \10071_b0 , \5854_b0 , w_25461 );
and ( w_25460 , w_25461 , \7192_b0 );
or ( \10072_b1 , \5819_b1 , \7190_b1 );
not ( \7190_b1 , w_25462 );
and ( \10072_b0 , \5819_b0 , w_25463 );
and ( w_25462 , w_25463 , \7190_b0 );
or ( \10073_b1 , \10071_b1 , w_25465 );
not ( w_25465 , w_25466 );
and ( \10073_b0 , \10071_b0 , w_25467 );
and ( w_25466 ,  , w_25467 );
buf ( w_25465 , \10072_b1 );
not ( w_25465 , w_25468 );
not (  , w_25469 );
and ( w_25468 , w_25469 , \10072_b0 );
or ( \10074_b1 , \10073_b1 , w_25470 );
xor ( \10074_b0 , \10073_b0 , w_25472 );
not ( w_25472 , w_25473 );
and ( w_25473 , w_25470 , w_25471 );
buf ( w_25470 , \7198_b1 );
not ( w_25470 , w_25474 );
not ( w_25471 , w_25475 );
and ( w_25474 , w_25475 , \7198_b0 );
or ( \10075_b1 , \10070_b1 , \10074_b1 );
xor ( \10075_b0 , \10070_b0 , w_25476 );
not ( w_25476 , w_25477 );
and ( w_25477 , \10074_b1 , \10074_b0 );
or ( \10076_b1 , \10061_b1 , \10075_b1 );
xor ( \10076_b0 , \10061_b0 , w_25478 );
not ( w_25478 , w_25479 );
and ( w_25479 , \10075_b1 , \10075_b0 );
buf ( \10077_b1 , \7105_b1 );
not ( \10077_b1 , w_25480 );
not ( \10077_b0 , w_25481 );
and ( w_25480 , w_25481 , \7105_b0 );
or ( \10078_b1 , \5770_b1 , \7117_b1 );
not ( \7117_b1 , w_25482 );
and ( \10078_b0 , \5770_b0 , w_25483 );
and ( w_25482 , w_25483 , \7117_b0 );
or ( \10079_b1 , \5737_b1 , \7115_b1 );
not ( \7115_b1 , w_25484 );
and ( \10079_b0 , \5737_b0 , w_25485 );
and ( w_25484 , w_25485 , \7115_b0 );
or ( \10080_b1 , \10078_b1 , w_25487 );
not ( w_25487 , w_25488 );
and ( \10080_b0 , \10078_b0 , w_25489 );
and ( w_25488 ,  , w_25489 );
buf ( w_25487 , \10079_b1 );
not ( w_25487 , w_25490 );
not (  , w_25491 );
and ( w_25490 , w_25491 , \10079_b0 );
or ( \10081_b1 , \10080_b1 , w_25492 );
xor ( \10081_b0 , \10080_b0 , w_25494 );
not ( w_25494 , w_25495 );
and ( w_25495 , w_25492 , w_25493 );
buf ( w_25492 , \7123_b1 );
not ( w_25492 , w_25496 );
not ( w_25493 , w_25497 );
and ( w_25496 , w_25497 , \7123_b0 );
or ( \10082_b1 , \10077_b1 , \10081_b1 );
xor ( \10082_b0 , \10077_b0 , w_25498 );
not ( w_25498 , w_25499 );
and ( w_25499 , \10081_b1 , \10081_b0 );
or ( \10083_b1 , \5792_b1 , \7140_b1 );
not ( \7140_b1 , w_25500 );
and ( \10083_b0 , \5792_b0 , w_25501 );
and ( w_25500 , w_25501 , \7140_b0 );
or ( \10084_b1 , \5758_b1 , \7138_b1 );
not ( \7138_b1 , w_25502 );
and ( \10084_b0 , \5758_b0 , w_25503 );
and ( w_25502 , w_25503 , \7138_b0 );
or ( \10085_b1 , \10083_b1 , w_25505 );
not ( w_25505 , w_25506 );
and ( \10085_b0 , \10083_b0 , w_25507 );
and ( w_25506 ,  , w_25507 );
buf ( w_25505 , \10084_b1 );
not ( w_25505 , w_25508 );
not (  , w_25509 );
and ( w_25508 , w_25509 , \10084_b0 );
or ( \10086_b1 , \10085_b1 , w_25510 );
xor ( \10086_b0 , \10085_b0 , w_25512 );
not ( w_25512 , w_25513 );
and ( w_25513 , w_25510 , w_25511 );
buf ( w_25510 , \7146_b1 );
not ( w_25510 , w_25514 );
not ( w_25511 , w_25515 );
and ( w_25514 , w_25515 , \7146_b0 );
or ( \10087_b1 , \10082_b1 , \10086_b1 );
xor ( \10087_b0 , \10082_b0 , w_25516 );
not ( w_25516 , w_25517 );
and ( w_25517 , \10086_b1 , \10086_b0 );
or ( \10088_b1 , \10076_b1 , \10087_b1 );
xor ( \10088_b0 , \10076_b0 , w_25518 );
not ( w_25518 , w_25519 );
and ( w_25519 , \10087_b1 , \10087_b0 );
or ( \10089_b1 , \10047_b1 , \10088_b1 );
xor ( \10089_b0 , \10047_b0 , w_25520 );
not ( w_25520 , w_25521 );
and ( w_25521 , \10088_b1 , \10088_b0 );
or ( \10090_b1 , \6057_b1 , \5916_b1 );
not ( \5916_b1 , w_25522 );
and ( \10090_b0 , \6057_b0 , w_25523 );
and ( w_25522 , w_25523 , \5916_b0 );
or ( \10091_b1 , \6029_b1 , \5914_b1 );
not ( \5914_b1 , w_25524 );
and ( \10091_b0 , \6029_b0 , w_25525 );
and ( w_25524 , w_25525 , \5914_b0 );
or ( \10092_b1 , \10090_b1 , w_25527 );
not ( w_25527 , w_25528 );
and ( \10092_b0 , \10090_b0 , w_25529 );
and ( w_25528 ,  , w_25529 );
buf ( w_25527 , \10091_b1 );
not ( w_25527 , w_25530 );
not (  , w_25531 );
and ( w_25530 , w_25531 , \10091_b0 );
or ( \10093_b1 , \10092_b1 , w_25532 );
xor ( \10093_b0 , \10092_b0 , w_25534 );
not ( w_25534 , w_25535 );
and ( w_25535 , w_25532 , w_25533 );
buf ( w_25532 , \5923_b1 );
not ( w_25532 , w_25536 );
not ( w_25533 , w_25537 );
and ( w_25536 , w_25537 , \5923_b0 );
or ( \10094_b1 , \6065_b1 , \5935_b1 );
not ( \5935_b1 , w_25538 );
and ( \10094_b0 , \6065_b0 , w_25539 );
and ( w_25538 , w_25539 , \5935_b0 );
or ( \10095_b1 , \6048_b1 , \5933_b1 );
not ( \5933_b1 , w_25540 );
and ( \10095_b0 , \6048_b0 , w_25541 );
and ( w_25540 , w_25541 , \5933_b0 );
or ( \10096_b1 , \10094_b1 , w_25543 );
not ( w_25543 , w_25544 );
and ( \10096_b0 , \10094_b0 , w_25545 );
and ( w_25544 ,  , w_25545 );
buf ( w_25543 , \10095_b1 );
not ( w_25543 , w_25546 );
not (  , w_25547 );
and ( w_25546 , w_25547 , \10095_b0 );
or ( \10097_b1 , \10096_b1 , w_25548 );
xor ( \10097_b0 , \10096_b0 , w_25550 );
not ( w_25550 , w_25551 );
and ( w_25551 , w_25548 , w_25549 );
buf ( w_25548 , \5942_b1 );
not ( w_25548 , w_25552 );
not ( w_25549 , w_25553 );
and ( w_25552 , w_25553 , \5942_b0 );
or ( \10098_b1 , \10093_b1 , \10097_b1 );
xor ( \10098_b0 , \10093_b0 , w_25554 );
not ( w_25554 , w_25555 );
and ( w_25555 , \10097_b1 , \10097_b0 );
or ( \10099_b1 , \5998_b1 , \5852_b1 );
not ( \5852_b1 , w_25556 );
and ( \10099_b0 , \5998_b0 , w_25557 );
and ( w_25556 , w_25557 , \5852_b0 );
or ( \10100_b1 , \5967_b1 , \5850_b1 );
not ( \5850_b1 , w_25558 );
and ( \10100_b0 , \5967_b0 , w_25559 );
and ( w_25558 , w_25559 , \5850_b0 );
or ( \10101_b1 , \10099_b1 , w_25561 );
not ( w_25561 , w_25562 );
and ( \10101_b0 , \10099_b0 , w_25563 );
and ( w_25562 ,  , w_25563 );
buf ( w_25561 , \10100_b1 );
not ( w_25561 , w_25564 );
not (  , w_25565 );
and ( w_25564 , w_25565 , \10100_b0 );
or ( \10102_b1 , \10101_b1 , w_25566 );
xor ( \10102_b0 , \10101_b0 , w_25568 );
not ( w_25568 , w_25569 );
and ( w_25569 , w_25566 , w_25567 );
buf ( w_25566 , \5859_b1 );
not ( w_25566 , w_25570 );
not ( w_25567 , w_25571 );
and ( w_25570 , w_25571 , \5859_b0 );
or ( \10103_b1 , \6018_b1 , \5871_b1 );
not ( \5871_b1 , w_25572 );
and ( \10103_b0 , \6018_b0 , w_25573 );
and ( w_25572 , w_25573 , \5871_b0 );
or ( \10104_b1 , \5986_b1 , \5869_b1 );
not ( \5869_b1 , w_25574 );
and ( \10104_b0 , \5986_b0 , w_25575 );
and ( w_25574 , w_25575 , \5869_b0 );
or ( \10105_b1 , \10103_b1 , w_25577 );
not ( w_25577 , w_25578 );
and ( \10105_b0 , \10103_b0 , w_25579 );
and ( w_25578 ,  , w_25579 );
buf ( w_25577 , \10104_b1 );
not ( w_25577 , w_25580 );
not (  , w_25581 );
and ( w_25580 , w_25581 , \10104_b0 );
or ( \10106_b1 , \10105_b1 , w_25582 );
xor ( \10106_b0 , \10105_b0 , w_25584 );
not ( w_25584 , w_25585 );
and ( w_25585 , w_25582 , w_25583 );
buf ( w_25582 , \5878_b1 );
not ( w_25582 , w_25586 );
not ( w_25583 , w_25587 );
and ( w_25586 , w_25587 , \5878_b0 );
or ( \10107_b1 , \10102_b1 , \10106_b1 );
xor ( \10107_b0 , \10102_b0 , w_25588 );
not ( w_25588 , w_25589 );
and ( w_25589 , \10106_b1 , \10106_b0 );
or ( \10108_b1 , \6041_b1 , \5891_b1 );
not ( \5891_b1 , w_25590 );
and ( \10108_b0 , \6041_b0 , w_25591 );
and ( w_25590 , w_25591 , \5891_b0 );
or ( \10109_b1 , \6006_b1 , \5889_b1 );
not ( \5889_b1 , w_25592 );
and ( \10109_b0 , \6006_b0 , w_25593 );
and ( w_25592 , w_25593 , \5889_b0 );
or ( \10110_b1 , \10108_b1 , w_25595 );
not ( w_25595 , w_25596 );
and ( \10110_b0 , \10108_b0 , w_25597 );
and ( w_25596 ,  , w_25597 );
buf ( w_25595 , \10109_b1 );
not ( w_25595 , w_25598 );
not (  , w_25599 );
and ( w_25598 , w_25599 , \10109_b0 );
or ( \10111_b1 , \10110_b1 , w_25600 );
xor ( \10111_b0 , \10110_b0 , w_25602 );
not ( w_25602 , w_25603 );
and ( w_25603 , w_25600 , w_25601 );
buf ( w_25600 , \5898_b1 );
not ( w_25600 , w_25604 );
not ( w_25601 , w_25605 );
and ( w_25604 , w_25605 , \5898_b0 );
or ( \10112_b1 , \10107_b1 , \10111_b1 );
xor ( \10112_b0 , \10107_b0 , w_25606 );
not ( w_25606 , w_25607 );
and ( w_25607 , \10111_b1 , \10111_b0 );
or ( \10113_b1 , \10098_b1 , \10112_b1 );
xor ( \10113_b0 , \10098_b0 , w_25608 );
not ( w_25608 , w_25609 );
and ( w_25609 , \10112_b1 , \10112_b0 );
or ( \10114_b1 , \5937_b1 , \5790_b1 );
not ( \5790_b1 , w_25610 );
and ( \10114_b0 , \5937_b0 , w_25611 );
and ( w_25610 , w_25611 , \5790_b0 );
or ( \10115_b1 , \5906_b1 , \5788_b1 );
not ( \5788_b1 , w_25612 );
and ( \10115_b0 , \5906_b0 , w_25613 );
and ( w_25612 , w_25613 , \5788_b0 );
or ( \10116_b1 , \10114_b1 , w_25615 );
not ( w_25615 , w_25616 );
and ( \10116_b0 , \10114_b0 , w_25617 );
and ( w_25616 ,  , w_25617 );
buf ( w_25615 , \10115_b1 );
not ( w_25615 , w_25618 );
not (  , w_25619 );
and ( w_25618 , w_25619 , \10115_b0 );
or ( \10117_b1 , \10116_b1 , w_25620 );
xor ( \10117_b0 , \10116_b0 , w_25622 );
not ( w_25622 , w_25623 );
and ( w_25623 , w_25620 , w_25621 );
buf ( w_25620 , \5797_b1 );
not ( w_25620 , w_25624 );
not ( w_25621 , w_25625 );
and ( w_25624 , w_25625 , \5797_b0 );
or ( \10118_b1 , \5957_b1 , \5809_b1 );
not ( \5809_b1 , w_25626 );
and ( \10118_b0 , \5957_b0 , w_25627 );
and ( w_25626 , w_25627 , \5809_b0 );
or ( \10119_b1 , \5925_b1 , \5807_b1 );
not ( \5807_b1 , w_25628 );
and ( \10119_b0 , \5925_b0 , w_25629 );
and ( w_25628 , w_25629 , \5807_b0 );
or ( \10120_b1 , \10118_b1 , w_25631 );
not ( w_25631 , w_25632 );
and ( \10120_b0 , \10118_b0 , w_25633 );
and ( w_25632 ,  , w_25633 );
buf ( w_25631 , \10119_b1 );
not ( w_25631 , w_25634 );
not (  , w_25635 );
and ( w_25634 , w_25635 , \10119_b0 );
or ( \10121_b1 , \10120_b1 , w_25636 );
xor ( \10121_b0 , \10120_b0 , w_25638 );
not ( w_25638 , w_25639 );
and ( w_25639 , w_25636 , w_25637 );
buf ( w_25636 , \5816_b1 );
not ( w_25636 , w_25640 );
not ( w_25637 , w_25641 );
and ( w_25640 , w_25641 , \5816_b0 );
or ( \10122_b1 , \10117_b1 , \10121_b1 );
xor ( \10122_b0 , \10117_b0 , w_25642 );
not ( w_25642 , w_25643 );
and ( w_25643 , \10121_b1 , \10121_b0 );
or ( \10123_b1 , \5979_b1 , \5829_b1 );
not ( \5829_b1 , w_25644 );
and ( \10123_b0 , \5979_b0 , w_25645 );
and ( w_25644 , w_25645 , \5829_b0 );
or ( \10124_b1 , \5945_b1 , \5827_b1 );
not ( \5827_b1 , w_25646 );
and ( \10124_b0 , \5945_b0 , w_25647 );
and ( w_25646 , w_25647 , \5827_b0 );
or ( \10125_b1 , \10123_b1 , w_25649 );
not ( w_25649 , w_25650 );
and ( \10125_b0 , \10123_b0 , w_25651 );
and ( w_25650 ,  , w_25651 );
buf ( w_25649 , \10124_b1 );
not ( w_25649 , w_25652 );
not (  , w_25653 );
and ( w_25652 , w_25653 , \10124_b0 );
or ( \10126_b1 , \10125_b1 , w_25654 );
xor ( \10126_b0 , \10125_b0 , w_25656 );
not ( w_25656 , w_25657 );
and ( w_25657 , w_25654 , w_25655 );
buf ( w_25654 , \5836_b1 );
not ( w_25654 , w_25658 );
not ( w_25655 , w_25659 );
and ( w_25658 , w_25659 , \5836_b0 );
or ( \10127_b1 , \10122_b1 , \10126_b1 );
xor ( \10127_b0 , \10122_b0 , w_25660 );
not ( w_25660 , w_25661 );
and ( w_25661 , \10126_b1 , \10126_b0 );
or ( \10128_b1 , \10113_b1 , \10127_b1 );
xor ( \10128_b0 , \10113_b0 , w_25662 );
not ( w_25662 , w_25663 );
and ( w_25663 , \10127_b1 , \10127_b0 );
or ( \10129_b1 , \10089_b1 , \10128_b1 );
xor ( \10129_b0 , \10089_b0 , w_25664 );
not ( w_25664 , w_25665 );
and ( w_25665 , \10128_b1 , \10128_b0 );
or ( \10130_b1 , \10043_b1 , \10129_b1 );
xor ( \10130_b0 , \10043_b0 , w_25666 );
not ( w_25666 , w_25667 );
and ( w_25667 , \10129_b1 , \10129_b0 );
or ( \10131_b1 , \9892_b1 , \9896_b1 );
not ( \9896_b1 , w_25668 );
and ( \10131_b0 , \9892_b0 , w_25669 );
and ( w_25668 , w_25669 , \9896_b0 );
or ( \10132_b1 , \9896_b1 , \9901_b1 );
not ( \9901_b1 , w_25670 );
and ( \10132_b0 , \9896_b0 , w_25671 );
and ( w_25670 , w_25671 , \9901_b0 );
or ( \10133_b1 , \9892_b1 , \9901_b1 );
not ( \9901_b1 , w_25672 );
and ( \10133_b0 , \9892_b0 , w_25673 );
and ( w_25672 , w_25673 , \9901_b0 );
or ( \10135_b1 , \9880_b1 , \9884_b1 );
not ( \9884_b1 , w_25674 );
and ( \10135_b0 , \9880_b0 , w_25675 );
and ( w_25674 , w_25675 , \9884_b0 );
or ( \10136_b1 , \9884_b1 , \9886_b1 );
not ( \9886_b1 , w_25676 );
and ( \10136_b0 , \9884_b0 , w_25677 );
and ( w_25676 , w_25677 , \9886_b0 );
or ( \10137_b1 , \9880_b1 , \9886_b1 );
not ( \9886_b1 , w_25678 );
and ( \10137_b0 , \9880_b0 , w_25679 );
and ( w_25678 , w_25679 , \9886_b0 );
or ( \10139_b1 , \10134_b1 , \10138_b1 );
xor ( \10139_b0 , \10134_b0 , w_25680 );
not ( w_25680 , w_25681 );
and ( w_25681 , \10138_b1 , \10138_b0 );
or ( \10140_b1 , \9861_b1 , w_25682 );
or ( \10140_b0 , \9861_b0 , \9875_b0 );
not ( \9875_b0 , w_25683 );
and ( w_25683 , w_25682 , \9875_b1 );
or ( \10141_b1 , \10139_b1 , \10140_b1 );
xor ( \10141_b0 , \10139_b0 , w_25684 );
not ( w_25684 , w_25685 );
and ( w_25685 , \10140_b1 , \10140_b0 );
or ( \10142_b1 , \10130_b1 , \10141_b1 );
xor ( \10142_b0 , \10130_b0 , w_25686 );
not ( w_25686 , w_25687 );
and ( w_25687 , \10141_b1 , \10141_b0 );
or ( \10143_b1 , \10014_b1 , \10142_b1 );
xor ( \10143_b0 , \10014_b0 , w_25688 );
not ( w_25688 , w_25689 );
and ( w_25689 , \10142_b1 , \10142_b0 );
or ( \10144_b1 , \10005_b1 , \10143_b1 );
xor ( \10144_b0 , \10005_b0 , w_25690 );
not ( w_25690 , w_25691 );
and ( w_25691 , \10143_b1 , \10143_b0 );
or ( \10145_b1 , \9828_b1 , \9839_b1 );
not ( \9839_b1 , w_25692 );
and ( \10145_b0 , \9828_b0 , w_25693 );
and ( w_25692 , w_25693 , \9839_b0 );
or ( \10146_b1 , \9839_b1 , \9979_b1 );
not ( \9979_b1 , w_25694 );
and ( \10146_b0 , \9839_b0 , w_25695 );
and ( w_25694 , w_25695 , \9979_b0 );
or ( \10147_b1 , \9828_b1 , \9979_b1 );
not ( \9979_b1 , w_25696 );
and ( \10147_b0 , \9828_b0 , w_25697 );
and ( w_25696 , w_25697 , \9979_b0 );
or ( \10149_b1 , \10144_b1 , w_25699 );
not ( w_25699 , w_25700 );
and ( \10149_b0 , \10144_b0 , w_25701 );
and ( w_25700 ,  , w_25701 );
buf ( w_25699 , \10148_b1 );
not ( w_25699 , w_25702 );
not (  , w_25703 );
and ( w_25702 , w_25703 , \10148_b0 );
or ( \10150_b1 , \10009_b1 , \10013_b1 );
not ( \10013_b1 , w_25704 );
and ( \10150_b0 , \10009_b0 , w_25705 );
and ( w_25704 , w_25705 , \10013_b0 );
or ( \10151_b1 , \10013_b1 , \10142_b1 );
not ( \10142_b1 , w_25706 );
and ( \10151_b0 , \10013_b0 , w_25707 );
and ( w_25706 , w_25707 , \10142_b0 );
or ( \10152_b1 , \10009_b1 , \10142_b1 );
not ( \10142_b1 , w_25708 );
and ( \10152_b0 , \10009_b0 , w_25709 );
and ( w_25708 , w_25709 , \10142_b0 );
or ( \10154_b1 , \10134_b1 , \10138_b1 );
not ( \10138_b1 , w_25710 );
and ( \10154_b0 , \10134_b0 , w_25711 );
and ( w_25710 , w_25711 , \10138_b0 );
or ( \10155_b1 , \10138_b1 , \10140_b1 );
not ( \10140_b1 , w_25712 );
and ( \10155_b0 , \10138_b0 , w_25713 );
and ( w_25712 , w_25713 , \10140_b0 );
or ( \10156_b1 , \10134_b1 , \10140_b1 );
not ( \10140_b1 , w_25714 );
and ( \10156_b0 , \10134_b0 , w_25715 );
and ( w_25714 , w_25715 , \10140_b0 );
or ( \10158_b1 , \10047_b1 , \10088_b1 );
not ( \10088_b1 , w_25716 );
and ( \10158_b0 , \10047_b0 , w_25717 );
and ( w_25716 , w_25717 , \10088_b0 );
or ( \10159_b1 , \10088_b1 , \10128_b1 );
not ( \10128_b1 , w_25718 );
and ( \10159_b0 , \10088_b0 , w_25719 );
and ( w_25718 , w_25719 , \10128_b0 );
or ( \10160_b1 , \10047_b1 , \10128_b1 );
not ( \10128_b1 , w_25720 );
and ( \10160_b0 , \10047_b0 , w_25721 );
and ( w_25720 , w_25721 , \10128_b0 );
or ( \10162_b1 , \10157_b1 , \10161_b1 );
xor ( \10162_b0 , \10157_b0 , w_25722 );
not ( w_25722 , w_25723 );
and ( w_25723 , \10161_b1 , \10161_b0 );
or ( \10163_b1 , \10028_b1 , \10042_b1 );
not ( \10042_b1 , w_25724 );
and ( \10163_b0 , \10028_b0 , w_25725 );
and ( w_25724 , w_25725 , \10042_b0 );
or ( \10164_b1 , \10162_b1 , \10163_b1 );
xor ( \10164_b0 , \10162_b0 , w_25726 );
not ( w_25726 , w_25727 );
and ( w_25727 , \10163_b1 , \10163_b0 );
or ( \10165_b1 , \10153_b1 , \10164_b1 );
xor ( \10165_b0 , \10153_b0 , w_25728 );
not ( w_25728 , w_25729 );
and ( w_25729 , \10164_b1 , \10164_b0 );
or ( \10166_b1 , \9994_b1 , \9998_b1 );
not ( \9998_b1 , w_25730 );
and ( \10166_b0 , \9994_b0 , w_25731 );
and ( w_25730 , w_25731 , \9998_b0 );
or ( \10167_b1 , \9998_b1 , \10003_b1 );
not ( \10003_b1 , w_25732 );
and ( \10167_b0 , \9998_b0 , w_25733 );
and ( w_25732 , w_25733 , \10003_b0 );
or ( \10168_b1 , \9994_b1 , \10003_b1 );
not ( \10003_b1 , w_25734 );
and ( \10168_b0 , \9994_b0 , w_25735 );
and ( w_25734 , w_25735 , \10003_b0 );
or ( \10170_b1 , \10043_b1 , \10129_b1 );
not ( \10129_b1 , w_25736 );
and ( \10170_b0 , \10043_b0 , w_25737 );
and ( w_25736 , w_25737 , \10129_b0 );
or ( \10171_b1 , \10129_b1 , \10141_b1 );
not ( \10141_b1 , w_25738 );
and ( \10171_b0 , \10129_b0 , w_25739 );
and ( w_25738 , w_25739 , \10141_b0 );
or ( \10172_b1 , \10043_b1 , \10141_b1 );
not ( \10141_b1 , w_25740 );
and ( \10172_b0 , \10043_b0 , w_25741 );
and ( w_25740 , w_25741 , \10141_b0 );
or ( \10174_b1 , \10169_b1 , \10173_b1 );
xor ( \10174_b0 , \10169_b0 , w_25742 );
not ( w_25742 , w_25743 );
and ( w_25743 , \10173_b1 , \10173_b0 );
or ( \10175_b1 , \6029_b1 , \5916_b1 );
not ( \5916_b1 , w_25744 );
and ( \10175_b0 , \6029_b0 , w_25745 );
and ( w_25744 , w_25745 , \5916_b0 );
or ( \10176_b1 , \6041_b1 , \5914_b1 );
not ( \5914_b1 , w_25746 );
and ( \10176_b0 , \6041_b0 , w_25747 );
and ( w_25746 , w_25747 , \5914_b0 );
or ( \10177_b1 , \10175_b1 , w_25749 );
not ( w_25749 , w_25750 );
and ( \10177_b0 , \10175_b0 , w_25751 );
and ( w_25750 ,  , w_25751 );
buf ( w_25749 , \10176_b1 );
not ( w_25749 , w_25752 );
not (  , w_25753 );
and ( w_25752 , w_25753 , \10176_b0 );
or ( \10178_b1 , \10177_b1 , w_25754 );
xor ( \10178_b0 , \10177_b0 , w_25756 );
not ( w_25756 , w_25757 );
and ( w_25757 , w_25754 , w_25755 );
buf ( w_25754 , \5923_b1 );
not ( w_25754 , w_25758 );
not ( w_25755 , w_25759 );
and ( w_25758 , w_25759 , \5923_b0 );
or ( \10179_b1 , \6048_b1 , \5935_b1 );
not ( \5935_b1 , w_25760 );
and ( \10179_b0 , \6048_b0 , w_25761 );
and ( w_25760 , w_25761 , \5935_b0 );
or ( \10180_b1 , \6057_b1 , \5933_b1 );
not ( \5933_b1 , w_25762 );
and ( \10180_b0 , \6057_b0 , w_25763 );
and ( w_25762 , w_25763 , \5933_b0 );
or ( \10181_b1 , \10179_b1 , w_25765 );
not ( w_25765 , w_25766 );
and ( \10181_b0 , \10179_b0 , w_25767 );
and ( w_25766 ,  , w_25767 );
buf ( w_25765 , \10180_b1 );
not ( w_25765 , w_25768 );
not (  , w_25769 );
and ( w_25768 , w_25769 , \10180_b0 );
or ( \10182_b1 , \10181_b1 , w_25770 );
xor ( \10182_b0 , \10181_b0 , w_25772 );
not ( w_25772 , w_25773 );
and ( w_25773 , w_25770 , w_25771 );
buf ( w_25770 , \5942_b1 );
not ( w_25770 , w_25774 );
not ( w_25771 , w_25775 );
and ( w_25774 , w_25775 , \5942_b0 );
or ( \10183_b1 , \10178_b1 , \10182_b1 );
xor ( \10183_b0 , \10178_b0 , w_25776 );
not ( w_25776 , w_25777 );
and ( w_25777 , \10182_b1 , \10182_b0 );
or ( \10184_b1 , \6065_b1 , w_25779 );
not ( w_25779 , w_25780 );
and ( \10184_b0 , \6065_b0 , w_25781 );
and ( w_25780 ,  , w_25781 );
buf ( w_25779 , \5953_b1 );
not ( w_25779 , w_25782 );
not (  , w_25783 );
and ( w_25782 , w_25783 , \5953_b0 );
or ( \10185_b1 , \10184_b1 , w_25784 );
xor ( \10185_b0 , \10184_b0 , w_25786 );
not ( w_25786 , w_25787 );
and ( w_25787 , w_25784 , w_25785 );
buf ( w_25784 , \5962_b1 );
not ( w_25784 , w_25788 );
not ( w_25785 , w_25789 );
and ( w_25788 , w_25789 , \5962_b0 );
or ( \10186_b1 , \10183_b1 , \10185_b1 );
xor ( \10186_b0 , \10183_b0 , w_25790 );
not ( w_25790 , w_25791 );
and ( w_25791 , \10185_b1 , \10185_b0 );
or ( \10187_b1 , \5967_b1 , \5852_b1 );
not ( \5852_b1 , w_25792 );
and ( \10187_b0 , \5967_b0 , w_25793 );
and ( w_25792 , w_25793 , \5852_b0 );
or ( \10188_b1 , \5979_b1 , \5850_b1 );
not ( \5850_b1 , w_25794 );
and ( \10188_b0 , \5979_b0 , w_25795 );
and ( w_25794 , w_25795 , \5850_b0 );
or ( \10189_b1 , \10187_b1 , w_25797 );
not ( w_25797 , w_25798 );
and ( \10189_b0 , \10187_b0 , w_25799 );
and ( w_25798 ,  , w_25799 );
buf ( w_25797 , \10188_b1 );
not ( w_25797 , w_25800 );
not (  , w_25801 );
and ( w_25800 , w_25801 , \10188_b0 );
or ( \10190_b1 , \10189_b1 , w_25802 );
xor ( \10190_b0 , \10189_b0 , w_25804 );
not ( w_25804 , w_25805 );
and ( w_25805 , w_25802 , w_25803 );
buf ( w_25802 , \5859_b1 );
not ( w_25802 , w_25806 );
not ( w_25803 , w_25807 );
and ( w_25806 , w_25807 , \5859_b0 );
or ( \10191_b1 , \5986_b1 , \5871_b1 );
not ( \5871_b1 , w_25808 );
and ( \10191_b0 , \5986_b0 , w_25809 );
and ( w_25808 , w_25809 , \5871_b0 );
or ( \10192_b1 , \5998_b1 , \5869_b1 );
not ( \5869_b1 , w_25810 );
and ( \10192_b0 , \5998_b0 , w_25811 );
and ( w_25810 , w_25811 , \5869_b0 );
or ( \10193_b1 , \10191_b1 , w_25813 );
not ( w_25813 , w_25814 );
and ( \10193_b0 , \10191_b0 , w_25815 );
and ( w_25814 ,  , w_25815 );
buf ( w_25813 , \10192_b1 );
not ( w_25813 , w_25816 );
not (  , w_25817 );
and ( w_25816 , w_25817 , \10192_b0 );
or ( \10194_b1 , \10193_b1 , w_25818 );
xor ( \10194_b0 , \10193_b0 , w_25820 );
not ( w_25820 , w_25821 );
and ( w_25821 , w_25818 , w_25819 );
buf ( w_25818 , \5878_b1 );
not ( w_25818 , w_25822 );
not ( w_25819 , w_25823 );
and ( w_25822 , w_25823 , \5878_b0 );
or ( \10195_b1 , \10190_b1 , \10194_b1 );
xor ( \10195_b0 , \10190_b0 , w_25824 );
not ( w_25824 , w_25825 );
and ( w_25825 , \10194_b1 , \10194_b0 );
or ( \10196_b1 , \6006_b1 , \5891_b1 );
not ( \5891_b1 , w_25826 );
and ( \10196_b0 , \6006_b0 , w_25827 );
and ( w_25826 , w_25827 , \5891_b0 );
or ( \10197_b1 , \6018_b1 , \5889_b1 );
not ( \5889_b1 , w_25828 );
and ( \10197_b0 , \6018_b0 , w_25829 );
and ( w_25828 , w_25829 , \5889_b0 );
or ( \10198_b1 , \10196_b1 , w_25831 );
not ( w_25831 , w_25832 );
and ( \10198_b0 , \10196_b0 , w_25833 );
and ( w_25832 ,  , w_25833 );
buf ( w_25831 , \10197_b1 );
not ( w_25831 , w_25834 );
not (  , w_25835 );
and ( w_25834 , w_25835 , \10197_b0 );
or ( \10199_b1 , \10198_b1 , w_25836 );
xor ( \10199_b0 , \10198_b0 , w_25838 );
not ( w_25838 , w_25839 );
and ( w_25839 , w_25836 , w_25837 );
buf ( w_25836 , \5898_b1 );
not ( w_25836 , w_25840 );
not ( w_25837 , w_25841 );
and ( w_25840 , w_25841 , \5898_b0 );
or ( \10200_b1 , \10195_b1 , \10199_b1 );
xor ( \10200_b0 , \10195_b0 , w_25842 );
not ( w_25842 , w_25843 );
and ( w_25843 , \10199_b1 , \10199_b0 );
or ( \10201_b1 , \10186_b1 , w_25844 );
xor ( \10201_b0 , \10186_b0 , w_25846 );
not ( w_25846 , w_25847 );
and ( w_25847 , w_25844 , w_25845 );
buf ( w_25844 , \10200_b1 );
not ( w_25844 , w_25848 );
not ( w_25845 , w_25849 );
and ( w_25848 , w_25849 , \10200_b0 );
or ( \10202_b1 , \10117_b1 , \10121_b1 );
not ( \10121_b1 , w_25850 );
and ( \10202_b0 , \10117_b0 , w_25851 );
and ( w_25850 , w_25851 , \10121_b0 );
or ( \10203_b1 , \10121_b1 , \10126_b1 );
not ( \10126_b1 , w_25852 );
and ( \10203_b0 , \10121_b0 , w_25853 );
and ( w_25852 , w_25853 , \10126_b0 );
or ( \10204_b1 , \10117_b1 , \10126_b1 );
not ( \10126_b1 , w_25854 );
and ( \10204_b0 , \10117_b0 , w_25855 );
and ( w_25854 , w_25855 , \10126_b0 );
or ( \10206_b1 , \10102_b1 , \10106_b1 );
not ( \10106_b1 , w_25856 );
and ( \10206_b0 , \10102_b0 , w_25857 );
and ( w_25856 , w_25857 , \10106_b0 );
or ( \10207_b1 , \10106_b1 , \10111_b1 );
not ( \10111_b1 , w_25858 );
and ( \10207_b0 , \10106_b0 , w_25859 );
and ( w_25858 , w_25859 , \10111_b0 );
or ( \10208_b1 , \10102_b1 , \10111_b1 );
not ( \10111_b1 , w_25860 );
and ( \10208_b0 , \10102_b0 , w_25861 );
and ( w_25860 , w_25861 , \10111_b0 );
or ( \10210_b1 , \10205_b1 , \10209_b1 );
xor ( \10210_b0 , \10205_b0 , w_25862 );
not ( w_25862 , w_25863 );
and ( w_25863 , \10209_b1 , \10209_b0 );
or ( \10211_b1 , \10093_b1 , \10097_b1 );
not ( \10097_b1 , w_25864 );
and ( \10211_b0 , \10093_b0 , w_25865 );
and ( w_25864 , w_25865 , \10097_b0 );
or ( \10212_b1 , \10210_b1 , \10211_b1 );
xor ( \10212_b0 , \10210_b0 , w_25866 );
not ( w_25866 , w_25867 );
and ( w_25867 , \10211_b1 , \10211_b0 );
or ( \10213_b1 , \10201_b1 , \10212_b1 );
xor ( \10213_b0 , \10201_b0 , w_25868 );
not ( w_25868 , w_25869 );
and ( w_25869 , \10212_b1 , \10212_b0 );
or ( \10214_b1 , \10077_b1 , \10081_b1 );
not ( \10081_b1 , w_25870 );
and ( \10214_b0 , \10077_b0 , w_25871 );
and ( w_25870 , w_25871 , \10081_b0 );
or ( \10215_b1 , \10081_b1 , \10086_b1 );
not ( \10086_b1 , w_25872 );
and ( \10215_b0 , \10081_b0 , w_25873 );
and ( w_25872 , w_25873 , \10086_b0 );
or ( \10216_b1 , \10077_b1 , \10086_b1 );
not ( \10086_b1 , w_25874 );
and ( \10216_b0 , \10077_b0 , w_25875 );
and ( w_25874 , w_25875 , \10086_b0 );
or ( \10218_b1 , \10065_b1 , \10069_b1 );
not ( \10069_b1 , w_25876 );
and ( \10218_b0 , \10065_b0 , w_25877 );
and ( w_25876 , w_25877 , \10069_b0 );
or ( \10219_b1 , \10069_b1 , \10074_b1 );
not ( \10074_b1 , w_25878 );
and ( \10219_b0 , \10069_b0 , w_25879 );
and ( w_25878 , w_25879 , \10074_b0 );
or ( \10220_b1 , \10065_b1 , \10074_b1 );
not ( \10074_b1 , w_25880 );
and ( \10220_b0 , \10065_b0 , w_25881 );
and ( w_25880 , w_25881 , \10074_b0 );
or ( \10222_b1 , \10217_b1 , \10221_b1 );
xor ( \10222_b0 , \10217_b0 , w_25882 );
not ( w_25882 , w_25883 );
and ( w_25883 , \10221_b1 , \10221_b0 );
or ( \10223_b1 , \10051_b1 , \10055_b1 );
not ( \10055_b1 , w_25884 );
and ( \10223_b0 , \10051_b0 , w_25885 );
and ( w_25884 , w_25885 , \10055_b0 );
or ( \10224_b1 , \10055_b1 , \10060_b1 );
not ( \10060_b1 , w_25886 );
and ( \10224_b0 , \10055_b0 , w_25887 );
and ( w_25886 , w_25887 , \10060_b0 );
or ( \10225_b1 , \10051_b1 , \10060_b1 );
not ( \10060_b1 , w_25888 );
and ( \10225_b0 , \10051_b0 , w_25889 );
and ( w_25888 , w_25889 , \10060_b0 );
or ( \10227_b1 , \10222_b1 , \10226_b1 );
xor ( \10227_b0 , \10222_b0 , w_25890 );
not ( w_25890 , w_25891 );
and ( w_25891 , \10226_b1 , \10226_b0 );
or ( \10228_b1 , \10213_b1 , \10227_b1 );
xor ( \10228_b0 , \10213_b0 , w_25892 );
not ( w_25892 , w_25893 );
and ( w_25893 , \10227_b1 , \10227_b0 );
or ( \10229_b1 , \10061_b1 , \10075_b1 );
not ( \10075_b1 , w_25894 );
and ( \10229_b0 , \10061_b0 , w_25895 );
and ( w_25894 , w_25895 , \10075_b0 );
or ( \10230_b1 , \10075_b1 , \10087_b1 );
not ( \10087_b1 , w_25896 );
and ( \10230_b0 , \10075_b0 , w_25897 );
and ( w_25896 , w_25897 , \10087_b0 );
or ( \10231_b1 , \10061_b1 , \10087_b1 );
not ( \10087_b1 , w_25898 );
and ( \10231_b0 , \10061_b0 , w_25899 );
and ( w_25898 , w_25899 , \10087_b0 );
or ( \10233_b1 , \5737_b1 , \7117_b1 );
not ( \7117_b1 , w_25900 );
and ( \10233_b0 , \5737_b0 , w_25901 );
and ( w_25900 , w_25901 , \7117_b0 );
buf ( \10234_b1 , \10233_b1 );
not ( \10234_b1 , w_25902 );
not ( \10234_b0 , w_25903 );
and ( w_25902 , w_25903 , \10233_b0 );
or ( \10235_b1 , \10234_b1 , w_25904 );
xor ( \10235_b0 , \10234_b0 , w_25906 );
not ( w_25906 , w_25907 );
and ( w_25907 , w_25904 , w_25905 );
buf ( w_25904 , \7123_b1 );
not ( w_25904 , w_25908 );
not ( w_25905 , w_25909 );
and ( w_25908 , w_25909 , \7123_b0 );
or ( \10236_b1 , \5962_b1 , \10235_b1 );
xor ( \10236_b0 , \5962_b0 , w_25910 );
not ( w_25910 , w_25911 );
and ( w_25911 , \10235_b1 , \10235_b0 );
or ( \10237_b1 , \5758_b1 , \7140_b1 );
not ( \7140_b1 , w_25912 );
and ( \10237_b0 , \5758_b0 , w_25913 );
and ( w_25912 , w_25913 , \7140_b0 );
or ( \10238_b1 , \5770_b1 , \7138_b1 );
not ( \7138_b1 , w_25914 );
and ( \10238_b0 , \5770_b0 , w_25915 );
and ( w_25914 , w_25915 , \7138_b0 );
or ( \10239_b1 , \10237_b1 , w_25917 );
not ( w_25917 , w_25918 );
and ( \10239_b0 , \10237_b0 , w_25919 );
and ( w_25918 ,  , w_25919 );
buf ( w_25917 , \10238_b1 );
not ( w_25917 , w_25920 );
not (  , w_25921 );
and ( w_25920 , w_25921 , \10238_b0 );
or ( \10240_b1 , \10239_b1 , w_25922 );
xor ( \10240_b0 , \10239_b0 , w_25924 );
not ( w_25924 , w_25925 );
and ( w_25925 , w_25922 , w_25923 );
buf ( w_25922 , \7146_b1 );
not ( w_25922 , w_25926 );
not ( w_25923 , w_25927 );
and ( w_25926 , w_25927 , \7146_b0 );
or ( \10241_b1 , \10236_b1 , \10240_b1 );
xor ( \10241_b0 , \10236_b0 , w_25928 );
not ( w_25928 , w_25929 );
and ( w_25929 , \10240_b1 , \10240_b0 );
or ( \10242_b1 , \10232_b1 , \10241_b1 );
xor ( \10242_b0 , \10232_b0 , w_25930 );
not ( w_25930 , w_25931 );
and ( w_25931 , \10241_b1 , \10241_b0 );
or ( \10243_b1 , \5906_b1 , \5790_b1 );
not ( \5790_b1 , w_25932 );
and ( \10243_b0 , \5906_b0 , w_25933 );
and ( w_25932 , w_25933 , \5790_b0 );
or ( \10244_b1 , \5918_b1 , \5788_b1 );
not ( \5788_b1 , w_25934 );
and ( \10244_b0 , \5918_b0 , w_25935 );
and ( w_25934 , w_25935 , \5788_b0 );
or ( \10245_b1 , \10243_b1 , w_25937 );
not ( w_25937 , w_25938 );
and ( \10245_b0 , \10243_b0 , w_25939 );
and ( w_25938 ,  , w_25939 );
buf ( w_25937 , \10244_b1 );
not ( w_25937 , w_25940 );
not (  , w_25941 );
and ( w_25940 , w_25941 , \10244_b0 );
or ( \10246_b1 , \10245_b1 , w_25942 );
xor ( \10246_b0 , \10245_b0 , w_25944 );
not ( w_25944 , w_25945 );
and ( w_25945 , w_25942 , w_25943 );
buf ( w_25942 , \5797_b1 );
not ( w_25942 , w_25946 );
not ( w_25943 , w_25947 );
and ( w_25946 , w_25947 , \5797_b0 );
or ( \10247_b1 , \5925_b1 , \5809_b1 );
not ( \5809_b1 , w_25948 );
and ( \10247_b0 , \5925_b0 , w_25949 );
and ( w_25948 , w_25949 , \5809_b0 );
or ( \10248_b1 , \5937_b1 , \5807_b1 );
not ( \5807_b1 , w_25950 );
and ( \10248_b0 , \5937_b0 , w_25951 );
and ( w_25950 , w_25951 , \5807_b0 );
or ( \10249_b1 , \10247_b1 , w_25953 );
not ( w_25953 , w_25954 );
and ( \10249_b0 , \10247_b0 , w_25955 );
and ( w_25954 ,  , w_25955 );
buf ( w_25953 , \10248_b1 );
not ( w_25953 , w_25956 );
not (  , w_25957 );
and ( w_25956 , w_25957 , \10248_b0 );
or ( \10250_b1 , \10249_b1 , w_25958 );
xor ( \10250_b0 , \10249_b0 , w_25960 );
not ( w_25960 , w_25961 );
and ( w_25961 , w_25958 , w_25959 );
buf ( w_25958 , \5816_b1 );
not ( w_25958 , w_25962 );
not ( w_25959 , w_25963 );
and ( w_25962 , w_25963 , \5816_b0 );
or ( \10251_b1 , \10246_b1 , \10250_b1 );
xor ( \10251_b0 , \10246_b0 , w_25964 );
not ( w_25964 , w_25965 );
and ( w_25965 , \10250_b1 , \10250_b0 );
or ( \10252_b1 , \5945_b1 , \5829_b1 );
not ( \5829_b1 , w_25966 );
and ( \10252_b0 , \5945_b0 , w_25967 );
and ( w_25966 , w_25967 , \5829_b0 );
or ( \10253_b1 , \5957_b1 , \5827_b1 );
not ( \5827_b1 , w_25968 );
and ( \10253_b0 , \5957_b0 , w_25969 );
and ( w_25968 , w_25969 , \5827_b0 );
or ( \10254_b1 , \10252_b1 , w_25971 );
not ( w_25971 , w_25972 );
and ( \10254_b0 , \10252_b0 , w_25973 );
and ( w_25972 ,  , w_25973 );
buf ( w_25971 , \10253_b1 );
not ( w_25971 , w_25974 );
not (  , w_25975 );
and ( w_25974 , w_25975 , \10253_b0 );
or ( \10255_b1 , \10254_b1 , w_25976 );
xor ( \10255_b0 , \10254_b0 , w_25978 );
not ( w_25978 , w_25979 );
and ( w_25979 , w_25976 , w_25977 );
buf ( w_25976 , \5836_b1 );
not ( w_25976 , w_25980 );
not ( w_25977 , w_25981 );
and ( w_25980 , w_25981 , \5836_b0 );
or ( \10256_b1 , \10251_b1 , \10255_b1 );
xor ( \10256_b0 , \10251_b0 , w_25982 );
not ( w_25982 , w_25983 );
and ( w_25983 , \10255_b1 , \10255_b0 );
or ( \10257_b1 , \5842_b1 , \7203_b1 );
not ( \7203_b1 , w_25984 );
and ( \10257_b0 , \5842_b0 , w_25985 );
and ( w_25984 , w_25985 , \7203_b0 );
or ( \10258_b1 , \5854_b1 , \7201_b1 );
not ( \7201_b1 , w_25986 );
and ( \10258_b0 , \5854_b0 , w_25987 );
and ( w_25986 , w_25987 , \7201_b0 );
or ( \10259_b1 , \10257_b1 , w_25989 );
not ( w_25989 , w_25990 );
and ( \10259_b0 , \10257_b0 , w_25991 );
and ( w_25990 ,  , w_25991 );
buf ( w_25989 , \10258_b1 );
not ( w_25989 , w_25992 );
not (  , w_25993 );
and ( w_25992 , w_25993 , \10258_b0 );
or ( \10260_b1 , \10259_b1 , w_25994 );
xor ( \10260_b0 , \10259_b0 , w_25996 );
not ( w_25996 , w_25997 );
and ( w_25997 , w_25994 , w_25995 );
buf ( w_25994 , \6824_b1 );
not ( w_25994 , w_25998 );
not ( w_25995 , w_25999 );
and ( w_25998 , w_25999 , \6824_b0 );
or ( \10261_b1 , \5861_b1 , \5750_b1 );
not ( \5750_b1 , w_26000 );
and ( \10261_b0 , \5861_b0 , w_26001 );
and ( w_26000 , w_26001 , \5750_b0 );
or ( \10262_b1 , \5873_b1 , \5748_b1 );
not ( \5748_b1 , w_26002 );
and ( \10262_b0 , \5873_b0 , w_26003 );
and ( w_26002 , w_26003 , \5748_b0 );
or ( \10263_b1 , \10261_b1 , w_26005 );
not ( w_26005 , w_26006 );
and ( \10263_b0 , \10261_b0 , w_26007 );
and ( w_26006 ,  , w_26007 );
buf ( w_26005 , \10262_b1 );
not ( w_26005 , w_26008 );
not (  , w_26009 );
and ( w_26008 , w_26009 , \10262_b0 );
or ( \10264_b1 , \10263_b1 , w_26010 );
xor ( \10264_b0 , \10263_b0 , w_26012 );
not ( w_26012 , w_26013 );
and ( w_26013 , w_26010 , w_26011 );
buf ( w_26010 , \5755_b1 );
not ( w_26010 , w_26014 );
not ( w_26011 , w_26015 );
and ( w_26014 , w_26015 , \5755_b0 );
or ( \10265_b1 , \10260_b1 , \10264_b1 );
xor ( \10265_b0 , \10260_b0 , w_26016 );
not ( w_26016 , w_26017 );
and ( w_26017 , \10264_b1 , \10264_b0 );
or ( \10266_b1 , \5881_b1 , \5768_b1 );
not ( \5768_b1 , w_26018 );
and ( \10266_b0 , \5881_b0 , w_26019 );
and ( w_26018 , w_26019 , \5768_b0 );
or ( \10267_b1 , \5893_b1 , \5766_b1 );
not ( \5766_b1 , w_26020 );
and ( \10267_b0 , \5893_b0 , w_26021 );
and ( w_26020 , w_26021 , \5766_b0 );
or ( \10268_b1 , \10266_b1 , w_26023 );
not ( w_26023 , w_26024 );
and ( \10268_b0 , \10266_b0 , w_26025 );
and ( w_26024 ,  , w_26025 );
buf ( w_26023 , \10267_b1 );
not ( w_26023 , w_26026 );
not (  , w_26027 );
and ( w_26026 , w_26027 , \10267_b0 );
or ( \10269_b1 , \10268_b1 , w_26028 );
xor ( \10269_b0 , \10268_b0 , w_26030 );
not ( w_26030 , w_26031 );
and ( w_26031 , w_26028 , w_26029 );
buf ( w_26028 , \5775_b1 );
not ( w_26028 , w_26032 );
not ( w_26029 , w_26033 );
and ( w_26032 , w_26033 , \5775_b0 );
or ( \10270_b1 , \10265_b1 , \10269_b1 );
xor ( \10270_b0 , \10265_b0 , w_26034 );
not ( w_26034 , w_26035 );
and ( w_26035 , \10269_b1 , \10269_b0 );
or ( \10271_b1 , \10256_b1 , \10270_b1 );
xor ( \10271_b0 , \10256_b0 , w_26036 );
not ( w_26036 , w_26037 );
and ( w_26037 , \10270_b1 , \10270_b0 );
or ( \10272_b1 , \5780_b1 , \7157_b1 );
not ( \7157_b1 , w_26038 );
and ( \10272_b0 , \5780_b0 , w_26039 );
and ( w_26038 , w_26039 , \7157_b0 );
or ( \10273_b1 , \5792_b1 , \7155_b1 );
not ( \7155_b1 , w_26040 );
and ( \10273_b0 , \5792_b0 , w_26041 );
and ( w_26040 , w_26041 , \7155_b0 );
or ( \10274_b1 , \10272_b1 , w_26043 );
not ( w_26043 , w_26044 );
and ( \10274_b0 , \10272_b0 , w_26045 );
and ( w_26044 ,  , w_26045 );
buf ( w_26043 , \10273_b1 );
not ( w_26043 , w_26046 );
not (  , w_26047 );
and ( w_26046 , w_26047 , \10273_b0 );
or ( \10275_b1 , \10274_b1 , w_26048 );
xor ( \10275_b0 , \10274_b0 , w_26050 );
not ( w_26050 , w_26051 );
and ( w_26051 , w_26048 , w_26049 );
buf ( w_26048 , \7163_b1 );
not ( w_26048 , w_26052 );
not ( w_26049 , w_26053 );
and ( w_26052 , w_26053 , \7163_b0 );
or ( \10276_b1 , \5799_b1 , \7175_b1 );
not ( \7175_b1 , w_26054 );
and ( \10276_b0 , \5799_b0 , w_26055 );
and ( w_26054 , w_26055 , \7175_b0 );
or ( \10277_b1 , \5811_b1 , \7173_b1 );
not ( \7173_b1 , w_26056 );
and ( \10277_b0 , \5811_b0 , w_26057 );
and ( w_26056 , w_26057 , \7173_b0 );
or ( \10278_b1 , \10276_b1 , w_26059 );
not ( w_26059 , w_26060 );
and ( \10278_b0 , \10276_b0 , w_26061 );
and ( w_26060 ,  , w_26061 );
buf ( w_26059 , \10277_b1 );
not ( w_26059 , w_26062 );
not (  , w_26063 );
and ( w_26062 , w_26063 , \10277_b0 );
or ( \10279_b1 , \10278_b1 , w_26064 );
xor ( \10279_b0 , \10278_b0 , w_26066 );
not ( w_26066 , w_26067 );
and ( w_26067 , w_26064 , w_26065 );
buf ( w_26064 , \7181_b1 );
not ( w_26064 , w_26068 );
not ( w_26065 , w_26069 );
and ( w_26068 , w_26069 , \7181_b0 );
or ( \10280_b1 , \10275_b1 , \10279_b1 );
xor ( \10280_b0 , \10275_b0 , w_26070 );
not ( w_26070 , w_26071 );
and ( w_26071 , \10279_b1 , \10279_b0 );
or ( \10281_b1 , \5819_b1 , \7192_b1 );
not ( \7192_b1 , w_26072 );
and ( \10281_b0 , \5819_b0 , w_26073 );
and ( w_26072 , w_26073 , \7192_b0 );
or ( \10282_b1 , \5831_b1 , \7190_b1 );
not ( \7190_b1 , w_26074 );
and ( \10282_b0 , \5831_b0 , w_26075 );
and ( w_26074 , w_26075 , \7190_b0 );
or ( \10283_b1 , \10281_b1 , w_26077 );
not ( w_26077 , w_26078 );
and ( \10283_b0 , \10281_b0 , w_26079 );
and ( w_26078 ,  , w_26079 );
buf ( w_26077 , \10282_b1 );
not ( w_26077 , w_26080 );
not (  , w_26081 );
and ( w_26080 , w_26081 , \10282_b0 );
or ( \10284_b1 , \10283_b1 , w_26082 );
xor ( \10284_b0 , \10283_b0 , w_26084 );
not ( w_26084 , w_26085 );
and ( w_26085 , w_26082 , w_26083 );
buf ( w_26082 , \7198_b1 );
not ( w_26082 , w_26086 );
not ( w_26083 , w_26087 );
and ( w_26086 , w_26087 , \7198_b0 );
or ( \10285_b1 , \10280_b1 , \10284_b1 );
xor ( \10285_b0 , \10280_b0 , w_26088 );
not ( w_26088 , w_26089 );
and ( w_26089 , \10284_b1 , \10284_b0 );
or ( \10286_b1 , \10271_b1 , \10285_b1 );
xor ( \10286_b0 , \10271_b0 , w_26090 );
not ( w_26090 , w_26091 );
and ( w_26091 , \10285_b1 , \10285_b0 );
or ( \10287_b1 , \10242_b1 , \10286_b1 );
xor ( \10287_b0 , \10242_b0 , w_26092 );
not ( w_26092 , w_26093 );
and ( w_26093 , \10286_b1 , \10286_b0 );
or ( \10288_b1 , \10228_b1 , \10287_b1 );
xor ( \10288_b0 , \10228_b0 , w_26094 );
not ( w_26094 , w_26095 );
and ( w_26095 , \10287_b1 , \10287_b0 );
or ( \10289_b1 , \10032_b1 , \10036_b1 );
not ( \10036_b1 , w_26096 );
and ( \10289_b0 , \10032_b0 , w_26097 );
and ( w_26096 , w_26097 , \10036_b0 );
or ( \10290_b1 , \10036_b1 , \10041_b1 );
not ( \10041_b1 , w_26098 );
and ( \10290_b0 , \10036_b0 , w_26099 );
and ( w_26098 , w_26099 , \10041_b0 );
or ( \10291_b1 , \10032_b1 , \10041_b1 );
not ( \10041_b1 , w_26100 );
and ( \10291_b0 , \10032_b0 , w_26101 );
and ( w_26100 , w_26101 , \10041_b0 );
or ( \10293_b1 , \10018_b1 , \10022_b1 );
not ( \10022_b1 , w_26102 );
and ( \10293_b0 , \10018_b0 , w_26103 );
and ( w_26102 , w_26103 , \10022_b0 );
or ( \10294_b1 , \10022_b1 , \10027_b1 );
not ( \10027_b1 , w_26104 );
and ( \10294_b0 , \10022_b0 , w_26105 );
and ( w_26104 , w_26105 , \10027_b0 );
or ( \10295_b1 , \10018_b1 , \10027_b1 );
not ( \10027_b1 , w_26106 );
and ( \10295_b0 , \10018_b0 , w_26107 );
and ( w_26106 , w_26107 , \10027_b0 );
or ( \10297_b1 , \10292_b1 , \10296_b1 );
xor ( \10297_b0 , \10292_b0 , w_26108 );
not ( w_26108 , w_26109 );
and ( w_26109 , \10296_b1 , \10296_b0 );
or ( \10298_b1 , \10098_b1 , \10112_b1 );
not ( \10112_b1 , w_26110 );
and ( \10298_b0 , \10098_b0 , w_26111 );
and ( w_26110 , w_26111 , \10112_b0 );
or ( \10299_b1 , \10112_b1 , \10127_b1 );
not ( \10127_b1 , w_26112 );
and ( \10299_b0 , \10112_b0 , w_26113 );
and ( w_26112 , w_26113 , \10127_b0 );
or ( \10300_b1 , \10098_b1 , \10127_b1 );
not ( \10127_b1 , w_26114 );
and ( \10300_b0 , \10098_b0 , w_26115 );
and ( w_26114 , w_26115 , \10127_b0 );
or ( \10302_b1 , \10297_b1 , \10301_b1 );
xor ( \10302_b0 , \10297_b0 , w_26116 );
not ( w_26116 , w_26117 );
and ( w_26117 , \10301_b1 , \10301_b0 );
or ( \10303_b1 , \10288_b1 , \10302_b1 );
xor ( \10303_b0 , \10288_b0 , w_26118 );
not ( w_26118 , w_26119 );
and ( w_26119 , \10302_b1 , \10302_b0 );
or ( \10304_b1 , \10174_b1 , \10303_b1 );
xor ( \10304_b0 , \10174_b0 , w_26120 );
not ( w_26120 , w_26121 );
and ( w_26121 , \10303_b1 , \10303_b0 );
or ( \10305_b1 , \10165_b1 , \10304_b1 );
xor ( \10305_b0 , \10165_b0 , w_26122 );
not ( w_26122 , w_26123 );
and ( w_26123 , \10304_b1 , \10304_b0 );
or ( \10306_b1 , \9990_b1 , \10004_b1 );
not ( \10004_b1 , w_26124 );
and ( \10306_b0 , \9990_b0 , w_26125 );
and ( w_26124 , w_26125 , \10004_b0 );
or ( \10307_b1 , \10004_b1 , \10143_b1 );
not ( \10143_b1 , w_26126 );
and ( \10307_b0 , \10004_b0 , w_26127 );
and ( w_26126 , w_26127 , \10143_b0 );
or ( \10308_b1 , \9990_b1 , \10143_b1 );
not ( \10143_b1 , w_26128 );
and ( \10308_b0 , \9990_b0 , w_26129 );
and ( w_26128 , w_26129 , \10143_b0 );
or ( \10310_b1 , \10305_b1 , w_26131 );
not ( w_26131 , w_26132 );
and ( \10310_b0 , \10305_b0 , w_26133 );
and ( w_26132 ,  , w_26133 );
buf ( w_26131 , \10309_b1 );
not ( w_26131 , w_26134 );
not (  , w_26135 );
and ( w_26134 , w_26135 , \10309_b0 );
or ( \10311_b1 , \10149_b1 , w_26137 );
not ( w_26137 , w_26138 );
and ( \10311_b0 , \10149_b0 , w_26139 );
and ( w_26138 ,  , w_26139 );
buf ( w_26137 , \10310_b1 );
not ( w_26137 , w_26140 );
not (  , w_26141 );
and ( w_26140 , w_26141 , \10310_b0 );
or ( \10312_b1 , \9986_b1 , w_26143 );
not ( w_26143 , w_26144 );
and ( \10312_b0 , \9986_b0 , w_26145 );
and ( w_26144 ,  , w_26145 );
buf ( w_26143 , \10311_b1 );
not ( w_26143 , w_26146 );
not (  , w_26147 );
and ( w_26146 , w_26147 , \10311_b0 );
or ( \10313_b1 , \9661_b1 , w_26149 );
not ( w_26149 , w_26150 );
and ( \10313_b0 , \9661_b0 , w_26151 );
and ( w_26150 ,  , w_26151 );
buf ( w_26149 , \10312_b1 );
not ( w_26149 , w_26152 );
not (  , w_26153 );
and ( w_26152 , w_26153 , \10312_b0 );
or ( \10314_b1 , \9010_b1 , w_26155 );
not ( w_26155 , w_26156 );
and ( \10314_b0 , \9010_b0 , w_26157 );
and ( w_26156 ,  , w_26157 );
buf ( w_26155 , \10313_b1 );
not ( w_26155 , w_26158 );
not (  , w_26159 );
and ( w_26158 , w_26159 , \10313_b0 );
or ( \10315_b1 , \10169_b1 , \10173_b1 );
not ( \10173_b1 , w_26160 );
and ( \10315_b0 , \10169_b0 , w_26161 );
and ( w_26160 , w_26161 , \10173_b0 );
or ( \10316_b1 , \10173_b1 , \10303_b1 );
not ( \10303_b1 , w_26162 );
and ( \10316_b0 , \10173_b0 , w_26163 );
and ( w_26162 , w_26163 , \10303_b0 );
or ( \10317_b1 , \10169_b1 , \10303_b1 );
not ( \10303_b1 , w_26164 );
and ( \10317_b0 , \10169_b0 , w_26165 );
and ( w_26164 , w_26165 , \10303_b0 );
or ( \10319_b1 , \10292_b1 , \10296_b1 );
not ( \10296_b1 , w_26166 );
and ( \10319_b0 , \10292_b0 , w_26167 );
and ( w_26166 , w_26167 , \10296_b0 );
or ( \10320_b1 , \10296_b1 , \10301_b1 );
not ( \10301_b1 , w_26168 );
and ( \10320_b0 , \10296_b0 , w_26169 );
and ( w_26168 , w_26169 , \10301_b0 );
or ( \10321_b1 , \10292_b1 , \10301_b1 );
not ( \10301_b1 , w_26170 );
and ( \10321_b0 , \10292_b0 , w_26171 );
and ( w_26170 , w_26171 , \10301_b0 );
or ( \10323_b1 , \10232_b1 , \10241_b1 );
not ( \10241_b1 , w_26172 );
and ( \10323_b0 , \10232_b0 , w_26173 );
and ( w_26172 , w_26173 , \10241_b0 );
or ( \10324_b1 , \10241_b1 , \10286_b1 );
not ( \10286_b1 , w_26174 );
and ( \10324_b0 , \10241_b0 , w_26175 );
and ( w_26174 , w_26175 , \10286_b0 );
or ( \10325_b1 , \10232_b1 , \10286_b1 );
not ( \10286_b1 , w_26176 );
and ( \10325_b0 , \10232_b0 , w_26177 );
and ( w_26176 , w_26177 , \10286_b0 );
or ( \10327_b1 , \10322_b1 , \10326_b1 );
xor ( \10327_b0 , \10322_b0 , w_26178 );
not ( w_26178 , w_26179 );
and ( w_26179 , \10326_b1 , \10326_b0 );
or ( \10328_b1 , \10201_b1 , \10212_b1 );
not ( \10212_b1 , w_26180 );
and ( \10328_b0 , \10201_b0 , w_26181 );
and ( w_26180 , w_26181 , \10212_b0 );
or ( \10329_b1 , \10212_b1 , \10227_b1 );
not ( \10227_b1 , w_26182 );
and ( \10329_b0 , \10212_b0 , w_26183 );
and ( w_26182 , w_26183 , \10227_b0 );
or ( \10330_b1 , \10201_b1 , \10227_b1 );
not ( \10227_b1 , w_26184 );
and ( \10330_b0 , \10201_b0 , w_26185 );
and ( w_26184 , w_26185 , \10227_b0 );
or ( \10332_b1 , \10327_b1 , \10331_b1 );
xor ( \10332_b0 , \10327_b0 , w_26186 );
not ( w_26186 , w_26187 );
and ( w_26187 , \10331_b1 , \10331_b0 );
or ( \10333_b1 , \10318_b1 , \10332_b1 );
xor ( \10333_b0 , \10318_b0 , w_26188 );
not ( w_26188 , w_26189 );
and ( w_26189 , \10332_b1 , \10332_b0 );
or ( \10334_b1 , \10157_b1 , \10161_b1 );
not ( \10161_b1 , w_26190 );
and ( \10334_b0 , \10157_b0 , w_26191 );
and ( w_26190 , w_26191 , \10161_b0 );
or ( \10335_b1 , \10161_b1 , \10163_b1 );
not ( \10163_b1 , w_26192 );
and ( \10335_b0 , \10161_b0 , w_26193 );
and ( w_26192 , w_26193 , \10163_b0 );
or ( \10336_b1 , \10157_b1 , \10163_b1 );
not ( \10163_b1 , w_26194 );
and ( \10336_b0 , \10157_b0 , w_26195 );
and ( w_26194 , w_26195 , \10163_b0 );
or ( \10338_b1 , \10228_b1 , \10287_b1 );
not ( \10287_b1 , w_26196 );
and ( \10338_b0 , \10228_b0 , w_26197 );
and ( w_26196 , w_26197 , \10287_b0 );
or ( \10339_b1 , \10287_b1 , \10302_b1 );
not ( \10302_b1 , w_26198 );
and ( \10339_b0 , \10287_b0 , w_26199 );
and ( w_26198 , w_26199 , \10302_b0 );
or ( \10340_b1 , \10228_b1 , \10302_b1 );
not ( \10302_b1 , w_26200 );
and ( \10340_b0 , \10228_b0 , w_26201 );
and ( w_26200 , w_26201 , \10302_b0 );
or ( \10342_b1 , \10337_b1 , \10341_b1 );
xor ( \10342_b0 , \10337_b0 , w_26202 );
not ( w_26202 , w_26203 );
and ( w_26203 , \10341_b1 , \10341_b0 );
or ( \10343_b1 , \10246_b1 , \10250_b1 );
not ( \10250_b1 , w_26204 );
and ( \10343_b0 , \10246_b0 , w_26205 );
and ( w_26204 , w_26205 , \10250_b0 );
or ( \10344_b1 , \10250_b1 , \10255_b1 );
not ( \10255_b1 , w_26206 );
and ( \10344_b0 , \10250_b0 , w_26207 );
and ( w_26206 , w_26207 , \10255_b0 );
or ( \10345_b1 , \10246_b1 , \10255_b1 );
not ( \10255_b1 , w_26208 );
and ( \10345_b0 , \10246_b0 , w_26209 );
and ( w_26208 , w_26209 , \10255_b0 );
or ( \10347_b1 , \10190_b1 , \10194_b1 );
not ( \10194_b1 , w_26210 );
and ( \10347_b0 , \10190_b0 , w_26211 );
and ( w_26210 , w_26211 , \10194_b0 );
or ( \10348_b1 , \10194_b1 , \10199_b1 );
not ( \10199_b1 , w_26212 );
and ( \10348_b0 , \10194_b0 , w_26213 );
and ( w_26212 , w_26213 , \10199_b0 );
or ( \10349_b1 , \10190_b1 , \10199_b1 );
not ( \10199_b1 , w_26214 );
and ( \10349_b0 , \10190_b0 , w_26215 );
and ( w_26214 , w_26215 , \10199_b0 );
or ( \10351_b1 , \10346_b1 , \10350_b1 );
xor ( \10351_b0 , \10346_b0 , w_26216 );
not ( w_26216 , w_26217 );
and ( w_26217 , \10350_b1 , \10350_b0 );
or ( \10352_b1 , \10178_b1 , \10182_b1 );
not ( \10182_b1 , w_26218 );
and ( \10352_b0 , \10178_b0 , w_26219 );
and ( w_26218 , w_26219 , \10182_b0 );
or ( \10353_b1 , \10182_b1 , \10185_b1 );
not ( \10185_b1 , w_26220 );
and ( \10353_b0 , \10182_b0 , w_26221 );
and ( w_26220 , w_26221 , \10185_b0 );
or ( \10354_b1 , \10178_b1 , \10185_b1 );
not ( \10185_b1 , w_26222 );
and ( \10354_b0 , \10178_b0 , w_26223 );
and ( w_26222 , w_26223 , \10185_b0 );
or ( \10356_b1 , \10351_b1 , \10355_b1 );
xor ( \10356_b0 , \10351_b0 , w_26224 );
not ( w_26224 , w_26225 );
and ( w_26225 , \10355_b1 , \10355_b0 );
or ( \10357_b1 , \5962_b1 , \10235_b1 );
not ( \10235_b1 , w_26226 );
and ( \10357_b0 , \5962_b0 , w_26227 );
and ( w_26226 , w_26227 , \10235_b0 );
or ( \10358_b1 , \10235_b1 , \10240_b1 );
not ( \10240_b1 , w_26228 );
and ( \10358_b0 , \10235_b0 , w_26229 );
and ( w_26228 , w_26229 , \10240_b0 );
or ( \10359_b1 , \5962_b1 , \10240_b1 );
not ( \10240_b1 , w_26230 );
and ( \10359_b0 , \5962_b0 , w_26231 );
and ( w_26230 , w_26231 , \10240_b0 );
or ( \10361_b1 , \10275_b1 , \10279_b1 );
not ( \10279_b1 , w_26232 );
and ( \10361_b0 , \10275_b0 , w_26233 );
and ( w_26232 , w_26233 , \10279_b0 );
or ( \10362_b1 , \10279_b1 , \10284_b1 );
not ( \10284_b1 , w_26234 );
and ( \10362_b0 , \10279_b0 , w_26235 );
and ( w_26234 , w_26235 , \10284_b0 );
or ( \10363_b1 , \10275_b1 , \10284_b1 );
not ( \10284_b1 , w_26236 );
and ( \10363_b0 , \10275_b0 , w_26237 );
and ( w_26236 , w_26237 , \10284_b0 );
or ( \10365_b1 , \10360_b1 , \10364_b1 );
xor ( \10365_b0 , \10360_b0 , w_26238 );
not ( w_26238 , w_26239 );
and ( w_26239 , \10364_b1 , \10364_b0 );
or ( \10366_b1 , \10260_b1 , \10264_b1 );
not ( \10264_b1 , w_26240 );
and ( \10366_b0 , \10260_b0 , w_26241 );
and ( w_26240 , w_26241 , \10264_b0 );
or ( \10367_b1 , \10264_b1 , \10269_b1 );
not ( \10269_b1 , w_26242 );
and ( \10367_b0 , \10264_b0 , w_26243 );
and ( w_26242 , w_26243 , \10269_b0 );
or ( \10368_b1 , \10260_b1 , \10269_b1 );
not ( \10269_b1 , w_26244 );
and ( \10368_b0 , \10260_b0 , w_26245 );
and ( w_26244 , w_26245 , \10269_b0 );
or ( \10370_b1 , \10365_b1 , \10369_b1 );
xor ( \10370_b0 , \10365_b0 , w_26246 );
not ( w_26246 , w_26247 );
and ( w_26247 , \10369_b1 , \10369_b0 );
or ( \10371_b1 , \10356_b1 , \10370_b1 );
xor ( \10371_b0 , \10356_b0 , w_26248 );
not ( w_26248 , w_26249 );
and ( w_26249 , \10370_b1 , \10370_b0 );
or ( \10372_b1 , \10256_b1 , \10270_b1 );
not ( \10270_b1 , w_26250 );
and ( \10372_b0 , \10256_b0 , w_26251 );
and ( w_26250 , w_26251 , \10270_b0 );
or ( \10373_b1 , \10270_b1 , \10285_b1 );
not ( \10285_b1 , w_26252 );
and ( \10373_b0 , \10270_b0 , w_26253 );
and ( w_26252 , w_26253 , \10285_b0 );
or ( \10374_b1 , \10256_b1 , \10285_b1 );
not ( \10285_b1 , w_26254 );
and ( \10374_b0 , \10256_b0 , w_26255 );
and ( w_26254 , w_26255 , \10285_b0 );
or ( \10376_b1 , \5873_b1 , \5750_b1 );
not ( \5750_b1 , w_26256 );
and ( \10376_b0 , \5873_b0 , w_26257 );
and ( w_26256 , w_26257 , \5750_b0 );
or ( \10377_b1 , \5842_b1 , \5748_b1 );
not ( \5748_b1 , w_26258 );
and ( \10377_b0 , \5842_b0 , w_26259 );
and ( w_26258 , w_26259 , \5748_b0 );
or ( \10378_b1 , \10376_b1 , w_26261 );
not ( w_26261 , w_26262 );
and ( \10378_b0 , \10376_b0 , w_26263 );
and ( w_26262 ,  , w_26263 );
buf ( w_26261 , \10377_b1 );
not ( w_26261 , w_26264 );
not (  , w_26265 );
and ( w_26264 , w_26265 , \10377_b0 );
or ( \10379_b1 , \10378_b1 , w_26266 );
xor ( \10379_b0 , \10378_b0 , w_26268 );
not ( w_26268 , w_26269 );
and ( w_26269 , w_26266 , w_26267 );
buf ( w_26266 , \5755_b1 );
not ( w_26266 , w_26270 );
not ( w_26267 , w_26271 );
and ( w_26270 , w_26271 , \5755_b0 );
or ( \10380_b1 , \5893_b1 , \5768_b1 );
not ( \5768_b1 , w_26272 );
and ( \10380_b0 , \5893_b0 , w_26273 );
and ( w_26272 , w_26273 , \5768_b0 );
or ( \10381_b1 , \5861_b1 , \5766_b1 );
not ( \5766_b1 , w_26274 );
and ( \10381_b0 , \5861_b0 , w_26275 );
and ( w_26274 , w_26275 , \5766_b0 );
or ( \10382_b1 , \10380_b1 , w_26277 );
not ( w_26277 , w_26278 );
and ( \10382_b0 , \10380_b0 , w_26279 );
and ( w_26278 ,  , w_26279 );
buf ( w_26277 , \10381_b1 );
not ( w_26277 , w_26280 );
not (  , w_26281 );
and ( w_26280 , w_26281 , \10381_b0 );
or ( \10383_b1 , \10382_b1 , w_26282 );
xor ( \10383_b0 , \10382_b0 , w_26284 );
not ( w_26284 , w_26285 );
and ( w_26285 , w_26282 , w_26283 );
buf ( w_26282 , \5775_b1 );
not ( w_26282 , w_26286 );
not ( w_26283 , w_26287 );
and ( w_26286 , w_26287 , \5775_b0 );
or ( \10384_b1 , \10379_b1 , \10383_b1 );
xor ( \10384_b0 , \10379_b0 , w_26288 );
not ( w_26288 , w_26289 );
and ( w_26289 , \10383_b1 , \10383_b0 );
or ( \10385_b1 , \5918_b1 , \5790_b1 );
not ( \5790_b1 , w_26290 );
and ( \10385_b0 , \5918_b0 , w_26291 );
and ( w_26290 , w_26291 , \5790_b0 );
or ( \10386_b1 , \5881_b1 , \5788_b1 );
not ( \5788_b1 , w_26292 );
and ( \10386_b0 , \5881_b0 , w_26293 );
and ( w_26292 , w_26293 , \5788_b0 );
or ( \10387_b1 , \10385_b1 , w_26295 );
not ( w_26295 , w_26296 );
and ( \10387_b0 , \10385_b0 , w_26297 );
and ( w_26296 ,  , w_26297 );
buf ( w_26295 , \10386_b1 );
not ( w_26295 , w_26298 );
not (  , w_26299 );
and ( w_26298 , w_26299 , \10386_b0 );
or ( \10388_b1 , \10387_b1 , w_26300 );
xor ( \10388_b0 , \10387_b0 , w_26302 );
not ( w_26302 , w_26303 );
and ( w_26303 , w_26300 , w_26301 );
buf ( w_26300 , \5797_b1 );
not ( w_26300 , w_26304 );
not ( w_26301 , w_26305 );
and ( w_26304 , w_26305 , \5797_b0 );
or ( \10389_b1 , \10384_b1 , \10388_b1 );
xor ( \10389_b0 , \10384_b0 , w_26306 );
not ( w_26306 , w_26307 );
and ( w_26307 , \10388_b1 , \10388_b0 );
or ( \10390_b1 , \5811_b1 , \7175_b1 );
not ( \7175_b1 , w_26308 );
and ( \10390_b0 , \5811_b0 , w_26309 );
and ( w_26308 , w_26309 , \7175_b0 );
or ( \10391_b1 , \5780_b1 , \7173_b1 );
not ( \7173_b1 , w_26310 );
and ( \10391_b0 , \5780_b0 , w_26311 );
and ( w_26310 , w_26311 , \7173_b0 );
or ( \10392_b1 , \10390_b1 , w_26313 );
not ( w_26313 , w_26314 );
and ( \10392_b0 , \10390_b0 , w_26315 );
and ( w_26314 ,  , w_26315 );
buf ( w_26313 , \10391_b1 );
not ( w_26313 , w_26316 );
not (  , w_26317 );
and ( w_26316 , w_26317 , \10391_b0 );
or ( \10393_b1 , \10392_b1 , w_26318 );
xor ( \10393_b0 , \10392_b0 , w_26320 );
not ( w_26320 , w_26321 );
and ( w_26321 , w_26318 , w_26319 );
buf ( w_26318 , \7181_b1 );
not ( w_26318 , w_26322 );
not ( w_26319 , w_26323 );
and ( w_26322 , w_26323 , \7181_b0 );
or ( \10394_b1 , \5831_b1 , \7192_b1 );
not ( \7192_b1 , w_26324 );
and ( \10394_b0 , \5831_b0 , w_26325 );
and ( w_26324 , w_26325 , \7192_b0 );
or ( \10395_b1 , \5799_b1 , \7190_b1 );
not ( \7190_b1 , w_26326 );
and ( \10395_b0 , \5799_b0 , w_26327 );
and ( w_26326 , w_26327 , \7190_b0 );
or ( \10396_b1 , \10394_b1 , w_26329 );
not ( w_26329 , w_26330 );
and ( \10396_b0 , \10394_b0 , w_26331 );
and ( w_26330 ,  , w_26331 );
buf ( w_26329 , \10395_b1 );
not ( w_26329 , w_26332 );
not (  , w_26333 );
and ( w_26332 , w_26333 , \10395_b0 );
or ( \10397_b1 , \10396_b1 , w_26334 );
xor ( \10397_b0 , \10396_b0 , w_26336 );
not ( w_26336 , w_26337 );
and ( w_26337 , w_26334 , w_26335 );
buf ( w_26334 , \7198_b1 );
not ( w_26334 , w_26338 );
not ( w_26335 , w_26339 );
and ( w_26338 , w_26339 , \7198_b0 );
or ( \10398_b1 , \10393_b1 , \10397_b1 );
xor ( \10398_b0 , \10393_b0 , w_26340 );
not ( w_26340 , w_26341 );
and ( w_26341 , \10397_b1 , \10397_b0 );
or ( \10399_b1 , \5854_b1 , \7203_b1 );
not ( \7203_b1 , w_26342 );
and ( \10399_b0 , \5854_b0 , w_26343 );
and ( w_26342 , w_26343 , \7203_b0 );
or ( \10400_b1 , \5819_b1 , \7201_b1 );
not ( \7201_b1 , w_26344 );
and ( \10400_b0 , \5819_b0 , w_26345 );
and ( w_26344 , w_26345 , \7201_b0 );
or ( \10401_b1 , \10399_b1 , w_26347 );
not ( w_26347 , w_26348 );
and ( \10401_b0 , \10399_b0 , w_26349 );
and ( w_26348 ,  , w_26349 );
buf ( w_26347 , \10400_b1 );
not ( w_26347 , w_26350 );
not (  , w_26351 );
and ( w_26350 , w_26351 , \10400_b0 );
or ( \10402_b1 , \10401_b1 , w_26352 );
xor ( \10402_b0 , \10401_b0 , w_26354 );
not ( w_26354 , w_26355 );
and ( w_26355 , w_26352 , w_26353 );
buf ( w_26352 , \6824_b1 );
not ( w_26352 , w_26356 );
not ( w_26353 , w_26357 );
and ( w_26356 , w_26357 , \6824_b0 );
or ( \10403_b1 , \10398_b1 , \10402_b1 );
xor ( \10403_b0 , \10398_b0 , w_26358 );
not ( w_26358 , w_26359 );
and ( w_26359 , \10402_b1 , \10402_b0 );
or ( \10404_b1 , \10389_b1 , \10403_b1 );
xor ( \10404_b0 , \10389_b0 , w_26360 );
not ( w_26360 , w_26361 );
and ( w_26361 , \10403_b1 , \10403_b0 );
buf ( \10405_b1 , \7123_b1 );
not ( \10405_b1 , w_26362 );
not ( \10405_b0 , w_26363 );
and ( w_26362 , w_26363 , \7123_b0 );
or ( \10406_b1 , \5770_b1 , \7140_b1 );
not ( \7140_b1 , w_26364 );
and ( \10406_b0 , \5770_b0 , w_26365 );
and ( w_26364 , w_26365 , \7140_b0 );
or ( \10407_b1 , \5737_b1 , \7138_b1 );
not ( \7138_b1 , w_26366 );
and ( \10407_b0 , \5737_b0 , w_26367 );
and ( w_26366 , w_26367 , \7138_b0 );
or ( \10408_b1 , \10406_b1 , w_26369 );
not ( w_26369 , w_26370 );
and ( \10408_b0 , \10406_b0 , w_26371 );
and ( w_26370 ,  , w_26371 );
buf ( w_26369 , \10407_b1 );
not ( w_26369 , w_26372 );
not (  , w_26373 );
and ( w_26372 , w_26373 , \10407_b0 );
or ( \10409_b1 , \10408_b1 , w_26374 );
xor ( \10409_b0 , \10408_b0 , w_26376 );
not ( w_26376 , w_26377 );
and ( w_26377 , w_26374 , w_26375 );
buf ( w_26374 , \7146_b1 );
not ( w_26374 , w_26378 );
not ( w_26375 , w_26379 );
and ( w_26378 , w_26379 , \7146_b0 );
or ( \10410_b1 , \10405_b1 , \10409_b1 );
xor ( \10410_b0 , \10405_b0 , w_26380 );
not ( w_26380 , w_26381 );
and ( w_26381 , \10409_b1 , \10409_b0 );
or ( \10411_b1 , \5792_b1 , \7157_b1 );
not ( \7157_b1 , w_26382 );
and ( \10411_b0 , \5792_b0 , w_26383 );
and ( w_26382 , w_26383 , \7157_b0 );
or ( \10412_b1 , \5758_b1 , \7155_b1 );
not ( \7155_b1 , w_26384 );
and ( \10412_b0 , \5758_b0 , w_26385 );
and ( w_26384 , w_26385 , \7155_b0 );
or ( \10413_b1 , \10411_b1 , w_26387 );
not ( w_26387 , w_26388 );
and ( \10413_b0 , \10411_b0 , w_26389 );
and ( w_26388 ,  , w_26389 );
buf ( w_26387 , \10412_b1 );
not ( w_26387 , w_26390 );
not (  , w_26391 );
and ( w_26390 , w_26391 , \10412_b0 );
or ( \10414_b1 , \10413_b1 , w_26392 );
xor ( \10414_b0 , \10413_b0 , w_26394 );
not ( w_26394 , w_26395 );
and ( w_26395 , w_26392 , w_26393 );
buf ( w_26392 , \7163_b1 );
not ( w_26392 , w_26396 );
not ( w_26393 , w_26397 );
and ( w_26396 , w_26397 , \7163_b0 );
or ( \10415_b1 , \10410_b1 , \10414_b1 );
xor ( \10415_b0 , \10410_b0 , w_26398 );
not ( w_26398 , w_26399 );
and ( w_26399 , \10414_b1 , \10414_b0 );
or ( \10416_b1 , \10404_b1 , \10415_b1 );
xor ( \10416_b0 , \10404_b0 , w_26400 );
not ( w_26400 , w_26401 );
and ( w_26401 , \10415_b1 , \10415_b0 );
or ( \10417_b1 , \10375_b1 , \10416_b1 );
xor ( \10417_b0 , \10375_b0 , w_26402 );
not ( w_26402 , w_26403 );
and ( w_26403 , \10416_b1 , \10416_b0 );
or ( \10418_b1 , \6057_b1 , \5935_b1 );
not ( \5935_b1 , w_26404 );
and ( \10418_b0 , \6057_b0 , w_26405 );
and ( w_26404 , w_26405 , \5935_b0 );
or ( \10419_b1 , \6029_b1 , \5933_b1 );
not ( \5933_b1 , w_26406 );
and ( \10419_b0 , \6029_b0 , w_26407 );
and ( w_26406 , w_26407 , \5933_b0 );
or ( \10420_b1 , \10418_b1 , w_26409 );
not ( w_26409 , w_26410 );
and ( \10420_b0 , \10418_b0 , w_26411 );
and ( w_26410 ,  , w_26411 );
buf ( w_26409 , \10419_b1 );
not ( w_26409 , w_26412 );
not (  , w_26413 );
and ( w_26412 , w_26413 , \10419_b0 );
or ( \10421_b1 , \10420_b1 , w_26414 );
xor ( \10421_b0 , \10420_b0 , w_26416 );
not ( w_26416 , w_26417 );
and ( w_26417 , w_26414 , w_26415 );
buf ( w_26414 , \5942_b1 );
not ( w_26414 , w_26418 );
not ( w_26415 , w_26419 );
and ( w_26418 , w_26419 , \5942_b0 );
or ( \10422_b1 , \6065_b1 , \5955_b1 );
not ( \5955_b1 , w_26420 );
and ( \10422_b0 , \6065_b0 , w_26421 );
and ( w_26420 , w_26421 , \5955_b0 );
or ( \10423_b1 , \6048_b1 , \5953_b1 );
not ( \5953_b1 , w_26422 );
and ( \10423_b0 , \6048_b0 , w_26423 );
and ( w_26422 , w_26423 , \5953_b0 );
or ( \10424_b1 , \10422_b1 , w_26425 );
not ( w_26425 , w_26426 );
and ( \10424_b0 , \10422_b0 , w_26427 );
and ( w_26426 ,  , w_26427 );
buf ( w_26425 , \10423_b1 );
not ( w_26425 , w_26428 );
not (  , w_26429 );
and ( w_26428 , w_26429 , \10423_b0 );
or ( \10425_b1 , \10424_b1 , w_26430 );
xor ( \10425_b0 , \10424_b0 , w_26432 );
not ( w_26432 , w_26433 );
and ( w_26433 , w_26430 , w_26431 );
buf ( w_26430 , \5962_b1 );
not ( w_26430 , w_26434 );
not ( w_26431 , w_26435 );
and ( w_26434 , w_26435 , \5962_b0 );
or ( \10426_b1 , \10421_b1 , \10425_b1 );
xor ( \10426_b0 , \10421_b0 , w_26436 );
not ( w_26436 , w_26437 );
and ( w_26437 , \10425_b1 , \10425_b0 );
or ( \10427_b1 , \5998_b1 , \5871_b1 );
not ( \5871_b1 , w_26438 );
and ( \10427_b0 , \5998_b0 , w_26439 );
and ( w_26438 , w_26439 , \5871_b0 );
or ( \10428_b1 , \5967_b1 , \5869_b1 );
not ( \5869_b1 , w_26440 );
and ( \10428_b0 , \5967_b0 , w_26441 );
and ( w_26440 , w_26441 , \5869_b0 );
or ( \10429_b1 , \10427_b1 , w_26443 );
not ( w_26443 , w_26444 );
and ( \10429_b0 , \10427_b0 , w_26445 );
and ( w_26444 ,  , w_26445 );
buf ( w_26443 , \10428_b1 );
not ( w_26443 , w_26446 );
not (  , w_26447 );
and ( w_26446 , w_26447 , \10428_b0 );
or ( \10430_b1 , \10429_b1 , w_26448 );
xor ( \10430_b0 , \10429_b0 , w_26450 );
not ( w_26450 , w_26451 );
and ( w_26451 , w_26448 , w_26449 );
buf ( w_26448 , \5878_b1 );
not ( w_26448 , w_26452 );
not ( w_26449 , w_26453 );
and ( w_26452 , w_26453 , \5878_b0 );
or ( \10431_b1 , \6018_b1 , \5891_b1 );
not ( \5891_b1 , w_26454 );
and ( \10431_b0 , \6018_b0 , w_26455 );
and ( w_26454 , w_26455 , \5891_b0 );
or ( \10432_b1 , \5986_b1 , \5889_b1 );
not ( \5889_b1 , w_26456 );
and ( \10432_b0 , \5986_b0 , w_26457 );
and ( w_26456 , w_26457 , \5889_b0 );
or ( \10433_b1 , \10431_b1 , w_26459 );
not ( w_26459 , w_26460 );
and ( \10433_b0 , \10431_b0 , w_26461 );
and ( w_26460 ,  , w_26461 );
buf ( w_26459 , \10432_b1 );
not ( w_26459 , w_26462 );
not (  , w_26463 );
and ( w_26462 , w_26463 , \10432_b0 );
or ( \10434_b1 , \10433_b1 , w_26464 );
xor ( \10434_b0 , \10433_b0 , w_26466 );
not ( w_26466 , w_26467 );
and ( w_26467 , w_26464 , w_26465 );
buf ( w_26464 , \5898_b1 );
not ( w_26464 , w_26468 );
not ( w_26465 , w_26469 );
and ( w_26468 , w_26469 , \5898_b0 );
or ( \10435_b1 , \10430_b1 , \10434_b1 );
xor ( \10435_b0 , \10430_b0 , w_26470 );
not ( w_26470 , w_26471 );
and ( w_26471 , \10434_b1 , \10434_b0 );
or ( \10436_b1 , \6041_b1 , \5916_b1 );
not ( \5916_b1 , w_26472 );
and ( \10436_b0 , \6041_b0 , w_26473 );
and ( w_26472 , w_26473 , \5916_b0 );
or ( \10437_b1 , \6006_b1 , \5914_b1 );
not ( \5914_b1 , w_26474 );
and ( \10437_b0 , \6006_b0 , w_26475 );
and ( w_26474 , w_26475 , \5914_b0 );
or ( \10438_b1 , \10436_b1 , w_26477 );
not ( w_26477 , w_26478 );
and ( \10438_b0 , \10436_b0 , w_26479 );
and ( w_26478 ,  , w_26479 );
buf ( w_26477 , \10437_b1 );
not ( w_26477 , w_26480 );
not (  , w_26481 );
and ( w_26480 , w_26481 , \10437_b0 );
or ( \10439_b1 , \10438_b1 , w_26482 );
xor ( \10439_b0 , \10438_b0 , w_26484 );
not ( w_26484 , w_26485 );
and ( w_26485 , w_26482 , w_26483 );
buf ( w_26482 , \5923_b1 );
not ( w_26482 , w_26486 );
not ( w_26483 , w_26487 );
and ( w_26486 , w_26487 , \5923_b0 );
or ( \10440_b1 , \10435_b1 , \10439_b1 );
xor ( \10440_b0 , \10435_b0 , w_26488 );
not ( w_26488 , w_26489 );
and ( w_26489 , \10439_b1 , \10439_b0 );
or ( \10441_b1 , \10426_b1 , \10440_b1 );
xor ( \10441_b0 , \10426_b0 , w_26490 );
not ( w_26490 , w_26491 );
and ( w_26491 , \10440_b1 , \10440_b0 );
or ( \10442_b1 , \5937_b1 , \5809_b1 );
not ( \5809_b1 , w_26492 );
and ( \10442_b0 , \5937_b0 , w_26493 );
and ( w_26492 , w_26493 , \5809_b0 );
or ( \10443_b1 , \5906_b1 , \5807_b1 );
not ( \5807_b1 , w_26494 );
and ( \10443_b0 , \5906_b0 , w_26495 );
and ( w_26494 , w_26495 , \5807_b0 );
or ( \10444_b1 , \10442_b1 , w_26497 );
not ( w_26497 , w_26498 );
and ( \10444_b0 , \10442_b0 , w_26499 );
and ( w_26498 ,  , w_26499 );
buf ( w_26497 , \10443_b1 );
not ( w_26497 , w_26500 );
not (  , w_26501 );
and ( w_26500 , w_26501 , \10443_b0 );
or ( \10445_b1 , \10444_b1 , w_26502 );
xor ( \10445_b0 , \10444_b0 , w_26504 );
not ( w_26504 , w_26505 );
and ( w_26505 , w_26502 , w_26503 );
buf ( w_26502 , \5816_b1 );
not ( w_26502 , w_26506 );
not ( w_26503 , w_26507 );
and ( w_26506 , w_26507 , \5816_b0 );
or ( \10446_b1 , \5957_b1 , \5829_b1 );
not ( \5829_b1 , w_26508 );
and ( \10446_b0 , \5957_b0 , w_26509 );
and ( w_26508 , w_26509 , \5829_b0 );
or ( \10447_b1 , \5925_b1 , \5827_b1 );
not ( \5827_b1 , w_26510 );
and ( \10447_b0 , \5925_b0 , w_26511 );
and ( w_26510 , w_26511 , \5827_b0 );
or ( \10448_b1 , \10446_b1 , w_26513 );
not ( w_26513 , w_26514 );
and ( \10448_b0 , \10446_b0 , w_26515 );
and ( w_26514 ,  , w_26515 );
buf ( w_26513 , \10447_b1 );
not ( w_26513 , w_26516 );
not (  , w_26517 );
and ( w_26516 , w_26517 , \10447_b0 );
or ( \10449_b1 , \10448_b1 , w_26518 );
xor ( \10449_b0 , \10448_b0 , w_26520 );
not ( w_26520 , w_26521 );
and ( w_26521 , w_26518 , w_26519 );
buf ( w_26518 , \5836_b1 );
not ( w_26518 , w_26522 );
not ( w_26519 , w_26523 );
and ( w_26522 , w_26523 , \5836_b0 );
or ( \10450_b1 , \10445_b1 , \10449_b1 );
xor ( \10450_b0 , \10445_b0 , w_26524 );
not ( w_26524 , w_26525 );
and ( w_26525 , \10449_b1 , \10449_b0 );
or ( \10451_b1 , \5979_b1 , \5852_b1 );
not ( \5852_b1 , w_26526 );
and ( \10451_b0 , \5979_b0 , w_26527 );
and ( w_26526 , w_26527 , \5852_b0 );
or ( \10452_b1 , \5945_b1 , \5850_b1 );
not ( \5850_b1 , w_26528 );
and ( \10452_b0 , \5945_b0 , w_26529 );
and ( w_26528 , w_26529 , \5850_b0 );
or ( \10453_b1 , \10451_b1 , w_26531 );
not ( w_26531 , w_26532 );
and ( \10453_b0 , \10451_b0 , w_26533 );
and ( w_26532 ,  , w_26533 );
buf ( w_26531 , \10452_b1 );
not ( w_26531 , w_26534 );
not (  , w_26535 );
and ( w_26534 , w_26535 , \10452_b0 );
or ( \10454_b1 , \10453_b1 , w_26536 );
xor ( \10454_b0 , \10453_b0 , w_26538 );
not ( w_26538 , w_26539 );
and ( w_26539 , w_26536 , w_26537 );
buf ( w_26536 , \5859_b1 );
not ( w_26536 , w_26540 );
not ( w_26537 , w_26541 );
and ( w_26540 , w_26541 , \5859_b0 );
or ( \10455_b1 , \10450_b1 , \10454_b1 );
xor ( \10455_b0 , \10450_b0 , w_26542 );
not ( w_26542 , w_26543 );
and ( w_26543 , \10454_b1 , \10454_b0 );
or ( \10456_b1 , \10441_b1 , \10455_b1 );
xor ( \10456_b0 , \10441_b0 , w_26544 );
not ( w_26544 , w_26545 );
and ( w_26545 , \10455_b1 , \10455_b0 );
or ( \10457_b1 , \10417_b1 , \10456_b1 );
xor ( \10457_b0 , \10417_b0 , w_26546 );
not ( w_26546 , w_26547 );
and ( w_26547 , \10456_b1 , \10456_b0 );
or ( \10458_b1 , \10371_b1 , \10457_b1 );
xor ( \10458_b0 , \10371_b0 , w_26548 );
not ( w_26548 , w_26549 );
and ( w_26549 , \10457_b1 , \10457_b0 );
or ( \10459_b1 , \10217_b1 , \10221_b1 );
not ( \10221_b1 , w_26550 );
and ( \10459_b0 , \10217_b0 , w_26551 );
and ( w_26550 , w_26551 , \10221_b0 );
or ( \10460_b1 , \10221_b1 , \10226_b1 );
not ( \10226_b1 , w_26552 );
and ( \10460_b0 , \10221_b0 , w_26553 );
and ( w_26552 , w_26553 , \10226_b0 );
or ( \10461_b1 , \10217_b1 , \10226_b1 );
not ( \10226_b1 , w_26554 );
and ( \10461_b0 , \10217_b0 , w_26555 );
and ( w_26554 , w_26555 , \10226_b0 );
or ( \10463_b1 , \10205_b1 , \10209_b1 );
not ( \10209_b1 , w_26556 );
and ( \10463_b0 , \10205_b0 , w_26557 );
and ( w_26556 , w_26557 , \10209_b0 );
or ( \10464_b1 , \10209_b1 , \10211_b1 );
not ( \10211_b1 , w_26558 );
and ( \10464_b0 , \10209_b0 , w_26559 );
and ( w_26558 , w_26559 , \10211_b0 );
or ( \10465_b1 , \10205_b1 , \10211_b1 );
not ( \10211_b1 , w_26560 );
and ( \10465_b0 , \10205_b0 , w_26561 );
and ( w_26560 , w_26561 , \10211_b0 );
or ( \10467_b1 , \10462_b1 , \10466_b1 );
xor ( \10467_b0 , \10462_b0 , w_26562 );
not ( w_26562 , w_26563 );
and ( w_26563 , \10466_b1 , \10466_b0 );
or ( \10468_b1 , \10186_b1 , w_26564 );
or ( \10468_b0 , \10186_b0 , \10200_b0 );
not ( \10200_b0 , w_26565 );
and ( w_26565 , w_26564 , \10200_b1 );
or ( \10469_b1 , \10467_b1 , \10468_b1 );
xor ( \10469_b0 , \10467_b0 , w_26566 );
not ( w_26566 , w_26567 );
and ( w_26567 , \10468_b1 , \10468_b0 );
or ( \10470_b1 , \10458_b1 , \10469_b1 );
xor ( \10470_b0 , \10458_b0 , w_26568 );
not ( w_26568 , w_26569 );
and ( w_26569 , \10469_b1 , \10469_b0 );
or ( \10471_b1 , \10342_b1 , \10470_b1 );
xor ( \10471_b0 , \10342_b0 , w_26570 );
not ( w_26570 , w_26571 );
and ( w_26571 , \10470_b1 , \10470_b0 );
or ( \10472_b1 , \10333_b1 , \10471_b1 );
xor ( \10472_b0 , \10333_b0 , w_26572 );
not ( w_26572 , w_26573 );
and ( w_26573 , \10471_b1 , \10471_b0 );
or ( \10473_b1 , \10153_b1 , \10164_b1 );
not ( \10164_b1 , w_26574 );
and ( \10473_b0 , \10153_b0 , w_26575 );
and ( w_26574 , w_26575 , \10164_b0 );
or ( \10474_b1 , \10164_b1 , \10304_b1 );
not ( \10304_b1 , w_26576 );
and ( \10474_b0 , \10164_b0 , w_26577 );
and ( w_26576 , w_26577 , \10304_b0 );
or ( \10475_b1 , \10153_b1 , \10304_b1 );
not ( \10304_b1 , w_26578 );
and ( \10475_b0 , \10153_b0 , w_26579 );
and ( w_26578 , w_26579 , \10304_b0 );
or ( \10477_b1 , \10472_b1 , w_26581 );
not ( w_26581 , w_26582 );
and ( \10477_b0 , \10472_b0 , w_26583 );
and ( w_26582 ,  , w_26583 );
buf ( w_26581 , \10476_b1 );
not ( w_26581 , w_26584 );
not (  , w_26585 );
and ( w_26584 , w_26585 , \10476_b0 );
or ( \10478_b1 , \10337_b1 , \10341_b1 );
not ( \10341_b1 , w_26586 );
and ( \10478_b0 , \10337_b0 , w_26587 );
and ( w_26586 , w_26587 , \10341_b0 );
or ( \10479_b1 , \10341_b1 , \10470_b1 );
not ( \10470_b1 , w_26588 );
and ( \10479_b0 , \10341_b0 , w_26589 );
and ( w_26588 , w_26589 , \10470_b0 );
or ( \10480_b1 , \10337_b1 , \10470_b1 );
not ( \10470_b1 , w_26590 );
and ( \10480_b0 , \10337_b0 , w_26591 );
and ( w_26590 , w_26591 , \10470_b0 );
or ( \10482_b1 , \10462_b1 , \10466_b1 );
not ( \10466_b1 , w_26592 );
and ( \10482_b0 , \10462_b0 , w_26593 );
and ( w_26592 , w_26593 , \10466_b0 );
or ( \10483_b1 , \10466_b1 , \10468_b1 );
not ( \10468_b1 , w_26594 );
and ( \10483_b0 , \10466_b0 , w_26595 );
and ( w_26594 , w_26595 , \10468_b0 );
or ( \10484_b1 , \10462_b1 , \10468_b1 );
not ( \10468_b1 , w_26596 );
and ( \10484_b0 , \10462_b0 , w_26597 );
and ( w_26596 , w_26597 , \10468_b0 );
or ( \10486_b1 , \10375_b1 , \10416_b1 );
not ( \10416_b1 , w_26598 );
and ( \10486_b0 , \10375_b0 , w_26599 );
and ( w_26598 , w_26599 , \10416_b0 );
or ( \10487_b1 , \10416_b1 , \10456_b1 );
not ( \10456_b1 , w_26600 );
and ( \10487_b0 , \10416_b0 , w_26601 );
and ( w_26600 , w_26601 , \10456_b0 );
or ( \10488_b1 , \10375_b1 , \10456_b1 );
not ( \10456_b1 , w_26602 );
and ( \10488_b0 , \10375_b0 , w_26603 );
and ( w_26602 , w_26603 , \10456_b0 );
or ( \10490_b1 , \10485_b1 , \10489_b1 );
xor ( \10490_b0 , \10485_b0 , w_26604 );
not ( w_26604 , w_26605 );
and ( w_26605 , \10489_b1 , \10489_b0 );
or ( \10491_b1 , \10356_b1 , \10370_b1 );
not ( \10370_b1 , w_26606 );
and ( \10491_b0 , \10356_b0 , w_26607 );
and ( w_26606 , w_26607 , \10370_b0 );
or ( \10492_b1 , \10490_b1 , \10491_b1 );
xor ( \10492_b0 , \10490_b0 , w_26608 );
not ( w_26608 , w_26609 );
and ( w_26609 , \10491_b1 , \10491_b0 );
or ( \10493_b1 , \10481_b1 , \10492_b1 );
xor ( \10493_b0 , \10481_b0 , w_26610 );
not ( w_26610 , w_26611 );
and ( w_26611 , \10492_b1 , \10492_b0 );
or ( \10494_b1 , \10322_b1 , \10326_b1 );
not ( \10326_b1 , w_26612 );
and ( \10494_b0 , \10322_b0 , w_26613 );
and ( w_26612 , w_26613 , \10326_b0 );
or ( \10495_b1 , \10326_b1 , \10331_b1 );
not ( \10331_b1 , w_26614 );
and ( \10495_b0 , \10326_b0 , w_26615 );
and ( w_26614 , w_26615 , \10331_b0 );
or ( \10496_b1 , \10322_b1 , \10331_b1 );
not ( \10331_b1 , w_26616 );
and ( \10496_b0 , \10322_b0 , w_26617 );
and ( w_26616 , w_26617 , \10331_b0 );
or ( \10498_b1 , \10371_b1 , \10457_b1 );
not ( \10457_b1 , w_26618 );
and ( \10498_b0 , \10371_b0 , w_26619 );
and ( w_26618 , w_26619 , \10457_b0 );
or ( \10499_b1 , \10457_b1 , \10469_b1 );
not ( \10469_b1 , w_26620 );
and ( \10499_b0 , \10457_b0 , w_26621 );
and ( w_26620 , w_26621 , \10469_b0 );
or ( \10500_b1 , \10371_b1 , \10469_b1 );
not ( \10469_b1 , w_26622 );
and ( \10500_b0 , \10371_b0 , w_26623 );
and ( w_26622 , w_26623 , \10469_b0 );
or ( \10502_b1 , \10497_b1 , \10501_b1 );
xor ( \10502_b0 , \10497_b0 , w_26624 );
not ( w_26624 , w_26625 );
and ( w_26625 , \10501_b1 , \10501_b0 );
or ( \10503_b1 , \6029_b1 , \5935_b1 );
not ( \5935_b1 , w_26626 );
and ( \10503_b0 , \6029_b0 , w_26627 );
and ( w_26626 , w_26627 , \5935_b0 );
or ( \10504_b1 , \6041_b1 , \5933_b1 );
not ( \5933_b1 , w_26628 );
and ( \10504_b0 , \6041_b0 , w_26629 );
and ( w_26628 , w_26629 , \5933_b0 );
or ( \10505_b1 , \10503_b1 , w_26631 );
not ( w_26631 , w_26632 );
and ( \10505_b0 , \10503_b0 , w_26633 );
and ( w_26632 ,  , w_26633 );
buf ( w_26631 , \10504_b1 );
not ( w_26631 , w_26634 );
not (  , w_26635 );
and ( w_26634 , w_26635 , \10504_b0 );
or ( \10506_b1 , \10505_b1 , w_26636 );
xor ( \10506_b0 , \10505_b0 , w_26638 );
not ( w_26638 , w_26639 );
and ( w_26639 , w_26636 , w_26637 );
buf ( w_26636 , \5942_b1 );
not ( w_26636 , w_26640 );
not ( w_26637 , w_26641 );
and ( w_26640 , w_26641 , \5942_b0 );
or ( \10507_b1 , \6048_b1 , \5955_b1 );
not ( \5955_b1 , w_26642 );
and ( \10507_b0 , \6048_b0 , w_26643 );
and ( w_26642 , w_26643 , \5955_b0 );
or ( \10508_b1 , \6057_b1 , \5953_b1 );
not ( \5953_b1 , w_26644 );
and ( \10508_b0 , \6057_b0 , w_26645 );
and ( w_26644 , w_26645 , \5953_b0 );
or ( \10509_b1 , \10507_b1 , w_26647 );
not ( w_26647 , w_26648 );
and ( \10509_b0 , \10507_b0 , w_26649 );
and ( w_26648 ,  , w_26649 );
buf ( w_26647 , \10508_b1 );
not ( w_26647 , w_26650 );
not (  , w_26651 );
and ( w_26650 , w_26651 , \10508_b0 );
or ( \10510_b1 , \10509_b1 , w_26652 );
xor ( \10510_b0 , \10509_b0 , w_26654 );
not ( w_26654 , w_26655 );
and ( w_26655 , w_26652 , w_26653 );
buf ( w_26652 , \5962_b1 );
not ( w_26652 , w_26656 );
not ( w_26653 , w_26657 );
and ( w_26656 , w_26657 , \5962_b0 );
or ( \10511_b1 , \10506_b1 , \10510_b1 );
xor ( \10511_b0 , \10506_b0 , w_26658 );
not ( w_26658 , w_26659 );
and ( w_26659 , \10510_b1 , \10510_b0 );
or ( \10512_b1 , \6065_b1 , w_26661 );
not ( w_26661 , w_26662 );
and ( \10512_b0 , \6065_b0 , w_26663 );
and ( w_26662 ,  , w_26663 );
buf ( w_26661 , \5975_b1 );
not ( w_26661 , w_26664 );
not (  , w_26665 );
and ( w_26664 , w_26665 , \5975_b0 );
or ( \10513_b1 , \10512_b1 , w_26666 );
xor ( \10513_b0 , \10512_b0 , w_26668 );
not ( w_26668 , w_26669 );
and ( w_26669 , w_26666 , w_26667 );
buf ( w_26666 , \5984_b1 );
not ( w_26666 , w_26670 );
not ( w_26667 , w_26671 );
and ( w_26670 , w_26671 , \5984_b0 );
or ( \10514_b1 , \10511_b1 , \10513_b1 );
xor ( \10514_b0 , \10511_b0 , w_26672 );
not ( w_26672 , w_26673 );
and ( w_26673 , \10513_b1 , \10513_b0 );
or ( \10515_b1 , \5967_b1 , \5871_b1 );
not ( \5871_b1 , w_26674 );
and ( \10515_b0 , \5967_b0 , w_26675 );
and ( w_26674 , w_26675 , \5871_b0 );
or ( \10516_b1 , \5979_b1 , \5869_b1 );
not ( \5869_b1 , w_26676 );
and ( \10516_b0 , \5979_b0 , w_26677 );
and ( w_26676 , w_26677 , \5869_b0 );
or ( \10517_b1 , \10515_b1 , w_26679 );
not ( w_26679 , w_26680 );
and ( \10517_b0 , \10515_b0 , w_26681 );
and ( w_26680 ,  , w_26681 );
buf ( w_26679 , \10516_b1 );
not ( w_26679 , w_26682 );
not (  , w_26683 );
and ( w_26682 , w_26683 , \10516_b0 );
or ( \10518_b1 , \10517_b1 , w_26684 );
xor ( \10518_b0 , \10517_b0 , w_26686 );
not ( w_26686 , w_26687 );
and ( w_26687 , w_26684 , w_26685 );
buf ( w_26684 , \5878_b1 );
not ( w_26684 , w_26688 );
not ( w_26685 , w_26689 );
and ( w_26688 , w_26689 , \5878_b0 );
or ( \10519_b1 , \5986_b1 , \5891_b1 );
not ( \5891_b1 , w_26690 );
and ( \10519_b0 , \5986_b0 , w_26691 );
and ( w_26690 , w_26691 , \5891_b0 );
or ( \10520_b1 , \5998_b1 , \5889_b1 );
not ( \5889_b1 , w_26692 );
and ( \10520_b0 , \5998_b0 , w_26693 );
and ( w_26692 , w_26693 , \5889_b0 );
or ( \10521_b1 , \10519_b1 , w_26695 );
not ( w_26695 , w_26696 );
and ( \10521_b0 , \10519_b0 , w_26697 );
and ( w_26696 ,  , w_26697 );
buf ( w_26695 , \10520_b1 );
not ( w_26695 , w_26698 );
not (  , w_26699 );
and ( w_26698 , w_26699 , \10520_b0 );
or ( \10522_b1 , \10521_b1 , w_26700 );
xor ( \10522_b0 , \10521_b0 , w_26702 );
not ( w_26702 , w_26703 );
and ( w_26703 , w_26700 , w_26701 );
buf ( w_26700 , \5898_b1 );
not ( w_26700 , w_26704 );
not ( w_26701 , w_26705 );
and ( w_26704 , w_26705 , \5898_b0 );
or ( \10523_b1 , \10518_b1 , \10522_b1 );
xor ( \10523_b0 , \10518_b0 , w_26706 );
not ( w_26706 , w_26707 );
and ( w_26707 , \10522_b1 , \10522_b0 );
or ( \10524_b1 , \6006_b1 , \5916_b1 );
not ( \5916_b1 , w_26708 );
and ( \10524_b0 , \6006_b0 , w_26709 );
and ( w_26708 , w_26709 , \5916_b0 );
or ( \10525_b1 , \6018_b1 , \5914_b1 );
not ( \5914_b1 , w_26710 );
and ( \10525_b0 , \6018_b0 , w_26711 );
and ( w_26710 , w_26711 , \5914_b0 );
or ( \10526_b1 , \10524_b1 , w_26713 );
not ( w_26713 , w_26714 );
and ( \10526_b0 , \10524_b0 , w_26715 );
and ( w_26714 ,  , w_26715 );
buf ( w_26713 , \10525_b1 );
not ( w_26713 , w_26716 );
not (  , w_26717 );
and ( w_26716 , w_26717 , \10525_b0 );
or ( \10527_b1 , \10526_b1 , w_26718 );
xor ( \10527_b0 , \10526_b0 , w_26720 );
not ( w_26720 , w_26721 );
and ( w_26721 , w_26718 , w_26719 );
buf ( w_26718 , \5923_b1 );
not ( w_26718 , w_26722 );
not ( w_26719 , w_26723 );
and ( w_26722 , w_26723 , \5923_b0 );
or ( \10528_b1 , \10523_b1 , \10527_b1 );
xor ( \10528_b0 , \10523_b0 , w_26724 );
not ( w_26724 , w_26725 );
and ( w_26725 , \10527_b1 , \10527_b0 );
or ( \10529_b1 , \10514_b1 , w_26726 );
xor ( \10529_b0 , \10514_b0 , w_26728 );
not ( w_26728 , w_26729 );
and ( w_26729 , w_26726 , w_26727 );
buf ( w_26726 , \10528_b1 );
not ( w_26726 , w_26730 );
not ( w_26727 , w_26731 );
and ( w_26730 , w_26731 , \10528_b0 );
or ( \10530_b1 , \10445_b1 , \10449_b1 );
not ( \10449_b1 , w_26732 );
and ( \10530_b0 , \10445_b0 , w_26733 );
and ( w_26732 , w_26733 , \10449_b0 );
or ( \10531_b1 , \10449_b1 , \10454_b1 );
not ( \10454_b1 , w_26734 );
and ( \10531_b0 , \10449_b0 , w_26735 );
and ( w_26734 , w_26735 , \10454_b0 );
or ( \10532_b1 , \10445_b1 , \10454_b1 );
not ( \10454_b1 , w_26736 );
and ( \10532_b0 , \10445_b0 , w_26737 );
and ( w_26736 , w_26737 , \10454_b0 );
or ( \10534_b1 , \10430_b1 , \10434_b1 );
not ( \10434_b1 , w_26738 );
and ( \10534_b0 , \10430_b0 , w_26739 );
and ( w_26738 , w_26739 , \10434_b0 );
or ( \10535_b1 , \10434_b1 , \10439_b1 );
not ( \10439_b1 , w_26740 );
and ( \10535_b0 , \10434_b0 , w_26741 );
and ( w_26740 , w_26741 , \10439_b0 );
or ( \10536_b1 , \10430_b1 , \10439_b1 );
not ( \10439_b1 , w_26742 );
and ( \10536_b0 , \10430_b0 , w_26743 );
and ( w_26742 , w_26743 , \10439_b0 );
or ( \10538_b1 , \10533_b1 , \10537_b1 );
xor ( \10538_b0 , \10533_b0 , w_26744 );
not ( w_26744 , w_26745 );
and ( w_26745 , \10537_b1 , \10537_b0 );
or ( \10539_b1 , \10421_b1 , \10425_b1 );
not ( \10425_b1 , w_26746 );
and ( \10539_b0 , \10421_b0 , w_26747 );
and ( w_26746 , w_26747 , \10425_b0 );
or ( \10540_b1 , \10538_b1 , \10539_b1 );
xor ( \10540_b0 , \10538_b0 , w_26748 );
not ( w_26748 , w_26749 );
and ( w_26749 , \10539_b1 , \10539_b0 );
or ( \10541_b1 , \10529_b1 , \10540_b1 );
xor ( \10541_b0 , \10529_b0 , w_26750 );
not ( w_26750 , w_26751 );
and ( w_26751 , \10540_b1 , \10540_b0 );
or ( \10542_b1 , \10405_b1 , \10409_b1 );
not ( \10409_b1 , w_26752 );
and ( \10542_b0 , \10405_b0 , w_26753 );
and ( w_26752 , w_26753 , \10409_b0 );
or ( \10543_b1 , \10409_b1 , \10414_b1 );
not ( \10414_b1 , w_26754 );
and ( \10543_b0 , \10409_b0 , w_26755 );
and ( w_26754 , w_26755 , \10414_b0 );
or ( \10544_b1 , \10405_b1 , \10414_b1 );
not ( \10414_b1 , w_26756 );
and ( \10544_b0 , \10405_b0 , w_26757 );
and ( w_26756 , w_26757 , \10414_b0 );
or ( \10546_b1 , \10393_b1 , \10397_b1 );
not ( \10397_b1 , w_26758 );
and ( \10546_b0 , \10393_b0 , w_26759 );
and ( w_26758 , w_26759 , \10397_b0 );
or ( \10547_b1 , \10397_b1 , \10402_b1 );
not ( \10402_b1 , w_26760 );
and ( \10547_b0 , \10397_b0 , w_26761 );
and ( w_26760 , w_26761 , \10402_b0 );
or ( \10548_b1 , \10393_b1 , \10402_b1 );
not ( \10402_b1 , w_26762 );
and ( \10548_b0 , \10393_b0 , w_26763 );
and ( w_26762 , w_26763 , \10402_b0 );
or ( \10550_b1 , \10545_b1 , \10549_b1 );
xor ( \10550_b0 , \10545_b0 , w_26764 );
not ( w_26764 , w_26765 );
and ( w_26765 , \10549_b1 , \10549_b0 );
or ( \10551_b1 , \10379_b1 , \10383_b1 );
not ( \10383_b1 , w_26766 );
and ( \10551_b0 , \10379_b0 , w_26767 );
and ( w_26766 , w_26767 , \10383_b0 );
or ( \10552_b1 , \10383_b1 , \10388_b1 );
not ( \10388_b1 , w_26768 );
and ( \10552_b0 , \10383_b0 , w_26769 );
and ( w_26768 , w_26769 , \10388_b0 );
or ( \10553_b1 , \10379_b1 , \10388_b1 );
not ( \10388_b1 , w_26770 );
and ( \10553_b0 , \10379_b0 , w_26771 );
and ( w_26770 , w_26771 , \10388_b0 );
or ( \10555_b1 , \10550_b1 , \10554_b1 );
xor ( \10555_b0 , \10550_b0 , w_26772 );
not ( w_26772 , w_26773 );
and ( w_26773 , \10554_b1 , \10554_b0 );
or ( \10556_b1 , \10541_b1 , \10555_b1 );
xor ( \10556_b0 , \10541_b0 , w_26774 );
not ( w_26774 , w_26775 );
and ( w_26775 , \10555_b1 , \10555_b0 );
or ( \10557_b1 , \10389_b1 , \10403_b1 );
not ( \10403_b1 , w_26776 );
and ( \10557_b0 , \10389_b0 , w_26777 );
and ( w_26776 , w_26777 , \10403_b0 );
or ( \10558_b1 , \10403_b1 , \10415_b1 );
not ( \10415_b1 , w_26778 );
and ( \10558_b0 , \10403_b0 , w_26779 );
and ( w_26778 , w_26779 , \10415_b0 );
or ( \10559_b1 , \10389_b1 , \10415_b1 );
not ( \10415_b1 , w_26780 );
and ( \10559_b0 , \10389_b0 , w_26781 );
and ( w_26780 , w_26781 , \10415_b0 );
or ( \10561_b1 , \5737_b1 , \7140_b1 );
not ( \7140_b1 , w_26782 );
and ( \10561_b0 , \5737_b0 , w_26783 );
and ( w_26782 , w_26783 , \7140_b0 );
buf ( \10562_b1 , \10561_b1 );
not ( \10562_b1 , w_26784 );
not ( \10562_b0 , w_26785 );
and ( w_26784 , w_26785 , \10561_b0 );
or ( \10563_b1 , \10562_b1 , w_26786 );
xor ( \10563_b0 , \10562_b0 , w_26788 );
not ( w_26788 , w_26789 );
and ( w_26789 , w_26786 , w_26787 );
buf ( w_26786 , \7146_b1 );
not ( w_26786 , w_26790 );
not ( w_26787 , w_26791 );
and ( w_26790 , w_26791 , \7146_b0 );
or ( \10564_b1 , \5984_b1 , \10563_b1 );
xor ( \10564_b0 , \5984_b0 , w_26792 );
not ( w_26792 , w_26793 );
and ( w_26793 , \10563_b1 , \10563_b0 );
or ( \10565_b1 , \5758_b1 , \7157_b1 );
not ( \7157_b1 , w_26794 );
and ( \10565_b0 , \5758_b0 , w_26795 );
and ( w_26794 , w_26795 , \7157_b0 );
or ( \10566_b1 , \5770_b1 , \7155_b1 );
not ( \7155_b1 , w_26796 );
and ( \10566_b0 , \5770_b0 , w_26797 );
and ( w_26796 , w_26797 , \7155_b0 );
or ( \10567_b1 , \10565_b1 , w_26799 );
not ( w_26799 , w_26800 );
and ( \10567_b0 , \10565_b0 , w_26801 );
and ( w_26800 ,  , w_26801 );
buf ( w_26799 , \10566_b1 );
not ( w_26799 , w_26802 );
not (  , w_26803 );
and ( w_26802 , w_26803 , \10566_b0 );
or ( \10568_b1 , \10567_b1 , w_26804 );
xor ( \10568_b0 , \10567_b0 , w_26806 );
not ( w_26806 , w_26807 );
and ( w_26807 , w_26804 , w_26805 );
buf ( w_26804 , \7163_b1 );
not ( w_26804 , w_26808 );
not ( w_26805 , w_26809 );
and ( w_26808 , w_26809 , \7163_b0 );
or ( \10569_b1 , \10564_b1 , \10568_b1 );
xor ( \10569_b0 , \10564_b0 , w_26810 );
not ( w_26810 , w_26811 );
and ( w_26811 , \10568_b1 , \10568_b0 );
or ( \10570_b1 , \10560_b1 , \10569_b1 );
xor ( \10570_b0 , \10560_b0 , w_26812 );
not ( w_26812 , w_26813 );
and ( w_26813 , \10569_b1 , \10569_b0 );
or ( \10571_b1 , \5906_b1 , \5809_b1 );
not ( \5809_b1 , w_26814 );
and ( \10571_b0 , \5906_b0 , w_26815 );
and ( w_26814 , w_26815 , \5809_b0 );
or ( \10572_b1 , \5918_b1 , \5807_b1 );
not ( \5807_b1 , w_26816 );
and ( \10572_b0 , \5918_b0 , w_26817 );
and ( w_26816 , w_26817 , \5807_b0 );
or ( \10573_b1 , \10571_b1 , w_26819 );
not ( w_26819 , w_26820 );
and ( \10573_b0 , \10571_b0 , w_26821 );
and ( w_26820 ,  , w_26821 );
buf ( w_26819 , \10572_b1 );
not ( w_26819 , w_26822 );
not (  , w_26823 );
and ( w_26822 , w_26823 , \10572_b0 );
or ( \10574_b1 , \10573_b1 , w_26824 );
xor ( \10574_b0 , \10573_b0 , w_26826 );
not ( w_26826 , w_26827 );
and ( w_26827 , w_26824 , w_26825 );
buf ( w_26824 , \5816_b1 );
not ( w_26824 , w_26828 );
not ( w_26825 , w_26829 );
and ( w_26828 , w_26829 , \5816_b0 );
or ( \10575_b1 , \5925_b1 , \5829_b1 );
not ( \5829_b1 , w_26830 );
and ( \10575_b0 , \5925_b0 , w_26831 );
and ( w_26830 , w_26831 , \5829_b0 );
or ( \10576_b1 , \5937_b1 , \5827_b1 );
not ( \5827_b1 , w_26832 );
and ( \10576_b0 , \5937_b0 , w_26833 );
and ( w_26832 , w_26833 , \5827_b0 );
or ( \10577_b1 , \10575_b1 , w_26835 );
not ( w_26835 , w_26836 );
and ( \10577_b0 , \10575_b0 , w_26837 );
and ( w_26836 ,  , w_26837 );
buf ( w_26835 , \10576_b1 );
not ( w_26835 , w_26838 );
not (  , w_26839 );
and ( w_26838 , w_26839 , \10576_b0 );
or ( \10578_b1 , \10577_b1 , w_26840 );
xor ( \10578_b0 , \10577_b0 , w_26842 );
not ( w_26842 , w_26843 );
and ( w_26843 , w_26840 , w_26841 );
buf ( w_26840 , \5836_b1 );
not ( w_26840 , w_26844 );
not ( w_26841 , w_26845 );
and ( w_26844 , w_26845 , \5836_b0 );
or ( \10579_b1 , \10574_b1 , \10578_b1 );
xor ( \10579_b0 , \10574_b0 , w_26846 );
not ( w_26846 , w_26847 );
and ( w_26847 , \10578_b1 , \10578_b0 );
or ( \10580_b1 , \5945_b1 , \5852_b1 );
not ( \5852_b1 , w_26848 );
and ( \10580_b0 , \5945_b0 , w_26849 );
and ( w_26848 , w_26849 , \5852_b0 );
or ( \10581_b1 , \5957_b1 , \5850_b1 );
not ( \5850_b1 , w_26850 );
and ( \10581_b0 , \5957_b0 , w_26851 );
and ( w_26850 , w_26851 , \5850_b0 );
or ( \10582_b1 , \10580_b1 , w_26853 );
not ( w_26853 , w_26854 );
and ( \10582_b0 , \10580_b0 , w_26855 );
and ( w_26854 ,  , w_26855 );
buf ( w_26853 , \10581_b1 );
not ( w_26853 , w_26856 );
not (  , w_26857 );
and ( w_26856 , w_26857 , \10581_b0 );
or ( \10583_b1 , \10582_b1 , w_26858 );
xor ( \10583_b0 , \10582_b0 , w_26860 );
not ( w_26860 , w_26861 );
and ( w_26861 , w_26858 , w_26859 );
buf ( w_26858 , \5859_b1 );
not ( w_26858 , w_26862 );
not ( w_26859 , w_26863 );
and ( w_26862 , w_26863 , \5859_b0 );
or ( \10584_b1 , \10579_b1 , \10583_b1 );
xor ( \10584_b0 , \10579_b0 , w_26864 );
not ( w_26864 , w_26865 );
and ( w_26865 , \10583_b1 , \10583_b0 );
or ( \10585_b1 , \5842_b1 , \5750_b1 );
not ( \5750_b1 , w_26866 );
and ( \10585_b0 , \5842_b0 , w_26867 );
and ( w_26866 , w_26867 , \5750_b0 );
or ( \10586_b1 , \5854_b1 , \5748_b1 );
not ( \5748_b1 , w_26868 );
and ( \10586_b0 , \5854_b0 , w_26869 );
and ( w_26868 , w_26869 , \5748_b0 );
or ( \10587_b1 , \10585_b1 , w_26871 );
not ( w_26871 , w_26872 );
and ( \10587_b0 , \10585_b0 , w_26873 );
and ( w_26872 ,  , w_26873 );
buf ( w_26871 , \10586_b1 );
not ( w_26871 , w_26874 );
not (  , w_26875 );
and ( w_26874 , w_26875 , \10586_b0 );
or ( \10588_b1 , \10587_b1 , w_26876 );
xor ( \10588_b0 , \10587_b0 , w_26878 );
not ( w_26878 , w_26879 );
and ( w_26879 , w_26876 , w_26877 );
buf ( w_26876 , \5755_b1 );
not ( w_26876 , w_26880 );
not ( w_26877 , w_26881 );
and ( w_26880 , w_26881 , \5755_b0 );
or ( \10589_b1 , \5861_b1 , \5768_b1 );
not ( \5768_b1 , w_26882 );
and ( \10589_b0 , \5861_b0 , w_26883 );
and ( w_26882 , w_26883 , \5768_b0 );
or ( \10590_b1 , \5873_b1 , \5766_b1 );
not ( \5766_b1 , w_26884 );
and ( \10590_b0 , \5873_b0 , w_26885 );
and ( w_26884 , w_26885 , \5766_b0 );
or ( \10591_b1 , \10589_b1 , w_26887 );
not ( w_26887 , w_26888 );
and ( \10591_b0 , \10589_b0 , w_26889 );
and ( w_26888 ,  , w_26889 );
buf ( w_26887 , \10590_b1 );
not ( w_26887 , w_26890 );
not (  , w_26891 );
and ( w_26890 , w_26891 , \10590_b0 );
or ( \10592_b1 , \10591_b1 , w_26892 );
xor ( \10592_b0 , \10591_b0 , w_26894 );
not ( w_26894 , w_26895 );
and ( w_26895 , w_26892 , w_26893 );
buf ( w_26892 , \5775_b1 );
not ( w_26892 , w_26896 );
not ( w_26893 , w_26897 );
and ( w_26896 , w_26897 , \5775_b0 );
or ( \10593_b1 , \10588_b1 , \10592_b1 );
xor ( \10593_b0 , \10588_b0 , w_26898 );
not ( w_26898 , w_26899 );
and ( w_26899 , \10592_b1 , \10592_b0 );
or ( \10594_b1 , \5881_b1 , \5790_b1 );
not ( \5790_b1 , w_26900 );
and ( \10594_b0 , \5881_b0 , w_26901 );
and ( w_26900 , w_26901 , \5790_b0 );
or ( \10595_b1 , \5893_b1 , \5788_b1 );
not ( \5788_b1 , w_26902 );
and ( \10595_b0 , \5893_b0 , w_26903 );
and ( w_26902 , w_26903 , \5788_b0 );
or ( \10596_b1 , \10594_b1 , w_26905 );
not ( w_26905 , w_26906 );
and ( \10596_b0 , \10594_b0 , w_26907 );
and ( w_26906 ,  , w_26907 );
buf ( w_26905 , \10595_b1 );
not ( w_26905 , w_26908 );
not (  , w_26909 );
and ( w_26908 , w_26909 , \10595_b0 );
or ( \10597_b1 , \10596_b1 , w_26910 );
xor ( \10597_b0 , \10596_b0 , w_26912 );
not ( w_26912 , w_26913 );
and ( w_26913 , w_26910 , w_26911 );
buf ( w_26910 , \5797_b1 );
not ( w_26910 , w_26914 );
not ( w_26911 , w_26915 );
and ( w_26914 , w_26915 , \5797_b0 );
or ( \10598_b1 , \10593_b1 , \10597_b1 );
xor ( \10598_b0 , \10593_b0 , w_26916 );
not ( w_26916 , w_26917 );
and ( w_26917 , \10597_b1 , \10597_b0 );
or ( \10599_b1 , \10584_b1 , \10598_b1 );
xor ( \10599_b0 , \10584_b0 , w_26918 );
not ( w_26918 , w_26919 );
and ( w_26919 , \10598_b1 , \10598_b0 );
or ( \10600_b1 , \5780_b1 , \7175_b1 );
not ( \7175_b1 , w_26920 );
and ( \10600_b0 , \5780_b0 , w_26921 );
and ( w_26920 , w_26921 , \7175_b0 );
or ( \10601_b1 , \5792_b1 , \7173_b1 );
not ( \7173_b1 , w_26922 );
and ( \10601_b0 , \5792_b0 , w_26923 );
and ( w_26922 , w_26923 , \7173_b0 );
or ( \10602_b1 , \10600_b1 , w_26925 );
not ( w_26925 , w_26926 );
and ( \10602_b0 , \10600_b0 , w_26927 );
and ( w_26926 ,  , w_26927 );
buf ( w_26925 , \10601_b1 );
not ( w_26925 , w_26928 );
not (  , w_26929 );
and ( w_26928 , w_26929 , \10601_b0 );
or ( \10603_b1 , \10602_b1 , w_26930 );
xor ( \10603_b0 , \10602_b0 , w_26932 );
not ( w_26932 , w_26933 );
and ( w_26933 , w_26930 , w_26931 );
buf ( w_26930 , \7181_b1 );
not ( w_26930 , w_26934 );
not ( w_26931 , w_26935 );
and ( w_26934 , w_26935 , \7181_b0 );
or ( \10604_b1 , \5799_b1 , \7192_b1 );
not ( \7192_b1 , w_26936 );
and ( \10604_b0 , \5799_b0 , w_26937 );
and ( w_26936 , w_26937 , \7192_b0 );
or ( \10605_b1 , \5811_b1 , \7190_b1 );
not ( \7190_b1 , w_26938 );
and ( \10605_b0 , \5811_b0 , w_26939 );
and ( w_26938 , w_26939 , \7190_b0 );
or ( \10606_b1 , \10604_b1 , w_26941 );
not ( w_26941 , w_26942 );
and ( \10606_b0 , \10604_b0 , w_26943 );
and ( w_26942 ,  , w_26943 );
buf ( w_26941 , \10605_b1 );
not ( w_26941 , w_26944 );
not (  , w_26945 );
and ( w_26944 , w_26945 , \10605_b0 );
or ( \10607_b1 , \10606_b1 , w_26946 );
xor ( \10607_b0 , \10606_b0 , w_26948 );
not ( w_26948 , w_26949 );
and ( w_26949 , w_26946 , w_26947 );
buf ( w_26946 , \7198_b1 );
not ( w_26946 , w_26950 );
not ( w_26947 , w_26951 );
and ( w_26950 , w_26951 , \7198_b0 );
or ( \10608_b1 , \10603_b1 , \10607_b1 );
xor ( \10608_b0 , \10603_b0 , w_26952 );
not ( w_26952 , w_26953 );
and ( w_26953 , \10607_b1 , \10607_b0 );
or ( \10609_b1 , \5819_b1 , \7203_b1 );
not ( \7203_b1 , w_26954 );
and ( \10609_b0 , \5819_b0 , w_26955 );
and ( w_26954 , w_26955 , \7203_b0 );
or ( \10610_b1 , \5831_b1 , \7201_b1 );
not ( \7201_b1 , w_26956 );
and ( \10610_b0 , \5831_b0 , w_26957 );
and ( w_26956 , w_26957 , \7201_b0 );
or ( \10611_b1 , \10609_b1 , w_26959 );
not ( w_26959 , w_26960 );
and ( \10611_b0 , \10609_b0 , w_26961 );
and ( w_26960 ,  , w_26961 );
buf ( w_26959 , \10610_b1 );
not ( w_26959 , w_26962 );
not (  , w_26963 );
and ( w_26962 , w_26963 , \10610_b0 );
or ( \10612_b1 , \10611_b1 , w_26964 );
xor ( \10612_b0 , \10611_b0 , w_26966 );
not ( w_26966 , w_26967 );
and ( w_26967 , w_26964 , w_26965 );
buf ( w_26964 , \6824_b1 );
not ( w_26964 , w_26968 );
not ( w_26965 , w_26969 );
and ( w_26968 , w_26969 , \6824_b0 );
or ( \10613_b1 , \10608_b1 , \10612_b1 );
xor ( \10613_b0 , \10608_b0 , w_26970 );
not ( w_26970 , w_26971 );
and ( w_26971 , \10612_b1 , \10612_b0 );
or ( \10614_b1 , \10599_b1 , \10613_b1 );
xor ( \10614_b0 , \10599_b0 , w_26972 );
not ( w_26972 , w_26973 );
and ( w_26973 , \10613_b1 , \10613_b0 );
or ( \10615_b1 , \10570_b1 , \10614_b1 );
xor ( \10615_b0 , \10570_b0 , w_26974 );
not ( w_26974 , w_26975 );
and ( w_26975 , \10614_b1 , \10614_b0 );
or ( \10616_b1 , \10556_b1 , \10615_b1 );
xor ( \10616_b0 , \10556_b0 , w_26976 );
not ( w_26976 , w_26977 );
and ( w_26977 , \10615_b1 , \10615_b0 );
or ( \10617_b1 , \10360_b1 , \10364_b1 );
not ( \10364_b1 , w_26978 );
and ( \10617_b0 , \10360_b0 , w_26979 );
and ( w_26978 , w_26979 , \10364_b0 );
or ( \10618_b1 , \10364_b1 , \10369_b1 );
not ( \10369_b1 , w_26980 );
and ( \10618_b0 , \10364_b0 , w_26981 );
and ( w_26980 , w_26981 , \10369_b0 );
or ( \10619_b1 , \10360_b1 , \10369_b1 );
not ( \10369_b1 , w_26982 );
and ( \10619_b0 , \10360_b0 , w_26983 );
and ( w_26982 , w_26983 , \10369_b0 );
or ( \10621_b1 , \10346_b1 , \10350_b1 );
not ( \10350_b1 , w_26984 );
and ( \10621_b0 , \10346_b0 , w_26985 );
and ( w_26984 , w_26985 , \10350_b0 );
or ( \10622_b1 , \10350_b1 , \10355_b1 );
not ( \10355_b1 , w_26986 );
and ( \10622_b0 , \10350_b0 , w_26987 );
and ( w_26986 , w_26987 , \10355_b0 );
or ( \10623_b1 , \10346_b1 , \10355_b1 );
not ( \10355_b1 , w_26988 );
and ( \10623_b0 , \10346_b0 , w_26989 );
and ( w_26988 , w_26989 , \10355_b0 );
or ( \10625_b1 , \10620_b1 , \10624_b1 );
xor ( \10625_b0 , \10620_b0 , w_26990 );
not ( w_26990 , w_26991 );
and ( w_26991 , \10624_b1 , \10624_b0 );
or ( \10626_b1 , \10426_b1 , \10440_b1 );
not ( \10440_b1 , w_26992 );
and ( \10626_b0 , \10426_b0 , w_26993 );
and ( w_26992 , w_26993 , \10440_b0 );
or ( \10627_b1 , \10440_b1 , \10455_b1 );
not ( \10455_b1 , w_26994 );
and ( \10627_b0 , \10440_b0 , w_26995 );
and ( w_26994 , w_26995 , \10455_b0 );
or ( \10628_b1 , \10426_b1 , \10455_b1 );
not ( \10455_b1 , w_26996 );
and ( \10628_b0 , \10426_b0 , w_26997 );
and ( w_26996 , w_26997 , \10455_b0 );
or ( \10630_b1 , \10625_b1 , \10629_b1 );
xor ( \10630_b0 , \10625_b0 , w_26998 );
not ( w_26998 , w_26999 );
and ( w_26999 , \10629_b1 , \10629_b0 );
or ( \10631_b1 , \10616_b1 , \10630_b1 );
xor ( \10631_b0 , \10616_b0 , w_27000 );
not ( w_27000 , w_27001 );
and ( w_27001 , \10630_b1 , \10630_b0 );
or ( \10632_b1 , \10502_b1 , \10631_b1 );
xor ( \10632_b0 , \10502_b0 , w_27002 );
not ( w_27002 , w_27003 );
and ( w_27003 , \10631_b1 , \10631_b0 );
or ( \10633_b1 , \10493_b1 , \10632_b1 );
xor ( \10633_b0 , \10493_b0 , w_27004 );
not ( w_27004 , w_27005 );
and ( w_27005 , \10632_b1 , \10632_b0 );
or ( \10634_b1 , \10318_b1 , \10332_b1 );
not ( \10332_b1 , w_27006 );
and ( \10634_b0 , \10318_b0 , w_27007 );
and ( w_27006 , w_27007 , \10332_b0 );
or ( \10635_b1 , \10332_b1 , \10471_b1 );
not ( \10471_b1 , w_27008 );
and ( \10635_b0 , \10332_b0 , w_27009 );
and ( w_27008 , w_27009 , \10471_b0 );
or ( \10636_b1 , \10318_b1 , \10471_b1 );
not ( \10471_b1 , w_27010 );
and ( \10636_b0 , \10318_b0 , w_27011 );
and ( w_27010 , w_27011 , \10471_b0 );
or ( \10638_b1 , \10633_b1 , w_27013 );
not ( w_27013 , w_27014 );
and ( \10638_b0 , \10633_b0 , w_27015 );
and ( w_27014 ,  , w_27015 );
buf ( w_27013 , \10637_b1 );
not ( w_27013 , w_27016 );
not (  , w_27017 );
and ( w_27016 , w_27017 , \10637_b0 );
or ( \10639_b1 , \10477_b1 , w_27019 );
not ( w_27019 , w_27020 );
and ( \10639_b0 , \10477_b0 , w_27021 );
and ( w_27020 ,  , w_27021 );
buf ( w_27019 , \10638_b1 );
not ( w_27019 , w_27022 );
not (  , w_27023 );
and ( w_27022 , w_27023 , \10638_b0 );
or ( \10640_b1 , \10497_b1 , \10501_b1 );
not ( \10501_b1 , w_27024 );
and ( \10640_b0 , \10497_b0 , w_27025 );
and ( w_27024 , w_27025 , \10501_b0 );
or ( \10641_b1 , \10501_b1 , \10631_b1 );
not ( \10631_b1 , w_27026 );
and ( \10641_b0 , \10501_b0 , w_27027 );
and ( w_27026 , w_27027 , \10631_b0 );
or ( \10642_b1 , \10497_b1 , \10631_b1 );
not ( \10631_b1 , w_27028 );
and ( \10642_b0 , \10497_b0 , w_27029 );
and ( w_27028 , w_27029 , \10631_b0 );
or ( \10644_b1 , \10620_b1 , \10624_b1 );
not ( \10624_b1 , w_27030 );
and ( \10644_b0 , \10620_b0 , w_27031 );
and ( w_27030 , w_27031 , \10624_b0 );
or ( \10645_b1 , \10624_b1 , \10629_b1 );
not ( \10629_b1 , w_27032 );
and ( \10645_b0 , \10624_b0 , w_27033 );
and ( w_27032 , w_27033 , \10629_b0 );
or ( \10646_b1 , \10620_b1 , \10629_b1 );
not ( \10629_b1 , w_27034 );
and ( \10646_b0 , \10620_b0 , w_27035 );
and ( w_27034 , w_27035 , \10629_b0 );
or ( \10648_b1 , \10560_b1 , \10569_b1 );
not ( \10569_b1 , w_27036 );
and ( \10648_b0 , \10560_b0 , w_27037 );
and ( w_27036 , w_27037 , \10569_b0 );
or ( \10649_b1 , \10569_b1 , \10614_b1 );
not ( \10614_b1 , w_27038 );
and ( \10649_b0 , \10569_b0 , w_27039 );
and ( w_27038 , w_27039 , \10614_b0 );
or ( \10650_b1 , \10560_b1 , \10614_b1 );
not ( \10614_b1 , w_27040 );
and ( \10650_b0 , \10560_b0 , w_27041 );
and ( w_27040 , w_27041 , \10614_b0 );
or ( \10652_b1 , \10647_b1 , \10651_b1 );
xor ( \10652_b0 , \10647_b0 , w_27042 );
not ( w_27042 , w_27043 );
and ( w_27043 , \10651_b1 , \10651_b0 );
or ( \10653_b1 , \10529_b1 , \10540_b1 );
not ( \10540_b1 , w_27044 );
and ( \10653_b0 , \10529_b0 , w_27045 );
and ( w_27044 , w_27045 , \10540_b0 );
or ( \10654_b1 , \10540_b1 , \10555_b1 );
not ( \10555_b1 , w_27046 );
and ( \10654_b0 , \10540_b0 , w_27047 );
and ( w_27046 , w_27047 , \10555_b0 );
or ( \10655_b1 , \10529_b1 , \10555_b1 );
not ( \10555_b1 , w_27048 );
and ( \10655_b0 , \10529_b0 , w_27049 );
and ( w_27048 , w_27049 , \10555_b0 );
or ( \10657_b1 , \10652_b1 , \10656_b1 );
xor ( \10657_b0 , \10652_b0 , w_27050 );
not ( w_27050 , w_27051 );
and ( w_27051 , \10656_b1 , \10656_b0 );
or ( \10658_b1 , \10643_b1 , \10657_b1 );
xor ( \10658_b0 , \10643_b0 , w_27052 );
not ( w_27052 , w_27053 );
and ( w_27053 , \10657_b1 , \10657_b0 );
or ( \10659_b1 , \10485_b1 , \10489_b1 );
not ( \10489_b1 , w_27054 );
and ( \10659_b0 , \10485_b0 , w_27055 );
and ( w_27054 , w_27055 , \10489_b0 );
or ( \10660_b1 , \10489_b1 , \10491_b1 );
not ( \10491_b1 , w_27056 );
and ( \10660_b0 , \10489_b0 , w_27057 );
and ( w_27056 , w_27057 , \10491_b0 );
or ( \10661_b1 , \10485_b1 , \10491_b1 );
not ( \10491_b1 , w_27058 );
and ( \10661_b0 , \10485_b0 , w_27059 );
and ( w_27058 , w_27059 , \10491_b0 );
or ( \10663_b1 , \10556_b1 , \10615_b1 );
not ( \10615_b1 , w_27060 );
and ( \10663_b0 , \10556_b0 , w_27061 );
and ( w_27060 , w_27061 , \10615_b0 );
or ( \10664_b1 , \10615_b1 , \10630_b1 );
not ( \10630_b1 , w_27062 );
and ( \10664_b0 , \10615_b0 , w_27063 );
and ( w_27062 , w_27063 , \10630_b0 );
or ( \10665_b1 , \10556_b1 , \10630_b1 );
not ( \10630_b1 , w_27064 );
and ( \10665_b0 , \10556_b0 , w_27065 );
and ( w_27064 , w_27065 , \10630_b0 );
or ( \10667_b1 , \10662_b1 , \10666_b1 );
xor ( \10667_b0 , \10662_b0 , w_27066 );
not ( w_27066 , w_27067 );
and ( w_27067 , \10666_b1 , \10666_b0 );
or ( \10668_b1 , \10574_b1 , \10578_b1 );
not ( \10578_b1 , w_27068 );
and ( \10668_b0 , \10574_b0 , w_27069 );
and ( w_27068 , w_27069 , \10578_b0 );
or ( \10669_b1 , \10578_b1 , \10583_b1 );
not ( \10583_b1 , w_27070 );
and ( \10669_b0 , \10578_b0 , w_27071 );
and ( w_27070 , w_27071 , \10583_b0 );
or ( \10670_b1 , \10574_b1 , \10583_b1 );
not ( \10583_b1 , w_27072 );
and ( \10670_b0 , \10574_b0 , w_27073 );
and ( w_27072 , w_27073 , \10583_b0 );
or ( \10672_b1 , \10518_b1 , \10522_b1 );
not ( \10522_b1 , w_27074 );
and ( \10672_b0 , \10518_b0 , w_27075 );
and ( w_27074 , w_27075 , \10522_b0 );
or ( \10673_b1 , \10522_b1 , \10527_b1 );
not ( \10527_b1 , w_27076 );
and ( \10673_b0 , \10522_b0 , w_27077 );
and ( w_27076 , w_27077 , \10527_b0 );
or ( \10674_b1 , \10518_b1 , \10527_b1 );
not ( \10527_b1 , w_27078 );
and ( \10674_b0 , \10518_b0 , w_27079 );
and ( w_27078 , w_27079 , \10527_b0 );
or ( \10676_b1 , \10671_b1 , \10675_b1 );
xor ( \10676_b0 , \10671_b0 , w_27080 );
not ( w_27080 , w_27081 );
and ( w_27081 , \10675_b1 , \10675_b0 );
or ( \10677_b1 , \10506_b1 , \10510_b1 );
not ( \10510_b1 , w_27082 );
and ( \10677_b0 , \10506_b0 , w_27083 );
and ( w_27082 , w_27083 , \10510_b0 );
or ( \10678_b1 , \10510_b1 , \10513_b1 );
not ( \10513_b1 , w_27084 );
and ( \10678_b0 , \10510_b0 , w_27085 );
and ( w_27084 , w_27085 , \10513_b0 );
or ( \10679_b1 , \10506_b1 , \10513_b1 );
not ( \10513_b1 , w_27086 );
and ( \10679_b0 , \10506_b0 , w_27087 );
and ( w_27086 , w_27087 , \10513_b0 );
or ( \10681_b1 , \10676_b1 , \10680_b1 );
xor ( \10681_b0 , \10676_b0 , w_27088 );
not ( w_27088 , w_27089 );
and ( w_27089 , \10680_b1 , \10680_b0 );
or ( \10682_b1 , \5984_b1 , \10563_b1 );
not ( \10563_b1 , w_27090 );
and ( \10682_b0 , \5984_b0 , w_27091 );
and ( w_27090 , w_27091 , \10563_b0 );
or ( \10683_b1 , \10563_b1 , \10568_b1 );
not ( \10568_b1 , w_27092 );
and ( \10683_b0 , \10563_b0 , w_27093 );
and ( w_27092 , w_27093 , \10568_b0 );
or ( \10684_b1 , \5984_b1 , \10568_b1 );
not ( \10568_b1 , w_27094 );
and ( \10684_b0 , \5984_b0 , w_27095 );
and ( w_27094 , w_27095 , \10568_b0 );
or ( \10686_b1 , \10603_b1 , \10607_b1 );
not ( \10607_b1 , w_27096 );
and ( \10686_b0 , \10603_b0 , w_27097 );
and ( w_27096 , w_27097 , \10607_b0 );
or ( \10687_b1 , \10607_b1 , \10612_b1 );
not ( \10612_b1 , w_27098 );
and ( \10687_b0 , \10607_b0 , w_27099 );
and ( w_27098 , w_27099 , \10612_b0 );
or ( \10688_b1 , \10603_b1 , \10612_b1 );
not ( \10612_b1 , w_27100 );
and ( \10688_b0 , \10603_b0 , w_27101 );
and ( w_27100 , w_27101 , \10612_b0 );
or ( \10690_b1 , \10685_b1 , \10689_b1 );
xor ( \10690_b0 , \10685_b0 , w_27102 );
not ( w_27102 , w_27103 );
and ( w_27103 , \10689_b1 , \10689_b0 );
or ( \10691_b1 , \10588_b1 , \10592_b1 );
not ( \10592_b1 , w_27104 );
and ( \10691_b0 , \10588_b0 , w_27105 );
and ( w_27104 , w_27105 , \10592_b0 );
or ( \10692_b1 , \10592_b1 , \10597_b1 );
not ( \10597_b1 , w_27106 );
and ( \10692_b0 , \10592_b0 , w_27107 );
and ( w_27106 , w_27107 , \10597_b0 );
or ( \10693_b1 , \10588_b1 , \10597_b1 );
not ( \10597_b1 , w_27108 );
and ( \10693_b0 , \10588_b0 , w_27109 );
and ( w_27108 , w_27109 , \10597_b0 );
or ( \10695_b1 , \10690_b1 , \10694_b1 );
xor ( \10695_b0 , \10690_b0 , w_27110 );
not ( w_27110 , w_27111 );
and ( w_27111 , \10694_b1 , \10694_b0 );
or ( \10696_b1 , \10681_b1 , \10695_b1 );
xor ( \10696_b0 , \10681_b0 , w_27112 );
not ( w_27112 , w_27113 );
and ( w_27113 , \10695_b1 , \10695_b0 );
or ( \10697_b1 , \10584_b1 , \10598_b1 );
not ( \10598_b1 , w_27114 );
and ( \10697_b0 , \10584_b0 , w_27115 );
and ( w_27114 , w_27115 , \10598_b0 );
or ( \10698_b1 , \10598_b1 , \10613_b1 );
not ( \10613_b1 , w_27116 );
and ( \10698_b0 , \10598_b0 , w_27117 );
and ( w_27116 , w_27117 , \10613_b0 );
or ( \10699_b1 , \10584_b1 , \10613_b1 );
not ( \10613_b1 , w_27118 );
and ( \10699_b0 , \10584_b0 , w_27119 );
and ( w_27118 , w_27119 , \10613_b0 );
or ( \10701_b1 , \5873_b1 , \5768_b1 );
not ( \5768_b1 , w_27120 );
and ( \10701_b0 , \5873_b0 , w_27121 );
and ( w_27120 , w_27121 , \5768_b0 );
or ( \10702_b1 , \5842_b1 , \5766_b1 );
not ( \5766_b1 , w_27122 );
and ( \10702_b0 , \5842_b0 , w_27123 );
and ( w_27122 , w_27123 , \5766_b0 );
or ( \10703_b1 , \10701_b1 , w_27125 );
not ( w_27125 , w_27126 );
and ( \10703_b0 , \10701_b0 , w_27127 );
and ( w_27126 ,  , w_27127 );
buf ( w_27125 , \10702_b1 );
not ( w_27125 , w_27128 );
not (  , w_27129 );
and ( w_27128 , w_27129 , \10702_b0 );
or ( \10704_b1 , \10703_b1 , w_27130 );
xor ( \10704_b0 , \10703_b0 , w_27132 );
not ( w_27132 , w_27133 );
and ( w_27133 , w_27130 , w_27131 );
buf ( w_27130 , \5775_b1 );
not ( w_27130 , w_27134 );
not ( w_27131 , w_27135 );
and ( w_27134 , w_27135 , \5775_b0 );
or ( \10705_b1 , \5893_b1 , \5790_b1 );
not ( \5790_b1 , w_27136 );
and ( \10705_b0 , \5893_b0 , w_27137 );
and ( w_27136 , w_27137 , \5790_b0 );
or ( \10706_b1 , \5861_b1 , \5788_b1 );
not ( \5788_b1 , w_27138 );
and ( \10706_b0 , \5861_b0 , w_27139 );
and ( w_27138 , w_27139 , \5788_b0 );
or ( \10707_b1 , \10705_b1 , w_27141 );
not ( w_27141 , w_27142 );
and ( \10707_b0 , \10705_b0 , w_27143 );
and ( w_27142 ,  , w_27143 );
buf ( w_27141 , \10706_b1 );
not ( w_27141 , w_27144 );
not (  , w_27145 );
and ( w_27144 , w_27145 , \10706_b0 );
or ( \10708_b1 , \10707_b1 , w_27146 );
xor ( \10708_b0 , \10707_b0 , w_27148 );
not ( w_27148 , w_27149 );
and ( w_27149 , w_27146 , w_27147 );
buf ( w_27146 , \5797_b1 );
not ( w_27146 , w_27150 );
not ( w_27147 , w_27151 );
and ( w_27150 , w_27151 , \5797_b0 );
or ( \10709_b1 , \10704_b1 , \10708_b1 );
xor ( \10709_b0 , \10704_b0 , w_27152 );
not ( w_27152 , w_27153 );
and ( w_27153 , \10708_b1 , \10708_b0 );
or ( \10710_b1 , \5918_b1 , \5809_b1 );
not ( \5809_b1 , w_27154 );
and ( \10710_b0 , \5918_b0 , w_27155 );
and ( w_27154 , w_27155 , \5809_b0 );
or ( \10711_b1 , \5881_b1 , \5807_b1 );
not ( \5807_b1 , w_27156 );
and ( \10711_b0 , \5881_b0 , w_27157 );
and ( w_27156 , w_27157 , \5807_b0 );
or ( \10712_b1 , \10710_b1 , w_27159 );
not ( w_27159 , w_27160 );
and ( \10712_b0 , \10710_b0 , w_27161 );
and ( w_27160 ,  , w_27161 );
buf ( w_27159 , \10711_b1 );
not ( w_27159 , w_27162 );
not (  , w_27163 );
and ( w_27162 , w_27163 , \10711_b0 );
or ( \10713_b1 , \10712_b1 , w_27164 );
xor ( \10713_b0 , \10712_b0 , w_27166 );
not ( w_27166 , w_27167 );
and ( w_27167 , w_27164 , w_27165 );
buf ( w_27164 , \5816_b1 );
not ( w_27164 , w_27168 );
not ( w_27165 , w_27169 );
and ( w_27168 , w_27169 , \5816_b0 );
or ( \10714_b1 , \10709_b1 , \10713_b1 );
xor ( \10714_b0 , \10709_b0 , w_27170 );
not ( w_27170 , w_27171 );
and ( w_27171 , \10713_b1 , \10713_b0 );
or ( \10715_b1 , \5811_b1 , \7192_b1 );
not ( \7192_b1 , w_27172 );
and ( \10715_b0 , \5811_b0 , w_27173 );
and ( w_27172 , w_27173 , \7192_b0 );
or ( \10716_b1 , \5780_b1 , \7190_b1 );
not ( \7190_b1 , w_27174 );
and ( \10716_b0 , \5780_b0 , w_27175 );
and ( w_27174 , w_27175 , \7190_b0 );
or ( \10717_b1 , \10715_b1 , w_27177 );
not ( w_27177 , w_27178 );
and ( \10717_b0 , \10715_b0 , w_27179 );
and ( w_27178 ,  , w_27179 );
buf ( w_27177 , \10716_b1 );
not ( w_27177 , w_27180 );
not (  , w_27181 );
and ( w_27180 , w_27181 , \10716_b0 );
or ( \10718_b1 , \10717_b1 , w_27182 );
xor ( \10718_b0 , \10717_b0 , w_27184 );
not ( w_27184 , w_27185 );
and ( w_27185 , w_27182 , w_27183 );
buf ( w_27182 , \7198_b1 );
not ( w_27182 , w_27186 );
not ( w_27183 , w_27187 );
and ( w_27186 , w_27187 , \7198_b0 );
or ( \10719_b1 , \5831_b1 , \7203_b1 );
not ( \7203_b1 , w_27188 );
and ( \10719_b0 , \5831_b0 , w_27189 );
and ( w_27188 , w_27189 , \7203_b0 );
or ( \10720_b1 , \5799_b1 , \7201_b1 );
not ( \7201_b1 , w_27190 );
and ( \10720_b0 , \5799_b0 , w_27191 );
and ( w_27190 , w_27191 , \7201_b0 );
or ( \10721_b1 , \10719_b1 , w_27193 );
not ( w_27193 , w_27194 );
and ( \10721_b0 , \10719_b0 , w_27195 );
and ( w_27194 ,  , w_27195 );
buf ( w_27193 , \10720_b1 );
not ( w_27193 , w_27196 );
not (  , w_27197 );
and ( w_27196 , w_27197 , \10720_b0 );
or ( \10722_b1 , \10721_b1 , w_27198 );
xor ( \10722_b0 , \10721_b0 , w_27200 );
not ( w_27200 , w_27201 );
and ( w_27201 , w_27198 , w_27199 );
buf ( w_27198 , \6824_b1 );
not ( w_27198 , w_27202 );
not ( w_27199 , w_27203 );
and ( w_27202 , w_27203 , \6824_b0 );
or ( \10723_b1 , \10718_b1 , \10722_b1 );
xor ( \10723_b0 , \10718_b0 , w_27204 );
not ( w_27204 , w_27205 );
and ( w_27205 , \10722_b1 , \10722_b0 );
or ( \10724_b1 , \5854_b1 , \5750_b1 );
not ( \5750_b1 , w_27206 );
and ( \10724_b0 , \5854_b0 , w_27207 );
and ( w_27206 , w_27207 , \5750_b0 );
or ( \10725_b1 , \5819_b1 , \5748_b1 );
not ( \5748_b1 , w_27208 );
and ( \10725_b0 , \5819_b0 , w_27209 );
and ( w_27208 , w_27209 , \5748_b0 );
or ( \10726_b1 , \10724_b1 , w_27211 );
not ( w_27211 , w_27212 );
and ( \10726_b0 , \10724_b0 , w_27213 );
and ( w_27212 ,  , w_27213 );
buf ( w_27211 , \10725_b1 );
not ( w_27211 , w_27214 );
not (  , w_27215 );
and ( w_27214 , w_27215 , \10725_b0 );
or ( \10727_b1 , \10726_b1 , w_27216 );
xor ( \10727_b0 , \10726_b0 , w_27218 );
not ( w_27218 , w_27219 );
and ( w_27219 , w_27216 , w_27217 );
buf ( w_27216 , \5755_b1 );
not ( w_27216 , w_27220 );
not ( w_27217 , w_27221 );
and ( w_27220 , w_27221 , \5755_b0 );
or ( \10728_b1 , \10723_b1 , \10727_b1 );
xor ( \10728_b0 , \10723_b0 , w_27222 );
not ( w_27222 , w_27223 );
and ( w_27223 , \10727_b1 , \10727_b0 );
or ( \10729_b1 , \10714_b1 , \10728_b1 );
xor ( \10729_b0 , \10714_b0 , w_27224 );
not ( w_27224 , w_27225 );
and ( w_27225 , \10728_b1 , \10728_b0 );
buf ( \10730_b1 , \7146_b1 );
not ( \10730_b1 , w_27226 );
not ( \10730_b0 , w_27227 );
and ( w_27226 , w_27227 , \7146_b0 );
or ( \10731_b1 , \5770_b1 , \7157_b1 );
not ( \7157_b1 , w_27228 );
and ( \10731_b0 , \5770_b0 , w_27229 );
and ( w_27228 , w_27229 , \7157_b0 );
or ( \10732_b1 , \5737_b1 , \7155_b1 );
not ( \7155_b1 , w_27230 );
and ( \10732_b0 , \5737_b0 , w_27231 );
and ( w_27230 , w_27231 , \7155_b0 );
or ( \10733_b1 , \10731_b1 , w_27233 );
not ( w_27233 , w_27234 );
and ( \10733_b0 , \10731_b0 , w_27235 );
and ( w_27234 ,  , w_27235 );
buf ( w_27233 , \10732_b1 );
not ( w_27233 , w_27236 );
not (  , w_27237 );
and ( w_27236 , w_27237 , \10732_b0 );
or ( \10734_b1 , \10733_b1 , w_27238 );
xor ( \10734_b0 , \10733_b0 , w_27240 );
not ( w_27240 , w_27241 );
and ( w_27241 , w_27238 , w_27239 );
buf ( w_27238 , \7163_b1 );
not ( w_27238 , w_27242 );
not ( w_27239 , w_27243 );
and ( w_27242 , w_27243 , \7163_b0 );
or ( \10735_b1 , \10730_b1 , \10734_b1 );
xor ( \10735_b0 , \10730_b0 , w_27244 );
not ( w_27244 , w_27245 );
and ( w_27245 , \10734_b1 , \10734_b0 );
or ( \10736_b1 , \5792_b1 , \7175_b1 );
not ( \7175_b1 , w_27246 );
and ( \10736_b0 , \5792_b0 , w_27247 );
and ( w_27246 , w_27247 , \7175_b0 );
or ( \10737_b1 , \5758_b1 , \7173_b1 );
not ( \7173_b1 , w_27248 );
and ( \10737_b0 , \5758_b0 , w_27249 );
and ( w_27248 , w_27249 , \7173_b0 );
or ( \10738_b1 , \10736_b1 , w_27251 );
not ( w_27251 , w_27252 );
and ( \10738_b0 , \10736_b0 , w_27253 );
and ( w_27252 ,  , w_27253 );
buf ( w_27251 , \10737_b1 );
not ( w_27251 , w_27254 );
not (  , w_27255 );
and ( w_27254 , w_27255 , \10737_b0 );
or ( \10739_b1 , \10738_b1 , w_27256 );
xor ( \10739_b0 , \10738_b0 , w_27258 );
not ( w_27258 , w_27259 );
and ( w_27259 , w_27256 , w_27257 );
buf ( w_27256 , \7181_b1 );
not ( w_27256 , w_27260 );
not ( w_27257 , w_27261 );
and ( w_27260 , w_27261 , \7181_b0 );
or ( \10740_b1 , \10735_b1 , \10739_b1 );
xor ( \10740_b0 , \10735_b0 , w_27262 );
not ( w_27262 , w_27263 );
and ( w_27263 , \10739_b1 , \10739_b0 );
or ( \10741_b1 , \10729_b1 , \10740_b1 );
xor ( \10741_b0 , \10729_b0 , w_27264 );
not ( w_27264 , w_27265 );
and ( w_27265 , \10740_b1 , \10740_b0 );
or ( \10742_b1 , \10700_b1 , \10741_b1 );
xor ( \10742_b0 , \10700_b0 , w_27266 );
not ( w_27266 , w_27267 );
and ( w_27267 , \10741_b1 , \10741_b0 );
or ( \10743_b1 , \6057_b1 , \5955_b1 );
not ( \5955_b1 , w_27268 );
and ( \10743_b0 , \6057_b0 , w_27269 );
and ( w_27268 , w_27269 , \5955_b0 );
or ( \10744_b1 , \6029_b1 , \5953_b1 );
not ( \5953_b1 , w_27270 );
and ( \10744_b0 , \6029_b0 , w_27271 );
and ( w_27270 , w_27271 , \5953_b0 );
or ( \10745_b1 , \10743_b1 , w_27273 );
not ( w_27273 , w_27274 );
and ( \10745_b0 , \10743_b0 , w_27275 );
and ( w_27274 ,  , w_27275 );
buf ( w_27273 , \10744_b1 );
not ( w_27273 , w_27276 );
not (  , w_27277 );
and ( w_27276 , w_27277 , \10744_b0 );
or ( \10746_b1 , \10745_b1 , w_27278 );
xor ( \10746_b0 , \10745_b0 , w_27280 );
not ( w_27280 , w_27281 );
and ( w_27281 , w_27278 , w_27279 );
buf ( w_27278 , \5962_b1 );
not ( w_27278 , w_27282 );
not ( w_27279 , w_27283 );
and ( w_27282 , w_27283 , \5962_b0 );
or ( \10747_b1 , \6065_b1 , \5977_b1 );
not ( \5977_b1 , w_27284 );
and ( \10747_b0 , \6065_b0 , w_27285 );
and ( w_27284 , w_27285 , \5977_b0 );
or ( \10748_b1 , \6048_b1 , \5975_b1 );
not ( \5975_b1 , w_27286 );
and ( \10748_b0 , \6048_b0 , w_27287 );
and ( w_27286 , w_27287 , \5975_b0 );
or ( \10749_b1 , \10747_b1 , w_27289 );
not ( w_27289 , w_27290 );
and ( \10749_b0 , \10747_b0 , w_27291 );
and ( w_27290 ,  , w_27291 );
buf ( w_27289 , \10748_b1 );
not ( w_27289 , w_27292 );
not (  , w_27293 );
and ( w_27292 , w_27293 , \10748_b0 );
or ( \10750_b1 , \10749_b1 , w_27294 );
xor ( \10750_b0 , \10749_b0 , w_27296 );
not ( w_27296 , w_27297 );
and ( w_27297 , w_27294 , w_27295 );
buf ( w_27294 , \5984_b1 );
not ( w_27294 , w_27298 );
not ( w_27295 , w_27299 );
and ( w_27298 , w_27299 , \5984_b0 );
or ( \10751_b1 , \10746_b1 , \10750_b1 );
xor ( \10751_b0 , \10746_b0 , w_27300 );
not ( w_27300 , w_27301 );
and ( w_27301 , \10750_b1 , \10750_b0 );
or ( \10752_b1 , \5998_b1 , \5891_b1 );
not ( \5891_b1 , w_27302 );
and ( \10752_b0 , \5998_b0 , w_27303 );
and ( w_27302 , w_27303 , \5891_b0 );
or ( \10753_b1 , \5967_b1 , \5889_b1 );
not ( \5889_b1 , w_27304 );
and ( \10753_b0 , \5967_b0 , w_27305 );
and ( w_27304 , w_27305 , \5889_b0 );
or ( \10754_b1 , \10752_b1 , w_27307 );
not ( w_27307 , w_27308 );
and ( \10754_b0 , \10752_b0 , w_27309 );
and ( w_27308 ,  , w_27309 );
buf ( w_27307 , \10753_b1 );
not ( w_27307 , w_27310 );
not (  , w_27311 );
and ( w_27310 , w_27311 , \10753_b0 );
or ( \10755_b1 , \10754_b1 , w_27312 );
xor ( \10755_b0 , \10754_b0 , w_27314 );
not ( w_27314 , w_27315 );
and ( w_27315 , w_27312 , w_27313 );
buf ( w_27312 , \5898_b1 );
not ( w_27312 , w_27316 );
not ( w_27313 , w_27317 );
and ( w_27316 , w_27317 , \5898_b0 );
or ( \10756_b1 , \6018_b1 , \5916_b1 );
not ( \5916_b1 , w_27318 );
and ( \10756_b0 , \6018_b0 , w_27319 );
and ( w_27318 , w_27319 , \5916_b0 );
or ( \10757_b1 , \5986_b1 , \5914_b1 );
not ( \5914_b1 , w_27320 );
and ( \10757_b0 , \5986_b0 , w_27321 );
and ( w_27320 , w_27321 , \5914_b0 );
or ( \10758_b1 , \10756_b1 , w_27323 );
not ( w_27323 , w_27324 );
and ( \10758_b0 , \10756_b0 , w_27325 );
and ( w_27324 ,  , w_27325 );
buf ( w_27323 , \10757_b1 );
not ( w_27323 , w_27326 );
not (  , w_27327 );
and ( w_27326 , w_27327 , \10757_b0 );
or ( \10759_b1 , \10758_b1 , w_27328 );
xor ( \10759_b0 , \10758_b0 , w_27330 );
not ( w_27330 , w_27331 );
and ( w_27331 , w_27328 , w_27329 );
buf ( w_27328 , \5923_b1 );
not ( w_27328 , w_27332 );
not ( w_27329 , w_27333 );
and ( w_27332 , w_27333 , \5923_b0 );
or ( \10760_b1 , \10755_b1 , \10759_b1 );
xor ( \10760_b0 , \10755_b0 , w_27334 );
not ( w_27334 , w_27335 );
and ( w_27335 , \10759_b1 , \10759_b0 );
or ( \10761_b1 , \6041_b1 , \5935_b1 );
not ( \5935_b1 , w_27336 );
and ( \10761_b0 , \6041_b0 , w_27337 );
and ( w_27336 , w_27337 , \5935_b0 );
or ( \10762_b1 , \6006_b1 , \5933_b1 );
not ( \5933_b1 , w_27338 );
and ( \10762_b0 , \6006_b0 , w_27339 );
and ( w_27338 , w_27339 , \5933_b0 );
or ( \10763_b1 , \10761_b1 , w_27341 );
not ( w_27341 , w_27342 );
and ( \10763_b0 , \10761_b0 , w_27343 );
and ( w_27342 ,  , w_27343 );
buf ( w_27341 , \10762_b1 );
not ( w_27341 , w_27344 );
not (  , w_27345 );
and ( w_27344 , w_27345 , \10762_b0 );
or ( \10764_b1 , \10763_b1 , w_27346 );
xor ( \10764_b0 , \10763_b0 , w_27348 );
not ( w_27348 , w_27349 );
and ( w_27349 , w_27346 , w_27347 );
buf ( w_27346 , \5942_b1 );
not ( w_27346 , w_27350 );
not ( w_27347 , w_27351 );
and ( w_27350 , w_27351 , \5942_b0 );
or ( \10765_b1 , \10760_b1 , \10764_b1 );
xor ( \10765_b0 , \10760_b0 , w_27352 );
not ( w_27352 , w_27353 );
and ( w_27353 , \10764_b1 , \10764_b0 );
or ( \10766_b1 , \10751_b1 , \10765_b1 );
xor ( \10766_b0 , \10751_b0 , w_27354 );
not ( w_27354 , w_27355 );
and ( w_27355 , \10765_b1 , \10765_b0 );
or ( \10767_b1 , \5937_b1 , \5829_b1 );
not ( \5829_b1 , w_27356 );
and ( \10767_b0 , \5937_b0 , w_27357 );
and ( w_27356 , w_27357 , \5829_b0 );
or ( \10768_b1 , \5906_b1 , \5827_b1 );
not ( \5827_b1 , w_27358 );
and ( \10768_b0 , \5906_b0 , w_27359 );
and ( w_27358 , w_27359 , \5827_b0 );
or ( \10769_b1 , \10767_b1 , w_27361 );
not ( w_27361 , w_27362 );
and ( \10769_b0 , \10767_b0 , w_27363 );
and ( w_27362 ,  , w_27363 );
buf ( w_27361 , \10768_b1 );
not ( w_27361 , w_27364 );
not (  , w_27365 );
and ( w_27364 , w_27365 , \10768_b0 );
or ( \10770_b1 , \10769_b1 , w_27366 );
xor ( \10770_b0 , \10769_b0 , w_27368 );
not ( w_27368 , w_27369 );
and ( w_27369 , w_27366 , w_27367 );
buf ( w_27366 , \5836_b1 );
not ( w_27366 , w_27370 );
not ( w_27367 , w_27371 );
and ( w_27370 , w_27371 , \5836_b0 );
or ( \10771_b1 , \5957_b1 , \5852_b1 );
not ( \5852_b1 , w_27372 );
and ( \10771_b0 , \5957_b0 , w_27373 );
and ( w_27372 , w_27373 , \5852_b0 );
or ( \10772_b1 , \5925_b1 , \5850_b1 );
not ( \5850_b1 , w_27374 );
and ( \10772_b0 , \5925_b0 , w_27375 );
and ( w_27374 , w_27375 , \5850_b0 );
or ( \10773_b1 , \10771_b1 , w_27377 );
not ( w_27377 , w_27378 );
and ( \10773_b0 , \10771_b0 , w_27379 );
and ( w_27378 ,  , w_27379 );
buf ( w_27377 , \10772_b1 );
not ( w_27377 , w_27380 );
not (  , w_27381 );
and ( w_27380 , w_27381 , \10772_b0 );
or ( \10774_b1 , \10773_b1 , w_27382 );
xor ( \10774_b0 , \10773_b0 , w_27384 );
not ( w_27384 , w_27385 );
and ( w_27385 , w_27382 , w_27383 );
buf ( w_27382 , \5859_b1 );
not ( w_27382 , w_27386 );
not ( w_27383 , w_27387 );
and ( w_27386 , w_27387 , \5859_b0 );
or ( \10775_b1 , \10770_b1 , \10774_b1 );
xor ( \10775_b0 , \10770_b0 , w_27388 );
not ( w_27388 , w_27389 );
and ( w_27389 , \10774_b1 , \10774_b0 );
or ( \10776_b1 , \5979_b1 , \5871_b1 );
not ( \5871_b1 , w_27390 );
and ( \10776_b0 , \5979_b0 , w_27391 );
and ( w_27390 , w_27391 , \5871_b0 );
or ( \10777_b1 , \5945_b1 , \5869_b1 );
not ( \5869_b1 , w_27392 );
and ( \10777_b0 , \5945_b0 , w_27393 );
and ( w_27392 , w_27393 , \5869_b0 );
or ( \10778_b1 , \10776_b1 , w_27395 );
not ( w_27395 , w_27396 );
and ( \10778_b0 , \10776_b0 , w_27397 );
and ( w_27396 ,  , w_27397 );
buf ( w_27395 , \10777_b1 );
not ( w_27395 , w_27398 );
not (  , w_27399 );
and ( w_27398 , w_27399 , \10777_b0 );
or ( \10779_b1 , \10778_b1 , w_27400 );
xor ( \10779_b0 , \10778_b0 , w_27402 );
not ( w_27402 , w_27403 );
and ( w_27403 , w_27400 , w_27401 );
buf ( w_27400 , \5878_b1 );
not ( w_27400 , w_27404 );
not ( w_27401 , w_27405 );
and ( w_27404 , w_27405 , \5878_b0 );
or ( \10780_b1 , \10775_b1 , \10779_b1 );
xor ( \10780_b0 , \10775_b0 , w_27406 );
not ( w_27406 , w_27407 );
and ( w_27407 , \10779_b1 , \10779_b0 );
or ( \10781_b1 , \10766_b1 , \10780_b1 );
xor ( \10781_b0 , \10766_b0 , w_27408 );
not ( w_27408 , w_27409 );
and ( w_27409 , \10780_b1 , \10780_b0 );
or ( \10782_b1 , \10742_b1 , \10781_b1 );
xor ( \10782_b0 , \10742_b0 , w_27410 );
not ( w_27410 , w_27411 );
and ( w_27411 , \10781_b1 , \10781_b0 );
or ( \10783_b1 , \10696_b1 , \10782_b1 );
xor ( \10783_b0 , \10696_b0 , w_27412 );
not ( w_27412 , w_27413 );
and ( w_27413 , \10782_b1 , \10782_b0 );
or ( \10784_b1 , \10545_b1 , \10549_b1 );
not ( \10549_b1 , w_27414 );
and ( \10784_b0 , \10545_b0 , w_27415 );
and ( w_27414 , w_27415 , \10549_b0 );
or ( \10785_b1 , \10549_b1 , \10554_b1 );
not ( \10554_b1 , w_27416 );
and ( \10785_b0 , \10549_b0 , w_27417 );
and ( w_27416 , w_27417 , \10554_b0 );
or ( \10786_b1 , \10545_b1 , \10554_b1 );
not ( \10554_b1 , w_27418 );
and ( \10786_b0 , \10545_b0 , w_27419 );
and ( w_27418 , w_27419 , \10554_b0 );
or ( \10788_b1 , \10533_b1 , \10537_b1 );
not ( \10537_b1 , w_27420 );
and ( \10788_b0 , \10533_b0 , w_27421 );
and ( w_27420 , w_27421 , \10537_b0 );
or ( \10789_b1 , \10537_b1 , \10539_b1 );
not ( \10539_b1 , w_27422 );
and ( \10789_b0 , \10537_b0 , w_27423 );
and ( w_27422 , w_27423 , \10539_b0 );
or ( \10790_b1 , \10533_b1 , \10539_b1 );
not ( \10539_b1 , w_27424 );
and ( \10790_b0 , \10533_b0 , w_27425 );
and ( w_27424 , w_27425 , \10539_b0 );
or ( \10792_b1 , \10787_b1 , \10791_b1 );
xor ( \10792_b0 , \10787_b0 , w_27426 );
not ( w_27426 , w_27427 );
and ( w_27427 , \10791_b1 , \10791_b0 );
or ( \10793_b1 , \10514_b1 , w_27428 );
or ( \10793_b0 , \10514_b0 , \10528_b0 );
not ( \10528_b0 , w_27429 );
and ( w_27429 , w_27428 , \10528_b1 );
or ( \10794_b1 , \10792_b1 , \10793_b1 );
xor ( \10794_b0 , \10792_b0 , w_27430 );
not ( w_27430 , w_27431 );
and ( w_27431 , \10793_b1 , \10793_b0 );
or ( \10795_b1 , \10783_b1 , \10794_b1 );
xor ( \10795_b0 , \10783_b0 , w_27432 );
not ( w_27432 , w_27433 );
and ( w_27433 , \10794_b1 , \10794_b0 );
or ( \10796_b1 , \10667_b1 , \10795_b1 );
xor ( \10796_b0 , \10667_b0 , w_27434 );
not ( w_27434 , w_27435 );
and ( w_27435 , \10795_b1 , \10795_b0 );
or ( \10797_b1 , \10658_b1 , \10796_b1 );
xor ( \10797_b0 , \10658_b0 , w_27436 );
not ( w_27436 , w_27437 );
and ( w_27437 , \10796_b1 , \10796_b0 );
or ( \10798_b1 , \10481_b1 , \10492_b1 );
not ( \10492_b1 , w_27438 );
and ( \10798_b0 , \10481_b0 , w_27439 );
and ( w_27438 , w_27439 , \10492_b0 );
or ( \10799_b1 , \10492_b1 , \10632_b1 );
not ( \10632_b1 , w_27440 );
and ( \10799_b0 , \10492_b0 , w_27441 );
and ( w_27440 , w_27441 , \10632_b0 );
or ( \10800_b1 , \10481_b1 , \10632_b1 );
not ( \10632_b1 , w_27442 );
and ( \10800_b0 , \10481_b0 , w_27443 );
and ( w_27442 , w_27443 , \10632_b0 );
or ( \10802_b1 , \10797_b1 , w_27445 );
not ( w_27445 , w_27446 );
and ( \10802_b0 , \10797_b0 , w_27447 );
and ( w_27446 ,  , w_27447 );
buf ( w_27445 , \10801_b1 );
not ( w_27445 , w_27448 );
not (  , w_27449 );
and ( w_27448 , w_27449 , \10801_b0 );
or ( \10803_b1 , \10662_b1 , \10666_b1 );
not ( \10666_b1 , w_27450 );
and ( \10803_b0 , \10662_b0 , w_27451 );
and ( w_27450 , w_27451 , \10666_b0 );
or ( \10804_b1 , \10666_b1 , \10795_b1 );
not ( \10795_b1 , w_27452 );
and ( \10804_b0 , \10666_b0 , w_27453 );
and ( w_27452 , w_27453 , \10795_b0 );
or ( \10805_b1 , \10662_b1 , \10795_b1 );
not ( \10795_b1 , w_27454 );
and ( \10805_b0 , \10662_b0 , w_27455 );
and ( w_27454 , w_27455 , \10795_b0 );
or ( \10807_b1 , \10787_b1 , \10791_b1 );
not ( \10791_b1 , w_27456 );
and ( \10807_b0 , \10787_b0 , w_27457 );
and ( w_27456 , w_27457 , \10791_b0 );
or ( \10808_b1 , \10791_b1 , \10793_b1 );
not ( \10793_b1 , w_27458 );
and ( \10808_b0 , \10791_b0 , w_27459 );
and ( w_27458 , w_27459 , \10793_b0 );
or ( \10809_b1 , \10787_b1 , \10793_b1 );
not ( \10793_b1 , w_27460 );
and ( \10809_b0 , \10787_b0 , w_27461 );
and ( w_27460 , w_27461 , \10793_b0 );
or ( \10811_b1 , \10700_b1 , \10741_b1 );
not ( \10741_b1 , w_27462 );
and ( \10811_b0 , \10700_b0 , w_27463 );
and ( w_27462 , w_27463 , \10741_b0 );
or ( \10812_b1 , \10741_b1 , \10781_b1 );
not ( \10781_b1 , w_27464 );
and ( \10812_b0 , \10741_b0 , w_27465 );
and ( w_27464 , w_27465 , \10781_b0 );
or ( \10813_b1 , \10700_b1 , \10781_b1 );
not ( \10781_b1 , w_27466 );
and ( \10813_b0 , \10700_b0 , w_27467 );
and ( w_27466 , w_27467 , \10781_b0 );
or ( \10815_b1 , \10810_b1 , \10814_b1 );
xor ( \10815_b0 , \10810_b0 , w_27468 );
not ( w_27468 , w_27469 );
and ( w_27469 , \10814_b1 , \10814_b0 );
or ( \10816_b1 , \10681_b1 , \10695_b1 );
not ( \10695_b1 , w_27470 );
and ( \10816_b0 , \10681_b0 , w_27471 );
and ( w_27470 , w_27471 , \10695_b0 );
or ( \10817_b1 , \10815_b1 , \10816_b1 );
xor ( \10817_b0 , \10815_b0 , w_27472 );
not ( w_27472 , w_27473 );
and ( w_27473 , \10816_b1 , \10816_b0 );
or ( \10818_b1 , \10806_b1 , \10817_b1 );
xor ( \10818_b0 , \10806_b0 , w_27474 );
not ( w_27474 , w_27475 );
and ( w_27475 , \10817_b1 , \10817_b0 );
or ( \10819_b1 , \10647_b1 , \10651_b1 );
not ( \10651_b1 , w_27476 );
and ( \10819_b0 , \10647_b0 , w_27477 );
and ( w_27476 , w_27477 , \10651_b0 );
or ( \10820_b1 , \10651_b1 , \10656_b1 );
not ( \10656_b1 , w_27478 );
and ( \10820_b0 , \10651_b0 , w_27479 );
and ( w_27478 , w_27479 , \10656_b0 );
or ( \10821_b1 , \10647_b1 , \10656_b1 );
not ( \10656_b1 , w_27480 );
and ( \10821_b0 , \10647_b0 , w_27481 );
and ( w_27480 , w_27481 , \10656_b0 );
or ( \10823_b1 , \10696_b1 , \10782_b1 );
not ( \10782_b1 , w_27482 );
and ( \10823_b0 , \10696_b0 , w_27483 );
and ( w_27482 , w_27483 , \10782_b0 );
or ( \10824_b1 , \10782_b1 , \10794_b1 );
not ( \10794_b1 , w_27484 );
and ( \10824_b0 , \10782_b0 , w_27485 );
and ( w_27484 , w_27485 , \10794_b0 );
or ( \10825_b1 , \10696_b1 , \10794_b1 );
not ( \10794_b1 , w_27486 );
and ( \10825_b0 , \10696_b0 , w_27487 );
and ( w_27486 , w_27487 , \10794_b0 );
or ( \10827_b1 , \10822_b1 , \10826_b1 );
xor ( \10827_b0 , \10822_b0 , w_27488 );
not ( w_27488 , w_27489 );
and ( w_27489 , \10826_b1 , \10826_b0 );
or ( \10828_b1 , \6029_b1 , \5955_b1 );
not ( \5955_b1 , w_27490 );
and ( \10828_b0 , \6029_b0 , w_27491 );
and ( w_27490 , w_27491 , \5955_b0 );
or ( \10829_b1 , \6041_b1 , \5953_b1 );
not ( \5953_b1 , w_27492 );
and ( \10829_b0 , \6041_b0 , w_27493 );
and ( w_27492 , w_27493 , \5953_b0 );
or ( \10830_b1 , \10828_b1 , w_27495 );
not ( w_27495 , w_27496 );
and ( \10830_b0 , \10828_b0 , w_27497 );
and ( w_27496 ,  , w_27497 );
buf ( w_27495 , \10829_b1 );
not ( w_27495 , w_27498 );
not (  , w_27499 );
and ( w_27498 , w_27499 , \10829_b0 );
or ( \10831_b1 , \10830_b1 , w_27500 );
xor ( \10831_b0 , \10830_b0 , w_27502 );
not ( w_27502 , w_27503 );
and ( w_27503 , w_27500 , w_27501 );
buf ( w_27500 , \5962_b1 );
not ( w_27500 , w_27504 );
not ( w_27501 , w_27505 );
and ( w_27504 , w_27505 , \5962_b0 );
or ( \10832_b1 , \6048_b1 , \5977_b1 );
not ( \5977_b1 , w_27506 );
and ( \10832_b0 , \6048_b0 , w_27507 );
and ( w_27506 , w_27507 , \5977_b0 );
or ( \10833_b1 , \6057_b1 , \5975_b1 );
not ( \5975_b1 , w_27508 );
and ( \10833_b0 , \6057_b0 , w_27509 );
and ( w_27508 , w_27509 , \5975_b0 );
or ( \10834_b1 , \10832_b1 , w_27511 );
not ( w_27511 , w_27512 );
and ( \10834_b0 , \10832_b0 , w_27513 );
and ( w_27512 ,  , w_27513 );
buf ( w_27511 , \10833_b1 );
not ( w_27511 , w_27514 );
not (  , w_27515 );
and ( w_27514 , w_27515 , \10833_b0 );
or ( \10835_b1 , \10834_b1 , w_27516 );
xor ( \10835_b0 , \10834_b0 , w_27518 );
not ( w_27518 , w_27519 );
and ( w_27519 , w_27516 , w_27517 );
buf ( w_27516 , \5984_b1 );
not ( w_27516 , w_27520 );
not ( w_27517 , w_27521 );
and ( w_27520 , w_27521 , \5984_b0 );
or ( \10836_b1 , \10831_b1 , \10835_b1 );
xor ( \10836_b0 , \10831_b0 , w_27522 );
not ( w_27522 , w_27523 );
and ( w_27523 , \10835_b1 , \10835_b0 );
or ( \10837_b1 , \6065_b1 , w_27525 );
not ( w_27525 , w_27526 );
and ( \10837_b0 , \6065_b0 , w_27527 );
and ( w_27526 ,  , w_27527 );
buf ( w_27525 , \5994_b1 );
not ( w_27525 , w_27528 );
not (  , w_27529 );
and ( w_27528 , w_27529 , \5994_b0 );
or ( \10838_b1 , \10837_b1 , w_27530 );
xor ( \10838_b0 , \10837_b0 , w_27532 );
not ( w_27532 , w_27533 );
and ( w_27533 , w_27530 , w_27531 );
buf ( w_27530 , \6003_b1 );
not ( w_27530 , w_27534 );
not ( w_27531 , w_27535 );
and ( w_27534 , w_27535 , \6003_b0 );
or ( \10839_b1 , \10836_b1 , \10838_b1 );
xor ( \10839_b0 , \10836_b0 , w_27536 );
not ( w_27536 , w_27537 );
and ( w_27537 , \10838_b1 , \10838_b0 );
or ( \10840_b1 , \5967_b1 , \5891_b1 );
not ( \5891_b1 , w_27538 );
and ( \10840_b0 , \5967_b0 , w_27539 );
and ( w_27538 , w_27539 , \5891_b0 );
or ( \10841_b1 , \5979_b1 , \5889_b1 );
not ( \5889_b1 , w_27540 );
and ( \10841_b0 , \5979_b0 , w_27541 );
and ( w_27540 , w_27541 , \5889_b0 );
or ( \10842_b1 , \10840_b1 , w_27543 );
not ( w_27543 , w_27544 );
and ( \10842_b0 , \10840_b0 , w_27545 );
and ( w_27544 ,  , w_27545 );
buf ( w_27543 , \10841_b1 );
not ( w_27543 , w_27546 );
not (  , w_27547 );
and ( w_27546 , w_27547 , \10841_b0 );
or ( \10843_b1 , \10842_b1 , w_27548 );
xor ( \10843_b0 , \10842_b0 , w_27550 );
not ( w_27550 , w_27551 );
and ( w_27551 , w_27548 , w_27549 );
buf ( w_27548 , \5898_b1 );
not ( w_27548 , w_27552 );
not ( w_27549 , w_27553 );
and ( w_27552 , w_27553 , \5898_b0 );
or ( \10844_b1 , \5986_b1 , \5916_b1 );
not ( \5916_b1 , w_27554 );
and ( \10844_b0 , \5986_b0 , w_27555 );
and ( w_27554 , w_27555 , \5916_b0 );
or ( \10845_b1 , \5998_b1 , \5914_b1 );
not ( \5914_b1 , w_27556 );
and ( \10845_b0 , \5998_b0 , w_27557 );
and ( w_27556 , w_27557 , \5914_b0 );
or ( \10846_b1 , \10844_b1 , w_27559 );
not ( w_27559 , w_27560 );
and ( \10846_b0 , \10844_b0 , w_27561 );
and ( w_27560 ,  , w_27561 );
buf ( w_27559 , \10845_b1 );
not ( w_27559 , w_27562 );
not (  , w_27563 );
and ( w_27562 , w_27563 , \10845_b0 );
or ( \10847_b1 , \10846_b1 , w_27564 );
xor ( \10847_b0 , \10846_b0 , w_27566 );
not ( w_27566 , w_27567 );
and ( w_27567 , w_27564 , w_27565 );
buf ( w_27564 , \5923_b1 );
not ( w_27564 , w_27568 );
not ( w_27565 , w_27569 );
and ( w_27568 , w_27569 , \5923_b0 );
or ( \10848_b1 , \10843_b1 , \10847_b1 );
xor ( \10848_b0 , \10843_b0 , w_27570 );
not ( w_27570 , w_27571 );
and ( w_27571 , \10847_b1 , \10847_b0 );
or ( \10849_b1 , \6006_b1 , \5935_b1 );
not ( \5935_b1 , w_27572 );
and ( \10849_b0 , \6006_b0 , w_27573 );
and ( w_27572 , w_27573 , \5935_b0 );
or ( \10850_b1 , \6018_b1 , \5933_b1 );
not ( \5933_b1 , w_27574 );
and ( \10850_b0 , \6018_b0 , w_27575 );
and ( w_27574 , w_27575 , \5933_b0 );
or ( \10851_b1 , \10849_b1 , w_27577 );
not ( w_27577 , w_27578 );
and ( \10851_b0 , \10849_b0 , w_27579 );
and ( w_27578 ,  , w_27579 );
buf ( w_27577 , \10850_b1 );
not ( w_27577 , w_27580 );
not (  , w_27581 );
and ( w_27580 , w_27581 , \10850_b0 );
or ( \10852_b1 , \10851_b1 , w_27582 );
xor ( \10852_b0 , \10851_b0 , w_27584 );
not ( w_27584 , w_27585 );
and ( w_27585 , w_27582 , w_27583 );
buf ( w_27582 , \5942_b1 );
not ( w_27582 , w_27586 );
not ( w_27583 , w_27587 );
and ( w_27586 , w_27587 , \5942_b0 );
or ( \10853_b1 , \10848_b1 , \10852_b1 );
xor ( \10853_b0 , \10848_b0 , w_27588 );
not ( w_27588 , w_27589 );
and ( w_27589 , \10852_b1 , \10852_b0 );
or ( \10854_b1 , \10839_b1 , w_27590 );
xor ( \10854_b0 , \10839_b0 , w_27592 );
not ( w_27592 , w_27593 );
and ( w_27593 , w_27590 , w_27591 );
buf ( w_27590 , \10853_b1 );
not ( w_27590 , w_27594 );
not ( w_27591 , w_27595 );
and ( w_27594 , w_27595 , \10853_b0 );
or ( \10855_b1 , \10770_b1 , \10774_b1 );
not ( \10774_b1 , w_27596 );
and ( \10855_b0 , \10770_b0 , w_27597 );
and ( w_27596 , w_27597 , \10774_b0 );
or ( \10856_b1 , \10774_b1 , \10779_b1 );
not ( \10779_b1 , w_27598 );
and ( \10856_b0 , \10774_b0 , w_27599 );
and ( w_27598 , w_27599 , \10779_b0 );
or ( \10857_b1 , \10770_b1 , \10779_b1 );
not ( \10779_b1 , w_27600 );
and ( \10857_b0 , \10770_b0 , w_27601 );
and ( w_27600 , w_27601 , \10779_b0 );
or ( \10859_b1 , \10755_b1 , \10759_b1 );
not ( \10759_b1 , w_27602 );
and ( \10859_b0 , \10755_b0 , w_27603 );
and ( w_27602 , w_27603 , \10759_b0 );
or ( \10860_b1 , \10759_b1 , \10764_b1 );
not ( \10764_b1 , w_27604 );
and ( \10860_b0 , \10759_b0 , w_27605 );
and ( w_27604 , w_27605 , \10764_b0 );
or ( \10861_b1 , \10755_b1 , \10764_b1 );
not ( \10764_b1 , w_27606 );
and ( \10861_b0 , \10755_b0 , w_27607 );
and ( w_27606 , w_27607 , \10764_b0 );
or ( \10863_b1 , \10858_b1 , \10862_b1 );
xor ( \10863_b0 , \10858_b0 , w_27608 );
not ( w_27608 , w_27609 );
and ( w_27609 , \10862_b1 , \10862_b0 );
or ( \10864_b1 , \10746_b1 , \10750_b1 );
not ( \10750_b1 , w_27610 );
and ( \10864_b0 , \10746_b0 , w_27611 );
and ( w_27610 , w_27611 , \10750_b0 );
or ( \10865_b1 , \10863_b1 , \10864_b1 );
xor ( \10865_b0 , \10863_b0 , w_27612 );
not ( w_27612 , w_27613 );
and ( w_27613 , \10864_b1 , \10864_b0 );
or ( \10866_b1 , \10854_b1 , \10865_b1 );
xor ( \10866_b0 , \10854_b0 , w_27614 );
not ( w_27614 , w_27615 );
and ( w_27615 , \10865_b1 , \10865_b0 );
or ( \10867_b1 , \10730_b1 , \10734_b1 );
not ( \10734_b1 , w_27616 );
and ( \10867_b0 , \10730_b0 , w_27617 );
and ( w_27616 , w_27617 , \10734_b0 );
or ( \10868_b1 , \10734_b1 , \10739_b1 );
not ( \10739_b1 , w_27618 );
and ( \10868_b0 , \10734_b0 , w_27619 );
and ( w_27618 , w_27619 , \10739_b0 );
or ( \10869_b1 , \10730_b1 , \10739_b1 );
not ( \10739_b1 , w_27620 );
and ( \10869_b0 , \10730_b0 , w_27621 );
and ( w_27620 , w_27621 , \10739_b0 );
or ( \10871_b1 , \10718_b1 , \10722_b1 );
not ( \10722_b1 , w_27622 );
and ( \10871_b0 , \10718_b0 , w_27623 );
and ( w_27622 , w_27623 , \10722_b0 );
or ( \10872_b1 , \10722_b1 , \10727_b1 );
not ( \10727_b1 , w_27624 );
and ( \10872_b0 , \10722_b0 , w_27625 );
and ( w_27624 , w_27625 , \10727_b0 );
or ( \10873_b1 , \10718_b1 , \10727_b1 );
not ( \10727_b1 , w_27626 );
and ( \10873_b0 , \10718_b0 , w_27627 );
and ( w_27626 , w_27627 , \10727_b0 );
or ( \10875_b1 , \10870_b1 , \10874_b1 );
xor ( \10875_b0 , \10870_b0 , w_27628 );
not ( w_27628 , w_27629 );
and ( w_27629 , \10874_b1 , \10874_b0 );
or ( \10876_b1 , \10704_b1 , \10708_b1 );
not ( \10708_b1 , w_27630 );
and ( \10876_b0 , \10704_b0 , w_27631 );
and ( w_27630 , w_27631 , \10708_b0 );
or ( \10877_b1 , \10708_b1 , \10713_b1 );
not ( \10713_b1 , w_27632 );
and ( \10877_b0 , \10708_b0 , w_27633 );
and ( w_27632 , w_27633 , \10713_b0 );
or ( \10878_b1 , \10704_b1 , \10713_b1 );
not ( \10713_b1 , w_27634 );
and ( \10878_b0 , \10704_b0 , w_27635 );
and ( w_27634 , w_27635 , \10713_b0 );
or ( \10880_b1 , \10875_b1 , \10879_b1 );
xor ( \10880_b0 , \10875_b0 , w_27636 );
not ( w_27636 , w_27637 );
and ( w_27637 , \10879_b1 , \10879_b0 );
or ( \10881_b1 , \10866_b1 , \10880_b1 );
xor ( \10881_b0 , \10866_b0 , w_27638 );
not ( w_27638 , w_27639 );
and ( w_27639 , \10880_b1 , \10880_b0 );
or ( \10882_b1 , \10714_b1 , \10728_b1 );
not ( \10728_b1 , w_27640 );
and ( \10882_b0 , \10714_b0 , w_27641 );
and ( w_27640 , w_27641 , \10728_b0 );
or ( \10883_b1 , \10728_b1 , \10740_b1 );
not ( \10740_b1 , w_27642 );
and ( \10883_b0 , \10728_b0 , w_27643 );
and ( w_27642 , w_27643 , \10740_b0 );
or ( \10884_b1 , \10714_b1 , \10740_b1 );
not ( \10740_b1 , w_27644 );
and ( \10884_b0 , \10714_b0 , w_27645 );
and ( w_27644 , w_27645 , \10740_b0 );
or ( \10886_b1 , \5737_b1 , \7157_b1 );
not ( \7157_b1 , w_27646 );
and ( \10886_b0 , \5737_b0 , w_27647 );
and ( w_27646 , w_27647 , \7157_b0 );
buf ( \10887_b1 , \10886_b1 );
not ( \10887_b1 , w_27648 );
not ( \10887_b0 , w_27649 );
and ( w_27648 , w_27649 , \10886_b0 );
or ( \10888_b1 , \10887_b1 , w_27650 );
xor ( \10888_b0 , \10887_b0 , w_27652 );
not ( w_27652 , w_27653 );
and ( w_27653 , w_27650 , w_27651 );
buf ( w_27650 , \7163_b1 );
not ( w_27650 , w_27654 );
not ( w_27651 , w_27655 );
and ( w_27654 , w_27655 , \7163_b0 );
or ( \10889_b1 , \6003_b1 , \10888_b1 );
xor ( \10889_b0 , \6003_b0 , w_27656 );
not ( w_27656 , w_27657 );
and ( w_27657 , \10888_b1 , \10888_b0 );
or ( \10890_b1 , \5758_b1 , \7175_b1 );
not ( \7175_b1 , w_27658 );
and ( \10890_b0 , \5758_b0 , w_27659 );
and ( w_27658 , w_27659 , \7175_b0 );
or ( \10891_b1 , \5770_b1 , \7173_b1 );
not ( \7173_b1 , w_27660 );
and ( \10891_b0 , \5770_b0 , w_27661 );
and ( w_27660 , w_27661 , \7173_b0 );
or ( \10892_b1 , \10890_b1 , w_27663 );
not ( w_27663 , w_27664 );
and ( \10892_b0 , \10890_b0 , w_27665 );
and ( w_27664 ,  , w_27665 );
buf ( w_27663 , \10891_b1 );
not ( w_27663 , w_27666 );
not (  , w_27667 );
and ( w_27666 , w_27667 , \10891_b0 );
or ( \10893_b1 , \10892_b1 , w_27668 );
xor ( \10893_b0 , \10892_b0 , w_27670 );
not ( w_27670 , w_27671 );
and ( w_27671 , w_27668 , w_27669 );
buf ( w_27668 , \7181_b1 );
not ( w_27668 , w_27672 );
not ( w_27669 , w_27673 );
and ( w_27672 , w_27673 , \7181_b0 );
or ( \10894_b1 , \10889_b1 , \10893_b1 );
xor ( \10894_b0 , \10889_b0 , w_27674 );
not ( w_27674 , w_27675 );
and ( w_27675 , \10893_b1 , \10893_b0 );
or ( \10895_b1 , \10885_b1 , \10894_b1 );
xor ( \10895_b0 , \10885_b0 , w_27676 );
not ( w_27676 , w_27677 );
and ( w_27677 , \10894_b1 , \10894_b0 );
or ( \10896_b1 , \5906_b1 , \5829_b1 );
not ( \5829_b1 , w_27678 );
and ( \10896_b0 , \5906_b0 , w_27679 );
and ( w_27678 , w_27679 , \5829_b0 );
or ( \10897_b1 , \5918_b1 , \5827_b1 );
not ( \5827_b1 , w_27680 );
and ( \10897_b0 , \5918_b0 , w_27681 );
and ( w_27680 , w_27681 , \5827_b0 );
or ( \10898_b1 , \10896_b1 , w_27683 );
not ( w_27683 , w_27684 );
and ( \10898_b0 , \10896_b0 , w_27685 );
and ( w_27684 ,  , w_27685 );
buf ( w_27683 , \10897_b1 );
not ( w_27683 , w_27686 );
not (  , w_27687 );
and ( w_27686 , w_27687 , \10897_b0 );
or ( \10899_b1 , \10898_b1 , w_27688 );
xor ( \10899_b0 , \10898_b0 , w_27690 );
not ( w_27690 , w_27691 );
and ( w_27691 , w_27688 , w_27689 );
buf ( w_27688 , \5836_b1 );
not ( w_27688 , w_27692 );
not ( w_27689 , w_27693 );
and ( w_27692 , w_27693 , \5836_b0 );
or ( \10900_b1 , \5925_b1 , \5852_b1 );
not ( \5852_b1 , w_27694 );
and ( \10900_b0 , \5925_b0 , w_27695 );
and ( w_27694 , w_27695 , \5852_b0 );
or ( \10901_b1 , \5937_b1 , \5850_b1 );
not ( \5850_b1 , w_27696 );
and ( \10901_b0 , \5937_b0 , w_27697 );
and ( w_27696 , w_27697 , \5850_b0 );
or ( \10902_b1 , \10900_b1 , w_27699 );
not ( w_27699 , w_27700 );
and ( \10902_b0 , \10900_b0 , w_27701 );
and ( w_27700 ,  , w_27701 );
buf ( w_27699 , \10901_b1 );
not ( w_27699 , w_27702 );
not (  , w_27703 );
and ( w_27702 , w_27703 , \10901_b0 );
or ( \10903_b1 , \10902_b1 , w_27704 );
xor ( \10903_b0 , \10902_b0 , w_27706 );
not ( w_27706 , w_27707 );
and ( w_27707 , w_27704 , w_27705 );
buf ( w_27704 , \5859_b1 );
not ( w_27704 , w_27708 );
not ( w_27705 , w_27709 );
and ( w_27708 , w_27709 , \5859_b0 );
or ( \10904_b1 , \10899_b1 , \10903_b1 );
xor ( \10904_b0 , \10899_b0 , w_27710 );
not ( w_27710 , w_27711 );
and ( w_27711 , \10903_b1 , \10903_b0 );
or ( \10905_b1 , \5945_b1 , \5871_b1 );
not ( \5871_b1 , w_27712 );
and ( \10905_b0 , \5945_b0 , w_27713 );
and ( w_27712 , w_27713 , \5871_b0 );
or ( \10906_b1 , \5957_b1 , \5869_b1 );
not ( \5869_b1 , w_27714 );
and ( \10906_b0 , \5957_b0 , w_27715 );
and ( w_27714 , w_27715 , \5869_b0 );
or ( \10907_b1 , \10905_b1 , w_27717 );
not ( w_27717 , w_27718 );
and ( \10907_b0 , \10905_b0 , w_27719 );
and ( w_27718 ,  , w_27719 );
buf ( w_27717 , \10906_b1 );
not ( w_27717 , w_27720 );
not (  , w_27721 );
and ( w_27720 , w_27721 , \10906_b0 );
or ( \10908_b1 , \10907_b1 , w_27722 );
xor ( \10908_b0 , \10907_b0 , w_27724 );
not ( w_27724 , w_27725 );
and ( w_27725 , w_27722 , w_27723 );
buf ( w_27722 , \5878_b1 );
not ( w_27722 , w_27726 );
not ( w_27723 , w_27727 );
and ( w_27726 , w_27727 , \5878_b0 );
or ( \10909_b1 , \10904_b1 , \10908_b1 );
xor ( \10909_b0 , \10904_b0 , w_27728 );
not ( w_27728 , w_27729 );
and ( w_27729 , \10908_b1 , \10908_b0 );
or ( \10910_b1 , \5842_b1 , \5768_b1 );
not ( \5768_b1 , w_27730 );
and ( \10910_b0 , \5842_b0 , w_27731 );
and ( w_27730 , w_27731 , \5768_b0 );
or ( \10911_b1 , \5854_b1 , \5766_b1 );
not ( \5766_b1 , w_27732 );
and ( \10911_b0 , \5854_b0 , w_27733 );
and ( w_27732 , w_27733 , \5766_b0 );
or ( \10912_b1 , \10910_b1 , w_27735 );
not ( w_27735 , w_27736 );
and ( \10912_b0 , \10910_b0 , w_27737 );
and ( w_27736 ,  , w_27737 );
buf ( w_27735 , \10911_b1 );
not ( w_27735 , w_27738 );
not (  , w_27739 );
and ( w_27738 , w_27739 , \10911_b0 );
or ( \10913_b1 , \10912_b1 , w_27740 );
xor ( \10913_b0 , \10912_b0 , w_27742 );
not ( w_27742 , w_27743 );
and ( w_27743 , w_27740 , w_27741 );
buf ( w_27740 , \5775_b1 );
not ( w_27740 , w_27744 );
not ( w_27741 , w_27745 );
and ( w_27744 , w_27745 , \5775_b0 );
or ( \10914_b1 , \5861_b1 , \5790_b1 );
not ( \5790_b1 , w_27746 );
and ( \10914_b0 , \5861_b0 , w_27747 );
and ( w_27746 , w_27747 , \5790_b0 );
or ( \10915_b1 , \5873_b1 , \5788_b1 );
not ( \5788_b1 , w_27748 );
and ( \10915_b0 , \5873_b0 , w_27749 );
and ( w_27748 , w_27749 , \5788_b0 );
or ( \10916_b1 , \10914_b1 , w_27751 );
not ( w_27751 , w_27752 );
and ( \10916_b0 , \10914_b0 , w_27753 );
and ( w_27752 ,  , w_27753 );
buf ( w_27751 , \10915_b1 );
not ( w_27751 , w_27754 );
not (  , w_27755 );
and ( w_27754 , w_27755 , \10915_b0 );
or ( \10917_b1 , \10916_b1 , w_27756 );
xor ( \10917_b0 , \10916_b0 , w_27758 );
not ( w_27758 , w_27759 );
and ( w_27759 , w_27756 , w_27757 );
buf ( w_27756 , \5797_b1 );
not ( w_27756 , w_27760 );
not ( w_27757 , w_27761 );
and ( w_27760 , w_27761 , \5797_b0 );
or ( \10918_b1 , \10913_b1 , \10917_b1 );
xor ( \10918_b0 , \10913_b0 , w_27762 );
not ( w_27762 , w_27763 );
and ( w_27763 , \10917_b1 , \10917_b0 );
or ( \10919_b1 , \5881_b1 , \5809_b1 );
not ( \5809_b1 , w_27764 );
and ( \10919_b0 , \5881_b0 , w_27765 );
and ( w_27764 , w_27765 , \5809_b0 );
or ( \10920_b1 , \5893_b1 , \5807_b1 );
not ( \5807_b1 , w_27766 );
and ( \10920_b0 , \5893_b0 , w_27767 );
and ( w_27766 , w_27767 , \5807_b0 );
or ( \10921_b1 , \10919_b1 , w_27769 );
not ( w_27769 , w_27770 );
and ( \10921_b0 , \10919_b0 , w_27771 );
and ( w_27770 ,  , w_27771 );
buf ( w_27769 , \10920_b1 );
not ( w_27769 , w_27772 );
not (  , w_27773 );
and ( w_27772 , w_27773 , \10920_b0 );
or ( \10922_b1 , \10921_b1 , w_27774 );
xor ( \10922_b0 , \10921_b0 , w_27776 );
not ( w_27776 , w_27777 );
and ( w_27777 , w_27774 , w_27775 );
buf ( w_27774 , \5816_b1 );
not ( w_27774 , w_27778 );
not ( w_27775 , w_27779 );
and ( w_27778 , w_27779 , \5816_b0 );
or ( \10923_b1 , \10918_b1 , \10922_b1 );
xor ( \10923_b0 , \10918_b0 , w_27780 );
not ( w_27780 , w_27781 );
and ( w_27781 , \10922_b1 , \10922_b0 );
or ( \10924_b1 , \10909_b1 , \10923_b1 );
xor ( \10924_b0 , \10909_b0 , w_27782 );
not ( w_27782 , w_27783 );
and ( w_27783 , \10923_b1 , \10923_b0 );
or ( \10925_b1 , \5780_b1 , \7192_b1 );
not ( \7192_b1 , w_27784 );
and ( \10925_b0 , \5780_b0 , w_27785 );
and ( w_27784 , w_27785 , \7192_b0 );
or ( \10926_b1 , \5792_b1 , \7190_b1 );
not ( \7190_b1 , w_27786 );
and ( \10926_b0 , \5792_b0 , w_27787 );
and ( w_27786 , w_27787 , \7190_b0 );
or ( \10927_b1 , \10925_b1 , w_27789 );
not ( w_27789 , w_27790 );
and ( \10927_b0 , \10925_b0 , w_27791 );
and ( w_27790 ,  , w_27791 );
buf ( w_27789 , \10926_b1 );
not ( w_27789 , w_27792 );
not (  , w_27793 );
and ( w_27792 , w_27793 , \10926_b0 );
or ( \10928_b1 , \10927_b1 , w_27794 );
xor ( \10928_b0 , \10927_b0 , w_27796 );
not ( w_27796 , w_27797 );
and ( w_27797 , w_27794 , w_27795 );
buf ( w_27794 , \7198_b1 );
not ( w_27794 , w_27798 );
not ( w_27795 , w_27799 );
and ( w_27798 , w_27799 , \7198_b0 );
or ( \10929_b1 , \5799_b1 , \7203_b1 );
not ( \7203_b1 , w_27800 );
and ( \10929_b0 , \5799_b0 , w_27801 );
and ( w_27800 , w_27801 , \7203_b0 );
or ( \10930_b1 , \5811_b1 , \7201_b1 );
not ( \7201_b1 , w_27802 );
and ( \10930_b0 , \5811_b0 , w_27803 );
and ( w_27802 , w_27803 , \7201_b0 );
or ( \10931_b1 , \10929_b1 , w_27805 );
not ( w_27805 , w_27806 );
and ( \10931_b0 , \10929_b0 , w_27807 );
and ( w_27806 ,  , w_27807 );
buf ( w_27805 , \10930_b1 );
not ( w_27805 , w_27808 );
not (  , w_27809 );
and ( w_27808 , w_27809 , \10930_b0 );
or ( \10932_b1 , \10931_b1 , w_27810 );
xor ( \10932_b0 , \10931_b0 , w_27812 );
not ( w_27812 , w_27813 );
and ( w_27813 , w_27810 , w_27811 );
buf ( w_27810 , \6824_b1 );
not ( w_27810 , w_27814 );
not ( w_27811 , w_27815 );
and ( w_27814 , w_27815 , \6824_b0 );
or ( \10933_b1 , \10928_b1 , \10932_b1 );
xor ( \10933_b0 , \10928_b0 , w_27816 );
not ( w_27816 , w_27817 );
and ( w_27817 , \10932_b1 , \10932_b0 );
or ( \10934_b1 , \5819_b1 , \5750_b1 );
not ( \5750_b1 , w_27818 );
and ( \10934_b0 , \5819_b0 , w_27819 );
and ( w_27818 , w_27819 , \5750_b0 );
or ( \10935_b1 , \5831_b1 , \5748_b1 );
not ( \5748_b1 , w_27820 );
and ( \10935_b0 , \5831_b0 , w_27821 );
and ( w_27820 , w_27821 , \5748_b0 );
or ( \10936_b1 , \10934_b1 , w_27823 );
not ( w_27823 , w_27824 );
and ( \10936_b0 , \10934_b0 , w_27825 );
and ( w_27824 ,  , w_27825 );
buf ( w_27823 , \10935_b1 );
not ( w_27823 , w_27826 );
not (  , w_27827 );
and ( w_27826 , w_27827 , \10935_b0 );
or ( \10937_b1 , \10936_b1 , w_27828 );
xor ( \10937_b0 , \10936_b0 , w_27830 );
not ( w_27830 , w_27831 );
and ( w_27831 , w_27828 , w_27829 );
buf ( w_27828 , \5755_b1 );
not ( w_27828 , w_27832 );
not ( w_27829 , w_27833 );
and ( w_27832 , w_27833 , \5755_b0 );
or ( \10938_b1 , \10933_b1 , \10937_b1 );
xor ( \10938_b0 , \10933_b0 , w_27834 );
not ( w_27834 , w_27835 );
and ( w_27835 , \10937_b1 , \10937_b0 );
or ( \10939_b1 , \10924_b1 , \10938_b1 );
xor ( \10939_b0 , \10924_b0 , w_27836 );
not ( w_27836 , w_27837 );
and ( w_27837 , \10938_b1 , \10938_b0 );
or ( \10940_b1 , \10895_b1 , \10939_b1 );
xor ( \10940_b0 , \10895_b0 , w_27838 );
not ( w_27838 , w_27839 );
and ( w_27839 , \10939_b1 , \10939_b0 );
or ( \10941_b1 , \10881_b1 , \10940_b1 );
xor ( \10941_b0 , \10881_b0 , w_27840 );
not ( w_27840 , w_27841 );
and ( w_27841 , \10940_b1 , \10940_b0 );
or ( \10942_b1 , \10685_b1 , \10689_b1 );
not ( \10689_b1 , w_27842 );
and ( \10942_b0 , \10685_b0 , w_27843 );
and ( w_27842 , w_27843 , \10689_b0 );
or ( \10943_b1 , \10689_b1 , \10694_b1 );
not ( \10694_b1 , w_27844 );
and ( \10943_b0 , \10689_b0 , w_27845 );
and ( w_27844 , w_27845 , \10694_b0 );
or ( \10944_b1 , \10685_b1 , \10694_b1 );
not ( \10694_b1 , w_27846 );
and ( \10944_b0 , \10685_b0 , w_27847 );
and ( w_27846 , w_27847 , \10694_b0 );
or ( \10946_b1 , \10671_b1 , \10675_b1 );
not ( \10675_b1 , w_27848 );
and ( \10946_b0 , \10671_b0 , w_27849 );
and ( w_27848 , w_27849 , \10675_b0 );
or ( \10947_b1 , \10675_b1 , \10680_b1 );
not ( \10680_b1 , w_27850 );
and ( \10947_b0 , \10675_b0 , w_27851 );
and ( w_27850 , w_27851 , \10680_b0 );
or ( \10948_b1 , \10671_b1 , \10680_b1 );
not ( \10680_b1 , w_27852 );
and ( \10948_b0 , \10671_b0 , w_27853 );
and ( w_27852 , w_27853 , \10680_b0 );
or ( \10950_b1 , \10945_b1 , \10949_b1 );
xor ( \10950_b0 , \10945_b0 , w_27854 );
not ( w_27854 , w_27855 );
and ( w_27855 , \10949_b1 , \10949_b0 );
or ( \10951_b1 , \10751_b1 , \10765_b1 );
not ( \10765_b1 , w_27856 );
and ( \10951_b0 , \10751_b0 , w_27857 );
and ( w_27856 , w_27857 , \10765_b0 );
or ( \10952_b1 , \10765_b1 , \10780_b1 );
not ( \10780_b1 , w_27858 );
and ( \10952_b0 , \10765_b0 , w_27859 );
and ( w_27858 , w_27859 , \10780_b0 );
or ( \10953_b1 , \10751_b1 , \10780_b1 );
not ( \10780_b1 , w_27860 );
and ( \10953_b0 , \10751_b0 , w_27861 );
and ( w_27860 , w_27861 , \10780_b0 );
or ( \10955_b1 , \10950_b1 , \10954_b1 );
xor ( \10955_b0 , \10950_b0 , w_27862 );
not ( w_27862 , w_27863 );
and ( w_27863 , \10954_b1 , \10954_b0 );
or ( \10956_b1 , \10941_b1 , \10955_b1 );
xor ( \10956_b0 , \10941_b0 , w_27864 );
not ( w_27864 , w_27865 );
and ( w_27865 , \10955_b1 , \10955_b0 );
or ( \10957_b1 , \10827_b1 , \10956_b1 );
xor ( \10957_b0 , \10827_b0 , w_27866 );
not ( w_27866 , w_27867 );
and ( w_27867 , \10956_b1 , \10956_b0 );
or ( \10958_b1 , \10818_b1 , \10957_b1 );
xor ( \10958_b0 , \10818_b0 , w_27868 );
not ( w_27868 , w_27869 );
and ( w_27869 , \10957_b1 , \10957_b0 );
or ( \10959_b1 , \10643_b1 , \10657_b1 );
not ( \10657_b1 , w_27870 );
and ( \10959_b0 , \10643_b0 , w_27871 );
and ( w_27870 , w_27871 , \10657_b0 );
or ( \10960_b1 , \10657_b1 , \10796_b1 );
not ( \10796_b1 , w_27872 );
and ( \10960_b0 , \10657_b0 , w_27873 );
and ( w_27872 , w_27873 , \10796_b0 );
or ( \10961_b1 , \10643_b1 , \10796_b1 );
not ( \10796_b1 , w_27874 );
and ( \10961_b0 , \10643_b0 , w_27875 );
and ( w_27874 , w_27875 , \10796_b0 );
or ( \10963_b1 , \10958_b1 , w_27877 );
not ( w_27877 , w_27878 );
and ( \10963_b0 , \10958_b0 , w_27879 );
and ( w_27878 ,  , w_27879 );
buf ( w_27877 , \10962_b1 );
not ( w_27877 , w_27880 );
not (  , w_27881 );
and ( w_27880 , w_27881 , \10962_b0 );
or ( \10964_b1 , \10802_b1 , w_27883 );
not ( w_27883 , w_27884 );
and ( \10964_b0 , \10802_b0 , w_27885 );
and ( w_27884 ,  , w_27885 );
buf ( w_27883 , \10963_b1 );
not ( w_27883 , w_27886 );
not (  , w_27887 );
and ( w_27886 , w_27887 , \10963_b0 );
or ( \10965_b1 , \10639_b1 , w_27889 );
not ( w_27889 , w_27890 );
and ( \10965_b0 , \10639_b0 , w_27891 );
and ( w_27890 ,  , w_27891 );
buf ( w_27889 , \10964_b1 );
not ( w_27889 , w_27892 );
not (  , w_27893 );
and ( w_27892 , w_27893 , \10964_b0 );
or ( \10966_b1 , \10822_b1 , \10826_b1 );
not ( \10826_b1 , w_27894 );
and ( \10966_b0 , \10822_b0 , w_27895 );
and ( w_27894 , w_27895 , \10826_b0 );
or ( \10967_b1 , \10826_b1 , \10956_b1 );
not ( \10956_b1 , w_27896 );
and ( \10967_b0 , \10826_b0 , w_27897 );
and ( w_27896 , w_27897 , \10956_b0 );
or ( \10968_b1 , \10822_b1 , \10956_b1 );
not ( \10956_b1 , w_27898 );
and ( \10968_b0 , \10822_b0 , w_27899 );
and ( w_27898 , w_27899 , \10956_b0 );
or ( \10970_b1 , \10945_b1 , \10949_b1 );
not ( \10949_b1 , w_27900 );
and ( \10970_b0 , \10945_b0 , w_27901 );
and ( w_27900 , w_27901 , \10949_b0 );
or ( \10971_b1 , \10949_b1 , \10954_b1 );
not ( \10954_b1 , w_27902 );
and ( \10971_b0 , \10949_b0 , w_27903 );
and ( w_27902 , w_27903 , \10954_b0 );
or ( \10972_b1 , \10945_b1 , \10954_b1 );
not ( \10954_b1 , w_27904 );
and ( \10972_b0 , \10945_b0 , w_27905 );
and ( w_27904 , w_27905 , \10954_b0 );
or ( \10974_b1 , \10885_b1 , \10894_b1 );
not ( \10894_b1 , w_27906 );
and ( \10974_b0 , \10885_b0 , w_27907 );
and ( w_27906 , w_27907 , \10894_b0 );
or ( \10975_b1 , \10894_b1 , \10939_b1 );
not ( \10939_b1 , w_27908 );
and ( \10975_b0 , \10894_b0 , w_27909 );
and ( w_27908 , w_27909 , \10939_b0 );
or ( \10976_b1 , \10885_b1 , \10939_b1 );
not ( \10939_b1 , w_27910 );
and ( \10976_b0 , \10885_b0 , w_27911 );
and ( w_27910 , w_27911 , \10939_b0 );
or ( \10978_b1 , \10973_b1 , \10977_b1 );
xor ( \10978_b0 , \10973_b0 , w_27912 );
not ( w_27912 , w_27913 );
and ( w_27913 , \10977_b1 , \10977_b0 );
or ( \10979_b1 , \10854_b1 , \10865_b1 );
not ( \10865_b1 , w_27914 );
and ( \10979_b0 , \10854_b0 , w_27915 );
and ( w_27914 , w_27915 , \10865_b0 );
or ( \10980_b1 , \10865_b1 , \10880_b1 );
not ( \10880_b1 , w_27916 );
and ( \10980_b0 , \10865_b0 , w_27917 );
and ( w_27916 , w_27917 , \10880_b0 );
or ( \10981_b1 , \10854_b1 , \10880_b1 );
not ( \10880_b1 , w_27918 );
and ( \10981_b0 , \10854_b0 , w_27919 );
and ( w_27918 , w_27919 , \10880_b0 );
or ( \10983_b1 , \10978_b1 , \10982_b1 );
xor ( \10983_b0 , \10978_b0 , w_27920 );
not ( w_27920 , w_27921 );
and ( w_27921 , \10982_b1 , \10982_b0 );
or ( \10984_b1 , \10969_b1 , \10983_b1 );
xor ( \10984_b0 , \10969_b0 , w_27922 );
not ( w_27922 , w_27923 );
and ( w_27923 , \10983_b1 , \10983_b0 );
or ( \10985_b1 , \10810_b1 , \10814_b1 );
not ( \10814_b1 , w_27924 );
and ( \10985_b0 , \10810_b0 , w_27925 );
and ( w_27924 , w_27925 , \10814_b0 );
or ( \10986_b1 , \10814_b1 , \10816_b1 );
not ( \10816_b1 , w_27926 );
and ( \10986_b0 , \10814_b0 , w_27927 );
and ( w_27926 , w_27927 , \10816_b0 );
or ( \10987_b1 , \10810_b1 , \10816_b1 );
not ( \10816_b1 , w_27928 );
and ( \10987_b0 , \10810_b0 , w_27929 );
and ( w_27928 , w_27929 , \10816_b0 );
or ( \10989_b1 , \10881_b1 , \10940_b1 );
not ( \10940_b1 , w_27930 );
and ( \10989_b0 , \10881_b0 , w_27931 );
and ( w_27930 , w_27931 , \10940_b0 );
or ( \10990_b1 , \10940_b1 , \10955_b1 );
not ( \10955_b1 , w_27932 );
and ( \10990_b0 , \10940_b0 , w_27933 );
and ( w_27932 , w_27933 , \10955_b0 );
or ( \10991_b1 , \10881_b1 , \10955_b1 );
not ( \10955_b1 , w_27934 );
and ( \10991_b0 , \10881_b0 , w_27935 );
and ( w_27934 , w_27935 , \10955_b0 );
or ( \10993_b1 , \10988_b1 , \10992_b1 );
xor ( \10993_b0 , \10988_b0 , w_27936 );
not ( w_27936 , w_27937 );
and ( w_27937 , \10992_b1 , \10992_b0 );
or ( \10994_b1 , \10899_b1 , \10903_b1 );
not ( \10903_b1 , w_27938 );
and ( \10994_b0 , \10899_b0 , w_27939 );
and ( w_27938 , w_27939 , \10903_b0 );
or ( \10995_b1 , \10903_b1 , \10908_b1 );
not ( \10908_b1 , w_27940 );
and ( \10995_b0 , \10903_b0 , w_27941 );
and ( w_27940 , w_27941 , \10908_b0 );
or ( \10996_b1 , \10899_b1 , \10908_b1 );
not ( \10908_b1 , w_27942 );
and ( \10996_b0 , \10899_b0 , w_27943 );
and ( w_27942 , w_27943 , \10908_b0 );
or ( \10998_b1 , \10843_b1 , \10847_b1 );
not ( \10847_b1 , w_27944 );
and ( \10998_b0 , \10843_b0 , w_27945 );
and ( w_27944 , w_27945 , \10847_b0 );
or ( \10999_b1 , \10847_b1 , \10852_b1 );
not ( \10852_b1 , w_27946 );
and ( \10999_b0 , \10847_b0 , w_27947 );
and ( w_27946 , w_27947 , \10852_b0 );
or ( \11000_b1 , \10843_b1 , \10852_b1 );
not ( \10852_b1 , w_27948 );
and ( \11000_b0 , \10843_b0 , w_27949 );
and ( w_27948 , w_27949 , \10852_b0 );
or ( \11002_b1 , \10997_b1 , \11001_b1 );
xor ( \11002_b0 , \10997_b0 , w_27950 );
not ( w_27950 , w_27951 );
and ( w_27951 , \11001_b1 , \11001_b0 );
or ( \11003_b1 , \10831_b1 , \10835_b1 );
not ( \10835_b1 , w_27952 );
and ( \11003_b0 , \10831_b0 , w_27953 );
and ( w_27952 , w_27953 , \10835_b0 );
or ( \11004_b1 , \10835_b1 , \10838_b1 );
not ( \10838_b1 , w_27954 );
and ( \11004_b0 , \10835_b0 , w_27955 );
and ( w_27954 , w_27955 , \10838_b0 );
or ( \11005_b1 , \10831_b1 , \10838_b1 );
not ( \10838_b1 , w_27956 );
and ( \11005_b0 , \10831_b0 , w_27957 );
and ( w_27956 , w_27957 , \10838_b0 );
or ( \11007_b1 , \11002_b1 , \11006_b1 );
xor ( \11007_b0 , \11002_b0 , w_27958 );
not ( w_27958 , w_27959 );
and ( w_27959 , \11006_b1 , \11006_b0 );
or ( \11008_b1 , \6003_b1 , \10888_b1 );
not ( \10888_b1 , w_27960 );
and ( \11008_b0 , \6003_b0 , w_27961 );
and ( w_27960 , w_27961 , \10888_b0 );
or ( \11009_b1 , \10888_b1 , \10893_b1 );
not ( \10893_b1 , w_27962 );
and ( \11009_b0 , \10888_b0 , w_27963 );
and ( w_27962 , w_27963 , \10893_b0 );
or ( \11010_b1 , \6003_b1 , \10893_b1 );
not ( \10893_b1 , w_27964 );
and ( \11010_b0 , \6003_b0 , w_27965 );
and ( w_27964 , w_27965 , \10893_b0 );
or ( \11012_b1 , \10928_b1 , \10932_b1 );
not ( \10932_b1 , w_27966 );
and ( \11012_b0 , \10928_b0 , w_27967 );
and ( w_27966 , w_27967 , \10932_b0 );
or ( \11013_b1 , \10932_b1 , \10937_b1 );
not ( \10937_b1 , w_27968 );
and ( \11013_b0 , \10932_b0 , w_27969 );
and ( w_27968 , w_27969 , \10937_b0 );
or ( \11014_b1 , \10928_b1 , \10937_b1 );
not ( \10937_b1 , w_27970 );
and ( \11014_b0 , \10928_b0 , w_27971 );
and ( w_27970 , w_27971 , \10937_b0 );
or ( \11016_b1 , \11011_b1 , \11015_b1 );
xor ( \11016_b0 , \11011_b0 , w_27972 );
not ( w_27972 , w_27973 );
and ( w_27973 , \11015_b1 , \11015_b0 );
or ( \11017_b1 , \10913_b1 , \10917_b1 );
not ( \10917_b1 , w_27974 );
and ( \11017_b0 , \10913_b0 , w_27975 );
and ( w_27974 , w_27975 , \10917_b0 );
or ( \11018_b1 , \10917_b1 , \10922_b1 );
not ( \10922_b1 , w_27976 );
and ( \11018_b0 , \10917_b0 , w_27977 );
and ( w_27976 , w_27977 , \10922_b0 );
or ( \11019_b1 , \10913_b1 , \10922_b1 );
not ( \10922_b1 , w_27978 );
and ( \11019_b0 , \10913_b0 , w_27979 );
and ( w_27978 , w_27979 , \10922_b0 );
or ( \11021_b1 , \11016_b1 , \11020_b1 );
xor ( \11021_b0 , \11016_b0 , w_27980 );
not ( w_27980 , w_27981 );
and ( w_27981 , \11020_b1 , \11020_b0 );
or ( \11022_b1 , \11007_b1 , \11021_b1 );
xor ( \11022_b0 , \11007_b0 , w_27982 );
not ( w_27982 , w_27983 );
and ( w_27983 , \11021_b1 , \11021_b0 );
or ( \11023_b1 , \10909_b1 , \10923_b1 );
not ( \10923_b1 , w_27984 );
and ( \11023_b0 , \10909_b0 , w_27985 );
and ( w_27984 , w_27985 , \10923_b0 );
or ( \11024_b1 , \10923_b1 , \10938_b1 );
not ( \10938_b1 , w_27986 );
and ( \11024_b0 , \10923_b0 , w_27987 );
and ( w_27986 , w_27987 , \10938_b0 );
or ( \11025_b1 , \10909_b1 , \10938_b1 );
not ( \10938_b1 , w_27988 );
and ( \11025_b0 , \10909_b0 , w_27989 );
and ( w_27988 , w_27989 , \10938_b0 );
or ( \11027_b1 , \5873_b1 , \5790_b1 );
not ( \5790_b1 , w_27990 );
and ( \11027_b0 , \5873_b0 , w_27991 );
and ( w_27990 , w_27991 , \5790_b0 );
or ( \11028_b1 , \5842_b1 , \5788_b1 );
not ( \5788_b1 , w_27992 );
and ( \11028_b0 , \5842_b0 , w_27993 );
and ( w_27992 , w_27993 , \5788_b0 );
or ( \11029_b1 , \11027_b1 , w_27995 );
not ( w_27995 , w_27996 );
and ( \11029_b0 , \11027_b0 , w_27997 );
and ( w_27996 ,  , w_27997 );
buf ( w_27995 , \11028_b1 );
not ( w_27995 , w_27998 );
not (  , w_27999 );
and ( w_27998 , w_27999 , \11028_b0 );
or ( \11030_b1 , \11029_b1 , w_28000 );
xor ( \11030_b0 , \11029_b0 , w_28002 );
not ( w_28002 , w_28003 );
and ( w_28003 , w_28000 , w_28001 );
buf ( w_28000 , \5797_b1 );
not ( w_28000 , w_28004 );
not ( w_28001 , w_28005 );
and ( w_28004 , w_28005 , \5797_b0 );
or ( \11031_b1 , \5893_b1 , \5809_b1 );
not ( \5809_b1 , w_28006 );
and ( \11031_b0 , \5893_b0 , w_28007 );
and ( w_28006 , w_28007 , \5809_b0 );
or ( \11032_b1 , \5861_b1 , \5807_b1 );
not ( \5807_b1 , w_28008 );
and ( \11032_b0 , \5861_b0 , w_28009 );
and ( w_28008 , w_28009 , \5807_b0 );
or ( \11033_b1 , \11031_b1 , w_28011 );
not ( w_28011 , w_28012 );
and ( \11033_b0 , \11031_b0 , w_28013 );
and ( w_28012 ,  , w_28013 );
buf ( w_28011 , \11032_b1 );
not ( w_28011 , w_28014 );
not (  , w_28015 );
and ( w_28014 , w_28015 , \11032_b0 );
or ( \11034_b1 , \11033_b1 , w_28016 );
xor ( \11034_b0 , \11033_b0 , w_28018 );
not ( w_28018 , w_28019 );
and ( w_28019 , w_28016 , w_28017 );
buf ( w_28016 , \5816_b1 );
not ( w_28016 , w_28020 );
not ( w_28017 , w_28021 );
and ( w_28020 , w_28021 , \5816_b0 );
or ( \11035_b1 , \11030_b1 , \11034_b1 );
xor ( \11035_b0 , \11030_b0 , w_28022 );
not ( w_28022 , w_28023 );
and ( w_28023 , \11034_b1 , \11034_b0 );
or ( \11036_b1 , \5918_b1 , \5829_b1 );
not ( \5829_b1 , w_28024 );
and ( \11036_b0 , \5918_b0 , w_28025 );
and ( w_28024 , w_28025 , \5829_b0 );
or ( \11037_b1 , \5881_b1 , \5827_b1 );
not ( \5827_b1 , w_28026 );
and ( \11037_b0 , \5881_b0 , w_28027 );
and ( w_28026 , w_28027 , \5827_b0 );
or ( \11038_b1 , \11036_b1 , w_28029 );
not ( w_28029 , w_28030 );
and ( \11038_b0 , \11036_b0 , w_28031 );
and ( w_28030 ,  , w_28031 );
buf ( w_28029 , \11037_b1 );
not ( w_28029 , w_28032 );
not (  , w_28033 );
and ( w_28032 , w_28033 , \11037_b0 );
or ( \11039_b1 , \11038_b1 , w_28034 );
xor ( \11039_b0 , \11038_b0 , w_28036 );
not ( w_28036 , w_28037 );
and ( w_28037 , w_28034 , w_28035 );
buf ( w_28034 , \5836_b1 );
not ( w_28034 , w_28038 );
not ( w_28035 , w_28039 );
and ( w_28038 , w_28039 , \5836_b0 );
or ( \11040_b1 , \11035_b1 , \11039_b1 );
xor ( \11040_b0 , \11035_b0 , w_28040 );
not ( w_28040 , w_28041 );
and ( w_28041 , \11039_b1 , \11039_b0 );
or ( \11041_b1 , \5811_b1 , \7203_b1 );
not ( \7203_b1 , w_28042 );
and ( \11041_b0 , \5811_b0 , w_28043 );
and ( w_28042 , w_28043 , \7203_b0 );
or ( \11042_b1 , \5780_b1 , \7201_b1 );
not ( \7201_b1 , w_28044 );
and ( \11042_b0 , \5780_b0 , w_28045 );
and ( w_28044 , w_28045 , \7201_b0 );
or ( \11043_b1 , \11041_b1 , w_28047 );
not ( w_28047 , w_28048 );
and ( \11043_b0 , \11041_b0 , w_28049 );
and ( w_28048 ,  , w_28049 );
buf ( w_28047 , \11042_b1 );
not ( w_28047 , w_28050 );
not (  , w_28051 );
and ( w_28050 , w_28051 , \11042_b0 );
or ( \11044_b1 , \11043_b1 , w_28052 );
xor ( \11044_b0 , \11043_b0 , w_28054 );
not ( w_28054 , w_28055 );
and ( w_28055 , w_28052 , w_28053 );
buf ( w_28052 , \6824_b1 );
not ( w_28052 , w_28056 );
not ( w_28053 , w_28057 );
and ( w_28056 , w_28057 , \6824_b0 );
or ( \11045_b1 , \5831_b1 , \5750_b1 );
not ( \5750_b1 , w_28058 );
and ( \11045_b0 , \5831_b0 , w_28059 );
and ( w_28058 , w_28059 , \5750_b0 );
or ( \11046_b1 , \5799_b1 , \5748_b1 );
not ( \5748_b1 , w_28060 );
and ( \11046_b0 , \5799_b0 , w_28061 );
and ( w_28060 , w_28061 , \5748_b0 );
or ( \11047_b1 , \11045_b1 , w_28063 );
not ( w_28063 , w_28064 );
and ( \11047_b0 , \11045_b0 , w_28065 );
and ( w_28064 ,  , w_28065 );
buf ( w_28063 , \11046_b1 );
not ( w_28063 , w_28066 );
not (  , w_28067 );
and ( w_28066 , w_28067 , \11046_b0 );
or ( \11048_b1 , \11047_b1 , w_28068 );
xor ( \11048_b0 , \11047_b0 , w_28070 );
not ( w_28070 , w_28071 );
and ( w_28071 , w_28068 , w_28069 );
buf ( w_28068 , \5755_b1 );
not ( w_28068 , w_28072 );
not ( w_28069 , w_28073 );
and ( w_28072 , w_28073 , \5755_b0 );
or ( \11049_b1 , \11044_b1 , \11048_b1 );
xor ( \11049_b0 , \11044_b0 , w_28074 );
not ( w_28074 , w_28075 );
and ( w_28075 , \11048_b1 , \11048_b0 );
or ( \11050_b1 , \5854_b1 , \5768_b1 );
not ( \5768_b1 , w_28076 );
and ( \11050_b0 , \5854_b0 , w_28077 );
and ( w_28076 , w_28077 , \5768_b0 );
or ( \11051_b1 , \5819_b1 , \5766_b1 );
not ( \5766_b1 , w_28078 );
and ( \11051_b0 , \5819_b0 , w_28079 );
and ( w_28078 , w_28079 , \5766_b0 );
or ( \11052_b1 , \11050_b1 , w_28081 );
not ( w_28081 , w_28082 );
and ( \11052_b0 , \11050_b0 , w_28083 );
and ( w_28082 ,  , w_28083 );
buf ( w_28081 , \11051_b1 );
not ( w_28081 , w_28084 );
not (  , w_28085 );
and ( w_28084 , w_28085 , \11051_b0 );
or ( \11053_b1 , \11052_b1 , w_28086 );
xor ( \11053_b0 , \11052_b0 , w_28088 );
not ( w_28088 , w_28089 );
and ( w_28089 , w_28086 , w_28087 );
buf ( w_28086 , \5775_b1 );
not ( w_28086 , w_28090 );
not ( w_28087 , w_28091 );
and ( w_28090 , w_28091 , \5775_b0 );
or ( \11054_b1 , \11049_b1 , \11053_b1 );
xor ( \11054_b0 , \11049_b0 , w_28092 );
not ( w_28092 , w_28093 );
and ( w_28093 , \11053_b1 , \11053_b0 );
or ( \11055_b1 , \11040_b1 , \11054_b1 );
xor ( \11055_b0 , \11040_b0 , w_28094 );
not ( w_28094 , w_28095 );
and ( w_28095 , \11054_b1 , \11054_b0 );
buf ( \11056_b1 , \7163_b1 );
not ( \11056_b1 , w_28096 );
not ( \11056_b0 , w_28097 );
and ( w_28096 , w_28097 , \7163_b0 );
or ( \11057_b1 , \5770_b1 , \7175_b1 );
not ( \7175_b1 , w_28098 );
and ( \11057_b0 , \5770_b0 , w_28099 );
and ( w_28098 , w_28099 , \7175_b0 );
or ( \11058_b1 , \5737_b1 , \7173_b1 );
not ( \7173_b1 , w_28100 );
and ( \11058_b0 , \5737_b0 , w_28101 );
and ( w_28100 , w_28101 , \7173_b0 );
or ( \11059_b1 , \11057_b1 , w_28103 );
not ( w_28103 , w_28104 );
and ( \11059_b0 , \11057_b0 , w_28105 );
and ( w_28104 ,  , w_28105 );
buf ( w_28103 , \11058_b1 );
not ( w_28103 , w_28106 );
not (  , w_28107 );
and ( w_28106 , w_28107 , \11058_b0 );
or ( \11060_b1 , \11059_b1 , w_28108 );
xor ( \11060_b0 , \11059_b0 , w_28110 );
not ( w_28110 , w_28111 );
and ( w_28111 , w_28108 , w_28109 );
buf ( w_28108 , \7181_b1 );
not ( w_28108 , w_28112 );
not ( w_28109 , w_28113 );
and ( w_28112 , w_28113 , \7181_b0 );
or ( \11061_b1 , \11056_b1 , \11060_b1 );
xor ( \11061_b0 , \11056_b0 , w_28114 );
not ( w_28114 , w_28115 );
and ( w_28115 , \11060_b1 , \11060_b0 );
or ( \11062_b1 , \5792_b1 , \7192_b1 );
not ( \7192_b1 , w_28116 );
and ( \11062_b0 , \5792_b0 , w_28117 );
and ( w_28116 , w_28117 , \7192_b0 );
or ( \11063_b1 , \5758_b1 , \7190_b1 );
not ( \7190_b1 , w_28118 );
and ( \11063_b0 , \5758_b0 , w_28119 );
and ( w_28118 , w_28119 , \7190_b0 );
or ( \11064_b1 , \11062_b1 , w_28121 );
not ( w_28121 , w_28122 );
and ( \11064_b0 , \11062_b0 , w_28123 );
and ( w_28122 ,  , w_28123 );
buf ( w_28121 , \11063_b1 );
not ( w_28121 , w_28124 );
not (  , w_28125 );
and ( w_28124 , w_28125 , \11063_b0 );
or ( \11065_b1 , \11064_b1 , w_28126 );
xor ( \11065_b0 , \11064_b0 , w_28128 );
not ( w_28128 , w_28129 );
and ( w_28129 , w_28126 , w_28127 );
buf ( w_28126 , \7198_b1 );
not ( w_28126 , w_28130 );
not ( w_28127 , w_28131 );
and ( w_28130 , w_28131 , \7198_b0 );
or ( \11066_b1 , \11061_b1 , \11065_b1 );
xor ( \11066_b0 , \11061_b0 , w_28132 );
not ( w_28132 , w_28133 );
and ( w_28133 , \11065_b1 , \11065_b0 );
or ( \11067_b1 , \11055_b1 , \11066_b1 );
xor ( \11067_b0 , \11055_b0 , w_28134 );
not ( w_28134 , w_28135 );
and ( w_28135 , \11066_b1 , \11066_b0 );
or ( \11068_b1 , \11026_b1 , \11067_b1 );
xor ( \11068_b0 , \11026_b0 , w_28136 );
not ( w_28136 , w_28137 );
and ( w_28137 , \11067_b1 , \11067_b0 );
or ( \11069_b1 , \6057_b1 , \5977_b1 );
not ( \5977_b1 , w_28138 );
and ( \11069_b0 , \6057_b0 , w_28139 );
and ( w_28138 , w_28139 , \5977_b0 );
or ( \11070_b1 , \6029_b1 , \5975_b1 );
not ( \5975_b1 , w_28140 );
and ( \11070_b0 , \6029_b0 , w_28141 );
and ( w_28140 , w_28141 , \5975_b0 );
or ( \11071_b1 , \11069_b1 , w_28143 );
not ( w_28143 , w_28144 );
and ( \11071_b0 , \11069_b0 , w_28145 );
and ( w_28144 ,  , w_28145 );
buf ( w_28143 , \11070_b1 );
not ( w_28143 , w_28146 );
not (  , w_28147 );
and ( w_28146 , w_28147 , \11070_b0 );
or ( \11072_b1 , \11071_b1 , w_28148 );
xor ( \11072_b0 , \11071_b0 , w_28150 );
not ( w_28150 , w_28151 );
and ( w_28151 , w_28148 , w_28149 );
buf ( w_28148 , \5984_b1 );
not ( w_28148 , w_28152 );
not ( w_28149 , w_28153 );
and ( w_28152 , w_28153 , \5984_b0 );
or ( \11073_b1 , \6065_b1 , \5996_b1 );
not ( \5996_b1 , w_28154 );
and ( \11073_b0 , \6065_b0 , w_28155 );
and ( w_28154 , w_28155 , \5996_b0 );
or ( \11074_b1 , \6048_b1 , \5994_b1 );
not ( \5994_b1 , w_28156 );
and ( \11074_b0 , \6048_b0 , w_28157 );
and ( w_28156 , w_28157 , \5994_b0 );
or ( \11075_b1 , \11073_b1 , w_28159 );
not ( w_28159 , w_28160 );
and ( \11075_b0 , \11073_b0 , w_28161 );
and ( w_28160 ,  , w_28161 );
buf ( w_28159 , \11074_b1 );
not ( w_28159 , w_28162 );
not (  , w_28163 );
and ( w_28162 , w_28163 , \11074_b0 );
or ( \11076_b1 , \11075_b1 , w_28164 );
xor ( \11076_b0 , \11075_b0 , w_28166 );
not ( w_28166 , w_28167 );
and ( w_28167 , w_28164 , w_28165 );
buf ( w_28164 , \6003_b1 );
not ( w_28164 , w_28168 );
not ( w_28165 , w_28169 );
and ( w_28168 , w_28169 , \6003_b0 );
or ( \11077_b1 , \11072_b1 , \11076_b1 );
xor ( \11077_b0 , \11072_b0 , w_28170 );
not ( w_28170 , w_28171 );
and ( w_28171 , \11076_b1 , \11076_b0 );
or ( \11078_b1 , \5998_b1 , \5916_b1 );
not ( \5916_b1 , w_28172 );
and ( \11078_b0 , \5998_b0 , w_28173 );
and ( w_28172 , w_28173 , \5916_b0 );
or ( \11079_b1 , \5967_b1 , \5914_b1 );
not ( \5914_b1 , w_28174 );
and ( \11079_b0 , \5967_b0 , w_28175 );
and ( w_28174 , w_28175 , \5914_b0 );
or ( \11080_b1 , \11078_b1 , w_28177 );
not ( w_28177 , w_28178 );
and ( \11080_b0 , \11078_b0 , w_28179 );
and ( w_28178 ,  , w_28179 );
buf ( w_28177 , \11079_b1 );
not ( w_28177 , w_28180 );
not (  , w_28181 );
and ( w_28180 , w_28181 , \11079_b0 );
or ( \11081_b1 , \11080_b1 , w_28182 );
xor ( \11081_b0 , \11080_b0 , w_28184 );
not ( w_28184 , w_28185 );
and ( w_28185 , w_28182 , w_28183 );
buf ( w_28182 , \5923_b1 );
not ( w_28182 , w_28186 );
not ( w_28183 , w_28187 );
and ( w_28186 , w_28187 , \5923_b0 );
or ( \11082_b1 , \6018_b1 , \5935_b1 );
not ( \5935_b1 , w_28188 );
and ( \11082_b0 , \6018_b0 , w_28189 );
and ( w_28188 , w_28189 , \5935_b0 );
or ( \11083_b1 , \5986_b1 , \5933_b1 );
not ( \5933_b1 , w_28190 );
and ( \11083_b0 , \5986_b0 , w_28191 );
and ( w_28190 , w_28191 , \5933_b0 );
or ( \11084_b1 , \11082_b1 , w_28193 );
not ( w_28193 , w_28194 );
and ( \11084_b0 , \11082_b0 , w_28195 );
and ( w_28194 ,  , w_28195 );
buf ( w_28193 , \11083_b1 );
not ( w_28193 , w_28196 );
not (  , w_28197 );
and ( w_28196 , w_28197 , \11083_b0 );
or ( \11085_b1 , \11084_b1 , w_28198 );
xor ( \11085_b0 , \11084_b0 , w_28200 );
not ( w_28200 , w_28201 );
and ( w_28201 , w_28198 , w_28199 );
buf ( w_28198 , \5942_b1 );
not ( w_28198 , w_28202 );
not ( w_28199 , w_28203 );
and ( w_28202 , w_28203 , \5942_b0 );
or ( \11086_b1 , \11081_b1 , \11085_b1 );
xor ( \11086_b0 , \11081_b0 , w_28204 );
not ( w_28204 , w_28205 );
and ( w_28205 , \11085_b1 , \11085_b0 );
or ( \11087_b1 , \6041_b1 , \5955_b1 );
not ( \5955_b1 , w_28206 );
and ( \11087_b0 , \6041_b0 , w_28207 );
and ( w_28206 , w_28207 , \5955_b0 );
or ( \11088_b1 , \6006_b1 , \5953_b1 );
not ( \5953_b1 , w_28208 );
and ( \11088_b0 , \6006_b0 , w_28209 );
and ( w_28208 , w_28209 , \5953_b0 );
or ( \11089_b1 , \11087_b1 , w_28211 );
not ( w_28211 , w_28212 );
and ( \11089_b0 , \11087_b0 , w_28213 );
and ( w_28212 ,  , w_28213 );
buf ( w_28211 , \11088_b1 );
not ( w_28211 , w_28214 );
not (  , w_28215 );
and ( w_28214 , w_28215 , \11088_b0 );
or ( \11090_b1 , \11089_b1 , w_28216 );
xor ( \11090_b0 , \11089_b0 , w_28218 );
not ( w_28218 , w_28219 );
and ( w_28219 , w_28216 , w_28217 );
buf ( w_28216 , \5962_b1 );
not ( w_28216 , w_28220 );
not ( w_28217 , w_28221 );
and ( w_28220 , w_28221 , \5962_b0 );
or ( \11091_b1 , \11086_b1 , \11090_b1 );
xor ( \11091_b0 , \11086_b0 , w_28222 );
not ( w_28222 , w_28223 );
and ( w_28223 , \11090_b1 , \11090_b0 );
or ( \11092_b1 , \11077_b1 , \11091_b1 );
xor ( \11092_b0 , \11077_b0 , w_28224 );
not ( w_28224 , w_28225 );
and ( w_28225 , \11091_b1 , \11091_b0 );
or ( \11093_b1 , \5937_b1 , \5852_b1 );
not ( \5852_b1 , w_28226 );
and ( \11093_b0 , \5937_b0 , w_28227 );
and ( w_28226 , w_28227 , \5852_b0 );
or ( \11094_b1 , \5906_b1 , \5850_b1 );
not ( \5850_b1 , w_28228 );
and ( \11094_b0 , \5906_b0 , w_28229 );
and ( w_28228 , w_28229 , \5850_b0 );
or ( \11095_b1 , \11093_b1 , w_28231 );
not ( w_28231 , w_28232 );
and ( \11095_b0 , \11093_b0 , w_28233 );
and ( w_28232 ,  , w_28233 );
buf ( w_28231 , \11094_b1 );
not ( w_28231 , w_28234 );
not (  , w_28235 );
and ( w_28234 , w_28235 , \11094_b0 );
or ( \11096_b1 , \11095_b1 , w_28236 );
xor ( \11096_b0 , \11095_b0 , w_28238 );
not ( w_28238 , w_28239 );
and ( w_28239 , w_28236 , w_28237 );
buf ( w_28236 , \5859_b1 );
not ( w_28236 , w_28240 );
not ( w_28237 , w_28241 );
and ( w_28240 , w_28241 , \5859_b0 );
or ( \11097_b1 , \5957_b1 , \5871_b1 );
not ( \5871_b1 , w_28242 );
and ( \11097_b0 , \5957_b0 , w_28243 );
and ( w_28242 , w_28243 , \5871_b0 );
or ( \11098_b1 , \5925_b1 , \5869_b1 );
not ( \5869_b1 , w_28244 );
and ( \11098_b0 , \5925_b0 , w_28245 );
and ( w_28244 , w_28245 , \5869_b0 );
or ( \11099_b1 , \11097_b1 , w_28247 );
not ( w_28247 , w_28248 );
and ( \11099_b0 , \11097_b0 , w_28249 );
and ( w_28248 ,  , w_28249 );
buf ( w_28247 , \11098_b1 );
not ( w_28247 , w_28250 );
not (  , w_28251 );
and ( w_28250 , w_28251 , \11098_b0 );
or ( \11100_b1 , \11099_b1 , w_28252 );
xor ( \11100_b0 , \11099_b0 , w_28254 );
not ( w_28254 , w_28255 );
and ( w_28255 , w_28252 , w_28253 );
buf ( w_28252 , \5878_b1 );
not ( w_28252 , w_28256 );
not ( w_28253 , w_28257 );
and ( w_28256 , w_28257 , \5878_b0 );
or ( \11101_b1 , \11096_b1 , \11100_b1 );
xor ( \11101_b0 , \11096_b0 , w_28258 );
not ( w_28258 , w_28259 );
and ( w_28259 , \11100_b1 , \11100_b0 );
or ( \11102_b1 , \5979_b1 , \5891_b1 );
not ( \5891_b1 , w_28260 );
and ( \11102_b0 , \5979_b0 , w_28261 );
and ( w_28260 , w_28261 , \5891_b0 );
or ( \11103_b1 , \5945_b1 , \5889_b1 );
not ( \5889_b1 , w_28262 );
and ( \11103_b0 , \5945_b0 , w_28263 );
and ( w_28262 , w_28263 , \5889_b0 );
or ( \11104_b1 , \11102_b1 , w_28265 );
not ( w_28265 , w_28266 );
and ( \11104_b0 , \11102_b0 , w_28267 );
and ( w_28266 ,  , w_28267 );
buf ( w_28265 , \11103_b1 );
not ( w_28265 , w_28268 );
not (  , w_28269 );
and ( w_28268 , w_28269 , \11103_b0 );
or ( \11105_b1 , \11104_b1 , w_28270 );
xor ( \11105_b0 , \11104_b0 , w_28272 );
not ( w_28272 , w_28273 );
and ( w_28273 , w_28270 , w_28271 );
buf ( w_28270 , \5898_b1 );
not ( w_28270 , w_28274 );
not ( w_28271 , w_28275 );
and ( w_28274 , w_28275 , \5898_b0 );
or ( \11106_b1 , \11101_b1 , \11105_b1 );
xor ( \11106_b0 , \11101_b0 , w_28276 );
not ( w_28276 , w_28277 );
and ( w_28277 , \11105_b1 , \11105_b0 );
or ( \11107_b1 , \11092_b1 , \11106_b1 );
xor ( \11107_b0 , \11092_b0 , w_28278 );
not ( w_28278 , w_28279 );
and ( w_28279 , \11106_b1 , \11106_b0 );
or ( \11108_b1 , \11068_b1 , \11107_b1 );
xor ( \11108_b0 , \11068_b0 , w_28280 );
not ( w_28280 , w_28281 );
and ( w_28281 , \11107_b1 , \11107_b0 );
or ( \11109_b1 , \11022_b1 , \11108_b1 );
xor ( \11109_b0 , \11022_b0 , w_28282 );
not ( w_28282 , w_28283 );
and ( w_28283 , \11108_b1 , \11108_b0 );
or ( \11110_b1 , \10870_b1 , \10874_b1 );
not ( \10874_b1 , w_28284 );
and ( \11110_b0 , \10870_b0 , w_28285 );
and ( w_28284 , w_28285 , \10874_b0 );
or ( \11111_b1 , \10874_b1 , \10879_b1 );
not ( \10879_b1 , w_28286 );
and ( \11111_b0 , \10874_b0 , w_28287 );
and ( w_28286 , w_28287 , \10879_b0 );
or ( \11112_b1 , \10870_b1 , \10879_b1 );
not ( \10879_b1 , w_28288 );
and ( \11112_b0 , \10870_b0 , w_28289 );
and ( w_28288 , w_28289 , \10879_b0 );
or ( \11114_b1 , \10858_b1 , \10862_b1 );
not ( \10862_b1 , w_28290 );
and ( \11114_b0 , \10858_b0 , w_28291 );
and ( w_28290 , w_28291 , \10862_b0 );
or ( \11115_b1 , \10862_b1 , \10864_b1 );
not ( \10864_b1 , w_28292 );
and ( \11115_b0 , \10862_b0 , w_28293 );
and ( w_28292 , w_28293 , \10864_b0 );
or ( \11116_b1 , \10858_b1 , \10864_b1 );
not ( \10864_b1 , w_28294 );
and ( \11116_b0 , \10858_b0 , w_28295 );
and ( w_28294 , w_28295 , \10864_b0 );
or ( \11118_b1 , \11113_b1 , \11117_b1 );
xor ( \11118_b0 , \11113_b0 , w_28296 );
not ( w_28296 , w_28297 );
and ( w_28297 , \11117_b1 , \11117_b0 );
or ( \11119_b1 , \10839_b1 , w_28298 );
or ( \11119_b0 , \10839_b0 , \10853_b0 );
not ( \10853_b0 , w_28299 );
and ( w_28299 , w_28298 , \10853_b1 );
or ( \11120_b1 , \11118_b1 , \11119_b1 );
xor ( \11120_b0 , \11118_b0 , w_28300 );
not ( w_28300 , w_28301 );
and ( w_28301 , \11119_b1 , \11119_b0 );
or ( \11121_b1 , \11109_b1 , \11120_b1 );
xor ( \11121_b0 , \11109_b0 , w_28302 );
not ( w_28302 , w_28303 );
and ( w_28303 , \11120_b1 , \11120_b0 );
or ( \11122_b1 , \10993_b1 , \11121_b1 );
xor ( \11122_b0 , \10993_b0 , w_28304 );
not ( w_28304 , w_28305 );
and ( w_28305 , \11121_b1 , \11121_b0 );
or ( \11123_b1 , \10984_b1 , \11122_b1 );
xor ( \11123_b0 , \10984_b0 , w_28306 );
not ( w_28306 , w_28307 );
and ( w_28307 , \11122_b1 , \11122_b0 );
or ( \11124_b1 , \10806_b1 , \10817_b1 );
not ( \10817_b1 , w_28308 );
and ( \11124_b0 , \10806_b0 , w_28309 );
and ( w_28308 , w_28309 , \10817_b0 );
or ( \11125_b1 , \10817_b1 , \10957_b1 );
not ( \10957_b1 , w_28310 );
and ( \11125_b0 , \10817_b0 , w_28311 );
and ( w_28310 , w_28311 , \10957_b0 );
or ( \11126_b1 , \10806_b1 , \10957_b1 );
not ( \10957_b1 , w_28312 );
and ( \11126_b0 , \10806_b0 , w_28313 );
and ( w_28312 , w_28313 , \10957_b0 );
or ( \11128_b1 , \11123_b1 , w_28315 );
not ( w_28315 , w_28316 );
and ( \11128_b0 , \11123_b0 , w_28317 );
and ( w_28316 ,  , w_28317 );
buf ( w_28315 , \11127_b1 );
not ( w_28315 , w_28318 );
not (  , w_28319 );
and ( w_28318 , w_28319 , \11127_b0 );
or ( \11129_b1 , \10988_b1 , \10992_b1 );
not ( \10992_b1 , w_28320 );
and ( \11129_b0 , \10988_b0 , w_28321 );
and ( w_28320 , w_28321 , \10992_b0 );
or ( \11130_b1 , \10992_b1 , \11121_b1 );
not ( \11121_b1 , w_28322 );
and ( \11130_b0 , \10992_b0 , w_28323 );
and ( w_28322 , w_28323 , \11121_b0 );
or ( \11131_b1 , \10988_b1 , \11121_b1 );
not ( \11121_b1 , w_28324 );
and ( \11131_b0 , \10988_b0 , w_28325 );
and ( w_28324 , w_28325 , \11121_b0 );
or ( \11133_b1 , \11113_b1 , \11117_b1 );
not ( \11117_b1 , w_28326 );
and ( \11133_b0 , \11113_b0 , w_28327 );
and ( w_28326 , w_28327 , \11117_b0 );
or ( \11134_b1 , \11117_b1 , \11119_b1 );
not ( \11119_b1 , w_28328 );
and ( \11134_b0 , \11117_b0 , w_28329 );
and ( w_28328 , w_28329 , \11119_b0 );
or ( \11135_b1 , \11113_b1 , \11119_b1 );
not ( \11119_b1 , w_28330 );
and ( \11135_b0 , \11113_b0 , w_28331 );
and ( w_28330 , w_28331 , \11119_b0 );
or ( \11137_b1 , \11026_b1 , \11067_b1 );
not ( \11067_b1 , w_28332 );
and ( \11137_b0 , \11026_b0 , w_28333 );
and ( w_28332 , w_28333 , \11067_b0 );
or ( \11138_b1 , \11067_b1 , \11107_b1 );
not ( \11107_b1 , w_28334 );
and ( \11138_b0 , \11067_b0 , w_28335 );
and ( w_28334 , w_28335 , \11107_b0 );
or ( \11139_b1 , \11026_b1 , \11107_b1 );
not ( \11107_b1 , w_28336 );
and ( \11139_b0 , \11026_b0 , w_28337 );
and ( w_28336 , w_28337 , \11107_b0 );
or ( \11141_b1 , \11136_b1 , \11140_b1 );
xor ( \11141_b0 , \11136_b0 , w_28338 );
not ( w_28338 , w_28339 );
and ( w_28339 , \11140_b1 , \11140_b0 );
or ( \11142_b1 , \11007_b1 , \11021_b1 );
not ( \11021_b1 , w_28340 );
and ( \11142_b0 , \11007_b0 , w_28341 );
and ( w_28340 , w_28341 , \11021_b0 );
or ( \11143_b1 , \11141_b1 , \11142_b1 );
xor ( \11143_b0 , \11141_b0 , w_28342 );
not ( w_28342 , w_28343 );
and ( w_28343 , \11142_b1 , \11142_b0 );
or ( \11144_b1 , \11132_b1 , \11143_b1 );
xor ( \11144_b0 , \11132_b0 , w_28344 );
not ( w_28344 , w_28345 );
and ( w_28345 , \11143_b1 , \11143_b0 );
or ( \11145_b1 , \10973_b1 , \10977_b1 );
not ( \10977_b1 , w_28346 );
and ( \11145_b0 , \10973_b0 , w_28347 );
and ( w_28346 , w_28347 , \10977_b0 );
or ( \11146_b1 , \10977_b1 , \10982_b1 );
not ( \10982_b1 , w_28348 );
and ( \11146_b0 , \10977_b0 , w_28349 );
and ( w_28348 , w_28349 , \10982_b0 );
or ( \11147_b1 , \10973_b1 , \10982_b1 );
not ( \10982_b1 , w_28350 );
and ( \11147_b0 , \10973_b0 , w_28351 );
and ( w_28350 , w_28351 , \10982_b0 );
or ( \11149_b1 , \11022_b1 , \11108_b1 );
not ( \11108_b1 , w_28352 );
and ( \11149_b0 , \11022_b0 , w_28353 );
and ( w_28352 , w_28353 , \11108_b0 );
or ( \11150_b1 , \11108_b1 , \11120_b1 );
not ( \11120_b1 , w_28354 );
and ( \11150_b0 , \11108_b0 , w_28355 );
and ( w_28354 , w_28355 , \11120_b0 );
or ( \11151_b1 , \11022_b1 , \11120_b1 );
not ( \11120_b1 , w_28356 );
and ( \11151_b0 , \11022_b0 , w_28357 );
and ( w_28356 , w_28357 , \11120_b0 );
or ( \11153_b1 , \11148_b1 , \11152_b1 );
xor ( \11153_b0 , \11148_b0 , w_28358 );
not ( w_28358 , w_28359 );
and ( w_28359 , \11152_b1 , \11152_b0 );
or ( \11154_b1 , \6029_b1 , \5977_b1 );
not ( \5977_b1 , w_28360 );
and ( \11154_b0 , \6029_b0 , w_28361 );
and ( w_28360 , w_28361 , \5977_b0 );
or ( \11155_b1 , \6041_b1 , \5975_b1 );
not ( \5975_b1 , w_28362 );
and ( \11155_b0 , \6041_b0 , w_28363 );
and ( w_28362 , w_28363 , \5975_b0 );
or ( \11156_b1 , \11154_b1 , w_28365 );
not ( w_28365 , w_28366 );
and ( \11156_b0 , \11154_b0 , w_28367 );
and ( w_28366 ,  , w_28367 );
buf ( w_28365 , \11155_b1 );
not ( w_28365 , w_28368 );
not (  , w_28369 );
and ( w_28368 , w_28369 , \11155_b0 );
or ( \11157_b1 , \11156_b1 , w_28370 );
xor ( \11157_b0 , \11156_b0 , w_28372 );
not ( w_28372 , w_28373 );
and ( w_28373 , w_28370 , w_28371 );
buf ( w_28370 , \5984_b1 );
not ( w_28370 , w_28374 );
not ( w_28371 , w_28375 );
and ( w_28374 , w_28375 , \5984_b0 );
or ( \11158_b1 , \6048_b1 , \5996_b1 );
not ( \5996_b1 , w_28376 );
and ( \11158_b0 , \6048_b0 , w_28377 );
and ( w_28376 , w_28377 , \5996_b0 );
or ( \11159_b1 , \6057_b1 , \5994_b1 );
not ( \5994_b1 , w_28378 );
and ( \11159_b0 , \6057_b0 , w_28379 );
and ( w_28378 , w_28379 , \5994_b0 );
or ( \11160_b1 , \11158_b1 , w_28381 );
not ( w_28381 , w_28382 );
and ( \11160_b0 , \11158_b0 , w_28383 );
and ( w_28382 ,  , w_28383 );
buf ( w_28381 , \11159_b1 );
not ( w_28381 , w_28384 );
not (  , w_28385 );
and ( w_28384 , w_28385 , \11159_b0 );
or ( \11161_b1 , \11160_b1 , w_28386 );
xor ( \11161_b0 , \11160_b0 , w_28388 );
not ( w_28388 , w_28389 );
and ( w_28389 , w_28386 , w_28387 );
buf ( w_28386 , \6003_b1 );
not ( w_28386 , w_28390 );
not ( w_28387 , w_28391 );
and ( w_28390 , w_28391 , \6003_b0 );
or ( \11162_b1 , \11157_b1 , \11161_b1 );
xor ( \11162_b0 , \11157_b0 , w_28392 );
not ( w_28392 , w_28393 );
and ( w_28393 , \11161_b1 , \11161_b0 );
or ( \11163_b1 , \6065_b1 , w_28395 );
not ( w_28395 , w_28396 );
and ( \11163_b0 , \6065_b0 , w_28397 );
and ( w_28396 ,  , w_28397 );
buf ( w_28395 , \6014_b1 );
not ( w_28395 , w_28398 );
not (  , w_28399 );
and ( w_28398 , w_28399 , \6014_b0 );
or ( \11164_b1 , \11163_b1 , w_28400 );
xor ( \11164_b0 , \11163_b0 , w_28402 );
not ( w_28402 , w_28403 );
and ( w_28403 , w_28400 , w_28401 );
buf ( w_28400 , \6023_b1 );
not ( w_28400 , w_28404 );
not ( w_28401 , w_28405 );
and ( w_28404 , w_28405 , \6023_b0 );
or ( \11165_b1 , \11162_b1 , \11164_b1 );
xor ( \11165_b0 , \11162_b0 , w_28406 );
not ( w_28406 , w_28407 );
and ( w_28407 , \11164_b1 , \11164_b0 );
or ( \11166_b1 , \5967_b1 , \5916_b1 );
not ( \5916_b1 , w_28408 );
and ( \11166_b0 , \5967_b0 , w_28409 );
and ( w_28408 , w_28409 , \5916_b0 );
or ( \11167_b1 , \5979_b1 , \5914_b1 );
not ( \5914_b1 , w_28410 );
and ( \11167_b0 , \5979_b0 , w_28411 );
and ( w_28410 , w_28411 , \5914_b0 );
or ( \11168_b1 , \11166_b1 , w_28413 );
not ( w_28413 , w_28414 );
and ( \11168_b0 , \11166_b0 , w_28415 );
and ( w_28414 ,  , w_28415 );
buf ( w_28413 , \11167_b1 );
not ( w_28413 , w_28416 );
not (  , w_28417 );
and ( w_28416 , w_28417 , \11167_b0 );
or ( \11169_b1 , \11168_b1 , w_28418 );
xor ( \11169_b0 , \11168_b0 , w_28420 );
not ( w_28420 , w_28421 );
and ( w_28421 , w_28418 , w_28419 );
buf ( w_28418 , \5923_b1 );
not ( w_28418 , w_28422 );
not ( w_28419 , w_28423 );
and ( w_28422 , w_28423 , \5923_b0 );
or ( \11170_b1 , \5986_b1 , \5935_b1 );
not ( \5935_b1 , w_28424 );
and ( \11170_b0 , \5986_b0 , w_28425 );
and ( w_28424 , w_28425 , \5935_b0 );
or ( \11171_b1 , \5998_b1 , \5933_b1 );
not ( \5933_b1 , w_28426 );
and ( \11171_b0 , \5998_b0 , w_28427 );
and ( w_28426 , w_28427 , \5933_b0 );
or ( \11172_b1 , \11170_b1 , w_28429 );
not ( w_28429 , w_28430 );
and ( \11172_b0 , \11170_b0 , w_28431 );
and ( w_28430 ,  , w_28431 );
buf ( w_28429 , \11171_b1 );
not ( w_28429 , w_28432 );
not (  , w_28433 );
and ( w_28432 , w_28433 , \11171_b0 );
or ( \11173_b1 , \11172_b1 , w_28434 );
xor ( \11173_b0 , \11172_b0 , w_28436 );
not ( w_28436 , w_28437 );
and ( w_28437 , w_28434 , w_28435 );
buf ( w_28434 , \5942_b1 );
not ( w_28434 , w_28438 );
not ( w_28435 , w_28439 );
and ( w_28438 , w_28439 , \5942_b0 );
or ( \11174_b1 , \11169_b1 , \11173_b1 );
xor ( \11174_b0 , \11169_b0 , w_28440 );
not ( w_28440 , w_28441 );
and ( w_28441 , \11173_b1 , \11173_b0 );
or ( \11175_b1 , \6006_b1 , \5955_b1 );
not ( \5955_b1 , w_28442 );
and ( \11175_b0 , \6006_b0 , w_28443 );
and ( w_28442 , w_28443 , \5955_b0 );
or ( \11176_b1 , \6018_b1 , \5953_b1 );
not ( \5953_b1 , w_28444 );
and ( \11176_b0 , \6018_b0 , w_28445 );
and ( w_28444 , w_28445 , \5953_b0 );
or ( \11177_b1 , \11175_b1 , w_28447 );
not ( w_28447 , w_28448 );
and ( \11177_b0 , \11175_b0 , w_28449 );
and ( w_28448 ,  , w_28449 );
buf ( w_28447 , \11176_b1 );
not ( w_28447 , w_28450 );
not (  , w_28451 );
and ( w_28450 , w_28451 , \11176_b0 );
or ( \11178_b1 , \11177_b1 , w_28452 );
xor ( \11178_b0 , \11177_b0 , w_28454 );
not ( w_28454 , w_28455 );
and ( w_28455 , w_28452 , w_28453 );
buf ( w_28452 , \5962_b1 );
not ( w_28452 , w_28456 );
not ( w_28453 , w_28457 );
and ( w_28456 , w_28457 , \5962_b0 );
or ( \11179_b1 , \11174_b1 , \11178_b1 );
xor ( \11179_b0 , \11174_b0 , w_28458 );
not ( w_28458 , w_28459 );
and ( w_28459 , \11178_b1 , \11178_b0 );
or ( \11180_b1 , \11165_b1 , w_28460 );
xor ( \11180_b0 , \11165_b0 , w_28462 );
not ( w_28462 , w_28463 );
and ( w_28463 , w_28460 , w_28461 );
buf ( w_28460 , \11179_b1 );
not ( w_28460 , w_28464 );
not ( w_28461 , w_28465 );
and ( w_28464 , w_28465 , \11179_b0 );
or ( \11181_b1 , \11096_b1 , \11100_b1 );
not ( \11100_b1 , w_28466 );
and ( \11181_b0 , \11096_b0 , w_28467 );
and ( w_28466 , w_28467 , \11100_b0 );
or ( \11182_b1 , \11100_b1 , \11105_b1 );
not ( \11105_b1 , w_28468 );
and ( \11182_b0 , \11100_b0 , w_28469 );
and ( w_28468 , w_28469 , \11105_b0 );
or ( \11183_b1 , \11096_b1 , \11105_b1 );
not ( \11105_b1 , w_28470 );
and ( \11183_b0 , \11096_b0 , w_28471 );
and ( w_28470 , w_28471 , \11105_b0 );
or ( \11185_b1 , \11081_b1 , \11085_b1 );
not ( \11085_b1 , w_28472 );
and ( \11185_b0 , \11081_b0 , w_28473 );
and ( w_28472 , w_28473 , \11085_b0 );
or ( \11186_b1 , \11085_b1 , \11090_b1 );
not ( \11090_b1 , w_28474 );
and ( \11186_b0 , \11085_b0 , w_28475 );
and ( w_28474 , w_28475 , \11090_b0 );
or ( \11187_b1 , \11081_b1 , \11090_b1 );
not ( \11090_b1 , w_28476 );
and ( \11187_b0 , \11081_b0 , w_28477 );
and ( w_28476 , w_28477 , \11090_b0 );
or ( \11189_b1 , \11184_b1 , \11188_b1 );
xor ( \11189_b0 , \11184_b0 , w_28478 );
not ( w_28478 , w_28479 );
and ( w_28479 , \11188_b1 , \11188_b0 );
or ( \11190_b1 , \11072_b1 , \11076_b1 );
not ( \11076_b1 , w_28480 );
and ( \11190_b0 , \11072_b0 , w_28481 );
and ( w_28480 , w_28481 , \11076_b0 );
or ( \11191_b1 , \11189_b1 , \11190_b1 );
xor ( \11191_b0 , \11189_b0 , w_28482 );
not ( w_28482 , w_28483 );
and ( w_28483 , \11190_b1 , \11190_b0 );
or ( \11192_b1 , \11180_b1 , \11191_b1 );
xor ( \11192_b0 , \11180_b0 , w_28484 );
not ( w_28484 , w_28485 );
and ( w_28485 , \11191_b1 , \11191_b0 );
or ( \11193_b1 , \11056_b1 , \11060_b1 );
not ( \11060_b1 , w_28486 );
and ( \11193_b0 , \11056_b0 , w_28487 );
and ( w_28486 , w_28487 , \11060_b0 );
or ( \11194_b1 , \11060_b1 , \11065_b1 );
not ( \11065_b1 , w_28488 );
and ( \11194_b0 , \11060_b0 , w_28489 );
and ( w_28488 , w_28489 , \11065_b0 );
or ( \11195_b1 , \11056_b1 , \11065_b1 );
not ( \11065_b1 , w_28490 );
and ( \11195_b0 , \11056_b0 , w_28491 );
and ( w_28490 , w_28491 , \11065_b0 );
or ( \11197_b1 , \11044_b1 , \11048_b1 );
not ( \11048_b1 , w_28492 );
and ( \11197_b0 , \11044_b0 , w_28493 );
and ( w_28492 , w_28493 , \11048_b0 );
or ( \11198_b1 , \11048_b1 , \11053_b1 );
not ( \11053_b1 , w_28494 );
and ( \11198_b0 , \11048_b0 , w_28495 );
and ( w_28494 , w_28495 , \11053_b0 );
or ( \11199_b1 , \11044_b1 , \11053_b1 );
not ( \11053_b1 , w_28496 );
and ( \11199_b0 , \11044_b0 , w_28497 );
and ( w_28496 , w_28497 , \11053_b0 );
or ( \11201_b1 , \11196_b1 , \11200_b1 );
xor ( \11201_b0 , \11196_b0 , w_28498 );
not ( w_28498 , w_28499 );
and ( w_28499 , \11200_b1 , \11200_b0 );
or ( \11202_b1 , \11030_b1 , \11034_b1 );
not ( \11034_b1 , w_28500 );
and ( \11202_b0 , \11030_b0 , w_28501 );
and ( w_28500 , w_28501 , \11034_b0 );
or ( \11203_b1 , \11034_b1 , \11039_b1 );
not ( \11039_b1 , w_28502 );
and ( \11203_b0 , \11034_b0 , w_28503 );
and ( w_28502 , w_28503 , \11039_b0 );
or ( \11204_b1 , \11030_b1 , \11039_b1 );
not ( \11039_b1 , w_28504 );
and ( \11204_b0 , \11030_b0 , w_28505 );
and ( w_28504 , w_28505 , \11039_b0 );
or ( \11206_b1 , \11201_b1 , \11205_b1 );
xor ( \11206_b0 , \11201_b0 , w_28506 );
not ( w_28506 , w_28507 );
and ( w_28507 , \11205_b1 , \11205_b0 );
or ( \11207_b1 , \11192_b1 , \11206_b1 );
xor ( \11207_b0 , \11192_b0 , w_28508 );
not ( w_28508 , w_28509 );
and ( w_28509 , \11206_b1 , \11206_b0 );
or ( \11208_b1 , \11040_b1 , \11054_b1 );
not ( \11054_b1 , w_28510 );
and ( \11208_b0 , \11040_b0 , w_28511 );
and ( w_28510 , w_28511 , \11054_b0 );
or ( \11209_b1 , \11054_b1 , \11066_b1 );
not ( \11066_b1 , w_28512 );
and ( \11209_b0 , \11054_b0 , w_28513 );
and ( w_28512 , w_28513 , \11066_b0 );
or ( \11210_b1 , \11040_b1 , \11066_b1 );
not ( \11066_b1 , w_28514 );
and ( \11210_b0 , \11040_b0 , w_28515 );
and ( w_28514 , w_28515 , \11066_b0 );
or ( \11212_b1 , \5737_b1 , \7175_b1 );
not ( \7175_b1 , w_28516 );
and ( \11212_b0 , \5737_b0 , w_28517 );
and ( w_28516 , w_28517 , \7175_b0 );
buf ( \11213_b1 , \11212_b1 );
not ( \11213_b1 , w_28518 );
not ( \11213_b0 , w_28519 );
and ( w_28518 , w_28519 , \11212_b0 );
or ( \11214_b1 , \11213_b1 , w_28520 );
xor ( \11214_b0 , \11213_b0 , w_28522 );
not ( w_28522 , w_28523 );
and ( w_28523 , w_28520 , w_28521 );
buf ( w_28520 , \7181_b1 );
not ( w_28520 , w_28524 );
not ( w_28521 , w_28525 );
and ( w_28524 , w_28525 , \7181_b0 );
or ( \11215_b1 , \6023_b1 , \11214_b1 );
xor ( \11215_b0 , \6023_b0 , w_28526 );
not ( w_28526 , w_28527 );
and ( w_28527 , \11214_b1 , \11214_b0 );
or ( \11216_b1 , \5758_b1 , \7192_b1 );
not ( \7192_b1 , w_28528 );
and ( \11216_b0 , \5758_b0 , w_28529 );
and ( w_28528 , w_28529 , \7192_b0 );
or ( \11217_b1 , \5770_b1 , \7190_b1 );
not ( \7190_b1 , w_28530 );
and ( \11217_b0 , \5770_b0 , w_28531 );
and ( w_28530 , w_28531 , \7190_b0 );
or ( \11218_b1 , \11216_b1 , w_28533 );
not ( w_28533 , w_28534 );
and ( \11218_b0 , \11216_b0 , w_28535 );
and ( w_28534 ,  , w_28535 );
buf ( w_28533 , \11217_b1 );
not ( w_28533 , w_28536 );
not (  , w_28537 );
and ( w_28536 , w_28537 , \11217_b0 );
or ( \11219_b1 , \11218_b1 , w_28538 );
xor ( \11219_b0 , \11218_b0 , w_28540 );
not ( w_28540 , w_28541 );
and ( w_28541 , w_28538 , w_28539 );
buf ( w_28538 , \7198_b1 );
not ( w_28538 , w_28542 );
not ( w_28539 , w_28543 );
and ( w_28542 , w_28543 , \7198_b0 );
or ( \11220_b1 , \11215_b1 , \11219_b1 );
xor ( \11220_b0 , \11215_b0 , w_28544 );
not ( w_28544 , w_28545 );
and ( w_28545 , \11219_b1 , \11219_b0 );
or ( \11221_b1 , \11211_b1 , \11220_b1 );
xor ( \11221_b0 , \11211_b0 , w_28546 );
not ( w_28546 , w_28547 );
and ( w_28547 , \11220_b1 , \11220_b0 );
or ( \11222_b1 , \5906_b1 , \5852_b1 );
not ( \5852_b1 , w_28548 );
and ( \11222_b0 , \5906_b0 , w_28549 );
and ( w_28548 , w_28549 , \5852_b0 );
or ( \11223_b1 , \5918_b1 , \5850_b1 );
not ( \5850_b1 , w_28550 );
and ( \11223_b0 , \5918_b0 , w_28551 );
and ( w_28550 , w_28551 , \5850_b0 );
or ( \11224_b1 , \11222_b1 , w_28553 );
not ( w_28553 , w_28554 );
and ( \11224_b0 , \11222_b0 , w_28555 );
and ( w_28554 ,  , w_28555 );
buf ( w_28553 , \11223_b1 );
not ( w_28553 , w_28556 );
not (  , w_28557 );
and ( w_28556 , w_28557 , \11223_b0 );
or ( \11225_b1 , \11224_b1 , w_28558 );
xor ( \11225_b0 , \11224_b0 , w_28560 );
not ( w_28560 , w_28561 );
and ( w_28561 , w_28558 , w_28559 );
buf ( w_28558 , \5859_b1 );
not ( w_28558 , w_28562 );
not ( w_28559 , w_28563 );
and ( w_28562 , w_28563 , \5859_b0 );
or ( \11226_b1 , \5925_b1 , \5871_b1 );
not ( \5871_b1 , w_28564 );
and ( \11226_b0 , \5925_b0 , w_28565 );
and ( w_28564 , w_28565 , \5871_b0 );
or ( \11227_b1 , \5937_b1 , \5869_b1 );
not ( \5869_b1 , w_28566 );
and ( \11227_b0 , \5937_b0 , w_28567 );
and ( w_28566 , w_28567 , \5869_b0 );
or ( \11228_b1 , \11226_b1 , w_28569 );
not ( w_28569 , w_28570 );
and ( \11228_b0 , \11226_b0 , w_28571 );
and ( w_28570 ,  , w_28571 );
buf ( w_28569 , \11227_b1 );
not ( w_28569 , w_28572 );
not (  , w_28573 );
and ( w_28572 , w_28573 , \11227_b0 );
or ( \11229_b1 , \11228_b1 , w_28574 );
xor ( \11229_b0 , \11228_b0 , w_28576 );
not ( w_28576 , w_28577 );
and ( w_28577 , w_28574 , w_28575 );
buf ( w_28574 , \5878_b1 );
not ( w_28574 , w_28578 );
not ( w_28575 , w_28579 );
and ( w_28578 , w_28579 , \5878_b0 );
or ( \11230_b1 , \11225_b1 , \11229_b1 );
xor ( \11230_b0 , \11225_b0 , w_28580 );
not ( w_28580 , w_28581 );
and ( w_28581 , \11229_b1 , \11229_b0 );
or ( \11231_b1 , \5945_b1 , \5891_b1 );
not ( \5891_b1 , w_28582 );
and ( \11231_b0 , \5945_b0 , w_28583 );
and ( w_28582 , w_28583 , \5891_b0 );
or ( \11232_b1 , \5957_b1 , \5889_b1 );
not ( \5889_b1 , w_28584 );
and ( \11232_b0 , \5957_b0 , w_28585 );
and ( w_28584 , w_28585 , \5889_b0 );
or ( \11233_b1 , \11231_b1 , w_28587 );
not ( w_28587 , w_28588 );
and ( \11233_b0 , \11231_b0 , w_28589 );
and ( w_28588 ,  , w_28589 );
buf ( w_28587 , \11232_b1 );
not ( w_28587 , w_28590 );
not (  , w_28591 );
and ( w_28590 , w_28591 , \11232_b0 );
or ( \11234_b1 , \11233_b1 , w_28592 );
xor ( \11234_b0 , \11233_b0 , w_28594 );
not ( w_28594 , w_28595 );
and ( w_28595 , w_28592 , w_28593 );
buf ( w_28592 , \5898_b1 );
not ( w_28592 , w_28596 );
not ( w_28593 , w_28597 );
and ( w_28596 , w_28597 , \5898_b0 );
or ( \11235_b1 , \11230_b1 , \11234_b1 );
xor ( \11235_b0 , \11230_b0 , w_28598 );
not ( w_28598 , w_28599 );
and ( w_28599 , \11234_b1 , \11234_b0 );
or ( \11236_b1 , \5842_b1 , \5790_b1 );
not ( \5790_b1 , w_28600 );
and ( \11236_b0 , \5842_b0 , w_28601 );
and ( w_28600 , w_28601 , \5790_b0 );
or ( \11237_b1 , \5854_b1 , \5788_b1 );
not ( \5788_b1 , w_28602 );
and ( \11237_b0 , \5854_b0 , w_28603 );
and ( w_28602 , w_28603 , \5788_b0 );
or ( \11238_b1 , \11236_b1 , w_28605 );
not ( w_28605 , w_28606 );
and ( \11238_b0 , \11236_b0 , w_28607 );
and ( w_28606 ,  , w_28607 );
buf ( w_28605 , \11237_b1 );
not ( w_28605 , w_28608 );
not (  , w_28609 );
and ( w_28608 , w_28609 , \11237_b0 );
or ( \11239_b1 , \11238_b1 , w_28610 );
xor ( \11239_b0 , \11238_b0 , w_28612 );
not ( w_28612 , w_28613 );
and ( w_28613 , w_28610 , w_28611 );
buf ( w_28610 , \5797_b1 );
not ( w_28610 , w_28614 );
not ( w_28611 , w_28615 );
and ( w_28614 , w_28615 , \5797_b0 );
or ( \11240_b1 , \5861_b1 , \5809_b1 );
not ( \5809_b1 , w_28616 );
and ( \11240_b0 , \5861_b0 , w_28617 );
and ( w_28616 , w_28617 , \5809_b0 );
or ( \11241_b1 , \5873_b1 , \5807_b1 );
not ( \5807_b1 , w_28618 );
and ( \11241_b0 , \5873_b0 , w_28619 );
and ( w_28618 , w_28619 , \5807_b0 );
or ( \11242_b1 , \11240_b1 , w_28621 );
not ( w_28621 , w_28622 );
and ( \11242_b0 , \11240_b0 , w_28623 );
and ( w_28622 ,  , w_28623 );
buf ( w_28621 , \11241_b1 );
not ( w_28621 , w_28624 );
not (  , w_28625 );
and ( w_28624 , w_28625 , \11241_b0 );
or ( \11243_b1 , \11242_b1 , w_28626 );
xor ( \11243_b0 , \11242_b0 , w_28628 );
not ( w_28628 , w_28629 );
and ( w_28629 , w_28626 , w_28627 );
buf ( w_28626 , \5816_b1 );
not ( w_28626 , w_28630 );
not ( w_28627 , w_28631 );
and ( w_28630 , w_28631 , \5816_b0 );
or ( \11244_b1 , \11239_b1 , \11243_b1 );
xor ( \11244_b0 , \11239_b0 , w_28632 );
not ( w_28632 , w_28633 );
and ( w_28633 , \11243_b1 , \11243_b0 );
or ( \11245_b1 , \5881_b1 , \5829_b1 );
not ( \5829_b1 , w_28634 );
and ( \11245_b0 , \5881_b0 , w_28635 );
and ( w_28634 , w_28635 , \5829_b0 );
or ( \11246_b1 , \5893_b1 , \5827_b1 );
not ( \5827_b1 , w_28636 );
and ( \11246_b0 , \5893_b0 , w_28637 );
and ( w_28636 , w_28637 , \5827_b0 );
or ( \11247_b1 , \11245_b1 , w_28639 );
not ( w_28639 , w_28640 );
and ( \11247_b0 , \11245_b0 , w_28641 );
and ( w_28640 ,  , w_28641 );
buf ( w_28639 , \11246_b1 );
not ( w_28639 , w_28642 );
not (  , w_28643 );
and ( w_28642 , w_28643 , \11246_b0 );
or ( \11248_b1 , \11247_b1 , w_28644 );
xor ( \11248_b0 , \11247_b0 , w_28646 );
not ( w_28646 , w_28647 );
and ( w_28647 , w_28644 , w_28645 );
buf ( w_28644 , \5836_b1 );
not ( w_28644 , w_28648 );
not ( w_28645 , w_28649 );
and ( w_28648 , w_28649 , \5836_b0 );
or ( \11249_b1 , \11244_b1 , \11248_b1 );
xor ( \11249_b0 , \11244_b0 , w_28650 );
not ( w_28650 , w_28651 );
and ( w_28651 , \11248_b1 , \11248_b0 );
or ( \11250_b1 , \11235_b1 , \11249_b1 );
xor ( \11250_b0 , \11235_b0 , w_28652 );
not ( w_28652 , w_28653 );
and ( w_28653 , \11249_b1 , \11249_b0 );
or ( \11251_b1 , \5780_b1 , \7203_b1 );
not ( \7203_b1 , w_28654 );
and ( \11251_b0 , \5780_b0 , w_28655 );
and ( w_28654 , w_28655 , \7203_b0 );
or ( \11252_b1 , \5792_b1 , \7201_b1 );
not ( \7201_b1 , w_28656 );
and ( \11252_b0 , \5792_b0 , w_28657 );
and ( w_28656 , w_28657 , \7201_b0 );
or ( \11253_b1 , \11251_b1 , w_28659 );
not ( w_28659 , w_28660 );
and ( \11253_b0 , \11251_b0 , w_28661 );
and ( w_28660 ,  , w_28661 );
buf ( w_28659 , \11252_b1 );
not ( w_28659 , w_28662 );
not (  , w_28663 );
and ( w_28662 , w_28663 , \11252_b0 );
or ( \11254_b1 , \11253_b1 , w_28664 );
xor ( \11254_b0 , \11253_b0 , w_28666 );
not ( w_28666 , w_28667 );
and ( w_28667 , w_28664 , w_28665 );
buf ( w_28664 , \6824_b1 );
not ( w_28664 , w_28668 );
not ( w_28665 , w_28669 );
and ( w_28668 , w_28669 , \6824_b0 );
or ( \11255_b1 , \5799_b1 , \5750_b1 );
not ( \5750_b1 , w_28670 );
and ( \11255_b0 , \5799_b0 , w_28671 );
and ( w_28670 , w_28671 , \5750_b0 );
or ( \11256_b1 , \5811_b1 , \5748_b1 );
not ( \5748_b1 , w_28672 );
and ( \11256_b0 , \5811_b0 , w_28673 );
and ( w_28672 , w_28673 , \5748_b0 );
or ( \11257_b1 , \11255_b1 , w_28675 );
not ( w_28675 , w_28676 );
and ( \11257_b0 , \11255_b0 , w_28677 );
and ( w_28676 ,  , w_28677 );
buf ( w_28675 , \11256_b1 );
not ( w_28675 , w_28678 );
not (  , w_28679 );
and ( w_28678 , w_28679 , \11256_b0 );
or ( \11258_b1 , \11257_b1 , w_28680 );
xor ( \11258_b0 , \11257_b0 , w_28682 );
not ( w_28682 , w_28683 );
and ( w_28683 , w_28680 , w_28681 );
buf ( w_28680 , \5755_b1 );
not ( w_28680 , w_28684 );
not ( w_28681 , w_28685 );
and ( w_28684 , w_28685 , \5755_b0 );
or ( \11259_b1 , \11254_b1 , \11258_b1 );
xor ( \11259_b0 , \11254_b0 , w_28686 );
not ( w_28686 , w_28687 );
and ( w_28687 , \11258_b1 , \11258_b0 );
or ( \11260_b1 , \5819_b1 , \5768_b1 );
not ( \5768_b1 , w_28688 );
and ( \11260_b0 , \5819_b0 , w_28689 );
and ( w_28688 , w_28689 , \5768_b0 );
or ( \11261_b1 , \5831_b1 , \5766_b1 );
not ( \5766_b1 , w_28690 );
and ( \11261_b0 , \5831_b0 , w_28691 );
and ( w_28690 , w_28691 , \5766_b0 );
or ( \11262_b1 , \11260_b1 , w_28693 );
not ( w_28693 , w_28694 );
and ( \11262_b0 , \11260_b0 , w_28695 );
and ( w_28694 ,  , w_28695 );
buf ( w_28693 , \11261_b1 );
not ( w_28693 , w_28696 );
not (  , w_28697 );
and ( w_28696 , w_28697 , \11261_b0 );
or ( \11263_b1 , \11262_b1 , w_28698 );
xor ( \11263_b0 , \11262_b0 , w_28700 );
not ( w_28700 , w_28701 );
and ( w_28701 , w_28698 , w_28699 );
buf ( w_28698 , \5775_b1 );
not ( w_28698 , w_28702 );
not ( w_28699 , w_28703 );
and ( w_28702 , w_28703 , \5775_b0 );
or ( \11264_b1 , \11259_b1 , \11263_b1 );
xor ( \11264_b0 , \11259_b0 , w_28704 );
not ( w_28704 , w_28705 );
and ( w_28705 , \11263_b1 , \11263_b0 );
or ( \11265_b1 , \11250_b1 , \11264_b1 );
xor ( \11265_b0 , \11250_b0 , w_28706 );
not ( w_28706 , w_28707 );
and ( w_28707 , \11264_b1 , \11264_b0 );
or ( \11266_b1 , \11221_b1 , \11265_b1 );
xor ( \11266_b0 , \11221_b0 , w_28708 );
not ( w_28708 , w_28709 );
and ( w_28709 , \11265_b1 , \11265_b0 );
or ( \11267_b1 , \11207_b1 , \11266_b1 );
xor ( \11267_b0 , \11207_b0 , w_28710 );
not ( w_28710 , w_28711 );
and ( w_28711 , \11266_b1 , \11266_b0 );
or ( \11268_b1 , \11011_b1 , \11015_b1 );
not ( \11015_b1 , w_28712 );
and ( \11268_b0 , \11011_b0 , w_28713 );
and ( w_28712 , w_28713 , \11015_b0 );
or ( \11269_b1 , \11015_b1 , \11020_b1 );
not ( \11020_b1 , w_28714 );
and ( \11269_b0 , \11015_b0 , w_28715 );
and ( w_28714 , w_28715 , \11020_b0 );
or ( \11270_b1 , \11011_b1 , \11020_b1 );
not ( \11020_b1 , w_28716 );
and ( \11270_b0 , \11011_b0 , w_28717 );
and ( w_28716 , w_28717 , \11020_b0 );
or ( \11272_b1 , \10997_b1 , \11001_b1 );
not ( \11001_b1 , w_28718 );
and ( \11272_b0 , \10997_b0 , w_28719 );
and ( w_28718 , w_28719 , \11001_b0 );
or ( \11273_b1 , \11001_b1 , \11006_b1 );
not ( \11006_b1 , w_28720 );
and ( \11273_b0 , \11001_b0 , w_28721 );
and ( w_28720 , w_28721 , \11006_b0 );
or ( \11274_b1 , \10997_b1 , \11006_b1 );
not ( \11006_b1 , w_28722 );
and ( \11274_b0 , \10997_b0 , w_28723 );
and ( w_28722 , w_28723 , \11006_b0 );
or ( \11276_b1 , \11271_b1 , \11275_b1 );
xor ( \11276_b0 , \11271_b0 , w_28724 );
not ( w_28724 , w_28725 );
and ( w_28725 , \11275_b1 , \11275_b0 );
or ( \11277_b1 , \11077_b1 , \11091_b1 );
not ( \11091_b1 , w_28726 );
and ( \11277_b0 , \11077_b0 , w_28727 );
and ( w_28726 , w_28727 , \11091_b0 );
or ( \11278_b1 , \11091_b1 , \11106_b1 );
not ( \11106_b1 , w_28728 );
and ( \11278_b0 , \11091_b0 , w_28729 );
and ( w_28728 , w_28729 , \11106_b0 );
or ( \11279_b1 , \11077_b1 , \11106_b1 );
not ( \11106_b1 , w_28730 );
and ( \11279_b0 , \11077_b0 , w_28731 );
and ( w_28730 , w_28731 , \11106_b0 );
or ( \11281_b1 , \11276_b1 , \11280_b1 );
xor ( \11281_b0 , \11276_b0 , w_28732 );
not ( w_28732 , w_28733 );
and ( w_28733 , \11280_b1 , \11280_b0 );
or ( \11282_b1 , \11267_b1 , \11281_b1 );
xor ( \11282_b0 , \11267_b0 , w_28734 );
not ( w_28734 , w_28735 );
and ( w_28735 , \11281_b1 , \11281_b0 );
or ( \11283_b1 , \11153_b1 , \11282_b1 );
xor ( \11283_b0 , \11153_b0 , w_28736 );
not ( w_28736 , w_28737 );
and ( w_28737 , \11282_b1 , \11282_b0 );
or ( \11284_b1 , \11144_b1 , \11283_b1 );
xor ( \11284_b0 , \11144_b0 , w_28738 );
not ( w_28738 , w_28739 );
and ( w_28739 , \11283_b1 , \11283_b0 );
or ( \11285_b1 , \10969_b1 , \10983_b1 );
not ( \10983_b1 , w_28740 );
and ( \11285_b0 , \10969_b0 , w_28741 );
and ( w_28740 , w_28741 , \10983_b0 );
or ( \11286_b1 , \10983_b1 , \11122_b1 );
not ( \11122_b1 , w_28742 );
and ( \11286_b0 , \10983_b0 , w_28743 );
and ( w_28742 , w_28743 , \11122_b0 );
or ( \11287_b1 , \10969_b1 , \11122_b1 );
not ( \11122_b1 , w_28744 );
and ( \11287_b0 , \10969_b0 , w_28745 );
and ( w_28744 , w_28745 , \11122_b0 );
or ( \11289_b1 , \11284_b1 , w_28747 );
not ( w_28747 , w_28748 );
and ( \11289_b0 , \11284_b0 , w_28749 );
and ( w_28748 ,  , w_28749 );
buf ( w_28747 , \11288_b1 );
not ( w_28747 , w_28750 );
not (  , w_28751 );
and ( w_28750 , w_28751 , \11288_b0 );
or ( \11290_b1 , \11128_b1 , w_28753 );
not ( w_28753 , w_28754 );
and ( \11290_b0 , \11128_b0 , w_28755 );
and ( w_28754 ,  , w_28755 );
buf ( w_28753 , \11289_b1 );
not ( w_28753 , w_28756 );
not (  , w_28757 );
and ( w_28756 , w_28757 , \11289_b0 );
or ( \11291_b1 , \11148_b1 , \11152_b1 );
not ( \11152_b1 , w_28758 );
and ( \11291_b0 , \11148_b0 , w_28759 );
and ( w_28758 , w_28759 , \11152_b0 );
or ( \11292_b1 , \11152_b1 , \11282_b1 );
not ( \11282_b1 , w_28760 );
and ( \11292_b0 , \11152_b0 , w_28761 );
and ( w_28760 , w_28761 , \11282_b0 );
or ( \11293_b1 , \11148_b1 , \11282_b1 );
not ( \11282_b1 , w_28762 );
and ( \11293_b0 , \11148_b0 , w_28763 );
and ( w_28762 , w_28763 , \11282_b0 );
or ( \11295_b1 , \11271_b1 , \11275_b1 );
not ( \11275_b1 , w_28764 );
and ( \11295_b0 , \11271_b0 , w_28765 );
and ( w_28764 , w_28765 , \11275_b0 );
or ( \11296_b1 , \11275_b1 , \11280_b1 );
not ( \11280_b1 , w_28766 );
and ( \11296_b0 , \11275_b0 , w_28767 );
and ( w_28766 , w_28767 , \11280_b0 );
or ( \11297_b1 , \11271_b1 , \11280_b1 );
not ( \11280_b1 , w_28768 );
and ( \11297_b0 , \11271_b0 , w_28769 );
and ( w_28768 , w_28769 , \11280_b0 );
or ( \11299_b1 , \11211_b1 , \11220_b1 );
not ( \11220_b1 , w_28770 );
and ( \11299_b0 , \11211_b0 , w_28771 );
and ( w_28770 , w_28771 , \11220_b0 );
or ( \11300_b1 , \11220_b1 , \11265_b1 );
not ( \11265_b1 , w_28772 );
and ( \11300_b0 , \11220_b0 , w_28773 );
and ( w_28772 , w_28773 , \11265_b0 );
or ( \11301_b1 , \11211_b1 , \11265_b1 );
not ( \11265_b1 , w_28774 );
and ( \11301_b0 , \11211_b0 , w_28775 );
and ( w_28774 , w_28775 , \11265_b0 );
or ( \11303_b1 , \11298_b1 , \11302_b1 );
xor ( \11303_b0 , \11298_b0 , w_28776 );
not ( w_28776 , w_28777 );
and ( w_28777 , \11302_b1 , \11302_b0 );
or ( \11304_b1 , \11180_b1 , \11191_b1 );
not ( \11191_b1 , w_28778 );
and ( \11304_b0 , \11180_b0 , w_28779 );
and ( w_28778 , w_28779 , \11191_b0 );
or ( \11305_b1 , \11191_b1 , \11206_b1 );
not ( \11206_b1 , w_28780 );
and ( \11305_b0 , \11191_b0 , w_28781 );
and ( w_28780 , w_28781 , \11206_b0 );
or ( \11306_b1 , \11180_b1 , \11206_b1 );
not ( \11206_b1 , w_28782 );
and ( \11306_b0 , \11180_b0 , w_28783 );
and ( w_28782 , w_28783 , \11206_b0 );
or ( \11308_b1 , \11303_b1 , \11307_b1 );
xor ( \11308_b0 , \11303_b0 , w_28784 );
not ( w_28784 , w_28785 );
and ( w_28785 , \11307_b1 , \11307_b0 );
or ( \11309_b1 , \11294_b1 , \11308_b1 );
xor ( \11309_b0 , \11294_b0 , w_28786 );
not ( w_28786 , w_28787 );
and ( w_28787 , \11308_b1 , \11308_b0 );
or ( \11310_b1 , \11136_b1 , \11140_b1 );
not ( \11140_b1 , w_28788 );
and ( \11310_b0 , \11136_b0 , w_28789 );
and ( w_28788 , w_28789 , \11140_b0 );
or ( \11311_b1 , \11140_b1 , \11142_b1 );
not ( \11142_b1 , w_28790 );
and ( \11311_b0 , \11140_b0 , w_28791 );
and ( w_28790 , w_28791 , \11142_b0 );
or ( \11312_b1 , \11136_b1 , \11142_b1 );
not ( \11142_b1 , w_28792 );
and ( \11312_b0 , \11136_b0 , w_28793 );
and ( w_28792 , w_28793 , \11142_b0 );
or ( \11314_b1 , \11207_b1 , \11266_b1 );
not ( \11266_b1 , w_28794 );
and ( \11314_b0 , \11207_b0 , w_28795 );
and ( w_28794 , w_28795 , \11266_b0 );
or ( \11315_b1 , \11266_b1 , \11281_b1 );
not ( \11281_b1 , w_28796 );
and ( \11315_b0 , \11266_b0 , w_28797 );
and ( w_28796 , w_28797 , \11281_b0 );
or ( \11316_b1 , \11207_b1 , \11281_b1 );
not ( \11281_b1 , w_28798 );
and ( \11316_b0 , \11207_b0 , w_28799 );
and ( w_28798 , w_28799 , \11281_b0 );
or ( \11318_b1 , \11313_b1 , \11317_b1 );
xor ( \11318_b0 , \11313_b0 , w_28800 );
not ( w_28800 , w_28801 );
and ( w_28801 , \11317_b1 , \11317_b0 );
or ( \11319_b1 , \11225_b1 , \11229_b1 );
not ( \11229_b1 , w_28802 );
and ( \11319_b0 , \11225_b0 , w_28803 );
and ( w_28802 , w_28803 , \11229_b0 );
or ( \11320_b1 , \11229_b1 , \11234_b1 );
not ( \11234_b1 , w_28804 );
and ( \11320_b0 , \11229_b0 , w_28805 );
and ( w_28804 , w_28805 , \11234_b0 );
or ( \11321_b1 , \11225_b1 , \11234_b1 );
not ( \11234_b1 , w_28806 );
and ( \11321_b0 , \11225_b0 , w_28807 );
and ( w_28806 , w_28807 , \11234_b0 );
or ( \11323_b1 , \11169_b1 , \11173_b1 );
not ( \11173_b1 , w_28808 );
and ( \11323_b0 , \11169_b0 , w_28809 );
and ( w_28808 , w_28809 , \11173_b0 );
or ( \11324_b1 , \11173_b1 , \11178_b1 );
not ( \11178_b1 , w_28810 );
and ( \11324_b0 , \11173_b0 , w_28811 );
and ( w_28810 , w_28811 , \11178_b0 );
or ( \11325_b1 , \11169_b1 , \11178_b1 );
not ( \11178_b1 , w_28812 );
and ( \11325_b0 , \11169_b0 , w_28813 );
and ( w_28812 , w_28813 , \11178_b0 );
or ( \11327_b1 , \11322_b1 , \11326_b1 );
xor ( \11327_b0 , \11322_b0 , w_28814 );
not ( w_28814 , w_28815 );
and ( w_28815 , \11326_b1 , \11326_b0 );
or ( \11328_b1 , \11157_b1 , \11161_b1 );
not ( \11161_b1 , w_28816 );
and ( \11328_b0 , \11157_b0 , w_28817 );
and ( w_28816 , w_28817 , \11161_b0 );
or ( \11329_b1 , \11161_b1 , \11164_b1 );
not ( \11164_b1 , w_28818 );
and ( \11329_b0 , \11161_b0 , w_28819 );
and ( w_28818 , w_28819 , \11164_b0 );
or ( \11330_b1 , \11157_b1 , \11164_b1 );
not ( \11164_b1 , w_28820 );
and ( \11330_b0 , \11157_b0 , w_28821 );
and ( w_28820 , w_28821 , \11164_b0 );
or ( \11332_b1 , \11327_b1 , \11331_b1 );
xor ( \11332_b0 , \11327_b0 , w_28822 );
not ( w_28822 , w_28823 );
and ( w_28823 , \11331_b1 , \11331_b0 );
or ( \11333_b1 , \6023_b1 , \11214_b1 );
not ( \11214_b1 , w_28824 );
and ( \11333_b0 , \6023_b0 , w_28825 );
and ( w_28824 , w_28825 , \11214_b0 );
or ( \11334_b1 , \11214_b1 , \11219_b1 );
not ( \11219_b1 , w_28826 );
and ( \11334_b0 , \11214_b0 , w_28827 );
and ( w_28826 , w_28827 , \11219_b0 );
or ( \11335_b1 , \6023_b1 , \11219_b1 );
not ( \11219_b1 , w_28828 );
and ( \11335_b0 , \6023_b0 , w_28829 );
and ( w_28828 , w_28829 , \11219_b0 );
or ( \11337_b1 , \11254_b1 , \11258_b1 );
not ( \11258_b1 , w_28830 );
and ( \11337_b0 , \11254_b0 , w_28831 );
and ( w_28830 , w_28831 , \11258_b0 );
or ( \11338_b1 , \11258_b1 , \11263_b1 );
not ( \11263_b1 , w_28832 );
and ( \11338_b0 , \11258_b0 , w_28833 );
and ( w_28832 , w_28833 , \11263_b0 );
or ( \11339_b1 , \11254_b1 , \11263_b1 );
not ( \11263_b1 , w_28834 );
and ( \11339_b0 , \11254_b0 , w_28835 );
and ( w_28834 , w_28835 , \11263_b0 );
or ( \11341_b1 , \11336_b1 , \11340_b1 );
xor ( \11341_b0 , \11336_b0 , w_28836 );
not ( w_28836 , w_28837 );
and ( w_28837 , \11340_b1 , \11340_b0 );
or ( \11342_b1 , \11239_b1 , \11243_b1 );
not ( \11243_b1 , w_28838 );
and ( \11342_b0 , \11239_b0 , w_28839 );
and ( w_28838 , w_28839 , \11243_b0 );
or ( \11343_b1 , \11243_b1 , \11248_b1 );
not ( \11248_b1 , w_28840 );
and ( \11343_b0 , \11243_b0 , w_28841 );
and ( w_28840 , w_28841 , \11248_b0 );
or ( \11344_b1 , \11239_b1 , \11248_b1 );
not ( \11248_b1 , w_28842 );
and ( \11344_b0 , \11239_b0 , w_28843 );
and ( w_28842 , w_28843 , \11248_b0 );
or ( \11346_b1 , \11341_b1 , \11345_b1 );
xor ( \11346_b0 , \11341_b0 , w_28844 );
not ( w_28844 , w_28845 );
and ( w_28845 , \11345_b1 , \11345_b0 );
or ( \11347_b1 , \11332_b1 , \11346_b1 );
xor ( \11347_b0 , \11332_b0 , w_28846 );
not ( w_28846 , w_28847 );
and ( w_28847 , \11346_b1 , \11346_b0 );
or ( \11348_b1 , \11235_b1 , \11249_b1 );
not ( \11249_b1 , w_28848 );
and ( \11348_b0 , \11235_b0 , w_28849 );
and ( w_28848 , w_28849 , \11249_b0 );
or ( \11349_b1 , \11249_b1 , \11264_b1 );
not ( \11264_b1 , w_28850 );
and ( \11349_b0 , \11249_b0 , w_28851 );
and ( w_28850 , w_28851 , \11264_b0 );
or ( \11350_b1 , \11235_b1 , \11264_b1 );
not ( \11264_b1 , w_28852 );
and ( \11350_b0 , \11235_b0 , w_28853 );
and ( w_28852 , w_28853 , \11264_b0 );
or ( \11352_b1 , \5873_b1 , \5809_b1 );
not ( \5809_b1 , w_28854 );
and ( \11352_b0 , \5873_b0 , w_28855 );
and ( w_28854 , w_28855 , \5809_b0 );
or ( \11353_b1 , \5842_b1 , \5807_b1 );
not ( \5807_b1 , w_28856 );
and ( \11353_b0 , \5842_b0 , w_28857 );
and ( w_28856 , w_28857 , \5807_b0 );
or ( \11354_b1 , \11352_b1 , w_28859 );
not ( w_28859 , w_28860 );
and ( \11354_b0 , \11352_b0 , w_28861 );
and ( w_28860 ,  , w_28861 );
buf ( w_28859 , \11353_b1 );
not ( w_28859 , w_28862 );
not (  , w_28863 );
and ( w_28862 , w_28863 , \11353_b0 );
or ( \11355_b1 , \11354_b1 , w_28864 );
xor ( \11355_b0 , \11354_b0 , w_28866 );
not ( w_28866 , w_28867 );
and ( w_28867 , w_28864 , w_28865 );
buf ( w_28864 , \5816_b1 );
not ( w_28864 , w_28868 );
not ( w_28865 , w_28869 );
and ( w_28868 , w_28869 , \5816_b0 );
or ( \11356_b1 , \5893_b1 , \5829_b1 );
not ( \5829_b1 , w_28870 );
and ( \11356_b0 , \5893_b0 , w_28871 );
and ( w_28870 , w_28871 , \5829_b0 );
or ( \11357_b1 , \5861_b1 , \5827_b1 );
not ( \5827_b1 , w_28872 );
and ( \11357_b0 , \5861_b0 , w_28873 );
and ( w_28872 , w_28873 , \5827_b0 );
or ( \11358_b1 , \11356_b1 , w_28875 );
not ( w_28875 , w_28876 );
and ( \11358_b0 , \11356_b0 , w_28877 );
and ( w_28876 ,  , w_28877 );
buf ( w_28875 , \11357_b1 );
not ( w_28875 , w_28878 );
not (  , w_28879 );
and ( w_28878 , w_28879 , \11357_b0 );
or ( \11359_b1 , \11358_b1 , w_28880 );
xor ( \11359_b0 , \11358_b0 , w_28882 );
not ( w_28882 , w_28883 );
and ( w_28883 , w_28880 , w_28881 );
buf ( w_28880 , \5836_b1 );
not ( w_28880 , w_28884 );
not ( w_28881 , w_28885 );
and ( w_28884 , w_28885 , \5836_b0 );
or ( \11360_b1 , \11355_b1 , \11359_b1 );
xor ( \11360_b0 , \11355_b0 , w_28886 );
not ( w_28886 , w_28887 );
and ( w_28887 , \11359_b1 , \11359_b0 );
or ( \11361_b1 , \5918_b1 , \5852_b1 );
not ( \5852_b1 , w_28888 );
and ( \11361_b0 , \5918_b0 , w_28889 );
and ( w_28888 , w_28889 , \5852_b0 );
or ( \11362_b1 , \5881_b1 , \5850_b1 );
not ( \5850_b1 , w_28890 );
and ( \11362_b0 , \5881_b0 , w_28891 );
and ( w_28890 , w_28891 , \5850_b0 );
or ( \11363_b1 , \11361_b1 , w_28893 );
not ( w_28893 , w_28894 );
and ( \11363_b0 , \11361_b0 , w_28895 );
and ( w_28894 ,  , w_28895 );
buf ( w_28893 , \11362_b1 );
not ( w_28893 , w_28896 );
not (  , w_28897 );
and ( w_28896 , w_28897 , \11362_b0 );
or ( \11364_b1 , \11363_b1 , w_28898 );
xor ( \11364_b0 , \11363_b0 , w_28900 );
not ( w_28900 , w_28901 );
and ( w_28901 , w_28898 , w_28899 );
buf ( w_28898 , \5859_b1 );
not ( w_28898 , w_28902 );
not ( w_28899 , w_28903 );
and ( w_28902 , w_28903 , \5859_b0 );
or ( \11365_b1 , \11360_b1 , \11364_b1 );
xor ( \11365_b0 , \11360_b0 , w_28904 );
not ( w_28904 , w_28905 );
and ( w_28905 , \11364_b1 , \11364_b0 );
or ( \11366_b1 , \5811_b1 , \5750_b1 );
not ( \5750_b1 , w_28906 );
and ( \11366_b0 , \5811_b0 , w_28907 );
and ( w_28906 , w_28907 , \5750_b0 );
or ( \11367_b1 , \5780_b1 , \5748_b1 );
not ( \5748_b1 , w_28908 );
and ( \11367_b0 , \5780_b0 , w_28909 );
and ( w_28908 , w_28909 , \5748_b0 );
or ( \11368_b1 , \11366_b1 , w_28911 );
not ( w_28911 , w_28912 );
and ( \11368_b0 , \11366_b0 , w_28913 );
and ( w_28912 ,  , w_28913 );
buf ( w_28911 , \11367_b1 );
not ( w_28911 , w_28914 );
not (  , w_28915 );
and ( w_28914 , w_28915 , \11367_b0 );
or ( \11369_b1 , \11368_b1 , w_28916 );
xor ( \11369_b0 , \11368_b0 , w_28918 );
not ( w_28918 , w_28919 );
and ( w_28919 , w_28916 , w_28917 );
buf ( w_28916 , \5755_b1 );
not ( w_28916 , w_28920 );
not ( w_28917 , w_28921 );
and ( w_28920 , w_28921 , \5755_b0 );
or ( \11370_b1 , \5831_b1 , \5768_b1 );
not ( \5768_b1 , w_28922 );
and ( \11370_b0 , \5831_b0 , w_28923 );
and ( w_28922 , w_28923 , \5768_b0 );
or ( \11371_b1 , \5799_b1 , \5766_b1 );
not ( \5766_b1 , w_28924 );
and ( \11371_b0 , \5799_b0 , w_28925 );
and ( w_28924 , w_28925 , \5766_b0 );
or ( \11372_b1 , \11370_b1 , w_28927 );
not ( w_28927 , w_28928 );
and ( \11372_b0 , \11370_b0 , w_28929 );
and ( w_28928 ,  , w_28929 );
buf ( w_28927 , \11371_b1 );
not ( w_28927 , w_28930 );
not (  , w_28931 );
and ( w_28930 , w_28931 , \11371_b0 );
or ( \11373_b1 , \11372_b1 , w_28932 );
xor ( \11373_b0 , \11372_b0 , w_28934 );
not ( w_28934 , w_28935 );
and ( w_28935 , w_28932 , w_28933 );
buf ( w_28932 , \5775_b1 );
not ( w_28932 , w_28936 );
not ( w_28933 , w_28937 );
and ( w_28936 , w_28937 , \5775_b0 );
or ( \11374_b1 , \11369_b1 , \11373_b1 );
xor ( \11374_b0 , \11369_b0 , w_28938 );
not ( w_28938 , w_28939 );
and ( w_28939 , \11373_b1 , \11373_b0 );
or ( \11375_b1 , \5854_b1 , \5790_b1 );
not ( \5790_b1 , w_28940 );
and ( \11375_b0 , \5854_b0 , w_28941 );
and ( w_28940 , w_28941 , \5790_b0 );
or ( \11376_b1 , \5819_b1 , \5788_b1 );
not ( \5788_b1 , w_28942 );
and ( \11376_b0 , \5819_b0 , w_28943 );
and ( w_28942 , w_28943 , \5788_b0 );
or ( \11377_b1 , \11375_b1 , w_28945 );
not ( w_28945 , w_28946 );
and ( \11377_b0 , \11375_b0 , w_28947 );
and ( w_28946 ,  , w_28947 );
buf ( w_28945 , \11376_b1 );
not ( w_28945 , w_28948 );
not (  , w_28949 );
and ( w_28948 , w_28949 , \11376_b0 );
or ( \11378_b1 , \11377_b1 , w_28950 );
xor ( \11378_b0 , \11377_b0 , w_28952 );
not ( w_28952 , w_28953 );
and ( w_28953 , w_28950 , w_28951 );
buf ( w_28950 , \5797_b1 );
not ( w_28950 , w_28954 );
not ( w_28951 , w_28955 );
and ( w_28954 , w_28955 , \5797_b0 );
or ( \11379_b1 , \11374_b1 , \11378_b1 );
xor ( \11379_b0 , \11374_b0 , w_28956 );
not ( w_28956 , w_28957 );
and ( w_28957 , \11378_b1 , \11378_b0 );
or ( \11380_b1 , \11365_b1 , \11379_b1 );
xor ( \11380_b0 , \11365_b0 , w_28958 );
not ( w_28958 , w_28959 );
and ( w_28959 , \11379_b1 , \11379_b0 );
buf ( \11381_b1 , \7181_b1 );
not ( \11381_b1 , w_28960 );
not ( \11381_b0 , w_28961 );
and ( w_28960 , w_28961 , \7181_b0 );
or ( \11382_b1 , \5770_b1 , \7192_b1 );
not ( \7192_b1 , w_28962 );
and ( \11382_b0 , \5770_b0 , w_28963 );
and ( w_28962 , w_28963 , \7192_b0 );
or ( \11383_b1 , \5737_b1 , \7190_b1 );
not ( \7190_b1 , w_28964 );
and ( \11383_b0 , \5737_b0 , w_28965 );
and ( w_28964 , w_28965 , \7190_b0 );
or ( \11384_b1 , \11382_b1 , w_28967 );
not ( w_28967 , w_28968 );
and ( \11384_b0 , \11382_b0 , w_28969 );
and ( w_28968 ,  , w_28969 );
buf ( w_28967 , \11383_b1 );
not ( w_28967 , w_28970 );
not (  , w_28971 );
and ( w_28970 , w_28971 , \11383_b0 );
or ( \11385_b1 , \11384_b1 , w_28972 );
xor ( \11385_b0 , \11384_b0 , w_28974 );
not ( w_28974 , w_28975 );
and ( w_28975 , w_28972 , w_28973 );
buf ( w_28972 , \7198_b1 );
not ( w_28972 , w_28976 );
not ( w_28973 , w_28977 );
and ( w_28976 , w_28977 , \7198_b0 );
or ( \11386_b1 , \11381_b1 , \11385_b1 );
xor ( \11386_b0 , \11381_b0 , w_28978 );
not ( w_28978 , w_28979 );
and ( w_28979 , \11385_b1 , \11385_b0 );
or ( \11387_b1 , \5792_b1 , \7203_b1 );
not ( \7203_b1 , w_28980 );
and ( \11387_b0 , \5792_b0 , w_28981 );
and ( w_28980 , w_28981 , \7203_b0 );
or ( \11388_b1 , \5758_b1 , \7201_b1 );
not ( \7201_b1 , w_28982 );
and ( \11388_b0 , \5758_b0 , w_28983 );
and ( w_28982 , w_28983 , \7201_b0 );
or ( \11389_b1 , \11387_b1 , w_28985 );
not ( w_28985 , w_28986 );
and ( \11389_b0 , \11387_b0 , w_28987 );
and ( w_28986 ,  , w_28987 );
buf ( w_28985 , \11388_b1 );
not ( w_28985 , w_28988 );
not (  , w_28989 );
and ( w_28988 , w_28989 , \11388_b0 );
or ( \11390_b1 , \11389_b1 , w_28990 );
xor ( \11390_b0 , \11389_b0 , w_28992 );
not ( w_28992 , w_28993 );
and ( w_28993 , w_28990 , w_28991 );
buf ( w_28990 , \6824_b1 );
not ( w_28990 , w_28994 );
not ( w_28991 , w_28995 );
and ( w_28994 , w_28995 , \6824_b0 );
or ( \11391_b1 , \11386_b1 , \11390_b1 );
xor ( \11391_b0 , \11386_b0 , w_28996 );
not ( w_28996 , w_28997 );
and ( w_28997 , \11390_b1 , \11390_b0 );
or ( \11392_b1 , \11380_b1 , \11391_b1 );
xor ( \11392_b0 , \11380_b0 , w_28998 );
not ( w_28998 , w_28999 );
and ( w_28999 , \11391_b1 , \11391_b0 );
or ( \11393_b1 , \11351_b1 , \11392_b1 );
xor ( \11393_b0 , \11351_b0 , w_29000 );
not ( w_29000 , w_29001 );
and ( w_29001 , \11392_b1 , \11392_b0 );
or ( \11394_b1 , \6057_b1 , \5996_b1 );
not ( \5996_b1 , w_29002 );
and ( \11394_b0 , \6057_b0 , w_29003 );
and ( w_29002 , w_29003 , \5996_b0 );
or ( \11395_b1 , \6029_b1 , \5994_b1 );
not ( \5994_b1 , w_29004 );
and ( \11395_b0 , \6029_b0 , w_29005 );
and ( w_29004 , w_29005 , \5994_b0 );
or ( \11396_b1 , \11394_b1 , w_29007 );
not ( w_29007 , w_29008 );
and ( \11396_b0 , \11394_b0 , w_29009 );
and ( w_29008 ,  , w_29009 );
buf ( w_29007 , \11395_b1 );
not ( w_29007 , w_29010 );
not (  , w_29011 );
and ( w_29010 , w_29011 , \11395_b0 );
or ( \11397_b1 , \11396_b1 , w_29012 );
xor ( \11397_b0 , \11396_b0 , w_29014 );
not ( w_29014 , w_29015 );
and ( w_29015 , w_29012 , w_29013 );
buf ( w_29012 , \6003_b1 );
not ( w_29012 , w_29016 );
not ( w_29013 , w_29017 );
and ( w_29016 , w_29017 , \6003_b0 );
or ( \11398_b1 , \6065_b1 , \6016_b1 );
not ( \6016_b1 , w_29018 );
and ( \11398_b0 , \6065_b0 , w_29019 );
and ( w_29018 , w_29019 , \6016_b0 );
or ( \11399_b1 , \6048_b1 , \6014_b1 );
not ( \6014_b1 , w_29020 );
and ( \11399_b0 , \6048_b0 , w_29021 );
and ( w_29020 , w_29021 , \6014_b0 );
or ( \11400_b1 , \11398_b1 , w_29023 );
not ( w_29023 , w_29024 );
and ( \11400_b0 , \11398_b0 , w_29025 );
and ( w_29024 ,  , w_29025 );
buf ( w_29023 , \11399_b1 );
not ( w_29023 , w_29026 );
not (  , w_29027 );
and ( w_29026 , w_29027 , \11399_b0 );
or ( \11401_b1 , \11400_b1 , w_29028 );
xor ( \11401_b0 , \11400_b0 , w_29030 );
not ( w_29030 , w_29031 );
and ( w_29031 , w_29028 , w_29029 );
buf ( w_29028 , \6023_b1 );
not ( w_29028 , w_29032 );
not ( w_29029 , w_29033 );
and ( w_29032 , w_29033 , \6023_b0 );
or ( \11402_b1 , \11397_b1 , \11401_b1 );
xor ( \11402_b0 , \11397_b0 , w_29034 );
not ( w_29034 , w_29035 );
and ( w_29035 , \11401_b1 , \11401_b0 );
or ( \11403_b1 , \5998_b1 , \5935_b1 );
not ( \5935_b1 , w_29036 );
and ( \11403_b0 , \5998_b0 , w_29037 );
and ( w_29036 , w_29037 , \5935_b0 );
or ( \11404_b1 , \5967_b1 , \5933_b1 );
not ( \5933_b1 , w_29038 );
and ( \11404_b0 , \5967_b0 , w_29039 );
and ( w_29038 , w_29039 , \5933_b0 );
or ( \11405_b1 , \11403_b1 , w_29041 );
not ( w_29041 , w_29042 );
and ( \11405_b0 , \11403_b0 , w_29043 );
and ( w_29042 ,  , w_29043 );
buf ( w_29041 , \11404_b1 );
not ( w_29041 , w_29044 );
not (  , w_29045 );
and ( w_29044 , w_29045 , \11404_b0 );
or ( \11406_b1 , \11405_b1 , w_29046 );
xor ( \11406_b0 , \11405_b0 , w_29048 );
not ( w_29048 , w_29049 );
and ( w_29049 , w_29046 , w_29047 );
buf ( w_29046 , \5942_b1 );
not ( w_29046 , w_29050 );
not ( w_29047 , w_29051 );
and ( w_29050 , w_29051 , \5942_b0 );
or ( \11407_b1 , \6018_b1 , \5955_b1 );
not ( \5955_b1 , w_29052 );
and ( \11407_b0 , \6018_b0 , w_29053 );
and ( w_29052 , w_29053 , \5955_b0 );
or ( \11408_b1 , \5986_b1 , \5953_b1 );
not ( \5953_b1 , w_29054 );
and ( \11408_b0 , \5986_b0 , w_29055 );
and ( w_29054 , w_29055 , \5953_b0 );
or ( \11409_b1 , \11407_b1 , w_29057 );
not ( w_29057 , w_29058 );
and ( \11409_b0 , \11407_b0 , w_29059 );
and ( w_29058 ,  , w_29059 );
buf ( w_29057 , \11408_b1 );
not ( w_29057 , w_29060 );
not (  , w_29061 );
and ( w_29060 , w_29061 , \11408_b0 );
or ( \11410_b1 , \11409_b1 , w_29062 );
xor ( \11410_b0 , \11409_b0 , w_29064 );
not ( w_29064 , w_29065 );
and ( w_29065 , w_29062 , w_29063 );
buf ( w_29062 , \5962_b1 );
not ( w_29062 , w_29066 );
not ( w_29063 , w_29067 );
and ( w_29066 , w_29067 , \5962_b0 );
or ( \11411_b1 , \11406_b1 , \11410_b1 );
xor ( \11411_b0 , \11406_b0 , w_29068 );
not ( w_29068 , w_29069 );
and ( w_29069 , \11410_b1 , \11410_b0 );
or ( \11412_b1 , \6041_b1 , \5977_b1 );
not ( \5977_b1 , w_29070 );
and ( \11412_b0 , \6041_b0 , w_29071 );
and ( w_29070 , w_29071 , \5977_b0 );
or ( \11413_b1 , \6006_b1 , \5975_b1 );
not ( \5975_b1 , w_29072 );
and ( \11413_b0 , \6006_b0 , w_29073 );
and ( w_29072 , w_29073 , \5975_b0 );
or ( \11414_b1 , \11412_b1 , w_29075 );
not ( w_29075 , w_29076 );
and ( \11414_b0 , \11412_b0 , w_29077 );
and ( w_29076 ,  , w_29077 );
buf ( w_29075 , \11413_b1 );
not ( w_29075 , w_29078 );
not (  , w_29079 );
and ( w_29078 , w_29079 , \11413_b0 );
or ( \11415_b1 , \11414_b1 , w_29080 );
xor ( \11415_b0 , \11414_b0 , w_29082 );
not ( w_29082 , w_29083 );
and ( w_29083 , w_29080 , w_29081 );
buf ( w_29080 , \5984_b1 );
not ( w_29080 , w_29084 );
not ( w_29081 , w_29085 );
and ( w_29084 , w_29085 , \5984_b0 );
or ( \11416_b1 , \11411_b1 , \11415_b1 );
xor ( \11416_b0 , \11411_b0 , w_29086 );
not ( w_29086 , w_29087 );
and ( w_29087 , \11415_b1 , \11415_b0 );
or ( \11417_b1 , \11402_b1 , \11416_b1 );
xor ( \11417_b0 , \11402_b0 , w_29088 );
not ( w_29088 , w_29089 );
and ( w_29089 , \11416_b1 , \11416_b0 );
or ( \11418_b1 , \5937_b1 , \5871_b1 );
not ( \5871_b1 , w_29090 );
and ( \11418_b0 , \5937_b0 , w_29091 );
and ( w_29090 , w_29091 , \5871_b0 );
or ( \11419_b1 , \5906_b1 , \5869_b1 );
not ( \5869_b1 , w_29092 );
and ( \11419_b0 , \5906_b0 , w_29093 );
and ( w_29092 , w_29093 , \5869_b0 );
or ( \11420_b1 , \11418_b1 , w_29095 );
not ( w_29095 , w_29096 );
and ( \11420_b0 , \11418_b0 , w_29097 );
and ( w_29096 ,  , w_29097 );
buf ( w_29095 , \11419_b1 );
not ( w_29095 , w_29098 );
not (  , w_29099 );
and ( w_29098 , w_29099 , \11419_b0 );
or ( \11421_b1 , \11420_b1 , w_29100 );
xor ( \11421_b0 , \11420_b0 , w_29102 );
not ( w_29102 , w_29103 );
and ( w_29103 , w_29100 , w_29101 );
buf ( w_29100 , \5878_b1 );
not ( w_29100 , w_29104 );
not ( w_29101 , w_29105 );
and ( w_29104 , w_29105 , \5878_b0 );
or ( \11422_b1 , \5957_b1 , \5891_b1 );
not ( \5891_b1 , w_29106 );
and ( \11422_b0 , \5957_b0 , w_29107 );
and ( w_29106 , w_29107 , \5891_b0 );
or ( \11423_b1 , \5925_b1 , \5889_b1 );
not ( \5889_b1 , w_29108 );
and ( \11423_b0 , \5925_b0 , w_29109 );
and ( w_29108 , w_29109 , \5889_b0 );
or ( \11424_b1 , \11422_b1 , w_29111 );
not ( w_29111 , w_29112 );
and ( \11424_b0 , \11422_b0 , w_29113 );
and ( w_29112 ,  , w_29113 );
buf ( w_29111 , \11423_b1 );
not ( w_29111 , w_29114 );
not (  , w_29115 );
and ( w_29114 , w_29115 , \11423_b0 );
or ( \11425_b1 , \11424_b1 , w_29116 );
xor ( \11425_b0 , \11424_b0 , w_29118 );
not ( w_29118 , w_29119 );
and ( w_29119 , w_29116 , w_29117 );
buf ( w_29116 , \5898_b1 );
not ( w_29116 , w_29120 );
not ( w_29117 , w_29121 );
and ( w_29120 , w_29121 , \5898_b0 );
or ( \11426_b1 , \11421_b1 , \11425_b1 );
xor ( \11426_b0 , \11421_b0 , w_29122 );
not ( w_29122 , w_29123 );
and ( w_29123 , \11425_b1 , \11425_b0 );
or ( \11427_b1 , \5979_b1 , \5916_b1 );
not ( \5916_b1 , w_29124 );
and ( \11427_b0 , \5979_b0 , w_29125 );
and ( w_29124 , w_29125 , \5916_b0 );
or ( \11428_b1 , \5945_b1 , \5914_b1 );
not ( \5914_b1 , w_29126 );
and ( \11428_b0 , \5945_b0 , w_29127 );
and ( w_29126 , w_29127 , \5914_b0 );
or ( \11429_b1 , \11427_b1 , w_29129 );
not ( w_29129 , w_29130 );
and ( \11429_b0 , \11427_b0 , w_29131 );
and ( w_29130 ,  , w_29131 );
buf ( w_29129 , \11428_b1 );
not ( w_29129 , w_29132 );
not (  , w_29133 );
and ( w_29132 , w_29133 , \11428_b0 );
or ( \11430_b1 , \11429_b1 , w_29134 );
xor ( \11430_b0 , \11429_b0 , w_29136 );
not ( w_29136 , w_29137 );
and ( w_29137 , w_29134 , w_29135 );
buf ( w_29134 , \5923_b1 );
not ( w_29134 , w_29138 );
not ( w_29135 , w_29139 );
and ( w_29138 , w_29139 , \5923_b0 );
or ( \11431_b1 , \11426_b1 , \11430_b1 );
xor ( \11431_b0 , \11426_b0 , w_29140 );
not ( w_29140 , w_29141 );
and ( w_29141 , \11430_b1 , \11430_b0 );
or ( \11432_b1 , \11417_b1 , \11431_b1 );
xor ( \11432_b0 , \11417_b0 , w_29142 );
not ( w_29142 , w_29143 );
and ( w_29143 , \11431_b1 , \11431_b0 );
or ( \11433_b1 , \11393_b1 , \11432_b1 );
xor ( \11433_b0 , \11393_b0 , w_29144 );
not ( w_29144 , w_29145 );
and ( w_29145 , \11432_b1 , \11432_b0 );
or ( \11434_b1 , \11347_b1 , \11433_b1 );
xor ( \11434_b0 , \11347_b0 , w_29146 );
not ( w_29146 , w_29147 );
and ( w_29147 , \11433_b1 , \11433_b0 );
or ( \11435_b1 , \11196_b1 , \11200_b1 );
not ( \11200_b1 , w_29148 );
and ( \11435_b0 , \11196_b0 , w_29149 );
and ( w_29148 , w_29149 , \11200_b0 );
or ( \11436_b1 , \11200_b1 , \11205_b1 );
not ( \11205_b1 , w_29150 );
and ( \11436_b0 , \11200_b0 , w_29151 );
and ( w_29150 , w_29151 , \11205_b0 );
or ( \11437_b1 , \11196_b1 , \11205_b1 );
not ( \11205_b1 , w_29152 );
and ( \11437_b0 , \11196_b0 , w_29153 );
and ( w_29152 , w_29153 , \11205_b0 );
or ( \11439_b1 , \11184_b1 , \11188_b1 );
not ( \11188_b1 , w_29154 );
and ( \11439_b0 , \11184_b0 , w_29155 );
and ( w_29154 , w_29155 , \11188_b0 );
or ( \11440_b1 , \11188_b1 , \11190_b1 );
not ( \11190_b1 , w_29156 );
and ( \11440_b0 , \11188_b0 , w_29157 );
and ( w_29156 , w_29157 , \11190_b0 );
or ( \11441_b1 , \11184_b1 , \11190_b1 );
not ( \11190_b1 , w_29158 );
and ( \11441_b0 , \11184_b0 , w_29159 );
and ( w_29158 , w_29159 , \11190_b0 );
or ( \11443_b1 , \11438_b1 , \11442_b1 );
xor ( \11443_b0 , \11438_b0 , w_29160 );
not ( w_29160 , w_29161 );
and ( w_29161 , \11442_b1 , \11442_b0 );
or ( \11444_b1 , \11165_b1 , w_29162 );
or ( \11444_b0 , \11165_b0 , \11179_b0 );
not ( \11179_b0 , w_29163 );
and ( w_29163 , w_29162 , \11179_b1 );
or ( \11445_b1 , \11443_b1 , \11444_b1 );
xor ( \11445_b0 , \11443_b0 , w_29164 );
not ( w_29164 , w_29165 );
and ( w_29165 , \11444_b1 , \11444_b0 );
or ( \11446_b1 , \11434_b1 , \11445_b1 );
xor ( \11446_b0 , \11434_b0 , w_29166 );
not ( w_29166 , w_29167 );
and ( w_29167 , \11445_b1 , \11445_b0 );
or ( \11447_b1 , \11318_b1 , \11446_b1 );
xor ( \11447_b0 , \11318_b0 , w_29168 );
not ( w_29168 , w_29169 );
and ( w_29169 , \11446_b1 , \11446_b0 );
or ( \11448_b1 , \11309_b1 , \11447_b1 );
xor ( \11448_b0 , \11309_b0 , w_29170 );
not ( w_29170 , w_29171 );
and ( w_29171 , \11447_b1 , \11447_b0 );
or ( \11449_b1 , \11132_b1 , \11143_b1 );
not ( \11143_b1 , w_29172 );
and ( \11449_b0 , \11132_b0 , w_29173 );
and ( w_29172 , w_29173 , \11143_b0 );
or ( \11450_b1 , \11143_b1 , \11283_b1 );
not ( \11283_b1 , w_29174 );
and ( \11450_b0 , \11143_b0 , w_29175 );
and ( w_29174 , w_29175 , \11283_b0 );
or ( \11451_b1 , \11132_b1 , \11283_b1 );
not ( \11283_b1 , w_29176 );
and ( \11451_b0 , \11132_b0 , w_29177 );
and ( w_29176 , w_29177 , \11283_b0 );
or ( \11453_b1 , \11448_b1 , w_29179 );
not ( w_29179 , w_29180 );
and ( \11453_b0 , \11448_b0 , w_29181 );
and ( w_29180 ,  , w_29181 );
buf ( w_29179 , \11452_b1 );
not ( w_29179 , w_29182 );
not (  , w_29183 );
and ( w_29182 , w_29183 , \11452_b0 );
or ( \11454_b1 , \11313_b1 , \11317_b1 );
not ( \11317_b1 , w_29184 );
and ( \11454_b0 , \11313_b0 , w_29185 );
and ( w_29184 , w_29185 , \11317_b0 );
or ( \11455_b1 , \11317_b1 , \11446_b1 );
not ( \11446_b1 , w_29186 );
and ( \11455_b0 , \11317_b0 , w_29187 );
and ( w_29186 , w_29187 , \11446_b0 );
or ( \11456_b1 , \11313_b1 , \11446_b1 );
not ( \11446_b1 , w_29188 );
and ( \11456_b0 , \11313_b0 , w_29189 );
and ( w_29188 , w_29189 , \11446_b0 );
or ( \11458_b1 , \11438_b1 , \11442_b1 );
not ( \11442_b1 , w_29190 );
and ( \11458_b0 , \11438_b0 , w_29191 );
and ( w_29190 , w_29191 , \11442_b0 );
or ( \11459_b1 , \11442_b1 , \11444_b1 );
not ( \11444_b1 , w_29192 );
and ( \11459_b0 , \11442_b0 , w_29193 );
and ( w_29192 , w_29193 , \11444_b0 );
or ( \11460_b1 , \11438_b1 , \11444_b1 );
not ( \11444_b1 , w_29194 );
and ( \11460_b0 , \11438_b0 , w_29195 );
and ( w_29194 , w_29195 , \11444_b0 );
or ( \11462_b1 , \11351_b1 , \11392_b1 );
not ( \11392_b1 , w_29196 );
and ( \11462_b0 , \11351_b0 , w_29197 );
and ( w_29196 , w_29197 , \11392_b0 );
or ( \11463_b1 , \11392_b1 , \11432_b1 );
not ( \11432_b1 , w_29198 );
and ( \11463_b0 , \11392_b0 , w_29199 );
and ( w_29198 , w_29199 , \11432_b0 );
or ( \11464_b1 , \11351_b1 , \11432_b1 );
not ( \11432_b1 , w_29200 );
and ( \11464_b0 , \11351_b0 , w_29201 );
and ( w_29200 , w_29201 , \11432_b0 );
or ( \11466_b1 , \11461_b1 , \11465_b1 );
xor ( \11466_b0 , \11461_b0 , w_29202 );
not ( w_29202 , w_29203 );
and ( w_29203 , \11465_b1 , \11465_b0 );
or ( \11467_b1 , \11332_b1 , \11346_b1 );
not ( \11346_b1 , w_29204 );
and ( \11467_b0 , \11332_b0 , w_29205 );
and ( w_29204 , w_29205 , \11346_b0 );
or ( \11468_b1 , \11466_b1 , \11467_b1 );
xor ( \11468_b0 , \11466_b0 , w_29206 );
not ( w_29206 , w_29207 );
and ( w_29207 , \11467_b1 , \11467_b0 );
or ( \11469_b1 , \11457_b1 , \11468_b1 );
xor ( \11469_b0 , \11457_b0 , w_29208 );
not ( w_29208 , w_29209 );
and ( w_29209 , \11468_b1 , \11468_b0 );
or ( \11470_b1 , \11298_b1 , \11302_b1 );
not ( \11302_b1 , w_29210 );
and ( \11470_b0 , \11298_b0 , w_29211 );
and ( w_29210 , w_29211 , \11302_b0 );
or ( \11471_b1 , \11302_b1 , \11307_b1 );
not ( \11307_b1 , w_29212 );
and ( \11471_b0 , \11302_b0 , w_29213 );
and ( w_29212 , w_29213 , \11307_b0 );
or ( \11472_b1 , \11298_b1 , \11307_b1 );
not ( \11307_b1 , w_29214 );
and ( \11472_b0 , \11298_b0 , w_29215 );
and ( w_29214 , w_29215 , \11307_b0 );
or ( \11474_b1 , \11347_b1 , \11433_b1 );
not ( \11433_b1 , w_29216 );
and ( \11474_b0 , \11347_b0 , w_29217 );
and ( w_29216 , w_29217 , \11433_b0 );
or ( \11475_b1 , \11433_b1 , \11445_b1 );
not ( \11445_b1 , w_29218 );
and ( \11475_b0 , \11433_b0 , w_29219 );
and ( w_29218 , w_29219 , \11445_b0 );
or ( \11476_b1 , \11347_b1 , \11445_b1 );
not ( \11445_b1 , w_29220 );
and ( \11476_b0 , \11347_b0 , w_29221 );
and ( w_29220 , w_29221 , \11445_b0 );
or ( \11478_b1 , \11473_b1 , \11477_b1 );
xor ( \11478_b0 , \11473_b0 , w_29222 );
not ( w_29222 , w_29223 );
and ( w_29223 , \11477_b1 , \11477_b0 );
or ( \11479_b1 , \6029_b1 , \5996_b1 );
not ( \5996_b1 , w_29224 );
and ( \11479_b0 , \6029_b0 , w_29225 );
and ( w_29224 , w_29225 , \5996_b0 );
or ( \11480_b1 , \6041_b1 , \5994_b1 );
not ( \5994_b1 , w_29226 );
and ( \11480_b0 , \6041_b0 , w_29227 );
and ( w_29226 , w_29227 , \5994_b0 );
or ( \11481_b1 , \11479_b1 , w_29229 );
not ( w_29229 , w_29230 );
and ( \11481_b0 , \11479_b0 , w_29231 );
and ( w_29230 ,  , w_29231 );
buf ( w_29229 , \11480_b1 );
not ( w_29229 , w_29232 );
not (  , w_29233 );
and ( w_29232 , w_29233 , \11480_b0 );
or ( \11482_b1 , \11481_b1 , w_29234 );
xor ( \11482_b0 , \11481_b0 , w_29236 );
not ( w_29236 , w_29237 );
and ( w_29237 , w_29234 , w_29235 );
buf ( w_29234 , \6003_b1 );
not ( w_29234 , w_29238 );
not ( w_29235 , w_29239 );
and ( w_29238 , w_29239 , \6003_b0 );
or ( \11483_b1 , \6048_b1 , \6016_b1 );
not ( \6016_b1 , w_29240 );
and ( \11483_b0 , \6048_b0 , w_29241 );
and ( w_29240 , w_29241 , \6016_b0 );
or ( \11484_b1 , \6057_b1 , \6014_b1 );
not ( \6014_b1 , w_29242 );
and ( \11484_b0 , \6057_b0 , w_29243 );
and ( w_29242 , w_29243 , \6014_b0 );
or ( \11485_b1 , \11483_b1 , w_29245 );
not ( w_29245 , w_29246 );
and ( \11485_b0 , \11483_b0 , w_29247 );
and ( w_29246 ,  , w_29247 );
buf ( w_29245 , \11484_b1 );
not ( w_29245 , w_29248 );
not (  , w_29249 );
and ( w_29248 , w_29249 , \11484_b0 );
or ( \11486_b1 , \11485_b1 , w_29250 );
xor ( \11486_b0 , \11485_b0 , w_29252 );
not ( w_29252 , w_29253 );
and ( w_29253 , w_29250 , w_29251 );
buf ( w_29250 , \6023_b1 );
not ( w_29250 , w_29254 );
not ( w_29251 , w_29255 );
and ( w_29254 , w_29255 , \6023_b0 );
or ( \11487_b1 , \11482_b1 , \11486_b1 );
xor ( \11487_b0 , \11482_b0 , w_29256 );
not ( w_29256 , w_29257 );
and ( w_29257 , \11486_b1 , \11486_b0 );
or ( \11488_b1 , \6065_b1 , w_29259 );
not ( w_29259 , w_29260 );
and ( \11488_b0 , \6065_b0 , w_29261 );
and ( w_29260 ,  , w_29261 );
buf ( w_29259 , \6037_b1 );
not ( w_29259 , w_29262 );
not (  , w_29263 );
and ( w_29262 , w_29263 , \6037_b0 );
or ( \11489_b1 , \11488_b1 , w_29264 );
xor ( \11489_b0 , \11488_b0 , w_29266 );
not ( w_29266 , w_29267 );
and ( w_29267 , w_29264 , w_29265 );
buf ( w_29264 , \6046_b1 );
not ( w_29264 , w_29268 );
not ( w_29265 , w_29269 );
and ( w_29268 , w_29269 , \6046_b0 );
or ( \11490_b1 , \11487_b1 , \11489_b1 );
xor ( \11490_b0 , \11487_b0 , w_29270 );
not ( w_29270 , w_29271 );
and ( w_29271 , \11489_b1 , \11489_b0 );
or ( \11491_b1 , \5967_b1 , \5935_b1 );
not ( \5935_b1 , w_29272 );
and ( \11491_b0 , \5967_b0 , w_29273 );
and ( w_29272 , w_29273 , \5935_b0 );
or ( \11492_b1 , \5979_b1 , \5933_b1 );
not ( \5933_b1 , w_29274 );
and ( \11492_b0 , \5979_b0 , w_29275 );
and ( w_29274 , w_29275 , \5933_b0 );
or ( \11493_b1 , \11491_b1 , w_29277 );
not ( w_29277 , w_29278 );
and ( \11493_b0 , \11491_b0 , w_29279 );
and ( w_29278 ,  , w_29279 );
buf ( w_29277 , \11492_b1 );
not ( w_29277 , w_29280 );
not (  , w_29281 );
and ( w_29280 , w_29281 , \11492_b0 );
or ( \11494_b1 , \11493_b1 , w_29282 );
xor ( \11494_b0 , \11493_b0 , w_29284 );
not ( w_29284 , w_29285 );
and ( w_29285 , w_29282 , w_29283 );
buf ( w_29282 , \5942_b1 );
not ( w_29282 , w_29286 );
not ( w_29283 , w_29287 );
and ( w_29286 , w_29287 , \5942_b0 );
or ( \11495_b1 , \5986_b1 , \5955_b1 );
not ( \5955_b1 , w_29288 );
and ( \11495_b0 , \5986_b0 , w_29289 );
and ( w_29288 , w_29289 , \5955_b0 );
or ( \11496_b1 , \5998_b1 , \5953_b1 );
not ( \5953_b1 , w_29290 );
and ( \11496_b0 , \5998_b0 , w_29291 );
and ( w_29290 , w_29291 , \5953_b0 );
or ( \11497_b1 , \11495_b1 , w_29293 );
not ( w_29293 , w_29294 );
and ( \11497_b0 , \11495_b0 , w_29295 );
and ( w_29294 ,  , w_29295 );
buf ( w_29293 , \11496_b1 );
not ( w_29293 , w_29296 );
not (  , w_29297 );
and ( w_29296 , w_29297 , \11496_b0 );
or ( \11498_b1 , \11497_b1 , w_29298 );
xor ( \11498_b0 , \11497_b0 , w_29300 );
not ( w_29300 , w_29301 );
and ( w_29301 , w_29298 , w_29299 );
buf ( w_29298 , \5962_b1 );
not ( w_29298 , w_29302 );
not ( w_29299 , w_29303 );
and ( w_29302 , w_29303 , \5962_b0 );
or ( \11499_b1 , \11494_b1 , \11498_b1 );
xor ( \11499_b0 , \11494_b0 , w_29304 );
not ( w_29304 , w_29305 );
and ( w_29305 , \11498_b1 , \11498_b0 );
or ( \11500_b1 , \6006_b1 , \5977_b1 );
not ( \5977_b1 , w_29306 );
and ( \11500_b0 , \6006_b0 , w_29307 );
and ( w_29306 , w_29307 , \5977_b0 );
or ( \11501_b1 , \6018_b1 , \5975_b1 );
not ( \5975_b1 , w_29308 );
and ( \11501_b0 , \6018_b0 , w_29309 );
and ( w_29308 , w_29309 , \5975_b0 );
or ( \11502_b1 , \11500_b1 , w_29311 );
not ( w_29311 , w_29312 );
and ( \11502_b0 , \11500_b0 , w_29313 );
and ( w_29312 ,  , w_29313 );
buf ( w_29311 , \11501_b1 );
not ( w_29311 , w_29314 );
not (  , w_29315 );
and ( w_29314 , w_29315 , \11501_b0 );
or ( \11503_b1 , \11502_b1 , w_29316 );
xor ( \11503_b0 , \11502_b0 , w_29318 );
not ( w_29318 , w_29319 );
and ( w_29319 , w_29316 , w_29317 );
buf ( w_29316 , \5984_b1 );
not ( w_29316 , w_29320 );
not ( w_29317 , w_29321 );
and ( w_29320 , w_29321 , \5984_b0 );
or ( \11504_b1 , \11499_b1 , \11503_b1 );
xor ( \11504_b0 , \11499_b0 , w_29322 );
not ( w_29322 , w_29323 );
and ( w_29323 , \11503_b1 , \11503_b0 );
or ( \11505_b1 , \11490_b1 , w_29324 );
xor ( \11505_b0 , \11490_b0 , w_29326 );
not ( w_29326 , w_29327 );
and ( w_29327 , w_29324 , w_29325 );
buf ( w_29324 , \11504_b1 );
not ( w_29324 , w_29328 );
not ( w_29325 , w_29329 );
and ( w_29328 , w_29329 , \11504_b0 );
or ( \11506_b1 , \11421_b1 , \11425_b1 );
not ( \11425_b1 , w_29330 );
and ( \11506_b0 , \11421_b0 , w_29331 );
and ( w_29330 , w_29331 , \11425_b0 );
or ( \11507_b1 , \11425_b1 , \11430_b1 );
not ( \11430_b1 , w_29332 );
and ( \11507_b0 , \11425_b0 , w_29333 );
and ( w_29332 , w_29333 , \11430_b0 );
or ( \11508_b1 , \11421_b1 , \11430_b1 );
not ( \11430_b1 , w_29334 );
and ( \11508_b0 , \11421_b0 , w_29335 );
and ( w_29334 , w_29335 , \11430_b0 );
or ( \11510_b1 , \11406_b1 , \11410_b1 );
not ( \11410_b1 , w_29336 );
and ( \11510_b0 , \11406_b0 , w_29337 );
and ( w_29336 , w_29337 , \11410_b0 );
or ( \11511_b1 , \11410_b1 , \11415_b1 );
not ( \11415_b1 , w_29338 );
and ( \11511_b0 , \11410_b0 , w_29339 );
and ( w_29338 , w_29339 , \11415_b0 );
or ( \11512_b1 , \11406_b1 , \11415_b1 );
not ( \11415_b1 , w_29340 );
and ( \11512_b0 , \11406_b0 , w_29341 );
and ( w_29340 , w_29341 , \11415_b0 );
or ( \11514_b1 , \11509_b1 , \11513_b1 );
xor ( \11514_b0 , \11509_b0 , w_29342 );
not ( w_29342 , w_29343 );
and ( w_29343 , \11513_b1 , \11513_b0 );
or ( \11515_b1 , \11397_b1 , \11401_b1 );
not ( \11401_b1 , w_29344 );
and ( \11515_b0 , \11397_b0 , w_29345 );
and ( w_29344 , w_29345 , \11401_b0 );
or ( \11516_b1 , \11514_b1 , \11515_b1 );
xor ( \11516_b0 , \11514_b0 , w_29346 );
not ( w_29346 , w_29347 );
and ( w_29347 , \11515_b1 , \11515_b0 );
or ( \11517_b1 , \11505_b1 , \11516_b1 );
xor ( \11517_b0 , \11505_b0 , w_29348 );
not ( w_29348 , w_29349 );
and ( w_29349 , \11516_b1 , \11516_b0 );
or ( \11518_b1 , \11381_b1 , \11385_b1 );
not ( \11385_b1 , w_29350 );
and ( \11518_b0 , \11381_b0 , w_29351 );
and ( w_29350 , w_29351 , \11385_b0 );
or ( \11519_b1 , \11385_b1 , \11390_b1 );
not ( \11390_b1 , w_29352 );
and ( \11519_b0 , \11385_b0 , w_29353 );
and ( w_29352 , w_29353 , \11390_b0 );
or ( \11520_b1 , \11381_b1 , \11390_b1 );
not ( \11390_b1 , w_29354 );
and ( \11520_b0 , \11381_b0 , w_29355 );
and ( w_29354 , w_29355 , \11390_b0 );
or ( \11522_b1 , \11369_b1 , \11373_b1 );
not ( \11373_b1 , w_29356 );
and ( \11522_b0 , \11369_b0 , w_29357 );
and ( w_29356 , w_29357 , \11373_b0 );
or ( \11523_b1 , \11373_b1 , \11378_b1 );
not ( \11378_b1 , w_29358 );
and ( \11523_b0 , \11373_b0 , w_29359 );
and ( w_29358 , w_29359 , \11378_b0 );
or ( \11524_b1 , \11369_b1 , \11378_b1 );
not ( \11378_b1 , w_29360 );
and ( \11524_b0 , \11369_b0 , w_29361 );
and ( w_29360 , w_29361 , \11378_b0 );
or ( \11526_b1 , \11521_b1 , \11525_b1 );
xor ( \11526_b0 , \11521_b0 , w_29362 );
not ( w_29362 , w_29363 );
and ( w_29363 , \11525_b1 , \11525_b0 );
or ( \11527_b1 , \11355_b1 , \11359_b1 );
not ( \11359_b1 , w_29364 );
and ( \11527_b0 , \11355_b0 , w_29365 );
and ( w_29364 , w_29365 , \11359_b0 );
or ( \11528_b1 , \11359_b1 , \11364_b1 );
not ( \11364_b1 , w_29366 );
and ( \11528_b0 , \11359_b0 , w_29367 );
and ( w_29366 , w_29367 , \11364_b0 );
or ( \11529_b1 , \11355_b1 , \11364_b1 );
not ( \11364_b1 , w_29368 );
and ( \11529_b0 , \11355_b0 , w_29369 );
and ( w_29368 , w_29369 , \11364_b0 );
or ( \11531_b1 , \11526_b1 , \11530_b1 );
xor ( \11531_b0 , \11526_b0 , w_29370 );
not ( w_29370 , w_29371 );
and ( w_29371 , \11530_b1 , \11530_b0 );
or ( \11532_b1 , \11517_b1 , \11531_b1 );
xor ( \11532_b0 , \11517_b0 , w_29372 );
not ( w_29372 , w_29373 );
and ( w_29373 , \11531_b1 , \11531_b0 );
or ( \11533_b1 , \11365_b1 , \11379_b1 );
not ( \11379_b1 , w_29374 );
and ( \11533_b0 , \11365_b0 , w_29375 );
and ( w_29374 , w_29375 , \11379_b0 );
or ( \11534_b1 , \11379_b1 , \11391_b1 );
not ( \11391_b1 , w_29376 );
and ( \11534_b0 , \11379_b0 , w_29377 );
and ( w_29376 , w_29377 , \11391_b0 );
or ( \11535_b1 , \11365_b1 , \11391_b1 );
not ( \11391_b1 , w_29378 );
and ( \11535_b0 , \11365_b0 , w_29379 );
and ( w_29378 , w_29379 , \11391_b0 );
or ( \11537_b1 , \5737_b1 , \7192_b1 );
not ( \7192_b1 , w_29380 );
and ( \11537_b0 , \5737_b0 , w_29381 );
and ( w_29380 , w_29381 , \7192_b0 );
buf ( \11538_b1 , \11537_b1 );
not ( \11538_b1 , w_29382 );
not ( \11538_b0 , w_29383 );
and ( w_29382 , w_29383 , \11537_b0 );
or ( \11539_b1 , \11538_b1 , w_29384 );
xor ( \11539_b0 , \11538_b0 , w_29386 );
not ( w_29386 , w_29387 );
and ( w_29387 , w_29384 , w_29385 );
buf ( w_29384 , \7198_b1 );
not ( w_29384 , w_29388 );
not ( w_29385 , w_29389 );
and ( w_29388 , w_29389 , \7198_b0 );
or ( \11540_b1 , \6046_b1 , \11539_b1 );
xor ( \11540_b0 , \6046_b0 , w_29390 );
not ( w_29390 , w_29391 );
and ( w_29391 , \11539_b1 , \11539_b0 );
or ( \11541_b1 , \5758_b1 , \7203_b1 );
not ( \7203_b1 , w_29392 );
and ( \11541_b0 , \5758_b0 , w_29393 );
and ( w_29392 , w_29393 , \7203_b0 );
or ( \11542_b1 , \5770_b1 , \7201_b1 );
not ( \7201_b1 , w_29394 );
and ( \11542_b0 , \5770_b0 , w_29395 );
and ( w_29394 , w_29395 , \7201_b0 );
or ( \11543_b1 , \11541_b1 , w_29397 );
not ( w_29397 , w_29398 );
and ( \11543_b0 , \11541_b0 , w_29399 );
and ( w_29398 ,  , w_29399 );
buf ( w_29397 , \11542_b1 );
not ( w_29397 , w_29400 );
not (  , w_29401 );
and ( w_29400 , w_29401 , \11542_b0 );
or ( \11544_b1 , \11543_b1 , w_29402 );
xor ( \11544_b0 , \11543_b0 , w_29404 );
not ( w_29404 , w_29405 );
and ( w_29405 , w_29402 , w_29403 );
buf ( w_29402 , \6824_b1 );
not ( w_29402 , w_29406 );
not ( w_29403 , w_29407 );
and ( w_29406 , w_29407 , \6824_b0 );
or ( \11545_b1 , \11540_b1 , \11544_b1 );
xor ( \11545_b0 , \11540_b0 , w_29408 );
not ( w_29408 , w_29409 );
and ( w_29409 , \11544_b1 , \11544_b0 );
or ( \11546_b1 , \11536_b1 , \11545_b1 );
xor ( \11546_b0 , \11536_b0 , w_29410 );
not ( w_29410 , w_29411 );
and ( w_29411 , \11545_b1 , \11545_b0 );
or ( \11547_b1 , \5906_b1 , \5871_b1 );
not ( \5871_b1 , w_29412 );
and ( \11547_b0 , \5906_b0 , w_29413 );
and ( w_29412 , w_29413 , \5871_b0 );
or ( \11548_b1 , \5918_b1 , \5869_b1 );
not ( \5869_b1 , w_29414 );
and ( \11548_b0 , \5918_b0 , w_29415 );
and ( w_29414 , w_29415 , \5869_b0 );
or ( \11549_b1 , \11547_b1 , w_29417 );
not ( w_29417 , w_29418 );
and ( \11549_b0 , \11547_b0 , w_29419 );
and ( w_29418 ,  , w_29419 );
buf ( w_29417 , \11548_b1 );
not ( w_29417 , w_29420 );
not (  , w_29421 );
and ( w_29420 , w_29421 , \11548_b0 );
or ( \11550_b1 , \11549_b1 , w_29422 );
xor ( \11550_b0 , \11549_b0 , w_29424 );
not ( w_29424 , w_29425 );
and ( w_29425 , w_29422 , w_29423 );
buf ( w_29422 , \5878_b1 );
not ( w_29422 , w_29426 );
not ( w_29423 , w_29427 );
and ( w_29426 , w_29427 , \5878_b0 );
or ( \11551_b1 , \5925_b1 , \5891_b1 );
not ( \5891_b1 , w_29428 );
and ( \11551_b0 , \5925_b0 , w_29429 );
and ( w_29428 , w_29429 , \5891_b0 );
or ( \11552_b1 , \5937_b1 , \5889_b1 );
not ( \5889_b1 , w_29430 );
and ( \11552_b0 , \5937_b0 , w_29431 );
and ( w_29430 , w_29431 , \5889_b0 );
or ( \11553_b1 , \11551_b1 , w_29433 );
not ( w_29433 , w_29434 );
and ( \11553_b0 , \11551_b0 , w_29435 );
and ( w_29434 ,  , w_29435 );
buf ( w_29433 , \11552_b1 );
not ( w_29433 , w_29436 );
not (  , w_29437 );
and ( w_29436 , w_29437 , \11552_b0 );
or ( \11554_b1 , \11553_b1 , w_29438 );
xor ( \11554_b0 , \11553_b0 , w_29440 );
not ( w_29440 , w_29441 );
and ( w_29441 , w_29438 , w_29439 );
buf ( w_29438 , \5898_b1 );
not ( w_29438 , w_29442 );
not ( w_29439 , w_29443 );
and ( w_29442 , w_29443 , \5898_b0 );
or ( \11555_b1 , \11550_b1 , \11554_b1 );
xor ( \11555_b0 , \11550_b0 , w_29444 );
not ( w_29444 , w_29445 );
and ( w_29445 , \11554_b1 , \11554_b0 );
or ( \11556_b1 , \5945_b1 , \5916_b1 );
not ( \5916_b1 , w_29446 );
and ( \11556_b0 , \5945_b0 , w_29447 );
and ( w_29446 , w_29447 , \5916_b0 );
or ( \11557_b1 , \5957_b1 , \5914_b1 );
not ( \5914_b1 , w_29448 );
and ( \11557_b0 , \5957_b0 , w_29449 );
and ( w_29448 , w_29449 , \5914_b0 );
or ( \11558_b1 , \11556_b1 , w_29451 );
not ( w_29451 , w_29452 );
and ( \11558_b0 , \11556_b0 , w_29453 );
and ( w_29452 ,  , w_29453 );
buf ( w_29451 , \11557_b1 );
not ( w_29451 , w_29454 );
not (  , w_29455 );
and ( w_29454 , w_29455 , \11557_b0 );
or ( \11559_b1 , \11558_b1 , w_29456 );
xor ( \11559_b0 , \11558_b0 , w_29458 );
not ( w_29458 , w_29459 );
and ( w_29459 , w_29456 , w_29457 );
buf ( w_29456 , \5923_b1 );
not ( w_29456 , w_29460 );
not ( w_29457 , w_29461 );
and ( w_29460 , w_29461 , \5923_b0 );
or ( \11560_b1 , \11555_b1 , \11559_b1 );
xor ( \11560_b0 , \11555_b0 , w_29462 );
not ( w_29462 , w_29463 );
and ( w_29463 , \11559_b1 , \11559_b0 );
or ( \11561_b1 , \5842_b1 , \5809_b1 );
not ( \5809_b1 , w_29464 );
and ( \11561_b0 , \5842_b0 , w_29465 );
and ( w_29464 , w_29465 , \5809_b0 );
or ( \11562_b1 , \5854_b1 , \5807_b1 );
not ( \5807_b1 , w_29466 );
and ( \11562_b0 , \5854_b0 , w_29467 );
and ( w_29466 , w_29467 , \5807_b0 );
or ( \11563_b1 , \11561_b1 , w_29469 );
not ( w_29469 , w_29470 );
and ( \11563_b0 , \11561_b0 , w_29471 );
and ( w_29470 ,  , w_29471 );
buf ( w_29469 , \11562_b1 );
not ( w_29469 , w_29472 );
not (  , w_29473 );
and ( w_29472 , w_29473 , \11562_b0 );
or ( \11564_b1 , \11563_b1 , w_29474 );
xor ( \11564_b0 , \11563_b0 , w_29476 );
not ( w_29476 , w_29477 );
and ( w_29477 , w_29474 , w_29475 );
buf ( w_29474 , \5816_b1 );
not ( w_29474 , w_29478 );
not ( w_29475 , w_29479 );
and ( w_29478 , w_29479 , \5816_b0 );
or ( \11565_b1 , \5861_b1 , \5829_b1 );
not ( \5829_b1 , w_29480 );
and ( \11565_b0 , \5861_b0 , w_29481 );
and ( w_29480 , w_29481 , \5829_b0 );
or ( \11566_b1 , \5873_b1 , \5827_b1 );
not ( \5827_b1 , w_29482 );
and ( \11566_b0 , \5873_b0 , w_29483 );
and ( w_29482 , w_29483 , \5827_b0 );
or ( \11567_b1 , \11565_b1 , w_29485 );
not ( w_29485 , w_29486 );
and ( \11567_b0 , \11565_b0 , w_29487 );
and ( w_29486 ,  , w_29487 );
buf ( w_29485 , \11566_b1 );
not ( w_29485 , w_29488 );
not (  , w_29489 );
and ( w_29488 , w_29489 , \11566_b0 );
or ( \11568_b1 , \11567_b1 , w_29490 );
xor ( \11568_b0 , \11567_b0 , w_29492 );
not ( w_29492 , w_29493 );
and ( w_29493 , w_29490 , w_29491 );
buf ( w_29490 , \5836_b1 );
not ( w_29490 , w_29494 );
not ( w_29491 , w_29495 );
and ( w_29494 , w_29495 , \5836_b0 );
or ( \11569_b1 , \11564_b1 , \11568_b1 );
xor ( \11569_b0 , \11564_b0 , w_29496 );
not ( w_29496 , w_29497 );
and ( w_29497 , \11568_b1 , \11568_b0 );
or ( \11570_b1 , \5881_b1 , \5852_b1 );
not ( \5852_b1 , w_29498 );
and ( \11570_b0 , \5881_b0 , w_29499 );
and ( w_29498 , w_29499 , \5852_b0 );
or ( \11571_b1 , \5893_b1 , \5850_b1 );
not ( \5850_b1 , w_29500 );
and ( \11571_b0 , \5893_b0 , w_29501 );
and ( w_29500 , w_29501 , \5850_b0 );
or ( \11572_b1 , \11570_b1 , w_29503 );
not ( w_29503 , w_29504 );
and ( \11572_b0 , \11570_b0 , w_29505 );
and ( w_29504 ,  , w_29505 );
buf ( w_29503 , \11571_b1 );
not ( w_29503 , w_29506 );
not (  , w_29507 );
and ( w_29506 , w_29507 , \11571_b0 );
or ( \11573_b1 , \11572_b1 , w_29508 );
xor ( \11573_b0 , \11572_b0 , w_29510 );
not ( w_29510 , w_29511 );
and ( w_29511 , w_29508 , w_29509 );
buf ( w_29508 , \5859_b1 );
not ( w_29508 , w_29512 );
not ( w_29509 , w_29513 );
and ( w_29512 , w_29513 , \5859_b0 );
or ( \11574_b1 , \11569_b1 , \11573_b1 );
xor ( \11574_b0 , \11569_b0 , w_29514 );
not ( w_29514 , w_29515 );
and ( w_29515 , \11573_b1 , \11573_b0 );
or ( \11575_b1 , \11560_b1 , \11574_b1 );
xor ( \11575_b0 , \11560_b0 , w_29516 );
not ( w_29516 , w_29517 );
and ( w_29517 , \11574_b1 , \11574_b0 );
or ( \11576_b1 , \5780_b1 , \5750_b1 );
not ( \5750_b1 , w_29518 );
and ( \11576_b0 , \5780_b0 , w_29519 );
and ( w_29518 , w_29519 , \5750_b0 );
or ( \11577_b1 , \5792_b1 , \5748_b1 );
not ( \5748_b1 , w_29520 );
and ( \11577_b0 , \5792_b0 , w_29521 );
and ( w_29520 , w_29521 , \5748_b0 );
or ( \11578_b1 , \11576_b1 , w_29523 );
not ( w_29523 , w_29524 );
and ( \11578_b0 , \11576_b0 , w_29525 );
and ( w_29524 ,  , w_29525 );
buf ( w_29523 , \11577_b1 );
not ( w_29523 , w_29526 );
not (  , w_29527 );
and ( w_29526 , w_29527 , \11577_b0 );
or ( \11579_b1 , \11578_b1 , w_29528 );
xor ( \11579_b0 , \11578_b0 , w_29530 );
not ( w_29530 , w_29531 );
and ( w_29531 , w_29528 , w_29529 );
buf ( w_29528 , \5755_b1 );
not ( w_29528 , w_29532 );
not ( w_29529 , w_29533 );
and ( w_29532 , w_29533 , \5755_b0 );
or ( \11580_b1 , \5799_b1 , \5768_b1 );
not ( \5768_b1 , w_29534 );
and ( \11580_b0 , \5799_b0 , w_29535 );
and ( w_29534 , w_29535 , \5768_b0 );
or ( \11581_b1 , \5811_b1 , \5766_b1 );
not ( \5766_b1 , w_29536 );
and ( \11581_b0 , \5811_b0 , w_29537 );
and ( w_29536 , w_29537 , \5766_b0 );
or ( \11582_b1 , \11580_b1 , w_29539 );
not ( w_29539 , w_29540 );
and ( \11582_b0 , \11580_b0 , w_29541 );
and ( w_29540 ,  , w_29541 );
buf ( w_29539 , \11581_b1 );
not ( w_29539 , w_29542 );
not (  , w_29543 );
and ( w_29542 , w_29543 , \11581_b0 );
or ( \11583_b1 , \11582_b1 , w_29544 );
xor ( \11583_b0 , \11582_b0 , w_29546 );
not ( w_29546 , w_29547 );
and ( w_29547 , w_29544 , w_29545 );
buf ( w_29544 , \5775_b1 );
not ( w_29544 , w_29548 );
not ( w_29545 , w_29549 );
and ( w_29548 , w_29549 , \5775_b0 );
or ( \11584_b1 , \11579_b1 , \11583_b1 );
xor ( \11584_b0 , \11579_b0 , w_29550 );
not ( w_29550 , w_29551 );
and ( w_29551 , \11583_b1 , \11583_b0 );
or ( \11585_b1 , \5819_b1 , \5790_b1 );
not ( \5790_b1 , w_29552 );
and ( \11585_b0 , \5819_b0 , w_29553 );
and ( w_29552 , w_29553 , \5790_b0 );
or ( \11586_b1 , \5831_b1 , \5788_b1 );
not ( \5788_b1 , w_29554 );
and ( \11586_b0 , \5831_b0 , w_29555 );
and ( w_29554 , w_29555 , \5788_b0 );
or ( \11587_b1 , \11585_b1 , w_29557 );
not ( w_29557 , w_29558 );
and ( \11587_b0 , \11585_b0 , w_29559 );
and ( w_29558 ,  , w_29559 );
buf ( w_29557 , \11586_b1 );
not ( w_29557 , w_29560 );
not (  , w_29561 );
and ( w_29560 , w_29561 , \11586_b0 );
or ( \11588_b1 , \11587_b1 , w_29562 );
xor ( \11588_b0 , \11587_b0 , w_29564 );
not ( w_29564 , w_29565 );
and ( w_29565 , w_29562 , w_29563 );
buf ( w_29562 , \5797_b1 );
not ( w_29562 , w_29566 );
not ( w_29563 , w_29567 );
and ( w_29566 , w_29567 , \5797_b0 );
or ( \11589_b1 , \11584_b1 , \11588_b1 );
xor ( \11589_b0 , \11584_b0 , w_29568 );
not ( w_29568 , w_29569 );
and ( w_29569 , \11588_b1 , \11588_b0 );
or ( \11590_b1 , \11575_b1 , \11589_b1 );
xor ( \11590_b0 , \11575_b0 , w_29570 );
not ( w_29570 , w_29571 );
and ( w_29571 , \11589_b1 , \11589_b0 );
or ( \11591_b1 , \11546_b1 , \11590_b1 );
xor ( \11591_b0 , \11546_b0 , w_29572 );
not ( w_29572 , w_29573 );
and ( w_29573 , \11590_b1 , \11590_b0 );
or ( \11592_b1 , \11532_b1 , \11591_b1 );
xor ( \11592_b0 , \11532_b0 , w_29574 );
not ( w_29574 , w_29575 );
and ( w_29575 , \11591_b1 , \11591_b0 );
or ( \11593_b1 , \11336_b1 , \11340_b1 );
not ( \11340_b1 , w_29576 );
and ( \11593_b0 , \11336_b0 , w_29577 );
and ( w_29576 , w_29577 , \11340_b0 );
or ( \11594_b1 , \11340_b1 , \11345_b1 );
not ( \11345_b1 , w_29578 );
and ( \11594_b0 , \11340_b0 , w_29579 );
and ( w_29578 , w_29579 , \11345_b0 );
or ( \11595_b1 , \11336_b1 , \11345_b1 );
not ( \11345_b1 , w_29580 );
and ( \11595_b0 , \11336_b0 , w_29581 );
and ( w_29580 , w_29581 , \11345_b0 );
or ( \11597_b1 , \11322_b1 , \11326_b1 );
not ( \11326_b1 , w_29582 );
and ( \11597_b0 , \11322_b0 , w_29583 );
and ( w_29582 , w_29583 , \11326_b0 );
or ( \11598_b1 , \11326_b1 , \11331_b1 );
not ( \11331_b1 , w_29584 );
and ( \11598_b0 , \11326_b0 , w_29585 );
and ( w_29584 , w_29585 , \11331_b0 );
or ( \11599_b1 , \11322_b1 , \11331_b1 );
not ( \11331_b1 , w_29586 );
and ( \11599_b0 , \11322_b0 , w_29587 );
and ( w_29586 , w_29587 , \11331_b0 );
or ( \11601_b1 , \11596_b1 , \11600_b1 );
xor ( \11601_b0 , \11596_b0 , w_29588 );
not ( w_29588 , w_29589 );
and ( w_29589 , \11600_b1 , \11600_b0 );
or ( \11602_b1 , \11402_b1 , \11416_b1 );
not ( \11416_b1 , w_29590 );
and ( \11602_b0 , \11402_b0 , w_29591 );
and ( w_29590 , w_29591 , \11416_b0 );
or ( \11603_b1 , \11416_b1 , \11431_b1 );
not ( \11431_b1 , w_29592 );
and ( \11603_b0 , \11416_b0 , w_29593 );
and ( w_29592 , w_29593 , \11431_b0 );
or ( \11604_b1 , \11402_b1 , \11431_b1 );
not ( \11431_b1 , w_29594 );
and ( \11604_b0 , \11402_b0 , w_29595 );
and ( w_29594 , w_29595 , \11431_b0 );
or ( \11606_b1 , \11601_b1 , \11605_b1 );
xor ( \11606_b0 , \11601_b0 , w_29596 );
not ( w_29596 , w_29597 );
and ( w_29597 , \11605_b1 , \11605_b0 );
or ( \11607_b1 , \11592_b1 , \11606_b1 );
xor ( \11607_b0 , \11592_b0 , w_29598 );
not ( w_29598 , w_29599 );
and ( w_29599 , \11606_b1 , \11606_b0 );
or ( \11608_b1 , \11478_b1 , \11607_b1 );
xor ( \11608_b0 , \11478_b0 , w_29600 );
not ( w_29600 , w_29601 );
and ( w_29601 , \11607_b1 , \11607_b0 );
or ( \11609_b1 , \11469_b1 , \11608_b1 );
xor ( \11609_b0 , \11469_b0 , w_29602 );
not ( w_29602 , w_29603 );
and ( w_29603 , \11608_b1 , \11608_b0 );
or ( \11610_b1 , \11294_b1 , \11308_b1 );
not ( \11308_b1 , w_29604 );
and ( \11610_b0 , \11294_b0 , w_29605 );
and ( w_29604 , w_29605 , \11308_b0 );
or ( \11611_b1 , \11308_b1 , \11447_b1 );
not ( \11447_b1 , w_29606 );
and ( \11611_b0 , \11308_b0 , w_29607 );
and ( w_29606 , w_29607 , \11447_b0 );
or ( \11612_b1 , \11294_b1 , \11447_b1 );
not ( \11447_b1 , w_29608 );
and ( \11612_b0 , \11294_b0 , w_29609 );
and ( w_29608 , w_29609 , \11447_b0 );
or ( \11614_b1 , \11609_b1 , w_29611 );
not ( w_29611 , w_29612 );
and ( \11614_b0 , \11609_b0 , w_29613 );
and ( w_29612 ,  , w_29613 );
buf ( w_29611 , \11613_b1 );
not ( w_29611 , w_29614 );
not (  , w_29615 );
and ( w_29614 , w_29615 , \11613_b0 );
or ( \11615_b1 , \11453_b1 , w_29617 );
not ( w_29617 , w_29618 );
and ( \11615_b0 , \11453_b0 , w_29619 );
and ( w_29618 ,  , w_29619 );
buf ( w_29617 , \11614_b1 );
not ( w_29617 , w_29620 );
not (  , w_29621 );
and ( w_29620 , w_29621 , \11614_b0 );
or ( \11616_b1 , \11290_b1 , w_29623 );
not ( w_29623 , w_29624 );
and ( \11616_b0 , \11290_b0 , w_29625 );
and ( w_29624 ,  , w_29625 );
buf ( w_29623 , \11615_b1 );
not ( w_29623 , w_29626 );
not (  , w_29627 );
and ( w_29626 , w_29627 , \11615_b0 );
or ( \11617_b1 , \10965_b1 , w_29629 );
not ( w_29629 , w_29630 );
and ( \11617_b0 , \10965_b0 , w_29631 );
and ( w_29630 ,  , w_29631 );
buf ( w_29629 , \11616_b1 );
not ( w_29629 , w_29632 );
not (  , w_29633 );
and ( w_29632 , w_29633 , \11616_b0 );
or ( \11618_b1 , \11473_b1 , \11477_b1 );
not ( \11477_b1 , w_29634 );
and ( \11618_b0 , \11473_b0 , w_29635 );
and ( w_29634 , w_29635 , \11477_b0 );
or ( \11619_b1 , \11477_b1 , \11607_b1 );
not ( \11607_b1 , w_29636 );
and ( \11619_b0 , \11477_b0 , w_29637 );
and ( w_29636 , w_29637 , \11607_b0 );
or ( \11620_b1 , \11473_b1 , \11607_b1 );
not ( \11607_b1 , w_29638 );
and ( \11620_b0 , \11473_b0 , w_29639 );
and ( w_29638 , w_29639 , \11607_b0 );
or ( \11622_b1 , \11596_b1 , \11600_b1 );
not ( \11600_b1 , w_29640 );
and ( \11622_b0 , \11596_b0 , w_29641 );
and ( w_29640 , w_29641 , \11600_b0 );
or ( \11623_b1 , \11600_b1 , \11605_b1 );
not ( \11605_b1 , w_29642 );
and ( \11623_b0 , \11600_b0 , w_29643 );
and ( w_29642 , w_29643 , \11605_b0 );
or ( \11624_b1 , \11596_b1 , \11605_b1 );
not ( \11605_b1 , w_29644 );
and ( \11624_b0 , \11596_b0 , w_29645 );
and ( w_29644 , w_29645 , \11605_b0 );
or ( \11626_b1 , \11536_b1 , \11545_b1 );
not ( \11545_b1 , w_29646 );
and ( \11626_b0 , \11536_b0 , w_29647 );
and ( w_29646 , w_29647 , \11545_b0 );
or ( \11627_b1 , \11545_b1 , \11590_b1 );
not ( \11590_b1 , w_29648 );
and ( \11627_b0 , \11545_b0 , w_29649 );
and ( w_29648 , w_29649 , \11590_b0 );
or ( \11628_b1 , \11536_b1 , \11590_b1 );
not ( \11590_b1 , w_29650 );
and ( \11628_b0 , \11536_b0 , w_29651 );
and ( w_29650 , w_29651 , \11590_b0 );
or ( \11630_b1 , \11625_b1 , \11629_b1 );
xor ( \11630_b0 , \11625_b0 , w_29652 );
not ( w_29652 , w_29653 );
and ( w_29653 , \11629_b1 , \11629_b0 );
or ( \11631_b1 , \11505_b1 , \11516_b1 );
not ( \11516_b1 , w_29654 );
and ( \11631_b0 , \11505_b0 , w_29655 );
and ( w_29654 , w_29655 , \11516_b0 );
or ( \11632_b1 , \11516_b1 , \11531_b1 );
not ( \11531_b1 , w_29656 );
and ( \11632_b0 , \11516_b0 , w_29657 );
and ( w_29656 , w_29657 , \11531_b0 );
or ( \11633_b1 , \11505_b1 , \11531_b1 );
not ( \11531_b1 , w_29658 );
and ( \11633_b0 , \11505_b0 , w_29659 );
and ( w_29658 , w_29659 , \11531_b0 );
or ( \11635_b1 , \11630_b1 , \11634_b1 );
xor ( \11635_b0 , \11630_b0 , w_29660 );
not ( w_29660 , w_29661 );
and ( w_29661 , \11634_b1 , \11634_b0 );
or ( \11636_b1 , \11621_b1 , \11635_b1 );
xor ( \11636_b0 , \11621_b0 , w_29662 );
not ( w_29662 , w_29663 );
and ( w_29663 , \11635_b1 , \11635_b0 );
or ( \11637_b1 , \11461_b1 , \11465_b1 );
not ( \11465_b1 , w_29664 );
and ( \11637_b0 , \11461_b0 , w_29665 );
and ( w_29664 , w_29665 , \11465_b0 );
or ( \11638_b1 , \11465_b1 , \11467_b1 );
not ( \11467_b1 , w_29666 );
and ( \11638_b0 , \11465_b0 , w_29667 );
and ( w_29666 , w_29667 , \11467_b0 );
or ( \11639_b1 , \11461_b1 , \11467_b1 );
not ( \11467_b1 , w_29668 );
and ( \11639_b0 , \11461_b0 , w_29669 );
and ( w_29668 , w_29669 , \11467_b0 );
or ( \11641_b1 , \11532_b1 , \11591_b1 );
not ( \11591_b1 , w_29670 );
and ( \11641_b0 , \11532_b0 , w_29671 );
and ( w_29670 , w_29671 , \11591_b0 );
or ( \11642_b1 , \11591_b1 , \11606_b1 );
not ( \11606_b1 , w_29672 );
and ( \11642_b0 , \11591_b0 , w_29673 );
and ( w_29672 , w_29673 , \11606_b0 );
or ( \11643_b1 , \11532_b1 , \11606_b1 );
not ( \11606_b1 , w_29674 );
and ( \11643_b0 , \11532_b0 , w_29675 );
and ( w_29674 , w_29675 , \11606_b0 );
or ( \11645_b1 , \11640_b1 , \11644_b1 );
xor ( \11645_b0 , \11640_b0 , w_29676 );
not ( w_29676 , w_29677 );
and ( w_29677 , \11644_b1 , \11644_b0 );
or ( \11646_b1 , \11550_b1 , \11554_b1 );
not ( \11554_b1 , w_29678 );
and ( \11646_b0 , \11550_b0 , w_29679 );
and ( w_29678 , w_29679 , \11554_b0 );
or ( \11647_b1 , \11554_b1 , \11559_b1 );
not ( \11559_b1 , w_29680 );
and ( \11647_b0 , \11554_b0 , w_29681 );
and ( w_29680 , w_29681 , \11559_b0 );
or ( \11648_b1 , \11550_b1 , \11559_b1 );
not ( \11559_b1 , w_29682 );
and ( \11648_b0 , \11550_b0 , w_29683 );
and ( w_29682 , w_29683 , \11559_b0 );
or ( \11650_b1 , \11494_b1 , \11498_b1 );
not ( \11498_b1 , w_29684 );
and ( \11650_b0 , \11494_b0 , w_29685 );
and ( w_29684 , w_29685 , \11498_b0 );
or ( \11651_b1 , \11498_b1 , \11503_b1 );
not ( \11503_b1 , w_29686 );
and ( \11651_b0 , \11498_b0 , w_29687 );
and ( w_29686 , w_29687 , \11503_b0 );
or ( \11652_b1 , \11494_b1 , \11503_b1 );
not ( \11503_b1 , w_29688 );
and ( \11652_b0 , \11494_b0 , w_29689 );
and ( w_29688 , w_29689 , \11503_b0 );
or ( \11654_b1 , \11649_b1 , \11653_b1 );
xor ( \11654_b0 , \11649_b0 , w_29690 );
not ( w_29690 , w_29691 );
and ( w_29691 , \11653_b1 , \11653_b0 );
or ( \11655_b1 , \11482_b1 , \11486_b1 );
not ( \11486_b1 , w_29692 );
and ( \11655_b0 , \11482_b0 , w_29693 );
and ( w_29692 , w_29693 , \11486_b0 );
or ( \11656_b1 , \11486_b1 , \11489_b1 );
not ( \11489_b1 , w_29694 );
and ( \11656_b0 , \11486_b0 , w_29695 );
and ( w_29694 , w_29695 , \11489_b0 );
or ( \11657_b1 , \11482_b1 , \11489_b1 );
not ( \11489_b1 , w_29696 );
and ( \11657_b0 , \11482_b0 , w_29697 );
and ( w_29696 , w_29697 , \11489_b0 );
or ( \11659_b1 , \11654_b1 , \11658_b1 );
xor ( \11659_b0 , \11654_b0 , w_29698 );
not ( w_29698 , w_29699 );
and ( w_29699 , \11658_b1 , \11658_b0 );
or ( \11660_b1 , \6046_b1 , \11539_b1 );
not ( \11539_b1 , w_29700 );
and ( \11660_b0 , \6046_b0 , w_29701 );
and ( w_29700 , w_29701 , \11539_b0 );
or ( \11661_b1 , \11539_b1 , \11544_b1 );
not ( \11544_b1 , w_29702 );
and ( \11661_b0 , \11539_b0 , w_29703 );
and ( w_29702 , w_29703 , \11544_b0 );
or ( \11662_b1 , \6046_b1 , \11544_b1 );
not ( \11544_b1 , w_29704 );
and ( \11662_b0 , \6046_b0 , w_29705 );
and ( w_29704 , w_29705 , \11544_b0 );
or ( \11664_b1 , \11579_b1 , \11583_b1 );
not ( \11583_b1 , w_29706 );
and ( \11664_b0 , \11579_b0 , w_29707 );
and ( w_29706 , w_29707 , \11583_b0 );
or ( \11665_b1 , \11583_b1 , \11588_b1 );
not ( \11588_b1 , w_29708 );
and ( \11665_b0 , \11583_b0 , w_29709 );
and ( w_29708 , w_29709 , \11588_b0 );
or ( \11666_b1 , \11579_b1 , \11588_b1 );
not ( \11588_b1 , w_29710 );
and ( \11666_b0 , \11579_b0 , w_29711 );
and ( w_29710 , w_29711 , \11588_b0 );
or ( \11668_b1 , \11663_b1 , \11667_b1 );
xor ( \11668_b0 , \11663_b0 , w_29712 );
not ( w_29712 , w_29713 );
and ( w_29713 , \11667_b1 , \11667_b0 );
or ( \11669_b1 , \11564_b1 , \11568_b1 );
not ( \11568_b1 , w_29714 );
and ( \11669_b0 , \11564_b0 , w_29715 );
and ( w_29714 , w_29715 , \11568_b0 );
or ( \11670_b1 , \11568_b1 , \11573_b1 );
not ( \11573_b1 , w_29716 );
and ( \11670_b0 , \11568_b0 , w_29717 );
and ( w_29716 , w_29717 , \11573_b0 );
or ( \11671_b1 , \11564_b1 , \11573_b1 );
not ( \11573_b1 , w_29718 );
and ( \11671_b0 , \11564_b0 , w_29719 );
and ( w_29718 , w_29719 , \11573_b0 );
or ( \11673_b1 , \11668_b1 , \11672_b1 );
xor ( \11673_b0 , \11668_b0 , w_29720 );
not ( w_29720 , w_29721 );
and ( w_29721 , \11672_b1 , \11672_b0 );
or ( \11674_b1 , \11659_b1 , \11673_b1 );
xor ( \11674_b0 , \11659_b0 , w_29722 );
not ( w_29722 , w_29723 );
and ( w_29723 , \11673_b1 , \11673_b0 );
or ( \11675_b1 , \11560_b1 , \11574_b1 );
not ( \11574_b1 , w_29724 );
and ( \11675_b0 , \11560_b0 , w_29725 );
and ( w_29724 , w_29725 , \11574_b0 );
or ( \11676_b1 , \11574_b1 , \11589_b1 );
not ( \11589_b1 , w_29726 );
and ( \11676_b0 , \11574_b0 , w_29727 );
and ( w_29726 , w_29727 , \11589_b0 );
or ( \11677_b1 , \11560_b1 , \11589_b1 );
not ( \11589_b1 , w_29728 );
and ( \11677_b0 , \11560_b0 , w_29729 );
and ( w_29728 , w_29729 , \11589_b0 );
or ( \11679_b1 , \5873_b1 , \5829_b1 );
not ( \5829_b1 , w_29730 );
and ( \11679_b0 , \5873_b0 , w_29731 );
and ( w_29730 , w_29731 , \5829_b0 );
or ( \11680_b1 , \5842_b1 , \5827_b1 );
not ( \5827_b1 , w_29732 );
and ( \11680_b0 , \5842_b0 , w_29733 );
and ( w_29732 , w_29733 , \5827_b0 );
or ( \11681_b1 , \11679_b1 , w_29735 );
not ( w_29735 , w_29736 );
and ( \11681_b0 , \11679_b0 , w_29737 );
and ( w_29736 ,  , w_29737 );
buf ( w_29735 , \11680_b1 );
not ( w_29735 , w_29738 );
not (  , w_29739 );
and ( w_29738 , w_29739 , \11680_b0 );
or ( \11682_b1 , \11681_b1 , w_29740 );
xor ( \11682_b0 , \11681_b0 , w_29742 );
not ( w_29742 , w_29743 );
and ( w_29743 , w_29740 , w_29741 );
buf ( w_29740 , \5836_b1 );
not ( w_29740 , w_29744 );
not ( w_29741 , w_29745 );
and ( w_29744 , w_29745 , \5836_b0 );
or ( \11683_b1 , \5893_b1 , \5852_b1 );
not ( \5852_b1 , w_29746 );
and ( \11683_b0 , \5893_b0 , w_29747 );
and ( w_29746 , w_29747 , \5852_b0 );
or ( \11684_b1 , \5861_b1 , \5850_b1 );
not ( \5850_b1 , w_29748 );
and ( \11684_b0 , \5861_b0 , w_29749 );
and ( w_29748 , w_29749 , \5850_b0 );
or ( \11685_b1 , \11683_b1 , w_29751 );
not ( w_29751 , w_29752 );
and ( \11685_b0 , \11683_b0 , w_29753 );
and ( w_29752 ,  , w_29753 );
buf ( w_29751 , \11684_b1 );
not ( w_29751 , w_29754 );
not (  , w_29755 );
and ( w_29754 , w_29755 , \11684_b0 );
or ( \11686_b1 , \11685_b1 , w_29756 );
xor ( \11686_b0 , \11685_b0 , w_29758 );
not ( w_29758 , w_29759 );
and ( w_29759 , w_29756 , w_29757 );
buf ( w_29756 , \5859_b1 );
not ( w_29756 , w_29760 );
not ( w_29757 , w_29761 );
and ( w_29760 , w_29761 , \5859_b0 );
or ( \11687_b1 , \11682_b1 , \11686_b1 );
xor ( \11687_b0 , \11682_b0 , w_29762 );
not ( w_29762 , w_29763 );
and ( w_29763 , \11686_b1 , \11686_b0 );
or ( \11688_b1 , \5918_b1 , \5871_b1 );
not ( \5871_b1 , w_29764 );
and ( \11688_b0 , \5918_b0 , w_29765 );
and ( w_29764 , w_29765 , \5871_b0 );
or ( \11689_b1 , \5881_b1 , \5869_b1 );
not ( \5869_b1 , w_29766 );
and ( \11689_b0 , \5881_b0 , w_29767 );
and ( w_29766 , w_29767 , \5869_b0 );
or ( \11690_b1 , \11688_b1 , w_29769 );
not ( w_29769 , w_29770 );
and ( \11690_b0 , \11688_b0 , w_29771 );
and ( w_29770 ,  , w_29771 );
buf ( w_29769 , \11689_b1 );
not ( w_29769 , w_29772 );
not (  , w_29773 );
and ( w_29772 , w_29773 , \11689_b0 );
or ( \11691_b1 , \11690_b1 , w_29774 );
xor ( \11691_b0 , \11690_b0 , w_29776 );
not ( w_29776 , w_29777 );
and ( w_29777 , w_29774 , w_29775 );
buf ( w_29774 , \5878_b1 );
not ( w_29774 , w_29778 );
not ( w_29775 , w_29779 );
and ( w_29778 , w_29779 , \5878_b0 );
or ( \11692_b1 , \11687_b1 , \11691_b1 );
xor ( \11692_b0 , \11687_b0 , w_29780 );
not ( w_29780 , w_29781 );
and ( w_29781 , \11691_b1 , \11691_b0 );
or ( \11693_b1 , \5811_b1 , \5768_b1 );
not ( \5768_b1 , w_29782 );
and ( \11693_b0 , \5811_b0 , w_29783 );
and ( w_29782 , w_29783 , \5768_b0 );
or ( \11694_b1 , \5780_b1 , \5766_b1 );
not ( \5766_b1 , w_29784 );
and ( \11694_b0 , \5780_b0 , w_29785 );
and ( w_29784 , w_29785 , \5766_b0 );
or ( \11695_b1 , \11693_b1 , w_29787 );
not ( w_29787 , w_29788 );
and ( \11695_b0 , \11693_b0 , w_29789 );
and ( w_29788 ,  , w_29789 );
buf ( w_29787 , \11694_b1 );
not ( w_29787 , w_29790 );
not (  , w_29791 );
and ( w_29790 , w_29791 , \11694_b0 );
or ( \11696_b1 , \11695_b1 , w_29792 );
xor ( \11696_b0 , \11695_b0 , w_29794 );
not ( w_29794 , w_29795 );
and ( w_29795 , w_29792 , w_29793 );
buf ( w_29792 , \5775_b1 );
not ( w_29792 , w_29796 );
not ( w_29793 , w_29797 );
and ( w_29796 , w_29797 , \5775_b0 );
or ( \11697_b1 , \5831_b1 , \5790_b1 );
not ( \5790_b1 , w_29798 );
and ( \11697_b0 , \5831_b0 , w_29799 );
and ( w_29798 , w_29799 , \5790_b0 );
or ( \11698_b1 , \5799_b1 , \5788_b1 );
not ( \5788_b1 , w_29800 );
and ( \11698_b0 , \5799_b0 , w_29801 );
and ( w_29800 , w_29801 , \5788_b0 );
or ( \11699_b1 , \11697_b1 , w_29803 );
not ( w_29803 , w_29804 );
and ( \11699_b0 , \11697_b0 , w_29805 );
and ( w_29804 ,  , w_29805 );
buf ( w_29803 , \11698_b1 );
not ( w_29803 , w_29806 );
not (  , w_29807 );
and ( w_29806 , w_29807 , \11698_b0 );
or ( \11700_b1 , \11699_b1 , w_29808 );
xor ( \11700_b0 , \11699_b0 , w_29810 );
not ( w_29810 , w_29811 );
and ( w_29811 , w_29808 , w_29809 );
buf ( w_29808 , \5797_b1 );
not ( w_29808 , w_29812 );
not ( w_29809 , w_29813 );
and ( w_29812 , w_29813 , \5797_b0 );
or ( \11701_b1 , \11696_b1 , \11700_b1 );
xor ( \11701_b0 , \11696_b0 , w_29814 );
not ( w_29814 , w_29815 );
and ( w_29815 , \11700_b1 , \11700_b0 );
or ( \11702_b1 , \5854_b1 , \5809_b1 );
not ( \5809_b1 , w_29816 );
and ( \11702_b0 , \5854_b0 , w_29817 );
and ( w_29816 , w_29817 , \5809_b0 );
or ( \11703_b1 , \5819_b1 , \5807_b1 );
not ( \5807_b1 , w_29818 );
and ( \11703_b0 , \5819_b0 , w_29819 );
and ( w_29818 , w_29819 , \5807_b0 );
or ( \11704_b1 , \11702_b1 , w_29821 );
not ( w_29821 , w_29822 );
and ( \11704_b0 , \11702_b0 , w_29823 );
and ( w_29822 ,  , w_29823 );
buf ( w_29821 , \11703_b1 );
not ( w_29821 , w_29824 );
not (  , w_29825 );
and ( w_29824 , w_29825 , \11703_b0 );
or ( \11705_b1 , \11704_b1 , w_29826 );
xor ( \11705_b0 , \11704_b0 , w_29828 );
not ( w_29828 , w_29829 );
and ( w_29829 , w_29826 , w_29827 );
buf ( w_29826 , \5816_b1 );
not ( w_29826 , w_29830 );
not ( w_29827 , w_29831 );
and ( w_29830 , w_29831 , \5816_b0 );
or ( \11706_b1 , \11701_b1 , \11705_b1 );
xor ( \11706_b0 , \11701_b0 , w_29832 );
not ( w_29832 , w_29833 );
and ( w_29833 , \11705_b1 , \11705_b0 );
or ( \11707_b1 , \11692_b1 , \11706_b1 );
xor ( \11707_b0 , \11692_b0 , w_29834 );
not ( w_29834 , w_29835 );
and ( w_29835 , \11706_b1 , \11706_b0 );
buf ( \11708_b1 , \7198_b1 );
not ( \11708_b1 , w_29836 );
not ( \11708_b0 , w_29837 );
and ( w_29836 , w_29837 , \7198_b0 );
or ( \11709_b1 , \5770_b1 , \7203_b1 );
not ( \7203_b1 , w_29838 );
and ( \11709_b0 , \5770_b0 , w_29839 );
and ( w_29838 , w_29839 , \7203_b0 );
or ( \11710_b1 , \5737_b1 , \7201_b1 );
not ( \7201_b1 , w_29840 );
and ( \11710_b0 , \5737_b0 , w_29841 );
and ( w_29840 , w_29841 , \7201_b0 );
or ( \11711_b1 , \11709_b1 , w_29843 );
not ( w_29843 , w_29844 );
and ( \11711_b0 , \11709_b0 , w_29845 );
and ( w_29844 ,  , w_29845 );
buf ( w_29843 , \11710_b1 );
not ( w_29843 , w_29846 );
not (  , w_29847 );
and ( w_29846 , w_29847 , \11710_b0 );
or ( \11712_b1 , \11711_b1 , w_29848 );
xor ( \11712_b0 , \11711_b0 , w_29850 );
not ( w_29850 , w_29851 );
and ( w_29851 , w_29848 , w_29849 );
buf ( w_29848 , \6824_b1 );
not ( w_29848 , w_29852 );
not ( w_29849 , w_29853 );
and ( w_29852 , w_29853 , \6824_b0 );
or ( \11713_b1 , \11708_b1 , \11712_b1 );
xor ( \11713_b0 , \11708_b0 , w_29854 );
not ( w_29854 , w_29855 );
and ( w_29855 , \11712_b1 , \11712_b0 );
or ( \11714_b1 , \5792_b1 , \5750_b1 );
not ( \5750_b1 , w_29856 );
and ( \11714_b0 , \5792_b0 , w_29857 );
and ( w_29856 , w_29857 , \5750_b0 );
or ( \11715_b1 , \5758_b1 , \5748_b1 );
not ( \5748_b1 , w_29858 );
and ( \11715_b0 , \5758_b0 , w_29859 );
and ( w_29858 , w_29859 , \5748_b0 );
or ( \11716_b1 , \11714_b1 , w_29861 );
not ( w_29861 , w_29862 );
and ( \11716_b0 , \11714_b0 , w_29863 );
and ( w_29862 ,  , w_29863 );
buf ( w_29861 , \11715_b1 );
not ( w_29861 , w_29864 );
not (  , w_29865 );
and ( w_29864 , w_29865 , \11715_b0 );
or ( \11717_b1 , \11716_b1 , w_29866 );
xor ( \11717_b0 , \11716_b0 , w_29868 );
not ( w_29868 , w_29869 );
and ( w_29869 , w_29866 , w_29867 );
buf ( w_29866 , \5755_b1 );
not ( w_29866 , w_29870 );
not ( w_29867 , w_29871 );
and ( w_29870 , w_29871 , \5755_b0 );
or ( \11718_b1 , \11713_b1 , \11717_b1 );
xor ( \11718_b0 , \11713_b0 , w_29872 );
not ( w_29872 , w_29873 );
and ( w_29873 , \11717_b1 , \11717_b0 );
or ( \11719_b1 , \11707_b1 , \11718_b1 );
xor ( \11719_b0 , \11707_b0 , w_29874 );
not ( w_29874 , w_29875 );
and ( w_29875 , \11718_b1 , \11718_b0 );
or ( \11720_b1 , \11678_b1 , \11719_b1 );
xor ( \11720_b0 , \11678_b0 , w_29876 );
not ( w_29876 , w_29877 );
and ( w_29877 , \11719_b1 , \11719_b0 );
or ( \11721_b1 , \6057_b1 , \6016_b1 );
not ( \6016_b1 , w_29878 );
and ( \11721_b0 , \6057_b0 , w_29879 );
and ( w_29878 , w_29879 , \6016_b0 );
or ( \11722_b1 , \6029_b1 , \6014_b1 );
not ( \6014_b1 , w_29880 );
and ( \11722_b0 , \6029_b0 , w_29881 );
and ( w_29880 , w_29881 , \6014_b0 );
or ( \11723_b1 , \11721_b1 , w_29883 );
not ( w_29883 , w_29884 );
and ( \11723_b0 , \11721_b0 , w_29885 );
and ( w_29884 ,  , w_29885 );
buf ( w_29883 , \11722_b1 );
not ( w_29883 , w_29886 );
not (  , w_29887 );
and ( w_29886 , w_29887 , \11722_b0 );
or ( \11724_b1 , \11723_b1 , w_29888 );
xor ( \11724_b0 , \11723_b0 , w_29890 );
not ( w_29890 , w_29891 );
and ( w_29891 , w_29888 , w_29889 );
buf ( w_29888 , \6023_b1 );
not ( w_29888 , w_29892 );
not ( w_29889 , w_29893 );
and ( w_29892 , w_29893 , \6023_b0 );
or ( \11725_b1 , \6065_b1 , \6039_b1 );
not ( \6039_b1 , w_29894 );
and ( \11725_b0 , \6065_b0 , w_29895 );
and ( w_29894 , w_29895 , \6039_b0 );
or ( \11726_b1 , \6048_b1 , \6037_b1 );
not ( \6037_b1 , w_29896 );
and ( \11726_b0 , \6048_b0 , w_29897 );
and ( w_29896 , w_29897 , \6037_b0 );
or ( \11727_b1 , \11725_b1 , w_29899 );
not ( w_29899 , w_29900 );
and ( \11727_b0 , \11725_b0 , w_29901 );
and ( w_29900 ,  , w_29901 );
buf ( w_29899 , \11726_b1 );
not ( w_29899 , w_29902 );
not (  , w_29903 );
and ( w_29902 , w_29903 , \11726_b0 );
or ( \11728_b1 , \11727_b1 , w_29904 );
xor ( \11728_b0 , \11727_b0 , w_29906 );
not ( w_29906 , w_29907 );
and ( w_29907 , w_29904 , w_29905 );
buf ( w_29904 , \6046_b1 );
not ( w_29904 , w_29908 );
not ( w_29905 , w_29909 );
and ( w_29908 , w_29909 , \6046_b0 );
or ( \11729_b1 , \11724_b1 , \11728_b1 );
xor ( \11729_b0 , \11724_b0 , w_29910 );
not ( w_29910 , w_29911 );
and ( w_29911 , \11728_b1 , \11728_b0 );
or ( \11730_b1 , \5998_b1 , \5955_b1 );
not ( \5955_b1 , w_29912 );
and ( \11730_b0 , \5998_b0 , w_29913 );
and ( w_29912 , w_29913 , \5955_b0 );
or ( \11731_b1 , \5967_b1 , \5953_b1 );
not ( \5953_b1 , w_29914 );
and ( \11731_b0 , \5967_b0 , w_29915 );
and ( w_29914 , w_29915 , \5953_b0 );
or ( \11732_b1 , \11730_b1 , w_29917 );
not ( w_29917 , w_29918 );
and ( \11732_b0 , \11730_b0 , w_29919 );
and ( w_29918 ,  , w_29919 );
buf ( w_29917 , \11731_b1 );
not ( w_29917 , w_29920 );
not (  , w_29921 );
and ( w_29920 , w_29921 , \11731_b0 );
or ( \11733_b1 , \11732_b1 , w_29922 );
xor ( \11733_b0 , \11732_b0 , w_29924 );
not ( w_29924 , w_29925 );
and ( w_29925 , w_29922 , w_29923 );
buf ( w_29922 , \5962_b1 );
not ( w_29922 , w_29926 );
not ( w_29923 , w_29927 );
and ( w_29926 , w_29927 , \5962_b0 );
or ( \11734_b1 , \6018_b1 , \5977_b1 );
not ( \5977_b1 , w_29928 );
and ( \11734_b0 , \6018_b0 , w_29929 );
and ( w_29928 , w_29929 , \5977_b0 );
or ( \11735_b1 , \5986_b1 , \5975_b1 );
not ( \5975_b1 , w_29930 );
and ( \11735_b0 , \5986_b0 , w_29931 );
and ( w_29930 , w_29931 , \5975_b0 );
or ( \11736_b1 , \11734_b1 , w_29933 );
not ( w_29933 , w_29934 );
and ( \11736_b0 , \11734_b0 , w_29935 );
and ( w_29934 ,  , w_29935 );
buf ( w_29933 , \11735_b1 );
not ( w_29933 , w_29936 );
not (  , w_29937 );
and ( w_29936 , w_29937 , \11735_b0 );
or ( \11737_b1 , \11736_b1 , w_29938 );
xor ( \11737_b0 , \11736_b0 , w_29940 );
not ( w_29940 , w_29941 );
and ( w_29941 , w_29938 , w_29939 );
buf ( w_29938 , \5984_b1 );
not ( w_29938 , w_29942 );
not ( w_29939 , w_29943 );
and ( w_29942 , w_29943 , \5984_b0 );
or ( \11738_b1 , \11733_b1 , \11737_b1 );
xor ( \11738_b0 , \11733_b0 , w_29944 );
not ( w_29944 , w_29945 );
and ( w_29945 , \11737_b1 , \11737_b0 );
or ( \11739_b1 , \6041_b1 , \5996_b1 );
not ( \5996_b1 , w_29946 );
and ( \11739_b0 , \6041_b0 , w_29947 );
and ( w_29946 , w_29947 , \5996_b0 );
or ( \11740_b1 , \6006_b1 , \5994_b1 );
not ( \5994_b1 , w_29948 );
and ( \11740_b0 , \6006_b0 , w_29949 );
and ( w_29948 , w_29949 , \5994_b0 );
or ( \11741_b1 , \11739_b1 , w_29951 );
not ( w_29951 , w_29952 );
and ( \11741_b0 , \11739_b0 , w_29953 );
and ( w_29952 ,  , w_29953 );
buf ( w_29951 , \11740_b1 );
not ( w_29951 , w_29954 );
not (  , w_29955 );
and ( w_29954 , w_29955 , \11740_b0 );
or ( \11742_b1 , \11741_b1 , w_29956 );
xor ( \11742_b0 , \11741_b0 , w_29958 );
not ( w_29958 , w_29959 );
and ( w_29959 , w_29956 , w_29957 );
buf ( w_29956 , \6003_b1 );
not ( w_29956 , w_29960 );
not ( w_29957 , w_29961 );
and ( w_29960 , w_29961 , \6003_b0 );
or ( \11743_b1 , \11738_b1 , \11742_b1 );
xor ( \11743_b0 , \11738_b0 , w_29962 );
not ( w_29962 , w_29963 );
and ( w_29963 , \11742_b1 , \11742_b0 );
or ( \11744_b1 , \11729_b1 , \11743_b1 );
xor ( \11744_b0 , \11729_b0 , w_29964 );
not ( w_29964 , w_29965 );
and ( w_29965 , \11743_b1 , \11743_b0 );
or ( \11745_b1 , \5937_b1 , \5891_b1 );
not ( \5891_b1 , w_29966 );
and ( \11745_b0 , \5937_b0 , w_29967 );
and ( w_29966 , w_29967 , \5891_b0 );
or ( \11746_b1 , \5906_b1 , \5889_b1 );
not ( \5889_b1 , w_29968 );
and ( \11746_b0 , \5906_b0 , w_29969 );
and ( w_29968 , w_29969 , \5889_b0 );
or ( \11747_b1 , \11745_b1 , w_29971 );
not ( w_29971 , w_29972 );
and ( \11747_b0 , \11745_b0 , w_29973 );
and ( w_29972 ,  , w_29973 );
buf ( w_29971 , \11746_b1 );
not ( w_29971 , w_29974 );
not (  , w_29975 );
and ( w_29974 , w_29975 , \11746_b0 );
or ( \11748_b1 , \11747_b1 , w_29976 );
xor ( \11748_b0 , \11747_b0 , w_29978 );
not ( w_29978 , w_29979 );
and ( w_29979 , w_29976 , w_29977 );
buf ( w_29976 , \5898_b1 );
not ( w_29976 , w_29980 );
not ( w_29977 , w_29981 );
and ( w_29980 , w_29981 , \5898_b0 );
or ( \11749_b1 , \5957_b1 , \5916_b1 );
not ( \5916_b1 , w_29982 );
and ( \11749_b0 , \5957_b0 , w_29983 );
and ( w_29982 , w_29983 , \5916_b0 );
or ( \11750_b1 , \5925_b1 , \5914_b1 );
not ( \5914_b1 , w_29984 );
and ( \11750_b0 , \5925_b0 , w_29985 );
and ( w_29984 , w_29985 , \5914_b0 );
or ( \11751_b1 , \11749_b1 , w_29987 );
not ( w_29987 , w_29988 );
and ( \11751_b0 , \11749_b0 , w_29989 );
and ( w_29988 ,  , w_29989 );
buf ( w_29987 , \11750_b1 );
not ( w_29987 , w_29990 );
not (  , w_29991 );
and ( w_29990 , w_29991 , \11750_b0 );
or ( \11752_b1 , \11751_b1 , w_29992 );
xor ( \11752_b0 , \11751_b0 , w_29994 );
not ( w_29994 , w_29995 );
and ( w_29995 , w_29992 , w_29993 );
buf ( w_29992 , \5923_b1 );
not ( w_29992 , w_29996 );
not ( w_29993 , w_29997 );
and ( w_29996 , w_29997 , \5923_b0 );
or ( \11753_b1 , \11748_b1 , \11752_b1 );
xor ( \11753_b0 , \11748_b0 , w_29998 );
not ( w_29998 , w_29999 );
and ( w_29999 , \11752_b1 , \11752_b0 );
or ( \11754_b1 , \5979_b1 , \5935_b1 );
not ( \5935_b1 , w_30000 );
and ( \11754_b0 , \5979_b0 , w_30001 );
and ( w_30000 , w_30001 , \5935_b0 );
or ( \11755_b1 , \5945_b1 , \5933_b1 );
not ( \5933_b1 , w_30002 );
and ( \11755_b0 , \5945_b0 , w_30003 );
and ( w_30002 , w_30003 , \5933_b0 );
or ( \11756_b1 , \11754_b1 , w_30005 );
not ( w_30005 , w_30006 );
and ( \11756_b0 , \11754_b0 , w_30007 );
and ( w_30006 ,  , w_30007 );
buf ( w_30005 , \11755_b1 );
not ( w_30005 , w_30008 );
not (  , w_30009 );
and ( w_30008 , w_30009 , \11755_b0 );
or ( \11757_b1 , \11756_b1 , w_30010 );
xor ( \11757_b0 , \11756_b0 , w_30012 );
not ( w_30012 , w_30013 );
and ( w_30013 , w_30010 , w_30011 );
buf ( w_30010 , \5942_b1 );
not ( w_30010 , w_30014 );
not ( w_30011 , w_30015 );
and ( w_30014 , w_30015 , \5942_b0 );
or ( \11758_b1 , \11753_b1 , \11757_b1 );
xor ( \11758_b0 , \11753_b0 , w_30016 );
not ( w_30016 , w_30017 );
and ( w_30017 , \11757_b1 , \11757_b0 );
or ( \11759_b1 , \11744_b1 , \11758_b1 );
xor ( \11759_b0 , \11744_b0 , w_30018 );
not ( w_30018 , w_30019 );
and ( w_30019 , \11758_b1 , \11758_b0 );
or ( \11760_b1 , \11720_b1 , \11759_b1 );
xor ( \11760_b0 , \11720_b0 , w_30020 );
not ( w_30020 , w_30021 );
and ( w_30021 , \11759_b1 , \11759_b0 );
or ( \11761_b1 , \11674_b1 , \11760_b1 );
xor ( \11761_b0 , \11674_b0 , w_30022 );
not ( w_30022 , w_30023 );
and ( w_30023 , \11760_b1 , \11760_b0 );
or ( \11762_b1 , \11521_b1 , \11525_b1 );
not ( \11525_b1 , w_30024 );
and ( \11762_b0 , \11521_b0 , w_30025 );
and ( w_30024 , w_30025 , \11525_b0 );
or ( \11763_b1 , \11525_b1 , \11530_b1 );
not ( \11530_b1 , w_30026 );
and ( \11763_b0 , \11525_b0 , w_30027 );
and ( w_30026 , w_30027 , \11530_b0 );
or ( \11764_b1 , \11521_b1 , \11530_b1 );
not ( \11530_b1 , w_30028 );
and ( \11764_b0 , \11521_b0 , w_30029 );
and ( w_30028 , w_30029 , \11530_b0 );
or ( \11766_b1 , \11509_b1 , \11513_b1 );
not ( \11513_b1 , w_30030 );
and ( \11766_b0 , \11509_b0 , w_30031 );
and ( w_30030 , w_30031 , \11513_b0 );
or ( \11767_b1 , \11513_b1 , \11515_b1 );
not ( \11515_b1 , w_30032 );
and ( \11767_b0 , \11513_b0 , w_30033 );
and ( w_30032 , w_30033 , \11515_b0 );
or ( \11768_b1 , \11509_b1 , \11515_b1 );
not ( \11515_b1 , w_30034 );
and ( \11768_b0 , \11509_b0 , w_30035 );
and ( w_30034 , w_30035 , \11515_b0 );
or ( \11770_b1 , \11765_b1 , \11769_b1 );
xor ( \11770_b0 , \11765_b0 , w_30036 );
not ( w_30036 , w_30037 );
and ( w_30037 , \11769_b1 , \11769_b0 );
or ( \11771_b1 , \11490_b1 , w_30038 );
or ( \11771_b0 , \11490_b0 , \11504_b0 );
not ( \11504_b0 , w_30039 );
and ( w_30039 , w_30038 , \11504_b1 );
or ( \11772_b1 , \11770_b1 , \11771_b1 );
xor ( \11772_b0 , \11770_b0 , w_30040 );
not ( w_30040 , w_30041 );
and ( w_30041 , \11771_b1 , \11771_b0 );
or ( \11773_b1 , \11761_b1 , \11772_b1 );
xor ( \11773_b0 , \11761_b0 , w_30042 );
not ( w_30042 , w_30043 );
and ( w_30043 , \11772_b1 , \11772_b0 );
or ( \11774_b1 , \11645_b1 , \11773_b1 );
xor ( \11774_b0 , \11645_b0 , w_30044 );
not ( w_30044 , w_30045 );
and ( w_30045 , \11773_b1 , \11773_b0 );
or ( \11775_b1 , \11636_b1 , \11774_b1 );
xor ( \11775_b0 , \11636_b0 , w_30046 );
not ( w_30046 , w_30047 );
and ( w_30047 , \11774_b1 , \11774_b0 );
or ( \11776_b1 , \11457_b1 , \11468_b1 );
not ( \11468_b1 , w_30048 );
and ( \11776_b0 , \11457_b0 , w_30049 );
and ( w_30048 , w_30049 , \11468_b0 );
or ( \11777_b1 , \11468_b1 , \11608_b1 );
not ( \11608_b1 , w_30050 );
and ( \11777_b0 , \11468_b0 , w_30051 );
and ( w_30050 , w_30051 , \11608_b0 );
or ( \11778_b1 , \11457_b1 , \11608_b1 );
not ( \11608_b1 , w_30052 );
and ( \11778_b0 , \11457_b0 , w_30053 );
and ( w_30052 , w_30053 , \11608_b0 );
or ( \11780_b1 , \11775_b1 , w_30055 );
not ( w_30055 , w_30056 );
and ( \11780_b0 , \11775_b0 , w_30057 );
and ( w_30056 ,  , w_30057 );
buf ( w_30055 , \11779_b1 );
not ( w_30055 , w_30058 );
not (  , w_30059 );
and ( w_30058 , w_30059 , \11779_b0 );
or ( \11781_b1 , \11640_b1 , \11644_b1 );
not ( \11644_b1 , w_30060 );
and ( \11781_b0 , \11640_b0 , w_30061 );
and ( w_30060 , w_30061 , \11644_b0 );
or ( \11782_b1 , \11644_b1 , \11773_b1 );
not ( \11773_b1 , w_30062 );
and ( \11782_b0 , \11644_b0 , w_30063 );
and ( w_30062 , w_30063 , \11773_b0 );
or ( \11783_b1 , \11640_b1 , \11773_b1 );
not ( \11773_b1 , w_30064 );
and ( \11783_b0 , \11640_b0 , w_30065 );
and ( w_30064 , w_30065 , \11773_b0 );
or ( \11785_b1 , \11765_b1 , \11769_b1 );
not ( \11769_b1 , w_30066 );
and ( \11785_b0 , \11765_b0 , w_30067 );
and ( w_30066 , w_30067 , \11769_b0 );
or ( \11786_b1 , \11769_b1 , \11771_b1 );
not ( \11771_b1 , w_30068 );
and ( \11786_b0 , \11769_b0 , w_30069 );
and ( w_30068 , w_30069 , \11771_b0 );
or ( \11787_b1 , \11765_b1 , \11771_b1 );
not ( \11771_b1 , w_30070 );
and ( \11787_b0 , \11765_b0 , w_30071 );
and ( w_30070 , w_30071 , \11771_b0 );
or ( \11789_b1 , \11678_b1 , \11719_b1 );
not ( \11719_b1 , w_30072 );
and ( \11789_b0 , \11678_b0 , w_30073 );
and ( w_30072 , w_30073 , \11719_b0 );
or ( \11790_b1 , \11719_b1 , \11759_b1 );
not ( \11759_b1 , w_30074 );
and ( \11790_b0 , \11719_b0 , w_30075 );
and ( w_30074 , w_30075 , \11759_b0 );
or ( \11791_b1 , \11678_b1 , \11759_b1 );
not ( \11759_b1 , w_30076 );
and ( \11791_b0 , \11678_b0 , w_30077 );
and ( w_30076 , w_30077 , \11759_b0 );
or ( \11793_b1 , \11788_b1 , \11792_b1 );
xor ( \11793_b0 , \11788_b0 , w_30078 );
not ( w_30078 , w_30079 );
and ( w_30079 , \11792_b1 , \11792_b0 );
or ( \11794_b1 , \11659_b1 , \11673_b1 );
not ( \11673_b1 , w_30080 );
and ( \11794_b0 , \11659_b0 , w_30081 );
and ( w_30080 , w_30081 , \11673_b0 );
or ( \11795_b1 , \11793_b1 , \11794_b1 );
xor ( \11795_b0 , \11793_b0 , w_30082 );
not ( w_30082 , w_30083 );
and ( w_30083 , \11794_b1 , \11794_b0 );
or ( \11796_b1 , \11784_b1 , \11795_b1 );
xor ( \11796_b0 , \11784_b0 , w_30084 );
not ( w_30084 , w_30085 );
and ( w_30085 , \11795_b1 , \11795_b0 );
or ( \11797_b1 , \11625_b1 , \11629_b1 );
not ( \11629_b1 , w_30086 );
and ( \11797_b0 , \11625_b0 , w_30087 );
and ( w_30086 , w_30087 , \11629_b0 );
or ( \11798_b1 , \11629_b1 , \11634_b1 );
not ( \11634_b1 , w_30088 );
and ( \11798_b0 , \11629_b0 , w_30089 );
and ( w_30088 , w_30089 , \11634_b0 );
or ( \11799_b1 , \11625_b1 , \11634_b1 );
not ( \11634_b1 , w_30090 );
and ( \11799_b0 , \11625_b0 , w_30091 );
and ( w_30090 , w_30091 , \11634_b0 );
or ( \11801_b1 , \11674_b1 , \11760_b1 );
not ( \11760_b1 , w_30092 );
and ( \11801_b0 , \11674_b0 , w_30093 );
and ( w_30092 , w_30093 , \11760_b0 );
or ( \11802_b1 , \11760_b1 , \11772_b1 );
not ( \11772_b1 , w_30094 );
and ( \11802_b0 , \11760_b0 , w_30095 );
and ( w_30094 , w_30095 , \11772_b0 );
or ( \11803_b1 , \11674_b1 , \11772_b1 );
not ( \11772_b1 , w_30096 );
and ( \11803_b0 , \11674_b0 , w_30097 );
and ( w_30096 , w_30097 , \11772_b0 );
or ( \11805_b1 , \11800_b1 , \11804_b1 );
xor ( \11805_b0 , \11800_b0 , w_30098 );
not ( w_30098 , w_30099 );
and ( w_30099 , \11804_b1 , \11804_b0 );
or ( \11806_b1 , \6029_b1 , \6016_b1 );
not ( \6016_b1 , w_30100 );
and ( \11806_b0 , \6029_b0 , w_30101 );
and ( w_30100 , w_30101 , \6016_b0 );
or ( \11807_b1 , \6041_b1 , \6014_b1 );
not ( \6014_b1 , w_30102 );
and ( \11807_b0 , \6041_b0 , w_30103 );
and ( w_30102 , w_30103 , \6014_b0 );
or ( \11808_b1 , \11806_b1 , w_30105 );
not ( w_30105 , w_30106 );
and ( \11808_b0 , \11806_b0 , w_30107 );
and ( w_30106 ,  , w_30107 );
buf ( w_30105 , \11807_b1 );
not ( w_30105 , w_30108 );
not (  , w_30109 );
and ( w_30108 , w_30109 , \11807_b0 );
or ( \11809_b1 , \11808_b1 , w_30110 );
xor ( \11809_b0 , \11808_b0 , w_30112 );
not ( w_30112 , w_30113 );
and ( w_30113 , w_30110 , w_30111 );
buf ( w_30110 , \6023_b1 );
not ( w_30110 , w_30114 );
not ( w_30111 , w_30115 );
and ( w_30114 , w_30115 , \6023_b0 );
or ( \11810_b1 , \6048_b1 , \6039_b1 );
not ( \6039_b1 , w_30116 );
and ( \11810_b0 , \6048_b0 , w_30117 );
and ( w_30116 , w_30117 , \6039_b0 );
or ( \11811_b1 , \6057_b1 , \6037_b1 );
not ( \6037_b1 , w_30118 );
and ( \11811_b0 , \6057_b0 , w_30119 );
and ( w_30118 , w_30119 , \6037_b0 );
or ( \11812_b1 , \11810_b1 , w_30121 );
not ( w_30121 , w_30122 );
and ( \11812_b0 , \11810_b0 , w_30123 );
and ( w_30122 ,  , w_30123 );
buf ( w_30121 , \11811_b1 );
not ( w_30121 , w_30124 );
not (  , w_30125 );
and ( w_30124 , w_30125 , \11811_b0 );
or ( \11813_b1 , \11812_b1 , w_30126 );
xor ( \11813_b0 , \11812_b0 , w_30128 );
not ( w_30128 , w_30129 );
and ( w_30129 , w_30126 , w_30127 );
buf ( w_30126 , \6046_b1 );
not ( w_30126 , w_30130 );
not ( w_30127 , w_30131 );
and ( w_30130 , w_30131 , \6046_b0 );
or ( \11814_b1 , \11809_b1 , \11813_b1 );
xor ( \11814_b0 , \11809_b0 , w_30132 );
not ( w_30132 , w_30133 );
and ( w_30133 , \11813_b1 , \11813_b0 );
or ( \11815_b1 , \6065_b1 , w_30135 );
not ( w_30135 , w_30136 );
and ( \11815_b0 , \6065_b0 , w_30137 );
and ( w_30136 ,  , w_30137 );
buf ( w_30135 , \6053_b1 );
not ( w_30135 , w_30138 );
not (  , w_30139 );
and ( w_30138 , w_30139 , \6053_b0 );
or ( \11816_b1 , \11815_b1 , w_30140 );
xor ( \11816_b0 , \11815_b0 , w_30142 );
not ( w_30142 , w_30143 );
and ( w_30143 , w_30140 , w_30141 );
buf ( w_30140 , \6062_b1 );
not ( w_30140 , w_30144 );
not ( w_30141 , w_30145 );
and ( w_30144 , w_30145 , \6062_b0 );
or ( \11817_b1 , \11814_b1 , \11816_b1 );
xor ( \11817_b0 , \11814_b0 , w_30146 );
not ( w_30146 , w_30147 );
and ( w_30147 , \11816_b1 , \11816_b0 );
or ( \11818_b1 , \5967_b1 , \5955_b1 );
not ( \5955_b1 , w_30148 );
and ( \11818_b0 , \5967_b0 , w_30149 );
and ( w_30148 , w_30149 , \5955_b0 );
or ( \11819_b1 , \5979_b1 , \5953_b1 );
not ( \5953_b1 , w_30150 );
and ( \11819_b0 , \5979_b0 , w_30151 );
and ( w_30150 , w_30151 , \5953_b0 );
or ( \11820_b1 , \11818_b1 , w_30153 );
not ( w_30153 , w_30154 );
and ( \11820_b0 , \11818_b0 , w_30155 );
and ( w_30154 ,  , w_30155 );
buf ( w_30153 , \11819_b1 );
not ( w_30153 , w_30156 );
not (  , w_30157 );
and ( w_30156 , w_30157 , \11819_b0 );
or ( \11821_b1 , \11820_b1 , w_30158 );
xor ( \11821_b0 , \11820_b0 , w_30160 );
not ( w_30160 , w_30161 );
and ( w_30161 , w_30158 , w_30159 );
buf ( w_30158 , \5962_b1 );
not ( w_30158 , w_30162 );
not ( w_30159 , w_30163 );
and ( w_30162 , w_30163 , \5962_b0 );
or ( \11822_b1 , \5986_b1 , \5977_b1 );
not ( \5977_b1 , w_30164 );
and ( \11822_b0 , \5986_b0 , w_30165 );
and ( w_30164 , w_30165 , \5977_b0 );
or ( \11823_b1 , \5998_b1 , \5975_b1 );
not ( \5975_b1 , w_30166 );
and ( \11823_b0 , \5998_b0 , w_30167 );
and ( w_30166 , w_30167 , \5975_b0 );
or ( \11824_b1 , \11822_b1 , w_30169 );
not ( w_30169 , w_30170 );
and ( \11824_b0 , \11822_b0 , w_30171 );
and ( w_30170 ,  , w_30171 );
buf ( w_30169 , \11823_b1 );
not ( w_30169 , w_30172 );
not (  , w_30173 );
and ( w_30172 , w_30173 , \11823_b0 );
or ( \11825_b1 , \11824_b1 , w_30174 );
xor ( \11825_b0 , \11824_b0 , w_30176 );
not ( w_30176 , w_30177 );
and ( w_30177 , w_30174 , w_30175 );
buf ( w_30174 , \5984_b1 );
not ( w_30174 , w_30178 );
not ( w_30175 , w_30179 );
and ( w_30178 , w_30179 , \5984_b0 );
or ( \11826_b1 , \11821_b1 , \11825_b1 );
xor ( \11826_b0 , \11821_b0 , w_30180 );
not ( w_30180 , w_30181 );
and ( w_30181 , \11825_b1 , \11825_b0 );
or ( \11827_b1 , \6006_b1 , \5996_b1 );
not ( \5996_b1 , w_30182 );
and ( \11827_b0 , \6006_b0 , w_30183 );
and ( w_30182 , w_30183 , \5996_b0 );
or ( \11828_b1 , \6018_b1 , \5994_b1 );
not ( \5994_b1 , w_30184 );
and ( \11828_b0 , \6018_b0 , w_30185 );
and ( w_30184 , w_30185 , \5994_b0 );
or ( \11829_b1 , \11827_b1 , w_30187 );
not ( w_30187 , w_30188 );
and ( \11829_b0 , \11827_b0 , w_30189 );
and ( w_30188 ,  , w_30189 );
buf ( w_30187 , \11828_b1 );
not ( w_30187 , w_30190 );
not (  , w_30191 );
and ( w_30190 , w_30191 , \11828_b0 );
or ( \11830_b1 , \11829_b1 , w_30192 );
xor ( \11830_b0 , \11829_b0 , w_30194 );
not ( w_30194 , w_30195 );
and ( w_30195 , w_30192 , w_30193 );
buf ( w_30192 , \6003_b1 );
not ( w_30192 , w_30196 );
not ( w_30193 , w_30197 );
and ( w_30196 , w_30197 , \6003_b0 );
or ( \11831_b1 , \11826_b1 , \11830_b1 );
xor ( \11831_b0 , \11826_b0 , w_30198 );
not ( w_30198 , w_30199 );
and ( w_30199 , \11830_b1 , \11830_b0 );
or ( \11832_b1 , \11817_b1 , w_30200 );
xor ( \11832_b0 , \11817_b0 , w_30202 );
not ( w_30202 , w_30203 );
and ( w_30203 , w_30200 , w_30201 );
buf ( w_30200 , \11831_b1 );
not ( w_30200 , w_30204 );
not ( w_30201 , w_30205 );
and ( w_30204 , w_30205 , \11831_b0 );
or ( \11833_b1 , \11748_b1 , \11752_b1 );
not ( \11752_b1 , w_30206 );
and ( \11833_b0 , \11748_b0 , w_30207 );
and ( w_30206 , w_30207 , \11752_b0 );
or ( \11834_b1 , \11752_b1 , \11757_b1 );
not ( \11757_b1 , w_30208 );
and ( \11834_b0 , \11752_b0 , w_30209 );
and ( w_30208 , w_30209 , \11757_b0 );
or ( \11835_b1 , \11748_b1 , \11757_b1 );
not ( \11757_b1 , w_30210 );
and ( \11835_b0 , \11748_b0 , w_30211 );
and ( w_30210 , w_30211 , \11757_b0 );
or ( \11837_b1 , \11733_b1 , \11737_b1 );
not ( \11737_b1 , w_30212 );
and ( \11837_b0 , \11733_b0 , w_30213 );
and ( w_30212 , w_30213 , \11737_b0 );
or ( \11838_b1 , \11737_b1 , \11742_b1 );
not ( \11742_b1 , w_30214 );
and ( \11838_b0 , \11737_b0 , w_30215 );
and ( w_30214 , w_30215 , \11742_b0 );
or ( \11839_b1 , \11733_b1 , \11742_b1 );
not ( \11742_b1 , w_30216 );
and ( \11839_b0 , \11733_b0 , w_30217 );
and ( w_30216 , w_30217 , \11742_b0 );
or ( \11841_b1 , \11836_b1 , \11840_b1 );
xor ( \11841_b0 , \11836_b0 , w_30218 );
not ( w_30218 , w_30219 );
and ( w_30219 , \11840_b1 , \11840_b0 );
or ( \11842_b1 , \11724_b1 , \11728_b1 );
not ( \11728_b1 , w_30220 );
and ( \11842_b0 , \11724_b0 , w_30221 );
and ( w_30220 , w_30221 , \11728_b0 );
or ( \11843_b1 , \11841_b1 , \11842_b1 );
xor ( \11843_b0 , \11841_b0 , w_30222 );
not ( w_30222 , w_30223 );
and ( w_30223 , \11842_b1 , \11842_b0 );
or ( \11844_b1 , \11832_b1 , \11843_b1 );
xor ( \11844_b0 , \11832_b0 , w_30224 );
not ( w_30224 , w_30225 );
and ( w_30225 , \11843_b1 , \11843_b0 );
or ( \11845_b1 , \11708_b1 , \11712_b1 );
not ( \11712_b1 , w_30226 );
and ( \11845_b0 , \11708_b0 , w_30227 );
and ( w_30226 , w_30227 , \11712_b0 );
or ( \11846_b1 , \11712_b1 , \11717_b1 );
not ( \11717_b1 , w_30228 );
and ( \11846_b0 , \11712_b0 , w_30229 );
and ( w_30228 , w_30229 , \11717_b0 );
or ( \11847_b1 , \11708_b1 , \11717_b1 );
not ( \11717_b1 , w_30230 );
and ( \11847_b0 , \11708_b0 , w_30231 );
and ( w_30230 , w_30231 , \11717_b0 );
or ( \11849_b1 , \11696_b1 , \11700_b1 );
not ( \11700_b1 , w_30232 );
and ( \11849_b0 , \11696_b0 , w_30233 );
and ( w_30232 , w_30233 , \11700_b0 );
or ( \11850_b1 , \11700_b1 , \11705_b1 );
not ( \11705_b1 , w_30234 );
and ( \11850_b0 , \11700_b0 , w_30235 );
and ( w_30234 , w_30235 , \11705_b0 );
or ( \11851_b1 , \11696_b1 , \11705_b1 );
not ( \11705_b1 , w_30236 );
and ( \11851_b0 , \11696_b0 , w_30237 );
and ( w_30236 , w_30237 , \11705_b0 );
or ( \11853_b1 , \11848_b1 , \11852_b1 );
xor ( \11853_b0 , \11848_b0 , w_30238 );
not ( w_30238 , w_30239 );
and ( w_30239 , \11852_b1 , \11852_b0 );
or ( \11854_b1 , \11682_b1 , \11686_b1 );
not ( \11686_b1 , w_30240 );
and ( \11854_b0 , \11682_b0 , w_30241 );
and ( w_30240 , w_30241 , \11686_b0 );
or ( \11855_b1 , \11686_b1 , \11691_b1 );
not ( \11691_b1 , w_30242 );
and ( \11855_b0 , \11686_b0 , w_30243 );
and ( w_30242 , w_30243 , \11691_b0 );
or ( \11856_b1 , \11682_b1 , \11691_b1 );
not ( \11691_b1 , w_30244 );
and ( \11856_b0 , \11682_b0 , w_30245 );
and ( w_30244 , w_30245 , \11691_b0 );
or ( \11858_b1 , \11853_b1 , \11857_b1 );
xor ( \11858_b0 , \11853_b0 , w_30246 );
not ( w_30246 , w_30247 );
and ( w_30247 , \11857_b1 , \11857_b0 );
or ( \11859_b1 , \11844_b1 , \11858_b1 );
xor ( \11859_b0 , \11844_b0 , w_30248 );
not ( w_30248 , w_30249 );
and ( w_30249 , \11858_b1 , \11858_b0 );
or ( \11860_b1 , \11692_b1 , \11706_b1 );
not ( \11706_b1 , w_30250 );
and ( \11860_b0 , \11692_b0 , w_30251 );
and ( w_30250 , w_30251 , \11706_b0 );
or ( \11861_b1 , \11706_b1 , \11718_b1 );
not ( \11718_b1 , w_30252 );
and ( \11861_b0 , \11706_b0 , w_30253 );
and ( w_30252 , w_30253 , \11718_b0 );
or ( \11862_b1 , \11692_b1 , \11718_b1 );
not ( \11718_b1 , w_30254 );
and ( \11862_b0 , \11692_b0 , w_30255 );
and ( w_30254 , w_30255 , \11718_b0 );
or ( \11864_b1 , \5737_b1 , \7203_b1 );
not ( \7203_b1 , w_30256 );
and ( \11864_b0 , \5737_b0 , w_30257 );
and ( w_30256 , w_30257 , \7203_b0 );
buf ( \11865_b1 , \11864_b1 );
not ( \11865_b1 , w_30258 );
not ( \11865_b0 , w_30259 );
and ( w_30258 , w_30259 , \11864_b0 );
or ( \11866_b1 , \11865_b1 , w_30260 );
xor ( \11866_b0 , \11865_b0 , w_30262 );
not ( w_30262 , w_30263 );
and ( w_30263 , w_30260 , w_30261 );
buf ( w_30260 , \6824_b1 );
not ( w_30260 , w_30264 );
not ( w_30261 , w_30265 );
and ( w_30264 , w_30265 , \6824_b0 );
or ( \11867_b1 , \6062_b1 , \11866_b1 );
xor ( \11867_b0 , \6062_b0 , w_30266 );
not ( w_30266 , w_30267 );
and ( w_30267 , \11866_b1 , \11866_b0 );
or ( \11868_b1 , \5758_b1 , \5750_b1 );
not ( \5750_b1 , w_30268 );
and ( \11868_b0 , \5758_b0 , w_30269 );
and ( w_30268 , w_30269 , \5750_b0 );
or ( \11869_b1 , \5770_b1 , \5748_b1 );
not ( \5748_b1 , w_30270 );
and ( \11869_b0 , \5770_b0 , w_30271 );
and ( w_30270 , w_30271 , \5748_b0 );
or ( \11870_b1 , \11868_b1 , w_30273 );
not ( w_30273 , w_30274 );
and ( \11870_b0 , \11868_b0 , w_30275 );
and ( w_30274 ,  , w_30275 );
buf ( w_30273 , \11869_b1 );
not ( w_30273 , w_30276 );
not (  , w_30277 );
and ( w_30276 , w_30277 , \11869_b0 );
or ( \11871_b1 , \11870_b1 , w_30278 );
xor ( \11871_b0 , \11870_b0 , w_30280 );
not ( w_30280 , w_30281 );
and ( w_30281 , w_30278 , w_30279 );
buf ( w_30278 , \5755_b1 );
not ( w_30278 , w_30282 );
not ( w_30279 , w_30283 );
and ( w_30282 , w_30283 , \5755_b0 );
or ( \11872_b1 , \11867_b1 , \11871_b1 );
xor ( \11872_b0 , \11867_b0 , w_30284 );
not ( w_30284 , w_30285 );
and ( w_30285 , \11871_b1 , \11871_b0 );
or ( \11873_b1 , \11863_b1 , \11872_b1 );
xor ( \11873_b0 , \11863_b0 , w_30286 );
not ( w_30286 , w_30287 );
and ( w_30287 , \11872_b1 , \11872_b0 );
or ( \11874_b1 , \5906_b1 , \5891_b1 );
not ( \5891_b1 , w_30288 );
and ( \11874_b0 , \5906_b0 , w_30289 );
and ( w_30288 , w_30289 , \5891_b0 );
or ( \11875_b1 , \5918_b1 , \5889_b1 );
not ( \5889_b1 , w_30290 );
and ( \11875_b0 , \5918_b0 , w_30291 );
and ( w_30290 , w_30291 , \5889_b0 );
or ( \11876_b1 , \11874_b1 , w_30293 );
not ( w_30293 , w_30294 );
and ( \11876_b0 , \11874_b0 , w_30295 );
and ( w_30294 ,  , w_30295 );
buf ( w_30293 , \11875_b1 );
not ( w_30293 , w_30296 );
not (  , w_30297 );
and ( w_30296 , w_30297 , \11875_b0 );
or ( \11877_b1 , \11876_b1 , w_30298 );
xor ( \11877_b0 , \11876_b0 , w_30300 );
not ( w_30300 , w_30301 );
and ( w_30301 , w_30298 , w_30299 );
buf ( w_30298 , \5898_b1 );
not ( w_30298 , w_30302 );
not ( w_30299 , w_30303 );
and ( w_30302 , w_30303 , \5898_b0 );
or ( \11878_b1 , \5925_b1 , \5916_b1 );
not ( \5916_b1 , w_30304 );
and ( \11878_b0 , \5925_b0 , w_30305 );
and ( w_30304 , w_30305 , \5916_b0 );
or ( \11879_b1 , \5937_b1 , \5914_b1 );
not ( \5914_b1 , w_30306 );
and ( \11879_b0 , \5937_b0 , w_30307 );
and ( w_30306 , w_30307 , \5914_b0 );
or ( \11880_b1 , \11878_b1 , w_30309 );
not ( w_30309 , w_30310 );
and ( \11880_b0 , \11878_b0 , w_30311 );
and ( w_30310 ,  , w_30311 );
buf ( w_30309 , \11879_b1 );
not ( w_30309 , w_30312 );
not (  , w_30313 );
and ( w_30312 , w_30313 , \11879_b0 );
or ( \11881_b1 , \11880_b1 , w_30314 );
xor ( \11881_b0 , \11880_b0 , w_30316 );
not ( w_30316 , w_30317 );
and ( w_30317 , w_30314 , w_30315 );
buf ( w_30314 , \5923_b1 );
not ( w_30314 , w_30318 );
not ( w_30315 , w_30319 );
and ( w_30318 , w_30319 , \5923_b0 );
or ( \11882_b1 , \11877_b1 , \11881_b1 );
xor ( \11882_b0 , \11877_b0 , w_30320 );
not ( w_30320 , w_30321 );
and ( w_30321 , \11881_b1 , \11881_b0 );
or ( \11883_b1 , \5945_b1 , \5935_b1 );
not ( \5935_b1 , w_30322 );
and ( \11883_b0 , \5945_b0 , w_30323 );
and ( w_30322 , w_30323 , \5935_b0 );
or ( \11884_b1 , \5957_b1 , \5933_b1 );
not ( \5933_b1 , w_30324 );
and ( \11884_b0 , \5957_b0 , w_30325 );
and ( w_30324 , w_30325 , \5933_b0 );
or ( \11885_b1 , \11883_b1 , w_30327 );
not ( w_30327 , w_30328 );
and ( \11885_b0 , \11883_b0 , w_30329 );
and ( w_30328 ,  , w_30329 );
buf ( w_30327 , \11884_b1 );
not ( w_30327 , w_30330 );
not (  , w_30331 );
and ( w_30330 , w_30331 , \11884_b0 );
or ( \11886_b1 , \11885_b1 , w_30332 );
xor ( \11886_b0 , \11885_b0 , w_30334 );
not ( w_30334 , w_30335 );
and ( w_30335 , w_30332 , w_30333 );
buf ( w_30332 , \5942_b1 );
not ( w_30332 , w_30336 );
not ( w_30333 , w_30337 );
and ( w_30336 , w_30337 , \5942_b0 );
or ( \11887_b1 , \11882_b1 , \11886_b1 );
xor ( \11887_b0 , \11882_b0 , w_30338 );
not ( w_30338 , w_30339 );
and ( w_30339 , \11886_b1 , \11886_b0 );
or ( \11888_b1 , \5842_b1 , \5829_b1 );
not ( \5829_b1 , w_30340 );
and ( \11888_b0 , \5842_b0 , w_30341 );
and ( w_30340 , w_30341 , \5829_b0 );
or ( \11889_b1 , \5854_b1 , \5827_b1 );
not ( \5827_b1 , w_30342 );
and ( \11889_b0 , \5854_b0 , w_30343 );
and ( w_30342 , w_30343 , \5827_b0 );
or ( \11890_b1 , \11888_b1 , w_30345 );
not ( w_30345 , w_30346 );
and ( \11890_b0 , \11888_b0 , w_30347 );
and ( w_30346 ,  , w_30347 );
buf ( w_30345 , \11889_b1 );
not ( w_30345 , w_30348 );
not (  , w_30349 );
and ( w_30348 , w_30349 , \11889_b0 );
or ( \11891_b1 , \11890_b1 , w_30350 );
xor ( \11891_b0 , \11890_b0 , w_30352 );
not ( w_30352 , w_30353 );
and ( w_30353 , w_30350 , w_30351 );
buf ( w_30350 , \5836_b1 );
not ( w_30350 , w_30354 );
not ( w_30351 , w_30355 );
and ( w_30354 , w_30355 , \5836_b0 );
or ( \11892_b1 , \5861_b1 , \5852_b1 );
not ( \5852_b1 , w_30356 );
and ( \11892_b0 , \5861_b0 , w_30357 );
and ( w_30356 , w_30357 , \5852_b0 );
or ( \11893_b1 , \5873_b1 , \5850_b1 );
not ( \5850_b1 , w_30358 );
and ( \11893_b0 , \5873_b0 , w_30359 );
and ( w_30358 , w_30359 , \5850_b0 );
or ( \11894_b1 , \11892_b1 , w_30361 );
not ( w_30361 , w_30362 );
and ( \11894_b0 , \11892_b0 , w_30363 );
and ( w_30362 ,  , w_30363 );
buf ( w_30361 , \11893_b1 );
not ( w_30361 , w_30364 );
not (  , w_30365 );
and ( w_30364 , w_30365 , \11893_b0 );
or ( \11895_b1 , \11894_b1 , w_30366 );
xor ( \11895_b0 , \11894_b0 , w_30368 );
not ( w_30368 , w_30369 );
and ( w_30369 , w_30366 , w_30367 );
buf ( w_30366 , \5859_b1 );
not ( w_30366 , w_30370 );
not ( w_30367 , w_30371 );
and ( w_30370 , w_30371 , \5859_b0 );
or ( \11896_b1 , \11891_b1 , \11895_b1 );
xor ( \11896_b0 , \11891_b0 , w_30372 );
not ( w_30372 , w_30373 );
and ( w_30373 , \11895_b1 , \11895_b0 );
or ( \11897_b1 , \5881_b1 , \5871_b1 );
not ( \5871_b1 , w_30374 );
and ( \11897_b0 , \5881_b0 , w_30375 );
and ( w_30374 , w_30375 , \5871_b0 );
or ( \11898_b1 , \5893_b1 , \5869_b1 );
not ( \5869_b1 , w_30376 );
and ( \11898_b0 , \5893_b0 , w_30377 );
and ( w_30376 , w_30377 , \5869_b0 );
or ( \11899_b1 , \11897_b1 , w_30379 );
not ( w_30379 , w_30380 );
and ( \11899_b0 , \11897_b0 , w_30381 );
and ( w_30380 ,  , w_30381 );
buf ( w_30379 , \11898_b1 );
not ( w_30379 , w_30382 );
not (  , w_30383 );
and ( w_30382 , w_30383 , \11898_b0 );
or ( \11900_b1 , \11899_b1 , w_30384 );
xor ( \11900_b0 , \11899_b0 , w_30386 );
not ( w_30386 , w_30387 );
and ( w_30387 , w_30384 , w_30385 );
buf ( w_30384 , \5878_b1 );
not ( w_30384 , w_30388 );
not ( w_30385 , w_30389 );
and ( w_30388 , w_30389 , \5878_b0 );
or ( \11901_b1 , \11896_b1 , \11900_b1 );
xor ( \11901_b0 , \11896_b0 , w_30390 );
not ( w_30390 , w_30391 );
and ( w_30391 , \11900_b1 , \11900_b0 );
or ( \11902_b1 , \11887_b1 , \11901_b1 );
xor ( \11902_b0 , \11887_b0 , w_30392 );
not ( w_30392 , w_30393 );
and ( w_30393 , \11901_b1 , \11901_b0 );
or ( \11903_b1 , \5780_b1 , \5768_b1 );
not ( \5768_b1 , w_30394 );
and ( \11903_b0 , \5780_b0 , w_30395 );
and ( w_30394 , w_30395 , \5768_b0 );
or ( \11904_b1 , \5792_b1 , \5766_b1 );
not ( \5766_b1 , w_30396 );
and ( \11904_b0 , \5792_b0 , w_30397 );
and ( w_30396 , w_30397 , \5766_b0 );
or ( \11905_b1 , \11903_b1 , w_30399 );
not ( w_30399 , w_30400 );
and ( \11905_b0 , \11903_b0 , w_30401 );
and ( w_30400 ,  , w_30401 );
buf ( w_30399 , \11904_b1 );
not ( w_30399 , w_30402 );
not (  , w_30403 );
and ( w_30402 , w_30403 , \11904_b0 );
or ( \11906_b1 , \11905_b1 , w_30404 );
xor ( \11906_b0 , \11905_b0 , w_30406 );
not ( w_30406 , w_30407 );
and ( w_30407 , w_30404 , w_30405 );
buf ( w_30404 , \5775_b1 );
not ( w_30404 , w_30408 );
not ( w_30405 , w_30409 );
and ( w_30408 , w_30409 , \5775_b0 );
or ( \11907_b1 , \5799_b1 , \5790_b1 );
not ( \5790_b1 , w_30410 );
and ( \11907_b0 , \5799_b0 , w_30411 );
and ( w_30410 , w_30411 , \5790_b0 );
or ( \11908_b1 , \5811_b1 , \5788_b1 );
not ( \5788_b1 , w_30412 );
and ( \11908_b0 , \5811_b0 , w_30413 );
and ( w_30412 , w_30413 , \5788_b0 );
or ( \11909_b1 , \11907_b1 , w_30415 );
not ( w_30415 , w_30416 );
and ( \11909_b0 , \11907_b0 , w_30417 );
and ( w_30416 ,  , w_30417 );
buf ( w_30415 , \11908_b1 );
not ( w_30415 , w_30418 );
not (  , w_30419 );
and ( w_30418 , w_30419 , \11908_b0 );
or ( \11910_b1 , \11909_b1 , w_30420 );
xor ( \11910_b0 , \11909_b0 , w_30422 );
not ( w_30422 , w_30423 );
and ( w_30423 , w_30420 , w_30421 );
buf ( w_30420 , \5797_b1 );
not ( w_30420 , w_30424 );
not ( w_30421 , w_30425 );
and ( w_30424 , w_30425 , \5797_b0 );
or ( \11911_b1 , \11906_b1 , \11910_b1 );
xor ( \11911_b0 , \11906_b0 , w_30426 );
not ( w_30426 , w_30427 );
and ( w_30427 , \11910_b1 , \11910_b0 );
or ( \11912_b1 , \5819_b1 , \5809_b1 );
not ( \5809_b1 , w_30428 );
and ( \11912_b0 , \5819_b0 , w_30429 );
and ( w_30428 , w_30429 , \5809_b0 );
or ( \11913_b1 , \5831_b1 , \5807_b1 );
not ( \5807_b1 , w_30430 );
and ( \11913_b0 , \5831_b0 , w_30431 );
and ( w_30430 , w_30431 , \5807_b0 );
or ( \11914_b1 , \11912_b1 , w_30433 );
not ( w_30433 , w_30434 );
and ( \11914_b0 , \11912_b0 , w_30435 );
and ( w_30434 ,  , w_30435 );
buf ( w_30433 , \11913_b1 );
not ( w_30433 , w_30436 );
not (  , w_30437 );
and ( w_30436 , w_30437 , \11913_b0 );
or ( \11915_b1 , \11914_b1 , w_30438 );
xor ( \11915_b0 , \11914_b0 , w_30440 );
not ( w_30440 , w_30441 );
and ( w_30441 , w_30438 , w_30439 );
buf ( w_30438 , \5816_b1 );
not ( w_30438 , w_30442 );
not ( w_30439 , w_30443 );
and ( w_30442 , w_30443 , \5816_b0 );
or ( \11916_b1 , \11911_b1 , \11915_b1 );
xor ( \11916_b0 , \11911_b0 , w_30444 );
not ( w_30444 , w_30445 );
and ( w_30445 , \11915_b1 , \11915_b0 );
or ( \11917_b1 , \11902_b1 , \11916_b1 );
xor ( \11917_b0 , \11902_b0 , w_30446 );
not ( w_30446 , w_30447 );
and ( w_30447 , \11916_b1 , \11916_b0 );
or ( \11918_b1 , \11873_b1 , \11917_b1 );
xor ( \11918_b0 , \11873_b0 , w_30448 );
not ( w_30448 , w_30449 );
and ( w_30449 , \11917_b1 , \11917_b0 );
or ( \11919_b1 , \11859_b1 , \11918_b1 );
xor ( \11919_b0 , \11859_b0 , w_30450 );
not ( w_30450 , w_30451 );
and ( w_30451 , \11918_b1 , \11918_b0 );
or ( \11920_b1 , \11663_b1 , \11667_b1 );
not ( \11667_b1 , w_30452 );
and ( \11920_b0 , \11663_b0 , w_30453 );
and ( w_30452 , w_30453 , \11667_b0 );
or ( \11921_b1 , \11667_b1 , \11672_b1 );
not ( \11672_b1 , w_30454 );
and ( \11921_b0 , \11667_b0 , w_30455 );
and ( w_30454 , w_30455 , \11672_b0 );
or ( \11922_b1 , \11663_b1 , \11672_b1 );
not ( \11672_b1 , w_30456 );
and ( \11922_b0 , \11663_b0 , w_30457 );
and ( w_30456 , w_30457 , \11672_b0 );
or ( \11924_b1 , \11649_b1 , \11653_b1 );
not ( \11653_b1 , w_30458 );
and ( \11924_b0 , \11649_b0 , w_30459 );
and ( w_30458 , w_30459 , \11653_b0 );
or ( \11925_b1 , \11653_b1 , \11658_b1 );
not ( \11658_b1 , w_30460 );
and ( \11925_b0 , \11653_b0 , w_30461 );
and ( w_30460 , w_30461 , \11658_b0 );
or ( \11926_b1 , \11649_b1 , \11658_b1 );
not ( \11658_b1 , w_30462 );
and ( \11926_b0 , \11649_b0 , w_30463 );
and ( w_30462 , w_30463 , \11658_b0 );
or ( \11928_b1 , \11923_b1 , \11927_b1 );
xor ( \11928_b0 , \11923_b0 , w_30464 );
not ( w_30464 , w_30465 );
and ( w_30465 , \11927_b1 , \11927_b0 );
or ( \11929_b1 , \11729_b1 , \11743_b1 );
not ( \11743_b1 , w_30466 );
and ( \11929_b0 , \11729_b0 , w_30467 );
and ( w_30466 , w_30467 , \11743_b0 );
or ( \11930_b1 , \11743_b1 , \11758_b1 );
not ( \11758_b1 , w_30468 );
and ( \11930_b0 , \11743_b0 , w_30469 );
and ( w_30468 , w_30469 , \11758_b0 );
or ( \11931_b1 , \11729_b1 , \11758_b1 );
not ( \11758_b1 , w_30470 );
and ( \11931_b0 , \11729_b0 , w_30471 );
and ( w_30470 , w_30471 , \11758_b0 );
or ( \11933_b1 , \11928_b1 , \11932_b1 );
xor ( \11933_b0 , \11928_b0 , w_30472 );
not ( w_30472 , w_30473 );
and ( w_30473 , \11932_b1 , \11932_b0 );
or ( \11934_b1 , \11919_b1 , \11933_b1 );
xor ( \11934_b0 , \11919_b0 , w_30474 );
not ( w_30474 , w_30475 );
and ( w_30475 , \11933_b1 , \11933_b0 );
or ( \11935_b1 , \11805_b1 , \11934_b1 );
xor ( \11935_b0 , \11805_b0 , w_30476 );
not ( w_30476 , w_30477 );
and ( w_30477 , \11934_b1 , \11934_b0 );
or ( \11936_b1 , \11796_b1 , \11935_b1 );
xor ( \11936_b0 , \11796_b0 , w_30478 );
not ( w_30478 , w_30479 );
and ( w_30479 , \11935_b1 , \11935_b0 );
or ( \11937_b1 , \11621_b1 , \11635_b1 );
not ( \11635_b1 , w_30480 );
and ( \11937_b0 , \11621_b0 , w_30481 );
and ( w_30480 , w_30481 , \11635_b0 );
or ( \11938_b1 , \11635_b1 , \11774_b1 );
not ( \11774_b1 , w_30482 );
and ( \11938_b0 , \11635_b0 , w_30483 );
and ( w_30482 , w_30483 , \11774_b0 );
or ( \11939_b1 , \11621_b1 , \11774_b1 );
not ( \11774_b1 , w_30484 );
and ( \11939_b0 , \11621_b0 , w_30485 );
and ( w_30484 , w_30485 , \11774_b0 );
or ( \11941_b1 , \11936_b1 , w_30487 );
not ( w_30487 , w_30488 );
and ( \11941_b0 , \11936_b0 , w_30489 );
and ( w_30488 ,  , w_30489 );
buf ( w_30487 , \11940_b1 );
not ( w_30487 , w_30490 );
not (  , w_30491 );
and ( w_30490 , w_30491 , \11940_b0 );
or ( \11942_b1 , \11780_b1 , w_30493 );
not ( w_30493 , w_30494 );
and ( \11942_b0 , \11780_b0 , w_30495 );
and ( w_30494 ,  , w_30495 );
buf ( w_30493 , \11941_b1 );
not ( w_30493 , w_30496 );
not (  , w_30497 );
and ( w_30496 , w_30497 , \11941_b0 );
or ( \11943_b1 , \11800_b1 , \11804_b1 );
not ( \11804_b1 , w_30498 );
and ( \11943_b0 , \11800_b0 , w_30499 );
and ( w_30498 , w_30499 , \11804_b0 );
or ( \11944_b1 , \11804_b1 , \11934_b1 );
not ( \11934_b1 , w_30500 );
and ( \11944_b0 , \11804_b0 , w_30501 );
and ( w_30500 , w_30501 , \11934_b0 );
or ( \11945_b1 , \11800_b1 , \11934_b1 );
not ( \11934_b1 , w_30502 );
and ( \11945_b0 , \11800_b0 , w_30503 );
and ( w_30502 , w_30503 , \11934_b0 );
or ( \11947_b1 , \11923_b1 , \11927_b1 );
not ( \11927_b1 , w_30504 );
and ( \11947_b0 , \11923_b0 , w_30505 );
and ( w_30504 , w_30505 , \11927_b0 );
or ( \11948_b1 , \11927_b1 , \11932_b1 );
not ( \11932_b1 , w_30506 );
and ( \11948_b0 , \11927_b0 , w_30507 );
and ( w_30506 , w_30507 , \11932_b0 );
or ( \11949_b1 , \11923_b1 , \11932_b1 );
not ( \11932_b1 , w_30508 );
and ( \11949_b0 , \11923_b0 , w_30509 );
and ( w_30508 , w_30509 , \11932_b0 );
or ( \11951_b1 , \11863_b1 , \11872_b1 );
not ( \11872_b1 , w_30510 );
and ( \11951_b0 , \11863_b0 , w_30511 );
and ( w_30510 , w_30511 , \11872_b0 );
or ( \11952_b1 , \11872_b1 , \11917_b1 );
not ( \11917_b1 , w_30512 );
and ( \11952_b0 , \11872_b0 , w_30513 );
and ( w_30512 , w_30513 , \11917_b0 );
or ( \11953_b1 , \11863_b1 , \11917_b1 );
not ( \11917_b1 , w_30514 );
and ( \11953_b0 , \11863_b0 , w_30515 );
and ( w_30514 , w_30515 , \11917_b0 );
or ( \11955_b1 , \11950_b1 , \11954_b1 );
xor ( \11955_b0 , \11950_b0 , w_30516 );
not ( w_30516 , w_30517 );
and ( w_30517 , \11954_b1 , \11954_b0 );
or ( \11956_b1 , \11832_b1 , \11843_b1 );
not ( \11843_b1 , w_30518 );
and ( \11956_b0 , \11832_b0 , w_30519 );
and ( w_30518 , w_30519 , \11843_b0 );
or ( \11957_b1 , \11843_b1 , \11858_b1 );
not ( \11858_b1 , w_30520 );
and ( \11957_b0 , \11843_b0 , w_30521 );
and ( w_30520 , w_30521 , \11858_b0 );
or ( \11958_b1 , \11832_b1 , \11858_b1 );
not ( \11858_b1 , w_30522 );
and ( \11958_b0 , \11832_b0 , w_30523 );
and ( w_30522 , w_30523 , \11858_b0 );
or ( \11960_b1 , \11955_b1 , \11959_b1 );
xor ( \11960_b0 , \11955_b0 , w_30524 );
not ( w_30524 , w_30525 );
and ( w_30525 , \11959_b1 , \11959_b0 );
or ( \11961_b1 , \11946_b1 , \11960_b1 );
xor ( \11961_b0 , \11946_b0 , w_30526 );
not ( w_30526 , w_30527 );
and ( w_30527 , \11960_b1 , \11960_b0 );
or ( \11962_b1 , \11788_b1 , \11792_b1 );
not ( \11792_b1 , w_30528 );
and ( \11962_b0 , \11788_b0 , w_30529 );
and ( w_30528 , w_30529 , \11792_b0 );
or ( \11963_b1 , \11792_b1 , \11794_b1 );
not ( \11794_b1 , w_30530 );
and ( \11963_b0 , \11792_b0 , w_30531 );
and ( w_30530 , w_30531 , \11794_b0 );
or ( \11964_b1 , \11788_b1 , \11794_b1 );
not ( \11794_b1 , w_30532 );
and ( \11964_b0 , \11788_b0 , w_30533 );
and ( w_30532 , w_30533 , \11794_b0 );
or ( \11966_b1 , \11859_b1 , \11918_b1 );
not ( \11918_b1 , w_30534 );
and ( \11966_b0 , \11859_b0 , w_30535 );
and ( w_30534 , w_30535 , \11918_b0 );
or ( \11967_b1 , \11918_b1 , \11933_b1 );
not ( \11933_b1 , w_30536 );
and ( \11967_b0 , \11918_b0 , w_30537 );
and ( w_30536 , w_30537 , \11933_b0 );
or ( \11968_b1 , \11859_b1 , \11933_b1 );
not ( \11933_b1 , w_30538 );
and ( \11968_b0 , \11859_b0 , w_30539 );
and ( w_30538 , w_30539 , \11933_b0 );
or ( \11970_b1 , \11965_b1 , \11969_b1 );
xor ( \11970_b0 , \11965_b0 , w_30540 );
not ( w_30540 , w_30541 );
and ( w_30541 , \11969_b1 , \11969_b0 );
or ( \11971_b1 , \11877_b1 , \11881_b1 );
not ( \11881_b1 , w_30542 );
and ( \11971_b0 , \11877_b0 , w_30543 );
and ( w_30542 , w_30543 , \11881_b0 );
or ( \11972_b1 , \11881_b1 , \11886_b1 );
not ( \11886_b1 , w_30544 );
and ( \11972_b0 , \11881_b0 , w_30545 );
and ( w_30544 , w_30545 , \11886_b0 );
or ( \11973_b1 , \11877_b1 , \11886_b1 );
not ( \11886_b1 , w_30546 );
and ( \11973_b0 , \11877_b0 , w_30547 );
and ( w_30546 , w_30547 , \11886_b0 );
or ( \11975_b1 , \11821_b1 , \11825_b1 );
not ( \11825_b1 , w_30548 );
and ( \11975_b0 , \11821_b0 , w_30549 );
and ( w_30548 , w_30549 , \11825_b0 );
or ( \11976_b1 , \11825_b1 , \11830_b1 );
not ( \11830_b1 , w_30550 );
and ( \11976_b0 , \11825_b0 , w_30551 );
and ( w_30550 , w_30551 , \11830_b0 );
or ( \11977_b1 , \11821_b1 , \11830_b1 );
not ( \11830_b1 , w_30552 );
and ( \11977_b0 , \11821_b0 , w_30553 );
and ( w_30552 , w_30553 , \11830_b0 );
or ( \11979_b1 , \11974_b1 , \11978_b1 );
xor ( \11979_b0 , \11974_b0 , w_30554 );
not ( w_30554 , w_30555 );
and ( w_30555 , \11978_b1 , \11978_b0 );
or ( \11980_b1 , \11809_b1 , \11813_b1 );
not ( \11813_b1 , w_30556 );
and ( \11980_b0 , \11809_b0 , w_30557 );
and ( w_30556 , w_30557 , \11813_b0 );
or ( \11981_b1 , \11813_b1 , \11816_b1 );
not ( \11816_b1 , w_30558 );
and ( \11981_b0 , \11813_b0 , w_30559 );
and ( w_30558 , w_30559 , \11816_b0 );
or ( \11982_b1 , \11809_b1 , \11816_b1 );
not ( \11816_b1 , w_30560 );
and ( \11982_b0 , \11809_b0 , w_30561 );
and ( w_30560 , w_30561 , \11816_b0 );
or ( \11984_b1 , \11979_b1 , \11983_b1 );
xor ( \11984_b0 , \11979_b0 , w_30562 );
not ( w_30562 , w_30563 );
and ( w_30563 , \11983_b1 , \11983_b0 );
or ( \11985_b1 , \6062_b1 , \11866_b1 );
not ( \11866_b1 , w_30564 );
and ( \11985_b0 , \6062_b0 , w_30565 );
and ( w_30564 , w_30565 , \11866_b0 );
or ( \11986_b1 , \11866_b1 , \11871_b1 );
not ( \11871_b1 , w_30566 );
and ( \11986_b0 , \11866_b0 , w_30567 );
and ( w_30566 , w_30567 , \11871_b0 );
or ( \11987_b1 , \6062_b1 , \11871_b1 );
not ( \11871_b1 , w_30568 );
and ( \11987_b0 , \6062_b0 , w_30569 );
and ( w_30568 , w_30569 , \11871_b0 );
or ( \11989_b1 , \11906_b1 , \11910_b1 );
not ( \11910_b1 , w_30570 );
and ( \11989_b0 , \11906_b0 , w_30571 );
and ( w_30570 , w_30571 , \11910_b0 );
or ( \11990_b1 , \11910_b1 , \11915_b1 );
not ( \11915_b1 , w_30572 );
and ( \11990_b0 , \11910_b0 , w_30573 );
and ( w_30572 , w_30573 , \11915_b0 );
or ( \11991_b1 , \11906_b1 , \11915_b1 );
not ( \11915_b1 , w_30574 );
and ( \11991_b0 , \11906_b0 , w_30575 );
and ( w_30574 , w_30575 , \11915_b0 );
or ( \11993_b1 , \11988_b1 , \11992_b1 );
xor ( \11993_b0 , \11988_b0 , w_30576 );
not ( w_30576 , w_30577 );
and ( w_30577 , \11992_b1 , \11992_b0 );
or ( \11994_b1 , \11891_b1 , \11895_b1 );
not ( \11895_b1 , w_30578 );
and ( \11994_b0 , \11891_b0 , w_30579 );
and ( w_30578 , w_30579 , \11895_b0 );
or ( \11995_b1 , \11895_b1 , \11900_b1 );
not ( \11900_b1 , w_30580 );
and ( \11995_b0 , \11895_b0 , w_30581 );
and ( w_30580 , w_30581 , \11900_b0 );
or ( \11996_b1 , \11891_b1 , \11900_b1 );
not ( \11900_b1 , w_30582 );
and ( \11996_b0 , \11891_b0 , w_30583 );
and ( w_30582 , w_30583 , \11900_b0 );
or ( \11998_b1 , \11993_b1 , \11997_b1 );
xor ( \11998_b0 , \11993_b0 , w_30584 );
not ( w_30584 , w_30585 );
and ( w_30585 , \11997_b1 , \11997_b0 );
or ( \11999_b1 , \11984_b1 , \11998_b1 );
xor ( \11999_b0 , \11984_b0 , w_30586 );
not ( w_30586 , w_30587 );
and ( w_30587 , \11998_b1 , \11998_b0 );
or ( \12000_b1 , \11887_b1 , \11901_b1 );
not ( \11901_b1 , w_30588 );
and ( \12000_b0 , \11887_b0 , w_30589 );
and ( w_30588 , w_30589 , \11901_b0 );
or ( \12001_b1 , \11901_b1 , \11916_b1 );
not ( \11916_b1 , w_30590 );
and ( \12001_b0 , \11901_b0 , w_30591 );
and ( w_30590 , w_30591 , \11916_b0 );
or ( \12002_b1 , \11887_b1 , \11916_b1 );
not ( \11916_b1 , w_30592 );
and ( \12002_b0 , \11887_b0 , w_30593 );
and ( w_30592 , w_30593 , \11916_b0 );
or ( \12004_b1 , \6858_b1 , \6862_b1 );
xor ( \12004_b0 , \6858_b0 , w_30594 );
not ( w_30594 , w_30595 );
and ( w_30595 , \6862_b1 , \6862_b0 );
or ( \12005_b1 , \12004_b1 , \6867_b1 );
xor ( \12005_b0 , \12004_b0 , w_30596 );
not ( w_30596 , w_30597 );
and ( w_30597 , \6867_b1 , \6867_b0 );
or ( \12006_b1 , \6841_b1 , \6845_b1 );
xor ( \12006_b0 , \6841_b0 , w_30598 );
not ( w_30598 , w_30599 );
and ( w_30599 , \6845_b1 , \6845_b0 );
or ( \12007_b1 , \12006_b1 , \6850_b1 );
xor ( \12007_b0 , \12006_b0 , w_30600 );
not ( w_30600 , w_30601 );
and ( w_30601 , \6850_b1 , \6850_b0 );
or ( \12008_b1 , \12005_b1 , \12007_b1 );
xor ( \12008_b0 , \12005_b0 , w_30602 );
not ( w_30602 , w_30603 );
and ( w_30603 , \12007_b1 , \12007_b0 );
or ( \12009_b1 , \6825_b1 , \6829_b1 );
xor ( \12009_b0 , \6825_b0 , w_30604 );
not ( w_30604 , w_30605 );
and ( w_30605 , \6829_b1 , \6829_b0 );
or ( \12010_b1 , \12009_b1 , \6834_b1 );
xor ( \12010_b0 , \12009_b0 , w_30606 );
not ( w_30606 , w_30607 );
and ( w_30607 , \6834_b1 , \6834_b0 );
or ( \12011_b1 , \12008_b1 , \12010_b1 );
xor ( \12011_b0 , \12008_b0 , w_30608 );
not ( w_30608 , w_30609 );
and ( w_30609 , \12010_b1 , \12010_b0 );
or ( \12012_b1 , \12003_b1 , \12011_b1 );
xor ( \12012_b0 , \12003_b0 , w_30610 );
not ( w_30610 , w_30611 );
and ( w_30611 , \12011_b1 , \12011_b0 );
or ( \12013_b1 , \6910_b1 , \6914_b1 );
xor ( \12013_b0 , \6910_b0 , w_30612 );
not ( w_30612 , w_30613 );
and ( w_30613 , \6914_b1 , \6914_b0 );
or ( \12014_b1 , \6893_b1 , \6897_b1 );
xor ( \12014_b0 , \6893_b0 , w_30614 );
not ( w_30614 , w_30615 );
and ( w_30615 , \6897_b1 , \6897_b0 );
or ( \12015_b1 , \12014_b1 , \6902_b1 );
xor ( \12015_b0 , \12014_b0 , w_30616 );
not ( w_30616 , w_30617 );
and ( w_30617 , \6902_b1 , \6902_b0 );
or ( \12016_b1 , \12013_b1 , \12015_b1 );
xor ( \12016_b0 , \12013_b0 , w_30618 );
not ( w_30618 , w_30619 );
and ( w_30619 , \12015_b1 , \12015_b0 );
or ( \12017_b1 , \6877_b1 , \6881_b1 );
xor ( \12017_b0 , \6877_b0 , w_30620 );
not ( w_30620 , w_30621 );
and ( w_30621 , \6881_b1 , \6881_b0 );
or ( \12018_b1 , \12017_b1 , \6886_b1 );
xor ( \12018_b0 , \12017_b0 , w_30622 );
not ( w_30622 , w_30623 );
and ( w_30623 , \6886_b1 , \6886_b0 );
or ( \12019_b1 , \12016_b1 , \12018_b1 );
xor ( \12019_b0 , \12016_b0 , w_30624 );
not ( w_30624 , w_30625 );
and ( w_30625 , \12018_b1 , \12018_b0 );
or ( \12020_b1 , \12012_b1 , \12019_b1 );
xor ( \12020_b0 , \12012_b0 , w_30626 );
not ( w_30626 , w_30627 );
and ( w_30627 , \12019_b1 , \12019_b0 );
or ( \12021_b1 , \11999_b1 , \12020_b1 );
xor ( \12021_b0 , \11999_b0 , w_30628 );
not ( w_30628 , w_30629 );
and ( w_30629 , \12020_b1 , \12020_b0 );
or ( \12022_b1 , \11848_b1 , \11852_b1 );
not ( \11852_b1 , w_30630 );
and ( \12022_b0 , \11848_b0 , w_30631 );
and ( w_30630 , w_30631 , \11852_b0 );
or ( \12023_b1 , \11852_b1 , \11857_b1 );
not ( \11857_b1 , w_30632 );
and ( \12023_b0 , \11852_b0 , w_30633 );
and ( w_30632 , w_30633 , \11857_b0 );
or ( \12024_b1 , \11848_b1 , \11857_b1 );
not ( \11857_b1 , w_30634 );
and ( \12024_b0 , \11848_b0 , w_30635 );
and ( w_30634 , w_30635 , \11857_b0 );
or ( \12026_b1 , \11836_b1 , \11840_b1 );
not ( \11840_b1 , w_30636 );
and ( \12026_b0 , \11836_b0 , w_30637 );
and ( w_30636 , w_30637 , \11840_b0 );
or ( \12027_b1 , \11840_b1 , \11842_b1 );
not ( \11842_b1 , w_30638 );
and ( \12027_b0 , \11840_b0 , w_30639 );
and ( w_30638 , w_30639 , \11842_b0 );
or ( \12028_b1 , \11836_b1 , \11842_b1 );
not ( \11842_b1 , w_30640 );
and ( \12028_b0 , \11836_b0 , w_30641 );
and ( w_30640 , w_30641 , \11842_b0 );
or ( \12030_b1 , \12025_b1 , \12029_b1 );
xor ( \12030_b0 , \12025_b0 , w_30642 );
not ( w_30642 , w_30643 );
and ( w_30643 , \12029_b1 , \12029_b0 );
or ( \12031_b1 , \11817_b1 , w_30644 );
or ( \12031_b0 , \11817_b0 , \11831_b0 );
not ( \11831_b0 , w_30645 );
and ( w_30645 , w_30644 , \11831_b1 );
or ( \12032_b1 , \12030_b1 , \12031_b1 );
xor ( \12032_b0 , \12030_b0 , w_30646 );
not ( w_30646 , w_30647 );
and ( w_30647 , \12031_b1 , \12031_b0 );
or ( \12033_b1 , \12021_b1 , \12032_b1 );
xor ( \12033_b0 , \12021_b0 , w_30648 );
not ( w_30648 , w_30649 );
and ( w_30649 , \12032_b1 , \12032_b0 );
or ( \12034_b1 , \11970_b1 , \12033_b1 );
xor ( \12034_b0 , \11970_b0 , w_30650 );
not ( w_30650 , w_30651 );
and ( w_30651 , \12033_b1 , \12033_b0 );
or ( \12035_b1 , \11961_b1 , \12034_b1 );
xor ( \12035_b0 , \11961_b0 , w_30652 );
not ( w_30652 , w_30653 );
and ( w_30653 , \12034_b1 , \12034_b0 );
or ( \12036_b1 , \11784_b1 , \11795_b1 );
not ( \11795_b1 , w_30654 );
and ( \12036_b0 , \11784_b0 , w_30655 );
and ( w_30654 , w_30655 , \11795_b0 );
or ( \12037_b1 , \11795_b1 , \11935_b1 );
not ( \11935_b1 , w_30656 );
and ( \12037_b0 , \11795_b0 , w_30657 );
and ( w_30656 , w_30657 , \11935_b0 );
or ( \12038_b1 , \11784_b1 , \11935_b1 );
not ( \11935_b1 , w_30658 );
and ( \12038_b0 , \11784_b0 , w_30659 );
and ( w_30658 , w_30659 , \11935_b0 );
or ( \12040_b1 , \12035_b1 , w_30661 );
not ( w_30661 , w_30662 );
and ( \12040_b0 , \12035_b0 , w_30663 );
and ( w_30662 ,  , w_30663 );
buf ( w_30661 , \12039_b1 );
not ( w_30661 , w_30664 );
not (  , w_30665 );
and ( w_30664 , w_30665 , \12039_b0 );
or ( \12041_b1 , \11965_b1 , \11969_b1 );
not ( \11969_b1 , w_30666 );
and ( \12041_b0 , \11965_b0 , w_30667 );
and ( w_30666 , w_30667 , \11969_b0 );
or ( \12042_b1 , \11969_b1 , \12033_b1 );
not ( \12033_b1 , w_30668 );
and ( \12042_b0 , \11969_b0 , w_30669 );
and ( w_30668 , w_30669 , \12033_b0 );
or ( \12043_b1 , \11965_b1 , \12033_b1 );
not ( \12033_b1 , w_30670 );
and ( \12043_b0 , \11965_b0 , w_30671 );
and ( w_30670 , w_30671 , \12033_b0 );
or ( \12045_b1 , \12025_b1 , \12029_b1 );
not ( \12029_b1 , w_30672 );
and ( \12045_b0 , \12025_b0 , w_30673 );
and ( w_30672 , w_30673 , \12029_b0 );
or ( \12046_b1 , \12029_b1 , \12031_b1 );
not ( \12031_b1 , w_30674 );
and ( \12046_b0 , \12029_b0 , w_30675 );
and ( w_30674 , w_30675 , \12031_b0 );
or ( \12047_b1 , \12025_b1 , \12031_b1 );
not ( \12031_b1 , w_30676 );
and ( \12047_b0 , \12025_b0 , w_30677 );
and ( w_30676 , w_30677 , \12031_b0 );
or ( \12049_b1 , \12003_b1 , \12011_b1 );
not ( \12011_b1 , w_30678 );
and ( \12049_b0 , \12003_b0 , w_30679 );
and ( w_30678 , w_30679 , \12011_b0 );
or ( \12050_b1 , \12011_b1 , \12019_b1 );
not ( \12019_b1 , w_30680 );
and ( \12050_b0 , \12011_b0 , w_30681 );
and ( w_30680 , w_30681 , \12019_b0 );
or ( \12051_b1 , \12003_b1 , \12019_b1 );
not ( \12019_b1 , w_30682 );
and ( \12051_b0 , \12003_b0 , w_30683 );
and ( w_30682 , w_30683 , \12019_b0 );
or ( \12053_b1 , \12048_b1 , \12052_b1 );
xor ( \12053_b0 , \12048_b0 , w_30684 );
not ( w_30684 , w_30685 );
and ( w_30685 , \12052_b1 , \12052_b0 );
or ( \12054_b1 , \11984_b1 , \11998_b1 );
not ( \11998_b1 , w_30686 );
and ( \12054_b0 , \11984_b0 , w_30687 );
and ( w_30686 , w_30687 , \11998_b0 );
or ( \12055_b1 , \12053_b1 , \12054_b1 );
xor ( \12055_b0 , \12053_b0 , w_30688 );
not ( w_30688 , w_30689 );
and ( w_30689 , \12054_b1 , \12054_b0 );
or ( \12056_b1 , \12044_b1 , \12055_b1 );
xor ( \12056_b0 , \12044_b0 , w_30690 );
not ( w_30690 , w_30691 );
and ( w_30691 , \12055_b1 , \12055_b0 );
or ( \12057_b1 , \11950_b1 , \11954_b1 );
not ( \11954_b1 , w_30692 );
and ( \12057_b0 , \11950_b0 , w_30693 );
and ( w_30692 , w_30693 , \11954_b0 );
or ( \12058_b1 , \11954_b1 , \11959_b1 );
not ( \11959_b1 , w_30694 );
and ( \12058_b0 , \11954_b0 , w_30695 );
and ( w_30694 , w_30695 , \11959_b0 );
or ( \12059_b1 , \11950_b1 , \11959_b1 );
not ( \11959_b1 , w_30696 );
and ( \12059_b0 , \11950_b0 , w_30697 );
and ( w_30696 , w_30697 , \11959_b0 );
or ( \12061_b1 , \11999_b1 , \12020_b1 );
not ( \12020_b1 , w_30698 );
and ( \12061_b0 , \11999_b0 , w_30699 );
and ( w_30698 , w_30699 , \12020_b0 );
or ( \12062_b1 , \12020_b1 , \12032_b1 );
not ( \12032_b1 , w_30700 );
and ( \12062_b0 , \12020_b0 , w_30701 );
and ( w_30700 , w_30701 , \12032_b0 );
or ( \12063_b1 , \11999_b1 , \12032_b1 );
not ( \12032_b1 , w_30702 );
and ( \12063_b0 , \11999_b0 , w_30703 );
and ( w_30702 , w_30703 , \12032_b0 );
or ( \12065_b1 , \12060_b1 , \12064_b1 );
xor ( \12065_b0 , \12060_b0 , w_30704 );
not ( w_30704 , w_30705 );
and ( w_30705 , \12064_b1 , \12064_b0 );
or ( \12066_b1 , \6921_b1 , w_30706 );
xor ( \12066_b0 , \6921_b0 , w_30708 );
not ( w_30708 , w_30709 );
and ( w_30709 , w_30706 , w_30707 );
buf ( w_30706 , \6923_b1 );
not ( w_30706 , w_30710 );
not ( w_30707 , w_30711 );
and ( w_30710 , w_30711 , \6923_b0 );
or ( \12067_b1 , \6889_b1 , \6905_b1 );
xor ( \12067_b0 , \6889_b0 , w_30712 );
not ( w_30712 , w_30713 );
and ( w_30713 , \6905_b1 , \6905_b0 );
or ( \12068_b1 , \12067_b1 , \6915_b1 );
xor ( \12068_b0 , \12067_b0 , w_30714 );
not ( w_30714 , w_30715 );
and ( w_30715 , \6915_b1 , \6915_b0 );
or ( \12069_b1 , \12066_b1 , \12068_b1 );
xor ( \12069_b0 , \12066_b0 , w_30716 );
not ( w_30716 , w_30717 );
and ( w_30717 , \12068_b1 , \12068_b0 );
or ( \12070_b1 , \6837_b1 , \6853_b1 );
xor ( \12070_b0 , \6837_b0 , w_30718 );
not ( w_30718 , w_30719 );
and ( w_30719 , \6853_b1 , \6853_b0 );
or ( \12071_b1 , \12070_b1 , \6870_b1 );
xor ( \12071_b0 , \12070_b0 , w_30720 );
not ( w_30720 , w_30721 );
and ( w_30721 , \6870_b1 , \6870_b0 );
or ( \12072_b1 , \12069_b1 , \12071_b1 );
xor ( \12072_b0 , \12069_b0 , w_30722 );
not ( w_30722 , w_30723 );
and ( w_30723 , \12071_b1 , \12071_b0 );
or ( \12073_b1 , \12005_b1 , \12007_b1 );
not ( \12007_b1 , w_30724 );
and ( \12073_b0 , \12005_b0 , w_30725 );
and ( w_30724 , w_30725 , \12007_b0 );
or ( \12074_b1 , \12007_b1 , \12010_b1 );
not ( \12010_b1 , w_30726 );
and ( \12074_b0 , \12007_b0 , w_30727 );
and ( w_30726 , w_30727 , \12010_b0 );
or ( \12075_b1 , \12005_b1 , \12010_b1 );
not ( \12010_b1 , w_30728 );
and ( \12075_b0 , \12005_b0 , w_30729 );
and ( w_30728 , w_30729 , \12010_b0 );
or ( \12077_b1 , \5736_b1 , \5756_b1 );
xor ( \12077_b0 , \5736_b0 , w_30730 );
not ( w_30730 , w_30731 );
and ( w_30731 , \5756_b1 , \5756_b0 );
or ( \12078_b1 , \12077_b1 , \5776_b1 );
xor ( \12078_b0 , \12077_b0 , w_30732 );
not ( w_30732 , w_30733 );
and ( w_30733 , \5776_b1 , \5776_b0 );
or ( \12079_b1 , \12076_b1 , \12078_b1 );
xor ( \12079_b0 , \12076_b0 , w_30734 );
not ( w_30734 , w_30735 );
and ( w_30735 , \12078_b1 , \12078_b0 );
or ( \12080_b1 , \6929_b1 , \6931_b1 );
xor ( \12080_b0 , \6929_b0 , w_30736 );
not ( w_30736 , w_30737 );
and ( w_30737 , \6931_b1 , \6931_b0 );
or ( \12081_b1 , \12080_b1 , \6934_b1 );
xor ( \12081_b0 , \12080_b0 , w_30738 );
not ( w_30738 , w_30739 );
and ( w_30739 , \6934_b1 , \6934_b0 );
or ( \12082_b1 , \12079_b1 , \12081_b1 );
xor ( \12082_b0 , \12079_b0 , w_30740 );
not ( w_30740 , w_30741 );
and ( w_30741 , \12081_b1 , \12081_b0 );
or ( \12083_b1 , \12072_b1 , \12082_b1 );
xor ( \12083_b0 , \12072_b0 , w_30742 );
not ( w_30742 , w_30743 );
and ( w_30743 , \12082_b1 , \12082_b0 );
or ( \12084_b1 , \11988_b1 , \11992_b1 );
not ( \11992_b1 , w_30744 );
and ( \12084_b0 , \11988_b0 , w_30745 );
and ( w_30744 , w_30745 , \11992_b0 );
or ( \12085_b1 , \11992_b1 , \11997_b1 );
not ( \11997_b1 , w_30746 );
and ( \12085_b0 , \11992_b0 , w_30747 );
and ( w_30746 , w_30747 , \11997_b0 );
or ( \12086_b1 , \11988_b1 , \11997_b1 );
not ( \11997_b1 , w_30748 );
and ( \12086_b0 , \11988_b0 , w_30749 );
and ( w_30748 , w_30749 , \11997_b0 );
or ( \12088_b1 , \11974_b1 , \11978_b1 );
not ( \11978_b1 , w_30750 );
and ( \12088_b0 , \11974_b0 , w_30751 );
and ( w_30750 , w_30751 , \11978_b0 );
or ( \12089_b1 , \11978_b1 , \11983_b1 );
not ( \11983_b1 , w_30752 );
and ( \12089_b0 , \11978_b0 , w_30753 );
and ( w_30752 , w_30753 , \11983_b0 );
or ( \12090_b1 , \11974_b1 , \11983_b1 );
not ( \11983_b1 , w_30754 );
and ( \12090_b0 , \11974_b0 , w_30755 );
and ( w_30754 , w_30755 , \11983_b0 );
or ( \12092_b1 , \12087_b1 , \12091_b1 );
xor ( \12092_b0 , \12087_b0 , w_30756 );
not ( w_30756 , w_30757 );
and ( w_30757 , \12091_b1 , \12091_b0 );
or ( \12093_b1 , \12013_b1 , \12015_b1 );
not ( \12015_b1 , w_30758 );
and ( \12093_b0 , \12013_b0 , w_30759 );
and ( w_30758 , w_30759 , \12015_b0 );
or ( \12094_b1 , \12015_b1 , \12018_b1 );
not ( \12018_b1 , w_30760 );
and ( \12094_b0 , \12015_b0 , w_30761 );
and ( w_30760 , w_30761 , \12018_b0 );
or ( \12095_b1 , \12013_b1 , \12018_b1 );
not ( \12018_b1 , w_30762 );
and ( \12095_b0 , \12013_b0 , w_30763 );
and ( w_30762 , w_30763 , \12018_b0 );
or ( \12097_b1 , \12092_b1 , \12096_b1 );
xor ( \12097_b0 , \12092_b0 , w_30764 );
not ( w_30764 , w_30765 );
and ( w_30765 , \12096_b1 , \12096_b0 );
or ( \12098_b1 , \12083_b1 , \12097_b1 );
xor ( \12098_b0 , \12083_b0 , w_30766 );
not ( w_30766 , w_30767 );
and ( w_30767 , \12097_b1 , \12097_b0 );
or ( \12099_b1 , \12065_b1 , \12098_b1 );
xor ( \12099_b0 , \12065_b0 , w_30768 );
not ( w_30768 , w_30769 );
and ( w_30769 , \12098_b1 , \12098_b0 );
or ( \12100_b1 , \12056_b1 , \12099_b1 );
xor ( \12100_b0 , \12056_b0 , w_30770 );
not ( w_30770 , w_30771 );
and ( w_30771 , \12099_b1 , \12099_b0 );
or ( \12101_b1 , \11946_b1 , \11960_b1 );
not ( \11960_b1 , w_30772 );
and ( \12101_b0 , \11946_b0 , w_30773 );
and ( w_30772 , w_30773 , \11960_b0 );
or ( \12102_b1 , \11960_b1 , \12034_b1 );
not ( \12034_b1 , w_30774 );
and ( \12102_b0 , \11960_b0 , w_30775 );
and ( w_30774 , w_30775 , \12034_b0 );
or ( \12103_b1 , \11946_b1 , \12034_b1 );
not ( \12034_b1 , w_30776 );
and ( \12103_b0 , \11946_b0 , w_30777 );
and ( w_30776 , w_30777 , \12034_b0 );
or ( \12105_b1 , \12100_b1 , w_30779 );
not ( w_30779 , w_30780 );
and ( \12105_b0 , \12100_b0 , w_30781 );
and ( w_30780 ,  , w_30781 );
buf ( w_30779 , \12104_b1 );
not ( w_30779 , w_30782 );
not (  , w_30783 );
and ( w_30782 , w_30783 , \12104_b0 );
or ( \12106_b1 , \12040_b1 , w_30785 );
not ( w_30785 , w_30786 );
and ( \12106_b0 , \12040_b0 , w_30787 );
and ( w_30786 ,  , w_30787 );
buf ( w_30785 , \12105_b1 );
not ( w_30785 , w_30788 );
not (  , w_30789 );
and ( w_30788 , w_30789 , \12105_b0 );
or ( \12107_b1 , \11942_b1 , w_30791 );
not ( w_30791 , w_30792 );
and ( \12107_b0 , \11942_b0 , w_30793 );
and ( w_30792 ,  , w_30793 );
buf ( w_30791 , \12106_b1 );
not ( w_30791 , w_30794 );
not (  , w_30795 );
and ( w_30794 , w_30795 , \12106_b0 );
or ( \12108_b1 , \12060_b1 , \12064_b1 );
not ( \12064_b1 , w_30796 );
and ( \12108_b0 , \12060_b0 , w_30797 );
and ( w_30796 , w_30797 , \12064_b0 );
or ( \12109_b1 , \12064_b1 , \12098_b1 );
not ( \12098_b1 , w_30798 );
and ( \12109_b0 , \12064_b0 , w_30799 );
and ( w_30798 , w_30799 , \12098_b0 );
or ( \12110_b1 , \12060_b1 , \12098_b1 );
not ( \12098_b1 , w_30800 );
and ( \12110_b0 , \12060_b0 , w_30801 );
and ( w_30800 , w_30801 , \12098_b0 );
or ( \12112_b1 , \12087_b1 , \12091_b1 );
not ( \12091_b1 , w_30802 );
and ( \12112_b0 , \12087_b0 , w_30803 );
and ( w_30802 , w_30803 , \12091_b0 );
or ( \12113_b1 , \12091_b1 , \12096_b1 );
not ( \12096_b1 , w_30804 );
and ( \12113_b0 , \12091_b0 , w_30805 );
and ( w_30804 , w_30805 , \12096_b0 );
or ( \12114_b1 , \12087_b1 , \12096_b1 );
not ( \12096_b1 , w_30806 );
and ( \12114_b0 , \12087_b0 , w_30807 );
and ( w_30806 , w_30807 , \12096_b0 );
or ( \12116_b1 , \12076_b1 , \12078_b1 );
not ( \12078_b1 , w_30808 );
and ( \12116_b0 , \12076_b0 , w_30809 );
and ( w_30808 , w_30809 , \12078_b0 );
or ( \12117_b1 , \12078_b1 , \12081_b1 );
not ( \12081_b1 , w_30810 );
and ( \12117_b0 , \12078_b0 , w_30811 );
and ( w_30810 , w_30811 , \12081_b0 );
or ( \12118_b1 , \12076_b1 , \12081_b1 );
not ( \12081_b1 , w_30812 );
and ( \12118_b0 , \12076_b0 , w_30813 );
and ( w_30812 , w_30813 , \12081_b0 );
or ( \12120_b1 , \12115_b1 , \12119_b1 );
xor ( \12120_b0 , \12115_b0 , w_30814 );
not ( w_30814 , w_30815 );
and ( w_30815 , \12119_b1 , \12119_b0 );
or ( \12121_b1 , \12066_b1 , \12068_b1 );
not ( \12068_b1 , w_30816 );
and ( \12121_b0 , \12066_b0 , w_30817 );
and ( w_30816 , w_30817 , \12068_b0 );
or ( \12122_b1 , \12068_b1 , \12071_b1 );
not ( \12071_b1 , w_30818 );
and ( \12122_b0 , \12068_b0 , w_30819 );
and ( w_30818 , w_30819 , \12071_b0 );
or ( \12123_b1 , \12066_b1 , \12071_b1 );
not ( \12071_b1 , w_30820 );
and ( \12123_b0 , \12066_b0 , w_30821 );
and ( w_30820 , w_30821 , \12071_b0 );
or ( \12125_b1 , \12120_b1 , \12124_b1 );
xor ( \12125_b0 , \12120_b0 , w_30822 );
not ( w_30822 , w_30823 );
and ( w_30823 , \12124_b1 , \12124_b0 );
or ( \12126_b1 , \12111_b1 , \12125_b1 );
xor ( \12126_b0 , \12111_b0 , w_30824 );
not ( w_30824 , w_30825 );
and ( w_30825 , \12125_b1 , \12125_b0 );
or ( \12127_b1 , \12048_b1 , \12052_b1 );
not ( \12052_b1 , w_30826 );
and ( \12127_b0 , \12048_b0 , w_30827 );
and ( w_30826 , w_30827 , \12052_b0 );
or ( \12128_b1 , \12052_b1 , \12054_b1 );
not ( \12054_b1 , w_30828 );
and ( \12128_b0 , \12052_b0 , w_30829 );
and ( w_30828 , w_30829 , \12054_b0 );
or ( \12129_b1 , \12048_b1 , \12054_b1 );
not ( \12054_b1 , w_30830 );
and ( \12129_b0 , \12048_b0 , w_30831 );
and ( w_30830 , w_30831 , \12054_b0 );
or ( \12131_b1 , \12072_b1 , \12082_b1 );
not ( \12082_b1 , w_30832 );
and ( \12131_b0 , \12072_b0 , w_30833 );
and ( w_30832 , w_30833 , \12082_b0 );
or ( \12132_b1 , \12082_b1 , \12097_b1 );
not ( \12097_b1 , w_30834 );
and ( \12132_b0 , \12082_b0 , w_30835 );
and ( w_30834 , w_30835 , \12097_b0 );
or ( \12133_b1 , \12072_b1 , \12097_b1 );
not ( \12097_b1 , w_30836 );
and ( \12133_b0 , \12072_b0 , w_30837 );
and ( w_30836 , w_30837 , \12097_b0 );
or ( \12135_b1 , \12130_b1 , \12134_b1 );
xor ( \12135_b0 , \12130_b0 , w_30838 );
not ( w_30838 , w_30839 );
and ( w_30839 , \12134_b1 , \12134_b0 );
or ( \12136_b1 , \6948_b1 , \6950_b1 );
xor ( \12136_b0 , \6948_b0 , w_30840 );
not ( w_30840 , w_30841 );
and ( w_30841 , \6950_b1 , \6950_b0 );
or ( \12137_b1 , \6937_b1 , \6939_b1 );
xor ( \12137_b0 , \6937_b0 , w_30842 );
not ( w_30842 , w_30843 );
and ( w_30843 , \6939_b1 , \6939_b0 );
or ( \12138_b1 , \12137_b1 , \6942_b1 );
xor ( \12138_b0 , \12137_b0 , w_30844 );
not ( w_30844 , w_30845 );
and ( w_30845 , \6942_b1 , \6942_b0 );
or ( \12139_b1 , \12136_b1 , \12138_b1 );
xor ( \12139_b0 , \12136_b0 , w_30846 );
not ( w_30846 , w_30847 );
and ( w_30847 , \12138_b1 , \12138_b0 );
or ( \12140_b1 , \6873_b1 , \6918_b1 );
xor ( \12140_b0 , \6873_b0 , w_30848 );
not ( w_30848 , w_30849 );
and ( w_30849 , \6918_b1 , \6918_b0 );
or ( \12141_b1 , \12140_b1 , \6924_b1 );
xor ( \12141_b0 , \12140_b0 , w_30850 );
not ( w_30850 , w_30851 );
and ( w_30851 , \6924_b1 , \6924_b0 );
or ( \12142_b1 , \12139_b1 , \12141_b1 );
xor ( \12142_b0 , \12139_b0 , w_30852 );
not ( w_30852 , w_30853 );
and ( w_30853 , \12141_b1 , \12141_b0 );
or ( \12143_b1 , \12135_b1 , \12142_b1 );
xor ( \12143_b0 , \12135_b0 , w_30854 );
not ( w_30854 , w_30855 );
and ( w_30855 , \12142_b1 , \12142_b0 );
or ( \12144_b1 , \12126_b1 , \12143_b1 );
xor ( \12144_b0 , \12126_b0 , w_30856 );
not ( w_30856 , w_30857 );
and ( w_30857 , \12143_b1 , \12143_b0 );
or ( \12145_b1 , \12044_b1 , \12055_b1 );
not ( \12055_b1 , w_30858 );
and ( \12145_b0 , \12044_b0 , w_30859 );
and ( w_30858 , w_30859 , \12055_b0 );
or ( \12146_b1 , \12055_b1 , \12099_b1 );
not ( \12099_b1 , w_30860 );
and ( \12146_b0 , \12055_b0 , w_30861 );
and ( w_30860 , w_30861 , \12099_b0 );
or ( \12147_b1 , \12044_b1 , \12099_b1 );
not ( \12099_b1 , w_30862 );
and ( \12147_b0 , \12044_b0 , w_30863 );
and ( w_30862 , w_30863 , \12099_b0 );
or ( \12149_b1 , \12144_b1 , w_30865 );
not ( w_30865 , w_30866 );
and ( \12149_b0 , \12144_b0 , w_30867 );
and ( w_30866 ,  , w_30867 );
buf ( w_30865 , \12148_b1 );
not ( w_30865 , w_30868 );
not (  , w_30869 );
and ( w_30868 , w_30869 , \12148_b0 );
or ( \12150_b1 , \12130_b1 , \12134_b1 );
not ( \12134_b1 , w_30870 );
and ( \12150_b0 , \12130_b0 , w_30871 );
and ( w_30870 , w_30871 , \12134_b0 );
or ( \12151_b1 , \12134_b1 , \12142_b1 );
not ( \12142_b1 , w_30872 );
and ( \12151_b0 , \12134_b0 , w_30873 );
and ( w_30872 , w_30873 , \12142_b0 );
or ( \12152_b1 , \12130_b1 , \12142_b1 );
not ( \12142_b1 , w_30874 );
and ( \12152_b0 , \12130_b0 , w_30875 );
and ( w_30874 , w_30875 , \12142_b0 );
or ( \12154_b1 , \6927_b1 , \6945_b1 );
xor ( \12154_b0 , \6927_b0 , w_30876 );
not ( w_30876 , w_30877 );
and ( w_30877 , \6945_b1 , \6945_b0 );
or ( \12155_b1 , \12154_b1 , \6951_b1 );
xor ( \12155_b0 , \12154_b0 , w_30878 );
not ( w_30878 , w_30879 );
and ( w_30879 , \6951_b1 , \6951_b0 );
or ( \12156_b1 , \12153_b1 , \12155_b1 );
xor ( \12156_b0 , \12153_b0 , w_30880 );
not ( w_30880 , w_30881 );
and ( w_30881 , \12155_b1 , \12155_b0 );
or ( \12157_b1 , \12115_b1 , \12119_b1 );
not ( \12119_b1 , w_30882 );
and ( \12157_b0 , \12115_b0 , w_30883 );
and ( w_30882 , w_30883 , \12119_b0 );
or ( \12158_b1 , \12119_b1 , \12124_b1 );
not ( \12124_b1 , w_30884 );
and ( \12158_b0 , \12119_b0 , w_30885 );
and ( w_30884 , w_30885 , \12124_b0 );
or ( \12159_b1 , \12115_b1 , \12124_b1 );
not ( \12124_b1 , w_30886 );
and ( \12159_b0 , \12115_b0 , w_30887 );
and ( w_30886 , w_30887 , \12124_b0 );
or ( \12161_b1 , \12136_b1 , \12138_b1 );
not ( \12138_b1 , w_30888 );
and ( \12161_b0 , \12136_b0 , w_30889 );
and ( w_30888 , w_30889 , \12138_b0 );
or ( \12162_b1 , \12138_b1 , \12141_b1 );
not ( \12141_b1 , w_30890 );
and ( \12162_b0 , \12138_b0 , w_30891 );
and ( w_30890 , w_30891 , \12141_b0 );
or ( \12163_b1 , \12136_b1 , \12141_b1 );
not ( \12141_b1 , w_30892 );
and ( \12163_b0 , \12136_b0 , w_30893 );
and ( w_30892 , w_30893 , \12141_b0 );
or ( \12165_b1 , \12160_b1 , \12164_b1 );
xor ( \12165_b0 , \12160_b0 , w_30894 );
not ( w_30894 , w_30895 );
and ( w_30895 , \12164_b1 , \12164_b0 );
or ( \12166_b1 , \6956_b1 , \6958_b1 );
xor ( \12166_b0 , \6956_b0 , w_30896 );
not ( w_30896 , w_30897 );
and ( w_30897 , \6958_b1 , \6958_b0 );
or ( \12167_b1 , \12166_b1 , \6961_b1 );
xor ( \12167_b0 , \12166_b0 , w_30898 );
not ( w_30898 , w_30899 );
and ( w_30899 , \6961_b1 , \6961_b0 );
or ( \12168_b1 , \12165_b1 , \12167_b1 );
xor ( \12168_b0 , \12165_b0 , w_30900 );
not ( w_30900 , w_30901 );
and ( w_30901 , \12167_b1 , \12167_b0 );
or ( \12169_b1 , \12156_b1 , \12168_b1 );
xor ( \12169_b0 , \12156_b0 , w_30902 );
not ( w_30902 , w_30903 );
and ( w_30903 , \12168_b1 , \12168_b0 );
or ( \12170_b1 , \12111_b1 , \12125_b1 );
not ( \12125_b1 , w_30904 );
and ( \12170_b0 , \12111_b0 , w_30905 );
and ( w_30904 , w_30905 , \12125_b0 );
or ( \12171_b1 , \12125_b1 , \12143_b1 );
not ( \12143_b1 , w_30906 );
and ( \12171_b0 , \12125_b0 , w_30907 );
and ( w_30906 , w_30907 , \12143_b0 );
or ( \12172_b1 , \12111_b1 , \12143_b1 );
not ( \12143_b1 , w_30908 );
and ( \12172_b0 , \12111_b0 , w_30909 );
and ( w_30908 , w_30909 , \12143_b0 );
or ( \12174_b1 , \12169_b1 , w_30911 );
not ( w_30911 , w_30912 );
and ( \12174_b0 , \12169_b0 , w_30913 );
and ( w_30912 ,  , w_30913 );
buf ( w_30911 , \12173_b1 );
not ( w_30911 , w_30914 );
not (  , w_30915 );
and ( w_30914 , w_30915 , \12173_b0 );
or ( \12175_b1 , \12149_b1 , w_30917 );
not ( w_30917 , w_30918 );
and ( \12175_b0 , \12149_b0 , w_30919 );
and ( w_30918 ,  , w_30919 );
buf ( w_30917 , \12174_b1 );
not ( w_30917 , w_30920 );
not (  , w_30921 );
and ( w_30920 , w_30921 , \12174_b0 );
or ( \12176_b1 , \12160_b1 , \12164_b1 );
not ( \12164_b1 , w_30922 );
and ( \12176_b0 , \12160_b0 , w_30923 );
and ( w_30922 , w_30923 , \12164_b0 );
or ( \12177_b1 , \12164_b1 , \12167_b1 );
not ( \12167_b1 , w_30924 );
and ( \12177_b0 , \12164_b0 , w_30925 );
and ( w_30924 , w_30925 , \12167_b0 );
or ( \12178_b1 , \12160_b1 , \12167_b1 );
not ( \12167_b1 , w_30926 );
and ( \12178_b0 , \12160_b0 , w_30927 );
and ( w_30926 , w_30927 , \12167_b0 );
or ( \12180_b1 , \6122_b1 , \6284_b1 );
xor ( \12180_b0 , \6122_b0 , w_30928 );
not ( w_30928 , w_30929 );
and ( w_30929 , \6284_b1 , \6284_b0 );
or ( \12181_b1 , \12180_b1 , \6342_b1 );
xor ( \12181_b0 , \12180_b0 , w_30930 );
not ( w_30930 , w_30931 );
and ( w_30931 , \6342_b1 , \6342_b0 );
or ( \12182_b1 , \12179_b1 , \12181_b1 );
xor ( \12182_b0 , \12179_b0 , w_30932 );
not ( w_30932 , w_30933 );
and ( w_30933 , \12181_b1 , \12181_b0 );
or ( \12183_b1 , \6954_b1 , \6964_b1 );
xor ( \12183_b0 , \6954_b0 , w_30934 );
not ( w_30934 , w_30935 );
and ( w_30935 , \6964_b1 , \6964_b0 );
or ( \12184_b1 , \12183_b1 , \6967_b1 );
xor ( \12184_b0 , \12183_b0 , w_30936 );
not ( w_30936 , w_30937 );
and ( w_30937 , \6967_b1 , \6967_b0 );
or ( \12185_b1 , \12182_b1 , \12184_b1 );
xor ( \12185_b0 , \12182_b0 , w_30938 );
not ( w_30938 , w_30939 );
and ( w_30939 , \12184_b1 , \12184_b0 );
or ( \12186_b1 , \12153_b1 , \12155_b1 );
not ( \12155_b1 , w_30940 );
and ( \12186_b0 , \12153_b0 , w_30941 );
and ( w_30940 , w_30941 , \12155_b0 );
or ( \12187_b1 , \12155_b1 , \12168_b1 );
not ( \12168_b1 , w_30942 );
and ( \12187_b0 , \12155_b0 , w_30943 );
and ( w_30942 , w_30943 , \12168_b0 );
or ( \12188_b1 , \12153_b1 , \12168_b1 );
not ( \12168_b1 , w_30944 );
and ( \12188_b0 , \12153_b0 , w_30945 );
and ( w_30944 , w_30945 , \12168_b0 );
or ( \12190_b1 , \12185_b1 , w_30947 );
not ( w_30947 , w_30948 );
and ( \12190_b0 , \12185_b0 , w_30949 );
and ( w_30948 ,  , w_30949 );
buf ( w_30947 , \12189_b1 );
not ( w_30947 , w_30950 );
not (  , w_30951 );
and ( w_30950 , w_30951 , \12189_b0 );
or ( \12191_b1 , \6970_b1 , \6972_b1 );
xor ( \12191_b0 , \6970_b0 , w_30952 );
not ( w_30952 , w_30953 );
and ( w_30953 , \6972_b1 , \6972_b0 );
or ( \12192_b1 , \12191_b1 , \6975_b1 );
xor ( \12192_b0 , \12191_b0 , w_30954 );
not ( w_30954 , w_30955 );
and ( w_30955 , \6975_b1 , \6975_b0 );
or ( \12193_b1 , \12179_b1 , \12181_b1 );
not ( \12181_b1 , w_30956 );
and ( \12193_b0 , \12179_b0 , w_30957 );
and ( w_30956 , w_30957 , \12181_b0 );
or ( \12194_b1 , \12181_b1 , \12184_b1 );
not ( \12184_b1 , w_30958 );
and ( \12194_b0 , \12181_b0 , w_30959 );
and ( w_30958 , w_30959 , \12184_b0 );
or ( \12195_b1 , \12179_b1 , \12184_b1 );
not ( \12184_b1 , w_30960 );
and ( \12195_b0 , \12179_b0 , w_30961 );
and ( w_30960 , w_30961 , \12184_b0 );
or ( \12197_b1 , \12192_b1 , w_30963 );
not ( w_30963 , w_30964 );
and ( \12197_b0 , \12192_b0 , w_30965 );
and ( w_30964 ,  , w_30965 );
buf ( w_30963 , \12196_b1 );
not ( w_30963 , w_30966 );
not (  , w_30967 );
and ( w_30966 , w_30967 , \12196_b0 );
or ( \12198_b1 , \12190_b1 , w_30969 );
not ( w_30969 , w_30970 );
and ( \12198_b0 , \12190_b0 , w_30971 );
and ( w_30970 ,  , w_30971 );
buf ( w_30969 , \12197_b1 );
not ( w_30969 , w_30972 );
not (  , w_30973 );
and ( w_30972 , w_30973 , \12197_b0 );
or ( \12199_b1 , \12175_b1 , w_30975 );
not ( w_30975 , w_30976 );
and ( \12199_b0 , \12175_b0 , w_30977 );
and ( w_30976 ,  , w_30977 );
buf ( w_30975 , \12198_b1 );
not ( w_30975 , w_30978 );
not (  , w_30979 );
and ( w_30978 , w_30979 , \12198_b0 );
or ( \12200_b1 , \12107_b1 , w_30981 );
not ( w_30981 , w_30982 );
and ( \12200_b0 , \12107_b0 , w_30983 );
and ( w_30982 ,  , w_30983 );
buf ( w_30981 , \12199_b1 );
not ( w_30981 , w_30984 );
not (  , w_30985 );
and ( w_30984 , w_30985 , \12199_b0 );
or ( \12201_b1 , \11617_b1 , w_30987 );
not ( w_30987 , w_30988 );
and ( \12201_b0 , \11617_b0 , w_30989 );
and ( w_30988 ,  , w_30989 );
buf ( w_30987 , \12200_b1 );
not ( w_30987 , w_30990 );
not (  , w_30991 );
and ( w_30990 , w_30991 , \12200_b0 );
or ( \12202_b1 , \10314_b1 , w_30993 );
not ( w_30993 , w_30994 );
and ( \12202_b0 , \10314_b0 , w_30995 );
and ( w_30994 ,  , w_30995 );
buf ( w_30993 , \12201_b1 );
not ( w_30993 , w_30996 );
not (  , w_30997 );
and ( w_30996 , w_30997 , \12201_b0 );
or ( \12203_b1 , \5945_b1 , \6991_b1 );
not ( \6991_b1 , w_30998 );
and ( \12203_b0 , \5945_b0 , w_30999 );
and ( w_30998 , w_30999 , \6991_b0 );
or ( \12204_b1 , \5957_b1 , \6988_b1 );
not ( \6988_b1 , w_31000 );
and ( \12204_b0 , \5957_b0 , w_31001 );
and ( w_31000 , w_31001 , \6988_b0 );
or ( \12205_b1 , \12203_b1 , w_31003 );
not ( w_31003 , w_31004 );
and ( \12205_b0 , \12203_b0 , w_31005 );
and ( w_31004 ,  , w_31005 );
buf ( w_31003 , \12204_b1 );
not ( w_31003 , w_31006 );
not (  , w_31007 );
and ( w_31006 , w_31007 , \12204_b0 );
or ( \12206_b1 , \12205_b1 , w_31008 );
xor ( \12206_b0 , \12205_b0 , w_31010 );
not ( w_31010 , w_31011 );
and ( w_31011 , w_31008 , w_31009 );
buf ( w_31008 , \6985_b1 );
not ( w_31008 , w_31012 );
not ( w_31009 , w_31013 );
and ( w_31012 , w_31013 , \6985_b0 );
or ( \12207_b1 , \7105_b1 , \12206_b1 );
not ( \12206_b1 , w_31014 );
and ( \12207_b0 , \7105_b0 , w_31015 );
and ( w_31014 , w_31015 , \12206_b0 );
or ( \12208_b1 , \5967_b1 , \7006_b1 );
not ( \7006_b1 , w_31016 );
and ( \12208_b0 , \5967_b0 , w_31017 );
and ( w_31016 , w_31017 , \7006_b0 );
or ( \12209_b1 , \5979_b1 , \7004_b1 );
not ( \7004_b1 , w_31018 );
and ( \12209_b0 , \5979_b0 , w_31019 );
and ( w_31018 , w_31019 , \7004_b0 );
or ( \12210_b1 , \12208_b1 , w_31021 );
not ( w_31021 , w_31022 );
and ( \12210_b0 , \12208_b0 , w_31023 );
and ( w_31022 ,  , w_31023 );
buf ( w_31021 , \12209_b1 );
not ( w_31021 , w_31024 );
not (  , w_31025 );
and ( w_31024 , w_31025 , \12209_b0 );
or ( \12211_b1 , \12210_b1 , w_31026 );
xor ( \12211_b0 , \12210_b0 , w_31028 );
not ( w_31028 , w_31029 );
and ( w_31029 , w_31026 , w_31027 );
buf ( w_31026 , \7012_b1 );
not ( w_31026 , w_31030 );
not ( w_31027 , w_31031 );
and ( w_31030 , w_31031 , \7012_b0 );
or ( \12212_b1 , \12206_b1 , \12211_b1 );
not ( \12211_b1 , w_31032 );
and ( \12212_b0 , \12206_b0 , w_31033 );
and ( w_31032 , w_31033 , \12211_b0 );
or ( \12213_b1 , \7105_b1 , \12211_b1 );
not ( \12211_b1 , w_31034 );
and ( \12213_b0 , \7105_b0 , w_31035 );
and ( w_31034 , w_31035 , \12211_b0 );
or ( \12215_b1 , \5986_b1 , \7026_b1 );
not ( \7026_b1 , w_31036 );
and ( \12215_b0 , \5986_b0 , w_31037 );
and ( w_31036 , w_31037 , \7026_b0 );
or ( \12216_b1 , \5998_b1 , \7024_b1 );
not ( \7024_b1 , w_31038 );
and ( \12216_b0 , \5998_b0 , w_31039 );
and ( w_31038 , w_31039 , \7024_b0 );
or ( \12217_b1 , \12215_b1 , w_31041 );
not ( w_31041 , w_31042 );
and ( \12217_b0 , \12215_b0 , w_31043 );
and ( w_31042 ,  , w_31043 );
buf ( w_31041 , \12216_b1 );
not ( w_31041 , w_31044 );
not (  , w_31045 );
and ( w_31044 , w_31045 , \12216_b0 );
or ( \12218_b1 , \12217_b1 , w_31046 );
xor ( \12218_b0 , \12217_b0 , w_31048 );
not ( w_31048 , w_31049 );
and ( w_31049 , w_31046 , w_31047 );
buf ( w_31046 , \7032_b1 );
not ( w_31046 , w_31050 );
not ( w_31047 , w_31051 );
and ( w_31050 , w_31051 , \7032_b0 );
or ( \12219_b1 , \6006_b1 , \7043_b1 );
not ( \7043_b1 , w_31052 );
and ( \12219_b0 , \6006_b0 , w_31053 );
and ( w_31052 , w_31053 , \7043_b0 );
or ( \12220_b1 , \6018_b1 , \7041_b1 );
not ( \7041_b1 , w_31054 );
and ( \12220_b0 , \6018_b0 , w_31055 );
and ( w_31054 , w_31055 , \7041_b0 );
or ( \12221_b1 , \12219_b1 , w_31057 );
not ( w_31057 , w_31058 );
and ( \12221_b0 , \12219_b0 , w_31059 );
and ( w_31058 ,  , w_31059 );
buf ( w_31057 , \12220_b1 );
not ( w_31057 , w_31060 );
not (  , w_31061 );
and ( w_31060 , w_31061 , \12220_b0 );
or ( \12222_b1 , \12221_b1 , w_31062 );
xor ( \12222_b0 , \12221_b0 , w_31064 );
not ( w_31064 , w_31065 );
and ( w_31065 , w_31062 , w_31063 );
buf ( w_31062 , \7049_b1 );
not ( w_31062 , w_31066 );
not ( w_31063 , w_31067 );
and ( w_31066 , w_31067 , \7049_b0 );
or ( \12223_b1 , \12218_b1 , \12222_b1 );
not ( \12222_b1 , w_31068 );
and ( \12223_b0 , \12218_b0 , w_31069 );
and ( w_31068 , w_31069 , \12222_b0 );
or ( \12224_b1 , \6029_b1 , \7061_b1 );
not ( \7061_b1 , w_31070 );
and ( \12224_b0 , \6029_b0 , w_31071 );
and ( w_31070 , w_31071 , \7061_b0 );
or ( \12225_b1 , \6041_b1 , \7059_b1 );
not ( \7059_b1 , w_31072 );
and ( \12225_b0 , \6041_b0 , w_31073 );
and ( w_31072 , w_31073 , \7059_b0 );
or ( \12226_b1 , \12224_b1 , w_31075 );
not ( w_31075 , w_31076 );
and ( \12226_b0 , \12224_b0 , w_31077 );
and ( w_31076 ,  , w_31077 );
buf ( w_31075 , \12225_b1 );
not ( w_31075 , w_31078 );
not (  , w_31079 );
and ( w_31078 , w_31079 , \12225_b0 );
or ( \12227_b1 , \12226_b1 , w_31080 );
xor ( \12227_b0 , \12226_b0 , w_31082 );
not ( w_31082 , w_31083 );
and ( w_31083 , w_31080 , w_31081 );
buf ( w_31080 , \7067_b1 );
not ( w_31080 , w_31084 );
not ( w_31081 , w_31085 );
and ( w_31084 , w_31085 , \7067_b0 );
or ( \12228_b1 , \12222_b1 , \12227_b1 );
not ( \12227_b1 , w_31086 );
and ( \12228_b0 , \12222_b0 , w_31087 );
and ( w_31086 , w_31087 , \12227_b0 );
or ( \12229_b1 , \12218_b1 , \12227_b1 );
not ( \12227_b1 , w_31088 );
and ( \12229_b0 , \12218_b0 , w_31089 );
and ( w_31088 , w_31089 , \12227_b0 );
or ( \12231_b1 , \12214_b1 , \12230_b1 );
not ( \12230_b1 , w_31090 );
and ( \12231_b0 , \12214_b0 , w_31091 );
and ( w_31090 , w_31091 , \12230_b0 );
or ( \12232_b1 , \6065_b1 , \7099_b1 );
not ( \7099_b1 , w_31092 );
and ( \12232_b0 , \6065_b0 , w_31093 );
and ( w_31092 , w_31093 , \7099_b0 );
or ( \12233_b1 , \6048_b1 , \7097_b1 );
not ( \7097_b1 , w_31094 );
and ( \12233_b0 , \6048_b0 , w_31095 );
and ( w_31094 , w_31095 , \7097_b0 );
or ( \12234_b1 , \12232_b1 , w_31097 );
not ( w_31097 , w_31098 );
and ( \12234_b0 , \12232_b0 , w_31099 );
and ( w_31098 ,  , w_31099 );
buf ( w_31097 , \12233_b1 );
not ( w_31097 , w_31100 );
not (  , w_31101 );
and ( w_31100 , w_31101 , \12233_b0 );
or ( \12235_b1 , \12234_b1 , w_31102 );
xor ( \12235_b0 , \12234_b0 , w_31104 );
not ( w_31104 , w_31105 );
and ( w_31105 , w_31102 , w_31103 );
buf ( w_31102 , \7105_b1 );
not ( w_31102 , w_31106 );
not ( w_31103 , w_31107 );
and ( w_31106 , w_31107 , \7105_b0 );
or ( \12236_b1 , \12230_b1 , \12235_b1 );
not ( \12235_b1 , w_31108 );
and ( \12236_b0 , \12230_b0 , w_31109 );
and ( w_31108 , w_31109 , \12235_b0 );
or ( \12237_b1 , \12214_b1 , \12235_b1 );
not ( \12235_b1 , w_31110 );
and ( \12237_b0 , \12214_b0 , w_31111 );
and ( w_31110 , w_31111 , \12235_b0 );
or ( \12239_b1 , \5967_b1 , \7026_b1 );
not ( \7026_b1 , w_31112 );
and ( \12239_b0 , \5967_b0 , w_31113 );
and ( w_31112 , w_31113 , \7026_b0 );
or ( \12240_b1 , \5979_b1 , \7024_b1 );
not ( \7024_b1 , w_31114 );
and ( \12240_b0 , \5979_b0 , w_31115 );
and ( w_31114 , w_31115 , \7024_b0 );
or ( \12241_b1 , \12239_b1 , w_31117 );
not ( w_31117 , w_31118 );
and ( \12241_b0 , \12239_b0 , w_31119 );
and ( w_31118 ,  , w_31119 );
buf ( w_31117 , \12240_b1 );
not ( w_31117 , w_31120 );
not (  , w_31121 );
and ( w_31120 , w_31121 , \12240_b0 );
or ( \12242_b1 , \12241_b1 , w_31122 );
xor ( \12242_b0 , \12241_b0 , w_31124 );
not ( w_31124 , w_31125 );
and ( w_31125 , w_31122 , w_31123 );
buf ( w_31122 , \7032_b1 );
not ( w_31122 , w_31126 );
not ( w_31123 , w_31127 );
and ( w_31126 , w_31127 , \7032_b0 );
or ( \12243_b1 , \5986_b1 , \7043_b1 );
not ( \7043_b1 , w_31128 );
and ( \12243_b0 , \5986_b0 , w_31129 );
and ( w_31128 , w_31129 , \7043_b0 );
or ( \12244_b1 , \5998_b1 , \7041_b1 );
not ( \7041_b1 , w_31130 );
and ( \12244_b0 , \5998_b0 , w_31131 );
and ( w_31130 , w_31131 , \7041_b0 );
or ( \12245_b1 , \12243_b1 , w_31133 );
not ( w_31133 , w_31134 );
and ( \12245_b0 , \12243_b0 , w_31135 );
and ( w_31134 ,  , w_31135 );
buf ( w_31133 , \12244_b1 );
not ( w_31133 , w_31136 );
not (  , w_31137 );
and ( w_31136 , w_31137 , \12244_b0 );
or ( \12246_b1 , \12245_b1 , w_31138 );
xor ( \12246_b0 , \12245_b0 , w_31140 );
not ( w_31140 , w_31141 );
and ( w_31141 , w_31138 , w_31139 );
buf ( w_31138 , \7049_b1 );
not ( w_31138 , w_31142 );
not ( w_31139 , w_31143 );
and ( w_31142 , w_31143 , \7049_b0 );
or ( \12247_b1 , \12242_b1 , \12246_b1 );
xor ( \12247_b0 , \12242_b0 , w_31144 );
not ( w_31144 , w_31145 );
and ( w_31145 , \12246_b1 , \12246_b0 );
or ( \12248_b1 , \6006_b1 , \7061_b1 );
not ( \7061_b1 , w_31146 );
and ( \12248_b0 , \6006_b0 , w_31147 );
and ( w_31146 , w_31147 , \7061_b0 );
or ( \12249_b1 , \6018_b1 , \7059_b1 );
not ( \7059_b1 , w_31148 );
and ( \12249_b0 , \6018_b0 , w_31149 );
and ( w_31148 , w_31149 , \7059_b0 );
or ( \12250_b1 , \12248_b1 , w_31151 );
not ( w_31151 , w_31152 );
and ( \12250_b0 , \12248_b0 , w_31153 );
and ( w_31152 ,  , w_31153 );
buf ( w_31151 , \12249_b1 );
not ( w_31151 , w_31154 );
not (  , w_31155 );
and ( w_31154 , w_31155 , \12249_b0 );
or ( \12251_b1 , \12250_b1 , w_31156 );
xor ( \12251_b0 , \12250_b0 , w_31158 );
not ( w_31158 , w_31159 );
and ( w_31159 , w_31156 , w_31157 );
buf ( w_31156 , \7067_b1 );
not ( w_31156 , w_31160 );
not ( w_31157 , w_31161 );
and ( w_31160 , w_31161 , \7067_b0 );
or ( \12252_b1 , \12247_b1 , \12251_b1 );
xor ( \12252_b0 , \12247_b0 , w_31162 );
not ( w_31162 , w_31163 );
and ( w_31163 , \12251_b1 , \12251_b0 );
or ( \12253_b1 , \5925_b1 , \6991_b1 );
not ( \6991_b1 , w_31164 );
and ( \12253_b0 , \5925_b0 , w_31165 );
and ( w_31164 , w_31165 , \6991_b0 );
or ( \12254_b1 , \5937_b1 , \6988_b1 );
not ( \6988_b1 , w_31166 );
and ( \12254_b0 , \5937_b0 , w_31167 );
and ( w_31166 , w_31167 , \6988_b0 );
or ( \12255_b1 , \12253_b1 , w_31169 );
not ( w_31169 , w_31170 );
and ( \12255_b0 , \12253_b0 , w_31171 );
and ( w_31170 ,  , w_31171 );
buf ( w_31169 , \12254_b1 );
not ( w_31169 , w_31172 );
not (  , w_31173 );
and ( w_31172 , w_31173 , \12254_b0 );
or ( \12256_b1 , \12255_b1 , w_31174 );
xor ( \12256_b0 , \12255_b0 , w_31176 );
not ( w_31176 , w_31177 );
and ( w_31177 , w_31174 , w_31175 );
buf ( w_31174 , \6985_b1 );
not ( w_31174 , w_31178 );
not ( w_31175 , w_31179 );
and ( w_31178 , w_31179 , \6985_b0 );
or ( \12257_b1 , \7123_b1 , \12256_b1 );
xor ( \12257_b0 , \7123_b0 , w_31180 );
not ( w_31180 , w_31181 );
and ( w_31181 , \12256_b1 , \12256_b0 );
or ( \12258_b1 , \5945_b1 , \7006_b1 );
not ( \7006_b1 , w_31182 );
and ( \12258_b0 , \5945_b0 , w_31183 );
and ( w_31182 , w_31183 , \7006_b0 );
or ( \12259_b1 , \5957_b1 , \7004_b1 );
not ( \7004_b1 , w_31184 );
and ( \12259_b0 , \5957_b0 , w_31185 );
and ( w_31184 , w_31185 , \7004_b0 );
or ( \12260_b1 , \12258_b1 , w_31187 );
not ( w_31187 , w_31188 );
and ( \12260_b0 , \12258_b0 , w_31189 );
and ( w_31188 ,  , w_31189 );
buf ( w_31187 , \12259_b1 );
not ( w_31187 , w_31190 );
not (  , w_31191 );
and ( w_31190 , w_31191 , \12259_b0 );
or ( \12261_b1 , \12260_b1 , w_31192 );
xor ( \12261_b0 , \12260_b0 , w_31194 );
not ( w_31194 , w_31195 );
and ( w_31195 , w_31192 , w_31193 );
buf ( w_31192 , \7012_b1 );
not ( w_31192 , w_31196 );
not ( w_31193 , w_31197 );
and ( w_31196 , w_31197 , \7012_b0 );
or ( \12262_b1 , \12257_b1 , \12261_b1 );
xor ( \12262_b0 , \12257_b0 , w_31198 );
not ( w_31198 , w_31199 );
and ( w_31199 , \12261_b1 , \12261_b0 );
or ( \12263_b1 , \12252_b1 , \12262_b1 );
xor ( \12263_b0 , \12252_b0 , w_31200 );
not ( w_31200 , w_31201 );
and ( w_31201 , \12262_b1 , \12262_b0 );
or ( \12264_b1 , \12238_b1 , \12263_b1 );
not ( \12263_b1 , w_31202 );
and ( \12264_b0 , \12238_b0 , w_31203 );
and ( w_31202 , w_31203 , \12263_b0 );
or ( \12265_b1 , \5957_b1 , \6991_b1 );
not ( \6991_b1 , w_31204 );
and ( \12265_b0 , \5957_b0 , w_31205 );
and ( w_31204 , w_31205 , \6991_b0 );
or ( \12266_b1 , \5925_b1 , \6988_b1 );
not ( \6988_b1 , w_31206 );
and ( \12266_b0 , \5925_b0 , w_31207 );
and ( w_31206 , w_31207 , \6988_b0 );
or ( \12267_b1 , \12265_b1 , w_31209 );
not ( w_31209 , w_31210 );
and ( \12267_b0 , \12265_b0 , w_31211 );
and ( w_31210 ,  , w_31211 );
buf ( w_31209 , \12266_b1 );
not ( w_31209 , w_31212 );
not (  , w_31213 );
and ( w_31212 , w_31213 , \12266_b0 );
or ( \12268_b1 , \12267_b1 , w_31214 );
xor ( \12268_b0 , \12267_b0 , w_31216 );
not ( w_31216 , w_31217 );
and ( w_31217 , w_31214 , w_31215 );
buf ( w_31214 , \6985_b1 );
not ( w_31214 , w_31218 );
not ( w_31215 , w_31219 );
and ( w_31218 , w_31219 , \6985_b0 );
or ( \12269_b1 , \5979_b1 , \7006_b1 );
not ( \7006_b1 , w_31220 );
and ( \12269_b0 , \5979_b0 , w_31221 );
and ( w_31220 , w_31221 , \7006_b0 );
or ( \12270_b1 , \5945_b1 , \7004_b1 );
not ( \7004_b1 , w_31222 );
and ( \12270_b0 , \5945_b0 , w_31223 );
and ( w_31222 , w_31223 , \7004_b0 );
or ( \12271_b1 , \12269_b1 , w_31225 );
not ( w_31225 , w_31226 );
and ( \12271_b0 , \12269_b0 , w_31227 );
and ( w_31226 ,  , w_31227 );
buf ( w_31225 , \12270_b1 );
not ( w_31225 , w_31228 );
not (  , w_31229 );
and ( w_31228 , w_31229 , \12270_b0 );
or ( \12272_b1 , \12271_b1 , w_31230 );
xor ( \12272_b0 , \12271_b0 , w_31232 );
not ( w_31232 , w_31233 );
and ( w_31233 , w_31230 , w_31231 );
buf ( w_31230 , \7012_b1 );
not ( w_31230 , w_31234 );
not ( w_31231 , w_31235 );
and ( w_31234 , w_31235 , \7012_b0 );
or ( \12273_b1 , \12268_b1 , \12272_b1 );
not ( \12272_b1 , w_31236 );
and ( \12273_b0 , \12268_b0 , w_31237 );
and ( w_31236 , w_31237 , \12272_b0 );
or ( \12274_b1 , \5998_b1 , \7026_b1 );
not ( \7026_b1 , w_31238 );
and ( \12274_b0 , \5998_b0 , w_31239 );
and ( w_31238 , w_31239 , \7026_b0 );
or ( \12275_b1 , \5967_b1 , \7024_b1 );
not ( \7024_b1 , w_31240 );
and ( \12275_b0 , \5967_b0 , w_31241 );
and ( w_31240 , w_31241 , \7024_b0 );
or ( \12276_b1 , \12274_b1 , w_31243 );
not ( w_31243 , w_31244 );
and ( \12276_b0 , \12274_b0 , w_31245 );
and ( w_31244 ,  , w_31245 );
buf ( w_31243 , \12275_b1 );
not ( w_31243 , w_31246 );
not (  , w_31247 );
and ( w_31246 , w_31247 , \12275_b0 );
or ( \12277_b1 , \12276_b1 , w_31248 );
xor ( \12277_b0 , \12276_b0 , w_31250 );
not ( w_31250 , w_31251 );
and ( w_31251 , w_31248 , w_31249 );
buf ( w_31248 , \7032_b1 );
not ( w_31248 , w_31252 );
not ( w_31249 , w_31253 );
and ( w_31252 , w_31253 , \7032_b0 );
or ( \12278_b1 , \12272_b1 , \12277_b1 );
not ( \12277_b1 , w_31254 );
and ( \12278_b0 , \12272_b0 , w_31255 );
and ( w_31254 , w_31255 , \12277_b0 );
or ( \12279_b1 , \12268_b1 , \12277_b1 );
not ( \12277_b1 , w_31256 );
and ( \12279_b0 , \12268_b0 , w_31257 );
and ( w_31256 , w_31257 , \12277_b0 );
or ( \12281_b1 , \6018_b1 , \7043_b1 );
not ( \7043_b1 , w_31258 );
and ( \12281_b0 , \6018_b0 , w_31259 );
and ( w_31258 , w_31259 , \7043_b0 );
or ( \12282_b1 , \5986_b1 , \7041_b1 );
not ( \7041_b1 , w_31260 );
and ( \12282_b0 , \5986_b0 , w_31261 );
and ( w_31260 , w_31261 , \7041_b0 );
or ( \12283_b1 , \12281_b1 , w_31263 );
not ( w_31263 , w_31264 );
and ( \12283_b0 , \12281_b0 , w_31265 );
and ( w_31264 ,  , w_31265 );
buf ( w_31263 , \12282_b1 );
not ( w_31263 , w_31266 );
not (  , w_31267 );
and ( w_31266 , w_31267 , \12282_b0 );
or ( \12284_b1 , \12283_b1 , w_31268 );
xor ( \12284_b0 , \12283_b0 , w_31270 );
not ( w_31270 , w_31271 );
and ( w_31271 , w_31268 , w_31269 );
buf ( w_31268 , \7049_b1 );
not ( w_31268 , w_31272 );
not ( w_31269 , w_31273 );
and ( w_31272 , w_31273 , \7049_b0 );
or ( \12285_b1 , \6041_b1 , \7061_b1 );
not ( \7061_b1 , w_31274 );
and ( \12285_b0 , \6041_b0 , w_31275 );
and ( w_31274 , w_31275 , \7061_b0 );
or ( \12286_b1 , \6006_b1 , \7059_b1 );
not ( \7059_b1 , w_31276 );
and ( \12286_b0 , \6006_b0 , w_31277 );
and ( w_31276 , w_31277 , \7059_b0 );
or ( \12287_b1 , \12285_b1 , w_31279 );
not ( w_31279 , w_31280 );
and ( \12287_b0 , \12285_b0 , w_31281 );
and ( w_31280 ,  , w_31281 );
buf ( w_31279 , \12286_b1 );
not ( w_31279 , w_31282 );
not (  , w_31283 );
and ( w_31282 , w_31283 , \12286_b0 );
or ( \12288_b1 , \12287_b1 , w_31284 );
xor ( \12288_b0 , \12287_b0 , w_31286 );
not ( w_31286 , w_31287 );
and ( w_31287 , w_31284 , w_31285 );
buf ( w_31284 , \7067_b1 );
not ( w_31284 , w_31288 );
not ( w_31285 , w_31289 );
and ( w_31288 , w_31289 , \7067_b0 );
or ( \12289_b1 , \12284_b1 , \12288_b1 );
not ( \12288_b1 , w_31290 );
and ( \12289_b0 , \12284_b0 , w_31291 );
and ( w_31290 , w_31291 , \12288_b0 );
or ( \12290_b1 , \6057_b1 , \7082_b1 );
not ( \7082_b1 , w_31292 );
and ( \12290_b0 , \6057_b0 , w_31293 );
and ( w_31292 , w_31293 , \7082_b0 );
or ( \12291_b1 , \6029_b1 , \7080_b1 );
not ( \7080_b1 , w_31294 );
and ( \12291_b0 , \6029_b0 , w_31295 );
and ( w_31294 , w_31295 , \7080_b0 );
or ( \12292_b1 , \12290_b1 , w_31297 );
not ( w_31297 , w_31298 );
and ( \12292_b0 , \12290_b0 , w_31299 );
and ( w_31298 ,  , w_31299 );
buf ( w_31297 , \12291_b1 );
not ( w_31297 , w_31300 );
not (  , w_31301 );
and ( w_31300 , w_31301 , \12291_b0 );
or ( \12293_b1 , \12292_b1 , w_31302 );
xor ( \12293_b0 , \12292_b0 , w_31304 );
not ( w_31304 , w_31305 );
and ( w_31305 , w_31302 , w_31303 );
buf ( w_31302 , \7088_b1 );
not ( w_31302 , w_31306 );
not ( w_31303 , w_31307 );
and ( w_31306 , w_31307 , \7088_b0 );
or ( \12294_b1 , \12288_b1 , \12293_b1 );
not ( \12293_b1 , w_31308 );
and ( \12294_b0 , \12288_b0 , w_31309 );
and ( w_31308 , w_31309 , \12293_b0 );
or ( \12295_b1 , \12284_b1 , \12293_b1 );
not ( \12293_b1 , w_31310 );
and ( \12295_b0 , \12284_b0 , w_31311 );
and ( w_31310 , w_31311 , \12293_b0 );
or ( \12297_b1 , \12280_b1 , \12296_b1 );
xor ( \12297_b0 , \12280_b0 , w_31312 );
not ( w_31312 , w_31313 );
and ( w_31313 , \12296_b1 , \12296_b0 );
or ( \12298_b1 , \6029_b1 , \7082_b1 );
not ( \7082_b1 , w_31314 );
and ( \12298_b0 , \6029_b0 , w_31315 );
and ( w_31314 , w_31315 , \7082_b0 );
or ( \12299_b1 , \6041_b1 , \7080_b1 );
not ( \7080_b1 , w_31316 );
and ( \12299_b0 , \6041_b0 , w_31317 );
and ( w_31316 , w_31317 , \7080_b0 );
or ( \12300_b1 , \12298_b1 , w_31319 );
not ( w_31319 , w_31320 );
and ( \12300_b0 , \12298_b0 , w_31321 );
and ( w_31320 ,  , w_31321 );
buf ( w_31319 , \12299_b1 );
not ( w_31319 , w_31322 );
not (  , w_31323 );
and ( w_31322 , w_31323 , \12299_b0 );
or ( \12301_b1 , \12300_b1 , w_31324 );
xor ( \12301_b0 , \12300_b0 , w_31326 );
not ( w_31326 , w_31327 );
and ( w_31327 , w_31324 , w_31325 );
buf ( w_31324 , \7088_b1 );
not ( w_31324 , w_31328 );
not ( w_31325 , w_31329 );
and ( w_31328 , w_31329 , \7088_b0 );
or ( \12302_b1 , \6048_b1 , \7099_b1 );
not ( \7099_b1 , w_31330 );
and ( \12302_b0 , \6048_b0 , w_31331 );
and ( w_31330 , w_31331 , \7099_b0 );
or ( \12303_b1 , \6057_b1 , \7097_b1 );
not ( \7097_b1 , w_31332 );
and ( \12303_b0 , \6057_b0 , w_31333 );
and ( w_31332 , w_31333 , \7097_b0 );
or ( \12304_b1 , \12302_b1 , w_31335 );
not ( w_31335 , w_31336 );
and ( \12304_b0 , \12302_b0 , w_31337 );
and ( w_31336 ,  , w_31337 );
buf ( w_31335 , \12303_b1 );
not ( w_31335 , w_31338 );
not (  , w_31339 );
and ( w_31338 , w_31339 , \12303_b0 );
or ( \12305_b1 , \12304_b1 , w_31340 );
xor ( \12305_b0 , \12304_b0 , w_31342 );
not ( w_31342 , w_31343 );
and ( w_31343 , w_31340 , w_31341 );
buf ( w_31340 , \7105_b1 );
not ( w_31340 , w_31344 );
not ( w_31341 , w_31345 );
and ( w_31344 , w_31345 , \7105_b0 );
or ( \12306_b1 , \12301_b1 , \12305_b1 );
xor ( \12306_b0 , \12301_b0 , w_31346 );
not ( w_31346 , w_31347 );
and ( w_31347 , \12305_b1 , \12305_b0 );
or ( \12307_b1 , \6065_b1 , w_31349 );
not ( w_31349 , w_31350 );
and ( \12307_b0 , \6065_b0 , w_31351 );
and ( w_31350 ,  , w_31351 );
buf ( w_31349 , \7115_b1 );
not ( w_31349 , w_31352 );
not (  , w_31353 );
and ( w_31352 , w_31353 , \7115_b0 );
or ( \12308_b1 , \12307_b1 , w_31354 );
xor ( \12308_b0 , \12307_b0 , w_31356 );
not ( w_31356 , w_31357 );
and ( w_31357 , w_31354 , w_31355 );
buf ( w_31354 , \7123_b1 );
not ( w_31354 , w_31358 );
not ( w_31355 , w_31359 );
and ( w_31358 , w_31359 , \7123_b0 );
or ( \12309_b1 , \12306_b1 , \12308_b1 );
xor ( \12309_b0 , \12306_b0 , w_31360 );
not ( w_31360 , w_31361 );
and ( w_31361 , \12308_b1 , \12308_b0 );
or ( \12310_b1 , \12297_b1 , \12309_b1 );
xor ( \12310_b0 , \12297_b0 , w_31362 );
not ( w_31362 , w_31363 );
and ( w_31363 , \12309_b1 , \12309_b0 );
or ( \12311_b1 , \12263_b1 , \12310_b1 );
not ( \12310_b1 , w_31364 );
and ( \12311_b0 , \12263_b0 , w_31365 );
and ( w_31364 , w_31365 , \12310_b0 );
or ( \12312_b1 , \12238_b1 , \12310_b1 );
not ( \12310_b1 , w_31366 );
and ( \12312_b0 , \12238_b0 , w_31367 );
and ( w_31366 , w_31367 , \12310_b0 );
or ( \12314_b1 , \7123_b1 , \12256_b1 );
not ( \12256_b1 , w_31368 );
and ( \12314_b0 , \7123_b0 , w_31369 );
and ( w_31368 , w_31369 , \12256_b0 );
or ( \12315_b1 , \12256_b1 , \12261_b1 );
not ( \12261_b1 , w_31370 );
and ( \12315_b0 , \12256_b0 , w_31371 );
and ( w_31370 , w_31371 , \12261_b0 );
or ( \12316_b1 , \7123_b1 , \12261_b1 );
not ( \12261_b1 , w_31372 );
and ( \12316_b0 , \7123_b0 , w_31373 );
and ( w_31372 , w_31373 , \12261_b0 );
or ( \12318_b1 , \12242_b1 , \12246_b1 );
not ( \12246_b1 , w_31374 );
and ( \12318_b0 , \12242_b0 , w_31375 );
and ( w_31374 , w_31375 , \12246_b0 );
or ( \12319_b1 , \12246_b1 , \12251_b1 );
not ( \12251_b1 , w_31376 );
and ( \12319_b0 , \12246_b0 , w_31377 );
and ( w_31376 , w_31377 , \12251_b0 );
or ( \12320_b1 , \12242_b1 , \12251_b1 );
not ( \12251_b1 , w_31378 );
and ( \12320_b0 , \12242_b0 , w_31379 );
and ( w_31378 , w_31379 , \12251_b0 );
or ( \12322_b1 , \12317_b1 , \12321_b1 );
xor ( \12322_b0 , \12317_b0 , w_31380 );
not ( w_31380 , w_31381 );
and ( w_31381 , \12321_b1 , \12321_b0 );
or ( \12323_b1 , \12301_b1 , \12305_b1 );
not ( \12305_b1 , w_31382 );
and ( \12323_b0 , \12301_b0 , w_31383 );
and ( w_31382 , w_31383 , \12305_b0 );
or ( \12324_b1 , \12305_b1 , \12308_b1 );
not ( \12308_b1 , w_31384 );
and ( \12324_b0 , \12305_b0 , w_31385 );
and ( w_31384 , w_31385 , \12308_b0 );
or ( \12325_b1 , \12301_b1 , \12308_b1 );
not ( \12308_b1 , w_31386 );
and ( \12325_b0 , \12301_b0 , w_31387 );
and ( w_31386 , w_31387 , \12308_b0 );
or ( \12327_b1 , \12322_b1 , \12326_b1 );
xor ( \12327_b0 , \12322_b0 , w_31388 );
not ( w_31388 , w_31389 );
and ( w_31389 , \12326_b1 , \12326_b0 );
or ( \12328_b1 , \12313_b1 , \12327_b1 );
xor ( \12328_b0 , \12313_b0 , w_31390 );
not ( w_31390 , w_31391 );
and ( w_31391 , \12327_b1 , \12327_b0 );
or ( \12329_b1 , \12280_b1 , \12296_b1 );
not ( \12296_b1 , w_31392 );
and ( \12329_b0 , \12280_b0 , w_31393 );
and ( w_31392 , w_31393 , \12296_b0 );
or ( \12330_b1 , \12296_b1 , \12309_b1 );
not ( \12309_b1 , w_31394 );
and ( \12330_b0 , \12296_b0 , w_31395 );
and ( w_31394 , w_31395 , \12309_b0 );
or ( \12331_b1 , \12280_b1 , \12309_b1 );
not ( \12309_b1 , w_31396 );
and ( \12331_b0 , \12280_b0 , w_31397 );
and ( w_31396 , w_31397 , \12309_b0 );
or ( \12333_b1 , \12252_b1 , \12262_b1 );
not ( \12262_b1 , w_31398 );
and ( \12333_b0 , \12252_b0 , w_31399 );
and ( w_31398 , w_31399 , \12262_b0 );
or ( \12334_b1 , \12332_b1 , \12333_b1 );
xor ( \12334_b0 , \12332_b0 , w_31400 );
not ( w_31400 , w_31401 );
and ( w_31401 , \12333_b1 , \12333_b0 );
or ( \12335_b1 , \6057_b1 , \7099_b1 );
not ( \7099_b1 , w_31402 );
and ( \12335_b0 , \6057_b0 , w_31403 );
and ( w_31402 , w_31403 , \7099_b0 );
or ( \12336_b1 , \6029_b1 , \7097_b1 );
not ( \7097_b1 , w_31404 );
and ( \12336_b0 , \6029_b0 , w_31405 );
and ( w_31404 , w_31405 , \7097_b0 );
or ( \12337_b1 , \12335_b1 , w_31407 );
not ( w_31407 , w_31408 );
and ( \12337_b0 , \12335_b0 , w_31409 );
and ( w_31408 ,  , w_31409 );
buf ( w_31407 , \12336_b1 );
not ( w_31407 , w_31410 );
not (  , w_31411 );
and ( w_31410 , w_31411 , \12336_b0 );
or ( \12338_b1 , \12337_b1 , w_31412 );
xor ( \12338_b0 , \12337_b0 , w_31414 );
not ( w_31414 , w_31415 );
and ( w_31415 , w_31412 , w_31413 );
buf ( w_31412 , \7105_b1 );
not ( w_31412 , w_31416 );
not ( w_31413 , w_31417 );
and ( w_31416 , w_31417 , \7105_b0 );
or ( \12339_b1 , \6065_b1 , \7117_b1 );
not ( \7117_b1 , w_31418 );
and ( \12339_b0 , \6065_b0 , w_31419 );
and ( w_31418 , w_31419 , \7117_b0 );
or ( \12340_b1 , \6048_b1 , \7115_b1 );
not ( \7115_b1 , w_31420 );
and ( \12340_b0 , \6048_b0 , w_31421 );
and ( w_31420 , w_31421 , \7115_b0 );
or ( \12341_b1 , \12339_b1 , w_31423 );
not ( w_31423 , w_31424 );
and ( \12341_b0 , \12339_b0 , w_31425 );
and ( w_31424 ,  , w_31425 );
buf ( w_31423 , \12340_b1 );
not ( w_31423 , w_31426 );
not (  , w_31427 );
and ( w_31426 , w_31427 , \12340_b0 );
or ( \12342_b1 , \12341_b1 , w_31428 );
xor ( \12342_b0 , \12341_b0 , w_31430 );
not ( w_31430 , w_31431 );
and ( w_31431 , w_31428 , w_31429 );
buf ( w_31428 , \7123_b1 );
not ( w_31428 , w_31432 );
not ( w_31429 , w_31433 );
and ( w_31432 , w_31433 , \7123_b0 );
or ( \12343_b1 , \12338_b1 , \12342_b1 );
xor ( \12343_b0 , \12338_b0 , w_31434 );
not ( w_31434 , w_31435 );
and ( w_31435 , \12342_b1 , \12342_b0 );
or ( \12344_b1 , \5998_b1 , \7043_b1 );
not ( \7043_b1 , w_31436 );
and ( \12344_b0 , \5998_b0 , w_31437 );
and ( w_31436 , w_31437 , \7043_b0 );
or ( \12345_b1 , \5967_b1 , \7041_b1 );
not ( \7041_b1 , w_31438 );
and ( \12345_b0 , \5967_b0 , w_31439 );
and ( w_31438 , w_31439 , \7041_b0 );
or ( \12346_b1 , \12344_b1 , w_31441 );
not ( w_31441 , w_31442 );
and ( \12346_b0 , \12344_b0 , w_31443 );
and ( w_31442 ,  , w_31443 );
buf ( w_31441 , \12345_b1 );
not ( w_31441 , w_31444 );
not (  , w_31445 );
and ( w_31444 , w_31445 , \12345_b0 );
or ( \12347_b1 , \12346_b1 , w_31446 );
xor ( \12347_b0 , \12346_b0 , w_31448 );
not ( w_31448 , w_31449 );
and ( w_31449 , w_31446 , w_31447 );
buf ( w_31446 , \7049_b1 );
not ( w_31446 , w_31450 );
not ( w_31447 , w_31451 );
and ( w_31450 , w_31451 , \7049_b0 );
or ( \12348_b1 , \6018_b1 , \7061_b1 );
not ( \7061_b1 , w_31452 );
and ( \12348_b0 , \6018_b0 , w_31453 );
and ( w_31452 , w_31453 , \7061_b0 );
or ( \12349_b1 , \5986_b1 , \7059_b1 );
not ( \7059_b1 , w_31454 );
and ( \12349_b0 , \5986_b0 , w_31455 );
and ( w_31454 , w_31455 , \7059_b0 );
or ( \12350_b1 , \12348_b1 , w_31457 );
not ( w_31457 , w_31458 );
and ( \12350_b0 , \12348_b0 , w_31459 );
and ( w_31458 ,  , w_31459 );
buf ( w_31457 , \12349_b1 );
not ( w_31457 , w_31460 );
not (  , w_31461 );
and ( w_31460 , w_31461 , \12349_b0 );
or ( \12351_b1 , \12350_b1 , w_31462 );
xor ( \12351_b0 , \12350_b0 , w_31464 );
not ( w_31464 , w_31465 );
and ( w_31465 , w_31462 , w_31463 );
buf ( w_31462 , \7067_b1 );
not ( w_31462 , w_31466 );
not ( w_31463 , w_31467 );
and ( w_31466 , w_31467 , \7067_b0 );
or ( \12352_b1 , \12347_b1 , \12351_b1 );
xor ( \12352_b0 , \12347_b0 , w_31468 );
not ( w_31468 , w_31469 );
and ( w_31469 , \12351_b1 , \12351_b0 );
or ( \12353_b1 , \6041_b1 , \7082_b1 );
not ( \7082_b1 , w_31470 );
and ( \12353_b0 , \6041_b0 , w_31471 );
and ( w_31470 , w_31471 , \7082_b0 );
or ( \12354_b1 , \6006_b1 , \7080_b1 );
not ( \7080_b1 , w_31472 );
and ( \12354_b0 , \6006_b0 , w_31473 );
and ( w_31472 , w_31473 , \7080_b0 );
or ( \12355_b1 , \12353_b1 , w_31475 );
not ( w_31475 , w_31476 );
and ( \12355_b0 , \12353_b0 , w_31477 );
and ( w_31476 ,  , w_31477 );
buf ( w_31475 , \12354_b1 );
not ( w_31475 , w_31478 );
not (  , w_31479 );
and ( w_31478 , w_31479 , \12354_b0 );
or ( \12356_b1 , \12355_b1 , w_31480 );
xor ( \12356_b0 , \12355_b0 , w_31482 );
not ( w_31482 , w_31483 );
and ( w_31483 , w_31480 , w_31481 );
buf ( w_31480 , \7088_b1 );
not ( w_31480 , w_31484 );
not ( w_31481 , w_31485 );
and ( w_31484 , w_31485 , \7088_b0 );
or ( \12357_b1 , \12352_b1 , \12356_b1 );
xor ( \12357_b0 , \12352_b0 , w_31486 );
not ( w_31486 , w_31487 );
and ( w_31487 , \12356_b1 , \12356_b0 );
or ( \12358_b1 , \12343_b1 , \12357_b1 );
xor ( \12358_b0 , \12343_b0 , w_31488 );
not ( w_31488 , w_31489 );
and ( w_31489 , \12357_b1 , \12357_b0 );
or ( \12359_b1 , \5937_b1 , \6991_b1 );
not ( \6991_b1 , w_31490 );
and ( \12359_b0 , \5937_b0 , w_31491 );
and ( w_31490 , w_31491 , \6991_b0 );
or ( \12360_b1 , \5906_b1 , \6988_b1 );
not ( \6988_b1 , w_31492 );
and ( \12360_b0 , \5906_b0 , w_31493 );
and ( w_31492 , w_31493 , \6988_b0 );
or ( \12361_b1 , \12359_b1 , w_31495 );
not ( w_31495 , w_31496 );
and ( \12361_b0 , \12359_b0 , w_31497 );
and ( w_31496 ,  , w_31497 );
buf ( w_31495 , \12360_b1 );
not ( w_31495 , w_31498 );
not (  , w_31499 );
and ( w_31498 , w_31499 , \12360_b0 );
or ( \12362_b1 , \12361_b1 , w_31500 );
xor ( \12362_b0 , \12361_b0 , w_31502 );
not ( w_31502 , w_31503 );
and ( w_31503 , w_31500 , w_31501 );
buf ( w_31500 , \6985_b1 );
not ( w_31500 , w_31504 );
not ( w_31501 , w_31505 );
and ( w_31504 , w_31505 , \6985_b0 );
or ( \12363_b1 , \5957_b1 , \7006_b1 );
not ( \7006_b1 , w_31506 );
and ( \12363_b0 , \5957_b0 , w_31507 );
and ( w_31506 , w_31507 , \7006_b0 );
or ( \12364_b1 , \5925_b1 , \7004_b1 );
not ( \7004_b1 , w_31508 );
and ( \12364_b0 , \5925_b0 , w_31509 );
and ( w_31508 , w_31509 , \7004_b0 );
or ( \12365_b1 , \12363_b1 , w_31511 );
not ( w_31511 , w_31512 );
and ( \12365_b0 , \12363_b0 , w_31513 );
and ( w_31512 ,  , w_31513 );
buf ( w_31511 , \12364_b1 );
not ( w_31511 , w_31514 );
not (  , w_31515 );
and ( w_31514 , w_31515 , \12364_b0 );
or ( \12366_b1 , \12365_b1 , w_31516 );
xor ( \12366_b0 , \12365_b0 , w_31518 );
not ( w_31518 , w_31519 );
and ( w_31519 , w_31516 , w_31517 );
buf ( w_31516 , \7012_b1 );
not ( w_31516 , w_31520 );
not ( w_31517 , w_31521 );
and ( w_31520 , w_31521 , \7012_b0 );
or ( \12367_b1 , \12362_b1 , \12366_b1 );
xor ( \12367_b0 , \12362_b0 , w_31522 );
not ( w_31522 , w_31523 );
and ( w_31523 , \12366_b1 , \12366_b0 );
or ( \12368_b1 , \5979_b1 , \7026_b1 );
not ( \7026_b1 , w_31524 );
and ( \12368_b0 , \5979_b0 , w_31525 );
and ( w_31524 , w_31525 , \7026_b0 );
or ( \12369_b1 , \5945_b1 , \7024_b1 );
not ( \7024_b1 , w_31526 );
and ( \12369_b0 , \5945_b0 , w_31527 );
and ( w_31526 , w_31527 , \7024_b0 );
or ( \12370_b1 , \12368_b1 , w_31529 );
not ( w_31529 , w_31530 );
and ( \12370_b0 , \12368_b0 , w_31531 );
and ( w_31530 ,  , w_31531 );
buf ( w_31529 , \12369_b1 );
not ( w_31529 , w_31532 );
not (  , w_31533 );
and ( w_31532 , w_31533 , \12369_b0 );
or ( \12371_b1 , \12370_b1 , w_31534 );
xor ( \12371_b0 , \12370_b0 , w_31536 );
not ( w_31536 , w_31537 );
and ( w_31537 , w_31534 , w_31535 );
buf ( w_31534 , \7032_b1 );
not ( w_31534 , w_31538 );
not ( w_31535 , w_31539 );
and ( w_31538 , w_31539 , \7032_b0 );
or ( \12372_b1 , \12367_b1 , \12371_b1 );
xor ( \12372_b0 , \12367_b0 , w_31540 );
not ( w_31540 , w_31541 );
and ( w_31541 , \12371_b1 , \12371_b0 );
or ( \12373_b1 , \12358_b1 , \12372_b1 );
xor ( \12373_b0 , \12358_b0 , w_31542 );
not ( w_31542 , w_31543 );
and ( w_31543 , \12372_b1 , \12372_b0 );
or ( \12374_b1 , \12334_b1 , \12373_b1 );
xor ( \12374_b0 , \12334_b0 , w_31544 );
not ( w_31544 , w_31545 );
and ( w_31545 , \12373_b1 , \12373_b0 );
or ( \12375_b1 , \12328_b1 , \12374_b1 );
xor ( \12375_b0 , \12328_b0 , w_31546 );
not ( w_31546 , w_31547 );
and ( w_31547 , \12374_b1 , \12374_b0 );
or ( \12376_b1 , \5979_b1 , \6991_b1 );
not ( \6991_b1 , w_31548 );
and ( \12376_b0 , \5979_b0 , w_31549 );
and ( w_31548 , w_31549 , \6991_b0 );
or ( \12377_b1 , \5945_b1 , \6988_b1 );
not ( \6988_b1 , w_31550 );
and ( \12377_b0 , \5945_b0 , w_31551 );
and ( w_31550 , w_31551 , \6988_b0 );
or ( \12378_b1 , \12376_b1 , w_31553 );
not ( w_31553 , w_31554 );
and ( \12378_b0 , \12376_b0 , w_31555 );
and ( w_31554 ,  , w_31555 );
buf ( w_31553 , \12377_b1 );
not ( w_31553 , w_31556 );
not (  , w_31557 );
and ( w_31556 , w_31557 , \12377_b0 );
or ( \12379_b1 , \12378_b1 , w_31558 );
xor ( \12379_b0 , \12378_b0 , w_31560 );
not ( w_31560 , w_31561 );
and ( w_31561 , w_31558 , w_31559 );
buf ( w_31558 , \6985_b1 );
not ( w_31558 , w_31562 );
not ( w_31559 , w_31563 );
and ( w_31562 , w_31563 , \6985_b0 );
or ( \12380_b1 , \5998_b1 , \7006_b1 );
not ( \7006_b1 , w_31564 );
and ( \12380_b0 , \5998_b0 , w_31565 );
and ( w_31564 , w_31565 , \7006_b0 );
or ( \12381_b1 , \5967_b1 , \7004_b1 );
not ( \7004_b1 , w_31566 );
and ( \12381_b0 , \5967_b0 , w_31567 );
and ( w_31566 , w_31567 , \7004_b0 );
or ( \12382_b1 , \12380_b1 , w_31569 );
not ( w_31569 , w_31570 );
and ( \12382_b0 , \12380_b0 , w_31571 );
and ( w_31570 ,  , w_31571 );
buf ( w_31569 , \12381_b1 );
not ( w_31569 , w_31572 );
not (  , w_31573 );
and ( w_31572 , w_31573 , \12381_b0 );
or ( \12383_b1 , \12382_b1 , w_31574 );
xor ( \12383_b0 , \12382_b0 , w_31576 );
not ( w_31576 , w_31577 );
and ( w_31577 , w_31574 , w_31575 );
buf ( w_31574 , \7012_b1 );
not ( w_31574 , w_31578 );
not ( w_31575 , w_31579 );
and ( w_31578 , w_31579 , \7012_b0 );
or ( \12384_b1 , \12379_b1 , \12383_b1 );
not ( \12383_b1 , w_31580 );
and ( \12384_b0 , \12379_b0 , w_31581 );
and ( w_31580 , w_31581 , \12383_b0 );
or ( \12385_b1 , \6018_b1 , \7026_b1 );
not ( \7026_b1 , w_31582 );
and ( \12385_b0 , \6018_b0 , w_31583 );
and ( w_31582 , w_31583 , \7026_b0 );
or ( \12386_b1 , \5986_b1 , \7024_b1 );
not ( \7024_b1 , w_31584 );
and ( \12386_b0 , \5986_b0 , w_31585 );
and ( w_31584 , w_31585 , \7024_b0 );
or ( \12387_b1 , \12385_b1 , w_31587 );
not ( w_31587 , w_31588 );
and ( \12387_b0 , \12385_b0 , w_31589 );
and ( w_31588 ,  , w_31589 );
buf ( w_31587 , \12386_b1 );
not ( w_31587 , w_31590 );
not (  , w_31591 );
and ( w_31590 , w_31591 , \12386_b0 );
or ( \12388_b1 , \12387_b1 , w_31592 );
xor ( \12388_b0 , \12387_b0 , w_31594 );
not ( w_31594 , w_31595 );
and ( w_31595 , w_31592 , w_31593 );
buf ( w_31592 , \7032_b1 );
not ( w_31592 , w_31596 );
not ( w_31593 , w_31597 );
and ( w_31596 , w_31597 , \7032_b0 );
or ( \12389_b1 , \12383_b1 , \12388_b1 );
not ( \12388_b1 , w_31598 );
and ( \12389_b0 , \12383_b0 , w_31599 );
and ( w_31598 , w_31599 , \12388_b0 );
or ( \12390_b1 , \12379_b1 , \12388_b1 );
not ( \12388_b1 , w_31600 );
and ( \12390_b0 , \12379_b0 , w_31601 );
and ( w_31600 , w_31601 , \12388_b0 );
or ( \12392_b1 , \6041_b1 , \7043_b1 );
not ( \7043_b1 , w_31602 );
and ( \12392_b0 , \6041_b0 , w_31603 );
and ( w_31602 , w_31603 , \7043_b0 );
or ( \12393_b1 , \6006_b1 , \7041_b1 );
not ( \7041_b1 , w_31604 );
and ( \12393_b0 , \6006_b0 , w_31605 );
and ( w_31604 , w_31605 , \7041_b0 );
or ( \12394_b1 , \12392_b1 , w_31607 );
not ( w_31607 , w_31608 );
and ( \12394_b0 , \12392_b0 , w_31609 );
and ( w_31608 ,  , w_31609 );
buf ( w_31607 , \12393_b1 );
not ( w_31607 , w_31610 );
not (  , w_31611 );
and ( w_31610 , w_31611 , \12393_b0 );
or ( \12395_b1 , \12394_b1 , w_31612 );
xor ( \12395_b0 , \12394_b0 , w_31614 );
not ( w_31614 , w_31615 );
and ( w_31615 , w_31612 , w_31613 );
buf ( w_31612 , \7049_b1 );
not ( w_31612 , w_31616 );
not ( w_31613 , w_31617 );
and ( w_31616 , w_31617 , \7049_b0 );
or ( \12396_b1 , \6057_b1 , \7061_b1 );
not ( \7061_b1 , w_31618 );
and ( \12396_b0 , \6057_b0 , w_31619 );
and ( w_31618 , w_31619 , \7061_b0 );
or ( \12397_b1 , \6029_b1 , \7059_b1 );
not ( \7059_b1 , w_31620 );
and ( \12397_b0 , \6029_b0 , w_31621 );
and ( w_31620 , w_31621 , \7059_b0 );
or ( \12398_b1 , \12396_b1 , w_31623 );
not ( w_31623 , w_31624 );
and ( \12398_b0 , \12396_b0 , w_31625 );
and ( w_31624 ,  , w_31625 );
buf ( w_31623 , \12397_b1 );
not ( w_31623 , w_31626 );
not (  , w_31627 );
and ( w_31626 , w_31627 , \12397_b0 );
or ( \12399_b1 , \12398_b1 , w_31628 );
xor ( \12399_b0 , \12398_b0 , w_31630 );
not ( w_31630 , w_31631 );
and ( w_31631 , w_31628 , w_31629 );
buf ( w_31628 , \7067_b1 );
not ( w_31628 , w_31632 );
not ( w_31629 , w_31633 );
and ( w_31632 , w_31633 , \7067_b0 );
or ( \12400_b1 , \12395_b1 , \12399_b1 );
not ( \12399_b1 , w_31634 );
and ( \12400_b0 , \12395_b0 , w_31635 );
and ( w_31634 , w_31635 , \12399_b0 );
or ( \12401_b1 , \6065_b1 , \7082_b1 );
not ( \7082_b1 , w_31636 );
and ( \12401_b0 , \6065_b0 , w_31637 );
and ( w_31636 , w_31637 , \7082_b0 );
or ( \12402_b1 , \6048_b1 , \7080_b1 );
not ( \7080_b1 , w_31638 );
and ( \12402_b0 , \6048_b0 , w_31639 );
and ( w_31638 , w_31639 , \7080_b0 );
or ( \12403_b1 , \12401_b1 , w_31641 );
not ( w_31641 , w_31642 );
and ( \12403_b0 , \12401_b0 , w_31643 );
and ( w_31642 ,  , w_31643 );
buf ( w_31641 , \12402_b1 );
not ( w_31641 , w_31644 );
not (  , w_31645 );
and ( w_31644 , w_31645 , \12402_b0 );
or ( \12404_b1 , \12403_b1 , w_31646 );
xor ( \12404_b0 , \12403_b0 , w_31648 );
not ( w_31648 , w_31649 );
and ( w_31649 , w_31646 , w_31647 );
buf ( w_31646 , \7088_b1 );
not ( w_31646 , w_31650 );
not ( w_31647 , w_31651 );
and ( w_31650 , w_31651 , \7088_b0 );
or ( \12405_b1 , \12399_b1 , \12404_b1 );
not ( \12404_b1 , w_31652 );
and ( \12405_b0 , \12399_b0 , w_31653 );
and ( w_31652 , w_31653 , \12404_b0 );
or ( \12406_b1 , \12395_b1 , \12404_b1 );
not ( \12404_b1 , w_31654 );
and ( \12406_b0 , \12395_b0 , w_31655 );
and ( w_31654 , w_31655 , \12404_b0 );
or ( \12408_b1 , \12391_b1 , \12407_b1 );
not ( \12407_b1 , w_31656 );
and ( \12408_b0 , \12391_b0 , w_31657 );
and ( w_31656 , w_31657 , \12407_b0 );
or ( \12409_b1 , \6048_b1 , \7082_b1 );
not ( \7082_b1 , w_31658 );
and ( \12409_b0 , \6048_b0 , w_31659 );
and ( w_31658 , w_31659 , \7082_b0 );
or ( \12410_b1 , \6057_b1 , \7080_b1 );
not ( \7080_b1 , w_31660 );
and ( \12410_b0 , \6057_b0 , w_31661 );
and ( w_31660 , w_31661 , \7080_b0 );
or ( \12411_b1 , \12409_b1 , w_31663 );
not ( w_31663 , w_31664 );
and ( \12411_b0 , \12409_b0 , w_31665 );
and ( w_31664 ,  , w_31665 );
buf ( w_31663 , \12410_b1 );
not ( w_31663 , w_31666 );
not (  , w_31667 );
and ( w_31666 , w_31667 , \12410_b0 );
or ( \12412_b1 , \12411_b1 , w_31668 );
xor ( \12412_b0 , \12411_b0 , w_31670 );
not ( w_31670 , w_31671 );
and ( w_31671 , w_31668 , w_31669 );
buf ( w_31668 , \7088_b1 );
not ( w_31668 , w_31672 );
not ( w_31669 , w_31673 );
and ( w_31672 , w_31673 , \7088_b0 );
or ( \12413_b1 , \12407_b1 , \12412_b1 );
not ( \12412_b1 , w_31674 );
and ( \12413_b0 , \12407_b0 , w_31675 );
and ( w_31674 , w_31675 , \12412_b0 );
or ( \12414_b1 , \12391_b1 , \12412_b1 );
not ( \12412_b1 , w_31676 );
and ( \12414_b0 , \12391_b0 , w_31677 );
and ( w_31676 , w_31677 , \12412_b0 );
or ( \12416_b1 , \6065_b1 , w_31679 );
not ( w_31679 , w_31680 );
and ( \12416_b0 , \6065_b0 , w_31681 );
and ( w_31680 ,  , w_31681 );
buf ( w_31679 , \7097_b1 );
not ( w_31679 , w_31682 );
not (  , w_31683 );
and ( w_31682 , w_31683 , \7097_b0 );
or ( \12417_b1 , \12416_b1 , w_31684 );
xor ( \12417_b0 , \12416_b0 , w_31686 );
not ( w_31686 , w_31687 );
and ( w_31687 , w_31684 , w_31685 );
buf ( w_31684 , \7105_b1 );
not ( w_31684 , w_31688 );
not ( w_31685 , w_31689 );
and ( w_31688 , w_31689 , \7105_b0 );
or ( \12418_b1 , \12218_b1 , \12222_b1 );
xor ( \12418_b0 , \12218_b0 , w_31690 );
not ( w_31690 , w_31691 );
and ( w_31691 , \12222_b1 , \12222_b0 );
or ( \12419_b1 , \12418_b1 , \12227_b1 );
xor ( \12419_b0 , \12418_b0 , w_31692 );
not ( w_31692 , w_31693 );
and ( w_31693 , \12227_b1 , \12227_b0 );
or ( \12420_b1 , \12417_b1 , \12419_b1 );
not ( \12419_b1 , w_31694 );
and ( \12420_b0 , \12417_b0 , w_31695 );
and ( w_31694 , w_31695 , \12419_b0 );
or ( \12421_b1 , \7105_b1 , \12206_b1 );
xor ( \12421_b0 , \7105_b0 , w_31696 );
not ( w_31696 , w_31697 );
and ( w_31697 , \12206_b1 , \12206_b0 );
or ( \12422_b1 , \12421_b1 , \12211_b1 );
xor ( \12422_b0 , \12421_b0 , w_31698 );
not ( w_31698 , w_31699 );
and ( w_31699 , \12211_b1 , \12211_b0 );
or ( \12423_b1 , \12419_b1 , \12422_b1 );
not ( \12422_b1 , w_31700 );
and ( \12423_b0 , \12419_b0 , w_31701 );
and ( w_31700 , w_31701 , \12422_b0 );
or ( \12424_b1 , \12417_b1 , \12422_b1 );
not ( \12422_b1 , w_31702 );
and ( \12424_b0 , \12417_b0 , w_31703 );
and ( w_31702 , w_31703 , \12422_b0 );
or ( \12426_b1 , \12415_b1 , \12425_b1 );
not ( \12425_b1 , w_31704 );
and ( \12426_b0 , \12415_b0 , w_31705 );
and ( w_31704 , w_31705 , \12425_b0 );
or ( \12427_b1 , \12284_b1 , \12288_b1 );
xor ( \12427_b0 , \12284_b0 , w_31706 );
not ( w_31706 , w_31707 );
and ( w_31707 , \12288_b1 , \12288_b0 );
or ( \12428_b1 , \12427_b1 , \12293_b1 );
xor ( \12428_b0 , \12427_b0 , w_31708 );
not ( w_31708 , w_31709 );
and ( w_31709 , \12293_b1 , \12293_b0 );
or ( \12429_b1 , \12425_b1 , \12428_b1 );
not ( \12428_b1 , w_31710 );
and ( \12429_b0 , \12425_b0 , w_31711 );
and ( w_31710 , w_31711 , \12428_b0 );
or ( \12430_b1 , \12415_b1 , \12428_b1 );
not ( \12428_b1 , w_31712 );
and ( \12430_b0 , \12415_b0 , w_31713 );
and ( w_31712 , w_31713 , \12428_b0 );
or ( \12432_b1 , \12268_b1 , \12272_b1 );
xor ( \12432_b0 , \12268_b0 , w_31714 );
not ( w_31714 , w_31715 );
and ( w_31715 , \12272_b1 , \12272_b0 );
or ( \12433_b1 , \12432_b1 , \12277_b1 );
xor ( \12433_b0 , \12432_b0 , w_31716 );
not ( w_31716 , w_31717 );
and ( w_31717 , \12277_b1 , \12277_b0 );
or ( \12434_b1 , \12214_b1 , \12230_b1 );
xor ( \12434_b0 , \12214_b0 , w_31718 );
not ( w_31718 , w_31719 );
and ( w_31719 , \12230_b1 , \12230_b0 );
or ( \12435_b1 , \12434_b1 , \12235_b1 );
xor ( \12435_b0 , \12434_b0 , w_31720 );
not ( w_31720 , w_31721 );
and ( w_31721 , \12235_b1 , \12235_b0 );
or ( \12436_b1 , \12433_b1 , \12435_b1 );
not ( \12435_b1 , w_31722 );
and ( \12436_b0 , \12433_b0 , w_31723 );
and ( w_31722 , w_31723 , \12435_b0 );
or ( \12437_b1 , \12431_b1 , \12436_b1 );
not ( \12436_b1 , w_31724 );
and ( \12437_b0 , \12431_b0 , w_31725 );
and ( w_31724 , w_31725 , \12436_b0 );
or ( \12438_b1 , \12238_b1 , \12263_b1 );
xor ( \12438_b0 , \12238_b0 , w_31726 );
not ( w_31726 , w_31727 );
and ( w_31727 , \12263_b1 , \12263_b0 );
or ( \12439_b1 , \12438_b1 , \12310_b1 );
xor ( \12439_b0 , \12438_b0 , w_31728 );
not ( w_31728 , w_31729 );
and ( w_31729 , \12310_b1 , \12310_b0 );
or ( \12440_b1 , \12436_b1 , \12439_b1 );
not ( \12439_b1 , w_31730 );
and ( \12440_b0 , \12436_b0 , w_31731 );
and ( w_31730 , w_31731 , \12439_b0 );
or ( \12441_b1 , \12431_b1 , \12439_b1 );
not ( \12439_b1 , w_31732 );
and ( \12441_b0 , \12431_b0 , w_31733 );
and ( w_31732 , w_31733 , \12439_b0 );
or ( \12443_b1 , \12375_b1 , w_31735 );
not ( w_31735 , w_31736 );
and ( \12443_b0 , \12375_b0 , w_31737 );
and ( w_31736 ,  , w_31737 );
buf ( w_31735 , \12442_b1 );
not ( w_31735 , w_31738 );
not (  , w_31739 );
and ( w_31738 , w_31739 , \12442_b0 );
or ( \12444_b1 , \12332_b1 , \12333_b1 );
not ( \12333_b1 , w_31740 );
and ( \12444_b0 , \12332_b0 , w_31741 );
and ( w_31740 , w_31741 , \12333_b0 );
or ( \12445_b1 , \12333_b1 , \12373_b1 );
not ( \12373_b1 , w_31742 );
and ( \12445_b0 , \12333_b0 , w_31743 );
and ( w_31742 , w_31743 , \12373_b0 );
or ( \12446_b1 , \12332_b1 , \12373_b1 );
not ( \12373_b1 , w_31744 );
and ( \12446_b0 , \12332_b0 , w_31745 );
and ( w_31744 , w_31745 , \12373_b0 );
or ( \12448_b1 , \6065_b1 , w_31747 );
not ( w_31747 , w_31748 );
and ( \12448_b0 , \6065_b0 , w_31749 );
and ( w_31748 ,  , w_31749 );
buf ( w_31747 , \7138_b1 );
not ( w_31747 , w_31750 );
not (  , w_31751 );
and ( w_31750 , w_31751 , \7138_b0 );
or ( \12449_b1 , \12448_b1 , w_31752 );
xor ( \12449_b0 , \12448_b0 , w_31754 );
not ( w_31754 , w_31755 );
and ( w_31755 , w_31752 , w_31753 );
buf ( w_31752 , \7146_b1 );
not ( w_31752 , w_31756 );
not ( w_31753 , w_31757 );
and ( w_31756 , w_31757 , \7146_b0 );
or ( \12450_b1 , \6006_b1 , \7082_b1 );
not ( \7082_b1 , w_31758 );
and ( \12450_b0 , \6006_b0 , w_31759 );
and ( w_31758 , w_31759 , \7082_b0 );
or ( \12451_b1 , \6018_b1 , \7080_b1 );
not ( \7080_b1 , w_31760 );
and ( \12451_b0 , \6018_b0 , w_31761 );
and ( w_31760 , w_31761 , \7080_b0 );
or ( \12452_b1 , \12450_b1 , w_31763 );
not ( w_31763 , w_31764 );
and ( \12452_b0 , \12450_b0 , w_31765 );
and ( w_31764 ,  , w_31765 );
buf ( w_31763 , \12451_b1 );
not ( w_31763 , w_31766 );
not (  , w_31767 );
and ( w_31766 , w_31767 , \12451_b0 );
or ( \12453_b1 , \12452_b1 , w_31768 );
xor ( \12453_b0 , \12452_b0 , w_31770 );
not ( w_31770 , w_31771 );
and ( w_31771 , w_31768 , w_31769 );
buf ( w_31768 , \7088_b1 );
not ( w_31768 , w_31772 );
not ( w_31769 , w_31773 );
and ( w_31772 , w_31773 , \7088_b0 );
or ( \12454_b1 , \6029_b1 , \7099_b1 );
not ( \7099_b1 , w_31774 );
and ( \12454_b0 , \6029_b0 , w_31775 );
and ( w_31774 , w_31775 , \7099_b0 );
or ( \12455_b1 , \6041_b1 , \7097_b1 );
not ( \7097_b1 , w_31776 );
and ( \12455_b0 , \6041_b0 , w_31777 );
and ( w_31776 , w_31777 , \7097_b0 );
or ( \12456_b1 , \12454_b1 , w_31779 );
not ( w_31779 , w_31780 );
and ( \12456_b0 , \12454_b0 , w_31781 );
and ( w_31780 ,  , w_31781 );
buf ( w_31779 , \12455_b1 );
not ( w_31779 , w_31782 );
not (  , w_31783 );
and ( w_31782 , w_31783 , \12455_b0 );
or ( \12457_b1 , \12456_b1 , w_31784 );
xor ( \12457_b0 , \12456_b0 , w_31786 );
not ( w_31786 , w_31787 );
and ( w_31787 , w_31784 , w_31785 );
buf ( w_31784 , \7105_b1 );
not ( w_31784 , w_31788 );
not ( w_31785 , w_31789 );
and ( w_31788 , w_31789 , \7105_b0 );
or ( \12458_b1 , \12453_b1 , \12457_b1 );
xor ( \12458_b0 , \12453_b0 , w_31790 );
not ( w_31790 , w_31791 );
and ( w_31791 , \12457_b1 , \12457_b0 );
or ( \12459_b1 , \6048_b1 , \7117_b1 );
not ( \7117_b1 , w_31792 );
and ( \12459_b0 , \6048_b0 , w_31793 );
and ( w_31792 , w_31793 , \7117_b0 );
or ( \12460_b1 , \6057_b1 , \7115_b1 );
not ( \7115_b1 , w_31794 );
and ( \12460_b0 , \6057_b0 , w_31795 );
and ( w_31794 , w_31795 , \7115_b0 );
or ( \12461_b1 , \12459_b1 , w_31797 );
not ( w_31797 , w_31798 );
and ( \12461_b0 , \12459_b0 , w_31799 );
and ( w_31798 ,  , w_31799 );
buf ( w_31797 , \12460_b1 );
not ( w_31797 , w_31800 );
not (  , w_31801 );
and ( w_31800 , w_31801 , \12460_b0 );
or ( \12462_b1 , \12461_b1 , w_31802 );
xor ( \12462_b0 , \12461_b0 , w_31804 );
not ( w_31804 , w_31805 );
and ( w_31805 , w_31802 , w_31803 );
buf ( w_31802 , \7123_b1 );
not ( w_31802 , w_31806 );
not ( w_31803 , w_31807 );
and ( w_31806 , w_31807 , \7123_b0 );
or ( \12463_b1 , \12458_b1 , \12462_b1 );
xor ( \12463_b0 , \12458_b0 , w_31808 );
not ( w_31808 , w_31809 );
and ( w_31809 , \12462_b1 , \12462_b0 );
or ( \12464_b1 , \12449_b1 , \12463_b1 );
xor ( \12464_b0 , \12449_b0 , w_31810 );
not ( w_31810 , w_31811 );
and ( w_31811 , \12463_b1 , \12463_b0 );
or ( \12465_b1 , \5945_b1 , \7026_b1 );
not ( \7026_b1 , w_31812 );
and ( \12465_b0 , \5945_b0 , w_31813 );
and ( w_31812 , w_31813 , \7026_b0 );
or ( \12466_b1 , \5957_b1 , \7024_b1 );
not ( \7024_b1 , w_31814 );
and ( \12466_b0 , \5957_b0 , w_31815 );
and ( w_31814 , w_31815 , \7024_b0 );
or ( \12467_b1 , \12465_b1 , w_31817 );
not ( w_31817 , w_31818 );
and ( \12467_b0 , \12465_b0 , w_31819 );
and ( w_31818 ,  , w_31819 );
buf ( w_31817 , \12466_b1 );
not ( w_31817 , w_31820 );
not (  , w_31821 );
and ( w_31820 , w_31821 , \12466_b0 );
or ( \12468_b1 , \12467_b1 , w_31822 );
xor ( \12468_b0 , \12467_b0 , w_31824 );
not ( w_31824 , w_31825 );
and ( w_31825 , w_31822 , w_31823 );
buf ( w_31822 , \7032_b1 );
not ( w_31822 , w_31826 );
not ( w_31823 , w_31827 );
and ( w_31826 , w_31827 , \7032_b0 );
or ( \12469_b1 , \5967_b1 , \7043_b1 );
not ( \7043_b1 , w_31828 );
and ( \12469_b0 , \5967_b0 , w_31829 );
and ( w_31828 , w_31829 , \7043_b0 );
or ( \12470_b1 , \5979_b1 , \7041_b1 );
not ( \7041_b1 , w_31830 );
and ( \12470_b0 , \5979_b0 , w_31831 );
and ( w_31830 , w_31831 , \7041_b0 );
or ( \12471_b1 , \12469_b1 , w_31833 );
not ( w_31833 , w_31834 );
and ( \12471_b0 , \12469_b0 , w_31835 );
and ( w_31834 ,  , w_31835 );
buf ( w_31833 , \12470_b1 );
not ( w_31833 , w_31836 );
not (  , w_31837 );
and ( w_31836 , w_31837 , \12470_b0 );
or ( \12472_b1 , \12471_b1 , w_31838 );
xor ( \12472_b0 , \12471_b0 , w_31840 );
not ( w_31840 , w_31841 );
and ( w_31841 , w_31838 , w_31839 );
buf ( w_31838 , \7049_b1 );
not ( w_31838 , w_31842 );
not ( w_31839 , w_31843 );
and ( w_31842 , w_31843 , \7049_b0 );
or ( \12473_b1 , \12468_b1 , \12472_b1 );
xor ( \12473_b0 , \12468_b0 , w_31844 );
not ( w_31844 , w_31845 );
and ( w_31845 , \12472_b1 , \12472_b0 );
or ( \12474_b1 , \5986_b1 , \7061_b1 );
not ( \7061_b1 , w_31846 );
and ( \12474_b0 , \5986_b0 , w_31847 );
and ( w_31846 , w_31847 , \7061_b0 );
or ( \12475_b1 , \5998_b1 , \7059_b1 );
not ( \7059_b1 , w_31848 );
and ( \12475_b0 , \5998_b0 , w_31849 );
and ( w_31848 , w_31849 , \7059_b0 );
or ( \12476_b1 , \12474_b1 , w_31851 );
not ( w_31851 , w_31852 );
and ( \12476_b0 , \12474_b0 , w_31853 );
and ( w_31852 ,  , w_31853 );
buf ( w_31851 , \12475_b1 );
not ( w_31851 , w_31854 );
not (  , w_31855 );
and ( w_31854 , w_31855 , \12475_b0 );
or ( \12477_b1 , \12476_b1 , w_31856 );
xor ( \12477_b0 , \12476_b0 , w_31858 );
not ( w_31858 , w_31859 );
and ( w_31859 , w_31856 , w_31857 );
buf ( w_31856 , \7067_b1 );
not ( w_31856 , w_31860 );
not ( w_31857 , w_31861 );
and ( w_31860 , w_31861 , \7067_b0 );
or ( \12478_b1 , \12473_b1 , \12477_b1 );
xor ( \12478_b0 , \12473_b0 , w_31862 );
not ( w_31862 , w_31863 );
and ( w_31863 , \12477_b1 , \12477_b0 );
or ( \12479_b1 , \12464_b1 , \12478_b1 );
xor ( \12479_b0 , \12464_b0 , w_31864 );
not ( w_31864 , w_31865 );
and ( w_31865 , \12478_b1 , \12478_b0 );
or ( \12480_b1 , \12362_b1 , \12366_b1 );
not ( \12366_b1 , w_31866 );
and ( \12480_b0 , \12362_b0 , w_31867 );
and ( w_31866 , w_31867 , \12366_b0 );
or ( \12481_b1 , \12366_b1 , \12371_b1 );
not ( \12371_b1 , w_31868 );
and ( \12481_b0 , \12366_b0 , w_31869 );
and ( w_31868 , w_31869 , \12371_b0 );
or ( \12482_b1 , \12362_b1 , \12371_b1 );
not ( \12371_b1 , w_31870 );
and ( \12482_b0 , \12362_b0 , w_31871 );
and ( w_31870 , w_31871 , \12371_b0 );
or ( \12484_b1 , \12347_b1 , \12351_b1 );
not ( \12351_b1 , w_31872 );
and ( \12484_b0 , \12347_b0 , w_31873 );
and ( w_31872 , w_31873 , \12351_b0 );
or ( \12485_b1 , \12351_b1 , \12356_b1 );
not ( \12356_b1 , w_31874 );
and ( \12485_b0 , \12351_b0 , w_31875 );
and ( w_31874 , w_31875 , \12356_b0 );
or ( \12486_b1 , \12347_b1 , \12356_b1 );
not ( \12356_b1 , w_31876 );
and ( \12486_b0 , \12347_b0 , w_31877 );
and ( w_31876 , w_31877 , \12356_b0 );
or ( \12488_b1 , \12483_b1 , \12487_b1 );
xor ( \12488_b0 , \12483_b0 , w_31878 );
not ( w_31878 , w_31879 );
and ( w_31879 , \12487_b1 , \12487_b0 );
or ( \12489_b1 , \12338_b1 , \12342_b1 );
not ( \12342_b1 , w_31880 );
and ( \12489_b0 , \12338_b0 , w_31881 );
and ( w_31880 , w_31881 , \12342_b0 );
or ( \12490_b1 , \12488_b1 , \12489_b1 );
xor ( \12490_b0 , \12488_b0 , w_31882 );
not ( w_31882 , w_31883 );
and ( w_31883 , \12489_b1 , \12489_b0 );
or ( \12491_b1 , \12479_b1 , \12490_b1 );
xor ( \12491_b0 , \12479_b0 , w_31884 );
not ( w_31884 , w_31885 );
and ( w_31885 , \12490_b1 , \12490_b0 );
or ( \12492_b1 , \12447_b1 , \12491_b1 );
xor ( \12492_b0 , \12447_b0 , w_31886 );
not ( w_31886 , w_31887 );
and ( w_31887 , \12491_b1 , \12491_b0 );
or ( \12493_b1 , \12317_b1 , \12321_b1 );
not ( \12321_b1 , w_31888 );
and ( \12493_b0 , \12317_b0 , w_31889 );
and ( w_31888 , w_31889 , \12321_b0 );
or ( \12494_b1 , \12321_b1 , \12326_b1 );
not ( \12326_b1 , w_31890 );
and ( \12494_b0 , \12321_b0 , w_31891 );
and ( w_31890 , w_31891 , \12326_b0 );
or ( \12495_b1 , \12317_b1 , \12326_b1 );
not ( \12326_b1 , w_31892 );
and ( \12495_b0 , \12317_b0 , w_31893 );
and ( w_31892 , w_31893 , \12326_b0 );
or ( \12497_b1 , \12343_b1 , \12357_b1 );
not ( \12357_b1 , w_31894 );
and ( \12497_b0 , \12343_b0 , w_31895 );
and ( w_31894 , w_31895 , \12357_b0 );
or ( \12498_b1 , \12357_b1 , \12372_b1 );
not ( \12372_b1 , w_31896 );
and ( \12498_b0 , \12357_b0 , w_31897 );
and ( w_31896 , w_31897 , \12372_b0 );
or ( \12499_b1 , \12343_b1 , \12372_b1 );
not ( \12372_b1 , w_31898 );
and ( \12499_b0 , \12343_b0 , w_31899 );
and ( w_31898 , w_31899 , \12372_b0 );
or ( \12501_b1 , \12496_b1 , \12500_b1 );
xor ( \12501_b0 , \12496_b0 , w_31900 );
not ( w_31900 , w_31901 );
and ( w_31901 , \12500_b1 , \12500_b0 );
or ( \12502_b1 , \5906_b1 , \6991_b1 );
not ( \6991_b1 , w_31902 );
and ( \12502_b0 , \5906_b0 , w_31903 );
and ( w_31902 , w_31903 , \6991_b0 );
or ( \12503_b1 , \5918_b1 , \6988_b1 );
not ( \6988_b1 , w_31904 );
and ( \12503_b0 , \5918_b0 , w_31905 );
and ( w_31904 , w_31905 , \6988_b0 );
or ( \12504_b1 , \12502_b1 , w_31907 );
not ( w_31907 , w_31908 );
and ( \12504_b0 , \12502_b0 , w_31909 );
and ( w_31908 ,  , w_31909 );
buf ( w_31907 , \12503_b1 );
not ( w_31907 , w_31910 );
not (  , w_31911 );
and ( w_31910 , w_31911 , \12503_b0 );
or ( \12505_b1 , \12504_b1 , w_31912 );
xor ( \12505_b0 , \12504_b0 , w_31914 );
not ( w_31914 , w_31915 );
and ( w_31915 , w_31912 , w_31913 );
buf ( w_31912 , \6985_b1 );
not ( w_31912 , w_31916 );
not ( w_31913 , w_31917 );
and ( w_31916 , w_31917 , \6985_b0 );
or ( \12506_b1 , \7146_b1 , \12505_b1 );
xor ( \12506_b0 , \7146_b0 , w_31918 );
not ( w_31918 , w_31919 );
and ( w_31919 , \12505_b1 , \12505_b0 );
or ( \12507_b1 , \5925_b1 , \7006_b1 );
not ( \7006_b1 , w_31920 );
and ( \12507_b0 , \5925_b0 , w_31921 );
and ( w_31920 , w_31921 , \7006_b0 );
or ( \12508_b1 , \5937_b1 , \7004_b1 );
not ( \7004_b1 , w_31922 );
and ( \12508_b0 , \5937_b0 , w_31923 );
and ( w_31922 , w_31923 , \7004_b0 );
or ( \12509_b1 , \12507_b1 , w_31925 );
not ( w_31925 , w_31926 );
and ( \12509_b0 , \12507_b0 , w_31927 );
and ( w_31926 ,  , w_31927 );
buf ( w_31925 , \12508_b1 );
not ( w_31925 , w_31928 );
not (  , w_31929 );
and ( w_31928 , w_31929 , \12508_b0 );
or ( \12510_b1 , \12509_b1 , w_31930 );
xor ( \12510_b0 , \12509_b0 , w_31932 );
not ( w_31932 , w_31933 );
and ( w_31933 , w_31930 , w_31931 );
buf ( w_31930 , \7012_b1 );
not ( w_31930 , w_31934 );
not ( w_31931 , w_31935 );
and ( w_31934 , w_31935 , \7012_b0 );
or ( \12511_b1 , \12506_b1 , \12510_b1 );
xor ( \12511_b0 , \12506_b0 , w_31936 );
not ( w_31936 , w_31937 );
and ( w_31937 , \12510_b1 , \12510_b0 );
or ( \12512_b1 , \12501_b1 , \12511_b1 );
xor ( \12512_b0 , \12501_b0 , w_31938 );
not ( w_31938 , w_31939 );
and ( w_31939 , \12511_b1 , \12511_b0 );
or ( \12513_b1 , \12492_b1 , \12512_b1 );
xor ( \12513_b0 , \12492_b0 , w_31940 );
not ( w_31940 , w_31941 );
and ( w_31941 , \12512_b1 , \12512_b0 );
or ( \12514_b1 , \12313_b1 , \12327_b1 );
not ( \12327_b1 , w_31942 );
and ( \12514_b0 , \12313_b0 , w_31943 );
and ( w_31942 , w_31943 , \12327_b0 );
or ( \12515_b1 , \12327_b1 , \12374_b1 );
not ( \12374_b1 , w_31944 );
and ( \12515_b0 , \12327_b0 , w_31945 );
and ( w_31944 , w_31945 , \12374_b0 );
or ( \12516_b1 , \12313_b1 , \12374_b1 );
not ( \12374_b1 , w_31946 );
and ( \12516_b0 , \12313_b0 , w_31947 );
and ( w_31946 , w_31947 , \12374_b0 );
or ( \12518_b1 , \12513_b1 , w_31949 );
not ( w_31949 , w_31950 );
and ( \12518_b0 , \12513_b0 , w_31951 );
and ( w_31950 ,  , w_31951 );
buf ( w_31949 , \12517_b1 );
not ( w_31949 , w_31952 );
not (  , w_31953 );
and ( w_31952 , w_31953 , \12517_b0 );
or ( \12519_b1 , \12443_b1 , w_31955 );
not ( w_31955 , w_31956 );
and ( \12519_b0 , \12443_b0 , w_31957 );
and ( w_31956 ,  , w_31957 );
buf ( w_31955 , \12518_b1 );
not ( w_31955 , w_31958 );
not (  , w_31959 );
and ( w_31958 , w_31959 , \12518_b0 );
or ( \12520_b1 , \12483_b1 , \12487_b1 );
not ( \12487_b1 , w_31960 );
and ( \12520_b0 , \12483_b0 , w_31961 );
and ( w_31960 , w_31961 , \12487_b0 );
or ( \12521_b1 , \12487_b1 , \12489_b1 );
not ( \12489_b1 , w_31962 );
and ( \12521_b0 , \12487_b0 , w_31963 );
and ( w_31962 , w_31963 , \12489_b0 );
or ( \12522_b1 , \12483_b1 , \12489_b1 );
not ( \12489_b1 , w_31964 );
and ( \12522_b0 , \12483_b0 , w_31965 );
and ( w_31964 , w_31965 , \12489_b0 );
or ( \12524_b1 , \12449_b1 , \12463_b1 );
not ( \12463_b1 , w_31966 );
and ( \12524_b0 , \12449_b0 , w_31967 );
and ( w_31966 , w_31967 , \12463_b0 );
or ( \12525_b1 , \12463_b1 , \12478_b1 );
not ( \12478_b1 , w_31968 );
and ( \12525_b0 , \12463_b0 , w_31969 );
and ( w_31968 , w_31969 , \12478_b0 );
or ( \12526_b1 , \12449_b1 , \12478_b1 );
not ( \12478_b1 , w_31970 );
and ( \12526_b0 , \12449_b0 , w_31971 );
and ( w_31970 , w_31971 , \12478_b0 );
or ( \12528_b1 , \12523_b1 , \12527_b1 );
xor ( \12528_b0 , \12523_b0 , w_31972 );
not ( w_31972 , w_31973 );
and ( w_31973 , \12527_b1 , \12527_b0 );
or ( \12529_b1 , \6041_b1 , \7099_b1 );
not ( \7099_b1 , w_31974 );
and ( \12529_b0 , \6041_b0 , w_31975 );
and ( w_31974 , w_31975 , \7099_b0 );
or ( \12530_b1 , \6006_b1 , \7097_b1 );
not ( \7097_b1 , w_31976 );
and ( \12530_b0 , \6006_b0 , w_31977 );
and ( w_31976 , w_31977 , \7097_b0 );
or ( \12531_b1 , \12529_b1 , w_31979 );
not ( w_31979 , w_31980 );
and ( \12531_b0 , \12529_b0 , w_31981 );
and ( w_31980 ,  , w_31981 );
buf ( w_31979 , \12530_b1 );
not ( w_31979 , w_31982 );
not (  , w_31983 );
and ( w_31982 , w_31983 , \12530_b0 );
or ( \12532_b1 , \12531_b1 , w_31984 );
xor ( \12532_b0 , \12531_b0 , w_31986 );
not ( w_31986 , w_31987 );
and ( w_31987 , w_31984 , w_31985 );
buf ( w_31984 , \7105_b1 );
not ( w_31984 , w_31988 );
not ( w_31985 , w_31989 );
and ( w_31988 , w_31989 , \7105_b0 );
or ( \12533_b1 , \6057_b1 , \7117_b1 );
not ( \7117_b1 , w_31990 );
and ( \12533_b0 , \6057_b0 , w_31991 );
and ( w_31990 , w_31991 , \7117_b0 );
or ( \12534_b1 , \6029_b1 , \7115_b1 );
not ( \7115_b1 , w_31992 );
and ( \12534_b0 , \6029_b0 , w_31993 );
and ( w_31992 , w_31993 , \7115_b0 );
or ( \12535_b1 , \12533_b1 , w_31995 );
not ( w_31995 , w_31996 );
and ( \12535_b0 , \12533_b0 , w_31997 );
and ( w_31996 ,  , w_31997 );
buf ( w_31995 , \12534_b1 );
not ( w_31995 , w_31998 );
not (  , w_31999 );
and ( w_31998 , w_31999 , \12534_b0 );
or ( \12536_b1 , \12535_b1 , w_32000 );
xor ( \12536_b0 , \12535_b0 , w_32002 );
not ( w_32002 , w_32003 );
and ( w_32003 , w_32000 , w_32001 );
buf ( w_32000 , \7123_b1 );
not ( w_32000 , w_32004 );
not ( w_32001 , w_32005 );
and ( w_32004 , w_32005 , \7123_b0 );
or ( \12537_b1 , \12532_b1 , \12536_b1 );
xor ( \12537_b0 , \12532_b0 , w_32006 );
not ( w_32006 , w_32007 );
and ( w_32007 , \12536_b1 , \12536_b0 );
or ( \12538_b1 , \6065_b1 , \7140_b1 );
not ( \7140_b1 , w_32008 );
and ( \12538_b0 , \6065_b0 , w_32009 );
and ( w_32008 , w_32009 , \7140_b0 );
or ( \12539_b1 , \6048_b1 , \7138_b1 );
not ( \7138_b1 , w_32010 );
and ( \12539_b0 , \6048_b0 , w_32011 );
and ( w_32010 , w_32011 , \7138_b0 );
or ( \12540_b1 , \12538_b1 , w_32013 );
not ( w_32013 , w_32014 );
and ( \12540_b0 , \12538_b0 , w_32015 );
and ( w_32014 ,  , w_32015 );
buf ( w_32013 , \12539_b1 );
not ( w_32013 , w_32016 );
not (  , w_32017 );
and ( w_32016 , w_32017 , \12539_b0 );
or ( \12541_b1 , \12540_b1 , w_32018 );
xor ( \12541_b0 , \12540_b0 , w_32020 );
not ( w_32020 , w_32021 );
and ( w_32021 , w_32018 , w_32019 );
buf ( w_32018 , \7146_b1 );
not ( w_32018 , w_32022 );
not ( w_32019 , w_32023 );
and ( w_32022 , w_32023 , \7146_b0 );
or ( \12542_b1 , \12537_b1 , \12541_b1 );
xor ( \12542_b0 , \12537_b0 , w_32024 );
not ( w_32024 , w_32025 );
and ( w_32025 , \12541_b1 , \12541_b0 );
or ( \12543_b1 , \5979_b1 , \7043_b1 );
not ( \7043_b1 , w_32026 );
and ( \12543_b0 , \5979_b0 , w_32027 );
and ( w_32026 , w_32027 , \7043_b0 );
or ( \12544_b1 , \5945_b1 , \7041_b1 );
not ( \7041_b1 , w_32028 );
and ( \12544_b0 , \5945_b0 , w_32029 );
and ( w_32028 , w_32029 , \7041_b0 );
or ( \12545_b1 , \12543_b1 , w_32031 );
not ( w_32031 , w_32032 );
and ( \12545_b0 , \12543_b0 , w_32033 );
and ( w_32032 ,  , w_32033 );
buf ( w_32031 , \12544_b1 );
not ( w_32031 , w_32034 );
not (  , w_32035 );
and ( w_32034 , w_32035 , \12544_b0 );
or ( \12546_b1 , \12545_b1 , w_32036 );
xor ( \12546_b0 , \12545_b0 , w_32038 );
not ( w_32038 , w_32039 );
and ( w_32039 , w_32036 , w_32037 );
buf ( w_32036 , \7049_b1 );
not ( w_32036 , w_32040 );
not ( w_32037 , w_32041 );
and ( w_32040 , w_32041 , \7049_b0 );
or ( \12547_b1 , \5998_b1 , \7061_b1 );
not ( \7061_b1 , w_32042 );
and ( \12547_b0 , \5998_b0 , w_32043 );
and ( w_32042 , w_32043 , \7061_b0 );
or ( \12548_b1 , \5967_b1 , \7059_b1 );
not ( \7059_b1 , w_32044 );
and ( \12548_b0 , \5967_b0 , w_32045 );
and ( w_32044 , w_32045 , \7059_b0 );
or ( \12549_b1 , \12547_b1 , w_32047 );
not ( w_32047 , w_32048 );
and ( \12549_b0 , \12547_b0 , w_32049 );
and ( w_32048 ,  , w_32049 );
buf ( w_32047 , \12548_b1 );
not ( w_32047 , w_32050 );
not (  , w_32051 );
and ( w_32050 , w_32051 , \12548_b0 );
or ( \12550_b1 , \12549_b1 , w_32052 );
xor ( \12550_b0 , \12549_b0 , w_32054 );
not ( w_32054 , w_32055 );
and ( w_32055 , w_32052 , w_32053 );
buf ( w_32052 , \7067_b1 );
not ( w_32052 , w_32056 );
not ( w_32053 , w_32057 );
and ( w_32056 , w_32057 , \7067_b0 );
or ( \12551_b1 , \12546_b1 , \12550_b1 );
xor ( \12551_b0 , \12546_b0 , w_32058 );
not ( w_32058 , w_32059 );
and ( w_32059 , \12550_b1 , \12550_b0 );
or ( \12552_b1 , \6018_b1 , \7082_b1 );
not ( \7082_b1 , w_32060 );
and ( \12552_b0 , \6018_b0 , w_32061 );
and ( w_32060 , w_32061 , \7082_b0 );
or ( \12553_b1 , \5986_b1 , \7080_b1 );
not ( \7080_b1 , w_32062 );
and ( \12553_b0 , \5986_b0 , w_32063 );
and ( w_32062 , w_32063 , \7080_b0 );
or ( \12554_b1 , \12552_b1 , w_32065 );
not ( w_32065 , w_32066 );
and ( \12554_b0 , \12552_b0 , w_32067 );
and ( w_32066 ,  , w_32067 );
buf ( w_32065 , \12553_b1 );
not ( w_32065 , w_32068 );
not (  , w_32069 );
and ( w_32068 , w_32069 , \12553_b0 );
or ( \12555_b1 , \12554_b1 , w_32070 );
xor ( \12555_b0 , \12554_b0 , w_32072 );
not ( w_32072 , w_32073 );
and ( w_32073 , w_32070 , w_32071 );
buf ( w_32070 , \7088_b1 );
not ( w_32070 , w_32074 );
not ( w_32071 , w_32075 );
and ( w_32074 , w_32075 , \7088_b0 );
or ( \12556_b1 , \12551_b1 , \12555_b1 );
xor ( \12556_b0 , \12551_b0 , w_32076 );
not ( w_32076 , w_32077 );
and ( w_32077 , \12555_b1 , \12555_b0 );
or ( \12557_b1 , \12542_b1 , \12556_b1 );
xor ( \12557_b0 , \12542_b0 , w_32078 );
not ( w_32078 , w_32079 );
and ( w_32079 , \12556_b1 , \12556_b0 );
or ( \12558_b1 , \5918_b1 , \6991_b1 );
not ( \6991_b1 , w_32080 );
and ( \12558_b0 , \5918_b0 , w_32081 );
and ( w_32080 , w_32081 , \6991_b0 );
or ( \12559_b1 , \5881_b1 , \6988_b1 );
not ( \6988_b1 , w_32082 );
and ( \12559_b0 , \5881_b0 , w_32083 );
and ( w_32082 , w_32083 , \6988_b0 );
or ( \12560_b1 , \12558_b1 , w_32085 );
not ( w_32085 , w_32086 );
and ( \12560_b0 , \12558_b0 , w_32087 );
and ( w_32086 ,  , w_32087 );
buf ( w_32085 , \12559_b1 );
not ( w_32085 , w_32088 );
not (  , w_32089 );
and ( w_32088 , w_32089 , \12559_b0 );
or ( \12561_b1 , \12560_b1 , w_32090 );
xor ( \12561_b0 , \12560_b0 , w_32092 );
not ( w_32092 , w_32093 );
and ( w_32093 , w_32090 , w_32091 );
buf ( w_32090 , \6985_b1 );
not ( w_32090 , w_32094 );
not ( w_32091 , w_32095 );
and ( w_32094 , w_32095 , \6985_b0 );
or ( \12562_b1 , \5937_b1 , \7006_b1 );
not ( \7006_b1 , w_32096 );
and ( \12562_b0 , \5937_b0 , w_32097 );
and ( w_32096 , w_32097 , \7006_b0 );
or ( \12563_b1 , \5906_b1 , \7004_b1 );
not ( \7004_b1 , w_32098 );
and ( \12563_b0 , \5906_b0 , w_32099 );
and ( w_32098 , w_32099 , \7004_b0 );
or ( \12564_b1 , \12562_b1 , w_32101 );
not ( w_32101 , w_32102 );
and ( \12564_b0 , \12562_b0 , w_32103 );
and ( w_32102 ,  , w_32103 );
buf ( w_32101 , \12563_b1 );
not ( w_32101 , w_32104 );
not (  , w_32105 );
and ( w_32104 , w_32105 , \12563_b0 );
or ( \12565_b1 , \12564_b1 , w_32106 );
xor ( \12565_b0 , \12564_b0 , w_32108 );
not ( w_32108 , w_32109 );
and ( w_32109 , w_32106 , w_32107 );
buf ( w_32106 , \7012_b1 );
not ( w_32106 , w_32110 );
not ( w_32107 , w_32111 );
and ( w_32110 , w_32111 , \7012_b0 );
or ( \12566_b1 , \12561_b1 , \12565_b1 );
xor ( \12566_b0 , \12561_b0 , w_32112 );
not ( w_32112 , w_32113 );
and ( w_32113 , \12565_b1 , \12565_b0 );
or ( \12567_b1 , \5957_b1 , \7026_b1 );
not ( \7026_b1 , w_32114 );
and ( \12567_b0 , \5957_b0 , w_32115 );
and ( w_32114 , w_32115 , \7026_b0 );
or ( \12568_b1 , \5925_b1 , \7024_b1 );
not ( \7024_b1 , w_32116 );
and ( \12568_b0 , \5925_b0 , w_32117 );
and ( w_32116 , w_32117 , \7024_b0 );
or ( \12569_b1 , \12567_b1 , w_32119 );
not ( w_32119 , w_32120 );
and ( \12569_b0 , \12567_b0 , w_32121 );
and ( w_32120 ,  , w_32121 );
buf ( w_32119 , \12568_b1 );
not ( w_32119 , w_32122 );
not (  , w_32123 );
and ( w_32122 , w_32123 , \12568_b0 );
or ( \12570_b1 , \12569_b1 , w_32124 );
xor ( \12570_b0 , \12569_b0 , w_32126 );
not ( w_32126 , w_32127 );
and ( w_32127 , w_32124 , w_32125 );
buf ( w_32124 , \7032_b1 );
not ( w_32124 , w_32128 );
not ( w_32125 , w_32129 );
and ( w_32128 , w_32129 , \7032_b0 );
or ( \12571_b1 , \12566_b1 , \12570_b1 );
xor ( \12571_b0 , \12566_b0 , w_32130 );
not ( w_32130 , w_32131 );
and ( w_32131 , \12570_b1 , \12570_b0 );
or ( \12572_b1 , \12557_b1 , \12571_b1 );
xor ( \12572_b0 , \12557_b0 , w_32132 );
not ( w_32132 , w_32133 );
and ( w_32133 , \12571_b1 , \12571_b0 );
or ( \12573_b1 , \12528_b1 , \12572_b1 );
xor ( \12573_b0 , \12528_b0 , w_32134 );
not ( w_32134 , w_32135 );
and ( w_32135 , \12572_b1 , \12572_b0 );
or ( \12574_b1 , \12496_b1 , \12500_b1 );
not ( \12500_b1 , w_32136 );
and ( \12574_b0 , \12496_b0 , w_32137 );
and ( w_32136 , w_32137 , \12500_b0 );
or ( \12575_b1 , \12500_b1 , \12511_b1 );
not ( \12511_b1 , w_32138 );
and ( \12575_b0 , \12500_b0 , w_32139 );
and ( w_32138 , w_32139 , \12511_b0 );
or ( \12576_b1 , \12496_b1 , \12511_b1 );
not ( \12511_b1 , w_32140 );
and ( \12576_b0 , \12496_b0 , w_32141 );
and ( w_32140 , w_32141 , \12511_b0 );
or ( \12578_b1 , \12479_b1 , \12490_b1 );
not ( \12490_b1 , w_32142 );
and ( \12578_b0 , \12479_b0 , w_32143 );
and ( w_32142 , w_32143 , \12490_b0 );
or ( \12579_b1 , \12577_b1 , \12578_b1 );
xor ( \12579_b0 , \12577_b0 , w_32144 );
not ( w_32144 , w_32145 );
and ( w_32145 , \12578_b1 , \12578_b0 );
or ( \12580_b1 , \7146_b1 , \12505_b1 );
not ( \12505_b1 , w_32146 );
and ( \12580_b0 , \7146_b0 , w_32147 );
and ( w_32146 , w_32147 , \12505_b0 );
or ( \12581_b1 , \12505_b1 , \12510_b1 );
not ( \12510_b1 , w_32148 );
and ( \12581_b0 , \12505_b0 , w_32149 );
and ( w_32148 , w_32149 , \12510_b0 );
or ( \12582_b1 , \7146_b1 , \12510_b1 );
not ( \12510_b1 , w_32150 );
and ( \12582_b0 , \7146_b0 , w_32151 );
and ( w_32150 , w_32151 , \12510_b0 );
or ( \12584_b1 , \12468_b1 , \12472_b1 );
not ( \12472_b1 , w_32152 );
and ( \12584_b0 , \12468_b0 , w_32153 );
and ( w_32152 , w_32153 , \12472_b0 );
or ( \12585_b1 , \12472_b1 , \12477_b1 );
not ( \12477_b1 , w_32154 );
and ( \12585_b0 , \12472_b0 , w_32155 );
and ( w_32154 , w_32155 , \12477_b0 );
or ( \12586_b1 , \12468_b1 , \12477_b1 );
not ( \12477_b1 , w_32156 );
and ( \12586_b0 , \12468_b0 , w_32157 );
and ( w_32156 , w_32157 , \12477_b0 );
or ( \12588_b1 , \12583_b1 , \12587_b1 );
xor ( \12588_b0 , \12583_b0 , w_32158 );
not ( w_32158 , w_32159 );
and ( w_32159 , \12587_b1 , \12587_b0 );
or ( \12589_b1 , \12453_b1 , \12457_b1 );
not ( \12457_b1 , w_32160 );
and ( \12589_b0 , \12453_b0 , w_32161 );
and ( w_32160 , w_32161 , \12457_b0 );
or ( \12590_b1 , \12457_b1 , \12462_b1 );
not ( \12462_b1 , w_32162 );
and ( \12590_b0 , \12457_b0 , w_32163 );
and ( w_32162 , w_32163 , \12462_b0 );
or ( \12591_b1 , \12453_b1 , \12462_b1 );
not ( \12462_b1 , w_32164 );
and ( \12591_b0 , \12453_b0 , w_32165 );
and ( w_32164 , w_32165 , \12462_b0 );
or ( \12593_b1 , \12588_b1 , \12592_b1 );
xor ( \12593_b0 , \12588_b0 , w_32166 );
not ( w_32166 , w_32167 );
and ( w_32167 , \12592_b1 , \12592_b0 );
or ( \12594_b1 , \12579_b1 , \12593_b1 );
xor ( \12594_b0 , \12579_b0 , w_32168 );
not ( w_32168 , w_32169 );
and ( w_32169 , \12593_b1 , \12593_b0 );
or ( \12595_b1 , \12573_b1 , \12594_b1 );
xor ( \12595_b0 , \12573_b0 , w_32170 );
not ( w_32170 , w_32171 );
and ( w_32171 , \12594_b1 , \12594_b0 );
or ( \12596_b1 , \12447_b1 , \12491_b1 );
not ( \12491_b1 , w_32172 );
and ( \12596_b0 , \12447_b0 , w_32173 );
and ( w_32172 , w_32173 , \12491_b0 );
or ( \12597_b1 , \12491_b1 , \12512_b1 );
not ( \12512_b1 , w_32174 );
and ( \12597_b0 , \12491_b0 , w_32175 );
and ( w_32174 , w_32175 , \12512_b0 );
or ( \12598_b1 , \12447_b1 , \12512_b1 );
not ( \12512_b1 , w_32176 );
and ( \12598_b0 , \12447_b0 , w_32177 );
and ( w_32176 , w_32177 , \12512_b0 );
or ( \12600_b1 , \12595_b1 , w_32179 );
not ( w_32179 , w_32180 );
and ( \12600_b0 , \12595_b0 , w_32181 );
and ( w_32180 ,  , w_32181 );
buf ( w_32179 , \12599_b1 );
not ( w_32179 , w_32182 );
not (  , w_32183 );
and ( w_32182 , w_32183 , \12599_b0 );
or ( \12601_b1 , \12577_b1 , \12578_b1 );
not ( \12578_b1 , w_32184 );
and ( \12601_b0 , \12577_b0 , w_32185 );
and ( w_32184 , w_32185 , \12578_b0 );
or ( \12602_b1 , \12578_b1 , \12593_b1 );
not ( \12593_b1 , w_32186 );
and ( \12602_b0 , \12578_b0 , w_32187 );
and ( w_32186 , w_32187 , \12593_b0 );
or ( \12603_b1 , \12577_b1 , \12593_b1 );
not ( \12593_b1 , w_32188 );
and ( \12603_b0 , \12577_b0 , w_32189 );
and ( w_32188 , w_32189 , \12593_b0 );
or ( \12605_b1 , \12523_b1 , \12527_b1 );
not ( \12527_b1 , w_32190 );
and ( \12605_b0 , \12523_b0 , w_32191 );
and ( w_32190 , w_32191 , \12527_b0 );
or ( \12606_b1 , \12527_b1 , \12572_b1 );
not ( \12572_b1 , w_32192 );
and ( \12606_b0 , \12527_b0 , w_32193 );
and ( w_32192 , w_32193 , \12572_b0 );
or ( \12607_b1 , \12523_b1 , \12572_b1 );
not ( \12572_b1 , w_32194 );
and ( \12607_b0 , \12523_b0 , w_32195 );
and ( w_32194 , w_32195 , \12572_b0 );
or ( \12609_b1 , \5881_b1 , \6991_b1 );
not ( \6991_b1 , w_32196 );
and ( \12609_b0 , \5881_b0 , w_32197 );
and ( w_32196 , w_32197 , \6991_b0 );
or ( \12610_b1 , \5893_b1 , \6988_b1 );
not ( \6988_b1 , w_32198 );
and ( \12610_b0 , \5893_b0 , w_32199 );
and ( w_32198 , w_32199 , \6988_b0 );
or ( \12611_b1 , \12609_b1 , w_32201 );
not ( w_32201 , w_32202 );
and ( \12611_b0 , \12609_b0 , w_32203 );
and ( w_32202 ,  , w_32203 );
buf ( w_32201 , \12610_b1 );
not ( w_32201 , w_32204 );
not (  , w_32205 );
and ( w_32204 , w_32205 , \12610_b0 );
or ( \12612_b1 , \12611_b1 , w_32206 );
xor ( \12612_b0 , \12611_b0 , w_32208 );
not ( w_32208 , w_32209 );
and ( w_32209 , w_32206 , w_32207 );
buf ( w_32206 , \6985_b1 );
not ( w_32206 , w_32210 );
not ( w_32207 , w_32211 );
and ( w_32210 , w_32211 , \6985_b0 );
or ( \12613_b1 , \7163_b1 , \12612_b1 );
xor ( \12613_b0 , \7163_b0 , w_32212 );
not ( w_32212 , w_32213 );
and ( w_32213 , \12612_b1 , \12612_b0 );
or ( \12614_b1 , \5906_b1 , \7006_b1 );
not ( \7006_b1 , w_32214 );
and ( \12614_b0 , \5906_b0 , w_32215 );
and ( w_32214 , w_32215 , \7006_b0 );
or ( \12615_b1 , \5918_b1 , \7004_b1 );
not ( \7004_b1 , w_32216 );
and ( \12615_b0 , \5918_b0 , w_32217 );
and ( w_32216 , w_32217 , \7004_b0 );
or ( \12616_b1 , \12614_b1 , w_32219 );
not ( w_32219 , w_32220 );
and ( \12616_b0 , \12614_b0 , w_32221 );
and ( w_32220 ,  , w_32221 );
buf ( w_32219 , \12615_b1 );
not ( w_32219 , w_32222 );
not (  , w_32223 );
and ( w_32222 , w_32223 , \12615_b0 );
or ( \12617_b1 , \12616_b1 , w_32224 );
xor ( \12617_b0 , \12616_b0 , w_32226 );
not ( w_32226 , w_32227 );
and ( w_32227 , w_32224 , w_32225 );
buf ( w_32224 , \7012_b1 );
not ( w_32224 , w_32228 );
not ( w_32225 , w_32229 );
and ( w_32228 , w_32229 , \7012_b0 );
or ( \12618_b1 , \12613_b1 , \12617_b1 );
xor ( \12618_b0 , \12613_b0 , w_32230 );
not ( w_32230 , w_32231 );
and ( w_32231 , \12617_b1 , \12617_b0 );
or ( \12619_b1 , \6048_b1 , \7140_b1 );
not ( \7140_b1 , w_32232 );
and ( \12619_b0 , \6048_b0 , w_32233 );
and ( w_32232 , w_32233 , \7140_b0 );
or ( \12620_b1 , \6057_b1 , \7138_b1 );
not ( \7138_b1 , w_32234 );
and ( \12620_b0 , \6057_b0 , w_32235 );
and ( w_32234 , w_32235 , \7138_b0 );
or ( \12621_b1 , \12619_b1 , w_32237 );
not ( w_32237 , w_32238 );
and ( \12621_b0 , \12619_b0 , w_32239 );
and ( w_32238 ,  , w_32239 );
buf ( w_32237 , \12620_b1 );
not ( w_32237 , w_32240 );
not (  , w_32241 );
and ( w_32240 , w_32241 , \12620_b0 );
or ( \12622_b1 , \12621_b1 , w_32242 );
xor ( \12622_b0 , \12621_b0 , w_32244 );
not ( w_32244 , w_32245 );
and ( w_32245 , w_32242 , w_32243 );
buf ( w_32242 , \7146_b1 );
not ( w_32242 , w_32246 );
not ( w_32243 , w_32247 );
and ( w_32246 , w_32247 , \7146_b0 );
or ( \12623_b1 , \6065_b1 , w_32249 );
not ( w_32249 , w_32250 );
and ( \12623_b0 , \6065_b0 , w_32251 );
and ( w_32250 ,  , w_32251 );
buf ( w_32249 , \7155_b1 );
not ( w_32249 , w_32252 );
not (  , w_32253 );
and ( w_32252 , w_32253 , \7155_b0 );
or ( \12624_b1 , \12623_b1 , w_32254 );
xor ( \12624_b0 , \12623_b0 , w_32256 );
not ( w_32256 , w_32257 );
and ( w_32257 , w_32254 , w_32255 );
buf ( w_32254 , \7163_b1 );
not ( w_32254 , w_32258 );
not ( w_32255 , w_32259 );
and ( w_32258 , w_32259 , \7163_b0 );
or ( \12625_b1 , \12622_b1 , \12624_b1 );
xor ( \12625_b0 , \12622_b0 , w_32260 );
not ( w_32260 , w_32261 );
and ( w_32261 , \12624_b1 , \12624_b0 );
or ( \12626_b1 , \5986_b1 , \7082_b1 );
not ( \7082_b1 , w_32262 );
and ( \12626_b0 , \5986_b0 , w_32263 );
and ( w_32262 , w_32263 , \7082_b0 );
or ( \12627_b1 , \5998_b1 , \7080_b1 );
not ( \7080_b1 , w_32264 );
and ( \12627_b0 , \5998_b0 , w_32265 );
and ( w_32264 , w_32265 , \7080_b0 );
or ( \12628_b1 , \12626_b1 , w_32267 );
not ( w_32267 , w_32268 );
and ( \12628_b0 , \12626_b0 , w_32269 );
and ( w_32268 ,  , w_32269 );
buf ( w_32267 , \12627_b1 );
not ( w_32267 , w_32270 );
not (  , w_32271 );
and ( w_32270 , w_32271 , \12627_b0 );
or ( \12629_b1 , \12628_b1 , w_32272 );
xor ( \12629_b0 , \12628_b0 , w_32274 );
not ( w_32274 , w_32275 );
and ( w_32275 , w_32272 , w_32273 );
buf ( w_32272 , \7088_b1 );
not ( w_32272 , w_32276 );
not ( w_32273 , w_32277 );
and ( w_32276 , w_32277 , \7088_b0 );
or ( \12630_b1 , \6006_b1 , \7099_b1 );
not ( \7099_b1 , w_32278 );
and ( \12630_b0 , \6006_b0 , w_32279 );
and ( w_32278 , w_32279 , \7099_b0 );
or ( \12631_b1 , \6018_b1 , \7097_b1 );
not ( \7097_b1 , w_32280 );
and ( \12631_b0 , \6018_b0 , w_32281 );
and ( w_32280 , w_32281 , \7097_b0 );
or ( \12632_b1 , \12630_b1 , w_32283 );
not ( w_32283 , w_32284 );
and ( \12632_b0 , \12630_b0 , w_32285 );
and ( w_32284 ,  , w_32285 );
buf ( w_32283 , \12631_b1 );
not ( w_32283 , w_32286 );
not (  , w_32287 );
and ( w_32286 , w_32287 , \12631_b0 );
or ( \12633_b1 , \12632_b1 , w_32288 );
xor ( \12633_b0 , \12632_b0 , w_32290 );
not ( w_32290 , w_32291 );
and ( w_32291 , w_32288 , w_32289 );
buf ( w_32288 , \7105_b1 );
not ( w_32288 , w_32292 );
not ( w_32289 , w_32293 );
and ( w_32292 , w_32293 , \7105_b0 );
or ( \12634_b1 , \12629_b1 , \12633_b1 );
xor ( \12634_b0 , \12629_b0 , w_32294 );
not ( w_32294 , w_32295 );
and ( w_32295 , \12633_b1 , \12633_b0 );
or ( \12635_b1 , \6029_b1 , \7117_b1 );
not ( \7117_b1 , w_32296 );
and ( \12635_b0 , \6029_b0 , w_32297 );
and ( w_32296 , w_32297 , \7117_b0 );
or ( \12636_b1 , \6041_b1 , \7115_b1 );
not ( \7115_b1 , w_32298 );
and ( \12636_b0 , \6041_b0 , w_32299 );
and ( w_32298 , w_32299 , \7115_b0 );
or ( \12637_b1 , \12635_b1 , w_32301 );
not ( w_32301 , w_32302 );
and ( \12637_b0 , \12635_b0 , w_32303 );
and ( w_32302 ,  , w_32303 );
buf ( w_32301 , \12636_b1 );
not ( w_32301 , w_32304 );
not (  , w_32305 );
and ( w_32304 , w_32305 , \12636_b0 );
or ( \12638_b1 , \12637_b1 , w_32306 );
xor ( \12638_b0 , \12637_b0 , w_32308 );
not ( w_32308 , w_32309 );
and ( w_32309 , w_32306 , w_32307 );
buf ( w_32306 , \7123_b1 );
not ( w_32306 , w_32310 );
not ( w_32307 , w_32311 );
and ( w_32310 , w_32311 , \7123_b0 );
or ( \12639_b1 , \12634_b1 , \12638_b1 );
xor ( \12639_b0 , \12634_b0 , w_32312 );
not ( w_32312 , w_32313 );
and ( w_32313 , \12638_b1 , \12638_b0 );
or ( \12640_b1 , \12625_b1 , \12639_b1 );
xor ( \12640_b0 , \12625_b0 , w_32314 );
not ( w_32314 , w_32315 );
and ( w_32315 , \12639_b1 , \12639_b0 );
or ( \12641_b1 , \12618_b1 , \12640_b1 );
xor ( \12641_b0 , \12618_b0 , w_32316 );
not ( w_32316 , w_32317 );
and ( w_32317 , \12640_b1 , \12640_b0 );
or ( \12642_b1 , \12561_b1 , \12565_b1 );
not ( \12565_b1 , w_32318 );
and ( \12642_b0 , \12561_b0 , w_32319 );
and ( w_32318 , w_32319 , \12565_b0 );
or ( \12643_b1 , \12565_b1 , \12570_b1 );
not ( \12570_b1 , w_32320 );
and ( \12643_b0 , \12565_b0 , w_32321 );
and ( w_32320 , w_32321 , \12570_b0 );
or ( \12644_b1 , \12561_b1 , \12570_b1 );
not ( \12570_b1 , w_32322 );
and ( \12644_b0 , \12561_b0 , w_32323 );
and ( w_32322 , w_32323 , \12570_b0 );
or ( \12646_b1 , \12546_b1 , \12550_b1 );
not ( \12550_b1 , w_32324 );
and ( \12646_b0 , \12546_b0 , w_32325 );
and ( w_32324 , w_32325 , \12550_b0 );
or ( \12647_b1 , \12550_b1 , \12555_b1 );
not ( \12555_b1 , w_32326 );
and ( \12647_b0 , \12550_b0 , w_32327 );
and ( w_32326 , w_32327 , \12555_b0 );
or ( \12648_b1 , \12546_b1 , \12555_b1 );
not ( \12555_b1 , w_32328 );
and ( \12648_b0 , \12546_b0 , w_32329 );
and ( w_32328 , w_32329 , \12555_b0 );
or ( \12650_b1 , \12645_b1 , \12649_b1 );
xor ( \12650_b0 , \12645_b0 , w_32330 );
not ( w_32330 , w_32331 );
and ( w_32331 , \12649_b1 , \12649_b0 );
or ( \12651_b1 , \12532_b1 , \12536_b1 );
not ( \12536_b1 , w_32332 );
and ( \12651_b0 , \12532_b0 , w_32333 );
and ( w_32332 , w_32333 , \12536_b0 );
or ( \12652_b1 , \12536_b1 , \12541_b1 );
not ( \12541_b1 , w_32334 );
and ( \12652_b0 , \12536_b0 , w_32335 );
and ( w_32334 , w_32335 , \12541_b0 );
or ( \12653_b1 , \12532_b1 , \12541_b1 );
not ( \12541_b1 , w_32336 );
and ( \12653_b0 , \12532_b0 , w_32337 );
and ( w_32336 , w_32337 , \12541_b0 );
or ( \12655_b1 , \12650_b1 , \12654_b1 );
xor ( \12655_b0 , \12650_b0 , w_32338 );
not ( w_32338 , w_32339 );
and ( w_32339 , \12654_b1 , \12654_b0 );
or ( \12656_b1 , \12641_b1 , \12655_b1 );
xor ( \12656_b0 , \12641_b0 , w_32340 );
not ( w_32340 , w_32341 );
and ( w_32341 , \12655_b1 , \12655_b0 );
or ( \12657_b1 , \12608_b1 , \12656_b1 );
xor ( \12657_b0 , \12608_b0 , w_32342 );
not ( w_32342 , w_32343 );
and ( w_32343 , \12656_b1 , \12656_b0 );
or ( \12658_b1 , \12583_b1 , \12587_b1 );
not ( \12587_b1 , w_32344 );
and ( \12658_b0 , \12583_b0 , w_32345 );
and ( w_32344 , w_32345 , \12587_b0 );
or ( \12659_b1 , \12587_b1 , \12592_b1 );
not ( \12592_b1 , w_32346 );
and ( \12659_b0 , \12587_b0 , w_32347 );
and ( w_32346 , w_32347 , \12592_b0 );
or ( \12660_b1 , \12583_b1 , \12592_b1 );
not ( \12592_b1 , w_32348 );
and ( \12660_b0 , \12583_b0 , w_32349 );
and ( w_32348 , w_32349 , \12592_b0 );
or ( \12662_b1 , \12542_b1 , \12556_b1 );
not ( \12556_b1 , w_32350 );
and ( \12662_b0 , \12542_b0 , w_32351 );
and ( w_32350 , w_32351 , \12556_b0 );
or ( \12663_b1 , \12556_b1 , \12571_b1 );
not ( \12571_b1 , w_32352 );
and ( \12663_b0 , \12556_b0 , w_32353 );
and ( w_32352 , w_32353 , \12571_b0 );
or ( \12664_b1 , \12542_b1 , \12571_b1 );
not ( \12571_b1 , w_32354 );
and ( \12664_b0 , \12542_b0 , w_32355 );
and ( w_32354 , w_32355 , \12571_b0 );
or ( \12666_b1 , \12661_b1 , \12665_b1 );
xor ( \12666_b0 , \12661_b0 , w_32356 );
not ( w_32356 , w_32357 );
and ( w_32357 , \12665_b1 , \12665_b0 );
or ( \12667_b1 , \5925_b1 , \7026_b1 );
not ( \7026_b1 , w_32358 );
and ( \12667_b0 , \5925_b0 , w_32359 );
and ( w_32358 , w_32359 , \7026_b0 );
or ( \12668_b1 , \5937_b1 , \7024_b1 );
not ( \7024_b1 , w_32360 );
and ( \12668_b0 , \5937_b0 , w_32361 );
and ( w_32360 , w_32361 , \7024_b0 );
or ( \12669_b1 , \12667_b1 , w_32363 );
not ( w_32363 , w_32364 );
and ( \12669_b0 , \12667_b0 , w_32365 );
and ( w_32364 ,  , w_32365 );
buf ( w_32363 , \12668_b1 );
not ( w_32363 , w_32366 );
not (  , w_32367 );
and ( w_32366 , w_32367 , \12668_b0 );
or ( \12670_b1 , \12669_b1 , w_32368 );
xor ( \12670_b0 , \12669_b0 , w_32370 );
not ( w_32370 , w_32371 );
and ( w_32371 , w_32368 , w_32369 );
buf ( w_32368 , \7032_b1 );
not ( w_32368 , w_32372 );
not ( w_32369 , w_32373 );
and ( w_32372 , w_32373 , \7032_b0 );
or ( \12671_b1 , \5945_b1 , \7043_b1 );
not ( \7043_b1 , w_32374 );
and ( \12671_b0 , \5945_b0 , w_32375 );
and ( w_32374 , w_32375 , \7043_b0 );
or ( \12672_b1 , \5957_b1 , \7041_b1 );
not ( \7041_b1 , w_32376 );
and ( \12672_b0 , \5957_b0 , w_32377 );
and ( w_32376 , w_32377 , \7041_b0 );
or ( \12673_b1 , \12671_b1 , w_32379 );
not ( w_32379 , w_32380 );
and ( \12673_b0 , \12671_b0 , w_32381 );
and ( w_32380 ,  , w_32381 );
buf ( w_32379 , \12672_b1 );
not ( w_32379 , w_32382 );
not (  , w_32383 );
and ( w_32382 , w_32383 , \12672_b0 );
or ( \12674_b1 , \12673_b1 , w_32384 );
xor ( \12674_b0 , \12673_b0 , w_32386 );
not ( w_32386 , w_32387 );
and ( w_32387 , w_32384 , w_32385 );
buf ( w_32384 , \7049_b1 );
not ( w_32384 , w_32388 );
not ( w_32385 , w_32389 );
and ( w_32388 , w_32389 , \7049_b0 );
or ( \12675_b1 , \12670_b1 , \12674_b1 );
xor ( \12675_b0 , \12670_b0 , w_32390 );
not ( w_32390 , w_32391 );
and ( w_32391 , \12674_b1 , \12674_b0 );
or ( \12676_b1 , \5967_b1 , \7061_b1 );
not ( \7061_b1 , w_32392 );
and ( \12676_b0 , \5967_b0 , w_32393 );
and ( w_32392 , w_32393 , \7061_b0 );
or ( \12677_b1 , \5979_b1 , \7059_b1 );
not ( \7059_b1 , w_32394 );
and ( \12677_b0 , \5979_b0 , w_32395 );
and ( w_32394 , w_32395 , \7059_b0 );
or ( \12678_b1 , \12676_b1 , w_32397 );
not ( w_32397 , w_32398 );
and ( \12678_b0 , \12676_b0 , w_32399 );
and ( w_32398 ,  , w_32399 );
buf ( w_32397 , \12677_b1 );
not ( w_32397 , w_32400 );
not (  , w_32401 );
and ( w_32400 , w_32401 , \12677_b0 );
or ( \12679_b1 , \12678_b1 , w_32402 );
xor ( \12679_b0 , \12678_b0 , w_32404 );
not ( w_32404 , w_32405 );
and ( w_32405 , w_32402 , w_32403 );
buf ( w_32402 , \7067_b1 );
not ( w_32402 , w_32406 );
not ( w_32403 , w_32407 );
and ( w_32406 , w_32407 , \7067_b0 );
or ( \12680_b1 , \12675_b1 , \12679_b1 );
xor ( \12680_b0 , \12675_b0 , w_32408 );
not ( w_32408 , w_32409 );
and ( w_32409 , \12679_b1 , \12679_b0 );
or ( \12681_b1 , \12666_b1 , \12680_b1 );
xor ( \12681_b0 , \12666_b0 , w_32410 );
not ( w_32410 , w_32411 );
and ( w_32411 , \12680_b1 , \12680_b0 );
or ( \12682_b1 , \12657_b1 , \12681_b1 );
xor ( \12682_b0 , \12657_b0 , w_32412 );
not ( w_32412 , w_32413 );
and ( w_32413 , \12681_b1 , \12681_b0 );
or ( \12683_b1 , \12604_b1 , \12682_b1 );
xor ( \12683_b0 , \12604_b0 , w_32414 );
not ( w_32414 , w_32415 );
and ( w_32415 , \12682_b1 , \12682_b0 );
or ( \12684_b1 , \12573_b1 , \12594_b1 );
not ( \12594_b1 , w_32416 );
and ( \12684_b0 , \12573_b0 , w_32417 );
and ( w_32416 , w_32417 , \12594_b0 );
or ( \12685_b1 , \12683_b1 , w_32419 );
not ( w_32419 , w_32420 );
and ( \12685_b0 , \12683_b0 , w_32421 );
and ( w_32420 ,  , w_32421 );
buf ( w_32419 , \12684_b1 );
not ( w_32419 , w_32422 );
not (  , w_32423 );
and ( w_32422 , w_32423 , \12684_b0 );
or ( \12686_b1 , \12600_b1 , w_32425 );
not ( w_32425 , w_32426 );
and ( \12686_b0 , \12600_b0 , w_32427 );
and ( w_32426 ,  , w_32427 );
buf ( w_32425 , \12685_b1 );
not ( w_32425 , w_32428 );
not (  , w_32429 );
and ( w_32428 , w_32429 , \12685_b0 );
or ( \12687_b1 , \12519_b1 , w_32431 );
not ( w_32431 , w_32432 );
and ( \12687_b0 , \12519_b0 , w_32433 );
and ( w_32432 ,  , w_32433 );
buf ( w_32431 , \12686_b1 );
not ( w_32431 , w_32434 );
not (  , w_32435 );
and ( w_32434 , w_32435 , \12686_b0 );
or ( \12688_b1 , \12608_b1 , \12656_b1 );
not ( \12656_b1 , w_32436 );
and ( \12688_b0 , \12608_b0 , w_32437 );
and ( w_32436 , w_32437 , \12656_b0 );
or ( \12689_b1 , \12656_b1 , \12681_b1 );
not ( \12681_b1 , w_32438 );
and ( \12689_b0 , \12656_b0 , w_32439 );
and ( w_32438 , w_32439 , \12681_b0 );
or ( \12690_b1 , \12608_b1 , \12681_b1 );
not ( \12681_b1 , w_32440 );
and ( \12690_b0 , \12608_b0 , w_32441 );
and ( w_32440 , w_32441 , \12681_b0 );
or ( \12692_b1 , \7163_b1 , \12612_b1 );
not ( \12612_b1 , w_32442 );
and ( \12692_b0 , \7163_b0 , w_32443 );
and ( w_32442 , w_32443 , \12612_b0 );
or ( \12693_b1 , \12612_b1 , \12617_b1 );
not ( \12617_b1 , w_32444 );
and ( \12693_b0 , \12612_b0 , w_32445 );
and ( w_32444 , w_32445 , \12617_b0 );
or ( \12694_b1 , \7163_b1 , \12617_b1 );
not ( \12617_b1 , w_32446 );
and ( \12694_b0 , \7163_b0 , w_32447 );
and ( w_32446 , w_32447 , \12617_b0 );
or ( \12696_b1 , \12670_b1 , \12674_b1 );
not ( \12674_b1 , w_32448 );
and ( \12696_b0 , \12670_b0 , w_32449 );
and ( w_32448 , w_32449 , \12674_b0 );
or ( \12697_b1 , \12674_b1 , \12679_b1 );
not ( \12679_b1 , w_32450 );
and ( \12697_b0 , \12674_b0 , w_32451 );
and ( w_32450 , w_32451 , \12679_b0 );
or ( \12698_b1 , \12670_b1 , \12679_b1 );
not ( \12679_b1 , w_32452 );
and ( \12698_b0 , \12670_b0 , w_32453 );
and ( w_32452 , w_32453 , \12679_b0 );
or ( \12700_b1 , \12695_b1 , \12699_b1 );
xor ( \12700_b0 , \12695_b0 , w_32454 );
not ( w_32454 , w_32455 );
and ( w_32455 , \12699_b1 , \12699_b0 );
or ( \12701_b1 , \12629_b1 , \12633_b1 );
not ( \12633_b1 , w_32456 );
and ( \12701_b0 , \12629_b0 , w_32457 );
and ( w_32456 , w_32457 , \12633_b0 );
or ( \12702_b1 , \12633_b1 , \12638_b1 );
not ( \12638_b1 , w_32458 );
and ( \12702_b0 , \12633_b0 , w_32459 );
and ( w_32458 , w_32459 , \12638_b0 );
or ( \12703_b1 , \12629_b1 , \12638_b1 );
not ( \12638_b1 , w_32460 );
and ( \12703_b0 , \12629_b0 , w_32461 );
and ( w_32460 , w_32461 , \12638_b0 );
or ( \12705_b1 , \12700_b1 , \12704_b1 );
xor ( \12705_b0 , \12700_b0 , w_32462 );
not ( w_32462 , w_32463 );
and ( w_32463 , \12704_b1 , \12704_b0 );
or ( \12706_b1 , \12645_b1 , \12649_b1 );
not ( \12649_b1 , w_32464 );
and ( \12706_b0 , \12645_b0 , w_32465 );
and ( w_32464 , w_32465 , \12649_b0 );
or ( \12707_b1 , \12649_b1 , \12654_b1 );
not ( \12654_b1 , w_32466 );
and ( \12707_b0 , \12649_b0 , w_32467 );
and ( w_32466 , w_32467 , \12654_b0 );
or ( \12708_b1 , \12645_b1 , \12654_b1 );
not ( \12654_b1 , w_32468 );
and ( \12708_b0 , \12645_b0 , w_32469 );
and ( w_32468 , w_32469 , \12654_b0 );
or ( \12710_b1 , \12622_b1 , \12624_b1 );
not ( \12624_b1 , w_32470 );
and ( \12710_b0 , \12622_b0 , w_32471 );
and ( w_32470 , w_32471 , \12624_b0 );
or ( \12711_b1 , \12624_b1 , \12639_b1 );
not ( \12639_b1 , w_32472 );
and ( \12711_b0 , \12624_b0 , w_32473 );
and ( w_32472 , w_32473 , \12639_b0 );
or ( \12712_b1 , \12622_b1 , \12639_b1 );
not ( \12639_b1 , w_32474 );
and ( \12712_b0 , \12622_b0 , w_32475 );
and ( w_32474 , w_32475 , \12639_b0 );
or ( \12714_b1 , \12709_b1 , \12713_b1 );
xor ( \12714_b0 , \12709_b0 , w_32476 );
not ( w_32476 , w_32477 );
and ( w_32477 , \12713_b1 , \12713_b0 );
or ( \12715_b1 , \5893_b1 , \6991_b1 );
not ( \6991_b1 , w_32478 );
and ( \12715_b0 , \5893_b0 , w_32479 );
and ( w_32478 , w_32479 , \6991_b0 );
or ( \12716_b1 , \5861_b1 , \6988_b1 );
not ( \6988_b1 , w_32480 );
and ( \12716_b0 , \5861_b0 , w_32481 );
and ( w_32480 , w_32481 , \6988_b0 );
or ( \12717_b1 , \12715_b1 , w_32483 );
not ( w_32483 , w_32484 );
and ( \12717_b0 , \12715_b0 , w_32485 );
and ( w_32484 ,  , w_32485 );
buf ( w_32483 , \12716_b1 );
not ( w_32483 , w_32486 );
not (  , w_32487 );
and ( w_32486 , w_32487 , \12716_b0 );
or ( \12718_b1 , \12717_b1 , w_32488 );
xor ( \12718_b0 , \12717_b0 , w_32490 );
not ( w_32490 , w_32491 );
and ( w_32491 , w_32488 , w_32489 );
buf ( w_32488 , \6985_b1 );
not ( w_32488 , w_32492 );
not ( w_32489 , w_32493 );
and ( w_32492 , w_32493 , \6985_b0 );
or ( \12719_b1 , \5918_b1 , \7006_b1 );
not ( \7006_b1 , w_32494 );
and ( \12719_b0 , \5918_b0 , w_32495 );
and ( w_32494 , w_32495 , \7006_b0 );
or ( \12720_b1 , \5881_b1 , \7004_b1 );
not ( \7004_b1 , w_32496 );
and ( \12720_b0 , \5881_b0 , w_32497 );
and ( w_32496 , w_32497 , \7004_b0 );
or ( \12721_b1 , \12719_b1 , w_32499 );
not ( w_32499 , w_32500 );
and ( \12721_b0 , \12719_b0 , w_32501 );
and ( w_32500 ,  , w_32501 );
buf ( w_32499 , \12720_b1 );
not ( w_32499 , w_32502 );
not (  , w_32503 );
and ( w_32502 , w_32503 , \12720_b0 );
or ( \12722_b1 , \12721_b1 , w_32504 );
xor ( \12722_b0 , \12721_b0 , w_32506 );
not ( w_32506 , w_32507 );
and ( w_32507 , w_32504 , w_32505 );
buf ( w_32504 , \7012_b1 );
not ( w_32504 , w_32508 );
not ( w_32505 , w_32509 );
and ( w_32508 , w_32509 , \7012_b0 );
or ( \12723_b1 , \12718_b1 , \12722_b1 );
xor ( \12723_b0 , \12718_b0 , w_32510 );
not ( w_32510 , w_32511 );
and ( w_32511 , \12722_b1 , \12722_b0 );
or ( \12724_b1 , \5937_b1 , \7026_b1 );
not ( \7026_b1 , w_32512 );
and ( \12724_b0 , \5937_b0 , w_32513 );
and ( w_32512 , w_32513 , \7026_b0 );
or ( \12725_b1 , \5906_b1 , \7024_b1 );
not ( \7024_b1 , w_32514 );
and ( \12725_b0 , \5906_b0 , w_32515 );
and ( w_32514 , w_32515 , \7024_b0 );
or ( \12726_b1 , \12724_b1 , w_32517 );
not ( w_32517 , w_32518 );
and ( \12726_b0 , \12724_b0 , w_32519 );
and ( w_32518 ,  , w_32519 );
buf ( w_32517 , \12725_b1 );
not ( w_32517 , w_32520 );
not (  , w_32521 );
and ( w_32520 , w_32521 , \12725_b0 );
or ( \12727_b1 , \12726_b1 , w_32522 );
xor ( \12727_b0 , \12726_b0 , w_32524 );
not ( w_32524 , w_32525 );
and ( w_32525 , w_32522 , w_32523 );
buf ( w_32522 , \7032_b1 );
not ( w_32522 , w_32526 );
not ( w_32523 , w_32527 );
and ( w_32526 , w_32527 , \7032_b0 );
or ( \12728_b1 , \12723_b1 , \12727_b1 );
xor ( \12728_b0 , \12723_b0 , w_32528 );
not ( w_32528 , w_32529 );
and ( w_32529 , \12727_b1 , \12727_b0 );
or ( \12729_b1 , \12714_b1 , \12728_b1 );
xor ( \12729_b0 , \12714_b0 , w_32530 );
not ( w_32530 , w_32531 );
and ( w_32531 , \12728_b1 , \12728_b0 );
or ( \12730_b1 , \12705_b1 , \12729_b1 );
xor ( \12730_b0 , \12705_b0 , w_32532 );
not ( w_32532 , w_32533 );
and ( w_32533 , \12729_b1 , \12729_b0 );
or ( \12731_b1 , \12691_b1 , \12730_b1 );
xor ( \12731_b0 , \12691_b0 , w_32534 );
not ( w_32534 , w_32535 );
and ( w_32535 , \12730_b1 , \12730_b0 );
or ( \12732_b1 , \12661_b1 , \12665_b1 );
not ( \12665_b1 , w_32536 );
and ( \12732_b0 , \12661_b0 , w_32537 );
and ( w_32536 , w_32537 , \12665_b0 );
or ( \12733_b1 , \12665_b1 , \12680_b1 );
not ( \12680_b1 , w_32538 );
and ( \12733_b0 , \12665_b0 , w_32539 );
and ( w_32538 , w_32539 , \12680_b0 );
or ( \12734_b1 , \12661_b1 , \12680_b1 );
not ( \12680_b1 , w_32540 );
and ( \12734_b0 , \12661_b0 , w_32541 );
and ( w_32540 , w_32541 , \12680_b0 );
or ( \12736_b1 , \12618_b1 , \12640_b1 );
not ( \12640_b1 , w_32542 );
and ( \12736_b0 , \12618_b0 , w_32543 );
and ( w_32542 , w_32543 , \12640_b0 );
or ( \12737_b1 , \12640_b1 , \12655_b1 );
not ( \12655_b1 , w_32544 );
and ( \12737_b0 , \12640_b0 , w_32545 );
and ( w_32544 , w_32545 , \12655_b0 );
or ( \12738_b1 , \12618_b1 , \12655_b1 );
not ( \12655_b1 , w_32546 );
and ( \12738_b0 , \12618_b0 , w_32547 );
and ( w_32546 , w_32547 , \12655_b0 );
or ( \12740_b1 , \12735_b1 , \12739_b1 );
xor ( \12740_b0 , \12735_b0 , w_32548 );
not ( w_32548 , w_32549 );
and ( w_32549 , \12739_b1 , \12739_b0 );
or ( \12741_b1 , \6065_b1 , \7157_b1 );
not ( \7157_b1 , w_32550 );
and ( \12741_b0 , \6065_b0 , w_32551 );
and ( w_32550 , w_32551 , \7157_b0 );
or ( \12742_b1 , \6048_b1 , \7155_b1 );
not ( \7155_b1 , w_32552 );
and ( \12742_b0 , \6048_b0 , w_32553 );
and ( w_32552 , w_32553 , \7155_b0 );
or ( \12743_b1 , \12741_b1 , w_32555 );
not ( w_32555 , w_32556 );
and ( \12743_b0 , \12741_b0 , w_32557 );
and ( w_32556 ,  , w_32557 );
buf ( w_32555 , \12742_b1 );
not ( w_32555 , w_32558 );
not (  , w_32559 );
and ( w_32558 , w_32559 , \12742_b0 );
or ( \12744_b1 , \12743_b1 , w_32560 );
xor ( \12744_b0 , \12743_b0 , w_32562 );
not ( w_32562 , w_32563 );
and ( w_32563 , w_32560 , w_32561 );
buf ( w_32560 , \7163_b1 );
not ( w_32560 , w_32564 );
not ( w_32561 , w_32565 );
and ( w_32564 , w_32565 , \7163_b0 );
or ( \12745_b1 , \6018_b1 , \7099_b1 );
not ( \7099_b1 , w_32566 );
and ( \12745_b0 , \6018_b0 , w_32567 );
and ( w_32566 , w_32567 , \7099_b0 );
or ( \12746_b1 , \5986_b1 , \7097_b1 );
not ( \7097_b1 , w_32568 );
and ( \12746_b0 , \5986_b0 , w_32569 );
and ( w_32568 , w_32569 , \7097_b0 );
or ( \12747_b1 , \12745_b1 , w_32571 );
not ( w_32571 , w_32572 );
and ( \12747_b0 , \12745_b0 , w_32573 );
and ( w_32572 ,  , w_32573 );
buf ( w_32571 , \12746_b1 );
not ( w_32571 , w_32574 );
not (  , w_32575 );
and ( w_32574 , w_32575 , \12746_b0 );
or ( \12748_b1 , \12747_b1 , w_32576 );
xor ( \12748_b0 , \12747_b0 , w_32578 );
not ( w_32578 , w_32579 );
and ( w_32579 , w_32576 , w_32577 );
buf ( w_32576 , \7105_b1 );
not ( w_32576 , w_32580 );
not ( w_32577 , w_32581 );
and ( w_32580 , w_32581 , \7105_b0 );
or ( \12749_b1 , \6041_b1 , \7117_b1 );
not ( \7117_b1 , w_32582 );
and ( \12749_b0 , \6041_b0 , w_32583 );
and ( w_32582 , w_32583 , \7117_b0 );
or ( \12750_b1 , \6006_b1 , \7115_b1 );
not ( \7115_b1 , w_32584 );
and ( \12750_b0 , \6006_b0 , w_32585 );
and ( w_32584 , w_32585 , \7115_b0 );
or ( \12751_b1 , \12749_b1 , w_32587 );
not ( w_32587 , w_32588 );
and ( \12751_b0 , \12749_b0 , w_32589 );
and ( w_32588 ,  , w_32589 );
buf ( w_32587 , \12750_b1 );
not ( w_32587 , w_32590 );
not (  , w_32591 );
and ( w_32590 , w_32591 , \12750_b0 );
or ( \12752_b1 , \12751_b1 , w_32592 );
xor ( \12752_b0 , \12751_b0 , w_32594 );
not ( w_32594 , w_32595 );
and ( w_32595 , w_32592 , w_32593 );
buf ( w_32592 , \7123_b1 );
not ( w_32592 , w_32596 );
not ( w_32593 , w_32597 );
and ( w_32596 , w_32597 , \7123_b0 );
or ( \12753_b1 , \12748_b1 , \12752_b1 );
xor ( \12753_b0 , \12748_b0 , w_32598 );
not ( w_32598 , w_32599 );
and ( w_32599 , \12752_b1 , \12752_b0 );
or ( \12754_b1 , \6057_b1 , \7140_b1 );
not ( \7140_b1 , w_32600 );
and ( \12754_b0 , \6057_b0 , w_32601 );
and ( w_32600 , w_32601 , \7140_b0 );
or ( \12755_b1 , \6029_b1 , \7138_b1 );
not ( \7138_b1 , w_32602 );
and ( \12755_b0 , \6029_b0 , w_32603 );
and ( w_32602 , w_32603 , \7138_b0 );
or ( \12756_b1 , \12754_b1 , w_32605 );
not ( w_32605 , w_32606 );
and ( \12756_b0 , \12754_b0 , w_32607 );
and ( w_32606 ,  , w_32607 );
buf ( w_32605 , \12755_b1 );
not ( w_32605 , w_32608 );
not (  , w_32609 );
and ( w_32608 , w_32609 , \12755_b0 );
or ( \12757_b1 , \12756_b1 , w_32610 );
xor ( \12757_b0 , \12756_b0 , w_32612 );
not ( w_32612 , w_32613 );
and ( w_32613 , w_32610 , w_32611 );
buf ( w_32610 , \7146_b1 );
not ( w_32610 , w_32614 );
not ( w_32611 , w_32615 );
and ( w_32614 , w_32615 , \7146_b0 );
or ( \12758_b1 , \12753_b1 , \12757_b1 );
xor ( \12758_b0 , \12753_b0 , w_32616 );
not ( w_32616 , w_32617 );
and ( w_32617 , \12757_b1 , \12757_b0 );
or ( \12759_b1 , \12744_b1 , \12758_b1 );
xor ( \12759_b0 , \12744_b0 , w_32618 );
not ( w_32618 , w_32619 );
and ( w_32619 , \12758_b1 , \12758_b0 );
or ( \12760_b1 , \5957_b1 , \7043_b1 );
not ( \7043_b1 , w_32620 );
and ( \12760_b0 , \5957_b0 , w_32621 );
and ( w_32620 , w_32621 , \7043_b0 );
or ( \12761_b1 , \5925_b1 , \7041_b1 );
not ( \7041_b1 , w_32622 );
and ( \12761_b0 , \5925_b0 , w_32623 );
and ( w_32622 , w_32623 , \7041_b0 );
or ( \12762_b1 , \12760_b1 , w_32625 );
not ( w_32625 , w_32626 );
and ( \12762_b0 , \12760_b0 , w_32627 );
and ( w_32626 ,  , w_32627 );
buf ( w_32625 , \12761_b1 );
not ( w_32625 , w_32628 );
not (  , w_32629 );
and ( w_32628 , w_32629 , \12761_b0 );
or ( \12763_b1 , \12762_b1 , w_32630 );
xor ( \12763_b0 , \12762_b0 , w_32632 );
not ( w_32632 , w_32633 );
and ( w_32633 , w_32630 , w_32631 );
buf ( w_32630 , \7049_b1 );
not ( w_32630 , w_32634 );
not ( w_32631 , w_32635 );
and ( w_32634 , w_32635 , \7049_b0 );
or ( \12764_b1 , \5979_b1 , \7061_b1 );
not ( \7061_b1 , w_32636 );
and ( \12764_b0 , \5979_b0 , w_32637 );
and ( w_32636 , w_32637 , \7061_b0 );
or ( \12765_b1 , \5945_b1 , \7059_b1 );
not ( \7059_b1 , w_32638 );
and ( \12765_b0 , \5945_b0 , w_32639 );
and ( w_32638 , w_32639 , \7059_b0 );
or ( \12766_b1 , \12764_b1 , w_32641 );
not ( w_32641 , w_32642 );
and ( \12766_b0 , \12764_b0 , w_32643 );
and ( w_32642 ,  , w_32643 );
buf ( w_32641 , \12765_b1 );
not ( w_32641 , w_32644 );
not (  , w_32645 );
and ( w_32644 , w_32645 , \12765_b0 );
or ( \12767_b1 , \12766_b1 , w_32646 );
xor ( \12767_b0 , \12766_b0 , w_32648 );
not ( w_32648 , w_32649 );
and ( w_32649 , w_32646 , w_32647 );
buf ( w_32646 , \7067_b1 );
not ( w_32646 , w_32650 );
not ( w_32647 , w_32651 );
and ( w_32650 , w_32651 , \7067_b0 );
or ( \12768_b1 , \12763_b1 , \12767_b1 );
xor ( \12768_b0 , \12763_b0 , w_32652 );
not ( w_32652 , w_32653 );
and ( w_32653 , \12767_b1 , \12767_b0 );
or ( \12769_b1 , \5998_b1 , \7082_b1 );
not ( \7082_b1 , w_32654 );
and ( \12769_b0 , \5998_b0 , w_32655 );
and ( w_32654 , w_32655 , \7082_b0 );
or ( \12770_b1 , \5967_b1 , \7080_b1 );
not ( \7080_b1 , w_32656 );
and ( \12770_b0 , \5967_b0 , w_32657 );
and ( w_32656 , w_32657 , \7080_b0 );
or ( \12771_b1 , \12769_b1 , w_32659 );
not ( w_32659 , w_32660 );
and ( \12771_b0 , \12769_b0 , w_32661 );
and ( w_32660 ,  , w_32661 );
buf ( w_32659 , \12770_b1 );
not ( w_32659 , w_32662 );
not (  , w_32663 );
and ( w_32662 , w_32663 , \12770_b0 );
or ( \12772_b1 , \12771_b1 , w_32664 );
xor ( \12772_b0 , \12771_b0 , w_32666 );
not ( w_32666 , w_32667 );
and ( w_32667 , w_32664 , w_32665 );
buf ( w_32664 , \7088_b1 );
not ( w_32664 , w_32668 );
not ( w_32665 , w_32669 );
and ( w_32668 , w_32669 , \7088_b0 );
or ( \12773_b1 , \12768_b1 , \12772_b1 );
xor ( \12773_b0 , \12768_b0 , w_32670 );
not ( w_32670 , w_32671 );
and ( w_32671 , \12772_b1 , \12772_b0 );
or ( \12774_b1 , \12759_b1 , \12773_b1 );
xor ( \12774_b0 , \12759_b0 , w_32672 );
not ( w_32672 , w_32673 );
and ( w_32673 , \12773_b1 , \12773_b0 );
or ( \12775_b1 , \12740_b1 , \12774_b1 );
xor ( \12775_b0 , \12740_b0 , w_32674 );
not ( w_32674 , w_32675 );
and ( w_32675 , \12774_b1 , \12774_b0 );
or ( \12776_b1 , \12731_b1 , \12775_b1 );
xor ( \12776_b0 , \12731_b0 , w_32676 );
not ( w_32676 , w_32677 );
and ( w_32677 , \12775_b1 , \12775_b0 );
or ( \12777_b1 , \12604_b1 , \12682_b1 );
not ( \12682_b1 , w_32678 );
and ( \12777_b0 , \12604_b0 , w_32679 );
and ( w_32678 , w_32679 , \12682_b0 );
or ( \12778_b1 , \12776_b1 , w_32681 );
not ( w_32681 , w_32682 );
and ( \12778_b0 , \12776_b0 , w_32683 );
and ( w_32682 ,  , w_32683 );
buf ( w_32681 , \12777_b1 );
not ( w_32681 , w_32684 );
not (  , w_32685 );
and ( w_32684 , w_32685 , \12777_b0 );
or ( \12779_b1 , \12735_b1 , \12739_b1 );
not ( \12739_b1 , w_32686 );
and ( \12779_b0 , \12735_b0 , w_32687 );
and ( w_32686 , w_32687 , \12739_b0 );
or ( \12780_b1 , \12739_b1 , \12774_b1 );
not ( \12774_b1 , w_32688 );
and ( \12780_b0 , \12739_b0 , w_32689 );
and ( w_32688 , w_32689 , \12774_b0 );
or ( \12781_b1 , \12735_b1 , \12774_b1 );
not ( \12774_b1 , w_32690 );
and ( \12781_b0 , \12735_b0 , w_32691 );
and ( w_32690 , w_32691 , \12774_b0 );
or ( \12783_b1 , \12705_b1 , \12729_b1 );
not ( \12729_b1 , w_32692 );
and ( \12783_b0 , \12705_b0 , w_32693 );
and ( w_32692 , w_32693 , \12729_b0 );
or ( \12784_b1 , \12782_b1 , \12783_b1 );
xor ( \12784_b0 , \12782_b0 , w_32694 );
not ( w_32694 , w_32695 );
and ( w_32695 , \12783_b1 , \12783_b0 );
or ( \12785_b1 , \12709_b1 , \12713_b1 );
not ( \12713_b1 , w_32696 );
and ( \12785_b0 , \12709_b0 , w_32697 );
and ( w_32696 , w_32697 , \12713_b0 );
or ( \12786_b1 , \12713_b1 , \12728_b1 );
not ( \12728_b1 , w_32698 );
and ( \12786_b0 , \12713_b0 , w_32699 );
and ( w_32698 , w_32699 , \12728_b0 );
or ( \12787_b1 , \12709_b1 , \12728_b1 );
not ( \12728_b1 , w_32700 );
and ( \12787_b0 , \12709_b0 , w_32701 );
and ( w_32700 , w_32701 , \12728_b0 );
or ( \12789_b1 , \6029_b1 , \7140_b1 );
not ( \7140_b1 , w_32702 );
and ( \12789_b0 , \6029_b0 , w_32703 );
and ( w_32702 , w_32703 , \7140_b0 );
or ( \12790_b1 , \6041_b1 , \7138_b1 );
not ( \7138_b1 , w_32704 );
and ( \12790_b0 , \6041_b0 , w_32705 );
and ( w_32704 , w_32705 , \7138_b0 );
or ( \12791_b1 , \12789_b1 , w_32707 );
not ( w_32707 , w_32708 );
and ( \12791_b0 , \12789_b0 , w_32709 );
and ( w_32708 ,  , w_32709 );
buf ( w_32707 , \12790_b1 );
not ( w_32707 , w_32710 );
not (  , w_32711 );
and ( w_32710 , w_32711 , \12790_b0 );
or ( \12792_b1 , \12791_b1 , w_32712 );
xor ( \12792_b0 , \12791_b0 , w_32714 );
not ( w_32714 , w_32715 );
and ( w_32715 , w_32712 , w_32713 );
buf ( w_32712 , \7146_b1 );
not ( w_32712 , w_32716 );
not ( w_32713 , w_32717 );
and ( w_32716 , w_32717 , \7146_b0 );
or ( \12793_b1 , \6048_b1 , \7157_b1 );
not ( \7157_b1 , w_32718 );
and ( \12793_b0 , \6048_b0 , w_32719 );
and ( w_32718 , w_32719 , \7157_b0 );
or ( \12794_b1 , \6057_b1 , \7155_b1 );
not ( \7155_b1 , w_32720 );
and ( \12794_b0 , \6057_b0 , w_32721 );
and ( w_32720 , w_32721 , \7155_b0 );
or ( \12795_b1 , \12793_b1 , w_32723 );
not ( w_32723 , w_32724 );
and ( \12795_b0 , \12793_b0 , w_32725 );
and ( w_32724 ,  , w_32725 );
buf ( w_32723 , \12794_b1 );
not ( w_32723 , w_32726 );
not (  , w_32727 );
and ( w_32726 , w_32727 , \12794_b0 );
or ( \12796_b1 , \12795_b1 , w_32728 );
xor ( \12796_b0 , \12795_b0 , w_32730 );
not ( w_32730 , w_32731 );
and ( w_32731 , w_32728 , w_32729 );
buf ( w_32728 , \7163_b1 );
not ( w_32728 , w_32732 );
not ( w_32729 , w_32733 );
and ( w_32732 , w_32733 , \7163_b0 );
or ( \12797_b1 , \12792_b1 , \12796_b1 );
xor ( \12797_b0 , \12792_b0 , w_32734 );
not ( w_32734 , w_32735 );
and ( w_32735 , \12796_b1 , \12796_b0 );
or ( \12798_b1 , \6065_b1 , w_32737 );
not ( w_32737 , w_32738 );
and ( \12798_b0 , \6065_b0 , w_32739 );
and ( w_32738 ,  , w_32739 );
buf ( w_32737 , \7173_b1 );
not ( w_32737 , w_32740 );
not (  , w_32741 );
and ( w_32740 , w_32741 , \7173_b0 );
or ( \12799_b1 , \12798_b1 , w_32742 );
xor ( \12799_b0 , \12798_b0 , w_32744 );
not ( w_32744 , w_32745 );
and ( w_32745 , w_32742 , w_32743 );
buf ( w_32742 , \7181_b1 );
not ( w_32742 , w_32746 );
not ( w_32743 , w_32747 );
and ( w_32746 , w_32747 , \7181_b0 );
or ( \12800_b1 , \12797_b1 , \12799_b1 );
xor ( \12800_b0 , \12797_b0 , w_32748 );
not ( w_32748 , w_32749 );
and ( w_32749 , \12799_b1 , \12799_b0 );
or ( \12801_b1 , \5967_b1 , \7082_b1 );
not ( \7082_b1 , w_32750 );
and ( \12801_b0 , \5967_b0 , w_32751 );
and ( w_32750 , w_32751 , \7082_b0 );
or ( \12802_b1 , \5979_b1 , \7080_b1 );
not ( \7080_b1 , w_32752 );
and ( \12802_b0 , \5979_b0 , w_32753 );
and ( w_32752 , w_32753 , \7080_b0 );
or ( \12803_b1 , \12801_b1 , w_32755 );
not ( w_32755 , w_32756 );
and ( \12803_b0 , \12801_b0 , w_32757 );
and ( w_32756 ,  , w_32757 );
buf ( w_32755 , \12802_b1 );
not ( w_32755 , w_32758 );
not (  , w_32759 );
and ( w_32758 , w_32759 , \12802_b0 );
or ( \12804_b1 , \12803_b1 , w_32760 );
xor ( \12804_b0 , \12803_b0 , w_32762 );
not ( w_32762 , w_32763 );
and ( w_32763 , w_32760 , w_32761 );
buf ( w_32760 , \7088_b1 );
not ( w_32760 , w_32764 );
not ( w_32761 , w_32765 );
and ( w_32764 , w_32765 , \7088_b0 );
or ( \12805_b1 , \5986_b1 , \7099_b1 );
not ( \7099_b1 , w_32766 );
and ( \12805_b0 , \5986_b0 , w_32767 );
and ( w_32766 , w_32767 , \7099_b0 );
or ( \12806_b1 , \5998_b1 , \7097_b1 );
not ( \7097_b1 , w_32768 );
and ( \12806_b0 , \5998_b0 , w_32769 );
and ( w_32768 , w_32769 , \7097_b0 );
or ( \12807_b1 , \12805_b1 , w_32771 );
not ( w_32771 , w_32772 );
and ( \12807_b0 , \12805_b0 , w_32773 );
and ( w_32772 ,  , w_32773 );
buf ( w_32771 , \12806_b1 );
not ( w_32771 , w_32774 );
not (  , w_32775 );
and ( w_32774 , w_32775 , \12806_b0 );
or ( \12808_b1 , \12807_b1 , w_32776 );
xor ( \12808_b0 , \12807_b0 , w_32778 );
not ( w_32778 , w_32779 );
and ( w_32779 , w_32776 , w_32777 );
buf ( w_32776 , \7105_b1 );
not ( w_32776 , w_32780 );
not ( w_32777 , w_32781 );
and ( w_32780 , w_32781 , \7105_b0 );
or ( \12809_b1 , \12804_b1 , \12808_b1 );
xor ( \12809_b0 , \12804_b0 , w_32782 );
not ( w_32782 , w_32783 );
and ( w_32783 , \12808_b1 , \12808_b0 );
or ( \12810_b1 , \6006_b1 , \7117_b1 );
not ( \7117_b1 , w_32784 );
and ( \12810_b0 , \6006_b0 , w_32785 );
and ( w_32784 , w_32785 , \7117_b0 );
or ( \12811_b1 , \6018_b1 , \7115_b1 );
not ( \7115_b1 , w_32786 );
and ( \12811_b0 , \6018_b0 , w_32787 );
and ( w_32786 , w_32787 , \7115_b0 );
or ( \12812_b1 , \12810_b1 , w_32789 );
not ( w_32789 , w_32790 );
and ( \12812_b0 , \12810_b0 , w_32791 );
and ( w_32790 ,  , w_32791 );
buf ( w_32789 , \12811_b1 );
not ( w_32789 , w_32792 );
not (  , w_32793 );
and ( w_32792 , w_32793 , \12811_b0 );
or ( \12813_b1 , \12812_b1 , w_32794 );
xor ( \12813_b0 , \12812_b0 , w_32796 );
not ( w_32796 , w_32797 );
and ( w_32797 , w_32794 , w_32795 );
buf ( w_32794 , \7123_b1 );
not ( w_32794 , w_32798 );
not ( w_32795 , w_32799 );
and ( w_32798 , w_32799 , \7123_b0 );
or ( \12814_b1 , \12809_b1 , \12813_b1 );
xor ( \12814_b0 , \12809_b0 , w_32800 );
not ( w_32800 , w_32801 );
and ( w_32801 , \12813_b1 , \12813_b0 );
or ( \12815_b1 , \12800_b1 , \12814_b1 );
xor ( \12815_b0 , \12800_b0 , w_32802 );
not ( w_32802 , w_32803 );
and ( w_32803 , \12814_b1 , \12814_b0 );
or ( \12816_b1 , \5906_b1 , \7026_b1 );
not ( \7026_b1 , w_32804 );
and ( \12816_b0 , \5906_b0 , w_32805 );
and ( w_32804 , w_32805 , \7026_b0 );
or ( \12817_b1 , \5918_b1 , \7024_b1 );
not ( \7024_b1 , w_32806 );
and ( \12817_b0 , \5918_b0 , w_32807 );
and ( w_32806 , w_32807 , \7024_b0 );
or ( \12818_b1 , \12816_b1 , w_32809 );
not ( w_32809 , w_32810 );
and ( \12818_b0 , \12816_b0 , w_32811 );
and ( w_32810 ,  , w_32811 );
buf ( w_32809 , \12817_b1 );
not ( w_32809 , w_32812 );
not (  , w_32813 );
and ( w_32812 , w_32813 , \12817_b0 );
or ( \12819_b1 , \12818_b1 , w_32814 );
xor ( \12819_b0 , \12818_b0 , w_32816 );
not ( w_32816 , w_32817 );
and ( w_32817 , w_32814 , w_32815 );
buf ( w_32814 , \7032_b1 );
not ( w_32814 , w_32818 );
not ( w_32815 , w_32819 );
and ( w_32818 , w_32819 , \7032_b0 );
or ( \12820_b1 , \5925_b1 , \7043_b1 );
not ( \7043_b1 , w_32820 );
and ( \12820_b0 , \5925_b0 , w_32821 );
and ( w_32820 , w_32821 , \7043_b0 );
or ( \12821_b1 , \5937_b1 , \7041_b1 );
not ( \7041_b1 , w_32822 );
and ( \12821_b0 , \5937_b0 , w_32823 );
and ( w_32822 , w_32823 , \7041_b0 );
or ( \12822_b1 , \12820_b1 , w_32825 );
not ( w_32825 , w_32826 );
and ( \12822_b0 , \12820_b0 , w_32827 );
and ( w_32826 ,  , w_32827 );
buf ( w_32825 , \12821_b1 );
not ( w_32825 , w_32828 );
not (  , w_32829 );
and ( w_32828 , w_32829 , \12821_b0 );
or ( \12823_b1 , \12822_b1 , w_32830 );
xor ( \12823_b0 , \12822_b0 , w_32832 );
not ( w_32832 , w_32833 );
and ( w_32833 , w_32830 , w_32831 );
buf ( w_32830 , \7049_b1 );
not ( w_32830 , w_32834 );
not ( w_32831 , w_32835 );
and ( w_32834 , w_32835 , \7049_b0 );
or ( \12824_b1 , \12819_b1 , \12823_b1 );
xor ( \12824_b0 , \12819_b0 , w_32836 );
not ( w_32836 , w_32837 );
and ( w_32837 , \12823_b1 , \12823_b0 );
or ( \12825_b1 , \5945_b1 , \7061_b1 );
not ( \7061_b1 , w_32838 );
and ( \12825_b0 , \5945_b0 , w_32839 );
and ( w_32838 , w_32839 , \7061_b0 );
or ( \12826_b1 , \5957_b1 , \7059_b1 );
not ( \7059_b1 , w_32840 );
and ( \12826_b0 , \5957_b0 , w_32841 );
and ( w_32840 , w_32841 , \7059_b0 );
or ( \12827_b1 , \12825_b1 , w_32843 );
not ( w_32843 , w_32844 );
and ( \12827_b0 , \12825_b0 , w_32845 );
and ( w_32844 ,  , w_32845 );
buf ( w_32843 , \12826_b1 );
not ( w_32843 , w_32846 );
not (  , w_32847 );
and ( w_32846 , w_32847 , \12826_b0 );
or ( \12828_b1 , \12827_b1 , w_32848 );
xor ( \12828_b0 , \12827_b0 , w_32850 );
not ( w_32850 , w_32851 );
and ( w_32851 , w_32848 , w_32849 );
buf ( w_32848 , \7067_b1 );
not ( w_32848 , w_32852 );
not ( w_32849 , w_32853 );
and ( w_32852 , w_32853 , \7067_b0 );
or ( \12829_b1 , \12824_b1 , \12828_b1 );
xor ( \12829_b0 , \12824_b0 , w_32854 );
not ( w_32854 , w_32855 );
and ( w_32855 , \12828_b1 , \12828_b0 );
or ( \12830_b1 , \12815_b1 , \12829_b1 );
xor ( \12830_b0 , \12815_b0 , w_32856 );
not ( w_32856 , w_32857 );
and ( w_32857 , \12829_b1 , \12829_b0 );
or ( \12831_b1 , \12718_b1 , \12722_b1 );
not ( \12722_b1 , w_32858 );
and ( \12831_b0 , \12718_b0 , w_32859 );
and ( w_32858 , w_32859 , \12722_b0 );
or ( \12832_b1 , \12722_b1 , \12727_b1 );
not ( \12727_b1 , w_32860 );
and ( \12832_b0 , \12722_b0 , w_32861 );
and ( w_32860 , w_32861 , \12727_b0 );
or ( \12833_b1 , \12718_b1 , \12727_b1 );
not ( \12727_b1 , w_32862 );
and ( \12833_b0 , \12718_b0 , w_32863 );
and ( w_32862 , w_32863 , \12727_b0 );
or ( \12835_b1 , \12763_b1 , \12767_b1 );
not ( \12767_b1 , w_32864 );
and ( \12835_b0 , \12763_b0 , w_32865 );
and ( w_32864 , w_32865 , \12767_b0 );
or ( \12836_b1 , \12767_b1 , \12772_b1 );
not ( \12772_b1 , w_32866 );
and ( \12836_b0 , \12767_b0 , w_32867 );
and ( w_32866 , w_32867 , \12772_b0 );
or ( \12837_b1 , \12763_b1 , \12772_b1 );
not ( \12772_b1 , w_32868 );
and ( \12837_b0 , \12763_b0 , w_32869 );
and ( w_32868 , w_32869 , \12772_b0 );
or ( \12839_b1 , \12834_b1 , \12838_b1 );
xor ( \12839_b0 , \12834_b0 , w_32870 );
not ( w_32870 , w_32871 );
and ( w_32871 , \12838_b1 , \12838_b0 );
or ( \12840_b1 , \12748_b1 , \12752_b1 );
not ( \12752_b1 , w_32872 );
and ( \12840_b0 , \12748_b0 , w_32873 );
and ( w_32872 , w_32873 , \12752_b0 );
or ( \12841_b1 , \12752_b1 , \12757_b1 );
not ( \12757_b1 , w_32874 );
and ( \12841_b0 , \12752_b0 , w_32875 );
and ( w_32874 , w_32875 , \12757_b0 );
or ( \12842_b1 , \12748_b1 , \12757_b1 );
not ( \12757_b1 , w_32876 );
and ( \12842_b0 , \12748_b0 , w_32877 );
and ( w_32876 , w_32877 , \12757_b0 );
or ( \12844_b1 , \12839_b1 , \12843_b1 );
xor ( \12844_b0 , \12839_b0 , w_32878 );
not ( w_32878 , w_32879 );
and ( w_32879 , \12843_b1 , \12843_b0 );
or ( \12845_b1 , \12830_b1 , \12844_b1 );
xor ( \12845_b0 , \12830_b0 , w_32880 );
not ( w_32880 , w_32881 );
and ( w_32881 , \12844_b1 , \12844_b0 );
or ( \12846_b1 , \12788_b1 , \12845_b1 );
xor ( \12846_b0 , \12788_b0 , w_32882 );
not ( w_32882 , w_32883 );
and ( w_32883 , \12845_b1 , \12845_b0 );
or ( \12847_b1 , \12695_b1 , \12699_b1 );
not ( \12699_b1 , w_32884 );
and ( \12847_b0 , \12695_b0 , w_32885 );
and ( w_32884 , w_32885 , \12699_b0 );
or ( \12848_b1 , \12699_b1 , \12704_b1 );
not ( \12704_b1 , w_32886 );
and ( \12848_b0 , \12699_b0 , w_32887 );
and ( w_32886 , w_32887 , \12704_b0 );
or ( \12849_b1 , \12695_b1 , \12704_b1 );
not ( \12704_b1 , w_32888 );
and ( \12849_b0 , \12695_b0 , w_32889 );
and ( w_32888 , w_32889 , \12704_b0 );
or ( \12851_b1 , \12744_b1 , \12758_b1 );
not ( \12758_b1 , w_32890 );
and ( \12851_b0 , \12744_b0 , w_32891 );
and ( w_32890 , w_32891 , \12758_b0 );
or ( \12852_b1 , \12758_b1 , \12773_b1 );
not ( \12773_b1 , w_32892 );
and ( \12852_b0 , \12758_b0 , w_32893 );
and ( w_32892 , w_32893 , \12773_b0 );
or ( \12853_b1 , \12744_b1 , \12773_b1 );
not ( \12773_b1 , w_32894 );
and ( \12853_b0 , \12744_b0 , w_32895 );
and ( w_32894 , w_32895 , \12773_b0 );
or ( \12855_b1 , \12850_b1 , \12854_b1 );
xor ( \12855_b0 , \12850_b0 , w_32896 );
not ( w_32896 , w_32897 );
and ( w_32897 , \12854_b1 , \12854_b0 );
or ( \12856_b1 , \5861_b1 , \6991_b1 );
not ( \6991_b1 , w_32898 );
and ( \12856_b0 , \5861_b0 , w_32899 );
and ( w_32898 , w_32899 , \6991_b0 );
or ( \12857_b1 , \5873_b1 , \6988_b1 );
not ( \6988_b1 , w_32900 );
and ( \12857_b0 , \5873_b0 , w_32901 );
and ( w_32900 , w_32901 , \6988_b0 );
or ( \12858_b1 , \12856_b1 , w_32903 );
not ( w_32903 , w_32904 );
and ( \12858_b0 , \12856_b0 , w_32905 );
and ( w_32904 ,  , w_32905 );
buf ( w_32903 , \12857_b1 );
not ( w_32903 , w_32906 );
not (  , w_32907 );
and ( w_32906 , w_32907 , \12857_b0 );
or ( \12859_b1 , \12858_b1 , w_32908 );
xor ( \12859_b0 , \12858_b0 , w_32910 );
not ( w_32910 , w_32911 );
and ( w_32911 , w_32908 , w_32909 );
buf ( w_32908 , \6985_b1 );
not ( w_32908 , w_32912 );
not ( w_32909 , w_32913 );
and ( w_32912 , w_32913 , \6985_b0 );
or ( \12860_b1 , \7181_b1 , \12859_b1 );
xor ( \12860_b0 , \7181_b0 , w_32914 );
not ( w_32914 , w_32915 );
and ( w_32915 , \12859_b1 , \12859_b0 );
or ( \12861_b1 , \5881_b1 , \7006_b1 );
not ( \7006_b1 , w_32916 );
and ( \12861_b0 , \5881_b0 , w_32917 );
and ( w_32916 , w_32917 , \7006_b0 );
or ( \12862_b1 , \5893_b1 , \7004_b1 );
not ( \7004_b1 , w_32918 );
and ( \12862_b0 , \5893_b0 , w_32919 );
and ( w_32918 , w_32919 , \7004_b0 );
or ( \12863_b1 , \12861_b1 , w_32921 );
not ( w_32921 , w_32922 );
and ( \12863_b0 , \12861_b0 , w_32923 );
and ( w_32922 ,  , w_32923 );
buf ( w_32921 , \12862_b1 );
not ( w_32921 , w_32924 );
not (  , w_32925 );
and ( w_32924 , w_32925 , \12862_b0 );
or ( \12864_b1 , \12863_b1 , w_32926 );
xor ( \12864_b0 , \12863_b0 , w_32928 );
not ( w_32928 , w_32929 );
and ( w_32929 , w_32926 , w_32927 );
buf ( w_32926 , \7012_b1 );
not ( w_32926 , w_32930 );
not ( w_32927 , w_32931 );
and ( w_32930 , w_32931 , \7012_b0 );
or ( \12865_b1 , \12860_b1 , \12864_b1 );
xor ( \12865_b0 , \12860_b0 , w_32932 );
not ( w_32932 , w_32933 );
and ( w_32933 , \12864_b1 , \12864_b0 );
or ( \12866_b1 , \12855_b1 , \12865_b1 );
xor ( \12866_b0 , \12855_b0 , w_32934 );
not ( w_32934 , w_32935 );
and ( w_32935 , \12865_b1 , \12865_b0 );
or ( \12867_b1 , \12846_b1 , \12866_b1 );
xor ( \12867_b0 , \12846_b0 , w_32936 );
not ( w_32936 , w_32937 );
and ( w_32937 , \12866_b1 , \12866_b0 );
or ( \12868_b1 , \12784_b1 , \12867_b1 );
xor ( \12868_b0 , \12784_b0 , w_32938 );
not ( w_32938 , w_32939 );
and ( w_32939 , \12867_b1 , \12867_b0 );
or ( \12869_b1 , \12691_b1 , \12730_b1 );
not ( \12730_b1 , w_32940 );
and ( \12869_b0 , \12691_b0 , w_32941 );
and ( w_32940 , w_32941 , \12730_b0 );
or ( \12870_b1 , \12730_b1 , \12775_b1 );
not ( \12775_b1 , w_32942 );
and ( \12870_b0 , \12730_b0 , w_32943 );
and ( w_32942 , w_32943 , \12775_b0 );
or ( \12871_b1 , \12691_b1 , \12775_b1 );
not ( \12775_b1 , w_32944 );
and ( \12871_b0 , \12691_b0 , w_32945 );
and ( w_32944 , w_32945 , \12775_b0 );
or ( \12873_b1 , \12868_b1 , w_32947 );
not ( w_32947 , w_32948 );
and ( \12873_b0 , \12868_b0 , w_32949 );
and ( w_32948 ,  , w_32949 );
buf ( w_32947 , \12872_b1 );
not ( w_32947 , w_32950 );
not (  , w_32951 );
and ( w_32950 , w_32951 , \12872_b0 );
or ( \12874_b1 , \12778_b1 , w_32953 );
not ( w_32953 , w_32954 );
and ( \12874_b0 , \12778_b0 , w_32955 );
and ( w_32954 ,  , w_32955 );
buf ( w_32953 , \12873_b1 );
not ( w_32953 , w_32956 );
not (  , w_32957 );
and ( w_32956 , w_32957 , \12873_b0 );
or ( \12875_b1 , \12788_b1 , \12845_b1 );
not ( \12845_b1 , w_32958 );
and ( \12875_b0 , \12788_b0 , w_32959 );
and ( w_32958 , w_32959 , \12845_b0 );
or ( \12876_b1 , \12845_b1 , \12866_b1 );
not ( \12866_b1 , w_32960 );
and ( \12876_b0 , \12845_b0 , w_32961 );
and ( w_32960 , w_32961 , \12866_b0 );
or ( \12877_b1 , \12788_b1 , \12866_b1 );
not ( \12866_b1 , w_32962 );
and ( \12877_b0 , \12788_b0 , w_32963 );
and ( w_32962 , w_32963 , \12866_b0 );
or ( \12879_b1 , \7181_b1 , \12859_b1 );
not ( \12859_b1 , w_32964 );
and ( \12879_b0 , \7181_b0 , w_32965 );
and ( w_32964 , w_32965 , \12859_b0 );
or ( \12880_b1 , \12859_b1 , \12864_b1 );
not ( \12864_b1 , w_32966 );
and ( \12880_b0 , \12859_b0 , w_32967 );
and ( w_32966 , w_32967 , \12864_b0 );
or ( \12881_b1 , \7181_b1 , \12864_b1 );
not ( \12864_b1 , w_32968 );
and ( \12881_b0 , \7181_b0 , w_32969 );
and ( w_32968 , w_32969 , \12864_b0 );
or ( \12883_b1 , \12819_b1 , \12823_b1 );
not ( \12823_b1 , w_32970 );
and ( \12883_b0 , \12819_b0 , w_32971 );
and ( w_32970 , w_32971 , \12823_b0 );
or ( \12884_b1 , \12823_b1 , \12828_b1 );
not ( \12828_b1 , w_32972 );
and ( \12884_b0 , \12823_b0 , w_32973 );
and ( w_32972 , w_32973 , \12828_b0 );
or ( \12885_b1 , \12819_b1 , \12828_b1 );
not ( \12828_b1 , w_32974 );
and ( \12885_b0 , \12819_b0 , w_32975 );
and ( w_32974 , w_32975 , \12828_b0 );
or ( \12887_b1 , \12882_b1 , \12886_b1 );
xor ( \12887_b0 , \12882_b0 , w_32976 );
not ( w_32976 , w_32977 );
and ( w_32977 , \12886_b1 , \12886_b0 );
or ( \12888_b1 , \12804_b1 , \12808_b1 );
not ( \12808_b1 , w_32978 );
and ( \12888_b0 , \12804_b0 , w_32979 );
and ( w_32978 , w_32979 , \12808_b0 );
or ( \12889_b1 , \12808_b1 , \12813_b1 );
not ( \12813_b1 , w_32980 );
and ( \12889_b0 , \12808_b0 , w_32981 );
and ( w_32980 , w_32981 , \12813_b0 );
or ( \12890_b1 , \12804_b1 , \12813_b1 );
not ( \12813_b1 , w_32982 );
and ( \12890_b0 , \12804_b0 , w_32983 );
and ( w_32982 , w_32983 , \12813_b0 );
or ( \12892_b1 , \12887_b1 , \12891_b1 );
xor ( \12892_b0 , \12887_b0 , w_32984 );
not ( w_32984 , w_32985 );
and ( w_32985 , \12891_b1 , \12891_b0 );
or ( \12893_b1 , \12834_b1 , \12838_b1 );
not ( \12838_b1 , w_32986 );
and ( \12893_b0 , \12834_b0 , w_32987 );
and ( w_32986 , w_32987 , \12838_b0 );
or ( \12894_b1 , \12838_b1 , \12843_b1 );
not ( \12843_b1 , w_32988 );
and ( \12894_b0 , \12838_b0 , w_32989 );
and ( w_32988 , w_32989 , \12843_b0 );
or ( \12895_b1 , \12834_b1 , \12843_b1 );
not ( \12843_b1 , w_32990 );
and ( \12895_b0 , \12834_b0 , w_32991 );
and ( w_32990 , w_32991 , \12843_b0 );
or ( \12897_b1 , \12800_b1 , \12814_b1 );
not ( \12814_b1 , w_32992 );
and ( \12897_b0 , \12800_b0 , w_32993 );
and ( w_32992 , w_32993 , \12814_b0 );
or ( \12898_b1 , \12814_b1 , \12829_b1 );
not ( \12829_b1 , w_32994 );
and ( \12898_b0 , \12814_b0 , w_32995 );
and ( w_32994 , w_32995 , \12829_b0 );
or ( \12899_b1 , \12800_b1 , \12829_b1 );
not ( \12829_b1 , w_32996 );
and ( \12899_b0 , \12800_b0 , w_32997 );
and ( w_32996 , w_32997 , \12829_b0 );
or ( \12901_b1 , \12896_b1 , \12900_b1 );
xor ( \12901_b0 , \12896_b0 , w_32998 );
not ( w_32998 , w_32999 );
and ( w_32999 , \12900_b1 , \12900_b0 );
or ( \12902_b1 , \5998_b1 , \7099_b1 );
not ( \7099_b1 , w_33000 );
and ( \12902_b0 , \5998_b0 , w_33001 );
and ( w_33000 , w_33001 , \7099_b0 );
or ( \12903_b1 , \5967_b1 , \7097_b1 );
not ( \7097_b1 , w_33002 );
and ( \12903_b0 , \5967_b0 , w_33003 );
and ( w_33002 , w_33003 , \7097_b0 );
or ( \12904_b1 , \12902_b1 , w_33005 );
not ( w_33005 , w_33006 );
and ( \12904_b0 , \12902_b0 , w_33007 );
and ( w_33006 ,  , w_33007 );
buf ( w_33005 , \12903_b1 );
not ( w_33005 , w_33008 );
not (  , w_33009 );
and ( w_33008 , w_33009 , \12903_b0 );
or ( \12905_b1 , \12904_b1 , w_33010 );
xor ( \12905_b0 , \12904_b0 , w_33012 );
not ( w_33012 , w_33013 );
and ( w_33013 , w_33010 , w_33011 );
buf ( w_33010 , \7105_b1 );
not ( w_33010 , w_33014 );
not ( w_33011 , w_33015 );
and ( w_33014 , w_33015 , \7105_b0 );
or ( \12906_b1 , \6018_b1 , \7117_b1 );
not ( \7117_b1 , w_33016 );
and ( \12906_b0 , \6018_b0 , w_33017 );
and ( w_33016 , w_33017 , \7117_b0 );
or ( \12907_b1 , \5986_b1 , \7115_b1 );
not ( \7115_b1 , w_33018 );
and ( \12907_b0 , \5986_b0 , w_33019 );
and ( w_33018 , w_33019 , \7115_b0 );
or ( \12908_b1 , \12906_b1 , w_33021 );
not ( w_33021 , w_33022 );
and ( \12908_b0 , \12906_b0 , w_33023 );
and ( w_33022 ,  , w_33023 );
buf ( w_33021 , \12907_b1 );
not ( w_33021 , w_33024 );
not (  , w_33025 );
and ( w_33024 , w_33025 , \12907_b0 );
or ( \12909_b1 , \12908_b1 , w_33026 );
xor ( \12909_b0 , \12908_b0 , w_33028 );
not ( w_33028 , w_33029 );
and ( w_33029 , w_33026 , w_33027 );
buf ( w_33026 , \7123_b1 );
not ( w_33026 , w_33030 );
not ( w_33027 , w_33031 );
and ( w_33030 , w_33031 , \7123_b0 );
or ( \12910_b1 , \12905_b1 , \12909_b1 );
xor ( \12910_b0 , \12905_b0 , w_33032 );
not ( w_33032 , w_33033 );
and ( w_33033 , \12909_b1 , \12909_b0 );
or ( \12911_b1 , \6041_b1 , \7140_b1 );
not ( \7140_b1 , w_33034 );
and ( \12911_b0 , \6041_b0 , w_33035 );
and ( w_33034 , w_33035 , \7140_b0 );
or ( \12912_b1 , \6006_b1 , \7138_b1 );
not ( \7138_b1 , w_33036 );
and ( \12912_b0 , \6006_b0 , w_33037 );
and ( w_33036 , w_33037 , \7138_b0 );
or ( \12913_b1 , \12911_b1 , w_33039 );
not ( w_33039 , w_33040 );
and ( \12913_b0 , \12911_b0 , w_33041 );
and ( w_33040 ,  , w_33041 );
buf ( w_33039 , \12912_b1 );
not ( w_33039 , w_33042 );
not (  , w_33043 );
and ( w_33042 , w_33043 , \12912_b0 );
or ( \12914_b1 , \12913_b1 , w_33044 );
xor ( \12914_b0 , \12913_b0 , w_33046 );
not ( w_33046 , w_33047 );
and ( w_33047 , w_33044 , w_33045 );
buf ( w_33044 , \7146_b1 );
not ( w_33044 , w_33048 );
not ( w_33045 , w_33049 );
and ( w_33048 , w_33049 , \7146_b0 );
or ( \12915_b1 , \12910_b1 , \12914_b1 );
xor ( \12915_b0 , \12910_b0 , w_33050 );
not ( w_33050 , w_33051 );
and ( w_33051 , \12914_b1 , \12914_b0 );
or ( \12916_b1 , \5937_b1 , \7043_b1 );
not ( \7043_b1 , w_33052 );
and ( \12916_b0 , \5937_b0 , w_33053 );
and ( w_33052 , w_33053 , \7043_b0 );
or ( \12917_b1 , \5906_b1 , \7041_b1 );
not ( \7041_b1 , w_33054 );
and ( \12917_b0 , \5906_b0 , w_33055 );
and ( w_33054 , w_33055 , \7041_b0 );
or ( \12918_b1 , \12916_b1 , w_33057 );
not ( w_33057 , w_33058 );
and ( \12918_b0 , \12916_b0 , w_33059 );
and ( w_33058 ,  , w_33059 );
buf ( w_33057 , \12917_b1 );
not ( w_33057 , w_33060 );
not (  , w_33061 );
and ( w_33060 , w_33061 , \12917_b0 );
or ( \12919_b1 , \12918_b1 , w_33062 );
xor ( \12919_b0 , \12918_b0 , w_33064 );
not ( w_33064 , w_33065 );
and ( w_33065 , w_33062 , w_33063 );
buf ( w_33062 , \7049_b1 );
not ( w_33062 , w_33066 );
not ( w_33063 , w_33067 );
and ( w_33066 , w_33067 , \7049_b0 );
or ( \12920_b1 , \5957_b1 , \7061_b1 );
not ( \7061_b1 , w_33068 );
and ( \12920_b0 , \5957_b0 , w_33069 );
and ( w_33068 , w_33069 , \7061_b0 );
or ( \12921_b1 , \5925_b1 , \7059_b1 );
not ( \7059_b1 , w_33070 );
and ( \12921_b0 , \5925_b0 , w_33071 );
and ( w_33070 , w_33071 , \7059_b0 );
or ( \12922_b1 , \12920_b1 , w_33073 );
not ( w_33073 , w_33074 );
and ( \12922_b0 , \12920_b0 , w_33075 );
and ( w_33074 ,  , w_33075 );
buf ( w_33073 , \12921_b1 );
not ( w_33073 , w_33076 );
not (  , w_33077 );
and ( w_33076 , w_33077 , \12921_b0 );
or ( \12923_b1 , \12922_b1 , w_33078 );
xor ( \12923_b0 , \12922_b0 , w_33080 );
not ( w_33080 , w_33081 );
and ( w_33081 , w_33078 , w_33079 );
buf ( w_33078 , \7067_b1 );
not ( w_33078 , w_33082 );
not ( w_33079 , w_33083 );
and ( w_33082 , w_33083 , \7067_b0 );
or ( \12924_b1 , \12919_b1 , \12923_b1 );
xor ( \12924_b0 , \12919_b0 , w_33084 );
not ( w_33084 , w_33085 );
and ( w_33085 , \12923_b1 , \12923_b0 );
or ( \12925_b1 , \5979_b1 , \7082_b1 );
not ( \7082_b1 , w_33086 );
and ( \12925_b0 , \5979_b0 , w_33087 );
and ( w_33086 , w_33087 , \7082_b0 );
or ( \12926_b1 , \5945_b1 , \7080_b1 );
not ( \7080_b1 , w_33088 );
and ( \12926_b0 , \5945_b0 , w_33089 );
and ( w_33088 , w_33089 , \7080_b0 );
or ( \12927_b1 , \12925_b1 , w_33091 );
not ( w_33091 , w_33092 );
and ( \12927_b0 , \12925_b0 , w_33093 );
and ( w_33092 ,  , w_33093 );
buf ( w_33091 , \12926_b1 );
not ( w_33091 , w_33094 );
not (  , w_33095 );
and ( w_33094 , w_33095 , \12926_b0 );
or ( \12928_b1 , \12927_b1 , w_33096 );
xor ( \12928_b0 , \12927_b0 , w_33098 );
not ( w_33098 , w_33099 );
and ( w_33099 , w_33096 , w_33097 );
buf ( w_33096 , \7088_b1 );
not ( w_33096 , w_33100 );
not ( w_33097 , w_33101 );
and ( w_33100 , w_33101 , \7088_b0 );
or ( \12929_b1 , \12924_b1 , \12928_b1 );
xor ( \12929_b0 , \12924_b0 , w_33102 );
not ( w_33102 , w_33103 );
and ( w_33103 , \12928_b1 , \12928_b0 );
or ( \12930_b1 , \12915_b1 , \12929_b1 );
xor ( \12930_b0 , \12915_b0 , w_33104 );
not ( w_33104 , w_33105 );
and ( w_33105 , \12929_b1 , \12929_b0 );
or ( \12931_b1 , \5873_b1 , \6991_b1 );
not ( \6991_b1 , w_33106 );
and ( \12931_b0 , \5873_b0 , w_33107 );
and ( w_33106 , w_33107 , \6991_b0 );
or ( \12932_b1 , \5842_b1 , \6988_b1 );
not ( \6988_b1 , w_33108 );
and ( \12932_b0 , \5842_b0 , w_33109 );
and ( w_33108 , w_33109 , \6988_b0 );
or ( \12933_b1 , \12931_b1 , w_33111 );
not ( w_33111 , w_33112 );
and ( \12933_b0 , \12931_b0 , w_33113 );
and ( w_33112 ,  , w_33113 );
buf ( w_33111 , \12932_b1 );
not ( w_33111 , w_33114 );
not (  , w_33115 );
and ( w_33114 , w_33115 , \12932_b0 );
or ( \12934_b1 , \12933_b1 , w_33116 );
xor ( \12934_b0 , \12933_b0 , w_33118 );
not ( w_33118 , w_33119 );
and ( w_33119 , w_33116 , w_33117 );
buf ( w_33116 , \6985_b1 );
not ( w_33116 , w_33120 );
not ( w_33117 , w_33121 );
and ( w_33120 , w_33121 , \6985_b0 );
or ( \12935_b1 , \5893_b1 , \7006_b1 );
not ( \7006_b1 , w_33122 );
and ( \12935_b0 , \5893_b0 , w_33123 );
and ( w_33122 , w_33123 , \7006_b0 );
or ( \12936_b1 , \5861_b1 , \7004_b1 );
not ( \7004_b1 , w_33124 );
and ( \12936_b0 , \5861_b0 , w_33125 );
and ( w_33124 , w_33125 , \7004_b0 );
or ( \12937_b1 , \12935_b1 , w_33127 );
not ( w_33127 , w_33128 );
and ( \12937_b0 , \12935_b0 , w_33129 );
and ( w_33128 ,  , w_33129 );
buf ( w_33127 , \12936_b1 );
not ( w_33127 , w_33130 );
not (  , w_33131 );
and ( w_33130 , w_33131 , \12936_b0 );
or ( \12938_b1 , \12937_b1 , w_33132 );
xor ( \12938_b0 , \12937_b0 , w_33134 );
not ( w_33134 , w_33135 );
and ( w_33135 , w_33132 , w_33133 );
buf ( w_33132 , \7012_b1 );
not ( w_33132 , w_33136 );
not ( w_33133 , w_33137 );
and ( w_33136 , w_33137 , \7012_b0 );
or ( \12939_b1 , \12934_b1 , \12938_b1 );
xor ( \12939_b0 , \12934_b0 , w_33138 );
not ( w_33138 , w_33139 );
and ( w_33139 , \12938_b1 , \12938_b0 );
or ( \12940_b1 , \5918_b1 , \7026_b1 );
not ( \7026_b1 , w_33140 );
and ( \12940_b0 , \5918_b0 , w_33141 );
and ( w_33140 , w_33141 , \7026_b0 );
or ( \12941_b1 , \5881_b1 , \7024_b1 );
not ( \7024_b1 , w_33142 );
and ( \12941_b0 , \5881_b0 , w_33143 );
and ( w_33142 , w_33143 , \7024_b0 );
or ( \12942_b1 , \12940_b1 , w_33145 );
not ( w_33145 , w_33146 );
and ( \12942_b0 , \12940_b0 , w_33147 );
and ( w_33146 ,  , w_33147 );
buf ( w_33145 , \12941_b1 );
not ( w_33145 , w_33148 );
not (  , w_33149 );
and ( w_33148 , w_33149 , \12941_b0 );
or ( \12943_b1 , \12942_b1 , w_33150 );
xor ( \12943_b0 , \12942_b0 , w_33152 );
not ( w_33152 , w_33153 );
and ( w_33153 , w_33150 , w_33151 );
buf ( w_33150 , \7032_b1 );
not ( w_33150 , w_33154 );
not ( w_33151 , w_33155 );
and ( w_33154 , w_33155 , \7032_b0 );
or ( \12944_b1 , \12939_b1 , \12943_b1 );
xor ( \12944_b0 , \12939_b0 , w_33156 );
not ( w_33156 , w_33157 );
and ( w_33157 , \12943_b1 , \12943_b0 );
or ( \12945_b1 , \12930_b1 , \12944_b1 );
xor ( \12945_b0 , \12930_b0 , w_33158 );
not ( w_33158 , w_33159 );
and ( w_33159 , \12944_b1 , \12944_b0 );
or ( \12946_b1 , \12901_b1 , \12945_b1 );
xor ( \12946_b0 , \12901_b0 , w_33160 );
not ( w_33160 , w_33161 );
and ( w_33161 , \12945_b1 , \12945_b0 );
or ( \12947_b1 , \12892_b1 , \12946_b1 );
xor ( \12947_b0 , \12892_b0 , w_33162 );
not ( w_33162 , w_33163 );
and ( w_33163 , \12946_b1 , \12946_b0 );
or ( \12948_b1 , \12878_b1 , \12947_b1 );
xor ( \12948_b0 , \12878_b0 , w_33164 );
not ( w_33164 , w_33165 );
and ( w_33165 , \12947_b1 , \12947_b0 );
or ( \12949_b1 , \12850_b1 , \12854_b1 );
not ( \12854_b1 , w_33166 );
and ( \12949_b0 , \12850_b0 , w_33167 );
and ( w_33166 , w_33167 , \12854_b0 );
or ( \12950_b1 , \12854_b1 , \12865_b1 );
not ( \12865_b1 , w_33168 );
and ( \12950_b0 , \12854_b0 , w_33169 );
and ( w_33168 , w_33169 , \12865_b0 );
or ( \12951_b1 , \12850_b1 , \12865_b1 );
not ( \12865_b1 , w_33170 );
and ( \12951_b0 , \12850_b0 , w_33171 );
and ( w_33170 , w_33171 , \12865_b0 );
or ( \12953_b1 , \12830_b1 , \12844_b1 );
not ( \12844_b1 , w_33172 );
and ( \12953_b0 , \12830_b0 , w_33173 );
and ( w_33172 , w_33173 , \12844_b0 );
or ( \12954_b1 , \12952_b1 , \12953_b1 );
xor ( \12954_b0 , \12952_b0 , w_33174 );
not ( w_33174 , w_33175 );
and ( w_33175 , \12953_b1 , \12953_b0 );
or ( \12955_b1 , \12792_b1 , \12796_b1 );
not ( \12796_b1 , w_33176 );
and ( \12955_b0 , \12792_b0 , w_33177 );
and ( w_33176 , w_33177 , \12796_b0 );
or ( \12956_b1 , \12796_b1 , \12799_b1 );
not ( \12799_b1 , w_33178 );
and ( \12956_b0 , \12796_b0 , w_33179 );
and ( w_33178 , w_33179 , \12799_b0 );
or ( \12957_b1 , \12792_b1 , \12799_b1 );
not ( \12799_b1 , w_33180 );
and ( \12957_b0 , \12792_b0 , w_33181 );
and ( w_33180 , w_33181 , \12799_b0 );
or ( \12959_b1 , \6057_b1 , \7157_b1 );
not ( \7157_b1 , w_33182 );
and ( \12959_b0 , \6057_b0 , w_33183 );
and ( w_33182 , w_33183 , \7157_b0 );
or ( \12960_b1 , \6029_b1 , \7155_b1 );
not ( \7155_b1 , w_33184 );
and ( \12960_b0 , \6029_b0 , w_33185 );
and ( w_33184 , w_33185 , \7155_b0 );
or ( \12961_b1 , \12959_b1 , w_33187 );
not ( w_33187 , w_33188 );
and ( \12961_b0 , \12959_b0 , w_33189 );
and ( w_33188 ,  , w_33189 );
buf ( w_33187 , \12960_b1 );
not ( w_33187 , w_33190 );
not (  , w_33191 );
and ( w_33190 , w_33191 , \12960_b0 );
or ( \12962_b1 , \12961_b1 , w_33192 );
xor ( \12962_b0 , \12961_b0 , w_33194 );
not ( w_33194 , w_33195 );
and ( w_33195 , w_33192 , w_33193 );
buf ( w_33192 , \7163_b1 );
not ( w_33192 , w_33196 );
not ( w_33193 , w_33197 );
and ( w_33196 , w_33197 , \7163_b0 );
or ( \12963_b1 , \12958_b1 , \12962_b1 );
xor ( \12963_b0 , \12958_b0 , w_33198 );
not ( w_33198 , w_33199 );
and ( w_33199 , \12962_b1 , \12962_b0 );
or ( \12964_b1 , \6065_b1 , \7175_b1 );
not ( \7175_b1 , w_33200 );
and ( \12964_b0 , \6065_b0 , w_33201 );
and ( w_33200 , w_33201 , \7175_b0 );
or ( \12965_b1 , \6048_b1 , \7173_b1 );
not ( \7173_b1 , w_33202 );
and ( \12965_b0 , \6048_b0 , w_33203 );
and ( w_33202 , w_33203 , \7173_b0 );
or ( \12966_b1 , \12964_b1 , w_33205 );
not ( w_33205 , w_33206 );
and ( \12966_b0 , \12964_b0 , w_33207 );
and ( w_33206 ,  , w_33207 );
buf ( w_33205 , \12965_b1 );
not ( w_33205 , w_33208 );
not (  , w_33209 );
and ( w_33208 , w_33209 , \12965_b0 );
or ( \12967_b1 , \12966_b1 , w_33210 );
xor ( \12967_b0 , \12966_b0 , w_33212 );
not ( w_33212 , w_33213 );
and ( w_33213 , w_33210 , w_33211 );
buf ( w_33210 , \7181_b1 );
not ( w_33210 , w_33214 );
not ( w_33211 , w_33215 );
and ( w_33214 , w_33215 , \7181_b0 );
or ( \12968_b1 , \12963_b1 , \12967_b1 );
xor ( \12968_b0 , \12963_b0 , w_33216 );
not ( w_33216 , w_33217 );
and ( w_33217 , \12967_b1 , \12967_b0 );
or ( \12969_b1 , \12954_b1 , \12968_b1 );
xor ( \12969_b0 , \12954_b0 , w_33218 );
not ( w_33218 , w_33219 );
and ( w_33219 , \12968_b1 , \12968_b0 );
or ( \12970_b1 , \12948_b1 , \12969_b1 );
xor ( \12970_b0 , \12948_b0 , w_33220 );
not ( w_33220 , w_33221 );
and ( w_33221 , \12969_b1 , \12969_b0 );
or ( \12971_b1 , \12782_b1 , \12783_b1 );
not ( \12783_b1 , w_33222 );
and ( \12971_b0 , \12782_b0 , w_33223 );
and ( w_33222 , w_33223 , \12783_b0 );
or ( \12972_b1 , \12783_b1 , \12867_b1 );
not ( \12867_b1 , w_33224 );
and ( \12972_b0 , \12783_b0 , w_33225 );
and ( w_33224 , w_33225 , \12867_b0 );
or ( \12973_b1 , \12782_b1 , \12867_b1 );
not ( \12867_b1 , w_33226 );
and ( \12973_b0 , \12782_b0 , w_33227 );
and ( w_33226 , w_33227 , \12867_b0 );
or ( \12975_b1 , \12970_b1 , w_33229 );
not ( w_33229 , w_33230 );
and ( \12975_b0 , \12970_b0 , w_33231 );
and ( w_33230 ,  , w_33231 );
buf ( w_33229 , \12974_b1 );
not ( w_33229 , w_33232 );
not (  , w_33233 );
and ( w_33232 , w_33233 , \12974_b0 );
or ( \12976_b1 , \12952_b1 , \12953_b1 );
not ( \12953_b1 , w_33234 );
and ( \12976_b0 , \12952_b0 , w_33235 );
and ( w_33234 , w_33235 , \12953_b0 );
or ( \12977_b1 , \12953_b1 , \12968_b1 );
not ( \12968_b1 , w_33236 );
and ( \12977_b0 , \12953_b0 , w_33237 );
and ( w_33236 , w_33237 , \12968_b0 );
or ( \12978_b1 , \12952_b1 , \12968_b1 );
not ( \12968_b1 , w_33238 );
and ( \12978_b0 , \12952_b0 , w_33239 );
and ( w_33238 , w_33239 , \12968_b0 );
or ( \12980_b1 , \12892_b1 , \12946_b1 );
not ( \12946_b1 , w_33240 );
and ( \12980_b0 , \12892_b0 , w_33241 );
and ( w_33240 , w_33241 , \12946_b0 );
or ( \12981_b1 , \12979_b1 , \12980_b1 );
xor ( \12981_b0 , \12979_b0 , w_33242 );
not ( w_33242 , w_33243 );
and ( w_33243 , \12980_b1 , \12980_b0 );
or ( \12982_b1 , \12896_b1 , \12900_b1 );
not ( \12900_b1 , w_33244 );
and ( \12982_b0 , \12896_b0 , w_33245 );
and ( w_33244 , w_33245 , \12900_b0 );
or ( \12983_b1 , \12900_b1 , \12945_b1 );
not ( \12945_b1 , w_33246 );
and ( \12983_b0 , \12900_b0 , w_33247 );
and ( w_33246 , w_33247 , \12945_b0 );
or ( \12984_b1 , \12896_b1 , \12945_b1 );
not ( \12945_b1 , w_33248 );
and ( \12984_b0 , \12896_b0 , w_33249 );
and ( w_33248 , w_33249 , \12945_b0 );
or ( \12986_b1 , \5881_b1 , \7026_b1 );
not ( \7026_b1 , w_33250 );
and ( \12986_b0 , \5881_b0 , w_33251 );
and ( w_33250 , w_33251 , \7026_b0 );
or ( \12987_b1 , \5893_b1 , \7024_b1 );
not ( \7024_b1 , w_33252 );
and ( \12987_b0 , \5893_b0 , w_33253 );
and ( w_33252 , w_33253 , \7024_b0 );
or ( \12988_b1 , \12986_b1 , w_33255 );
not ( w_33255 , w_33256 );
and ( \12988_b0 , \12986_b0 , w_33257 );
and ( w_33256 ,  , w_33257 );
buf ( w_33255 , \12987_b1 );
not ( w_33255 , w_33258 );
not (  , w_33259 );
and ( w_33258 , w_33259 , \12987_b0 );
or ( \12989_b1 , \12988_b1 , w_33260 );
xor ( \12989_b0 , \12988_b0 , w_33262 );
not ( w_33262 , w_33263 );
and ( w_33263 , w_33260 , w_33261 );
buf ( w_33260 , \7032_b1 );
not ( w_33260 , w_33264 );
not ( w_33261 , w_33265 );
and ( w_33264 , w_33265 , \7032_b0 );
or ( \12990_b1 , \5906_b1 , \7043_b1 );
not ( \7043_b1 , w_33266 );
and ( \12990_b0 , \5906_b0 , w_33267 );
and ( w_33266 , w_33267 , \7043_b0 );
or ( \12991_b1 , \5918_b1 , \7041_b1 );
not ( \7041_b1 , w_33268 );
and ( \12991_b0 , \5918_b0 , w_33269 );
and ( w_33268 , w_33269 , \7041_b0 );
or ( \12992_b1 , \12990_b1 , w_33271 );
not ( w_33271 , w_33272 );
and ( \12992_b0 , \12990_b0 , w_33273 );
and ( w_33272 ,  , w_33273 );
buf ( w_33271 , \12991_b1 );
not ( w_33271 , w_33274 );
not (  , w_33275 );
and ( w_33274 , w_33275 , \12991_b0 );
or ( \12993_b1 , \12992_b1 , w_33276 );
xor ( \12993_b0 , \12992_b0 , w_33278 );
not ( w_33278 , w_33279 );
and ( w_33279 , w_33276 , w_33277 );
buf ( w_33276 , \7049_b1 );
not ( w_33276 , w_33280 );
not ( w_33277 , w_33281 );
and ( w_33280 , w_33281 , \7049_b0 );
or ( \12994_b1 , \12989_b1 , \12993_b1 );
xor ( \12994_b0 , \12989_b0 , w_33282 );
not ( w_33282 , w_33283 );
and ( w_33283 , \12993_b1 , \12993_b0 );
or ( \12995_b1 , \5925_b1 , \7061_b1 );
not ( \7061_b1 , w_33284 );
and ( \12995_b0 , \5925_b0 , w_33285 );
and ( w_33284 , w_33285 , \7061_b0 );
or ( \12996_b1 , \5937_b1 , \7059_b1 );
not ( \7059_b1 , w_33286 );
and ( \12996_b0 , \5937_b0 , w_33287 );
and ( w_33286 , w_33287 , \7059_b0 );
or ( \12997_b1 , \12995_b1 , w_33289 );
not ( w_33289 , w_33290 );
and ( \12997_b0 , \12995_b0 , w_33291 );
and ( w_33290 ,  , w_33291 );
buf ( w_33289 , \12996_b1 );
not ( w_33289 , w_33292 );
not (  , w_33293 );
and ( w_33292 , w_33293 , \12996_b0 );
or ( \12998_b1 , \12997_b1 , w_33294 );
xor ( \12998_b0 , \12997_b0 , w_33296 );
not ( w_33296 , w_33297 );
and ( w_33297 , w_33294 , w_33295 );
buf ( w_33294 , \7067_b1 );
not ( w_33294 , w_33298 );
not ( w_33295 , w_33299 );
and ( w_33298 , w_33299 , \7067_b0 );
or ( \12999_b1 , \12994_b1 , \12998_b1 );
xor ( \12999_b0 , \12994_b0 , w_33300 );
not ( w_33300 , w_33301 );
and ( w_33301 , \12998_b1 , \12998_b0 );
or ( \13000_b1 , \5842_b1 , \6991_b1 );
not ( \6991_b1 , w_33302 );
and ( \13000_b0 , \5842_b0 , w_33303 );
and ( w_33302 , w_33303 , \6991_b0 );
or ( \13001_b1 , \5854_b1 , \6988_b1 );
not ( \6988_b1 , w_33304 );
and ( \13001_b0 , \5854_b0 , w_33305 );
and ( w_33304 , w_33305 , \6988_b0 );
or ( \13002_b1 , \13000_b1 , w_33307 );
not ( w_33307 , w_33308 );
and ( \13002_b0 , \13000_b0 , w_33309 );
and ( w_33308 ,  , w_33309 );
buf ( w_33307 , \13001_b1 );
not ( w_33307 , w_33310 );
not (  , w_33311 );
and ( w_33310 , w_33311 , \13001_b0 );
or ( \13003_b1 , \13002_b1 , w_33312 );
xor ( \13003_b0 , \13002_b0 , w_33314 );
not ( w_33314 , w_33315 );
and ( w_33315 , w_33312 , w_33313 );
buf ( w_33312 , \6985_b1 );
not ( w_33312 , w_33316 );
not ( w_33313 , w_33317 );
and ( w_33316 , w_33317 , \6985_b0 );
or ( \13004_b1 , \7198_b1 , \13003_b1 );
xor ( \13004_b0 , \7198_b0 , w_33318 );
not ( w_33318 , w_33319 );
and ( w_33319 , \13003_b1 , \13003_b0 );
or ( \13005_b1 , \5861_b1 , \7006_b1 );
not ( \7006_b1 , w_33320 );
and ( \13005_b0 , \5861_b0 , w_33321 );
and ( w_33320 , w_33321 , \7006_b0 );
or ( \13006_b1 , \5873_b1 , \7004_b1 );
not ( \7004_b1 , w_33322 );
and ( \13006_b0 , \5873_b0 , w_33323 );
and ( w_33322 , w_33323 , \7004_b0 );
or ( \13007_b1 , \13005_b1 , w_33325 );
not ( w_33325 , w_33326 );
and ( \13007_b0 , \13005_b0 , w_33327 );
and ( w_33326 ,  , w_33327 );
buf ( w_33325 , \13006_b1 );
not ( w_33325 , w_33328 );
not (  , w_33329 );
and ( w_33328 , w_33329 , \13006_b0 );
or ( \13008_b1 , \13007_b1 , w_33330 );
xor ( \13008_b0 , \13007_b0 , w_33332 );
not ( w_33332 , w_33333 );
and ( w_33333 , w_33330 , w_33331 );
buf ( w_33330 , \7012_b1 );
not ( w_33330 , w_33334 );
not ( w_33331 , w_33335 );
and ( w_33334 , w_33335 , \7012_b0 );
or ( \13009_b1 , \13004_b1 , \13008_b1 );
xor ( \13009_b0 , \13004_b0 , w_33336 );
not ( w_33336 , w_33337 );
and ( w_33337 , \13008_b1 , \13008_b0 );
or ( \13010_b1 , \12999_b1 , \13009_b1 );
xor ( \13010_b0 , \12999_b0 , w_33338 );
not ( w_33338 , w_33339 );
and ( w_33339 , \13009_b1 , \13009_b0 );
or ( \13011_b1 , \6065_b1 , w_33341 );
not ( w_33341 , w_33342 );
and ( \13011_b0 , \6065_b0 , w_33343 );
and ( w_33342 ,  , w_33343 );
buf ( w_33341 , \7190_b1 );
not ( w_33341 , w_33344 );
not (  , w_33345 );
and ( w_33344 , w_33345 , \7190_b0 );
or ( \13012_b1 , \13011_b1 , w_33346 );
xor ( \13012_b0 , \13011_b0 , w_33348 );
not ( w_33348 , w_33349 );
and ( w_33349 , w_33346 , w_33347 );
buf ( w_33346 , \7198_b1 );
not ( w_33346 , w_33350 );
not ( w_33347 , w_33351 );
and ( w_33350 , w_33351 , \7198_b0 );
or ( \13013_b1 , \6006_b1 , \7140_b1 );
not ( \7140_b1 , w_33352 );
and ( \13013_b0 , \6006_b0 , w_33353 );
and ( w_33352 , w_33353 , \7140_b0 );
or ( \13014_b1 , \6018_b1 , \7138_b1 );
not ( \7138_b1 , w_33354 );
and ( \13014_b0 , \6018_b0 , w_33355 );
and ( w_33354 , w_33355 , \7138_b0 );
or ( \13015_b1 , \13013_b1 , w_33357 );
not ( w_33357 , w_33358 );
and ( \13015_b0 , \13013_b0 , w_33359 );
and ( w_33358 ,  , w_33359 );
buf ( w_33357 , \13014_b1 );
not ( w_33357 , w_33360 );
not (  , w_33361 );
and ( w_33360 , w_33361 , \13014_b0 );
or ( \13016_b1 , \13015_b1 , w_33362 );
xor ( \13016_b0 , \13015_b0 , w_33364 );
not ( w_33364 , w_33365 );
and ( w_33365 , w_33362 , w_33363 );
buf ( w_33362 , \7146_b1 );
not ( w_33362 , w_33366 );
not ( w_33363 , w_33367 );
and ( w_33366 , w_33367 , \7146_b0 );
or ( \13017_b1 , \6029_b1 , \7157_b1 );
not ( \7157_b1 , w_33368 );
and ( \13017_b0 , \6029_b0 , w_33369 );
and ( w_33368 , w_33369 , \7157_b0 );
or ( \13018_b1 , \6041_b1 , \7155_b1 );
not ( \7155_b1 , w_33370 );
and ( \13018_b0 , \6041_b0 , w_33371 );
and ( w_33370 , w_33371 , \7155_b0 );
or ( \13019_b1 , \13017_b1 , w_33373 );
not ( w_33373 , w_33374 );
and ( \13019_b0 , \13017_b0 , w_33375 );
and ( w_33374 ,  , w_33375 );
buf ( w_33373 , \13018_b1 );
not ( w_33373 , w_33376 );
not (  , w_33377 );
and ( w_33376 , w_33377 , \13018_b0 );
or ( \13020_b1 , \13019_b1 , w_33378 );
xor ( \13020_b0 , \13019_b0 , w_33380 );
not ( w_33380 , w_33381 );
and ( w_33381 , w_33378 , w_33379 );
buf ( w_33378 , \7163_b1 );
not ( w_33378 , w_33382 );
not ( w_33379 , w_33383 );
and ( w_33382 , w_33383 , \7163_b0 );
or ( \13021_b1 , \13016_b1 , \13020_b1 );
xor ( \13021_b0 , \13016_b0 , w_33384 );
not ( w_33384 , w_33385 );
and ( w_33385 , \13020_b1 , \13020_b0 );
or ( \13022_b1 , \6048_b1 , \7175_b1 );
not ( \7175_b1 , w_33386 );
and ( \13022_b0 , \6048_b0 , w_33387 );
and ( w_33386 , w_33387 , \7175_b0 );
or ( \13023_b1 , \6057_b1 , \7173_b1 );
not ( \7173_b1 , w_33388 );
and ( \13023_b0 , \6057_b0 , w_33389 );
and ( w_33388 , w_33389 , \7173_b0 );
or ( \13024_b1 , \13022_b1 , w_33391 );
not ( w_33391 , w_33392 );
and ( \13024_b0 , \13022_b0 , w_33393 );
and ( w_33392 ,  , w_33393 );
buf ( w_33391 , \13023_b1 );
not ( w_33391 , w_33394 );
not (  , w_33395 );
and ( w_33394 , w_33395 , \13023_b0 );
or ( \13025_b1 , \13024_b1 , w_33396 );
xor ( \13025_b0 , \13024_b0 , w_33398 );
not ( w_33398 , w_33399 );
and ( w_33399 , w_33396 , w_33397 );
buf ( w_33396 , \7181_b1 );
not ( w_33396 , w_33400 );
not ( w_33397 , w_33401 );
and ( w_33400 , w_33401 , \7181_b0 );
or ( \13026_b1 , \13021_b1 , \13025_b1 );
xor ( \13026_b0 , \13021_b0 , w_33402 );
not ( w_33402 , w_33403 );
and ( w_33403 , \13025_b1 , \13025_b0 );
or ( \13027_b1 , \13012_b1 , \13026_b1 );
xor ( \13027_b0 , \13012_b0 , w_33404 );
not ( w_33404 , w_33405 );
and ( w_33405 , \13026_b1 , \13026_b0 );
or ( \13028_b1 , \5945_b1 , \7082_b1 );
not ( \7082_b1 , w_33406 );
and ( \13028_b0 , \5945_b0 , w_33407 );
and ( w_33406 , w_33407 , \7082_b0 );
or ( \13029_b1 , \5957_b1 , \7080_b1 );
not ( \7080_b1 , w_33408 );
and ( \13029_b0 , \5957_b0 , w_33409 );
and ( w_33408 , w_33409 , \7080_b0 );
or ( \13030_b1 , \13028_b1 , w_33411 );
not ( w_33411 , w_33412 );
and ( \13030_b0 , \13028_b0 , w_33413 );
and ( w_33412 ,  , w_33413 );
buf ( w_33411 , \13029_b1 );
not ( w_33411 , w_33414 );
not (  , w_33415 );
and ( w_33414 , w_33415 , \13029_b0 );
or ( \13031_b1 , \13030_b1 , w_33416 );
xor ( \13031_b0 , \13030_b0 , w_33418 );
not ( w_33418 , w_33419 );
and ( w_33419 , w_33416 , w_33417 );
buf ( w_33416 , \7088_b1 );
not ( w_33416 , w_33420 );
not ( w_33417 , w_33421 );
and ( w_33420 , w_33421 , \7088_b0 );
or ( \13032_b1 , \5967_b1 , \7099_b1 );
not ( \7099_b1 , w_33422 );
and ( \13032_b0 , \5967_b0 , w_33423 );
and ( w_33422 , w_33423 , \7099_b0 );
or ( \13033_b1 , \5979_b1 , \7097_b1 );
not ( \7097_b1 , w_33424 );
and ( \13033_b0 , \5979_b0 , w_33425 );
and ( w_33424 , w_33425 , \7097_b0 );
or ( \13034_b1 , \13032_b1 , w_33427 );
not ( w_33427 , w_33428 );
and ( \13034_b0 , \13032_b0 , w_33429 );
and ( w_33428 ,  , w_33429 );
buf ( w_33427 , \13033_b1 );
not ( w_33427 , w_33430 );
not (  , w_33431 );
and ( w_33430 , w_33431 , \13033_b0 );
or ( \13035_b1 , \13034_b1 , w_33432 );
xor ( \13035_b0 , \13034_b0 , w_33434 );
not ( w_33434 , w_33435 );
and ( w_33435 , w_33432 , w_33433 );
buf ( w_33432 , \7105_b1 );
not ( w_33432 , w_33436 );
not ( w_33433 , w_33437 );
and ( w_33436 , w_33437 , \7105_b0 );
or ( \13036_b1 , \13031_b1 , \13035_b1 );
xor ( \13036_b0 , \13031_b0 , w_33438 );
not ( w_33438 , w_33439 );
and ( w_33439 , \13035_b1 , \13035_b0 );
or ( \13037_b1 , \5986_b1 , \7117_b1 );
not ( \7117_b1 , w_33440 );
and ( \13037_b0 , \5986_b0 , w_33441 );
and ( w_33440 , w_33441 , \7117_b0 );
or ( \13038_b1 , \5998_b1 , \7115_b1 );
not ( \7115_b1 , w_33442 );
and ( \13038_b0 , \5998_b0 , w_33443 );
and ( w_33442 , w_33443 , \7115_b0 );
or ( \13039_b1 , \13037_b1 , w_33445 );
not ( w_33445 , w_33446 );
and ( \13039_b0 , \13037_b0 , w_33447 );
and ( w_33446 ,  , w_33447 );
buf ( w_33445 , \13038_b1 );
not ( w_33445 , w_33448 );
not (  , w_33449 );
and ( w_33448 , w_33449 , \13038_b0 );
or ( \13040_b1 , \13039_b1 , w_33450 );
xor ( \13040_b0 , \13039_b0 , w_33452 );
not ( w_33452 , w_33453 );
and ( w_33453 , w_33450 , w_33451 );
buf ( w_33450 , \7123_b1 );
not ( w_33450 , w_33454 );
not ( w_33451 , w_33455 );
and ( w_33454 , w_33455 , \7123_b0 );
or ( \13041_b1 , \13036_b1 , \13040_b1 );
xor ( \13041_b0 , \13036_b0 , w_33456 );
not ( w_33456 , w_33457 );
and ( w_33457 , \13040_b1 , \13040_b0 );
or ( \13042_b1 , \13027_b1 , \13041_b1 );
xor ( \13042_b0 , \13027_b0 , w_33458 );
not ( w_33458 , w_33459 );
and ( w_33459 , \13041_b1 , \13041_b0 );
or ( \13043_b1 , \13010_b1 , \13042_b1 );
xor ( \13043_b0 , \13010_b0 , w_33460 );
not ( w_33460 , w_33461 );
and ( w_33461 , \13042_b1 , \13042_b0 );
or ( \13044_b1 , \12934_b1 , \12938_b1 );
not ( \12938_b1 , w_33462 );
and ( \13044_b0 , \12934_b0 , w_33463 );
and ( w_33462 , w_33463 , \12938_b0 );
or ( \13045_b1 , \12938_b1 , \12943_b1 );
not ( \12943_b1 , w_33464 );
and ( \13045_b0 , \12938_b0 , w_33465 );
and ( w_33464 , w_33465 , \12943_b0 );
or ( \13046_b1 , \12934_b1 , \12943_b1 );
not ( \12943_b1 , w_33466 );
and ( \13046_b0 , \12934_b0 , w_33467 );
and ( w_33466 , w_33467 , \12943_b0 );
or ( \13048_b1 , \12919_b1 , \12923_b1 );
not ( \12923_b1 , w_33468 );
and ( \13048_b0 , \12919_b0 , w_33469 );
and ( w_33468 , w_33469 , \12923_b0 );
or ( \13049_b1 , \12923_b1 , \12928_b1 );
not ( \12928_b1 , w_33470 );
and ( \13049_b0 , \12923_b0 , w_33471 );
and ( w_33470 , w_33471 , \12928_b0 );
or ( \13050_b1 , \12919_b1 , \12928_b1 );
not ( \12928_b1 , w_33472 );
and ( \13050_b0 , \12919_b0 , w_33473 );
and ( w_33472 , w_33473 , \12928_b0 );
or ( \13052_b1 , \13047_b1 , \13051_b1 );
xor ( \13052_b0 , \13047_b0 , w_33474 );
not ( w_33474 , w_33475 );
and ( w_33475 , \13051_b1 , \13051_b0 );
or ( \13053_b1 , \12905_b1 , \12909_b1 );
not ( \12909_b1 , w_33476 );
and ( \13053_b0 , \12905_b0 , w_33477 );
and ( w_33476 , w_33477 , \12909_b0 );
or ( \13054_b1 , \12909_b1 , \12914_b1 );
not ( \12914_b1 , w_33478 );
and ( \13054_b0 , \12909_b0 , w_33479 );
and ( w_33478 , w_33479 , \12914_b0 );
or ( \13055_b1 , \12905_b1 , \12914_b1 );
not ( \12914_b1 , w_33480 );
and ( \13055_b0 , \12905_b0 , w_33481 );
and ( w_33480 , w_33481 , \12914_b0 );
or ( \13057_b1 , \13052_b1 , \13056_b1 );
xor ( \13057_b0 , \13052_b0 , w_33482 );
not ( w_33482 , w_33483 );
and ( w_33483 , \13056_b1 , \13056_b0 );
or ( \13058_b1 , \13043_b1 , \13057_b1 );
xor ( \13058_b0 , \13043_b0 , w_33484 );
not ( w_33484 , w_33485 );
and ( w_33485 , \13057_b1 , \13057_b0 );
or ( \13059_b1 , \12985_b1 , \13058_b1 );
xor ( \13059_b0 , \12985_b0 , w_33486 );
not ( w_33486 , w_33487 );
and ( w_33487 , \13058_b1 , \13058_b0 );
or ( \13060_b1 , \12882_b1 , \12886_b1 );
not ( \12886_b1 , w_33488 );
and ( \13060_b0 , \12882_b0 , w_33489 );
and ( w_33488 , w_33489 , \12886_b0 );
or ( \13061_b1 , \12886_b1 , \12891_b1 );
not ( \12891_b1 , w_33490 );
and ( \13061_b0 , \12886_b0 , w_33491 );
and ( w_33490 , w_33491 , \12891_b0 );
or ( \13062_b1 , \12882_b1 , \12891_b1 );
not ( \12891_b1 , w_33492 );
and ( \13062_b0 , \12882_b0 , w_33493 );
and ( w_33492 , w_33493 , \12891_b0 );
or ( \13064_b1 , \12958_b1 , \12962_b1 );
not ( \12962_b1 , w_33494 );
and ( \13064_b0 , \12958_b0 , w_33495 );
and ( w_33494 , w_33495 , \12962_b0 );
or ( \13065_b1 , \12962_b1 , \12967_b1 );
not ( \12967_b1 , w_33496 );
and ( \13065_b0 , \12962_b0 , w_33497 );
and ( w_33496 , w_33497 , \12967_b0 );
or ( \13066_b1 , \12958_b1 , \12967_b1 );
not ( \12967_b1 , w_33498 );
and ( \13066_b0 , \12958_b0 , w_33499 );
and ( w_33498 , w_33499 , \12967_b0 );
or ( \13068_b1 , \13063_b1 , \13067_b1 );
xor ( \13068_b0 , \13063_b0 , w_33500 );
not ( w_33500 , w_33501 );
and ( w_33501 , \13067_b1 , \13067_b0 );
or ( \13069_b1 , \12915_b1 , \12929_b1 );
not ( \12929_b1 , w_33502 );
and ( \13069_b0 , \12915_b0 , w_33503 );
and ( w_33502 , w_33503 , \12929_b0 );
or ( \13070_b1 , \12929_b1 , \12944_b1 );
not ( \12944_b1 , w_33504 );
and ( \13070_b0 , \12929_b0 , w_33505 );
and ( w_33504 , w_33505 , \12944_b0 );
or ( \13071_b1 , \12915_b1 , \12944_b1 );
not ( \12944_b1 , w_33506 );
and ( \13071_b0 , \12915_b0 , w_33507 );
and ( w_33506 , w_33507 , \12944_b0 );
or ( \13073_b1 , \13068_b1 , \13072_b1 );
xor ( \13073_b0 , \13068_b0 , w_33508 );
not ( w_33508 , w_33509 );
and ( w_33509 , \13072_b1 , \13072_b0 );
or ( \13074_b1 , \13059_b1 , \13073_b1 );
xor ( \13074_b0 , \13059_b0 , w_33510 );
not ( w_33510 , w_33511 );
and ( w_33511 , \13073_b1 , \13073_b0 );
or ( \13075_b1 , \12981_b1 , \13074_b1 );
xor ( \13075_b0 , \12981_b0 , w_33512 );
not ( w_33512 , w_33513 );
and ( w_33513 , \13074_b1 , \13074_b0 );
or ( \13076_b1 , \12878_b1 , \12947_b1 );
not ( \12947_b1 , w_33514 );
and ( \13076_b0 , \12878_b0 , w_33515 );
and ( w_33514 , w_33515 , \12947_b0 );
or ( \13077_b1 , \12947_b1 , \12969_b1 );
not ( \12969_b1 , w_33516 );
and ( \13077_b0 , \12947_b0 , w_33517 );
and ( w_33516 , w_33517 , \12969_b0 );
or ( \13078_b1 , \12878_b1 , \12969_b1 );
not ( \12969_b1 , w_33518 );
and ( \13078_b0 , \12878_b0 , w_33519 );
and ( w_33518 , w_33519 , \12969_b0 );
or ( \13080_b1 , \13075_b1 , w_33521 );
not ( w_33521 , w_33522 );
and ( \13080_b0 , \13075_b0 , w_33523 );
and ( w_33522 ,  , w_33523 );
buf ( w_33521 , \13079_b1 );
not ( w_33521 , w_33524 );
not (  , w_33525 );
and ( w_33524 , w_33525 , \13079_b0 );
or ( \13081_b1 , \12975_b1 , w_33527 );
not ( w_33527 , w_33528 );
and ( \13081_b0 , \12975_b0 , w_33529 );
and ( w_33528 ,  , w_33529 );
buf ( w_33527 , \13080_b1 );
not ( w_33527 , w_33530 );
not (  , w_33531 );
and ( w_33530 , w_33531 , \13080_b0 );
or ( \13082_b1 , \12874_b1 , w_33533 );
not ( w_33533 , w_33534 );
and ( \13082_b0 , \12874_b0 , w_33535 );
and ( w_33534 ,  , w_33535 );
buf ( w_33533 , \13081_b1 );
not ( w_33533 , w_33536 );
not (  , w_33537 );
and ( w_33536 , w_33537 , \13081_b0 );
or ( \13083_b1 , \12687_b1 , w_33539 );
not ( w_33539 , w_33540 );
and ( \13083_b0 , \12687_b0 , w_33541 );
and ( w_33540 ,  , w_33541 );
buf ( w_33539 , \13082_b1 );
not ( w_33539 , w_33542 );
not (  , w_33543 );
and ( w_33542 , w_33543 , \13082_b0 );
or ( \13084_b1 , \12985_b1 , \13058_b1 );
not ( \13058_b1 , w_33544 );
and ( \13084_b0 , \12985_b0 , w_33545 );
and ( w_33544 , w_33545 , \13058_b0 );
or ( \13085_b1 , \13058_b1 , \13073_b1 );
not ( \13073_b1 , w_33546 );
and ( \13085_b0 , \13058_b0 , w_33547 );
and ( w_33546 , w_33547 , \13073_b0 );
or ( \13086_b1 , \12985_b1 , \13073_b1 );
not ( \13073_b1 , w_33548 );
and ( \13086_b0 , \12985_b0 , w_33549 );
and ( w_33548 , w_33549 , \13073_b0 );
or ( \13088_b1 , \13047_b1 , \13051_b1 );
not ( \13051_b1 , w_33550 );
and ( \13088_b0 , \13047_b0 , w_33551 );
and ( w_33550 , w_33551 , \13051_b0 );
or ( \13089_b1 , \13051_b1 , \13056_b1 );
not ( \13056_b1 , w_33552 );
and ( \13089_b0 , \13051_b0 , w_33553 );
and ( w_33552 , w_33553 , \13056_b0 );
or ( \13090_b1 , \13047_b1 , \13056_b1 );
not ( \13056_b1 , w_33554 );
and ( \13090_b0 , \13047_b0 , w_33555 );
and ( w_33554 , w_33555 , \13056_b0 );
or ( \13092_b1 , \13012_b1 , \13026_b1 );
not ( \13026_b1 , w_33556 );
and ( \13092_b0 , \13012_b0 , w_33557 );
and ( w_33556 , w_33557 , \13026_b0 );
or ( \13093_b1 , \13026_b1 , \13041_b1 );
not ( \13041_b1 , w_33558 );
and ( \13093_b0 , \13026_b0 , w_33559 );
and ( w_33558 , w_33559 , \13041_b0 );
or ( \13094_b1 , \13012_b1 , \13041_b1 );
not ( \13041_b1 , w_33560 );
and ( \13094_b0 , \13012_b0 , w_33561 );
and ( w_33560 , w_33561 , \13041_b0 );
or ( \13096_b1 , \13091_b1 , \13095_b1 );
xor ( \13096_b0 , \13091_b0 , w_33562 );
not ( w_33562 , w_33563 );
and ( w_33563 , \13095_b1 , \13095_b0 );
or ( \13097_b1 , \12999_b1 , \13009_b1 );
not ( \13009_b1 , w_33564 );
and ( \13097_b0 , \12999_b0 , w_33565 );
and ( w_33564 , w_33565 , \13009_b0 );
or ( \13098_b1 , \13096_b1 , \13097_b1 );
xor ( \13098_b0 , \13096_b0 , w_33566 );
not ( w_33566 , w_33567 );
and ( w_33567 , \13097_b1 , \13097_b0 );
or ( \13099_b1 , \13087_b1 , \13098_b1 );
xor ( \13099_b0 , \13087_b0 , w_33568 );
not ( w_33568 , w_33569 );
and ( w_33569 , \13098_b1 , \13098_b0 );
or ( \13100_b1 , \13063_b1 , \13067_b1 );
not ( \13067_b1 , w_33570 );
and ( \13100_b0 , \13063_b0 , w_33571 );
and ( w_33570 , w_33571 , \13067_b0 );
or ( \13101_b1 , \13067_b1 , \13072_b1 );
not ( \13072_b1 , w_33572 );
and ( \13101_b0 , \13067_b0 , w_33573 );
and ( w_33572 , w_33573 , \13072_b0 );
or ( \13102_b1 , \13063_b1 , \13072_b1 );
not ( \13072_b1 , w_33574 );
and ( \13102_b0 , \13063_b0 , w_33575 );
and ( w_33574 , w_33575 , \13072_b0 );
or ( \13104_b1 , \13010_b1 , \13042_b1 );
not ( \13042_b1 , w_33576 );
and ( \13104_b0 , \13010_b0 , w_33577 );
and ( w_33576 , w_33577 , \13042_b0 );
or ( \13105_b1 , \13042_b1 , \13057_b1 );
not ( \13057_b1 , w_33578 );
and ( \13105_b0 , \13042_b0 , w_33579 );
and ( w_33578 , w_33579 , \13057_b0 );
or ( \13106_b1 , \13010_b1 , \13057_b1 );
not ( \13057_b1 , w_33580 );
and ( \13106_b0 , \13010_b0 , w_33581 );
and ( w_33580 , w_33581 , \13057_b0 );
or ( \13108_b1 , \13103_b1 , \13107_b1 );
xor ( \13108_b0 , \13103_b0 , w_33582 );
not ( w_33582 , w_33583 );
and ( w_33583 , \13107_b1 , \13107_b0 );
or ( \13109_b1 , \5918_b1 , \7043_b1 );
not ( \7043_b1 , w_33584 );
and ( \13109_b0 , \5918_b0 , w_33585 );
and ( w_33584 , w_33585 , \7043_b0 );
or ( \13110_b1 , \5881_b1 , \7041_b1 );
not ( \7041_b1 , w_33586 );
and ( \13110_b0 , \5881_b0 , w_33587 );
and ( w_33586 , w_33587 , \7041_b0 );
or ( \13111_b1 , \13109_b1 , w_33589 );
not ( w_33589 , w_33590 );
and ( \13111_b0 , \13109_b0 , w_33591 );
and ( w_33590 ,  , w_33591 );
buf ( w_33589 , \13110_b1 );
not ( w_33589 , w_33592 );
not (  , w_33593 );
and ( w_33592 , w_33593 , \13110_b0 );
or ( \13112_b1 , \13111_b1 , w_33594 );
xor ( \13112_b0 , \13111_b0 , w_33596 );
not ( w_33596 , w_33597 );
and ( w_33597 , w_33594 , w_33595 );
buf ( w_33594 , \7049_b1 );
not ( w_33594 , w_33598 );
not ( w_33595 , w_33599 );
and ( w_33598 , w_33599 , \7049_b0 );
or ( \13113_b1 , \5937_b1 , \7061_b1 );
not ( \7061_b1 , w_33600 );
and ( \13113_b0 , \5937_b0 , w_33601 );
and ( w_33600 , w_33601 , \7061_b0 );
or ( \13114_b1 , \5906_b1 , \7059_b1 );
not ( \7059_b1 , w_33602 );
and ( \13114_b0 , \5906_b0 , w_33603 );
and ( w_33602 , w_33603 , \7059_b0 );
or ( \13115_b1 , \13113_b1 , w_33605 );
not ( w_33605 , w_33606 );
and ( \13115_b0 , \13113_b0 , w_33607 );
and ( w_33606 ,  , w_33607 );
buf ( w_33605 , \13114_b1 );
not ( w_33605 , w_33608 );
not (  , w_33609 );
and ( w_33608 , w_33609 , \13114_b0 );
or ( \13116_b1 , \13115_b1 , w_33610 );
xor ( \13116_b0 , \13115_b0 , w_33612 );
not ( w_33612 , w_33613 );
and ( w_33613 , w_33610 , w_33611 );
buf ( w_33610 , \7067_b1 );
not ( w_33610 , w_33614 );
not ( w_33611 , w_33615 );
and ( w_33614 , w_33615 , \7067_b0 );
or ( \13117_b1 , \13112_b1 , \13116_b1 );
xor ( \13117_b0 , \13112_b0 , w_33616 );
not ( w_33616 , w_33617 );
and ( w_33617 , \13116_b1 , \13116_b0 );
or ( \13118_b1 , \5957_b1 , \7082_b1 );
not ( \7082_b1 , w_33618 );
and ( \13118_b0 , \5957_b0 , w_33619 );
and ( w_33618 , w_33619 , \7082_b0 );
or ( \13119_b1 , \5925_b1 , \7080_b1 );
not ( \7080_b1 , w_33620 );
and ( \13119_b0 , \5925_b0 , w_33621 );
and ( w_33620 , w_33621 , \7080_b0 );
or ( \13120_b1 , \13118_b1 , w_33623 );
not ( w_33623 , w_33624 );
and ( \13120_b0 , \13118_b0 , w_33625 );
and ( w_33624 ,  , w_33625 );
buf ( w_33623 , \13119_b1 );
not ( w_33623 , w_33626 );
not (  , w_33627 );
and ( w_33626 , w_33627 , \13119_b0 );
or ( \13121_b1 , \13120_b1 , w_33628 );
xor ( \13121_b0 , \13120_b0 , w_33630 );
not ( w_33630 , w_33631 );
and ( w_33631 , w_33628 , w_33629 );
buf ( w_33628 , \7088_b1 );
not ( w_33628 , w_33632 );
not ( w_33629 , w_33633 );
and ( w_33632 , w_33633 , \7088_b0 );
or ( \13122_b1 , \13117_b1 , \13121_b1 );
xor ( \13122_b0 , \13117_b0 , w_33634 );
not ( w_33634 , w_33635 );
and ( w_33635 , \13121_b1 , \13121_b0 );
or ( \13123_b1 , \5854_b1 , \6991_b1 );
not ( \6991_b1 , w_33636 );
and ( \13123_b0 , \5854_b0 , w_33637 );
and ( w_33636 , w_33637 , \6991_b0 );
or ( \13124_b1 , \5819_b1 , \6988_b1 );
not ( \6988_b1 , w_33638 );
and ( \13124_b0 , \5819_b0 , w_33639 );
and ( w_33638 , w_33639 , \6988_b0 );
or ( \13125_b1 , \13123_b1 , w_33641 );
not ( w_33641 , w_33642 );
and ( \13125_b0 , \13123_b0 , w_33643 );
and ( w_33642 ,  , w_33643 );
buf ( w_33641 , \13124_b1 );
not ( w_33641 , w_33644 );
not (  , w_33645 );
and ( w_33644 , w_33645 , \13124_b0 );
or ( \13126_b1 , \13125_b1 , w_33646 );
xor ( \13126_b0 , \13125_b0 , w_33648 );
not ( w_33648 , w_33649 );
and ( w_33649 , w_33646 , w_33647 );
buf ( w_33646 , \6985_b1 );
not ( w_33646 , w_33650 );
not ( w_33647 , w_33651 );
and ( w_33650 , w_33651 , \6985_b0 );
or ( \13127_b1 , \5873_b1 , \7006_b1 );
not ( \7006_b1 , w_33652 );
and ( \13127_b0 , \5873_b0 , w_33653 );
and ( w_33652 , w_33653 , \7006_b0 );
or ( \13128_b1 , \5842_b1 , \7004_b1 );
not ( \7004_b1 , w_33654 );
and ( \13128_b0 , \5842_b0 , w_33655 );
and ( w_33654 , w_33655 , \7004_b0 );
or ( \13129_b1 , \13127_b1 , w_33657 );
not ( w_33657 , w_33658 );
and ( \13129_b0 , \13127_b0 , w_33659 );
and ( w_33658 ,  , w_33659 );
buf ( w_33657 , \13128_b1 );
not ( w_33657 , w_33660 );
not (  , w_33661 );
and ( w_33660 , w_33661 , \13128_b0 );
or ( \13130_b1 , \13129_b1 , w_33662 );
xor ( \13130_b0 , \13129_b0 , w_33664 );
not ( w_33664 , w_33665 );
and ( w_33665 , w_33662 , w_33663 );
buf ( w_33662 , \7012_b1 );
not ( w_33662 , w_33666 );
not ( w_33663 , w_33667 );
and ( w_33666 , w_33667 , \7012_b0 );
or ( \13131_b1 , \13126_b1 , \13130_b1 );
xor ( \13131_b0 , \13126_b0 , w_33668 );
not ( w_33668 , w_33669 );
and ( w_33669 , \13130_b1 , \13130_b0 );
or ( \13132_b1 , \5893_b1 , \7026_b1 );
not ( \7026_b1 , w_33670 );
and ( \13132_b0 , \5893_b0 , w_33671 );
and ( w_33670 , w_33671 , \7026_b0 );
or ( \13133_b1 , \5861_b1 , \7024_b1 );
not ( \7024_b1 , w_33672 );
and ( \13133_b0 , \5861_b0 , w_33673 );
and ( w_33672 , w_33673 , \7024_b0 );
or ( \13134_b1 , \13132_b1 , w_33675 );
not ( w_33675 , w_33676 );
and ( \13134_b0 , \13132_b0 , w_33677 );
and ( w_33676 ,  , w_33677 );
buf ( w_33675 , \13133_b1 );
not ( w_33675 , w_33678 );
not (  , w_33679 );
and ( w_33678 , w_33679 , \13133_b0 );
or ( \13135_b1 , \13134_b1 , w_33680 );
xor ( \13135_b0 , \13134_b0 , w_33682 );
not ( w_33682 , w_33683 );
and ( w_33683 , w_33680 , w_33681 );
buf ( w_33680 , \7032_b1 );
not ( w_33680 , w_33684 );
not ( w_33681 , w_33685 );
and ( w_33684 , w_33685 , \7032_b0 );
or ( \13136_b1 , \13131_b1 , \13135_b1 );
xor ( \13136_b0 , \13131_b0 , w_33686 );
not ( w_33686 , w_33687 );
and ( w_33687 , \13135_b1 , \13135_b0 );
or ( \13137_b1 , \13122_b1 , \13136_b1 );
xor ( \13137_b0 , \13122_b0 , w_33688 );
not ( w_33688 , w_33689 );
and ( w_33689 , \13136_b1 , \13136_b0 );
or ( \13138_b1 , \13016_b1 , \13020_b1 );
not ( \13020_b1 , w_33690 );
and ( \13138_b0 , \13016_b0 , w_33691 );
and ( w_33690 , w_33691 , \13020_b0 );
or ( \13139_b1 , \13020_b1 , \13025_b1 );
not ( \13025_b1 , w_33692 );
and ( \13139_b0 , \13020_b0 , w_33693 );
and ( w_33692 , w_33693 , \13025_b0 );
or ( \13140_b1 , \13016_b1 , \13025_b1 );
not ( \13025_b1 , w_33694 );
and ( \13140_b0 , \13016_b0 , w_33695 );
and ( w_33694 , w_33695 , \13025_b0 );
or ( \13142_b1 , \6041_b1 , \7157_b1 );
not ( \7157_b1 , w_33696 );
and ( \13142_b0 , \6041_b0 , w_33697 );
and ( w_33696 , w_33697 , \7157_b0 );
or ( \13143_b1 , \6006_b1 , \7155_b1 );
not ( \7155_b1 , w_33698 );
and ( \13143_b0 , \6006_b0 , w_33699 );
and ( w_33698 , w_33699 , \7155_b0 );
or ( \13144_b1 , \13142_b1 , w_33701 );
not ( w_33701 , w_33702 );
and ( \13144_b0 , \13142_b0 , w_33703 );
and ( w_33702 ,  , w_33703 );
buf ( w_33701 , \13143_b1 );
not ( w_33701 , w_33704 );
not (  , w_33705 );
and ( w_33704 , w_33705 , \13143_b0 );
or ( \13145_b1 , \13144_b1 , w_33706 );
xor ( \13145_b0 , \13144_b0 , w_33708 );
not ( w_33708 , w_33709 );
and ( w_33709 , w_33706 , w_33707 );
buf ( w_33706 , \7163_b1 );
not ( w_33706 , w_33710 );
not ( w_33707 , w_33711 );
and ( w_33710 , w_33711 , \7163_b0 );
or ( \13146_b1 , \6057_b1 , \7175_b1 );
not ( \7175_b1 , w_33712 );
and ( \13146_b0 , \6057_b0 , w_33713 );
and ( w_33712 , w_33713 , \7175_b0 );
or ( \13147_b1 , \6029_b1 , \7173_b1 );
not ( \7173_b1 , w_33714 );
and ( \13147_b0 , \6029_b0 , w_33715 );
and ( w_33714 , w_33715 , \7173_b0 );
or ( \13148_b1 , \13146_b1 , w_33717 );
not ( w_33717 , w_33718 );
and ( \13148_b0 , \13146_b0 , w_33719 );
and ( w_33718 ,  , w_33719 );
buf ( w_33717 , \13147_b1 );
not ( w_33717 , w_33720 );
not (  , w_33721 );
and ( w_33720 , w_33721 , \13147_b0 );
or ( \13149_b1 , \13148_b1 , w_33722 );
xor ( \13149_b0 , \13148_b0 , w_33724 );
not ( w_33724 , w_33725 );
and ( w_33725 , w_33722 , w_33723 );
buf ( w_33722 , \7181_b1 );
not ( w_33722 , w_33726 );
not ( w_33723 , w_33727 );
and ( w_33726 , w_33727 , \7181_b0 );
or ( \13150_b1 , \13145_b1 , \13149_b1 );
xor ( \13150_b0 , \13145_b0 , w_33728 );
not ( w_33728 , w_33729 );
and ( w_33729 , \13149_b1 , \13149_b0 );
or ( \13151_b1 , \6065_b1 , \7192_b1 );
not ( \7192_b1 , w_33730 );
and ( \13151_b0 , \6065_b0 , w_33731 );
and ( w_33730 , w_33731 , \7192_b0 );
or ( \13152_b1 , \6048_b1 , \7190_b1 );
not ( \7190_b1 , w_33732 );
and ( \13152_b0 , \6048_b0 , w_33733 );
and ( w_33732 , w_33733 , \7190_b0 );
or ( \13153_b1 , \13151_b1 , w_33735 );
not ( w_33735 , w_33736 );
and ( \13153_b0 , \13151_b0 , w_33737 );
and ( w_33736 ,  , w_33737 );
buf ( w_33735 , \13152_b1 );
not ( w_33735 , w_33738 );
not (  , w_33739 );
and ( w_33738 , w_33739 , \13152_b0 );
or ( \13154_b1 , \13153_b1 , w_33740 );
xor ( \13154_b0 , \13153_b0 , w_33742 );
not ( w_33742 , w_33743 );
and ( w_33743 , w_33740 , w_33741 );
buf ( w_33740 , \7198_b1 );
not ( w_33740 , w_33744 );
not ( w_33741 , w_33745 );
and ( w_33744 , w_33745 , \7198_b0 );
or ( \13155_b1 , \13150_b1 , \13154_b1 );
xor ( \13155_b0 , \13150_b0 , w_33746 );
not ( w_33746 , w_33747 );
and ( w_33747 , \13154_b1 , \13154_b0 );
or ( \13156_b1 , \13141_b1 , \13155_b1 );
xor ( \13156_b0 , \13141_b0 , w_33748 );
not ( w_33748 , w_33749 );
and ( w_33749 , \13155_b1 , \13155_b0 );
or ( \13157_b1 , \5979_b1 , \7099_b1 );
not ( \7099_b1 , w_33750 );
and ( \13157_b0 , \5979_b0 , w_33751 );
and ( w_33750 , w_33751 , \7099_b0 );
or ( \13158_b1 , \5945_b1 , \7097_b1 );
not ( \7097_b1 , w_33752 );
and ( \13158_b0 , \5945_b0 , w_33753 );
and ( w_33752 , w_33753 , \7097_b0 );
or ( \13159_b1 , \13157_b1 , w_33755 );
not ( w_33755 , w_33756 );
and ( \13159_b0 , \13157_b0 , w_33757 );
and ( w_33756 ,  , w_33757 );
buf ( w_33755 , \13158_b1 );
not ( w_33755 , w_33758 );
not (  , w_33759 );
and ( w_33758 , w_33759 , \13158_b0 );
or ( \13160_b1 , \13159_b1 , w_33760 );
xor ( \13160_b0 , \13159_b0 , w_33762 );
not ( w_33762 , w_33763 );
and ( w_33763 , w_33760 , w_33761 );
buf ( w_33760 , \7105_b1 );
not ( w_33760 , w_33764 );
not ( w_33761 , w_33765 );
and ( w_33764 , w_33765 , \7105_b0 );
or ( \13161_b1 , \5998_b1 , \7117_b1 );
not ( \7117_b1 , w_33766 );
and ( \13161_b0 , \5998_b0 , w_33767 );
and ( w_33766 , w_33767 , \7117_b0 );
or ( \13162_b1 , \5967_b1 , \7115_b1 );
not ( \7115_b1 , w_33768 );
and ( \13162_b0 , \5967_b0 , w_33769 );
and ( w_33768 , w_33769 , \7115_b0 );
or ( \13163_b1 , \13161_b1 , w_33771 );
not ( w_33771 , w_33772 );
and ( \13163_b0 , \13161_b0 , w_33773 );
and ( w_33772 ,  , w_33773 );
buf ( w_33771 , \13162_b1 );
not ( w_33771 , w_33774 );
not (  , w_33775 );
and ( w_33774 , w_33775 , \13162_b0 );
or ( \13164_b1 , \13163_b1 , w_33776 );
xor ( \13164_b0 , \13163_b0 , w_33778 );
not ( w_33778 , w_33779 );
and ( w_33779 , w_33776 , w_33777 );
buf ( w_33776 , \7123_b1 );
not ( w_33776 , w_33780 );
not ( w_33777 , w_33781 );
and ( w_33780 , w_33781 , \7123_b0 );
or ( \13165_b1 , \13160_b1 , \13164_b1 );
xor ( \13165_b0 , \13160_b0 , w_33782 );
not ( w_33782 , w_33783 );
and ( w_33783 , \13164_b1 , \13164_b0 );
or ( \13166_b1 , \6018_b1 , \7140_b1 );
not ( \7140_b1 , w_33784 );
and ( \13166_b0 , \6018_b0 , w_33785 );
and ( w_33784 , w_33785 , \7140_b0 );
or ( \13167_b1 , \5986_b1 , \7138_b1 );
not ( \7138_b1 , w_33786 );
and ( \13167_b0 , \5986_b0 , w_33787 );
and ( w_33786 , w_33787 , \7138_b0 );
or ( \13168_b1 , \13166_b1 , w_33789 );
not ( w_33789 , w_33790 );
and ( \13168_b0 , \13166_b0 , w_33791 );
and ( w_33790 ,  , w_33791 );
buf ( w_33789 , \13167_b1 );
not ( w_33789 , w_33792 );
not (  , w_33793 );
and ( w_33792 , w_33793 , \13167_b0 );
or ( \13169_b1 , \13168_b1 , w_33794 );
xor ( \13169_b0 , \13168_b0 , w_33796 );
not ( w_33796 , w_33797 );
and ( w_33797 , w_33794 , w_33795 );
buf ( w_33794 , \7146_b1 );
not ( w_33794 , w_33798 );
not ( w_33795 , w_33799 );
and ( w_33798 , w_33799 , \7146_b0 );
or ( \13170_b1 , \13165_b1 , \13169_b1 );
xor ( \13170_b0 , \13165_b0 , w_33800 );
not ( w_33800 , w_33801 );
and ( w_33801 , \13169_b1 , \13169_b0 );
or ( \13171_b1 , \13156_b1 , \13170_b1 );
xor ( \13171_b0 , \13156_b0 , w_33802 );
not ( w_33802 , w_33803 );
and ( w_33803 , \13170_b1 , \13170_b0 );
or ( \13172_b1 , \13137_b1 , \13171_b1 );
xor ( \13172_b0 , \13137_b0 , w_33804 );
not ( w_33804 , w_33805 );
and ( w_33805 , \13171_b1 , \13171_b0 );
or ( \13173_b1 , \7198_b1 , \13003_b1 );
not ( \13003_b1 , w_33806 );
and ( \13173_b0 , \7198_b0 , w_33807 );
and ( w_33806 , w_33807 , \13003_b0 );
or ( \13174_b1 , \13003_b1 , \13008_b1 );
not ( \13008_b1 , w_33808 );
and ( \13174_b0 , \13003_b0 , w_33809 );
and ( w_33808 , w_33809 , \13008_b0 );
or ( \13175_b1 , \7198_b1 , \13008_b1 );
not ( \13008_b1 , w_33810 );
and ( \13175_b0 , \7198_b0 , w_33811 );
and ( w_33810 , w_33811 , \13008_b0 );
or ( \13177_b1 , \12989_b1 , \12993_b1 );
not ( \12993_b1 , w_33812 );
and ( \13177_b0 , \12989_b0 , w_33813 );
and ( w_33812 , w_33813 , \12993_b0 );
or ( \13178_b1 , \12993_b1 , \12998_b1 );
not ( \12998_b1 , w_33814 );
and ( \13178_b0 , \12993_b0 , w_33815 );
and ( w_33814 , w_33815 , \12998_b0 );
or ( \13179_b1 , \12989_b1 , \12998_b1 );
not ( \12998_b1 , w_33816 );
and ( \13179_b0 , \12989_b0 , w_33817 );
and ( w_33816 , w_33817 , \12998_b0 );
or ( \13181_b1 , \13176_b1 , \13180_b1 );
xor ( \13181_b0 , \13176_b0 , w_33818 );
not ( w_33818 , w_33819 );
and ( w_33819 , \13180_b1 , \13180_b0 );
or ( \13182_b1 , \13031_b1 , \13035_b1 );
not ( \13035_b1 , w_33820 );
and ( \13182_b0 , \13031_b0 , w_33821 );
and ( w_33820 , w_33821 , \13035_b0 );
or ( \13183_b1 , \13035_b1 , \13040_b1 );
not ( \13040_b1 , w_33822 );
and ( \13183_b0 , \13035_b0 , w_33823 );
and ( w_33822 , w_33823 , \13040_b0 );
or ( \13184_b1 , \13031_b1 , \13040_b1 );
not ( \13040_b1 , w_33824 );
and ( \13184_b0 , \13031_b0 , w_33825 );
and ( w_33824 , w_33825 , \13040_b0 );
or ( \13186_b1 , \13181_b1 , \13185_b1 );
xor ( \13186_b0 , \13181_b0 , w_33826 );
not ( w_33826 , w_33827 );
and ( w_33827 , \13185_b1 , \13185_b0 );
or ( \13187_b1 , \13172_b1 , \13186_b1 );
xor ( \13187_b0 , \13172_b0 , w_33828 );
not ( w_33828 , w_33829 );
and ( w_33829 , \13186_b1 , \13186_b0 );
or ( \13188_b1 , \13108_b1 , \13187_b1 );
xor ( \13188_b0 , \13108_b0 , w_33830 );
not ( w_33830 , w_33831 );
and ( w_33831 , \13187_b1 , \13187_b0 );
or ( \13189_b1 , \13099_b1 , \13188_b1 );
xor ( \13189_b0 , \13099_b0 , w_33832 );
not ( w_33832 , w_33833 );
and ( w_33833 , \13188_b1 , \13188_b0 );
or ( \13190_b1 , \12979_b1 , \12980_b1 );
not ( \12980_b1 , w_33834 );
and ( \13190_b0 , \12979_b0 , w_33835 );
and ( w_33834 , w_33835 , \12980_b0 );
or ( \13191_b1 , \12980_b1 , \13074_b1 );
not ( \13074_b1 , w_33836 );
and ( \13191_b0 , \12980_b0 , w_33837 );
and ( w_33836 , w_33837 , \13074_b0 );
or ( \13192_b1 , \12979_b1 , \13074_b1 );
not ( \13074_b1 , w_33838 );
and ( \13192_b0 , \12979_b0 , w_33839 );
and ( w_33838 , w_33839 , \13074_b0 );
or ( \13194_b1 , \13189_b1 , w_33841 );
not ( w_33841 , w_33842 );
and ( \13194_b0 , \13189_b0 , w_33843 );
and ( w_33842 ,  , w_33843 );
buf ( w_33841 , \13193_b1 );
not ( w_33841 , w_33844 );
not (  , w_33845 );
and ( w_33844 , w_33845 , \13193_b0 );
or ( \13195_b1 , \13103_b1 , \13107_b1 );
not ( \13107_b1 , w_33846 );
and ( \13195_b0 , \13103_b0 , w_33847 );
and ( w_33846 , w_33847 , \13107_b0 );
or ( \13196_b1 , \13107_b1 , \13187_b1 );
not ( \13187_b1 , w_33848 );
and ( \13196_b0 , \13107_b0 , w_33849 );
and ( w_33848 , w_33849 , \13187_b0 );
or ( \13197_b1 , \13103_b1 , \13187_b1 );
not ( \13187_b1 , w_33850 );
and ( \13197_b0 , \13103_b0 , w_33851 );
and ( w_33850 , w_33851 , \13187_b0 );
or ( \13199_b1 , \13176_b1 , \13180_b1 );
not ( \13180_b1 , w_33852 );
and ( \13199_b0 , \13176_b0 , w_33853 );
and ( w_33852 , w_33853 , \13180_b0 );
or ( \13200_b1 , \13180_b1 , \13185_b1 );
not ( \13185_b1 , w_33854 );
and ( \13200_b0 , \13180_b0 , w_33855 );
and ( w_33854 , w_33855 , \13185_b0 );
or ( \13201_b1 , \13176_b1 , \13185_b1 );
not ( \13185_b1 , w_33856 );
and ( \13201_b0 , \13176_b0 , w_33857 );
and ( w_33856 , w_33857 , \13185_b0 );
or ( \13203_b1 , \13141_b1 , \13155_b1 );
not ( \13155_b1 , w_33858 );
and ( \13203_b0 , \13141_b0 , w_33859 );
and ( w_33858 , w_33859 , \13155_b0 );
or ( \13204_b1 , \13155_b1 , \13170_b1 );
not ( \13170_b1 , w_33860 );
and ( \13204_b0 , \13155_b0 , w_33861 );
and ( w_33860 , w_33861 , \13170_b0 );
or ( \13205_b1 , \13141_b1 , \13170_b1 );
not ( \13170_b1 , w_33862 );
and ( \13205_b0 , \13141_b0 , w_33863 );
and ( w_33862 , w_33863 , \13170_b0 );
or ( \13207_b1 , \13202_b1 , \13206_b1 );
xor ( \13207_b0 , \13202_b0 , w_33864 );
not ( w_33864 , w_33865 );
and ( w_33865 , \13206_b1 , \13206_b0 );
or ( \13208_b1 , \13122_b1 , \13136_b1 );
not ( \13136_b1 , w_33866 );
and ( \13208_b0 , \13122_b0 , w_33867 );
and ( w_33866 , w_33867 , \13136_b0 );
or ( \13209_b1 , \13207_b1 , \13208_b1 );
xor ( \13209_b0 , \13207_b0 , w_33868 );
not ( w_33868 , w_33869 );
and ( w_33869 , \13208_b1 , \13208_b0 );
or ( \13210_b1 , \13198_b1 , \13209_b1 );
xor ( \13210_b0 , \13198_b0 , w_33870 );
not ( w_33870 , w_33871 );
and ( w_33871 , \13209_b1 , \13209_b0 );
or ( \13211_b1 , \13091_b1 , \13095_b1 );
not ( \13095_b1 , w_33872 );
and ( \13211_b0 , \13091_b0 , w_33873 );
and ( w_33872 , w_33873 , \13095_b0 );
or ( \13212_b1 , \13095_b1 , \13097_b1 );
not ( \13097_b1 , w_33874 );
and ( \13212_b0 , \13095_b0 , w_33875 );
and ( w_33874 , w_33875 , \13097_b0 );
or ( \13213_b1 , \13091_b1 , \13097_b1 );
not ( \13097_b1 , w_33876 );
and ( \13213_b0 , \13091_b0 , w_33877 );
and ( w_33876 , w_33877 , \13097_b0 );
or ( \13215_b1 , \13137_b1 , \13171_b1 );
not ( \13171_b1 , w_33878 );
and ( \13215_b0 , \13137_b0 , w_33879 );
and ( w_33878 , w_33879 , \13171_b0 );
or ( \13216_b1 , \13171_b1 , \13186_b1 );
not ( \13186_b1 , w_33880 );
and ( \13216_b0 , \13171_b0 , w_33881 );
and ( w_33880 , w_33881 , \13186_b0 );
or ( \13217_b1 , \13137_b1 , \13186_b1 );
not ( \13186_b1 , w_33882 );
and ( \13217_b0 , \13137_b0 , w_33883 );
and ( w_33882 , w_33883 , \13186_b0 );
or ( \13219_b1 , \13214_b1 , \13218_b1 );
xor ( \13219_b0 , \13214_b0 , w_33884 );
not ( w_33884 , w_33885 );
and ( w_33885 , \13218_b1 , \13218_b0 );
or ( \13220_b1 , \5925_b1 , \7082_b1 );
not ( \7082_b1 , w_33886 );
and ( \13220_b0 , \5925_b0 , w_33887 );
and ( w_33886 , w_33887 , \7082_b0 );
or ( \13221_b1 , \5937_b1 , \7080_b1 );
not ( \7080_b1 , w_33888 );
and ( \13221_b0 , \5937_b0 , w_33889 );
and ( w_33888 , w_33889 , \7080_b0 );
or ( \13222_b1 , \13220_b1 , w_33891 );
not ( w_33891 , w_33892 );
and ( \13222_b0 , \13220_b0 , w_33893 );
and ( w_33892 ,  , w_33893 );
buf ( w_33891 , \13221_b1 );
not ( w_33891 , w_33894 );
not (  , w_33895 );
and ( w_33894 , w_33895 , \13221_b0 );
or ( \13223_b1 , \13222_b1 , w_33896 );
xor ( \13223_b0 , \13222_b0 , w_33898 );
not ( w_33898 , w_33899 );
and ( w_33899 , w_33896 , w_33897 );
buf ( w_33896 , \7088_b1 );
not ( w_33896 , w_33900 );
not ( w_33897 , w_33901 );
and ( w_33900 , w_33901 , \7088_b0 );
or ( \13224_b1 , \5945_b1 , \7099_b1 );
not ( \7099_b1 , w_33902 );
and ( \13224_b0 , \5945_b0 , w_33903 );
and ( w_33902 , w_33903 , \7099_b0 );
or ( \13225_b1 , \5957_b1 , \7097_b1 );
not ( \7097_b1 , w_33904 );
and ( \13225_b0 , \5957_b0 , w_33905 );
and ( w_33904 , w_33905 , \7097_b0 );
or ( \13226_b1 , \13224_b1 , w_33907 );
not ( w_33907 , w_33908 );
and ( \13226_b0 , \13224_b0 , w_33909 );
and ( w_33908 ,  , w_33909 );
buf ( w_33907 , \13225_b1 );
not ( w_33907 , w_33910 );
not (  , w_33911 );
and ( w_33910 , w_33911 , \13225_b0 );
or ( \13227_b1 , \13226_b1 , w_33912 );
xor ( \13227_b0 , \13226_b0 , w_33914 );
not ( w_33914 , w_33915 );
and ( w_33915 , w_33912 , w_33913 );
buf ( w_33912 , \7105_b1 );
not ( w_33912 , w_33916 );
not ( w_33913 , w_33917 );
and ( w_33916 , w_33917 , \7105_b0 );
or ( \13228_b1 , \13223_b1 , \13227_b1 );
xor ( \13228_b0 , \13223_b0 , w_33918 );
not ( w_33918 , w_33919 );
and ( w_33919 , \13227_b1 , \13227_b0 );
or ( \13229_b1 , \5967_b1 , \7117_b1 );
not ( \7117_b1 , w_33920 );
and ( \13229_b0 , \5967_b0 , w_33921 );
and ( w_33920 , w_33921 , \7117_b0 );
or ( \13230_b1 , \5979_b1 , \7115_b1 );
not ( \7115_b1 , w_33922 );
and ( \13230_b0 , \5979_b0 , w_33923 );
and ( w_33922 , w_33923 , \7115_b0 );
or ( \13231_b1 , \13229_b1 , w_33925 );
not ( w_33925 , w_33926 );
and ( \13231_b0 , \13229_b0 , w_33927 );
and ( w_33926 ,  , w_33927 );
buf ( w_33925 , \13230_b1 );
not ( w_33925 , w_33928 );
not (  , w_33929 );
and ( w_33928 , w_33929 , \13230_b0 );
or ( \13232_b1 , \13231_b1 , w_33930 );
xor ( \13232_b0 , \13231_b0 , w_33932 );
not ( w_33932 , w_33933 );
and ( w_33933 , w_33930 , w_33931 );
buf ( w_33930 , \7123_b1 );
not ( w_33930 , w_33934 );
not ( w_33931 , w_33935 );
and ( w_33934 , w_33935 , \7123_b0 );
or ( \13233_b1 , \13228_b1 , \13232_b1 );
xor ( \13233_b0 , \13228_b0 , w_33936 );
not ( w_33936 , w_33937 );
and ( w_33937 , \13232_b1 , \13232_b0 );
or ( \13234_b1 , \5861_b1 , \7026_b1 );
not ( \7026_b1 , w_33938 );
and ( \13234_b0 , \5861_b0 , w_33939 );
and ( w_33938 , w_33939 , \7026_b0 );
or ( \13235_b1 , \5873_b1 , \7024_b1 );
not ( \7024_b1 , w_33940 );
and ( \13235_b0 , \5873_b0 , w_33941 );
and ( w_33940 , w_33941 , \7024_b0 );
or ( \13236_b1 , \13234_b1 , w_33943 );
not ( w_33943 , w_33944 );
and ( \13236_b0 , \13234_b0 , w_33945 );
and ( w_33944 ,  , w_33945 );
buf ( w_33943 , \13235_b1 );
not ( w_33943 , w_33946 );
not (  , w_33947 );
and ( w_33946 , w_33947 , \13235_b0 );
or ( \13237_b1 , \13236_b1 , w_33948 );
xor ( \13237_b0 , \13236_b0 , w_33950 );
not ( w_33950 , w_33951 );
and ( w_33951 , w_33948 , w_33949 );
buf ( w_33948 , \7032_b1 );
not ( w_33948 , w_33952 );
not ( w_33949 , w_33953 );
and ( w_33952 , w_33953 , \7032_b0 );
or ( \13238_b1 , \5881_b1 , \7043_b1 );
not ( \7043_b1 , w_33954 );
and ( \13238_b0 , \5881_b0 , w_33955 );
and ( w_33954 , w_33955 , \7043_b0 );
or ( \13239_b1 , \5893_b1 , \7041_b1 );
not ( \7041_b1 , w_33956 );
and ( \13239_b0 , \5893_b0 , w_33957 );
and ( w_33956 , w_33957 , \7041_b0 );
or ( \13240_b1 , \13238_b1 , w_33959 );
not ( w_33959 , w_33960 );
and ( \13240_b0 , \13238_b0 , w_33961 );
and ( w_33960 ,  , w_33961 );
buf ( w_33959 , \13239_b1 );
not ( w_33959 , w_33962 );
not (  , w_33963 );
and ( w_33962 , w_33963 , \13239_b0 );
or ( \13241_b1 , \13240_b1 , w_33964 );
xor ( \13241_b0 , \13240_b0 , w_33966 );
not ( w_33966 , w_33967 );
and ( w_33967 , w_33964 , w_33965 );
buf ( w_33964 , \7049_b1 );
not ( w_33964 , w_33968 );
not ( w_33965 , w_33969 );
and ( w_33968 , w_33969 , \7049_b0 );
or ( \13242_b1 , \13237_b1 , \13241_b1 );
xor ( \13242_b0 , \13237_b0 , w_33970 );
not ( w_33970 , w_33971 );
and ( w_33971 , \13241_b1 , \13241_b0 );
or ( \13243_b1 , \5906_b1 , \7061_b1 );
not ( \7061_b1 , w_33972 );
and ( \13243_b0 , \5906_b0 , w_33973 );
and ( w_33972 , w_33973 , \7061_b0 );
or ( \13244_b1 , \5918_b1 , \7059_b1 );
not ( \7059_b1 , w_33974 );
and ( \13244_b0 , \5918_b0 , w_33975 );
and ( w_33974 , w_33975 , \7059_b0 );
or ( \13245_b1 , \13243_b1 , w_33977 );
not ( w_33977 , w_33978 );
and ( \13245_b0 , \13243_b0 , w_33979 );
and ( w_33978 ,  , w_33979 );
buf ( w_33977 , \13244_b1 );
not ( w_33977 , w_33980 );
not (  , w_33981 );
and ( w_33980 , w_33981 , \13244_b0 );
or ( \13246_b1 , \13245_b1 , w_33982 );
xor ( \13246_b0 , \13245_b0 , w_33984 );
not ( w_33984 , w_33985 );
and ( w_33985 , w_33982 , w_33983 );
buf ( w_33982 , \7067_b1 );
not ( w_33982 , w_33986 );
not ( w_33983 , w_33987 );
and ( w_33986 , w_33987 , \7067_b0 );
or ( \13247_b1 , \13242_b1 , \13246_b1 );
xor ( \13247_b0 , \13242_b0 , w_33988 );
not ( w_33988 , w_33989 );
and ( w_33989 , \13246_b1 , \13246_b0 );
or ( \13248_b1 , \13233_b1 , \13247_b1 );
xor ( \13248_b0 , \13233_b0 , w_33990 );
not ( w_33990 , w_33991 );
and ( w_33991 , \13247_b1 , \13247_b0 );
or ( \13249_b1 , \5819_b1 , \6991_b1 );
not ( \6991_b1 , w_33992 );
and ( \13249_b0 , \5819_b0 , w_33993 );
and ( w_33992 , w_33993 , \6991_b0 );
or ( \13250_b1 , \5831_b1 , \6988_b1 );
not ( \6988_b1 , w_33994 );
and ( \13250_b0 , \5831_b0 , w_33995 );
and ( w_33994 , w_33995 , \6988_b0 );
or ( \13251_b1 , \13249_b1 , w_33997 );
not ( w_33997 , w_33998 );
and ( \13251_b0 , \13249_b0 , w_33999 );
and ( w_33998 ,  , w_33999 );
buf ( w_33997 , \13250_b1 );
not ( w_33997 , w_34000 );
not (  , w_34001 );
and ( w_34000 , w_34001 , \13250_b0 );
or ( \13252_b1 , \13251_b1 , w_34002 );
xor ( \13252_b0 , \13251_b0 , w_34004 );
not ( w_34004 , w_34005 );
and ( w_34005 , w_34002 , w_34003 );
buf ( w_34002 , \6985_b1 );
not ( w_34002 , w_34006 );
not ( w_34003 , w_34007 );
and ( w_34006 , w_34007 , \6985_b0 );
or ( \13253_b1 , \6824_b1 , \13252_b1 );
xor ( \13253_b0 , \6824_b0 , w_34008 );
not ( w_34008 , w_34009 );
and ( w_34009 , \13252_b1 , \13252_b0 );
or ( \13254_b1 , \5842_b1 , \7006_b1 );
not ( \7006_b1 , w_34010 );
and ( \13254_b0 , \5842_b0 , w_34011 );
and ( w_34010 , w_34011 , \7006_b0 );
or ( \13255_b1 , \5854_b1 , \7004_b1 );
not ( \7004_b1 , w_34012 );
and ( \13255_b0 , \5854_b0 , w_34013 );
and ( w_34012 , w_34013 , \7004_b0 );
or ( \13256_b1 , \13254_b1 , w_34015 );
not ( w_34015 , w_34016 );
and ( \13256_b0 , \13254_b0 , w_34017 );
and ( w_34016 ,  , w_34017 );
buf ( w_34015 , \13255_b1 );
not ( w_34015 , w_34018 );
not (  , w_34019 );
and ( w_34018 , w_34019 , \13255_b0 );
or ( \13257_b1 , \13256_b1 , w_34020 );
xor ( \13257_b0 , \13256_b0 , w_34022 );
not ( w_34022 , w_34023 );
and ( w_34023 , w_34020 , w_34021 );
buf ( w_34020 , \7012_b1 );
not ( w_34020 , w_34024 );
not ( w_34021 , w_34025 );
and ( w_34024 , w_34025 , \7012_b0 );
or ( \13258_b1 , \13253_b1 , \13257_b1 );
xor ( \13258_b0 , \13253_b0 , w_34026 );
not ( w_34026 , w_34027 );
and ( w_34027 , \13257_b1 , \13257_b0 );
or ( \13259_b1 , \13248_b1 , \13258_b1 );
xor ( \13259_b0 , \13248_b0 , w_34028 );
not ( w_34028 , w_34029 );
and ( w_34029 , \13258_b1 , \13258_b0 );
or ( \13260_b1 , \13145_b1 , \13149_b1 );
not ( \13149_b1 , w_34030 );
and ( \13260_b0 , \13145_b0 , w_34031 );
and ( w_34030 , w_34031 , \13149_b0 );
or ( \13261_b1 , \13149_b1 , \13154_b1 );
not ( \13154_b1 , w_34032 );
and ( \13261_b0 , \13149_b0 , w_34033 );
and ( w_34032 , w_34033 , \13154_b0 );
or ( \13262_b1 , \13145_b1 , \13154_b1 );
not ( \13154_b1 , w_34034 );
and ( \13262_b0 , \13145_b0 , w_34035 );
and ( w_34034 , w_34035 , \13154_b0 );
or ( \13264_b1 , \6048_b1 , \7192_b1 );
not ( \7192_b1 , w_34036 );
and ( \13264_b0 , \6048_b0 , w_34037 );
and ( w_34036 , w_34037 , \7192_b0 );
or ( \13265_b1 , \6057_b1 , \7190_b1 );
not ( \7190_b1 , w_34038 );
and ( \13265_b0 , \6057_b0 , w_34039 );
and ( w_34038 , w_34039 , \7190_b0 );
or ( \13266_b1 , \13264_b1 , w_34041 );
not ( w_34041 , w_34042 );
and ( \13266_b0 , \13264_b0 , w_34043 );
and ( w_34042 ,  , w_34043 );
buf ( w_34041 , \13265_b1 );
not ( w_34041 , w_34044 );
not (  , w_34045 );
and ( w_34044 , w_34045 , \13265_b0 );
or ( \13267_b1 , \13266_b1 , w_34046 );
xor ( \13267_b0 , \13266_b0 , w_34048 );
not ( w_34048 , w_34049 );
and ( w_34049 , w_34046 , w_34047 );
buf ( w_34046 , \7198_b1 );
not ( w_34046 , w_34050 );
not ( w_34047 , w_34051 );
and ( w_34050 , w_34051 , \7198_b0 );
or ( \13268_b1 , \6065_b1 , w_34053 );
not ( w_34053 , w_34054 );
and ( \13268_b0 , \6065_b0 , w_34055 );
and ( w_34054 ,  , w_34055 );
buf ( w_34053 , \7201_b1 );
not ( w_34053 , w_34056 );
not (  , w_34057 );
and ( w_34056 , w_34057 , \7201_b0 );
or ( \13269_b1 , \13268_b1 , w_34058 );
xor ( \13269_b0 , \13268_b0 , w_34060 );
not ( w_34060 , w_34061 );
and ( w_34061 , w_34058 , w_34059 );
buf ( w_34058 , \6824_b1 );
not ( w_34058 , w_34062 );
not ( w_34059 , w_34063 );
and ( w_34062 , w_34063 , \6824_b0 );
or ( \13270_b1 , \13267_b1 , \13269_b1 );
xor ( \13270_b0 , \13267_b0 , w_34064 );
not ( w_34064 , w_34065 );
and ( w_34065 , \13269_b1 , \13269_b0 );
or ( \13271_b1 , \13263_b1 , \13270_b1 );
xor ( \13271_b0 , \13263_b0 , w_34066 );
not ( w_34066 , w_34067 );
and ( w_34067 , \13270_b1 , \13270_b0 );
or ( \13272_b1 , \5986_b1 , \7140_b1 );
not ( \7140_b1 , w_34068 );
and ( \13272_b0 , \5986_b0 , w_34069 );
and ( w_34068 , w_34069 , \7140_b0 );
or ( \13273_b1 , \5998_b1 , \7138_b1 );
not ( \7138_b1 , w_34070 );
and ( \13273_b0 , \5998_b0 , w_34071 );
and ( w_34070 , w_34071 , \7138_b0 );
or ( \13274_b1 , \13272_b1 , w_34073 );
not ( w_34073 , w_34074 );
and ( \13274_b0 , \13272_b0 , w_34075 );
and ( w_34074 ,  , w_34075 );
buf ( w_34073 , \13273_b1 );
not ( w_34073 , w_34076 );
not (  , w_34077 );
and ( w_34076 , w_34077 , \13273_b0 );
or ( \13275_b1 , \13274_b1 , w_34078 );
xor ( \13275_b0 , \13274_b0 , w_34080 );
not ( w_34080 , w_34081 );
and ( w_34081 , w_34078 , w_34079 );
buf ( w_34078 , \7146_b1 );
not ( w_34078 , w_34082 );
not ( w_34079 , w_34083 );
and ( w_34082 , w_34083 , \7146_b0 );
or ( \13276_b1 , \6006_b1 , \7157_b1 );
not ( \7157_b1 , w_34084 );
and ( \13276_b0 , \6006_b0 , w_34085 );
and ( w_34084 , w_34085 , \7157_b0 );
or ( \13277_b1 , \6018_b1 , \7155_b1 );
not ( \7155_b1 , w_34086 );
and ( \13277_b0 , \6018_b0 , w_34087 );
and ( w_34086 , w_34087 , \7155_b0 );
or ( \13278_b1 , \13276_b1 , w_34089 );
not ( w_34089 , w_34090 );
and ( \13278_b0 , \13276_b0 , w_34091 );
and ( w_34090 ,  , w_34091 );
buf ( w_34089 , \13277_b1 );
not ( w_34089 , w_34092 );
not (  , w_34093 );
and ( w_34092 , w_34093 , \13277_b0 );
or ( \13279_b1 , \13278_b1 , w_34094 );
xor ( \13279_b0 , \13278_b0 , w_34096 );
not ( w_34096 , w_34097 );
and ( w_34097 , w_34094 , w_34095 );
buf ( w_34094 , \7163_b1 );
not ( w_34094 , w_34098 );
not ( w_34095 , w_34099 );
and ( w_34098 , w_34099 , \7163_b0 );
or ( \13280_b1 , \13275_b1 , \13279_b1 );
xor ( \13280_b0 , \13275_b0 , w_34100 );
not ( w_34100 , w_34101 );
and ( w_34101 , \13279_b1 , \13279_b0 );
or ( \13281_b1 , \6029_b1 , \7175_b1 );
not ( \7175_b1 , w_34102 );
and ( \13281_b0 , \6029_b0 , w_34103 );
and ( w_34102 , w_34103 , \7175_b0 );
or ( \13282_b1 , \6041_b1 , \7173_b1 );
not ( \7173_b1 , w_34104 );
and ( \13282_b0 , \6041_b0 , w_34105 );
and ( w_34104 , w_34105 , \7173_b0 );
or ( \13283_b1 , \13281_b1 , w_34107 );
not ( w_34107 , w_34108 );
and ( \13283_b0 , \13281_b0 , w_34109 );
and ( w_34108 ,  , w_34109 );
buf ( w_34107 , \13282_b1 );
not ( w_34107 , w_34110 );
not (  , w_34111 );
and ( w_34110 , w_34111 , \13282_b0 );
or ( \13284_b1 , \13283_b1 , w_34112 );
xor ( \13284_b0 , \13283_b0 , w_34114 );
not ( w_34114 , w_34115 );
and ( w_34115 , w_34112 , w_34113 );
buf ( w_34112 , \7181_b1 );
not ( w_34112 , w_34116 );
not ( w_34113 , w_34117 );
and ( w_34116 , w_34117 , \7181_b0 );
or ( \13285_b1 , \13280_b1 , \13284_b1 );
xor ( \13285_b0 , \13280_b0 , w_34118 );
not ( w_34118 , w_34119 );
and ( w_34119 , \13284_b1 , \13284_b0 );
or ( \13286_b1 , \13271_b1 , \13285_b1 );
xor ( \13286_b0 , \13271_b0 , w_34120 );
not ( w_34120 , w_34121 );
and ( w_34121 , \13285_b1 , \13285_b0 );
or ( \13287_b1 , \13259_b1 , \13286_b1 );
xor ( \13287_b0 , \13259_b0 , w_34122 );
not ( w_34122 , w_34123 );
and ( w_34123 , \13286_b1 , \13286_b0 );
or ( \13288_b1 , \13126_b1 , \13130_b1 );
not ( \13130_b1 , w_34124 );
and ( \13288_b0 , \13126_b0 , w_34125 );
and ( w_34124 , w_34125 , \13130_b0 );
or ( \13289_b1 , \13130_b1 , \13135_b1 );
not ( \13135_b1 , w_34126 );
and ( \13289_b0 , \13130_b0 , w_34127 );
and ( w_34126 , w_34127 , \13135_b0 );
or ( \13290_b1 , \13126_b1 , \13135_b1 );
not ( \13135_b1 , w_34128 );
and ( \13290_b0 , \13126_b0 , w_34129 );
and ( w_34128 , w_34129 , \13135_b0 );
or ( \13292_b1 , \13112_b1 , \13116_b1 );
not ( \13116_b1 , w_34130 );
and ( \13292_b0 , \13112_b0 , w_34131 );
and ( w_34130 , w_34131 , \13116_b0 );
or ( \13293_b1 , \13116_b1 , \13121_b1 );
not ( \13121_b1 , w_34132 );
and ( \13293_b0 , \13116_b0 , w_34133 );
and ( w_34132 , w_34133 , \13121_b0 );
or ( \13294_b1 , \13112_b1 , \13121_b1 );
not ( \13121_b1 , w_34134 );
and ( \13294_b0 , \13112_b0 , w_34135 );
and ( w_34134 , w_34135 , \13121_b0 );
or ( \13296_b1 , \13291_b1 , \13295_b1 );
xor ( \13296_b0 , \13291_b0 , w_34136 );
not ( w_34136 , w_34137 );
and ( w_34137 , \13295_b1 , \13295_b0 );
or ( \13297_b1 , \13160_b1 , \13164_b1 );
not ( \13164_b1 , w_34138 );
and ( \13297_b0 , \13160_b0 , w_34139 );
and ( w_34138 , w_34139 , \13164_b0 );
or ( \13298_b1 , \13164_b1 , \13169_b1 );
not ( \13169_b1 , w_34140 );
and ( \13298_b0 , \13164_b0 , w_34141 );
and ( w_34140 , w_34141 , \13169_b0 );
or ( \13299_b1 , \13160_b1 , \13169_b1 );
not ( \13169_b1 , w_34142 );
and ( \13299_b0 , \13160_b0 , w_34143 );
and ( w_34142 , w_34143 , \13169_b0 );
or ( \13301_b1 , \13296_b1 , \13300_b1 );
xor ( \13301_b0 , \13296_b0 , w_34144 );
not ( w_34144 , w_34145 );
and ( w_34145 , \13300_b1 , \13300_b0 );
or ( \13302_b1 , \13287_b1 , \13301_b1 );
xor ( \13302_b0 , \13287_b0 , w_34146 );
not ( w_34146 , w_34147 );
and ( w_34147 , \13301_b1 , \13301_b0 );
or ( \13303_b1 , \13219_b1 , \13302_b1 );
xor ( \13303_b0 , \13219_b0 , w_34148 );
not ( w_34148 , w_34149 );
and ( w_34149 , \13302_b1 , \13302_b0 );
or ( \13304_b1 , \13210_b1 , \13303_b1 );
xor ( \13304_b0 , \13210_b0 , w_34150 );
not ( w_34150 , w_34151 );
and ( w_34151 , \13303_b1 , \13303_b0 );
or ( \13305_b1 , \13087_b1 , \13098_b1 );
not ( \13098_b1 , w_34152 );
and ( \13305_b0 , \13087_b0 , w_34153 );
and ( w_34152 , w_34153 , \13098_b0 );
or ( \13306_b1 , \13098_b1 , \13188_b1 );
not ( \13188_b1 , w_34154 );
and ( \13306_b0 , \13098_b0 , w_34155 );
and ( w_34154 , w_34155 , \13188_b0 );
or ( \13307_b1 , \13087_b1 , \13188_b1 );
not ( \13188_b1 , w_34156 );
and ( \13307_b0 , \13087_b0 , w_34157 );
and ( w_34156 , w_34157 , \13188_b0 );
or ( \13309_b1 , \13304_b1 , w_34159 );
not ( w_34159 , w_34160 );
and ( \13309_b0 , \13304_b0 , w_34161 );
and ( w_34160 ,  , w_34161 );
buf ( w_34159 , \13308_b1 );
not ( w_34159 , w_34162 );
not (  , w_34163 );
and ( w_34162 , w_34163 , \13308_b0 );
or ( \13310_b1 , \13194_b1 , w_34165 );
not ( w_34165 , w_34166 );
and ( \13310_b0 , \13194_b0 , w_34167 );
and ( w_34166 ,  , w_34167 );
buf ( w_34165 , \13309_b1 );
not ( w_34165 , w_34168 );
not (  , w_34169 );
and ( w_34168 , w_34169 , \13309_b0 );
or ( \13311_b1 , \13214_b1 , \13218_b1 );
not ( \13218_b1 , w_34170 );
and ( \13311_b0 , \13214_b0 , w_34171 );
and ( w_34170 , w_34171 , \13218_b0 );
or ( \13312_b1 , \13218_b1 , \13302_b1 );
not ( \13302_b1 , w_34172 );
and ( \13312_b0 , \13218_b0 , w_34173 );
and ( w_34172 , w_34173 , \13302_b0 );
or ( \13313_b1 , \13214_b1 , \13302_b1 );
not ( \13302_b1 , w_34174 );
and ( \13313_b0 , \13214_b0 , w_34175 );
and ( w_34174 , w_34175 , \13302_b0 );
or ( \13315_b1 , \7770_b1 , \7774_b1 );
xor ( \13315_b0 , \7770_b0 , w_34176 );
not ( w_34176 , w_34177 );
and ( w_34177 , \7774_b1 , \7774_b0 );
or ( \13316_b1 , \13315_b1 , \7779_b1 );
xor ( \13316_b0 , \13315_b0 , w_34178 );
not ( w_34178 , w_34179 );
and ( w_34179 , \7779_b1 , \7779_b0 );
or ( \13317_b1 , \7822_b1 , \7826_b1 );
xor ( \13317_b0 , \7822_b0 , w_34180 );
not ( w_34180 , w_34181 );
and ( w_34181 , \7826_b1 , \7826_b0 );
or ( \13318_b1 , \13317_b1 , \7831_b1 );
xor ( \13318_b0 , \13317_b0 , w_34182 );
not ( w_34182 , w_34183 );
and ( w_34183 , \7831_b1 , \7831_b0 );
or ( \13319_b1 , \7803_b1 , \7807_b1 );
xor ( \13319_b0 , \7803_b0 , w_34184 );
not ( w_34184 , w_34185 );
and ( w_34185 , \7807_b1 , \7807_b0 );
or ( \13320_b1 , \13319_b1 , \7812_b1 );
xor ( \13320_b0 , \13319_b0 , w_34186 );
not ( w_34186 , w_34187 );
and ( w_34187 , \7812_b1 , \7812_b0 );
or ( \13321_b1 , \13318_b1 , \13320_b1 );
xor ( \13321_b0 , \13318_b0 , w_34188 );
not ( w_34188 , w_34189 );
and ( w_34189 , \13320_b1 , \13320_b0 );
or ( \13322_b1 , \7786_b1 , \7790_b1 );
xor ( \13322_b0 , \7786_b0 , w_34190 );
not ( w_34190 , w_34191 );
and ( w_34191 , \7790_b1 , \7790_b0 );
or ( \13323_b1 , \13322_b1 , \7795_b1 );
xor ( \13323_b0 , \13322_b0 , w_34192 );
not ( w_34192 , w_34193 );
and ( w_34193 , \7795_b1 , \7795_b0 );
or ( \13324_b1 , \13321_b1 , \13323_b1 );
xor ( \13324_b0 , \13321_b0 , w_34194 );
not ( w_34194 , w_34195 );
and ( w_34195 , \13323_b1 , \13323_b0 );
or ( \13325_b1 , \13316_b1 , \13324_b1 );
xor ( \13325_b0 , \13316_b0 , w_34196 );
not ( w_34196 , w_34197 );
and ( w_34197 , \13324_b1 , \13324_b0 );
or ( \13326_b1 , \13275_b1 , \13279_b1 );
not ( \13279_b1 , w_34198 );
and ( \13326_b0 , \13275_b0 , w_34199 );
and ( w_34198 , w_34199 , \13279_b0 );
or ( \13327_b1 , \13279_b1 , \13284_b1 );
not ( \13284_b1 , w_34200 );
and ( \13327_b0 , \13279_b0 , w_34201 );
and ( w_34200 , w_34201 , \13284_b0 );
or ( \13328_b1 , \13275_b1 , \13284_b1 );
not ( \13284_b1 , w_34202 );
and ( \13328_b0 , \13275_b0 , w_34203 );
and ( w_34202 , w_34203 , \13284_b0 );
or ( \13330_b1 , \13267_b1 , \13269_b1 );
not ( \13269_b1 , w_34204 );
and ( \13330_b0 , \13267_b0 , w_34205 );
and ( w_34204 , w_34205 , \13269_b0 );
or ( \13331_b1 , \13329_b1 , \13330_b1 );
xor ( \13331_b0 , \13329_b0 , w_34206 );
not ( w_34206 , w_34207 );
and ( w_34207 , \13330_b1 , \13330_b0 );
or ( \13332_b1 , \6065_b1 , \7203_b1 );
not ( \7203_b1 , w_34208 );
and ( \13332_b0 , \6065_b0 , w_34209 );
and ( w_34208 , w_34209 , \7203_b0 );
or ( \13333_b1 , \6048_b1 , \7201_b1 );
not ( \7201_b1 , w_34210 );
and ( \13333_b0 , \6048_b0 , w_34211 );
and ( w_34210 , w_34211 , \7201_b0 );
or ( \13334_b1 , \13332_b1 , w_34213 );
not ( w_34213 , w_34214 );
and ( \13334_b0 , \13332_b0 , w_34215 );
and ( w_34214 ,  , w_34215 );
buf ( w_34213 , \13333_b1 );
not ( w_34213 , w_34216 );
not (  , w_34217 );
and ( w_34216 , w_34217 , \13333_b0 );
or ( \13335_b1 , \13334_b1 , w_34218 );
xor ( \13335_b0 , \13334_b0 , w_34220 );
not ( w_34220 , w_34221 );
and ( w_34221 , w_34218 , w_34219 );
buf ( w_34218 , \6824_b1 );
not ( w_34218 , w_34222 );
not ( w_34219 , w_34223 );
and ( w_34222 , w_34223 , \6824_b0 );
or ( \13336_b1 , \13331_b1 , \13335_b1 );
xor ( \13336_b0 , \13331_b0 , w_34224 );
not ( w_34224 , w_34225 );
and ( w_34225 , \13335_b1 , \13335_b0 );
or ( \13337_b1 , \13325_b1 , \13336_b1 );
xor ( \13337_b0 , \13325_b0 , w_34226 );
not ( w_34226 , w_34227 );
and ( w_34227 , \13336_b1 , \13336_b0 );
or ( \13338_b1 , \13291_b1 , \13295_b1 );
not ( \13295_b1 , w_34228 );
and ( \13338_b0 , \13291_b0 , w_34229 );
and ( w_34228 , w_34229 , \13295_b0 );
or ( \13339_b1 , \13295_b1 , \13300_b1 );
not ( \13300_b1 , w_34230 );
and ( \13339_b0 , \13295_b0 , w_34231 );
and ( w_34230 , w_34231 , \13300_b0 );
or ( \13340_b1 , \13291_b1 , \13300_b1 );
not ( \13300_b1 , w_34232 );
and ( \13340_b0 , \13291_b0 , w_34233 );
and ( w_34232 , w_34233 , \13300_b0 );
or ( \13342_b1 , \13263_b1 , \13270_b1 );
not ( \13270_b1 , w_34234 );
and ( \13342_b0 , \13263_b0 , w_34235 );
and ( w_34234 , w_34235 , \13270_b0 );
or ( \13343_b1 , \13270_b1 , \13285_b1 );
not ( \13285_b1 , w_34236 );
and ( \13343_b0 , \13270_b0 , w_34237 );
and ( w_34236 , w_34237 , \13285_b0 );
or ( \13344_b1 , \13263_b1 , \13285_b1 );
not ( \13285_b1 , w_34238 );
and ( \13344_b0 , \13263_b0 , w_34239 );
and ( w_34238 , w_34239 , \13285_b0 );
or ( \13346_b1 , \13341_b1 , \13345_b1 );
xor ( \13346_b0 , \13341_b0 , w_34240 );
not ( w_34240 , w_34241 );
and ( w_34241 , \13345_b1 , \13345_b0 );
or ( \13347_b1 , \13233_b1 , \13247_b1 );
not ( \13247_b1 , w_34242 );
and ( \13347_b0 , \13233_b0 , w_34243 );
and ( w_34242 , w_34243 , \13247_b0 );
or ( \13348_b1 , \13247_b1 , \13258_b1 );
not ( \13258_b1 , w_34244 );
and ( \13348_b0 , \13247_b0 , w_34245 );
and ( w_34244 , w_34245 , \13258_b0 );
or ( \13349_b1 , \13233_b1 , \13258_b1 );
not ( \13258_b1 , w_34246 );
and ( \13349_b0 , \13233_b0 , w_34247 );
and ( w_34246 , w_34247 , \13258_b0 );
or ( \13351_b1 , \13346_b1 , \13350_b1 );
xor ( \13351_b0 , \13346_b0 , w_34248 );
not ( w_34248 , w_34249 );
and ( w_34249 , \13350_b1 , \13350_b0 );
or ( \13352_b1 , \13337_b1 , \13351_b1 );
xor ( \13352_b0 , \13337_b0 , w_34250 );
not ( w_34250 , w_34251 );
and ( w_34251 , \13351_b1 , \13351_b0 );
or ( \13353_b1 , \13314_b1 , \13352_b1 );
xor ( \13353_b0 , \13314_b0 , w_34252 );
not ( w_34252 , w_34253 );
and ( w_34253 , \13352_b1 , \13352_b0 );
or ( \13354_b1 , \13202_b1 , \13206_b1 );
not ( \13206_b1 , w_34254 );
and ( \13354_b0 , \13202_b0 , w_34255 );
and ( w_34254 , w_34255 , \13206_b0 );
or ( \13355_b1 , \13206_b1 , \13208_b1 );
not ( \13208_b1 , w_34256 );
and ( \13355_b0 , \13206_b0 , w_34257 );
and ( w_34256 , w_34257 , \13208_b0 );
or ( \13356_b1 , \13202_b1 , \13208_b1 );
not ( \13208_b1 , w_34258 );
and ( \13356_b0 , \13202_b0 , w_34259 );
and ( w_34258 , w_34259 , \13208_b0 );
or ( \13358_b1 , \13259_b1 , \13286_b1 );
not ( \13286_b1 , w_34260 );
and ( \13358_b0 , \13259_b0 , w_34261 );
and ( w_34260 , w_34261 , \13286_b0 );
or ( \13359_b1 , \13286_b1 , \13301_b1 );
not ( \13301_b1 , w_34262 );
and ( \13359_b0 , \13286_b0 , w_34263 );
and ( w_34262 , w_34263 , \13301_b0 );
or ( \13360_b1 , \13259_b1 , \13301_b1 );
not ( \13301_b1 , w_34264 );
and ( \13360_b0 , \13259_b0 , w_34265 );
and ( w_34264 , w_34265 , \13301_b0 );
or ( \13362_b1 , \13357_b1 , \13361_b1 );
xor ( \13362_b0 , \13357_b0 , w_34266 );
not ( w_34266 , w_34267 );
and ( w_34267 , \13361_b1 , \13361_b0 );
or ( \13363_b1 , \6824_b1 , \13252_b1 );
not ( \13252_b1 , w_34268 );
and ( \13363_b0 , \6824_b0 , w_34269 );
and ( w_34268 , w_34269 , \13252_b0 );
or ( \13364_b1 , \13252_b1 , \13257_b1 );
not ( \13257_b1 , w_34270 );
and ( \13364_b0 , \13252_b0 , w_34271 );
and ( w_34270 , w_34271 , \13257_b0 );
or ( \13365_b1 , \6824_b1 , \13257_b1 );
not ( \13257_b1 , w_34272 );
and ( \13365_b0 , \6824_b0 , w_34273 );
and ( w_34272 , w_34273 , \13257_b0 );
or ( \13367_b1 , \13237_b1 , \13241_b1 );
not ( \13241_b1 , w_34274 );
and ( \13367_b0 , \13237_b0 , w_34275 );
and ( w_34274 , w_34275 , \13241_b0 );
or ( \13368_b1 , \13241_b1 , \13246_b1 );
not ( \13246_b1 , w_34276 );
and ( \13368_b0 , \13241_b0 , w_34277 );
and ( w_34276 , w_34277 , \13246_b0 );
or ( \13369_b1 , \13237_b1 , \13246_b1 );
not ( \13246_b1 , w_34278 );
and ( \13369_b0 , \13237_b0 , w_34279 );
and ( w_34278 , w_34279 , \13246_b0 );
or ( \13371_b1 , \13366_b1 , \13370_b1 );
xor ( \13371_b0 , \13366_b0 , w_34280 );
not ( w_34280 , w_34281 );
and ( w_34281 , \13370_b1 , \13370_b0 );
or ( \13372_b1 , \13223_b1 , \13227_b1 );
not ( \13227_b1 , w_34282 );
and ( \13372_b0 , \13223_b0 , w_34283 );
and ( w_34282 , w_34283 , \13227_b0 );
or ( \13373_b1 , \13227_b1 , \13232_b1 );
not ( \13232_b1 , w_34284 );
and ( \13373_b0 , \13227_b0 , w_34285 );
and ( w_34284 , w_34285 , \13232_b0 );
or ( \13374_b1 , \13223_b1 , \13232_b1 );
not ( \13232_b1 , w_34286 );
and ( \13374_b0 , \13223_b0 , w_34287 );
and ( w_34286 , w_34287 , \13232_b0 );
or ( \13376_b1 , \13371_b1 , \13375_b1 );
xor ( \13376_b0 , \13371_b0 , w_34288 );
not ( w_34288 , w_34289 );
and ( w_34289 , \13375_b1 , \13375_b0 );
or ( \13377_b1 , \13362_b1 , \13376_b1 );
xor ( \13377_b0 , \13362_b0 , w_34290 );
not ( w_34290 , w_34291 );
and ( w_34291 , \13376_b1 , \13376_b0 );
or ( \13378_b1 , \13353_b1 , \13377_b1 );
xor ( \13378_b0 , \13353_b0 , w_34292 );
not ( w_34292 , w_34293 );
and ( w_34293 , \13377_b1 , \13377_b0 );
or ( \13379_b1 , \13198_b1 , \13209_b1 );
not ( \13209_b1 , w_34294 );
and ( \13379_b0 , \13198_b0 , w_34295 );
and ( w_34294 , w_34295 , \13209_b0 );
or ( \13380_b1 , \13209_b1 , \13303_b1 );
not ( \13303_b1 , w_34296 );
and ( \13380_b0 , \13209_b0 , w_34297 );
and ( w_34296 , w_34297 , \13303_b0 );
or ( \13381_b1 , \13198_b1 , \13303_b1 );
not ( \13303_b1 , w_34298 );
and ( \13381_b0 , \13198_b0 , w_34299 );
and ( w_34298 , w_34299 , \13303_b0 );
or ( \13383_b1 , \13378_b1 , w_34301 );
not ( w_34301 , w_34302 );
and ( \13383_b0 , \13378_b0 , w_34303 );
and ( w_34302 ,  , w_34303 );
buf ( w_34301 , \13382_b1 );
not ( w_34301 , w_34304 );
not (  , w_34305 );
and ( w_34304 , w_34305 , \13382_b0 );
or ( \13384_b1 , \13341_b1 , \13345_b1 );
not ( \13345_b1 , w_34306 );
and ( \13384_b0 , \13341_b0 , w_34307 );
and ( w_34306 , w_34307 , \13345_b0 );
or ( \13385_b1 , \13345_b1 , \13350_b1 );
not ( \13350_b1 , w_34308 );
and ( \13385_b0 , \13345_b0 , w_34309 );
and ( w_34308 , w_34309 , \13350_b0 );
or ( \13386_b1 , \13341_b1 , \13350_b1 );
not ( \13350_b1 , w_34310 );
and ( \13386_b0 , \13341_b0 , w_34311 );
and ( w_34310 , w_34311 , \13350_b0 );
or ( \13388_b1 , \13316_b1 , \13324_b1 );
not ( \13324_b1 , w_34312 );
and ( \13388_b0 , \13316_b0 , w_34313 );
and ( w_34312 , w_34313 , \13324_b0 );
or ( \13389_b1 , \13324_b1 , \13336_b1 );
not ( \13336_b1 , w_34314 );
and ( \13389_b0 , \13324_b0 , w_34315 );
and ( w_34314 , w_34315 , \13336_b0 );
or ( \13390_b1 , \13316_b1 , \13336_b1 );
not ( \13336_b1 , w_34316 );
and ( \13390_b0 , \13316_b0 , w_34317 );
and ( w_34316 , w_34317 , \13336_b0 );
or ( \13392_b1 , \13387_b1 , \13391_b1 );
xor ( \13392_b0 , \13387_b0 , w_34318 );
not ( w_34318 , w_34319 );
and ( w_34319 , \13391_b1 , \13391_b0 );
or ( \13393_b1 , \7845_b1 , \7847_b1 );
xor ( \13393_b0 , \7845_b0 , w_34320 );
not ( w_34320 , w_34321 );
and ( w_34321 , \7847_b1 , \7847_b0 );
or ( \13394_b1 , \13393_b1 , \7850_b1 );
xor ( \13394_b0 , \13393_b0 , w_34322 );
not ( w_34322 , w_34323 );
and ( w_34323 , \7850_b1 , \7850_b0 );
or ( \13395_b1 , \7834_b1 , \7836_b1 );
xor ( \13395_b0 , \7834_b0 , w_34324 );
not ( w_34324 , w_34325 );
and ( w_34325 , \7836_b1 , \7836_b0 );
or ( \13396_b1 , \13395_b1 , \7839_b1 );
xor ( \13396_b0 , \13395_b0 , w_34326 );
not ( w_34326 , w_34327 );
and ( w_34327 , \7839_b1 , \7839_b0 );
or ( \13397_b1 , \13394_b1 , \13396_b1 );
xor ( \13397_b0 , \13394_b0 , w_34328 );
not ( w_34328 , w_34329 );
and ( w_34329 , \13396_b1 , \13396_b0 );
or ( \13398_b1 , \7782_b1 , \7798_b1 );
xor ( \13398_b0 , \7782_b0 , w_34330 );
not ( w_34330 , w_34331 );
and ( w_34331 , \7798_b1 , \7798_b0 );
or ( \13399_b1 , \13398_b1 , \7815_b1 );
xor ( \13399_b0 , \13398_b0 , w_34332 );
not ( w_34332 , w_34333 );
and ( w_34333 , \7815_b1 , \7815_b0 );
or ( \13400_b1 , \13397_b1 , \13399_b1 );
xor ( \13400_b0 , \13397_b0 , w_34334 );
not ( w_34334 , w_34335 );
and ( w_34335 , \13399_b1 , \13399_b0 );
or ( \13401_b1 , \13392_b1 , \13400_b1 );
xor ( \13401_b0 , \13392_b0 , w_34336 );
not ( w_34336 , w_34337 );
and ( w_34337 , \13400_b1 , \13400_b0 );
or ( \13402_b1 , \13357_b1 , \13361_b1 );
not ( \13361_b1 , w_34338 );
and ( \13402_b0 , \13357_b0 , w_34339 );
and ( w_34338 , w_34339 , \13361_b0 );
or ( \13403_b1 , \13361_b1 , \13376_b1 );
not ( \13376_b1 , w_34340 );
and ( \13403_b0 , \13361_b0 , w_34341 );
and ( w_34340 , w_34341 , \13376_b0 );
or ( \13404_b1 , \13357_b1 , \13376_b1 );
not ( \13376_b1 , w_34342 );
and ( \13404_b0 , \13357_b0 , w_34343 );
and ( w_34342 , w_34343 , \13376_b0 );
or ( \13406_b1 , \13337_b1 , \13351_b1 );
not ( \13351_b1 , w_34344 );
and ( \13406_b0 , \13337_b0 , w_34345 );
and ( w_34344 , w_34345 , \13351_b0 );
or ( \13407_b1 , \13405_b1 , \13406_b1 );
xor ( \13407_b0 , \13405_b0 , w_34346 );
not ( w_34346 , w_34347 );
and ( w_34347 , \13406_b1 , \13406_b0 );
or ( \13408_b1 , \13366_b1 , \13370_b1 );
not ( \13370_b1 , w_34348 );
and ( \13408_b0 , \13366_b0 , w_34349 );
and ( w_34348 , w_34349 , \13370_b0 );
or ( \13409_b1 , \13370_b1 , \13375_b1 );
not ( \13375_b1 , w_34350 );
and ( \13409_b0 , \13370_b0 , w_34351 );
and ( w_34350 , w_34351 , \13375_b0 );
or ( \13410_b1 , \13366_b1 , \13375_b1 );
not ( \13375_b1 , w_34352 );
and ( \13410_b0 , \13366_b0 , w_34353 );
and ( w_34352 , w_34353 , \13375_b0 );
or ( \13412_b1 , \13329_b1 , \13330_b1 );
not ( \13330_b1 , w_34354 );
and ( \13412_b0 , \13329_b0 , w_34355 );
and ( w_34354 , w_34355 , \13330_b0 );
or ( \13413_b1 , \13330_b1 , \13335_b1 );
not ( \13335_b1 , w_34356 );
and ( \13413_b0 , \13330_b0 , w_34357 );
and ( w_34356 , w_34357 , \13335_b0 );
or ( \13414_b1 , \13329_b1 , \13335_b1 );
not ( \13335_b1 , w_34358 );
and ( \13414_b0 , \13329_b0 , w_34359 );
and ( w_34358 , w_34359 , \13335_b0 );
or ( \13416_b1 , \13411_b1 , \13415_b1 );
xor ( \13416_b0 , \13411_b0 , w_34360 );
not ( w_34360 , w_34361 );
and ( w_34361 , \13415_b1 , \13415_b0 );
or ( \13417_b1 , \13318_b1 , \13320_b1 );
not ( \13320_b1 , w_34362 );
and ( \13417_b0 , \13318_b0 , w_34363 );
and ( w_34362 , w_34363 , \13320_b0 );
or ( \13418_b1 , \13320_b1 , \13323_b1 );
not ( \13323_b1 , w_34364 );
and ( \13418_b0 , \13320_b0 , w_34365 );
and ( w_34364 , w_34365 , \13323_b0 );
or ( \13419_b1 , \13318_b1 , \13323_b1 );
not ( \13323_b1 , w_34366 );
and ( \13419_b0 , \13318_b0 , w_34367 );
and ( w_34366 , w_34367 , \13323_b0 );
or ( \13421_b1 , \13416_b1 , \13420_b1 );
xor ( \13421_b0 , \13416_b0 , w_34368 );
not ( w_34368 , w_34369 );
and ( w_34369 , \13420_b1 , \13420_b0 );
or ( \13422_b1 , \13407_b1 , \13421_b1 );
xor ( \13422_b0 , \13407_b0 , w_34370 );
not ( w_34370 , w_34371 );
and ( w_34371 , \13421_b1 , \13421_b0 );
or ( \13423_b1 , \13401_b1 , \13422_b1 );
xor ( \13423_b0 , \13401_b0 , w_34372 );
not ( w_34372 , w_34373 );
and ( w_34373 , \13422_b1 , \13422_b0 );
or ( \13424_b1 , \13314_b1 , \13352_b1 );
not ( \13352_b1 , w_34374 );
and ( \13424_b0 , \13314_b0 , w_34375 );
and ( w_34374 , w_34375 , \13352_b0 );
or ( \13425_b1 , \13352_b1 , \13377_b1 );
not ( \13377_b1 , w_34376 );
and ( \13425_b0 , \13352_b0 , w_34377 );
and ( w_34376 , w_34377 , \13377_b0 );
or ( \13426_b1 , \13314_b1 , \13377_b1 );
not ( \13377_b1 , w_34378 );
and ( \13426_b0 , \13314_b0 , w_34379 );
and ( w_34378 , w_34379 , \13377_b0 );
or ( \13428_b1 , \13423_b1 , w_34381 );
not ( w_34381 , w_34382 );
and ( \13428_b0 , \13423_b0 , w_34383 );
and ( w_34382 ,  , w_34383 );
buf ( w_34381 , \13427_b1 );
not ( w_34381 , w_34384 );
not (  , w_34385 );
and ( w_34384 , w_34385 , \13427_b0 );
or ( \13429_b1 , \13383_b1 , w_34387 );
not ( w_34387 , w_34388 );
and ( \13429_b0 , \13383_b0 , w_34389 );
and ( w_34388 ,  , w_34389 );
buf ( w_34387 , \13428_b1 );
not ( w_34387 , w_34390 );
not (  , w_34391 );
and ( w_34390 , w_34391 , \13428_b0 );
or ( \13430_b1 , \13310_b1 , w_34393 );
not ( w_34393 , w_34394 );
and ( \13430_b0 , \13310_b0 , w_34395 );
and ( w_34394 ,  , w_34395 );
buf ( w_34393 , \13429_b1 );
not ( w_34393 , w_34396 );
not (  , w_34397 );
and ( w_34396 , w_34397 , \13429_b0 );
or ( \13431_b1 , \13405_b1 , \13406_b1 );
not ( \13406_b1 , w_34398 );
and ( \13431_b0 , \13405_b0 , w_34399 );
and ( w_34398 , w_34399 , \13406_b0 );
or ( \13432_b1 , \13406_b1 , \13421_b1 );
not ( \13421_b1 , w_34400 );
and ( \13432_b0 , \13406_b0 , w_34401 );
and ( w_34400 , w_34401 , \13421_b0 );
or ( \13433_b1 , \13405_b1 , \13421_b1 );
not ( \13421_b1 , w_34402 );
and ( \13433_b0 , \13405_b0 , w_34403 );
and ( w_34402 , w_34403 , \13421_b0 );
or ( \13435_b1 , \13387_b1 , \13391_b1 );
not ( \13391_b1 , w_34404 );
and ( \13435_b0 , \13387_b0 , w_34405 );
and ( w_34404 , w_34405 , \13391_b0 );
or ( \13436_b1 , \13391_b1 , \13400_b1 );
not ( \13400_b1 , w_34406 );
and ( \13436_b0 , \13391_b0 , w_34407 );
and ( w_34406 , w_34407 , \13400_b0 );
or ( \13437_b1 , \13387_b1 , \13400_b1 );
not ( \13400_b1 , w_34408 );
and ( \13437_b0 , \13387_b0 , w_34409 );
and ( w_34408 , w_34409 , \13400_b0 );
or ( \13439_b1 , \7016_b1 , \7071_b1 );
xor ( \13439_b0 , \7016_b0 , w_34410 );
not ( w_34410 , w_34411 );
and ( w_34411 , \7071_b1 , \7071_b0 );
or ( \13440_b1 , \13439_b1 , \7127_b1 );
xor ( \13440_b0 , \13439_b0 , w_34412 );
not ( w_34412 , w_34413 );
and ( w_34413 , \7127_b1 , \7127_b0 );
or ( \13441_b1 , \7858_b1 , \7860_b1 );
xor ( \13441_b0 , \7858_b0 , w_34414 );
not ( w_34414 , w_34415 );
and ( w_34415 , \7860_b1 , \7860_b0 );
or ( \13442_b1 , \13441_b1 , \7863_b1 );
xor ( \13442_b0 , \13441_b0 , w_34416 );
not ( w_34416 , w_34417 );
and ( w_34417 , \7863_b1 , \7863_b0 );
or ( \13443_b1 , \13440_b1 , \13442_b1 );
xor ( \13443_b0 , \13440_b0 , w_34418 );
not ( w_34418 , w_34419 );
and ( w_34419 , \13442_b1 , \13442_b0 );
or ( \13444_b1 , \7818_b1 , \7842_b1 );
xor ( \13444_b0 , \7818_b0 , w_34420 );
not ( w_34420 , w_34421 );
and ( w_34421 , \7842_b1 , \7842_b0 );
or ( \13445_b1 , \13444_b1 , \7853_b1 );
xor ( \13445_b0 , \13444_b0 , w_34422 );
not ( w_34422 , w_34423 );
and ( w_34423 , \7853_b1 , \7853_b0 );
or ( \13446_b1 , \13443_b1 , \13445_b1 );
xor ( \13446_b0 , \13443_b0 , w_34424 );
not ( w_34424 , w_34425 );
and ( w_34425 , \13445_b1 , \13445_b0 );
or ( \13447_b1 , \13438_b1 , \13446_b1 );
xor ( \13447_b0 , \13438_b0 , w_34426 );
not ( w_34426 , w_34427 );
and ( w_34427 , \13446_b1 , \13446_b0 );
or ( \13448_b1 , \13411_b1 , \13415_b1 );
not ( \13415_b1 , w_34428 );
and ( \13448_b0 , \13411_b0 , w_34429 );
and ( w_34428 , w_34429 , \13415_b0 );
or ( \13449_b1 , \13415_b1 , \13420_b1 );
not ( \13420_b1 , w_34430 );
and ( \13449_b0 , \13415_b0 , w_34431 );
and ( w_34430 , w_34431 , \13420_b0 );
or ( \13450_b1 , \13411_b1 , \13420_b1 );
not ( \13420_b1 , w_34432 );
and ( \13450_b0 , \13411_b0 , w_34433 );
and ( w_34432 , w_34433 , \13420_b0 );
or ( \13452_b1 , \13394_b1 , \13396_b1 );
not ( \13396_b1 , w_34434 );
and ( \13452_b0 , \13394_b0 , w_34435 );
and ( w_34434 , w_34435 , \13396_b0 );
or ( \13453_b1 , \13396_b1 , \13399_b1 );
not ( \13399_b1 , w_34436 );
and ( \13453_b0 , \13396_b0 , w_34437 );
and ( w_34436 , w_34437 , \13399_b0 );
or ( \13454_b1 , \13394_b1 , \13399_b1 );
not ( \13399_b1 , w_34438 );
and ( \13454_b0 , \13394_b0 , w_34439 );
and ( w_34438 , w_34439 , \13399_b0 );
or ( \13456_b1 , \13451_b1 , \13455_b1 );
xor ( \13456_b0 , \13451_b0 , w_34440 );
not ( w_34440 , w_34441 );
and ( w_34441 , \13455_b1 , \13455_b0 );
or ( \13457_b1 , \7185_b1 , \7213_b1 );
xor ( \13457_b0 , \7185_b0 , w_34442 );
not ( w_34442 , w_34443 );
and ( w_34443 , \7213_b1 , \7213_b0 );
or ( \13458_b1 , \13457_b1 , \7218_b1 );
xor ( \13458_b0 , \13457_b0 , w_34444 );
not ( w_34444 , w_34445 );
and ( w_34445 , \7218_b1 , \7218_b0 );
or ( \13459_b1 , \13456_b1 , \13458_b1 );
xor ( \13459_b0 , \13456_b0 , w_34446 );
not ( w_34446 , w_34447 );
and ( w_34447 , \13458_b1 , \13458_b0 );
or ( \13460_b1 , \13447_b1 , \13459_b1 );
xor ( \13460_b0 , \13447_b0 , w_34448 );
not ( w_34448 , w_34449 );
and ( w_34449 , \13459_b1 , \13459_b0 );
or ( \13461_b1 , \13434_b1 , \13460_b1 );
xor ( \13461_b0 , \13434_b0 , w_34450 );
not ( w_34450 , w_34451 );
and ( w_34451 , \13460_b1 , \13460_b0 );
or ( \13462_b1 , \13401_b1 , \13422_b1 );
not ( \13422_b1 , w_34452 );
and ( \13462_b0 , \13401_b0 , w_34453 );
and ( w_34452 , w_34453 , \13422_b0 );
or ( \13463_b1 , \13461_b1 , w_34455 );
not ( w_34455 , w_34456 );
and ( \13463_b0 , \13461_b0 , w_34457 );
and ( w_34456 ,  , w_34457 );
buf ( w_34455 , \13462_b1 );
not ( w_34455 , w_34458 );
not (  , w_34459 );
and ( w_34458 , w_34459 , \13462_b0 );
or ( \13464_b1 , \13438_b1 , \13446_b1 );
not ( \13446_b1 , w_34460 );
and ( \13464_b0 , \13438_b0 , w_34461 );
and ( w_34460 , w_34461 , \13446_b0 );
or ( \13465_b1 , \13446_b1 , \13459_b1 );
not ( \13459_b1 , w_34462 );
and ( \13465_b0 , \13446_b0 , w_34463 );
and ( w_34462 , w_34463 , \13459_b0 );
or ( \13466_b1 , \13438_b1 , \13459_b1 );
not ( \13459_b1 , w_34464 );
and ( \13466_b0 , \13438_b0 , w_34465 );
and ( w_34464 , w_34465 , \13459_b0 );
or ( \13468_b1 , \7130_b1 , \7221_b1 );
xor ( \13468_b0 , \7130_b0 , w_34466 );
not ( w_34466 , w_34467 );
and ( w_34467 , \7221_b1 , \7221_b0 );
or ( \13469_b1 , \13468_b1 , \7258_b1 );
xor ( \13469_b0 , \13468_b0 , w_34468 );
not ( w_34468 , w_34469 );
and ( w_34469 , \7258_b1 , \7258_b0 );
or ( \13470_b1 , \7856_b1 , \7866_b1 );
xor ( \13470_b0 , \7856_b0 , w_34470 );
not ( w_34470 , w_34471 );
and ( w_34471 , \7866_b1 , \7866_b0 );
or ( \13471_b1 , \13470_b1 , \7869_b1 );
xor ( \13471_b0 , \13470_b0 , w_34472 );
not ( w_34472 , w_34473 );
and ( w_34473 , \7869_b1 , \7869_b0 );
or ( \13472_b1 , \13469_b1 , \13471_b1 );
xor ( \13472_b0 , \13469_b0 , w_34474 );
not ( w_34474 , w_34475 );
and ( w_34475 , \13471_b1 , \13471_b0 );
or ( \13473_b1 , \13467_b1 , \13472_b1 );
xor ( \13473_b0 , \13467_b0 , w_34476 );
not ( w_34476 , w_34477 );
and ( w_34477 , \13472_b1 , \13472_b0 );
or ( \13474_b1 , \13451_b1 , \13455_b1 );
not ( \13455_b1 , w_34478 );
and ( \13474_b0 , \13451_b0 , w_34479 );
and ( w_34478 , w_34479 , \13455_b0 );
or ( \13475_b1 , \13455_b1 , \13458_b1 );
not ( \13458_b1 , w_34480 );
and ( \13475_b0 , \13455_b0 , w_34481 );
and ( w_34480 , w_34481 , \13458_b0 );
or ( \13476_b1 , \13451_b1 , \13458_b1 );
not ( \13458_b1 , w_34482 );
and ( \13476_b0 , \13451_b0 , w_34483 );
and ( w_34482 , w_34483 , \13458_b0 );
or ( \13478_b1 , \13440_b1 , \13442_b1 );
not ( \13442_b1 , w_34484 );
and ( \13478_b0 , \13440_b0 , w_34485 );
and ( w_34484 , w_34485 , \13442_b0 );
or ( \13479_b1 , \13442_b1 , \13445_b1 );
not ( \13445_b1 , w_34486 );
and ( \13479_b0 , \13442_b0 , w_34487 );
and ( w_34486 , w_34487 , \13445_b0 );
or ( \13480_b1 , \13440_b1 , \13445_b1 );
not ( \13445_b1 , w_34488 );
and ( \13480_b0 , \13440_b0 , w_34489 );
and ( w_34488 , w_34489 , \13445_b0 );
or ( \13482_b1 , \13477_b1 , \13481_b1 );
xor ( \13482_b0 , \13477_b0 , w_34490 );
not ( w_34490 , w_34491 );
and ( w_34491 , \13481_b1 , \13481_b0 );
or ( \13483_b1 , \7271_b1 , \7315_b1 );
xor ( \13483_b0 , \7271_b0 , w_34492 );
not ( w_34492 , w_34493 );
and ( w_34493 , \7315_b1 , \7315_b0 );
or ( \13484_b1 , \13483_b1 , \7338_b1 );
xor ( \13484_b0 , \13483_b0 , w_34494 );
not ( w_34494 , w_34495 );
and ( w_34495 , \7338_b1 , \7338_b0 );
or ( \13485_b1 , \13482_b1 , \13484_b1 );
xor ( \13485_b0 , \13482_b0 , w_34496 );
not ( w_34496 , w_34497 );
and ( w_34497 , \13484_b1 , \13484_b0 );
or ( \13486_b1 , \13473_b1 , \13485_b1 );
xor ( \13486_b0 , \13473_b0 , w_34498 );
not ( w_34498 , w_34499 );
and ( w_34499 , \13485_b1 , \13485_b0 );
or ( \13487_b1 , \13434_b1 , \13460_b1 );
not ( \13460_b1 , w_34500 );
and ( \13487_b0 , \13434_b0 , w_34501 );
and ( w_34500 , w_34501 , \13460_b0 );
or ( \13488_b1 , \13486_b1 , w_34503 );
not ( w_34503 , w_34504 );
and ( \13488_b0 , \13486_b0 , w_34505 );
and ( w_34504 ,  , w_34505 );
buf ( w_34503 , \13487_b1 );
not ( w_34503 , w_34506 );
not (  , w_34507 );
and ( w_34506 , w_34507 , \13487_b0 );
or ( \13489_b1 , \13463_b1 , w_34509 );
not ( w_34509 , w_34510 );
and ( \13489_b0 , \13463_b0 , w_34511 );
and ( w_34510 ,  , w_34511 );
buf ( w_34509 , \13488_b1 );
not ( w_34509 , w_34512 );
not (  , w_34513 );
and ( w_34512 , w_34513 , \13488_b0 );
or ( \13490_b1 , \13477_b1 , \13481_b1 );
not ( \13481_b1 , w_34514 );
and ( \13490_b0 , \13477_b0 , w_34515 );
and ( w_34514 , w_34515 , \13481_b0 );
or ( \13491_b1 , \13481_b1 , \13484_b1 );
not ( \13484_b1 , w_34516 );
and ( \13491_b0 , \13481_b0 , w_34517 );
and ( w_34516 , w_34517 , \13484_b0 );
or ( \13492_b1 , \13477_b1 , \13484_b1 );
not ( \13484_b1 , w_34518 );
and ( \13492_b0 , \13477_b0 , w_34519 );
and ( w_34518 , w_34519 , \13484_b0 );
or ( \13494_b1 , \13469_b1 , \13471_b1 );
not ( \13471_b1 , w_34520 );
and ( \13494_b0 , \13469_b0 , w_34521 );
and ( w_34520 , w_34521 , \13471_b0 );
or ( \13495_b1 , \13493_b1 , \13494_b1 );
xor ( \13495_b0 , \13493_b0 , w_34522 );
not ( w_34522 , w_34523 );
and ( w_34523 , \13494_b1 , \13494_b0 );
or ( \13496_b1 , \7872_b1 , \7873_b1 );
xor ( \13496_b0 , \7872_b0 , w_34524 );
not ( w_34524 , w_34525 );
and ( w_34525 , \7873_b1 , \7873_b0 );
or ( \13497_b1 , \13496_b1 , \7876_b1 );
xor ( \13497_b0 , \13496_b0 , w_34526 );
not ( w_34526 , w_34527 );
and ( w_34527 , \7876_b1 , \7876_b0 );
or ( \13498_b1 , \13495_b1 , \13497_b1 );
xor ( \13498_b0 , \13495_b0 , w_34528 );
not ( w_34528 , w_34529 );
and ( w_34529 , \13497_b1 , \13497_b0 );
or ( \13499_b1 , \13467_b1 , \13472_b1 );
not ( \13472_b1 , w_34530 );
and ( \13499_b0 , \13467_b0 , w_34531 );
and ( w_34530 , w_34531 , \13472_b0 );
or ( \13500_b1 , \13472_b1 , \13485_b1 );
not ( \13485_b1 , w_34532 );
and ( \13500_b0 , \13472_b0 , w_34533 );
and ( w_34532 , w_34533 , \13485_b0 );
or ( \13501_b1 , \13467_b1 , \13485_b1 );
not ( \13485_b1 , w_34534 );
and ( \13501_b0 , \13467_b0 , w_34535 );
and ( w_34534 , w_34535 , \13485_b0 );
or ( \13503_b1 , \13498_b1 , w_34537 );
not ( w_34537 , w_34538 );
and ( \13503_b0 , \13498_b0 , w_34539 );
and ( w_34538 ,  , w_34539 );
buf ( w_34537 , \13502_b1 );
not ( w_34537 , w_34540 );
not (  , w_34541 );
and ( w_34540 , w_34541 , \13502_b0 );
or ( \13504_b1 , \7879_b1 , \7880_b1 );
xor ( \13504_b0 , \7879_b0 , w_34542 );
not ( w_34542 , w_34543 );
and ( w_34543 , \7880_b1 , \7880_b0 );
or ( \13505_b1 , \13504_b1 , \7883_b1 );
xor ( \13505_b0 , \13504_b0 , w_34544 );
not ( w_34544 , w_34545 );
and ( w_34545 , \7883_b1 , \7883_b0 );
or ( \13506_b1 , \13493_b1 , \13494_b1 );
not ( \13494_b1 , w_34546 );
and ( \13506_b0 , \13493_b0 , w_34547 );
and ( w_34546 , w_34547 , \13494_b0 );
or ( \13507_b1 , \13494_b1 , \13497_b1 );
not ( \13497_b1 , w_34548 );
and ( \13507_b0 , \13494_b0 , w_34549 );
and ( w_34548 , w_34549 , \13497_b0 );
or ( \13508_b1 , \13493_b1 , \13497_b1 );
not ( \13497_b1 , w_34550 );
and ( \13508_b0 , \13493_b0 , w_34551 );
and ( w_34550 , w_34551 , \13497_b0 );
or ( \13510_b1 , \13505_b1 , w_34553 );
not ( w_34553 , w_34554 );
and ( \13510_b0 , \13505_b0 , w_34555 );
and ( w_34554 ,  , w_34555 );
buf ( w_34553 , \13509_b1 );
not ( w_34553 , w_34556 );
not (  , w_34557 );
and ( w_34556 , w_34557 , \13509_b0 );
or ( \13511_b1 , \13503_b1 , w_34559 );
not ( w_34559 , w_34560 );
and ( \13511_b0 , \13503_b0 , w_34561 );
and ( w_34560 ,  , w_34561 );
buf ( w_34559 , \13510_b1 );
not ( w_34559 , w_34562 );
not (  , w_34563 );
and ( w_34562 , w_34563 , \13510_b0 );
or ( \13512_b1 , \13489_b1 , w_34565 );
not ( w_34565 , w_34566 );
and ( \13512_b0 , \13489_b0 , w_34567 );
and ( w_34566 ,  , w_34567 );
buf ( w_34565 , \13511_b1 );
not ( w_34565 , w_34568 );
not (  , w_34569 );
and ( w_34568 , w_34569 , \13511_b0 );
or ( \13513_b1 , \13430_b1 , w_34571 );
not ( w_34571 , w_34572 );
and ( \13513_b0 , \13430_b0 , w_34573 );
and ( w_34572 ,  , w_34573 );
buf ( w_34571 , \13512_b1 );
not ( w_34571 , w_34574 );
not (  , w_34575 );
and ( w_34574 , w_34575 , \13512_b0 );
or ( \13514_b1 , \13083_b1 , w_34577 );
not ( w_34577 , w_34578 );
and ( \13514_b0 , \13083_b0 , w_34579 );
and ( w_34578 ,  , w_34579 );
buf ( w_34577 , \13513_b1 );
not ( w_34577 , w_34580 );
not (  , w_34581 );
and ( w_34580 , w_34581 , \13513_b0 );
or ( \13515_b1 , \6018_b1 , \6991_b1 );
not ( \6991_b1 , w_34582 );
and ( \13515_b0 , \6018_b0 , w_34583 );
and ( w_34582 , w_34583 , \6991_b0 );
or ( \13516_b1 , \5986_b1 , \6988_b1 );
not ( \6988_b1 , w_34584 );
and ( \13516_b0 , \5986_b0 , w_34585 );
and ( w_34584 , w_34585 , \6988_b0 );
or ( \13517_b1 , \13515_b1 , w_34587 );
not ( w_34587 , w_34588 );
and ( \13517_b0 , \13515_b0 , w_34589 );
and ( w_34588 ,  , w_34589 );
buf ( w_34587 , \13516_b1 );
not ( w_34587 , w_34590 );
not (  , w_34591 );
and ( w_34590 , w_34591 , \13516_b0 );
or ( \13518_b1 , \13517_b1 , w_34592 );
xor ( \13518_b0 , \13517_b0 , w_34594 );
not ( w_34594 , w_34595 );
and ( w_34595 , w_34592 , w_34593 );
buf ( w_34592 , \6985_b1 );
not ( w_34592 , w_34596 );
not ( w_34593 , w_34597 );
and ( w_34596 , w_34597 , \6985_b0 );
or ( \13519_b1 , \6041_b1 , \7006_b1 );
not ( \7006_b1 , w_34598 );
and ( \13519_b0 , \6041_b0 , w_34599 );
and ( w_34598 , w_34599 , \7006_b0 );
or ( \13520_b1 , \6006_b1 , \7004_b1 );
not ( \7004_b1 , w_34600 );
and ( \13520_b0 , \6006_b0 , w_34601 );
and ( w_34600 , w_34601 , \7004_b0 );
or ( \13521_b1 , \13519_b1 , w_34603 );
not ( w_34603 , w_34604 );
and ( \13521_b0 , \13519_b0 , w_34605 );
and ( w_34604 ,  , w_34605 );
buf ( w_34603 , \13520_b1 );
not ( w_34603 , w_34606 );
not (  , w_34607 );
and ( w_34606 , w_34607 , \13520_b0 );
or ( \13522_b1 , \13521_b1 , w_34608 );
xor ( \13522_b0 , \13521_b0 , w_34610 );
not ( w_34610 , w_34611 );
and ( w_34611 , w_34608 , w_34609 );
buf ( w_34608 , \7012_b1 );
not ( w_34608 , w_34612 );
not ( w_34609 , w_34613 );
and ( w_34612 , w_34613 , \7012_b0 );
or ( \13523_b1 , \13518_b1 , \13522_b1 );
xor ( \13523_b0 , \13518_b0 , w_34614 );
not ( w_34614 , w_34615 );
and ( w_34615 , \13522_b1 , \13522_b0 );
or ( \13524_b1 , \6057_b1 , \7026_b1 );
not ( \7026_b1 , w_34616 );
and ( \13524_b0 , \6057_b0 , w_34617 );
and ( w_34616 , w_34617 , \7026_b0 );
or ( \13525_b1 , \6029_b1 , \7024_b1 );
not ( \7024_b1 , w_34618 );
and ( \13525_b0 , \6029_b0 , w_34619 );
and ( w_34618 , w_34619 , \7024_b0 );
or ( \13526_b1 , \13524_b1 , w_34621 );
not ( w_34621 , w_34622 );
and ( \13526_b0 , \13524_b0 , w_34623 );
and ( w_34622 ,  , w_34623 );
buf ( w_34621 , \13525_b1 );
not ( w_34621 , w_34624 );
not (  , w_34625 );
and ( w_34624 , w_34625 , \13525_b0 );
or ( \13527_b1 , \13526_b1 , w_34626 );
xor ( \13527_b0 , \13526_b0 , w_34628 );
not ( w_34628 , w_34629 );
and ( w_34629 , w_34626 , w_34627 );
buf ( w_34626 , \7032_b1 );
not ( w_34626 , w_34630 );
not ( w_34627 , w_34631 );
and ( w_34630 , w_34631 , \7032_b0 );
or ( \13528_b1 , \13523_b1 , \13527_b1 );
xor ( \13528_b0 , \13523_b0 , w_34632 );
not ( w_34632 , w_34633 );
and ( w_34633 , \13527_b1 , \13527_b0 );
or ( \13529_b1 , \6006_b1 , \6991_b1 );
not ( \6991_b1 , w_34634 );
and ( \13529_b0 , \6006_b0 , w_34635 );
and ( w_34634 , w_34635 , \6991_b0 );
or ( \13530_b1 , \6018_b1 , \6988_b1 );
not ( \6988_b1 , w_34636 );
and ( \13530_b0 , \6018_b0 , w_34637 );
and ( w_34636 , w_34637 , \6988_b0 );
or ( \13531_b1 , \13529_b1 , w_34639 );
not ( w_34639 , w_34640 );
and ( \13531_b0 , \13529_b0 , w_34641 );
and ( w_34640 ,  , w_34641 );
buf ( w_34639 , \13530_b1 );
not ( w_34639 , w_34642 );
not (  , w_34643 );
and ( w_34642 , w_34643 , \13530_b0 );
or ( \13532_b1 , \13531_b1 , w_34644 );
xor ( \13532_b0 , \13531_b0 , w_34646 );
not ( w_34646 , w_34647 );
and ( w_34647 , w_34644 , w_34645 );
buf ( w_34644 , \6985_b1 );
not ( w_34644 , w_34648 );
not ( w_34645 , w_34649 );
and ( w_34648 , w_34649 , \6985_b0 );
or ( \13533_b1 , \7049_b1 , \13532_b1 );
not ( \13532_b1 , w_34650 );
and ( \13533_b0 , \7049_b0 , w_34651 );
and ( w_34650 , w_34651 , \13532_b0 );
or ( \13534_b1 , \6029_b1 , \7006_b1 );
not ( \7006_b1 , w_34652 );
and ( \13534_b0 , \6029_b0 , w_34653 );
and ( w_34652 , w_34653 , \7006_b0 );
or ( \13535_b1 , \6041_b1 , \7004_b1 );
not ( \7004_b1 , w_34654 );
and ( \13535_b0 , \6041_b0 , w_34655 );
and ( w_34654 , w_34655 , \7004_b0 );
or ( \13536_b1 , \13534_b1 , w_34657 );
not ( w_34657 , w_34658 );
and ( \13536_b0 , \13534_b0 , w_34659 );
and ( w_34658 ,  , w_34659 );
buf ( w_34657 , \13535_b1 );
not ( w_34657 , w_34660 );
not (  , w_34661 );
and ( w_34660 , w_34661 , \13535_b0 );
or ( \13537_b1 , \13536_b1 , w_34662 );
xor ( \13537_b0 , \13536_b0 , w_34664 );
not ( w_34664 , w_34665 );
and ( w_34665 , w_34662 , w_34663 );
buf ( w_34662 , \7012_b1 );
not ( w_34662 , w_34666 );
not ( w_34663 , w_34667 );
and ( w_34666 , w_34667 , \7012_b0 );
or ( \13538_b1 , \13532_b1 , \13537_b1 );
not ( \13537_b1 , w_34668 );
and ( \13538_b0 , \13532_b0 , w_34669 );
and ( w_34668 , w_34669 , \13537_b0 );
or ( \13539_b1 , \7049_b1 , \13537_b1 );
not ( \13537_b1 , w_34670 );
and ( \13539_b0 , \7049_b0 , w_34671 );
and ( w_34670 , w_34671 , \13537_b0 );
or ( \13541_b1 , \6048_b1 , \7026_b1 );
not ( \7026_b1 , w_34672 );
and ( \13541_b0 , \6048_b0 , w_34673 );
and ( w_34672 , w_34673 , \7026_b0 );
or ( \13542_b1 , \6057_b1 , \7024_b1 );
not ( \7024_b1 , w_34674 );
and ( \13542_b0 , \6057_b0 , w_34675 );
and ( w_34674 , w_34675 , \7024_b0 );
or ( \13543_b1 , \13541_b1 , w_34677 );
not ( w_34677 , w_34678 );
and ( \13543_b0 , \13541_b0 , w_34679 );
and ( w_34678 ,  , w_34679 );
buf ( w_34677 , \13542_b1 );
not ( w_34677 , w_34680 );
not (  , w_34681 );
and ( w_34680 , w_34681 , \13542_b0 );
or ( \13544_b1 , \13543_b1 , w_34682 );
xor ( \13544_b0 , \13543_b0 , w_34684 );
not ( w_34684 , w_34685 );
and ( w_34685 , w_34682 , w_34683 );
buf ( w_34682 , \7032_b1 );
not ( w_34682 , w_34686 );
not ( w_34683 , w_34687 );
and ( w_34686 , w_34687 , \7032_b0 );
or ( \13545_b1 , \6065_b1 , w_34689 );
not ( w_34689 , w_34690 );
and ( \13545_b0 , \6065_b0 , w_34691 );
and ( w_34690 ,  , w_34691 );
buf ( w_34689 , \7041_b1 );
not ( w_34689 , w_34692 );
not (  , w_34693 );
and ( w_34692 , w_34693 , \7041_b0 );
or ( \13546_b1 , \13545_b1 , w_34694 );
xor ( \13546_b0 , \13545_b0 , w_34696 );
not ( w_34696 , w_34697 );
and ( w_34697 , w_34694 , w_34695 );
buf ( w_34694 , \7049_b1 );
not ( w_34694 , w_34698 );
not ( w_34695 , w_34699 );
and ( w_34698 , w_34699 , \7049_b0 );
or ( \13547_b1 , \13544_b1 , \13546_b1 );
not ( \13546_b1 , w_34700 );
and ( \13547_b0 , \13544_b0 , w_34701 );
and ( w_34700 , w_34701 , \13546_b0 );
or ( \13548_b1 , \13540_b1 , \13547_b1 );
xor ( \13548_b0 , \13540_b0 , w_34702 );
not ( w_34702 , w_34703 );
and ( w_34703 , \13547_b1 , \13547_b0 );
or ( \13549_b1 , \6065_b1 , \7043_b1 );
not ( \7043_b1 , w_34704 );
and ( \13549_b0 , \6065_b0 , w_34705 );
and ( w_34704 , w_34705 , \7043_b0 );
or ( \13550_b1 , \6048_b1 , \7041_b1 );
not ( \7041_b1 , w_34706 );
and ( \13550_b0 , \6048_b0 , w_34707 );
and ( w_34706 , w_34707 , \7041_b0 );
or ( \13551_b1 , \13549_b1 , w_34709 );
not ( w_34709 , w_34710 );
and ( \13551_b0 , \13549_b0 , w_34711 );
and ( w_34710 ,  , w_34711 );
buf ( w_34709 , \13550_b1 );
not ( w_34709 , w_34712 );
not (  , w_34713 );
and ( w_34712 , w_34713 , \13550_b0 );
or ( \13552_b1 , \13551_b1 , w_34714 );
xor ( \13552_b0 , \13551_b0 , w_34716 );
not ( w_34716 , w_34717 );
and ( w_34717 , w_34714 , w_34715 );
buf ( w_34714 , \7049_b1 );
not ( w_34714 , w_34718 );
not ( w_34715 , w_34719 );
and ( w_34718 , w_34719 , \7049_b0 );
or ( \13553_b1 , \13548_b1 , \13552_b1 );
xor ( \13553_b0 , \13548_b0 , w_34720 );
not ( w_34720 , w_34721 );
and ( w_34721 , \13552_b1 , \13552_b0 );
or ( \13554_b1 , \13528_b1 , \13553_b1 );
xor ( \13554_b0 , \13528_b0 , w_34722 );
not ( w_34722 , w_34723 );
and ( w_34723 , \13553_b1 , \13553_b0 );
or ( \13555_b1 , \6041_b1 , \6991_b1 );
not ( \6991_b1 , w_34724 );
and ( \13555_b0 , \6041_b0 , w_34725 );
and ( w_34724 , w_34725 , \6991_b0 );
or ( \13556_b1 , \6006_b1 , \6988_b1 );
not ( \6988_b1 , w_34726 );
and ( \13556_b0 , \6006_b0 , w_34727 );
and ( w_34726 , w_34727 , \6988_b0 );
or ( \13557_b1 , \13555_b1 , w_34729 );
not ( w_34729 , w_34730 );
and ( \13557_b0 , \13555_b0 , w_34731 );
and ( w_34730 ,  , w_34731 );
buf ( w_34729 , \13556_b1 );
not ( w_34729 , w_34732 );
not (  , w_34733 );
and ( w_34732 , w_34733 , \13556_b0 );
or ( \13558_b1 , \13557_b1 , w_34734 );
xor ( \13558_b0 , \13557_b0 , w_34736 );
not ( w_34736 , w_34737 );
and ( w_34737 , w_34734 , w_34735 );
buf ( w_34734 , \6985_b1 );
not ( w_34734 , w_34738 );
not ( w_34735 , w_34739 );
and ( w_34738 , w_34739 , \6985_b0 );
or ( \13559_b1 , \6057_b1 , \7006_b1 );
not ( \7006_b1 , w_34740 );
and ( \13559_b0 , \6057_b0 , w_34741 );
and ( w_34740 , w_34741 , \7006_b0 );
or ( \13560_b1 , \6029_b1 , \7004_b1 );
not ( \7004_b1 , w_34742 );
and ( \13560_b0 , \6029_b0 , w_34743 );
and ( w_34742 , w_34743 , \7004_b0 );
or ( \13561_b1 , \13559_b1 , w_34745 );
not ( w_34745 , w_34746 );
and ( \13561_b0 , \13559_b0 , w_34747 );
and ( w_34746 ,  , w_34747 );
buf ( w_34745 , \13560_b1 );
not ( w_34745 , w_34748 );
not (  , w_34749 );
and ( w_34748 , w_34749 , \13560_b0 );
or ( \13562_b1 , \13561_b1 , w_34750 );
xor ( \13562_b0 , \13561_b0 , w_34752 );
not ( w_34752 , w_34753 );
and ( w_34753 , w_34750 , w_34751 );
buf ( w_34750 , \7012_b1 );
not ( w_34750 , w_34754 );
not ( w_34751 , w_34755 );
and ( w_34754 , w_34755 , \7012_b0 );
or ( \13563_b1 , \13558_b1 , \13562_b1 );
not ( \13562_b1 , w_34756 );
and ( \13563_b0 , \13558_b0 , w_34757 );
and ( w_34756 , w_34757 , \13562_b0 );
or ( \13564_b1 , \6065_b1 , \7026_b1 );
not ( \7026_b1 , w_34758 );
and ( \13564_b0 , \6065_b0 , w_34759 );
and ( w_34758 , w_34759 , \7026_b0 );
or ( \13565_b1 , \6048_b1 , \7024_b1 );
not ( \7024_b1 , w_34760 );
and ( \13565_b0 , \6048_b0 , w_34761 );
and ( w_34760 , w_34761 , \7024_b0 );
or ( \13566_b1 , \13564_b1 , w_34763 );
not ( w_34763 , w_34764 );
and ( \13566_b0 , \13564_b0 , w_34765 );
and ( w_34764 ,  , w_34765 );
buf ( w_34763 , \13565_b1 );
not ( w_34763 , w_34766 );
not (  , w_34767 );
and ( w_34766 , w_34767 , \13565_b0 );
or ( \13567_b1 , \13566_b1 , w_34768 );
xor ( \13567_b0 , \13566_b0 , w_34770 );
not ( w_34770 , w_34771 );
and ( w_34771 , w_34768 , w_34769 );
buf ( w_34768 , \7032_b1 );
not ( w_34768 , w_34772 );
not ( w_34769 , w_34773 );
and ( w_34772 , w_34773 , \7032_b0 );
or ( \13568_b1 , \13562_b1 , \13567_b1 );
not ( \13567_b1 , w_34774 );
and ( \13568_b0 , \13562_b0 , w_34775 );
and ( w_34774 , w_34775 , \13567_b0 );
or ( \13569_b1 , \13558_b1 , \13567_b1 );
not ( \13567_b1 , w_34776 );
and ( \13569_b0 , \13558_b0 , w_34777 );
and ( w_34776 , w_34777 , \13567_b0 );
or ( \13571_b1 , \13544_b1 , \13546_b1 );
xor ( \13571_b0 , \13544_b0 , w_34778 );
not ( w_34778 , w_34779 );
and ( w_34779 , \13546_b1 , \13546_b0 );
or ( \13572_b1 , \13570_b1 , \13571_b1 );
not ( \13571_b1 , w_34780 );
and ( \13572_b0 , \13570_b0 , w_34781 );
and ( w_34780 , w_34781 , \13571_b0 );
or ( \13573_b1 , \7049_b1 , \13532_b1 );
xor ( \13573_b0 , \7049_b0 , w_34782 );
not ( w_34782 , w_34783 );
and ( w_34783 , \13532_b1 , \13532_b0 );
or ( \13574_b1 , \13573_b1 , \13537_b1 );
xor ( \13574_b0 , \13573_b0 , w_34784 );
not ( w_34784 , w_34785 );
and ( w_34785 , \13537_b1 , \13537_b0 );
or ( \13575_b1 , \13571_b1 , \13574_b1 );
not ( \13574_b1 , w_34786 );
and ( \13575_b0 , \13571_b0 , w_34787 );
and ( w_34786 , w_34787 , \13574_b0 );
or ( \13576_b1 , \13570_b1 , \13574_b1 );
not ( \13574_b1 , w_34788 );
and ( \13576_b0 , \13570_b0 , w_34789 );
and ( w_34788 , w_34789 , \13574_b0 );
or ( \13578_b1 , \13554_b1 , w_34791 );
not ( w_34791 , w_34792 );
and ( \13578_b0 , \13554_b0 , w_34793 );
and ( w_34792 ,  , w_34793 );
buf ( w_34791 , \13577_b1 );
not ( w_34791 , w_34794 );
not (  , w_34795 );
and ( w_34794 , w_34795 , \13577_b0 );
or ( \13579_b1 , \13540_b1 , \13547_b1 );
not ( \13547_b1 , w_34796 );
and ( \13579_b0 , \13540_b0 , w_34797 );
and ( w_34796 , w_34797 , \13547_b0 );
or ( \13580_b1 , \13547_b1 , \13552_b1 );
not ( \13552_b1 , w_34798 );
and ( \13580_b0 , \13547_b0 , w_34799 );
and ( w_34798 , w_34799 , \13552_b0 );
or ( \13581_b1 , \13540_b1 , \13552_b1 );
not ( \13552_b1 , w_34800 );
and ( \13581_b0 , \13540_b0 , w_34801 );
and ( w_34800 , w_34801 , \13552_b0 );
or ( \13583_b1 , \13518_b1 , \13522_b1 );
not ( \13522_b1 , w_34802 );
and ( \13583_b0 , \13518_b0 , w_34803 );
and ( w_34802 , w_34803 , \13522_b0 );
or ( \13584_b1 , \13522_b1 , \13527_b1 );
not ( \13527_b1 , w_34804 );
and ( \13584_b0 , \13522_b0 , w_34805 );
and ( w_34804 , w_34805 , \13527_b0 );
or ( \13585_b1 , \13518_b1 , \13527_b1 );
not ( \13527_b1 , w_34806 );
and ( \13585_b0 , \13518_b0 , w_34807 );
and ( w_34806 , w_34807 , \13527_b0 );
or ( \13587_b1 , \6029_b1 , \7026_b1 );
not ( \7026_b1 , w_34808 );
and ( \13587_b0 , \6029_b0 , w_34809 );
and ( w_34808 , w_34809 , \7026_b0 );
or ( \13588_b1 , \6041_b1 , \7024_b1 );
not ( \7024_b1 , w_34810 );
and ( \13588_b0 , \6041_b0 , w_34811 );
and ( w_34810 , w_34811 , \7024_b0 );
or ( \13589_b1 , \13587_b1 , w_34813 );
not ( w_34813 , w_34814 );
and ( \13589_b0 , \13587_b0 , w_34815 );
and ( w_34814 ,  , w_34815 );
buf ( w_34813 , \13588_b1 );
not ( w_34813 , w_34816 );
not (  , w_34817 );
and ( w_34816 , w_34817 , \13588_b0 );
or ( \13590_b1 , \13589_b1 , w_34818 );
xor ( \13590_b0 , \13589_b0 , w_34820 );
not ( w_34820 , w_34821 );
and ( w_34821 , w_34818 , w_34819 );
buf ( w_34818 , \7032_b1 );
not ( w_34818 , w_34822 );
not ( w_34819 , w_34823 );
and ( w_34822 , w_34823 , \7032_b0 );
or ( \13591_b1 , \6048_b1 , \7043_b1 );
not ( \7043_b1 , w_34824 );
and ( \13591_b0 , \6048_b0 , w_34825 );
and ( w_34824 , w_34825 , \7043_b0 );
or ( \13592_b1 , \6057_b1 , \7041_b1 );
not ( \7041_b1 , w_34826 );
and ( \13592_b0 , \6057_b0 , w_34827 );
and ( w_34826 , w_34827 , \7041_b0 );
or ( \13593_b1 , \13591_b1 , w_34829 );
not ( w_34829 , w_34830 );
and ( \13593_b0 , \13591_b0 , w_34831 );
and ( w_34830 ,  , w_34831 );
buf ( w_34829 , \13592_b1 );
not ( w_34829 , w_34832 );
not (  , w_34833 );
and ( w_34832 , w_34833 , \13592_b0 );
or ( \13594_b1 , \13593_b1 , w_34834 );
xor ( \13594_b0 , \13593_b0 , w_34836 );
not ( w_34836 , w_34837 );
and ( w_34837 , w_34834 , w_34835 );
buf ( w_34834 , \7049_b1 );
not ( w_34834 , w_34838 );
not ( w_34835 , w_34839 );
and ( w_34838 , w_34839 , \7049_b0 );
or ( \13595_b1 , \13590_b1 , \13594_b1 );
xor ( \13595_b0 , \13590_b0 , w_34840 );
not ( w_34840 , w_34841 );
and ( w_34841 , \13594_b1 , \13594_b0 );
or ( \13596_b1 , \6065_b1 , w_34843 );
not ( w_34843 , w_34844 );
and ( \13596_b0 , \6065_b0 , w_34845 );
and ( w_34844 ,  , w_34845 );
buf ( w_34843 , \7059_b1 );
not ( w_34843 , w_34846 );
not (  , w_34847 );
and ( w_34846 , w_34847 , \7059_b0 );
or ( \13597_b1 , \13596_b1 , w_34848 );
xor ( \13597_b0 , \13596_b0 , w_34850 );
not ( w_34850 , w_34851 );
and ( w_34851 , w_34848 , w_34849 );
buf ( w_34848 , \7067_b1 );
not ( w_34848 , w_34852 );
not ( w_34849 , w_34853 );
and ( w_34852 , w_34853 , \7067_b0 );
or ( \13598_b1 , \13595_b1 , \13597_b1 );
xor ( \13598_b0 , \13595_b0 , w_34854 );
not ( w_34854 , w_34855 );
and ( w_34855 , \13597_b1 , \13597_b0 );
or ( \13599_b1 , \13586_b1 , \13598_b1 );
xor ( \13599_b0 , \13586_b0 , w_34856 );
not ( w_34856 , w_34857 );
and ( w_34857 , \13598_b1 , \13598_b0 );
or ( \13600_b1 , \5986_b1 , \6991_b1 );
not ( \6991_b1 , w_34858 );
and ( \13600_b0 , \5986_b0 , w_34859 );
and ( w_34858 , w_34859 , \6991_b0 );
or ( \13601_b1 , \5998_b1 , \6988_b1 );
not ( \6988_b1 , w_34860 );
and ( \13601_b0 , \5998_b0 , w_34861 );
and ( w_34860 , w_34861 , \6988_b0 );
or ( \13602_b1 , \13600_b1 , w_34863 );
not ( w_34863 , w_34864 );
and ( \13602_b0 , \13600_b0 , w_34865 );
and ( w_34864 ,  , w_34865 );
buf ( w_34863 , \13601_b1 );
not ( w_34863 , w_34866 );
not (  , w_34867 );
and ( w_34866 , w_34867 , \13601_b0 );
or ( \13603_b1 , \13602_b1 , w_34868 );
xor ( \13603_b0 , \13602_b0 , w_34870 );
not ( w_34870 , w_34871 );
and ( w_34871 , w_34868 , w_34869 );
buf ( w_34868 , \6985_b1 );
not ( w_34868 , w_34872 );
not ( w_34869 , w_34873 );
and ( w_34872 , w_34873 , \6985_b0 );
or ( \13604_b1 , \7067_b1 , \13603_b1 );
xor ( \13604_b0 , \7067_b0 , w_34874 );
not ( w_34874 , w_34875 );
and ( w_34875 , \13603_b1 , \13603_b0 );
or ( \13605_b1 , \6006_b1 , \7006_b1 );
not ( \7006_b1 , w_34876 );
and ( \13605_b0 , \6006_b0 , w_34877 );
and ( w_34876 , w_34877 , \7006_b0 );
or ( \13606_b1 , \6018_b1 , \7004_b1 );
not ( \7004_b1 , w_34878 );
and ( \13606_b0 , \6018_b0 , w_34879 );
and ( w_34878 , w_34879 , \7004_b0 );
or ( \13607_b1 , \13605_b1 , w_34881 );
not ( w_34881 , w_34882 );
and ( \13607_b0 , \13605_b0 , w_34883 );
and ( w_34882 ,  , w_34883 );
buf ( w_34881 , \13606_b1 );
not ( w_34881 , w_34884 );
not (  , w_34885 );
and ( w_34884 , w_34885 , \13606_b0 );
or ( \13608_b1 , \13607_b1 , w_34886 );
xor ( \13608_b0 , \13607_b0 , w_34888 );
not ( w_34888 , w_34889 );
and ( w_34889 , w_34886 , w_34887 );
buf ( w_34886 , \7012_b1 );
not ( w_34886 , w_34890 );
not ( w_34887 , w_34891 );
and ( w_34890 , w_34891 , \7012_b0 );
or ( \13609_b1 , \13604_b1 , \13608_b1 );
xor ( \13609_b0 , \13604_b0 , w_34892 );
not ( w_34892 , w_34893 );
and ( w_34893 , \13608_b1 , \13608_b0 );
or ( \13610_b1 , \13599_b1 , \13609_b1 );
xor ( \13610_b0 , \13599_b0 , w_34894 );
not ( w_34894 , w_34895 );
and ( w_34895 , \13609_b1 , \13609_b0 );
or ( \13611_b1 , \13582_b1 , \13610_b1 );
xor ( \13611_b0 , \13582_b0 , w_34896 );
not ( w_34896 , w_34897 );
and ( w_34897 , \13610_b1 , \13610_b0 );
or ( \13612_b1 , \13528_b1 , \13553_b1 );
not ( \13553_b1 , w_34898 );
and ( \13612_b0 , \13528_b0 , w_34899 );
and ( w_34898 , w_34899 , \13553_b0 );
or ( \13613_b1 , \13611_b1 , w_34901 );
not ( w_34901 , w_34902 );
and ( \13613_b0 , \13611_b0 , w_34903 );
and ( w_34902 ,  , w_34903 );
buf ( w_34901 , \13612_b1 );
not ( w_34901 , w_34904 );
not (  , w_34905 );
and ( w_34904 , w_34905 , \13612_b0 );
or ( \13614_b1 , \13578_b1 , w_34907 );
not ( w_34907 , w_34908 );
and ( \13614_b0 , \13578_b0 , w_34909 );
and ( w_34908 ,  , w_34909 );
buf ( w_34907 , \13613_b1 );
not ( w_34907 , w_34910 );
not (  , w_34911 );
and ( w_34910 , w_34911 , \13613_b0 );
or ( \13615_b1 , \13586_b1 , \13598_b1 );
not ( \13598_b1 , w_34912 );
and ( \13615_b0 , \13586_b0 , w_34913 );
and ( w_34912 , w_34913 , \13598_b0 );
or ( \13616_b1 , \13598_b1 , \13609_b1 );
not ( \13609_b1 , w_34914 );
and ( \13616_b0 , \13598_b0 , w_34915 );
and ( w_34914 , w_34915 , \13609_b0 );
or ( \13617_b1 , \13586_b1 , \13609_b1 );
not ( \13609_b1 , w_34916 );
and ( \13617_b0 , \13586_b0 , w_34917 );
and ( w_34916 , w_34917 , \13609_b0 );
or ( \13619_b1 , \6065_b1 , \7061_b1 );
not ( \7061_b1 , w_34918 );
and ( \13619_b0 , \6065_b0 , w_34919 );
and ( w_34918 , w_34919 , \7061_b0 );
or ( \13620_b1 , \6048_b1 , \7059_b1 );
not ( \7059_b1 , w_34920 );
and ( \13620_b0 , \6048_b0 , w_34921 );
and ( w_34920 , w_34921 , \7059_b0 );
or ( \13621_b1 , \13619_b1 , w_34923 );
not ( w_34923 , w_34924 );
and ( \13621_b0 , \13619_b0 , w_34925 );
and ( w_34924 ,  , w_34925 );
buf ( w_34923 , \13620_b1 );
not ( w_34923 , w_34926 );
not (  , w_34927 );
and ( w_34926 , w_34927 , \13620_b0 );
or ( \13622_b1 , \13621_b1 , w_34928 );
xor ( \13622_b0 , \13621_b0 , w_34930 );
not ( w_34930 , w_34931 );
and ( w_34931 , w_34928 , w_34929 );
buf ( w_34928 , \7067_b1 );
not ( w_34928 , w_34932 );
not ( w_34929 , w_34933 );
and ( w_34932 , w_34933 , \7067_b0 );
or ( \13623_b1 , \5998_b1 , \6991_b1 );
not ( \6991_b1 , w_34934 );
and ( \13623_b0 , \5998_b0 , w_34935 );
and ( w_34934 , w_34935 , \6991_b0 );
or ( \13624_b1 , \5967_b1 , \6988_b1 );
not ( \6988_b1 , w_34936 );
and ( \13624_b0 , \5967_b0 , w_34937 );
and ( w_34936 , w_34937 , \6988_b0 );
or ( \13625_b1 , \13623_b1 , w_34939 );
not ( w_34939 , w_34940 );
and ( \13625_b0 , \13623_b0 , w_34941 );
and ( w_34940 ,  , w_34941 );
buf ( w_34939 , \13624_b1 );
not ( w_34939 , w_34942 );
not (  , w_34943 );
and ( w_34942 , w_34943 , \13624_b0 );
or ( \13626_b1 , \13625_b1 , w_34944 );
xor ( \13626_b0 , \13625_b0 , w_34946 );
not ( w_34946 , w_34947 );
and ( w_34947 , w_34944 , w_34945 );
buf ( w_34944 , \6985_b1 );
not ( w_34944 , w_34948 );
not ( w_34945 , w_34949 );
and ( w_34948 , w_34949 , \6985_b0 );
or ( \13627_b1 , \6018_b1 , \7006_b1 );
not ( \7006_b1 , w_34950 );
and ( \13627_b0 , \6018_b0 , w_34951 );
and ( w_34950 , w_34951 , \7006_b0 );
or ( \13628_b1 , \5986_b1 , \7004_b1 );
not ( \7004_b1 , w_34952 );
and ( \13628_b0 , \5986_b0 , w_34953 );
and ( w_34952 , w_34953 , \7004_b0 );
or ( \13629_b1 , \13627_b1 , w_34955 );
not ( w_34955 , w_34956 );
and ( \13629_b0 , \13627_b0 , w_34957 );
and ( w_34956 ,  , w_34957 );
buf ( w_34955 , \13628_b1 );
not ( w_34955 , w_34958 );
not (  , w_34959 );
and ( w_34958 , w_34959 , \13628_b0 );
or ( \13630_b1 , \13629_b1 , w_34960 );
xor ( \13630_b0 , \13629_b0 , w_34962 );
not ( w_34962 , w_34963 );
and ( w_34963 , w_34960 , w_34961 );
buf ( w_34960 , \7012_b1 );
not ( w_34960 , w_34964 );
not ( w_34961 , w_34965 );
and ( w_34964 , w_34965 , \7012_b0 );
or ( \13631_b1 , \13626_b1 , \13630_b1 );
xor ( \13631_b0 , \13626_b0 , w_34966 );
not ( w_34966 , w_34967 );
and ( w_34967 , \13630_b1 , \13630_b0 );
or ( \13632_b1 , \6041_b1 , \7026_b1 );
not ( \7026_b1 , w_34968 );
and ( \13632_b0 , \6041_b0 , w_34969 );
and ( w_34968 , w_34969 , \7026_b0 );
or ( \13633_b1 , \6006_b1 , \7024_b1 );
not ( \7024_b1 , w_34970 );
and ( \13633_b0 , \6006_b0 , w_34971 );
and ( w_34970 , w_34971 , \7024_b0 );
or ( \13634_b1 , \13632_b1 , w_34973 );
not ( w_34973 , w_34974 );
and ( \13634_b0 , \13632_b0 , w_34975 );
and ( w_34974 ,  , w_34975 );
buf ( w_34973 , \13633_b1 );
not ( w_34973 , w_34976 );
not (  , w_34977 );
and ( w_34976 , w_34977 , \13633_b0 );
or ( \13635_b1 , \13634_b1 , w_34978 );
xor ( \13635_b0 , \13634_b0 , w_34980 );
not ( w_34980 , w_34981 );
and ( w_34981 , w_34978 , w_34979 );
buf ( w_34978 , \7032_b1 );
not ( w_34978 , w_34982 );
not ( w_34979 , w_34983 );
and ( w_34982 , w_34983 , \7032_b0 );
or ( \13636_b1 , \13631_b1 , \13635_b1 );
xor ( \13636_b0 , \13631_b0 , w_34984 );
not ( w_34984 , w_34985 );
and ( w_34985 , \13635_b1 , \13635_b0 );
or ( \13637_b1 , \13622_b1 , \13636_b1 );
xor ( \13637_b0 , \13622_b0 , w_34986 );
not ( w_34986 , w_34987 );
and ( w_34987 , \13636_b1 , \13636_b0 );
or ( \13638_b1 , \13618_b1 , \13637_b1 );
xor ( \13638_b0 , \13618_b0 , w_34988 );
not ( w_34988 , w_34989 );
and ( w_34989 , \13637_b1 , \13637_b0 );
or ( \13639_b1 , \7067_b1 , \13603_b1 );
not ( \13603_b1 , w_34990 );
and ( \13639_b0 , \7067_b0 , w_34991 );
and ( w_34990 , w_34991 , \13603_b0 );
or ( \13640_b1 , \13603_b1 , \13608_b1 );
not ( \13608_b1 , w_34992 );
and ( \13640_b0 , \13603_b0 , w_34993 );
and ( w_34992 , w_34993 , \13608_b0 );
or ( \13641_b1 , \7067_b1 , \13608_b1 );
not ( \13608_b1 , w_34994 );
and ( \13641_b0 , \7067_b0 , w_34995 );
and ( w_34994 , w_34995 , \13608_b0 );
or ( \13643_b1 , \13590_b1 , \13594_b1 );
not ( \13594_b1 , w_34996 );
and ( \13643_b0 , \13590_b0 , w_34997 );
and ( w_34996 , w_34997 , \13594_b0 );
or ( \13644_b1 , \13594_b1 , \13597_b1 );
not ( \13597_b1 , w_34998 );
and ( \13644_b0 , \13594_b0 , w_34999 );
and ( w_34998 , w_34999 , \13597_b0 );
or ( \13645_b1 , \13590_b1 , \13597_b1 );
not ( \13597_b1 , w_35000 );
and ( \13645_b0 , \13590_b0 , w_35001 );
and ( w_35000 , w_35001 , \13597_b0 );
or ( \13647_b1 , \13642_b1 , \13646_b1 );
xor ( \13647_b0 , \13642_b0 , w_35002 );
not ( w_35002 , w_35003 );
and ( w_35003 , \13646_b1 , \13646_b0 );
or ( \13648_b1 , \6057_b1 , \7043_b1 );
not ( \7043_b1 , w_35004 );
and ( \13648_b0 , \6057_b0 , w_35005 );
and ( w_35004 , w_35005 , \7043_b0 );
or ( \13649_b1 , \6029_b1 , \7041_b1 );
not ( \7041_b1 , w_35006 );
and ( \13649_b0 , \6029_b0 , w_35007 );
and ( w_35006 , w_35007 , \7041_b0 );
or ( \13650_b1 , \13648_b1 , w_35009 );
not ( w_35009 , w_35010 );
and ( \13650_b0 , \13648_b0 , w_35011 );
and ( w_35010 ,  , w_35011 );
buf ( w_35009 , \13649_b1 );
not ( w_35009 , w_35012 );
not (  , w_35013 );
and ( w_35012 , w_35013 , \13649_b0 );
or ( \13651_b1 , \13650_b1 , w_35014 );
xor ( \13651_b0 , \13650_b0 , w_35016 );
not ( w_35016 , w_35017 );
and ( w_35017 , w_35014 , w_35015 );
buf ( w_35014 , \7049_b1 );
not ( w_35014 , w_35018 );
not ( w_35015 , w_35019 );
and ( w_35018 , w_35019 , \7049_b0 );
or ( \13652_b1 , \13647_b1 , \13651_b1 );
xor ( \13652_b0 , \13647_b0 , w_35020 );
not ( w_35020 , w_35021 );
and ( w_35021 , \13651_b1 , \13651_b0 );
or ( \13653_b1 , \13638_b1 , \13652_b1 );
xor ( \13653_b0 , \13638_b0 , w_35022 );
not ( w_35022 , w_35023 );
and ( w_35023 , \13652_b1 , \13652_b0 );
or ( \13654_b1 , \13582_b1 , \13610_b1 );
not ( \13610_b1 , w_35024 );
and ( \13654_b0 , \13582_b0 , w_35025 );
and ( w_35024 , w_35025 , \13610_b0 );
or ( \13655_b1 , \13653_b1 , w_35027 );
not ( w_35027 , w_35028 );
and ( \13655_b0 , \13653_b0 , w_35029 );
and ( w_35028 ,  , w_35029 );
buf ( w_35027 , \13654_b1 );
not ( w_35027 , w_35030 );
not (  , w_35031 );
and ( w_35030 , w_35031 , \13654_b0 );
or ( \13656_b1 , \13626_b1 , \13630_b1 );
not ( \13630_b1 , w_35032 );
and ( \13656_b0 , \13626_b0 , w_35033 );
and ( w_35032 , w_35033 , \13630_b0 );
or ( \13657_b1 , \13630_b1 , \13635_b1 );
not ( \13635_b1 , w_35034 );
and ( \13657_b0 , \13630_b0 , w_35035 );
and ( w_35034 , w_35035 , \13635_b0 );
or ( \13658_b1 , \13626_b1 , \13635_b1 );
not ( \13635_b1 , w_35036 );
and ( \13658_b0 , \13626_b0 , w_35037 );
and ( w_35036 , w_35037 , \13635_b0 );
or ( \13660_b1 , \6065_b1 , w_35039 );
not ( w_35039 , w_35040 );
and ( \13660_b0 , \6065_b0 , w_35041 );
and ( w_35040 ,  , w_35041 );
buf ( w_35039 , \7080_b1 );
not ( w_35039 , w_35042 );
not (  , w_35043 );
and ( w_35042 , w_35043 , \7080_b0 );
or ( \13661_b1 , \13660_b1 , w_35044 );
xor ( \13661_b0 , \13660_b0 , w_35046 );
not ( w_35046 , w_35047 );
and ( w_35047 , w_35044 , w_35045 );
buf ( w_35044 , \7088_b1 );
not ( w_35044 , w_35048 );
not ( w_35045 , w_35049 );
and ( w_35048 , w_35049 , \7088_b0 );
or ( \13662_b1 , \13659_b1 , \13661_b1 );
xor ( \13662_b0 , \13659_b0 , w_35050 );
not ( w_35050 , w_35051 );
and ( w_35051 , \13661_b1 , \13661_b0 );
or ( \13663_b1 , \6006_b1 , \7026_b1 );
not ( \7026_b1 , w_35052 );
and ( \13663_b0 , \6006_b0 , w_35053 );
and ( w_35052 , w_35053 , \7026_b0 );
or ( \13664_b1 , \6018_b1 , \7024_b1 );
not ( \7024_b1 , w_35054 );
and ( \13664_b0 , \6018_b0 , w_35055 );
and ( w_35054 , w_35055 , \7024_b0 );
or ( \13665_b1 , \13663_b1 , w_35057 );
not ( w_35057 , w_35058 );
and ( \13665_b0 , \13663_b0 , w_35059 );
and ( w_35058 ,  , w_35059 );
buf ( w_35057 , \13664_b1 );
not ( w_35057 , w_35060 );
not (  , w_35061 );
and ( w_35060 , w_35061 , \13664_b0 );
or ( \13666_b1 , \13665_b1 , w_35062 );
xor ( \13666_b0 , \13665_b0 , w_35064 );
not ( w_35064 , w_35065 );
and ( w_35065 , w_35062 , w_35063 );
buf ( w_35062 , \7032_b1 );
not ( w_35062 , w_35066 );
not ( w_35063 , w_35067 );
and ( w_35066 , w_35067 , \7032_b0 );
or ( \13667_b1 , \6029_b1 , \7043_b1 );
not ( \7043_b1 , w_35068 );
and ( \13667_b0 , \6029_b0 , w_35069 );
and ( w_35068 , w_35069 , \7043_b0 );
or ( \13668_b1 , \6041_b1 , \7041_b1 );
not ( \7041_b1 , w_35070 );
and ( \13668_b0 , \6041_b0 , w_35071 );
and ( w_35070 , w_35071 , \7041_b0 );
or ( \13669_b1 , \13667_b1 , w_35073 );
not ( w_35073 , w_35074 );
and ( \13669_b0 , \13667_b0 , w_35075 );
and ( w_35074 ,  , w_35075 );
buf ( w_35073 , \13668_b1 );
not ( w_35073 , w_35076 );
not (  , w_35077 );
and ( w_35076 , w_35077 , \13668_b0 );
or ( \13670_b1 , \13669_b1 , w_35078 );
xor ( \13670_b0 , \13669_b0 , w_35080 );
not ( w_35080 , w_35081 );
and ( w_35081 , w_35078 , w_35079 );
buf ( w_35078 , \7049_b1 );
not ( w_35078 , w_35082 );
not ( w_35079 , w_35083 );
and ( w_35082 , w_35083 , \7049_b0 );
or ( \13671_b1 , \13666_b1 , \13670_b1 );
xor ( \13671_b0 , \13666_b0 , w_35084 );
not ( w_35084 , w_35085 );
and ( w_35085 , \13670_b1 , \13670_b0 );
or ( \13672_b1 , \6048_b1 , \7061_b1 );
not ( \7061_b1 , w_35086 );
and ( \13672_b0 , \6048_b0 , w_35087 );
and ( w_35086 , w_35087 , \7061_b0 );
or ( \13673_b1 , \6057_b1 , \7059_b1 );
not ( \7059_b1 , w_35088 );
and ( \13673_b0 , \6057_b0 , w_35089 );
and ( w_35088 , w_35089 , \7059_b0 );
or ( \13674_b1 , \13672_b1 , w_35091 );
not ( w_35091 , w_35092 );
and ( \13674_b0 , \13672_b0 , w_35093 );
and ( w_35092 ,  , w_35093 );
buf ( w_35091 , \13673_b1 );
not ( w_35091 , w_35094 );
not (  , w_35095 );
and ( w_35094 , w_35095 , \13673_b0 );
or ( \13675_b1 , \13674_b1 , w_35096 );
xor ( \13675_b0 , \13674_b0 , w_35098 );
not ( w_35098 , w_35099 );
and ( w_35099 , w_35096 , w_35097 );
buf ( w_35096 , \7067_b1 );
not ( w_35096 , w_35100 );
not ( w_35097 , w_35101 );
and ( w_35100 , w_35101 , \7067_b0 );
or ( \13676_b1 , \13671_b1 , \13675_b1 );
xor ( \13676_b0 , \13671_b0 , w_35102 );
not ( w_35102 , w_35103 );
and ( w_35103 , \13675_b1 , \13675_b0 );
or ( \13677_b1 , \13662_b1 , \13676_b1 );
xor ( \13677_b0 , \13662_b0 , w_35104 );
not ( w_35104 , w_35105 );
and ( w_35105 , \13676_b1 , \13676_b0 );
or ( \13678_b1 , \13642_b1 , \13646_b1 );
not ( \13646_b1 , w_35106 );
and ( \13678_b0 , \13642_b0 , w_35107 );
and ( w_35106 , w_35107 , \13646_b0 );
or ( \13679_b1 , \13646_b1 , \13651_b1 );
not ( \13651_b1 , w_35108 );
and ( \13679_b0 , \13646_b0 , w_35109 );
and ( w_35108 , w_35109 , \13651_b0 );
or ( \13680_b1 , \13642_b1 , \13651_b1 );
not ( \13651_b1 , w_35110 );
and ( \13680_b0 , \13642_b0 , w_35111 );
and ( w_35110 , w_35111 , \13651_b0 );
or ( \13682_b1 , \13622_b1 , \13636_b1 );
not ( \13636_b1 , w_35112 );
and ( \13682_b0 , \13622_b0 , w_35113 );
and ( w_35112 , w_35113 , \13636_b0 );
or ( \13683_b1 , \13681_b1 , \13682_b1 );
xor ( \13683_b0 , \13681_b0 , w_35114 );
not ( w_35114 , w_35115 );
and ( w_35115 , \13682_b1 , \13682_b0 );
or ( \13684_b1 , \5967_b1 , \6991_b1 );
not ( \6991_b1 , w_35116 );
and ( \13684_b0 , \5967_b0 , w_35117 );
and ( w_35116 , w_35117 , \6991_b0 );
or ( \13685_b1 , \5979_b1 , \6988_b1 );
not ( \6988_b1 , w_35118 );
and ( \13685_b0 , \5979_b0 , w_35119 );
and ( w_35118 , w_35119 , \6988_b0 );
or ( \13686_b1 , \13684_b1 , w_35121 );
not ( w_35121 , w_35122 );
and ( \13686_b0 , \13684_b0 , w_35123 );
and ( w_35122 ,  , w_35123 );
buf ( w_35121 , \13685_b1 );
not ( w_35121 , w_35124 );
not (  , w_35125 );
and ( w_35124 , w_35125 , \13685_b0 );
or ( \13687_b1 , \13686_b1 , w_35126 );
xor ( \13687_b0 , \13686_b0 , w_35128 );
not ( w_35128 , w_35129 );
and ( w_35129 , w_35126 , w_35127 );
buf ( w_35126 , \6985_b1 );
not ( w_35126 , w_35130 );
not ( w_35127 , w_35131 );
and ( w_35130 , w_35131 , \6985_b0 );
or ( \13688_b1 , \7088_b1 , \13687_b1 );
xor ( \13688_b0 , \7088_b0 , w_35132 );
not ( w_35132 , w_35133 );
and ( w_35133 , \13687_b1 , \13687_b0 );
or ( \13689_b1 , \5986_b1 , \7006_b1 );
not ( \7006_b1 , w_35134 );
and ( \13689_b0 , \5986_b0 , w_35135 );
and ( w_35134 , w_35135 , \7006_b0 );
or ( \13690_b1 , \5998_b1 , \7004_b1 );
not ( \7004_b1 , w_35136 );
and ( \13690_b0 , \5998_b0 , w_35137 );
and ( w_35136 , w_35137 , \7004_b0 );
or ( \13691_b1 , \13689_b1 , w_35139 );
not ( w_35139 , w_35140 );
and ( \13691_b0 , \13689_b0 , w_35141 );
and ( w_35140 ,  , w_35141 );
buf ( w_35139 , \13690_b1 );
not ( w_35139 , w_35142 );
not (  , w_35143 );
and ( w_35142 , w_35143 , \13690_b0 );
or ( \13692_b1 , \13691_b1 , w_35144 );
xor ( \13692_b0 , \13691_b0 , w_35146 );
not ( w_35146 , w_35147 );
and ( w_35147 , w_35144 , w_35145 );
buf ( w_35144 , \7012_b1 );
not ( w_35144 , w_35148 );
not ( w_35145 , w_35149 );
and ( w_35148 , w_35149 , \7012_b0 );
or ( \13693_b1 , \13688_b1 , \13692_b1 );
xor ( \13693_b0 , \13688_b0 , w_35150 );
not ( w_35150 , w_35151 );
and ( w_35151 , \13692_b1 , \13692_b0 );
or ( \13694_b1 , \13683_b1 , \13693_b1 );
xor ( \13694_b0 , \13683_b0 , w_35152 );
not ( w_35152 , w_35153 );
and ( w_35153 , \13693_b1 , \13693_b0 );
or ( \13695_b1 , \13677_b1 , \13694_b1 );
xor ( \13695_b0 , \13677_b0 , w_35154 );
not ( w_35154 , w_35155 );
and ( w_35155 , \13694_b1 , \13694_b0 );
or ( \13696_b1 , \13618_b1 , \13637_b1 );
not ( \13637_b1 , w_35156 );
and ( \13696_b0 , \13618_b0 , w_35157 );
and ( w_35156 , w_35157 , \13637_b0 );
or ( \13697_b1 , \13637_b1 , \13652_b1 );
not ( \13652_b1 , w_35158 );
and ( \13697_b0 , \13637_b0 , w_35159 );
and ( w_35158 , w_35159 , \13652_b0 );
or ( \13698_b1 , \13618_b1 , \13652_b1 );
not ( \13652_b1 , w_35160 );
and ( \13698_b0 , \13618_b0 , w_35161 );
and ( w_35160 , w_35161 , \13652_b0 );
or ( \13700_b1 , \13695_b1 , w_35163 );
not ( w_35163 , w_35164 );
and ( \13700_b0 , \13695_b0 , w_35165 );
and ( w_35164 ,  , w_35165 );
buf ( w_35163 , \13699_b1 );
not ( w_35163 , w_35166 );
not (  , w_35167 );
and ( w_35166 , w_35167 , \13699_b0 );
or ( \13701_b1 , \13655_b1 , w_35169 );
not ( w_35169 , w_35170 );
and ( \13701_b0 , \13655_b0 , w_35171 );
and ( w_35170 ,  , w_35171 );
buf ( w_35169 , \13700_b1 );
not ( w_35169 , w_35172 );
not (  , w_35173 );
and ( w_35172 , w_35173 , \13700_b0 );
or ( \13702_b1 , \13614_b1 , w_35175 );
not ( w_35175 , w_35176 );
and ( \13702_b0 , \13614_b0 , w_35177 );
and ( w_35176 ,  , w_35177 );
buf ( w_35175 , \13701_b1 );
not ( w_35175 , w_35178 );
not (  , w_35179 );
and ( w_35178 , w_35179 , \13701_b0 );
or ( \13703_b1 , \13681_b1 , \13682_b1 );
not ( \13682_b1 , w_35180 );
and ( \13703_b0 , \13681_b0 , w_35181 );
and ( w_35180 , w_35181 , \13682_b0 );
or ( \13704_b1 , \13682_b1 , \13693_b1 );
not ( \13693_b1 , w_35182 );
and ( \13704_b0 , \13682_b0 , w_35183 );
and ( w_35182 , w_35183 , \13693_b0 );
or ( \13705_b1 , \13681_b1 , \13693_b1 );
not ( \13693_b1 , w_35184 );
and ( \13705_b0 , \13681_b0 , w_35185 );
and ( w_35184 , w_35185 , \13693_b0 );
or ( \13707_b1 , \13659_b1 , \13661_b1 );
not ( \13661_b1 , w_35186 );
and ( \13707_b0 , \13659_b0 , w_35187 );
and ( w_35186 , w_35187 , \13661_b0 );
or ( \13708_b1 , \13661_b1 , \13676_b1 );
not ( \13676_b1 , w_35188 );
and ( \13708_b0 , \13661_b0 , w_35189 );
and ( w_35188 , w_35189 , \13676_b0 );
or ( \13709_b1 , \13659_b1 , \13676_b1 );
not ( \13676_b1 , w_35190 );
and ( \13709_b0 , \13659_b0 , w_35191 );
and ( w_35190 , w_35191 , \13676_b0 );
or ( \13711_b1 , \12379_b1 , \12383_b1 );
xor ( \13711_b0 , \12379_b0 , w_35192 );
not ( w_35192 , w_35193 );
and ( w_35193 , \12383_b1 , \12383_b0 );
or ( \13712_b1 , \13711_b1 , \12388_b1 );
xor ( \13712_b0 , \13711_b0 , w_35194 );
not ( w_35194 , w_35195 );
and ( w_35195 , \12388_b1 , \12388_b0 );
or ( \13713_b1 , \13710_b1 , \13712_b1 );
xor ( \13713_b0 , \13710_b0 , w_35196 );
not ( w_35196 , w_35197 );
and ( w_35197 , \13712_b1 , \13712_b0 );
or ( \13714_b1 , \7088_b1 , \13687_b1 );
not ( \13687_b1 , w_35198 );
and ( \13714_b0 , \7088_b0 , w_35199 );
and ( w_35198 , w_35199 , \13687_b0 );
or ( \13715_b1 , \13687_b1 , \13692_b1 );
not ( \13692_b1 , w_35200 );
and ( \13715_b0 , \13687_b0 , w_35201 );
and ( w_35200 , w_35201 , \13692_b0 );
or ( \13716_b1 , \7088_b1 , \13692_b1 );
not ( \13692_b1 , w_35202 );
and ( \13716_b0 , \7088_b0 , w_35203 );
and ( w_35202 , w_35203 , \13692_b0 );
or ( \13718_b1 , \13666_b1 , \13670_b1 );
not ( \13670_b1 , w_35204 );
and ( \13718_b0 , \13666_b0 , w_35205 );
and ( w_35204 , w_35205 , \13670_b0 );
or ( \13719_b1 , \13670_b1 , \13675_b1 );
not ( \13675_b1 , w_35206 );
and ( \13719_b0 , \13670_b0 , w_35207 );
and ( w_35206 , w_35207 , \13675_b0 );
or ( \13720_b1 , \13666_b1 , \13675_b1 );
not ( \13675_b1 , w_35208 );
and ( \13720_b0 , \13666_b0 , w_35209 );
and ( w_35208 , w_35209 , \13675_b0 );
or ( \13722_b1 , \13717_b1 , \13721_b1 );
xor ( \13722_b0 , \13717_b0 , w_35210 );
not ( w_35210 , w_35211 );
and ( w_35211 , \13721_b1 , \13721_b0 );
or ( \13723_b1 , \12395_b1 , \12399_b1 );
xor ( \13723_b0 , \12395_b0 , w_35212 );
not ( w_35212 , w_35213 );
and ( w_35213 , \12399_b1 , \12399_b0 );
or ( \13724_b1 , \13723_b1 , \12404_b1 );
xor ( \13724_b0 , \13723_b0 , w_35214 );
not ( w_35214 , w_35215 );
and ( w_35215 , \12404_b1 , \12404_b0 );
or ( \13725_b1 , \13722_b1 , \13724_b1 );
xor ( \13725_b0 , \13722_b0 , w_35216 );
not ( w_35216 , w_35217 );
and ( w_35217 , \13724_b1 , \13724_b0 );
or ( \13726_b1 , \13713_b1 , \13725_b1 );
xor ( \13726_b0 , \13713_b0 , w_35218 );
not ( w_35218 , w_35219 );
and ( w_35219 , \13725_b1 , \13725_b0 );
or ( \13727_b1 , \13706_b1 , \13726_b1 );
xor ( \13727_b0 , \13706_b0 , w_35220 );
not ( w_35220 , w_35221 );
and ( w_35221 , \13726_b1 , \13726_b0 );
or ( \13728_b1 , \13677_b1 , \13694_b1 );
not ( \13694_b1 , w_35222 );
and ( \13728_b0 , \13677_b0 , w_35223 );
and ( w_35222 , w_35223 , \13694_b0 );
or ( \13729_b1 , \13727_b1 , w_35225 );
not ( w_35225 , w_35226 );
and ( \13729_b0 , \13727_b0 , w_35227 );
and ( w_35226 ,  , w_35227 );
buf ( w_35225 , \13728_b1 );
not ( w_35225 , w_35228 );
not (  , w_35229 );
and ( w_35228 , w_35229 , \13728_b0 );
or ( \13730_b1 , \13710_b1 , \13712_b1 );
not ( \13712_b1 , w_35230 );
and ( \13730_b0 , \13710_b0 , w_35231 );
and ( w_35230 , w_35231 , \13712_b0 );
or ( \13731_b1 , \13712_b1 , \13725_b1 );
not ( \13725_b1 , w_35232 );
and ( \13731_b0 , \13712_b0 , w_35233 );
and ( w_35232 , w_35233 , \13725_b0 );
or ( \13732_b1 , \13710_b1 , \13725_b1 );
not ( \13725_b1 , w_35234 );
and ( \13732_b0 , \13710_b0 , w_35235 );
and ( w_35234 , w_35235 , \13725_b0 );
or ( \13734_b1 , \13717_b1 , \13721_b1 );
not ( \13721_b1 , w_35236 );
and ( \13734_b0 , \13717_b0 , w_35237 );
and ( w_35236 , w_35237 , \13721_b0 );
or ( \13735_b1 , \13721_b1 , \13724_b1 );
not ( \13724_b1 , w_35238 );
and ( \13735_b0 , \13721_b0 , w_35239 );
and ( w_35238 , w_35239 , \13724_b0 );
or ( \13736_b1 , \13717_b1 , \13724_b1 );
not ( \13724_b1 , w_35240 );
and ( \13736_b0 , \13717_b0 , w_35241 );
and ( w_35240 , w_35241 , \13724_b0 );
or ( \13738_b1 , \12417_b1 , \12419_b1 );
xor ( \13738_b0 , \12417_b0 , w_35242 );
not ( w_35242 , w_35243 );
and ( w_35243 , \12419_b1 , \12419_b0 );
or ( \13739_b1 , \13738_b1 , \12422_b1 );
xor ( \13739_b0 , \13738_b0 , w_35244 );
not ( w_35244 , w_35245 );
and ( w_35245 , \12422_b1 , \12422_b0 );
or ( \13740_b1 , \13737_b1 , \13739_b1 );
xor ( \13740_b0 , \13737_b0 , w_35246 );
not ( w_35246 , w_35247 );
and ( w_35247 , \13739_b1 , \13739_b0 );
or ( \13741_b1 , \12391_b1 , \12407_b1 );
xor ( \13741_b0 , \12391_b0 , w_35248 );
not ( w_35248 , w_35249 );
and ( w_35249 , \12407_b1 , \12407_b0 );
or ( \13742_b1 , \13741_b1 , \12412_b1 );
xor ( \13742_b0 , \13741_b0 , w_35250 );
not ( w_35250 , w_35251 );
and ( w_35251 , \12412_b1 , \12412_b0 );
or ( \13743_b1 , \13740_b1 , \13742_b1 );
xor ( \13743_b0 , \13740_b0 , w_35252 );
not ( w_35252 , w_35253 );
and ( w_35253 , \13742_b1 , \13742_b0 );
or ( \13744_b1 , \13733_b1 , \13743_b1 );
xor ( \13744_b0 , \13733_b0 , w_35254 );
not ( w_35254 , w_35255 );
and ( w_35255 , \13743_b1 , \13743_b0 );
or ( \13745_b1 , \13706_b1 , \13726_b1 );
not ( \13726_b1 , w_35256 );
and ( \13745_b0 , \13706_b0 , w_35257 );
and ( w_35256 , w_35257 , \13726_b0 );
or ( \13746_b1 , \13744_b1 , w_35259 );
not ( w_35259 , w_35260 );
and ( \13746_b0 , \13744_b0 , w_35261 );
and ( w_35260 ,  , w_35261 );
buf ( w_35259 , \13745_b1 );
not ( w_35259 , w_35262 );
not (  , w_35263 );
and ( w_35262 , w_35263 , \13745_b0 );
or ( \13747_b1 , \13729_b1 , w_35265 );
not ( w_35265 , w_35266 );
and ( \13747_b0 , \13729_b0 , w_35267 );
and ( w_35266 ,  , w_35267 );
buf ( w_35265 , \13746_b1 );
not ( w_35265 , w_35268 );
not (  , w_35269 );
and ( w_35268 , w_35269 , \13746_b0 );
or ( \13748_b1 , \13737_b1 , \13739_b1 );
not ( \13739_b1 , w_35270 );
and ( \13748_b0 , \13737_b0 , w_35271 );
and ( w_35270 , w_35271 , \13739_b0 );
or ( \13749_b1 , \13739_b1 , \13742_b1 );
not ( \13742_b1 , w_35272 );
and ( \13749_b0 , \13739_b0 , w_35273 );
and ( w_35272 , w_35273 , \13742_b0 );
or ( \13750_b1 , \13737_b1 , \13742_b1 );
not ( \13742_b1 , w_35274 );
and ( \13750_b0 , \13737_b0 , w_35275 );
and ( w_35274 , w_35275 , \13742_b0 );
or ( \13752_b1 , \12433_b1 , \12435_b1 );
xor ( \13752_b0 , \12433_b0 , w_35276 );
not ( w_35276 , w_35277 );
and ( w_35277 , \12435_b1 , \12435_b0 );
or ( \13753_b1 , \13751_b1 , \13752_b1 );
xor ( \13753_b0 , \13751_b0 , w_35278 );
not ( w_35278 , w_35279 );
and ( w_35279 , \13752_b1 , \13752_b0 );
or ( \13754_b1 , \12415_b1 , \12425_b1 );
xor ( \13754_b0 , \12415_b0 , w_35280 );
not ( w_35280 , w_35281 );
and ( w_35281 , \12425_b1 , \12425_b0 );
or ( \13755_b1 , \13754_b1 , \12428_b1 );
xor ( \13755_b0 , \13754_b0 , w_35282 );
not ( w_35282 , w_35283 );
and ( w_35283 , \12428_b1 , \12428_b0 );
or ( \13756_b1 , \13753_b1 , \13755_b1 );
xor ( \13756_b0 , \13753_b0 , w_35284 );
not ( w_35284 , w_35285 );
and ( w_35285 , \13755_b1 , \13755_b0 );
or ( \13757_b1 , \13733_b1 , \13743_b1 );
not ( \13743_b1 , w_35286 );
and ( \13757_b0 , \13733_b0 , w_35287 );
and ( w_35286 , w_35287 , \13743_b0 );
or ( \13758_b1 , \13756_b1 , w_35289 );
not ( w_35289 , w_35290 );
and ( \13758_b0 , \13756_b0 , w_35291 );
and ( w_35290 ,  , w_35291 );
buf ( w_35289 , \13757_b1 );
not ( w_35289 , w_35292 );
not (  , w_35293 );
and ( w_35292 , w_35293 , \13757_b0 );
or ( \13759_b1 , \12431_b1 , \12436_b1 );
xor ( \13759_b0 , \12431_b0 , w_35294 );
not ( w_35294 , w_35295 );
and ( w_35295 , \12436_b1 , \12436_b0 );
or ( \13760_b1 , \13759_b1 , \12439_b1 );
xor ( \13760_b0 , \13759_b0 , w_35296 );
not ( w_35296 , w_35297 );
and ( w_35297 , \12439_b1 , \12439_b0 );
or ( \13761_b1 , \13751_b1 , \13752_b1 );
not ( \13752_b1 , w_35298 );
and ( \13761_b0 , \13751_b0 , w_35299 );
and ( w_35298 , w_35299 , \13752_b0 );
or ( \13762_b1 , \13752_b1 , \13755_b1 );
not ( \13755_b1 , w_35300 );
and ( \13762_b0 , \13752_b0 , w_35301 );
and ( w_35300 , w_35301 , \13755_b0 );
or ( \13763_b1 , \13751_b1 , \13755_b1 );
not ( \13755_b1 , w_35302 );
and ( \13763_b0 , \13751_b0 , w_35303 );
and ( w_35302 , w_35303 , \13755_b0 );
or ( \13765_b1 , \13760_b1 , w_35305 );
not ( w_35305 , w_35306 );
and ( \13765_b0 , \13760_b0 , w_35307 );
and ( w_35306 ,  , w_35307 );
buf ( w_35305 , \13764_b1 );
not ( w_35305 , w_35308 );
not (  , w_35309 );
and ( w_35308 , w_35309 , \13764_b0 );
or ( \13766_b1 , \13758_b1 , w_35311 );
not ( w_35311 , w_35312 );
and ( \13766_b0 , \13758_b0 , w_35313 );
and ( w_35312 ,  , w_35313 );
buf ( w_35311 , \13765_b1 );
not ( w_35311 , w_35314 );
not (  , w_35315 );
and ( w_35314 , w_35315 , \13765_b0 );
or ( \13767_b1 , \13747_b1 , w_35317 );
not ( w_35317 , w_35318 );
and ( \13767_b0 , \13747_b0 , w_35319 );
and ( w_35318 ,  , w_35319 );
buf ( w_35317 , \13766_b1 );
not ( w_35317 , w_35320 );
not (  , w_35321 );
and ( w_35320 , w_35321 , \13766_b0 );
or ( \13768_b1 , \13702_b1 , w_35323 );
not ( w_35323 , w_35324 );
and ( \13768_b0 , \13702_b0 , w_35325 );
and ( w_35324 ,  , w_35325 );
buf ( w_35323 , \13767_b1 );
not ( w_35323 , w_35326 );
not (  , w_35327 );
and ( w_35326 , w_35327 , \13767_b0 );
or ( \13769_b1 , \6057_b1 , \6991_b1 );
not ( \6991_b1 , w_35328 );
and ( \13769_b0 , \6057_b0 , w_35329 );
and ( w_35328 , w_35329 , \6991_b0 );
or ( \13770_b1 , \6029_b1 , \6988_b1 );
not ( \6988_b1 , w_35330 );
and ( \13770_b0 , \6029_b0 , w_35331 );
and ( w_35330 , w_35331 , \6988_b0 );
or ( \13771_b1 , \13769_b1 , w_35333 );
not ( w_35333 , w_35334 );
and ( \13771_b0 , \13769_b0 , w_35335 );
and ( w_35334 ,  , w_35335 );
buf ( w_35333 , \13770_b1 );
not ( w_35333 , w_35336 );
not (  , w_35337 );
and ( w_35336 , w_35337 , \13770_b0 );
or ( \13772_b1 , \13771_b1 , w_35338 );
xor ( \13772_b0 , \13771_b0 , w_35340 );
not ( w_35340 , w_35341 );
and ( w_35341 , w_35338 , w_35339 );
buf ( w_35338 , \6985_b1 );
not ( w_35338 , w_35342 );
not ( w_35339 , w_35343 );
and ( w_35342 , w_35343 , \6985_b0 );
or ( \13773_b1 , \6065_b1 , \7006_b1 );
not ( \7006_b1 , w_35344 );
and ( \13773_b0 , \6065_b0 , w_35345 );
and ( w_35344 , w_35345 , \7006_b0 );
or ( \13774_b1 , \6048_b1 , \7004_b1 );
not ( \7004_b1 , w_35346 );
and ( \13774_b0 , \6048_b0 , w_35347 );
and ( w_35346 , w_35347 , \7004_b0 );
or ( \13775_b1 , \13773_b1 , w_35349 );
not ( w_35349 , w_35350 );
and ( \13775_b0 , \13773_b0 , w_35351 );
and ( w_35350 ,  , w_35351 );
buf ( w_35349 , \13774_b1 );
not ( w_35349 , w_35352 );
not (  , w_35353 );
and ( w_35352 , w_35353 , \13774_b0 );
or ( \13776_b1 , \13775_b1 , w_35354 );
xor ( \13776_b0 , \13775_b0 , w_35356 );
not ( w_35356 , w_35357 );
and ( w_35357 , w_35354 , w_35355 );
buf ( w_35354 , \7012_b1 );
not ( w_35354 , w_35358 );
not ( w_35355 , w_35359 );
and ( w_35358 , w_35359 , \7012_b0 );
or ( \13777_b1 , \13772_b1 , \13776_b1 );
xor ( \13777_b0 , \13772_b0 , w_35360 );
not ( w_35360 , w_35361 );
and ( w_35361 , \13776_b1 , \13776_b0 );
or ( \13778_b1 , \6048_b1 , \6991_b1 );
not ( \6991_b1 , w_35362 );
and ( \13778_b0 , \6048_b0 , w_35363 );
and ( w_35362 , w_35363 , \6991_b0 );
or ( \13779_b1 , \6057_b1 , \6988_b1 );
not ( \6988_b1 , w_35364 );
and ( \13779_b0 , \6057_b0 , w_35365 );
and ( w_35364 , w_35365 , \6988_b0 );
or ( \13780_b1 , \13778_b1 , w_35367 );
not ( w_35367 , w_35368 );
and ( \13780_b0 , \13778_b0 , w_35369 );
and ( w_35368 ,  , w_35369 );
buf ( w_35367 , \13779_b1 );
not ( w_35367 , w_35370 );
not (  , w_35371 );
and ( w_35370 , w_35371 , \13779_b0 );
or ( \13781_b1 , \13780_b1 , w_35372 );
xor ( \13781_b0 , \13780_b0 , w_35374 );
not ( w_35374 , w_35375 );
and ( w_35375 , w_35372 , w_35373 );
buf ( w_35372 , \6985_b1 );
not ( w_35372 , w_35376 );
not ( w_35373 , w_35377 );
and ( w_35376 , w_35377 , \6985_b0 );
or ( \13782_b1 , \13781_b1 , \7012_b1 );
not ( \7012_b1 , w_35378 );
and ( \13782_b0 , \13781_b0 , w_35379 );
and ( w_35378 , w_35379 , \7012_b0 );
or ( \13783_b1 , \13777_b1 , w_35381 );
not ( w_35381 , w_35382 );
and ( \13783_b0 , \13777_b0 , w_35383 );
and ( w_35382 ,  , w_35383 );
buf ( w_35381 , \13782_b1 );
not ( w_35381 , w_35384 );
not (  , w_35385 );
and ( w_35384 , w_35385 , \13782_b0 );
or ( \13784_b1 , \6065_b1 , w_35387 );
not ( w_35387 , w_35388 );
and ( \13784_b0 , \6065_b0 , w_35389 );
and ( w_35388 ,  , w_35389 );
buf ( w_35387 , \7024_b1 );
not ( w_35387 , w_35390 );
not (  , w_35391 );
and ( w_35390 , w_35391 , \7024_b0 );
or ( \13785_b1 , \13784_b1 , w_35392 );
xor ( \13785_b0 , \13784_b0 , w_35394 );
not ( w_35394 , w_35395 );
and ( w_35395 , w_35392 , w_35393 );
buf ( w_35392 , \7032_b1 );
not ( w_35392 , w_35396 );
not ( w_35393 , w_35397 );
and ( w_35396 , w_35397 , \7032_b0 );
or ( \13786_b1 , \6029_b1 , \6991_b1 );
not ( \6991_b1 , w_35398 );
and ( \13786_b0 , \6029_b0 , w_35399 );
and ( w_35398 , w_35399 , \6991_b0 );
or ( \13787_b1 , \6041_b1 , \6988_b1 );
not ( \6988_b1 , w_35400 );
and ( \13787_b0 , \6041_b0 , w_35401 );
and ( w_35400 , w_35401 , \6988_b0 );
or ( \13788_b1 , \13786_b1 , w_35403 );
not ( w_35403 , w_35404 );
and ( \13788_b0 , \13786_b0 , w_35405 );
and ( w_35404 ,  , w_35405 );
buf ( w_35403 , \13787_b1 );
not ( w_35403 , w_35406 );
not (  , w_35407 );
and ( w_35406 , w_35407 , \13787_b0 );
or ( \13789_b1 , \13788_b1 , w_35408 );
xor ( \13789_b0 , \13788_b0 , w_35410 );
not ( w_35410 , w_35411 );
and ( w_35411 , w_35408 , w_35409 );
buf ( w_35408 , \6985_b1 );
not ( w_35408 , w_35412 );
not ( w_35409 , w_35413 );
and ( w_35412 , w_35413 , \6985_b0 );
or ( \13790_b1 , \7032_b1 , \13789_b1 );
xor ( \13790_b0 , \7032_b0 , w_35414 );
not ( w_35414 , w_35415 );
and ( w_35415 , \13789_b1 , \13789_b0 );
or ( \13791_b1 , \6048_b1 , \7006_b1 );
not ( \7006_b1 , w_35416 );
and ( \13791_b0 , \6048_b0 , w_35417 );
and ( w_35416 , w_35417 , \7006_b0 );
or ( \13792_b1 , \6057_b1 , \7004_b1 );
not ( \7004_b1 , w_35418 );
and ( \13792_b0 , \6057_b0 , w_35419 );
and ( w_35418 , w_35419 , \7004_b0 );
or ( \13793_b1 , \13791_b1 , w_35421 );
not ( w_35421 , w_35422 );
and ( \13793_b0 , \13791_b0 , w_35423 );
and ( w_35422 ,  , w_35423 );
buf ( w_35421 , \13792_b1 );
not ( w_35421 , w_35424 );
not (  , w_35425 );
and ( w_35424 , w_35425 , \13792_b0 );
or ( \13794_b1 , \13793_b1 , w_35426 );
xor ( \13794_b0 , \13793_b0 , w_35428 );
not ( w_35428 , w_35429 );
and ( w_35429 , w_35426 , w_35427 );
buf ( w_35426 , \7012_b1 );
not ( w_35426 , w_35430 );
not ( w_35427 , w_35431 );
and ( w_35430 , w_35431 , \7012_b0 );
or ( \13795_b1 , \13790_b1 , \13794_b1 );
xor ( \13795_b0 , \13790_b0 , w_35432 );
not ( w_35432 , w_35433 );
and ( w_35433 , \13794_b1 , \13794_b0 );
or ( \13796_b1 , \13785_b1 , \13795_b1 );
xor ( \13796_b0 , \13785_b0 , w_35434 );
not ( w_35434 , w_35435 );
and ( w_35435 , \13795_b1 , \13795_b0 );
or ( \13797_b1 , \13772_b1 , \13776_b1 );
not ( \13776_b1 , w_35436 );
and ( \13797_b0 , \13772_b0 , w_35437 );
and ( w_35436 , w_35437 , \13776_b0 );
or ( \13798_b1 , \13796_b1 , w_35439 );
not ( w_35439 , w_35440 );
and ( \13798_b0 , \13796_b0 , w_35441 );
and ( w_35440 ,  , w_35441 );
buf ( w_35439 , \13797_b1 );
not ( w_35439 , w_35442 );
not (  , w_35443 );
and ( w_35442 , w_35443 , \13797_b0 );
or ( \13799_b1 , \13783_b1 , w_35445 );
not ( w_35445 , w_35446 );
and ( \13799_b0 , \13783_b0 , w_35447 );
and ( w_35446 ,  , w_35447 );
buf ( w_35445 , \13798_b1 );
not ( w_35445 , w_35448 );
not (  , w_35449 );
and ( w_35448 , w_35449 , \13798_b0 );
or ( \13800_b1 , \7032_b1 , \13789_b1 );
not ( \13789_b1 , w_35450 );
and ( \13800_b0 , \7032_b0 , w_35451 );
and ( w_35450 , w_35451 , \13789_b0 );
or ( \13801_b1 , \13789_b1 , \13794_b1 );
not ( \13794_b1 , w_35452 );
and ( \13801_b0 , \13789_b0 , w_35453 );
and ( w_35452 , w_35453 , \13794_b0 );
or ( \13802_b1 , \7032_b1 , \13794_b1 );
not ( \13794_b1 , w_35454 );
and ( \13802_b0 , \7032_b0 , w_35455 );
and ( w_35454 , w_35455 , \13794_b0 );
or ( \13804_b1 , \13558_b1 , \13562_b1 );
xor ( \13804_b0 , \13558_b0 , w_35456 );
not ( w_35456 , w_35457 );
and ( w_35457 , \13562_b1 , \13562_b0 );
or ( \13805_b1 , \13804_b1 , \13567_b1 );
xor ( \13805_b0 , \13804_b0 , w_35458 );
not ( w_35458 , w_35459 );
and ( w_35459 , \13567_b1 , \13567_b0 );
or ( \13806_b1 , \13803_b1 , \13805_b1 );
xor ( \13806_b0 , \13803_b0 , w_35460 );
not ( w_35460 , w_35461 );
and ( w_35461 , \13805_b1 , \13805_b0 );
or ( \13807_b1 , \13785_b1 , \13795_b1 );
not ( \13795_b1 , w_35462 );
and ( \13807_b0 , \13785_b0 , w_35463 );
and ( w_35462 , w_35463 , \13795_b0 );
or ( \13808_b1 , \13806_b1 , w_35465 );
not ( w_35465 , w_35466 );
and ( \13808_b0 , \13806_b0 , w_35467 );
and ( w_35466 ,  , w_35467 );
buf ( w_35465 , \13807_b1 );
not ( w_35465 , w_35468 );
not (  , w_35469 );
and ( w_35468 , w_35469 , \13807_b0 );
or ( \13809_b1 , \13570_b1 , \13571_b1 );
xor ( \13809_b0 , \13570_b0 , w_35470 );
not ( w_35470 , w_35471 );
and ( w_35471 , \13571_b1 , \13571_b0 );
or ( \13810_b1 , \13809_b1 , \13574_b1 );
xor ( \13810_b0 , \13809_b0 , w_35472 );
not ( w_35472 , w_35473 );
and ( w_35473 , \13574_b1 , \13574_b0 );
or ( \13811_b1 , \13803_b1 , \13805_b1 );
not ( \13805_b1 , w_35474 );
and ( \13811_b0 , \13803_b0 , w_35475 );
and ( w_35474 , w_35475 , \13805_b0 );
or ( \13812_b1 , \13810_b1 , w_35477 );
not ( w_35477 , w_35478 );
and ( \13812_b0 , \13810_b0 , w_35479 );
and ( w_35478 ,  , w_35479 );
buf ( w_35477 , \13811_b1 );
not ( w_35477 , w_35480 );
not (  , w_35481 );
and ( w_35480 , w_35481 , \13811_b0 );
or ( \13813_b1 , \13808_b1 , w_35483 );
not ( w_35483 , w_35484 );
and ( \13813_b0 , \13808_b0 , w_35485 );
and ( w_35484 ,  , w_35485 );
buf ( w_35483 , \13812_b1 );
not ( w_35483 , w_35486 );
not (  , w_35487 );
and ( w_35486 , w_35487 , \13812_b0 );
or ( \13814_b1 , \13799_b1 , w_35489 );
not ( w_35489 , w_35490 );
and ( \13814_b0 , \13799_b0 , w_35491 );
and ( w_35490 ,  , w_35491 );
buf ( w_35489 , \13813_b1 );
not ( w_35489 , w_35492 );
not (  , w_35493 );
and ( w_35492 , w_35493 , \13813_b0 );
or ( \13815_b1 , \13781_b1 , \7012_b1 );
xor ( \13815_b0 , \13781_b0 , w_35494 );
not ( w_35494 , w_35495 );
and ( w_35495 , \7012_b1 , \7012_b0 );
or ( \13816_b1 , \6065_b1 , w_35497 );
not ( w_35497 , w_35498 );
and ( \13816_b0 , \6065_b0 , w_35499 );
and ( w_35498 ,  , w_35499 );
buf ( w_35497 , \7004_b1 );
not ( w_35497 , w_35500 );
not (  , w_35501 );
and ( w_35500 , w_35501 , \7004_b0 );
or ( \13817_b1 , \13816_b1 , w_35502 );
xor ( \13817_b0 , \13816_b0 , w_35504 );
not ( w_35504 , w_35505 );
and ( w_35505 , w_35502 , w_35503 );
buf ( w_35502 , \7012_b1 );
not ( w_35502 , w_35506 );
not ( w_35503 , w_35507 );
and ( w_35506 , w_35507 , \7012_b0 );
or ( \13818_b1 , \13815_b1 , w_35509 );
not ( w_35509 , w_35510 );
and ( \13818_b0 , \13815_b0 , w_35511 );
and ( w_35510 ,  , w_35511 );
buf ( w_35509 , \13817_b1 );
not ( w_35509 , w_35512 );
not (  , w_35513 );
and ( w_35512 , w_35513 , \13817_b0 );
or ( \13819_b1 , \6065_b1 , \6991_b1 );
not ( \6991_b1 , w_35514 );
and ( \13819_b0 , \6065_b0 , w_35515 );
and ( w_35514 , w_35515 , \6991_b0 );
or ( \13820_b1 , \6048_b1 , \6988_b1 );
not ( \6988_b1 , w_35516 );
and ( \13820_b0 , \6048_b0 , w_35517 );
and ( w_35516 , w_35517 , \6988_b0 );
or ( \13821_b1 , \13819_b1 , w_35519 );
not ( w_35519 , w_35520 );
and ( \13821_b0 , \13819_b0 , w_35521 );
and ( w_35520 ,  , w_35521 );
buf ( w_35519 , \13820_b1 );
not ( w_35519 , w_35522 );
not (  , w_35523 );
and ( w_35522 , w_35523 , \13820_b0 );
or ( \13822_b1 , \13821_b1 , w_35524 );
xor ( \13822_b0 , \13821_b0 , w_35526 );
not ( w_35526 , w_35527 );
and ( w_35527 , w_35524 , w_35525 );
buf ( w_35524 , \6985_b1 );
not ( w_35524 , w_35528 );
not ( w_35525 , w_35529 );
and ( w_35528 , w_35529 , \6985_b0 );
or ( \13823_b1 , \6065_b1 , w_35531 );
not ( w_35531 , w_35532 );
and ( \13823_b0 , \6065_b0 , w_35533 );
and ( w_35532 ,  , w_35533 );
buf ( w_35531 , \6988_b1 );
not ( w_35531 , w_35534 );
not (  , w_35535 );
and ( w_35534 , w_35535 , \6988_b0 );
or ( \13824_b1 , \13823_b1 , w_35536 );
xor ( \13824_b0 , \13823_b0 , w_35538 );
not ( w_35538 , w_35539 );
and ( w_35539 , w_35536 , w_35537 );
buf ( w_35536 , \6985_b1 );
not ( w_35536 , w_35540 );
not ( w_35537 , w_35541 );
and ( w_35540 , w_35541 , \6985_b0 );
or ( \13825_b1 , \13824_b1 , \6985_b1 );
not ( \6985_b1 , w_35542 );
and ( \13825_b0 , \13824_b0 , w_35543 );
and ( w_35542 , w_35543 , \6985_b0 );
or ( \13826_b1 , \13822_b1 , w_35545 );
not ( w_35545 , w_35546 );
and ( \13826_b0 , \13822_b0 , w_35547 );
and ( w_35546 ,  , w_35547 );
buf ( w_35545 , \13825_b1 );
not ( w_35545 , w_35548 );
not (  , w_35549 );
and ( w_35548 , w_35549 , \13825_b0 );
or ( \13827_b1 , \13818_b1 , w_35550 );
or ( \13827_b0 , \13818_b0 , \13826_b0 );
not ( \13826_b0 , w_35551 );
and ( w_35551 , w_35550 , \13826_b1 );
or ( \13828_b1 , \13815_b1 , w_35553 );
not ( w_35553 , w_35554 );
and ( \13828_b0 , \13815_b0 , w_35555 );
and ( w_35554 ,  , w_35555 );
buf ( w_35553 , \13817_b1 );
not ( w_35553 , w_35556 );
not (  , w_35557 );
and ( w_35556 , w_35557 , \13817_b0 );
or ( \13829_b1 , \13827_b1 , w_35559 );
not ( w_35559 , w_35560 );
and ( \13829_b0 , \13827_b0 , w_35561 );
and ( w_35560 ,  , w_35561 );
buf ( w_35559 , \13828_b1 );
not ( w_35559 , w_35562 );
not (  , w_35563 );
and ( w_35562 , w_35563 , \13828_b0 );
buf ( \13830_b1 , \13829_b1 );
not ( \13830_b1 , w_35564 );
not ( \13830_b0 , w_35565 );
and ( w_35564 , w_35565 , \13829_b0 );
or ( \13831_b1 , \13814_b1 , w_35566 );
or ( \13831_b0 , \13814_b0 , \13830_b0 );
not ( \13830_b0 , w_35567 );
and ( w_35567 , w_35566 , \13830_b1 );
or ( \13832_b1 , \13777_b1 , w_35569 );
not ( w_35569 , w_35570 );
and ( \13832_b0 , \13777_b0 , w_35571 );
and ( w_35570 ,  , w_35571 );
buf ( w_35569 , \13782_b1 );
not ( w_35569 , w_35572 );
not (  , w_35573 );
and ( w_35572 , w_35573 , \13782_b0 );
or ( \13833_b1 , \13798_b1 , w_35574 );
or ( \13833_b0 , \13798_b0 , \13832_b0 );
not ( \13832_b0 , w_35575 );
and ( w_35575 , w_35574 , \13832_b1 );
or ( \13834_b1 , \13796_b1 , w_35577 );
not ( w_35577 , w_35578 );
and ( \13834_b0 , \13796_b0 , w_35579 );
and ( w_35578 ,  , w_35579 );
buf ( w_35577 , \13797_b1 );
not ( w_35577 , w_35580 );
not (  , w_35581 );
and ( w_35580 , w_35581 , \13797_b0 );
or ( \13835_b1 , \13833_b1 , w_35583 );
not ( w_35583 , w_35584 );
and ( \13835_b0 , \13833_b0 , w_35585 );
and ( w_35584 ,  , w_35585 );
buf ( w_35583 , \13834_b1 );
not ( w_35583 , w_35586 );
not (  , w_35587 );
and ( w_35586 , w_35587 , \13834_b0 );
or ( \13836_b1 , \13813_b1 , \13835_b1 );
not ( \13835_b1 , w_35588 );
and ( \13836_b0 , \13813_b0 , w_35589 );
and ( w_35588 , w_35589 , \13835_b0 );
or ( \13837_b1 , \13806_b1 , w_35591 );
not ( w_35591 , w_35592 );
and ( \13837_b0 , \13806_b0 , w_35593 );
and ( w_35592 ,  , w_35593 );
buf ( w_35591 , \13807_b1 );
not ( w_35591 , w_35594 );
not (  , w_35595 );
and ( w_35594 , w_35595 , \13807_b0 );
or ( \13838_b1 , \13812_b1 , w_35596 );
or ( \13838_b0 , \13812_b0 , \13837_b0 );
not ( \13837_b0 , w_35597 );
and ( w_35597 , w_35596 , \13837_b1 );
or ( \13839_b1 , \13810_b1 , w_35599 );
not ( w_35599 , w_35600 );
and ( \13839_b0 , \13810_b0 , w_35601 );
and ( w_35600 ,  , w_35601 );
buf ( w_35599 , \13811_b1 );
not ( w_35599 , w_35602 );
not (  , w_35603 );
and ( w_35602 , w_35603 , \13811_b0 );
or ( \13840_b1 , \13838_b1 , w_35605 );
not ( w_35605 , w_35606 );
and ( \13840_b0 , \13838_b0 , w_35607 );
and ( w_35606 ,  , w_35607 );
buf ( w_35605 , \13839_b1 );
not ( w_35605 , w_35608 );
not (  , w_35609 );
and ( w_35608 , w_35609 , \13839_b0 );
or ( \13841_b1 , \13836_b1 , w_35611 );
not ( w_35611 , w_35612 );
and ( \13841_b0 , \13836_b0 , w_35613 );
and ( w_35612 ,  , w_35613 );
buf ( w_35611 , \13840_b1 );
not ( w_35611 , w_35614 );
not (  , w_35615 );
and ( w_35614 , w_35615 , \13840_b0 );
or ( \13842_b1 , \13831_b1 , w_35617 );
not ( w_35617 , w_35618 );
and ( \13842_b0 , \13831_b0 , w_35619 );
and ( w_35618 ,  , w_35619 );
buf ( w_35617 , \13841_b1 );
not ( w_35617 , w_35620 );
not (  , w_35621 );
and ( w_35620 , w_35621 , \13841_b0 );
or ( \13843_b1 , \13768_b1 , \13842_b1 );
not ( \13842_b1 , w_35622 );
and ( \13843_b0 , \13768_b0 , w_35623 );
and ( w_35622 , w_35623 , \13842_b0 );
or ( \13844_b1 , \13554_b1 , w_35625 );
not ( w_35625 , w_35626 );
and ( \13844_b0 , \13554_b0 , w_35627 );
and ( w_35626 ,  , w_35627 );
buf ( w_35625 , \13577_b1 );
not ( w_35625 , w_35628 );
not (  , w_35629 );
and ( w_35628 , w_35629 , \13577_b0 );
or ( \13845_b1 , \13613_b1 , w_35630 );
or ( \13845_b0 , \13613_b0 , \13844_b0 );
not ( \13844_b0 , w_35631 );
and ( w_35631 , w_35630 , \13844_b1 );
or ( \13846_b1 , \13611_b1 , w_35633 );
not ( w_35633 , w_35634 );
and ( \13846_b0 , \13611_b0 , w_35635 );
and ( w_35634 ,  , w_35635 );
buf ( w_35633 , \13612_b1 );
not ( w_35633 , w_35636 );
not (  , w_35637 );
and ( w_35636 , w_35637 , \13612_b0 );
or ( \13847_b1 , \13845_b1 , w_35639 );
not ( w_35639 , w_35640 );
and ( \13847_b0 , \13845_b0 , w_35641 );
and ( w_35640 ,  , w_35641 );
buf ( w_35639 , \13846_b1 );
not ( w_35639 , w_35642 );
not (  , w_35643 );
and ( w_35642 , w_35643 , \13846_b0 );
or ( \13848_b1 , \13701_b1 , \13847_b1 );
not ( \13847_b1 , w_35644 );
and ( \13848_b0 , \13701_b0 , w_35645 );
and ( w_35644 , w_35645 , \13847_b0 );
or ( \13849_b1 , \13653_b1 , w_35647 );
not ( w_35647 , w_35648 );
and ( \13849_b0 , \13653_b0 , w_35649 );
and ( w_35648 ,  , w_35649 );
buf ( w_35647 , \13654_b1 );
not ( w_35647 , w_35650 );
not (  , w_35651 );
and ( w_35650 , w_35651 , \13654_b0 );
or ( \13850_b1 , \13700_b1 , w_35652 );
or ( \13850_b0 , \13700_b0 , \13849_b0 );
not ( \13849_b0 , w_35653 );
and ( w_35653 , w_35652 , \13849_b1 );
or ( \13851_b1 , \13695_b1 , w_35655 );
not ( w_35655 , w_35656 );
and ( \13851_b0 , \13695_b0 , w_35657 );
and ( w_35656 ,  , w_35657 );
buf ( w_35655 , \13699_b1 );
not ( w_35655 , w_35658 );
not (  , w_35659 );
and ( w_35658 , w_35659 , \13699_b0 );
or ( \13852_b1 , \13850_b1 , w_35661 );
not ( w_35661 , w_35662 );
and ( \13852_b0 , \13850_b0 , w_35663 );
and ( w_35662 ,  , w_35663 );
buf ( w_35661 , \13851_b1 );
not ( w_35661 , w_35664 );
not (  , w_35665 );
and ( w_35664 , w_35665 , \13851_b0 );
or ( \13853_b1 , \13848_b1 , w_35667 );
not ( w_35667 , w_35668 );
and ( \13853_b0 , \13848_b0 , w_35669 );
and ( w_35668 ,  , w_35669 );
buf ( w_35667 , \13852_b1 );
not ( w_35667 , w_35670 );
not (  , w_35671 );
and ( w_35670 , w_35671 , \13852_b0 );
or ( \13854_b1 , \13767_b1 , w_35672 );
or ( \13854_b0 , \13767_b0 , \13853_b0 );
not ( \13853_b0 , w_35673 );
and ( w_35673 , w_35672 , \13853_b1 );
or ( \13855_b1 , \13727_b1 , w_35675 );
not ( w_35675 , w_35676 );
and ( \13855_b0 , \13727_b0 , w_35677 );
and ( w_35676 ,  , w_35677 );
buf ( w_35675 , \13728_b1 );
not ( w_35675 , w_35678 );
not (  , w_35679 );
and ( w_35678 , w_35679 , \13728_b0 );
or ( \13856_b1 , \13746_b1 , w_35680 );
or ( \13856_b0 , \13746_b0 , \13855_b0 );
not ( \13855_b0 , w_35681 );
and ( w_35681 , w_35680 , \13855_b1 );
or ( \13857_b1 , \13744_b1 , w_35683 );
not ( w_35683 , w_35684 );
and ( \13857_b0 , \13744_b0 , w_35685 );
and ( w_35684 ,  , w_35685 );
buf ( w_35683 , \13745_b1 );
not ( w_35683 , w_35686 );
not (  , w_35687 );
and ( w_35686 , w_35687 , \13745_b0 );
or ( \13858_b1 , \13856_b1 , w_35689 );
not ( w_35689 , w_35690 );
and ( \13858_b0 , \13856_b0 , w_35691 );
and ( w_35690 ,  , w_35691 );
buf ( w_35689 , \13857_b1 );
not ( w_35689 , w_35692 );
not (  , w_35693 );
and ( w_35692 , w_35693 , \13857_b0 );
or ( \13859_b1 , \13766_b1 , \13858_b1 );
not ( \13858_b1 , w_35694 );
and ( \13859_b0 , \13766_b0 , w_35695 );
and ( w_35694 , w_35695 , \13858_b0 );
or ( \13860_b1 , \13756_b1 , w_35697 );
not ( w_35697 , w_35698 );
and ( \13860_b0 , \13756_b0 , w_35699 );
and ( w_35698 ,  , w_35699 );
buf ( w_35697 , \13757_b1 );
not ( w_35697 , w_35700 );
not (  , w_35701 );
and ( w_35700 , w_35701 , \13757_b0 );
or ( \13861_b1 , \13765_b1 , w_35702 );
or ( \13861_b0 , \13765_b0 , \13860_b0 );
not ( \13860_b0 , w_35703 );
and ( w_35703 , w_35702 , \13860_b1 );
or ( \13862_b1 , \13760_b1 , w_35705 );
not ( w_35705 , w_35706 );
and ( \13862_b0 , \13760_b0 , w_35707 );
and ( w_35706 ,  , w_35707 );
buf ( w_35705 , \13764_b1 );
not ( w_35705 , w_35708 );
not (  , w_35709 );
and ( w_35708 , w_35709 , \13764_b0 );
or ( \13863_b1 , \13861_b1 , w_35711 );
not ( w_35711 , w_35712 );
and ( \13863_b0 , \13861_b0 , w_35713 );
and ( w_35712 ,  , w_35713 );
buf ( w_35711 , \13862_b1 );
not ( w_35711 , w_35714 );
not (  , w_35715 );
and ( w_35714 , w_35715 , \13862_b0 );
or ( \13864_b1 , \13859_b1 , w_35717 );
not ( w_35717 , w_35718 );
and ( \13864_b0 , \13859_b0 , w_35719 );
and ( w_35718 ,  , w_35719 );
buf ( w_35717 , \13863_b1 );
not ( w_35717 , w_35720 );
not (  , w_35721 );
and ( w_35720 , w_35721 , \13863_b0 );
or ( \13865_b1 , \13854_b1 , w_35723 );
not ( w_35723 , w_35724 );
and ( \13865_b0 , \13854_b0 , w_35725 );
and ( w_35724 ,  , w_35725 );
buf ( w_35723 , \13864_b1 );
not ( w_35723 , w_35726 );
not (  , w_35727 );
and ( w_35726 , w_35727 , \13864_b0 );
or ( \13866_b1 , \13843_b1 , w_35729 );
not ( w_35729 , w_35730 );
and ( \13866_b0 , \13843_b0 , w_35731 );
and ( w_35730 ,  , w_35731 );
buf ( w_35729 , \13865_b1 );
not ( w_35729 , w_35732 );
not (  , w_35733 );
and ( w_35732 , w_35733 , \13865_b0 );
or ( \13867_b1 , \13514_b1 , w_35734 );
or ( \13867_b0 , \13514_b0 , \13866_b0 );
not ( \13866_b0 , w_35735 );
and ( w_35735 , w_35734 , \13866_b1 );
or ( \13868_b1 , \12375_b1 , w_35737 );
not ( w_35737 , w_35738 );
and ( \13868_b0 , \12375_b0 , w_35739 );
and ( w_35738 ,  , w_35739 );
buf ( w_35737 , \12442_b1 );
not ( w_35737 , w_35740 );
not (  , w_35741 );
and ( w_35740 , w_35741 , \12442_b0 );
or ( \13869_b1 , \12518_b1 , w_35742 );
or ( \13869_b0 , \12518_b0 , \13868_b0 );
not ( \13868_b0 , w_35743 );
and ( w_35743 , w_35742 , \13868_b1 );
or ( \13870_b1 , \12513_b1 , w_35745 );
not ( w_35745 , w_35746 );
and ( \13870_b0 , \12513_b0 , w_35747 );
and ( w_35746 ,  , w_35747 );
buf ( w_35745 , \12517_b1 );
not ( w_35745 , w_35748 );
not (  , w_35749 );
and ( w_35748 , w_35749 , \12517_b0 );
or ( \13871_b1 , \13869_b1 , w_35751 );
not ( w_35751 , w_35752 );
and ( \13871_b0 , \13869_b0 , w_35753 );
and ( w_35752 ,  , w_35753 );
buf ( w_35751 , \13870_b1 );
not ( w_35751 , w_35754 );
not (  , w_35755 );
and ( w_35754 , w_35755 , \13870_b0 );
or ( \13872_b1 , \12686_b1 , \13871_b1 );
not ( \13871_b1 , w_35756 );
and ( \13872_b0 , \12686_b0 , w_35757 );
and ( w_35756 , w_35757 , \13871_b0 );
or ( \13873_b1 , \12595_b1 , w_35759 );
not ( w_35759 , w_35760 );
and ( \13873_b0 , \12595_b0 , w_35761 );
and ( w_35760 ,  , w_35761 );
buf ( w_35759 , \12599_b1 );
not ( w_35759 , w_35762 );
not (  , w_35763 );
and ( w_35762 , w_35763 , \12599_b0 );
or ( \13874_b1 , \12685_b1 , w_35764 );
or ( \13874_b0 , \12685_b0 , \13873_b0 );
not ( \13873_b0 , w_35765 );
and ( w_35765 , w_35764 , \13873_b1 );
or ( \13875_b1 , \12683_b1 , w_35767 );
not ( w_35767 , w_35768 );
and ( \13875_b0 , \12683_b0 , w_35769 );
and ( w_35768 ,  , w_35769 );
buf ( w_35767 , \12684_b1 );
not ( w_35767 , w_35770 );
not (  , w_35771 );
and ( w_35770 , w_35771 , \12684_b0 );
or ( \13876_b1 , \13874_b1 , w_35773 );
not ( w_35773 , w_35774 );
and ( \13876_b0 , \13874_b0 , w_35775 );
and ( w_35774 ,  , w_35775 );
buf ( w_35773 , \13875_b1 );
not ( w_35773 , w_35776 );
not (  , w_35777 );
and ( w_35776 , w_35777 , \13875_b0 );
or ( \13877_b1 , \13872_b1 , w_35779 );
not ( w_35779 , w_35780 );
and ( \13877_b0 , \13872_b0 , w_35781 );
and ( w_35780 ,  , w_35781 );
buf ( w_35779 , \13876_b1 );
not ( w_35779 , w_35782 );
not (  , w_35783 );
and ( w_35782 , w_35783 , \13876_b0 );
or ( \13878_b1 , \13082_b1 , w_35784 );
or ( \13878_b0 , \13082_b0 , \13877_b0 );
not ( \13877_b0 , w_35785 );
and ( w_35785 , w_35784 , \13877_b1 );
or ( \13879_b1 , \12776_b1 , w_35787 );
not ( w_35787 , w_35788 );
and ( \13879_b0 , \12776_b0 , w_35789 );
and ( w_35788 ,  , w_35789 );
buf ( w_35787 , \12777_b1 );
not ( w_35787 , w_35790 );
not (  , w_35791 );
and ( w_35790 , w_35791 , \12777_b0 );
or ( \13880_b1 , \12873_b1 , w_35792 );
or ( \13880_b0 , \12873_b0 , \13879_b0 );
not ( \13879_b0 , w_35793 );
and ( w_35793 , w_35792 , \13879_b1 );
or ( \13881_b1 , \12868_b1 , w_35795 );
not ( w_35795 , w_35796 );
and ( \13881_b0 , \12868_b0 , w_35797 );
and ( w_35796 ,  , w_35797 );
buf ( w_35795 , \12872_b1 );
not ( w_35795 , w_35798 );
not (  , w_35799 );
and ( w_35798 , w_35799 , \12872_b0 );
or ( \13882_b1 , \13880_b1 , w_35801 );
not ( w_35801 , w_35802 );
and ( \13882_b0 , \13880_b0 , w_35803 );
and ( w_35802 ,  , w_35803 );
buf ( w_35801 , \13881_b1 );
not ( w_35801 , w_35804 );
not (  , w_35805 );
and ( w_35804 , w_35805 , \13881_b0 );
or ( \13883_b1 , \13081_b1 , \13882_b1 );
not ( \13882_b1 , w_35806 );
and ( \13883_b0 , \13081_b0 , w_35807 );
and ( w_35806 , w_35807 , \13882_b0 );
or ( \13884_b1 , \12970_b1 , w_35809 );
not ( w_35809 , w_35810 );
and ( \13884_b0 , \12970_b0 , w_35811 );
and ( w_35810 ,  , w_35811 );
buf ( w_35809 , \12974_b1 );
not ( w_35809 , w_35812 );
not (  , w_35813 );
and ( w_35812 , w_35813 , \12974_b0 );
or ( \13885_b1 , \13080_b1 , w_35814 );
or ( \13885_b0 , \13080_b0 , \13884_b0 );
not ( \13884_b0 , w_35815 );
and ( w_35815 , w_35814 , \13884_b1 );
or ( \13886_b1 , \13075_b1 , w_35817 );
not ( w_35817 , w_35818 );
and ( \13886_b0 , \13075_b0 , w_35819 );
and ( w_35818 ,  , w_35819 );
buf ( w_35817 , \13079_b1 );
not ( w_35817 , w_35820 );
not (  , w_35821 );
and ( w_35820 , w_35821 , \13079_b0 );
or ( \13887_b1 , \13885_b1 , w_35823 );
not ( w_35823 , w_35824 );
and ( \13887_b0 , \13885_b0 , w_35825 );
and ( w_35824 ,  , w_35825 );
buf ( w_35823 , \13886_b1 );
not ( w_35823 , w_35826 );
not (  , w_35827 );
and ( w_35826 , w_35827 , \13886_b0 );
or ( \13888_b1 , \13883_b1 , w_35829 );
not ( w_35829 , w_35830 );
and ( \13888_b0 , \13883_b0 , w_35831 );
and ( w_35830 ,  , w_35831 );
buf ( w_35829 , \13887_b1 );
not ( w_35829 , w_35832 );
not (  , w_35833 );
and ( w_35832 , w_35833 , \13887_b0 );
or ( \13889_b1 , \13878_b1 , w_35835 );
not ( w_35835 , w_35836 );
and ( \13889_b0 , \13878_b0 , w_35837 );
and ( w_35836 ,  , w_35837 );
buf ( w_35835 , \13888_b1 );
not ( w_35835 , w_35838 );
not (  , w_35839 );
and ( w_35838 , w_35839 , \13888_b0 );
or ( \13890_b1 , \13513_b1 , \13889_b1 );
not ( \13889_b1 , w_35840 );
and ( \13890_b0 , \13513_b0 , w_35841 );
and ( w_35840 , w_35841 , \13889_b0 );
or ( \13891_b1 , \13189_b1 , w_35843 );
not ( w_35843 , w_35844 );
and ( \13891_b0 , \13189_b0 , w_35845 );
and ( w_35844 ,  , w_35845 );
buf ( w_35843 , \13193_b1 );
not ( w_35843 , w_35846 );
not (  , w_35847 );
and ( w_35846 , w_35847 , \13193_b0 );
or ( \13892_b1 , \13309_b1 , w_35848 );
or ( \13892_b0 , \13309_b0 , \13891_b0 );
not ( \13891_b0 , w_35849 );
and ( w_35849 , w_35848 , \13891_b1 );
or ( \13893_b1 , \13304_b1 , w_35851 );
not ( w_35851 , w_35852 );
and ( \13893_b0 , \13304_b0 , w_35853 );
and ( w_35852 ,  , w_35853 );
buf ( w_35851 , \13308_b1 );
not ( w_35851 , w_35854 );
not (  , w_35855 );
and ( w_35854 , w_35855 , \13308_b0 );
or ( \13894_b1 , \13892_b1 , w_35857 );
not ( w_35857 , w_35858 );
and ( \13894_b0 , \13892_b0 , w_35859 );
and ( w_35858 ,  , w_35859 );
buf ( w_35857 , \13893_b1 );
not ( w_35857 , w_35860 );
not (  , w_35861 );
and ( w_35860 , w_35861 , \13893_b0 );
or ( \13895_b1 , \13429_b1 , \13894_b1 );
not ( \13894_b1 , w_35862 );
and ( \13895_b0 , \13429_b0 , w_35863 );
and ( w_35862 , w_35863 , \13894_b0 );
or ( \13896_b1 , \13378_b1 , w_35865 );
not ( w_35865 , w_35866 );
and ( \13896_b0 , \13378_b0 , w_35867 );
and ( w_35866 ,  , w_35867 );
buf ( w_35865 , \13382_b1 );
not ( w_35865 , w_35868 );
not (  , w_35869 );
and ( w_35868 , w_35869 , \13382_b0 );
or ( \13897_b1 , \13428_b1 , w_35870 );
or ( \13897_b0 , \13428_b0 , \13896_b0 );
not ( \13896_b0 , w_35871 );
and ( w_35871 , w_35870 , \13896_b1 );
or ( \13898_b1 , \13423_b1 , w_35873 );
not ( w_35873 , w_35874 );
and ( \13898_b0 , \13423_b0 , w_35875 );
and ( w_35874 ,  , w_35875 );
buf ( w_35873 , \13427_b1 );
not ( w_35873 , w_35876 );
not (  , w_35877 );
and ( w_35876 , w_35877 , \13427_b0 );
or ( \13899_b1 , \13897_b1 , w_35879 );
not ( w_35879 , w_35880 );
and ( \13899_b0 , \13897_b0 , w_35881 );
and ( w_35880 ,  , w_35881 );
buf ( w_35879 , \13898_b1 );
not ( w_35879 , w_35882 );
not (  , w_35883 );
and ( w_35882 , w_35883 , \13898_b0 );
or ( \13900_b1 , \13895_b1 , w_35885 );
not ( w_35885 , w_35886 );
and ( \13900_b0 , \13895_b0 , w_35887 );
and ( w_35886 ,  , w_35887 );
buf ( w_35885 , \13899_b1 );
not ( w_35885 , w_35888 );
not (  , w_35889 );
and ( w_35888 , w_35889 , \13899_b0 );
or ( \13901_b1 , \13512_b1 , w_35890 );
or ( \13901_b0 , \13512_b0 , \13900_b0 );
not ( \13900_b0 , w_35891 );
and ( w_35891 , w_35890 , \13900_b1 );
or ( \13902_b1 , \13461_b1 , w_35893 );
not ( w_35893 , w_35894 );
and ( \13902_b0 , \13461_b0 , w_35895 );
and ( w_35894 ,  , w_35895 );
buf ( w_35893 , \13462_b1 );
not ( w_35893 , w_35896 );
not (  , w_35897 );
and ( w_35896 , w_35897 , \13462_b0 );
or ( \13903_b1 , \13488_b1 , w_35898 );
or ( \13903_b0 , \13488_b0 , \13902_b0 );
not ( \13902_b0 , w_35899 );
and ( w_35899 , w_35898 , \13902_b1 );
or ( \13904_b1 , \13486_b1 , w_35901 );
not ( w_35901 , w_35902 );
and ( \13904_b0 , \13486_b0 , w_35903 );
and ( w_35902 ,  , w_35903 );
buf ( w_35901 , \13487_b1 );
not ( w_35901 , w_35904 );
not (  , w_35905 );
and ( w_35904 , w_35905 , \13487_b0 );
or ( \13905_b1 , \13903_b1 , w_35907 );
not ( w_35907 , w_35908 );
and ( \13905_b0 , \13903_b0 , w_35909 );
and ( w_35908 ,  , w_35909 );
buf ( w_35907 , \13904_b1 );
not ( w_35907 , w_35910 );
not (  , w_35911 );
and ( w_35910 , w_35911 , \13904_b0 );
or ( \13906_b1 , \13511_b1 , \13905_b1 );
not ( \13905_b1 , w_35912 );
and ( \13906_b0 , \13511_b0 , w_35913 );
and ( w_35912 , w_35913 , \13905_b0 );
or ( \13907_b1 , \13498_b1 , w_35915 );
not ( w_35915 , w_35916 );
and ( \13907_b0 , \13498_b0 , w_35917 );
and ( w_35916 ,  , w_35917 );
buf ( w_35915 , \13502_b1 );
not ( w_35915 , w_35918 );
not (  , w_35919 );
and ( w_35918 , w_35919 , \13502_b0 );
or ( \13908_b1 , \13510_b1 , w_35920 );
or ( \13908_b0 , \13510_b0 , \13907_b0 );
not ( \13907_b0 , w_35921 );
and ( w_35921 , w_35920 , \13907_b1 );
or ( \13909_b1 , \13505_b1 , w_35923 );
not ( w_35923 , w_35924 );
and ( \13909_b0 , \13505_b0 , w_35925 );
and ( w_35924 ,  , w_35925 );
buf ( w_35923 , \13509_b1 );
not ( w_35923 , w_35926 );
not (  , w_35927 );
and ( w_35926 , w_35927 , \13509_b0 );
or ( \13910_b1 , \13908_b1 , w_35929 );
not ( w_35929 , w_35930 );
and ( \13910_b0 , \13908_b0 , w_35931 );
and ( w_35930 ,  , w_35931 );
buf ( w_35929 , \13909_b1 );
not ( w_35929 , w_35932 );
not (  , w_35933 );
and ( w_35932 , w_35933 , \13909_b0 );
or ( \13911_b1 , \13906_b1 , w_35935 );
not ( w_35935 , w_35936 );
and ( \13911_b0 , \13906_b0 , w_35937 );
and ( w_35936 ,  , w_35937 );
buf ( w_35935 , \13910_b1 );
not ( w_35935 , w_35938 );
not (  , w_35939 );
and ( w_35938 , w_35939 , \13910_b0 );
or ( \13912_b1 , \13901_b1 , w_35941 );
not ( w_35941 , w_35942 );
and ( \13912_b0 , \13901_b0 , w_35943 );
and ( w_35942 ,  , w_35943 );
buf ( w_35941 , \13911_b1 );
not ( w_35941 , w_35944 );
not (  , w_35945 );
and ( w_35944 , w_35945 , \13911_b0 );
or ( \13913_b1 , \13890_b1 , w_35947 );
not ( w_35947 , w_35948 );
and ( \13913_b0 , \13890_b0 , w_35949 );
and ( w_35948 ,  , w_35949 );
buf ( w_35947 , \13912_b1 );
not ( w_35947 , w_35950 );
not (  , w_35951 );
and ( w_35950 , w_35951 , \13912_b0 );
or ( \13914_b1 , \13867_b1 , w_35953 );
not ( w_35953 , w_35954 );
and ( \13914_b0 , \13867_b0 , w_35955 );
and ( w_35954 ,  , w_35955 );
buf ( w_35953 , \13913_b1 );
not ( w_35953 , w_35956 );
not (  , w_35957 );
and ( w_35956 , w_35957 , \13913_b0 );
or ( \13915_b1 , \12202_b1 , \13914_b1 );
not ( \13914_b1 , w_35958 );
and ( \13915_b0 , \12202_b0 , w_35959 );
and ( w_35958 , w_35959 , \13914_b0 );
or ( \13916_b1 , \7766_b1 , w_35961 );
not ( w_35961 , w_35962 );
and ( \13916_b0 , \7766_b0 , w_35963 );
and ( w_35962 ,  , w_35963 );
buf ( w_35961 , \7886_b1 );
not ( w_35961 , w_35964 );
not (  , w_35965 );
and ( w_35964 , w_35965 , \7886_b0 );
or ( \13917_b1 , \8041_b1 , w_35966 );
or ( \13917_b0 , \8041_b0 , \13916_b0 );
not ( \13916_b0 , w_35967 );
and ( w_35967 , w_35966 , \13916_b1 );
or ( \13918_b1 , \8036_b1 , w_35969 );
not ( w_35969 , w_35970 );
and ( \13918_b0 , \8036_b0 , w_35971 );
and ( w_35970 ,  , w_35971 );
buf ( w_35969 , \8040_b1 );
not ( w_35969 , w_35972 );
not (  , w_35973 );
and ( w_35972 , w_35973 , \8040_b0 );
or ( \13919_b1 , \13917_b1 , w_35975 );
not ( w_35975 , w_35976 );
and ( \13919_b0 , \13917_b0 , w_35977 );
and ( w_35976 ,  , w_35977 );
buf ( w_35975 , \13918_b1 );
not ( w_35975 , w_35978 );
not (  , w_35979 );
and ( w_35978 , w_35979 , \13918_b0 );
or ( \13920_b1 , \8360_b1 , \13919_b1 );
not ( \13919_b1 , w_35980 );
and ( \13920_b0 , \8360_b0 , w_35981 );
and ( w_35980 , w_35981 , \13919_b0 );
or ( \13921_b1 , \8195_b1 , w_35983 );
not ( w_35983 , w_35984 );
and ( \13921_b0 , \8195_b0 , w_35985 );
and ( w_35984 ,  , w_35985 );
buf ( w_35983 , \8199_b1 );
not ( w_35983 , w_35986 );
not (  , w_35987 );
and ( w_35986 , w_35987 , \8199_b0 );
or ( \13922_b1 , \8359_b1 , w_35988 );
or ( \13922_b0 , \8359_b0 , \13921_b0 );
not ( \13921_b0 , w_35989 );
and ( w_35989 , w_35988 , \13921_b1 );
or ( \13923_b1 , \8354_b1 , w_35991 );
not ( w_35991 , w_35992 );
and ( \13923_b0 , \8354_b0 , w_35993 );
and ( w_35992 ,  , w_35993 );
buf ( w_35991 , \8358_b1 );
not ( w_35991 , w_35994 );
not (  , w_35995 );
and ( w_35994 , w_35995 , \8358_b0 );
or ( \13924_b1 , \13922_b1 , w_35997 );
not ( w_35997 , w_35998 );
and ( \13924_b0 , \13922_b0 , w_35999 );
and ( w_35998 ,  , w_35999 );
buf ( w_35997 , \13923_b1 );
not ( w_35997 , w_36000 );
not (  , w_36001 );
and ( w_36000 , w_36001 , \13923_b0 );
or ( \13925_b1 , \13920_b1 , w_36003 );
not ( w_36003 , w_36004 );
and ( \13925_b0 , \13920_b0 , w_36005 );
and ( w_36004 ,  , w_36005 );
buf ( w_36003 , \13924_b1 );
not ( w_36003 , w_36006 );
not (  , w_36007 );
and ( w_36006 , w_36007 , \13924_b0 );
or ( \13926_b1 , \9009_b1 , w_36008 );
or ( \13926_b0 , \9009_b0 , \13925_b0 );
not ( \13925_b0 , w_36009 );
and ( w_36009 , w_36008 , \13925_b1 );
or ( \13927_b1 , \8516_b1 , w_36011 );
not ( w_36011 , w_36012 );
and ( \13927_b0 , \8516_b0 , w_36013 );
and ( w_36012 ,  , w_36013 );
buf ( w_36011 , \8520_b1 );
not ( w_36011 , w_36014 );
not (  , w_36015 );
and ( w_36014 , w_36015 , \8520_b0 );
or ( \13928_b1 , \8682_b1 , w_36016 );
or ( \13928_b0 , \8682_b0 , \13927_b0 );
not ( \13927_b0 , w_36017 );
and ( w_36017 , w_36016 , \13927_b1 );
or ( \13929_b1 , \8677_b1 , w_36019 );
not ( w_36019 , w_36020 );
and ( \13929_b0 , \8677_b0 , w_36021 );
and ( w_36020 ,  , w_36021 );
buf ( w_36019 , \8681_b1 );
not ( w_36019 , w_36022 );
not (  , w_36023 );
and ( w_36022 , w_36023 , \8681_b0 );
or ( \13930_b1 , \13928_b1 , w_36025 );
not ( w_36025 , w_36026 );
and ( \13930_b0 , \13928_b0 , w_36027 );
and ( w_36026 ,  , w_36027 );
buf ( w_36025 , \13929_b1 );
not ( w_36025 , w_36028 );
not (  , w_36029 );
and ( w_36028 , w_36029 , \13929_b0 );
or ( \13931_b1 , \9008_b1 , \13930_b1 );
not ( \13930_b1 , w_36030 );
and ( \13931_b0 , \9008_b0 , w_36031 );
and ( w_36030 , w_36031 , \13930_b0 );
or ( \13932_b1 , \8841_b1 , w_36033 );
not ( w_36033 , w_36034 );
and ( \13932_b0 , \8841_b0 , w_36035 );
and ( w_36034 ,  , w_36035 );
buf ( w_36033 , \8845_b1 );
not ( w_36033 , w_36036 );
not (  , w_36037 );
and ( w_36036 , w_36037 , \8845_b0 );
or ( \13933_b1 , \9007_b1 , w_36038 );
or ( \13933_b0 , \9007_b0 , \13932_b0 );
not ( \13932_b0 , w_36039 );
and ( w_36039 , w_36038 , \13932_b1 );
or ( \13934_b1 , \9002_b1 , w_36041 );
not ( w_36041 , w_36042 );
and ( \13934_b0 , \9002_b0 , w_36043 );
and ( w_36042 ,  , w_36043 );
buf ( w_36041 , \9006_b1 );
not ( w_36041 , w_36044 );
not (  , w_36045 );
and ( w_36044 , w_36045 , \9006_b0 );
or ( \13935_b1 , \13933_b1 , w_36047 );
not ( w_36047 , w_36048 );
and ( \13935_b0 , \13933_b0 , w_36049 );
and ( w_36048 ,  , w_36049 );
buf ( w_36047 , \13934_b1 );
not ( w_36047 , w_36050 );
not (  , w_36051 );
and ( w_36050 , w_36051 , \13934_b0 );
or ( \13936_b1 , \13931_b1 , w_36053 );
not ( w_36053 , w_36054 );
and ( \13936_b0 , \13931_b0 , w_36055 );
and ( w_36054 ,  , w_36055 );
buf ( w_36053 , \13935_b1 );
not ( w_36053 , w_36056 );
not (  , w_36057 );
and ( w_36056 , w_36057 , \13935_b0 );
or ( \13937_b1 , \13926_b1 , w_36059 );
not ( w_36059 , w_36060 );
and ( \13937_b0 , \13926_b0 , w_36061 );
and ( w_36060 ,  , w_36061 );
buf ( w_36059 , \13936_b1 );
not ( w_36059 , w_36062 );
not (  , w_36063 );
and ( w_36062 , w_36063 , \13936_b0 );
or ( \13938_b1 , \10313_b1 , \13937_b1 );
not ( \13937_b1 , w_36064 );
and ( \13938_b0 , \10313_b0 , w_36065 );
and ( w_36064 , w_36065 , \13937_b0 );
or ( \13939_b1 , \9168_b1 , w_36067 );
not ( w_36067 , w_36068 );
and ( \13939_b0 , \9168_b0 , w_36069 );
and ( w_36068 ,  , w_36069 );
buf ( w_36067 , \9172_b1 );
not ( w_36067 , w_36070 );
not (  , w_36071 );
and ( w_36070 , w_36071 , \9172_b0 );
or ( \13940_b1 , \9334_b1 , w_36072 );
or ( \13940_b0 , \9334_b0 , \13939_b0 );
not ( \13939_b0 , w_36073 );
and ( w_36073 , w_36072 , \13939_b1 );
or ( \13941_b1 , \9329_b1 , w_36075 );
not ( w_36075 , w_36076 );
and ( \13941_b0 , \9329_b0 , w_36077 );
and ( w_36076 ,  , w_36077 );
buf ( w_36075 , \9333_b1 );
not ( w_36075 , w_36078 );
not (  , w_36079 );
and ( w_36078 , w_36079 , \9333_b0 );
or ( \13942_b1 , \13940_b1 , w_36081 );
not ( w_36081 , w_36082 );
and ( \13942_b0 , \13940_b0 , w_36083 );
and ( w_36082 ,  , w_36083 );
buf ( w_36081 , \13941_b1 );
not ( w_36081 , w_36084 );
not (  , w_36085 );
and ( w_36084 , w_36085 , \13941_b0 );
or ( \13943_b1 , \9660_b1 , \13942_b1 );
not ( \13942_b1 , w_36086 );
and ( \13943_b0 , \9660_b0 , w_36087 );
and ( w_36086 , w_36087 , \13942_b0 );
or ( \13944_b1 , \9493_b1 , w_36089 );
not ( w_36089 , w_36090 );
and ( \13944_b0 , \9493_b0 , w_36091 );
and ( w_36090 ,  , w_36091 );
buf ( w_36089 , \9497_b1 );
not ( w_36089 , w_36092 );
not (  , w_36093 );
and ( w_36092 , w_36093 , \9497_b0 );
or ( \13945_b1 , \9659_b1 , w_36094 );
or ( \13945_b0 , \9659_b0 , \13944_b0 );
not ( \13944_b0 , w_36095 );
and ( w_36095 , w_36094 , \13944_b1 );
or ( \13946_b1 , \9654_b1 , w_36097 );
not ( w_36097 , w_36098 );
and ( \13946_b0 , \9654_b0 , w_36099 );
and ( w_36098 ,  , w_36099 );
buf ( w_36097 , \9658_b1 );
not ( w_36097 , w_36100 );
not (  , w_36101 );
and ( w_36100 , w_36101 , \9658_b0 );
or ( \13947_b1 , \13945_b1 , w_36103 );
not ( w_36103 , w_36104 );
and ( \13947_b0 , \13945_b0 , w_36105 );
and ( w_36104 ,  , w_36105 );
buf ( w_36103 , \13946_b1 );
not ( w_36103 , w_36106 );
not (  , w_36107 );
and ( w_36106 , w_36107 , \13946_b0 );
or ( \13948_b1 , \13943_b1 , w_36109 );
not ( w_36109 , w_36110 );
and ( \13948_b0 , \13943_b0 , w_36111 );
and ( w_36110 ,  , w_36111 );
buf ( w_36109 , \13947_b1 );
not ( w_36109 , w_36112 );
not (  , w_36113 );
and ( w_36112 , w_36113 , \13947_b0 );
or ( \13949_b1 , \10312_b1 , w_36114 );
or ( \13949_b0 , \10312_b0 , \13948_b0 );
not ( \13948_b0 , w_36115 );
and ( w_36115 , w_36114 , \13948_b1 );
or ( \13950_b1 , \9819_b1 , w_36117 );
not ( w_36117 , w_36118 );
and ( \13950_b0 , \9819_b0 , w_36119 );
and ( w_36118 ,  , w_36119 );
buf ( w_36117 , \9823_b1 );
not ( w_36117 , w_36120 );
not (  , w_36121 );
and ( w_36120 , w_36121 , \9823_b0 );
or ( \13951_b1 , \9985_b1 , w_36122 );
or ( \13951_b0 , \9985_b0 , \13950_b0 );
not ( \13950_b0 , w_36123 );
and ( w_36123 , w_36122 , \13950_b1 );
or ( \13952_b1 , \9980_b1 , w_36125 );
not ( w_36125 , w_36126 );
and ( \13952_b0 , \9980_b0 , w_36127 );
and ( w_36126 ,  , w_36127 );
buf ( w_36125 , \9984_b1 );
not ( w_36125 , w_36128 );
not (  , w_36129 );
and ( w_36128 , w_36129 , \9984_b0 );
or ( \13953_b1 , \13951_b1 , w_36131 );
not ( w_36131 , w_36132 );
and ( \13953_b0 , \13951_b0 , w_36133 );
and ( w_36132 ,  , w_36133 );
buf ( w_36131 , \13952_b1 );
not ( w_36131 , w_36134 );
not (  , w_36135 );
and ( w_36134 , w_36135 , \13952_b0 );
or ( \13954_b1 , \10311_b1 , \13953_b1 );
not ( \13953_b1 , w_36136 );
and ( \13954_b0 , \10311_b0 , w_36137 );
and ( w_36136 , w_36137 , \13953_b0 );
or ( \13955_b1 , \10144_b1 , w_36139 );
not ( w_36139 , w_36140 );
and ( \13955_b0 , \10144_b0 , w_36141 );
and ( w_36140 ,  , w_36141 );
buf ( w_36139 , \10148_b1 );
not ( w_36139 , w_36142 );
not (  , w_36143 );
and ( w_36142 , w_36143 , \10148_b0 );
or ( \13956_b1 , \10310_b1 , w_36144 );
or ( \13956_b0 , \10310_b0 , \13955_b0 );
not ( \13955_b0 , w_36145 );
and ( w_36145 , w_36144 , \13955_b1 );
or ( \13957_b1 , \10305_b1 , w_36147 );
not ( w_36147 , w_36148 );
and ( \13957_b0 , \10305_b0 , w_36149 );
and ( w_36148 ,  , w_36149 );
buf ( w_36147 , \10309_b1 );
not ( w_36147 , w_36150 );
not (  , w_36151 );
and ( w_36150 , w_36151 , \10309_b0 );
or ( \13958_b1 , \13956_b1 , w_36153 );
not ( w_36153 , w_36154 );
and ( \13958_b0 , \13956_b0 , w_36155 );
and ( w_36154 ,  , w_36155 );
buf ( w_36153 , \13957_b1 );
not ( w_36153 , w_36156 );
not (  , w_36157 );
and ( w_36156 , w_36157 , \13957_b0 );
or ( \13959_b1 , \13954_b1 , w_36159 );
not ( w_36159 , w_36160 );
and ( \13959_b0 , \13954_b0 , w_36161 );
and ( w_36160 ,  , w_36161 );
buf ( w_36159 , \13958_b1 );
not ( w_36159 , w_36162 );
not (  , w_36163 );
and ( w_36162 , w_36163 , \13958_b0 );
or ( \13960_b1 , \13949_b1 , w_36165 );
not ( w_36165 , w_36166 );
and ( \13960_b0 , \13949_b0 , w_36167 );
and ( w_36166 ,  , w_36167 );
buf ( w_36165 , \13959_b1 );
not ( w_36165 , w_36168 );
not (  , w_36169 );
and ( w_36168 , w_36169 , \13959_b0 );
or ( \13961_b1 , \13938_b1 , w_36171 );
not ( w_36171 , w_36172 );
and ( \13961_b0 , \13938_b0 , w_36173 );
and ( w_36172 ,  , w_36173 );
buf ( w_36171 , \13960_b1 );
not ( w_36171 , w_36174 );
not (  , w_36175 );
and ( w_36174 , w_36175 , \13960_b0 );
or ( \13962_b1 , \12201_b1 , w_36176 );
or ( \13962_b0 , \12201_b0 , \13961_b0 );
not ( \13961_b0 , w_36177 );
and ( w_36177 , w_36176 , \13961_b1 );
or ( \13963_b1 , \10472_b1 , w_36179 );
not ( w_36179 , w_36180 );
and ( \13963_b0 , \10472_b0 , w_36181 );
and ( w_36180 ,  , w_36181 );
buf ( w_36179 , \10476_b1 );
not ( w_36179 , w_36182 );
not (  , w_36183 );
and ( w_36182 , w_36183 , \10476_b0 );
or ( \13964_b1 , \10638_b1 , w_36184 );
or ( \13964_b0 , \10638_b0 , \13963_b0 );
not ( \13963_b0 , w_36185 );
and ( w_36185 , w_36184 , \13963_b1 );
or ( \13965_b1 , \10633_b1 , w_36187 );
not ( w_36187 , w_36188 );
and ( \13965_b0 , \10633_b0 , w_36189 );
and ( w_36188 ,  , w_36189 );
buf ( w_36187 , \10637_b1 );
not ( w_36187 , w_36190 );
not (  , w_36191 );
and ( w_36190 , w_36191 , \10637_b0 );
or ( \13966_b1 , \13964_b1 , w_36193 );
not ( w_36193 , w_36194 );
and ( \13966_b0 , \13964_b0 , w_36195 );
and ( w_36194 ,  , w_36195 );
buf ( w_36193 , \13965_b1 );
not ( w_36193 , w_36196 );
not (  , w_36197 );
and ( w_36196 , w_36197 , \13965_b0 );
or ( \13967_b1 , \10964_b1 , \13966_b1 );
not ( \13966_b1 , w_36198 );
and ( \13967_b0 , \10964_b0 , w_36199 );
and ( w_36198 , w_36199 , \13966_b0 );
or ( \13968_b1 , \10797_b1 , w_36201 );
not ( w_36201 , w_36202 );
and ( \13968_b0 , \10797_b0 , w_36203 );
and ( w_36202 ,  , w_36203 );
buf ( w_36201 , \10801_b1 );
not ( w_36201 , w_36204 );
not (  , w_36205 );
and ( w_36204 , w_36205 , \10801_b0 );
or ( \13969_b1 , \10963_b1 , w_36206 );
or ( \13969_b0 , \10963_b0 , \13968_b0 );
not ( \13968_b0 , w_36207 );
and ( w_36207 , w_36206 , \13968_b1 );
or ( \13970_b1 , \10958_b1 , w_36209 );
not ( w_36209 , w_36210 );
and ( \13970_b0 , \10958_b0 , w_36211 );
and ( w_36210 ,  , w_36211 );
buf ( w_36209 , \10962_b1 );
not ( w_36209 , w_36212 );
not (  , w_36213 );
and ( w_36212 , w_36213 , \10962_b0 );
or ( \13971_b1 , \13969_b1 , w_36215 );
not ( w_36215 , w_36216 );
and ( \13971_b0 , \13969_b0 , w_36217 );
and ( w_36216 ,  , w_36217 );
buf ( w_36215 , \13970_b1 );
not ( w_36215 , w_36218 );
not (  , w_36219 );
and ( w_36218 , w_36219 , \13970_b0 );
or ( \13972_b1 , \13967_b1 , w_36221 );
not ( w_36221 , w_36222 );
and ( \13972_b0 , \13967_b0 , w_36223 );
and ( w_36222 ,  , w_36223 );
buf ( w_36221 , \13971_b1 );
not ( w_36221 , w_36224 );
not (  , w_36225 );
and ( w_36224 , w_36225 , \13971_b0 );
or ( \13973_b1 , \11616_b1 , w_36226 );
or ( \13973_b0 , \11616_b0 , \13972_b0 );
not ( \13972_b0 , w_36227 );
and ( w_36227 , w_36226 , \13972_b1 );
or ( \13974_b1 , \11123_b1 , w_36229 );
not ( w_36229 , w_36230 );
and ( \13974_b0 , \11123_b0 , w_36231 );
and ( w_36230 ,  , w_36231 );
buf ( w_36229 , \11127_b1 );
not ( w_36229 , w_36232 );
not (  , w_36233 );
and ( w_36232 , w_36233 , \11127_b0 );
or ( \13975_b1 , \11289_b1 , w_36234 );
or ( \13975_b0 , \11289_b0 , \13974_b0 );
not ( \13974_b0 , w_36235 );
and ( w_36235 , w_36234 , \13974_b1 );
or ( \13976_b1 , \11284_b1 , w_36237 );
not ( w_36237 , w_36238 );
and ( \13976_b0 , \11284_b0 , w_36239 );
and ( w_36238 ,  , w_36239 );
buf ( w_36237 , \11288_b1 );
not ( w_36237 , w_36240 );
not (  , w_36241 );
and ( w_36240 , w_36241 , \11288_b0 );
or ( \13977_b1 , \13975_b1 , w_36243 );
not ( w_36243 , w_36244 );
and ( \13977_b0 , \13975_b0 , w_36245 );
and ( w_36244 ,  , w_36245 );
buf ( w_36243 , \13976_b1 );
not ( w_36243 , w_36246 );
not (  , w_36247 );
and ( w_36246 , w_36247 , \13976_b0 );
or ( \13978_b1 , \11615_b1 , \13977_b1 );
not ( \13977_b1 , w_36248 );
and ( \13978_b0 , \11615_b0 , w_36249 );
and ( w_36248 , w_36249 , \13977_b0 );
or ( \13979_b1 , \11448_b1 , w_36251 );
not ( w_36251 , w_36252 );
and ( \13979_b0 , \11448_b0 , w_36253 );
and ( w_36252 ,  , w_36253 );
buf ( w_36251 , \11452_b1 );
not ( w_36251 , w_36254 );
not (  , w_36255 );
and ( w_36254 , w_36255 , \11452_b0 );
or ( \13980_b1 , \11614_b1 , w_36256 );
or ( \13980_b0 , \11614_b0 , \13979_b0 );
not ( \13979_b0 , w_36257 );
and ( w_36257 , w_36256 , \13979_b1 );
or ( \13981_b1 , \11609_b1 , w_36259 );
not ( w_36259 , w_36260 );
and ( \13981_b0 , \11609_b0 , w_36261 );
and ( w_36260 ,  , w_36261 );
buf ( w_36259 , \11613_b1 );
not ( w_36259 , w_36262 );
not (  , w_36263 );
and ( w_36262 , w_36263 , \11613_b0 );
or ( \13982_b1 , \13980_b1 , w_36265 );
not ( w_36265 , w_36266 );
and ( \13982_b0 , \13980_b0 , w_36267 );
and ( w_36266 ,  , w_36267 );
buf ( w_36265 , \13981_b1 );
not ( w_36265 , w_36268 );
not (  , w_36269 );
and ( w_36268 , w_36269 , \13981_b0 );
or ( \13983_b1 , \13978_b1 , w_36271 );
not ( w_36271 , w_36272 );
and ( \13983_b0 , \13978_b0 , w_36273 );
and ( w_36272 ,  , w_36273 );
buf ( w_36271 , \13982_b1 );
not ( w_36271 , w_36274 );
not (  , w_36275 );
and ( w_36274 , w_36275 , \13982_b0 );
or ( \13984_b1 , \13973_b1 , w_36277 );
not ( w_36277 , w_36278 );
and ( \13984_b0 , \13973_b0 , w_36279 );
and ( w_36278 ,  , w_36279 );
buf ( w_36277 , \13983_b1 );
not ( w_36277 , w_36280 );
not (  , w_36281 );
and ( w_36280 , w_36281 , \13983_b0 );
or ( \13985_b1 , \12200_b1 , \13984_b1 );
not ( \13984_b1 , w_36282 );
and ( \13985_b0 , \12200_b0 , w_36283 );
and ( w_36282 , w_36283 , \13984_b0 );
or ( \13986_b1 , \11775_b1 , w_36285 );
not ( w_36285 , w_36286 );
and ( \13986_b0 , \11775_b0 , w_36287 );
and ( w_36286 ,  , w_36287 );
buf ( w_36285 , \11779_b1 );
not ( w_36285 , w_36288 );
not (  , w_36289 );
and ( w_36288 , w_36289 , \11779_b0 );
or ( \13987_b1 , \11941_b1 , w_36290 );
or ( \13987_b0 , \11941_b0 , \13986_b0 );
not ( \13986_b0 , w_36291 );
and ( w_36291 , w_36290 , \13986_b1 );
or ( \13988_b1 , \11936_b1 , w_36293 );
not ( w_36293 , w_36294 );
and ( \13988_b0 , \11936_b0 , w_36295 );
and ( w_36294 ,  , w_36295 );
buf ( w_36293 , \11940_b1 );
not ( w_36293 , w_36296 );
not (  , w_36297 );
and ( w_36296 , w_36297 , \11940_b0 );
or ( \13989_b1 , \13987_b1 , w_36299 );
not ( w_36299 , w_36300 );
and ( \13989_b0 , \13987_b0 , w_36301 );
and ( w_36300 ,  , w_36301 );
buf ( w_36299 , \13988_b1 );
not ( w_36299 , w_36302 );
not (  , w_36303 );
and ( w_36302 , w_36303 , \13988_b0 );
or ( \13990_b1 , \12106_b1 , \13989_b1 );
not ( \13989_b1 , w_36304 );
and ( \13990_b0 , \12106_b0 , w_36305 );
and ( w_36304 , w_36305 , \13989_b0 );
or ( \13991_b1 , \12035_b1 , w_36307 );
not ( w_36307 , w_36308 );
and ( \13991_b0 , \12035_b0 , w_36309 );
and ( w_36308 ,  , w_36309 );
buf ( w_36307 , \12039_b1 );
not ( w_36307 , w_36310 );
not (  , w_36311 );
and ( w_36310 , w_36311 , \12039_b0 );
or ( \13992_b1 , \12105_b1 , w_36312 );
or ( \13992_b0 , \12105_b0 , \13991_b0 );
not ( \13991_b0 , w_36313 );
and ( w_36313 , w_36312 , \13991_b1 );
or ( \13993_b1 , \12100_b1 , w_36315 );
not ( w_36315 , w_36316 );
and ( \13993_b0 , \12100_b0 , w_36317 );
and ( w_36316 ,  , w_36317 );
buf ( w_36315 , \12104_b1 );
not ( w_36315 , w_36318 );
not (  , w_36319 );
and ( w_36318 , w_36319 , \12104_b0 );
or ( \13994_b1 , \13992_b1 , w_36321 );
not ( w_36321 , w_36322 );
and ( \13994_b0 , \13992_b0 , w_36323 );
and ( w_36322 ,  , w_36323 );
buf ( w_36321 , \13993_b1 );
not ( w_36321 , w_36324 );
not (  , w_36325 );
and ( w_36324 , w_36325 , \13993_b0 );
or ( \13995_b1 , \13990_b1 , w_36327 );
not ( w_36327 , w_36328 );
and ( \13995_b0 , \13990_b0 , w_36329 );
and ( w_36328 ,  , w_36329 );
buf ( w_36327 , \13994_b1 );
not ( w_36327 , w_36330 );
not (  , w_36331 );
and ( w_36330 , w_36331 , \13994_b0 );
or ( \13996_b1 , \12199_b1 , w_36332 );
or ( \13996_b0 , \12199_b0 , \13995_b0 );
not ( \13995_b0 , w_36333 );
and ( w_36333 , w_36332 , \13995_b1 );
or ( \13997_b1 , \12144_b1 , w_36335 );
not ( w_36335 , w_36336 );
and ( \13997_b0 , \12144_b0 , w_36337 );
and ( w_36336 ,  , w_36337 );
buf ( w_36335 , \12148_b1 );
not ( w_36335 , w_36338 );
not (  , w_36339 );
and ( w_36338 , w_36339 , \12148_b0 );
or ( \13998_b1 , \12174_b1 , w_36340 );
or ( \13998_b0 , \12174_b0 , \13997_b0 );
not ( \13997_b0 , w_36341 );
and ( w_36341 , w_36340 , \13997_b1 );
or ( \13999_b1 , \12169_b1 , w_36343 );
not ( w_36343 , w_36344 );
and ( \13999_b0 , \12169_b0 , w_36345 );
and ( w_36344 ,  , w_36345 );
buf ( w_36343 , \12173_b1 );
not ( w_36343 , w_36346 );
not (  , w_36347 );
and ( w_36346 , w_36347 , \12173_b0 );
or ( \14000_b1 , \13998_b1 , w_36349 );
not ( w_36349 , w_36350 );
and ( \14000_b0 , \13998_b0 , w_36351 );
and ( w_36350 ,  , w_36351 );
buf ( w_36349 , \13999_b1 );
not ( w_36349 , w_36352 );
not (  , w_36353 );
and ( w_36352 , w_36353 , \13999_b0 );
or ( \14001_b1 , \12198_b1 , \14000_b1 );
not ( \14000_b1 , w_36354 );
and ( \14001_b0 , \12198_b0 , w_36355 );
and ( w_36354 , w_36355 , \14000_b0 );
or ( \14002_b1 , \12185_b1 , w_36357 );
not ( w_36357 , w_36358 );
and ( \14002_b0 , \12185_b0 , w_36359 );
and ( w_36358 ,  , w_36359 );
buf ( w_36357 , \12189_b1 );
not ( w_36357 , w_36360 );
not (  , w_36361 );
and ( w_36360 , w_36361 , \12189_b0 );
or ( \14003_b1 , \12197_b1 , w_36362 );
or ( \14003_b0 , \12197_b0 , \14002_b0 );
not ( \14002_b0 , w_36363 );
and ( w_36363 , w_36362 , \14002_b1 );
or ( \14004_b1 , \12192_b1 , w_36365 );
not ( w_36365 , w_36366 );
and ( \14004_b0 , \12192_b0 , w_36367 );
and ( w_36366 ,  , w_36367 );
buf ( w_36365 , \12196_b1 );
not ( w_36365 , w_36368 );
not (  , w_36369 );
and ( w_36368 , w_36369 , \12196_b0 );
or ( \14005_b1 , \14003_b1 , w_36371 );
not ( w_36371 , w_36372 );
and ( \14005_b0 , \14003_b0 , w_36373 );
and ( w_36372 ,  , w_36373 );
buf ( w_36371 , \14004_b1 );
not ( w_36371 , w_36374 );
not (  , w_36375 );
and ( w_36374 , w_36375 , \14004_b0 );
or ( \14006_b1 , \14001_b1 , w_36377 );
not ( w_36377 , w_36378 );
and ( \14006_b0 , \14001_b0 , w_36379 );
and ( w_36378 ,  , w_36379 );
buf ( w_36377 , \14005_b1 );
not ( w_36377 , w_36380 );
not (  , w_36381 );
and ( w_36380 , w_36381 , \14005_b0 );
or ( \14007_b1 , \13996_b1 , w_36383 );
not ( w_36383 , w_36384 );
and ( \14007_b0 , \13996_b0 , w_36385 );
and ( w_36384 ,  , w_36385 );
buf ( w_36383 , \14006_b1 );
not ( w_36383 , w_36386 );
not (  , w_36387 );
and ( w_36386 , w_36387 , \14006_b0 );
or ( \14008_b1 , \13985_b1 , w_36389 );
not ( w_36389 , w_36390 );
and ( \14008_b0 , \13985_b0 , w_36391 );
and ( w_36390 ,  , w_36391 );
buf ( w_36389 , \14007_b1 );
not ( w_36389 , w_36392 );
not (  , w_36393 );
and ( w_36392 , w_36393 , \14007_b0 );
or ( \14009_b1 , \13962_b1 , w_36395 );
not ( w_36395 , w_36396 );
and ( \14009_b0 , \13962_b0 , w_36397 );
and ( w_36396 ,  , w_36397 );
buf ( w_36395 , \14008_b1 );
not ( w_36395 , w_36398 );
not (  , w_36399 );
and ( w_36398 , w_36399 , \14008_b0 );
or ( \14010_b1 , \13915_b1 , w_36401 );
not ( w_36401 , w_36402 );
and ( \14010_b0 , \13915_b0 , w_36403 );
and ( w_36402 ,  , w_36403 );
buf ( w_36401 , \14009_b1 );
not ( w_36401 , w_36404 );
not (  , w_36405 );
and ( w_36404 , w_36405 , \14009_b0 );
buf ( \14011_b1 , \14010_b1 );
not ( \14011_b1 , w_36406 );
not ( \14011_b0 , w_36407 );
and ( w_36406 , w_36407 , \14010_b0 );
or ( \14012_b1 , \6982_b1 , w_36408 );
xor ( \14012_b0 , \6982_b0 , w_36410 );
not ( w_36410 , w_36411 );
and ( w_36411 , w_36408 , w_36409 );
buf ( w_36408 , \14011_b1 );
not ( w_36408 , w_36412 );
not ( w_36409 , w_36413 );
and ( w_36412 , w_36413 , \14011_b0 );
buf ( \14013_b1 , \14012_b1 );
buf ( \14013_b0 , \14012_b0 );
buf ( \14014_b1 , \14013_b1 );
buf ( \14014_b0 , \14013_b0 );
buf ( \14015_b1 , \12197_b1 );
not ( \14015_b1 , w_36414 );
not ( \14015_b0 , w_36415 );
and ( w_36414 , w_36415 , \12197_b0 );
or ( \14016_b1 , \14004_b1 , w_36417 );
not ( w_36417 , w_36418 );
and ( \14016_b0 , \14004_b0 , w_36419 );
and ( w_36418 ,  , w_36419 );
buf ( w_36417 , \14015_b1 );
not ( w_36417 , w_36420 );
not (  , w_36421 );
and ( w_36420 , w_36421 , \14015_b0 );
or ( \14017_b1 , \13510_b1 , w_36423 );
not ( w_36423 , w_36424 );
and ( \14017_b0 , \13510_b0 , w_36425 );
and ( w_36424 ,  , w_36425 );
buf ( w_36423 , \7887_b1 );
not ( w_36423 , w_36426 );
not (  , w_36427 );
and ( w_36426 , w_36427 , \7887_b0 );
or ( \14018_b1 , \8041_b1 , w_36429 );
not ( w_36429 , w_36430 );
and ( \14018_b0 , \8041_b0 , w_36431 );
and ( w_36430 ,  , w_36431 );
buf ( w_36429 , \8200_b1 );
not ( w_36429 , w_36432 );
not (  , w_36433 );
and ( w_36432 , w_36433 , \8200_b0 );
or ( \14019_b1 , \14017_b1 , w_36435 );
not ( w_36435 , w_36436 );
and ( \14019_b0 , \14017_b0 , w_36437 );
and ( w_36436 ,  , w_36437 );
buf ( w_36435 , \14018_b1 );
not ( w_36435 , w_36438 );
not (  , w_36439 );
and ( w_36438 , w_36439 , \14018_b0 );
or ( \14020_b1 , \8359_b1 , w_36441 );
not ( w_36441 , w_36442 );
and ( \14020_b0 , \8359_b0 , w_36443 );
and ( w_36442 ,  , w_36443 );
buf ( w_36441 , \8521_b1 );
not ( w_36441 , w_36444 );
not (  , w_36445 );
and ( w_36444 , w_36445 , \8521_b0 );
or ( \14021_b1 , \8682_b1 , w_36447 );
not ( w_36447 , w_36448 );
and ( \14021_b0 , \8682_b0 , w_36449 );
and ( w_36448 ,  , w_36449 );
buf ( w_36447 , \8846_b1 );
not ( w_36447 , w_36450 );
not (  , w_36451 );
and ( w_36450 , w_36451 , \8846_b0 );
or ( \14022_b1 , \14020_b1 , w_36453 );
not ( w_36453 , w_36454 );
and ( \14022_b0 , \14020_b0 , w_36455 );
and ( w_36454 ,  , w_36455 );
buf ( w_36453 , \14021_b1 );
not ( w_36453 , w_36456 );
not (  , w_36457 );
and ( w_36456 , w_36457 , \14021_b0 );
or ( \14023_b1 , \14019_b1 , w_36459 );
not ( w_36459 , w_36460 );
and ( \14023_b0 , \14019_b0 , w_36461 );
and ( w_36460 ,  , w_36461 );
buf ( w_36459 , \14022_b1 );
not ( w_36459 , w_36462 );
not (  , w_36463 );
and ( w_36462 , w_36463 , \14022_b0 );
or ( \14024_b1 , \9007_b1 , w_36465 );
not ( w_36465 , w_36466 );
and ( \14024_b0 , \9007_b0 , w_36467 );
and ( w_36466 ,  , w_36467 );
buf ( w_36465 , \9173_b1 );
not ( w_36465 , w_36468 );
not (  , w_36469 );
and ( w_36468 , w_36469 , \9173_b0 );
or ( \14025_b1 , \9334_b1 , w_36471 );
not ( w_36471 , w_36472 );
and ( \14025_b0 , \9334_b0 , w_36473 );
and ( w_36472 ,  , w_36473 );
buf ( w_36471 , \9498_b1 );
not ( w_36471 , w_36474 );
not (  , w_36475 );
and ( w_36474 , w_36475 , \9498_b0 );
or ( \14026_b1 , \14024_b1 , w_36477 );
not ( w_36477 , w_36478 );
and ( \14026_b0 , \14024_b0 , w_36479 );
and ( w_36478 ,  , w_36479 );
buf ( w_36477 , \14025_b1 );
not ( w_36477 , w_36480 );
not (  , w_36481 );
and ( w_36480 , w_36481 , \14025_b0 );
or ( \14027_b1 , \9659_b1 , w_36483 );
not ( w_36483 , w_36484 );
and ( \14027_b0 , \9659_b0 , w_36485 );
and ( w_36484 ,  , w_36485 );
buf ( w_36483 , \9824_b1 );
not ( w_36483 , w_36486 );
not (  , w_36487 );
and ( w_36486 , w_36487 , \9824_b0 );
or ( \14028_b1 , \9985_b1 , w_36489 );
not ( w_36489 , w_36490 );
and ( \14028_b0 , \9985_b0 , w_36491 );
and ( w_36490 ,  , w_36491 );
buf ( w_36489 , \10149_b1 );
not ( w_36489 , w_36492 );
not (  , w_36493 );
and ( w_36492 , w_36493 , \10149_b0 );
or ( \14029_b1 , \14027_b1 , w_36495 );
not ( w_36495 , w_36496 );
and ( \14029_b0 , \14027_b0 , w_36497 );
and ( w_36496 ,  , w_36497 );
buf ( w_36495 , \14028_b1 );
not ( w_36495 , w_36498 );
not (  , w_36499 );
and ( w_36498 , w_36499 , \14028_b0 );
or ( \14030_b1 , \14026_b1 , w_36501 );
not ( w_36501 , w_36502 );
and ( \14030_b0 , \14026_b0 , w_36503 );
and ( w_36502 ,  , w_36503 );
buf ( w_36501 , \14029_b1 );
not ( w_36501 , w_36504 );
not (  , w_36505 );
and ( w_36504 , w_36505 , \14029_b0 );
or ( \14031_b1 , \14023_b1 , w_36507 );
not ( w_36507 , w_36508 );
and ( \14031_b0 , \14023_b0 , w_36509 );
and ( w_36508 ,  , w_36509 );
buf ( w_36507 , \14030_b1 );
not ( w_36507 , w_36510 );
not (  , w_36511 );
and ( w_36510 , w_36511 , \14030_b0 );
or ( \14032_b1 , \10310_b1 , w_36513 );
not ( w_36513 , w_36514 );
and ( \14032_b0 , \10310_b0 , w_36515 );
and ( w_36514 ,  , w_36515 );
buf ( w_36513 , \10477_b1 );
not ( w_36513 , w_36516 );
not (  , w_36517 );
and ( w_36516 , w_36517 , \10477_b0 );
or ( \14033_b1 , \10638_b1 , w_36519 );
not ( w_36519 , w_36520 );
and ( \14033_b0 , \10638_b0 , w_36521 );
and ( w_36520 ,  , w_36521 );
buf ( w_36519 , \10802_b1 );
not ( w_36519 , w_36522 );
not (  , w_36523 );
and ( w_36522 , w_36523 , \10802_b0 );
or ( \14034_b1 , \14032_b1 , w_36525 );
not ( w_36525 , w_36526 );
and ( \14034_b0 , \14032_b0 , w_36527 );
and ( w_36526 ,  , w_36527 );
buf ( w_36525 , \14033_b1 );
not ( w_36525 , w_36528 );
not (  , w_36529 );
and ( w_36528 , w_36529 , \14033_b0 );
or ( \14035_b1 , \10963_b1 , w_36531 );
not ( w_36531 , w_36532 );
and ( \14035_b0 , \10963_b0 , w_36533 );
and ( w_36532 ,  , w_36533 );
buf ( w_36531 , \11128_b1 );
not ( w_36531 , w_36534 );
not (  , w_36535 );
and ( w_36534 , w_36535 , \11128_b0 );
or ( \14036_b1 , \11289_b1 , w_36537 );
not ( w_36537 , w_36538 );
and ( \14036_b0 , \11289_b0 , w_36539 );
and ( w_36538 ,  , w_36539 );
buf ( w_36537 , \11453_b1 );
not ( w_36537 , w_36540 );
not (  , w_36541 );
and ( w_36540 , w_36541 , \11453_b0 );
or ( \14037_b1 , \14035_b1 , w_36543 );
not ( w_36543 , w_36544 );
and ( \14037_b0 , \14035_b0 , w_36545 );
and ( w_36544 ,  , w_36545 );
buf ( w_36543 , \14036_b1 );
not ( w_36543 , w_36546 );
not (  , w_36547 );
and ( w_36546 , w_36547 , \14036_b0 );
or ( \14038_b1 , \14034_b1 , w_36549 );
not ( w_36549 , w_36550 );
and ( \14038_b0 , \14034_b0 , w_36551 );
and ( w_36550 ,  , w_36551 );
buf ( w_36549 , \14037_b1 );
not ( w_36549 , w_36552 );
not (  , w_36553 );
and ( w_36552 , w_36553 , \14037_b0 );
or ( \14039_b1 , \11614_b1 , w_36555 );
not ( w_36555 , w_36556 );
and ( \14039_b0 , \11614_b0 , w_36557 );
and ( w_36556 ,  , w_36557 );
buf ( w_36555 , \11780_b1 );
not ( w_36555 , w_36558 );
not (  , w_36559 );
and ( w_36558 , w_36559 , \11780_b0 );
or ( \14040_b1 , \11941_b1 , w_36561 );
not ( w_36561 , w_36562 );
and ( \14040_b0 , \11941_b0 , w_36563 );
and ( w_36562 ,  , w_36563 );
buf ( w_36561 , \12040_b1 );
not ( w_36561 , w_36564 );
not (  , w_36565 );
and ( w_36564 , w_36565 , \12040_b0 );
or ( \14041_b1 , \14039_b1 , w_36567 );
not ( w_36567 , w_36568 );
and ( \14041_b0 , \14039_b0 , w_36569 );
and ( w_36568 ,  , w_36569 );
buf ( w_36567 , \14040_b1 );
not ( w_36567 , w_36570 );
not (  , w_36571 );
and ( w_36570 , w_36571 , \14040_b0 );
or ( \14042_b1 , \12105_b1 , w_36573 );
not ( w_36573 , w_36574 );
and ( \14042_b0 , \12105_b0 , w_36575 );
and ( w_36574 ,  , w_36575 );
buf ( w_36573 , \12149_b1 );
not ( w_36573 , w_36576 );
not (  , w_36577 );
and ( w_36576 , w_36577 , \12149_b0 );
or ( \14043_b1 , \12174_b1 , w_36579 );
not ( w_36579 , w_36580 );
and ( \14043_b0 , \12174_b0 , w_36581 );
and ( w_36580 ,  , w_36581 );
buf ( w_36579 , \12190_b1 );
not ( w_36579 , w_36582 );
not (  , w_36583 );
and ( w_36582 , w_36583 , \12190_b0 );
or ( \14044_b1 , \14042_b1 , w_36585 );
not ( w_36585 , w_36586 );
and ( \14044_b0 , \14042_b0 , w_36587 );
and ( w_36586 ,  , w_36587 );
buf ( w_36585 , \14043_b1 );
not ( w_36585 , w_36588 );
not (  , w_36589 );
and ( w_36588 , w_36589 , \14043_b0 );
or ( \14045_b1 , \14041_b1 , w_36591 );
not ( w_36591 , w_36592 );
and ( \14045_b0 , \14041_b0 , w_36593 );
and ( w_36592 ,  , w_36593 );
buf ( w_36591 , \14044_b1 );
not ( w_36591 , w_36594 );
not (  , w_36595 );
and ( w_36594 , w_36595 , \14044_b0 );
or ( \14046_b1 , \14038_b1 , w_36597 );
not ( w_36597 , w_36598 );
and ( \14046_b0 , \14038_b0 , w_36599 );
and ( w_36598 ,  , w_36599 );
buf ( w_36597 , \14045_b1 );
not ( w_36597 , w_36600 );
not (  , w_36601 );
and ( w_36600 , w_36601 , \14045_b0 );
or ( \14047_b1 , \14031_b1 , w_36603 );
not ( w_36603 , w_36604 );
and ( \14047_b0 , \14031_b0 , w_36605 );
and ( w_36604 ,  , w_36605 );
buf ( w_36603 , \14046_b1 );
not ( w_36603 , w_36606 );
not (  , w_36607 );
and ( w_36606 , w_36607 , \14046_b0 );
or ( \14048_b1 , \13765_b1 , w_36609 );
not ( w_36609 , w_36610 );
and ( \14048_b0 , \13765_b0 , w_36611 );
and ( w_36610 ,  , w_36611 );
buf ( w_36609 , \12443_b1 );
not ( w_36609 , w_36612 );
not (  , w_36613 );
and ( w_36612 , w_36613 , \12443_b0 );
or ( \14049_b1 , \12518_b1 , w_36615 );
not ( w_36615 , w_36616 );
and ( \14049_b0 , \12518_b0 , w_36617 );
and ( w_36616 ,  , w_36617 );
buf ( w_36615 , \12600_b1 );
not ( w_36615 , w_36618 );
not (  , w_36619 );
and ( w_36618 , w_36619 , \12600_b0 );
or ( \14050_b1 , \14048_b1 , w_36621 );
not ( w_36621 , w_36622 );
and ( \14050_b0 , \14048_b0 , w_36623 );
and ( w_36622 ,  , w_36623 );
buf ( w_36621 , \14049_b1 );
not ( w_36621 , w_36624 );
not (  , w_36625 );
and ( w_36624 , w_36625 , \14049_b0 );
or ( \14051_b1 , \12685_b1 , w_36627 );
not ( w_36627 , w_36628 );
and ( \14051_b0 , \12685_b0 , w_36629 );
and ( w_36628 ,  , w_36629 );
buf ( w_36627 , \12778_b1 );
not ( w_36627 , w_36630 );
not (  , w_36631 );
and ( w_36630 , w_36631 , \12778_b0 );
or ( \14052_b1 , \12873_b1 , w_36633 );
not ( w_36633 , w_36634 );
and ( \14052_b0 , \12873_b0 , w_36635 );
and ( w_36634 ,  , w_36635 );
buf ( w_36633 , \12975_b1 );
not ( w_36633 , w_36636 );
not (  , w_36637 );
and ( w_36636 , w_36637 , \12975_b0 );
or ( \14053_b1 , \14051_b1 , w_36639 );
not ( w_36639 , w_36640 );
and ( \14053_b0 , \14051_b0 , w_36641 );
and ( w_36640 ,  , w_36641 );
buf ( w_36639 , \14052_b1 );
not ( w_36639 , w_36642 );
not (  , w_36643 );
and ( w_36642 , w_36643 , \14052_b0 );
or ( \14054_b1 , \14050_b1 , w_36645 );
not ( w_36645 , w_36646 );
and ( \14054_b0 , \14050_b0 , w_36647 );
and ( w_36646 ,  , w_36647 );
buf ( w_36645 , \14053_b1 );
not ( w_36645 , w_36648 );
not (  , w_36649 );
and ( w_36648 , w_36649 , \14053_b0 );
or ( \14055_b1 , \13080_b1 , w_36651 );
not ( w_36651 , w_36652 );
and ( \14055_b0 , \13080_b0 , w_36653 );
and ( w_36652 ,  , w_36653 );
buf ( w_36651 , \13194_b1 );
not ( w_36651 , w_36654 );
not (  , w_36655 );
and ( w_36654 , w_36655 , \13194_b0 );
or ( \14056_b1 , \13309_b1 , w_36657 );
not ( w_36657 , w_36658 );
and ( \14056_b0 , \13309_b0 , w_36659 );
and ( w_36658 ,  , w_36659 );
buf ( w_36657 , \13383_b1 );
not ( w_36657 , w_36660 );
not (  , w_36661 );
and ( w_36660 , w_36661 , \13383_b0 );
or ( \14057_b1 , \14055_b1 , w_36663 );
not ( w_36663 , w_36664 );
and ( \14057_b0 , \14055_b0 , w_36665 );
and ( w_36664 ,  , w_36665 );
buf ( w_36663 , \14056_b1 );
not ( w_36663 , w_36666 );
not (  , w_36667 );
and ( w_36666 , w_36667 , \14056_b0 );
or ( \14058_b1 , \13428_b1 , w_36669 );
not ( w_36669 , w_36670 );
and ( \14058_b0 , \13428_b0 , w_36671 );
and ( w_36670 ,  , w_36671 );
buf ( w_36669 , \13463_b1 );
not ( w_36669 , w_36672 );
not (  , w_36673 );
and ( w_36672 , w_36673 , \13463_b0 );
or ( \14059_b1 , \13488_b1 , w_36675 );
not ( w_36675 , w_36676 );
and ( \14059_b0 , \13488_b0 , w_36677 );
and ( w_36676 ,  , w_36677 );
buf ( w_36675 , \13503_b1 );
not ( w_36675 , w_36678 );
not (  , w_36679 );
and ( w_36678 , w_36679 , \13503_b0 );
or ( \14060_b1 , \14058_b1 , w_36681 );
not ( w_36681 , w_36682 );
and ( \14060_b0 , \14058_b0 , w_36683 );
and ( w_36682 ,  , w_36683 );
buf ( w_36681 , \14059_b1 );
not ( w_36681 , w_36684 );
not (  , w_36685 );
and ( w_36684 , w_36685 , \14059_b0 );
or ( \14061_b1 , \14057_b1 , w_36687 );
not ( w_36687 , w_36688 );
and ( \14061_b0 , \14057_b0 , w_36689 );
and ( w_36688 ,  , w_36689 );
buf ( w_36687 , \14060_b1 );
not ( w_36687 , w_36690 );
not (  , w_36691 );
and ( w_36690 , w_36691 , \14060_b0 );
or ( \14062_b1 , \14054_b1 , w_36693 );
not ( w_36693 , w_36694 );
and ( \14062_b0 , \14054_b0 , w_36695 );
and ( w_36694 ,  , w_36695 );
buf ( w_36693 , \14061_b1 );
not ( w_36693 , w_36696 );
not (  , w_36697 );
and ( w_36696 , w_36697 , \14061_b0 );
or ( \14063_b1 , \13812_b1 , w_36699 );
not ( w_36699 , w_36700 );
and ( \14063_b0 , \13812_b0 , w_36701 );
and ( w_36700 ,  , w_36701 );
buf ( w_36699 , \13578_b1 );
not ( w_36699 , w_36702 );
not (  , w_36703 );
and ( w_36702 , w_36703 , \13578_b0 );
or ( \14064_b1 , \13613_b1 , w_36705 );
not ( w_36705 , w_36706 );
and ( \14064_b0 , \13613_b0 , w_36707 );
and ( w_36706 ,  , w_36707 );
buf ( w_36705 , \13655_b1 );
not ( w_36705 , w_36708 );
not (  , w_36709 );
and ( w_36708 , w_36709 , \13655_b0 );
or ( \14065_b1 , \14063_b1 , w_36711 );
not ( w_36711 , w_36712 );
and ( \14065_b0 , \14063_b0 , w_36713 );
and ( w_36712 ,  , w_36713 );
buf ( w_36711 , \14064_b1 );
not ( w_36711 , w_36714 );
not (  , w_36715 );
and ( w_36714 , w_36715 , \14064_b0 );
or ( \14066_b1 , \13700_b1 , w_36717 );
not ( w_36717 , w_36718 );
and ( \14066_b0 , \13700_b0 , w_36719 );
and ( w_36718 ,  , w_36719 );
buf ( w_36717 , \13729_b1 );
not ( w_36717 , w_36720 );
not (  , w_36721 );
and ( w_36720 , w_36721 , \13729_b0 );
or ( \14067_b1 , \13746_b1 , w_36723 );
not ( w_36723 , w_36724 );
and ( \14067_b0 , \13746_b0 , w_36725 );
and ( w_36724 ,  , w_36725 );
buf ( w_36723 , \13758_b1 );
not ( w_36723 , w_36726 );
not (  , w_36727 );
and ( w_36726 , w_36727 , \13758_b0 );
or ( \14068_b1 , \14066_b1 , w_36729 );
not ( w_36729 , w_36730 );
and ( \14068_b0 , \14066_b0 , w_36731 );
and ( w_36730 ,  , w_36731 );
buf ( w_36729 , \14067_b1 );
not ( w_36729 , w_36732 );
not (  , w_36733 );
and ( w_36732 , w_36733 , \14067_b0 );
or ( \14069_b1 , \14065_b1 , w_36735 );
not ( w_36735 , w_36736 );
and ( \14069_b0 , \14065_b0 , w_36737 );
and ( w_36736 ,  , w_36737 );
buf ( w_36735 , \14068_b1 );
not ( w_36735 , w_36738 );
not (  , w_36739 );
and ( w_36738 , w_36739 , \14068_b0 );
or ( \14070_b1 , \13818_b1 , w_36741 );
not ( w_36741 , w_36742 );
and ( \14070_b0 , \13818_b0 , w_36743 );
and ( w_36742 ,  , w_36743 );
buf ( w_36741 , \13783_b1 );
not ( w_36741 , w_36744 );
not (  , w_36745 );
and ( w_36744 , w_36745 , \13783_b0 );
or ( \14071_b1 , \13798_b1 , w_36747 );
not ( w_36747 , w_36748 );
and ( \14071_b0 , \13798_b0 , w_36749 );
and ( w_36748 ,  , w_36749 );
buf ( w_36747 , \13808_b1 );
not ( w_36747 , w_36750 );
not (  , w_36751 );
and ( w_36750 , w_36751 , \13808_b0 );
or ( \14072_b1 , \14070_b1 , w_36753 );
not ( w_36753 , w_36754 );
and ( \14072_b0 , \14070_b0 , w_36755 );
and ( w_36754 ,  , w_36755 );
buf ( w_36753 , \14071_b1 );
not ( w_36753 , w_36756 );
not (  , w_36757 );
and ( w_36756 , w_36757 , \14071_b0 );
or ( \14073_b1 , \14072_b1 , w_36758 );
or ( \14073_b0 , \14072_b0 , \13826_b0 );
not ( \13826_b0 , w_36759 );
and ( w_36759 , w_36758 , \13826_b1 );
or ( \14074_b1 , \13783_b1 , w_36760 );
or ( \14074_b0 , \13783_b0 , \13828_b0 );
not ( \13828_b0 , w_36761 );
and ( w_36761 , w_36760 , \13828_b1 );
or ( \14075_b1 , \14074_b1 , w_36763 );
not ( w_36763 , w_36764 );
and ( \14075_b0 , \14074_b0 , w_36765 );
and ( w_36764 ,  , w_36765 );
buf ( w_36763 , \13832_b1 );
not ( w_36763 , w_36766 );
not (  , w_36767 );
and ( w_36766 , w_36767 , \13832_b0 );
or ( \14076_b1 , \14071_b1 , \14075_b1 );
not ( \14075_b1 , w_36768 );
and ( \14076_b0 , \14071_b0 , w_36769 );
and ( w_36768 , w_36769 , \14075_b0 );
or ( \14077_b1 , \13808_b1 , w_36770 );
or ( \14077_b0 , \13808_b0 , \13834_b0 );
not ( \13834_b0 , w_36771 );
and ( w_36771 , w_36770 , \13834_b1 );
or ( \14078_b1 , \14077_b1 , w_36773 );
not ( w_36773 , w_36774 );
and ( \14078_b0 , \14077_b0 , w_36775 );
and ( w_36774 ,  , w_36775 );
buf ( w_36773 , \13837_b1 );
not ( w_36773 , w_36776 );
not (  , w_36777 );
and ( w_36776 , w_36777 , \13837_b0 );
or ( \14079_b1 , \14076_b1 , w_36779 );
not ( w_36779 , w_36780 );
and ( \14079_b0 , \14076_b0 , w_36781 );
and ( w_36780 ,  , w_36781 );
buf ( w_36779 , \14078_b1 );
not ( w_36779 , w_36782 );
not (  , w_36783 );
and ( w_36782 , w_36783 , \14078_b0 );
or ( \14080_b1 , \14073_b1 , w_36785 );
not ( w_36785 , w_36786 );
and ( \14080_b0 , \14073_b0 , w_36787 );
and ( w_36786 ,  , w_36787 );
buf ( w_36785 , \14079_b1 );
not ( w_36785 , w_36788 );
not (  , w_36789 );
and ( w_36788 , w_36789 , \14079_b0 );
or ( \14081_b1 , \14069_b1 , \14080_b1 );
not ( \14080_b1 , w_36790 );
and ( \14081_b0 , \14069_b0 , w_36791 );
and ( w_36790 , w_36791 , \14080_b0 );
or ( \14082_b1 , \13578_b1 , w_36792 );
or ( \14082_b0 , \13578_b0 , \13839_b0 );
not ( \13839_b0 , w_36793 );
and ( w_36793 , w_36792 , \13839_b1 );
or ( \14083_b1 , \14082_b1 , w_36795 );
not ( w_36795 , w_36796 );
and ( \14083_b0 , \14082_b0 , w_36797 );
and ( w_36796 ,  , w_36797 );
buf ( w_36795 , \13844_b1 );
not ( w_36795 , w_36798 );
not (  , w_36799 );
and ( w_36798 , w_36799 , \13844_b0 );
or ( \14084_b1 , \14064_b1 , \14083_b1 );
not ( \14083_b1 , w_36800 );
and ( \14084_b0 , \14064_b0 , w_36801 );
and ( w_36800 , w_36801 , \14083_b0 );
or ( \14085_b1 , \13655_b1 , w_36802 );
or ( \14085_b0 , \13655_b0 , \13846_b0 );
not ( \13846_b0 , w_36803 );
and ( w_36803 , w_36802 , \13846_b1 );
or ( \14086_b1 , \14085_b1 , w_36805 );
not ( w_36805 , w_36806 );
and ( \14086_b0 , \14085_b0 , w_36807 );
and ( w_36806 ,  , w_36807 );
buf ( w_36805 , \13849_b1 );
not ( w_36805 , w_36808 );
not (  , w_36809 );
and ( w_36808 , w_36809 , \13849_b0 );
or ( \14087_b1 , \14084_b1 , w_36811 );
not ( w_36811 , w_36812 );
and ( \14087_b0 , \14084_b0 , w_36813 );
and ( w_36812 ,  , w_36813 );
buf ( w_36811 , \14086_b1 );
not ( w_36811 , w_36814 );
not (  , w_36815 );
and ( w_36814 , w_36815 , \14086_b0 );
or ( \14088_b1 , \14068_b1 , w_36816 );
or ( \14088_b0 , \14068_b0 , \14087_b0 );
not ( \14087_b0 , w_36817 );
and ( w_36817 , w_36816 , \14087_b1 );
or ( \14089_b1 , \13729_b1 , w_36818 );
or ( \14089_b0 , \13729_b0 , \13851_b0 );
not ( \13851_b0 , w_36819 );
and ( w_36819 , w_36818 , \13851_b1 );
or ( \14090_b1 , \14089_b1 , w_36821 );
not ( w_36821 , w_36822 );
and ( \14090_b0 , \14089_b0 , w_36823 );
and ( w_36822 ,  , w_36823 );
buf ( w_36821 , \13855_b1 );
not ( w_36821 , w_36824 );
not (  , w_36825 );
and ( w_36824 , w_36825 , \13855_b0 );
or ( \14091_b1 , \14067_b1 , \14090_b1 );
not ( \14090_b1 , w_36826 );
and ( \14091_b0 , \14067_b0 , w_36827 );
and ( w_36826 , w_36827 , \14090_b0 );
or ( \14092_b1 , \13758_b1 , w_36828 );
or ( \14092_b0 , \13758_b0 , \13857_b0 );
not ( \13857_b0 , w_36829 );
and ( w_36829 , w_36828 , \13857_b1 );
or ( \14093_b1 , \14092_b1 , w_36831 );
not ( w_36831 , w_36832 );
and ( \14093_b0 , \14092_b0 , w_36833 );
and ( w_36832 ,  , w_36833 );
buf ( w_36831 , \13860_b1 );
not ( w_36831 , w_36834 );
not (  , w_36835 );
and ( w_36834 , w_36835 , \13860_b0 );
or ( \14094_b1 , \14091_b1 , w_36837 );
not ( w_36837 , w_36838 );
and ( \14094_b0 , \14091_b0 , w_36839 );
and ( w_36838 ,  , w_36839 );
buf ( w_36837 , \14093_b1 );
not ( w_36837 , w_36840 );
not (  , w_36841 );
and ( w_36840 , w_36841 , \14093_b0 );
or ( \14095_b1 , \14088_b1 , w_36843 );
not ( w_36843 , w_36844 );
and ( \14095_b0 , \14088_b0 , w_36845 );
and ( w_36844 ,  , w_36845 );
buf ( w_36843 , \14094_b1 );
not ( w_36843 , w_36846 );
not (  , w_36847 );
and ( w_36846 , w_36847 , \14094_b0 );
or ( \14096_b1 , \14081_b1 , w_36849 );
not ( w_36849 , w_36850 );
and ( \14096_b0 , \14081_b0 , w_36851 );
and ( w_36850 ,  , w_36851 );
buf ( w_36849 , \14095_b1 );
not ( w_36849 , w_36852 );
not (  , w_36853 );
and ( w_36852 , w_36853 , \14095_b0 );
or ( \14097_b1 , \14062_b1 , w_36854 );
or ( \14097_b0 , \14062_b0 , \14096_b0 );
not ( \14096_b0 , w_36855 );
and ( w_36855 , w_36854 , \14096_b1 );
or ( \14098_b1 , \12443_b1 , w_36856 );
or ( \14098_b0 , \12443_b0 , \13862_b0 );
not ( \13862_b0 , w_36857 );
and ( w_36857 , w_36856 , \13862_b1 );
or ( \14099_b1 , \14098_b1 , w_36859 );
not ( w_36859 , w_36860 );
and ( \14099_b0 , \14098_b0 , w_36861 );
and ( w_36860 ,  , w_36861 );
buf ( w_36859 , \13868_b1 );
not ( w_36859 , w_36862 );
not (  , w_36863 );
and ( w_36862 , w_36863 , \13868_b0 );
or ( \14100_b1 , \14049_b1 , \14099_b1 );
not ( \14099_b1 , w_36864 );
and ( \14100_b0 , \14049_b0 , w_36865 );
and ( w_36864 , w_36865 , \14099_b0 );
or ( \14101_b1 , \12600_b1 , w_36866 );
or ( \14101_b0 , \12600_b0 , \13870_b0 );
not ( \13870_b0 , w_36867 );
and ( w_36867 , w_36866 , \13870_b1 );
or ( \14102_b1 , \14101_b1 , w_36869 );
not ( w_36869 , w_36870 );
and ( \14102_b0 , \14101_b0 , w_36871 );
and ( w_36870 ,  , w_36871 );
buf ( w_36869 , \13873_b1 );
not ( w_36869 , w_36872 );
not (  , w_36873 );
and ( w_36872 , w_36873 , \13873_b0 );
or ( \14103_b1 , \14100_b1 , w_36875 );
not ( w_36875 , w_36876 );
and ( \14103_b0 , \14100_b0 , w_36877 );
and ( w_36876 ,  , w_36877 );
buf ( w_36875 , \14102_b1 );
not ( w_36875 , w_36878 );
not (  , w_36879 );
and ( w_36878 , w_36879 , \14102_b0 );
or ( \14104_b1 , \14053_b1 , w_36880 );
or ( \14104_b0 , \14053_b0 , \14103_b0 );
not ( \14103_b0 , w_36881 );
and ( w_36881 , w_36880 , \14103_b1 );
or ( \14105_b1 , \12778_b1 , w_36882 );
or ( \14105_b0 , \12778_b0 , \13875_b0 );
not ( \13875_b0 , w_36883 );
and ( w_36883 , w_36882 , \13875_b1 );
or ( \14106_b1 , \14105_b1 , w_36885 );
not ( w_36885 , w_36886 );
and ( \14106_b0 , \14105_b0 , w_36887 );
and ( w_36886 ,  , w_36887 );
buf ( w_36885 , \13879_b1 );
not ( w_36885 , w_36888 );
not (  , w_36889 );
and ( w_36888 , w_36889 , \13879_b0 );
or ( \14107_b1 , \14052_b1 , \14106_b1 );
not ( \14106_b1 , w_36890 );
and ( \14107_b0 , \14052_b0 , w_36891 );
and ( w_36890 , w_36891 , \14106_b0 );
or ( \14108_b1 , \12975_b1 , w_36892 );
or ( \14108_b0 , \12975_b0 , \13881_b0 );
not ( \13881_b0 , w_36893 );
and ( w_36893 , w_36892 , \13881_b1 );
or ( \14109_b1 , \14108_b1 , w_36895 );
not ( w_36895 , w_36896 );
and ( \14109_b0 , \14108_b0 , w_36897 );
and ( w_36896 ,  , w_36897 );
buf ( w_36895 , \13884_b1 );
not ( w_36895 , w_36898 );
not (  , w_36899 );
and ( w_36898 , w_36899 , \13884_b0 );
or ( \14110_b1 , \14107_b1 , w_36901 );
not ( w_36901 , w_36902 );
and ( \14110_b0 , \14107_b0 , w_36903 );
and ( w_36902 ,  , w_36903 );
buf ( w_36901 , \14109_b1 );
not ( w_36901 , w_36904 );
not (  , w_36905 );
and ( w_36904 , w_36905 , \14109_b0 );
or ( \14111_b1 , \14104_b1 , w_36907 );
not ( w_36907 , w_36908 );
and ( \14111_b0 , \14104_b0 , w_36909 );
and ( w_36908 ,  , w_36909 );
buf ( w_36907 , \14110_b1 );
not ( w_36907 , w_36910 );
not (  , w_36911 );
and ( w_36910 , w_36911 , \14110_b0 );
or ( \14112_b1 , \14061_b1 , \14111_b1 );
not ( \14111_b1 , w_36912 );
and ( \14112_b0 , \14061_b0 , w_36913 );
and ( w_36912 , w_36913 , \14111_b0 );
or ( \14113_b1 , \13194_b1 , w_36914 );
or ( \14113_b0 , \13194_b0 , \13886_b0 );
not ( \13886_b0 , w_36915 );
and ( w_36915 , w_36914 , \13886_b1 );
or ( \14114_b1 , \14113_b1 , w_36917 );
not ( w_36917 , w_36918 );
and ( \14114_b0 , \14113_b0 , w_36919 );
and ( w_36918 ,  , w_36919 );
buf ( w_36917 , \13891_b1 );
not ( w_36917 , w_36920 );
not (  , w_36921 );
and ( w_36920 , w_36921 , \13891_b0 );
or ( \14115_b1 , \14056_b1 , \14114_b1 );
not ( \14114_b1 , w_36922 );
and ( \14115_b0 , \14056_b0 , w_36923 );
and ( w_36922 , w_36923 , \14114_b0 );
or ( \14116_b1 , \13383_b1 , w_36924 );
or ( \14116_b0 , \13383_b0 , \13893_b0 );
not ( \13893_b0 , w_36925 );
and ( w_36925 , w_36924 , \13893_b1 );
or ( \14117_b1 , \14116_b1 , w_36927 );
not ( w_36927 , w_36928 );
and ( \14117_b0 , \14116_b0 , w_36929 );
and ( w_36928 ,  , w_36929 );
buf ( w_36927 , \13896_b1 );
not ( w_36927 , w_36930 );
not (  , w_36931 );
and ( w_36930 , w_36931 , \13896_b0 );
or ( \14118_b1 , \14115_b1 , w_36933 );
not ( w_36933 , w_36934 );
and ( \14118_b0 , \14115_b0 , w_36935 );
and ( w_36934 ,  , w_36935 );
buf ( w_36933 , \14117_b1 );
not ( w_36933 , w_36936 );
not (  , w_36937 );
and ( w_36936 , w_36937 , \14117_b0 );
or ( \14119_b1 , \14060_b1 , w_36938 );
or ( \14119_b0 , \14060_b0 , \14118_b0 );
not ( \14118_b0 , w_36939 );
and ( w_36939 , w_36938 , \14118_b1 );
or ( \14120_b1 , \13463_b1 , w_36940 );
or ( \14120_b0 , \13463_b0 , \13898_b0 );
not ( \13898_b0 , w_36941 );
and ( w_36941 , w_36940 , \13898_b1 );
or ( \14121_b1 , \14120_b1 , w_36943 );
not ( w_36943 , w_36944 );
and ( \14121_b0 , \14120_b0 , w_36945 );
and ( w_36944 ,  , w_36945 );
buf ( w_36943 , \13902_b1 );
not ( w_36943 , w_36946 );
not (  , w_36947 );
and ( w_36946 , w_36947 , \13902_b0 );
or ( \14122_b1 , \14059_b1 , \14121_b1 );
not ( \14121_b1 , w_36948 );
and ( \14122_b0 , \14059_b0 , w_36949 );
and ( w_36948 , w_36949 , \14121_b0 );
or ( \14123_b1 , \13503_b1 , w_36950 );
or ( \14123_b0 , \13503_b0 , \13904_b0 );
not ( \13904_b0 , w_36951 );
and ( w_36951 , w_36950 , \13904_b1 );
or ( \14124_b1 , \14123_b1 , w_36953 );
not ( w_36953 , w_36954 );
and ( \14124_b0 , \14123_b0 , w_36955 );
and ( w_36954 ,  , w_36955 );
buf ( w_36953 , \13907_b1 );
not ( w_36953 , w_36956 );
not (  , w_36957 );
and ( w_36956 , w_36957 , \13907_b0 );
or ( \14125_b1 , \14122_b1 , w_36959 );
not ( w_36959 , w_36960 );
and ( \14125_b0 , \14122_b0 , w_36961 );
and ( w_36960 ,  , w_36961 );
buf ( w_36959 , \14124_b1 );
not ( w_36959 , w_36962 );
not (  , w_36963 );
and ( w_36962 , w_36963 , \14124_b0 );
or ( \14126_b1 , \14119_b1 , w_36965 );
not ( w_36965 , w_36966 );
and ( \14126_b0 , \14119_b0 , w_36967 );
and ( w_36966 ,  , w_36967 );
buf ( w_36965 , \14125_b1 );
not ( w_36965 , w_36968 );
not (  , w_36969 );
and ( w_36968 , w_36969 , \14125_b0 );
or ( \14127_b1 , \14112_b1 , w_36971 );
not ( w_36971 , w_36972 );
and ( \14127_b0 , \14112_b0 , w_36973 );
and ( w_36972 ,  , w_36973 );
buf ( w_36971 , \14126_b1 );
not ( w_36971 , w_36974 );
not (  , w_36975 );
and ( w_36974 , w_36975 , \14126_b0 );
or ( \14128_b1 , \14097_b1 , w_36977 );
not ( w_36977 , w_36978 );
and ( \14128_b0 , \14097_b0 , w_36979 );
and ( w_36978 ,  , w_36979 );
buf ( w_36977 , \14127_b1 );
not ( w_36977 , w_36980 );
not (  , w_36981 );
and ( w_36980 , w_36981 , \14127_b0 );
or ( \14129_b1 , \14047_b1 , \14128_b1 );
not ( \14128_b1 , w_36982 );
and ( \14129_b0 , \14047_b0 , w_36983 );
and ( w_36982 , w_36983 , \14128_b0 );
or ( \14130_b1 , \7887_b1 , w_36984 );
or ( \14130_b0 , \7887_b0 , \13909_b0 );
not ( \13909_b0 , w_36985 );
and ( w_36985 , w_36984 , \13909_b1 );
or ( \14131_b1 , \14130_b1 , w_36987 );
not ( w_36987 , w_36988 );
and ( \14131_b0 , \14130_b0 , w_36989 );
and ( w_36988 ,  , w_36989 );
buf ( w_36987 , \13916_b1 );
not ( w_36987 , w_36990 );
not (  , w_36991 );
and ( w_36990 , w_36991 , \13916_b0 );
or ( \14132_b1 , \14018_b1 , \14131_b1 );
not ( \14131_b1 , w_36992 );
and ( \14132_b0 , \14018_b0 , w_36993 );
and ( w_36992 , w_36993 , \14131_b0 );
or ( \14133_b1 , \8200_b1 , w_36994 );
or ( \14133_b0 , \8200_b0 , \13918_b0 );
not ( \13918_b0 , w_36995 );
and ( w_36995 , w_36994 , \13918_b1 );
or ( \14134_b1 , \14133_b1 , w_36997 );
not ( w_36997 , w_36998 );
and ( \14134_b0 , \14133_b0 , w_36999 );
and ( w_36998 ,  , w_36999 );
buf ( w_36997 , \13921_b1 );
not ( w_36997 , w_37000 );
not (  , w_37001 );
and ( w_37000 , w_37001 , \13921_b0 );
or ( \14135_b1 , \14132_b1 , w_37003 );
not ( w_37003 , w_37004 );
and ( \14135_b0 , \14132_b0 , w_37005 );
and ( w_37004 ,  , w_37005 );
buf ( w_37003 , \14134_b1 );
not ( w_37003 , w_37006 );
not (  , w_37007 );
and ( w_37006 , w_37007 , \14134_b0 );
or ( \14136_b1 , \14022_b1 , w_37008 );
or ( \14136_b0 , \14022_b0 , \14135_b0 );
not ( \14135_b0 , w_37009 );
and ( w_37009 , w_37008 , \14135_b1 );
or ( \14137_b1 , \8521_b1 , w_37010 );
or ( \14137_b0 , \8521_b0 , \13923_b0 );
not ( \13923_b0 , w_37011 );
and ( w_37011 , w_37010 , \13923_b1 );
or ( \14138_b1 , \14137_b1 , w_37013 );
not ( w_37013 , w_37014 );
and ( \14138_b0 , \14137_b0 , w_37015 );
and ( w_37014 ,  , w_37015 );
buf ( w_37013 , \13927_b1 );
not ( w_37013 , w_37016 );
not (  , w_37017 );
and ( w_37016 , w_37017 , \13927_b0 );
or ( \14139_b1 , \14021_b1 , \14138_b1 );
not ( \14138_b1 , w_37018 );
and ( \14139_b0 , \14021_b0 , w_37019 );
and ( w_37018 , w_37019 , \14138_b0 );
or ( \14140_b1 , \8846_b1 , w_37020 );
or ( \14140_b0 , \8846_b0 , \13929_b0 );
not ( \13929_b0 , w_37021 );
and ( w_37021 , w_37020 , \13929_b1 );
or ( \14141_b1 , \14140_b1 , w_37023 );
not ( w_37023 , w_37024 );
and ( \14141_b0 , \14140_b0 , w_37025 );
and ( w_37024 ,  , w_37025 );
buf ( w_37023 , \13932_b1 );
not ( w_37023 , w_37026 );
not (  , w_37027 );
and ( w_37026 , w_37027 , \13932_b0 );
or ( \14142_b1 , \14139_b1 , w_37029 );
not ( w_37029 , w_37030 );
and ( \14142_b0 , \14139_b0 , w_37031 );
and ( w_37030 ,  , w_37031 );
buf ( w_37029 , \14141_b1 );
not ( w_37029 , w_37032 );
not (  , w_37033 );
and ( w_37032 , w_37033 , \14141_b0 );
or ( \14143_b1 , \14136_b1 , w_37035 );
not ( w_37035 , w_37036 );
and ( \14143_b0 , \14136_b0 , w_37037 );
and ( w_37036 ,  , w_37037 );
buf ( w_37035 , \14142_b1 );
not ( w_37035 , w_37038 );
not (  , w_37039 );
and ( w_37038 , w_37039 , \14142_b0 );
or ( \14144_b1 , \14030_b1 , \14143_b1 );
not ( \14143_b1 , w_37040 );
and ( \14144_b0 , \14030_b0 , w_37041 );
and ( w_37040 , w_37041 , \14143_b0 );
or ( \14145_b1 , \9173_b1 , w_37042 );
or ( \14145_b0 , \9173_b0 , \13934_b0 );
not ( \13934_b0 , w_37043 );
and ( w_37043 , w_37042 , \13934_b1 );
or ( \14146_b1 , \14145_b1 , w_37045 );
not ( w_37045 , w_37046 );
and ( \14146_b0 , \14145_b0 , w_37047 );
and ( w_37046 ,  , w_37047 );
buf ( w_37045 , \13939_b1 );
not ( w_37045 , w_37048 );
not (  , w_37049 );
and ( w_37048 , w_37049 , \13939_b0 );
or ( \14147_b1 , \14025_b1 , \14146_b1 );
not ( \14146_b1 , w_37050 );
and ( \14147_b0 , \14025_b0 , w_37051 );
and ( w_37050 , w_37051 , \14146_b0 );
or ( \14148_b1 , \9498_b1 , w_37052 );
or ( \14148_b0 , \9498_b0 , \13941_b0 );
not ( \13941_b0 , w_37053 );
and ( w_37053 , w_37052 , \13941_b1 );
or ( \14149_b1 , \14148_b1 , w_37055 );
not ( w_37055 , w_37056 );
and ( \14149_b0 , \14148_b0 , w_37057 );
and ( w_37056 ,  , w_37057 );
buf ( w_37055 , \13944_b1 );
not ( w_37055 , w_37058 );
not (  , w_37059 );
and ( w_37058 , w_37059 , \13944_b0 );
or ( \14150_b1 , \14147_b1 , w_37061 );
not ( w_37061 , w_37062 );
and ( \14150_b0 , \14147_b0 , w_37063 );
and ( w_37062 ,  , w_37063 );
buf ( w_37061 , \14149_b1 );
not ( w_37061 , w_37064 );
not (  , w_37065 );
and ( w_37064 , w_37065 , \14149_b0 );
or ( \14151_b1 , \14029_b1 , w_37066 );
or ( \14151_b0 , \14029_b0 , \14150_b0 );
not ( \14150_b0 , w_37067 );
and ( w_37067 , w_37066 , \14150_b1 );
or ( \14152_b1 , \9824_b1 , w_37068 );
or ( \14152_b0 , \9824_b0 , \13946_b0 );
not ( \13946_b0 , w_37069 );
and ( w_37069 , w_37068 , \13946_b1 );
or ( \14153_b1 , \14152_b1 , w_37071 );
not ( w_37071 , w_37072 );
and ( \14153_b0 , \14152_b0 , w_37073 );
and ( w_37072 ,  , w_37073 );
buf ( w_37071 , \13950_b1 );
not ( w_37071 , w_37074 );
not (  , w_37075 );
and ( w_37074 , w_37075 , \13950_b0 );
or ( \14154_b1 , \14028_b1 , \14153_b1 );
not ( \14153_b1 , w_37076 );
and ( \14154_b0 , \14028_b0 , w_37077 );
and ( w_37076 , w_37077 , \14153_b0 );
or ( \14155_b1 , \10149_b1 , w_37078 );
or ( \14155_b0 , \10149_b0 , \13952_b0 );
not ( \13952_b0 , w_37079 );
and ( w_37079 , w_37078 , \13952_b1 );
or ( \14156_b1 , \14155_b1 , w_37081 );
not ( w_37081 , w_37082 );
and ( \14156_b0 , \14155_b0 , w_37083 );
and ( w_37082 ,  , w_37083 );
buf ( w_37081 , \13955_b1 );
not ( w_37081 , w_37084 );
not (  , w_37085 );
and ( w_37084 , w_37085 , \13955_b0 );
or ( \14157_b1 , \14154_b1 , w_37087 );
not ( w_37087 , w_37088 );
and ( \14157_b0 , \14154_b0 , w_37089 );
and ( w_37088 ,  , w_37089 );
buf ( w_37087 , \14156_b1 );
not ( w_37087 , w_37090 );
not (  , w_37091 );
and ( w_37090 , w_37091 , \14156_b0 );
or ( \14158_b1 , \14151_b1 , w_37093 );
not ( w_37093 , w_37094 );
and ( \14158_b0 , \14151_b0 , w_37095 );
and ( w_37094 ,  , w_37095 );
buf ( w_37093 , \14157_b1 );
not ( w_37093 , w_37096 );
not (  , w_37097 );
and ( w_37096 , w_37097 , \14157_b0 );
or ( \14159_b1 , \14144_b1 , w_37099 );
not ( w_37099 , w_37100 );
and ( \14159_b0 , \14144_b0 , w_37101 );
and ( w_37100 ,  , w_37101 );
buf ( w_37099 , \14158_b1 );
not ( w_37099 , w_37102 );
not (  , w_37103 );
and ( w_37102 , w_37103 , \14158_b0 );
or ( \14160_b1 , \14046_b1 , w_37104 );
or ( \14160_b0 , \14046_b0 , \14159_b0 );
not ( \14159_b0 , w_37105 );
and ( w_37105 , w_37104 , \14159_b1 );
or ( \14161_b1 , \10477_b1 , w_37106 );
or ( \14161_b0 , \10477_b0 , \13957_b0 );
not ( \13957_b0 , w_37107 );
and ( w_37107 , w_37106 , \13957_b1 );
or ( \14162_b1 , \14161_b1 , w_37109 );
not ( w_37109 , w_37110 );
and ( \14162_b0 , \14161_b0 , w_37111 );
and ( w_37110 ,  , w_37111 );
buf ( w_37109 , \13963_b1 );
not ( w_37109 , w_37112 );
not (  , w_37113 );
and ( w_37112 , w_37113 , \13963_b0 );
or ( \14163_b1 , \14033_b1 , \14162_b1 );
not ( \14162_b1 , w_37114 );
and ( \14163_b0 , \14033_b0 , w_37115 );
and ( w_37114 , w_37115 , \14162_b0 );
or ( \14164_b1 , \10802_b1 , w_37116 );
or ( \14164_b0 , \10802_b0 , \13965_b0 );
not ( \13965_b0 , w_37117 );
and ( w_37117 , w_37116 , \13965_b1 );
or ( \14165_b1 , \14164_b1 , w_37119 );
not ( w_37119 , w_37120 );
and ( \14165_b0 , \14164_b0 , w_37121 );
and ( w_37120 ,  , w_37121 );
buf ( w_37119 , \13968_b1 );
not ( w_37119 , w_37122 );
not (  , w_37123 );
and ( w_37122 , w_37123 , \13968_b0 );
or ( \14166_b1 , \14163_b1 , w_37125 );
not ( w_37125 , w_37126 );
and ( \14166_b0 , \14163_b0 , w_37127 );
and ( w_37126 ,  , w_37127 );
buf ( w_37125 , \14165_b1 );
not ( w_37125 , w_37128 );
not (  , w_37129 );
and ( w_37128 , w_37129 , \14165_b0 );
or ( \14167_b1 , \14037_b1 , w_37130 );
or ( \14167_b0 , \14037_b0 , \14166_b0 );
not ( \14166_b0 , w_37131 );
and ( w_37131 , w_37130 , \14166_b1 );
or ( \14168_b1 , \11128_b1 , w_37132 );
or ( \14168_b0 , \11128_b0 , \13970_b0 );
not ( \13970_b0 , w_37133 );
and ( w_37133 , w_37132 , \13970_b1 );
or ( \14169_b1 , \14168_b1 , w_37135 );
not ( w_37135 , w_37136 );
and ( \14169_b0 , \14168_b0 , w_37137 );
and ( w_37136 ,  , w_37137 );
buf ( w_37135 , \13974_b1 );
not ( w_37135 , w_37138 );
not (  , w_37139 );
and ( w_37138 , w_37139 , \13974_b0 );
or ( \14170_b1 , \14036_b1 , \14169_b1 );
not ( \14169_b1 , w_37140 );
and ( \14170_b0 , \14036_b0 , w_37141 );
and ( w_37140 , w_37141 , \14169_b0 );
or ( \14171_b1 , \11453_b1 , w_37142 );
or ( \14171_b0 , \11453_b0 , \13976_b0 );
not ( \13976_b0 , w_37143 );
and ( w_37143 , w_37142 , \13976_b1 );
or ( \14172_b1 , \14171_b1 , w_37145 );
not ( w_37145 , w_37146 );
and ( \14172_b0 , \14171_b0 , w_37147 );
and ( w_37146 ,  , w_37147 );
buf ( w_37145 , \13979_b1 );
not ( w_37145 , w_37148 );
not (  , w_37149 );
and ( w_37148 , w_37149 , \13979_b0 );
or ( \14173_b1 , \14170_b1 , w_37151 );
not ( w_37151 , w_37152 );
and ( \14173_b0 , \14170_b0 , w_37153 );
and ( w_37152 ,  , w_37153 );
buf ( w_37151 , \14172_b1 );
not ( w_37151 , w_37154 );
not (  , w_37155 );
and ( w_37154 , w_37155 , \14172_b0 );
or ( \14174_b1 , \14167_b1 , w_37157 );
not ( w_37157 , w_37158 );
and ( \14174_b0 , \14167_b0 , w_37159 );
and ( w_37158 ,  , w_37159 );
buf ( w_37157 , \14173_b1 );
not ( w_37157 , w_37160 );
not (  , w_37161 );
and ( w_37160 , w_37161 , \14173_b0 );
or ( \14175_b1 , \14045_b1 , \14174_b1 );
not ( \14174_b1 , w_37162 );
and ( \14175_b0 , \14045_b0 , w_37163 );
and ( w_37162 , w_37163 , \14174_b0 );
or ( \14176_b1 , \11780_b1 , w_37164 );
or ( \14176_b0 , \11780_b0 , \13981_b0 );
not ( \13981_b0 , w_37165 );
and ( w_37165 , w_37164 , \13981_b1 );
or ( \14177_b1 , \14176_b1 , w_37167 );
not ( w_37167 , w_37168 );
and ( \14177_b0 , \14176_b0 , w_37169 );
and ( w_37168 ,  , w_37169 );
buf ( w_37167 , \13986_b1 );
not ( w_37167 , w_37170 );
not (  , w_37171 );
and ( w_37170 , w_37171 , \13986_b0 );
or ( \14178_b1 , \14040_b1 , \14177_b1 );
not ( \14177_b1 , w_37172 );
and ( \14178_b0 , \14040_b0 , w_37173 );
and ( w_37172 , w_37173 , \14177_b0 );
or ( \14179_b1 , \12040_b1 , w_37174 );
or ( \14179_b0 , \12040_b0 , \13988_b0 );
not ( \13988_b0 , w_37175 );
and ( w_37175 , w_37174 , \13988_b1 );
or ( \14180_b1 , \14179_b1 , w_37177 );
not ( w_37177 , w_37178 );
and ( \14180_b0 , \14179_b0 , w_37179 );
and ( w_37178 ,  , w_37179 );
buf ( w_37177 , \13991_b1 );
not ( w_37177 , w_37180 );
not (  , w_37181 );
and ( w_37180 , w_37181 , \13991_b0 );
or ( \14181_b1 , \14178_b1 , w_37183 );
not ( w_37183 , w_37184 );
and ( \14181_b0 , \14178_b0 , w_37185 );
and ( w_37184 ,  , w_37185 );
buf ( w_37183 , \14180_b1 );
not ( w_37183 , w_37186 );
not (  , w_37187 );
and ( w_37186 , w_37187 , \14180_b0 );
or ( \14182_b1 , \14044_b1 , w_37188 );
or ( \14182_b0 , \14044_b0 , \14181_b0 );
not ( \14181_b0 , w_37189 );
and ( w_37189 , w_37188 , \14181_b1 );
or ( \14183_b1 , \12149_b1 , w_37190 );
or ( \14183_b0 , \12149_b0 , \13993_b0 );
not ( \13993_b0 , w_37191 );
and ( w_37191 , w_37190 , \13993_b1 );
or ( \14184_b1 , \14183_b1 , w_37193 );
not ( w_37193 , w_37194 );
and ( \14184_b0 , \14183_b0 , w_37195 );
and ( w_37194 ,  , w_37195 );
buf ( w_37193 , \13997_b1 );
not ( w_37193 , w_37196 );
not (  , w_37197 );
and ( w_37196 , w_37197 , \13997_b0 );
or ( \14185_b1 , \14043_b1 , \14184_b1 );
not ( \14184_b1 , w_37198 );
and ( \14185_b0 , \14043_b0 , w_37199 );
and ( w_37198 , w_37199 , \14184_b0 );
or ( \14186_b1 , \12190_b1 , w_37200 );
or ( \14186_b0 , \12190_b0 , \13999_b0 );
not ( \13999_b0 , w_37201 );
and ( w_37201 , w_37200 , \13999_b1 );
or ( \14187_b1 , \14186_b1 , w_37203 );
not ( w_37203 , w_37204 );
and ( \14187_b0 , \14186_b0 , w_37205 );
and ( w_37204 ,  , w_37205 );
buf ( w_37203 , \14002_b1 );
not ( w_37203 , w_37206 );
not (  , w_37207 );
and ( w_37206 , w_37207 , \14002_b0 );
or ( \14188_b1 , \14185_b1 , w_37209 );
not ( w_37209 , w_37210 );
and ( \14188_b0 , \14185_b0 , w_37211 );
and ( w_37210 ,  , w_37211 );
buf ( w_37209 , \14187_b1 );
not ( w_37209 , w_37212 );
not (  , w_37213 );
and ( w_37212 , w_37213 , \14187_b0 );
or ( \14189_b1 , \14182_b1 , w_37215 );
not ( w_37215 , w_37216 );
and ( \14189_b0 , \14182_b0 , w_37217 );
and ( w_37216 ,  , w_37217 );
buf ( w_37215 , \14188_b1 );
not ( w_37215 , w_37218 );
not (  , w_37219 );
and ( w_37218 , w_37219 , \14188_b0 );
or ( \14190_b1 , \14175_b1 , w_37221 );
not ( w_37221 , w_37222 );
and ( \14190_b0 , \14175_b0 , w_37223 );
and ( w_37222 ,  , w_37223 );
buf ( w_37221 , \14189_b1 );
not ( w_37221 , w_37224 );
not (  , w_37225 );
and ( w_37224 , w_37225 , \14189_b0 );
or ( \14191_b1 , \14160_b1 , w_37227 );
not ( w_37227 , w_37228 );
and ( \14191_b0 , \14160_b0 , w_37229 );
and ( w_37228 ,  , w_37229 );
buf ( w_37227 , \14190_b1 );
not ( w_37227 , w_37230 );
not (  , w_37231 );
and ( w_37230 , w_37231 , \14190_b0 );
or ( \14192_b1 , \14129_b1 , w_37233 );
not ( w_37233 , w_37234 );
and ( \14192_b0 , \14129_b0 , w_37235 );
and ( w_37234 ,  , w_37235 );
buf ( w_37233 , \14191_b1 );
not ( w_37233 , w_37236 );
not (  , w_37237 );
and ( w_37236 , w_37237 , \14191_b0 );
buf ( \14193_b1 , \14192_b1 );
not ( \14193_b1 , w_37238 );
not ( \14193_b0 , w_37239 );
and ( w_37238 , w_37239 , \14192_b0 );
or ( \14194_b1 , \14016_b1 , w_37240 );
xor ( \14194_b0 , \14016_b0 , w_37242 );
not ( w_37242 , w_37243 );
and ( w_37243 , w_37240 , w_37241 );
buf ( w_37240 , \14193_b1 );
not ( w_37240 , w_37244 );
not ( w_37241 , w_37245 );
and ( w_37244 , w_37245 , \14193_b0 );
buf ( \14195_b1 , \14194_b1 );
buf ( \14195_b0 , \14194_b0 );
buf ( \14196_b1 , \14195_b1 );
buf ( \14196_b0 , \14195_b0 );
buf ( \14197_b1 , \12190_b1 );
not ( \14197_b1 , w_37246 );
not ( \14197_b0 , w_37247 );
and ( w_37246 , w_37247 , \12190_b0 );
or ( \14198_b1 , \14002_b1 , w_37249 );
not ( w_37249 , w_37250 );
and ( \14198_b0 , \14002_b0 , w_37251 );
and ( w_37250 ,  , w_37251 );
buf ( w_37249 , \14197_b1 );
not ( w_37249 , w_37252 );
not (  , w_37253 );
and ( w_37252 , w_37253 , \14197_b0 );
or ( \14199_b1 , \13511_b1 , w_37255 );
not ( w_37255 , w_37256 );
and ( \14199_b0 , \13511_b0 , w_37257 );
and ( w_37256 ,  , w_37257 );
buf ( w_37255 , \8042_b1 );
not ( w_37255 , w_37258 );
not (  , w_37259 );
and ( w_37258 , w_37259 , \8042_b0 );
or ( \14200_b1 , \8360_b1 , w_37261 );
not ( w_37261 , w_37262 );
and ( \14200_b0 , \8360_b0 , w_37263 );
and ( w_37262 ,  , w_37263 );
buf ( w_37261 , \8683_b1 );
not ( w_37261 , w_37264 );
not (  , w_37265 );
and ( w_37264 , w_37265 , \8683_b0 );
or ( \14201_b1 , \14199_b1 , w_37267 );
not ( w_37267 , w_37268 );
and ( \14201_b0 , \14199_b0 , w_37269 );
and ( w_37268 ,  , w_37269 );
buf ( w_37267 , \14200_b1 );
not ( w_37267 , w_37270 );
not (  , w_37271 );
and ( w_37270 , w_37271 , \14200_b0 );
or ( \14202_b1 , \9008_b1 , w_37273 );
not ( w_37273 , w_37274 );
and ( \14202_b0 , \9008_b0 , w_37275 );
and ( w_37274 ,  , w_37275 );
buf ( w_37273 , \9335_b1 );
not ( w_37273 , w_37276 );
not (  , w_37277 );
and ( w_37276 , w_37277 , \9335_b0 );
or ( \14203_b1 , \9660_b1 , w_37279 );
not ( w_37279 , w_37280 );
and ( \14203_b0 , \9660_b0 , w_37281 );
and ( w_37280 ,  , w_37281 );
buf ( w_37279 , \9986_b1 );
not ( w_37279 , w_37282 );
not (  , w_37283 );
and ( w_37282 , w_37283 , \9986_b0 );
or ( \14204_b1 , \14202_b1 , w_37285 );
not ( w_37285 , w_37286 );
and ( \14204_b0 , \14202_b0 , w_37287 );
and ( w_37286 ,  , w_37287 );
buf ( w_37285 , \14203_b1 );
not ( w_37285 , w_37288 );
not (  , w_37289 );
and ( w_37288 , w_37289 , \14203_b0 );
or ( \14205_b1 , \14201_b1 , w_37291 );
not ( w_37291 , w_37292 );
and ( \14205_b0 , \14201_b0 , w_37293 );
and ( w_37292 ,  , w_37293 );
buf ( w_37291 , \14204_b1 );
not ( w_37291 , w_37294 );
not (  , w_37295 );
and ( w_37294 , w_37295 , \14204_b0 );
or ( \14206_b1 , \10311_b1 , w_37297 );
not ( w_37297 , w_37298 );
and ( \14206_b0 , \10311_b0 , w_37299 );
and ( w_37298 ,  , w_37299 );
buf ( w_37297 , \10639_b1 );
not ( w_37297 , w_37300 );
not (  , w_37301 );
and ( w_37300 , w_37301 , \10639_b0 );
or ( \14207_b1 , \10964_b1 , w_37303 );
not ( w_37303 , w_37304 );
and ( \14207_b0 , \10964_b0 , w_37305 );
and ( w_37304 ,  , w_37305 );
buf ( w_37303 , \11290_b1 );
not ( w_37303 , w_37306 );
not (  , w_37307 );
and ( w_37306 , w_37307 , \11290_b0 );
or ( \14208_b1 , \14206_b1 , w_37309 );
not ( w_37309 , w_37310 );
and ( \14208_b0 , \14206_b0 , w_37311 );
and ( w_37310 ,  , w_37311 );
buf ( w_37309 , \14207_b1 );
not ( w_37309 , w_37312 );
not (  , w_37313 );
and ( w_37312 , w_37313 , \14207_b0 );
or ( \14209_b1 , \11615_b1 , w_37315 );
not ( w_37315 , w_37316 );
and ( \14209_b0 , \11615_b0 , w_37317 );
and ( w_37316 ,  , w_37317 );
buf ( w_37315 , \11942_b1 );
not ( w_37315 , w_37318 );
not (  , w_37319 );
and ( w_37318 , w_37319 , \11942_b0 );
or ( \14210_b1 , \12106_b1 , w_37321 );
not ( w_37321 , w_37322 );
and ( \14210_b0 , \12106_b0 , w_37323 );
and ( w_37322 ,  , w_37323 );
buf ( w_37321 , \12175_b1 );
not ( w_37321 , w_37324 );
not (  , w_37325 );
and ( w_37324 , w_37325 , \12175_b0 );
or ( \14211_b1 , \14209_b1 , w_37327 );
not ( w_37327 , w_37328 );
and ( \14211_b0 , \14209_b0 , w_37329 );
and ( w_37328 ,  , w_37329 );
buf ( w_37327 , \14210_b1 );
not ( w_37327 , w_37330 );
not (  , w_37331 );
and ( w_37330 , w_37331 , \14210_b0 );
or ( \14212_b1 , \14208_b1 , w_37333 );
not ( w_37333 , w_37334 );
and ( \14212_b0 , \14208_b0 , w_37335 );
and ( w_37334 ,  , w_37335 );
buf ( w_37333 , \14211_b1 );
not ( w_37333 , w_37336 );
not (  , w_37337 );
and ( w_37336 , w_37337 , \14211_b0 );
or ( \14213_b1 , \14205_b1 , w_37339 );
not ( w_37339 , w_37340 );
and ( \14213_b0 , \14205_b0 , w_37341 );
and ( w_37340 ,  , w_37341 );
buf ( w_37339 , \14212_b1 );
not ( w_37339 , w_37342 );
not (  , w_37343 );
and ( w_37342 , w_37343 , \14212_b0 );
or ( \14214_b1 , \13766_b1 , w_37345 );
not ( w_37345 , w_37346 );
and ( \14214_b0 , \13766_b0 , w_37347 );
and ( w_37346 ,  , w_37347 );
buf ( w_37345 , \12519_b1 );
not ( w_37345 , w_37348 );
not (  , w_37349 );
and ( w_37348 , w_37349 , \12519_b0 );
or ( \14215_b1 , \12686_b1 , w_37351 );
not ( w_37351 , w_37352 );
and ( \14215_b0 , \12686_b0 , w_37353 );
and ( w_37352 ,  , w_37353 );
buf ( w_37351 , \12874_b1 );
not ( w_37351 , w_37354 );
not (  , w_37355 );
and ( w_37354 , w_37355 , \12874_b0 );
or ( \14216_b1 , \14214_b1 , w_37357 );
not ( w_37357 , w_37358 );
and ( \14216_b0 , \14214_b0 , w_37359 );
and ( w_37358 ,  , w_37359 );
buf ( w_37357 , \14215_b1 );
not ( w_37357 , w_37360 );
not (  , w_37361 );
and ( w_37360 , w_37361 , \14215_b0 );
or ( \14217_b1 , \13081_b1 , w_37363 );
not ( w_37363 , w_37364 );
and ( \14217_b0 , \13081_b0 , w_37365 );
and ( w_37364 ,  , w_37365 );
buf ( w_37363 , \13310_b1 );
not ( w_37363 , w_37366 );
not (  , w_37367 );
and ( w_37366 , w_37367 , \13310_b0 );
or ( \14218_b1 , \13429_b1 , w_37369 );
not ( w_37369 , w_37370 );
and ( \14218_b0 , \13429_b0 , w_37371 );
and ( w_37370 ,  , w_37371 );
buf ( w_37369 , \13489_b1 );
not ( w_37369 , w_37372 );
not (  , w_37373 );
and ( w_37372 , w_37373 , \13489_b0 );
or ( \14219_b1 , \14217_b1 , w_37375 );
not ( w_37375 , w_37376 );
and ( \14219_b0 , \14217_b0 , w_37377 );
and ( w_37376 ,  , w_37377 );
buf ( w_37375 , \14218_b1 );
not ( w_37375 , w_37378 );
not (  , w_37379 );
and ( w_37378 , w_37379 , \14218_b0 );
or ( \14220_b1 , \14216_b1 , w_37381 );
not ( w_37381 , w_37382 );
and ( \14220_b0 , \14216_b0 , w_37383 );
and ( w_37382 ,  , w_37383 );
buf ( w_37381 , \14219_b1 );
not ( w_37381 , w_37384 );
not (  , w_37385 );
and ( w_37384 , w_37385 , \14219_b0 );
or ( \14221_b1 , \13813_b1 , w_37387 );
not ( w_37387 , w_37388 );
and ( \14221_b0 , \13813_b0 , w_37389 );
and ( w_37388 ,  , w_37389 );
buf ( w_37387 , \13614_b1 );
not ( w_37387 , w_37390 );
not (  , w_37391 );
and ( w_37390 , w_37391 , \13614_b0 );
or ( \14222_b1 , \13701_b1 , w_37393 );
not ( w_37393 , w_37394 );
and ( \14222_b0 , \13701_b0 , w_37395 );
and ( w_37394 ,  , w_37395 );
buf ( w_37393 , \13747_b1 );
not ( w_37393 , w_37396 );
not (  , w_37397 );
and ( w_37396 , w_37397 , \13747_b0 );
or ( \14223_b1 , \14221_b1 , w_37399 );
not ( w_37399 , w_37400 );
and ( \14223_b0 , \14221_b0 , w_37401 );
and ( w_37400 ,  , w_37401 );
buf ( w_37399 , \14222_b1 );
not ( w_37399 , w_37402 );
not (  , w_37403 );
and ( w_37402 , w_37403 , \14222_b0 );
or ( \14224_b1 , \13799_b1 , \13829_b1 );
not ( \13829_b1 , w_37404 );
and ( \14224_b0 , \13799_b0 , w_37405 );
and ( w_37404 , w_37405 , \13829_b0 );
or ( \14225_b1 , \14224_b1 , w_37407 );
not ( w_37407 , w_37408 );
and ( \14225_b0 , \14224_b0 , w_37409 );
and ( w_37408 ,  , w_37409 );
buf ( w_37407 , \13835_b1 );
not ( w_37407 , w_37410 );
not (  , w_37411 );
and ( w_37410 , w_37411 , \13835_b0 );
buf ( \14226_b1 , \14225_b1 );
not ( \14226_b1 , w_37412 );
not ( \14226_b0 , w_37413 );
and ( w_37412 , w_37413 , \14225_b0 );
or ( \14227_b1 , \14223_b1 , \14226_b1 );
not ( \14226_b1 , w_37414 );
and ( \14227_b0 , \14223_b0 , w_37415 );
and ( w_37414 , w_37415 , \14226_b0 );
or ( \14228_b1 , \13614_b1 , \13840_b1 );
not ( \13840_b1 , w_37416 );
and ( \14228_b0 , \13614_b0 , w_37417 );
and ( w_37416 , w_37417 , \13840_b0 );
or ( \14229_b1 , \14228_b1 , w_37419 );
not ( w_37419 , w_37420 );
and ( \14229_b0 , \14228_b0 , w_37421 );
and ( w_37420 ,  , w_37421 );
buf ( w_37419 , \13847_b1 );
not ( w_37419 , w_37422 );
not (  , w_37423 );
and ( w_37422 , w_37423 , \13847_b0 );
or ( \14230_b1 , \14222_b1 , w_37424 );
or ( \14230_b0 , \14222_b0 , \14229_b0 );
not ( \14229_b0 , w_37425 );
and ( w_37425 , w_37424 , \14229_b1 );
or ( \14231_b1 , \13747_b1 , \13852_b1 );
not ( \13852_b1 , w_37426 );
and ( \14231_b0 , \13747_b0 , w_37427 );
and ( w_37426 , w_37427 , \13852_b0 );
or ( \14232_b1 , \14231_b1 , w_37429 );
not ( w_37429 , w_37430 );
and ( \14232_b0 , \14231_b0 , w_37431 );
and ( w_37430 ,  , w_37431 );
buf ( w_37429 , \13858_b1 );
not ( w_37429 , w_37432 );
not (  , w_37433 );
and ( w_37432 , w_37433 , \13858_b0 );
or ( \14233_b1 , \14230_b1 , w_37435 );
not ( w_37435 , w_37436 );
and ( \14233_b0 , \14230_b0 , w_37437 );
and ( w_37436 ,  , w_37437 );
buf ( w_37435 , \14232_b1 );
not ( w_37435 , w_37438 );
not (  , w_37439 );
and ( w_37438 , w_37439 , \14232_b0 );
or ( \14234_b1 , \14227_b1 , w_37441 );
not ( w_37441 , w_37442 );
and ( \14234_b0 , \14227_b0 , w_37443 );
and ( w_37442 ,  , w_37443 );
buf ( w_37441 , \14233_b1 );
not ( w_37441 , w_37444 );
not (  , w_37445 );
and ( w_37444 , w_37445 , \14233_b0 );
or ( \14235_b1 , \14220_b1 , w_37446 );
or ( \14235_b0 , \14220_b0 , \14234_b0 );
not ( \14234_b0 , w_37447 );
and ( w_37447 , w_37446 , \14234_b1 );
or ( \14236_b1 , \12519_b1 , \13863_b1 );
not ( \13863_b1 , w_37448 );
and ( \14236_b0 , \12519_b0 , w_37449 );
and ( w_37448 , w_37449 , \13863_b0 );
or ( \14237_b1 , \14236_b1 , w_37451 );
not ( w_37451 , w_37452 );
and ( \14237_b0 , \14236_b0 , w_37453 );
and ( w_37452 ,  , w_37453 );
buf ( w_37451 , \13871_b1 );
not ( w_37451 , w_37454 );
not (  , w_37455 );
and ( w_37454 , w_37455 , \13871_b0 );
or ( \14238_b1 , \14215_b1 , w_37456 );
or ( \14238_b0 , \14215_b0 , \14237_b0 );
not ( \14237_b0 , w_37457 );
and ( w_37457 , w_37456 , \14237_b1 );
or ( \14239_b1 , \12874_b1 , \13876_b1 );
not ( \13876_b1 , w_37458 );
and ( \14239_b0 , \12874_b0 , w_37459 );
and ( w_37458 , w_37459 , \13876_b0 );
or ( \14240_b1 , \14239_b1 , w_37461 );
not ( w_37461 , w_37462 );
and ( \14240_b0 , \14239_b0 , w_37463 );
and ( w_37462 ,  , w_37463 );
buf ( w_37461 , \13882_b1 );
not ( w_37461 , w_37464 );
not (  , w_37465 );
and ( w_37464 , w_37465 , \13882_b0 );
or ( \14241_b1 , \14238_b1 , w_37467 );
not ( w_37467 , w_37468 );
and ( \14241_b0 , \14238_b0 , w_37469 );
and ( w_37468 ,  , w_37469 );
buf ( w_37467 , \14240_b1 );
not ( w_37467 , w_37470 );
not (  , w_37471 );
and ( w_37470 , w_37471 , \14240_b0 );
or ( \14242_b1 , \14219_b1 , \14241_b1 );
not ( \14241_b1 , w_37472 );
and ( \14242_b0 , \14219_b0 , w_37473 );
and ( w_37472 , w_37473 , \14241_b0 );
or ( \14243_b1 , \13310_b1 , \13887_b1 );
not ( \13887_b1 , w_37474 );
and ( \14243_b0 , \13310_b0 , w_37475 );
and ( w_37474 , w_37475 , \13887_b0 );
or ( \14244_b1 , \14243_b1 , w_37477 );
not ( w_37477 , w_37478 );
and ( \14244_b0 , \14243_b0 , w_37479 );
and ( w_37478 ,  , w_37479 );
buf ( w_37477 , \13894_b1 );
not ( w_37477 , w_37480 );
not (  , w_37481 );
and ( w_37480 , w_37481 , \13894_b0 );
or ( \14245_b1 , \14218_b1 , w_37482 );
or ( \14245_b0 , \14218_b0 , \14244_b0 );
not ( \14244_b0 , w_37483 );
and ( w_37483 , w_37482 , \14244_b1 );
or ( \14246_b1 , \13489_b1 , \13899_b1 );
not ( \13899_b1 , w_37484 );
and ( \14246_b0 , \13489_b0 , w_37485 );
and ( w_37484 , w_37485 , \13899_b0 );
or ( \14247_b1 , \14246_b1 , w_37487 );
not ( w_37487 , w_37488 );
and ( \14247_b0 , \14246_b0 , w_37489 );
and ( w_37488 ,  , w_37489 );
buf ( w_37487 , \13905_b1 );
not ( w_37487 , w_37490 );
not (  , w_37491 );
and ( w_37490 , w_37491 , \13905_b0 );
or ( \14248_b1 , \14245_b1 , w_37493 );
not ( w_37493 , w_37494 );
and ( \14248_b0 , \14245_b0 , w_37495 );
and ( w_37494 ,  , w_37495 );
buf ( w_37493 , \14247_b1 );
not ( w_37493 , w_37496 );
not (  , w_37497 );
and ( w_37496 , w_37497 , \14247_b0 );
or ( \14249_b1 , \14242_b1 , w_37499 );
not ( w_37499 , w_37500 );
and ( \14249_b0 , \14242_b0 , w_37501 );
and ( w_37500 ,  , w_37501 );
buf ( w_37499 , \14248_b1 );
not ( w_37499 , w_37502 );
not (  , w_37503 );
and ( w_37502 , w_37503 , \14248_b0 );
or ( \14250_b1 , \14235_b1 , w_37505 );
not ( w_37505 , w_37506 );
and ( \14250_b0 , \14235_b0 , w_37507 );
and ( w_37506 ,  , w_37507 );
buf ( w_37505 , \14249_b1 );
not ( w_37505 , w_37508 );
not (  , w_37509 );
and ( w_37508 , w_37509 , \14249_b0 );
or ( \14251_b1 , \14213_b1 , \14250_b1 );
not ( \14250_b1 , w_37510 );
and ( \14251_b0 , \14213_b0 , w_37511 );
and ( w_37510 , w_37511 , \14250_b0 );
or ( \14252_b1 , \8042_b1 , \13910_b1 );
not ( \13910_b1 , w_37512 );
and ( \14252_b0 , \8042_b0 , w_37513 );
and ( w_37512 , w_37513 , \13910_b0 );
or ( \14253_b1 , \14252_b1 , w_37515 );
not ( w_37515 , w_37516 );
and ( \14253_b0 , \14252_b0 , w_37517 );
and ( w_37516 ,  , w_37517 );
buf ( w_37515 , \13919_b1 );
not ( w_37515 , w_37518 );
not (  , w_37519 );
and ( w_37518 , w_37519 , \13919_b0 );
or ( \14254_b1 , \14200_b1 , w_37520 );
or ( \14254_b0 , \14200_b0 , \14253_b0 );
not ( \14253_b0 , w_37521 );
and ( w_37521 , w_37520 , \14253_b1 );
or ( \14255_b1 , \8683_b1 , \13924_b1 );
not ( \13924_b1 , w_37522 );
and ( \14255_b0 , \8683_b0 , w_37523 );
and ( w_37522 , w_37523 , \13924_b0 );
or ( \14256_b1 , \14255_b1 , w_37525 );
not ( w_37525 , w_37526 );
and ( \14256_b0 , \14255_b0 , w_37527 );
and ( w_37526 ,  , w_37527 );
buf ( w_37525 , \13930_b1 );
not ( w_37525 , w_37528 );
not (  , w_37529 );
and ( w_37528 , w_37529 , \13930_b0 );
or ( \14257_b1 , \14254_b1 , w_37531 );
not ( w_37531 , w_37532 );
and ( \14257_b0 , \14254_b0 , w_37533 );
and ( w_37532 ,  , w_37533 );
buf ( w_37531 , \14256_b1 );
not ( w_37531 , w_37534 );
not (  , w_37535 );
and ( w_37534 , w_37535 , \14256_b0 );
or ( \14258_b1 , \14204_b1 , \14257_b1 );
not ( \14257_b1 , w_37536 );
and ( \14258_b0 , \14204_b0 , w_37537 );
and ( w_37536 , w_37537 , \14257_b0 );
or ( \14259_b1 , \9335_b1 , \13935_b1 );
not ( \13935_b1 , w_37538 );
and ( \14259_b0 , \9335_b0 , w_37539 );
and ( w_37538 , w_37539 , \13935_b0 );
or ( \14260_b1 , \14259_b1 , w_37541 );
not ( w_37541 , w_37542 );
and ( \14260_b0 , \14259_b0 , w_37543 );
and ( w_37542 ,  , w_37543 );
buf ( w_37541 , \13942_b1 );
not ( w_37541 , w_37544 );
not (  , w_37545 );
and ( w_37544 , w_37545 , \13942_b0 );
or ( \14261_b1 , \14203_b1 , w_37546 );
or ( \14261_b0 , \14203_b0 , \14260_b0 );
not ( \14260_b0 , w_37547 );
and ( w_37547 , w_37546 , \14260_b1 );
or ( \14262_b1 , \9986_b1 , \13947_b1 );
not ( \13947_b1 , w_37548 );
and ( \14262_b0 , \9986_b0 , w_37549 );
and ( w_37548 , w_37549 , \13947_b0 );
or ( \14263_b1 , \14262_b1 , w_37551 );
not ( w_37551 , w_37552 );
and ( \14263_b0 , \14262_b0 , w_37553 );
and ( w_37552 ,  , w_37553 );
buf ( w_37551 , \13953_b1 );
not ( w_37551 , w_37554 );
not (  , w_37555 );
and ( w_37554 , w_37555 , \13953_b0 );
or ( \14264_b1 , \14261_b1 , w_37557 );
not ( w_37557 , w_37558 );
and ( \14264_b0 , \14261_b0 , w_37559 );
and ( w_37558 ,  , w_37559 );
buf ( w_37557 , \14263_b1 );
not ( w_37557 , w_37560 );
not (  , w_37561 );
and ( w_37560 , w_37561 , \14263_b0 );
or ( \14265_b1 , \14258_b1 , w_37563 );
not ( w_37563 , w_37564 );
and ( \14265_b0 , \14258_b0 , w_37565 );
and ( w_37564 ,  , w_37565 );
buf ( w_37563 , \14264_b1 );
not ( w_37563 , w_37566 );
not (  , w_37567 );
and ( w_37566 , w_37567 , \14264_b0 );
or ( \14266_b1 , \14212_b1 , w_37568 );
or ( \14266_b0 , \14212_b0 , \14265_b0 );
not ( \14265_b0 , w_37569 );
and ( w_37569 , w_37568 , \14265_b1 );
or ( \14267_b1 , \10639_b1 , \13958_b1 );
not ( \13958_b1 , w_37570 );
and ( \14267_b0 , \10639_b0 , w_37571 );
and ( w_37570 , w_37571 , \13958_b0 );
or ( \14268_b1 , \14267_b1 , w_37573 );
not ( w_37573 , w_37574 );
and ( \14268_b0 , \14267_b0 , w_37575 );
and ( w_37574 ,  , w_37575 );
buf ( w_37573 , \13966_b1 );
not ( w_37573 , w_37576 );
not (  , w_37577 );
and ( w_37576 , w_37577 , \13966_b0 );
or ( \14269_b1 , \14207_b1 , w_37578 );
or ( \14269_b0 , \14207_b0 , \14268_b0 );
not ( \14268_b0 , w_37579 );
and ( w_37579 , w_37578 , \14268_b1 );
or ( \14270_b1 , \11290_b1 , \13971_b1 );
not ( \13971_b1 , w_37580 );
and ( \14270_b0 , \11290_b0 , w_37581 );
and ( w_37580 , w_37581 , \13971_b0 );
or ( \14271_b1 , \14270_b1 , w_37583 );
not ( w_37583 , w_37584 );
and ( \14271_b0 , \14270_b0 , w_37585 );
and ( w_37584 ,  , w_37585 );
buf ( w_37583 , \13977_b1 );
not ( w_37583 , w_37586 );
not (  , w_37587 );
and ( w_37586 , w_37587 , \13977_b0 );
or ( \14272_b1 , \14269_b1 , w_37589 );
not ( w_37589 , w_37590 );
and ( \14272_b0 , \14269_b0 , w_37591 );
and ( w_37590 ,  , w_37591 );
buf ( w_37589 , \14271_b1 );
not ( w_37589 , w_37592 );
not (  , w_37593 );
and ( w_37592 , w_37593 , \14271_b0 );
or ( \14273_b1 , \14211_b1 , \14272_b1 );
not ( \14272_b1 , w_37594 );
and ( \14273_b0 , \14211_b0 , w_37595 );
and ( w_37594 , w_37595 , \14272_b0 );
or ( \14274_b1 , \11942_b1 , \13982_b1 );
not ( \13982_b1 , w_37596 );
and ( \14274_b0 , \11942_b0 , w_37597 );
and ( w_37596 , w_37597 , \13982_b0 );
or ( \14275_b1 , \14274_b1 , w_37599 );
not ( w_37599 , w_37600 );
and ( \14275_b0 , \14274_b0 , w_37601 );
and ( w_37600 ,  , w_37601 );
buf ( w_37599 , \13989_b1 );
not ( w_37599 , w_37602 );
not (  , w_37603 );
and ( w_37602 , w_37603 , \13989_b0 );
or ( \14276_b1 , \14210_b1 , w_37604 );
or ( \14276_b0 , \14210_b0 , \14275_b0 );
not ( \14275_b0 , w_37605 );
and ( w_37605 , w_37604 , \14275_b1 );
or ( \14277_b1 , \12175_b1 , \13994_b1 );
not ( \13994_b1 , w_37606 );
and ( \14277_b0 , \12175_b0 , w_37607 );
and ( w_37606 , w_37607 , \13994_b0 );
or ( \14278_b1 , \14277_b1 , w_37609 );
not ( w_37609 , w_37610 );
and ( \14278_b0 , \14277_b0 , w_37611 );
and ( w_37610 ,  , w_37611 );
buf ( w_37609 , \14000_b1 );
not ( w_37609 , w_37612 );
not (  , w_37613 );
and ( w_37612 , w_37613 , \14000_b0 );
or ( \14279_b1 , \14276_b1 , w_37615 );
not ( w_37615 , w_37616 );
and ( \14279_b0 , \14276_b0 , w_37617 );
and ( w_37616 ,  , w_37617 );
buf ( w_37615 , \14278_b1 );
not ( w_37615 , w_37618 );
not (  , w_37619 );
and ( w_37618 , w_37619 , \14278_b0 );
or ( \14280_b1 , \14273_b1 , w_37621 );
not ( w_37621 , w_37622 );
and ( \14280_b0 , \14273_b0 , w_37623 );
and ( w_37622 ,  , w_37623 );
buf ( w_37621 , \14279_b1 );
not ( w_37621 , w_37624 );
not (  , w_37625 );
and ( w_37624 , w_37625 , \14279_b0 );
or ( \14281_b1 , \14266_b1 , w_37627 );
not ( w_37627 , w_37628 );
and ( \14281_b0 , \14266_b0 , w_37629 );
and ( w_37628 ,  , w_37629 );
buf ( w_37627 , \14280_b1 );
not ( w_37627 , w_37630 );
not (  , w_37631 );
and ( w_37630 , w_37631 , \14280_b0 );
or ( \14282_b1 , \14251_b1 , w_37633 );
not ( w_37633 , w_37634 );
and ( \14282_b0 , \14251_b0 , w_37635 );
and ( w_37634 ,  , w_37635 );
buf ( w_37633 , \14281_b1 );
not ( w_37633 , w_37636 );
not (  , w_37637 );
and ( w_37636 , w_37637 , \14281_b0 );
buf ( \14283_b1 , \14282_b1 );
not ( \14283_b1 , w_37638 );
not ( \14283_b0 , w_37639 );
and ( w_37638 , w_37639 , \14282_b0 );
or ( \14284_b1 , \14198_b1 , w_37640 );
xor ( \14284_b0 , \14198_b0 , w_37642 );
not ( w_37642 , w_37643 );
and ( w_37643 , w_37640 , w_37641 );
buf ( w_37640 , \14283_b1 );
not ( w_37640 , w_37644 );
not ( w_37641 , w_37645 );
and ( w_37644 , w_37645 , \14283_b0 );
buf ( \14285_b1 , \14284_b1 );
buf ( \14285_b0 , \14284_b0 );
buf ( \14286_b1 , \14285_b1 );
buf ( \14286_b0 , \14285_b0 );
buf ( \14287_b1 , \12174_b1 );
not ( \14287_b1 , w_37646 );
not ( \14287_b0 , w_37647 );
and ( w_37646 , w_37647 , \12174_b0 );
or ( \14288_b1 , \13999_b1 , w_37649 );
not ( w_37649 , w_37650 );
and ( \14288_b0 , \13999_b0 , w_37651 );
and ( w_37650 ,  , w_37651 );
buf ( w_37649 , \14287_b1 );
not ( w_37649 , w_37652 );
not (  , w_37653 );
and ( w_37652 , w_37653 , \14287_b0 );
or ( \14289_b1 , \14059_b1 , w_37655 );
not ( w_37655 , w_37656 );
and ( \14289_b0 , \14059_b0 , w_37657 );
and ( w_37656 ,  , w_37657 );
buf ( w_37655 , \14017_b1 );
not ( w_37655 , w_37658 );
not (  , w_37659 );
and ( w_37658 , w_37659 , \14017_b0 );
or ( \14290_b1 , \14018_b1 , w_37661 );
not ( w_37661 , w_37662 );
and ( \14290_b0 , \14018_b0 , w_37663 );
and ( w_37662 ,  , w_37663 );
buf ( w_37661 , \14020_b1 );
not ( w_37661 , w_37664 );
not (  , w_37665 );
and ( w_37664 , w_37665 , \14020_b0 );
or ( \14291_b1 , \14289_b1 , w_37667 );
not ( w_37667 , w_37668 );
and ( \14291_b0 , \14289_b0 , w_37669 );
and ( w_37668 ,  , w_37669 );
buf ( w_37667 , \14290_b1 );
not ( w_37667 , w_37670 );
not (  , w_37671 );
and ( w_37670 , w_37671 , \14290_b0 );
or ( \14292_b1 , \14021_b1 , w_37673 );
not ( w_37673 , w_37674 );
and ( \14292_b0 , \14021_b0 , w_37675 );
and ( w_37674 ,  , w_37675 );
buf ( w_37673 , \14024_b1 );
not ( w_37673 , w_37676 );
not (  , w_37677 );
and ( w_37676 , w_37677 , \14024_b0 );
or ( \14293_b1 , \14025_b1 , w_37679 );
not ( w_37679 , w_37680 );
and ( \14293_b0 , \14025_b0 , w_37681 );
and ( w_37680 ,  , w_37681 );
buf ( w_37679 , \14027_b1 );
not ( w_37679 , w_37682 );
not (  , w_37683 );
and ( w_37682 , w_37683 , \14027_b0 );
or ( \14294_b1 , \14292_b1 , w_37685 );
not ( w_37685 , w_37686 );
and ( \14294_b0 , \14292_b0 , w_37687 );
and ( w_37686 ,  , w_37687 );
buf ( w_37685 , \14293_b1 );
not ( w_37685 , w_37688 );
not (  , w_37689 );
and ( w_37688 , w_37689 , \14293_b0 );
or ( \14295_b1 , \14291_b1 , w_37691 );
not ( w_37691 , w_37692 );
and ( \14295_b0 , \14291_b0 , w_37693 );
and ( w_37692 ,  , w_37693 );
buf ( w_37691 , \14294_b1 );
not ( w_37691 , w_37694 );
not (  , w_37695 );
and ( w_37694 , w_37695 , \14294_b0 );
or ( \14296_b1 , \14028_b1 , w_37697 );
not ( w_37697 , w_37698 );
and ( \14296_b0 , \14028_b0 , w_37699 );
and ( w_37698 ,  , w_37699 );
buf ( w_37697 , \14032_b1 );
not ( w_37697 , w_37700 );
not (  , w_37701 );
and ( w_37700 , w_37701 , \14032_b0 );
or ( \14297_b1 , \14033_b1 , w_37703 );
not ( w_37703 , w_37704 );
and ( \14297_b0 , \14033_b0 , w_37705 );
and ( w_37704 ,  , w_37705 );
buf ( w_37703 , \14035_b1 );
not ( w_37703 , w_37706 );
not (  , w_37707 );
and ( w_37706 , w_37707 , \14035_b0 );
or ( \14298_b1 , \14296_b1 , w_37709 );
not ( w_37709 , w_37710 );
and ( \14298_b0 , \14296_b0 , w_37711 );
and ( w_37710 ,  , w_37711 );
buf ( w_37709 , \14297_b1 );
not ( w_37709 , w_37712 );
not (  , w_37713 );
and ( w_37712 , w_37713 , \14297_b0 );
or ( \14299_b1 , \14036_b1 , w_37715 );
not ( w_37715 , w_37716 );
and ( \14299_b0 , \14036_b0 , w_37717 );
and ( w_37716 ,  , w_37717 );
buf ( w_37715 , \14039_b1 );
not ( w_37715 , w_37718 );
not (  , w_37719 );
and ( w_37718 , w_37719 , \14039_b0 );
or ( \14300_b1 , \14040_b1 , w_37721 );
not ( w_37721 , w_37722 );
and ( \14300_b0 , \14040_b0 , w_37723 );
and ( w_37722 ,  , w_37723 );
buf ( w_37721 , \14042_b1 );
not ( w_37721 , w_37724 );
not (  , w_37725 );
and ( w_37724 , w_37725 , \14042_b0 );
or ( \14301_b1 , \14299_b1 , w_37727 );
not ( w_37727 , w_37728 );
and ( \14301_b0 , \14299_b0 , w_37729 );
and ( w_37728 ,  , w_37729 );
buf ( w_37727 , \14300_b1 );
not ( w_37727 , w_37730 );
not (  , w_37731 );
and ( w_37730 , w_37731 , \14300_b0 );
or ( \14302_b1 , \14298_b1 , w_37733 );
not ( w_37733 , w_37734 );
and ( \14302_b0 , \14298_b0 , w_37735 );
and ( w_37734 ,  , w_37735 );
buf ( w_37733 , \14301_b1 );
not ( w_37733 , w_37736 );
not (  , w_37737 );
and ( w_37736 , w_37737 , \14301_b0 );
or ( \14303_b1 , \14295_b1 , w_37739 );
not ( w_37739 , w_37740 );
and ( \14303_b0 , \14295_b0 , w_37741 );
and ( w_37740 ,  , w_37741 );
buf ( w_37739 , \14302_b1 );
not ( w_37739 , w_37742 );
not (  , w_37743 );
and ( w_37742 , w_37743 , \14302_b0 );
or ( \14304_b1 , \14067_b1 , w_37745 );
not ( w_37745 , w_37746 );
and ( \14304_b0 , \14067_b0 , w_37747 );
and ( w_37746 ,  , w_37747 );
buf ( w_37745 , \14048_b1 );
not ( w_37745 , w_37748 );
not (  , w_37749 );
and ( w_37748 , w_37749 , \14048_b0 );
or ( \14305_b1 , \14049_b1 , w_37751 );
not ( w_37751 , w_37752 );
and ( \14305_b0 , \14049_b0 , w_37753 );
and ( w_37752 ,  , w_37753 );
buf ( w_37751 , \14051_b1 );
not ( w_37751 , w_37754 );
not (  , w_37755 );
and ( w_37754 , w_37755 , \14051_b0 );
or ( \14306_b1 , \14304_b1 , w_37757 );
not ( w_37757 , w_37758 );
and ( \14306_b0 , \14304_b0 , w_37759 );
and ( w_37758 ,  , w_37759 );
buf ( w_37757 , \14305_b1 );
not ( w_37757 , w_37760 );
not (  , w_37761 );
and ( w_37760 , w_37761 , \14305_b0 );
or ( \14307_b1 , \14052_b1 , w_37763 );
not ( w_37763 , w_37764 );
and ( \14307_b0 , \14052_b0 , w_37765 );
and ( w_37764 ,  , w_37765 );
buf ( w_37763 , \14055_b1 );
not ( w_37763 , w_37766 );
not (  , w_37767 );
and ( w_37766 , w_37767 , \14055_b0 );
or ( \14308_b1 , \14056_b1 , w_37769 );
not ( w_37769 , w_37770 );
and ( \14308_b0 , \14056_b0 , w_37771 );
and ( w_37770 ,  , w_37771 );
buf ( w_37769 , \14058_b1 );
not ( w_37769 , w_37772 );
not (  , w_37773 );
and ( w_37772 , w_37773 , \14058_b0 );
or ( \14309_b1 , \14307_b1 , w_37775 );
not ( w_37775 , w_37776 );
and ( \14309_b0 , \14307_b0 , w_37777 );
and ( w_37776 ,  , w_37777 );
buf ( w_37775 , \14308_b1 );
not ( w_37775 , w_37778 );
not (  , w_37779 );
and ( w_37778 , w_37779 , \14308_b0 );
or ( \14310_b1 , \14306_b1 , w_37781 );
not ( w_37781 , w_37782 );
and ( \14310_b0 , \14306_b0 , w_37783 );
and ( w_37782 ,  , w_37783 );
buf ( w_37781 , \14309_b1 );
not ( w_37781 , w_37784 );
not (  , w_37785 );
and ( w_37784 , w_37785 , \14309_b0 );
or ( \14311_b1 , \14071_b1 , w_37787 );
not ( w_37787 , w_37788 );
and ( \14311_b0 , \14071_b0 , w_37789 );
and ( w_37788 ,  , w_37789 );
buf ( w_37787 , \14063_b1 );
not ( w_37787 , w_37790 );
not (  , w_37791 );
and ( w_37790 , w_37791 , \14063_b0 );
or ( \14312_b1 , \14064_b1 , w_37793 );
not ( w_37793 , w_37794 );
and ( \14312_b0 , \14064_b0 , w_37795 );
and ( w_37794 ,  , w_37795 );
buf ( w_37793 , \14066_b1 );
not ( w_37793 , w_37796 );
not (  , w_37797 );
and ( w_37796 , w_37797 , \14066_b0 );
or ( \14313_b1 , \14311_b1 , w_37799 );
not ( w_37799 , w_37800 );
and ( \14313_b0 , \14311_b0 , w_37801 );
and ( w_37800 ,  , w_37801 );
buf ( w_37799 , \14312_b1 );
not ( w_37799 , w_37802 );
not (  , w_37803 );
and ( w_37802 , w_37803 , \14312_b0 );
buf ( \14314_b1 , \13826_b1 );
not ( \14314_b1 , w_37804 );
not ( \14314_b0 , w_37805 );
and ( w_37804 , w_37805 , \13826_b0 );
or ( \14315_b1 , \14070_b1 , \14314_b1 );
not ( \14314_b1 , w_37806 );
and ( \14315_b0 , \14070_b0 , w_37807 );
and ( w_37806 , w_37807 , \14314_b0 );
or ( \14316_b1 , \14315_b1 , w_37809 );
not ( w_37809 , w_37810 );
and ( \14316_b0 , \14315_b0 , w_37811 );
and ( w_37810 ,  , w_37811 );
buf ( w_37809 , \14075_b1 );
not ( w_37809 , w_37812 );
not (  , w_37813 );
and ( w_37812 , w_37813 , \14075_b0 );
buf ( \14317_b1 , \14316_b1 );
not ( \14317_b1 , w_37814 );
not ( \14317_b0 , w_37815 );
and ( w_37814 , w_37815 , \14316_b0 );
or ( \14318_b1 , \14313_b1 , \14317_b1 );
not ( \14317_b1 , w_37816 );
and ( \14318_b0 , \14313_b0 , w_37817 );
and ( w_37816 , w_37817 , \14317_b0 );
or ( \14319_b1 , \14063_b1 , \14078_b1 );
not ( \14078_b1 , w_37818 );
and ( \14319_b0 , \14063_b0 , w_37819 );
and ( w_37818 , w_37819 , \14078_b0 );
or ( \14320_b1 , \14319_b1 , w_37821 );
not ( w_37821 , w_37822 );
and ( \14320_b0 , \14319_b0 , w_37823 );
and ( w_37822 ,  , w_37823 );
buf ( w_37821 , \14083_b1 );
not ( w_37821 , w_37824 );
not (  , w_37825 );
and ( w_37824 , w_37825 , \14083_b0 );
or ( \14321_b1 , \14312_b1 , w_37826 );
or ( \14321_b0 , \14312_b0 , \14320_b0 );
not ( \14320_b0 , w_37827 );
and ( w_37827 , w_37826 , \14320_b1 );
or ( \14322_b1 , \14066_b1 , \14086_b1 );
not ( \14086_b1 , w_37828 );
and ( \14322_b0 , \14066_b0 , w_37829 );
and ( w_37828 , w_37829 , \14086_b0 );
or ( \14323_b1 , \14322_b1 , w_37831 );
not ( w_37831 , w_37832 );
and ( \14323_b0 , \14322_b0 , w_37833 );
and ( w_37832 ,  , w_37833 );
buf ( w_37831 , \14090_b1 );
not ( w_37831 , w_37834 );
not (  , w_37835 );
and ( w_37834 , w_37835 , \14090_b0 );
or ( \14324_b1 , \14321_b1 , w_37837 );
not ( w_37837 , w_37838 );
and ( \14324_b0 , \14321_b0 , w_37839 );
and ( w_37838 ,  , w_37839 );
buf ( w_37837 , \14323_b1 );
not ( w_37837 , w_37840 );
not (  , w_37841 );
and ( w_37840 , w_37841 , \14323_b0 );
or ( \14325_b1 , \14318_b1 , w_37843 );
not ( w_37843 , w_37844 );
and ( \14325_b0 , \14318_b0 , w_37845 );
and ( w_37844 ,  , w_37845 );
buf ( w_37843 , \14324_b1 );
not ( w_37843 , w_37846 );
not (  , w_37847 );
and ( w_37846 , w_37847 , \14324_b0 );
or ( \14326_b1 , \14310_b1 , w_37848 );
or ( \14326_b0 , \14310_b0 , \14325_b0 );
not ( \14325_b0 , w_37849 );
and ( w_37849 , w_37848 , \14325_b1 );
or ( \14327_b1 , \14048_b1 , \14093_b1 );
not ( \14093_b1 , w_37850 );
and ( \14327_b0 , \14048_b0 , w_37851 );
and ( w_37850 , w_37851 , \14093_b0 );
or ( \14328_b1 , \14327_b1 , w_37853 );
not ( w_37853 , w_37854 );
and ( \14328_b0 , \14327_b0 , w_37855 );
and ( w_37854 ,  , w_37855 );
buf ( w_37853 , \14099_b1 );
not ( w_37853 , w_37856 );
not (  , w_37857 );
and ( w_37856 , w_37857 , \14099_b0 );
or ( \14329_b1 , \14305_b1 , w_37858 );
or ( \14329_b0 , \14305_b0 , \14328_b0 );
not ( \14328_b0 , w_37859 );
and ( w_37859 , w_37858 , \14328_b1 );
or ( \14330_b1 , \14051_b1 , \14102_b1 );
not ( \14102_b1 , w_37860 );
and ( \14330_b0 , \14051_b0 , w_37861 );
and ( w_37860 , w_37861 , \14102_b0 );
or ( \14331_b1 , \14330_b1 , w_37863 );
not ( w_37863 , w_37864 );
and ( \14331_b0 , \14330_b0 , w_37865 );
and ( w_37864 ,  , w_37865 );
buf ( w_37863 , \14106_b1 );
not ( w_37863 , w_37866 );
not (  , w_37867 );
and ( w_37866 , w_37867 , \14106_b0 );
or ( \14332_b1 , \14329_b1 , w_37869 );
not ( w_37869 , w_37870 );
and ( \14332_b0 , \14329_b0 , w_37871 );
and ( w_37870 ,  , w_37871 );
buf ( w_37869 , \14331_b1 );
not ( w_37869 , w_37872 );
not (  , w_37873 );
and ( w_37872 , w_37873 , \14331_b0 );
or ( \14333_b1 , \14309_b1 , \14332_b1 );
not ( \14332_b1 , w_37874 );
and ( \14333_b0 , \14309_b0 , w_37875 );
and ( w_37874 , w_37875 , \14332_b0 );
or ( \14334_b1 , \14055_b1 , \14109_b1 );
not ( \14109_b1 , w_37876 );
and ( \14334_b0 , \14055_b0 , w_37877 );
and ( w_37876 , w_37877 , \14109_b0 );
or ( \14335_b1 , \14334_b1 , w_37879 );
not ( w_37879 , w_37880 );
and ( \14335_b0 , \14334_b0 , w_37881 );
and ( w_37880 ,  , w_37881 );
buf ( w_37879 , \14114_b1 );
not ( w_37879 , w_37882 );
not (  , w_37883 );
and ( w_37882 , w_37883 , \14114_b0 );
or ( \14336_b1 , \14308_b1 , w_37884 );
or ( \14336_b0 , \14308_b0 , \14335_b0 );
not ( \14335_b0 , w_37885 );
and ( w_37885 , w_37884 , \14335_b1 );
or ( \14337_b1 , \14058_b1 , \14117_b1 );
not ( \14117_b1 , w_37886 );
and ( \14337_b0 , \14058_b0 , w_37887 );
and ( w_37886 , w_37887 , \14117_b0 );
or ( \14338_b1 , \14337_b1 , w_37889 );
not ( w_37889 , w_37890 );
and ( \14338_b0 , \14337_b0 , w_37891 );
and ( w_37890 ,  , w_37891 );
buf ( w_37889 , \14121_b1 );
not ( w_37889 , w_37892 );
not (  , w_37893 );
and ( w_37892 , w_37893 , \14121_b0 );
or ( \14339_b1 , \14336_b1 , w_37895 );
not ( w_37895 , w_37896 );
and ( \14339_b0 , \14336_b0 , w_37897 );
and ( w_37896 ,  , w_37897 );
buf ( w_37895 , \14338_b1 );
not ( w_37895 , w_37898 );
not (  , w_37899 );
and ( w_37898 , w_37899 , \14338_b0 );
or ( \14340_b1 , \14333_b1 , w_37901 );
not ( w_37901 , w_37902 );
and ( \14340_b0 , \14333_b0 , w_37903 );
and ( w_37902 ,  , w_37903 );
buf ( w_37901 , \14339_b1 );
not ( w_37901 , w_37904 );
not (  , w_37905 );
and ( w_37904 , w_37905 , \14339_b0 );
or ( \14341_b1 , \14326_b1 , w_37907 );
not ( w_37907 , w_37908 );
and ( \14341_b0 , \14326_b0 , w_37909 );
and ( w_37908 ,  , w_37909 );
buf ( w_37907 , \14340_b1 );
not ( w_37907 , w_37910 );
not (  , w_37911 );
and ( w_37910 , w_37911 , \14340_b0 );
or ( \14342_b1 , \14303_b1 , \14341_b1 );
not ( \14341_b1 , w_37912 );
and ( \14342_b0 , \14303_b0 , w_37913 );
and ( w_37912 , w_37913 , \14341_b0 );
or ( \14343_b1 , \14017_b1 , \14124_b1 );
not ( \14124_b1 , w_37914 );
and ( \14343_b0 , \14017_b0 , w_37915 );
and ( w_37914 , w_37915 , \14124_b0 );
or ( \14344_b1 , \14343_b1 , w_37917 );
not ( w_37917 , w_37918 );
and ( \14344_b0 , \14343_b0 , w_37919 );
and ( w_37918 ,  , w_37919 );
buf ( w_37917 , \14131_b1 );
not ( w_37917 , w_37920 );
not (  , w_37921 );
and ( w_37920 , w_37921 , \14131_b0 );
or ( \14345_b1 , \14290_b1 , w_37922 );
or ( \14345_b0 , \14290_b0 , \14344_b0 );
not ( \14344_b0 , w_37923 );
and ( w_37923 , w_37922 , \14344_b1 );
or ( \14346_b1 , \14020_b1 , \14134_b1 );
not ( \14134_b1 , w_37924 );
and ( \14346_b0 , \14020_b0 , w_37925 );
and ( w_37924 , w_37925 , \14134_b0 );
or ( \14347_b1 , \14346_b1 , w_37927 );
not ( w_37927 , w_37928 );
and ( \14347_b0 , \14346_b0 , w_37929 );
and ( w_37928 ,  , w_37929 );
buf ( w_37927 , \14138_b1 );
not ( w_37927 , w_37930 );
not (  , w_37931 );
and ( w_37930 , w_37931 , \14138_b0 );
or ( \14348_b1 , \14345_b1 , w_37933 );
not ( w_37933 , w_37934 );
and ( \14348_b0 , \14345_b0 , w_37935 );
and ( w_37934 ,  , w_37935 );
buf ( w_37933 , \14347_b1 );
not ( w_37933 , w_37936 );
not (  , w_37937 );
and ( w_37936 , w_37937 , \14347_b0 );
or ( \14349_b1 , \14294_b1 , \14348_b1 );
not ( \14348_b1 , w_37938 );
and ( \14349_b0 , \14294_b0 , w_37939 );
and ( w_37938 , w_37939 , \14348_b0 );
or ( \14350_b1 , \14024_b1 , \14141_b1 );
not ( \14141_b1 , w_37940 );
and ( \14350_b0 , \14024_b0 , w_37941 );
and ( w_37940 , w_37941 , \14141_b0 );
or ( \14351_b1 , \14350_b1 , w_37943 );
not ( w_37943 , w_37944 );
and ( \14351_b0 , \14350_b0 , w_37945 );
and ( w_37944 ,  , w_37945 );
buf ( w_37943 , \14146_b1 );
not ( w_37943 , w_37946 );
not (  , w_37947 );
and ( w_37946 , w_37947 , \14146_b0 );
or ( \14352_b1 , \14293_b1 , w_37948 );
or ( \14352_b0 , \14293_b0 , \14351_b0 );
not ( \14351_b0 , w_37949 );
and ( w_37949 , w_37948 , \14351_b1 );
or ( \14353_b1 , \14027_b1 , \14149_b1 );
not ( \14149_b1 , w_37950 );
and ( \14353_b0 , \14027_b0 , w_37951 );
and ( w_37950 , w_37951 , \14149_b0 );
or ( \14354_b1 , \14353_b1 , w_37953 );
not ( w_37953 , w_37954 );
and ( \14354_b0 , \14353_b0 , w_37955 );
and ( w_37954 ,  , w_37955 );
buf ( w_37953 , \14153_b1 );
not ( w_37953 , w_37956 );
not (  , w_37957 );
and ( w_37956 , w_37957 , \14153_b0 );
or ( \14355_b1 , \14352_b1 , w_37959 );
not ( w_37959 , w_37960 );
and ( \14355_b0 , \14352_b0 , w_37961 );
and ( w_37960 ,  , w_37961 );
buf ( w_37959 , \14354_b1 );
not ( w_37959 , w_37962 );
not (  , w_37963 );
and ( w_37962 , w_37963 , \14354_b0 );
or ( \14356_b1 , \14349_b1 , w_37965 );
not ( w_37965 , w_37966 );
and ( \14356_b0 , \14349_b0 , w_37967 );
and ( w_37966 ,  , w_37967 );
buf ( w_37965 , \14355_b1 );
not ( w_37965 , w_37968 );
not (  , w_37969 );
and ( w_37968 , w_37969 , \14355_b0 );
or ( \14357_b1 , \14302_b1 , w_37970 );
or ( \14357_b0 , \14302_b0 , \14356_b0 );
not ( \14356_b0 , w_37971 );
and ( w_37971 , w_37970 , \14356_b1 );
or ( \14358_b1 , \14032_b1 , \14156_b1 );
not ( \14156_b1 , w_37972 );
and ( \14358_b0 , \14032_b0 , w_37973 );
and ( w_37972 , w_37973 , \14156_b0 );
or ( \14359_b1 , \14358_b1 , w_37975 );
not ( w_37975 , w_37976 );
and ( \14359_b0 , \14358_b0 , w_37977 );
and ( w_37976 ,  , w_37977 );
buf ( w_37975 , \14162_b1 );
not ( w_37975 , w_37978 );
not (  , w_37979 );
and ( w_37978 , w_37979 , \14162_b0 );
or ( \14360_b1 , \14297_b1 , w_37980 );
or ( \14360_b0 , \14297_b0 , \14359_b0 );
not ( \14359_b0 , w_37981 );
and ( w_37981 , w_37980 , \14359_b1 );
or ( \14361_b1 , \14035_b1 , \14165_b1 );
not ( \14165_b1 , w_37982 );
and ( \14361_b0 , \14035_b0 , w_37983 );
and ( w_37982 , w_37983 , \14165_b0 );
or ( \14362_b1 , \14361_b1 , w_37985 );
not ( w_37985 , w_37986 );
and ( \14362_b0 , \14361_b0 , w_37987 );
and ( w_37986 ,  , w_37987 );
buf ( w_37985 , \14169_b1 );
not ( w_37985 , w_37988 );
not (  , w_37989 );
and ( w_37988 , w_37989 , \14169_b0 );
or ( \14363_b1 , \14360_b1 , w_37991 );
not ( w_37991 , w_37992 );
and ( \14363_b0 , \14360_b0 , w_37993 );
and ( w_37992 ,  , w_37993 );
buf ( w_37991 , \14362_b1 );
not ( w_37991 , w_37994 );
not (  , w_37995 );
and ( w_37994 , w_37995 , \14362_b0 );
or ( \14364_b1 , \14301_b1 , \14363_b1 );
not ( \14363_b1 , w_37996 );
and ( \14364_b0 , \14301_b0 , w_37997 );
and ( w_37996 , w_37997 , \14363_b0 );
or ( \14365_b1 , \14039_b1 , \14172_b1 );
not ( \14172_b1 , w_37998 );
and ( \14365_b0 , \14039_b0 , w_37999 );
and ( w_37998 , w_37999 , \14172_b0 );
or ( \14366_b1 , \14365_b1 , w_38001 );
not ( w_38001 , w_38002 );
and ( \14366_b0 , \14365_b0 , w_38003 );
and ( w_38002 ,  , w_38003 );
buf ( w_38001 , \14177_b1 );
not ( w_38001 , w_38004 );
not (  , w_38005 );
and ( w_38004 , w_38005 , \14177_b0 );
or ( \14367_b1 , \14300_b1 , w_38006 );
or ( \14367_b0 , \14300_b0 , \14366_b0 );
not ( \14366_b0 , w_38007 );
and ( w_38007 , w_38006 , \14366_b1 );
or ( \14368_b1 , \14042_b1 , \14180_b1 );
not ( \14180_b1 , w_38008 );
and ( \14368_b0 , \14042_b0 , w_38009 );
and ( w_38008 , w_38009 , \14180_b0 );
or ( \14369_b1 , \14368_b1 , w_38011 );
not ( w_38011 , w_38012 );
and ( \14369_b0 , \14368_b0 , w_38013 );
and ( w_38012 ,  , w_38013 );
buf ( w_38011 , \14184_b1 );
not ( w_38011 , w_38014 );
not (  , w_38015 );
and ( w_38014 , w_38015 , \14184_b0 );
or ( \14370_b1 , \14367_b1 , w_38017 );
not ( w_38017 , w_38018 );
and ( \14370_b0 , \14367_b0 , w_38019 );
and ( w_38018 ,  , w_38019 );
buf ( w_38017 , \14369_b1 );
not ( w_38017 , w_38020 );
not (  , w_38021 );
and ( w_38020 , w_38021 , \14369_b0 );
or ( \14371_b1 , \14364_b1 , w_38023 );
not ( w_38023 , w_38024 );
and ( \14371_b0 , \14364_b0 , w_38025 );
and ( w_38024 ,  , w_38025 );
buf ( w_38023 , \14370_b1 );
not ( w_38023 , w_38026 );
not (  , w_38027 );
and ( w_38026 , w_38027 , \14370_b0 );
or ( \14372_b1 , \14357_b1 , w_38029 );
not ( w_38029 , w_38030 );
and ( \14372_b0 , \14357_b0 , w_38031 );
and ( w_38030 ,  , w_38031 );
buf ( w_38029 , \14371_b1 );
not ( w_38029 , w_38032 );
not (  , w_38033 );
and ( w_38032 , w_38033 , \14371_b0 );
or ( \14373_b1 , \14342_b1 , w_38035 );
not ( w_38035 , w_38036 );
and ( \14373_b0 , \14342_b0 , w_38037 );
and ( w_38036 ,  , w_38037 );
buf ( w_38035 , \14372_b1 );
not ( w_38035 , w_38038 );
not (  , w_38039 );
and ( w_38038 , w_38039 , \14372_b0 );
buf ( \14374_b1 , \14373_b1 );
not ( \14374_b1 , w_38040 );
not ( \14374_b0 , w_38041 );
and ( w_38040 , w_38041 , \14373_b0 );
or ( \14375_b1 , \14288_b1 , w_38042 );
xor ( \14375_b0 , \14288_b0 , w_38044 );
not ( w_38044 , w_38045 );
and ( w_38045 , w_38042 , w_38043 );
buf ( w_38042 , \14374_b1 );
not ( w_38042 , w_38046 );
not ( w_38043 , w_38047 );
and ( w_38046 , w_38047 , \14374_b0 );
buf ( \14376_b1 , \14375_b1 );
buf ( \14376_b0 , \14375_b0 );
buf ( \14377_b1 , \14376_b1 );
buf ( \14377_b0 , \14376_b0 );
buf ( \14378_b1 , \12149_b1 );
not ( \14378_b1 , w_38048 );
not ( \14378_b0 , w_38049 );
and ( w_38048 , w_38049 , \12149_b0 );
or ( \14379_b1 , \13997_b1 , w_38051 );
not ( w_38051 , w_38052 );
and ( \14379_b0 , \13997_b0 , w_38053 );
and ( w_38052 ,  , w_38053 );
buf ( w_38051 , \14378_b1 );
not ( w_38051 , w_38054 );
not (  , w_38055 );
and ( w_38054 , w_38055 , \14378_b0 );
or ( \14380_b1 , \13512_b1 , w_38057 );
not ( w_38057 , w_38058 );
and ( \14380_b0 , \13512_b0 , w_38059 );
and ( w_38058 ,  , w_38059 );
buf ( w_38057 , \8361_b1 );
not ( w_38057 , w_38060 );
not (  , w_38061 );
and ( w_38060 , w_38061 , \8361_b0 );
or ( \14381_b1 , \9009_b1 , w_38063 );
not ( w_38063 , w_38064 );
and ( \14381_b0 , \9009_b0 , w_38065 );
and ( w_38064 ,  , w_38065 );
buf ( w_38063 , \9661_b1 );
not ( w_38063 , w_38066 );
not (  , w_38067 );
and ( w_38066 , w_38067 , \9661_b0 );
or ( \14382_b1 , \14380_b1 , w_38069 );
not ( w_38069 , w_38070 );
and ( \14382_b0 , \14380_b0 , w_38071 );
and ( w_38070 ,  , w_38071 );
buf ( w_38069 , \14381_b1 );
not ( w_38069 , w_38072 );
not (  , w_38073 );
and ( w_38072 , w_38073 , \14381_b0 );
or ( \14383_b1 , \10312_b1 , w_38075 );
not ( w_38075 , w_38076 );
and ( \14383_b0 , \10312_b0 , w_38077 );
and ( w_38076 ,  , w_38077 );
buf ( w_38075 , \10965_b1 );
not ( w_38075 , w_38078 );
not (  , w_38079 );
and ( w_38078 , w_38079 , \10965_b0 );
or ( \14384_b1 , \11616_b1 , w_38081 );
not ( w_38081 , w_38082 );
and ( \14384_b0 , \11616_b0 , w_38083 );
and ( w_38082 ,  , w_38083 );
buf ( w_38081 , \12107_b1 );
not ( w_38081 , w_38084 );
not (  , w_38085 );
and ( w_38084 , w_38085 , \12107_b0 );
or ( \14385_b1 , \14383_b1 , w_38087 );
not ( w_38087 , w_38088 );
and ( \14385_b0 , \14383_b0 , w_38089 );
and ( w_38088 ,  , w_38089 );
buf ( w_38087 , \14384_b1 );
not ( w_38087 , w_38090 );
not (  , w_38091 );
and ( w_38090 , w_38091 , \14384_b0 );
or ( \14386_b1 , \14382_b1 , w_38093 );
not ( w_38093 , w_38094 );
and ( \14386_b0 , \14382_b0 , w_38095 );
and ( w_38094 ,  , w_38095 );
buf ( w_38093 , \14385_b1 );
not ( w_38093 , w_38096 );
not (  , w_38097 );
and ( w_38096 , w_38097 , \14385_b0 );
or ( \14387_b1 , \13767_b1 , w_38099 );
not ( w_38099 , w_38100 );
and ( \14387_b0 , \13767_b0 , w_38101 );
and ( w_38100 ,  , w_38101 );
buf ( w_38099 , \12687_b1 );
not ( w_38099 , w_38102 );
not (  , w_38103 );
and ( w_38102 , w_38103 , \12687_b0 );
or ( \14388_b1 , \13082_b1 , w_38105 );
not ( w_38105 , w_38106 );
and ( \14388_b0 , \13082_b0 , w_38107 );
and ( w_38106 ,  , w_38107 );
buf ( w_38105 , \13430_b1 );
not ( w_38105 , w_38108 );
not (  , w_38109 );
and ( w_38108 , w_38109 , \13430_b0 );
or ( \14389_b1 , \14387_b1 , w_38111 );
not ( w_38111 , w_38112 );
and ( \14389_b0 , \14387_b0 , w_38113 );
and ( w_38112 ,  , w_38113 );
buf ( w_38111 , \14388_b1 );
not ( w_38111 , w_38114 );
not (  , w_38115 );
and ( w_38114 , w_38115 , \14388_b0 );
or ( \14390_b1 , \13814_b1 , w_38117 );
not ( w_38117 , w_38118 );
and ( \14390_b0 , \13814_b0 , w_38119 );
and ( w_38118 ,  , w_38119 );
buf ( w_38117 , \13702_b1 );
not ( w_38117 , w_38120 );
not (  , w_38121 );
and ( w_38120 , w_38121 , \13702_b0 );
or ( \14391_b1 , \14390_b1 , \13829_b1 );
not ( \13829_b1 , w_38122 );
and ( \14391_b0 , \14390_b0 , w_38123 );
and ( w_38122 , w_38123 , \13829_b0 );
or ( \14392_b1 , \13702_b1 , w_38124 );
or ( \14392_b0 , \13702_b0 , \13841_b0 );
not ( \13841_b0 , w_38125 );
and ( w_38125 , w_38124 , \13841_b1 );
or ( \14393_b1 , \14392_b1 , w_38127 );
not ( w_38127 , w_38128 );
and ( \14393_b0 , \14392_b0 , w_38129 );
and ( w_38128 ,  , w_38129 );
buf ( w_38127 , \13853_b1 );
not ( w_38127 , w_38130 );
not (  , w_38131 );
and ( w_38130 , w_38131 , \13853_b0 );
or ( \14394_b1 , \14391_b1 , w_38133 );
not ( w_38133 , w_38134 );
and ( \14394_b0 , \14391_b0 , w_38135 );
and ( w_38134 ,  , w_38135 );
buf ( w_38133 , \14393_b1 );
not ( w_38133 , w_38136 );
not (  , w_38137 );
and ( w_38136 , w_38137 , \14393_b0 );
or ( \14395_b1 , \14389_b1 , w_38138 );
or ( \14395_b0 , \14389_b0 , \14394_b0 );
not ( \14394_b0 , w_38139 );
and ( w_38139 , w_38138 , \14394_b1 );
or ( \14396_b1 , \12687_b1 , w_38140 );
or ( \14396_b0 , \12687_b0 , \13864_b0 );
not ( \13864_b0 , w_38141 );
and ( w_38141 , w_38140 , \13864_b1 );
or ( \14397_b1 , \14396_b1 , w_38143 );
not ( w_38143 , w_38144 );
and ( \14397_b0 , \14396_b0 , w_38145 );
and ( w_38144 ,  , w_38145 );
buf ( w_38143 , \13877_b1 );
not ( w_38143 , w_38146 );
not (  , w_38147 );
and ( w_38146 , w_38147 , \13877_b0 );
or ( \14398_b1 , \14388_b1 , \14397_b1 );
not ( \14397_b1 , w_38148 );
and ( \14398_b0 , \14388_b0 , w_38149 );
and ( w_38148 , w_38149 , \14397_b0 );
or ( \14399_b1 , \13430_b1 , w_38150 );
or ( \14399_b0 , \13430_b0 , \13888_b0 );
not ( \13888_b0 , w_38151 );
and ( w_38151 , w_38150 , \13888_b1 );
or ( \14400_b1 , \14399_b1 , w_38153 );
not ( w_38153 , w_38154 );
and ( \14400_b0 , \14399_b0 , w_38155 );
and ( w_38154 ,  , w_38155 );
buf ( w_38153 , \13900_b1 );
not ( w_38153 , w_38156 );
not (  , w_38157 );
and ( w_38156 , w_38157 , \13900_b0 );
or ( \14401_b1 , \14398_b1 , w_38159 );
not ( w_38159 , w_38160 );
and ( \14401_b0 , \14398_b0 , w_38161 );
and ( w_38160 ,  , w_38161 );
buf ( w_38159 , \14400_b1 );
not ( w_38159 , w_38162 );
not (  , w_38163 );
and ( w_38162 , w_38163 , \14400_b0 );
or ( \14402_b1 , \14395_b1 , w_38165 );
not ( w_38165 , w_38166 );
and ( \14402_b0 , \14395_b0 , w_38167 );
and ( w_38166 ,  , w_38167 );
buf ( w_38165 , \14401_b1 );
not ( w_38165 , w_38168 );
not (  , w_38169 );
and ( w_38168 , w_38169 , \14401_b0 );
or ( \14403_b1 , \14386_b1 , \14402_b1 );
not ( \14402_b1 , w_38170 );
and ( \14403_b0 , \14386_b0 , w_38171 );
and ( w_38170 , w_38171 , \14402_b0 );
or ( \14404_b1 , \8361_b1 , w_38172 );
or ( \14404_b0 , \8361_b0 , \13911_b0 );
not ( \13911_b0 , w_38173 );
and ( w_38173 , w_38172 , \13911_b1 );
or ( \14405_b1 , \14404_b1 , w_38175 );
not ( w_38175 , w_38176 );
and ( \14405_b0 , \14404_b0 , w_38177 );
and ( w_38176 ,  , w_38177 );
buf ( w_38175 , \13925_b1 );
not ( w_38175 , w_38178 );
not (  , w_38179 );
and ( w_38178 , w_38179 , \13925_b0 );
or ( \14406_b1 , \14381_b1 , \14405_b1 );
not ( \14405_b1 , w_38180 );
and ( \14406_b0 , \14381_b0 , w_38181 );
and ( w_38180 , w_38181 , \14405_b0 );
or ( \14407_b1 , \9661_b1 , w_38182 );
or ( \14407_b0 , \9661_b0 , \13936_b0 );
not ( \13936_b0 , w_38183 );
and ( w_38183 , w_38182 , \13936_b1 );
or ( \14408_b1 , \14407_b1 , w_38185 );
not ( w_38185 , w_38186 );
and ( \14408_b0 , \14407_b0 , w_38187 );
and ( w_38186 ,  , w_38187 );
buf ( w_38185 , \13948_b1 );
not ( w_38185 , w_38188 );
not (  , w_38189 );
and ( w_38188 , w_38189 , \13948_b0 );
or ( \14409_b1 , \14406_b1 , w_38191 );
not ( w_38191 , w_38192 );
and ( \14409_b0 , \14406_b0 , w_38193 );
and ( w_38192 ,  , w_38193 );
buf ( w_38191 , \14408_b1 );
not ( w_38191 , w_38194 );
not (  , w_38195 );
and ( w_38194 , w_38195 , \14408_b0 );
or ( \14410_b1 , \14385_b1 , w_38196 );
or ( \14410_b0 , \14385_b0 , \14409_b0 );
not ( \14409_b0 , w_38197 );
and ( w_38197 , w_38196 , \14409_b1 );
or ( \14411_b1 , \10965_b1 , w_38198 );
or ( \14411_b0 , \10965_b0 , \13959_b0 );
not ( \13959_b0 , w_38199 );
and ( w_38199 , w_38198 , \13959_b1 );
or ( \14412_b1 , \14411_b1 , w_38201 );
not ( w_38201 , w_38202 );
and ( \14412_b0 , \14411_b0 , w_38203 );
and ( w_38202 ,  , w_38203 );
buf ( w_38201 , \13972_b1 );
not ( w_38201 , w_38204 );
not (  , w_38205 );
and ( w_38204 , w_38205 , \13972_b0 );
or ( \14413_b1 , \14384_b1 , \14412_b1 );
not ( \14412_b1 , w_38206 );
and ( \14413_b0 , \14384_b0 , w_38207 );
and ( w_38206 , w_38207 , \14412_b0 );
or ( \14414_b1 , \12107_b1 , w_38208 );
or ( \14414_b0 , \12107_b0 , \13983_b0 );
not ( \13983_b0 , w_38209 );
and ( w_38209 , w_38208 , \13983_b1 );
or ( \14415_b1 , \14414_b1 , w_38211 );
not ( w_38211 , w_38212 );
and ( \14415_b0 , \14414_b0 , w_38213 );
and ( w_38212 ,  , w_38213 );
buf ( w_38211 , \13995_b1 );
not ( w_38211 , w_38214 );
not (  , w_38215 );
and ( w_38214 , w_38215 , \13995_b0 );
or ( \14416_b1 , \14413_b1 , w_38217 );
not ( w_38217 , w_38218 );
and ( \14416_b0 , \14413_b0 , w_38219 );
and ( w_38218 ,  , w_38219 );
buf ( w_38217 , \14415_b1 );
not ( w_38217 , w_38220 );
not (  , w_38221 );
and ( w_38220 , w_38221 , \14415_b0 );
or ( \14417_b1 , \14410_b1 , w_38223 );
not ( w_38223 , w_38224 );
and ( \14417_b0 , \14410_b0 , w_38225 );
and ( w_38224 ,  , w_38225 );
buf ( w_38223 , \14416_b1 );
not ( w_38223 , w_38226 );
not (  , w_38227 );
and ( w_38226 , w_38227 , \14416_b0 );
or ( \14418_b1 , \14403_b1 , w_38229 );
not ( w_38229 , w_38230 );
and ( \14418_b0 , \14403_b0 , w_38231 );
and ( w_38230 ,  , w_38231 );
buf ( w_38229 , \14417_b1 );
not ( w_38229 , w_38232 );
not (  , w_38233 );
and ( w_38232 , w_38233 , \14417_b0 );
buf ( \14419_b1 , \14418_b1 );
not ( \14419_b1 , w_38234 );
not ( \14419_b0 , w_38235 );
and ( w_38234 , w_38235 , \14418_b0 );
or ( \14420_b1 , \14379_b1 , w_38236 );
xor ( \14420_b0 , \14379_b0 , w_38238 );
not ( w_38238 , w_38239 );
and ( w_38239 , w_38236 , w_38237 );
buf ( w_38236 , \14419_b1 );
not ( w_38236 , w_38240 );
not ( w_38237 , w_38241 );
and ( w_38240 , w_38241 , \14419_b0 );
buf ( \14421_b1 , \14420_b1 );
buf ( \14421_b0 , \14420_b0 );
buf ( \14422_b1 , \14421_b1 );
buf ( \14422_b0 , \14421_b0 );
buf ( \14423_b1 , \12105_b1 );
not ( \14423_b1 , w_38242 );
not ( \14423_b0 , w_38243 );
and ( w_38242 , w_38243 , \12105_b0 );
or ( \14424_b1 , \13993_b1 , w_38245 );
not ( w_38245 , w_38246 );
and ( \14424_b0 , \13993_b0 , w_38247 );
and ( w_38246 ,  , w_38247 );
buf ( w_38245 , \14423_b1 );
not ( w_38245 , w_38248 );
not (  , w_38249 );
and ( w_38248 , w_38249 , \14423_b0 );
or ( \14425_b1 , \14060_b1 , w_38251 );
not ( w_38251 , w_38252 );
and ( \14425_b0 , \14060_b0 , w_38253 );
and ( w_38252 ,  , w_38253 );
buf ( w_38251 , \14019_b1 );
not ( w_38251 , w_38254 );
not (  , w_38255 );
and ( w_38254 , w_38255 , \14019_b0 );
or ( \14426_b1 , \14022_b1 , w_38257 );
not ( w_38257 , w_38258 );
and ( \14426_b0 , \14022_b0 , w_38259 );
and ( w_38258 ,  , w_38259 );
buf ( w_38257 , \14026_b1 );
not ( w_38257 , w_38260 );
not (  , w_38261 );
and ( w_38260 , w_38261 , \14026_b0 );
or ( \14427_b1 , \14425_b1 , w_38263 );
not ( w_38263 , w_38264 );
and ( \14427_b0 , \14425_b0 , w_38265 );
and ( w_38264 ,  , w_38265 );
buf ( w_38263 , \14426_b1 );
not ( w_38263 , w_38266 );
not (  , w_38267 );
and ( w_38266 , w_38267 , \14426_b0 );
or ( \14428_b1 , \14029_b1 , w_38269 );
not ( w_38269 , w_38270 );
and ( \14428_b0 , \14029_b0 , w_38271 );
and ( w_38270 ,  , w_38271 );
buf ( w_38269 , \14034_b1 );
not ( w_38269 , w_38272 );
not (  , w_38273 );
and ( w_38272 , w_38273 , \14034_b0 );
or ( \14429_b1 , \14037_b1 , w_38275 );
not ( w_38275 , w_38276 );
and ( \14429_b0 , \14037_b0 , w_38277 );
and ( w_38276 ,  , w_38277 );
buf ( w_38275 , \14041_b1 );
not ( w_38275 , w_38278 );
not (  , w_38279 );
and ( w_38278 , w_38279 , \14041_b0 );
or ( \14430_b1 , \14428_b1 , w_38281 );
not ( w_38281 , w_38282 );
and ( \14430_b0 , \14428_b0 , w_38283 );
and ( w_38282 ,  , w_38283 );
buf ( w_38281 , \14429_b1 );
not ( w_38281 , w_38284 );
not (  , w_38285 );
and ( w_38284 , w_38285 , \14429_b0 );
or ( \14431_b1 , \14427_b1 , w_38287 );
not ( w_38287 , w_38288 );
and ( \14431_b0 , \14427_b0 , w_38289 );
and ( w_38288 ,  , w_38289 );
buf ( w_38287 , \14430_b1 );
not ( w_38287 , w_38290 );
not (  , w_38291 );
and ( w_38290 , w_38291 , \14430_b0 );
or ( \14432_b1 , \14068_b1 , w_38293 );
not ( w_38293 , w_38294 );
and ( \14432_b0 , \14068_b0 , w_38295 );
and ( w_38294 ,  , w_38295 );
buf ( w_38293 , \14050_b1 );
not ( w_38293 , w_38296 );
not (  , w_38297 );
and ( w_38296 , w_38297 , \14050_b0 );
or ( \14433_b1 , \14053_b1 , w_38299 );
not ( w_38299 , w_38300 );
and ( \14433_b0 , \14053_b0 , w_38301 );
and ( w_38300 ,  , w_38301 );
buf ( w_38299 , \14057_b1 );
not ( w_38299 , w_38302 );
not (  , w_38303 );
and ( w_38302 , w_38303 , \14057_b0 );
or ( \14434_b1 , \14432_b1 , w_38305 );
not ( w_38305 , w_38306 );
and ( \14434_b0 , \14432_b0 , w_38307 );
and ( w_38306 ,  , w_38307 );
buf ( w_38305 , \14433_b1 );
not ( w_38305 , w_38308 );
not (  , w_38309 );
and ( w_38308 , w_38309 , \14433_b0 );
or ( \14435_b1 , \14072_b1 , w_38311 );
not ( w_38311 , w_38312 );
and ( \14435_b0 , \14072_b0 , w_38313 );
and ( w_38312 ,  , w_38313 );
buf ( w_38311 , \14065_b1 );
not ( w_38311 , w_38314 );
not (  , w_38315 );
and ( w_38314 , w_38315 , \14065_b0 );
or ( \14436_b1 , \14435_b1 , \14314_b1 );
not ( \14314_b1 , w_38316 );
and ( \14436_b0 , \14435_b0 , w_38317 );
and ( w_38316 , w_38317 , \14314_b0 );
or ( \14437_b1 , \14065_b1 , w_38318 );
or ( \14437_b0 , \14065_b0 , \14079_b0 );
not ( \14079_b0 , w_38319 );
and ( w_38319 , w_38318 , \14079_b1 );
or ( \14438_b1 , \14437_b1 , w_38321 );
not ( w_38321 , w_38322 );
and ( \14438_b0 , \14437_b0 , w_38323 );
and ( w_38322 ,  , w_38323 );
buf ( w_38321 , \14087_b1 );
not ( w_38321 , w_38324 );
not (  , w_38325 );
and ( w_38324 , w_38325 , \14087_b0 );
or ( \14439_b1 , \14436_b1 , w_38327 );
not ( w_38327 , w_38328 );
and ( \14439_b0 , \14436_b0 , w_38329 );
and ( w_38328 ,  , w_38329 );
buf ( w_38327 , \14438_b1 );
not ( w_38327 , w_38330 );
not (  , w_38331 );
and ( w_38330 , w_38331 , \14438_b0 );
or ( \14440_b1 , \14434_b1 , w_38332 );
or ( \14440_b0 , \14434_b0 , \14439_b0 );
not ( \14439_b0 , w_38333 );
and ( w_38333 , w_38332 , \14439_b1 );
or ( \14441_b1 , \14050_b1 , w_38334 );
or ( \14441_b0 , \14050_b0 , \14094_b0 );
not ( \14094_b0 , w_38335 );
and ( w_38335 , w_38334 , \14094_b1 );
or ( \14442_b1 , \14441_b1 , w_38337 );
not ( w_38337 , w_38338 );
and ( \14442_b0 , \14441_b0 , w_38339 );
and ( w_38338 ,  , w_38339 );
buf ( w_38337 , \14103_b1 );
not ( w_38337 , w_38340 );
not (  , w_38341 );
and ( w_38340 , w_38341 , \14103_b0 );
or ( \14443_b1 , \14433_b1 , \14442_b1 );
not ( \14442_b1 , w_38342 );
and ( \14443_b0 , \14433_b0 , w_38343 );
and ( w_38342 , w_38343 , \14442_b0 );
or ( \14444_b1 , \14057_b1 , w_38344 );
or ( \14444_b0 , \14057_b0 , \14110_b0 );
not ( \14110_b0 , w_38345 );
and ( w_38345 , w_38344 , \14110_b1 );
or ( \14445_b1 , \14444_b1 , w_38347 );
not ( w_38347 , w_38348 );
and ( \14445_b0 , \14444_b0 , w_38349 );
and ( w_38348 ,  , w_38349 );
buf ( w_38347 , \14118_b1 );
not ( w_38347 , w_38350 );
not (  , w_38351 );
and ( w_38350 , w_38351 , \14118_b0 );
or ( \14446_b1 , \14443_b1 , w_38353 );
not ( w_38353 , w_38354 );
and ( \14446_b0 , \14443_b0 , w_38355 );
and ( w_38354 ,  , w_38355 );
buf ( w_38353 , \14445_b1 );
not ( w_38353 , w_38356 );
not (  , w_38357 );
and ( w_38356 , w_38357 , \14445_b0 );
or ( \14447_b1 , \14440_b1 , w_38359 );
not ( w_38359 , w_38360 );
and ( \14447_b0 , \14440_b0 , w_38361 );
and ( w_38360 ,  , w_38361 );
buf ( w_38359 , \14446_b1 );
not ( w_38359 , w_38362 );
not (  , w_38363 );
and ( w_38362 , w_38363 , \14446_b0 );
or ( \14448_b1 , \14431_b1 , \14447_b1 );
not ( \14447_b1 , w_38364 );
and ( \14448_b0 , \14431_b0 , w_38365 );
and ( w_38364 , w_38365 , \14447_b0 );
or ( \14449_b1 , \14019_b1 , w_38366 );
or ( \14449_b0 , \14019_b0 , \14125_b0 );
not ( \14125_b0 , w_38367 );
and ( w_38367 , w_38366 , \14125_b1 );
or ( \14450_b1 , \14449_b1 , w_38369 );
not ( w_38369 , w_38370 );
and ( \14450_b0 , \14449_b0 , w_38371 );
and ( w_38370 ,  , w_38371 );
buf ( w_38369 , \14135_b1 );
not ( w_38369 , w_38372 );
not (  , w_38373 );
and ( w_38372 , w_38373 , \14135_b0 );
or ( \14451_b1 , \14426_b1 , \14450_b1 );
not ( \14450_b1 , w_38374 );
and ( \14451_b0 , \14426_b0 , w_38375 );
and ( w_38374 , w_38375 , \14450_b0 );
or ( \14452_b1 , \14026_b1 , w_38376 );
or ( \14452_b0 , \14026_b0 , \14142_b0 );
not ( \14142_b0 , w_38377 );
and ( w_38377 , w_38376 , \14142_b1 );
or ( \14453_b1 , \14452_b1 , w_38379 );
not ( w_38379 , w_38380 );
and ( \14453_b0 , \14452_b0 , w_38381 );
and ( w_38380 ,  , w_38381 );
buf ( w_38379 , \14150_b1 );
not ( w_38379 , w_38382 );
not (  , w_38383 );
and ( w_38382 , w_38383 , \14150_b0 );
or ( \14454_b1 , \14451_b1 , w_38385 );
not ( w_38385 , w_38386 );
and ( \14454_b0 , \14451_b0 , w_38387 );
and ( w_38386 ,  , w_38387 );
buf ( w_38385 , \14453_b1 );
not ( w_38385 , w_38388 );
not (  , w_38389 );
and ( w_38388 , w_38389 , \14453_b0 );
or ( \14455_b1 , \14430_b1 , w_38390 );
or ( \14455_b0 , \14430_b0 , \14454_b0 );
not ( \14454_b0 , w_38391 );
and ( w_38391 , w_38390 , \14454_b1 );
or ( \14456_b1 , \14034_b1 , w_38392 );
or ( \14456_b0 , \14034_b0 , \14157_b0 );
not ( \14157_b0 , w_38393 );
and ( w_38393 , w_38392 , \14157_b1 );
or ( \14457_b1 , \14456_b1 , w_38395 );
not ( w_38395 , w_38396 );
and ( \14457_b0 , \14456_b0 , w_38397 );
and ( w_38396 ,  , w_38397 );
buf ( w_38395 , \14166_b1 );
not ( w_38395 , w_38398 );
not (  , w_38399 );
and ( w_38398 , w_38399 , \14166_b0 );
or ( \14458_b1 , \14429_b1 , \14457_b1 );
not ( \14457_b1 , w_38400 );
and ( \14458_b0 , \14429_b0 , w_38401 );
and ( w_38400 , w_38401 , \14457_b0 );
or ( \14459_b1 , \14041_b1 , w_38402 );
or ( \14459_b0 , \14041_b0 , \14173_b0 );
not ( \14173_b0 , w_38403 );
and ( w_38403 , w_38402 , \14173_b1 );
or ( \14460_b1 , \14459_b1 , w_38405 );
not ( w_38405 , w_38406 );
and ( \14460_b0 , \14459_b0 , w_38407 );
and ( w_38406 ,  , w_38407 );
buf ( w_38405 , \14181_b1 );
not ( w_38405 , w_38408 );
not (  , w_38409 );
and ( w_38408 , w_38409 , \14181_b0 );
or ( \14461_b1 , \14458_b1 , w_38411 );
not ( w_38411 , w_38412 );
and ( \14461_b0 , \14458_b0 , w_38413 );
and ( w_38412 ,  , w_38413 );
buf ( w_38411 , \14460_b1 );
not ( w_38411 , w_38414 );
not (  , w_38415 );
and ( w_38414 , w_38415 , \14460_b0 );
or ( \14462_b1 , \14455_b1 , w_38417 );
not ( w_38417 , w_38418 );
and ( \14462_b0 , \14455_b0 , w_38419 );
and ( w_38418 ,  , w_38419 );
buf ( w_38417 , \14461_b1 );
not ( w_38417 , w_38420 );
not (  , w_38421 );
and ( w_38420 , w_38421 , \14461_b0 );
or ( \14463_b1 , \14448_b1 , w_38423 );
not ( w_38423 , w_38424 );
and ( \14463_b0 , \14448_b0 , w_38425 );
and ( w_38424 ,  , w_38425 );
buf ( w_38423 , \14462_b1 );
not ( w_38423 , w_38426 );
not (  , w_38427 );
and ( w_38426 , w_38427 , \14462_b0 );
buf ( \14464_b1 , \14463_b1 );
not ( \14464_b1 , w_38428 );
not ( \14464_b0 , w_38429 );
and ( w_38428 , w_38429 , \14463_b0 );
or ( \14465_b1 , \14424_b1 , w_38430 );
xor ( \14465_b0 , \14424_b0 , w_38432 );
not ( w_38432 , w_38433 );
and ( w_38433 , w_38430 , w_38431 );
buf ( w_38430 , \14464_b1 );
not ( w_38430 , w_38434 );
not ( w_38431 , w_38435 );
and ( w_38434 , w_38435 , \14464_b0 );
buf ( \14466_b1 , \14465_b1 );
buf ( \14466_b0 , \14465_b0 );
buf ( \14467_b1 , \14466_b1 );
buf ( \14467_b0 , \14466_b0 );
buf ( \14468_b1 , \12040_b1 );
not ( \14468_b1 , w_38436 );
not ( \14468_b0 , w_38437 );
and ( w_38436 , w_38437 , \12040_b0 );
or ( \14469_b1 , \13991_b1 , w_38439 );
not ( w_38439 , w_38440 );
and ( \14469_b0 , \13991_b0 , w_38441 );
and ( w_38440 ,  , w_38441 );
buf ( w_38439 , \14468_b1 );
not ( w_38439 , w_38442 );
not (  , w_38443 );
and ( w_38442 , w_38443 , \14468_b0 );
or ( \14470_b1 , \14218_b1 , w_38445 );
not ( w_38445 , w_38446 );
and ( \14470_b0 , \14218_b0 , w_38447 );
and ( w_38446 ,  , w_38447 );
buf ( w_38445 , \14199_b1 );
not ( w_38445 , w_38448 );
not (  , w_38449 );
and ( w_38448 , w_38449 , \14199_b0 );
or ( \14471_b1 , \14200_b1 , w_38451 );
not ( w_38451 , w_38452 );
and ( \14471_b0 , \14200_b0 , w_38453 );
and ( w_38452 ,  , w_38453 );
buf ( w_38451 , \14202_b1 );
not ( w_38451 , w_38454 );
not (  , w_38455 );
and ( w_38454 , w_38455 , \14202_b0 );
or ( \14472_b1 , \14470_b1 , w_38457 );
not ( w_38457 , w_38458 );
and ( \14472_b0 , \14470_b0 , w_38459 );
and ( w_38458 ,  , w_38459 );
buf ( w_38457 , \14471_b1 );
not ( w_38457 , w_38460 );
not (  , w_38461 );
and ( w_38460 , w_38461 , \14471_b0 );
or ( \14473_b1 , \14203_b1 , w_38463 );
not ( w_38463 , w_38464 );
and ( \14473_b0 , \14203_b0 , w_38465 );
and ( w_38464 ,  , w_38465 );
buf ( w_38463 , \14206_b1 );
not ( w_38463 , w_38466 );
not (  , w_38467 );
and ( w_38466 , w_38467 , \14206_b0 );
or ( \14474_b1 , \14207_b1 , w_38469 );
not ( w_38469 , w_38470 );
and ( \14474_b0 , \14207_b0 , w_38471 );
and ( w_38470 ,  , w_38471 );
buf ( w_38469 , \14209_b1 );
not ( w_38469 , w_38472 );
not (  , w_38473 );
and ( w_38472 , w_38473 , \14209_b0 );
or ( \14475_b1 , \14473_b1 , w_38475 );
not ( w_38475 , w_38476 );
and ( \14475_b0 , \14473_b0 , w_38477 );
and ( w_38476 ,  , w_38477 );
buf ( w_38475 , \14474_b1 );
not ( w_38475 , w_38478 );
not (  , w_38479 );
and ( w_38478 , w_38479 , \14474_b0 );
or ( \14476_b1 , \14472_b1 , w_38481 );
not ( w_38481 , w_38482 );
and ( \14476_b0 , \14472_b0 , w_38483 );
and ( w_38482 ,  , w_38483 );
buf ( w_38481 , \14475_b1 );
not ( w_38481 , w_38484 );
not (  , w_38485 );
and ( w_38484 , w_38485 , \14475_b0 );
or ( \14477_b1 , \14222_b1 , w_38487 );
not ( w_38487 , w_38488 );
and ( \14477_b0 , \14222_b0 , w_38489 );
and ( w_38488 ,  , w_38489 );
buf ( w_38487 , \14214_b1 );
not ( w_38487 , w_38490 );
not (  , w_38491 );
and ( w_38490 , w_38491 , \14214_b0 );
or ( \14478_b1 , \14215_b1 , w_38493 );
not ( w_38493 , w_38494 );
and ( \14478_b0 , \14215_b0 , w_38495 );
and ( w_38494 ,  , w_38495 );
buf ( w_38493 , \14217_b1 );
not ( w_38493 , w_38496 );
not (  , w_38497 );
and ( w_38496 , w_38497 , \14217_b0 );
or ( \14479_b1 , \14477_b1 , w_38499 );
not ( w_38499 , w_38500 );
and ( \14479_b0 , \14477_b0 , w_38501 );
and ( w_38500 ,  , w_38501 );
buf ( w_38499 , \14478_b1 );
not ( w_38499 , w_38502 );
not (  , w_38503 );
and ( w_38502 , w_38503 , \14478_b0 );
or ( \14480_b1 , \14221_b1 , w_38504 );
or ( \14480_b0 , \14221_b0 , \14225_b0 );
not ( \14225_b0 , w_38505 );
and ( w_38505 , w_38504 , \14225_b1 );
or ( \14481_b1 , \14480_b1 , w_38507 );
not ( w_38507 , w_38508 );
and ( \14481_b0 , \14480_b0 , w_38509 );
and ( w_38508 ,  , w_38509 );
buf ( w_38507 , \14229_b1 );
not ( w_38507 , w_38510 );
not (  , w_38511 );
and ( w_38510 , w_38511 , \14229_b0 );
buf ( \14482_b1 , \14481_b1 );
not ( \14482_b1 , w_38512 );
not ( \14482_b0 , w_38513 );
and ( w_38512 , w_38513 , \14481_b0 );
or ( \14483_b1 , \14479_b1 , w_38514 );
or ( \14483_b0 , \14479_b0 , \14482_b0 );
not ( \14482_b0 , w_38515 );
and ( w_38515 , w_38514 , \14482_b1 );
or ( \14484_b1 , \14214_b1 , w_38516 );
or ( \14484_b0 , \14214_b0 , \14232_b0 );
not ( \14232_b0 , w_38517 );
and ( w_38517 , w_38516 , \14232_b1 );
or ( \14485_b1 , \14484_b1 , w_38519 );
not ( w_38519 , w_38520 );
and ( \14485_b0 , \14484_b0 , w_38521 );
and ( w_38520 ,  , w_38521 );
buf ( w_38519 , \14237_b1 );
not ( w_38519 , w_38522 );
not (  , w_38523 );
and ( w_38522 , w_38523 , \14237_b0 );
or ( \14486_b1 , \14478_b1 , \14485_b1 );
not ( \14485_b1 , w_38524 );
and ( \14486_b0 , \14478_b0 , w_38525 );
and ( w_38524 , w_38525 , \14485_b0 );
or ( \14487_b1 , \14217_b1 , w_38526 );
or ( \14487_b0 , \14217_b0 , \14240_b0 );
not ( \14240_b0 , w_38527 );
and ( w_38527 , w_38526 , \14240_b1 );
or ( \14488_b1 , \14487_b1 , w_38529 );
not ( w_38529 , w_38530 );
and ( \14488_b0 , \14487_b0 , w_38531 );
and ( w_38530 ,  , w_38531 );
buf ( w_38529 , \14244_b1 );
not ( w_38529 , w_38532 );
not (  , w_38533 );
and ( w_38532 , w_38533 , \14244_b0 );
or ( \14489_b1 , \14486_b1 , w_38535 );
not ( w_38535 , w_38536 );
and ( \14489_b0 , \14486_b0 , w_38537 );
and ( w_38536 ,  , w_38537 );
buf ( w_38535 , \14488_b1 );
not ( w_38535 , w_38538 );
not (  , w_38539 );
and ( w_38538 , w_38539 , \14488_b0 );
or ( \14490_b1 , \14483_b1 , w_38541 );
not ( w_38541 , w_38542 );
and ( \14490_b0 , \14483_b0 , w_38543 );
and ( w_38542 ,  , w_38543 );
buf ( w_38541 , \14489_b1 );
not ( w_38541 , w_38544 );
not (  , w_38545 );
and ( w_38544 , w_38545 , \14489_b0 );
or ( \14491_b1 , \14476_b1 , \14490_b1 );
not ( \14490_b1 , w_38546 );
and ( \14491_b0 , \14476_b0 , w_38547 );
and ( w_38546 , w_38547 , \14490_b0 );
or ( \14492_b1 , \14199_b1 , w_38548 );
or ( \14492_b0 , \14199_b0 , \14247_b0 );
not ( \14247_b0 , w_38549 );
and ( w_38549 , w_38548 , \14247_b1 );
or ( \14493_b1 , \14492_b1 , w_38551 );
not ( w_38551 , w_38552 );
and ( \14493_b0 , \14492_b0 , w_38553 );
and ( w_38552 ,  , w_38553 );
buf ( w_38551 , \14253_b1 );
not ( w_38551 , w_38554 );
not (  , w_38555 );
and ( w_38554 , w_38555 , \14253_b0 );
or ( \14494_b1 , \14471_b1 , \14493_b1 );
not ( \14493_b1 , w_38556 );
and ( \14494_b0 , \14471_b0 , w_38557 );
and ( w_38556 , w_38557 , \14493_b0 );
or ( \14495_b1 , \14202_b1 , w_38558 );
or ( \14495_b0 , \14202_b0 , \14256_b0 );
not ( \14256_b0 , w_38559 );
and ( w_38559 , w_38558 , \14256_b1 );
or ( \14496_b1 , \14495_b1 , w_38561 );
not ( w_38561 , w_38562 );
and ( \14496_b0 , \14495_b0 , w_38563 );
and ( w_38562 ,  , w_38563 );
buf ( w_38561 , \14260_b1 );
not ( w_38561 , w_38564 );
not (  , w_38565 );
and ( w_38564 , w_38565 , \14260_b0 );
or ( \14497_b1 , \14494_b1 , w_38567 );
not ( w_38567 , w_38568 );
and ( \14497_b0 , \14494_b0 , w_38569 );
and ( w_38568 ,  , w_38569 );
buf ( w_38567 , \14496_b1 );
not ( w_38567 , w_38570 );
not (  , w_38571 );
and ( w_38570 , w_38571 , \14496_b0 );
or ( \14498_b1 , \14475_b1 , w_38572 );
or ( \14498_b0 , \14475_b0 , \14497_b0 );
not ( \14497_b0 , w_38573 );
and ( w_38573 , w_38572 , \14497_b1 );
or ( \14499_b1 , \14206_b1 , w_38574 );
or ( \14499_b0 , \14206_b0 , \14263_b0 );
not ( \14263_b0 , w_38575 );
and ( w_38575 , w_38574 , \14263_b1 );
or ( \14500_b1 , \14499_b1 , w_38577 );
not ( w_38577 , w_38578 );
and ( \14500_b0 , \14499_b0 , w_38579 );
and ( w_38578 ,  , w_38579 );
buf ( w_38577 , \14268_b1 );
not ( w_38577 , w_38580 );
not (  , w_38581 );
and ( w_38580 , w_38581 , \14268_b0 );
or ( \14501_b1 , \14474_b1 , \14500_b1 );
not ( \14500_b1 , w_38582 );
and ( \14501_b0 , \14474_b0 , w_38583 );
and ( w_38582 , w_38583 , \14500_b0 );
or ( \14502_b1 , \14209_b1 , w_38584 );
or ( \14502_b0 , \14209_b0 , \14271_b0 );
not ( \14271_b0 , w_38585 );
and ( w_38585 , w_38584 , \14271_b1 );
or ( \14503_b1 , \14502_b1 , w_38587 );
not ( w_38587 , w_38588 );
and ( \14503_b0 , \14502_b0 , w_38589 );
and ( w_38588 ,  , w_38589 );
buf ( w_38587 , \14275_b1 );
not ( w_38587 , w_38590 );
not (  , w_38591 );
and ( w_38590 , w_38591 , \14275_b0 );
or ( \14504_b1 , \14501_b1 , w_38593 );
not ( w_38593 , w_38594 );
and ( \14504_b0 , \14501_b0 , w_38595 );
and ( w_38594 ,  , w_38595 );
buf ( w_38593 , \14503_b1 );
not ( w_38593 , w_38596 );
not (  , w_38597 );
and ( w_38596 , w_38597 , \14503_b0 );
or ( \14505_b1 , \14498_b1 , w_38599 );
not ( w_38599 , w_38600 );
and ( \14505_b0 , \14498_b0 , w_38601 );
and ( w_38600 ,  , w_38601 );
buf ( w_38599 , \14504_b1 );
not ( w_38599 , w_38602 );
not (  , w_38603 );
and ( w_38602 , w_38603 , \14504_b0 );
or ( \14506_b1 , \14491_b1 , w_38605 );
not ( w_38605 , w_38606 );
and ( \14506_b0 , \14491_b0 , w_38607 );
and ( w_38606 ,  , w_38607 );
buf ( w_38605 , \14505_b1 );
not ( w_38605 , w_38608 );
not (  , w_38609 );
and ( w_38608 , w_38609 , \14505_b0 );
buf ( \14507_b1 , \14506_b1 );
not ( \14507_b1 , w_38610 );
not ( \14507_b0 , w_38611 );
and ( w_38610 , w_38611 , \14506_b0 );
or ( \14508_b1 , \14469_b1 , w_38612 );
xor ( \14508_b0 , \14469_b0 , w_38614 );
not ( w_38614 , w_38615 );
and ( w_38615 , w_38612 , w_38613 );
buf ( w_38612 , \14507_b1 );
not ( w_38612 , w_38616 );
not ( w_38613 , w_38617 );
and ( w_38616 , w_38617 , \14507_b0 );
buf ( \14509_b1 , \14508_b1 );
buf ( \14509_b0 , \14508_b0 );
buf ( \14510_b1 , \14509_b1 );
buf ( \14510_b0 , \14509_b0 );
buf ( \14511_b1 , \11941_b1 );
not ( \14511_b1 , w_38618 );
not ( \14511_b0 , w_38619 );
and ( w_38618 , w_38619 , \11941_b0 );
or ( \14512_b1 , \13988_b1 , w_38621 );
not ( w_38621 , w_38622 );
and ( \14512_b0 , \13988_b0 , w_38623 );
and ( w_38622 ,  , w_38623 );
buf ( w_38621 , \14511_b1 );
not ( w_38621 , w_38624 );
not (  , w_38625 );
and ( w_38624 , w_38625 , \14511_b0 );
or ( \14513_b1 , \14308_b1 , w_38627 );
not ( w_38627 , w_38628 );
and ( \14513_b0 , \14308_b0 , w_38629 );
and ( w_38628 ,  , w_38629 );
buf ( w_38627 , \14289_b1 );
not ( w_38627 , w_38630 );
not (  , w_38631 );
and ( w_38630 , w_38631 , \14289_b0 );
or ( \14514_b1 , \14290_b1 , w_38633 );
not ( w_38633 , w_38634 );
and ( \14514_b0 , \14290_b0 , w_38635 );
and ( w_38634 ,  , w_38635 );
buf ( w_38633 , \14292_b1 );
not ( w_38633 , w_38636 );
not (  , w_38637 );
and ( w_38636 , w_38637 , \14292_b0 );
or ( \14515_b1 , \14513_b1 , w_38639 );
not ( w_38639 , w_38640 );
and ( \14515_b0 , \14513_b0 , w_38641 );
and ( w_38640 ,  , w_38641 );
buf ( w_38639 , \14514_b1 );
not ( w_38639 , w_38642 );
not (  , w_38643 );
and ( w_38642 , w_38643 , \14514_b0 );
or ( \14516_b1 , \14293_b1 , w_38645 );
not ( w_38645 , w_38646 );
and ( \14516_b0 , \14293_b0 , w_38647 );
and ( w_38646 ,  , w_38647 );
buf ( w_38645 , \14296_b1 );
not ( w_38645 , w_38648 );
not (  , w_38649 );
and ( w_38648 , w_38649 , \14296_b0 );
or ( \14517_b1 , \14297_b1 , w_38651 );
not ( w_38651 , w_38652 );
and ( \14517_b0 , \14297_b0 , w_38653 );
and ( w_38652 ,  , w_38653 );
buf ( w_38651 , \14299_b1 );
not ( w_38651 , w_38654 );
not (  , w_38655 );
and ( w_38654 , w_38655 , \14299_b0 );
or ( \14518_b1 , \14516_b1 , w_38657 );
not ( w_38657 , w_38658 );
and ( \14518_b0 , \14516_b0 , w_38659 );
and ( w_38658 ,  , w_38659 );
buf ( w_38657 , \14517_b1 );
not ( w_38657 , w_38660 );
not (  , w_38661 );
and ( w_38660 , w_38661 , \14517_b0 );
or ( \14519_b1 , \14515_b1 , w_38663 );
not ( w_38663 , w_38664 );
and ( \14519_b0 , \14515_b0 , w_38665 );
and ( w_38664 ,  , w_38665 );
buf ( w_38663 , \14518_b1 );
not ( w_38663 , w_38666 );
not (  , w_38667 );
and ( w_38666 , w_38667 , \14518_b0 );
or ( \14520_b1 , \14312_b1 , w_38669 );
not ( w_38669 , w_38670 );
and ( \14520_b0 , \14312_b0 , w_38671 );
and ( w_38670 ,  , w_38671 );
buf ( w_38669 , \14304_b1 );
not ( w_38669 , w_38672 );
not (  , w_38673 );
and ( w_38672 , w_38673 , \14304_b0 );
or ( \14521_b1 , \14305_b1 , w_38675 );
not ( w_38675 , w_38676 );
and ( \14521_b0 , \14305_b0 , w_38677 );
and ( w_38676 ,  , w_38677 );
buf ( w_38675 , \14307_b1 );
not ( w_38675 , w_38678 );
not (  , w_38679 );
and ( w_38678 , w_38679 , \14307_b0 );
or ( \14522_b1 , \14520_b1 , w_38681 );
not ( w_38681 , w_38682 );
and ( \14522_b0 , \14520_b0 , w_38683 );
and ( w_38682 ,  , w_38683 );
buf ( w_38681 , \14521_b1 );
not ( w_38681 , w_38684 );
not (  , w_38685 );
and ( w_38684 , w_38685 , \14521_b0 );
or ( \14523_b1 , \14311_b1 , w_38686 );
or ( \14523_b0 , \14311_b0 , \14316_b0 );
not ( \14316_b0 , w_38687 );
and ( w_38687 , w_38686 , \14316_b1 );
or ( \14524_b1 , \14523_b1 , w_38689 );
not ( w_38689 , w_38690 );
and ( \14524_b0 , \14523_b0 , w_38691 );
and ( w_38690 ,  , w_38691 );
buf ( w_38689 , \14320_b1 );
not ( w_38689 , w_38692 );
not (  , w_38693 );
and ( w_38692 , w_38693 , \14320_b0 );
buf ( \14525_b1 , \14524_b1 );
not ( \14525_b1 , w_38694 );
not ( \14525_b0 , w_38695 );
and ( w_38694 , w_38695 , \14524_b0 );
or ( \14526_b1 , \14522_b1 , w_38696 );
or ( \14526_b0 , \14522_b0 , \14525_b0 );
not ( \14525_b0 , w_38697 );
and ( w_38697 , w_38696 , \14525_b1 );
or ( \14527_b1 , \14304_b1 , w_38698 );
or ( \14527_b0 , \14304_b0 , \14323_b0 );
not ( \14323_b0 , w_38699 );
and ( w_38699 , w_38698 , \14323_b1 );
or ( \14528_b1 , \14527_b1 , w_38701 );
not ( w_38701 , w_38702 );
and ( \14528_b0 , \14527_b0 , w_38703 );
and ( w_38702 ,  , w_38703 );
buf ( w_38701 , \14328_b1 );
not ( w_38701 , w_38704 );
not (  , w_38705 );
and ( w_38704 , w_38705 , \14328_b0 );
or ( \14529_b1 , \14521_b1 , \14528_b1 );
not ( \14528_b1 , w_38706 );
and ( \14529_b0 , \14521_b0 , w_38707 );
and ( w_38706 , w_38707 , \14528_b0 );
or ( \14530_b1 , \14307_b1 , w_38708 );
or ( \14530_b0 , \14307_b0 , \14331_b0 );
not ( \14331_b0 , w_38709 );
and ( w_38709 , w_38708 , \14331_b1 );
or ( \14531_b1 , \14530_b1 , w_38711 );
not ( w_38711 , w_38712 );
and ( \14531_b0 , \14530_b0 , w_38713 );
and ( w_38712 ,  , w_38713 );
buf ( w_38711 , \14335_b1 );
not ( w_38711 , w_38714 );
not (  , w_38715 );
and ( w_38714 , w_38715 , \14335_b0 );
or ( \14532_b1 , \14529_b1 , w_38717 );
not ( w_38717 , w_38718 );
and ( \14532_b0 , \14529_b0 , w_38719 );
and ( w_38718 ,  , w_38719 );
buf ( w_38717 , \14531_b1 );
not ( w_38717 , w_38720 );
not (  , w_38721 );
and ( w_38720 , w_38721 , \14531_b0 );
or ( \14533_b1 , \14526_b1 , w_38723 );
not ( w_38723 , w_38724 );
and ( \14533_b0 , \14526_b0 , w_38725 );
and ( w_38724 ,  , w_38725 );
buf ( w_38723 , \14532_b1 );
not ( w_38723 , w_38726 );
not (  , w_38727 );
and ( w_38726 , w_38727 , \14532_b0 );
or ( \14534_b1 , \14519_b1 , \14533_b1 );
not ( \14533_b1 , w_38728 );
and ( \14534_b0 , \14519_b0 , w_38729 );
and ( w_38728 , w_38729 , \14533_b0 );
or ( \14535_b1 , \14289_b1 , w_38730 );
or ( \14535_b0 , \14289_b0 , \14338_b0 );
not ( \14338_b0 , w_38731 );
and ( w_38731 , w_38730 , \14338_b1 );
or ( \14536_b1 , \14535_b1 , w_38733 );
not ( w_38733 , w_38734 );
and ( \14536_b0 , \14535_b0 , w_38735 );
and ( w_38734 ,  , w_38735 );
buf ( w_38733 , \14344_b1 );
not ( w_38733 , w_38736 );
not (  , w_38737 );
and ( w_38736 , w_38737 , \14344_b0 );
or ( \14537_b1 , \14514_b1 , \14536_b1 );
not ( \14536_b1 , w_38738 );
and ( \14537_b0 , \14514_b0 , w_38739 );
and ( w_38738 , w_38739 , \14536_b0 );
or ( \14538_b1 , \14292_b1 , w_38740 );
or ( \14538_b0 , \14292_b0 , \14347_b0 );
not ( \14347_b0 , w_38741 );
and ( w_38741 , w_38740 , \14347_b1 );
or ( \14539_b1 , \14538_b1 , w_38743 );
not ( w_38743 , w_38744 );
and ( \14539_b0 , \14538_b0 , w_38745 );
and ( w_38744 ,  , w_38745 );
buf ( w_38743 , \14351_b1 );
not ( w_38743 , w_38746 );
not (  , w_38747 );
and ( w_38746 , w_38747 , \14351_b0 );
or ( \14540_b1 , \14537_b1 , w_38749 );
not ( w_38749 , w_38750 );
and ( \14540_b0 , \14537_b0 , w_38751 );
and ( w_38750 ,  , w_38751 );
buf ( w_38749 , \14539_b1 );
not ( w_38749 , w_38752 );
not (  , w_38753 );
and ( w_38752 , w_38753 , \14539_b0 );
or ( \14541_b1 , \14518_b1 , w_38754 );
or ( \14541_b0 , \14518_b0 , \14540_b0 );
not ( \14540_b0 , w_38755 );
and ( w_38755 , w_38754 , \14540_b1 );
or ( \14542_b1 , \14296_b1 , w_38756 );
or ( \14542_b0 , \14296_b0 , \14354_b0 );
not ( \14354_b0 , w_38757 );
and ( w_38757 , w_38756 , \14354_b1 );
or ( \14543_b1 , \14542_b1 , w_38759 );
not ( w_38759 , w_38760 );
and ( \14543_b0 , \14542_b0 , w_38761 );
and ( w_38760 ,  , w_38761 );
buf ( w_38759 , \14359_b1 );
not ( w_38759 , w_38762 );
not (  , w_38763 );
and ( w_38762 , w_38763 , \14359_b0 );
or ( \14544_b1 , \14517_b1 , \14543_b1 );
not ( \14543_b1 , w_38764 );
and ( \14544_b0 , \14517_b0 , w_38765 );
and ( w_38764 , w_38765 , \14543_b0 );
or ( \14545_b1 , \14299_b1 , w_38766 );
or ( \14545_b0 , \14299_b0 , \14362_b0 );
not ( \14362_b0 , w_38767 );
and ( w_38767 , w_38766 , \14362_b1 );
or ( \14546_b1 , \14545_b1 , w_38769 );
not ( w_38769 , w_38770 );
and ( \14546_b0 , \14545_b0 , w_38771 );
and ( w_38770 ,  , w_38771 );
buf ( w_38769 , \14366_b1 );
not ( w_38769 , w_38772 );
not (  , w_38773 );
and ( w_38772 , w_38773 , \14366_b0 );
or ( \14547_b1 , \14544_b1 , w_38775 );
not ( w_38775 , w_38776 );
and ( \14547_b0 , \14544_b0 , w_38777 );
and ( w_38776 ,  , w_38777 );
buf ( w_38775 , \14546_b1 );
not ( w_38775 , w_38778 );
not (  , w_38779 );
and ( w_38778 , w_38779 , \14546_b0 );
or ( \14548_b1 , \14541_b1 , w_38781 );
not ( w_38781 , w_38782 );
and ( \14548_b0 , \14541_b0 , w_38783 );
and ( w_38782 ,  , w_38783 );
buf ( w_38781 , \14547_b1 );
not ( w_38781 , w_38784 );
not (  , w_38785 );
and ( w_38784 , w_38785 , \14547_b0 );
or ( \14549_b1 , \14534_b1 , w_38787 );
not ( w_38787 , w_38788 );
and ( \14549_b0 , \14534_b0 , w_38789 );
and ( w_38788 ,  , w_38789 );
buf ( w_38787 , \14548_b1 );
not ( w_38787 , w_38790 );
not (  , w_38791 );
and ( w_38790 , w_38791 , \14548_b0 );
buf ( \14550_b1 , \14549_b1 );
not ( \14550_b1 , w_38792 );
not ( \14550_b0 , w_38793 );
and ( w_38792 , w_38793 , \14549_b0 );
or ( \14551_b1 , \14512_b1 , w_38794 );
xor ( \14551_b0 , \14512_b0 , w_38796 );
not ( w_38796 , w_38797 );
and ( w_38797 , w_38794 , w_38795 );
buf ( w_38794 , \14550_b1 );
not ( w_38794 , w_38798 );
not ( w_38795 , w_38799 );
and ( w_38798 , w_38799 , \14550_b0 );
buf ( \14552_b1 , \14551_b1 );
buf ( \14552_b0 , \14551_b0 );
buf ( \14553_b1 , \14552_b1 );
buf ( \14553_b0 , \14552_b0 );
buf ( \14554_b1 , \11780_b1 );
not ( \14554_b1 , w_38800 );
not ( \14554_b0 , w_38801 );
and ( w_38800 , w_38801 , \11780_b0 );
or ( \14555_b1 , \13986_b1 , w_38803 );
not ( w_38803 , w_38804 );
and ( \14555_b0 , \13986_b0 , w_38805 );
and ( w_38804 ,  , w_38805 );
buf ( w_38803 , \14554_b1 );
not ( w_38803 , w_38806 );
not (  , w_38807 );
and ( w_38806 , w_38807 , \14554_b0 );
or ( \14556_b1 , \13513_b1 , w_38809 );
not ( w_38809 , w_38810 );
and ( \14556_b0 , \13513_b0 , w_38811 );
and ( w_38810 ,  , w_38811 );
buf ( w_38809 , \9010_b1 );
not ( w_38809 , w_38812 );
not (  , w_38813 );
and ( w_38812 , w_38813 , \9010_b0 );
or ( \14557_b1 , \10313_b1 , w_38815 );
not ( w_38815 , w_38816 );
and ( \14557_b0 , \10313_b0 , w_38817 );
and ( w_38816 ,  , w_38817 );
buf ( w_38815 , \11617_b1 );
not ( w_38815 , w_38818 );
not (  , w_38819 );
and ( w_38818 , w_38819 , \11617_b0 );
or ( \14558_b1 , \14556_b1 , w_38821 );
not ( w_38821 , w_38822 );
and ( \14558_b0 , \14556_b0 , w_38823 );
and ( w_38822 ,  , w_38823 );
buf ( w_38821 , \14557_b1 );
not ( w_38821 , w_38824 );
not (  , w_38825 );
and ( w_38824 , w_38825 , \14557_b0 );
or ( \14559_b1 , \13768_b1 , w_38827 );
not ( w_38827 , w_38828 );
and ( \14559_b0 , \13768_b0 , w_38829 );
and ( w_38828 ,  , w_38829 );
buf ( w_38827 , \13083_b1 );
not ( w_38827 , w_38830 );
not (  , w_38831 );
and ( w_38830 , w_38831 , \13083_b0 );
buf ( \14560_b1 , \13842_b1 );
not ( \14560_b1 , w_38832 );
not ( \14560_b0 , w_38833 );
and ( w_38832 , w_38833 , \13842_b0 );
or ( \14561_b1 , \14559_b1 , w_38834 );
or ( \14561_b0 , \14559_b0 , \14560_b0 );
not ( \14560_b0 , w_38835 );
and ( w_38835 , w_38834 , \14560_b1 );
or ( \14562_b1 , \13083_b1 , \13865_b1 );
not ( \13865_b1 , w_38836 );
and ( \14562_b0 , \13083_b0 , w_38837 );
and ( w_38836 , w_38837 , \13865_b0 );
or ( \14563_b1 , \14562_b1 , w_38839 );
not ( w_38839 , w_38840 );
and ( \14563_b0 , \14562_b0 , w_38841 );
and ( w_38840 ,  , w_38841 );
buf ( w_38839 , \13889_b1 );
not ( w_38839 , w_38842 );
not (  , w_38843 );
and ( w_38842 , w_38843 , \13889_b0 );
or ( \14564_b1 , \14561_b1 , w_38845 );
not ( w_38845 , w_38846 );
and ( \14564_b0 , \14561_b0 , w_38847 );
and ( w_38846 ,  , w_38847 );
buf ( w_38845 , \14563_b1 );
not ( w_38845 , w_38848 );
not (  , w_38849 );
and ( w_38848 , w_38849 , \14563_b0 );
or ( \14565_b1 , \14558_b1 , \14564_b1 );
not ( \14564_b1 , w_38850 );
and ( \14565_b0 , \14558_b0 , w_38851 );
and ( w_38850 , w_38851 , \14564_b0 );
or ( \14566_b1 , \9010_b1 , \13912_b1 );
not ( \13912_b1 , w_38852 );
and ( \14566_b0 , \9010_b0 , w_38853 );
and ( w_38852 , w_38853 , \13912_b0 );
or ( \14567_b1 , \14566_b1 , w_38855 );
not ( w_38855 , w_38856 );
and ( \14567_b0 , \14566_b0 , w_38857 );
and ( w_38856 ,  , w_38857 );
buf ( w_38855 , \13937_b1 );
not ( w_38855 , w_38858 );
not (  , w_38859 );
and ( w_38858 , w_38859 , \13937_b0 );
or ( \14568_b1 , \14557_b1 , w_38860 );
or ( \14568_b0 , \14557_b0 , \14567_b0 );
not ( \14567_b0 , w_38861 );
and ( w_38861 , w_38860 , \14567_b1 );
or ( \14569_b1 , \11617_b1 , \13960_b1 );
not ( \13960_b1 , w_38862 );
and ( \14569_b0 , \11617_b0 , w_38863 );
and ( w_38862 , w_38863 , \13960_b0 );
or ( \14570_b1 , \14569_b1 , w_38865 );
not ( w_38865 , w_38866 );
and ( \14570_b0 , \14569_b0 , w_38867 );
and ( w_38866 ,  , w_38867 );
buf ( w_38865 , \13984_b1 );
not ( w_38865 , w_38868 );
not (  , w_38869 );
and ( w_38868 , w_38869 , \13984_b0 );
or ( \14571_b1 , \14568_b1 , w_38871 );
not ( w_38871 , w_38872 );
and ( \14571_b0 , \14568_b0 , w_38873 );
and ( w_38872 ,  , w_38873 );
buf ( w_38871 , \14570_b1 );
not ( w_38871 , w_38874 );
not (  , w_38875 );
and ( w_38874 , w_38875 , \14570_b0 );
or ( \14572_b1 , \14565_b1 , w_38877 );
not ( w_38877 , w_38878 );
and ( \14572_b0 , \14565_b0 , w_38879 );
and ( w_38878 ,  , w_38879 );
buf ( w_38877 , \14571_b1 );
not ( w_38877 , w_38880 );
not (  , w_38881 );
and ( w_38880 , w_38881 , \14571_b0 );
buf ( \14573_b1 , \14572_b1 );
not ( \14573_b1 , w_38882 );
not ( \14573_b0 , w_38883 );
and ( w_38882 , w_38883 , \14572_b0 );
or ( \14574_b1 , \14555_b1 , w_38884 );
xor ( \14574_b0 , \14555_b0 , w_38886 );
not ( w_38886 , w_38887 );
and ( w_38887 , w_38884 , w_38885 );
buf ( w_38884 , \14573_b1 );
not ( w_38884 , w_38888 );
not ( w_38885 , w_38889 );
and ( w_38888 , w_38889 , \14573_b0 );
buf ( \14575_b1 , \14574_b1 );
buf ( \14575_b0 , \14574_b0 );
buf ( \14576_b1 , \14575_b1 );
buf ( \14576_b0 , \14575_b0 );
buf ( \14577_b1 , \11614_b1 );
not ( \14577_b1 , w_38890 );
not ( \14577_b0 , w_38891 );
and ( w_38890 , w_38891 , \11614_b0 );
or ( \14578_b1 , \13981_b1 , w_38893 );
not ( w_38893 , w_38894 );
and ( \14578_b0 , \13981_b0 , w_38895 );
and ( w_38894 ,  , w_38895 );
buf ( w_38893 , \14577_b1 );
not ( w_38893 , w_38896 );
not (  , w_38897 );
and ( w_38896 , w_38897 , \14577_b0 );
or ( \14579_b1 , \14061_b1 , w_38899 );
not ( w_38899 , w_38900 );
and ( \14579_b0 , \14061_b0 , w_38901 );
and ( w_38900 ,  , w_38901 );
buf ( w_38899 , \14023_b1 );
not ( w_38899 , w_38902 );
not (  , w_38903 );
and ( w_38902 , w_38903 , \14023_b0 );
or ( \14580_b1 , \14030_b1 , w_38905 );
not ( w_38905 , w_38906 );
and ( \14580_b0 , \14030_b0 , w_38907 );
and ( w_38906 ,  , w_38907 );
buf ( w_38905 , \14038_b1 );
not ( w_38905 , w_38908 );
not (  , w_38909 );
and ( w_38908 , w_38909 , \14038_b0 );
or ( \14581_b1 , \14579_b1 , w_38911 );
not ( w_38911 , w_38912 );
and ( \14581_b0 , \14579_b0 , w_38913 );
and ( w_38912 ,  , w_38913 );
buf ( w_38911 , \14580_b1 );
not ( w_38911 , w_38914 );
not (  , w_38915 );
and ( w_38914 , w_38915 , \14580_b0 );
or ( \14582_b1 , \14069_b1 , w_38917 );
not ( w_38917 , w_38918 );
and ( \14582_b0 , \14069_b0 , w_38919 );
and ( w_38918 ,  , w_38919 );
buf ( w_38917 , \14054_b1 );
not ( w_38917 , w_38920 );
not (  , w_38921 );
and ( w_38920 , w_38921 , \14054_b0 );
buf ( \14583_b1 , \14080_b1 );
not ( \14583_b1 , w_38922 );
not ( \14583_b0 , w_38923 );
and ( w_38922 , w_38923 , \14080_b0 );
or ( \14584_b1 , \14582_b1 , w_38924 );
or ( \14584_b0 , \14582_b0 , \14583_b0 );
not ( \14583_b0 , w_38925 );
and ( w_38925 , w_38924 , \14583_b1 );
or ( \14585_b1 , \14054_b1 , \14095_b1 );
not ( \14095_b1 , w_38926 );
and ( \14585_b0 , \14054_b0 , w_38927 );
and ( w_38926 , w_38927 , \14095_b0 );
or ( \14586_b1 , \14585_b1 , w_38929 );
not ( w_38929 , w_38930 );
and ( \14586_b0 , \14585_b0 , w_38931 );
and ( w_38930 ,  , w_38931 );
buf ( w_38929 , \14111_b1 );
not ( w_38929 , w_38932 );
not (  , w_38933 );
and ( w_38932 , w_38933 , \14111_b0 );
or ( \14587_b1 , \14584_b1 , w_38935 );
not ( w_38935 , w_38936 );
and ( \14587_b0 , \14584_b0 , w_38937 );
and ( w_38936 ,  , w_38937 );
buf ( w_38935 , \14586_b1 );
not ( w_38935 , w_38938 );
not (  , w_38939 );
and ( w_38938 , w_38939 , \14586_b0 );
or ( \14588_b1 , \14581_b1 , \14587_b1 );
not ( \14587_b1 , w_38940 );
and ( \14588_b0 , \14581_b0 , w_38941 );
and ( w_38940 , w_38941 , \14587_b0 );
or ( \14589_b1 , \14023_b1 , \14126_b1 );
not ( \14126_b1 , w_38942 );
and ( \14589_b0 , \14023_b0 , w_38943 );
and ( w_38942 , w_38943 , \14126_b0 );
or ( \14590_b1 , \14589_b1 , w_38945 );
not ( w_38945 , w_38946 );
and ( \14590_b0 , \14589_b0 , w_38947 );
and ( w_38946 ,  , w_38947 );
buf ( w_38945 , \14143_b1 );
not ( w_38945 , w_38948 );
not (  , w_38949 );
and ( w_38948 , w_38949 , \14143_b0 );
or ( \14591_b1 , \14580_b1 , w_38950 );
or ( \14591_b0 , \14580_b0 , \14590_b0 );
not ( \14590_b0 , w_38951 );
and ( w_38951 , w_38950 , \14590_b1 );
or ( \14592_b1 , \14038_b1 , \14158_b1 );
not ( \14158_b1 , w_38952 );
and ( \14592_b0 , \14038_b0 , w_38953 );
and ( w_38952 , w_38953 , \14158_b0 );
or ( \14593_b1 , \14592_b1 , w_38955 );
not ( w_38955 , w_38956 );
and ( \14593_b0 , \14592_b0 , w_38957 );
and ( w_38956 ,  , w_38957 );
buf ( w_38955 , \14174_b1 );
not ( w_38955 , w_38958 );
not (  , w_38959 );
and ( w_38958 , w_38959 , \14174_b0 );
or ( \14594_b1 , \14591_b1 , w_38961 );
not ( w_38961 , w_38962 );
and ( \14594_b0 , \14591_b0 , w_38963 );
and ( w_38962 ,  , w_38963 );
buf ( w_38961 , \14593_b1 );
not ( w_38961 , w_38964 );
not (  , w_38965 );
and ( w_38964 , w_38965 , \14593_b0 );
or ( \14595_b1 , \14588_b1 , w_38967 );
not ( w_38967 , w_38968 );
and ( \14595_b0 , \14588_b0 , w_38969 );
and ( w_38968 ,  , w_38969 );
buf ( w_38967 , \14594_b1 );
not ( w_38967 , w_38970 );
not (  , w_38971 );
and ( w_38970 , w_38971 , \14594_b0 );
buf ( \14596_b1 , \14595_b1 );
not ( \14596_b1 , w_38972 );
not ( \14596_b0 , w_38973 );
and ( w_38972 , w_38973 , \14595_b0 );
or ( \14597_b1 , \14578_b1 , w_38974 );
xor ( \14597_b0 , \14578_b0 , w_38976 );
not ( w_38976 , w_38977 );
and ( w_38977 , w_38974 , w_38975 );
buf ( w_38974 , \14596_b1 );
not ( w_38974 , w_38978 );
not ( w_38975 , w_38979 );
and ( w_38978 , w_38979 , \14596_b0 );
buf ( \14598_b1 , \14597_b1 );
buf ( \14598_b0 , \14597_b0 );
buf ( \14599_b1 , \14598_b1 );
buf ( \14599_b0 , \14598_b0 );
buf ( \14600_b1 , \11453_b1 );
not ( \14600_b1 , w_38980 );
not ( \14600_b0 , w_38981 );
and ( w_38980 , w_38981 , \11453_b0 );
or ( \14601_b1 , \13979_b1 , w_38983 );
not ( w_38983 , w_38984 );
and ( \14601_b0 , \13979_b0 , w_38985 );
and ( w_38984 ,  , w_38985 );
buf ( w_38983 , \14600_b1 );
not ( w_38983 , w_38986 );
not (  , w_38987 );
and ( w_38986 , w_38987 , \14600_b0 );
or ( \14602_b1 , \14219_b1 , w_38989 );
not ( w_38989 , w_38990 );
and ( \14602_b0 , \14219_b0 , w_38991 );
and ( w_38990 ,  , w_38991 );
buf ( w_38989 , \14201_b1 );
not ( w_38989 , w_38992 );
not (  , w_38993 );
and ( w_38992 , w_38993 , \14201_b0 );
or ( \14603_b1 , \14204_b1 , w_38995 );
not ( w_38995 , w_38996 );
and ( \14603_b0 , \14204_b0 , w_38997 );
and ( w_38996 ,  , w_38997 );
buf ( w_38995 , \14208_b1 );
not ( w_38995 , w_38998 );
not (  , w_38999 );
and ( w_38998 , w_38999 , \14208_b0 );
or ( \14604_b1 , \14602_b1 , w_39001 );
not ( w_39001 , w_39002 );
and ( \14604_b0 , \14602_b0 , w_39003 );
and ( w_39002 ,  , w_39003 );
buf ( w_39001 , \14603_b1 );
not ( w_39001 , w_39004 );
not (  , w_39005 );
and ( w_39004 , w_39005 , \14603_b0 );
or ( \14605_b1 , \14223_b1 , w_39007 );
not ( w_39007 , w_39008 );
and ( \14605_b0 , \14223_b0 , w_39009 );
and ( w_39008 ,  , w_39009 );
buf ( w_39007 , \14216_b1 );
not ( w_39007 , w_39010 );
not (  , w_39011 );
and ( w_39010 , w_39011 , \14216_b0 );
or ( \14606_b1 , \14605_b1 , w_39012 );
or ( \14606_b0 , \14605_b0 , \14225_b0 );
not ( \14225_b0 , w_39013 );
and ( w_39013 , w_39012 , \14225_b1 );
or ( \14607_b1 , \14216_b1 , \14233_b1 );
not ( \14233_b1 , w_39014 );
and ( \14607_b0 , \14216_b0 , w_39015 );
and ( w_39014 , w_39015 , \14233_b0 );
or ( \14608_b1 , \14607_b1 , w_39017 );
not ( w_39017 , w_39018 );
and ( \14608_b0 , \14607_b0 , w_39019 );
and ( w_39018 ,  , w_39019 );
buf ( w_39017 , \14241_b1 );
not ( w_39017 , w_39020 );
not (  , w_39021 );
and ( w_39020 , w_39021 , \14241_b0 );
or ( \14609_b1 , \14606_b1 , w_39023 );
not ( w_39023 , w_39024 );
and ( \14609_b0 , \14606_b0 , w_39025 );
and ( w_39024 ,  , w_39025 );
buf ( w_39023 , \14608_b1 );
not ( w_39023 , w_39026 );
not (  , w_39027 );
and ( w_39026 , w_39027 , \14608_b0 );
or ( \14610_b1 , \14604_b1 , \14609_b1 );
not ( \14609_b1 , w_39028 );
and ( \14610_b0 , \14604_b0 , w_39029 );
and ( w_39028 , w_39029 , \14609_b0 );
or ( \14611_b1 , \14201_b1 , \14248_b1 );
not ( \14248_b1 , w_39030 );
and ( \14611_b0 , \14201_b0 , w_39031 );
and ( w_39030 , w_39031 , \14248_b0 );
or ( \14612_b1 , \14611_b1 , w_39033 );
not ( w_39033 , w_39034 );
and ( \14612_b0 , \14611_b0 , w_39035 );
and ( w_39034 ,  , w_39035 );
buf ( w_39033 , \14257_b1 );
not ( w_39033 , w_39036 );
not (  , w_39037 );
and ( w_39036 , w_39037 , \14257_b0 );
or ( \14613_b1 , \14603_b1 , w_39038 );
or ( \14613_b0 , \14603_b0 , \14612_b0 );
not ( \14612_b0 , w_39039 );
and ( w_39039 , w_39038 , \14612_b1 );
or ( \14614_b1 , \14208_b1 , \14264_b1 );
not ( \14264_b1 , w_39040 );
and ( \14614_b0 , \14208_b0 , w_39041 );
and ( w_39040 , w_39041 , \14264_b0 );
or ( \14615_b1 , \14614_b1 , w_39043 );
not ( w_39043 , w_39044 );
and ( \14615_b0 , \14614_b0 , w_39045 );
and ( w_39044 ,  , w_39045 );
buf ( w_39043 , \14272_b1 );
not ( w_39043 , w_39046 );
not (  , w_39047 );
and ( w_39046 , w_39047 , \14272_b0 );
or ( \14616_b1 , \14613_b1 , w_39049 );
not ( w_39049 , w_39050 );
and ( \14616_b0 , \14613_b0 , w_39051 );
and ( w_39050 ,  , w_39051 );
buf ( w_39049 , \14615_b1 );
not ( w_39049 , w_39052 );
not (  , w_39053 );
and ( w_39052 , w_39053 , \14615_b0 );
or ( \14617_b1 , \14610_b1 , w_39055 );
not ( w_39055 , w_39056 );
and ( \14617_b0 , \14610_b0 , w_39057 );
and ( w_39056 ,  , w_39057 );
buf ( w_39055 , \14616_b1 );
not ( w_39055 , w_39058 );
not (  , w_39059 );
and ( w_39058 , w_39059 , \14616_b0 );
buf ( \14618_b1 , \14617_b1 );
not ( \14618_b1 , w_39060 );
not ( \14618_b0 , w_39061 );
and ( w_39060 , w_39061 , \14617_b0 );
or ( \14619_b1 , \14601_b1 , w_39062 );
xor ( \14619_b0 , \14601_b0 , w_39064 );
not ( w_39064 , w_39065 );
and ( w_39065 , w_39062 , w_39063 );
buf ( w_39062 , \14618_b1 );
not ( w_39062 , w_39066 );
not ( w_39063 , w_39067 );
and ( w_39066 , w_39067 , \14618_b0 );
buf ( \14620_b1 , \14619_b1 );
buf ( \14620_b0 , \14619_b0 );
buf ( \14621_b1 , \14620_b1 );
buf ( \14621_b0 , \14620_b0 );
buf ( \14622_b1 , \11289_b1 );
not ( \14622_b1 , w_39068 );
not ( \14622_b0 , w_39069 );
and ( w_39068 , w_39069 , \11289_b0 );
or ( \14623_b1 , \13976_b1 , w_39071 );
not ( w_39071 , w_39072 );
and ( \14623_b0 , \13976_b0 , w_39073 );
and ( w_39072 ,  , w_39073 );
buf ( w_39071 , \14622_b1 );
not ( w_39071 , w_39074 );
not (  , w_39075 );
and ( w_39074 , w_39075 , \14622_b0 );
or ( \14624_b1 , \14309_b1 , w_39077 );
not ( w_39077 , w_39078 );
and ( \14624_b0 , \14309_b0 , w_39079 );
and ( w_39078 ,  , w_39079 );
buf ( w_39077 , \14291_b1 );
not ( w_39077 , w_39080 );
not (  , w_39081 );
and ( w_39080 , w_39081 , \14291_b0 );
or ( \14625_b1 , \14294_b1 , w_39083 );
not ( w_39083 , w_39084 );
and ( \14625_b0 , \14294_b0 , w_39085 );
and ( w_39084 ,  , w_39085 );
buf ( w_39083 , \14298_b1 );
not ( w_39083 , w_39086 );
not (  , w_39087 );
and ( w_39086 , w_39087 , \14298_b0 );
or ( \14626_b1 , \14624_b1 , w_39089 );
not ( w_39089 , w_39090 );
and ( \14626_b0 , \14624_b0 , w_39091 );
and ( w_39090 ,  , w_39091 );
buf ( w_39089 , \14625_b1 );
not ( w_39089 , w_39092 );
not (  , w_39093 );
and ( w_39092 , w_39093 , \14625_b0 );
or ( \14627_b1 , \14313_b1 , w_39095 );
not ( w_39095 , w_39096 );
and ( \14627_b0 , \14313_b0 , w_39097 );
and ( w_39096 ,  , w_39097 );
buf ( w_39095 , \14306_b1 );
not ( w_39095 , w_39098 );
not (  , w_39099 );
and ( w_39098 , w_39099 , \14306_b0 );
or ( \14628_b1 , \14627_b1 , w_39100 );
or ( \14628_b0 , \14627_b0 , \14316_b0 );
not ( \14316_b0 , w_39101 );
and ( w_39101 , w_39100 , \14316_b1 );
or ( \14629_b1 , \14306_b1 , \14324_b1 );
not ( \14324_b1 , w_39102 );
and ( \14629_b0 , \14306_b0 , w_39103 );
and ( w_39102 , w_39103 , \14324_b0 );
or ( \14630_b1 , \14629_b1 , w_39105 );
not ( w_39105 , w_39106 );
and ( \14630_b0 , \14629_b0 , w_39107 );
and ( w_39106 ,  , w_39107 );
buf ( w_39105 , \14332_b1 );
not ( w_39105 , w_39108 );
not (  , w_39109 );
and ( w_39108 , w_39109 , \14332_b0 );
or ( \14631_b1 , \14628_b1 , w_39111 );
not ( w_39111 , w_39112 );
and ( \14631_b0 , \14628_b0 , w_39113 );
and ( w_39112 ,  , w_39113 );
buf ( w_39111 , \14630_b1 );
not ( w_39111 , w_39114 );
not (  , w_39115 );
and ( w_39114 , w_39115 , \14630_b0 );
or ( \14632_b1 , \14626_b1 , \14631_b1 );
not ( \14631_b1 , w_39116 );
and ( \14632_b0 , \14626_b0 , w_39117 );
and ( w_39116 , w_39117 , \14631_b0 );
or ( \14633_b1 , \14291_b1 , \14339_b1 );
not ( \14339_b1 , w_39118 );
and ( \14633_b0 , \14291_b0 , w_39119 );
and ( w_39118 , w_39119 , \14339_b0 );
or ( \14634_b1 , \14633_b1 , w_39121 );
not ( w_39121 , w_39122 );
and ( \14634_b0 , \14633_b0 , w_39123 );
and ( w_39122 ,  , w_39123 );
buf ( w_39121 , \14348_b1 );
not ( w_39121 , w_39124 );
not (  , w_39125 );
and ( w_39124 , w_39125 , \14348_b0 );
or ( \14635_b1 , \14625_b1 , w_39126 );
or ( \14635_b0 , \14625_b0 , \14634_b0 );
not ( \14634_b0 , w_39127 );
and ( w_39127 , w_39126 , \14634_b1 );
or ( \14636_b1 , \14298_b1 , \14355_b1 );
not ( \14355_b1 , w_39128 );
and ( \14636_b0 , \14298_b0 , w_39129 );
and ( w_39128 , w_39129 , \14355_b0 );
or ( \14637_b1 , \14636_b1 , w_39131 );
not ( w_39131 , w_39132 );
and ( \14637_b0 , \14636_b0 , w_39133 );
and ( w_39132 ,  , w_39133 );
buf ( w_39131 , \14363_b1 );
not ( w_39131 , w_39134 );
not (  , w_39135 );
and ( w_39134 , w_39135 , \14363_b0 );
or ( \14638_b1 , \14635_b1 , w_39137 );
not ( w_39137 , w_39138 );
and ( \14638_b0 , \14635_b0 , w_39139 );
and ( w_39138 ,  , w_39139 );
buf ( w_39137 , \14637_b1 );
not ( w_39137 , w_39140 );
not (  , w_39141 );
and ( w_39140 , w_39141 , \14637_b0 );
or ( \14639_b1 , \14632_b1 , w_39143 );
not ( w_39143 , w_39144 );
and ( \14639_b0 , \14632_b0 , w_39145 );
and ( w_39144 ,  , w_39145 );
buf ( w_39143 , \14638_b1 );
not ( w_39143 , w_39146 );
not (  , w_39147 );
and ( w_39146 , w_39147 , \14638_b0 );
buf ( \14640_b1 , \14639_b1 );
not ( \14640_b1 , w_39148 );
not ( \14640_b0 , w_39149 );
and ( w_39148 , w_39149 , \14639_b0 );
or ( \14641_b1 , \14623_b1 , w_39150 );
xor ( \14641_b0 , \14623_b0 , w_39152 );
not ( w_39152 , w_39153 );
and ( w_39153 , w_39150 , w_39151 );
buf ( w_39150 , \14640_b1 );
not ( w_39150 , w_39154 );
not ( w_39151 , w_39155 );
and ( w_39154 , w_39155 , \14640_b0 );
buf ( \14642_b1 , \14641_b1 );
buf ( \14642_b0 , \14641_b0 );
buf ( \14643_b1 , \14642_b1 );
buf ( \14643_b0 , \14642_b0 );
buf ( \14644_b1 , \11128_b1 );
not ( \14644_b1 , w_39156 );
not ( \14644_b0 , w_39157 );
and ( w_39156 , w_39157 , \11128_b0 );
or ( \14645_b1 , \13974_b1 , w_39159 );
not ( w_39159 , w_39160 );
and ( \14645_b0 , \13974_b0 , w_39161 );
and ( w_39160 ,  , w_39161 );
buf ( w_39159 , \14644_b1 );
not ( w_39159 , w_39162 );
not (  , w_39163 );
and ( w_39162 , w_39163 , \14644_b0 );
or ( \14646_b1 , \14388_b1 , w_39165 );
not ( w_39165 , w_39166 );
and ( \14646_b0 , \14388_b0 , w_39167 );
and ( w_39166 ,  , w_39167 );
buf ( w_39165 , \14380_b1 );
not ( w_39165 , w_39168 );
not (  , w_39169 );
and ( w_39168 , w_39169 , \14380_b0 );
or ( \14647_b1 , \14381_b1 , w_39171 );
not ( w_39171 , w_39172 );
and ( \14647_b0 , \14381_b0 , w_39173 );
and ( w_39172 ,  , w_39173 );
buf ( w_39171 , \14383_b1 );
not ( w_39171 , w_39174 );
not (  , w_39175 );
and ( w_39174 , w_39175 , \14383_b0 );
or ( \14648_b1 , \14646_b1 , w_39177 );
not ( w_39177 , w_39178 );
and ( \14648_b0 , \14646_b0 , w_39179 );
and ( w_39178 ,  , w_39179 );
buf ( w_39177 , \14647_b1 );
not ( w_39177 , w_39180 );
not (  , w_39181 );
and ( w_39180 , w_39181 , \14647_b0 );
or ( \14649_b1 , \14390_b1 , w_39183 );
not ( w_39183 , w_39184 );
and ( \14649_b0 , \14390_b0 , w_39185 );
and ( w_39184 ,  , w_39185 );
buf ( w_39183 , \14387_b1 );
not ( w_39183 , w_39186 );
not (  , w_39187 );
and ( w_39186 , w_39187 , \14387_b0 );
or ( \14650_b1 , \14649_b1 , w_39188 );
or ( \14650_b0 , \14649_b0 , \13830_b0 );
not ( \13830_b0 , w_39189 );
and ( w_39189 , w_39188 , \13830_b1 );
or ( \14651_b1 , \14387_b1 , \14393_b1 );
not ( \14393_b1 , w_39190 );
and ( \14651_b0 , \14387_b0 , w_39191 );
and ( w_39190 , w_39191 , \14393_b0 );
or ( \14652_b1 , \14651_b1 , w_39193 );
not ( w_39193 , w_39194 );
and ( \14652_b0 , \14651_b0 , w_39195 );
and ( w_39194 ,  , w_39195 );
buf ( w_39193 , \14397_b1 );
not ( w_39193 , w_39196 );
not (  , w_39197 );
and ( w_39196 , w_39197 , \14397_b0 );
or ( \14653_b1 , \14650_b1 , w_39199 );
not ( w_39199 , w_39200 );
and ( \14653_b0 , \14650_b0 , w_39201 );
and ( w_39200 ,  , w_39201 );
buf ( w_39199 , \14652_b1 );
not ( w_39199 , w_39202 );
not (  , w_39203 );
and ( w_39202 , w_39203 , \14652_b0 );
or ( \14654_b1 , \14648_b1 , \14653_b1 );
not ( \14653_b1 , w_39204 );
and ( \14654_b0 , \14648_b0 , w_39205 );
and ( w_39204 , w_39205 , \14653_b0 );
or ( \14655_b1 , \14380_b1 , \14400_b1 );
not ( \14400_b1 , w_39206 );
and ( \14655_b0 , \14380_b0 , w_39207 );
and ( w_39206 , w_39207 , \14400_b0 );
or ( \14656_b1 , \14655_b1 , w_39209 );
not ( w_39209 , w_39210 );
and ( \14656_b0 , \14655_b0 , w_39211 );
and ( w_39210 ,  , w_39211 );
buf ( w_39209 , \14405_b1 );
not ( w_39209 , w_39212 );
not (  , w_39213 );
and ( w_39212 , w_39213 , \14405_b0 );
or ( \14657_b1 , \14647_b1 , w_39214 );
or ( \14657_b0 , \14647_b0 , \14656_b0 );
not ( \14656_b0 , w_39215 );
and ( w_39215 , w_39214 , \14656_b1 );
or ( \14658_b1 , \14383_b1 , \14408_b1 );
not ( \14408_b1 , w_39216 );
and ( \14658_b0 , \14383_b0 , w_39217 );
and ( w_39216 , w_39217 , \14408_b0 );
or ( \14659_b1 , \14658_b1 , w_39219 );
not ( w_39219 , w_39220 );
and ( \14659_b0 , \14658_b0 , w_39221 );
and ( w_39220 ,  , w_39221 );
buf ( w_39219 , \14412_b1 );
not ( w_39219 , w_39222 );
not (  , w_39223 );
and ( w_39222 , w_39223 , \14412_b0 );
or ( \14660_b1 , \14657_b1 , w_39225 );
not ( w_39225 , w_39226 );
and ( \14660_b0 , \14657_b0 , w_39227 );
and ( w_39226 ,  , w_39227 );
buf ( w_39225 , \14659_b1 );
not ( w_39225 , w_39228 );
not (  , w_39229 );
and ( w_39228 , w_39229 , \14659_b0 );
or ( \14661_b1 , \14654_b1 , w_39231 );
not ( w_39231 , w_39232 );
and ( \14661_b0 , \14654_b0 , w_39233 );
and ( w_39232 ,  , w_39233 );
buf ( w_39231 , \14660_b1 );
not ( w_39231 , w_39234 );
not (  , w_39235 );
and ( w_39234 , w_39235 , \14660_b0 );
buf ( \14662_b1 , \14661_b1 );
not ( \14662_b1 , w_39236 );
not ( \14662_b0 , w_39237 );
and ( w_39236 , w_39237 , \14661_b0 );
or ( \14663_b1 , \14645_b1 , w_39238 );
xor ( \14663_b0 , \14645_b0 , w_39240 );
not ( w_39240 , w_39241 );
and ( w_39241 , w_39238 , w_39239 );
buf ( w_39238 , \14662_b1 );
not ( w_39238 , w_39242 );
not ( w_39239 , w_39243 );
and ( w_39242 , w_39243 , \14662_b0 );
buf ( \14664_b1 , \14663_b1 );
buf ( \14664_b0 , \14663_b0 );
buf ( \14665_b1 , \14664_b1 );
buf ( \14665_b0 , \14664_b0 );
buf ( \14666_b1 , \10963_b1 );
not ( \14666_b1 , w_39244 );
not ( \14666_b0 , w_39245 );
and ( w_39244 , w_39245 , \10963_b0 );
or ( \14667_b1 , \13970_b1 , w_39247 );
not ( w_39247 , w_39248 );
and ( \14667_b0 , \13970_b0 , w_39249 );
and ( w_39248 ,  , w_39249 );
buf ( w_39247 , \14666_b1 );
not ( w_39247 , w_39250 );
not (  , w_39251 );
and ( w_39250 , w_39251 , \14666_b0 );
or ( \14668_b1 , \14433_b1 , w_39253 );
not ( w_39253 , w_39254 );
and ( \14668_b0 , \14433_b0 , w_39255 );
and ( w_39254 ,  , w_39255 );
buf ( w_39253 , \14425_b1 );
not ( w_39253 , w_39256 );
not (  , w_39257 );
and ( w_39256 , w_39257 , \14425_b0 );
or ( \14669_b1 , \14426_b1 , w_39259 );
not ( w_39259 , w_39260 );
and ( \14669_b0 , \14426_b0 , w_39261 );
and ( w_39260 ,  , w_39261 );
buf ( w_39259 , \14428_b1 );
not ( w_39259 , w_39262 );
not (  , w_39263 );
and ( w_39262 , w_39263 , \14428_b0 );
or ( \14670_b1 , \14668_b1 , w_39265 );
not ( w_39265 , w_39266 );
and ( \14670_b0 , \14668_b0 , w_39267 );
and ( w_39266 ,  , w_39267 );
buf ( w_39265 , \14669_b1 );
not ( w_39265 , w_39268 );
not (  , w_39269 );
and ( w_39268 , w_39269 , \14669_b0 );
or ( \14671_b1 , \14435_b1 , w_39271 );
not ( w_39271 , w_39272 );
and ( \14671_b0 , \14435_b0 , w_39273 );
and ( w_39272 ,  , w_39273 );
buf ( w_39271 , \14432_b1 );
not ( w_39271 , w_39274 );
not (  , w_39275 );
and ( w_39274 , w_39275 , \14432_b0 );
or ( \14672_b1 , \14671_b1 , w_39276 );
or ( \14672_b0 , \14671_b0 , \13826_b0 );
not ( \13826_b0 , w_39277 );
and ( w_39277 , w_39276 , \13826_b1 );
or ( \14673_b1 , \14432_b1 , \14438_b1 );
not ( \14438_b1 , w_39278 );
and ( \14673_b0 , \14432_b0 , w_39279 );
and ( w_39278 , w_39279 , \14438_b0 );
or ( \14674_b1 , \14673_b1 , w_39281 );
not ( w_39281 , w_39282 );
and ( \14674_b0 , \14673_b0 , w_39283 );
and ( w_39282 ,  , w_39283 );
buf ( w_39281 , \14442_b1 );
not ( w_39281 , w_39284 );
not (  , w_39285 );
and ( w_39284 , w_39285 , \14442_b0 );
or ( \14675_b1 , \14672_b1 , w_39287 );
not ( w_39287 , w_39288 );
and ( \14675_b0 , \14672_b0 , w_39289 );
and ( w_39288 ,  , w_39289 );
buf ( w_39287 , \14674_b1 );
not ( w_39287 , w_39290 );
not (  , w_39291 );
and ( w_39290 , w_39291 , \14674_b0 );
or ( \14676_b1 , \14670_b1 , \14675_b1 );
not ( \14675_b1 , w_39292 );
and ( \14676_b0 , \14670_b0 , w_39293 );
and ( w_39292 , w_39293 , \14675_b0 );
or ( \14677_b1 , \14425_b1 , \14445_b1 );
not ( \14445_b1 , w_39294 );
and ( \14677_b0 , \14425_b0 , w_39295 );
and ( w_39294 , w_39295 , \14445_b0 );
or ( \14678_b1 , \14677_b1 , w_39297 );
not ( w_39297 , w_39298 );
and ( \14678_b0 , \14677_b0 , w_39299 );
and ( w_39298 ,  , w_39299 );
buf ( w_39297 , \14450_b1 );
not ( w_39297 , w_39300 );
not (  , w_39301 );
and ( w_39300 , w_39301 , \14450_b0 );
or ( \14679_b1 , \14669_b1 , w_39302 );
or ( \14679_b0 , \14669_b0 , \14678_b0 );
not ( \14678_b0 , w_39303 );
and ( w_39303 , w_39302 , \14678_b1 );
or ( \14680_b1 , \14428_b1 , \14453_b1 );
not ( \14453_b1 , w_39304 );
and ( \14680_b0 , \14428_b0 , w_39305 );
and ( w_39304 , w_39305 , \14453_b0 );
or ( \14681_b1 , \14680_b1 , w_39307 );
not ( w_39307 , w_39308 );
and ( \14681_b0 , \14680_b0 , w_39309 );
and ( w_39308 ,  , w_39309 );
buf ( w_39307 , \14457_b1 );
not ( w_39307 , w_39310 );
not (  , w_39311 );
and ( w_39310 , w_39311 , \14457_b0 );
or ( \14682_b1 , \14679_b1 , w_39313 );
not ( w_39313 , w_39314 );
and ( \14682_b0 , \14679_b0 , w_39315 );
and ( w_39314 ,  , w_39315 );
buf ( w_39313 , \14681_b1 );
not ( w_39313 , w_39316 );
not (  , w_39317 );
and ( w_39316 , w_39317 , \14681_b0 );
or ( \14683_b1 , \14676_b1 , w_39319 );
not ( w_39319 , w_39320 );
and ( \14683_b0 , \14676_b0 , w_39321 );
and ( w_39320 ,  , w_39321 );
buf ( w_39319 , \14682_b1 );
not ( w_39319 , w_39322 );
not (  , w_39323 );
and ( w_39322 , w_39323 , \14682_b0 );
buf ( \14684_b1 , \14683_b1 );
not ( \14684_b1 , w_39324 );
not ( \14684_b0 , w_39325 );
and ( w_39324 , w_39325 , \14683_b0 );
or ( \14685_b1 , \14667_b1 , w_39326 );
xor ( \14685_b0 , \14667_b0 , w_39328 );
not ( w_39328 , w_39329 );
and ( w_39329 , w_39326 , w_39327 );
buf ( w_39326 , \14684_b1 );
not ( w_39326 , w_39330 );
not ( w_39327 , w_39331 );
and ( w_39330 , w_39331 , \14684_b0 );
buf ( \14686_b1 , \14685_b1 );
buf ( \14686_b0 , \14685_b0 );
buf ( \14687_b1 , \14686_b1 );
buf ( \14687_b0 , \14686_b0 );
buf ( \14688_b1 , \10802_b1 );
not ( \14688_b1 , w_39332 );
not ( \14688_b0 , w_39333 );
and ( w_39332 , w_39333 , \10802_b0 );
or ( \14689_b1 , \13968_b1 , w_39335 );
not ( w_39335 , w_39336 );
and ( \14689_b0 , \13968_b0 , w_39337 );
and ( w_39336 ,  , w_39337 );
buf ( w_39335 , \14688_b1 );
not ( w_39335 , w_39338 );
not (  , w_39339 );
and ( w_39338 , w_39339 , \14688_b0 );
or ( \14690_b1 , \14478_b1 , w_39341 );
not ( w_39341 , w_39342 );
and ( \14690_b0 , \14478_b0 , w_39343 );
and ( w_39342 ,  , w_39343 );
buf ( w_39341 , \14470_b1 );
not ( w_39341 , w_39344 );
not (  , w_39345 );
and ( w_39344 , w_39345 , \14470_b0 );
or ( \14691_b1 , \14471_b1 , w_39347 );
not ( w_39347 , w_39348 );
and ( \14691_b0 , \14471_b0 , w_39349 );
and ( w_39348 ,  , w_39349 );
buf ( w_39347 , \14473_b1 );
not ( w_39347 , w_39350 );
not (  , w_39351 );
and ( w_39350 , w_39351 , \14473_b0 );
or ( \14692_b1 , \14690_b1 , w_39353 );
not ( w_39353 , w_39354 );
and ( \14692_b0 , \14690_b0 , w_39355 );
and ( w_39354 ,  , w_39355 );
buf ( w_39353 , \14691_b1 );
not ( w_39353 , w_39356 );
not (  , w_39357 );
and ( w_39356 , w_39357 , \14691_b0 );
or ( \14693_b1 , \14477_b1 , \14481_b1 );
not ( \14481_b1 , w_39358 );
and ( \14693_b0 , \14477_b0 , w_39359 );
and ( w_39358 , w_39359 , \14481_b0 );
or ( \14694_b1 , \14693_b1 , w_39361 );
not ( w_39361 , w_39362 );
and ( \14694_b0 , \14693_b0 , w_39363 );
and ( w_39362 ,  , w_39363 );
buf ( w_39361 , \14485_b1 );
not ( w_39361 , w_39364 );
not (  , w_39365 );
and ( w_39364 , w_39365 , \14485_b0 );
buf ( \14695_b1 , \14694_b1 );
not ( \14695_b1 , w_39366 );
not ( \14695_b0 , w_39367 );
and ( w_39366 , w_39367 , \14694_b0 );
or ( \14696_b1 , \14692_b1 , \14695_b1 );
not ( \14695_b1 , w_39368 );
and ( \14696_b0 , \14692_b0 , w_39369 );
and ( w_39368 , w_39369 , \14695_b0 );
or ( \14697_b1 , \14470_b1 , \14488_b1 );
not ( \14488_b1 , w_39370 );
and ( \14697_b0 , \14470_b0 , w_39371 );
and ( w_39370 , w_39371 , \14488_b0 );
or ( \14698_b1 , \14697_b1 , w_39373 );
not ( w_39373 , w_39374 );
and ( \14698_b0 , \14697_b0 , w_39375 );
and ( w_39374 ,  , w_39375 );
buf ( w_39373 , \14493_b1 );
not ( w_39373 , w_39376 );
not (  , w_39377 );
and ( w_39376 , w_39377 , \14493_b0 );
or ( \14699_b1 , \14691_b1 , w_39378 );
or ( \14699_b0 , \14691_b0 , \14698_b0 );
not ( \14698_b0 , w_39379 );
and ( w_39379 , w_39378 , \14698_b1 );
or ( \14700_b1 , \14473_b1 , \14496_b1 );
not ( \14496_b1 , w_39380 );
and ( \14700_b0 , \14473_b0 , w_39381 );
and ( w_39380 , w_39381 , \14496_b0 );
or ( \14701_b1 , \14700_b1 , w_39383 );
not ( w_39383 , w_39384 );
and ( \14701_b0 , \14700_b0 , w_39385 );
and ( w_39384 ,  , w_39385 );
buf ( w_39383 , \14500_b1 );
not ( w_39383 , w_39386 );
not (  , w_39387 );
and ( w_39386 , w_39387 , \14500_b0 );
or ( \14702_b1 , \14699_b1 , w_39389 );
not ( w_39389 , w_39390 );
and ( \14702_b0 , \14699_b0 , w_39391 );
and ( w_39390 ,  , w_39391 );
buf ( w_39389 , \14701_b1 );
not ( w_39389 , w_39392 );
not (  , w_39393 );
and ( w_39392 , w_39393 , \14701_b0 );
or ( \14703_b1 , \14696_b1 , w_39395 );
not ( w_39395 , w_39396 );
and ( \14703_b0 , \14696_b0 , w_39397 );
and ( w_39396 ,  , w_39397 );
buf ( w_39395 , \14702_b1 );
not ( w_39395 , w_39398 );
not (  , w_39399 );
and ( w_39398 , w_39399 , \14702_b0 );
buf ( \14704_b1 , \14703_b1 );
not ( \14704_b1 , w_39400 );
not ( \14704_b0 , w_39401 );
and ( w_39400 , w_39401 , \14703_b0 );
or ( \14705_b1 , \14689_b1 , w_39402 );
xor ( \14705_b0 , \14689_b0 , w_39404 );
not ( w_39404 , w_39405 );
and ( w_39405 , w_39402 , w_39403 );
buf ( w_39402 , \14704_b1 );
not ( w_39402 , w_39406 );
not ( w_39403 , w_39407 );
and ( w_39406 , w_39407 , \14704_b0 );
buf ( \14706_b1 , \14705_b1 );
buf ( \14706_b0 , \14705_b0 );
buf ( \14707_b1 , \14706_b1 );
buf ( \14707_b0 , \14706_b0 );
buf ( \14708_b1 , \10638_b1 );
not ( \14708_b1 , w_39408 );
not ( \14708_b0 , w_39409 );
and ( w_39408 , w_39409 , \10638_b0 );
or ( \14709_b1 , \13965_b1 , w_39411 );
not ( w_39411 , w_39412 );
and ( \14709_b0 , \13965_b0 , w_39413 );
and ( w_39412 ,  , w_39413 );
buf ( w_39411 , \14708_b1 );
not ( w_39411 , w_39414 );
not (  , w_39415 );
and ( w_39414 , w_39415 , \14708_b0 );
or ( \14710_b1 , \14521_b1 , w_39417 );
not ( w_39417 , w_39418 );
and ( \14710_b0 , \14521_b0 , w_39419 );
and ( w_39418 ,  , w_39419 );
buf ( w_39417 , \14513_b1 );
not ( w_39417 , w_39420 );
not (  , w_39421 );
and ( w_39420 , w_39421 , \14513_b0 );
or ( \14711_b1 , \14514_b1 , w_39423 );
not ( w_39423 , w_39424 );
and ( \14711_b0 , \14514_b0 , w_39425 );
and ( w_39424 ,  , w_39425 );
buf ( w_39423 , \14516_b1 );
not ( w_39423 , w_39426 );
not (  , w_39427 );
and ( w_39426 , w_39427 , \14516_b0 );
or ( \14712_b1 , \14710_b1 , w_39429 );
not ( w_39429 , w_39430 );
and ( \14712_b0 , \14710_b0 , w_39431 );
and ( w_39430 ,  , w_39431 );
buf ( w_39429 , \14711_b1 );
not ( w_39429 , w_39432 );
not (  , w_39433 );
and ( w_39432 , w_39433 , \14711_b0 );
or ( \14713_b1 , \14520_b1 , \14524_b1 );
not ( \14524_b1 , w_39434 );
and ( \14713_b0 , \14520_b0 , w_39435 );
and ( w_39434 , w_39435 , \14524_b0 );
or ( \14714_b1 , \14713_b1 , w_39437 );
not ( w_39437 , w_39438 );
and ( \14714_b0 , \14713_b0 , w_39439 );
and ( w_39438 ,  , w_39439 );
buf ( w_39437 , \14528_b1 );
not ( w_39437 , w_39440 );
not (  , w_39441 );
and ( w_39440 , w_39441 , \14528_b0 );
buf ( \14715_b1 , \14714_b1 );
not ( \14715_b1 , w_39442 );
not ( \14715_b0 , w_39443 );
and ( w_39442 , w_39443 , \14714_b0 );
or ( \14716_b1 , \14712_b1 , \14715_b1 );
not ( \14715_b1 , w_39444 );
and ( \14716_b0 , \14712_b0 , w_39445 );
and ( w_39444 , w_39445 , \14715_b0 );
or ( \14717_b1 , \14513_b1 , \14531_b1 );
not ( \14531_b1 , w_39446 );
and ( \14717_b0 , \14513_b0 , w_39447 );
and ( w_39446 , w_39447 , \14531_b0 );
or ( \14718_b1 , \14717_b1 , w_39449 );
not ( w_39449 , w_39450 );
and ( \14718_b0 , \14717_b0 , w_39451 );
and ( w_39450 ,  , w_39451 );
buf ( w_39449 , \14536_b1 );
not ( w_39449 , w_39452 );
not (  , w_39453 );
and ( w_39452 , w_39453 , \14536_b0 );
or ( \14719_b1 , \14711_b1 , w_39454 );
or ( \14719_b0 , \14711_b0 , \14718_b0 );
not ( \14718_b0 , w_39455 );
and ( w_39455 , w_39454 , \14718_b1 );
or ( \14720_b1 , \14516_b1 , \14539_b1 );
not ( \14539_b1 , w_39456 );
and ( \14720_b0 , \14516_b0 , w_39457 );
and ( w_39456 , w_39457 , \14539_b0 );
or ( \14721_b1 , \14720_b1 , w_39459 );
not ( w_39459 , w_39460 );
and ( \14721_b0 , \14720_b0 , w_39461 );
and ( w_39460 ,  , w_39461 );
buf ( w_39459 , \14543_b1 );
not ( w_39459 , w_39462 );
not (  , w_39463 );
and ( w_39462 , w_39463 , \14543_b0 );
or ( \14722_b1 , \14719_b1 , w_39465 );
not ( w_39465 , w_39466 );
and ( \14722_b0 , \14719_b0 , w_39467 );
and ( w_39466 ,  , w_39467 );
buf ( w_39465 , \14721_b1 );
not ( w_39465 , w_39468 );
not (  , w_39469 );
and ( w_39468 , w_39469 , \14721_b0 );
or ( \14723_b1 , \14716_b1 , w_39471 );
not ( w_39471 , w_39472 );
and ( \14723_b0 , \14716_b0 , w_39473 );
and ( w_39472 ,  , w_39473 );
buf ( w_39471 , \14722_b1 );
not ( w_39471 , w_39474 );
not (  , w_39475 );
and ( w_39474 , w_39475 , \14722_b0 );
buf ( \14724_b1 , \14723_b1 );
not ( \14724_b1 , w_39476 );
not ( \14724_b0 , w_39477 );
and ( w_39476 , w_39477 , \14723_b0 );
or ( \14725_b1 , \14709_b1 , w_39478 );
xor ( \14725_b0 , \14709_b0 , w_39480 );
not ( w_39480 , w_39481 );
and ( w_39481 , w_39478 , w_39479 );
buf ( w_39478 , \14724_b1 );
not ( w_39478 , w_39482 );
not ( w_39479 , w_39483 );
and ( w_39482 , w_39483 , \14724_b0 );
buf ( \14726_b1 , \14725_b1 );
buf ( \14726_b0 , \14725_b0 );
buf ( \14727_b1 , \14726_b1 );
buf ( \14727_b0 , \14726_b0 );
buf ( \14728_b1 , \10477_b1 );
not ( \14728_b1 , w_39484 );
not ( \14728_b0 , w_39485 );
and ( w_39484 , w_39485 , \10477_b0 );
or ( \14729_b1 , \13963_b1 , w_39487 );
not ( w_39487 , w_39488 );
and ( \14729_b0 , \13963_b0 , w_39489 );
and ( w_39488 ,  , w_39489 );
buf ( w_39487 , \14728_b1 );
not ( w_39487 , w_39490 );
not (  , w_39491 );
and ( w_39490 , w_39491 , \14728_b0 );
or ( \14730_b1 , \13514_b1 , w_39493 );
not ( w_39493 , w_39494 );
and ( \14730_b0 , \13514_b0 , w_39495 );
and ( w_39494 ,  , w_39495 );
buf ( w_39493 , \10314_b1 );
not ( w_39493 , w_39496 );
not (  , w_39497 );
and ( w_39496 , w_39497 , \10314_b0 );
buf ( \14731_b1 , \13866_b1 );
not ( \14731_b1 , w_39498 );
not ( \14731_b0 , w_39499 );
and ( w_39498 , w_39499 , \13866_b0 );
or ( \14732_b1 , \14730_b1 , \14731_b1 );
not ( \14731_b1 , w_39500 );
and ( \14732_b0 , \14730_b0 , w_39501 );
and ( w_39500 , w_39501 , \14731_b0 );
or ( \14733_b1 , \10314_b1 , w_39502 );
or ( \14733_b0 , \10314_b0 , \13913_b0 );
not ( \13913_b0 , w_39503 );
and ( w_39503 , w_39502 , \13913_b1 );
or ( \14734_b1 , \14733_b1 , w_39505 );
not ( w_39505 , w_39506 );
and ( \14734_b0 , \14733_b0 , w_39507 );
and ( w_39506 ,  , w_39507 );
buf ( w_39505 , \13961_b1 );
not ( w_39505 , w_39508 );
not (  , w_39509 );
and ( w_39508 , w_39509 , \13961_b0 );
or ( \14735_b1 , \14732_b1 , w_39511 );
not ( w_39511 , w_39512 );
and ( \14735_b0 , \14732_b0 , w_39513 );
and ( w_39512 ,  , w_39513 );
buf ( w_39511 , \14734_b1 );
not ( w_39511 , w_39514 );
not (  , w_39515 );
and ( w_39514 , w_39515 , \14734_b0 );
buf ( \14736_b1 , \14735_b1 );
not ( \14736_b1 , w_39516 );
not ( \14736_b0 , w_39517 );
and ( w_39516 , w_39517 , \14735_b0 );
or ( \14737_b1 , \14729_b1 , w_39518 );
xor ( \14737_b0 , \14729_b0 , w_39520 );
not ( w_39520 , w_39521 );
and ( w_39521 , w_39518 , w_39519 );
buf ( w_39518 , \14736_b1 );
not ( w_39518 , w_39522 );
not ( w_39519 , w_39523 );
and ( w_39522 , w_39523 , \14736_b0 );
buf ( \14738_b1 , \14737_b1 );
buf ( \14738_b0 , \14737_b0 );
buf ( \14739_b1 , \14738_b1 );
buf ( \14739_b0 , \14738_b0 );
buf ( \14740_b1 , \10310_b1 );
not ( \14740_b1 , w_39524 );
not ( \14740_b0 , w_39525 );
and ( w_39524 , w_39525 , \10310_b0 );
or ( \14741_b1 , \13957_b1 , w_39527 );
not ( w_39527 , w_39528 );
and ( \14741_b0 , \13957_b0 , w_39529 );
and ( w_39528 ,  , w_39529 );
buf ( w_39527 , \14740_b1 );
not ( w_39527 , w_39530 );
not (  , w_39531 );
and ( w_39530 , w_39531 , \14740_b0 );
or ( \14742_b1 , \14062_b1 , w_39533 );
not ( w_39533 , w_39534 );
and ( \14742_b0 , \14062_b0 , w_39535 );
and ( w_39534 ,  , w_39535 );
buf ( w_39533 , \14031_b1 );
not ( w_39533 , w_39536 );
not (  , w_39537 );
and ( w_39536 , w_39537 , \14031_b0 );
buf ( \14743_b1 , \14096_b1 );
not ( \14743_b1 , w_39538 );
not ( \14743_b0 , w_39539 );
and ( w_39538 , w_39539 , \14096_b0 );
or ( \14744_b1 , \14742_b1 , \14743_b1 );
not ( \14743_b1 , w_39540 );
and ( \14744_b0 , \14742_b0 , w_39541 );
and ( w_39540 , w_39541 , \14743_b0 );
or ( \14745_b1 , \14031_b1 , w_39542 );
or ( \14745_b0 , \14031_b0 , \14127_b0 );
not ( \14127_b0 , w_39543 );
and ( w_39543 , w_39542 , \14127_b1 );
or ( \14746_b1 , \14745_b1 , w_39545 );
not ( w_39545 , w_39546 );
and ( \14746_b0 , \14745_b0 , w_39547 );
and ( w_39546 ,  , w_39547 );
buf ( w_39545 , \14159_b1 );
not ( w_39545 , w_39548 );
not (  , w_39549 );
and ( w_39548 , w_39549 , \14159_b0 );
or ( \14747_b1 , \14744_b1 , w_39551 );
not ( w_39551 , w_39552 );
and ( \14747_b0 , \14744_b0 , w_39553 );
and ( w_39552 ,  , w_39553 );
buf ( w_39551 , \14746_b1 );
not ( w_39551 , w_39554 );
not (  , w_39555 );
and ( w_39554 , w_39555 , \14746_b0 );
buf ( \14748_b1 , \14747_b1 );
not ( \14748_b1 , w_39556 );
not ( \14748_b0 , w_39557 );
and ( w_39556 , w_39557 , \14747_b0 );
or ( \14749_b1 , \14741_b1 , w_39558 );
xor ( \14749_b0 , \14741_b0 , w_39560 );
not ( w_39560 , w_39561 );
and ( w_39561 , w_39558 , w_39559 );
buf ( w_39558 , \14748_b1 );
not ( w_39558 , w_39562 );
not ( w_39559 , w_39563 );
and ( w_39562 , w_39563 , \14748_b0 );
buf ( \14750_b1 , \14749_b1 );
buf ( \14750_b0 , \14749_b0 );
buf ( \14751_b1 , \14750_b1 );
buf ( \14751_b0 , \14750_b0 );
buf ( \14752_b1 , \10149_b1 );
not ( \14752_b1 , w_39564 );
not ( \14752_b0 , w_39565 );
and ( w_39564 , w_39565 , \10149_b0 );
or ( \14753_b1 , \13955_b1 , w_39567 );
not ( w_39567 , w_39568 );
and ( \14753_b0 , \13955_b0 , w_39569 );
and ( w_39568 ,  , w_39569 );
buf ( w_39567 , \14752_b1 );
not ( w_39567 , w_39570 );
not (  , w_39571 );
and ( w_39570 , w_39571 , \14752_b0 );
or ( \14754_b1 , \14220_b1 , w_39573 );
not ( w_39573 , w_39574 );
and ( \14754_b0 , \14220_b0 , w_39575 );
and ( w_39574 ,  , w_39575 );
buf ( w_39573 , \14205_b1 );
not ( w_39573 , w_39576 );
not (  , w_39577 );
and ( w_39576 , w_39577 , \14205_b0 );
buf ( \14755_b1 , \14234_b1 );
not ( \14755_b1 , w_39578 );
not ( \14755_b0 , w_39579 );
and ( w_39578 , w_39579 , \14234_b0 );
or ( \14756_b1 , \14754_b1 , \14755_b1 );
not ( \14755_b1 , w_39580 );
and ( \14756_b0 , \14754_b0 , w_39581 );
and ( w_39580 , w_39581 , \14755_b0 );
or ( \14757_b1 , \14205_b1 , w_39582 );
or ( \14757_b0 , \14205_b0 , \14249_b0 );
not ( \14249_b0 , w_39583 );
and ( w_39583 , w_39582 , \14249_b1 );
or ( \14758_b1 , \14757_b1 , w_39585 );
not ( w_39585 , w_39586 );
and ( \14758_b0 , \14757_b0 , w_39587 );
and ( w_39586 ,  , w_39587 );
buf ( w_39585 , \14265_b1 );
not ( w_39585 , w_39588 );
not (  , w_39589 );
and ( w_39588 , w_39589 , \14265_b0 );
or ( \14759_b1 , \14756_b1 , w_39591 );
not ( w_39591 , w_39592 );
and ( \14759_b0 , \14756_b0 , w_39593 );
and ( w_39592 ,  , w_39593 );
buf ( w_39591 , \14758_b1 );
not ( w_39591 , w_39594 );
not (  , w_39595 );
and ( w_39594 , w_39595 , \14758_b0 );
buf ( \14760_b1 , \14759_b1 );
not ( \14760_b1 , w_39596 );
not ( \14760_b0 , w_39597 );
and ( w_39596 , w_39597 , \14759_b0 );
or ( \14761_b1 , \14753_b1 , w_39598 );
xor ( \14761_b0 , \14753_b0 , w_39600 );
not ( w_39600 , w_39601 );
and ( w_39601 , w_39598 , w_39599 );
buf ( w_39598 , \14760_b1 );
not ( w_39598 , w_39602 );
not ( w_39599 , w_39603 );
and ( w_39602 , w_39603 , \14760_b0 );
buf ( \14762_b1 , \14761_b1 );
buf ( \14762_b0 , \14761_b0 );
buf ( \14763_b1 , \14762_b1 );
buf ( \14763_b0 , \14762_b0 );
buf ( \14764_b1 , \9985_b1 );
not ( \14764_b1 , w_39604 );
not ( \14764_b0 , w_39605 );
and ( w_39604 , w_39605 , \9985_b0 );
or ( \14765_b1 , \13952_b1 , w_39607 );
not ( w_39607 , w_39608 );
and ( \14765_b0 , \13952_b0 , w_39609 );
and ( w_39608 ,  , w_39609 );
buf ( w_39607 , \14764_b1 );
not ( w_39607 , w_39610 );
not (  , w_39611 );
and ( w_39610 , w_39611 , \14764_b0 );
or ( \14766_b1 , \14310_b1 , w_39613 );
not ( w_39613 , w_39614 );
and ( \14766_b0 , \14310_b0 , w_39615 );
and ( w_39614 ,  , w_39615 );
buf ( w_39613 , \14295_b1 );
not ( w_39613 , w_39616 );
not (  , w_39617 );
and ( w_39616 , w_39617 , \14295_b0 );
buf ( \14767_b1 , \14325_b1 );
not ( \14767_b1 , w_39618 );
not ( \14767_b0 , w_39619 );
and ( w_39618 , w_39619 , \14325_b0 );
or ( \14768_b1 , \14766_b1 , \14767_b1 );
not ( \14767_b1 , w_39620 );
and ( \14768_b0 , \14766_b0 , w_39621 );
and ( w_39620 , w_39621 , \14767_b0 );
or ( \14769_b1 , \14295_b1 , w_39622 );
or ( \14769_b0 , \14295_b0 , \14340_b0 );
not ( \14340_b0 , w_39623 );
and ( w_39623 , w_39622 , \14340_b1 );
or ( \14770_b1 , \14769_b1 , w_39625 );
not ( w_39625 , w_39626 );
and ( \14770_b0 , \14769_b0 , w_39627 );
and ( w_39626 ,  , w_39627 );
buf ( w_39625 , \14356_b1 );
not ( w_39625 , w_39628 );
not (  , w_39629 );
and ( w_39628 , w_39629 , \14356_b0 );
or ( \14771_b1 , \14768_b1 , w_39631 );
not ( w_39631 , w_39632 );
and ( \14771_b0 , \14768_b0 , w_39633 );
and ( w_39632 ,  , w_39633 );
buf ( w_39631 , \14770_b1 );
not ( w_39631 , w_39634 );
not (  , w_39635 );
and ( w_39634 , w_39635 , \14770_b0 );
buf ( \14772_b1 , \14771_b1 );
not ( \14772_b1 , w_39636 );
not ( \14772_b0 , w_39637 );
and ( w_39636 , w_39637 , \14771_b0 );
or ( \14773_b1 , \14765_b1 , w_39638 );
xor ( \14773_b0 , \14765_b0 , w_39640 );
not ( w_39640 , w_39641 );
and ( w_39641 , w_39638 , w_39639 );
buf ( w_39638 , \14772_b1 );
not ( w_39638 , w_39642 );
not ( w_39639 , w_39643 );
and ( w_39642 , w_39643 , \14772_b0 );
buf ( \14774_b1 , \14773_b1 );
buf ( \14774_b0 , \14773_b0 );
buf ( \14775_b1 , \14774_b1 );
buf ( \14775_b0 , \14774_b0 );
buf ( \14776_b1 , \9824_b1 );
not ( \14776_b1 , w_39644 );
not ( \14776_b0 , w_39645 );
and ( w_39644 , w_39645 , \9824_b0 );
or ( \14777_b1 , \13950_b1 , w_39647 );
not ( w_39647 , w_39648 );
and ( \14777_b0 , \13950_b0 , w_39649 );
and ( w_39648 ,  , w_39649 );
buf ( w_39647 , \14776_b1 );
not ( w_39647 , w_39650 );
not (  , w_39651 );
and ( w_39650 , w_39651 , \14776_b0 );
or ( \14778_b1 , \14389_b1 , w_39653 );
not ( w_39653 , w_39654 );
and ( \14778_b0 , \14389_b0 , w_39655 );
and ( w_39654 ,  , w_39655 );
buf ( w_39653 , \14382_b1 );
not ( w_39653 , w_39656 );
not (  , w_39657 );
and ( w_39656 , w_39657 , \14382_b0 );
buf ( \14779_b1 , \14394_b1 );
not ( \14779_b1 , w_39658 );
not ( \14779_b0 , w_39659 );
and ( w_39658 , w_39659 , \14394_b0 );
or ( \14780_b1 , \14778_b1 , \14779_b1 );
not ( \14779_b1 , w_39660 );
and ( \14780_b0 , \14778_b0 , w_39661 );
and ( w_39660 , w_39661 , \14779_b0 );
or ( \14781_b1 , \14382_b1 , w_39662 );
or ( \14781_b0 , \14382_b0 , \14401_b0 );
not ( \14401_b0 , w_39663 );
and ( w_39663 , w_39662 , \14401_b1 );
or ( \14782_b1 , \14781_b1 , w_39665 );
not ( w_39665 , w_39666 );
and ( \14782_b0 , \14781_b0 , w_39667 );
and ( w_39666 ,  , w_39667 );
buf ( w_39665 , \14409_b1 );
not ( w_39665 , w_39668 );
not (  , w_39669 );
and ( w_39668 , w_39669 , \14409_b0 );
or ( \14783_b1 , \14780_b1 , w_39671 );
not ( w_39671 , w_39672 );
and ( \14783_b0 , \14780_b0 , w_39673 );
and ( w_39672 ,  , w_39673 );
buf ( w_39671 , \14782_b1 );
not ( w_39671 , w_39674 );
not (  , w_39675 );
and ( w_39674 , w_39675 , \14782_b0 );
buf ( \14784_b1 , \14783_b1 );
not ( \14784_b1 , w_39676 );
not ( \14784_b0 , w_39677 );
and ( w_39676 , w_39677 , \14783_b0 );
or ( \14785_b1 , \14777_b1 , w_39678 );
xor ( \14785_b0 , \14777_b0 , w_39680 );
not ( w_39680 , w_39681 );
and ( w_39681 , w_39678 , w_39679 );
buf ( w_39678 , \14784_b1 );
not ( w_39678 , w_39682 );
not ( w_39679 , w_39683 );
and ( w_39682 , w_39683 , \14784_b0 );
buf ( \14786_b1 , \14785_b1 );
buf ( \14786_b0 , \14785_b0 );
buf ( \14787_b1 , \14786_b1 );
buf ( \14787_b0 , \14786_b0 );
buf ( \14788_b1 , \9659_b1 );
not ( \14788_b1 , w_39684 );
not ( \14788_b0 , w_39685 );
and ( w_39684 , w_39685 , \9659_b0 );
or ( \14789_b1 , \13946_b1 , w_39687 );
not ( w_39687 , w_39688 );
and ( \14789_b0 , \13946_b0 , w_39689 );
and ( w_39688 ,  , w_39689 );
buf ( w_39687 , \14788_b1 );
not ( w_39687 , w_39690 );
not (  , w_39691 );
and ( w_39690 , w_39691 , \14788_b0 );
or ( \14790_b1 , \14434_b1 , w_39693 );
not ( w_39693 , w_39694 );
and ( \14790_b0 , \14434_b0 , w_39695 );
and ( w_39694 ,  , w_39695 );
buf ( w_39693 , \14427_b1 );
not ( w_39693 , w_39696 );
not (  , w_39697 );
and ( w_39696 , w_39697 , \14427_b0 );
buf ( \14791_b1 , \14439_b1 );
not ( \14791_b1 , w_39698 );
not ( \14791_b0 , w_39699 );
and ( w_39698 , w_39699 , \14439_b0 );
or ( \14792_b1 , \14790_b1 , \14791_b1 );
not ( \14791_b1 , w_39700 );
and ( \14792_b0 , \14790_b0 , w_39701 );
and ( w_39700 , w_39701 , \14791_b0 );
or ( \14793_b1 , \14427_b1 , w_39702 );
or ( \14793_b0 , \14427_b0 , \14446_b0 );
not ( \14446_b0 , w_39703 );
and ( w_39703 , w_39702 , \14446_b1 );
or ( \14794_b1 , \14793_b1 , w_39705 );
not ( w_39705 , w_39706 );
and ( \14794_b0 , \14793_b0 , w_39707 );
and ( w_39706 ,  , w_39707 );
buf ( w_39705 , \14454_b1 );
not ( w_39705 , w_39708 );
not (  , w_39709 );
and ( w_39708 , w_39709 , \14454_b0 );
or ( \14795_b1 , \14792_b1 , w_39711 );
not ( w_39711 , w_39712 );
and ( \14795_b0 , \14792_b0 , w_39713 );
and ( w_39712 ,  , w_39713 );
buf ( w_39711 , \14794_b1 );
not ( w_39711 , w_39714 );
not (  , w_39715 );
and ( w_39714 , w_39715 , \14794_b0 );
buf ( \14796_b1 , \14795_b1 );
not ( \14796_b1 , w_39716 );
not ( \14796_b0 , w_39717 );
and ( w_39716 , w_39717 , \14795_b0 );
or ( \14797_b1 , \14789_b1 , w_39718 );
xor ( \14797_b0 , \14789_b0 , w_39720 );
not ( w_39720 , w_39721 );
and ( w_39721 , w_39718 , w_39719 );
buf ( w_39718 , \14796_b1 );
not ( w_39718 , w_39722 );
not ( w_39719 , w_39723 );
and ( w_39722 , w_39723 , \14796_b0 );
buf ( \14798_b1 , \14797_b1 );
buf ( \14798_b0 , \14797_b0 );
buf ( \14799_b1 , \14798_b1 );
buf ( \14799_b0 , \14798_b0 );
buf ( \14800_b1 , \9498_b1 );
not ( \14800_b1 , w_39724 );
not ( \14800_b0 , w_39725 );
and ( w_39724 , w_39725 , \9498_b0 );
or ( \14801_b1 , \13944_b1 , w_39727 );
not ( w_39727 , w_39728 );
and ( \14801_b0 , \13944_b0 , w_39729 );
and ( w_39728 ,  , w_39729 );
buf ( w_39727 , \14800_b1 );
not ( w_39727 , w_39730 );
not (  , w_39731 );
and ( w_39730 , w_39731 , \14800_b0 );
or ( \14802_b1 , \14479_b1 , w_39733 );
not ( w_39733 , w_39734 );
and ( \14802_b0 , \14479_b0 , w_39735 );
and ( w_39734 ,  , w_39735 );
buf ( w_39733 , \14472_b1 );
not ( w_39733 , w_39736 );
not (  , w_39737 );
and ( w_39736 , w_39737 , \14472_b0 );
or ( \14803_b1 , \14802_b1 , \14481_b1 );
not ( \14481_b1 , w_39738 );
and ( \14803_b0 , \14802_b0 , w_39739 );
and ( w_39738 , w_39739 , \14481_b0 );
or ( \14804_b1 , \14472_b1 , w_39740 );
or ( \14804_b0 , \14472_b0 , \14489_b0 );
not ( \14489_b0 , w_39741 );
and ( w_39741 , w_39740 , \14489_b1 );
or ( \14805_b1 , \14804_b1 , w_39743 );
not ( w_39743 , w_39744 );
and ( \14805_b0 , \14804_b0 , w_39745 );
and ( w_39744 ,  , w_39745 );
buf ( w_39743 , \14497_b1 );
not ( w_39743 , w_39746 );
not (  , w_39747 );
and ( w_39746 , w_39747 , \14497_b0 );
or ( \14806_b1 , \14803_b1 , w_39749 );
not ( w_39749 , w_39750 );
and ( \14806_b0 , \14803_b0 , w_39751 );
and ( w_39750 ,  , w_39751 );
buf ( w_39749 , \14805_b1 );
not ( w_39749 , w_39752 );
not (  , w_39753 );
and ( w_39752 , w_39753 , \14805_b0 );
buf ( \14807_b1 , \14806_b1 );
not ( \14807_b1 , w_39754 );
not ( \14807_b0 , w_39755 );
and ( w_39754 , w_39755 , \14806_b0 );
or ( \14808_b1 , \14801_b1 , w_39756 );
xor ( \14808_b0 , \14801_b0 , w_39758 );
not ( w_39758 , w_39759 );
and ( w_39759 , w_39756 , w_39757 );
buf ( w_39756 , \14807_b1 );
not ( w_39756 , w_39760 );
not ( w_39757 , w_39761 );
and ( w_39760 , w_39761 , \14807_b0 );
buf ( \14809_b1 , \14808_b1 );
buf ( \14809_b0 , \14808_b0 );
buf ( \14810_b1 , \14809_b1 );
buf ( \14810_b0 , \14809_b0 );
buf ( \14811_b1 , \9334_b1 );
not ( \14811_b1 , w_39762 );
not ( \14811_b0 , w_39763 );
and ( w_39762 , w_39763 , \9334_b0 );
or ( \14812_b1 , \13941_b1 , w_39765 );
not ( w_39765 , w_39766 );
and ( \14812_b0 , \13941_b0 , w_39767 );
and ( w_39766 ,  , w_39767 );
buf ( w_39765 , \14811_b1 );
not ( w_39765 , w_39768 );
not (  , w_39769 );
and ( w_39768 , w_39769 , \14811_b0 );
or ( \14813_b1 , \14522_b1 , w_39771 );
not ( w_39771 , w_39772 );
and ( \14813_b0 , \14522_b0 , w_39773 );
and ( w_39772 ,  , w_39773 );
buf ( w_39771 , \14515_b1 );
not ( w_39771 , w_39774 );
not (  , w_39775 );
and ( w_39774 , w_39775 , \14515_b0 );
or ( \14814_b1 , \14813_b1 , \14524_b1 );
not ( \14524_b1 , w_39776 );
and ( \14814_b0 , \14813_b0 , w_39777 );
and ( w_39776 , w_39777 , \14524_b0 );
or ( \14815_b1 , \14515_b1 , w_39778 );
or ( \14815_b0 , \14515_b0 , \14532_b0 );
not ( \14532_b0 , w_39779 );
and ( w_39779 , w_39778 , \14532_b1 );
or ( \14816_b1 , \14815_b1 , w_39781 );
not ( w_39781 , w_39782 );
and ( \14816_b0 , \14815_b0 , w_39783 );
and ( w_39782 ,  , w_39783 );
buf ( w_39781 , \14540_b1 );
not ( w_39781 , w_39784 );
not (  , w_39785 );
and ( w_39784 , w_39785 , \14540_b0 );
or ( \14817_b1 , \14814_b1 , w_39787 );
not ( w_39787 , w_39788 );
and ( \14817_b0 , \14814_b0 , w_39789 );
and ( w_39788 ,  , w_39789 );
buf ( w_39787 , \14816_b1 );
not ( w_39787 , w_39790 );
not (  , w_39791 );
and ( w_39790 , w_39791 , \14816_b0 );
buf ( \14818_b1 , \14817_b1 );
not ( \14818_b1 , w_39792 );
not ( \14818_b0 , w_39793 );
and ( w_39792 , w_39793 , \14817_b0 );
or ( \14819_b1 , \14812_b1 , w_39794 );
xor ( \14819_b0 , \14812_b0 , w_39796 );
not ( w_39796 , w_39797 );
and ( w_39797 , w_39794 , w_39795 );
buf ( w_39794 , \14818_b1 );
not ( w_39794 , w_39798 );
not ( w_39795 , w_39799 );
and ( w_39798 , w_39799 , \14818_b0 );
buf ( \14820_b1 , \14819_b1 );
buf ( \14820_b0 , \14819_b0 );
buf ( \14821_b1 , \14820_b1 );
buf ( \14821_b0 , \14820_b0 );
buf ( \14822_b1 , \9173_b1 );
not ( \14822_b1 , w_39800 );
not ( \14822_b0 , w_39801 );
and ( w_39800 , w_39801 , \9173_b0 );
or ( \14823_b1 , \13939_b1 , w_39803 );
not ( w_39803 , w_39804 );
and ( \14823_b0 , \13939_b0 , w_39805 );
and ( w_39804 ,  , w_39805 );
buf ( w_39803 , \14822_b1 );
not ( w_39803 , w_39806 );
not (  , w_39807 );
and ( w_39806 , w_39807 , \14822_b0 );
or ( \14824_b1 , \14559_b1 , w_39809 );
not ( w_39809 , w_39810 );
and ( \14824_b0 , \14559_b0 , w_39811 );
and ( w_39810 ,  , w_39811 );
buf ( w_39809 , \14556_b1 );
not ( w_39809 , w_39812 );
not (  , w_39813 );
and ( w_39812 , w_39813 , \14556_b0 );
or ( \14825_b1 , \14824_b1 , \13842_b1 );
not ( \13842_b1 , w_39814 );
and ( \14825_b0 , \14824_b0 , w_39815 );
and ( w_39814 , w_39815 , \13842_b0 );
or ( \14826_b1 , \14556_b1 , w_39816 );
or ( \14826_b0 , \14556_b0 , \14563_b0 );
not ( \14563_b0 , w_39817 );
and ( w_39817 , w_39816 , \14563_b1 );
or ( \14827_b1 , \14826_b1 , w_39819 );
not ( w_39819 , w_39820 );
and ( \14827_b0 , \14826_b0 , w_39821 );
and ( w_39820 ,  , w_39821 );
buf ( w_39819 , \14567_b1 );
not ( w_39819 , w_39822 );
not (  , w_39823 );
and ( w_39822 , w_39823 , \14567_b0 );
or ( \14828_b1 , \14825_b1 , w_39825 );
not ( w_39825 , w_39826 );
and ( \14828_b0 , \14825_b0 , w_39827 );
and ( w_39826 ,  , w_39827 );
buf ( w_39825 , \14827_b1 );
not ( w_39825 , w_39828 );
not (  , w_39829 );
and ( w_39828 , w_39829 , \14827_b0 );
buf ( \14829_b1 , \14828_b1 );
not ( \14829_b1 , w_39830 );
not ( \14829_b0 , w_39831 );
and ( w_39830 , w_39831 , \14828_b0 );
or ( \14830_b1 , \14823_b1 , w_39832 );
xor ( \14830_b0 , \14823_b0 , w_39834 );
not ( w_39834 , w_39835 );
and ( w_39835 , w_39832 , w_39833 );
buf ( w_39832 , \14829_b1 );
not ( w_39832 , w_39836 );
not ( w_39833 , w_39837 );
and ( w_39836 , w_39837 , \14829_b0 );
buf ( \14831_b1 , \14830_b1 );
buf ( \14831_b0 , \14830_b0 );
buf ( \14832_b1 , \14831_b1 );
buf ( \14832_b0 , \14831_b0 );
buf ( \14833_b1 , \9007_b1 );
not ( \14833_b1 , w_39838 );
not ( \14833_b0 , w_39839 );
and ( w_39838 , w_39839 , \9007_b0 );
or ( \14834_b1 , \13934_b1 , w_39841 );
not ( w_39841 , w_39842 );
and ( \14834_b0 , \13934_b0 , w_39843 );
and ( w_39842 ,  , w_39843 );
buf ( w_39841 , \14833_b1 );
not ( w_39841 , w_39844 );
not (  , w_39845 );
and ( w_39844 , w_39845 , \14833_b0 );
or ( \14835_b1 , \14582_b1 , w_39847 );
not ( w_39847 , w_39848 );
and ( \14835_b0 , \14582_b0 , w_39849 );
and ( w_39848 ,  , w_39849 );
buf ( w_39847 , \14579_b1 );
not ( w_39847 , w_39850 );
not (  , w_39851 );
and ( w_39850 , w_39851 , \14579_b0 );
or ( \14836_b1 , \14835_b1 , \14080_b1 );
not ( \14080_b1 , w_39852 );
and ( \14836_b0 , \14835_b0 , w_39853 );
and ( w_39852 , w_39853 , \14080_b0 );
or ( \14837_b1 , \14579_b1 , w_39854 );
or ( \14837_b0 , \14579_b0 , \14586_b0 );
not ( \14586_b0 , w_39855 );
and ( w_39855 , w_39854 , \14586_b1 );
or ( \14838_b1 , \14837_b1 , w_39857 );
not ( w_39857 , w_39858 );
and ( \14838_b0 , \14837_b0 , w_39859 );
and ( w_39858 ,  , w_39859 );
buf ( w_39857 , \14590_b1 );
not ( w_39857 , w_39860 );
not (  , w_39861 );
and ( w_39860 , w_39861 , \14590_b0 );
or ( \14839_b1 , \14836_b1 , w_39863 );
not ( w_39863 , w_39864 );
and ( \14839_b0 , \14836_b0 , w_39865 );
and ( w_39864 ,  , w_39865 );
buf ( w_39863 , \14838_b1 );
not ( w_39863 , w_39866 );
not (  , w_39867 );
and ( w_39866 , w_39867 , \14838_b0 );
buf ( \14840_b1 , \14839_b1 );
not ( \14840_b1 , w_39868 );
not ( \14840_b0 , w_39869 );
and ( w_39868 , w_39869 , \14839_b0 );
or ( \14841_b1 , \14834_b1 , w_39870 );
xor ( \14841_b0 , \14834_b0 , w_39872 );
not ( w_39872 , w_39873 );
and ( w_39873 , w_39870 , w_39871 );
buf ( w_39870 , \14840_b1 );
not ( w_39870 , w_39874 );
not ( w_39871 , w_39875 );
and ( w_39874 , w_39875 , \14840_b0 );
buf ( \14842_b1 , \14841_b1 );
buf ( \14842_b0 , \14841_b0 );
buf ( \14843_b1 , \14842_b1 );
buf ( \14843_b0 , \14842_b0 );
buf ( \14844_b1 , \8846_b1 );
not ( \14844_b1 , w_39876 );
not ( \14844_b0 , w_39877 );
and ( w_39876 , w_39877 , \8846_b0 );
or ( \14845_b1 , \13932_b1 , w_39879 );
not ( w_39879 , w_39880 );
and ( \14845_b0 , \13932_b0 , w_39881 );
and ( w_39880 ,  , w_39881 );
buf ( w_39879 , \14844_b1 );
not ( w_39879 , w_39882 );
not (  , w_39883 );
and ( w_39882 , w_39883 , \14844_b0 );
or ( \14846_b1 , \14605_b1 , w_39885 );
not ( w_39885 , w_39886 );
and ( \14846_b0 , \14605_b0 , w_39887 );
and ( w_39886 ,  , w_39887 );
buf ( w_39885 , \14602_b1 );
not ( w_39885 , w_39888 );
not (  , w_39889 );
and ( w_39888 , w_39889 , \14602_b0 );
or ( \14847_b1 , \14846_b1 , \14226_b1 );
not ( \14226_b1 , w_39890 );
and ( \14847_b0 , \14846_b0 , w_39891 );
and ( w_39890 , w_39891 , \14226_b0 );
or ( \14848_b1 , \14602_b1 , w_39892 );
or ( \14848_b0 , \14602_b0 , \14608_b0 );
not ( \14608_b0 , w_39893 );
and ( w_39893 , w_39892 , \14608_b1 );
or ( \14849_b1 , \14848_b1 , w_39895 );
not ( w_39895 , w_39896 );
and ( \14849_b0 , \14848_b0 , w_39897 );
and ( w_39896 ,  , w_39897 );
buf ( w_39895 , \14612_b1 );
not ( w_39895 , w_39898 );
not (  , w_39899 );
and ( w_39898 , w_39899 , \14612_b0 );
or ( \14850_b1 , \14847_b1 , w_39901 );
not ( w_39901 , w_39902 );
and ( \14850_b0 , \14847_b0 , w_39903 );
and ( w_39902 ,  , w_39903 );
buf ( w_39901 , \14849_b1 );
not ( w_39901 , w_39904 );
not (  , w_39905 );
and ( w_39904 , w_39905 , \14849_b0 );
buf ( \14851_b1 , \14850_b1 );
not ( \14851_b1 , w_39906 );
not ( \14851_b0 , w_39907 );
and ( w_39906 , w_39907 , \14850_b0 );
or ( \14852_b1 , \14845_b1 , w_39908 );
xor ( \14852_b0 , \14845_b0 , w_39910 );
not ( w_39910 , w_39911 );
and ( w_39911 , w_39908 , w_39909 );
buf ( w_39908 , \14851_b1 );
not ( w_39908 , w_39912 );
not ( w_39909 , w_39913 );
and ( w_39912 , w_39913 , \14851_b0 );
buf ( \14853_b1 , \14852_b1 );
buf ( \14853_b0 , \14852_b0 );
buf ( \14854_b1 , \14853_b1 );
buf ( \14854_b0 , \14853_b0 );
buf ( \14855_b1 , \8682_b1 );
not ( \14855_b1 , w_39914 );
not ( \14855_b0 , w_39915 );
and ( w_39914 , w_39915 , \8682_b0 );
or ( \14856_b1 , \13929_b1 , w_39917 );
not ( w_39917 , w_39918 );
and ( \14856_b0 , \13929_b0 , w_39919 );
and ( w_39918 ,  , w_39919 );
buf ( w_39917 , \14855_b1 );
not ( w_39917 , w_39920 );
not (  , w_39921 );
and ( w_39920 , w_39921 , \14855_b0 );
or ( \14857_b1 , \14627_b1 , w_39923 );
not ( w_39923 , w_39924 );
and ( \14857_b0 , \14627_b0 , w_39925 );
and ( w_39924 ,  , w_39925 );
buf ( w_39923 , \14624_b1 );
not ( w_39923 , w_39926 );
not (  , w_39927 );
and ( w_39926 , w_39927 , \14624_b0 );
or ( \14858_b1 , \14857_b1 , \14317_b1 );
not ( \14317_b1 , w_39928 );
and ( \14858_b0 , \14857_b0 , w_39929 );
and ( w_39928 , w_39929 , \14317_b0 );
or ( \14859_b1 , \14624_b1 , w_39930 );
or ( \14859_b0 , \14624_b0 , \14630_b0 );
not ( \14630_b0 , w_39931 );
and ( w_39931 , w_39930 , \14630_b1 );
or ( \14860_b1 , \14859_b1 , w_39933 );
not ( w_39933 , w_39934 );
and ( \14860_b0 , \14859_b0 , w_39935 );
and ( w_39934 ,  , w_39935 );
buf ( w_39933 , \14634_b1 );
not ( w_39933 , w_39936 );
not (  , w_39937 );
and ( w_39936 , w_39937 , \14634_b0 );
or ( \14861_b1 , \14858_b1 , w_39939 );
not ( w_39939 , w_39940 );
and ( \14861_b0 , \14858_b0 , w_39941 );
and ( w_39940 ,  , w_39941 );
buf ( w_39939 , \14860_b1 );
not ( w_39939 , w_39942 );
not (  , w_39943 );
and ( w_39942 , w_39943 , \14860_b0 );
buf ( \14862_b1 , \14861_b1 );
not ( \14862_b1 , w_39944 );
not ( \14862_b0 , w_39945 );
and ( w_39944 , w_39945 , \14861_b0 );
or ( \14863_b1 , \14856_b1 , w_39946 );
xor ( \14863_b0 , \14856_b0 , w_39948 );
not ( w_39948 , w_39949 );
and ( w_39949 , w_39946 , w_39947 );
buf ( w_39946 , \14862_b1 );
not ( w_39946 , w_39950 );
not ( w_39947 , w_39951 );
and ( w_39950 , w_39951 , \14862_b0 );
buf ( \14864_b1 , \14863_b1 );
buf ( \14864_b0 , \14863_b0 );
buf ( \14865_b1 , \14864_b1 );
buf ( \14865_b0 , \14864_b0 );
buf ( \14866_b1 , \8521_b1 );
not ( \14866_b1 , w_39952 );
not ( \14866_b0 , w_39953 );
and ( w_39952 , w_39953 , \8521_b0 );
or ( \14867_b1 , \13927_b1 , w_39955 );
not ( w_39955 , w_39956 );
and ( \14867_b0 , \13927_b0 , w_39957 );
and ( w_39956 ,  , w_39957 );
buf ( w_39955 , \14866_b1 );
not ( w_39955 , w_39958 );
not (  , w_39959 );
and ( w_39958 , w_39959 , \14866_b0 );
or ( \14868_b1 , \14649_b1 , w_39961 );
not ( w_39961 , w_39962 );
and ( \14868_b0 , \14649_b0 , w_39963 );
and ( w_39962 ,  , w_39963 );
buf ( w_39961 , \14646_b1 );
not ( w_39961 , w_39964 );
not (  , w_39965 );
and ( w_39964 , w_39965 , \14646_b0 );
or ( \14869_b1 , \14868_b1 , \13829_b1 );
not ( \13829_b1 , w_39966 );
and ( \14869_b0 , \14868_b0 , w_39967 );
and ( w_39966 , w_39967 , \13829_b0 );
or ( \14870_b1 , \14646_b1 , w_39968 );
or ( \14870_b0 , \14646_b0 , \14652_b0 );
not ( \14652_b0 , w_39969 );
and ( w_39969 , w_39968 , \14652_b1 );
or ( \14871_b1 , \14870_b1 , w_39971 );
not ( w_39971 , w_39972 );
and ( \14871_b0 , \14870_b0 , w_39973 );
and ( w_39972 ,  , w_39973 );
buf ( w_39971 , \14656_b1 );
not ( w_39971 , w_39974 );
not (  , w_39975 );
and ( w_39974 , w_39975 , \14656_b0 );
or ( \14872_b1 , \14869_b1 , w_39977 );
not ( w_39977 , w_39978 );
and ( \14872_b0 , \14869_b0 , w_39979 );
and ( w_39978 ,  , w_39979 );
buf ( w_39977 , \14871_b1 );
not ( w_39977 , w_39980 );
not (  , w_39981 );
and ( w_39980 , w_39981 , \14871_b0 );
buf ( \14873_b1 , \14872_b1 );
not ( \14873_b1 , w_39982 );
not ( \14873_b0 , w_39983 );
and ( w_39982 , w_39983 , \14872_b0 );
or ( \14874_b1 , \14867_b1 , w_39984 );
xor ( \14874_b0 , \14867_b0 , w_39986 );
not ( w_39986 , w_39987 );
and ( w_39987 , w_39984 , w_39985 );
buf ( w_39984 , \14873_b1 );
not ( w_39984 , w_39988 );
not ( w_39985 , w_39989 );
and ( w_39988 , w_39989 , \14873_b0 );
buf ( \14875_b1 , \14874_b1 );
buf ( \14875_b0 , \14874_b0 );
buf ( \14876_b1 , \14875_b1 );
buf ( \14876_b0 , \14875_b0 );
buf ( \14877_b1 , \8359_b1 );
not ( \14877_b1 , w_39990 );
not ( \14877_b0 , w_39991 );
and ( w_39990 , w_39991 , \8359_b0 );
or ( \14878_b1 , \13923_b1 , w_39993 );
not ( w_39993 , w_39994 );
and ( \14878_b0 , \13923_b0 , w_39995 );
and ( w_39994 ,  , w_39995 );
buf ( w_39993 , \14877_b1 );
not ( w_39993 , w_39996 );
not (  , w_39997 );
and ( w_39996 , w_39997 , \14877_b0 );
or ( \14879_b1 , \14671_b1 , w_39999 );
not ( w_39999 , w_40000 );
and ( \14879_b0 , \14671_b0 , w_40001 );
and ( w_40000 ,  , w_40001 );
buf ( w_39999 , \14668_b1 );
not ( w_39999 , w_40002 );
not (  , w_40003 );
and ( w_40002 , w_40003 , \14668_b0 );
or ( \14880_b1 , \14879_b1 , \14314_b1 );
not ( \14314_b1 , w_40004 );
and ( \14880_b0 , \14879_b0 , w_40005 );
and ( w_40004 , w_40005 , \14314_b0 );
or ( \14881_b1 , \14668_b1 , w_40006 );
or ( \14881_b0 , \14668_b0 , \14674_b0 );
not ( \14674_b0 , w_40007 );
and ( w_40007 , w_40006 , \14674_b1 );
or ( \14882_b1 , \14881_b1 , w_40009 );
not ( w_40009 , w_40010 );
and ( \14882_b0 , \14881_b0 , w_40011 );
and ( w_40010 ,  , w_40011 );
buf ( w_40009 , \14678_b1 );
not ( w_40009 , w_40012 );
not (  , w_40013 );
and ( w_40012 , w_40013 , \14678_b0 );
or ( \14883_b1 , \14880_b1 , w_40015 );
not ( w_40015 , w_40016 );
and ( \14883_b0 , \14880_b0 , w_40017 );
and ( w_40016 ,  , w_40017 );
buf ( w_40015 , \14882_b1 );
not ( w_40015 , w_40018 );
not (  , w_40019 );
and ( w_40018 , w_40019 , \14882_b0 );
buf ( \14884_b1 , \14883_b1 );
not ( \14884_b1 , w_40020 );
not ( \14884_b0 , w_40021 );
and ( w_40020 , w_40021 , \14883_b0 );
or ( \14885_b1 , \14878_b1 , w_40022 );
xor ( \14885_b0 , \14878_b0 , w_40024 );
not ( w_40024 , w_40025 );
and ( w_40025 , w_40022 , w_40023 );
buf ( w_40022 , \14884_b1 );
not ( w_40022 , w_40026 );
not ( w_40023 , w_40027 );
and ( w_40026 , w_40027 , \14884_b0 );
buf ( \14886_b1 , \14885_b1 );
buf ( \14886_b0 , \14885_b0 );
buf ( \14887_b1 , \14886_b1 );
buf ( \14887_b0 , \14886_b0 );
buf ( \14888_b1 , \8200_b1 );
not ( \14888_b1 , w_40028 );
not ( \14888_b0 , w_40029 );
and ( w_40028 , w_40029 , \8200_b0 );
or ( \14889_b1 , \13921_b1 , w_40031 );
not ( w_40031 , w_40032 );
and ( \14889_b0 , \13921_b0 , w_40033 );
and ( w_40032 ,  , w_40033 );
buf ( w_40031 , \14888_b1 );
not ( w_40031 , w_40034 );
not (  , w_40035 );
and ( w_40034 , w_40035 , \14888_b0 );
or ( \14890_b1 , \14690_b1 , w_40036 );
or ( \14890_b0 , \14690_b0 , \14694_b0 );
not ( \14694_b0 , w_40037 );
and ( w_40037 , w_40036 , \14694_b1 );
or ( \14891_b1 , \14890_b1 , w_40039 );
not ( w_40039 , w_40040 );
and ( \14891_b0 , \14890_b0 , w_40041 );
and ( w_40040 ,  , w_40041 );
buf ( w_40039 , \14698_b1 );
not ( w_40039 , w_40042 );
not (  , w_40043 );
and ( w_40042 , w_40043 , \14698_b0 );
or ( \14892_b1 , \14889_b1 , w_40044 );
xor ( \14892_b0 , \14889_b0 , w_40046 );
not ( w_40046 , w_40047 );
and ( w_40047 , w_40044 , w_40045 );
buf ( w_40044 , \14891_b1 );
not ( w_40044 , w_40048 );
not ( w_40045 , w_40049 );
and ( w_40048 , w_40049 , \14891_b0 );
buf ( \14893_b1 , \14892_b1 );
buf ( \14893_b0 , \14892_b0 );
buf ( \14894_b1 , \14893_b1 );
buf ( \14894_b0 , \14893_b0 );
buf ( \14895_b1 , \8041_b1 );
not ( \14895_b1 , w_40050 );
not ( \14895_b0 , w_40051 );
and ( w_40050 , w_40051 , \8041_b0 );
or ( \14896_b1 , \13918_b1 , w_40053 );
not ( w_40053 , w_40054 );
and ( \14896_b0 , \13918_b0 , w_40055 );
and ( w_40054 ,  , w_40055 );
buf ( w_40053 , \14895_b1 );
not ( w_40053 , w_40056 );
not (  , w_40057 );
and ( w_40056 , w_40057 , \14895_b0 );
or ( \14897_b1 , \14710_b1 , w_40058 );
or ( \14897_b0 , \14710_b0 , \14714_b0 );
not ( \14714_b0 , w_40059 );
and ( w_40059 , w_40058 , \14714_b1 );
or ( \14898_b1 , \14897_b1 , w_40061 );
not ( w_40061 , w_40062 );
and ( \14898_b0 , \14897_b0 , w_40063 );
and ( w_40062 ,  , w_40063 );
buf ( w_40061 , \14718_b1 );
not ( w_40061 , w_40064 );
not (  , w_40065 );
and ( w_40064 , w_40065 , \14718_b0 );
or ( \14899_b1 , \14896_b1 , w_40066 );
xor ( \14899_b0 , \14896_b0 , w_40068 );
not ( w_40068 , w_40069 );
and ( w_40069 , w_40066 , w_40067 );
buf ( w_40066 , \14898_b1 );
not ( w_40066 , w_40070 );
not ( w_40067 , w_40071 );
and ( w_40070 , w_40071 , \14898_b0 );
buf ( \14900_b1 , \14899_b1 );
buf ( \14900_b0 , \14899_b0 );
buf ( \14901_b1 , \14900_b1 );
buf ( \14901_b0 , \14900_b0 );
buf ( \14902_b1 , \7887_b1 );
not ( \14902_b1 , w_40072 );
not ( \14902_b0 , w_40073 );
and ( w_40072 , w_40073 , \7887_b0 );
or ( \14903_b1 , \13916_b1 , w_40075 );
not ( w_40075 , w_40076 );
and ( \14903_b0 , \13916_b0 , w_40077 );
and ( w_40076 ,  , w_40077 );
buf ( w_40075 , \14902_b1 );
not ( w_40075 , w_40078 );
not (  , w_40079 );
and ( w_40078 , w_40079 , \14902_b0 );
or ( \14904_b1 , \14903_b1 , w_40080 );
xor ( \14904_b0 , \14903_b0 , w_40082 );
not ( w_40082 , w_40083 );
and ( w_40083 , w_40080 , w_40081 );
buf ( w_40080 , \13914_b1 );
not ( w_40080 , w_40084 );
not ( w_40081 , w_40085 );
and ( w_40084 , w_40085 , \13914_b0 );
buf ( \14905_b1 , \14904_b1 );
buf ( \14905_b0 , \14904_b0 );
buf ( \14906_b1 , \14905_b1 );
buf ( \14906_b0 , \14905_b0 );
buf ( \14907_b1 , \13510_b1 );
not ( \14907_b1 , w_40086 );
not ( \14907_b0 , w_40087 );
and ( w_40086 , w_40087 , \13510_b0 );
or ( \14908_b1 , \13909_b1 , w_40089 );
not ( w_40089 , w_40090 );
and ( \14908_b0 , \13909_b0 , w_40091 );
and ( w_40090 ,  , w_40091 );
buf ( w_40089 , \14907_b1 );
not ( w_40089 , w_40092 );
not (  , w_40093 );
and ( w_40092 , w_40093 , \14907_b0 );
or ( \14909_b1 , \14908_b1 , w_40094 );
xor ( \14909_b0 , \14908_b0 , w_40096 );
not ( w_40096 , w_40097 );
and ( w_40097 , w_40094 , w_40095 );
buf ( w_40094 , \14128_b1 );
not ( w_40094 , w_40098 );
not ( w_40095 , w_40099 );
and ( w_40098 , w_40099 , \14128_b0 );
buf ( \14910_b1 , \14909_b1 );
buf ( \14910_b0 , \14909_b0 );
buf ( \14911_b1 , \14910_b1 );
buf ( \14911_b0 , \14910_b0 );
buf ( \14912_b1 , \13503_b1 );
not ( \14912_b1 , w_40100 );
not ( \14912_b0 , w_40101 );
and ( w_40100 , w_40101 , \13503_b0 );
or ( \14913_b1 , \13907_b1 , w_40103 );
not ( w_40103 , w_40104 );
and ( \14913_b0 , \13907_b0 , w_40105 );
and ( w_40104 ,  , w_40105 );
buf ( w_40103 , \14912_b1 );
not ( w_40103 , w_40106 );
not (  , w_40107 );
and ( w_40106 , w_40107 , \14912_b0 );
or ( \14914_b1 , \14913_b1 , w_40108 );
xor ( \14914_b0 , \14913_b0 , w_40110 );
not ( w_40110 , w_40111 );
and ( w_40111 , w_40108 , w_40109 );
buf ( w_40108 , \14250_b1 );
not ( w_40108 , w_40112 );
not ( w_40109 , w_40113 );
and ( w_40112 , w_40113 , \14250_b0 );
buf ( \14915_b1 , \14914_b1 );
buf ( \14915_b0 , \14914_b0 );
buf ( \14916_b1 , \14915_b1 );
buf ( \14916_b0 , \14915_b0 );
buf ( \14917_b1 , \13488_b1 );
not ( \14917_b1 , w_40114 );
not ( \14917_b0 , w_40115 );
and ( w_40114 , w_40115 , \13488_b0 );
or ( \14918_b1 , \13904_b1 , w_40117 );
not ( w_40117 , w_40118 );
and ( \14918_b0 , \13904_b0 , w_40119 );
and ( w_40118 ,  , w_40119 );
buf ( w_40117 , \14917_b1 );
not ( w_40117 , w_40120 );
not (  , w_40121 );
and ( w_40120 , w_40121 , \14917_b0 );
or ( \14919_b1 , \14918_b1 , w_40122 );
xor ( \14919_b0 , \14918_b0 , w_40124 );
not ( w_40124 , w_40125 );
and ( w_40125 , w_40122 , w_40123 );
buf ( w_40122 , \14341_b1 );
not ( w_40122 , w_40126 );
not ( w_40123 , w_40127 );
and ( w_40126 , w_40127 , \14341_b0 );
buf ( \14920_b1 , \14919_b1 );
buf ( \14920_b0 , \14919_b0 );
buf ( \14921_b1 , \14920_b1 );
buf ( \14921_b0 , \14920_b0 );
buf ( \14922_b1 , \13463_b1 );
not ( \14922_b1 , w_40128 );
not ( \14922_b0 , w_40129 );
and ( w_40128 , w_40129 , \13463_b0 );
or ( \14923_b1 , \13902_b1 , w_40131 );
not ( w_40131 , w_40132 );
and ( \14923_b0 , \13902_b0 , w_40133 );
and ( w_40132 ,  , w_40133 );
buf ( w_40131 , \14922_b1 );
not ( w_40131 , w_40134 );
not (  , w_40135 );
and ( w_40134 , w_40135 , \14922_b0 );
or ( \14924_b1 , \14923_b1 , w_40136 );
xor ( \14924_b0 , \14923_b0 , w_40138 );
not ( w_40138 , w_40139 );
and ( w_40139 , w_40136 , w_40137 );
buf ( w_40136 , \14402_b1 );
not ( w_40136 , w_40140 );
not ( w_40137 , w_40141 );
and ( w_40140 , w_40141 , \14402_b0 );
buf ( \14925_b1 , \14924_b1 );
buf ( \14925_b0 , \14924_b0 );
buf ( \14926_b1 , \14925_b1 );
buf ( \14926_b0 , \14925_b0 );
buf ( \14927_b1 , \13428_b1 );
not ( \14927_b1 , w_40142 );
not ( \14927_b0 , w_40143 );
and ( w_40142 , w_40143 , \13428_b0 );
or ( \14928_b1 , \13898_b1 , w_40145 );
not ( w_40145 , w_40146 );
and ( \14928_b0 , \13898_b0 , w_40147 );
and ( w_40146 ,  , w_40147 );
buf ( w_40145 , \14927_b1 );
not ( w_40145 , w_40148 );
not (  , w_40149 );
and ( w_40148 , w_40149 , \14927_b0 );
or ( \14929_b1 , \14928_b1 , w_40150 );
xor ( \14929_b0 , \14928_b0 , w_40152 );
not ( w_40152 , w_40153 );
and ( w_40153 , w_40150 , w_40151 );
buf ( w_40150 , \14447_b1 );
not ( w_40150 , w_40154 );
not ( w_40151 , w_40155 );
and ( w_40154 , w_40155 , \14447_b0 );
buf ( \14930_b1 , \14929_b1 );
buf ( \14930_b0 , \14929_b0 );
buf ( \14931_b1 , \14930_b1 );
buf ( \14931_b0 , \14930_b0 );
buf ( \14932_b1 , \13383_b1 );
not ( \14932_b1 , w_40156 );
not ( \14932_b0 , w_40157 );
and ( w_40156 , w_40157 , \13383_b0 );
or ( \14933_b1 , \13896_b1 , w_40159 );
not ( w_40159 , w_40160 );
and ( \14933_b0 , \13896_b0 , w_40161 );
and ( w_40160 ,  , w_40161 );
buf ( w_40159 , \14932_b1 );
not ( w_40159 , w_40162 );
not (  , w_40163 );
and ( w_40162 , w_40163 , \14932_b0 );
or ( \14934_b1 , \14933_b1 , w_40164 );
xor ( \14934_b0 , \14933_b0 , w_40166 );
not ( w_40166 , w_40167 );
and ( w_40167 , w_40164 , w_40165 );
buf ( w_40164 , \14490_b1 );
not ( w_40164 , w_40168 );
not ( w_40165 , w_40169 );
and ( w_40168 , w_40169 , \14490_b0 );
buf ( \14935_b1 , \14934_b1 );
buf ( \14935_b0 , \14934_b0 );
buf ( \14936_b1 , \14935_b1 );
buf ( \14936_b0 , \14935_b0 );
buf ( \14937_b1 , \13309_b1 );
not ( \14937_b1 , w_40170 );
not ( \14937_b0 , w_40171 );
and ( w_40170 , w_40171 , \13309_b0 );
or ( \14938_b1 , \13893_b1 , w_40173 );
not ( w_40173 , w_40174 );
and ( \14938_b0 , \13893_b0 , w_40175 );
and ( w_40174 ,  , w_40175 );
buf ( w_40173 , \14937_b1 );
not ( w_40173 , w_40176 );
not (  , w_40177 );
and ( w_40176 , w_40177 , \14937_b0 );
or ( \14939_b1 , \14938_b1 , w_40178 );
xor ( \14939_b0 , \14938_b0 , w_40180 );
not ( w_40180 , w_40181 );
and ( w_40181 , w_40178 , w_40179 );
buf ( w_40178 , \14533_b1 );
not ( w_40178 , w_40182 );
not ( w_40179 , w_40183 );
and ( w_40182 , w_40183 , \14533_b0 );
buf ( \14940_b1 , \14939_b1 );
buf ( \14940_b0 , \14939_b0 );
buf ( \14941_b1 , \14940_b1 );
buf ( \14941_b0 , \14940_b0 );
buf ( \14942_b1 , \13194_b1 );
not ( \14942_b1 , w_40184 );
not ( \14942_b0 , w_40185 );
and ( w_40184 , w_40185 , \13194_b0 );
or ( \14943_b1 , \13891_b1 , w_40187 );
not ( w_40187 , w_40188 );
and ( \14943_b0 , \13891_b0 , w_40189 );
and ( w_40188 ,  , w_40189 );
buf ( w_40187 , \14942_b1 );
not ( w_40187 , w_40190 );
not (  , w_40191 );
and ( w_40190 , w_40191 , \14942_b0 );
or ( \14944_b1 , \14943_b1 , w_40192 );
xor ( \14944_b0 , \14943_b0 , w_40194 );
not ( w_40194 , w_40195 );
and ( w_40195 , w_40192 , w_40193 );
buf ( w_40192 , \14564_b1 );
not ( w_40192 , w_40196 );
not ( w_40193 , w_40197 );
and ( w_40196 , w_40197 , \14564_b0 );
buf ( \14945_b1 , \14944_b1 );
buf ( \14945_b0 , \14944_b0 );
buf ( \14946_b1 , \14945_b1 );
buf ( \14946_b0 , \14945_b0 );
buf ( \14947_b1 , \13080_b1 );
not ( \14947_b1 , w_40198 );
not ( \14947_b0 , w_40199 );
and ( w_40198 , w_40199 , \13080_b0 );
or ( \14948_b1 , \13886_b1 , w_40201 );
not ( w_40201 , w_40202 );
and ( \14948_b0 , \13886_b0 , w_40203 );
and ( w_40202 ,  , w_40203 );
buf ( w_40201 , \14947_b1 );
not ( w_40201 , w_40204 );
not (  , w_40205 );
and ( w_40204 , w_40205 , \14947_b0 );
or ( \14949_b1 , \14948_b1 , w_40206 );
xor ( \14949_b0 , \14948_b0 , w_40208 );
not ( w_40208 , w_40209 );
and ( w_40209 , w_40206 , w_40207 );
buf ( w_40206 , \14587_b1 );
not ( w_40206 , w_40210 );
not ( w_40207 , w_40211 );
and ( w_40210 , w_40211 , \14587_b0 );
buf ( \14950_b1 , \14949_b1 );
buf ( \14950_b0 , \14949_b0 );
buf ( \14951_b1 , \14950_b1 );
buf ( \14951_b0 , \14950_b0 );
buf ( \14952_b1 , \12975_b1 );
not ( \14952_b1 , w_40212 );
not ( \14952_b0 , w_40213 );
and ( w_40212 , w_40213 , \12975_b0 );
or ( \14953_b1 , \13884_b1 , w_40215 );
not ( w_40215 , w_40216 );
and ( \14953_b0 , \13884_b0 , w_40217 );
and ( w_40216 ,  , w_40217 );
buf ( w_40215 , \14952_b1 );
not ( w_40215 , w_40218 );
not (  , w_40219 );
and ( w_40218 , w_40219 , \14952_b0 );
or ( \14954_b1 , \14953_b1 , w_40220 );
xor ( \14954_b0 , \14953_b0 , w_40222 );
not ( w_40222 , w_40223 );
and ( w_40223 , w_40220 , w_40221 );
buf ( w_40220 , \14609_b1 );
not ( w_40220 , w_40224 );
not ( w_40221 , w_40225 );
and ( w_40224 , w_40225 , \14609_b0 );
buf ( \14955_b1 , \14954_b1 );
buf ( \14955_b0 , \14954_b0 );
buf ( \14956_b1 , \14955_b1 );
buf ( \14956_b0 , \14955_b0 );
buf ( \14957_b1 , \12873_b1 );
not ( \14957_b1 , w_40226 );
not ( \14957_b0 , w_40227 );
and ( w_40226 , w_40227 , \12873_b0 );
or ( \14958_b1 , \13881_b1 , w_40229 );
not ( w_40229 , w_40230 );
and ( \14958_b0 , \13881_b0 , w_40231 );
and ( w_40230 ,  , w_40231 );
buf ( w_40229 , \14957_b1 );
not ( w_40229 , w_40232 );
not (  , w_40233 );
and ( w_40232 , w_40233 , \14957_b0 );
or ( \14959_b1 , \14958_b1 , w_40234 );
xor ( \14959_b0 , \14958_b0 , w_40236 );
not ( w_40236 , w_40237 );
and ( w_40237 , w_40234 , w_40235 );
buf ( w_40234 , \14631_b1 );
not ( w_40234 , w_40238 );
not ( w_40235 , w_40239 );
and ( w_40238 , w_40239 , \14631_b0 );
buf ( \14960_b1 , \14959_b1 );
buf ( \14960_b0 , \14959_b0 );
buf ( \14961_b1 , \14960_b1 );
buf ( \14961_b0 , \14960_b0 );
buf ( \14962_b1 , \12778_b1 );
not ( \14962_b1 , w_40240 );
not ( \14962_b0 , w_40241 );
and ( w_40240 , w_40241 , \12778_b0 );
or ( \14963_b1 , \13879_b1 , w_40243 );
not ( w_40243 , w_40244 );
and ( \14963_b0 , \13879_b0 , w_40245 );
and ( w_40244 ,  , w_40245 );
buf ( w_40243 , \14962_b1 );
not ( w_40243 , w_40246 );
not (  , w_40247 );
and ( w_40246 , w_40247 , \14962_b0 );
or ( \14964_b1 , \14963_b1 , w_40248 );
xor ( \14964_b0 , \14963_b0 , w_40250 );
not ( w_40250 , w_40251 );
and ( w_40251 , w_40248 , w_40249 );
buf ( w_40248 , \14653_b1 );
not ( w_40248 , w_40252 );
not ( w_40249 , w_40253 );
and ( w_40252 , w_40253 , \14653_b0 );
buf ( \14965_b1 , \14964_b1 );
buf ( \14965_b0 , \14964_b0 );
buf ( \14966_b1 , \14965_b1 );
buf ( \14966_b0 , \14965_b0 );
buf ( \14967_b1 , \12685_b1 );
not ( \14967_b1 , w_40254 );
not ( \14967_b0 , w_40255 );
and ( w_40254 , w_40255 , \12685_b0 );
or ( \14968_b1 , \13875_b1 , w_40257 );
not ( w_40257 , w_40258 );
and ( \14968_b0 , \13875_b0 , w_40259 );
and ( w_40258 ,  , w_40259 );
buf ( w_40257 , \14967_b1 );
not ( w_40257 , w_40260 );
not (  , w_40261 );
and ( w_40260 , w_40261 , \14967_b0 );
or ( \14969_b1 , \14968_b1 , w_40262 );
xor ( \14969_b0 , \14968_b0 , w_40264 );
not ( w_40264 , w_40265 );
and ( w_40265 , w_40262 , w_40263 );
buf ( w_40262 , \14675_b1 );
not ( w_40262 , w_40266 );
not ( w_40263 , w_40267 );
and ( w_40266 , w_40267 , \14675_b0 );
buf ( \14970_b1 , \14969_b1 );
buf ( \14970_b0 , \14969_b0 );
buf ( \14971_b1 , \14970_b1 );
buf ( \14971_b0 , \14970_b0 );
buf ( \14972_b1 , \12600_b1 );
not ( \14972_b1 , w_40268 );
not ( \14972_b0 , w_40269 );
and ( w_40268 , w_40269 , \12600_b0 );
or ( \14973_b1 , \13873_b1 , w_40271 );
not ( w_40271 , w_40272 );
and ( \14973_b0 , \13873_b0 , w_40273 );
and ( w_40272 ,  , w_40273 );
buf ( w_40271 , \14972_b1 );
not ( w_40271 , w_40274 );
not (  , w_40275 );
and ( w_40274 , w_40275 , \14972_b0 );
or ( \14974_b1 , \14973_b1 , w_40276 );
xor ( \14974_b0 , \14973_b0 , w_40278 );
not ( w_40278 , w_40279 );
and ( w_40279 , w_40276 , w_40277 );
buf ( w_40276 , \14695_b1 );
not ( w_40276 , w_40280 );
not ( w_40277 , w_40281 );
and ( w_40280 , w_40281 , \14695_b0 );
buf ( \14975_b1 , \14974_b1 );
buf ( \14975_b0 , \14974_b0 );
buf ( \14976_b1 , \14975_b1 );
buf ( \14976_b0 , \14975_b0 );
buf ( \14977_b1 , \12518_b1 );
not ( \14977_b1 , w_40282 );
not ( \14977_b0 , w_40283 );
and ( w_40282 , w_40283 , \12518_b0 );
or ( \14978_b1 , \13870_b1 , w_40285 );
not ( w_40285 , w_40286 );
and ( \14978_b0 , \13870_b0 , w_40287 );
and ( w_40286 ,  , w_40287 );
buf ( w_40285 , \14977_b1 );
not ( w_40285 , w_40288 );
not (  , w_40289 );
and ( w_40288 , w_40289 , \14977_b0 );
or ( \14979_b1 , \14978_b1 , w_40290 );
xor ( \14979_b0 , \14978_b0 , w_40292 );
not ( w_40292 , w_40293 );
and ( w_40293 , w_40290 , w_40291 );
buf ( w_40290 , \14715_b1 );
not ( w_40290 , w_40294 );
not ( w_40291 , w_40295 );
and ( w_40294 , w_40295 , \14715_b0 );
buf ( \14980_b1 , \14979_b1 );
buf ( \14980_b0 , \14979_b0 );
buf ( \14981_b1 , \14980_b1 );
buf ( \14981_b0 , \14980_b0 );
buf ( \14982_b1 , \12443_b1 );
not ( \14982_b1 , w_40296 );
not ( \14982_b0 , w_40297 );
and ( w_40296 , w_40297 , \12443_b0 );
or ( \14983_b1 , \13868_b1 , w_40299 );
not ( w_40299 , w_40300 );
and ( \14983_b0 , \13868_b0 , w_40301 );
and ( w_40300 ,  , w_40301 );
buf ( w_40299 , \14982_b1 );
not ( w_40299 , w_40302 );
not (  , w_40303 );
and ( w_40302 , w_40303 , \14982_b0 );
or ( \14984_b1 , \14983_b1 , w_40304 );
xor ( \14984_b0 , \14983_b0 , w_40306 );
not ( w_40306 , w_40307 );
and ( w_40307 , w_40304 , w_40305 );
buf ( w_40304 , \14731_b1 );
not ( w_40304 , w_40308 );
not ( w_40305 , w_40309 );
and ( w_40308 , w_40309 , \14731_b0 );
buf ( \14985_b1 , \14984_b1 );
buf ( \14985_b0 , \14984_b0 );
buf ( \14986_b1 , \14985_b1 );
buf ( \14986_b0 , \14985_b0 );
buf ( \14987_b1 , \13765_b1 );
not ( \14987_b1 , w_40310 );
not ( \14987_b0 , w_40311 );
and ( w_40310 , w_40311 , \13765_b0 );
or ( \14988_b1 , \13862_b1 , w_40313 );
not ( w_40313 , w_40314 );
and ( \14988_b0 , \13862_b0 , w_40315 );
and ( w_40314 ,  , w_40315 );
buf ( w_40313 , \14987_b1 );
not ( w_40313 , w_40316 );
not (  , w_40317 );
and ( w_40316 , w_40317 , \14987_b0 );
or ( \14989_b1 , \14988_b1 , w_40318 );
xor ( \14989_b0 , \14988_b0 , w_40320 );
not ( w_40320 , w_40321 );
and ( w_40321 , w_40318 , w_40319 );
buf ( w_40318 , \14743_b1 );
not ( w_40318 , w_40322 );
not ( w_40319 , w_40323 );
and ( w_40322 , w_40323 , \14743_b0 );
buf ( \14990_b1 , \14989_b1 );
buf ( \14990_b0 , \14989_b0 );
buf ( \14991_b1 , \14990_b1 );
buf ( \14991_b0 , \14990_b0 );
buf ( \14992_b1 , \13758_b1 );
not ( \14992_b1 , w_40324 );
not ( \14992_b0 , w_40325 );
and ( w_40324 , w_40325 , \13758_b0 );
or ( \14993_b1 , \13860_b1 , w_40327 );
not ( w_40327 , w_40328 );
and ( \14993_b0 , \13860_b0 , w_40329 );
and ( w_40328 ,  , w_40329 );
buf ( w_40327 , \14992_b1 );
not ( w_40327 , w_40330 );
not (  , w_40331 );
and ( w_40330 , w_40331 , \14992_b0 );
or ( \14994_b1 , \14993_b1 , w_40332 );
xor ( \14994_b0 , \14993_b0 , w_40334 );
not ( w_40334 , w_40335 );
and ( w_40335 , w_40332 , w_40333 );
buf ( w_40332 , \14755_b1 );
not ( w_40332 , w_40336 );
not ( w_40333 , w_40337 );
and ( w_40336 , w_40337 , \14755_b0 );
buf ( \14995_b1 , \14994_b1 );
buf ( \14995_b0 , \14994_b0 );
buf ( \14996_b1 , \14995_b1 );
buf ( \14996_b0 , \14995_b0 );
buf ( \14997_b1 , \13746_b1 );
not ( \14997_b1 , w_40338 );
not ( \14997_b0 , w_40339 );
and ( w_40338 , w_40339 , \13746_b0 );
or ( \14998_b1 , \13857_b1 , w_40341 );
not ( w_40341 , w_40342 );
and ( \14998_b0 , \13857_b0 , w_40343 );
and ( w_40342 ,  , w_40343 );
buf ( w_40341 , \14997_b1 );
not ( w_40341 , w_40344 );
not (  , w_40345 );
and ( w_40344 , w_40345 , \14997_b0 );
or ( \14999_b1 , \14998_b1 , w_40346 );
xor ( \14999_b0 , \14998_b0 , w_40348 );
not ( w_40348 , w_40349 );
and ( w_40349 , w_40346 , w_40347 );
buf ( w_40346 , \14767_b1 );
not ( w_40346 , w_40350 );
not ( w_40347 , w_40351 );
and ( w_40350 , w_40351 , \14767_b0 );
buf ( \15000_b1 , \14999_b1 );
buf ( \15000_b0 , \14999_b0 );
buf ( \15001_b1 , \15000_b1 );
buf ( \15001_b0 , \15000_b0 );
buf ( \15002_b1 , \13729_b1 );
not ( \15002_b1 , w_40352 );
not ( \15002_b0 , w_40353 );
and ( w_40352 , w_40353 , \13729_b0 );
or ( \15003_b1 , \13855_b1 , w_40355 );
not ( w_40355 , w_40356 );
and ( \15003_b0 , \13855_b0 , w_40357 );
and ( w_40356 ,  , w_40357 );
buf ( w_40355 , \15002_b1 );
not ( w_40355 , w_40358 );
not (  , w_40359 );
and ( w_40358 , w_40359 , \15002_b0 );
or ( \15004_b1 , \15003_b1 , w_40360 );
xor ( \15004_b0 , \15003_b0 , w_40362 );
not ( w_40362 , w_40363 );
and ( w_40363 , w_40360 , w_40361 );
buf ( w_40360 , \14779_b1 );
not ( w_40360 , w_40364 );
not ( w_40361 , w_40365 );
and ( w_40364 , w_40365 , \14779_b0 );
buf ( \15005_b1 , \15004_b1 );
buf ( \15005_b0 , \15004_b0 );
buf ( \15006_b1 , \15005_b1 );
buf ( \15006_b0 , \15005_b0 );
buf ( \15007_b1 , \13700_b1 );
not ( \15007_b1 , w_40366 );
not ( \15007_b0 , w_40367 );
and ( w_40366 , w_40367 , \13700_b0 );
or ( \15008_b1 , \13851_b1 , w_40369 );
not ( w_40369 , w_40370 );
and ( \15008_b0 , \13851_b0 , w_40371 );
and ( w_40370 ,  , w_40371 );
buf ( w_40369 , \15007_b1 );
not ( w_40369 , w_40372 );
not (  , w_40373 );
and ( w_40372 , w_40373 , \15007_b0 );
or ( \15009_b1 , \15008_b1 , w_40374 );
xor ( \15009_b0 , \15008_b0 , w_40376 );
not ( w_40376 , w_40377 );
and ( w_40377 , w_40374 , w_40375 );
buf ( w_40374 , \14791_b1 );
not ( w_40374 , w_40378 );
not ( w_40375 , w_40379 );
and ( w_40378 , w_40379 , \14791_b0 );
buf ( \15010_b1 , \15009_b1 );
buf ( \15010_b0 , \15009_b0 );
buf ( \15011_b1 , \15010_b1 );
buf ( \15011_b0 , \15010_b0 );
buf ( \15012_b1 , \13655_b1 );
not ( \15012_b1 , w_40380 );
not ( \15012_b0 , w_40381 );
and ( w_40380 , w_40381 , \13655_b0 );
or ( \15013_b1 , \13849_b1 , w_40383 );
not ( w_40383 , w_40384 );
and ( \15013_b0 , \13849_b0 , w_40385 );
and ( w_40384 ,  , w_40385 );
buf ( w_40383 , \15012_b1 );
not ( w_40383 , w_40386 );
not (  , w_40387 );
and ( w_40386 , w_40387 , \15012_b0 );
or ( \15014_b1 , \15013_b1 , w_40388 );
xor ( \15014_b0 , \15013_b0 , w_40390 );
not ( w_40390 , w_40391 );
and ( w_40391 , w_40388 , w_40389 );
buf ( w_40388 , \14481_b1 );
not ( w_40388 , w_40392 );
not ( w_40389 , w_40393 );
and ( w_40392 , w_40393 , \14481_b0 );
buf ( \15015_b1 , \15014_b1 );
buf ( \15015_b0 , \15014_b0 );
buf ( \15016_b1 , \15015_b1 );
buf ( \15016_b0 , \15015_b0 );
buf ( \15017_b1 , \13613_b1 );
not ( \15017_b1 , w_40394 );
not ( \15017_b0 , w_40395 );
and ( w_40394 , w_40395 , \13613_b0 );
or ( \15018_b1 , \13846_b1 , w_40397 );
not ( w_40397 , w_40398 );
and ( \15018_b0 , \13846_b0 , w_40399 );
and ( w_40398 ,  , w_40399 );
buf ( w_40397 , \15017_b1 );
not ( w_40397 , w_40400 );
not (  , w_40401 );
and ( w_40400 , w_40401 , \15017_b0 );
or ( \15019_b1 , \15018_b1 , w_40402 );
xor ( \15019_b0 , \15018_b0 , w_40404 );
not ( w_40404 , w_40405 );
and ( w_40405 , w_40402 , w_40403 );
buf ( w_40402 , \14524_b1 );
not ( w_40402 , w_40406 );
not ( w_40403 , w_40407 );
and ( w_40406 , w_40407 , \14524_b0 );
buf ( \15020_b1 , \15019_b1 );
buf ( \15020_b0 , \15019_b0 );
buf ( \15021_b1 , \15020_b1 );
buf ( \15021_b0 , \15020_b0 );
buf ( \15022_b1 , \13578_b1 );
not ( \15022_b1 , w_40408 );
not ( \15022_b0 , w_40409 );
and ( w_40408 , w_40409 , \13578_b0 );
or ( \15023_b1 , \13844_b1 , w_40411 );
not ( w_40411 , w_40412 );
and ( \15023_b0 , \13844_b0 , w_40413 );
and ( w_40412 ,  , w_40413 );
buf ( w_40411 , \15022_b1 );
not ( w_40411 , w_40414 );
not (  , w_40415 );
and ( w_40414 , w_40415 , \15022_b0 );
or ( \15024_b1 , \15023_b1 , w_40416 );
xor ( \15024_b0 , \15023_b0 , w_40418 );
not ( w_40418 , w_40419 );
and ( w_40419 , w_40416 , w_40417 );
buf ( w_40416 , \13842_b1 );
not ( w_40416 , w_40420 );
not ( w_40417 , w_40421 );
and ( w_40420 , w_40421 , \13842_b0 );
buf ( \15025_b1 , \15024_b1 );
buf ( \15025_b0 , \15024_b0 );
buf ( \15026_b1 , \15025_b1 );
buf ( \15026_b0 , \15025_b0 );
buf ( \15027_b1 , \13812_b1 );
not ( \15027_b1 , w_40422 );
not ( \15027_b0 , w_40423 );
and ( w_40422 , w_40423 , \13812_b0 );
or ( \15028_b1 , \13839_b1 , w_40425 );
not ( w_40425 , w_40426 );
and ( \15028_b0 , \13839_b0 , w_40427 );
and ( w_40426 ,  , w_40427 );
buf ( w_40425 , \15027_b1 );
not ( w_40425 , w_40428 );
not (  , w_40429 );
and ( w_40428 , w_40429 , \15027_b0 );
or ( \15029_b1 , \15028_b1 , w_40430 );
xor ( \15029_b0 , \15028_b0 , w_40432 );
not ( w_40432 , w_40433 );
and ( w_40433 , w_40430 , w_40431 );
buf ( w_40430 , \14080_b1 );
not ( w_40430 , w_40434 );
not ( w_40431 , w_40435 );
and ( w_40434 , w_40435 , \14080_b0 );
buf ( \15030_b1 , \15029_b1 );
buf ( \15030_b0 , \15029_b0 );
buf ( \15031_b1 , \15030_b1 );
buf ( \15031_b0 , \15030_b0 );
or ( \342_b1 , \322_b1 , w_40438 );
or ( \342_b0 , \322_b0 , w_40437 );
not ( w_40437 , w_40439 );
and ( w_40439 , w_40438 , w_40436 );
or ( w_40436 , \340_b1 , w_40440 );
or ( w_40437 , \340_b0 , \341_b0 );
not ( \341_b0 , w_40441 );
and ( w_40441 , w_40440 , \341_b1 );
or ( \370_b1 , \363_b1 , w_40444 );
or ( \370_b0 , \363_b0 , w_40443 );
not ( w_40443 , w_40445 );
and ( w_40445 , w_40444 , w_40442 );
or ( w_40442 , \368_b1 , w_40446 );
or ( w_40443 , \368_b0 , \369_b0 );
not ( \369_b0 , w_40447 );
and ( w_40447 , w_40446 , \369_b1 );
or ( \388_b1 , \385_b1 , w_40450 );
or ( \388_b0 , \385_b0 , w_40449 );
not ( w_40449 , w_40451 );
and ( w_40451 , w_40450 , w_40448 );
or ( w_40448 , \386_b1 , w_40452 );
or ( w_40449 , \386_b0 , \387_b0 );
not ( \387_b0 , w_40453 );
and ( w_40453 , w_40452 , \387_b1 );
or ( \408_b1 , \384_b1 , w_40456 );
or ( \408_b0 , \384_b0 , w_40455 );
not ( w_40455 , w_40457 );
and ( w_40457 , w_40456 , w_40454 );
or ( w_40454 , \406_b1 , w_40458 );
or ( w_40455 , \406_b0 , \407_b0 );
not ( \407_b0 , w_40459 );
and ( w_40459 , w_40458 , \407_b1 );
or ( \412_b1 , \409_b1 , w_40462 );
or ( \412_b0 , \409_b0 , w_40461 );
not ( w_40461 , w_40463 );
and ( w_40463 , w_40462 , w_40460 );
or ( w_40460 , \410_b1 , w_40464 );
or ( w_40461 , \410_b0 , \411_b0 );
not ( \411_b0 , w_40465 );
and ( w_40465 , w_40464 , \411_b1 );
or ( \428_b1 , \425_b1 , w_40468 );
or ( \428_b0 , \425_b0 , w_40467 );
not ( w_40467 , w_40469 );
and ( w_40469 , w_40468 , w_40466 );
or ( w_40466 , \426_b1 , w_40470 );
or ( w_40467 , \426_b0 , \427_b0 );
not ( \427_b0 , w_40471 );
and ( w_40471 , w_40470 , \427_b1 );
or ( \448_b1 , \443_b1 , w_40474 );
or ( \448_b0 , \443_b0 , w_40473 );
not ( w_40473 , w_40475 );
and ( w_40475 , w_40474 , w_40472 );
or ( w_40472 , \446_b1 , w_40476 );
or ( w_40473 , \446_b0 , \447_b0 );
not ( \447_b0 , w_40477 );
and ( w_40477 , w_40476 , \447_b1 );
or ( \468_b1 , \461_b1 , w_40480 );
or ( \468_b0 , \461_b0 , w_40479 );
not ( w_40479 , w_40481 );
and ( w_40481 , w_40480 , w_40478 );
or ( w_40478 , \466_b1 , w_40482 );
or ( w_40479 , \466_b0 , \467_b0 );
not ( \467_b0 , w_40483 );
and ( w_40483 , w_40482 , \467_b1 );
or ( \473_b1 , \469_b1 , w_40486 );
or ( \473_b0 , \469_b0 , w_40485 );
not ( w_40485 , w_40487 );
and ( w_40487 , w_40486 , w_40484 );
or ( w_40484 , \471_b1 , w_40488 );
or ( w_40485 , \471_b0 , \472_b0 );
not ( \472_b0 , w_40489 );
and ( w_40489 , w_40488 , \472_b1 );
or ( \480_b1 , \476_b1 , w_40492 );
or ( \480_b0 , \476_b0 , w_40491 );
not ( w_40491 , w_40493 );
and ( w_40493 , w_40492 , w_40490 );
or ( w_40490 , \478_b1 , w_40494 );
or ( w_40491 , \478_b0 , \479_b0 );
not ( \479_b0 , w_40495 );
and ( w_40495 , w_40494 , \479_b1 );
or ( \499_b1 , \494_b1 , w_40498 );
or ( \499_b0 , \494_b0 , w_40497 );
not ( w_40497 , w_40499 );
and ( w_40499 , w_40498 , w_40496 );
or ( w_40496 , \497_b1 , w_40500 );
or ( w_40497 , \497_b0 , \498_b0 );
not ( \498_b0 , w_40501 );
and ( w_40501 , w_40500 , \498_b1 );
or ( \518_b1 , \511_b1 , w_40504 );
or ( \518_b0 , \511_b0 , w_40503 );
not ( w_40503 , w_40505 );
and ( w_40505 , w_40504 , w_40502 );
or ( w_40502 , \516_b1 , w_40506 );
or ( w_40503 , \516_b0 , \517_b0 );
not ( \517_b0 , w_40507 );
and ( w_40507 , w_40506 , \517_b1 );
or ( \524_b1 , \519_b1 , w_40510 );
or ( \524_b0 , \519_b0 , w_40509 );
not ( w_40509 , w_40511 );
and ( w_40511 , w_40510 , w_40508 );
or ( w_40508 , \522_b1 , w_40512 );
or ( w_40509 , \522_b0 , \523_b0 );
not ( \523_b0 , w_40513 );
and ( w_40513 , w_40512 , \523_b1 );
or ( \532_b1 , \527_b1 , w_40516 );
or ( \532_b0 , \527_b0 , w_40515 );
not ( w_40515 , w_40517 );
and ( w_40517 , w_40516 , w_40514 );
or ( w_40514 , \530_b1 , w_40518 );
or ( w_40515 , \530_b0 , \531_b0 );
not ( \531_b0 , w_40519 );
and ( w_40519 , w_40518 , \531_b1 );
or ( \554_b1 , \547_b1 , w_40522 );
or ( \554_b0 , \547_b0 , w_40521 );
not ( w_40521 , w_40523 );
and ( w_40523 , w_40522 , w_40520 );
or ( w_40520 , \552_b1 , w_40524 );
or ( w_40521 , \552_b0 , \553_b0 );
not ( \553_b0 , w_40525 );
and ( w_40525 , w_40524 , \553_b1 );
or ( \574_b1 , \567_b1 , w_40528 );
or ( \574_b0 , \567_b0 , w_40527 );
not ( w_40527 , w_40529 );
and ( w_40529 , w_40528 , w_40526 );
or ( w_40526 , \572_b1 , w_40530 );
or ( w_40527 , \572_b0 , \573_b0 );
not ( \573_b0 , w_40531 );
and ( w_40531 , w_40530 , \573_b1 );
or ( \583_b1 , \578_b1 , w_40534 );
or ( \583_b0 , \578_b0 , w_40533 );
not ( w_40533 , w_40535 );
and ( w_40535 , w_40534 , w_40532 );
or ( w_40532 , \581_b1 , w_40536 );
or ( w_40533 , \581_b0 , \582_b0 );
not ( \582_b0 , w_40537 );
and ( w_40537 , w_40536 , \582_b1 );
or ( \600_b1 , \592_b1 , w_40540 );
or ( \600_b0 , \592_b0 , w_40539 );
not ( w_40539 , w_40541 );
and ( w_40541 , w_40540 , w_40538 );
or ( w_40538 , \598_b1 , w_40542 );
or ( w_40539 , \598_b0 , \599_b0 );
not ( \599_b0 , w_40543 );
and ( w_40543 , w_40542 , \599_b1 );
or ( \619_b1 , \612_b1 , w_40546 );
or ( \619_b0 , \612_b0 , w_40545 );
not ( w_40545 , w_40547 );
and ( w_40547 , w_40546 , w_40544 );
or ( w_40544 , \617_b1 , w_40548 );
or ( w_40545 , \617_b0 , \618_b0 );
not ( \618_b0 , w_40549 );
and ( w_40549 , w_40548 , \618_b1 );
or ( \626_b1 , \620_b1 , w_40552 );
or ( \626_b0 , \620_b0 , w_40551 );
not ( w_40551 , w_40553 );
and ( w_40553 , w_40552 , w_40550 );
or ( w_40550 , \624_b1 , w_40554 );
or ( w_40551 , \624_b0 , \625_b0 );
not ( \625_b0 , w_40555 );
and ( w_40555 , w_40554 , \625_b1 );
or ( \635_b1 , \630_b1 , w_40558 );
or ( \635_b0 , \630_b0 , w_40557 );
not ( w_40557 , w_40559 );
and ( w_40559 , w_40558 , w_40556 );
or ( w_40556 , \633_b1 , w_40560 );
or ( w_40557 , \633_b0 , \634_b0 );
not ( \634_b0 , w_40561 );
and ( w_40561 , w_40560 , \634_b1 );
or ( \641_b1 , \636_b1 , w_40564 );
or ( \641_b0 , \636_b0 , w_40563 );
not ( w_40563 , w_40565 );
and ( w_40565 , w_40564 , w_40562 );
or ( w_40562 , \639_b1 , w_40566 );
or ( w_40563 , \639_b0 , \640_b0 );
not ( \640_b0 , w_40567 );
and ( w_40567 , w_40566 , \640_b1 );
or ( \651_b1 , \646_b1 , w_40570 );
or ( \651_b0 , \646_b0 , w_40569 );
not ( w_40569 , w_40571 );
and ( w_40571 , w_40570 , w_40568 );
or ( w_40568 , \649_b1 , w_40572 );
or ( w_40569 , \649_b0 , \650_b0 );
not ( \650_b0 , w_40573 );
and ( w_40573 , w_40572 , \650_b1 );
or ( \657_b1 , \652_b1 , w_40576 );
or ( \657_b0 , \652_b0 , w_40575 );
not ( w_40575 , w_40577 );
and ( w_40577 , w_40576 , w_40574 );
or ( w_40574 , \655_b1 , w_40578 );
or ( w_40575 , \655_b0 , \656_b0 );
not ( \656_b0 , w_40579 );
and ( w_40579 , w_40578 , \656_b1 );
or ( \681_b1 , \674_b1 , w_40582 );
or ( \681_b0 , \674_b0 , w_40581 );
not ( w_40581 , w_40583 );
and ( w_40583 , w_40582 , w_40580 );
or ( w_40580 , \679_b1 , w_40584 );
or ( w_40581 , \679_b0 , \680_b0 );
not ( \680_b0 , w_40585 );
and ( w_40585 , w_40584 , \680_b1 );
or ( \697_b1 , \690_b1 , w_40588 );
or ( \697_b0 , \690_b0 , w_40587 );
not ( w_40587 , w_40589 );
and ( w_40589 , w_40588 , w_40586 );
or ( w_40586 , \695_b1 , w_40590 );
or ( w_40587 , \695_b0 , \696_b0 );
not ( \696_b0 , w_40591 );
and ( w_40591 , w_40590 , \696_b1 );
or ( \708_b1 , \698_b1 , w_40594 );
or ( \708_b0 , \698_b0 , w_40593 );
not ( w_40593 , w_40595 );
and ( w_40595 , w_40594 , w_40592 );
or ( w_40592 , \706_b1 , w_40596 );
or ( w_40593 , \706_b0 , \707_b0 );
not ( \707_b0 , w_40597 );
and ( w_40597 , w_40596 , \707_b1 );
or ( \717_b1 , \713_b1 , w_40600 );
or ( \717_b0 , \713_b0 , w_40599 );
not ( w_40599 , w_40601 );
and ( w_40601 , w_40600 , w_40598 );
or ( w_40598 , \715_b1 , w_40602 );
or ( w_40599 , \715_b0 , \716_b0 );
not ( \716_b0 , w_40603 );
and ( w_40603 , w_40602 , \716_b1 );
or ( \723_b1 , \718_b1 , w_40606 );
or ( \723_b0 , \718_b0 , w_40605 );
not ( w_40605 , w_40607 );
and ( w_40607 , w_40606 , w_40604 );
or ( w_40604 , \721_b1 , w_40608 );
or ( w_40605 , \721_b0 , \722_b0 );
not ( \722_b0 , w_40609 );
and ( w_40609 , w_40608 , \722_b1 );
or ( \730_b1 , \726_b1 , w_40612 );
or ( \730_b0 , \726_b0 , w_40611 );
not ( w_40611 , w_40613 );
and ( w_40613 , w_40612 , w_40610 );
or ( w_40610 , \728_b1 , w_40614 );
or ( w_40611 , \728_b0 , \729_b0 );
not ( \729_b0 , w_40615 );
and ( w_40615 , w_40614 , \729_b1 );
or ( \755_b1 , \748_b1 , w_40618 );
or ( \755_b0 , \748_b0 , w_40617 );
not ( w_40617 , w_40619 );
and ( w_40619 , w_40618 , w_40616 );
or ( w_40616 , \753_b1 , w_40620 );
or ( w_40617 , \753_b0 , \754_b0 );
not ( \754_b0 , w_40621 );
and ( w_40621 , w_40620 , \754_b1 );
or ( \771_b1 , \764_b1 , w_40624 );
or ( \771_b0 , \764_b0 , w_40623 );
not ( w_40623 , w_40625 );
and ( w_40625 , w_40624 , w_40622 );
or ( w_40622 , \769_b1 , w_40626 );
or ( w_40623 , \769_b0 , \770_b0 );
not ( \770_b0 , w_40627 );
and ( w_40627 , w_40626 , \770_b1 );
or ( \782_b1 , \772_b1 , w_40630 );
or ( \782_b0 , \772_b0 , w_40629 );
not ( w_40629 , w_40631 );
and ( w_40631 , w_40630 , w_40628 );
or ( w_40628 , \780_b1 , w_40632 );
or ( w_40629 , \780_b0 , \781_b0 );
not ( \781_b0 , w_40633 );
and ( w_40633 , w_40632 , \781_b1 );
or ( \791_b1 , \787_b1 , w_40636 );
or ( \791_b0 , \787_b0 , w_40635 );
not ( w_40635 , w_40637 );
and ( w_40637 , w_40636 , w_40634 );
or ( w_40634 , \789_b1 , w_40638 );
or ( w_40635 , \789_b0 , \790_b0 );
not ( \790_b0 , w_40639 );
and ( w_40639 , w_40638 , \790_b1 );
or ( \797_b1 , \792_b1 , w_40642 );
or ( \797_b0 , \792_b0 , w_40641 );
not ( w_40641 , w_40643 );
and ( w_40643 , w_40642 , w_40640 );
or ( w_40640 , \795_b1 , w_40644 );
or ( w_40641 , \795_b0 , \796_b0 );
not ( \796_b0 , w_40645 );
and ( w_40645 , w_40644 , \796_b1 );
or ( \805_b1 , \800_b1 , w_40648 );
or ( \805_b0 , \800_b0 , w_40647 );
not ( w_40647 , w_40649 );
and ( w_40649 , w_40648 , w_40646 );
or ( w_40646 , \803_b1 , w_40650 );
or ( w_40647 , \803_b0 , \804_b0 );
not ( \804_b0 , w_40651 );
and ( w_40651 , w_40650 , \804_b1 );
or ( \831_b1 , \824_b1 , w_40654 );
or ( \831_b0 , \824_b0 , w_40653 );
not ( w_40653 , w_40655 );
and ( w_40655 , w_40654 , w_40652 );
or ( w_40652 , \829_b1 , w_40656 );
or ( w_40653 , \829_b0 , \830_b0 );
not ( \830_b0 , w_40657 );
and ( w_40657 , w_40656 , \830_b1 );
or ( \845_b1 , \840_b1 , w_40660 );
or ( \845_b0 , \840_b0 , w_40659 );
not ( w_40659 , w_40661 );
and ( w_40661 , w_40660 , w_40658 );
or ( w_40658 , \843_b1 , w_40662 );
or ( w_40659 , \843_b0 , \844_b0 );
not ( \844_b0 , w_40663 );
and ( w_40663 , w_40662 , \844_b1 );
or ( \862_b1 , \855_b1 , w_40666 );
or ( \862_b0 , \855_b0 , w_40665 );
not ( w_40665 , w_40667 );
and ( w_40667 , w_40666 , w_40664 );
or ( w_40664 , \860_b1 , w_40668 );
or ( w_40665 , \860_b0 , \861_b0 );
not ( \861_b0 , w_40669 );
and ( w_40669 , w_40668 , \861_b1 );
or ( \865_b1 , \846_b1 , w_40672 );
or ( \865_b0 , \846_b0 , w_40671 );
not ( w_40671 , w_40673 );
and ( w_40673 , w_40672 , w_40670 );
or ( w_40670 , \863_b1 , w_40674 );
or ( w_40671 , \863_b0 , \864_b0 );
not ( \864_b0 , w_40675 );
and ( w_40675 , w_40674 , \864_b1 );
or ( \874_b1 , \870_b1 , w_40678 );
or ( \874_b0 , \870_b0 , w_40677 );
not ( w_40677 , w_40679 );
and ( w_40679 , w_40678 , w_40676 );
or ( w_40676 , \872_b1 , w_40680 );
or ( w_40677 , \872_b0 , \873_b0 );
not ( \873_b0 , w_40681 );
and ( w_40681 , w_40680 , \873_b1 );
or ( \880_b1 , \875_b1 , w_40684 );
or ( \880_b0 , \875_b0 , w_40683 );
not ( w_40683 , w_40685 );
and ( w_40685 , w_40684 , w_40682 );
or ( w_40682 , \878_b1 , w_40686 );
or ( w_40683 , \878_b0 , \879_b0 );
not ( \879_b0 , w_40687 );
and ( w_40687 , w_40686 , \879_b1 );
or ( \888_b1 , \883_b1 , w_40690 );
or ( \888_b0 , \883_b0 , w_40689 );
not ( w_40689 , w_40691 );
and ( w_40691 , w_40690 , w_40688 );
or ( w_40688 , \886_b1 , w_40692 );
or ( w_40689 , \886_b0 , \887_b0 );
not ( \887_b0 , w_40693 );
and ( w_40693 , w_40692 , \887_b1 );
or ( \908_b1 , \903_b1 , w_40696 );
or ( \908_b0 , \903_b0 , w_40695 );
not ( w_40695 , w_40697 );
and ( w_40697 , w_40696 , w_40694 );
or ( w_40694 , \906_b1 , w_40698 );
or ( w_40695 , \906_b0 , \907_b0 );
not ( \907_b0 , w_40699 );
and ( w_40699 , w_40698 , \907_b1 );
or ( \927_b1 , \920_b1 , w_40702 );
or ( \927_b0 , \920_b0 , w_40701 );
not ( w_40701 , w_40703 );
and ( w_40703 , w_40702 , w_40700 );
or ( w_40700 , \925_b1 , w_40704 );
or ( w_40701 , \925_b0 , \926_b0 );
not ( \926_b0 , w_40705 );
and ( w_40705 , w_40704 , \926_b1 );
or ( \944_b1 , \937_b1 , w_40708 );
or ( \944_b0 , \937_b0 , w_40707 );
not ( w_40707 , w_40709 );
and ( w_40709 , w_40708 , w_40706 );
or ( w_40706 , \942_b1 , w_40710 );
or ( w_40707 , \942_b0 , \943_b0 );
not ( \943_b0 , w_40711 );
and ( w_40711 , w_40710 , \943_b1 );
or ( \947_b1 , \928_b1 , w_40714 );
or ( \947_b0 , \928_b0 , w_40713 );
not ( w_40713 , w_40715 );
and ( w_40715 , w_40714 , w_40712 );
or ( w_40712 , \945_b1 , w_40716 );
or ( w_40713 , \945_b0 , \946_b0 );
not ( \946_b0 , w_40717 );
and ( w_40717 , w_40716 , \946_b1 );
or ( \957_b1 , \952_b1 , w_40720 );
or ( \957_b0 , \952_b0 , w_40719 );
not ( w_40719 , w_40721 );
and ( w_40721 , w_40720 , w_40718 );
or ( w_40718 , \955_b1 , w_40722 );
or ( w_40719 , \955_b0 , \956_b0 );
not ( \956_b0 , w_40723 );
and ( w_40723 , w_40722 , \956_b1 );
or ( \963_b1 , \958_b1 , w_40726 );
or ( \963_b0 , \958_b0 , w_40725 );
not ( w_40725 , w_40727 );
and ( w_40727 , w_40726 , w_40724 );
or ( w_40724 , \961_b1 , w_40728 );
or ( w_40725 , \961_b0 , \962_b0 );
not ( \962_b0 , w_40729 );
and ( w_40729 , w_40728 , \962_b1 );
or ( \971_b1 , \966_b1 , w_40732 );
or ( \971_b0 , \966_b0 , w_40731 );
not ( w_40731 , w_40733 );
and ( w_40733 , w_40732 , w_40730 );
or ( w_40730 , \969_b1 , w_40734 );
or ( w_40731 , \969_b0 , \970_b0 );
not ( \970_b0 , w_40735 );
and ( w_40735 , w_40734 , \970_b1 );
or ( \997_b1 , \990_b1 , w_40738 );
or ( \997_b0 , \990_b0 , w_40737 );
not ( w_40737 , w_40739 );
and ( w_40739 , w_40738 , w_40736 );
or ( w_40736 , \995_b1 , w_40740 );
or ( w_40737 , \995_b0 , \996_b0 );
not ( \996_b0 , w_40741 );
and ( w_40741 , w_40740 , \996_b1 );
or ( \1013_b1 , \1006_b1 , w_40744 );
or ( \1013_b0 , \1006_b0 , w_40743 );
not ( w_40743 , w_40745 );
and ( w_40745 , w_40744 , w_40742 );
or ( w_40742 , \1011_b1 , w_40746 );
or ( w_40743 , \1011_b0 , \1012_b0 );
not ( \1012_b0 , w_40747 );
and ( w_40747 , w_40746 , \1012_b1 );
or ( \1030_b1 , \1023_b1 , w_40750 );
or ( \1030_b0 , \1023_b0 , w_40749 );
not ( w_40749 , w_40751 );
and ( w_40751 , w_40750 , w_40748 );
or ( w_40748 , \1028_b1 , w_40752 );
or ( w_40749 , \1028_b0 , \1029_b0 );
not ( \1029_b0 , w_40753 );
and ( w_40753 , w_40752 , \1029_b1 );
or ( \1033_b1 , \1014_b1 , w_40756 );
or ( \1033_b0 , \1014_b0 , w_40755 );
not ( w_40755 , w_40757 );
and ( w_40757 , w_40756 , w_40754 );
or ( w_40754 , \1031_b1 , w_40758 );
or ( w_40755 , \1031_b0 , \1032_b0 );
not ( \1032_b0 , w_40759 );
and ( w_40759 , w_40758 , \1032_b1 );
or ( \1044_b1 , \1039_b1 , w_40762 );
or ( \1044_b0 , \1039_b0 , w_40761 );
not ( w_40761 , w_40763 );
and ( w_40763 , w_40762 , w_40760 );
or ( w_40760 , \1042_b1 , w_40764 );
or ( w_40761 , \1042_b0 , \1043_b0 );
not ( \1043_b0 , w_40765 );
and ( w_40765 , w_40764 , \1043_b1 );
or ( \1052_b1 , \1047_b1 , w_40768 );
or ( \1052_b0 , \1047_b0 , w_40767 );
not ( w_40767 , w_40769 );
and ( w_40769 , w_40768 , w_40766 );
or ( w_40766 , \1050_b1 , w_40770 );
or ( w_40767 , \1050_b0 , \1051_b0 );
not ( \1051_b0 , w_40771 );
and ( w_40771 , w_40770 , \1051_b1 );
or ( \1077_b1 , \1070_b1 , w_40774 );
or ( \1077_b0 , \1070_b0 , w_40773 );
not ( w_40773 , w_40775 );
and ( w_40775 , w_40774 , w_40772 );
or ( w_40772 , \1075_b1 , w_40776 );
or ( w_40773 , \1075_b0 , \1076_b0 );
not ( \1076_b0 , w_40777 );
and ( w_40777 , w_40776 , \1076_b1 );
or ( \1093_b1 , \1086_b1 , w_40780 );
or ( \1093_b0 , \1086_b0 , w_40779 );
not ( w_40779 , w_40781 );
and ( w_40781 , w_40780 , w_40778 );
or ( w_40778 , \1091_b1 , w_40782 );
or ( w_40779 , \1091_b0 , \1092_b0 );
not ( \1092_b0 , w_40783 );
and ( w_40783 , w_40782 , \1092_b1 );
or ( \1111_b1 , \1103_b1 , w_40786 );
or ( \1111_b0 , \1103_b0 , w_40785 );
not ( w_40785 , w_40787 );
and ( w_40787 , w_40786 , w_40784 );
or ( w_40784 , \1109_b1 , w_40788 );
or ( w_40785 , \1109_b0 , \1110_b0 );
not ( \1110_b0 , w_40789 );
and ( w_40789 , w_40788 , \1110_b1 );
or ( \1114_b1 , \1094_b1 , w_40792 );
or ( \1114_b0 , \1094_b0 , w_40791 );
not ( w_40791 , w_40793 );
and ( w_40793 , w_40792 , w_40790 );
or ( w_40790 , \1112_b1 , w_40794 );
or ( w_40791 , \1112_b0 , \1113_b0 );
not ( \1113_b0 , w_40795 );
and ( w_40795 , w_40794 , \1113_b1 );
or ( \1123_b1 , \1118_b1 , w_40798 );
or ( \1123_b0 , \1118_b0 , w_40797 );
not ( w_40797 , w_40799 );
and ( w_40799 , w_40798 , w_40796 );
or ( w_40796 , \1121_b1 , w_40800 );
or ( w_40797 , \1121_b0 , \1122_b0 );
not ( \1122_b0 , w_40801 );
and ( w_40801 , w_40800 , \1122_b1 );
or ( \1129_b1 , \1124_b1 , w_40804 );
or ( \1129_b0 , \1124_b0 , w_40803 );
not ( w_40803 , w_40805 );
and ( w_40805 , w_40804 , w_40802 );
or ( w_40802 , \1127_b1 , w_40806 );
or ( w_40803 , \1127_b0 , \1128_b0 );
not ( \1128_b0 , w_40807 );
and ( w_40807 , w_40806 , \1128_b1 );
or ( \1137_b1 , \1132_b1 , w_40810 );
or ( \1137_b0 , \1132_b0 , w_40809 );
not ( w_40809 , w_40811 );
and ( w_40811 , w_40810 , w_40808 );
or ( w_40808 , \1135_b1 , w_40812 );
or ( w_40809 , \1135_b0 , \1136_b0 );
not ( \1136_b0 , w_40813 );
and ( w_40813 , w_40812 , \1136_b1 );
or ( \1153_b1 , \1146_b1 , w_40816 );
or ( \1153_b0 , \1146_b0 , w_40815 );
not ( w_40815 , w_40817 );
and ( w_40817 , w_40816 , w_40814 );
or ( w_40814 , \1151_b1 , w_40818 );
or ( w_40815 , \1151_b0 , \1152_b0 );
not ( \1152_b0 , w_40819 );
and ( w_40819 , w_40818 , \1152_b1 );
or ( \1169_b1 , \1162_b1 , w_40822 );
or ( \1169_b0 , \1162_b0 , w_40821 );
not ( w_40821 , w_40823 );
and ( w_40823 , w_40822 , w_40820 );
or ( w_40820 , \1167_b1 , w_40824 );
or ( w_40821 , \1167_b0 , \1168_b0 );
not ( \1168_b0 , w_40825 );
and ( w_40825 , w_40824 , \1168_b1 );
or ( \1190_b1 , \1183_b1 , w_40828 );
or ( \1190_b0 , \1183_b0 , w_40827 );
not ( w_40827 , w_40829 );
and ( w_40829 , w_40828 , w_40826 );
or ( w_40826 , \1188_b1 , w_40830 );
or ( w_40827 , \1188_b0 , \1189_b0 );
not ( \1189_b0 , w_40831 );
and ( w_40831 , w_40830 , \1189_b1 );
or ( \1193_b1 , \1170_b1 , w_40834 );
or ( \1193_b0 , \1170_b0 , w_40833 );
not ( w_40833 , w_40835 );
and ( w_40835 , w_40834 , w_40832 );
or ( w_40832 , \1191_b1 , w_40836 );
or ( w_40833 , \1191_b0 , \1192_b0 );
not ( \1192_b0 , w_40837 );
and ( w_40837 , w_40836 , \1192_b1 );
or ( \1207_b1 , \1199_b1 , w_40840 );
or ( \1207_b0 , \1199_b0 , w_40839 );
not ( w_40839 , w_40841 );
and ( w_40841 , w_40840 , w_40838 );
or ( w_40838 , \1205_b1 , w_40842 );
or ( w_40839 , \1205_b0 , \1206_b0 );
not ( \1206_b0 , w_40843 );
and ( w_40843 , w_40842 , \1206_b1 );
or ( \1217_b1 , \1212_b1 , w_40846 );
or ( \1217_b0 , \1212_b0 , w_40845 );
not ( w_40845 , w_40847 );
and ( w_40847 , w_40846 , w_40844 );
or ( w_40844 , \1215_b1 , w_40848 );
or ( w_40845 , \1215_b0 , \1216_b0 );
not ( \1216_b0 , w_40849 );
and ( w_40849 , w_40848 , \1216_b1 );
or ( \1222_b1 , \1218_b1 , w_40852 );
or ( \1222_b0 , \1218_b0 , w_40851 );
not ( w_40851 , w_40853 );
and ( w_40853 , w_40852 , w_40850 );
or ( w_40850 , \1220_b1 , w_40854 );
or ( w_40851 , \1220_b0 , \1221_b0 );
not ( \1221_b0 , w_40855 );
and ( w_40855 , w_40854 , \1221_b1 );
or ( \1233_b1 , \1228_b1 , w_40858 );
or ( \1233_b0 , \1228_b0 , w_40857 );
not ( w_40857 , w_40859 );
and ( w_40859 , w_40858 , w_40856 );
or ( w_40856 , \1231_b1 , w_40860 );
or ( w_40857 , \1231_b0 , \1232_b0 );
not ( \1232_b0 , w_40861 );
and ( w_40861 , w_40860 , \1232_b1 );
or ( \1239_b1 , \1234_b1 , w_40864 );
or ( \1239_b0 , \1234_b0 , w_40863 );
not ( w_40863 , w_40865 );
and ( w_40865 , w_40864 , w_40862 );
or ( w_40862 , \1237_b1 , w_40866 );
or ( w_40863 , \1237_b0 , \1238_b0 );
not ( \1238_b0 , w_40867 );
and ( w_40867 , w_40866 , \1238_b1 );
or ( \1259_b1 , \1252_b1 , w_40870 );
or ( \1259_b0 , \1252_b0 , w_40869 );
not ( w_40869 , w_40871 );
and ( w_40871 , w_40870 , w_40868 );
or ( w_40868 , \1257_b1 , w_40872 );
or ( w_40869 , \1257_b0 , \1258_b0 );
not ( \1258_b0 , w_40873 );
and ( w_40873 , w_40872 , \1258_b1 );
or ( \1275_b1 , \1268_b1 , w_40876 );
or ( \1275_b0 , \1268_b0 , w_40875 );
not ( w_40875 , w_40877 );
and ( w_40877 , w_40876 , w_40874 );
or ( w_40874 , \1273_b1 , w_40878 );
or ( w_40875 , \1273_b0 , \1274_b0 );
not ( \1274_b0 , w_40879 );
and ( w_40879 , w_40878 , \1274_b1 );
or ( \1295_b1 , \1288_b1 , w_40882 );
or ( \1295_b0 , \1288_b0 , w_40881 );
not ( w_40881 , w_40883 );
and ( w_40883 , w_40882 , w_40880 );
or ( w_40880 , \1293_b1 , w_40884 );
or ( w_40881 , \1293_b0 , \1294_b0 );
not ( \1294_b0 , w_40885 );
and ( w_40885 , w_40884 , \1294_b1 );
or ( \1298_b1 , \1276_b1 , w_40888 );
or ( \1298_b0 , \1276_b0 , w_40887 );
not ( w_40887 , w_40889 );
and ( w_40889 , w_40888 , w_40886 );
or ( w_40886 , \1296_b1 , w_40890 );
or ( w_40887 , \1296_b0 , \1297_b0 );
not ( \1297_b0 , w_40891 );
and ( w_40891 , w_40890 , \1297_b1 );
or ( \1315_b1 , \1311_b1 , w_40894 );
or ( \1315_b0 , \1311_b0 , w_40893 );
not ( w_40893 , w_40895 );
and ( w_40895 , w_40894 , w_40892 );
or ( w_40892 , \1313_b1 , w_40896 );
or ( w_40893 , \1313_b0 , \1314_b0 );
not ( \1314_b0 , w_40897 );
and ( w_40897 , w_40896 , \1314_b1 );
or ( \1326_b1 , \1321_b1 , w_40900 );
or ( \1326_b0 , \1321_b0 , w_40899 );
not ( w_40899 , w_40901 );
and ( w_40901 , w_40900 , w_40898 );
or ( w_40898 , \1324_b1 , w_40902 );
or ( w_40899 , \1324_b0 , \1325_b0 );
not ( \1325_b0 , w_40903 );
and ( w_40903 , w_40902 , \1325_b1 );
or ( \1329_b1 , \1316_b1 , w_40906 );
or ( \1329_b0 , \1316_b0 , w_40905 );
not ( w_40905 , w_40907 );
and ( w_40907 , w_40906 , w_40904 );
or ( w_40904 , \1327_b1 , w_40908 );
or ( w_40905 , \1327_b0 , \1328_b0 );
not ( \1328_b0 , w_40909 );
and ( w_40909 , w_40908 , \1328_b1 );
or ( \1337_b1 , \1333_b1 , w_40912 );
or ( \1337_b0 , \1333_b0 , w_40911 );
not ( w_40911 , w_40913 );
and ( w_40913 , w_40912 , w_40910 );
or ( w_40910 , \1335_b1 , w_40914 );
or ( w_40911 , \1335_b0 , \1336_b0 );
not ( \1336_b0 , w_40915 );
and ( w_40915 , w_40914 , \1336_b1 );
or ( \1343_b1 , \1338_b1 , w_40918 );
or ( \1343_b0 , \1338_b0 , w_40917 );
not ( w_40917 , w_40919 );
and ( w_40919 , w_40918 , w_40916 );
or ( w_40916 , \1341_b1 , w_40920 );
or ( w_40917 , \1341_b0 , \1342_b0 );
not ( \1342_b0 , w_40921 );
and ( w_40921 , w_40920 , \1342_b1 );
or ( \1350_b1 , \1346_b1 , w_40924 );
or ( \1350_b0 , \1346_b0 , w_40923 );
not ( w_40923 , w_40925 );
and ( w_40925 , w_40924 , w_40922 );
or ( w_40922 , \1348_b1 , w_40926 );
or ( w_40923 , \1348_b0 , \1349_b0 );
not ( \1349_b0 , w_40927 );
and ( w_40927 , w_40926 , \1349_b1 );
or ( \1376_b1 , \1369_b1 , w_40930 );
or ( \1376_b0 , \1369_b0 , w_40929 );
not ( w_40929 , w_40931 );
and ( w_40931 , w_40930 , w_40928 );
or ( w_40928 , \1374_b1 , w_40932 );
or ( w_40929 , \1374_b0 , \1375_b0 );
not ( \1375_b0 , w_40933 );
and ( w_40933 , w_40932 , \1375_b1 );
or ( \1392_b1 , \1385_b1 , w_40936 );
or ( \1392_b0 , \1385_b0 , w_40935 );
not ( w_40935 , w_40937 );
and ( w_40937 , w_40936 , w_40934 );
or ( w_40934 , \1390_b1 , w_40938 );
or ( w_40935 , \1390_b0 , \1391_b0 );
not ( \1391_b0 , w_40939 );
and ( w_40939 , w_40938 , \1391_b1 );
or ( \1409_b1 , \1402_b1 , w_40942 );
or ( \1409_b0 , \1402_b0 , w_40941 );
not ( w_40941 , w_40943 );
and ( w_40943 , w_40942 , w_40940 );
or ( w_40940 , \1407_b1 , w_40944 );
or ( w_40941 , \1407_b0 , \1408_b0 );
not ( \1408_b0 , w_40945 );
and ( w_40945 , w_40944 , \1408_b1 );
or ( \1412_b1 , \1393_b1 , w_40948 );
or ( \1412_b0 , \1393_b0 , w_40947 );
not ( w_40947 , w_40949 );
and ( w_40949 , w_40948 , w_40946 );
or ( w_40946 , \1410_b1 , w_40950 );
or ( w_40947 , \1410_b0 , \1411_b0 );
not ( \1411_b0 , w_40951 );
and ( w_40951 , w_40950 , \1411_b1 );
or ( \1426_b1 , \1421_b1 , w_40954 );
or ( \1426_b0 , \1421_b0 , w_40953 );
not ( w_40953 , w_40955 );
and ( w_40955 , w_40954 , w_40952 );
or ( w_40952 , \1424_b1 , w_40956 );
or ( w_40953 , \1424_b0 , \1425_b0 );
not ( \1425_b0 , w_40957 );
and ( w_40957 , w_40956 , \1425_b1 );
or ( \1433_b1 , \1429_b1 , w_40960 );
or ( \1433_b0 , \1429_b0 , w_40959 );
not ( w_40959 , w_40961 );
and ( w_40961 , w_40960 , w_40958 );
or ( w_40958 , \1431_b1 , w_40962 );
or ( w_40959 , \1431_b0 , \1432_b0 );
not ( \1432_b0 , w_40963 );
and ( w_40963 , w_40962 , \1432_b1 );
or ( \1442_b1 , \1434_b1 , w_40966 );
or ( \1442_b0 , \1434_b0 , w_40965 );
not ( w_40965 , w_40967 );
and ( w_40967 , w_40966 , w_40964 );
or ( w_40964 , \1440_b1 , w_40968 );
or ( w_40965 , \1440_b0 , \1441_b0 );
not ( \1441_b0 , w_40969 );
and ( w_40969 , w_40968 , \1441_b1 );
or ( \1452_b1 , \1447_b1 , w_40972 );
or ( \1452_b0 , \1447_b0 , w_40971 );
not ( w_40971 , w_40973 );
and ( w_40973 , w_40972 , w_40970 );
or ( w_40970 , \1450_b1 , w_40974 );
or ( w_40971 , \1450_b0 , \1451_b0 );
not ( \1451_b0 , w_40975 );
and ( w_40975 , w_40974 , \1451_b1 );
or ( \1458_b1 , \1453_b1 , w_40978 );
or ( \1458_b0 , \1453_b0 , w_40977 );
not ( w_40977 , w_40979 );
and ( w_40979 , w_40978 , w_40976 );
or ( w_40976 , \1456_b1 , w_40980 );
or ( w_40977 , \1456_b0 , \1457_b0 );
not ( \1457_b0 , w_40981 );
and ( w_40981 , w_40980 , \1457_b1 );
or ( \1466_b1 , \1461_b1 , w_40984 );
or ( \1466_b0 , \1461_b0 , w_40983 );
not ( w_40983 , w_40985 );
and ( w_40985 , w_40984 , w_40982 );
or ( w_40982 , \1464_b1 , w_40986 );
or ( w_40983 , \1464_b0 , \1465_b0 );
not ( \1465_b0 , w_40987 );
and ( w_40987 , w_40986 , \1465_b1 );
or ( \1491_b1 , \1484_b1 , w_40990 );
or ( \1491_b0 , \1484_b0 , w_40989 );
not ( w_40989 , w_40991 );
and ( w_40991 , w_40990 , w_40988 );
or ( w_40988 , \1489_b1 , w_40992 );
or ( w_40989 , \1489_b0 , \1490_b0 );
not ( \1490_b0 , w_40993 );
and ( w_40993 , w_40992 , \1490_b1 );
or ( \1507_b1 , \1500_b1 , w_40996 );
or ( \1507_b0 , \1500_b0 , w_40995 );
not ( w_40995 , w_40997 );
and ( w_40997 , w_40996 , w_40994 );
or ( w_40994 , \1505_b1 , w_40998 );
or ( w_40995 , \1505_b0 , \1506_b0 );
not ( \1506_b0 , w_40999 );
and ( w_40999 , w_40998 , \1506_b1 );
or ( \1524_b1 , \1517_b1 , w_41002 );
or ( \1524_b0 , \1517_b0 , w_41001 );
not ( w_41001 , w_41003 );
and ( w_41003 , w_41002 , w_41000 );
or ( w_41000 , \1522_b1 , w_41004 );
or ( w_41001 , \1522_b0 , \1523_b0 );
not ( \1523_b0 , w_41005 );
and ( w_41005 , w_41004 , \1523_b1 );
or ( \1527_b1 , \1508_b1 , w_41008 );
or ( \1527_b0 , \1508_b0 , w_41007 );
not ( w_41007 , w_41009 );
and ( w_41009 , w_41008 , w_41006 );
or ( w_41006 , \1525_b1 , w_41010 );
or ( w_41007 , \1525_b0 , \1526_b0 );
not ( \1526_b0 , w_41011 );
and ( w_41011 , w_41010 , \1526_b1 );
or ( \1541_b1 , \1536_b1 , w_41014 );
or ( \1541_b0 , \1536_b0 , w_41013 );
not ( w_41013 , w_41015 );
and ( w_41015 , w_41014 , w_41012 );
or ( w_41012 , \1539_b1 , w_41016 );
or ( w_41013 , \1539_b0 , \1540_b0 );
not ( \1540_b0 , w_41017 );
and ( w_41017 , w_41016 , \1540_b1 );
or ( \1549_b1 , \1544_b1 , w_41020 );
or ( \1549_b0 , \1544_b0 , w_41019 );
not ( w_41019 , w_41021 );
and ( w_41021 , w_41020 , w_41018 );
or ( w_41018 , \1547_b1 , w_41022 );
or ( w_41019 , \1547_b0 , \1548_b0 );
not ( \1548_b0 , w_41023 );
and ( w_41023 , w_41022 , \1548_b1 );
or ( \1558_b1 , \1550_b1 , w_41026 );
or ( \1558_b0 , \1550_b0 , w_41025 );
not ( w_41025 , w_41027 );
and ( w_41027 , w_41026 , w_41024 );
or ( w_41024 , \1556_b1 , w_41028 );
or ( w_41025 , \1556_b0 , \1557_b0 );
not ( \1557_b0 , w_41029 );
and ( w_41029 , w_41028 , \1557_b1 );
or ( \1567_b1 , \1563_b1 , w_41032 );
or ( \1567_b0 , \1563_b0 , w_41031 );
not ( w_41031 , w_41033 );
and ( w_41033 , w_41032 , w_41030 );
or ( w_41030 , \1565_b1 , w_41034 );
or ( w_41031 , \1565_b0 , \1566_b0 );
not ( \1566_b0 , w_41035 );
and ( w_41035 , w_41034 , \1566_b1 );
or ( \1573_b1 , \1568_b1 , w_41038 );
or ( \1573_b0 , \1568_b0 , w_41037 );
not ( w_41037 , w_41039 );
and ( w_41039 , w_41038 , w_41036 );
or ( w_41036 , \1571_b1 , w_41040 );
or ( w_41037 , \1571_b0 , \1572_b0 );
not ( \1572_b0 , w_41041 );
and ( w_41041 , w_41040 , \1572_b1 );
or ( \1581_b1 , \1576_b1 , w_41044 );
or ( \1581_b0 , \1576_b0 , w_41043 );
not ( w_41043 , w_41045 );
and ( w_41045 , w_41044 , w_41042 );
or ( w_41042 , \1579_b1 , w_41046 );
or ( w_41043 , \1579_b0 , \1580_b0 );
not ( \1580_b0 , w_41047 );
and ( w_41047 , w_41046 , \1580_b1 );
or ( \1603_b1 , \1596_b1 , w_41050 );
or ( \1603_b0 , \1596_b0 , w_41049 );
not ( w_41049 , w_41051 );
and ( w_41051 , w_41050 , w_41048 );
or ( w_41048 , \1601_b1 , w_41052 );
or ( w_41049 , \1601_b0 , \1602_b0 );
not ( \1602_b0 , w_41053 );
and ( w_41053 , w_41052 , \1602_b1 );
or ( \1623_b1 , \1616_b1 , w_41056 );
or ( \1623_b0 , \1616_b0 , w_41055 );
not ( w_41055 , w_41057 );
and ( w_41057 , w_41056 , w_41054 );
or ( w_41054 , \1621_b1 , w_41058 );
or ( w_41055 , \1621_b0 , \1622_b0 );
not ( \1622_b0 , w_41059 );
and ( w_41059 , w_41058 , \1622_b1 );
or ( \1640_b1 , \1633_b1 , w_41062 );
or ( \1640_b0 , \1633_b0 , w_41061 );
not ( w_41061 , w_41063 );
and ( w_41063 , w_41062 , w_41060 );
or ( w_41060 , \1638_b1 , w_41064 );
or ( w_41061 , \1638_b0 , \1639_b0 );
not ( \1639_b0 , w_41065 );
and ( w_41065 , w_41064 , \1639_b1 );
or ( \1643_b1 , \1624_b1 , w_41068 );
or ( \1643_b0 , \1624_b0 , w_41067 );
not ( w_41067 , w_41069 );
and ( w_41069 , w_41068 , w_41066 );
or ( w_41066 , \1641_b1 , w_41070 );
or ( w_41067 , \1641_b0 , \1642_b0 );
not ( \1642_b0 , w_41071 );
and ( w_41071 , w_41070 , \1642_b1 );
or ( \1653_b1 , \1648_b1 , w_41074 );
or ( \1653_b0 , \1648_b0 , w_41073 );
not ( w_41073 , w_41075 );
and ( w_41075 , w_41074 , w_41072 );
or ( w_41072 , \1651_b1 , w_41076 );
or ( w_41073 , \1651_b0 , \1652_b0 );
not ( \1652_b0 , w_41077 );
and ( w_41077 , w_41076 , \1652_b1 );
or ( \1670_b1 , \1663_b1 , w_41080 );
or ( \1670_b0 , \1663_b0 , w_41079 );
not ( w_41079 , w_41081 );
and ( w_41081 , w_41080 , w_41078 );
or ( w_41078 , \1668_b1 , w_41082 );
or ( w_41079 , \1668_b0 , \1669_b0 );
not ( \1669_b0 , w_41083 );
and ( w_41083 , w_41082 , \1669_b1 );
or ( \1676_b1 , \1654_b1 , w_41086 );
or ( \1676_b0 , \1654_b0 , w_41085 );
not ( w_41085 , w_41087 );
and ( w_41087 , w_41086 , w_41084 );
or ( w_41084 , \1674_b1 , w_41088 );
or ( w_41085 , \1674_b0 , \1675_b0 );
not ( \1675_b0 , w_41089 );
and ( w_41089 , w_41088 , \1675_b1 );
or ( \1685_b1 , \1681_b1 , w_41092 );
or ( \1685_b0 , \1681_b0 , w_41091 );
not ( w_41091 , w_41093 );
and ( w_41093 , w_41092 , w_41090 );
or ( w_41090 , \1683_b1 , w_41094 );
or ( w_41091 , \1683_b0 , \1684_b0 );
not ( \1684_b0 , w_41095 );
and ( w_41095 , w_41094 , \1684_b1 );
or ( \1691_b1 , \1686_b1 , w_41098 );
or ( \1691_b0 , \1686_b0 , w_41097 );
not ( w_41097 , w_41099 );
and ( w_41099 , w_41098 , w_41096 );
or ( w_41096 , \1689_b1 , w_41100 );
or ( w_41097 , \1689_b0 , \1690_b0 );
not ( \1690_b0 , w_41101 );
and ( w_41101 , w_41100 , \1690_b1 );
or ( \1699_b1 , \1694_b1 , w_41104 );
or ( \1699_b0 , \1694_b0 , w_41103 );
not ( w_41103 , w_41105 );
and ( w_41105 , w_41104 , w_41102 );
or ( w_41102 , \1697_b1 , w_41106 );
or ( w_41103 , \1697_b0 , \1698_b0 );
not ( \1698_b0 , w_41107 );
and ( w_41107 , w_41106 , \1698_b1 );
or ( \1721_b1 , \1714_b1 , w_41110 );
or ( \1721_b0 , \1714_b0 , w_41109 );
not ( w_41109 , w_41111 );
and ( w_41111 , w_41110 , w_41108 );
or ( w_41108 , \1719_b1 , w_41112 );
or ( w_41109 , \1719_b0 , \1720_b0 );
not ( \1720_b0 , w_41113 );
and ( w_41113 , w_41112 , \1720_b1 );
or ( \1737_b1 , \1730_b1 , w_41116 );
or ( \1737_b0 , \1730_b0 , w_41115 );
not ( w_41115 , w_41117 );
and ( w_41117 , w_41116 , w_41114 );
or ( w_41114 , \1735_b1 , w_41118 );
or ( w_41115 , \1735_b0 , \1736_b0 );
not ( \1736_b0 , w_41119 );
and ( w_41119 , w_41118 , \1736_b1 );
or ( \1757_b1 , \1750_b1 , w_41122 );
or ( \1757_b0 , \1750_b0 , w_41121 );
not ( w_41121 , w_41123 );
and ( w_41123 , w_41122 , w_41120 );
or ( w_41120 , \1755_b1 , w_41124 );
or ( w_41121 , \1755_b0 , \1756_b0 );
not ( \1756_b0 , w_41125 );
and ( w_41125 , w_41124 , \1756_b1 );
or ( \1760_b1 , \1738_b1 , w_41128 );
or ( \1760_b0 , \1738_b0 , w_41127 );
not ( w_41127 , w_41129 );
and ( w_41129 , w_41128 , w_41126 );
or ( w_41126 , \1758_b1 , w_41130 );
or ( w_41127 , \1758_b0 , \1759_b0 );
not ( \1759_b0 , w_41131 );
and ( w_41131 , w_41130 , \1759_b1 );
or ( \1777_b1 , \1769_b1 , w_41134 );
or ( \1777_b0 , \1769_b0 , w_41133 );
not ( w_41133 , w_41135 );
and ( w_41135 , w_41134 , w_41132 );
or ( w_41132 , \1775_b1 , w_41136 );
or ( w_41133 , \1775_b0 , \1776_b0 );
not ( \1776_b0 , w_41137 );
and ( w_41137 , w_41136 , \1776_b1 );
or ( \1785_b1 , \1781_b1 , w_41140 );
or ( \1785_b0 , \1781_b0 , w_41139 );
not ( w_41139 , w_41141 );
and ( w_41141 , w_41140 , w_41138 );
or ( w_41138 , \1783_b1 , w_41142 );
or ( w_41139 , \1783_b0 , \1784_b0 );
not ( \1784_b0 , w_41143 );
and ( w_41143 , w_41142 , \1784_b1 );
or ( \1796_b1 , \1791_b1 , w_41146 );
or ( \1796_b0 , \1791_b0 , w_41145 );
not ( w_41145 , w_41147 );
and ( w_41147 , w_41146 , w_41144 );
or ( w_41144 , \1794_b1 , w_41148 );
or ( w_41145 , \1794_b0 , \1795_b0 );
not ( \1795_b0 , w_41149 );
and ( w_41149 , w_41148 , \1795_b1 );
or ( \1799_b1 , \1786_b1 , w_41152 );
or ( \1799_b0 , \1786_b0 , w_41151 );
not ( w_41151 , w_41153 );
and ( w_41153 , w_41152 , w_41150 );
or ( w_41150 , \1797_b1 , w_41154 );
or ( w_41151 , \1797_b0 , \1798_b0 );
not ( \1798_b0 , w_41155 );
and ( w_41155 , w_41154 , \1798_b1 );
or ( \1808_b1 , \1804_b1 , w_41158 );
or ( \1808_b0 , \1804_b0 , w_41157 );
not ( w_41157 , w_41159 );
and ( w_41159 , w_41158 , w_41156 );
or ( w_41156 , \1806_b1 , w_41160 );
or ( w_41157 , \1806_b0 , \1807_b0 );
not ( \1807_b0 , w_41161 );
and ( w_41161 , w_41160 , \1807_b1 );
or ( \1814_b1 , \1809_b1 , w_41164 );
or ( \1814_b0 , \1809_b0 , w_41163 );
not ( w_41163 , w_41165 );
and ( w_41165 , w_41164 , w_41162 );
or ( w_41162 , \1812_b1 , w_41166 );
or ( w_41163 , \1812_b0 , \1813_b0 );
not ( \1813_b0 , w_41167 );
and ( w_41167 , w_41166 , \1813_b1 );
or ( \1822_b1 , \1817_b1 , w_41170 );
or ( \1822_b0 , \1817_b0 , w_41169 );
not ( w_41169 , w_41171 );
and ( w_41171 , w_41170 , w_41168 );
or ( w_41168 , \1820_b1 , w_41172 );
or ( w_41169 , \1820_b0 , \1821_b0 );
not ( \1821_b0 , w_41173 );
and ( w_41173 , w_41172 , \1821_b1 );
or ( \1848_b1 , \1841_b1 , w_41176 );
or ( \1848_b0 , \1841_b0 , w_41175 );
not ( w_41175 , w_41177 );
and ( w_41177 , w_41176 , w_41174 );
or ( w_41174 , \1846_b1 , w_41178 );
or ( w_41175 , \1846_b0 , \1847_b0 );
not ( \1847_b0 , w_41179 );
and ( w_41179 , w_41178 , \1847_b1 );
or ( \1864_b1 , \1857_b1 , w_41182 );
or ( \1864_b0 , \1857_b0 , w_41181 );
not ( w_41181 , w_41183 );
and ( w_41183 , w_41182 , w_41180 );
or ( w_41180 , \1862_b1 , w_41184 );
or ( w_41181 , \1862_b0 , \1863_b0 );
not ( \1863_b0 , w_41185 );
and ( w_41185 , w_41184 , \1863_b1 );
or ( \1881_b1 , \1874_b1 , w_41188 );
or ( \1881_b0 , \1874_b0 , w_41187 );
not ( w_41187 , w_41189 );
and ( w_41189 , w_41188 , w_41186 );
or ( w_41186 , \1879_b1 , w_41190 );
or ( w_41187 , \1879_b0 , \1880_b0 );
not ( \1880_b0 , w_41191 );
and ( w_41191 , w_41190 , \1880_b1 );
or ( \1884_b1 , \1865_b1 , w_41194 );
or ( \1884_b0 , \1865_b0 , w_41193 );
not ( w_41193 , w_41195 );
and ( w_41195 , w_41194 , w_41192 );
or ( w_41192 , \1882_b1 , w_41196 );
or ( w_41193 , \1882_b0 , \1883_b0 );
not ( \1883_b0 , w_41197 );
and ( w_41197 , w_41196 , \1883_b1 );
or ( \1894_b1 , \1889_b1 , w_41200 );
or ( \1894_b0 , \1889_b0 , w_41199 );
not ( w_41199 , w_41201 );
and ( w_41201 , w_41200 , w_41198 );
or ( w_41198 , \1892_b1 , w_41202 );
or ( w_41199 , \1892_b0 , \1893_b0 );
not ( \1893_b0 , w_41203 );
and ( w_41203 , w_41202 , \1893_b1 );
or ( \1911_b1 , \1904_b1 , w_41206 );
or ( \1911_b0 , \1904_b0 , w_41205 );
not ( w_41205 , w_41207 );
and ( w_41207 , w_41206 , w_41204 );
or ( w_41204 , \1909_b1 , w_41208 );
or ( w_41205 , \1909_b0 , \1910_b0 );
not ( \1910_b0 , w_41209 );
and ( w_41209 , w_41208 , \1910_b1 );
or ( \1918_b1 , \1914_b1 , w_41212 );
or ( \1918_b0 , \1914_b0 , w_41211 );
not ( w_41211 , w_41213 );
and ( w_41213 , w_41212 , w_41210 );
or ( w_41210 , \1916_b1 , w_41214 );
or ( w_41211 , \1916_b0 , \1917_b0 );
not ( \1917_b0 , w_41215 );
and ( w_41215 , w_41214 , \1917_b1 );
or ( \1921_b1 , \1895_b1 , w_41218 );
or ( \1921_b0 , \1895_b0 , w_41217 );
not ( w_41217 , w_41219 );
and ( w_41219 , w_41218 , w_41216 );
or ( w_41216 , \1919_b1 , w_41220 );
or ( w_41217 , \1919_b0 , \1920_b0 );
not ( \1920_b0 , w_41221 );
and ( w_41221 , w_41220 , \1920_b1 );
or ( \1931_b1 , \1926_b1 , w_41224 );
or ( \1931_b0 , \1926_b0 , w_41223 );
not ( w_41223 , w_41225 );
and ( w_41225 , w_41224 , w_41222 );
or ( w_41222 , \1929_b1 , w_41226 );
or ( w_41223 , \1929_b0 , \1930_b0 );
not ( \1930_b0 , w_41227 );
and ( w_41227 , w_41226 , \1930_b1 );
or ( \1937_b1 , \1932_b1 , w_41230 );
or ( \1937_b0 , \1932_b0 , w_41229 );
not ( w_41229 , w_41231 );
and ( w_41231 , w_41230 , w_41228 );
or ( w_41228 , \1935_b1 , w_41232 );
or ( w_41229 , \1935_b0 , \1936_b0 );
not ( \1936_b0 , w_41233 );
and ( w_41233 , w_41232 , \1936_b1 );
or ( \1945_b1 , \1940_b1 , w_41236 );
or ( \1945_b0 , \1940_b0 , w_41235 );
not ( w_41235 , w_41237 );
and ( w_41237 , w_41236 , w_41234 );
or ( w_41234 , \1943_b1 , w_41238 );
or ( w_41235 , \1943_b0 , \1944_b0 );
not ( \1944_b0 , w_41239 );
and ( w_41239 , w_41238 , \1944_b1 );
or ( \1970_b1 , \1963_b1 , w_41242 );
or ( \1970_b0 , \1963_b0 , w_41241 );
not ( w_41241 , w_41243 );
and ( w_41243 , w_41242 , w_41240 );
or ( w_41240 , \1968_b1 , w_41244 );
or ( w_41241 , \1968_b0 , \1969_b0 );
not ( \1969_b0 , w_41245 );
and ( w_41245 , w_41244 , \1969_b1 );
or ( \1986_b1 , \1979_b1 , w_41248 );
or ( \1986_b0 , \1979_b0 , w_41247 );
not ( w_41247 , w_41249 );
and ( w_41249 , w_41248 , w_41246 );
or ( w_41246 , \1984_b1 , w_41250 );
or ( w_41247 , \1984_b0 , \1985_b0 );
not ( \1985_b0 , w_41251 );
and ( w_41251 , w_41250 , \1985_b1 );
or ( \2003_b1 , \1996_b1 , w_41254 );
or ( \2003_b0 , \1996_b0 , w_41253 );
not ( w_41253 , w_41255 );
and ( w_41255 , w_41254 , w_41252 );
or ( w_41252 , \2001_b1 , w_41256 );
or ( w_41253 , \2001_b0 , \2002_b0 );
not ( \2002_b0 , w_41257 );
and ( w_41257 , w_41256 , \2002_b1 );
or ( \2006_b1 , \1987_b1 , w_41260 );
or ( \2006_b0 , \1987_b0 , w_41259 );
not ( w_41259 , w_41261 );
and ( w_41261 , w_41260 , w_41258 );
or ( w_41258 , \2004_b1 , w_41262 );
or ( w_41259 , \2004_b0 , \2005_b0 );
not ( \2005_b0 , w_41263 );
and ( w_41263 , w_41262 , \2005_b1 );
or ( \2022_b1 , \2015_b1 , w_41266 );
or ( \2022_b0 , \2015_b0 , w_41265 );
not ( w_41265 , w_41267 );
and ( w_41267 , w_41266 , w_41264 );
or ( w_41264 , \2020_b1 , w_41268 );
or ( w_41265 , \2020_b0 , \2021_b0 );
not ( \2021_b0 , w_41269 );
and ( w_41269 , w_41268 , \2021_b1 );
or ( \2038_b1 , \2031_b1 , w_41272 );
or ( \2038_b0 , \2031_b0 , w_41271 );
not ( w_41271 , w_41273 );
and ( w_41273 , w_41272 , w_41270 );
or ( w_41270 , \2036_b1 , w_41274 );
or ( w_41271 , \2036_b0 , \2037_b0 );
not ( \2037_b0 , w_41275 );
and ( w_41275 , w_41274 , \2037_b1 );
or ( \2048_b1 , \2043_b1 , w_41278 );
or ( \2048_b0 , \2043_b0 , w_41277 );
not ( w_41277 , w_41279 );
and ( w_41279 , w_41278 , w_41276 );
or ( w_41276 , \2046_b1 , w_41280 );
or ( w_41277 , \2046_b0 , \2047_b0 );
not ( \2047_b0 , w_41281 );
and ( w_41281 , w_41280 , \2047_b1 );
or ( \2051_b1 , \2039_b1 , w_41284 );
or ( \2051_b0 , \2039_b0 , w_41283 );
not ( w_41283 , w_41285 );
and ( w_41285 , w_41284 , w_41282 );
or ( w_41282 , \2049_b1 , w_41286 );
or ( w_41283 , \2049_b0 , \2050_b0 );
not ( \2050_b0 , w_41287 );
and ( w_41287 , w_41286 , \2050_b1 );
or ( \2061_b1 , \2056_b1 , w_41290 );
or ( \2061_b0 , \2056_b0 , w_41289 );
not ( w_41289 , w_41291 );
and ( w_41291 , w_41290 , w_41288 );
or ( w_41288 , \2059_b1 , w_41292 );
or ( w_41289 , \2059_b0 , \2060_b0 );
not ( \2060_b0 , w_41293 );
and ( w_41293 , w_41292 , \2060_b1 );
or ( \2067_b1 , \2062_b1 , w_41296 );
or ( \2067_b0 , \2062_b0 , w_41295 );
not ( w_41295 , w_41297 );
and ( w_41297 , w_41296 , w_41294 );
or ( w_41294 , \2065_b1 , w_41298 );
or ( w_41295 , \2065_b0 , \2066_b0 );
not ( \2066_b0 , w_41299 );
and ( w_41299 , w_41298 , \2066_b1 );
or ( \2078_b1 , \2073_b1 , w_41302 );
or ( \2078_b0 , \2073_b0 , w_41301 );
not ( w_41301 , w_41303 );
and ( w_41303 , w_41302 , w_41300 );
or ( w_41300 , \2076_b1 , w_41304 );
or ( w_41301 , \2076_b0 , \2077_b0 );
not ( \2077_b0 , w_41305 );
and ( w_41305 , w_41304 , \2077_b1 );
or ( \2100_b1 , \2093_b1 , w_41308 );
or ( \2100_b0 , \2093_b0 , w_41307 );
not ( w_41307 , w_41309 );
and ( w_41309 , w_41308 , w_41306 );
or ( w_41306 , \2098_b1 , w_41310 );
or ( w_41307 , \2098_b0 , \2099_b0 );
not ( \2099_b0 , w_41311 );
and ( w_41311 , w_41310 , \2099_b1 );
or ( \2116_b1 , \2109_b1 , w_41314 );
or ( \2116_b0 , \2109_b0 , w_41313 );
not ( w_41313 , w_41315 );
and ( w_41315 , w_41314 , w_41312 );
or ( w_41312 , \2114_b1 , w_41316 );
or ( w_41313 , \2114_b0 , \2115_b0 );
not ( \2115_b0 , w_41317 );
and ( w_41317 , w_41316 , \2115_b1 );
or ( \2137_b1 , \2130_b1 , w_41320 );
or ( \2137_b0 , \2130_b0 , w_41319 );
not ( w_41319 , w_41321 );
and ( w_41321 , w_41320 , w_41318 );
or ( w_41318 , \2135_b1 , w_41322 );
or ( w_41319 , \2135_b0 , \2136_b0 );
not ( \2136_b0 , w_41323 );
and ( w_41323 , w_41322 , \2136_b1 );
or ( \2140_b1 , \2117_b1 , w_41326 );
or ( \2140_b0 , \2117_b0 , w_41325 );
not ( w_41325 , w_41327 );
and ( w_41327 , w_41326 , w_41324 );
or ( w_41324 , \2138_b1 , w_41328 );
or ( w_41325 , \2138_b0 , \2139_b0 );
not ( \2139_b0 , w_41329 );
and ( w_41329 , w_41328 , \2139_b1 );
or ( \2150_b1 , \2145_b1 , w_41332 );
or ( \2150_b0 , \2145_b0 , w_41331 );
not ( w_41331 , w_41333 );
and ( w_41333 , w_41332 , w_41330 );
or ( w_41330 , \2148_b1 , w_41334 );
or ( w_41331 , \2148_b0 , \2149_b0 );
not ( \2149_b0 , w_41335 );
and ( w_41335 , w_41334 , \2149_b1 );
or ( \2165_b1 , \2160_b1 , w_41338 );
or ( \2165_b0 , \2160_b0 , w_41337 );
not ( w_41337 , w_41339 );
and ( w_41339 , w_41338 , w_41336 );
or ( w_41336 , \2163_b1 , w_41340 );
or ( w_41337 , \2163_b0 , \2164_b0 );
not ( \2164_b0 , w_41341 );
and ( w_41341 , w_41340 , \2164_b1 );
or ( \2181_b1 , \2174_b1 , w_41344 );
or ( \2181_b0 , \2174_b0 , w_41343 );
not ( w_41343 , w_41345 );
and ( w_41345 , w_41344 , w_41342 );
or ( w_41342 , \2179_b1 , w_41346 );
or ( w_41343 , \2179_b0 , \2180_b0 );
not ( \2180_b0 , w_41347 );
and ( w_41347 , w_41346 , \2180_b1 );
or ( \2186_b1 , \2182_b1 , w_41350 );
or ( \2186_b0 , \2182_b0 , w_41349 );
not ( w_41349 , w_41351 );
and ( w_41351 , w_41350 , w_41348 );
or ( w_41348 , \2184_b1 , w_41352 );
or ( w_41349 , \2184_b0 , \2185_b0 );
not ( \2185_b0 , w_41353 );
and ( w_41353 , w_41352 , \2185_b1 );
or ( \2189_b1 , \2151_b1 , w_41356 );
or ( \2189_b0 , \2151_b0 , w_41355 );
not ( w_41355 , w_41357 );
and ( w_41357 , w_41356 , w_41354 );
or ( w_41354 , \2187_b1 , w_41358 );
or ( w_41355 , \2187_b0 , \2188_b0 );
not ( \2188_b0 , w_41359 );
and ( w_41359 , w_41358 , \2188_b1 );
or ( \2199_b1 , \2194_b1 , w_41362 );
or ( \2199_b0 , \2194_b0 , w_41361 );
not ( w_41361 , w_41363 );
and ( w_41363 , w_41362 , w_41360 );
or ( w_41360 , \2197_b1 , w_41364 );
or ( w_41361 , \2197_b0 , \2198_b0 );
not ( \2198_b0 , w_41365 );
and ( w_41365 , w_41364 , \2198_b1 );
or ( \2205_b1 , \2200_b1 , w_41368 );
or ( \2205_b0 , \2200_b0 , w_41367 );
not ( w_41367 , w_41369 );
and ( w_41369 , w_41368 , w_41366 );
or ( w_41366 , \2203_b1 , w_41370 );
or ( w_41367 , \2203_b0 , \2204_b0 );
not ( \2204_b0 , w_41371 );
and ( w_41371 , w_41370 , \2204_b1 );
or ( \2212_b1 , \2208_b1 , w_41374 );
or ( \2212_b0 , \2208_b0 , w_41373 );
not ( w_41373 , w_41375 );
and ( w_41375 , w_41374 , w_41372 );
or ( w_41372 , \2210_b1 , w_41376 );
or ( w_41373 , \2210_b0 , \2211_b0 );
not ( \2211_b0 , w_41377 );
and ( w_41377 , w_41376 , \2211_b1 );
or ( \2220_b1 , \2215_b1 , w_41380 );
or ( \2220_b0 , \2215_b0 , w_41379 );
not ( w_41379 , w_41381 );
and ( w_41381 , w_41380 , w_41378 );
or ( w_41378 , \2218_b1 , w_41382 );
or ( w_41379 , \2218_b0 , \2219_b0 );
not ( \2219_b0 , w_41383 );
and ( w_41383 , w_41382 , \2219_b1 );
or ( \2240_b1 , \2233_b1 , w_41386 );
or ( \2240_b0 , \2233_b0 , w_41385 );
not ( w_41385 , w_41387 );
and ( w_41387 , w_41386 , w_41384 );
or ( w_41384 , \2238_b1 , w_41388 );
or ( w_41385 , \2238_b0 , \2239_b0 );
not ( \2239_b0 , w_41389 );
and ( w_41389 , w_41388 , \2239_b1 );
or ( \2256_b1 , \2249_b1 , w_41392 );
or ( \2256_b0 , \2249_b0 , w_41391 );
not ( w_41391 , w_41393 );
and ( w_41393 , w_41392 , w_41390 );
or ( w_41390 , \2254_b1 , w_41394 );
or ( w_41391 , \2254_b0 , \2255_b0 );
not ( \2255_b0 , w_41395 );
and ( w_41395 , w_41394 , \2255_b1 );
or ( \2276_b1 , \2269_b1 , w_41398 );
or ( \2276_b0 , \2269_b0 , w_41397 );
not ( w_41397 , w_41399 );
and ( w_41399 , w_41398 , w_41396 );
or ( w_41396 , \2274_b1 , w_41400 );
or ( w_41397 , \2274_b0 , \2275_b0 );
not ( \2275_b0 , w_41401 );
and ( w_41401 , w_41400 , \2275_b1 );
or ( \2279_b1 , \2257_b1 , w_41404 );
or ( \2279_b0 , \2257_b0 , w_41403 );
not ( w_41403 , w_41405 );
and ( w_41405 , w_41404 , w_41402 );
or ( w_41402 , \2277_b1 , w_41406 );
or ( w_41403 , \2277_b0 , \2278_b0 );
not ( \2278_b0 , w_41407 );
and ( w_41407 , w_41406 , \2278_b1 );
or ( \2295_b1 , \2288_b1 , w_41410 );
or ( \2295_b0 , \2288_b0 , w_41409 );
not ( w_41409 , w_41411 );
and ( w_41411 , w_41410 , w_41408 );
or ( w_41408 , \2293_b1 , w_41412 );
or ( w_41409 , \2293_b0 , \2294_b0 );
not ( \2294_b0 , w_41413 );
and ( w_41413 , w_41412 , \2294_b1 );
or ( \2309_b1 , \2304_b1 , w_41416 );
or ( \2309_b0 , \2304_b0 , w_41415 );
not ( w_41415 , w_41417 );
and ( w_41417 , w_41416 , w_41414 );
or ( w_41414 , \2307_b1 , w_41418 );
or ( w_41415 , \2307_b0 , \2308_b0 );
not ( \2308_b0 , w_41419 );
and ( w_41419 , w_41418 , \2308_b1 );
or ( \2315_b1 , \2310_b1 , w_41422 );
or ( \2315_b0 , \2310_b0 , w_41421 );
not ( w_41421 , w_41423 );
and ( w_41423 , w_41422 , w_41420 );
or ( w_41420 , \2313_b1 , w_41424 );
or ( w_41421 , \2313_b0 , \2314_b0 );
not ( \2314_b0 , w_41425 );
and ( w_41425 , w_41424 , \2314_b1 );
or ( \2326_b1 , \2321_b1 , w_41428 );
or ( \2326_b0 , \2321_b0 , w_41427 );
not ( w_41427 , w_41429 );
and ( w_41429 , w_41428 , w_41426 );
or ( w_41426 , \2324_b1 , w_41430 );
or ( w_41427 , \2324_b0 , \2325_b0 );
not ( \2325_b0 , w_41431 );
and ( w_41431 , w_41430 , \2325_b1 );
or ( \2329_b1 , \2316_b1 , w_41434 );
or ( \2329_b0 , \2316_b0 , w_41433 );
not ( w_41433 , w_41435 );
and ( w_41435 , w_41434 , w_41432 );
or ( w_41432 , \2327_b1 , w_41436 );
or ( w_41433 , \2327_b0 , \2328_b0 );
not ( \2328_b0 , w_41437 );
and ( w_41437 , w_41436 , \2328_b1 );
or ( \2339_b1 , \2334_b1 , w_41440 );
or ( \2339_b0 , \2334_b0 , w_41439 );
not ( w_41439 , w_41441 );
and ( w_41441 , w_41440 , w_41438 );
or ( w_41438 , \2337_b1 , w_41442 );
or ( w_41439 , \2337_b0 , \2338_b0 );
not ( \2338_b0 , w_41443 );
and ( w_41443 , w_41442 , \2338_b1 );
or ( \2345_b1 , \2340_b1 , w_41446 );
or ( \2345_b0 , \2340_b0 , w_41445 );
not ( w_41445 , w_41447 );
and ( w_41447 , w_41446 , w_41444 );
or ( w_41444 , \2343_b1 , w_41448 );
or ( w_41445 , \2343_b0 , \2344_b0 );
not ( \2344_b0 , w_41449 );
and ( w_41449 , w_41448 , \2344_b1 );
or ( \2355_b1 , \2350_b1 , w_41452 );
or ( \2355_b0 , \2350_b0 , w_41451 );
not ( w_41451 , w_41453 );
and ( w_41453 , w_41452 , w_41450 );
or ( w_41450 , \2353_b1 , w_41454 );
or ( w_41451 , \2353_b0 , \2354_b0 );
not ( \2354_b0 , w_41455 );
and ( w_41455 , w_41454 , \2354_b1 );
or ( \2361_b1 , \2356_b1 , w_41458 );
or ( \2361_b0 , \2356_b0 , w_41457 );
not ( w_41457 , w_41459 );
and ( w_41459 , w_41458 , w_41456 );
or ( w_41456 , \2359_b1 , w_41460 );
or ( w_41457 , \2359_b0 , \2360_b0 );
not ( \2360_b0 , w_41461 );
and ( w_41461 , w_41460 , \2360_b1 );
or ( \2387_b1 , \2380_b1 , w_41464 );
or ( \2387_b0 , \2380_b0 , w_41463 );
not ( w_41463 , w_41465 );
and ( w_41465 , w_41464 , w_41462 );
or ( w_41462 , \2385_b1 , w_41466 );
or ( w_41463 , \2385_b0 , \2386_b0 );
not ( \2386_b0 , w_41467 );
and ( w_41467 , w_41466 , \2386_b1 );
or ( \2403_b1 , \2396_b1 , w_41470 );
or ( \2403_b0 , \2396_b0 , w_41469 );
not ( w_41469 , w_41471 );
and ( w_41471 , w_41470 , w_41468 );
or ( w_41468 , \2401_b1 , w_41472 );
or ( w_41469 , \2401_b0 , \2402_b0 );
not ( \2402_b0 , w_41473 );
and ( w_41473 , w_41472 , \2402_b1 );
or ( \2420_b1 , \2413_b1 , w_41476 );
or ( \2420_b0 , \2413_b0 , w_41475 );
not ( w_41475 , w_41477 );
and ( w_41477 , w_41476 , w_41474 );
or ( w_41474 , \2418_b1 , w_41478 );
or ( w_41475 , \2418_b0 , \2419_b0 );
not ( \2419_b0 , w_41479 );
and ( w_41479 , w_41478 , \2419_b1 );
or ( \2423_b1 , \2404_b1 , w_41482 );
or ( \2423_b0 , \2404_b0 , w_41481 );
not ( w_41481 , w_41483 );
and ( w_41483 , w_41482 , w_41480 );
or ( w_41480 , \2421_b1 , w_41484 );
or ( w_41481 , \2421_b0 , \2422_b0 );
not ( \2422_b0 , w_41485 );
and ( w_41485 , w_41484 , \2422_b1 );
or ( \2433_b1 , \2428_b1 , w_41488 );
or ( \2433_b0 , \2428_b0 , w_41487 );
not ( w_41487 , w_41489 );
and ( w_41489 , w_41488 , w_41486 );
or ( w_41486 , \2431_b1 , w_41490 );
or ( w_41487 , \2431_b0 , \2432_b0 );
not ( \2432_b0 , w_41491 );
and ( w_41491 , w_41490 , \2432_b1 );
or ( \2450_b1 , \2443_b1 , w_41494 );
or ( \2450_b0 , \2443_b0 , w_41493 );
not ( w_41493 , w_41495 );
and ( w_41495 , w_41494 , w_41492 );
or ( w_41492 , \2448_b1 , w_41496 );
or ( w_41493 , \2448_b0 , \2449_b0 );
not ( \2449_b0 , w_41497 );
and ( w_41497 , w_41496 , \2449_b1 );
or ( \2466_b1 , \2459_b1 , w_41500 );
or ( \2466_b0 , \2459_b0 , w_41499 );
not ( w_41499 , w_41501 );
and ( w_41501 , w_41500 , w_41498 );
or ( w_41498 , \2464_b1 , w_41502 );
or ( w_41499 , \2464_b0 , \2465_b0 );
not ( \2465_b0 , w_41503 );
and ( w_41503 , w_41502 , \2465_b1 );
or ( \2470_b1 , \2434_b1 , w_41506 );
or ( \2470_b0 , \2434_b0 , w_41505 );
not ( w_41505 , w_41507 );
and ( w_41507 , w_41506 , w_41504 );
or ( w_41504 , \2468_b1 , w_41508 );
or ( w_41505 , \2468_b0 , \2469_b0 );
not ( \2469_b0 , w_41509 );
and ( w_41509 , w_41508 , \2469_b1 );
or ( \2480_b1 , \2475_b1 , w_41512 );
or ( \2480_b0 , \2475_b0 , w_41511 );
not ( w_41511 , w_41513 );
and ( w_41513 , w_41512 , w_41510 );
or ( w_41510 , \2478_b1 , w_41514 );
or ( w_41511 , \2478_b0 , \2479_b0 );
not ( \2479_b0 , w_41515 );
and ( w_41515 , w_41514 , \2479_b1 );
or ( \2486_b1 , \2481_b1 , w_41518 );
or ( \2486_b0 , \2481_b0 , w_41517 );
not ( w_41517 , w_41519 );
and ( w_41519 , w_41518 , w_41516 );
or ( w_41516 , \2484_b1 , w_41520 );
or ( w_41517 , \2484_b0 , \2485_b0 );
not ( \2485_b0 , w_41521 );
and ( w_41521 , w_41520 , \2485_b1 );
or ( \2494_b1 , \2489_b1 , w_41524 );
or ( \2494_b0 , \2489_b0 , w_41523 );
not ( w_41523 , w_41525 );
and ( w_41525 , w_41524 , w_41522 );
or ( w_41522 , \2492_b1 , w_41526 );
or ( w_41523 , \2492_b0 , \2493_b0 );
not ( \2493_b0 , w_41527 );
and ( w_41527 , w_41526 , \2493_b1 );
or ( \2502_b1 , \2497_b1 , w_41530 );
or ( \2502_b0 , \2497_b0 , w_41529 );
not ( w_41529 , w_41531 );
and ( w_41531 , w_41530 , w_41528 );
or ( w_41528 , \2500_b1 , w_41532 );
or ( w_41529 , \2500_b0 , \2501_b0 );
not ( \2501_b0 , w_41533 );
and ( w_41533 , w_41532 , \2501_b1 );
or ( \2522_b1 , \2515_b1 , w_41536 );
or ( \2522_b0 , \2515_b0 , w_41535 );
not ( w_41535 , w_41537 );
and ( w_41537 , w_41536 , w_41534 );
or ( w_41534 , \2520_b1 , w_41538 );
or ( w_41535 , \2520_b0 , \2521_b0 );
not ( \2521_b0 , w_41539 );
and ( w_41539 , w_41538 , \2521_b1 );
or ( \2539_b1 , \2531_b1 , w_41542 );
or ( \2539_b0 , \2531_b0 , w_41541 );
not ( w_41541 , w_41543 );
and ( w_41543 , w_41542 , w_41540 );
or ( w_41540 , \2537_b1 , w_41544 );
or ( w_41541 , \2537_b0 , \2538_b0 );
not ( \2538_b0 , w_41545 );
and ( w_41545 , w_41544 , \2538_b1 );
or ( \2546_b1 , \2540_b1 , w_41548 );
or ( \2546_b0 , \2540_b0 , w_41547 );
not ( w_41547 , w_41549 );
and ( w_41549 , w_41548 , w_41546 );
or ( w_41546 , \2544_b1 , w_41550 );
or ( w_41547 , \2544_b0 , \2545_b0 );
not ( \2545_b0 , w_41551 );
and ( w_41551 , w_41550 , \2545_b1 );
or ( \2565_b1 , \2558_b1 , w_41554 );
or ( \2565_b0 , \2558_b0 , w_41553 );
not ( w_41553 , w_41555 );
and ( w_41555 , w_41554 , w_41552 );
or ( w_41552 , \2563_b1 , w_41556 );
or ( w_41553 , \2563_b0 , \2564_b0 );
not ( \2564_b0 , w_41557 );
and ( w_41557 , w_41556 , \2564_b1 );
or ( \2581_b1 , \2574_b1 , w_41560 );
or ( \2581_b0 , \2574_b0 , w_41559 );
not ( w_41559 , w_41561 );
and ( w_41561 , w_41560 , w_41558 );
or ( w_41558 , \2579_b1 , w_41562 );
or ( w_41559 , \2579_b0 , \2580_b0 );
not ( \2580_b0 , w_41563 );
and ( w_41563 , w_41562 , \2580_b1 );
or ( \2598_b1 , \2591_b1 , w_41566 );
or ( \2598_b0 , \2591_b0 , w_41565 );
not ( w_41565 , w_41567 );
and ( w_41567 , w_41566 , w_41564 );
or ( w_41564 , \2596_b1 , w_41568 );
or ( w_41565 , \2596_b0 , \2597_b0 );
not ( \2597_b0 , w_41569 );
and ( w_41569 , w_41568 , \2597_b1 );
or ( \2601_b1 , \2582_b1 , w_41572 );
or ( \2601_b0 , \2582_b0 , w_41571 );
not ( w_41571 , w_41573 );
and ( w_41573 , w_41572 , w_41570 );
or ( w_41570 , \2599_b1 , w_41574 );
or ( w_41571 , \2599_b0 , \2600_b0 );
not ( \2600_b0 , w_41575 );
and ( w_41575 , w_41574 , \2600_b1 );
or ( \2611_b1 , \2606_b1 , w_41578 );
or ( \2611_b0 , \2606_b0 , w_41577 );
not ( w_41577 , w_41579 );
and ( w_41579 , w_41578 , w_41576 );
or ( w_41576 , \2609_b1 , w_41580 );
or ( w_41577 , \2609_b0 , \2610_b0 );
not ( \2610_b0 , w_41581 );
and ( w_41581 , w_41580 , \2610_b1 );
or ( \2614_b1 , \2602_b1 , w_41584 );
or ( \2614_b0 , \2602_b0 , w_41583 );
not ( w_41583 , w_41585 );
and ( w_41585 , w_41584 , w_41582 );
or ( w_41582 , \2612_b1 , w_41586 );
or ( w_41583 , \2612_b0 , \2613_b0 );
not ( \2613_b0 , w_41587 );
and ( w_41587 , w_41586 , \2613_b1 );
or ( \2624_b1 , \2619_b1 , w_41590 );
or ( \2624_b0 , \2619_b0 , w_41589 );
not ( w_41589 , w_41591 );
and ( w_41591 , w_41590 , w_41588 );
or ( w_41588 , \2622_b1 , w_41592 );
or ( w_41589 , \2622_b0 , \2623_b0 );
not ( \2623_b0 , w_41593 );
and ( w_41593 , w_41592 , \2623_b1 );
or ( \2632_b1 , \2627_b1 , w_41596 );
or ( \2632_b0 , \2627_b0 , w_41595 );
not ( w_41595 , w_41597 );
and ( w_41597 , w_41596 , w_41594 );
or ( w_41594 , \2630_b1 , w_41598 );
or ( w_41595 , \2630_b0 , \2631_b0 );
not ( \2631_b0 , w_41599 );
and ( w_41599 , w_41598 , \2631_b1 );
or ( \2642_b1 , \2638_b1 , w_41602 );
or ( \2642_b0 , \2638_b0 , w_41601 );
not ( w_41601 , w_41603 );
and ( w_41603 , w_41602 , w_41600 );
or ( w_41600 , \2640_b1 , w_41604 );
or ( w_41601 , \2640_b0 , \2641_b0 );
not ( \2641_b0 , w_41605 );
and ( w_41605 , w_41604 , \2641_b1 );
or ( \2645_b1 , \2633_b1 , w_41608 );
or ( \2645_b0 , \2633_b0 , w_41607 );
not ( w_41607 , w_41609 );
and ( w_41609 , w_41608 , w_41606 );
or ( w_41606 , \2643_b1 , w_41610 );
or ( w_41607 , \2643_b0 , \2644_b0 );
not ( \2644_b0 , w_41611 );
and ( w_41611 , w_41610 , \2644_b1 );
or ( \2655_b1 , \2650_b1 , w_41614 );
or ( \2655_b0 , \2650_b0 , w_41613 );
not ( w_41613 , w_41615 );
and ( w_41615 , w_41614 , w_41612 );
or ( w_41612 , \2653_b1 , w_41616 );
or ( w_41613 , \2653_b0 , \2654_b0 );
not ( \2654_b0 , w_41617 );
and ( w_41617 , w_41616 , \2654_b1 );
or ( \2661_b1 , \2656_b1 , w_41620 );
or ( \2661_b0 , \2656_b0 , w_41619 );
not ( w_41619 , w_41621 );
and ( w_41621 , w_41620 , w_41618 );
or ( w_41618 , \2659_b1 , w_41622 );
or ( w_41619 , \2659_b0 , \2660_b0 );
not ( \2660_b0 , w_41623 );
and ( w_41623 , w_41622 , \2660_b1 );
or ( \2672_b1 , \2667_b1 , w_41626 );
or ( \2672_b0 , \2667_b0 , w_41625 );
not ( w_41625 , w_41627 );
and ( w_41627 , w_41626 , w_41624 );
or ( w_41624 , \2670_b1 , w_41628 );
or ( w_41625 , \2670_b0 , \2671_b0 );
not ( \2671_b0 , w_41629 );
and ( w_41629 , w_41628 , \2671_b1 );
or ( \2692_b1 , \2685_b1 , w_41632 );
or ( \2692_b0 , \2685_b0 , w_41631 );
not ( w_41631 , w_41633 );
and ( w_41633 , w_41632 , w_41630 );
or ( w_41630 , \2690_b1 , w_41634 );
or ( w_41631 , \2690_b0 , \2691_b0 );
not ( \2691_b0 , w_41635 );
and ( w_41635 , w_41634 , \2691_b1 );
or ( \2705_b1 , \2698_b1 , w_41638 );
or ( \2705_b0 , \2698_b0 , w_41637 );
not ( w_41637 , w_41639 );
and ( w_41639 , w_41638 , w_41636 );
or ( w_41636 , \2703_b1 , w_41640 );
or ( w_41637 , \2703_b0 , \2704_b0 );
not ( \2704_b0 , w_41641 );
and ( w_41641 , w_41640 , \2704_b1 );
or ( \2722_b1 , \2715_b1 , w_41644 );
or ( \2722_b0 , \2715_b0 , w_41643 );
not ( w_41643 , w_41645 );
and ( w_41645 , w_41644 , w_41642 );
or ( w_41642 , \2720_b1 , w_41646 );
or ( w_41643 , \2720_b0 , \2721_b0 );
not ( \2721_b0 , w_41647 );
and ( w_41647 , w_41646 , \2721_b1 );
or ( \2725_b1 , \2706_b1 , w_41650 );
or ( \2725_b0 , \2706_b0 , w_41649 );
not ( w_41649 , w_41651 );
and ( w_41651 , w_41650 , w_41648 );
or ( w_41648 , \2723_b1 , w_41652 );
or ( w_41649 , \2723_b0 , \2724_b0 );
not ( \2724_b0 , w_41653 );
and ( w_41653 , w_41652 , \2724_b1 );
or ( \2741_b1 , \2734_b1 , w_41656 );
or ( \2741_b0 , \2734_b0 , w_41655 );
not ( w_41655 , w_41657 );
and ( w_41657 , w_41656 , w_41654 );
or ( w_41654 , \2739_b1 , w_41658 );
or ( w_41655 , \2739_b0 , \2740_b0 );
not ( \2740_b0 , w_41659 );
and ( w_41659 , w_41658 , \2740_b1 );
or ( \2757_b1 , \2750_b1 , w_41662 );
or ( \2757_b0 , \2750_b0 , w_41661 );
not ( w_41661 , w_41663 );
and ( w_41663 , w_41662 , w_41660 );
or ( w_41660 , \2755_b1 , w_41664 );
or ( w_41661 , \2755_b0 , \2756_b0 );
not ( \2756_b0 , w_41665 );
and ( w_41665 , w_41664 , \2756_b1 );
or ( \2768_b1 , \2758_b1 , w_41668 );
or ( \2768_b0 , \2758_b0 , w_41667 );
not ( w_41667 , w_41669 );
and ( w_41669 , w_41668 , w_41666 );
or ( w_41666 , \2766_b1 , w_41670 );
or ( w_41667 , \2766_b0 , \2767_b0 );
not ( \2767_b0 , w_41671 );
and ( w_41671 , w_41670 , \2767_b1 );
or ( \2778_b1 , \2774_b1 , w_41674 );
or ( \2778_b0 , \2774_b0 , w_41673 );
not ( w_41673 , w_41675 );
and ( w_41675 , w_41674 , w_41672 );
or ( w_41672 , \2776_b1 , w_41676 );
or ( w_41673 , \2776_b0 , \2777_b0 );
not ( \2777_b0 , w_41677 );
and ( w_41677 , w_41676 , \2777_b1 );
or ( \2781_b1 , \2769_b1 , w_41680 );
or ( \2781_b0 , \2769_b0 , w_41679 );
not ( w_41679 , w_41681 );
and ( w_41681 , w_41680 , w_41678 );
or ( w_41678 , \2779_b1 , w_41682 );
or ( w_41679 , \2779_b0 , \2780_b0 );
not ( \2780_b0 , w_41683 );
and ( w_41683 , w_41682 , \2780_b1 );
or ( \2791_b1 , \2786_b1 , w_41686 );
or ( \2791_b0 , \2786_b0 , w_41685 );
not ( w_41685 , w_41687 );
and ( w_41687 , w_41686 , w_41684 );
or ( w_41684 , \2789_b1 , w_41688 );
or ( w_41685 , \2789_b0 , \2790_b0 );
not ( \2790_b0 , w_41689 );
and ( w_41689 , w_41688 , \2790_b1 );
or ( \2799_b1 , \2794_b1 , w_41692 );
or ( \2799_b0 , \2794_b0 , w_41691 );
not ( w_41691 , w_41693 );
and ( w_41693 , w_41692 , w_41690 );
or ( w_41690 , \2797_b1 , w_41694 );
or ( w_41691 , \2797_b0 , \2798_b0 );
not ( \2798_b0 , w_41695 );
and ( w_41695 , w_41694 , \2798_b1 );
or ( \2805_b1 , \2800_b1 , w_41698 );
or ( \2805_b0 , \2800_b0 , w_41697 );
not ( w_41697 , w_41699 );
and ( w_41699 , w_41698 , w_41696 );
or ( w_41696 , \2803_b1 , w_41700 );
or ( w_41697 , \2803_b0 , \2804_b0 );
not ( \2804_b0 , w_41701 );
and ( w_41701 , w_41700 , \2804_b1 );
or ( \2813_b1 , \2808_b1 , w_41704 );
or ( \2813_b0 , \2808_b0 , w_41703 );
not ( w_41703 , w_41705 );
and ( w_41705 , w_41704 , w_41702 );
or ( w_41702 , \2811_b1 , w_41706 );
or ( w_41703 , \2811_b0 , \2812_b0 );
not ( \2812_b0 , w_41707 );
and ( w_41707 , w_41706 , \2812_b1 );
or ( \2820_b1 , \2816_b1 , w_41710 );
or ( \2820_b0 , \2816_b0 , w_41709 );
not ( w_41709 , w_41711 );
and ( w_41711 , w_41710 , w_41708 );
or ( w_41708 , \2818_b1 , w_41712 );
or ( w_41709 , \2818_b0 , \2819_b0 );
not ( \2819_b0 , w_41713 );
and ( w_41713 , w_41712 , \2819_b1 );
or ( \2840_b1 , \2833_b1 , w_41716 );
or ( \2840_b0 , \2833_b0 , w_41715 );
not ( w_41715 , w_41717 );
and ( w_41717 , w_41716 , w_41714 );
or ( w_41714 , \2838_b1 , w_41718 );
or ( w_41715 , \2838_b0 , \2839_b0 );
not ( \2839_b0 , w_41719 );
and ( w_41719 , w_41718 , \2839_b1 );
or ( \2855_b1 , \2849_b1 , w_41722 );
or ( \2855_b0 , \2849_b0 , w_41721 );
not ( w_41721 , w_41723 );
and ( w_41723 , w_41722 , w_41720 );
or ( w_41720 , \2853_b1 , w_41724 );
or ( w_41721 , \2853_b0 , \2854_b0 );
not ( \2854_b0 , w_41725 );
and ( w_41725 , w_41724 , \2854_b1 );
or ( \2872_b1 , \2865_b1 , w_41728 );
or ( \2872_b0 , \2865_b0 , w_41727 );
not ( w_41727 , w_41729 );
and ( w_41729 , w_41728 , w_41726 );
or ( w_41726 , \2870_b1 , w_41730 );
or ( w_41727 , \2870_b0 , \2871_b0 );
not ( \2871_b0 , w_41731 );
and ( w_41731 , w_41730 , \2871_b1 );
or ( \2875_b1 , \2856_b1 , w_41734 );
or ( \2875_b0 , \2856_b0 , w_41733 );
not ( w_41733 , w_41735 );
and ( w_41735 , w_41734 , w_41732 );
or ( w_41732 , \2873_b1 , w_41736 );
or ( w_41733 , \2873_b0 , \2874_b0 );
not ( \2874_b0 , w_41737 );
and ( w_41737 , w_41736 , \2874_b1 );
or ( \2891_b1 , \2884_b1 , w_41740 );
or ( \2891_b0 , \2884_b0 , w_41739 );
not ( w_41739 , w_41741 );
and ( w_41741 , w_41740 , w_41738 );
or ( w_41738 , \2889_b1 , w_41742 );
or ( w_41739 , \2889_b0 , \2890_b0 );
not ( \2890_b0 , w_41743 );
and ( w_41743 , w_41742 , \2890_b1 );
or ( \2907_b1 , \2900_b1 , w_41746 );
or ( \2907_b0 , \2900_b0 , w_41745 );
not ( w_41745 , w_41747 );
and ( w_41747 , w_41746 , w_41744 );
or ( w_41744 , \2905_b1 , w_41748 );
or ( w_41745 , \2905_b0 , \2906_b0 );
not ( \2906_b0 , w_41749 );
and ( w_41749 , w_41748 , \2906_b1 );
or ( \2924_b1 , \2908_b1 , w_41752 );
or ( \2924_b0 , \2908_b0 , w_41751 );
not ( w_41751 , w_41753 );
and ( w_41753 , w_41752 , w_41750 );
or ( w_41750 , \2922_b1 , w_41754 );
or ( w_41751 , \2922_b0 , \2923_b0 );
not ( \2923_b0 , w_41755 );
and ( w_41755 , w_41754 , \2923_b1 );
or ( \2934_b1 , \2930_b1 , w_41758 );
or ( \2934_b0 , \2930_b0 , w_41757 );
not ( w_41757 , w_41759 );
and ( w_41759 , w_41758 , w_41756 );
or ( w_41756 , \2932_b1 , w_41760 );
or ( w_41757 , \2932_b0 , \2933_b0 );
not ( \2933_b0 , w_41761 );
and ( w_41761 , w_41760 , \2933_b1 );
or ( \2937_b1 , \2925_b1 , w_41764 );
or ( \2937_b0 , \2925_b0 , w_41763 );
not ( w_41763 , w_41765 );
and ( w_41765 , w_41764 , w_41762 );
or ( w_41762 , \2935_b1 , w_41766 );
or ( w_41763 , \2935_b0 , \2936_b0 );
not ( \2936_b0 , w_41767 );
and ( w_41767 , w_41766 , \2936_b1 );
or ( \2947_b1 , \2942_b1 , w_41770 );
or ( \2947_b0 , \2942_b0 , w_41769 );
not ( w_41769 , w_41771 );
and ( w_41771 , w_41770 , w_41768 );
or ( w_41768 , \2945_b1 , w_41772 );
or ( w_41769 , \2945_b0 , \2946_b0 );
not ( \2946_b0 , w_41773 );
and ( w_41773 , w_41772 , \2946_b1 );
or ( \2955_b1 , \2950_b1 , w_41776 );
or ( \2955_b0 , \2950_b0 , w_41775 );
not ( w_41775 , w_41777 );
and ( w_41777 , w_41776 , w_41774 );
or ( w_41774 , \2953_b1 , w_41778 );
or ( w_41775 , \2953_b0 , \2954_b0 );
not ( \2954_b0 , w_41779 );
and ( w_41779 , w_41778 , \2954_b1 );
or ( \2961_b1 , \2956_b1 , w_41782 );
or ( \2961_b0 , \2956_b0 , w_41781 );
not ( w_41781 , w_41783 );
and ( w_41783 , w_41782 , w_41780 );
or ( w_41780 , \2959_b1 , w_41784 );
or ( w_41781 , \2959_b0 , \2960_b0 );
not ( \2960_b0 , w_41785 );
and ( w_41785 , w_41784 , \2960_b1 );
or ( \2971_b1 , \2966_b1 , w_41788 );
or ( \2971_b0 , \2966_b0 , w_41787 );
not ( w_41787 , w_41789 );
and ( w_41789 , w_41788 , w_41786 );
or ( w_41786 , \2969_b1 , w_41790 );
or ( w_41787 , \2969_b0 , \2970_b0 );
not ( \2970_b0 , w_41791 );
and ( w_41791 , w_41790 , \2970_b1 );
or ( \2977_b1 , \2972_b1 , w_41794 );
or ( \2977_b0 , \2972_b0 , w_41793 );
not ( w_41793 , w_41795 );
and ( w_41795 , w_41794 , w_41792 );
or ( w_41792 , \2975_b1 , w_41796 );
or ( w_41793 , \2975_b0 , \2976_b0 );
not ( \2976_b0 , w_41797 );
and ( w_41797 , w_41796 , \2976_b1 );
or ( \2988_b1 , \2983_b1 , w_41800 );
or ( \2988_b0 , \2983_b0 , w_41799 );
not ( w_41799 , w_41801 );
and ( w_41801 , w_41800 , w_41798 );
or ( w_41798 , \2986_b1 , w_41802 );
or ( w_41799 , \2986_b0 , \2987_b0 );
not ( \2987_b0 , w_41803 );
and ( w_41803 , w_41802 , \2987_b1 );
or ( \3008_b1 , \3001_b1 , w_41806 );
or ( \3008_b0 , \3001_b0 , w_41805 );
not ( w_41805 , w_41807 );
and ( w_41807 , w_41806 , w_41804 );
or ( w_41804 , \3006_b1 , w_41808 );
or ( w_41805 , \3006_b0 , \3007_b0 );
not ( \3007_b0 , w_41809 );
and ( w_41809 , w_41808 , \3007_b1 );
or ( \3024_b1 , \3017_b1 , w_41812 );
or ( \3024_b0 , \3017_b0 , w_41811 );
not ( w_41811 , w_41813 );
and ( w_41813 , w_41812 , w_41810 );
or ( w_41810 , \3022_b1 , w_41814 );
or ( w_41811 , \3022_b0 , \3023_b0 );
not ( \3023_b0 , w_41815 );
and ( w_41815 , w_41814 , \3023_b1 );
or ( \3041_b1 , \3034_b1 , w_41818 );
or ( \3041_b0 , \3034_b0 , w_41817 );
not ( w_41817 , w_41819 );
and ( w_41819 , w_41818 , w_41816 );
or ( w_41816 , \3039_b1 , w_41820 );
or ( w_41817 , \3039_b0 , \3040_b0 );
not ( \3040_b0 , w_41821 );
and ( w_41821 , w_41820 , \3040_b1 );
or ( \3044_b1 , \3025_b1 , w_41824 );
or ( \3044_b0 , \3025_b0 , w_41823 );
not ( w_41823 , w_41825 );
and ( w_41825 , w_41824 , w_41822 );
or ( w_41822 , \3042_b1 , w_41826 );
or ( w_41823 , \3042_b0 , \3043_b0 );
not ( \3043_b0 , w_41827 );
and ( w_41827 , w_41826 , \3043_b1 );
or ( \3054_b1 , \3049_b1 , w_41830 );
or ( \3054_b0 , \3049_b0 , w_41829 );
not ( w_41829 , w_41831 );
and ( w_41831 , w_41830 , w_41828 );
or ( w_41828 , \3052_b1 , w_41832 );
or ( w_41829 , \3052_b0 , \3053_b0 );
not ( \3053_b0 , w_41833 );
and ( w_41833 , w_41832 , \3053_b1 );
or ( \3071_b1 , \3064_b1 , w_41836 );
or ( \3071_b0 , \3064_b0 , w_41835 );
not ( w_41835 , w_41837 );
and ( w_41837 , w_41836 , w_41834 );
or ( w_41834 , \3069_b1 , w_41838 );
or ( w_41835 , \3069_b0 , \3070_b0 );
not ( \3070_b0 , w_41839 );
and ( w_41839 , w_41838 , \3070_b1 );
or ( \3087_b1 , \3080_b1 , w_41842 );
or ( \3087_b0 , \3080_b0 , w_41841 );
not ( w_41841 , w_41843 );
and ( w_41843 , w_41842 , w_41840 );
or ( w_41840 , \3085_b1 , w_41844 );
or ( w_41841 , \3085_b0 , \3086_b0 );
not ( \3086_b0 , w_41845 );
and ( w_41845 , w_41844 , \3086_b1 );
or ( \3093_b1 , \3088_b1 , w_41848 );
or ( \3093_b0 , \3088_b0 , w_41847 );
not ( w_41847 , w_41849 );
and ( w_41849 , w_41848 , w_41846 );
or ( w_41846 , \3091_b1 , w_41850 );
or ( w_41847 , \3091_b0 , \3092_b0 );
not ( \3092_b0 , w_41851 );
and ( w_41851 , w_41850 , \3092_b1 );
or ( \3096_b1 , \3055_b1 , w_41854 );
or ( \3096_b0 , \3055_b0 , w_41853 );
not ( w_41853 , w_41855 );
and ( w_41855 , w_41854 , w_41852 );
or ( w_41852 , \3094_b1 , w_41856 );
or ( w_41853 , \3094_b0 , \3095_b0 );
not ( \3095_b0 , w_41857 );
and ( w_41857 , w_41856 , \3095_b1 );
or ( \3106_b1 , \3101_b1 , w_41860 );
or ( \3106_b0 , \3101_b0 , w_41859 );
not ( w_41859 , w_41861 );
and ( w_41861 , w_41860 , w_41858 );
or ( w_41858 , \3104_b1 , w_41862 );
or ( w_41859 , \3104_b0 , \3105_b0 );
not ( \3105_b0 , w_41863 );
and ( w_41863 , w_41862 , \3105_b1 );
or ( \3112_b1 , \3107_b1 , w_41866 );
or ( \3112_b0 , \3107_b0 , w_41865 );
not ( w_41865 , w_41867 );
and ( w_41867 , w_41866 , w_41864 );
or ( w_41864 , \3110_b1 , w_41868 );
or ( w_41865 , \3110_b0 , \3111_b0 );
not ( \3111_b0 , w_41869 );
and ( w_41869 , w_41868 , \3111_b1 );
or ( \3122_b1 , \3117_b1 , w_41872 );
or ( \3122_b0 , \3117_b0 , w_41871 );
not ( w_41871 , w_41873 );
and ( w_41873 , w_41872 , w_41870 );
or ( w_41870 , \3120_b1 , w_41874 );
or ( w_41871 , \3120_b0 , \3121_b0 );
not ( \3121_b0 , w_41875 );
and ( w_41875 , w_41874 , \3121_b1 );
or ( \3128_b1 , \3123_b1 , w_41878 );
or ( \3128_b0 , \3123_b0 , w_41877 );
not ( w_41877 , w_41879 );
and ( w_41879 , w_41878 , w_41876 );
or ( w_41876 , \3126_b1 , w_41880 );
or ( w_41877 , \3126_b0 , \3127_b0 );
not ( \3127_b0 , w_41881 );
and ( w_41881 , w_41880 , \3127_b1 );
or ( \3135_b1 , \3131_b1 , w_41884 );
or ( \3135_b0 , \3131_b0 , w_41883 );
not ( w_41883 , w_41885 );
and ( w_41885 , w_41884 , w_41882 );
or ( w_41882 , \3133_b1 , w_41886 );
or ( w_41883 , \3133_b0 , \3134_b0 );
not ( \3134_b0 , w_41887 );
and ( w_41887 , w_41886 , \3134_b1 );
or ( \3155_b1 , \3148_b1 , w_41890 );
or ( \3155_b0 , \3148_b0 , w_41889 );
not ( w_41889 , w_41891 );
and ( w_41891 , w_41890 , w_41888 );
or ( w_41888 , \3153_b1 , w_41892 );
or ( w_41889 , \3153_b0 , \3154_b0 );
not ( \3154_b0 , w_41893 );
and ( w_41893 , w_41892 , \3154_b1 );
or ( \3171_b1 , \3164_b1 , w_41896 );
or ( \3171_b0 , \3164_b0 , w_41895 );
not ( w_41895 , w_41897 );
and ( w_41897 , w_41896 , w_41894 );
or ( w_41894 , \3169_b1 , w_41898 );
or ( w_41895 , \3169_b0 , \3170_b0 );
not ( \3170_b0 , w_41899 );
and ( w_41899 , w_41898 , \3170_b1 );
or ( \3184_b1 , \3181_b1 , w_41902 );
or ( \3184_b0 , \3181_b0 , w_41901 );
not ( w_41901 , w_41903 );
and ( w_41903 , w_41902 , w_41900 );
or ( w_41900 , \3182_b1 , w_41904 );
or ( w_41901 , \3182_b0 , \3183_b0 );
not ( \3183_b0 , w_41905 );
and ( w_41905 , w_41904 , \3183_b1 );
or ( \3187_b1 , \3172_b1 , w_41908 );
or ( \3187_b0 , \3172_b0 , w_41907 );
not ( w_41907 , w_41909 );
and ( w_41909 , w_41908 , w_41906 );
or ( w_41906 , \3185_b1 , w_41910 );
or ( w_41907 , \3185_b0 , \3186_b0 );
not ( \3186_b0 , w_41911 );
and ( w_41911 , w_41910 , \3186_b1 );
or ( \3203_b1 , \3196_b1 , w_41914 );
or ( \3203_b0 , \3196_b0 , w_41913 );
not ( w_41913 , w_41915 );
and ( w_41915 , w_41914 , w_41912 );
or ( w_41912 , \3201_b1 , w_41916 );
or ( w_41913 , \3201_b0 , \3202_b0 );
not ( \3202_b0 , w_41917 );
and ( w_41917 , w_41916 , \3202_b1 );
or ( \3219_b1 , \3212_b1 , w_41920 );
or ( \3219_b0 , \3212_b0 , w_41919 );
not ( w_41919 , w_41921 );
and ( w_41921 , w_41920 , w_41918 );
or ( w_41918 , \3217_b1 , w_41922 );
or ( w_41919 , \3217_b0 , \3218_b0 );
not ( \3218_b0 , w_41923 );
and ( w_41923 , w_41922 , \3218_b1 );
or ( \3227_b1 , \3220_b1 , w_41926 );
or ( \3227_b0 , \3220_b0 , w_41925 );
not ( w_41925 , w_41927 );
and ( w_41927 , w_41926 , w_41924 );
or ( w_41924 , \3225_b1 , w_41928 );
or ( w_41925 , \3225_b0 , \3226_b0 );
not ( \3226_b0 , w_41929 );
and ( w_41929 , w_41928 , \3226_b1 );
or ( \3238_b1 , \3233_b1 , w_41932 );
or ( \3238_b0 , \3233_b0 , w_41931 );
not ( w_41931 , w_41933 );
and ( w_41933 , w_41932 , w_41930 );
or ( w_41930 , \3236_b1 , w_41934 );
or ( w_41931 , \3236_b0 , \3237_b0 );
not ( \3237_b0 , w_41935 );
and ( w_41935 , w_41934 , \3237_b1 );
or ( \3241_b1 , \3228_b1 , w_41938 );
or ( \3241_b0 , \3228_b0 , w_41937 );
not ( w_41937 , w_41939 );
and ( w_41939 , w_41938 , w_41936 );
or ( w_41936 , \3239_b1 , w_41940 );
or ( w_41937 , \3239_b0 , \3240_b0 );
not ( \3240_b0 , w_41941 );
and ( w_41941 , w_41940 , \3240_b1 );
or ( \3250_b1 , \3246_b1 , w_41944 );
or ( \3250_b0 , \3246_b0 , w_41943 );
not ( w_41943 , w_41945 );
and ( w_41945 , w_41944 , w_41942 );
or ( w_41942 , \3248_b1 , w_41946 );
or ( w_41943 , \3248_b0 , \3249_b0 );
not ( \3249_b0 , w_41947 );
and ( w_41947 , w_41946 , \3249_b1 );
or ( \3259_b1 , \3251_b1 , w_41950 );
or ( \3259_b0 , \3251_b0 , w_41949 );
not ( w_41949 , w_41951 );
and ( w_41951 , w_41950 , w_41948 );
or ( w_41948 , \3257_b1 , w_41952 );
or ( w_41949 , \3257_b0 , \3258_b0 );
not ( \3258_b0 , w_41953 );
and ( w_41953 , w_41952 , \3258_b1 );
or ( \3269_b1 , \3264_b1 , w_41956 );
or ( \3269_b0 , \3264_b0 , w_41955 );
not ( w_41955 , w_41957 );
and ( w_41957 , w_41956 , w_41954 );
or ( w_41954 , \3267_b1 , w_41958 );
or ( w_41955 , \3267_b0 , \3268_b0 );
not ( \3268_b0 , w_41959 );
and ( w_41959 , w_41958 , \3268_b1 );
or ( \3275_b1 , \3270_b1 , w_41962 );
or ( \3275_b0 , \3270_b0 , w_41961 );
not ( w_41961 , w_41963 );
and ( w_41963 , w_41962 , w_41960 );
or ( w_41960 , \3273_b1 , w_41964 );
or ( w_41961 , \3273_b0 , \3274_b0 );
not ( \3274_b0 , w_41965 );
and ( w_41965 , w_41964 , \3274_b1 );
or ( \3283_b1 , \3278_b1 , w_41968 );
or ( \3283_b0 , \3278_b0 , w_41967 );
not ( w_41967 , w_41969 );
and ( w_41969 , w_41968 , w_41966 );
or ( w_41966 , \3281_b1 , w_41970 );
or ( w_41967 , \3281_b0 , \3282_b0 );
not ( \3282_b0 , w_41971 );
and ( w_41971 , w_41970 , \3282_b1 );
or ( \3303_b1 , \3296_b1 , w_41974 );
or ( \3303_b0 , \3296_b0 , w_41973 );
not ( w_41973 , w_41975 );
and ( w_41975 , w_41974 , w_41972 );
or ( w_41972 , \3301_b1 , w_41976 );
or ( w_41973 , \3301_b0 , \3302_b0 );
not ( \3302_b0 , w_41977 );
and ( w_41977 , w_41976 , \3302_b1 );
or ( \3319_b1 , \3312_b1 , w_41980 );
or ( \3319_b0 , \3312_b0 , w_41979 );
not ( w_41979 , w_41981 );
and ( w_41981 , w_41980 , w_41978 );
or ( w_41978 , \3317_b1 , w_41982 );
or ( w_41979 , \3317_b0 , \3318_b0 );
not ( \3318_b0 , w_41983 );
and ( w_41983 , w_41982 , \3318_b1 );
or ( \3336_b1 , \3329_b1 , w_41986 );
or ( \3336_b0 , \3329_b0 , w_41985 );
not ( w_41985 , w_41987 );
and ( w_41987 , w_41986 , w_41984 );
or ( w_41984 , \3334_b1 , w_41988 );
or ( w_41985 , \3334_b0 , \3335_b0 );
not ( \3335_b0 , w_41989 );
and ( w_41989 , w_41988 , \3335_b1 );
or ( \3339_b1 , \3320_b1 , w_41992 );
or ( \3339_b0 , \3320_b0 , w_41991 );
not ( w_41991 , w_41993 );
and ( w_41993 , w_41992 , w_41990 );
or ( w_41990 , \3337_b1 , w_41994 );
or ( w_41991 , \3337_b0 , \3338_b0 );
not ( \3338_b0 , w_41995 );
and ( w_41995 , w_41994 , \3338_b1 );
or ( \3355_b1 , \3348_b1 , w_41998 );
or ( \3355_b0 , \3348_b0 , w_41997 );
not ( w_41997 , w_41999 );
and ( w_41999 , w_41998 , w_41996 );
or ( w_41996 , \3353_b1 , w_42000 );
or ( w_41997 , \3353_b0 , \3354_b0 );
not ( \3354_b0 , w_42001 );
and ( w_42001 , w_42000 , \3354_b1 );
or ( \3371_b1 , \3364_b1 , w_42004 );
or ( \3371_b0 , \3364_b0 , w_42003 );
not ( w_42003 , w_42005 );
and ( w_42005 , w_42004 , w_42002 );
or ( w_42002 , \3369_b1 , w_42006 );
or ( w_42003 , \3369_b0 , \3370_b0 );
not ( \3370_b0 , w_42007 );
and ( w_42007 , w_42006 , \3370_b1 );
or ( \3379_b1 , \3372_b1 , w_42010 );
or ( \3379_b0 , \3372_b0 , w_42009 );
not ( w_42009 , w_42011 );
and ( w_42011 , w_42010 , w_42008 );
or ( w_42008 , \3377_b1 , w_42012 );
or ( w_42009 , \3377_b0 , \3378_b0 );
not ( \3378_b0 , w_42013 );
and ( w_42013 , w_42012 , \3378_b1 );
or ( \3390_b1 , \3385_b1 , w_42016 );
or ( \3390_b0 , \3385_b0 , w_42015 );
not ( w_42015 , w_42017 );
and ( w_42017 , w_42016 , w_42014 );
or ( w_42014 , \3388_b1 , w_42018 );
or ( w_42015 , \3388_b0 , \3389_b0 );
not ( \3389_b0 , w_42019 );
and ( w_42019 , w_42018 , \3389_b1 );
or ( \3393_b1 , \3380_b1 , w_42022 );
or ( \3393_b0 , \3380_b0 , w_42021 );
not ( w_42021 , w_42023 );
and ( w_42023 , w_42022 , w_42020 );
or ( w_42020 , \3391_b1 , w_42024 );
or ( w_42021 , \3391_b0 , \3392_b0 );
not ( \3392_b0 , w_42025 );
and ( w_42025 , w_42024 , \3392_b1 );
or ( \3403_b1 , \3398_b1 , w_42028 );
or ( \3403_b0 , \3398_b0 , w_42027 );
not ( w_42027 , w_42029 );
and ( w_42029 , w_42028 , w_42026 );
or ( w_42026 , \3401_b1 , w_42030 );
or ( w_42027 , \3401_b0 , \3402_b0 );
not ( \3402_b0 , w_42031 );
and ( w_42031 , w_42030 , \3402_b1 );
or ( \3411_b1 , \3406_b1 , w_42034 );
or ( \3411_b0 , \3406_b0 , w_42033 );
not ( w_42033 , w_42035 );
and ( w_42035 , w_42034 , w_42032 );
or ( w_42032 , \3409_b1 , w_42036 );
or ( w_42033 , \3409_b0 , \3410_b0 );
not ( \3410_b0 , w_42037 );
and ( w_42037 , w_42036 , \3410_b1 );
or ( \3422_b1 , \3417_b1 , w_42040 );
or ( \3422_b0 , \3417_b0 , w_42039 );
not ( w_42039 , w_42041 );
and ( w_42041 , w_42040 , w_42038 );
or ( w_42038 , \3420_b1 , w_42042 );
or ( w_42039 , \3420_b0 , \3421_b0 );
not ( \3421_b0 , w_42043 );
and ( w_42043 , w_42042 , \3421_b1 );
or ( \3425_b1 , \3412_b1 , w_42046 );
or ( \3425_b0 , \3412_b0 , w_42045 );
not ( w_42045 , w_42047 );
and ( w_42047 , w_42046 , w_42044 );
or ( w_42044 , \3423_b1 , w_42048 );
or ( w_42045 , \3423_b0 , \3424_b0 );
not ( \3424_b0 , w_42049 );
and ( w_42049 , w_42048 , \3424_b1 );
or ( \3434_b1 , \3430_b1 , w_42052 );
or ( \3434_b0 , \3430_b0 , w_42051 );
not ( w_42051 , w_42053 );
and ( w_42053 , w_42052 , w_42050 );
or ( w_42050 , \3432_b1 , w_42054 );
or ( w_42051 , \3432_b0 , \3433_b0 );
not ( \3433_b0 , w_42055 );
and ( w_42055 , w_42054 , \3433_b1 );
or ( \3440_b1 , \3435_b1 , w_42058 );
or ( \3440_b0 , \3435_b0 , w_42057 );
not ( w_42057 , w_42059 );
and ( w_42059 , w_42058 , w_42056 );
or ( w_42056 , \3438_b1 , w_42060 );
or ( w_42057 , \3438_b0 , \3439_b0 );
not ( \3439_b0 , w_42061 );
and ( w_42061 , w_42060 , \3439_b1 );
or ( \3448_b1 , \3443_b1 , w_42064 );
or ( \3448_b0 , \3443_b0 , w_42063 );
not ( w_42063 , w_42065 );
and ( w_42065 , w_42064 , w_42062 );
or ( w_42062 , \3446_b1 , w_42066 );
or ( w_42063 , \3446_b0 , \3447_b0 );
not ( \3447_b0 , w_42067 );
and ( w_42067 , w_42066 , \3447_b1 );
or ( \3468_b1 , \3461_b1 , w_42070 );
or ( \3468_b0 , \3461_b0 , w_42069 );
not ( w_42069 , w_42071 );
and ( w_42071 , w_42070 , w_42068 );
or ( w_42068 , \3466_b1 , w_42072 );
or ( w_42069 , \3466_b0 , \3467_b0 );
not ( \3467_b0 , w_42073 );
and ( w_42073 , w_42072 , \3467_b1 );
or ( \3484_b1 , \3477_b1 , w_42076 );
or ( \3484_b0 , \3477_b0 , w_42075 );
not ( w_42075 , w_42077 );
and ( w_42077 , w_42076 , w_42074 );
or ( w_42074 , \3482_b1 , w_42078 );
or ( w_42075 , \3482_b0 , \3483_b0 );
not ( \3483_b0 , w_42079 );
and ( w_42079 , w_42078 , \3483_b1 );
or ( \3497_b1 , \3494_b1 , w_42082 );
or ( \3497_b0 , \3494_b0 , w_42081 );
not ( w_42081 , w_42083 );
and ( w_42083 , w_42082 , w_42080 );
or ( w_42080 , \3495_b1 , w_42084 );
or ( w_42081 , \3495_b0 , \3496_b0 );
not ( \3496_b0 , w_42085 );
and ( w_42085 , w_42084 , \3496_b1 );
or ( \3500_b1 , \3485_b1 , w_42088 );
or ( \3500_b0 , \3485_b0 , w_42087 );
not ( w_42087 , w_42089 );
and ( w_42089 , w_42088 , w_42086 );
or ( w_42086 , \3498_b1 , w_42090 );
or ( w_42087 , \3498_b0 , \3499_b0 );
not ( \3499_b0 , w_42091 );
and ( w_42091 , w_42090 , \3499_b1 );
or ( \3516_b1 , \3509_b1 , w_42094 );
or ( \3516_b0 , \3509_b0 , w_42093 );
not ( w_42093 , w_42095 );
and ( w_42095 , w_42094 , w_42092 );
or ( w_42092 , \3514_b1 , w_42096 );
or ( w_42093 , \3514_b0 , \3515_b0 );
not ( \3515_b0 , w_42097 );
and ( w_42097 , w_42096 , \3515_b1 );
or ( \3532_b1 , \3525_b1 , w_42100 );
or ( \3532_b0 , \3525_b0 , w_42099 );
not ( w_42099 , w_42101 );
and ( w_42101 , w_42100 , w_42098 );
or ( w_42098 , \3530_b1 , w_42102 );
or ( w_42099 , \3530_b0 , \3531_b0 );
not ( \3531_b0 , w_42103 );
and ( w_42103 , w_42102 , \3531_b1 );
or ( \3538_b1 , \3533_b1 , w_42106 );
or ( \3538_b0 , \3533_b0 , w_42105 );
not ( w_42105 , w_42107 );
and ( w_42107 , w_42106 , w_42104 );
or ( w_42104 , \3536_b1 , w_42108 );
or ( w_42105 , \3536_b0 , \3537_b0 );
not ( \3537_b0 , w_42109 );
and ( w_42109 , w_42108 , \3537_b1 );
or ( \3549_b1 , \3544_b1 , w_42112 );
or ( \3549_b0 , \3544_b0 , w_42111 );
not ( w_42111 , w_42113 );
and ( w_42113 , w_42112 , w_42110 );
or ( w_42110 , \3547_b1 , w_42114 );
or ( w_42111 , \3547_b0 , \3548_b0 );
not ( \3548_b0 , w_42115 );
and ( w_42115 , w_42114 , \3548_b1 );
or ( \3552_b1 , \3539_b1 , w_42118 );
or ( \3552_b0 , \3539_b0 , w_42117 );
not ( w_42117 , w_42119 );
and ( w_42119 , w_42118 , w_42116 );
or ( w_42116 , \3550_b1 , w_42120 );
or ( w_42117 , \3550_b0 , \3551_b0 );
not ( \3551_b0 , w_42121 );
and ( w_42121 , w_42120 , \3551_b1 );
or ( \3562_b1 , \3557_b1 , w_42124 );
or ( \3562_b0 , \3557_b0 , w_42123 );
not ( w_42123 , w_42125 );
and ( w_42125 , w_42124 , w_42122 );
or ( w_42122 , \3560_b1 , w_42126 );
or ( w_42123 , \3560_b0 , \3561_b0 );
not ( \3561_b0 , w_42127 );
and ( w_42127 , w_42126 , \3561_b1 );
or ( \3568_b1 , \3563_b1 , w_42130 );
or ( \3568_b0 , \3563_b0 , w_42129 );
not ( w_42129 , w_42131 );
and ( w_42131 , w_42130 , w_42128 );
or ( w_42128 , \3566_b1 , w_42132 );
or ( w_42129 , \3566_b0 , \3567_b0 );
not ( \3567_b0 , w_42133 );
and ( w_42133 , w_42132 , \3567_b1 );
or ( \3579_b1 , \3574_b1 , w_42136 );
or ( \3579_b0 , \3574_b0 , w_42135 );
not ( w_42135 , w_42137 );
and ( w_42137 , w_42136 , w_42134 );
or ( w_42134 , \3577_b1 , w_42138 );
or ( w_42135 , \3577_b0 , \3578_b0 );
not ( \3578_b0 , w_42139 );
and ( w_42139 , w_42138 , \3578_b1 );
or ( \3587_b1 , \3582_b1 , w_42142 );
or ( \3587_b0 , \3582_b0 , w_42141 );
not ( w_42141 , w_42143 );
and ( w_42143 , w_42142 , w_42140 );
or ( w_42140 , \3585_b1 , w_42144 );
or ( w_42141 , \3585_b0 , \3586_b0 );
not ( \3586_b0 , w_42145 );
and ( w_42145 , w_42144 , \3586_b1 );
or ( \3607_b1 , \3600_b1 , w_42148 );
or ( \3607_b0 , \3600_b0 , w_42147 );
not ( w_42147 , w_42149 );
and ( w_42149 , w_42148 , w_42146 );
or ( w_42146 , \3605_b1 , w_42150 );
or ( w_42147 , \3605_b0 , \3606_b0 );
not ( \3606_b0 , w_42151 );
and ( w_42151 , w_42150 , \3606_b1 );
or ( \3623_b1 , \3616_b1 , w_42154 );
or ( \3623_b0 , \3616_b0 , w_42153 );
not ( w_42153 , w_42155 );
and ( w_42155 , w_42154 , w_42152 );
or ( w_42152 , \3621_b1 , w_42156 );
or ( w_42153 , \3621_b0 , \3622_b0 );
not ( \3622_b0 , w_42157 );
and ( w_42157 , w_42156 , \3622_b1 );
or ( \3640_b1 , \3633_b1 , w_42160 );
or ( \3640_b0 , \3633_b0 , w_42159 );
not ( w_42159 , w_42161 );
and ( w_42161 , w_42160 , w_42158 );
or ( w_42158 , \3638_b1 , w_42162 );
or ( w_42159 , \3638_b0 , \3639_b0 );
not ( \3639_b0 , w_42163 );
and ( w_42163 , w_42162 , \3639_b1 );
or ( \3643_b1 , \3624_b1 , w_42166 );
or ( \3643_b0 , \3624_b0 , w_42165 );
not ( w_42165 , w_42167 );
and ( w_42167 , w_42166 , w_42164 );
or ( w_42164 , \3641_b1 , w_42168 );
or ( w_42165 , \3641_b0 , \3642_b0 );
not ( \3642_b0 , w_42169 );
and ( w_42169 , w_42168 , \3642_b1 );
or ( \3653_b1 , \3648_b1 , w_42172 );
or ( \3653_b0 , \3648_b0 , w_42171 );
not ( w_42171 , w_42173 );
and ( w_42173 , w_42172 , w_42170 );
or ( w_42170 , \3651_b1 , w_42174 );
or ( w_42171 , \3651_b0 , \3652_b0 );
not ( \3652_b0 , w_42175 );
and ( w_42175 , w_42174 , \3652_b1 );
or ( \3670_b1 , \3663_b1 , w_42178 );
or ( \3670_b0 , \3663_b0 , w_42177 );
not ( w_42177 , w_42179 );
and ( w_42179 , w_42178 , w_42176 );
or ( w_42176 , \3668_b1 , w_42180 );
or ( w_42177 , \3668_b0 , \3669_b0 );
not ( \3669_b0 , w_42181 );
and ( w_42181 , w_42180 , \3669_b1 );
or ( \3678_b1 , \3673_b1 , w_42184 );
or ( \3678_b0 , \3673_b0 , w_42183 );
not ( w_42183 , w_42185 );
and ( w_42185 , w_42184 , w_42182 );
or ( w_42182 , \3676_b1 , w_42186 );
or ( w_42183 , \3676_b0 , \3677_b0 );
not ( \3677_b0 , w_42187 );
and ( w_42187 , w_42186 , \3677_b1 );
or ( \3681_b1 , \3654_b1 , w_42190 );
or ( \3681_b0 , \3654_b0 , w_42189 );
not ( w_42189 , w_42191 );
and ( w_42191 , w_42190 , w_42188 );
or ( w_42188 , \3679_b1 , w_42192 );
or ( w_42189 , \3679_b0 , \3680_b0 );
not ( \3680_b0 , w_42193 );
and ( w_42193 , w_42192 , \3680_b1 );
or ( \3691_b1 , \3686_b1 , w_42196 );
or ( \3691_b0 , \3686_b0 , w_42195 );
not ( w_42195 , w_42197 );
and ( w_42197 , w_42196 , w_42194 );
or ( w_42194 , \3689_b1 , w_42198 );
or ( w_42195 , \3689_b0 , \3690_b0 );
not ( \3690_b0 , w_42199 );
and ( w_42199 , w_42198 , \3690_b1 );
or ( \3697_b1 , \3692_b1 , w_42202 );
or ( \3697_b0 , \3692_b0 , w_42201 );
not ( w_42201 , w_42203 );
and ( w_42203 , w_42202 , w_42200 );
or ( w_42200 , \3695_b1 , w_42204 );
or ( w_42201 , \3695_b0 , \3696_b0 );
not ( \3696_b0 , w_42205 );
and ( w_42205 , w_42204 , \3696_b1 );
or ( \3704_b1 , \3700_b1 , w_42208 );
or ( \3704_b0 , \3700_b0 , w_42207 );
not ( w_42207 , w_42209 );
and ( w_42209 , w_42208 , w_42206 );
or ( w_42206 , \3702_b1 , w_42210 );
or ( w_42207 , \3702_b0 , \3703_b0 );
not ( \3703_b0 , w_42211 );
and ( w_42211 , w_42210 , \3703_b1 );
or ( \3712_b1 , \3707_b1 , w_42214 );
or ( \3712_b0 , \3707_b0 , w_42213 );
not ( w_42213 , w_42215 );
and ( w_42215 , w_42214 , w_42212 );
or ( w_42212 , \3710_b1 , w_42216 );
or ( w_42213 , \3710_b0 , \3711_b0 );
not ( \3711_b0 , w_42217 );
and ( w_42217 , w_42216 , \3711_b1 );
or ( \3732_b1 , \3725_b1 , w_42220 );
or ( \3732_b0 , \3725_b0 , w_42219 );
not ( w_42219 , w_42221 );
and ( w_42221 , w_42220 , w_42218 );
or ( w_42218 , \3730_b1 , w_42222 );
or ( w_42219 , \3730_b0 , \3731_b0 );
not ( \3731_b0 , w_42223 );
and ( w_42223 , w_42222 , \3731_b1 );
or ( \3746_b1 , \3741_b1 , w_42226 );
or ( \3746_b0 , \3741_b0 , w_42225 );
not ( w_42225 , w_42227 );
and ( w_42227 , w_42226 , w_42224 );
or ( w_42224 , \3744_b1 , w_42228 );
or ( w_42225 , \3744_b0 , \3745_b0 );
not ( \3745_b0 , w_42229 );
and ( w_42229 , w_42228 , \3745_b1 );
or ( \3754_b1 , \3747_b1 , w_42232 );
or ( \3754_b0 , \3747_b0 , w_42231 );
not ( w_42231 , w_42233 );
and ( w_42233 , w_42232 , w_42230 );
or ( w_42230 , \3752_b1 , w_42234 );
or ( w_42231 , \3752_b0 , \3753_b0 );
not ( \3753_b0 , w_42235 );
and ( w_42235 , w_42234 , \3753_b1 );
or ( \3770_b1 , \3763_b1 , w_42238 );
or ( \3770_b0 , \3763_b0 , w_42237 );
not ( w_42237 , w_42239 );
and ( w_42239 , w_42238 , w_42236 );
or ( w_42236 , \3768_b1 , w_42240 );
or ( w_42237 , \3768_b0 , \3769_b0 );
not ( \3769_b0 , w_42241 );
and ( w_42241 , w_42240 , \3769_b1 );
or ( \3782_b1 , \3779_b1 , w_42244 );
or ( \3782_b0 , \3779_b0 , w_42243 );
not ( w_42243 , w_42245 );
and ( w_42245 , w_42244 , w_42242 );
or ( w_42242 , \3780_b1 , w_42246 );
or ( w_42243 , \3780_b0 , \3781_b0 );
not ( \3781_b0 , w_42247 );
and ( w_42247 , w_42246 , \3781_b1 );
or ( \3799_b1 , \3792_b1 , w_42250 );
or ( \3799_b0 , \3792_b0 , w_42249 );
not ( w_42249 , w_42251 );
and ( w_42251 , w_42250 , w_42248 );
or ( w_42248 , \3797_b1 , w_42252 );
or ( w_42249 , \3797_b0 , \3798_b0 );
not ( \3798_b0 , w_42253 );
and ( w_42253 , w_42252 , \3798_b1 );
or ( \3802_b1 , \3783_b1 , w_42256 );
or ( \3802_b0 , \3783_b0 , w_42255 );
not ( w_42255 , w_42257 );
and ( w_42257 , w_42256 , w_42254 );
or ( w_42254 , \3800_b1 , w_42258 );
or ( w_42255 , \3800_b0 , \3801_b0 );
not ( \3801_b0 , w_42259 );
and ( w_42259 , w_42258 , \3801_b1 );
or ( \3815_b1 , \3810_b1 , w_42262 );
or ( \3815_b0 , \3810_b0 , w_42261 );
not ( w_42261 , w_42263 );
and ( w_42263 , w_42262 , w_42260 );
or ( w_42260 , \3813_b1 , w_42264 );
or ( w_42261 , \3813_b0 , \3814_b0 );
not ( \3814_b0 , w_42265 );
and ( w_42265 , w_42264 , \3814_b1 );
or ( \3818_b1 , \3803_b1 , w_42268 );
or ( \3818_b0 , \3803_b0 , w_42267 );
not ( w_42267 , w_42269 );
and ( w_42269 , w_42268 , w_42266 );
or ( w_42266 , \3816_b1 , w_42270 );
or ( w_42267 , \3816_b0 , \3817_b0 );
not ( \3817_b0 , w_42271 );
and ( w_42271 , w_42270 , \3817_b1 );
or ( \3828_b1 , \3823_b1 , w_42274 );
or ( \3828_b0 , \3823_b0 , w_42273 );
not ( w_42273 , w_42275 );
and ( w_42275 , w_42274 , w_42272 );
or ( w_42272 , \3826_b1 , w_42276 );
or ( w_42273 , \3826_b0 , \3827_b0 );
not ( \3827_b0 , w_42277 );
and ( w_42277 , w_42276 , \3827_b1 );
or ( \3834_b1 , \3829_b1 , w_42280 );
or ( \3834_b0 , \3829_b0 , w_42279 );
not ( w_42279 , w_42281 );
and ( w_42281 , w_42280 , w_42278 );
or ( w_42278 , \3832_b1 , w_42282 );
or ( w_42279 , \3832_b0 , \3833_b0 );
not ( \3833_b0 , w_42283 );
and ( w_42283 , w_42282 , \3833_b1 );
or ( \3845_b1 , \3840_b1 , w_42286 );
or ( \3845_b0 , \3840_b0 , w_42285 );
not ( w_42285 , w_42287 );
and ( w_42287 , w_42286 , w_42284 );
or ( w_42284 , \3843_b1 , w_42288 );
or ( w_42285 , \3843_b0 , \3844_b0 );
not ( \3844_b0 , w_42289 );
and ( w_42289 , w_42288 , \3844_b1 );
or ( \3856_b1 , \3851_b1 , w_42292 );
or ( \3856_b0 , \3851_b0 , w_42291 );
not ( w_42291 , w_42293 );
and ( w_42293 , w_42292 , w_42290 );
or ( w_42290 , \3854_b1 , w_42294 );
or ( w_42291 , \3854_b0 , \3855_b0 );
not ( \3855_b0 , w_42295 );
and ( w_42295 , w_42294 , \3855_b1 );
or ( \3876_b1 , \3869_b1 , w_42298 );
or ( \3876_b0 , \3869_b0 , w_42297 );
not ( w_42297 , w_42299 );
and ( w_42299 , w_42298 , w_42296 );
or ( w_42296 , \3874_b1 , w_42300 );
or ( w_42297 , \3874_b0 , \3875_b0 );
not ( \3875_b0 , w_42301 );
and ( w_42301 , w_42300 , \3875_b1 );
or ( \3892_b1 , \3885_b1 , w_42304 );
or ( \3892_b0 , \3885_b0 , w_42303 );
not ( w_42303 , w_42305 );
and ( w_42305 , w_42304 , w_42302 );
or ( w_42302 , \3890_b1 , w_42306 );
or ( w_42303 , \3890_b0 , \3891_b0 );
not ( \3891_b0 , w_42307 );
and ( w_42307 , w_42306 , \3891_b1 );
or ( \3909_b1 , \3902_b1 , w_42310 );
or ( \3909_b0 , \3902_b0 , w_42309 );
not ( w_42309 , w_42311 );
and ( w_42311 , w_42310 , w_42308 );
or ( w_42308 , \3907_b1 , w_42312 );
or ( w_42309 , \3907_b0 , \3908_b0 );
not ( \3908_b0 , w_42313 );
and ( w_42313 , w_42312 , \3908_b1 );
or ( \3912_b1 , \3893_b1 , w_42316 );
or ( \3912_b0 , \3893_b0 , w_42315 );
not ( w_42315 , w_42317 );
and ( w_42317 , w_42316 , w_42314 );
or ( w_42314 , \3910_b1 , w_42318 );
or ( w_42315 , \3910_b0 , \3911_b0 );
not ( \3911_b0 , w_42319 );
and ( w_42319 , w_42318 , \3911_b1 );
or ( \3922_b1 , \3917_b1 , w_42322 );
or ( \3922_b0 , \3917_b0 , w_42321 );
not ( w_42321 , w_42323 );
and ( w_42323 , w_42322 , w_42320 );
or ( w_42320 , \3920_b1 , w_42324 );
or ( w_42321 , \3920_b0 , \3921_b0 );
not ( \3921_b0 , w_42325 );
and ( w_42325 , w_42324 , \3921_b1 );
or ( \3939_b1 , \3932_b1 , w_42328 );
or ( \3939_b0 , \3932_b0 , w_42327 );
not ( w_42327 , w_42329 );
and ( w_42329 , w_42328 , w_42326 );
or ( w_42326 , \3937_b1 , w_42330 );
or ( w_42327 , \3937_b0 , \3938_b0 );
not ( \3938_b0 , w_42331 );
and ( w_42331 , w_42330 , \3938_b1 );
or ( \3947_b1 , \3942_b1 , w_42334 );
or ( \3947_b0 , \3942_b0 , w_42333 );
not ( w_42333 , w_42335 );
and ( w_42335 , w_42334 , w_42332 );
or ( w_42332 , \3945_b1 , w_42336 );
or ( w_42333 , \3945_b0 , \3946_b0 );
not ( \3946_b0 , w_42337 );
and ( w_42337 , w_42336 , \3946_b1 );
or ( \3950_b1 , \3923_b1 , w_42340 );
or ( \3950_b0 , \3923_b0 , w_42339 );
not ( w_42339 , w_42341 );
and ( w_42341 , w_42340 , w_42338 );
or ( w_42338 , \3948_b1 , w_42342 );
or ( w_42339 , \3948_b0 , \3949_b0 );
not ( \3949_b0 , w_42343 );
and ( w_42343 , w_42342 , \3949_b1 );
or ( \3960_b1 , \3955_b1 , w_42346 );
or ( \3960_b0 , \3955_b0 , w_42345 );
not ( w_42345 , w_42347 );
and ( w_42347 , w_42346 , w_42344 );
or ( w_42344 , \3958_b1 , w_42348 );
or ( w_42345 , \3958_b0 , \3959_b0 );
not ( \3959_b0 , w_42349 );
and ( w_42349 , w_42348 , \3959_b1 );
or ( \3966_b1 , \3961_b1 , w_42352 );
or ( \3966_b0 , \3961_b0 , w_42351 );
not ( w_42351 , w_42353 );
and ( w_42353 , w_42352 , w_42350 );
or ( w_42350 , \3964_b1 , w_42354 );
or ( w_42351 , \3964_b0 , \3965_b0 );
not ( \3965_b0 , w_42355 );
and ( w_42355 , w_42354 , \3965_b1 );
or ( \3973_b1 , \3969_b1 , w_42358 );
or ( \3973_b0 , \3969_b0 , w_42357 );
not ( w_42357 , w_42359 );
and ( w_42359 , w_42358 , w_42356 );
or ( w_42356 , \3971_b1 , w_42360 );
or ( w_42357 , \3971_b0 , \3972_b0 );
not ( \3972_b0 , w_42361 );
and ( w_42361 , w_42360 , \3972_b1 );
or ( \3980_b1 , \3976_b1 , w_42364 );
or ( \3980_b0 , \3976_b0 , w_42363 );
not ( w_42363 , w_42365 );
and ( w_42365 , w_42364 , w_42362 );
or ( w_42362 , \3978_b1 , w_42366 );
or ( w_42363 , \3978_b0 , \3979_b0 );
not ( \3979_b0 , w_42367 );
and ( w_42367 , w_42366 , \3979_b1 );
or ( \4000_b1 , \3993_b1 , w_42370 );
or ( \4000_b0 , \3993_b0 , w_42369 );
not ( w_42369 , w_42371 );
and ( w_42371 , w_42370 , w_42368 );
or ( w_42368 , \3998_b1 , w_42372 );
or ( w_42369 , \3998_b0 , \3999_b0 );
not ( \3999_b0 , w_42373 );
and ( w_42373 , w_42372 , \3999_b1 );
or ( \4012_b1 , \4009_b1 , w_42376 );
or ( \4012_b0 , \4009_b0 , w_42375 );
not ( w_42375 , w_42377 );
and ( w_42377 , w_42376 , w_42374 );
or ( w_42374 , \4010_b1 , w_42378 );
or ( w_42375 , \4010_b0 , \4011_b0 );
not ( \4011_b0 , w_42379 );
and ( w_42379 , w_42378 , \4011_b1 );
or ( \4029_b1 , \4022_b1 , w_42382 );
or ( \4029_b0 , \4022_b0 , w_42381 );
not ( w_42381 , w_42383 );
and ( w_42383 , w_42382 , w_42380 );
or ( w_42380 , \4027_b1 , w_42384 );
or ( w_42381 , \4027_b0 , \4028_b0 );
not ( \4028_b0 , w_42385 );
and ( w_42385 , w_42384 , \4028_b1 );
or ( \4032_b1 , \4013_b1 , w_42388 );
or ( \4032_b0 , \4013_b0 , w_42387 );
not ( w_42387 , w_42389 );
and ( w_42389 , w_42388 , w_42386 );
or ( w_42386 , \4030_b1 , w_42390 );
or ( w_42387 , \4030_b0 , \4031_b0 );
not ( \4031_b0 , w_42391 );
and ( w_42391 , w_42390 , \4031_b1 );
or ( \4048_b1 , \4041_b1 , w_42394 );
or ( \4048_b0 , \4041_b0 , w_42393 );
not ( w_42393 , w_42395 );
and ( w_42395 , w_42394 , w_42392 );
or ( w_42392 , \4046_b1 , w_42396 );
or ( w_42393 , \4046_b0 , \4047_b0 );
not ( \4047_b0 , w_42397 );
and ( w_42397 , w_42396 , \4047_b1 );
or ( \4063_b1 , \4056_b1 , w_42400 );
or ( \4063_b0 , \4056_b0 , w_42399 );
not ( w_42399 , w_42401 );
and ( w_42401 , w_42400 , w_42398 );
or ( w_42398 , \4061_b1 , w_42402 );
or ( w_42399 , \4061_b0 , \4062_b0 );
not ( \4062_b0 , w_42403 );
and ( w_42403 , w_42402 , \4062_b1 );
or ( \4074_b1 , \4069_b1 , w_42406 );
or ( \4074_b0 , \4069_b0 , w_42405 );
not ( w_42405 , w_42407 );
and ( w_42407 , w_42406 , w_42404 );
or ( w_42404 , \4072_b1 , w_42408 );
or ( w_42405 , \4072_b0 , \4073_b0 );
not ( \4073_b0 , w_42409 );
and ( w_42409 , w_42408 , \4073_b1 );
or ( \4077_b1 , \4064_b1 , w_42412 );
or ( \4077_b0 , \4064_b0 , w_42411 );
not ( w_42411 , w_42413 );
and ( w_42413 , w_42412 , w_42410 );
or ( w_42410 , \4075_b1 , w_42414 );
or ( w_42411 , \4075_b0 , \4076_b0 );
not ( \4076_b0 , w_42415 );
and ( w_42415 , w_42414 , \4076_b1 );
or ( \4087_b1 , \4082_b1 , w_42418 );
or ( \4087_b0 , \4082_b0 , w_42417 );
not ( w_42417 , w_42419 );
and ( w_42419 , w_42418 , w_42416 );
or ( w_42416 , \4085_b1 , w_42420 );
or ( w_42417 , \4085_b0 , \4086_b0 );
not ( \4086_b0 , w_42421 );
and ( w_42421 , w_42420 , \4086_b1 );
or ( \4093_b1 , \4088_b1 , w_42424 );
or ( \4093_b0 , \4088_b0 , w_42423 );
not ( w_42423 , w_42425 );
and ( w_42425 , w_42424 , w_42422 );
or ( w_42422 , \4091_b1 , w_42426 );
or ( w_42423 , \4091_b0 , \4092_b0 );
not ( \4092_b0 , w_42427 );
and ( w_42427 , w_42426 , \4092_b1 );
or ( \4103_b1 , \4098_b1 , w_42430 );
or ( \4103_b0 , \4098_b0 , w_42429 );
not ( w_42429 , w_42431 );
and ( w_42431 , w_42430 , w_42428 );
or ( w_42428 , \4101_b1 , w_42432 );
or ( w_42429 , \4101_b0 , \4102_b0 );
not ( \4102_b0 , w_42433 );
and ( w_42433 , w_42432 , \4102_b1 );
or ( \4109_b1 , \4104_b1 , w_42436 );
or ( \4109_b0 , \4104_b0 , w_42435 );
not ( w_42435 , w_42437 );
and ( w_42437 , w_42436 , w_42434 );
or ( w_42434 , \4107_b1 , w_42438 );
or ( w_42435 , \4107_b0 , \4108_b0 );
not ( \4108_b0 , w_42439 );
and ( w_42439 , w_42438 , \4108_b1 );
or ( \4120_b1 , \4115_b1 , w_42442 );
or ( \4120_b0 , \4115_b0 , w_42441 );
not ( w_42441 , w_42443 );
and ( w_42443 , w_42442 , w_42440 );
or ( w_42440 , \4118_b1 , w_42444 );
or ( w_42441 , \4118_b0 , \4119_b0 );
not ( \4119_b0 , w_42445 );
and ( w_42445 , w_42444 , \4119_b1 );
or ( \4140_b1 , \4133_b1 , w_42448 );
or ( \4140_b0 , \4133_b0 , w_42447 );
not ( w_42447 , w_42449 );
and ( w_42449 , w_42448 , w_42446 );
or ( w_42446 , \4138_b1 , w_42450 );
or ( w_42447 , \4138_b0 , \4139_b0 );
not ( \4139_b0 , w_42451 );
and ( w_42451 , w_42450 , \4139_b1 );
or ( \4156_b1 , \4149_b1 , w_42454 );
or ( \4156_b0 , \4149_b0 , w_42453 );
not ( w_42453 , w_42455 );
and ( w_42455 , w_42454 , w_42452 );
or ( w_42452 , \4154_b1 , w_42456 );
or ( w_42453 , \4154_b0 , \4155_b0 );
not ( \4155_b0 , w_42457 );
and ( w_42457 , w_42456 , \4155_b1 );
or ( \4173_b1 , \4166_b1 , w_42460 );
or ( \4173_b0 , \4166_b0 , w_42459 );
not ( w_42459 , w_42461 );
and ( w_42461 , w_42460 , w_42458 );
or ( w_42458 , \4171_b1 , w_42462 );
or ( w_42459 , \4171_b0 , \4172_b0 );
not ( \4172_b0 , w_42463 );
and ( w_42463 , w_42462 , \4172_b1 );
or ( \4176_b1 , \4157_b1 , w_42466 );
or ( \4176_b0 , \4157_b0 , w_42465 );
not ( w_42465 , w_42467 );
and ( w_42467 , w_42466 , w_42464 );
or ( w_42464 , \4174_b1 , w_42468 );
or ( w_42465 , \4174_b0 , \4175_b0 );
not ( \4175_b0 , w_42469 );
and ( w_42469 , w_42468 , \4175_b1 );
or ( \4186_b1 , \4181_b1 , w_42472 );
or ( \4186_b0 , \4181_b0 , w_42471 );
not ( w_42471 , w_42473 );
and ( w_42473 , w_42472 , w_42470 );
or ( w_42470 , \4184_b1 , w_42474 );
or ( w_42471 , \4184_b0 , \4185_b0 );
not ( \4185_b0 , w_42475 );
and ( w_42475 , w_42474 , \4185_b1 );
or ( \4203_b1 , \4196_b1 , w_42478 );
or ( \4203_b0 , \4196_b0 , w_42477 );
not ( w_42477 , w_42479 );
and ( w_42479 , w_42478 , w_42476 );
or ( w_42476 , \4201_b1 , w_42480 );
or ( w_42477 , \4201_b0 , \4202_b0 );
not ( \4202_b0 , w_42481 );
and ( w_42481 , w_42480 , \4202_b1 );
or ( \4210_b1 , \4206_b1 , w_42484 );
or ( \4210_b0 , \4206_b0 , w_42483 );
not ( w_42483 , w_42485 );
and ( w_42485 , w_42484 , w_42482 );
or ( w_42482 , \4208_b1 , w_42486 );
or ( w_42483 , \4208_b0 , \4209_b0 );
not ( \4209_b0 , w_42487 );
and ( w_42487 , w_42486 , \4209_b1 );
or ( \4213_b1 , \4187_b1 , w_42490 );
or ( \4213_b0 , \4187_b0 , w_42489 );
not ( w_42489 , w_42491 );
and ( w_42491 , w_42490 , w_42488 );
or ( w_42488 , \4211_b1 , w_42492 );
or ( w_42489 , \4211_b0 , \4212_b0 );
not ( \4212_b0 , w_42493 );
and ( w_42493 , w_42492 , \4212_b1 );
or ( \4223_b1 , \4218_b1 , w_42496 );
or ( \4223_b0 , \4218_b0 , w_42495 );
not ( w_42495 , w_42497 );
and ( w_42497 , w_42496 , w_42494 );
or ( w_42494 , \4221_b1 , w_42498 );
or ( w_42495 , \4221_b0 , \4222_b0 );
not ( \4222_b0 , w_42499 );
and ( w_42499 , w_42498 , \4222_b1 );
or ( \4229_b1 , \4224_b1 , w_42502 );
or ( \4229_b0 , \4224_b0 , w_42501 );
not ( w_42501 , w_42503 );
and ( w_42503 , w_42502 , w_42500 );
or ( w_42500 , \4227_b1 , w_42504 );
or ( w_42501 , \4227_b0 , \4228_b0 );
not ( \4228_b0 , w_42505 );
and ( w_42505 , w_42504 , \4228_b1 );
or ( \4237_b1 , \4232_b1 , w_42508 );
or ( \4237_b0 , \4232_b0 , w_42507 );
not ( w_42507 , w_42509 );
and ( w_42509 , w_42508 , w_42506 );
or ( w_42506 , \4235_b1 , w_42510 );
or ( w_42507 , \4235_b0 , \4236_b0 );
not ( \4236_b0 , w_42511 );
and ( w_42511 , w_42510 , \4236_b1 );
or ( \4244_b1 , \4240_b1 , w_42514 );
or ( \4244_b0 , \4240_b0 , w_42513 );
not ( w_42513 , w_42515 );
and ( w_42515 , w_42514 , w_42512 );
or ( w_42512 , \4242_b1 , w_42516 );
or ( w_42513 , \4242_b0 , \4243_b0 );
not ( \4243_b0 , w_42517 );
and ( w_42517 , w_42516 , \4243_b1 );
or ( \4264_b1 , \4257_b1 , w_42520 );
or ( \4264_b0 , \4257_b0 , w_42519 );
not ( w_42519 , w_42521 );
and ( w_42521 , w_42520 , w_42518 );
or ( w_42518 , \4262_b1 , w_42522 );
or ( w_42519 , \4262_b0 , \4263_b0 );
not ( \4263_b0 , w_42523 );
and ( w_42523 , w_42522 , \4263_b1 );
or ( \4280_b1 , \4273_b1 , w_42526 );
or ( \4280_b0 , \4273_b0 , w_42525 );
not ( w_42525 , w_42527 );
and ( w_42527 , w_42526 , w_42524 );
or ( w_42524 , \4278_b1 , w_42528 );
or ( w_42525 , \4278_b0 , \4279_b0 );
not ( \4279_b0 , w_42529 );
and ( w_42529 , w_42528 , \4279_b1 );
or ( \4293_b1 , \4290_b1 , w_42532 );
or ( \4293_b0 , \4290_b0 , w_42531 );
not ( w_42531 , w_42533 );
and ( w_42533 , w_42532 , w_42530 );
or ( w_42530 , \4291_b1 , w_42534 );
or ( w_42531 , \4291_b0 , \4292_b0 );
not ( \4292_b0 , w_42535 );
and ( w_42535 , w_42534 , \4292_b1 );
or ( \4296_b1 , \4281_b1 , w_42538 );
or ( \4296_b0 , \4281_b0 , w_42537 );
not ( w_42537 , w_42539 );
and ( w_42539 , w_42538 , w_42536 );
or ( w_42536 , \4294_b1 , w_42540 );
or ( w_42537 , \4294_b0 , \4295_b0 );
not ( \4295_b0 , w_42541 );
and ( w_42541 , w_42540 , \4295_b1 );
or ( \4312_b1 , \4305_b1 , w_42544 );
or ( \4312_b0 , \4305_b0 , w_42543 );
not ( w_42543 , w_42545 );
and ( w_42545 , w_42544 , w_42542 );
or ( w_42542 , \4310_b1 , w_42546 );
or ( w_42543 , \4310_b0 , \4311_b0 );
not ( \4311_b0 , w_42547 );
and ( w_42547 , w_42546 , \4311_b1 );
or ( \4320_b1 , \4315_b1 , w_42550 );
or ( \4320_b0 , \4315_b0 , w_42549 );
not ( w_42549 , w_42551 );
and ( w_42551 , w_42550 , w_42548 );
or ( w_42548 , \4318_b1 , w_42552 );
or ( w_42549 , \4318_b0 , \4319_b0 );
not ( \4319_b0 , w_42553 );
and ( w_42553 , w_42552 , \4319_b1 );
or ( \4329_b1 , \4321_b1 , w_42556 );
or ( \4329_b0 , \4321_b0 , w_42555 );
not ( w_42555 , w_42557 );
and ( w_42557 , w_42556 , w_42554 );
or ( w_42554 , \4327_b1 , w_42558 );
or ( w_42555 , \4327_b0 , \4328_b0 );
not ( \4328_b0 , w_42559 );
and ( w_42559 , w_42558 , \4328_b1 );
or ( \4339_b1 , \4334_b1 , w_42562 );
or ( \4339_b0 , \4334_b0 , w_42561 );
not ( w_42561 , w_42563 );
and ( w_42563 , w_42562 , w_42560 );
or ( w_42560 , \4337_b1 , w_42564 );
or ( w_42561 , \4337_b0 , \4338_b0 );
not ( \4338_b0 , w_42565 );
and ( w_42565 , w_42564 , \4338_b1 );
or ( \4345_b1 , \4340_b1 , w_42568 );
or ( \4345_b0 , \4340_b0 , w_42567 );
not ( w_42567 , w_42569 );
and ( w_42569 , w_42568 , w_42566 );
or ( w_42566 , \4343_b1 , w_42570 );
or ( w_42567 , \4343_b0 , \4344_b0 );
not ( \4344_b0 , w_42571 );
and ( w_42571 , w_42570 , \4344_b1 );
or ( \4356_b1 , \4351_b1 , w_42574 );
or ( \4356_b0 , \4351_b0 , w_42573 );
not ( w_42573 , w_42575 );
and ( w_42575 , w_42574 , w_42572 );
or ( w_42572 , \4354_b1 , w_42576 );
or ( w_42573 , \4354_b0 , \4355_b0 );
not ( \4355_b0 , w_42577 );
and ( w_42577 , w_42576 , \4355_b1 );
or ( \4386_b1 , \4379_b1 , w_42580 );
or ( \4386_b0 , \4379_b0 , w_42579 );
not ( w_42579 , w_42581 );
and ( w_42581 , w_42580 , w_42578 );
or ( w_42578 , \4384_b1 , w_42582 );
or ( w_42579 , \4384_b0 , \4385_b0 );
not ( \4385_b0 , w_42583 );
and ( w_42583 , w_42582 , \4385_b1 );
or ( \4402_b1 , \4395_b1 , w_42586 );
or ( \4402_b0 , \4395_b0 , w_42585 );
not ( w_42585 , w_42587 );
and ( w_42587 , w_42586 , w_42584 );
or ( w_42584 , \4400_b1 , w_42588 );
or ( w_42585 , \4400_b0 , \4401_b0 );
not ( \4401_b0 , w_42589 );
and ( w_42589 , w_42588 , \4401_b1 );
or ( \4419_b1 , \4412_b1 , w_42592 );
or ( \4419_b0 , \4412_b0 , w_42591 );
not ( w_42591 , w_42593 );
and ( w_42593 , w_42592 , w_42590 );
or ( w_42590 , \4417_b1 , w_42594 );
or ( w_42591 , \4417_b0 , \4418_b0 );
not ( \4418_b0 , w_42595 );
and ( w_42595 , w_42594 , \4418_b1 );
or ( \4422_b1 , \4403_b1 , w_42598 );
or ( \4422_b0 , \4403_b0 , w_42597 );
not ( w_42597 , w_42599 );
and ( w_42599 , w_42598 , w_42596 );
or ( w_42596 , \4420_b1 , w_42600 );
or ( w_42597 , \4420_b0 , \4421_b0 );
not ( \4421_b0 , w_42601 );
and ( w_42601 , w_42600 , \4421_b1 );
or ( \4432_b1 , \4427_b1 , w_42604 );
or ( \4432_b0 , \4427_b0 , w_42603 );
not ( w_42603 , w_42605 );
and ( w_42605 , w_42604 , w_42602 );
or ( w_42602 , \4430_b1 , w_42606 );
or ( w_42603 , \4430_b0 , \4431_b0 );
not ( \4431_b0 , w_42607 );
and ( w_42607 , w_42606 , \4431_b1 );
or ( \4441_b1 , \4433_b1 , w_42610 );
or ( \4441_b0 , \4433_b0 , w_42609 );
not ( w_42609 , w_42611 );
and ( w_42611 , w_42610 , w_42608 );
or ( w_42608 , \4439_b1 , w_42612 );
or ( w_42609 , \4439_b0 , \4440_b0 );
not ( \4440_b0 , w_42613 );
and ( w_42613 , w_42612 , \4440_b1 );
or ( \4450_b1 , \4446_b1 , w_42616 );
or ( \4450_b0 , \4446_b0 , w_42615 );
not ( w_42615 , w_42617 );
and ( w_42617 , w_42616 , w_42614 );
or ( w_42614 , \4448_b1 , w_42618 );
or ( w_42615 , \4448_b0 , \4449_b0 );
not ( \4449_b0 , w_42619 );
and ( w_42619 , w_42618 , \4449_b1 );
or ( \4456_b1 , \4451_b1 , w_42622 );
or ( \4456_b0 , \4451_b0 , w_42621 );
not ( w_42621 , w_42623 );
and ( w_42623 , w_42622 , w_42620 );
or ( w_42620 , \4454_b1 , w_42624 );
or ( w_42621 , \4454_b0 , \4455_b0 );
not ( \4455_b0 , w_42625 );
and ( w_42625 , w_42624 , \4455_b1 );
or ( \4463_b1 , \4459_b1 , w_42628 );
or ( \4463_b0 , \4459_b0 , w_42627 );
not ( w_42627 , w_42629 );
and ( w_42629 , w_42628 , w_42626 );
or ( w_42626 , \4461_b1 , w_42630 );
or ( w_42627 , \4461_b0 , \4462_b0 );
not ( \4462_b0 , w_42631 );
and ( w_42631 , w_42630 , \4462_b1 );
or ( \4481_b1 , \4476_b1 , w_42634 );
or ( \4481_b0 , \4476_b0 , w_42633 );
not ( w_42633 , w_42635 );
and ( w_42635 , w_42634 , w_42632 );
or ( w_42632 , \4479_b1 , w_42636 );
or ( w_42633 , \4479_b0 , \4480_b0 );
not ( \4480_b0 , w_42637 );
and ( w_42637 , w_42636 , \4480_b1 );
or ( \4493_b1 , \4486_b1 , w_42640 );
or ( \4493_b0 , \4486_b0 , w_42639 );
not ( w_42639 , w_42641 );
and ( w_42641 , w_42640 , w_42638 );
or ( w_42638 , \4491_b1 , w_42642 );
or ( w_42639 , \4491_b0 , \4492_b0 );
not ( \4492_b0 , w_42643 );
and ( w_42643 , w_42642 , \4492_b1 );
or ( \4505_b1 , \4502_b1 , w_42646 );
or ( \4505_b0 , \4502_b0 , w_42645 );
not ( w_42645 , w_42647 );
and ( w_42647 , w_42646 , w_42644 );
or ( w_42644 , \4503_b1 , w_42648 );
or ( w_42645 , \4503_b0 , \4504_b0 );
not ( \4504_b0 , w_42649 );
and ( w_42649 , w_42648 , \4504_b1 );
or ( \4521_b1 , \4514_b1 , w_42652 );
or ( \4521_b0 , \4514_b0 , w_42651 );
not ( w_42651 , w_42653 );
and ( w_42653 , w_42652 , w_42650 );
or ( w_42650 , \4519_b1 , w_42654 );
or ( w_42651 , \4519_b0 , \4520_b0 );
not ( \4520_b0 , w_42655 );
and ( w_42655 , w_42654 , \4520_b1 );
or ( \4538_b1 , \4531_b1 , w_42658 );
or ( \4538_b0 , \4531_b0 , w_42657 );
not ( w_42657 , w_42659 );
and ( w_42659 , w_42658 , w_42656 );
or ( w_42656 , \4536_b1 , w_42660 );
or ( w_42657 , \4536_b0 , \4537_b0 );
not ( \4537_b0 , w_42661 );
and ( w_42661 , w_42660 , \4537_b1 );
or ( \4541_b1 , \4522_b1 , w_42664 );
or ( \4541_b0 , \4522_b0 , w_42663 );
not ( w_42663 , w_42665 );
and ( w_42665 , w_42664 , w_42662 );
or ( w_42662 , \4539_b1 , w_42666 );
or ( w_42663 , \4539_b0 , \4540_b0 );
not ( \4540_b0 , w_42667 );
and ( w_42667 , w_42666 , \4540_b1 );
or ( \4552_b1 , \4547_b1 , w_42670 );
or ( \4552_b0 , \4547_b0 , w_42669 );
not ( w_42669 , w_42671 );
and ( w_42671 , w_42670 , w_42668 );
or ( w_42668 , \4550_b1 , w_42672 );
or ( w_42669 , \4550_b0 , \4551_b0 );
not ( \4551_b0 , w_42673 );
and ( w_42673 , w_42672 , \4551_b1 );
or ( \4555_b1 , \4542_b1 , w_42676 );
or ( \4555_b0 , \4542_b0 , w_42675 );
not ( w_42675 , w_42677 );
and ( w_42677 , w_42676 , w_42674 );
or ( w_42674 , \4553_b1 , w_42678 );
or ( w_42675 , \4553_b0 , \4554_b0 );
not ( \4554_b0 , w_42679 );
and ( w_42679 , w_42678 , \4554_b1 );
or ( \4564_b1 , \4560_b1 , w_42682 );
or ( \4564_b0 , \4560_b0 , w_42681 );
not ( w_42681 , w_42683 );
and ( w_42683 , w_42682 , w_42680 );
or ( w_42680 , \4562_b1 , w_42684 );
or ( w_42681 , \4562_b0 , \4563_b0 );
not ( \4563_b0 , w_42685 );
and ( w_42685 , w_42684 , \4563_b1 );
or ( \4570_b1 , \4565_b1 , w_42688 );
or ( \4570_b0 , \4565_b0 , w_42687 );
not ( w_42687 , w_42689 );
and ( w_42689 , w_42688 , w_42686 );
or ( w_42686 , \4568_b1 , w_42690 );
or ( w_42687 , \4568_b0 , \4569_b0 );
not ( \4569_b0 , w_42691 );
and ( w_42691 , w_42690 , \4569_b1 );
or ( \4578_b1 , \4573_b1 , w_42694 );
or ( \4578_b0 , \4573_b0 , w_42693 );
not ( w_42693 , w_42695 );
and ( w_42695 , w_42694 , w_42692 );
or ( w_42692 , \4576_b1 , w_42696 );
or ( w_42693 , \4576_b0 , \4577_b0 );
not ( \4577_b0 , w_42697 );
and ( w_42697 , w_42696 , \4577_b1 );
or ( \4598_b1 , \4591_b1 , w_42700 );
or ( \4598_b0 , \4591_b0 , w_42699 );
not ( w_42699 , w_42701 );
and ( w_42701 , w_42700 , w_42698 );
or ( w_42698 , \4596_b1 , w_42702 );
or ( w_42699 , \4596_b0 , \4597_b0 );
not ( \4597_b0 , w_42703 );
and ( w_42703 , w_42702 , \4597_b1 );
or ( \4614_b1 , \4607_b1 , w_42706 );
or ( \4614_b0 , \4607_b0 , w_42705 );
not ( w_42705 , w_42707 );
and ( w_42707 , w_42706 , w_42704 );
or ( w_42704 , \4612_b1 , w_42708 );
or ( w_42705 , \4612_b0 , \4613_b0 );
not ( \4613_b0 , w_42709 );
and ( w_42709 , w_42708 , \4613_b1 );
or ( \4631_b1 , \4624_b1 , w_42712 );
or ( \4631_b0 , \4624_b0 , w_42711 );
not ( w_42711 , w_42713 );
and ( w_42713 , w_42712 , w_42710 );
or ( w_42710 , \4629_b1 , w_42714 );
or ( w_42711 , \4629_b0 , \4630_b0 );
not ( \4630_b0 , w_42715 );
and ( w_42715 , w_42714 , \4630_b1 );
or ( \4634_b1 , \4615_b1 , w_42718 );
or ( \4634_b0 , \4615_b0 , w_42717 );
not ( w_42717 , w_42719 );
and ( w_42719 , w_42718 , w_42716 );
or ( w_42716 , \4632_b1 , w_42720 );
or ( w_42717 , \4632_b0 , \4633_b0 );
not ( \4633_b0 , w_42721 );
and ( w_42721 , w_42720 , \4633_b1 );
or ( \4644_b1 , \4639_b1 , w_42724 );
or ( \4644_b0 , \4639_b0 , w_42723 );
not ( w_42723 , w_42725 );
and ( w_42725 , w_42724 , w_42722 );
or ( w_42722 , \4642_b1 , w_42726 );
or ( w_42723 , \4642_b0 , \4643_b0 );
not ( \4643_b0 , w_42727 );
and ( w_42727 , w_42726 , \4643_b1 );
or ( \4650_b1 , \4645_b1 , w_42730 );
or ( \4650_b0 , \4645_b0 , w_42729 );
not ( w_42729 , w_42731 );
and ( w_42731 , w_42730 , w_42728 );
or ( w_42728 , \4648_b1 , w_42732 );
or ( w_42729 , \4648_b0 , \4649_b0 );
not ( \4649_b0 , w_42733 );
and ( w_42733 , w_42732 , \4649_b1 );
or ( \4658_b1 , \4653_b1 , w_42736 );
or ( \4658_b0 , \4653_b0 , w_42735 );
not ( w_42735 , w_42737 );
and ( w_42737 , w_42736 , w_42734 );
or ( w_42734 , \4656_b1 , w_42738 );
or ( w_42735 , \4656_b0 , \4657_b0 );
not ( \4657_b0 , w_42739 );
and ( w_42739 , w_42738 , \4657_b1 );
or ( \4666_b1 , \4661_b1 , w_42742 );
or ( \4666_b0 , \4661_b0 , w_42741 );
not ( w_42741 , w_42743 );
and ( w_42743 , w_42742 , w_42740 );
or ( w_42740 , \4664_b1 , w_42744 );
or ( w_42741 , \4664_b0 , \4665_b0 );
not ( \4665_b0 , w_42745 );
and ( w_42745 , w_42744 , \4665_b1 );
or ( \4682_b1 , \4679_b1 , w_42748 );
or ( \4682_b0 , \4679_b0 , w_42747 );
not ( w_42747 , w_42749 );
and ( w_42749 , w_42748 , w_42746 );
or ( w_42746 , \4680_b1 , w_42750 );
or ( w_42747 , \4680_b0 , \4681_b0 );
not ( \4681_b0 , w_42751 );
and ( w_42751 , w_42750 , \4681_b1 );
or ( \4698_b1 , \4691_b1 , w_42754 );
or ( \4698_b0 , \4691_b0 , w_42753 );
not ( w_42753 , w_42755 );
and ( w_42755 , w_42754 , w_42752 );
or ( w_42752 , \4696_b1 , w_42756 );
or ( w_42753 , \4696_b0 , \4697_b0 );
not ( \4697_b0 , w_42757 );
and ( w_42757 , w_42756 , \4697_b1 );
or ( \4715_b1 , \4708_b1 , w_42760 );
or ( \4715_b0 , \4708_b0 , w_42759 );
not ( w_42759 , w_42761 );
and ( w_42761 , w_42760 , w_42758 );
or ( w_42758 , \4713_b1 , w_42762 );
or ( w_42759 , \4713_b0 , \4714_b0 );
not ( \4714_b0 , w_42763 );
and ( w_42763 , w_42762 , \4714_b1 );
or ( \4718_b1 , \4699_b1 , w_42766 );
or ( \4718_b0 , \4699_b0 , w_42765 );
not ( w_42765 , w_42767 );
and ( w_42767 , w_42766 , w_42764 );
or ( w_42764 , \4716_b1 , w_42768 );
or ( w_42765 , \4716_b0 , \4717_b0 );
not ( \4717_b0 , w_42769 );
and ( w_42769 , w_42768 , \4717_b1 );
or ( \4730_b1 , \4725_b1 , w_42772 );
or ( \4730_b0 , \4725_b0 , w_42771 );
not ( w_42771 , w_42773 );
and ( w_42773 , w_42772 , w_42770 );
or ( w_42770 , \4728_b1 , w_42774 );
or ( w_42771 , \4728_b0 , \4729_b0 );
not ( \4729_b0 , w_42775 );
and ( w_42775 , w_42774 , \4729_b1 );
or ( \4736_b1 , \4731_b1 , w_42778 );
or ( \4736_b0 , \4731_b0 , w_42777 );
not ( w_42777 , w_42779 );
and ( w_42779 , w_42778 , w_42776 );
or ( w_42776 , \4734_b1 , w_42780 );
or ( w_42777 , \4734_b0 , \4735_b0 );
not ( \4735_b0 , w_42781 );
and ( w_42781 , w_42780 , \4735_b1 );
or ( \4747_b1 , \4742_b1 , w_42784 );
or ( \4747_b0 , \4742_b0 , w_42783 );
not ( w_42783 , w_42785 );
and ( w_42785 , w_42784 , w_42782 );
or ( w_42782 , \4745_b1 , w_42786 );
or ( w_42783 , \4745_b0 , \4746_b0 );
not ( \4746_b0 , w_42787 );
and ( w_42787 , w_42786 , \4746_b1 );
or ( \4758_b1 , \4753_b1 , w_42790 );
or ( \4758_b0 , \4753_b0 , w_42789 );
not ( w_42789 , w_42791 );
and ( w_42791 , w_42790 , w_42788 );
or ( w_42788 , \4756_b1 , w_42792 );
or ( w_42789 , \4756_b0 , \4757_b0 );
not ( \4757_b0 , w_42793 );
and ( w_42793 , w_42792 , \4757_b1 );
or ( \4778_b1 , \4771_b1 , w_42796 );
or ( \4778_b0 , \4771_b0 , w_42795 );
not ( w_42795 , w_42797 );
and ( w_42797 , w_42796 , w_42794 );
or ( w_42794 , \4776_b1 , w_42798 );
or ( w_42795 , \4776_b0 , \4777_b0 );
not ( \4777_b0 , w_42799 );
and ( w_42799 , w_42798 , \4777_b1 );
or ( \4794_b1 , \4787_b1 , w_42802 );
or ( \4794_b0 , \4787_b0 , w_42801 );
not ( w_42801 , w_42803 );
and ( w_42803 , w_42802 , w_42800 );
or ( w_42800 , \4792_b1 , w_42804 );
or ( w_42801 , \4792_b0 , \4793_b0 );
not ( \4793_b0 , w_42805 );
and ( w_42805 , w_42804 , \4793_b1 );
or ( \4811_b1 , \4804_b1 , w_42808 );
or ( \4811_b0 , \4804_b0 , w_42807 );
not ( w_42807 , w_42809 );
and ( w_42809 , w_42808 , w_42806 );
or ( w_42806 , \4809_b1 , w_42810 );
or ( w_42807 , \4809_b0 , \4810_b0 );
not ( \4810_b0 , w_42811 );
and ( w_42811 , w_42810 , \4810_b1 );
or ( \4814_b1 , \4795_b1 , w_42814 );
or ( \4814_b0 , \4795_b0 , w_42813 );
not ( w_42813 , w_42815 );
and ( w_42815 , w_42814 , w_42812 );
or ( w_42812 , \4812_b1 , w_42816 );
or ( w_42813 , \4812_b0 , \4813_b0 );
not ( \4813_b0 , w_42817 );
and ( w_42817 , w_42816 , \4813_b1 );
or ( \4826_b1 , \4821_b1 , w_42820 );
or ( \4826_b0 , \4821_b0 , w_42819 );
not ( w_42819 , w_42821 );
and ( w_42821 , w_42820 , w_42818 );
or ( w_42818 , \4824_b1 , w_42822 );
or ( w_42819 , \4824_b0 , \4825_b0 );
not ( \4825_b0 , w_42823 );
and ( w_42823 , w_42822 , \4825_b1 );
or ( \4832_b1 , \4827_b1 , w_42826 );
or ( \4832_b0 , \4827_b0 , w_42825 );
not ( w_42825 , w_42827 );
and ( w_42827 , w_42826 , w_42824 );
or ( w_42824 , \4830_b1 , w_42828 );
or ( w_42825 , \4830_b0 , \4831_b0 );
not ( \4831_b0 , w_42829 );
and ( w_42829 , w_42828 , \4831_b1 );
or ( \4839_b1 , \4835_b1 , w_42832 );
or ( \4839_b0 , \4835_b0 , w_42831 );
not ( w_42831 , w_42833 );
and ( w_42833 , w_42832 , w_42830 );
or ( w_42830 , \4837_b1 , w_42834 );
or ( w_42831 , \4837_b0 , \4838_b0 );
not ( \4838_b0 , w_42835 );
and ( w_42835 , w_42834 , \4838_b1 );
or ( \4846_b1 , \4842_b1 , w_42838 );
or ( \4846_b0 , \4842_b0 , w_42837 );
not ( w_42837 , w_42839 );
and ( w_42839 , w_42838 , w_42836 );
or ( w_42836 , \4844_b1 , w_42840 );
or ( w_42837 , \4844_b0 , \4845_b0 );
not ( \4845_b0 , w_42841 );
and ( w_42841 , w_42840 , \4845_b1 );
or ( \4866_b1 , \4859_b1 , w_42844 );
or ( \4866_b0 , \4859_b0 , w_42843 );
not ( w_42843 , w_42845 );
and ( w_42845 , w_42844 , w_42842 );
or ( w_42842 , \4864_b1 , w_42846 );
or ( w_42843 , \4864_b0 , \4865_b0 );
not ( \4865_b0 , w_42847 );
and ( w_42847 , w_42846 , \4865_b1 );
or ( \4878_b1 , \4875_b1 , w_42850 );
or ( \4878_b0 , \4875_b0 , w_42849 );
not ( w_42849 , w_42851 );
and ( w_42851 , w_42850 , w_42848 );
or ( w_42848 , \4876_b1 , w_42852 );
or ( w_42849 , \4876_b0 , \4877_b0 );
not ( \4877_b0 , w_42853 );
and ( w_42853 , w_42852 , \4877_b1 );
or ( \4895_b1 , \4888_b1 , w_42856 );
or ( \4895_b0 , \4888_b0 , w_42855 );
not ( w_42855 , w_42857 );
and ( w_42857 , w_42856 , w_42854 );
or ( w_42854 , \4893_b1 , w_42858 );
or ( w_42855 , \4893_b0 , \4894_b0 );
not ( \4894_b0 , w_42859 );
and ( w_42859 , w_42858 , \4894_b1 );
or ( \4898_b1 , \4879_b1 , w_42862 );
or ( \4898_b0 , \4879_b0 , w_42861 );
not ( w_42861 , w_42863 );
and ( w_42863 , w_42862 , w_42860 );
or ( w_42860 , \4896_b1 , w_42864 );
or ( w_42861 , \4896_b0 , \4897_b0 );
not ( \4897_b0 , w_42865 );
and ( w_42865 , w_42864 , \4897_b1 );
or ( \4908_b1 , \4903_b1 , w_42868 );
or ( \4908_b0 , \4903_b0 , w_42867 );
not ( w_42867 , w_42869 );
and ( w_42869 , w_42868 , w_42866 );
or ( w_42866 , \4906_b1 , w_42870 );
or ( w_42867 , \4906_b0 , \4907_b0 );
not ( \4907_b0 , w_42871 );
and ( w_42871 , w_42870 , \4907_b1 );
or ( \4914_b1 , \4909_b1 , w_42874 );
or ( \4914_b0 , \4909_b0 , w_42873 );
not ( w_42873 , w_42875 );
and ( w_42875 , w_42874 , w_42872 );
or ( w_42872 , \4912_b1 , w_42876 );
or ( w_42873 , \4912_b0 , \4913_b0 );
not ( \4913_b0 , w_42877 );
and ( w_42877 , w_42876 , \4913_b1 );
or ( \4924_b1 , \4919_b1 , w_42880 );
or ( \4924_b0 , \4919_b0 , w_42879 );
not ( w_42879 , w_42881 );
and ( w_42881 , w_42880 , w_42878 );
or ( w_42878 , \4922_b1 , w_42882 );
or ( w_42879 , \4922_b0 , \4923_b0 );
not ( \4923_b0 , w_42883 );
and ( w_42883 , w_42882 , \4923_b1 );
or ( \4930_b1 , \4925_b1 , w_42886 );
or ( \4930_b0 , \4925_b0 , w_42885 );
not ( w_42885 , w_42887 );
and ( w_42887 , w_42886 , w_42884 );
or ( w_42884 , \4928_b1 , w_42888 );
or ( w_42885 , \4928_b0 , \4929_b0 );
not ( \4929_b0 , w_42889 );
and ( w_42889 , w_42888 , \4929_b1 );
or ( \4941_b1 , \4936_b1 , w_42892 );
or ( \4941_b0 , \4936_b0 , w_42891 );
not ( w_42891 , w_42893 );
and ( w_42893 , w_42892 , w_42890 );
or ( w_42890 , \4939_b1 , w_42894 );
or ( w_42891 , \4939_b0 , \4940_b0 );
not ( \4940_b0 , w_42895 );
and ( w_42895 , w_42894 , \4940_b1 );
or ( \4961_b1 , \4954_b1 , w_42898 );
or ( \4961_b0 , \4954_b0 , w_42897 );
not ( w_42897 , w_42899 );
and ( w_42899 , w_42898 , w_42896 );
or ( w_42896 , \4959_b1 , w_42900 );
or ( w_42897 , \4959_b0 , \4960_b0 );
not ( \4960_b0 , w_42901 );
and ( w_42901 , w_42900 , \4960_b1 );
or ( \4977_b1 , \4970_b1 , w_42904 );
or ( \4977_b0 , \4970_b0 , w_42903 );
not ( w_42903 , w_42905 );
and ( w_42905 , w_42904 , w_42902 );
or ( w_42902 , \4975_b1 , w_42906 );
or ( w_42903 , \4975_b0 , \4976_b0 );
not ( \4976_b0 , w_42907 );
and ( w_42907 , w_42906 , \4976_b1 );
or ( \4990_b1 , \4978_b1 , w_42910 );
or ( \4990_b0 , \4978_b0 , w_42909 );
not ( w_42909 , w_42911 );
and ( w_42911 , w_42910 , w_42908 );
or ( w_42908 , \4988_b1 , w_42912 );
or ( w_42909 , \4988_b0 , \4989_b0 );
not ( \4989_b0 , w_42913 );
and ( w_42913 , w_42912 , \4989_b1 );
or ( \5000_b1 , \4995_b1 , w_42916 );
or ( \5000_b0 , \4995_b0 , w_42915 );
not ( w_42915 , w_42917 );
and ( w_42917 , w_42916 , w_42914 );
or ( w_42914 , \4998_b1 , w_42918 );
or ( w_42915 , \4998_b0 , \4999_b0 );
not ( \4999_b0 , w_42919 );
and ( w_42919 , w_42918 , \4999_b1 );
or ( \5006_b1 , \5001_b1 , w_42922 );
or ( \5006_b0 , \5001_b0 , w_42921 );
not ( w_42921 , w_42923 );
and ( w_42923 , w_42922 , w_42920 );
or ( w_42920 , \5004_b1 , w_42924 );
or ( w_42921 , \5004_b0 , \5005_b0 );
not ( \5005_b0 , w_42925 );
and ( w_42925 , w_42924 , \5005_b1 );
or ( \5014_b1 , \5009_b1 , w_42928 );
or ( \5014_b0 , \5009_b0 , w_42927 );
not ( w_42927 , w_42929 );
and ( w_42929 , w_42928 , w_42926 );
or ( w_42926 , \5012_b1 , w_42930 );
or ( w_42927 , \5012_b0 , \5013_b0 );
not ( \5013_b0 , w_42931 );
and ( w_42931 , w_42930 , \5013_b1 );
or ( \5021_b1 , \5017_b1 , w_42934 );
or ( \5021_b0 , \5017_b0 , w_42933 );
not ( w_42933 , w_42935 );
and ( w_42935 , w_42934 , w_42932 );
or ( w_42932 , \5019_b1 , w_42936 );
or ( w_42933 , \5019_b0 , \5020_b0 );
not ( \5020_b0 , w_42937 );
and ( w_42937 , w_42936 , \5020_b1 );
or ( \5039_b1 , \5034_b1 , w_42940 );
or ( \5039_b0 , \5034_b0 , w_42939 );
not ( w_42939 , w_42941 );
and ( w_42941 , w_42940 , w_42938 );
or ( w_42938 , \5037_b1 , w_42942 );
or ( w_42939 , \5037_b0 , \5038_b0 );
not ( \5038_b0 , w_42943 );
and ( w_42943 , w_42942 , \5038_b1 );
or ( \5051_b1 , \5048_b1 , w_42946 );
or ( \5051_b0 , \5048_b0 , w_42945 );
not ( w_42945 , w_42947 );
and ( w_42947 , w_42946 , w_42944 );
or ( w_42944 , \5049_b1 , w_42948 );
or ( w_42945 , \5049_b0 , \5050_b0 );
not ( \5050_b0 , w_42949 );
and ( w_42949 , w_42948 , \5050_b1 );
or ( \5068_b1 , \5061_b1 , w_42952 );
or ( \5068_b0 , \5061_b0 , w_42951 );
not ( w_42951 , w_42953 );
and ( w_42953 , w_42952 , w_42950 );
or ( w_42950 , \5066_b1 , w_42954 );
or ( w_42951 , \5066_b0 , \5067_b0 );
not ( \5067_b0 , w_42955 );
and ( w_42955 , w_42954 , \5067_b1 );
or ( \5071_b1 , \5052_b1 , w_42958 );
or ( \5071_b0 , \5052_b0 , w_42957 );
not ( w_42957 , w_42959 );
and ( w_42959 , w_42958 , w_42956 );
or ( w_42956 , \5069_b1 , w_42960 );
or ( w_42957 , \5069_b0 , \5070_b0 );
not ( \5070_b0 , w_42961 );
and ( w_42961 , w_42960 , \5070_b1 );
or ( \5080_b1 , \5076_b1 , w_42964 );
or ( \5080_b0 , \5076_b0 , w_42963 );
not ( w_42963 , w_42965 );
and ( w_42965 , w_42964 , w_42962 );
or ( w_42962 , \5078_b1 , w_42966 );
or ( w_42963 , \5078_b0 , \5079_b0 );
not ( \5079_b0 , w_42967 );
and ( w_42967 , w_42966 , \5079_b1 );
or ( \5086_b1 , \5081_b1 , w_42970 );
or ( \5086_b0 , \5081_b0 , w_42969 );
not ( w_42969 , w_42971 );
and ( w_42971 , w_42970 , w_42968 );
or ( w_42968 , \5084_b1 , w_42972 );
or ( w_42969 , \5084_b0 , \5085_b0 );
not ( \5085_b0 , w_42973 );
and ( w_42973 , w_42972 , \5085_b1 );
or ( \5097_b1 , \5092_b1 , w_42976 );
or ( \5097_b0 , \5092_b0 , w_42975 );
not ( w_42975 , w_42977 );
and ( w_42977 , w_42976 , w_42974 );
or ( w_42974 , \5095_b1 , w_42978 );
or ( w_42975 , \5095_b0 , \5096_b0 );
not ( \5096_b0 , w_42979 );
and ( w_42979 , w_42978 , \5096_b1 );
or ( \5127_b1 , \5120_b1 , w_42982 );
or ( \5127_b0 , \5120_b0 , w_42981 );
not ( w_42981 , w_42983 );
and ( w_42983 , w_42982 , w_42980 );
or ( w_42980 , \5125_b1 , w_42984 );
or ( w_42981 , \5125_b0 , \5126_b0 );
not ( \5126_b0 , w_42985 );
and ( w_42985 , w_42984 , \5126_b1 );
or ( \5143_b1 , \5136_b1 , w_42988 );
or ( \5143_b0 , \5136_b0 , w_42987 );
not ( w_42987 , w_42989 );
and ( w_42989 , w_42988 , w_42986 );
or ( w_42986 , \5141_b1 , w_42990 );
or ( w_42987 , \5141_b0 , \5142_b0 );
not ( \5142_b0 , w_42991 );
and ( w_42991 , w_42990 , \5142_b1 );
or ( \5149_b1 , \5144_b1 , w_42994 );
or ( \5149_b0 , \5144_b0 , w_42993 );
not ( w_42993 , w_42995 );
and ( w_42995 , w_42994 , w_42992 );
or ( w_42992 , \5147_b1 , w_42996 );
or ( w_42993 , \5147_b0 , \5148_b0 );
not ( \5148_b0 , w_42997 );
and ( w_42997 , w_42996 , \5148_b1 );
or ( \5160_b1 , \5155_b1 , w_43000 );
or ( \5160_b0 , \5155_b0 , w_42999 );
not ( w_42999 , w_43001 );
and ( w_43001 , w_43000 , w_42998 );
or ( w_42998 , \5158_b1 , w_43002 );
or ( w_42999 , \5158_b0 , \5159_b0 );
not ( \5159_b0 , w_43003 );
and ( w_43003 , w_43002 , \5159_b1 );
or ( \5167_b1 , \5163_b1 , w_43006 );
or ( \5167_b0 , \5163_b0 , w_43005 );
not ( w_43005 , w_43007 );
and ( w_43007 , w_43006 , w_43004 );
or ( w_43004 , \5165_b1 , w_43008 );
or ( w_43005 , \5165_b0 , \5166_b0 );
not ( \5166_b0 , w_43009 );
and ( w_43009 , w_43008 , \5166_b1 );
or ( \5183_b1 , \5180_b1 , w_43012 );
or ( \5183_b0 , \5180_b0 , w_43011 );
not ( w_43011 , w_43013 );
and ( w_43013 , w_43012 , w_43010 );
or ( w_43010 , \5181_b1 , w_43014 );
or ( w_43011 , \5181_b0 , \5182_b0 );
not ( \5182_b0 , w_43015 );
and ( w_43015 , w_43014 , \5182_b1 );
or ( \5199_b1 , \5192_b1 , w_43018 );
or ( \5199_b0 , \5192_b0 , w_43017 );
not ( w_43017 , w_43019 );
and ( w_43019 , w_43018 , w_43016 );
or ( w_43016 , \5197_b1 , w_43020 );
or ( w_43017 , \5197_b0 , \5198_b0 );
not ( \5198_b0 , w_43021 );
and ( w_43021 , w_43020 , \5198_b1 );
or ( \5207_b1 , \5200_b1 , w_43024 );
or ( \5207_b0 , \5200_b0 , w_43023 );
not ( w_43023 , w_43025 );
and ( w_43025 , w_43024 , w_43022 );
or ( w_43022 , \5205_b1 , w_43026 );
or ( w_43023 , \5205_b0 , \5206_b0 );
not ( \5206_b0 , w_43027 );
and ( w_43027 , w_43026 , \5206_b1 );
or ( \5214_b1 , \5210_b1 , w_43030 );
or ( \5214_b0 , \5210_b0 , w_43029 );
not ( w_43029 , w_43031 );
and ( w_43031 , w_43030 , w_43028 );
or ( w_43028 , \5212_b1 , w_43032 );
or ( w_43029 , \5212_b0 , \5213_b0 );
not ( \5213_b0 , w_43033 );
and ( w_43033 , w_43032 , \5213_b1 );
or ( \5222_b1 , \5217_b1 , w_43036 );
or ( \5222_b0 , \5217_b0 , w_43035 );
not ( w_43035 , w_43037 );
and ( w_43037 , w_43036 , w_43034 );
or ( w_43034 , \5220_b1 , w_43038 );
or ( w_43035 , \5220_b0 , \5221_b0 );
not ( \5221_b0 , w_43039 );
and ( w_43039 , w_43038 , \5221_b1 );
or ( \5242_b1 , \5235_b1 , w_43042 );
or ( \5242_b0 , \5235_b0 , w_43041 );
not ( w_43041 , w_43043 );
and ( w_43043 , w_43042 , w_43040 );
or ( w_43040 , \5240_b1 , w_43044 );
or ( w_43041 , \5240_b0 , \5241_b0 );
not ( \5241_b0 , w_43045 );
and ( w_43045 , w_43044 , \5241_b1 );
or ( \5258_b1 , \5251_b1 , w_43048 );
or ( \5258_b0 , \5251_b0 , w_43047 );
not ( w_43047 , w_43049 );
and ( w_43049 , w_43048 , w_43046 );
or ( w_43046 , \5256_b1 , w_43050 );
or ( w_43047 , \5256_b0 , \5257_b0 );
not ( \5257_b0 , w_43051 );
and ( w_43051 , w_43050 , \5257_b1 );
or ( \5266_b1 , \5259_b1 , w_43054 );
or ( \5266_b0 , \5259_b0 , w_43053 );
not ( w_43053 , w_43055 );
and ( w_43055 , w_43054 , w_43052 );
or ( w_43052 , \5264_b1 , w_43056 );
or ( w_43053 , \5264_b0 , \5265_b0 );
not ( \5265_b0 , w_43057 );
and ( w_43057 , w_43056 , \5265_b1 );
or ( \5276_b1 , \5271_b1 , w_43060 );
or ( \5276_b0 , \5271_b0 , w_43059 );
not ( w_43059 , w_43061 );
and ( w_43061 , w_43060 , w_43058 );
or ( w_43058 , \5274_b1 , w_43062 );
or ( w_43059 , \5274_b0 , \5275_b0 );
not ( \5275_b0 , w_43063 );
and ( w_43063 , w_43062 , \5275_b1 );
or ( \5282_b1 , \5277_b1 , w_43066 );
or ( \5282_b0 , \5277_b0 , w_43065 );
not ( w_43065 , w_43067 );
and ( w_43067 , w_43066 , w_43064 );
or ( w_43064 , \5280_b1 , w_43068 );
or ( w_43065 , \5280_b0 , \5281_b0 );
not ( \5281_b0 , w_43069 );
and ( w_43069 , w_43068 , \5281_b1 );
or ( \5293_b1 , \5288_b1 , w_43072 );
or ( \5293_b0 , \5288_b0 , w_43071 );
not ( w_43071 , w_43073 );
and ( w_43073 , w_43072 , w_43070 );
or ( w_43070 , \5291_b1 , w_43074 );
or ( w_43071 , \5291_b0 , \5292_b0 );
not ( \5292_b0 , w_43075 );
and ( w_43075 , w_43074 , \5292_b1 );
or ( \5313_b1 , \5306_b1 , w_43078 );
or ( \5313_b0 , \5306_b0 , w_43077 );
not ( w_43077 , w_43079 );
and ( w_43079 , w_43078 , w_43076 );
or ( w_43076 , \5311_b1 , w_43080 );
or ( w_43077 , \5311_b0 , \5312_b0 );
not ( \5312_b0 , w_43081 );
and ( w_43081 , w_43080 , \5312_b1 );
or ( \5325_b1 , \5322_b1 , w_43084 );
or ( \5325_b0 , \5322_b0 , w_43083 );
not ( w_43083 , w_43085 );
and ( w_43085 , w_43084 , w_43082 );
or ( w_43082 , \5323_b1 , w_43086 );
or ( w_43083 , \5323_b0 , \5324_b0 );
not ( \5324_b0 , w_43087 );
and ( w_43087 , w_43086 , \5324_b1 );
or ( \5331_b1 , \5326_b1 , w_43090 );
or ( \5331_b0 , \5326_b0 , w_43089 );
not ( w_43089 , w_43091 );
and ( w_43091 , w_43090 , w_43088 );
or ( w_43088 , \5329_b1 , w_43092 );
or ( w_43089 , \5329_b0 , \5330_b0 );
not ( \5330_b0 , w_43093 );
and ( w_43093 , w_43092 , \5330_b1 );
or ( \5339_b1 , \5334_b1 , w_43096 );
or ( \5339_b0 , \5334_b0 , w_43095 );
not ( w_43095 , w_43097 );
and ( w_43097 , w_43096 , w_43094 );
or ( w_43094 , \5337_b1 , w_43098 );
or ( w_43095 , \5337_b0 , \5338_b0 );
not ( \5338_b0 , w_43099 );
and ( w_43099 , w_43098 , \5338_b1 );
or ( \5346_b1 , \5342_b1 , w_43102 );
or ( \5346_b0 , \5342_b0 , w_43101 );
not ( w_43101 , w_43103 );
and ( w_43103 , w_43102 , w_43100 );
or ( w_43100 , \5344_b1 , w_43104 );
or ( w_43101 , \5344_b0 , \5345_b0 );
not ( \5345_b0 , w_43105 );
and ( w_43105 , w_43104 , \5345_b1 );
or ( \5366_b1 , \5359_b1 , w_43108 );
or ( \5366_b0 , \5359_b0 , w_43107 );
not ( w_43107 , w_43109 );
and ( w_43109 , w_43108 , w_43106 );
or ( w_43106 , \5364_b1 , w_43110 );
or ( w_43107 , \5364_b0 , \5365_b0 );
not ( \5365_b0 , w_43111 );
and ( w_43111 , w_43110 , \5365_b1 );
or ( \5374_b1 , \5369_b1 , w_43114 );
or ( \5374_b0 , \5369_b0 , w_43113 );
not ( w_43113 , w_43115 );
and ( w_43115 , w_43114 , w_43112 );
or ( w_43112 , \5372_b1 , w_43116 );
or ( w_43113 , \5372_b0 , \5373_b0 );
not ( \5373_b0 , w_43117 );
and ( w_43117 , w_43116 , \5373_b1 );
or ( \5382_b1 , \5377_b1 , w_43120 );
or ( \5382_b0 , \5377_b0 , w_43119 );
not ( w_43119 , w_43121 );
and ( w_43121 , w_43120 , w_43118 );
or ( w_43118 , \5380_b1 , w_43122 );
or ( w_43119 , \5380_b0 , \5381_b0 );
not ( \5381_b0 , w_43123 );
and ( w_43123 , w_43122 , \5381_b1 );
or ( \5402_b1 , \5397_b1 , w_43126 );
or ( \5402_b0 , \5397_b0 , w_43125 );
not ( w_43125 , w_43127 );
and ( w_43127 , w_43126 , w_43124 );
or ( w_43124 , \5400_b1 , w_43128 );
or ( w_43125 , \5400_b0 , \5401_b0 );
not ( \5401_b0 , w_43129 );
and ( w_43129 , w_43128 , \5401_b1 );
or ( \5414_b1 , \5411_b1 , w_43132 );
or ( \5414_b0 , \5411_b0 , w_43131 );
not ( w_43131 , w_43133 );
and ( w_43133 , w_43132 , w_43130 );
or ( w_43130 , \5412_b1 , w_43134 );
or ( w_43131 , \5412_b0 , \5413_b0 );
not ( \5413_b0 , w_43135 );
and ( w_43135 , w_43134 , \5413_b1 );
or ( \5422_b1 , \5415_b1 , w_43138 );
or ( \5422_b0 , \5415_b0 , w_43137 );
not ( w_43137 , w_43139 );
and ( w_43139 , w_43138 , w_43136 );
or ( w_43136 , \5420_b1 , w_43140 );
or ( w_43137 , \5420_b0 , \5421_b0 );
not ( \5421_b0 , w_43141 );
and ( w_43141 , w_43140 , \5421_b1 );
or ( \5435_b1 , \5430_b1 , w_43144 );
or ( \5435_b0 , \5430_b0 , w_43143 );
not ( w_43143 , w_43145 );
and ( w_43145 , w_43144 , w_43142 );
or ( w_43142 , \5433_b1 , w_43146 );
or ( w_43143 , \5433_b0 , \5434_b0 );
not ( \5434_b0 , w_43147 );
and ( w_43147 , w_43146 , \5434_b1 );
or ( \5465_b1 , \5458_b1 , w_43150 );
or ( \5465_b0 , \5458_b0 , w_43149 );
not ( w_43149 , w_43151 );
and ( w_43151 , w_43150 , w_43148 );
or ( w_43148 , \5463_b1 , w_43152 );
or ( w_43149 , \5463_b0 , \5464_b0 );
not ( \5464_b0 , w_43153 );
and ( w_43153 , w_43152 , \5464_b1 );
or ( \5473_b1 , \5468_b1 , w_43156 );
or ( \5473_b0 , \5468_b0 , w_43155 );
not ( w_43155 , w_43157 );
and ( w_43157 , w_43156 , w_43154 );
or ( w_43154 , \5471_b1 , w_43158 );
or ( w_43155 , \5471_b0 , \5472_b0 );
not ( \5472_b0 , w_43159 );
and ( w_43159 , w_43158 , \5472_b1 );
or ( \5480_b1 , \5476_b1 , w_43162 );
or ( \5480_b0 , \5476_b0 , w_43161 );
not ( w_43161 , w_43163 );
and ( w_43163 , w_43162 , w_43160 );
or ( w_43160 , \5478_b1 , w_43164 );
or ( w_43161 , \5478_b0 , \5479_b0 );
not ( \5479_b0 , w_43165 );
and ( w_43165 , w_43164 , \5479_b1 );
or ( \5496_b1 , \5493_b1 , w_43168 );
or ( \5496_b0 , \5493_b0 , w_43167 );
not ( w_43167 , w_43169 );
and ( w_43169 , w_43168 , w_43166 );
or ( w_43166 , \5494_b1 , w_43170 );
or ( w_43167 , \5494_b0 , \5495_b0 );
not ( \5495_b0 , w_43171 );
and ( w_43171 , w_43170 , \5495_b1 );
or ( \5511_b1 , \5504_b1 , w_43174 );
or ( \5511_b0 , \5504_b0 , w_43173 );
not ( w_43173 , w_43175 );
and ( w_43175 , w_43174 , w_43172 );
or ( w_43172 , \5509_b1 , w_43176 );
or ( w_43173 , \5509_b0 , \5510_b0 );
not ( \5510_b0 , w_43177 );
and ( w_43177 , w_43176 , \5510_b1 );
or ( \5541_b1 , \5534_b1 , w_43180 );
or ( \5541_b0 , \5534_b0 , w_43179 );
not ( w_43179 , w_43181 );
and ( w_43181 , w_43180 , w_43178 );
or ( w_43178 , \5539_b1 , w_43182 );
or ( w_43179 , \5539_b0 , \5540_b0 );
not ( \5540_b0 , w_43183 );
and ( w_43183 , w_43182 , \5540_b1 );
or ( \5548_b1 , \5544_b1 , w_43186 );
or ( \5548_b0 , \5544_b0 , w_43185 );
not ( w_43185 , w_43187 );
and ( w_43187 , w_43186 , w_43184 );
or ( w_43184 , \5546_b1 , w_43188 );
or ( w_43185 , \5546_b0 , \5547_b0 );
not ( \5547_b0 , w_43189 );
and ( w_43189 , w_43188 , \5547_b1 );
or ( \5564_b1 , \5561_b1 , w_43192 );
or ( \5564_b0 , \5561_b0 , w_43191 );
not ( w_43191 , w_43193 );
and ( w_43193 , w_43192 , w_43190 );
or ( w_43190 , \5562_b1 , w_43194 );
or ( w_43191 , \5562_b0 , \5563_b0 );
not ( \5563_b0 , w_43195 );
and ( w_43195 , w_43194 , \5563_b1 );
or ( \5779_b1 , \5757_b1 , w_43198 );
or ( \5779_b0 , \5757_b0 , w_43197 );
not ( w_43197 , w_43199 );
and ( w_43199 , w_43198 , w_43196 );
or ( w_43196 , \5777_b1 , w_43200 );
or ( w_43197 , \5777_b0 , \5778_b0 );
not ( \5778_b0 , w_43201 );
and ( w_43201 , w_43200 , \5778_b1 );
or ( \5840_b1 , \5818_b1 , w_43204 );
or ( \5840_b0 , \5818_b0 , w_43203 );
not ( w_43203 , w_43205 );
and ( w_43205 , w_43204 , w_43202 );
or ( w_43202 , \5838_b1 , w_43206 );
or ( w_43203 , \5838_b0 , \5839_b0 );
not ( \5839_b0 , w_43207 );
and ( w_43207 , w_43206 , \5839_b1 );
or ( \5902_b1 , \5880_b1 , w_43210 );
or ( \5902_b0 , \5880_b0 , w_43209 );
not ( w_43209 , w_43211 );
and ( w_43211 , w_43210 , w_43208 );
or ( w_43208 , \5900_b1 , w_43212 );
or ( w_43209 , \5900_b0 , \5901_b0 );
not ( \5901_b0 , w_43213 );
and ( w_43213 , w_43212 , \5901_b1 );
or ( \5905_b1 , \5841_b1 , w_43216 );
or ( \5905_b0 , \5841_b0 , w_43215 );
not ( w_43215 , w_43217 );
and ( w_43217 , w_43216 , w_43214 );
or ( w_43214 , \5903_b1 , w_43218 );
or ( w_43215 , \5903_b0 , \5904_b0 );
not ( \5904_b0 , w_43219 );
and ( w_43219 , w_43218 , \5904_b1 );
or ( \5966_b1 , \5944_b1 , w_43222 );
or ( \5966_b0 , \5944_b0 , w_43221 );
not ( w_43221 , w_43223 );
and ( w_43223 , w_43222 , w_43220 );
or ( w_43220 , \5964_b1 , w_43224 );
or ( w_43221 , \5964_b0 , \5965_b0 );
not ( \5965_b0 , w_43225 );
and ( w_43225 , w_43224 , \5965_b1 );
or ( \6027_b1 , \6005_b1 , w_43228 );
or ( \6027_b0 , \6005_b0 , w_43227 );
not ( w_43227 , w_43229 );
and ( w_43229 , w_43228 , w_43226 );
or ( w_43226 , \6025_b1 , w_43230 );
or ( w_43227 , \6025_b0 , \6026_b0 );
not ( \6026_b0 , w_43231 );
and ( w_43231 , w_43230 , \6026_b1 );
or ( \6071_b1 , \6064_b1 , w_43234 );
or ( \6071_b0 , \6064_b0 , w_43233 );
not ( w_43233 , w_43235 );
and ( w_43235 , w_43234 , w_43232 );
or ( w_43232 , \6069_b1 , w_43236 );
or ( w_43233 , \6069_b0 , \6070_b0 );
not ( \6070_b0 , w_43237 );
and ( w_43237 , w_43236 , \6070_b1 );
or ( \6074_b1 , \6028_b1 , w_43240 );
or ( \6074_b0 , \6028_b0 , w_43239 );
not ( w_43239 , w_43241 );
and ( w_43241 , w_43240 , w_43238 );
or ( w_43238 , \6072_b1 , w_43242 );
or ( w_43239 , \6072_b0 , \6073_b0 );
not ( \6073_b0 , w_43243 );
and ( w_43243 , w_43242 , \6073_b1 );
or ( \6119_b1 , \6102_b1 , w_43246 );
or ( \6119_b0 , \6102_b0 , w_43245 );
not ( w_43245 , w_43247 );
and ( w_43247 , w_43246 , w_43244 );
or ( w_43244 , \6117_b1 , w_43248 );
or ( w_43245 , \6117_b0 , \6118_b0 );
not ( \6118_b0 , w_43249 );
and ( w_43249 , w_43248 , \6118_b1 );
or ( \6122_b1 , \6075_b1 , w_43252 );
or ( \6122_b0 , \6075_b0 , w_43251 );
not ( w_43251 , w_43253 );
and ( w_43253 , w_43252 , w_43250 );
or ( w_43250 , \6120_b1 , w_43254 );
or ( w_43251 , \6120_b0 , \6121_b0 );
not ( \6121_b0 , w_43255 );
and ( w_43255 , w_43254 , \6121_b1 );
or ( \6165_b1 , \6151_b1 , w_43258 );
or ( \6165_b0 , \6151_b0 , w_43257 );
not ( w_43257 , w_43259 );
and ( w_43259 , w_43258 , w_43256 );
or ( w_43256 , \6163_b1 , w_43260 );
or ( w_43257 , \6163_b0 , \6164_b0 );
not ( \6164_b0 , w_43261 );
and ( w_43261 , w_43260 , \6164_b1 );
or ( \6177_b1 , \6173_b1 , w_43264 );
or ( \6177_b0 , \6173_b0 , w_43263 );
not ( w_43263 , w_43265 );
and ( w_43265 , w_43264 , w_43262 );
or ( w_43262 , \6175_b1 , w_43266 );
or ( w_43263 , \6175_b0 , \6176_b0 );
not ( \6176_b0 , w_43267 );
and ( w_43267 , w_43266 , \6176_b1 );
or ( \6181_b1 , \6178_b1 , w_43270 );
or ( \6181_b0 , \6178_b0 , w_43269 );
not ( w_43269 , w_43271 );
and ( w_43271 , w_43270 , w_43268 );
or ( w_43268 , \6179_b1 , w_43272 );
or ( w_43269 , \6179_b0 , \6180_b0 );
not ( \6180_b0 , w_43273 );
and ( w_43273 , w_43272 , \6180_b1 );
or ( \6198_b1 , \6195_b1 , w_43276 );
or ( \6198_b0 , \6195_b0 , w_43275 );
not ( w_43275 , w_43277 );
and ( w_43277 , w_43276 , w_43274 );
or ( w_43274 , \6196_b1 , w_43278 );
or ( w_43275 , \6196_b0 , \6197_b0 );
not ( \6197_b0 , w_43279 );
and ( w_43279 , w_43278 , \6197_b1 );
or ( \6202_b1 , \6199_b1 , w_43282 );
or ( \6202_b0 , \6199_b0 , w_43281 );
not ( w_43281 , w_43283 );
and ( w_43283 , w_43282 , w_43280 );
or ( w_43280 , \6200_b1 , w_43284 );
or ( w_43281 , \6200_b0 , \6201_b0 );
not ( \6201_b0 , w_43285 );
and ( w_43285 , w_43284 , \6201_b1 );
or ( \6207_b1 , \6203_b1 , w_43288 );
or ( \6207_b0 , \6203_b0 , w_43287 );
not ( w_43287 , w_43289 );
and ( w_43289 , w_43288 , w_43286 );
or ( w_43286 , \6205_b1 , w_43290 );
or ( w_43287 , \6205_b0 , \6206_b0 );
not ( \6206_b0 , w_43291 );
and ( w_43291 , w_43290 , \6206_b1 );
or ( \6284_b1 , \6237_b1 , w_43294 );
or ( \6284_b0 , \6237_b0 , w_43293 );
not ( w_43293 , w_43295 );
and ( w_43295 , w_43294 , w_43292 );
or ( w_43292 , \6282_b1 , w_43296 );
or ( w_43293 , \6282_b0 , \6283_b0 );
not ( \6283_b0 , w_43297 );
and ( w_43297 , w_43296 , \6283_b1 );
or ( \6317_b1 , \6314_b1 , w_43300 );
or ( \6317_b0 , \6314_b0 , w_43299 );
not ( w_43299 , w_43301 );
and ( w_43301 , w_43300 , w_43298 );
or ( w_43298 , \6315_b1 , w_43302 );
or ( w_43299 , \6315_b0 , \6316_b0 );
not ( \6316_b0 , w_43303 );
and ( w_43303 , w_43302 , \6316_b1 );
or ( \6321_b1 , \6318_b1 , w_43306 );
or ( \6321_b0 , \6318_b0 , w_43305 );
not ( w_43305 , w_43307 );
and ( w_43307 , w_43306 , w_43304 );
or ( w_43304 , \6319_b1 , w_43308 );
or ( w_43305 , \6319_b0 , \6320_b0 );
not ( \6320_b0 , w_43309 );
and ( w_43309 , w_43308 , \6320_b1 );
or ( \6329_b1 , \6326_b1 , w_43312 );
or ( \6329_b0 , \6326_b0 , w_43311 );
not ( w_43311 , w_43313 );
and ( w_43313 , w_43312 , w_43310 );
or ( w_43310 , \6327_b1 , w_43314 );
or ( w_43311 , \6327_b0 , \6328_b0 );
not ( \6328_b0 , w_43315 );
and ( w_43315 , w_43314 , \6328_b1 );
or ( \6333_b1 , \6330_b1 , w_43318 );
or ( \6333_b0 , \6330_b0 , w_43317 );
not ( w_43317 , w_43319 );
and ( w_43319 , w_43318 , w_43316 );
or ( w_43316 , \6331_b1 , w_43320 );
or ( w_43317 , \6331_b0 , \6332_b0 );
not ( \6332_b0 , w_43321 );
and ( w_43321 , w_43320 , \6332_b1 );
or ( \6338_b1 , \6335_b1 , w_43324 );
or ( \6338_b0 , \6335_b0 , w_43323 );
not ( w_43323 , w_43325 );
and ( w_43325 , w_43324 , w_43322 );
or ( w_43322 , \6336_b1 , w_43326 );
or ( w_43323 , \6336_b0 , \6337_b0 );
not ( \6337_b0 , w_43327 );
and ( w_43327 , w_43326 , \6337_b1 );
or ( \6342_b1 , \6325_b1 , w_43330 );
or ( \6342_b0 , \6325_b0 , w_43329 );
not ( w_43329 , w_43331 );
and ( w_43331 , w_43330 , w_43328 );
or ( w_43328 , \6340_b1 , w_43332 );
or ( w_43329 , \6340_b0 , \6341_b0 );
not ( \6341_b0 , w_43333 );
and ( w_43333 , w_43332 , \6341_b1 );
or ( \6345_b1 , \6285_b1 , w_43336 );
or ( \6345_b0 , \6285_b0 , w_43335 );
not ( w_43335 , w_43337 );
and ( w_43337 , w_43336 , w_43334 );
or ( w_43334 , \6343_b1 , w_43338 );
or ( w_43335 , \6343_b0 , \6344_b0 );
not ( \6344_b0 , w_43339 );
and ( w_43339 , w_43338 , \6344_b1 );
or ( \6349_b1 , \6346_b1 , w_43342 );
or ( \6349_b0 , \6346_b0 , w_43341 );
not ( w_43341 , w_43343 );
and ( w_43343 , w_43342 , w_43340 );
or ( w_43340 , \6347_b1 , w_43344 );
or ( w_43341 , \6347_b0 , \6348_b0 );
not ( \6348_b0 , w_43345 );
and ( w_43345 , w_43344 , \6348_b1 );
or ( \6353_b1 , \6350_b1 , w_43348 );
or ( \6353_b0 , \6350_b0 , w_43347 );
not ( w_43347 , w_43349 );
and ( w_43349 , w_43348 , w_43346 );
or ( w_43346 , \6351_b1 , w_43350 );
or ( w_43347 , \6351_b0 , \6352_b0 );
not ( \6352_b0 , w_43351 );
and ( w_43351 , w_43350 , \6352_b1 );
or ( \6358_b1 , \6355_b1 , w_43354 );
or ( \6358_b0 , \6355_b0 , w_43353 );
not ( w_43353 , w_43355 );
and ( w_43355 , w_43354 , w_43352 );
or ( w_43352 , \6356_b1 , w_43356 );
or ( w_43353 , \6356_b0 , \6357_b0 );
not ( \6357_b0 , w_43357 );
and ( w_43357 , w_43356 , \6357_b1 );
or ( \6363_b1 , \6360_b1 , w_43360 );
or ( \6363_b0 , \6360_b0 , w_43359 );
not ( w_43359 , w_43361 );
and ( w_43361 , w_43360 , w_43358 );
or ( w_43358 , \6361_b1 , w_43362 );
or ( w_43359 , \6361_b0 , \6362_b0 );
not ( \6362_b0 , w_43363 );
and ( w_43363 , w_43362 , \6362_b1 );
or ( \6367_b1 , \6364_b1 , w_43366 );
or ( \6367_b0 , \6364_b0 , w_43365 );
not ( w_43365 , w_43367 );
and ( w_43367 , w_43366 , w_43364 );
or ( w_43364 , \6365_b1 , w_43368 );
or ( w_43365 , \6365_b0 , \6366_b0 );
not ( \6366_b0 , w_43369 );
and ( w_43369 , w_43368 , \6366_b1 );
or ( \6372_b1 , \6369_b1 , w_43372 );
or ( \6372_b0 , \6369_b0 , w_43371 );
not ( w_43371 , w_43373 );
and ( w_43373 , w_43372 , w_43370 );
or ( w_43370 , \6370_b1 , w_43374 );
or ( w_43371 , \6370_b0 , \6371_b0 );
not ( \6371_b0 , w_43375 );
and ( w_43375 , w_43374 , \6371_b1 );
or ( \6378_b1 , \6375_b1 , w_43378 );
or ( \6378_b0 , \6375_b0 , w_43377 );
not ( w_43377 , w_43379 );
and ( w_43379 , w_43378 , w_43376 );
or ( w_43376 , \6376_b1 , w_43380 );
or ( w_43377 , \6376_b0 , \6377_b0 );
not ( \6377_b0 , w_43381 );
and ( w_43381 , w_43380 , \6377_b1 );
or ( \6468_b1 , \6465_b1 , w_43384 );
or ( \6468_b0 , \6465_b0 , w_43383 );
not ( w_43383 , w_43385 );
and ( w_43385 , w_43384 , w_43382 );
or ( w_43382 , \6466_b1 , w_43386 );
or ( w_43383 , \6466_b0 , \6467_b0 );
not ( \6467_b0 , w_43387 );
and ( w_43387 , w_43386 , \6467_b1 );
or ( \6472_b1 , \6469_b1 , w_43390 );
or ( \6472_b0 , \6469_b0 , w_43389 );
not ( w_43389 , w_43391 );
and ( w_43391 , w_43390 , w_43388 );
or ( w_43388 , \6470_b1 , w_43392 );
or ( w_43389 , \6470_b0 , \6471_b0 );
not ( \6471_b0 , w_43393 );
and ( w_43393 , w_43392 , \6471_b1 );
or ( \6478_b1 , \6464_b1 , w_43396 );
or ( \6478_b0 , \6464_b0 , w_43395 );
not ( w_43395 , w_43397 );
and ( w_43397 , w_43396 , w_43394 );
or ( w_43394 , \6476_b1 , w_43398 );
or ( w_43395 , \6476_b0 , \6477_b0 );
not ( \6477_b0 , w_43399 );
and ( w_43399 , w_43398 , \6477_b1 );
or ( \6492_b1 , \6489_b1 , w_43402 );
or ( \6492_b0 , \6489_b0 , w_43401 );
not ( w_43401 , w_43403 );
and ( w_43403 , w_43402 , w_43400 );
or ( w_43400 , \6490_b1 , w_43404 );
or ( w_43401 , \6490_b0 , \6491_b0 );
not ( \6491_b0 , w_43405 );
and ( w_43405 , w_43404 , \6491_b1 );
or ( \6502_b1 , \6499_b1 , w_43408 );
or ( \6502_b0 , \6499_b0 , w_43407 );
not ( w_43407 , w_43409 );
and ( w_43409 , w_43408 , w_43406 );
or ( w_43406 , \6500_b1 , w_43410 );
or ( w_43407 , \6500_b0 , \6501_b0 );
not ( \6501_b0 , w_43411 );
and ( w_43411 , w_43410 , \6501_b1 );
or ( \6548_b1 , \6545_b1 , w_43414 );
or ( \6548_b0 , \6545_b0 , w_43413 );
not ( w_43413 , w_43415 );
and ( w_43415 , w_43414 , w_43412 );
or ( w_43412 , \6546_b1 , w_43416 );
or ( w_43413 , \6546_b0 , \6547_b0 );
not ( \6547_b0 , w_43417 );
and ( w_43417 , w_43416 , \6547_b1 );
or ( \6552_b1 , \6549_b1 , w_43420 );
or ( \6552_b0 , \6549_b0 , w_43419 );
not ( w_43419 , w_43421 );
and ( w_43421 , w_43420 , w_43418 );
or ( w_43418 , \6550_b1 , w_43422 );
or ( w_43419 , \6550_b0 , \6551_b0 );
not ( \6551_b0 , w_43423 );
and ( w_43423 , w_43422 , \6551_b1 );
or ( \6560_b1 , \6557_b1 , w_43426 );
or ( \6560_b0 , \6557_b0 , w_43425 );
not ( w_43425 , w_43427 );
and ( w_43427 , w_43426 , w_43424 );
or ( w_43424 , \6558_b1 , w_43428 );
or ( w_43425 , \6558_b0 , \6559_b0 );
not ( \6559_b0 , w_43429 );
and ( w_43429 , w_43428 , \6559_b1 );
or ( \6564_b1 , \6561_b1 , w_43432 );
or ( \6564_b0 , \6561_b0 , w_43431 );
not ( w_43431 , w_43433 );
and ( w_43433 , w_43432 , w_43430 );
or ( w_43430 , \6562_b1 , w_43434 );
or ( w_43431 , \6562_b0 , \6563_b0 );
not ( \6563_b0 , w_43435 );
and ( w_43435 , w_43434 , \6563_b1 );
or ( \6569_b1 , \6566_b1 , w_43438 );
or ( \6569_b0 , \6566_b0 , w_43437 );
not ( w_43437 , w_43439 );
and ( w_43439 , w_43438 , w_43436 );
or ( w_43436 , \6567_b1 , w_43440 );
or ( w_43437 , \6567_b0 , \6568_b0 );
not ( \6568_b0 , w_43441 );
and ( w_43441 , w_43440 , \6568_b1 );
or ( \6575_b1 , \6572_b1 , w_43444 );
or ( \6575_b0 , \6572_b0 , w_43443 );
not ( w_43443 , w_43445 );
and ( w_43445 , w_43444 , w_43442 );
or ( w_43442 , \6573_b1 , w_43446 );
or ( w_43443 , \6573_b0 , \6574_b0 );
not ( \6574_b0 , w_43447 );
and ( w_43447 , w_43446 , \6574_b1 );
or ( \6635_b1 , \6632_b1 , w_43450 );
or ( \6635_b0 , \6632_b0 , w_43449 );
not ( w_43449 , w_43451 );
and ( w_43451 , w_43450 , w_43448 );
or ( w_43448 , \6633_b1 , w_43452 );
or ( w_43449 , \6633_b0 , \6634_b0 );
not ( \6634_b0 , w_43453 );
and ( w_43453 , w_43452 , \6634_b1 );
or ( \6639_b1 , \6636_b1 , w_43456 );
or ( \6639_b0 , \6636_b0 , w_43455 );
not ( w_43455 , w_43457 );
and ( w_43457 , w_43456 , w_43454 );
or ( w_43454 , \6637_b1 , w_43458 );
or ( w_43455 , \6637_b0 , \6638_b0 );
not ( \6638_b0 , w_43459 );
and ( w_43459 , w_43458 , \6638_b1 );
or ( \6644_b1 , \6641_b1 , w_43462 );
or ( \6644_b0 , \6641_b0 , w_43461 );
not ( w_43461 , w_43463 );
and ( w_43463 , w_43462 , w_43460 );
or ( w_43460 , \6642_b1 , w_43464 );
or ( w_43461 , \6642_b0 , \6643_b0 );
not ( \6643_b0 , w_43465 );
and ( w_43465 , w_43464 , \6643_b1 );
or ( \6649_b1 , \6479_b1 , w_43468 );
or ( \6649_b0 , \6479_b0 , w_43467 );
not ( w_43467 , w_43469 );
and ( w_43469 , w_43468 , w_43466 );
or ( w_43466 , \6647_b1 , w_43470 );
or ( w_43467 , \6647_b0 , \6648_b0 );
not ( \6648_b0 , w_43471 );
and ( w_43471 , w_43470 , \6648_b1 );
or ( \6653_b1 , \6650_b1 , w_43474 );
or ( \6653_b0 , \6650_b0 , w_43473 );
not ( w_43473 , w_43475 );
and ( w_43475 , w_43474 , w_43472 );
or ( w_43472 , \6651_b1 , w_43476 );
or ( w_43473 , \6651_b0 , \6652_b0 );
not ( \6652_b0 , w_43477 );
and ( w_43477 , w_43476 , \6652_b1 );
or ( \6657_b1 , \6654_b1 , w_43480 );
or ( \6657_b0 , \6654_b0 , w_43479 );
not ( w_43479 , w_43481 );
and ( w_43481 , w_43480 , w_43478 );
or ( w_43478 , \6655_b1 , w_43482 );
or ( w_43479 , \6655_b0 , \6656_b0 );
not ( \6656_b0 , w_43483 );
and ( w_43483 , w_43482 , \6656_b1 );
or ( \6662_b1 , \6659_b1 , w_43486 );
or ( \6662_b0 , \6659_b0 , w_43485 );
not ( w_43485 , w_43487 );
and ( w_43487 , w_43486 , w_43484 );
or ( w_43484 , \6660_b1 , w_43488 );
or ( w_43485 , \6660_b0 , \6661_b0 );
not ( \6661_b0 , w_43489 );
and ( w_43489 , w_43488 , \6661_b1 );
or ( \6668_b1 , \6665_b1 , w_43492 );
or ( \6668_b0 , \6665_b0 , w_43491 );
not ( w_43491 , w_43493 );
and ( w_43493 , w_43492 , w_43490 );
or ( w_43490 , \6666_b1 , w_43494 );
or ( w_43491 , \6666_b0 , \6667_b0 );
not ( \6667_b0 , w_43495 );
and ( w_43495 , w_43494 , \6667_b1 );
or ( \6672_b1 , \6669_b1 , w_43498 );
or ( \6672_b0 , \6669_b0 , w_43497 );
not ( w_43497 , w_43499 );
and ( w_43499 , w_43498 , w_43496 );
or ( w_43496 , \6670_b1 , w_43500 );
or ( w_43497 , \6670_b0 , \6671_b0 );
not ( \6671_b0 , w_43501 );
and ( w_43501 , w_43500 , \6671_b1 );
or ( \6677_b1 , \6673_b1 , w_43504 );
or ( \6677_b0 , \6673_b0 , w_43503 );
not ( w_43503 , w_43505 );
and ( w_43505 , w_43504 , w_43502 );
or ( w_43502 , \6675_b1 , w_43506 );
or ( w_43503 , \6675_b0 , \6676_b0 );
not ( \6676_b0 , w_43507 );
and ( w_43507 , w_43506 , \6676_b1 );
or ( \6681_b1 , \6678_b1 , w_43510 );
or ( \6681_b0 , \6678_b0 , w_43509 );
not ( w_43509 , w_43511 );
and ( w_43511 , w_43510 , w_43508 );
or ( w_43508 , \6679_b1 , w_43512 );
or ( w_43509 , \6679_b0 , \6680_b0 );
not ( \6680_b0 , w_43513 );
and ( w_43513 , w_43512 , \6680_b1 );
or ( \6686_b1 , \6683_b1 , w_43516 );
or ( \6686_b0 , \6683_b0 , w_43515 );
not ( w_43515 , w_43517 );
and ( w_43517 , w_43516 , w_43514 );
or ( w_43514 , \6684_b1 , w_43518 );
or ( w_43515 , \6684_b0 , \6685_b0 );
not ( \6685_b0 , w_43519 );
and ( w_43519 , w_43518 , \6685_b1 );
or ( \6690_b1 , \6687_b1 , w_43522 );
or ( \6690_b0 , \6687_b0 , w_43521 );
not ( w_43521 , w_43523 );
and ( w_43523 , w_43522 , w_43520 );
or ( w_43520 , \6688_b1 , w_43524 );
or ( w_43521 , \6688_b0 , \6689_b0 );
not ( \6689_b0 , w_43525 );
and ( w_43525 , w_43524 , \6689_b1 );
or ( \6695_b1 , \6692_b1 , w_43528 );
or ( \6695_b0 , \6692_b0 , w_43527 );
not ( w_43527 , w_43529 );
and ( w_43529 , w_43528 , w_43526 );
or ( w_43526 , \6693_b1 , w_43530 );
or ( w_43527 , \6693_b0 , \6694_b0 );
not ( \6694_b0 , w_43531 );
and ( w_43531 , w_43530 , \6694_b1 );
or ( \6700_b1 , \6697_b1 , w_43534 );
or ( \6700_b0 , \6697_b0 , w_43533 );
not ( w_43533 , w_43535 );
and ( w_43535 , w_43534 , w_43532 );
or ( w_43532 , \6698_b1 , w_43536 );
or ( w_43533 , \6698_b0 , \6699_b0 );
not ( \6699_b0 , w_43537 );
and ( w_43537 , w_43536 , \6699_b1 );
or ( \6704_b1 , \6701_b1 , w_43540 );
or ( \6704_b0 , \6701_b0 , w_43539 );
not ( w_43539 , w_43541 );
and ( w_43541 , w_43540 , w_43538 );
or ( w_43538 , \6702_b1 , w_43542 );
or ( w_43539 , \6702_b0 , \6703_b0 );
not ( \6703_b0 , w_43543 );
and ( w_43543 , w_43542 , \6703_b1 );
or ( \6709_b1 , \6706_b1 , w_43546 );
or ( \6709_b0 , \6706_b0 , w_43545 );
not ( w_43545 , w_43547 );
and ( w_43547 , w_43546 , w_43544 );
or ( w_43544 , \6707_b1 , w_43548 );
or ( w_43545 , \6707_b0 , \6708_b0 );
not ( \6708_b0 , w_43549 );
and ( w_43549 , w_43548 , \6708_b1 );
or ( \6715_b1 , \6712_b1 , w_43552 );
or ( \6715_b0 , \6712_b0 , w_43551 );
not ( w_43551 , w_43553 );
and ( w_43553 , w_43552 , w_43550 );
or ( w_43550 , \6713_b1 , w_43554 );
or ( w_43551 , \6713_b0 , \6714_b0 );
not ( \6714_b0 , w_43555 );
and ( w_43555 , w_43554 , \6714_b1 );
or ( \6805_b1 , \6802_b1 , w_43558 );
or ( \6805_b0 , \6802_b0 , w_43557 );
not ( w_43557 , w_43559 );
and ( w_43559 , w_43558 , w_43556 );
or ( w_43556 , \6803_b1 , w_43560 );
or ( w_43557 , \6803_b0 , \6804_b0 );
not ( \6804_b0 , w_43561 );
and ( w_43561 , w_43560 , \6804_b1 );
or ( \6809_b1 , \6806_b1 , w_43564 );
or ( \6809_b0 , \6806_b0 , w_43563 );
not ( w_43563 , w_43565 );
and ( w_43565 , w_43564 , w_43562 );
or ( w_43562 , \6807_b1 , w_43566 );
or ( w_43563 , \6807_b0 , \6808_b0 );
not ( \6808_b0 , w_43567 );
and ( w_43567 , w_43566 , \6808_b1 );
or ( \6837_b1 , \6830_b1 , w_43570 );
or ( \6837_b0 , \6830_b0 , w_43569 );
not ( w_43569 , w_43571 );
and ( w_43571 , w_43570 , w_43568 );
or ( w_43568 , \6835_b1 , w_43572 );
or ( w_43569 , \6835_b0 , \6836_b0 );
not ( \6836_b0 , w_43573 );
and ( w_43573 , w_43572 , \6836_b1 );
or ( \6853_b1 , \6846_b1 , w_43576 );
or ( \6853_b0 , \6846_b0 , w_43575 );
not ( w_43575 , w_43577 );
and ( w_43577 , w_43576 , w_43574 );
or ( w_43574 , \6851_b1 , w_43578 );
or ( w_43575 , \6851_b0 , \6852_b0 );
not ( \6852_b0 , w_43579 );
and ( w_43579 , w_43578 , \6852_b1 );
or ( \6870_b1 , \6863_b1 , w_43582 );
or ( \6870_b0 , \6863_b0 , w_43581 );
not ( w_43581 , w_43583 );
and ( w_43583 , w_43582 , w_43580 );
or ( w_43580 , \6868_b1 , w_43584 );
or ( w_43581 , \6868_b0 , \6869_b0 );
not ( \6869_b0 , w_43585 );
and ( w_43585 , w_43584 , \6869_b1 );
or ( \6873_b1 , \6854_b1 , w_43588 );
or ( \6873_b0 , \6854_b0 , w_43587 );
not ( w_43587 , w_43589 );
and ( w_43589 , w_43588 , w_43586 );
or ( w_43586 , \6871_b1 , w_43590 );
or ( w_43587 , \6871_b0 , \6872_b0 );
not ( \6872_b0 , w_43591 );
and ( w_43591 , w_43590 , \6872_b1 );
or ( \6889_b1 , \6882_b1 , w_43594 );
or ( \6889_b0 , \6882_b0 , w_43593 );
not ( w_43593 , w_43595 );
and ( w_43595 , w_43594 , w_43592 );
or ( w_43592 , \6887_b1 , w_43596 );
or ( w_43593 , \6887_b0 , \6888_b0 );
not ( \6888_b0 , w_43597 );
and ( w_43597 , w_43596 , \6888_b1 );
or ( \6905_b1 , \6898_b1 , w_43600 );
or ( \6905_b0 , \6898_b0 , w_43599 );
not ( w_43599 , w_43601 );
and ( w_43601 , w_43600 , w_43598 );
or ( w_43598 , \6903_b1 , w_43602 );
or ( w_43599 , \6903_b0 , \6904_b0 );
not ( \6904_b0 , w_43603 );
and ( w_43603 , w_43602 , \6904_b1 );
or ( \6918_b1 , \6906_b1 , w_43606 );
or ( \6918_b0 , \6906_b0 , w_43605 );
not ( w_43605 , w_43607 );
and ( w_43607 , w_43606 , w_43604 );
or ( w_43604 , \6916_b1 , w_43608 );
or ( w_43605 , \6916_b0 , \6917_b0 );
not ( \6917_b0 , w_43609 );
and ( w_43609 , w_43608 , \6917_b1 );
or ( \6927_b1 , \6919_b1 , w_43612 );
or ( \6927_b0 , \6919_b0 , w_43611 );
not ( w_43611 , w_43613 );
and ( w_43613 , w_43612 , w_43610 );
or ( w_43610 , \6925_b1 , w_43614 );
or ( w_43611 , \6925_b0 , \6926_b0 );
not ( \6926_b0 , w_43615 );
and ( w_43615 , w_43614 , \6926_b1 );
or ( \6937_b1 , \6932_b1 , w_43618 );
or ( \6937_b0 , \6932_b0 , w_43617 );
not ( w_43617 , w_43619 );
and ( w_43619 , w_43618 , w_43616 );
or ( w_43616 , \6935_b1 , w_43620 );
or ( w_43617 , \6935_b0 , \6936_b0 );
not ( \6936_b0 , w_43621 );
and ( w_43621 , w_43620 , \6936_b1 );
or ( \6945_b1 , \6940_b1 , w_43624 );
or ( \6945_b0 , \6940_b0 , w_43623 );
not ( w_43623 , w_43625 );
and ( w_43625 , w_43624 , w_43622 );
or ( w_43622 , \6943_b1 , w_43626 );
or ( w_43623 , \6943_b0 , \6944_b0 );
not ( \6944_b0 , w_43627 );
and ( w_43627 , w_43626 , \6944_b1 );
or ( \6954_b1 , \6946_b1 , w_43630 );
or ( \6954_b0 , \6946_b0 , w_43629 );
not ( w_43629 , w_43631 );
and ( w_43631 , w_43630 , w_43628 );
or ( w_43628 , \6952_b1 , w_43632 );
or ( w_43629 , \6952_b0 , \6953_b0 );
not ( \6953_b0 , w_43633 );
and ( w_43633 , w_43632 , \6953_b1 );
or ( \6964_b1 , \6959_b1 , w_43636 );
or ( \6964_b0 , \6959_b0 , w_43635 );
not ( w_43635 , w_43637 );
and ( w_43637 , w_43636 , w_43634 );
or ( w_43634 , \6962_b1 , w_43638 );
or ( w_43635 , \6962_b0 , \6963_b0 );
not ( \6963_b0 , w_43639 );
and ( w_43639 , w_43638 , \6963_b1 );
or ( \6970_b1 , \6965_b1 , w_43642 );
or ( \6970_b0 , \6965_b0 , w_43641 );
not ( w_43641 , w_43643 );
and ( w_43643 , w_43642 , w_43640 );
or ( w_43640 , \6968_b1 , w_43644 );
or ( w_43641 , \6968_b0 , \6969_b0 );
not ( \6969_b0 , w_43645 );
and ( w_43645 , w_43644 , \6969_b1 );
or ( \6978_b1 , \6973_b1 , w_43648 );
or ( \6978_b0 , \6973_b0 , w_43647 );
not ( w_43647 , w_43649 );
and ( w_43649 , w_43648 , w_43646 );
or ( w_43646 , \6976_b1 , w_43650 );
or ( w_43647 , \6976_b0 , \6977_b0 );
not ( \6977_b0 , w_43651 );
and ( w_43651 , w_43650 , \6977_b1 );
or ( \7016_b1 , \6996_b1 , w_43654 );
or ( \7016_b0 , \6996_b0 , w_43653 );
not ( w_43653 , w_43655 );
and ( w_43655 , w_43654 , w_43652 );
or ( w_43652 , \7014_b1 , w_43656 );
or ( w_43653 , \7014_b0 , \7015_b0 );
not ( \7015_b0 , w_43657 );
and ( w_43657 , w_43656 , \7015_b1 );
or ( \7071_b1 , \7051_b1 , w_43660 );
or ( \7071_b0 , \7051_b0 , w_43659 );
not ( w_43659 , w_43661 );
and ( w_43661 , w_43660 , w_43658 );
or ( w_43658 , \7069_b1 , w_43662 );
or ( w_43659 , \7069_b0 , \7070_b0 );
not ( \7070_b0 , w_43663 );
and ( w_43663 , w_43662 , \7070_b1 );
or ( \7127_b1 , \7107_b1 , w_43666 );
or ( \7127_b0 , \7107_b0 , w_43665 );
not ( w_43665 , w_43667 );
and ( w_43667 , w_43666 , w_43664 );
or ( w_43664 , \7125_b1 , w_43668 );
or ( w_43665 , \7125_b0 , \7126_b0 );
not ( \7126_b0 , w_43669 );
and ( w_43669 , w_43668 , \7126_b1 );
or ( \7130_b1 , \7072_b1 , w_43672 );
or ( \7130_b0 , \7072_b0 , w_43671 );
not ( w_43671 , w_43673 );
and ( w_43673 , w_43672 , w_43670 );
or ( w_43670 , \7128_b1 , w_43674 );
or ( w_43671 , \7128_b0 , \7129_b0 );
not ( \7129_b0 , w_43675 );
and ( w_43675 , w_43674 , \7129_b1 );
or ( \7185_b1 , \7165_b1 , w_43678 );
or ( \7185_b0 , \7165_b0 , w_43677 );
not ( w_43677 , w_43679 );
and ( w_43679 , w_43678 , w_43676 );
or ( w_43676 , \7183_b1 , w_43680 );
or ( w_43677 , \7183_b0 , \7184_b0 );
not ( \7184_b0 , w_43681 );
and ( w_43681 , w_43680 , \7184_b1 );
or ( \7213_b1 , \7208_b1 , w_43684 );
or ( \7213_b0 , \7208_b0 , w_43683 );
not ( w_43683 , w_43685 );
and ( w_43685 , w_43684 , w_43682 );
or ( w_43682 , \7211_b1 , w_43686 );
or ( w_43683 , \7211_b0 , \7212_b0 );
not ( \7212_b0 , w_43687 );
and ( w_43687 , w_43686 , \7212_b1 );
or ( \7221_b1 , \7214_b1 , w_43690 );
or ( \7221_b0 , \7214_b0 , w_43689 );
not ( w_43689 , w_43691 );
and ( w_43691 , w_43690 , w_43688 );
or ( w_43688 , \7219_b1 , w_43692 );
or ( w_43689 , \7219_b0 , \7220_b0 );
not ( \7220_b0 , w_43693 );
and ( w_43693 , w_43692 , \7220_b1 );
or ( \7258_b1 , \7241_b1 , w_43696 );
or ( \7258_b0 , \7241_b0 , w_43695 );
not ( w_43695 , w_43697 );
and ( w_43697 , w_43696 , w_43694 );
or ( w_43694 , \7256_b1 , w_43698 );
or ( w_43695 , \7256_b0 , \7257_b0 );
not ( \7257_b0 , w_43699 );
and ( w_43699 , w_43698 , \7257_b1 );
or ( \7261_b1 , \7222_b1 , w_43702 );
or ( \7261_b0 , \7222_b0 , w_43701 );
not ( w_43701 , w_43703 );
and ( w_43703 , w_43702 , w_43700 );
or ( w_43700 , \7259_b1 , w_43704 );
or ( w_43701 , \7259_b0 , \7260_b0 );
not ( \7260_b0 , w_43705 );
and ( w_43705 , w_43704 , \7260_b1 );
or ( \7320_b1 , \7317_b1 , w_43708 );
or ( \7320_b0 , \7317_b0 , w_43707 );
not ( w_43707 , w_43709 );
and ( w_43709 , w_43708 , w_43706 );
or ( w_43706 , \7318_b1 , w_43710 );
or ( w_43707 , \7318_b0 , \7319_b0 );
not ( \7319_b0 , w_43711 );
and ( w_43711 , w_43710 , \7319_b1 );
or ( \7341_b1 , \7316_b1 , w_43714 );
or ( \7341_b0 , \7316_b0 , w_43713 );
not ( w_43713 , w_43715 );
and ( w_43715 , w_43714 , w_43712 );
or ( w_43712 , \7339_b1 , w_43716 );
or ( w_43713 , \7339_b0 , \7340_b0 );
not ( \7340_b0 , w_43717 );
and ( w_43717 , w_43716 , \7340_b1 );
or ( \7346_b1 , \7343_b1 , w_43720 );
or ( \7346_b0 , \7343_b0 , w_43719 );
not ( w_43719 , w_43721 );
and ( w_43721 , w_43720 , w_43718 );
or ( w_43718 , \7344_b1 , w_43722 );
or ( w_43719 , \7344_b0 , \7345_b0 );
not ( \7345_b0 , w_43723 );
and ( w_43723 , w_43722 , \7345_b1 );
or ( \7350_b1 , \7347_b1 , w_43726 );
or ( \7350_b0 , \7347_b0 , w_43725 );
not ( w_43725 , w_43727 );
and ( w_43727 , w_43726 , w_43724 );
or ( w_43724 , \7348_b1 , w_43728 );
or ( w_43725 , \7348_b0 , \7349_b0 );
not ( \7349_b0 , w_43729 );
and ( w_43729 , w_43728 , \7349_b1 );
or ( \7355_b1 , \7352_b1 , w_43732 );
or ( \7355_b0 , \7352_b0 , w_43731 );
not ( w_43731 , w_43733 );
and ( w_43733 , w_43732 , w_43730 );
or ( w_43730 , \7353_b1 , w_43734 );
or ( w_43731 , \7353_b0 , \7354_b0 );
not ( \7354_b0 , w_43735 );
and ( w_43735 , w_43734 , \7354_b1 );
or ( \7359_b1 , \7342_b1 , w_43738 );
or ( \7359_b0 , \7342_b0 , w_43737 );
not ( w_43737 , w_43739 );
and ( w_43739 , w_43738 , w_43736 );
or ( w_43736 , \7357_b1 , w_43740 );
or ( w_43737 , \7357_b0 , \7358_b0 );
not ( \7358_b0 , w_43741 );
and ( w_43741 , w_43740 , \7358_b1 );
or ( \7422_b1 , \7419_b1 , w_43744 );
or ( \7422_b0 , \7419_b0 , w_43743 );
not ( w_43743 , w_43745 );
and ( w_43745 , w_43744 , w_43742 );
or ( w_43742 , \7420_b1 , w_43746 );
or ( w_43743 , \7420_b0 , \7421_b0 );
not ( \7421_b0 , w_43747 );
and ( w_43747 , w_43746 , \7421_b1 );
or ( \7426_b1 , \7423_b1 , w_43750 );
or ( \7426_b0 , \7423_b0 , w_43749 );
not ( w_43749 , w_43751 );
and ( w_43751 , w_43750 , w_43748 );
or ( w_43748 , \7424_b1 , w_43752 );
or ( w_43749 , \7424_b0 , \7425_b0 );
not ( \7425_b0 , w_43753 );
and ( w_43753 , w_43752 , \7425_b1 );
or ( \7459_b1 , \7452_b1 , w_43756 );
or ( \7459_b0 , \7452_b0 , w_43755 );
not ( w_43755 , w_43757 );
and ( w_43757 , w_43756 , w_43754 );
or ( w_43754 , \7457_b1 , w_43758 );
or ( w_43755 , \7457_b0 , \7458_b0 );
not ( \7458_b0 , w_43759 );
and ( w_43759 , w_43758 , \7458_b1 );
or ( \7475_b1 , \7468_b1 , w_43762 );
or ( \7475_b0 , \7468_b0 , w_43761 );
not ( w_43761 , w_43763 );
and ( w_43763 , w_43762 , w_43760 );
or ( w_43760 , \7473_b1 , w_43764 );
or ( w_43761 , \7473_b0 , \7474_b0 );
not ( \7474_b0 , w_43765 );
and ( w_43765 , w_43764 , \7474_b1 );
or ( \7480_b1 , \7477_b1 , w_43768 );
or ( \7480_b0 , \7477_b0 , w_43767 );
not ( w_43767 , w_43769 );
and ( w_43769 , w_43768 , w_43766 );
or ( w_43766 , \7478_b1 , w_43770 );
or ( w_43767 , \7478_b0 , \7479_b0 );
not ( \7479_b0 , w_43771 );
and ( w_43771 , w_43770 , \7479_b1 );
or ( \7483_b1 , \7476_b1 , w_43774 );
or ( \7483_b0 , \7476_b0 , w_43773 );
not ( w_43773 , w_43775 );
and ( w_43775 , w_43774 , w_43772 );
or ( w_43772 , \7481_b1 , w_43776 );
or ( w_43773 , \7481_b0 , \7482_b0 );
not ( \7482_b0 , w_43777 );
and ( w_43777 , w_43776 , \7482_b1 );
or ( \7487_b1 , \7484_b1 , w_43780 );
or ( \7487_b0 , \7484_b0 , w_43779 );
not ( w_43779 , w_43781 );
and ( w_43781 , w_43780 , w_43778 );
or ( w_43778 , \7485_b1 , w_43782 );
or ( w_43779 , \7485_b0 , \7486_b0 );
not ( \7486_b0 , w_43783 );
and ( w_43783 , w_43782 , \7486_b1 );
or ( \7492_b1 , \7489_b1 , w_43786 );
or ( \7492_b0 , \7489_b0 , w_43785 );
not ( w_43785 , w_43787 );
and ( w_43787 , w_43786 , w_43784 );
or ( w_43784 , \7490_b1 , w_43788 );
or ( w_43785 , \7490_b0 , \7491_b0 );
not ( \7491_b0 , w_43789 );
and ( w_43789 , w_43788 , \7491_b1 );
or ( \7572_b1 , \7569_b1 , w_43792 );
or ( \7572_b0 , \7569_b0 , w_43791 );
not ( w_43791 , w_43793 );
and ( w_43793 , w_43792 , w_43790 );
or ( w_43790 , \7570_b1 , w_43794 );
or ( w_43791 , \7570_b0 , \7571_b0 );
not ( \7571_b0 , w_43795 );
and ( w_43795 , w_43794 , \7571_b1 );
or ( \7576_b1 , \7573_b1 , w_43798 );
or ( \7576_b0 , \7573_b0 , w_43797 );
not ( w_43797 , w_43799 );
and ( w_43799 , w_43798 , w_43796 );
or ( w_43796 , \7574_b1 , w_43800 );
or ( w_43797 , \7574_b0 , \7575_b0 );
not ( \7575_b0 , w_43801 );
and ( w_43801 , w_43800 , \7575_b1 );
or ( \7586_b1 , \7495_b1 , w_43804 );
or ( \7586_b0 , \7495_b0 , w_43803 );
not ( w_43803 , w_43805 );
and ( w_43805 , w_43804 , w_43802 );
or ( w_43802 , \7584_b1 , w_43806 );
or ( w_43803 , \7584_b0 , \7585_b0 );
not ( \7585_b0 , w_43807 );
and ( w_43807 , w_43806 , \7585_b1 );
or ( \7590_b1 , \7587_b1 , w_43810 );
or ( \7590_b0 , \7587_b0 , w_43809 );
not ( w_43809 , w_43811 );
and ( w_43811 , w_43810 , w_43808 );
or ( w_43808 , \7588_b1 , w_43812 );
or ( w_43809 , \7588_b0 , \7589_b0 );
not ( \7589_b0 , w_43813 );
and ( w_43813 , w_43812 , \7589_b1 );
or ( \7594_b1 , \7591_b1 , w_43816 );
or ( \7594_b0 , \7591_b0 , w_43815 );
not ( w_43815 , w_43817 );
and ( w_43817 , w_43816 , w_43814 );
or ( w_43814 , \7592_b1 , w_43818 );
or ( w_43815 , \7592_b0 , \7593_b0 );
not ( \7593_b0 , w_43819 );
and ( w_43819 , w_43818 , \7593_b1 );
or ( \7599_b1 , \7596_b1 , w_43822 );
or ( \7599_b0 , \7596_b0 , w_43821 );
not ( w_43821 , w_43823 );
and ( w_43823 , w_43822 , w_43820 );
or ( w_43820 , \7597_b1 , w_43824 );
or ( w_43821 , \7597_b0 , \7598_b0 );
not ( \7598_b0 , w_43825 );
and ( w_43825 , w_43824 , \7598_b1 );
or ( \7604_b1 , \7601_b1 , w_43828 );
or ( \7604_b0 , \7601_b0 , w_43827 );
not ( w_43827 , w_43829 );
and ( w_43829 , w_43828 , w_43826 );
or ( w_43826 , \7602_b1 , w_43830 );
or ( w_43827 , \7602_b0 , \7603_b0 );
not ( \7603_b0 , w_43831 );
and ( w_43831 , w_43830 , \7603_b1 );
or ( \7608_b1 , \7605_b1 , w_43834 );
or ( \7608_b0 , \7605_b0 , w_43833 );
not ( w_43833 , w_43835 );
and ( w_43835 , w_43834 , w_43832 );
or ( w_43832 , \7606_b1 , w_43836 );
or ( w_43833 , \7606_b0 , \7607_b0 );
not ( \7607_b0 , w_43837 );
and ( w_43837 , w_43836 , \7607_b1 );
or ( \7613_b1 , \7610_b1 , w_43840 );
or ( \7613_b0 , \7610_b0 , w_43839 );
not ( w_43839 , w_43841 );
and ( w_43841 , w_43840 , w_43838 );
or ( w_43838 , \7611_b1 , w_43842 );
or ( w_43839 , \7611_b0 , \7612_b0 );
not ( \7612_b0 , w_43843 );
and ( w_43843 , w_43842 , \7612_b1 );
or ( \7617_b1 , \7614_b1 , w_43846 );
or ( \7617_b0 , \7614_b0 , w_43845 );
not ( w_43845 , w_43847 );
and ( w_43847 , w_43846 , w_43844 );
or ( w_43844 , \7615_b1 , w_43848 );
or ( w_43845 , \7615_b0 , \7616_b0 );
not ( \7616_b0 , w_43849 );
and ( w_43849 , w_43848 , \7616_b1 );
or ( \7622_b1 , \7619_b1 , w_43852 );
or ( \7622_b0 , \7619_b0 , w_43851 );
not ( w_43851 , w_43853 );
and ( w_43853 , w_43852 , w_43850 );
or ( w_43850 , \7620_b1 , w_43854 );
or ( w_43851 , \7620_b0 , \7621_b0 );
not ( \7621_b0 , w_43855 );
and ( w_43855 , w_43854 , \7621_b1 );
or ( \7630_b1 , \7627_b1 , w_43858 );
or ( \7630_b0 , \7627_b0 , w_43857 );
not ( w_43857 , w_43859 );
and ( w_43859 , w_43858 , w_43856 );
or ( w_43856 , \7628_b1 , w_43860 );
or ( w_43857 , \7628_b0 , \7629_b0 );
not ( \7629_b0 , w_43861 );
and ( w_43861 , w_43860 , \7629_b1 );
or ( \7634_b1 , \7631_b1 , w_43864 );
or ( \7634_b0 , \7631_b0 , w_43863 );
not ( w_43863 , w_43865 );
and ( w_43865 , w_43864 , w_43862 );
or ( w_43862 , \7632_b1 , w_43866 );
or ( w_43863 , \7632_b0 , \7633_b0 );
not ( \7633_b0 , w_43867 );
and ( w_43867 , w_43866 , \7633_b1 );
or ( \7668_b1 , \7665_b1 , w_43870 );
or ( \7668_b0 , \7665_b0 , w_43869 );
not ( w_43869 , w_43871 );
and ( w_43871 , w_43870 , w_43868 );
or ( w_43868 , \7666_b1 , w_43872 );
or ( w_43869 , \7666_b0 , \7667_b0 );
not ( \7667_b0 , w_43873 );
and ( w_43873 , w_43872 , \7667_b1 );
or ( \7672_b1 , \7669_b1 , w_43876 );
or ( \7672_b0 , \7669_b0 , w_43875 );
not ( w_43875 , w_43877 );
and ( w_43877 , w_43876 , w_43874 );
or ( w_43874 , \7670_b1 , w_43878 );
or ( w_43875 , \7670_b0 , \7671_b0 );
not ( \7671_b0 , w_43879 );
and ( w_43879 , w_43878 , \7671_b1 );
or ( \7677_b1 , \7674_b1 , w_43882 );
or ( \7677_b0 , \7674_b0 , w_43881 );
not ( w_43881 , w_43883 );
and ( w_43883 , w_43882 , w_43880 );
or ( w_43880 , \7675_b1 , w_43884 );
or ( w_43881 , \7675_b0 , \7676_b0 );
not ( \7676_b0 , w_43885 );
and ( w_43885 , w_43884 , \7676_b1 );
or ( \7684_b1 , \7681_b1 , w_43888 );
or ( \7684_b0 , \7681_b0 , w_43887 );
not ( w_43887 , w_43889 );
and ( w_43889 , w_43888 , w_43886 );
or ( w_43886 , \7682_b1 , w_43890 );
or ( w_43887 , \7682_b0 , \7683_b0 );
not ( \7683_b0 , w_43891 );
and ( w_43891 , w_43890 , \7683_b1 );
or ( \7688_b1 , \7685_b1 , w_43894 );
or ( \7688_b0 , \7685_b0 , w_43893 );
not ( w_43893 , w_43895 );
and ( w_43895 , w_43894 , w_43892 );
or ( w_43892 , \7686_b1 , w_43896 );
or ( w_43893 , \7686_b0 , \7687_b0 );
not ( \7687_b0 , w_43897 );
and ( w_43897 , w_43896 , \7687_b1 );
or ( \7737_b1 , \7734_b1 , w_43900 );
or ( \7737_b0 , \7734_b0 , w_43899 );
not ( w_43899 , w_43901 );
and ( w_43901 , w_43900 , w_43898 );
or ( w_43898 , \7735_b1 , w_43902 );
or ( w_43899 , \7735_b0 , \7736_b0 );
not ( \7736_b0 , w_43903 );
and ( w_43903 , w_43902 , \7736_b1 );
or ( \7741_b1 , \7738_b1 , w_43906 );
or ( \7741_b0 , \7738_b0 , w_43905 );
not ( w_43905 , w_43907 );
and ( w_43907 , w_43906 , w_43904 );
or ( w_43904 , \7739_b1 , w_43908 );
or ( w_43905 , \7739_b0 , \7740_b0 );
not ( \7740_b0 , w_43909 );
and ( w_43909 , w_43908 , \7740_b1 );
or ( \7752_b1 , \7749_b1 , w_43912 );
or ( \7752_b0 , \7749_b0 , w_43911 );
not ( w_43911 , w_43913 );
and ( w_43913 , w_43912 , w_43910 );
or ( w_43910 , \7750_b1 , w_43914 );
or ( w_43911 , \7750_b0 , \7751_b0 );
not ( \7751_b0 , w_43915 );
and ( w_43915 , w_43914 , \7751_b1 );
or ( \7756_b1 , \7753_b1 , w_43918 );
or ( \7756_b0 , \7753_b0 , w_43917 );
not ( w_43917 , w_43919 );
and ( w_43919 , w_43918 , w_43916 );
or ( w_43916 , \7754_b1 , w_43920 );
or ( w_43917 , \7754_b0 , \7755_b0 );
not ( \7755_b0 , w_43921 );
and ( w_43921 , w_43920 , \7755_b1 );
or ( \7761_b1 , \7758_b1 , w_43924 );
or ( \7761_b0 , \7758_b0 , w_43923 );
not ( w_43923 , w_43925 );
and ( w_43925 , w_43924 , w_43922 );
or ( w_43922 , \7759_b1 , w_43926 );
or ( w_43923 , \7759_b0 , \7760_b0 );
not ( \7760_b0 , w_43927 );
and ( w_43927 , w_43926 , \7760_b1 );
or ( \7782_b1 , \7775_b1 , w_43930 );
or ( \7782_b0 , \7775_b0 , w_43929 );
not ( w_43929 , w_43931 );
and ( w_43931 , w_43930 , w_43928 );
or ( w_43928 , \7780_b1 , w_43932 );
or ( w_43929 , \7780_b0 , \7781_b0 );
not ( \7781_b0 , w_43933 );
and ( w_43933 , w_43932 , \7781_b1 );
or ( \7798_b1 , \7791_b1 , w_43936 );
or ( \7798_b0 , \7791_b0 , w_43935 );
not ( w_43935 , w_43937 );
and ( w_43937 , w_43936 , w_43934 );
or ( w_43934 , \7796_b1 , w_43938 );
or ( w_43935 , \7796_b0 , \7797_b0 );
not ( \7797_b0 , w_43939 );
and ( w_43939 , w_43938 , \7797_b1 );
or ( \7815_b1 , \7808_b1 , w_43942 );
or ( \7815_b0 , \7808_b0 , w_43941 );
not ( w_43941 , w_43943 );
and ( w_43943 , w_43942 , w_43940 );
or ( w_43940 , \7813_b1 , w_43944 );
or ( w_43941 , \7813_b0 , \7814_b0 );
not ( \7814_b0 , w_43945 );
and ( w_43945 , w_43944 , \7814_b1 );
or ( \7818_b1 , \7799_b1 , w_43948 );
or ( \7818_b0 , \7799_b0 , w_43947 );
not ( w_43947 , w_43949 );
and ( w_43949 , w_43948 , w_43946 );
or ( w_43946 , \7816_b1 , w_43950 );
or ( w_43947 , \7816_b0 , \7817_b0 );
not ( \7817_b0 , w_43951 );
and ( w_43951 , w_43950 , \7817_b1 );
or ( \7834_b1 , \7827_b1 , w_43954 );
or ( \7834_b0 , \7827_b0 , w_43953 );
not ( w_43953 , w_43955 );
and ( w_43955 , w_43954 , w_43952 );
or ( w_43952 , \7832_b1 , w_43956 );
or ( w_43953 , \7832_b0 , \7833_b0 );
not ( \7833_b0 , w_43957 );
and ( w_43957 , w_43956 , \7833_b1 );
or ( \7842_b1 , \7837_b1 , w_43960 );
or ( \7842_b0 , \7837_b0 , w_43959 );
not ( w_43959 , w_43961 );
and ( w_43961 , w_43960 , w_43958 );
or ( w_43958 , \7840_b1 , w_43962 );
or ( w_43959 , \7840_b0 , \7841_b0 );
not ( \7841_b0 , w_43963 );
and ( w_43963 , w_43962 , \7841_b1 );
or ( \7853_b1 , \7848_b1 , w_43966 );
or ( \7853_b0 , \7848_b0 , w_43965 );
not ( w_43965 , w_43967 );
and ( w_43967 , w_43966 , w_43964 );
or ( w_43964 , \7851_b1 , w_43968 );
or ( w_43965 , \7851_b0 , \7852_b0 );
not ( \7852_b0 , w_43969 );
and ( w_43969 , w_43968 , \7852_b1 );
or ( \7856_b1 , \7843_b1 , w_43972 );
or ( \7856_b0 , \7843_b0 , w_43971 );
not ( w_43971 , w_43973 );
and ( w_43973 , w_43972 , w_43970 );
or ( w_43970 , \7854_b1 , w_43974 );
or ( w_43971 , \7854_b0 , \7855_b0 );
not ( \7855_b0 , w_43975 );
and ( w_43975 , w_43974 , \7855_b1 );
or ( \7866_b1 , \7861_b1 , w_43978 );
or ( \7866_b0 , \7861_b0 , w_43977 );
not ( w_43977 , w_43979 );
and ( w_43979 , w_43978 , w_43976 );
or ( w_43976 , \7864_b1 , w_43980 );
or ( w_43977 , \7864_b0 , \7865_b0 );
not ( \7865_b0 , w_43981 );
and ( w_43981 , w_43980 , \7865_b1 );
or ( \7872_b1 , \7867_b1 , w_43984 );
or ( \7872_b0 , \7867_b0 , w_43983 );
not ( w_43983 , w_43985 );
and ( w_43985 , w_43984 , w_43982 );
or ( w_43982 , \7870_b1 , w_43986 );
or ( w_43983 , \7870_b0 , \7871_b0 );
not ( \7871_b0 , w_43987 );
and ( w_43987 , w_43986 , \7871_b1 );
or ( \7879_b1 , \7874_b1 , w_43990 );
or ( \7879_b0 , \7874_b0 , w_43989 );
not ( w_43989 , w_43991 );
and ( w_43991 , w_43990 , w_43988 );
or ( w_43988 , \7877_b1 , w_43992 );
or ( w_43989 , \7877_b0 , \7878_b0 );
not ( \7878_b0 , w_43993 );
and ( w_43993 , w_43992 , \7878_b1 );
or ( \7886_b1 , \7881_b1 , w_43996 );
or ( \7886_b0 , \7881_b0 , w_43995 );
not ( w_43995 , w_43997 );
and ( w_43997 , w_43996 , w_43994 );
or ( w_43994 , \7884_b1 , w_43998 );
or ( w_43995 , \7884_b0 , \7885_b0 );
not ( \7885_b0 , w_43999 );
and ( w_43999 , w_43998 , \7885_b1 );
or ( \7891_b1 , \7888_b1 , w_44002 );
or ( \7891_b0 , \7888_b0 , w_44001 );
not ( w_44001 , w_44003 );
and ( w_44003 , w_44002 , w_44000 );
or ( w_44000 , \7889_b1 , w_44004 );
or ( w_44001 , \7889_b0 , \7890_b0 );
not ( \7890_b0 , w_44005 );
and ( w_44005 , w_44004 , \7890_b1 );
or ( \7895_b1 , \7892_b1 , w_44008 );
or ( \7895_b0 , \7892_b0 , w_44007 );
not ( w_44007 , w_44009 );
and ( w_44009 , w_44008 , w_44006 );
or ( w_44006 , \7893_b1 , w_44010 );
or ( w_44007 , \7893_b0 , \7894_b0 );
not ( \7894_b0 , w_44011 );
and ( w_44011 , w_44010 , \7894_b1 );
or ( \7899_b1 , \7896_b1 , w_44014 );
or ( \7899_b0 , \7896_b0 , w_44013 );
not ( w_44013 , w_44015 );
and ( w_44015 , w_44014 , w_44012 );
or ( w_44012 , \7897_b1 , w_44016 );
or ( w_44013 , \7897_b0 , \7898_b0 );
not ( \7898_b0 , w_44017 );
and ( w_44017 , w_44016 , \7898_b1 );
or ( \7904_b1 , \7901_b1 , w_44020 );
or ( \7904_b0 , \7901_b0 , w_44019 );
not ( w_44019 , w_44021 );
and ( w_44021 , w_44020 , w_44018 );
or ( w_44018 , \7902_b1 , w_44022 );
or ( w_44019 , \7902_b0 , \7903_b0 );
not ( \7903_b0 , w_44023 );
and ( w_44023 , w_44022 , \7903_b1 );
or ( \7910_b1 , \7907_b1 , w_44026 );
or ( \7910_b0 , \7907_b0 , w_44025 );
not ( w_44025 , w_44027 );
and ( w_44027 , w_44026 , w_44024 );
or ( w_44024 , \7908_b1 , w_44028 );
or ( w_44025 , \7908_b0 , \7909_b0 );
not ( \7909_b0 , w_44029 );
and ( w_44029 , w_44028 , \7909_b1 );
or ( \7916_b1 , \7913_b1 , w_44032 );
or ( \7916_b0 , \7913_b0 , w_44031 );
not ( w_44031 , w_44033 );
and ( w_44033 , w_44032 , w_44030 );
or ( w_44030 , \7914_b1 , w_44034 );
or ( w_44031 , \7914_b0 , \7915_b0 );
not ( \7915_b0 , w_44035 );
and ( w_44035 , w_44034 , \7915_b1 );
or ( \7920_b1 , \7917_b1 , w_44038 );
or ( \7920_b0 , \7917_b0 , w_44037 );
not ( w_44037 , w_44039 );
and ( w_44039 , w_44038 , w_44036 );
or ( w_44036 , \7918_b1 , w_44040 );
or ( w_44037 , \7918_b0 , \7919_b0 );
not ( \7919_b0 , w_44041 );
and ( w_44041 , w_44040 , \7919_b1 );
or ( \7938_b1 , \7935_b1 , w_44044 );
or ( \7938_b0 , \7935_b0 , w_44043 );
not ( w_44043 , w_44045 );
and ( w_44045 , w_44044 , w_44042 );
or ( w_44042 , \7936_b1 , w_44046 );
or ( w_44043 , \7936_b0 , \7937_b0 );
not ( \7937_b0 , w_44047 );
and ( w_44047 , w_44046 , \7937_b1 );
or ( \7942_b1 , \7939_b1 , w_44050 );
or ( \7942_b0 , \7939_b0 , w_44049 );
not ( w_44049 , w_44051 );
and ( w_44051 , w_44050 , w_44048 );
or ( w_44048 , \7940_b1 , w_44052 );
or ( w_44049 , \7940_b0 , \7941_b0 );
not ( \7941_b0 , w_44053 );
and ( w_44053 , w_44052 , \7941_b1 );
or ( \7947_b1 , \7944_b1 , w_44056 );
or ( \7947_b0 , \7944_b0 , w_44055 );
not ( w_44055 , w_44057 );
and ( w_44057 , w_44056 , w_44054 );
or ( w_44054 , \7945_b1 , w_44058 );
or ( w_44055 , \7945_b0 , \7946_b0 );
not ( \7946_b0 , w_44059 );
and ( w_44059 , w_44058 , \7946_b1 );
or ( \8023_b1 , \8020_b1 , w_44062 );
or ( \8023_b0 , \8020_b0 , w_44061 );
not ( w_44061 , w_44063 );
and ( w_44063 , w_44062 , w_44060 );
or ( w_44060 , \8021_b1 , w_44064 );
or ( w_44061 , \8021_b0 , \8022_b0 );
not ( \8022_b0 , w_44065 );
and ( w_44065 , w_44064 , \8022_b1 );
or ( \8027_b1 , \8024_b1 , w_44068 );
or ( \8027_b0 , \8024_b0 , w_44067 );
not ( w_44067 , w_44069 );
and ( w_44069 , w_44068 , w_44066 );
or ( w_44066 , \8025_b1 , w_44070 );
or ( w_44067 , \8025_b0 , \8026_b0 );
not ( \8026_b0 , w_44071 );
and ( w_44071 , w_44070 , \8026_b1 );
or ( \8032_b1 , \8029_b1 , w_44074 );
or ( \8032_b0 , \8029_b0 , w_44073 );
not ( w_44073 , w_44075 );
and ( w_44075 , w_44074 , w_44072 );
or ( w_44072 , \8030_b1 , w_44076 );
or ( w_44073 , \8030_b0 , \8031_b0 );
not ( \8031_b0 , w_44077 );
and ( w_44077 , w_44076 , \8031_b1 );
or ( \8040_b1 , \8037_b1 , w_44080 );
or ( \8040_b0 , \8037_b0 , w_44079 );
not ( w_44079 , w_44081 );
and ( w_44081 , w_44080 , w_44078 );
or ( w_44078 , \8038_b1 , w_44082 );
or ( w_44079 , \8038_b0 , \8039_b0 );
not ( \8039_b0 , w_44083 );
and ( w_44083 , w_44082 , \8039_b1 );
or ( \8046_b1 , \8043_b1 , w_44086 );
or ( \8046_b0 , \8043_b0 , w_44085 );
not ( w_44085 , w_44087 );
and ( w_44087 , w_44086 , w_44084 );
or ( w_44084 , \8044_b1 , w_44088 );
or ( w_44085 , \8044_b0 , \8045_b0 );
not ( \8045_b0 , w_44089 );
and ( w_44089 , w_44088 , \8045_b1 );
or ( \8050_b1 , \8047_b1 , w_44092 );
or ( \8050_b0 , \8047_b0 , w_44091 );
not ( w_44091 , w_44093 );
and ( w_44093 , w_44092 , w_44090 );
or ( w_44090 , \8048_b1 , w_44094 );
or ( w_44091 , \8048_b0 , \8049_b0 );
not ( \8049_b0 , w_44095 );
and ( w_44095 , w_44094 , \8049_b1 );
or ( \8054_b1 , \8051_b1 , w_44098 );
or ( \8054_b0 , \8051_b0 , w_44097 );
not ( w_44097 , w_44099 );
and ( w_44099 , w_44098 , w_44096 );
or ( w_44096 , \8052_b1 , w_44100 );
or ( w_44097 , \8052_b0 , \8053_b0 );
not ( \8053_b0 , w_44101 );
and ( w_44101 , w_44100 , \8053_b1 );
or ( \8062_b1 , \8059_b1 , w_44104 );
or ( \8062_b0 , \8059_b0 , w_44103 );
not ( w_44103 , w_44105 );
and ( w_44105 , w_44104 , w_44102 );
or ( w_44102 , \8060_b1 , w_44106 );
or ( w_44103 , \8060_b0 , \8061_b0 );
not ( \8061_b0 , w_44107 );
and ( w_44107 , w_44106 , \8061_b1 );
or ( \8066_b1 , \8063_b1 , w_44110 );
or ( \8066_b0 , \8063_b0 , w_44109 );
not ( w_44109 , w_44111 );
and ( w_44111 , w_44110 , w_44108 );
or ( w_44108 , \8064_b1 , w_44112 );
or ( w_44109 , \8064_b0 , \8065_b0 );
not ( \8065_b0 , w_44113 );
and ( w_44113 , w_44112 , \8065_b1 );
or ( \8071_b1 , \8068_b1 , w_44116 );
or ( \8071_b0 , \8068_b0 , w_44115 );
not ( w_44115 , w_44117 );
and ( w_44117 , w_44116 , w_44114 );
or ( w_44114 , \8069_b1 , w_44118 );
or ( w_44115 , \8069_b0 , \8070_b0 );
not ( \8070_b0 , w_44119 );
and ( w_44119 , w_44118 , \8070_b1 );
or ( \8075_b1 , \8072_b1 , w_44122 );
or ( \8075_b0 , \8072_b0 , w_44121 );
not ( w_44121 , w_44123 );
and ( w_44123 , w_44122 , w_44120 );
or ( w_44120 , \8073_b1 , w_44124 );
or ( w_44121 , \8073_b0 , \8074_b0 );
not ( \8074_b0 , w_44125 );
and ( w_44125 , w_44124 , \8074_b1 );
or ( \8080_b1 , \8077_b1 , w_44128 );
or ( \8080_b0 , \8077_b0 , w_44127 );
not ( w_44127 , w_44129 );
and ( w_44129 , w_44128 , w_44126 );
or ( w_44126 , \8078_b1 , w_44130 );
or ( w_44127 , \8078_b0 , \8079_b0 );
not ( \8079_b0 , w_44131 );
and ( w_44131 , w_44130 , \8079_b1 );
or ( \8166_b1 , \8163_b1 , w_44134 );
or ( \8166_b0 , \8163_b0 , w_44133 );
not ( w_44133 , w_44135 );
and ( w_44135 , w_44134 , w_44132 );
or ( w_44132 , \8164_b1 , w_44136 );
or ( w_44133 , \8164_b0 , \8165_b0 );
not ( \8165_b0 , w_44137 );
and ( w_44137 , w_44136 , \8165_b1 );
or ( \8170_b1 , \8167_b1 , w_44140 );
or ( \8170_b0 , \8167_b0 , w_44139 );
not ( w_44139 , w_44141 );
and ( w_44141 , w_44140 , w_44138 );
or ( w_44138 , \8168_b1 , w_44142 );
or ( w_44139 , \8168_b0 , \8169_b0 );
not ( \8169_b0 , w_44143 );
and ( w_44143 , w_44142 , \8169_b1 );
or ( \8175_b1 , \8172_b1 , w_44146 );
or ( \8175_b0 , \8172_b0 , w_44145 );
not ( w_44145 , w_44147 );
and ( w_44147 , w_44146 , w_44144 );
or ( w_44144 , \8173_b1 , w_44148 );
or ( w_44145 , \8173_b0 , \8174_b0 );
not ( \8174_b0 , w_44149 );
and ( w_44149 , w_44148 , \8174_b1 );
or ( \8182_b1 , \8179_b1 , w_44152 );
or ( \8182_b0 , \8179_b0 , w_44151 );
not ( w_44151 , w_44153 );
and ( w_44153 , w_44152 , w_44150 );
or ( w_44150 , \8180_b1 , w_44154 );
or ( w_44151 , \8180_b0 , \8181_b0 );
not ( \8181_b0 , w_44155 );
and ( w_44155 , w_44154 , \8181_b1 );
or ( \8186_b1 , \8183_b1 , w_44158 );
or ( \8186_b0 , \8183_b0 , w_44157 );
not ( w_44157 , w_44159 );
and ( w_44159 , w_44158 , w_44156 );
or ( w_44156 , \8184_b1 , w_44160 );
or ( w_44157 , \8184_b0 , \8185_b0 );
not ( \8185_b0 , w_44161 );
and ( w_44161 , w_44160 , \8185_b1 );
or ( \8191_b1 , \8188_b1 , w_44164 );
or ( \8191_b0 , \8188_b0 , w_44163 );
not ( w_44163 , w_44165 );
and ( w_44165 , w_44164 , w_44162 );
or ( w_44162 , \8189_b1 , w_44166 );
or ( w_44163 , \8189_b0 , \8190_b0 );
not ( \8190_b0 , w_44167 );
and ( w_44167 , w_44166 , \8190_b1 );
or ( \8199_b1 , \8196_b1 , w_44170 );
or ( \8199_b0 , \8196_b0 , w_44169 );
not ( w_44169 , w_44171 );
and ( w_44171 , w_44170 , w_44168 );
or ( w_44168 , \8197_b1 , w_44172 );
or ( w_44169 , \8197_b0 , \8198_b0 );
not ( \8198_b0 , w_44173 );
and ( w_44173 , w_44172 , \8198_b1 );
or ( \8204_b1 , \8201_b1 , w_44176 );
or ( \8204_b0 , \8201_b0 , w_44175 );
not ( w_44175 , w_44177 );
and ( w_44177 , w_44176 , w_44174 );
or ( w_44174 , \8202_b1 , w_44178 );
or ( w_44175 , \8202_b0 , \8203_b0 );
not ( \8203_b0 , w_44179 );
and ( w_44179 , w_44178 , \8203_b1 );
or ( \8208_b1 , \8205_b1 , w_44182 );
or ( \8208_b0 , \8205_b0 , w_44181 );
not ( w_44181 , w_44183 );
and ( w_44183 , w_44182 , w_44180 );
or ( w_44180 , \8206_b1 , w_44184 );
or ( w_44181 , \8206_b0 , \8207_b0 );
not ( \8207_b0 , w_44185 );
and ( w_44185 , w_44184 , \8207_b1 );
or ( \8212_b1 , \8209_b1 , w_44188 );
or ( \8212_b0 , \8209_b0 , w_44187 );
not ( w_44187 , w_44189 );
and ( w_44189 , w_44188 , w_44186 );
or ( w_44186 , \8210_b1 , w_44190 );
or ( w_44187 , \8210_b0 , \8211_b0 );
not ( \8211_b0 , w_44191 );
and ( w_44191 , w_44190 , \8211_b1 );
or ( \8217_b1 , \8214_b1 , w_44194 );
or ( \8217_b0 , \8214_b0 , w_44193 );
not ( w_44193 , w_44195 );
and ( w_44195 , w_44194 , w_44192 );
or ( w_44192 , \8215_b1 , w_44196 );
or ( w_44193 , \8215_b0 , \8216_b0 );
not ( \8216_b0 , w_44197 );
and ( w_44197 , w_44196 , \8216_b1 );
or ( \8222_b1 , \8219_b1 , w_44200 );
or ( \8222_b0 , \8219_b0 , w_44199 );
not ( w_44199 , w_44201 );
and ( w_44201 , w_44200 , w_44198 );
or ( w_44198 , \8220_b1 , w_44202 );
or ( w_44199 , \8220_b0 , \8221_b0 );
not ( \8221_b0 , w_44203 );
and ( w_44203 , w_44202 , \8221_b1 );
or ( \8226_b1 , \8223_b1 , w_44206 );
or ( \8226_b0 , \8223_b0 , w_44205 );
not ( w_44205 , w_44207 );
and ( w_44207 , w_44206 , w_44204 );
or ( w_44204 , \8224_b1 , w_44208 );
or ( w_44205 , \8224_b0 , \8225_b0 );
not ( \8225_b0 , w_44209 );
and ( w_44209 , w_44208 , \8225_b1 );
or ( \8258_b1 , \8255_b1 , w_44212 );
or ( \8258_b0 , \8255_b0 , w_44211 );
not ( w_44211 , w_44213 );
and ( w_44213 , w_44212 , w_44210 );
or ( w_44210 , \8256_b1 , w_44214 );
or ( w_44211 , \8256_b0 , \8257_b0 );
not ( \8257_b0 , w_44215 );
and ( w_44215 , w_44214 , \8257_b1 );
or ( \8262_b1 , \8259_b1 , w_44218 );
or ( \8262_b0 , \8259_b0 , w_44217 );
not ( w_44217 , w_44219 );
and ( w_44219 , w_44218 , w_44216 );
or ( w_44216 , \8260_b1 , w_44220 );
or ( w_44217 , \8260_b0 , \8261_b0 );
not ( \8261_b0 , w_44221 );
and ( w_44221 , w_44220 , \8261_b1 );
or ( \8270_b1 , \8267_b1 , w_44224 );
or ( \8270_b0 , \8267_b0 , w_44223 );
not ( w_44223 , w_44225 );
and ( w_44225 , w_44224 , w_44222 );
or ( w_44222 , \8268_b1 , w_44226 );
or ( w_44223 , \8268_b0 , \8269_b0 );
not ( \8269_b0 , w_44227 );
and ( w_44227 , w_44226 , \8269_b1 );
or ( \8274_b1 , \8271_b1 , w_44230 );
or ( \8274_b0 , \8271_b0 , w_44229 );
not ( w_44229 , w_44231 );
and ( w_44231 , w_44230 , w_44228 );
or ( w_44228 , \8272_b1 , w_44232 );
or ( w_44229 , \8272_b0 , \8273_b0 );
not ( \8273_b0 , w_44233 );
and ( w_44233 , w_44232 , \8273_b1 );
or ( \8279_b1 , \8276_b1 , w_44236 );
or ( \8279_b0 , \8276_b0 , w_44235 );
not ( w_44235 , w_44237 );
and ( w_44237 , w_44236 , w_44234 );
or ( w_44234 , \8277_b1 , w_44238 );
or ( w_44235 , \8277_b0 , \8278_b0 );
not ( \8278_b0 , w_44239 );
and ( w_44239 , w_44238 , \8278_b1 );
or ( \8288_b1 , \8285_b1 , w_44242 );
or ( \8288_b0 , \8285_b0 , w_44241 );
not ( w_44241 , w_44243 );
and ( w_44243 , w_44242 , w_44240 );
or ( w_44240 , \8286_b1 , w_44244 );
or ( w_44241 , \8286_b0 , \8287_b0 );
not ( \8287_b0 , w_44245 );
and ( w_44245 , w_44244 , \8287_b1 );
or ( \8292_b1 , \8289_b1 , w_44248 );
or ( \8292_b0 , \8289_b0 , w_44247 );
not ( w_44247 , w_44249 );
and ( w_44249 , w_44248 , w_44246 );
or ( w_44246 , \8290_b1 , w_44250 );
or ( w_44247 , \8290_b0 , \8291_b0 );
not ( \8291_b0 , w_44251 );
and ( w_44251 , w_44250 , \8291_b1 );
or ( \8297_b1 , \8294_b1 , w_44254 );
or ( \8297_b0 , \8294_b0 , w_44253 );
not ( w_44253 , w_44255 );
and ( w_44255 , w_44254 , w_44252 );
or ( w_44252 , \8295_b1 , w_44256 );
or ( w_44253 , \8295_b0 , \8296_b0 );
not ( \8296_b0 , w_44257 );
and ( w_44257 , w_44256 , \8296_b1 );
or ( \8358_b1 , \8355_b1 , w_44260 );
or ( \8358_b0 , \8355_b0 , w_44259 );
not ( w_44259 , w_44261 );
and ( w_44261 , w_44260 , w_44258 );
or ( w_44258 , \8356_b1 , w_44262 );
or ( w_44259 , \8356_b0 , \8357_b0 );
not ( \8357_b0 , w_44263 );
and ( w_44263 , w_44262 , \8357_b1 );
or ( \8365_b1 , \8362_b1 , w_44266 );
or ( \8365_b0 , \8362_b0 , w_44265 );
not ( w_44265 , w_44267 );
and ( w_44267 , w_44266 , w_44264 );
or ( w_44264 , \8363_b1 , w_44268 );
or ( w_44265 , \8363_b0 , \8364_b0 );
not ( \8364_b0 , w_44269 );
and ( w_44269 , w_44268 , \8364_b1 );
or ( \8371_b1 , \8368_b1 , w_44272 );
or ( \8371_b0 , \8368_b0 , w_44271 );
not ( w_44271 , w_44273 );
and ( w_44273 , w_44272 , w_44270 );
or ( w_44270 , \8369_b1 , w_44274 );
or ( w_44271 , \8369_b0 , \8370_b0 );
not ( \8370_b0 , w_44275 );
and ( w_44275 , w_44274 , \8370_b1 );
or ( \8375_b1 , \8372_b1 , w_44278 );
or ( \8375_b0 , \8372_b0 , w_44277 );
not ( w_44277 , w_44279 );
and ( w_44279 , w_44278 , w_44276 );
or ( w_44276 , \8373_b1 , w_44280 );
or ( w_44277 , \8373_b0 , \8374_b0 );
not ( \8374_b0 , w_44281 );
and ( w_44281 , w_44280 , \8374_b1 );
or ( \8379_b1 , \8376_b1 , w_44284 );
or ( \8379_b0 , \8376_b0 , w_44283 );
not ( w_44283 , w_44285 );
and ( w_44285 , w_44284 , w_44282 );
or ( w_44282 , \8377_b1 , w_44286 );
or ( w_44283 , \8377_b0 , \8378_b0 );
not ( \8378_b0 , w_44287 );
and ( w_44287 , w_44286 , \8378_b1 );
or ( \8384_b1 , \8381_b1 , w_44290 );
or ( \8384_b0 , \8381_b0 , w_44289 );
not ( w_44289 , w_44291 );
and ( w_44291 , w_44290 , w_44288 );
or ( w_44288 , \8382_b1 , w_44292 );
or ( w_44289 , \8382_b0 , \8383_b0 );
not ( \8383_b0 , w_44293 );
and ( w_44293 , w_44292 , \8383_b1 );
or ( \8389_b1 , \8386_b1 , w_44296 );
or ( \8389_b0 , \8386_b0 , w_44295 );
not ( w_44295 , w_44297 );
and ( w_44297 , w_44296 , w_44294 );
or ( w_44294 , \8387_b1 , w_44298 );
or ( w_44295 , \8387_b0 , \8388_b0 );
not ( \8388_b0 , w_44299 );
and ( w_44299 , w_44298 , \8388_b1 );
or ( \8393_b1 , \8390_b1 , w_44302 );
or ( \8393_b0 , \8390_b0 , w_44301 );
not ( w_44301 , w_44303 );
and ( w_44303 , w_44302 , w_44300 );
or ( w_44300 , \8391_b1 , w_44304 );
or ( w_44301 , \8391_b0 , \8392_b0 );
not ( \8392_b0 , w_44305 );
and ( w_44305 , w_44304 , \8392_b1 );
or ( \8398_b1 , \8395_b1 , w_44308 );
or ( \8398_b0 , \8395_b0 , w_44307 );
not ( w_44307 , w_44309 );
and ( w_44309 , w_44308 , w_44306 );
or ( w_44306 , \8396_b1 , w_44310 );
or ( w_44307 , \8396_b0 , \8397_b0 );
not ( \8397_b0 , w_44311 );
and ( w_44311 , w_44310 , \8397_b1 );
or ( \8404_b1 , \8401_b1 , w_44314 );
or ( \8404_b0 , \8401_b0 , w_44313 );
not ( w_44313 , w_44315 );
and ( w_44315 , w_44314 , w_44312 );
or ( w_44312 , \8402_b1 , w_44316 );
or ( w_44313 , \8402_b0 , \8403_b0 );
not ( \8403_b0 , w_44317 );
and ( w_44317 , w_44316 , \8403_b1 );
or ( \8491_b1 , \8488_b1 , w_44320 );
or ( \8491_b0 , \8488_b0 , w_44319 );
not ( w_44319 , w_44321 );
and ( w_44321 , w_44320 , w_44318 );
or ( w_44318 , \8489_b1 , w_44322 );
or ( w_44319 , \8489_b0 , \8490_b0 );
not ( \8490_b0 , w_44323 );
and ( w_44323 , w_44322 , \8490_b1 );
or ( \8495_b1 , \8492_b1 , w_44326 );
or ( \8495_b0 , \8492_b0 , w_44325 );
not ( w_44325 , w_44327 );
and ( w_44327 , w_44326 , w_44324 );
or ( w_44324 , \8493_b1 , w_44328 );
or ( w_44325 , \8493_b0 , \8494_b0 );
not ( \8494_b0 , w_44329 );
and ( w_44329 , w_44328 , \8494_b1 );
or ( \8504_b1 , \8501_b1 , w_44332 );
or ( \8504_b0 , \8501_b0 , w_44331 );
not ( w_44331 , w_44333 );
and ( w_44333 , w_44332 , w_44330 );
or ( w_44330 , \8502_b1 , w_44334 );
or ( w_44331 , \8502_b0 , \8503_b0 );
not ( \8503_b0 , w_44335 );
and ( w_44335 , w_44334 , \8503_b1 );
or ( \8508_b1 , \8505_b1 , w_44338 );
or ( \8508_b0 , \8505_b0 , w_44337 );
not ( w_44337 , w_44339 );
and ( w_44339 , w_44338 , w_44336 );
or ( w_44336 , \8506_b1 , w_44340 );
or ( w_44337 , \8506_b0 , \8507_b0 );
not ( \8507_b0 , w_44341 );
and ( w_44341 , w_44340 , \8507_b1 );
or ( \8513_b1 , \8510_b1 , w_44344 );
or ( \8513_b0 , \8510_b0 , w_44343 );
not ( w_44343 , w_44345 );
and ( w_44345 , w_44344 , w_44342 );
or ( w_44342 , \8511_b1 , w_44346 );
or ( w_44343 , \8511_b0 , \8512_b0 );
not ( \8512_b0 , w_44347 );
and ( w_44347 , w_44346 , \8512_b1 );
or ( \8520_b1 , \8517_b1 , w_44350 );
or ( \8520_b0 , \8517_b0 , w_44349 );
not ( w_44349 , w_44351 );
and ( w_44351 , w_44350 , w_44348 );
or ( w_44348 , \8518_b1 , w_44352 );
or ( w_44349 , \8518_b0 , \8519_b0 );
not ( \8519_b0 , w_44353 );
and ( w_44353 , w_44352 , \8519_b1 );
or ( \8525_b1 , \8522_b1 , w_44356 );
or ( \8525_b0 , \8522_b0 , w_44355 );
not ( w_44355 , w_44357 );
and ( w_44357 , w_44356 , w_44354 );
or ( w_44354 , \8523_b1 , w_44358 );
or ( w_44355 , \8523_b0 , \8524_b0 );
not ( \8524_b0 , w_44359 );
and ( w_44359 , w_44358 , \8524_b1 );
or ( \8529_b1 , \8526_b1 , w_44362 );
or ( \8529_b0 , \8526_b0 , w_44361 );
not ( w_44361 , w_44363 );
and ( w_44363 , w_44362 , w_44360 );
or ( w_44360 , \8527_b1 , w_44364 );
or ( w_44361 , \8527_b0 , \8528_b0 );
not ( \8528_b0 , w_44365 );
and ( w_44365 , w_44364 , \8528_b1 );
or ( \8533_b1 , \8530_b1 , w_44368 );
or ( \8533_b0 , \8530_b0 , w_44367 );
not ( w_44367 , w_44369 );
and ( w_44369 , w_44368 , w_44366 );
or ( w_44366 , \8531_b1 , w_44370 );
or ( w_44367 , \8531_b0 , \8532_b0 );
not ( \8532_b0 , w_44371 );
and ( w_44371 , w_44370 , \8532_b1 );
or ( \8541_b1 , \8538_b1 , w_44374 );
or ( \8541_b0 , \8538_b0 , w_44373 );
not ( w_44373 , w_44375 );
and ( w_44375 , w_44374 , w_44372 );
or ( w_44372 , \8539_b1 , w_44376 );
or ( w_44373 , \8539_b0 , \8540_b0 );
not ( \8540_b0 , w_44377 );
and ( w_44377 , w_44376 , \8540_b1 );
or ( \8545_b1 , \8542_b1 , w_44380 );
or ( \8545_b0 , \8542_b0 , w_44379 );
not ( w_44379 , w_44381 );
and ( w_44381 , w_44380 , w_44378 );
or ( w_44378 , \8543_b1 , w_44382 );
or ( w_44379 , \8543_b0 , \8544_b0 );
not ( \8544_b0 , w_44383 );
and ( w_44383 , w_44382 , \8544_b1 );
or ( \8577_b1 , \8574_b1 , w_44386 );
or ( \8577_b0 , \8574_b0 , w_44385 );
not ( w_44385 , w_44387 );
and ( w_44387 , w_44386 , w_44384 );
or ( w_44384 , \8575_b1 , w_44388 );
or ( w_44385 , \8575_b0 , \8576_b0 );
not ( \8576_b0 , w_44389 );
and ( w_44389 , w_44388 , \8576_b1 );
or ( \8581_b1 , \8578_b1 , w_44392 );
or ( \8581_b0 , \8578_b0 , w_44391 );
not ( w_44391 , w_44393 );
and ( w_44393 , w_44392 , w_44390 );
or ( w_44390 , \8579_b1 , w_44394 );
or ( w_44391 , \8579_b0 , \8580_b0 );
not ( \8580_b0 , w_44395 );
and ( w_44395 , w_44394 , \8580_b1 );
or ( \8589_b1 , \8586_b1 , w_44398 );
or ( \8589_b0 , \8586_b0 , w_44397 );
not ( w_44397 , w_44399 );
and ( w_44399 , w_44398 , w_44396 );
or ( w_44396 , \8587_b1 , w_44400 );
or ( w_44397 , \8587_b0 , \8588_b0 );
not ( \8588_b0 , w_44401 );
and ( w_44401 , w_44400 , \8588_b1 );
or ( \8593_b1 , \8590_b1 , w_44404 );
or ( \8593_b0 , \8590_b0 , w_44403 );
not ( w_44403 , w_44405 );
and ( w_44405 , w_44404 , w_44402 );
or ( w_44402 , \8591_b1 , w_44406 );
or ( w_44403 , \8591_b0 , \8592_b0 );
not ( \8592_b0 , w_44407 );
and ( w_44407 , w_44406 , \8592_b1 );
or ( \8598_b1 , \8595_b1 , w_44410 );
or ( \8598_b0 , \8595_b0 , w_44409 );
not ( w_44409 , w_44411 );
and ( w_44411 , w_44410 , w_44408 );
or ( w_44408 , \8596_b1 , w_44412 );
or ( w_44409 , \8596_b0 , \8597_b0 );
not ( \8597_b0 , w_44413 );
and ( w_44413 , w_44412 , \8597_b1 );
or ( \8604_b1 , \8601_b1 , w_44416 );
or ( \8604_b0 , \8601_b0 , w_44415 );
not ( w_44415 , w_44417 );
and ( w_44417 , w_44416 , w_44414 );
or ( w_44414 , \8602_b1 , w_44418 );
or ( w_44415 , \8602_b0 , \8603_b0 );
not ( \8603_b0 , w_44419 );
and ( w_44419 , w_44418 , \8603_b1 );
or ( \8664_b1 , \8661_b1 , w_44422 );
or ( \8664_b0 , \8661_b0 , w_44421 );
not ( w_44421 , w_44423 );
and ( w_44423 , w_44422 , w_44420 );
or ( w_44420 , \8662_b1 , w_44424 );
or ( w_44421 , \8662_b0 , \8663_b0 );
not ( \8663_b0 , w_44425 );
and ( w_44425 , w_44424 , \8663_b1 );
or ( \8668_b1 , \8665_b1 , w_44428 );
or ( \8668_b0 , \8665_b0 , w_44427 );
not ( w_44427 , w_44429 );
and ( w_44429 , w_44428 , w_44426 );
or ( w_44426 , \8666_b1 , w_44430 );
or ( w_44427 , \8666_b0 , \8667_b0 );
not ( \8667_b0 , w_44431 );
and ( w_44431 , w_44430 , \8667_b1 );
or ( \8673_b1 , \8670_b1 , w_44434 );
or ( \8673_b0 , \8670_b0 , w_44433 );
not ( w_44433 , w_44435 );
and ( w_44435 , w_44434 , w_44432 );
or ( w_44432 , \8671_b1 , w_44436 );
or ( w_44433 , \8671_b0 , \8672_b0 );
not ( \8672_b0 , w_44437 );
and ( w_44437 , w_44436 , \8672_b1 );
or ( \8681_b1 , \8678_b1 , w_44440 );
or ( \8681_b0 , \8678_b0 , w_44439 );
not ( w_44439 , w_44441 );
and ( w_44441 , w_44440 , w_44438 );
or ( w_44438 , \8679_b1 , w_44442 );
or ( w_44439 , \8679_b0 , \8680_b0 );
not ( \8680_b0 , w_44443 );
and ( w_44443 , w_44442 , \8680_b1 );
or ( \8687_b1 , \8684_b1 , w_44446 );
or ( \8687_b0 , \8684_b0 , w_44445 );
not ( w_44445 , w_44447 );
and ( w_44447 , w_44446 , w_44444 );
or ( w_44444 , \8685_b1 , w_44448 );
or ( w_44445 , \8685_b0 , \8686_b0 );
not ( \8686_b0 , w_44449 );
and ( w_44449 , w_44448 , \8686_b1 );
or ( \8691_b1 , \8688_b1 , w_44452 );
or ( \8691_b0 , \8688_b0 , w_44451 );
not ( w_44451 , w_44453 );
and ( w_44453 , w_44452 , w_44450 );
or ( w_44450 , \8689_b1 , w_44454 );
or ( w_44451 , \8689_b0 , \8690_b0 );
not ( \8690_b0 , w_44455 );
and ( w_44455 , w_44454 , \8690_b1 );
or ( \8695_b1 , \8692_b1 , w_44458 );
or ( \8695_b0 , \8692_b0 , w_44457 );
not ( w_44457 , w_44459 );
and ( w_44459 , w_44458 , w_44456 );
or ( w_44456 , \8693_b1 , w_44460 );
or ( w_44457 , \8693_b0 , \8694_b0 );
not ( \8694_b0 , w_44461 );
and ( w_44461 , w_44460 , \8694_b1 );
or ( \8700_b1 , \8697_b1 , w_44464 );
or ( \8700_b0 , \8697_b0 , w_44463 );
not ( w_44463 , w_44465 );
and ( w_44465 , w_44464 , w_44462 );
or ( w_44462 , \8698_b1 , w_44466 );
or ( w_44463 , \8698_b0 , \8699_b0 );
not ( \8699_b0 , w_44467 );
and ( w_44467 , w_44466 , \8699_b1 );
or ( \8706_b1 , \8703_b1 , w_44470 );
or ( \8706_b0 , \8703_b0 , w_44469 );
not ( w_44469 , w_44471 );
and ( w_44471 , w_44470 , w_44468 );
or ( w_44468 , \8704_b1 , w_44472 );
or ( w_44469 , \8704_b0 , \8705_b0 );
not ( \8705_b0 , w_44473 );
and ( w_44473 , w_44472 , \8705_b1 );
or ( \8710_b1 , \8707_b1 , w_44476 );
or ( \8710_b0 , \8707_b0 , w_44475 );
not ( w_44475 , w_44477 );
and ( w_44477 , w_44476 , w_44474 );
or ( w_44474 , \8708_b1 , w_44478 );
or ( w_44475 , \8708_b0 , \8709_b0 );
not ( \8709_b0 , w_44479 );
and ( w_44479 , w_44478 , \8709_b1 );
or ( \8715_b1 , \8712_b1 , w_44482 );
or ( \8715_b0 , \8712_b0 , w_44481 );
not ( w_44481 , w_44483 );
and ( w_44483 , w_44482 , w_44480 );
or ( w_44480 , \8713_b1 , w_44484 );
or ( w_44481 , \8713_b0 , \8714_b0 );
not ( \8714_b0 , w_44485 );
and ( w_44485 , w_44484 , \8714_b1 );
or ( \8719_b1 , \8716_b1 , w_44488 );
or ( \8719_b0 , \8716_b0 , w_44487 );
not ( w_44487 , w_44489 );
and ( w_44489 , w_44488 , w_44486 );
or ( w_44486 , \8717_b1 , w_44490 );
or ( w_44487 , \8717_b0 , \8718_b0 );
not ( \8718_b0 , w_44491 );
and ( w_44491 , w_44490 , \8718_b1 );
or ( \8724_b1 , \8721_b1 , w_44494 );
or ( \8724_b0 , \8721_b0 , w_44493 );
not ( w_44493 , w_44495 );
and ( w_44495 , w_44494 , w_44492 );
or ( w_44492 , \8722_b1 , w_44496 );
or ( w_44493 , \8722_b0 , \8723_b0 );
not ( \8723_b0 , w_44497 );
and ( w_44497 , w_44496 , \8723_b1 );
or ( \8729_b1 , \8726_b1 , w_44500 );
or ( \8729_b0 , \8726_b0 , w_44499 );
not ( w_44499 , w_44501 );
and ( w_44501 , w_44500 , w_44498 );
or ( w_44498 , \8727_b1 , w_44502 );
or ( w_44499 , \8727_b0 , \8728_b0 );
not ( \8728_b0 , w_44503 );
and ( w_44503 , w_44502 , \8728_b1 );
or ( \8733_b1 , \8730_b1 , w_44506 );
or ( \8733_b0 , \8730_b0 , w_44505 );
not ( w_44505 , w_44507 );
and ( w_44507 , w_44506 , w_44504 );
or ( w_44504 , \8731_b1 , w_44508 );
or ( w_44505 , \8731_b0 , \8732_b0 );
not ( \8732_b0 , w_44509 );
and ( w_44509 , w_44508 , \8732_b1 );
or ( \8738_b1 , \8735_b1 , w_44512 );
or ( \8738_b0 , \8735_b0 , w_44511 );
not ( w_44511 , w_44513 );
and ( w_44513 , w_44512 , w_44510 );
or ( w_44510 , \8736_b1 , w_44514 );
or ( w_44511 , \8736_b0 , \8737_b0 );
not ( \8737_b0 , w_44515 );
and ( w_44515 , w_44514 , \8737_b1 );
or ( \8744_b1 , \8741_b1 , w_44518 );
or ( \8744_b0 , \8741_b0 , w_44517 );
not ( w_44517 , w_44519 );
and ( w_44519 , w_44518 , w_44516 );
or ( w_44516 , \8742_b1 , w_44520 );
or ( w_44517 , \8742_b0 , \8743_b0 );
not ( \8743_b0 , w_44521 );
and ( w_44521 , w_44520 , \8743_b1 );
or ( \8831_b1 , \8828_b1 , w_44524 );
or ( \8831_b0 , \8828_b0 , w_44523 );
not ( w_44523 , w_44525 );
and ( w_44525 , w_44524 , w_44522 );
or ( w_44522 , \8829_b1 , w_44526 );
or ( w_44523 , \8829_b0 , \8830_b0 );
not ( \8830_b0 , w_44527 );
and ( w_44527 , w_44526 , \8830_b1 );
or ( \8835_b1 , \8832_b1 , w_44530 );
or ( \8835_b0 , \8832_b0 , w_44529 );
not ( w_44529 , w_44531 );
and ( w_44531 , w_44530 , w_44528 );
or ( w_44528 , \8833_b1 , w_44532 );
or ( w_44529 , \8833_b0 , \8834_b0 );
not ( \8834_b0 , w_44533 );
and ( w_44533 , w_44532 , \8834_b1 );
or ( \8845_b1 , \8842_b1 , w_44536 );
or ( \8845_b0 , \8842_b0 , w_44535 );
not ( w_44535 , w_44537 );
and ( w_44537 , w_44536 , w_44534 );
or ( w_44534 , \8843_b1 , w_44538 );
or ( w_44535 , \8843_b0 , \8844_b0 );
not ( \8844_b0 , w_44539 );
and ( w_44539 , w_44538 , \8844_b1 );
or ( \8850_b1 , \8847_b1 , w_44542 );
or ( \8850_b0 , \8847_b0 , w_44541 );
not ( w_44541 , w_44543 );
and ( w_44543 , w_44542 , w_44540 );
or ( w_44540 , \8848_b1 , w_44544 );
or ( w_44541 , \8848_b0 , \8849_b0 );
not ( \8849_b0 , w_44545 );
and ( w_44545 , w_44544 , \8849_b1 );
or ( \8854_b1 , \8851_b1 , w_44548 );
or ( \8854_b0 , \8851_b0 , w_44547 );
not ( w_44547 , w_44549 );
and ( w_44549 , w_44548 , w_44546 );
or ( w_44546 , \8852_b1 , w_44550 );
or ( w_44547 , \8852_b0 , \8853_b0 );
not ( \8853_b0 , w_44551 );
and ( w_44551 , w_44550 , \8853_b1 );
or ( \8858_b1 , \8855_b1 , w_44554 );
or ( \8858_b0 , \8855_b0 , w_44553 );
not ( w_44553 , w_44555 );
and ( w_44555 , w_44554 , w_44552 );
or ( w_44552 , \8856_b1 , w_44556 );
or ( w_44553 , \8856_b0 , \8857_b0 );
not ( \8857_b0 , w_44557 );
and ( w_44557 , w_44556 , \8857_b1 );
or ( \8866_b1 , \8863_b1 , w_44560 );
or ( \8866_b0 , \8863_b0 , w_44559 );
not ( w_44559 , w_44561 );
and ( w_44561 , w_44560 , w_44558 );
or ( w_44558 , \8864_b1 , w_44562 );
or ( w_44559 , \8864_b0 , \8865_b0 );
not ( \8865_b0 , w_44563 );
and ( w_44563 , w_44562 , \8865_b1 );
or ( \8870_b1 , \8867_b1 , w_44566 );
or ( \8870_b0 , \8867_b0 , w_44565 );
not ( w_44565 , w_44567 );
and ( w_44567 , w_44566 , w_44564 );
or ( w_44564 , \8868_b1 , w_44568 );
or ( w_44565 , \8868_b0 , \8869_b0 );
not ( \8869_b0 , w_44569 );
and ( w_44569 , w_44568 , \8869_b1 );
or ( \8902_b1 , \8899_b1 , w_44572 );
or ( \8902_b0 , \8899_b0 , w_44571 );
not ( w_44571 , w_44573 );
and ( w_44573 , w_44572 , w_44570 );
or ( w_44570 , \8900_b1 , w_44574 );
or ( w_44571 , \8900_b0 , \8901_b0 );
not ( \8901_b0 , w_44575 );
and ( w_44575 , w_44574 , \8901_b1 );
or ( \8906_b1 , \8903_b1 , w_44578 );
or ( \8906_b0 , \8903_b0 , w_44577 );
not ( w_44577 , w_44579 );
and ( w_44579 , w_44578 , w_44576 );
or ( w_44576 , \8904_b1 , w_44580 );
or ( w_44577 , \8904_b0 , \8905_b0 );
not ( \8905_b0 , w_44581 );
and ( w_44581 , w_44580 , \8905_b1 );
or ( \8914_b1 , \8911_b1 , w_44584 );
or ( \8914_b0 , \8911_b0 , w_44583 );
not ( w_44583 , w_44585 );
and ( w_44585 , w_44584 , w_44582 );
or ( w_44582 , \8912_b1 , w_44586 );
or ( w_44583 , \8912_b0 , \8913_b0 );
not ( \8913_b0 , w_44587 );
and ( w_44587 , w_44586 , \8913_b1 );
or ( \8918_b1 , \8915_b1 , w_44590 );
or ( \8918_b0 , \8915_b0 , w_44589 );
not ( w_44589 , w_44591 );
and ( w_44591 , w_44590 , w_44588 );
or ( w_44588 , \8916_b1 , w_44592 );
or ( w_44589 , \8916_b0 , \8917_b0 );
not ( \8917_b0 , w_44593 );
and ( w_44593 , w_44592 , \8917_b1 );
or ( \8923_b1 , \8920_b1 , w_44596 );
or ( \8923_b0 , \8920_b0 , w_44595 );
not ( w_44595 , w_44597 );
and ( w_44597 , w_44596 , w_44594 );
or ( w_44594 , \8921_b1 , w_44598 );
or ( w_44595 , \8921_b0 , \8922_b0 );
not ( \8922_b0 , w_44599 );
and ( w_44599 , w_44598 , \8922_b1 );
or ( \8929_b1 , \8926_b1 , w_44602 );
or ( \8929_b0 , \8926_b0 , w_44601 );
not ( w_44601 , w_44603 );
and ( w_44603 , w_44602 , w_44600 );
or ( w_44600 , \8927_b1 , w_44604 );
or ( w_44601 , \8927_b0 , \8928_b0 );
not ( \8928_b0 , w_44605 );
and ( w_44605 , w_44604 , \8928_b1 );
or ( \8989_b1 , \8986_b1 , w_44608 );
or ( \8989_b0 , \8986_b0 , w_44607 );
not ( w_44607 , w_44609 );
and ( w_44609 , w_44608 , w_44606 );
or ( w_44606 , \8987_b1 , w_44610 );
or ( w_44607 , \8987_b0 , \8988_b0 );
not ( \8988_b0 , w_44611 );
and ( w_44611 , w_44610 , \8988_b1 );
or ( \8993_b1 , \8990_b1 , w_44614 );
or ( \8993_b0 , \8990_b0 , w_44613 );
not ( w_44613 , w_44615 );
and ( w_44615 , w_44614 , w_44612 );
or ( w_44612 , \8991_b1 , w_44616 );
or ( w_44613 , \8991_b0 , \8992_b0 );
not ( \8992_b0 , w_44617 );
and ( w_44617 , w_44616 , \8992_b1 );
or ( \8998_b1 , \8995_b1 , w_44620 );
or ( \8998_b0 , \8995_b0 , w_44619 );
not ( w_44619 , w_44621 );
and ( w_44621 , w_44620 , w_44618 );
or ( w_44618 , \8996_b1 , w_44622 );
or ( w_44619 , \8996_b0 , \8997_b0 );
not ( \8997_b0 , w_44623 );
and ( w_44623 , w_44622 , \8997_b1 );
or ( \9006_b1 , \9003_b1 , w_44626 );
or ( \9006_b0 , \9003_b0 , w_44625 );
not ( w_44625 , w_44627 );
and ( w_44627 , w_44626 , w_44624 );
or ( w_44624 , \9004_b1 , w_44628 );
or ( w_44625 , \9004_b0 , \9005_b0 );
not ( \9005_b0 , w_44629 );
and ( w_44629 , w_44628 , \9005_b1 );
or ( \9014_b1 , \9011_b1 , w_44632 );
or ( \9014_b0 , \9011_b0 , w_44631 );
not ( w_44631 , w_44633 );
and ( w_44633 , w_44632 , w_44630 );
or ( w_44630 , \9012_b1 , w_44634 );
or ( w_44631 , \9012_b0 , \9013_b0 );
not ( \9013_b0 , w_44635 );
and ( w_44635 , w_44634 , \9013_b1 );
or ( \9018_b1 , \9015_b1 , w_44638 );
or ( \9018_b0 , \9015_b0 , w_44637 );
not ( w_44637 , w_44639 );
and ( w_44639 , w_44638 , w_44636 );
or ( w_44636 , \9016_b1 , w_44640 );
or ( w_44637 , \9016_b0 , \9017_b0 );
not ( \9017_b0 , w_44641 );
and ( w_44641 , w_44640 , \9017_b1 );
or ( \9022_b1 , \9019_b1 , w_44644 );
or ( \9022_b0 , \9019_b0 , w_44643 );
not ( w_44643 , w_44645 );
and ( w_44645 , w_44644 , w_44642 );
or ( w_44642 , \9020_b1 , w_44646 );
or ( w_44643 , \9020_b0 , \9021_b0 );
not ( \9021_b0 , w_44647 );
and ( w_44647 , w_44646 , \9021_b1 );
or ( \9027_b1 , \9024_b1 , w_44650 );
or ( \9027_b0 , \9024_b0 , w_44649 );
not ( w_44649 , w_44651 );
and ( w_44651 , w_44650 , w_44648 );
or ( w_44648 , \9025_b1 , w_44652 );
or ( w_44649 , \9025_b0 , \9026_b0 );
not ( \9026_b0 , w_44653 );
and ( w_44653 , w_44652 , \9026_b1 );
or ( \9033_b1 , \9030_b1 , w_44656 );
or ( \9033_b0 , \9030_b0 , w_44655 );
not ( w_44655 , w_44657 );
and ( w_44657 , w_44656 , w_44654 );
or ( w_44654 , \9031_b1 , w_44658 );
or ( w_44655 , \9031_b0 , \9032_b0 );
not ( \9032_b0 , w_44659 );
and ( w_44659 , w_44658 , \9032_b1 );
or ( \9037_b1 , \9034_b1 , w_44662 );
or ( \9037_b0 , \9034_b0 , w_44661 );
not ( w_44661 , w_44663 );
and ( w_44663 , w_44662 , w_44660 );
or ( w_44660 , \9035_b1 , w_44664 );
or ( w_44661 , \9035_b0 , \9036_b0 );
not ( \9036_b0 , w_44665 );
and ( w_44665 , w_44664 , \9036_b1 );
or ( \9042_b1 , \9039_b1 , w_44668 );
or ( \9042_b0 , \9039_b0 , w_44667 );
not ( w_44667 , w_44669 );
and ( w_44669 , w_44668 , w_44666 );
or ( w_44666 , \9040_b1 , w_44670 );
or ( w_44667 , \9040_b0 , \9041_b0 );
not ( \9041_b0 , w_44671 );
and ( w_44671 , w_44670 , \9041_b1 );
or ( \9046_b1 , \9043_b1 , w_44674 );
or ( \9046_b0 , \9043_b0 , w_44673 );
not ( w_44673 , w_44675 );
and ( w_44675 , w_44674 , w_44672 );
or ( w_44672 , \9044_b1 , w_44676 );
or ( w_44673 , \9044_b0 , \9045_b0 );
not ( \9045_b0 , w_44677 );
and ( w_44677 , w_44676 , \9045_b1 );
or ( \9051_b1 , \9048_b1 , w_44680 );
or ( \9051_b0 , \9048_b0 , w_44679 );
not ( w_44679 , w_44681 );
and ( w_44681 , w_44680 , w_44678 );
or ( w_44678 , \9049_b1 , w_44682 );
or ( w_44679 , \9049_b0 , \9050_b0 );
not ( \9050_b0 , w_44683 );
and ( w_44683 , w_44682 , \9050_b1 );
or ( \9056_b1 , \9053_b1 , w_44686 );
or ( \9056_b0 , \9053_b0 , w_44685 );
not ( w_44685 , w_44687 );
and ( w_44687 , w_44686 , w_44684 );
or ( w_44684 , \9054_b1 , w_44688 );
or ( w_44685 , \9054_b0 , \9055_b0 );
not ( \9055_b0 , w_44689 );
and ( w_44689 , w_44688 , \9055_b1 );
or ( \9060_b1 , \9057_b1 , w_44692 );
or ( \9060_b0 , \9057_b0 , w_44691 );
not ( w_44691 , w_44693 );
and ( w_44693 , w_44692 , w_44690 );
or ( w_44690 , \9058_b1 , w_44694 );
or ( w_44691 , \9058_b0 , \9059_b0 );
not ( \9059_b0 , w_44695 );
and ( w_44695 , w_44694 , \9059_b1 );
or ( \9065_b1 , \9062_b1 , w_44698 );
or ( \9065_b0 , \9062_b0 , w_44697 );
not ( w_44697 , w_44699 );
and ( w_44699 , w_44698 , w_44696 );
or ( w_44696 , \9063_b1 , w_44700 );
or ( w_44697 , \9063_b0 , \9064_b0 );
not ( \9064_b0 , w_44701 );
and ( w_44701 , w_44700 , \9064_b1 );
or ( \9071_b1 , \9068_b1 , w_44704 );
or ( \9071_b0 , \9068_b0 , w_44703 );
not ( w_44703 , w_44705 );
and ( w_44705 , w_44704 , w_44702 );
or ( w_44702 , \9069_b1 , w_44706 );
or ( w_44703 , \9069_b0 , \9070_b0 );
not ( \9070_b0 , w_44707 );
and ( w_44707 , w_44706 , \9070_b1 );
or ( \9158_b1 , \9155_b1 , w_44710 );
or ( \9158_b0 , \9155_b0 , w_44709 );
not ( w_44709 , w_44711 );
and ( w_44711 , w_44710 , w_44708 );
or ( w_44708 , \9156_b1 , w_44712 );
or ( w_44709 , \9156_b0 , \9157_b0 );
not ( \9157_b0 , w_44713 );
and ( w_44713 , w_44712 , \9157_b1 );
or ( \9162_b1 , \9159_b1 , w_44716 );
or ( \9162_b0 , \9159_b0 , w_44715 );
not ( w_44715 , w_44717 );
and ( w_44717 , w_44716 , w_44714 );
or ( w_44714 , \9160_b1 , w_44718 );
or ( w_44715 , \9160_b0 , \9161_b0 );
not ( \9161_b0 , w_44719 );
and ( w_44719 , w_44718 , \9161_b1 );
or ( \9172_b1 , \9169_b1 , w_44722 );
or ( \9172_b0 , \9169_b0 , w_44721 );
not ( w_44721 , w_44723 );
and ( w_44723 , w_44722 , w_44720 );
or ( w_44720 , \9170_b1 , w_44724 );
or ( w_44721 , \9170_b0 , \9171_b0 );
not ( \9171_b0 , w_44725 );
and ( w_44725 , w_44724 , \9171_b1 );
or ( \9177_b1 , \9174_b1 , w_44728 );
or ( \9177_b0 , \9174_b0 , w_44727 );
not ( w_44727 , w_44729 );
and ( w_44729 , w_44728 , w_44726 );
or ( w_44726 , \9175_b1 , w_44730 );
or ( w_44727 , \9175_b0 , \9176_b0 );
not ( \9176_b0 , w_44731 );
and ( w_44731 , w_44730 , \9176_b1 );
or ( \9181_b1 , \9178_b1 , w_44734 );
or ( \9181_b0 , \9178_b0 , w_44733 );
not ( w_44733 , w_44735 );
and ( w_44735 , w_44734 , w_44732 );
or ( w_44732 , \9179_b1 , w_44736 );
or ( w_44733 , \9179_b0 , \9180_b0 );
not ( \9180_b0 , w_44737 );
and ( w_44737 , w_44736 , \9180_b1 );
or ( \9185_b1 , \9182_b1 , w_44740 );
or ( \9185_b0 , \9182_b0 , w_44739 );
not ( w_44739 , w_44741 );
and ( w_44741 , w_44740 , w_44738 );
or ( w_44738 , \9183_b1 , w_44742 );
or ( w_44739 , \9183_b0 , \9184_b0 );
not ( \9184_b0 , w_44743 );
and ( w_44743 , w_44742 , \9184_b1 );
or ( \9193_b1 , \9190_b1 , w_44746 );
or ( \9193_b0 , \9190_b0 , w_44745 );
not ( w_44745 , w_44747 );
and ( w_44747 , w_44746 , w_44744 );
or ( w_44744 , \9191_b1 , w_44748 );
or ( w_44745 , \9191_b0 , \9192_b0 );
not ( \9192_b0 , w_44749 );
and ( w_44749 , w_44748 , \9192_b1 );
or ( \9197_b1 , \9194_b1 , w_44752 );
or ( \9197_b0 , \9194_b0 , w_44751 );
not ( w_44751 , w_44753 );
and ( w_44753 , w_44752 , w_44750 );
or ( w_44750 , \9195_b1 , w_44754 );
or ( w_44751 , \9195_b0 , \9196_b0 );
not ( \9196_b0 , w_44755 );
and ( w_44755 , w_44754 , \9196_b1 );
or ( \9229_b1 , \9226_b1 , w_44758 );
or ( \9229_b0 , \9226_b0 , w_44757 );
not ( w_44757 , w_44759 );
and ( w_44759 , w_44758 , w_44756 );
or ( w_44756 , \9227_b1 , w_44760 );
or ( w_44757 , \9227_b0 , \9228_b0 );
not ( \9228_b0 , w_44761 );
and ( w_44761 , w_44760 , \9228_b1 );
or ( \9233_b1 , \9230_b1 , w_44764 );
or ( \9233_b0 , \9230_b0 , w_44763 );
not ( w_44763 , w_44765 );
and ( w_44765 , w_44764 , w_44762 );
or ( w_44762 , \9231_b1 , w_44766 );
or ( w_44763 , \9231_b0 , \9232_b0 );
not ( \9232_b0 , w_44767 );
and ( w_44767 , w_44766 , \9232_b1 );
or ( \9241_b1 , \9238_b1 , w_44770 );
or ( \9241_b0 , \9238_b0 , w_44769 );
not ( w_44769 , w_44771 );
and ( w_44771 , w_44770 , w_44768 );
or ( w_44768 , \9239_b1 , w_44772 );
or ( w_44769 , \9239_b0 , \9240_b0 );
not ( \9240_b0 , w_44773 );
and ( w_44773 , w_44772 , \9240_b1 );
or ( \9245_b1 , \9242_b1 , w_44776 );
or ( \9245_b0 , \9242_b0 , w_44775 );
not ( w_44775 , w_44777 );
and ( w_44777 , w_44776 , w_44774 );
or ( w_44774 , \9243_b1 , w_44778 );
or ( w_44775 , \9243_b0 , \9244_b0 );
not ( \9244_b0 , w_44779 );
and ( w_44779 , w_44778 , \9244_b1 );
or ( \9250_b1 , \9247_b1 , w_44782 );
or ( \9250_b0 , \9247_b0 , w_44781 );
not ( w_44781 , w_44783 );
and ( w_44783 , w_44782 , w_44780 );
or ( w_44780 , \9248_b1 , w_44784 );
or ( w_44781 , \9248_b0 , \9249_b0 );
not ( \9249_b0 , w_44785 );
and ( w_44785 , w_44784 , \9249_b1 );
or ( \9256_b1 , \9253_b1 , w_44788 );
or ( \9256_b0 , \9253_b0 , w_44787 );
not ( w_44787 , w_44789 );
and ( w_44789 , w_44788 , w_44786 );
or ( w_44786 , \9254_b1 , w_44790 );
or ( w_44787 , \9254_b0 , \9255_b0 );
not ( \9255_b0 , w_44791 );
and ( w_44791 , w_44790 , \9255_b1 );
or ( \9316_b1 , \9313_b1 , w_44794 );
or ( \9316_b0 , \9313_b0 , w_44793 );
not ( w_44793 , w_44795 );
and ( w_44795 , w_44794 , w_44792 );
or ( w_44792 , \9314_b1 , w_44796 );
or ( w_44793 , \9314_b0 , \9315_b0 );
not ( \9315_b0 , w_44797 );
and ( w_44797 , w_44796 , \9315_b1 );
or ( \9320_b1 , \9317_b1 , w_44800 );
or ( \9320_b0 , \9317_b0 , w_44799 );
not ( w_44799 , w_44801 );
and ( w_44801 , w_44800 , w_44798 );
or ( w_44798 , \9318_b1 , w_44802 );
or ( w_44799 , \9318_b0 , \9319_b0 );
not ( \9319_b0 , w_44803 );
and ( w_44803 , w_44802 , \9319_b1 );
or ( \9325_b1 , \9322_b1 , w_44806 );
or ( \9325_b0 , \9322_b0 , w_44805 );
not ( w_44805 , w_44807 );
and ( w_44807 , w_44806 , w_44804 );
or ( w_44804 , \9323_b1 , w_44808 );
or ( w_44805 , \9323_b0 , \9324_b0 );
not ( \9324_b0 , w_44809 );
and ( w_44809 , w_44808 , \9324_b1 );
or ( \9333_b1 , \9330_b1 , w_44812 );
or ( \9333_b0 , \9330_b0 , w_44811 );
not ( w_44811 , w_44813 );
and ( w_44813 , w_44812 , w_44810 );
or ( w_44810 , \9331_b1 , w_44814 );
or ( w_44811 , \9331_b0 , \9332_b0 );
not ( \9332_b0 , w_44815 );
and ( w_44815 , w_44814 , \9332_b1 );
or ( \9339_b1 , \9336_b1 , w_44818 );
or ( \9339_b0 , \9336_b0 , w_44817 );
not ( w_44817 , w_44819 );
and ( w_44819 , w_44818 , w_44816 );
or ( w_44816 , \9337_b1 , w_44820 );
or ( w_44817 , \9337_b0 , \9338_b0 );
not ( \9338_b0 , w_44821 );
and ( w_44821 , w_44820 , \9338_b1 );
or ( \9343_b1 , \9340_b1 , w_44824 );
or ( \9343_b0 , \9340_b0 , w_44823 );
not ( w_44823 , w_44825 );
and ( w_44825 , w_44824 , w_44822 );
or ( w_44822 , \9341_b1 , w_44826 );
or ( w_44823 , \9341_b0 , \9342_b0 );
not ( \9342_b0 , w_44827 );
and ( w_44827 , w_44826 , \9342_b1 );
or ( \9347_b1 , \9344_b1 , w_44830 );
or ( \9347_b0 , \9344_b0 , w_44829 );
not ( w_44829 , w_44831 );
and ( w_44831 , w_44830 , w_44828 );
or ( w_44828 , \9345_b1 , w_44832 );
or ( w_44829 , \9345_b0 , \9346_b0 );
not ( \9346_b0 , w_44833 );
and ( w_44833 , w_44832 , \9346_b1 );
or ( \9352_b1 , \9349_b1 , w_44836 );
or ( \9352_b0 , \9349_b0 , w_44835 );
not ( w_44835 , w_44837 );
and ( w_44837 , w_44836 , w_44834 );
or ( w_44834 , \9350_b1 , w_44838 );
or ( w_44835 , \9350_b0 , \9351_b0 );
not ( \9351_b0 , w_44839 );
and ( w_44839 , w_44838 , \9351_b1 );
or ( \9358_b1 , \9355_b1 , w_44842 );
or ( \9358_b0 , \9355_b0 , w_44841 );
not ( w_44841 , w_44843 );
and ( w_44843 , w_44842 , w_44840 );
or ( w_44840 , \9356_b1 , w_44844 );
or ( w_44841 , \9356_b0 , \9357_b0 );
not ( \9357_b0 , w_44845 );
and ( w_44845 , w_44844 , \9357_b1 );
or ( \9362_b1 , \9359_b1 , w_44848 );
or ( \9362_b0 , \9359_b0 , w_44847 );
not ( w_44847 , w_44849 );
and ( w_44849 , w_44848 , w_44846 );
or ( w_44846 , \9360_b1 , w_44850 );
or ( w_44847 , \9360_b0 , \9361_b0 );
not ( \9361_b0 , w_44851 );
and ( w_44851 , w_44850 , \9361_b1 );
or ( \9367_b1 , \9364_b1 , w_44854 );
or ( \9367_b0 , \9364_b0 , w_44853 );
not ( w_44853 , w_44855 );
and ( w_44855 , w_44854 , w_44852 );
or ( w_44852 , \9365_b1 , w_44856 );
or ( w_44853 , \9365_b0 , \9366_b0 );
not ( \9366_b0 , w_44857 );
and ( w_44857 , w_44856 , \9366_b1 );
or ( \9371_b1 , \9368_b1 , w_44860 );
or ( \9371_b0 , \9368_b0 , w_44859 );
not ( w_44859 , w_44861 );
and ( w_44861 , w_44860 , w_44858 );
or ( w_44858 , \9369_b1 , w_44862 );
or ( w_44859 , \9369_b0 , \9370_b0 );
not ( \9370_b0 , w_44863 );
and ( w_44863 , w_44862 , \9370_b1 );
or ( \9376_b1 , \9373_b1 , w_44866 );
or ( \9376_b0 , \9373_b0 , w_44865 );
not ( w_44865 , w_44867 );
and ( w_44867 , w_44866 , w_44864 );
or ( w_44864 , \9374_b1 , w_44868 );
or ( w_44865 , \9374_b0 , \9375_b0 );
not ( \9375_b0 , w_44869 );
and ( w_44869 , w_44868 , \9375_b1 );
or ( \9381_b1 , \9378_b1 , w_44872 );
or ( \9381_b0 , \9378_b0 , w_44871 );
not ( w_44871 , w_44873 );
and ( w_44873 , w_44872 , w_44870 );
or ( w_44870 , \9379_b1 , w_44874 );
or ( w_44871 , \9379_b0 , \9380_b0 );
not ( \9380_b0 , w_44875 );
and ( w_44875 , w_44874 , \9380_b1 );
or ( \9385_b1 , \9382_b1 , w_44878 );
or ( \9385_b0 , \9382_b0 , w_44877 );
not ( w_44877 , w_44879 );
and ( w_44879 , w_44878 , w_44876 );
or ( w_44876 , \9383_b1 , w_44880 );
or ( w_44877 , \9383_b0 , \9384_b0 );
not ( \9384_b0 , w_44881 );
and ( w_44881 , w_44880 , \9384_b1 );
or ( \9390_b1 , \9387_b1 , w_44884 );
or ( \9390_b0 , \9387_b0 , w_44883 );
not ( w_44883 , w_44885 );
and ( w_44885 , w_44884 , w_44882 );
or ( w_44882 , \9388_b1 , w_44886 );
or ( w_44883 , \9388_b0 , \9389_b0 );
not ( \9389_b0 , w_44887 );
and ( w_44887 , w_44886 , \9389_b1 );
or ( \9396_b1 , \9393_b1 , w_44890 );
or ( \9396_b0 , \9393_b0 , w_44889 );
not ( w_44889 , w_44891 );
and ( w_44891 , w_44890 , w_44888 );
or ( w_44888 , \9394_b1 , w_44892 );
or ( w_44889 , \9394_b0 , \9395_b0 );
not ( \9395_b0 , w_44893 );
and ( w_44893 , w_44892 , \9395_b1 );
or ( \9483_b1 , \9480_b1 , w_44896 );
or ( \9483_b0 , \9480_b0 , w_44895 );
not ( w_44895 , w_44897 );
and ( w_44897 , w_44896 , w_44894 );
or ( w_44894 , \9481_b1 , w_44898 );
or ( w_44895 , \9481_b0 , \9482_b0 );
not ( \9482_b0 , w_44899 );
and ( w_44899 , w_44898 , \9482_b1 );
or ( \9487_b1 , \9484_b1 , w_44902 );
or ( \9487_b0 , \9484_b0 , w_44901 );
not ( w_44901 , w_44903 );
and ( w_44903 , w_44902 , w_44900 );
or ( w_44900 , \9485_b1 , w_44904 );
or ( w_44901 , \9485_b0 , \9486_b0 );
not ( \9486_b0 , w_44905 );
and ( w_44905 , w_44904 , \9486_b1 );
or ( \9497_b1 , \9494_b1 , w_44908 );
or ( \9497_b0 , \9494_b0 , w_44907 );
not ( w_44907 , w_44909 );
and ( w_44909 , w_44908 , w_44906 );
or ( w_44906 , \9495_b1 , w_44910 );
or ( w_44907 , \9495_b0 , \9496_b0 );
not ( \9496_b0 , w_44911 );
and ( w_44911 , w_44910 , \9496_b1 );
or ( \9502_b1 , \9499_b1 , w_44914 );
or ( \9502_b0 , \9499_b0 , w_44913 );
not ( w_44913 , w_44915 );
and ( w_44915 , w_44914 , w_44912 );
or ( w_44912 , \9500_b1 , w_44916 );
or ( w_44913 , \9500_b0 , \9501_b0 );
not ( \9501_b0 , w_44917 );
and ( w_44917 , w_44916 , \9501_b1 );
or ( \9506_b1 , \9503_b1 , w_44920 );
or ( \9506_b0 , \9503_b0 , w_44919 );
not ( w_44919 , w_44921 );
and ( w_44921 , w_44920 , w_44918 );
or ( w_44918 , \9504_b1 , w_44922 );
or ( w_44919 , \9504_b0 , \9505_b0 );
not ( \9505_b0 , w_44923 );
and ( w_44923 , w_44922 , \9505_b1 );
or ( \9510_b1 , \9507_b1 , w_44926 );
or ( \9510_b0 , \9507_b0 , w_44925 );
not ( w_44925 , w_44927 );
and ( w_44927 , w_44926 , w_44924 );
or ( w_44924 , \9508_b1 , w_44928 );
or ( w_44925 , \9508_b0 , \9509_b0 );
not ( \9509_b0 , w_44929 );
and ( w_44929 , w_44928 , \9509_b1 );
or ( \9518_b1 , \9515_b1 , w_44932 );
or ( \9518_b0 , \9515_b0 , w_44931 );
not ( w_44931 , w_44933 );
and ( w_44933 , w_44932 , w_44930 );
or ( w_44930 , \9516_b1 , w_44934 );
or ( w_44931 , \9516_b0 , \9517_b0 );
not ( \9517_b0 , w_44935 );
and ( w_44935 , w_44934 , \9517_b1 );
or ( \9522_b1 , \9519_b1 , w_44938 );
or ( \9522_b0 , \9519_b0 , w_44937 );
not ( w_44937 , w_44939 );
and ( w_44939 , w_44938 , w_44936 );
or ( w_44936 , \9520_b1 , w_44940 );
or ( w_44937 , \9520_b0 , \9521_b0 );
not ( \9521_b0 , w_44941 );
and ( w_44941 , w_44940 , \9521_b1 );
or ( \9554_b1 , \9551_b1 , w_44944 );
or ( \9554_b0 , \9551_b0 , w_44943 );
not ( w_44943 , w_44945 );
and ( w_44945 , w_44944 , w_44942 );
or ( w_44942 , \9552_b1 , w_44946 );
or ( w_44943 , \9552_b0 , \9553_b0 );
not ( \9553_b0 , w_44947 );
and ( w_44947 , w_44946 , \9553_b1 );
or ( \9558_b1 , \9555_b1 , w_44950 );
or ( \9558_b0 , \9555_b0 , w_44949 );
not ( w_44949 , w_44951 );
and ( w_44951 , w_44950 , w_44948 );
or ( w_44948 , \9556_b1 , w_44952 );
or ( w_44949 , \9556_b0 , \9557_b0 );
not ( \9557_b0 , w_44953 );
and ( w_44953 , w_44952 , \9557_b1 );
or ( \9566_b1 , \9563_b1 , w_44956 );
or ( \9566_b0 , \9563_b0 , w_44955 );
not ( w_44955 , w_44957 );
and ( w_44957 , w_44956 , w_44954 );
or ( w_44954 , \9564_b1 , w_44958 );
or ( w_44955 , \9564_b0 , \9565_b0 );
not ( \9565_b0 , w_44959 );
and ( w_44959 , w_44958 , \9565_b1 );
or ( \9570_b1 , \9567_b1 , w_44962 );
or ( \9570_b0 , \9567_b0 , w_44961 );
not ( w_44961 , w_44963 );
and ( w_44963 , w_44962 , w_44960 );
or ( w_44960 , \9568_b1 , w_44964 );
or ( w_44961 , \9568_b0 , \9569_b0 );
not ( \9569_b0 , w_44965 );
and ( w_44965 , w_44964 , \9569_b1 );
or ( \9575_b1 , \9572_b1 , w_44968 );
or ( \9575_b0 , \9572_b0 , w_44967 );
not ( w_44967 , w_44969 );
and ( w_44969 , w_44968 , w_44966 );
or ( w_44966 , \9573_b1 , w_44970 );
or ( w_44967 , \9573_b0 , \9574_b0 );
not ( \9574_b0 , w_44971 );
and ( w_44971 , w_44970 , \9574_b1 );
or ( \9581_b1 , \9578_b1 , w_44974 );
or ( \9581_b0 , \9578_b0 , w_44973 );
not ( w_44973 , w_44975 );
and ( w_44975 , w_44974 , w_44972 );
or ( w_44972 , \9579_b1 , w_44976 );
or ( w_44973 , \9579_b0 , \9580_b0 );
not ( \9580_b0 , w_44977 );
and ( w_44977 , w_44976 , \9580_b1 );
or ( \9641_b1 , \9638_b1 , w_44980 );
or ( \9641_b0 , \9638_b0 , w_44979 );
not ( w_44979 , w_44981 );
and ( w_44981 , w_44980 , w_44978 );
or ( w_44978 , \9639_b1 , w_44982 );
or ( w_44979 , \9639_b0 , \9640_b0 );
not ( \9640_b0 , w_44983 );
and ( w_44983 , w_44982 , \9640_b1 );
or ( \9645_b1 , \9642_b1 , w_44986 );
or ( \9645_b0 , \9642_b0 , w_44985 );
not ( w_44985 , w_44987 );
and ( w_44987 , w_44986 , w_44984 );
or ( w_44984 , \9643_b1 , w_44988 );
or ( w_44985 , \9643_b0 , \9644_b0 );
not ( \9644_b0 , w_44989 );
and ( w_44989 , w_44988 , \9644_b1 );
or ( \9650_b1 , \9647_b1 , w_44992 );
or ( \9650_b0 , \9647_b0 , w_44991 );
not ( w_44991 , w_44993 );
and ( w_44993 , w_44992 , w_44990 );
or ( w_44990 , \9648_b1 , w_44994 );
or ( w_44991 , \9648_b0 , \9649_b0 );
not ( \9649_b0 , w_44995 );
and ( w_44995 , w_44994 , \9649_b1 );
or ( \9658_b1 , \9655_b1 , w_44998 );
or ( \9658_b0 , \9655_b0 , w_44997 );
not ( w_44997 , w_44999 );
and ( w_44999 , w_44998 , w_44996 );
or ( w_44996 , \9656_b1 , w_45000 );
or ( w_44997 , \9656_b0 , \9657_b0 );
not ( \9657_b0 , w_45001 );
and ( w_45001 , w_45000 , \9657_b1 );
or ( \9665_b1 , \9662_b1 , w_45004 );
or ( \9665_b0 , \9662_b0 , w_45003 );
not ( w_45003 , w_45005 );
and ( w_45005 , w_45004 , w_45002 );
or ( w_45002 , \9663_b1 , w_45006 );
or ( w_45003 , \9663_b0 , \9664_b0 );
not ( \9664_b0 , w_45007 );
and ( w_45007 , w_45006 , \9664_b1 );
or ( \9669_b1 , \9666_b1 , w_45010 );
or ( \9669_b0 , \9666_b0 , w_45009 );
not ( w_45009 , w_45011 );
and ( w_45011 , w_45010 , w_45008 );
or ( w_45008 , \9667_b1 , w_45012 );
or ( w_45009 , \9667_b0 , \9668_b0 );
not ( \9668_b0 , w_45013 );
and ( w_45013 , w_45012 , \9668_b1 );
or ( \9673_b1 , \9670_b1 , w_45016 );
or ( \9673_b0 , \9670_b0 , w_45015 );
not ( w_45015 , w_45017 );
and ( w_45017 , w_45016 , w_45014 );
or ( w_45014 , \9671_b1 , w_45018 );
or ( w_45015 , \9671_b0 , \9672_b0 );
not ( \9672_b0 , w_45019 );
and ( w_45019 , w_45018 , \9672_b1 );
or ( \9678_b1 , \9675_b1 , w_45022 );
or ( \9678_b0 , \9675_b0 , w_45021 );
not ( w_45021 , w_45023 );
and ( w_45023 , w_45022 , w_45020 );
or ( w_45020 , \9676_b1 , w_45024 );
or ( w_45021 , \9676_b0 , \9677_b0 );
not ( \9677_b0 , w_45025 );
and ( w_45025 , w_45024 , \9677_b1 );
or ( \9684_b1 , \9681_b1 , w_45028 );
or ( \9684_b0 , \9681_b0 , w_45027 );
not ( w_45027 , w_45029 );
and ( w_45029 , w_45028 , w_45026 );
or ( w_45026 , \9682_b1 , w_45030 );
or ( w_45027 , \9682_b0 , \9683_b0 );
not ( \9683_b0 , w_45031 );
and ( w_45031 , w_45030 , \9683_b1 );
or ( \9688_b1 , \9685_b1 , w_45034 );
or ( \9688_b0 , \9685_b0 , w_45033 );
not ( w_45033 , w_45035 );
and ( w_45035 , w_45034 , w_45032 );
or ( w_45032 , \9686_b1 , w_45036 );
or ( w_45033 , \9686_b0 , \9687_b0 );
not ( \9687_b0 , w_45037 );
and ( w_45037 , w_45036 , \9687_b1 );
or ( \9693_b1 , \9690_b1 , w_45040 );
or ( \9693_b0 , \9690_b0 , w_45039 );
not ( w_45039 , w_45041 );
and ( w_45041 , w_45040 , w_45038 );
or ( w_45038 , \9691_b1 , w_45042 );
or ( w_45039 , \9691_b0 , \9692_b0 );
not ( \9692_b0 , w_45043 );
and ( w_45043 , w_45042 , \9692_b1 );
or ( \9697_b1 , \9694_b1 , w_45046 );
or ( \9697_b0 , \9694_b0 , w_45045 );
not ( w_45045 , w_45047 );
and ( w_45047 , w_45046 , w_45044 );
or ( w_45044 , \9695_b1 , w_45048 );
or ( w_45045 , \9695_b0 , \9696_b0 );
not ( \9696_b0 , w_45049 );
and ( w_45049 , w_45048 , \9696_b1 );
or ( \9702_b1 , \9699_b1 , w_45052 );
or ( \9702_b0 , \9699_b0 , w_45051 );
not ( w_45051 , w_45053 );
and ( w_45053 , w_45052 , w_45050 );
or ( w_45050 , \9700_b1 , w_45054 );
or ( w_45051 , \9700_b0 , \9701_b0 );
not ( \9701_b0 , w_45055 );
and ( w_45055 , w_45054 , \9701_b1 );
or ( \9707_b1 , \9704_b1 , w_45058 );
or ( \9707_b0 , \9704_b0 , w_45057 );
not ( w_45057 , w_45059 );
and ( w_45059 , w_45058 , w_45056 );
or ( w_45056 , \9705_b1 , w_45060 );
or ( w_45057 , \9705_b0 , \9706_b0 );
not ( \9706_b0 , w_45061 );
and ( w_45061 , w_45060 , \9706_b1 );
or ( \9711_b1 , \9708_b1 , w_45064 );
or ( \9711_b0 , \9708_b0 , w_45063 );
not ( w_45063 , w_45065 );
and ( w_45065 , w_45064 , w_45062 );
or ( w_45062 , \9709_b1 , w_45066 );
or ( w_45063 , \9709_b0 , \9710_b0 );
not ( \9710_b0 , w_45067 );
and ( w_45067 , w_45066 , \9710_b1 );
or ( \9716_b1 , \9713_b1 , w_45070 );
or ( \9716_b0 , \9713_b0 , w_45069 );
not ( w_45069 , w_45071 );
and ( w_45071 , w_45070 , w_45068 );
or ( w_45068 , \9714_b1 , w_45072 );
or ( w_45069 , \9714_b0 , \9715_b0 );
not ( \9715_b0 , w_45073 );
and ( w_45073 , w_45072 , \9715_b1 );
or ( \9722_b1 , \9719_b1 , w_45076 );
or ( \9722_b0 , \9719_b0 , w_45075 );
not ( w_45075 , w_45077 );
and ( w_45077 , w_45076 , w_45074 );
or ( w_45074 , \9720_b1 , w_45078 );
or ( w_45075 , \9720_b0 , \9721_b0 );
not ( \9721_b0 , w_45079 );
and ( w_45079 , w_45078 , \9721_b1 );
or ( \9809_b1 , \9806_b1 , w_45082 );
or ( \9809_b0 , \9806_b0 , w_45081 );
not ( w_45081 , w_45083 );
and ( w_45083 , w_45082 , w_45080 );
or ( w_45080 , \9807_b1 , w_45084 );
or ( w_45081 , \9807_b0 , \9808_b0 );
not ( \9808_b0 , w_45085 );
and ( w_45085 , w_45084 , \9808_b1 );
or ( \9813_b1 , \9810_b1 , w_45088 );
or ( \9813_b0 , \9810_b0 , w_45087 );
not ( w_45087 , w_45089 );
and ( w_45089 , w_45088 , w_45086 );
or ( w_45086 , \9811_b1 , w_45090 );
or ( w_45087 , \9811_b0 , \9812_b0 );
not ( \9812_b0 , w_45091 );
and ( w_45091 , w_45090 , \9812_b1 );
or ( \9823_b1 , \9820_b1 , w_45094 );
or ( \9823_b0 , \9820_b0 , w_45093 );
not ( w_45093 , w_45095 );
and ( w_45095 , w_45094 , w_45092 );
or ( w_45092 , \9821_b1 , w_45096 );
or ( w_45093 , \9821_b0 , \9822_b0 );
not ( \9822_b0 , w_45097 );
and ( w_45097 , w_45096 , \9822_b1 );
or ( \9828_b1 , \9825_b1 , w_45100 );
or ( \9828_b0 , \9825_b0 , w_45099 );
not ( w_45099 , w_45101 );
and ( w_45101 , w_45100 , w_45098 );
or ( w_45098 , \9826_b1 , w_45102 );
or ( w_45099 , \9826_b0 , \9827_b0 );
not ( \9827_b0 , w_45103 );
and ( w_45103 , w_45102 , \9827_b1 );
or ( \9832_b1 , \9829_b1 , w_45106 );
or ( \9832_b0 , \9829_b0 , w_45105 );
not ( w_45105 , w_45107 );
and ( w_45107 , w_45106 , w_45104 );
or ( w_45104 , \9830_b1 , w_45108 );
or ( w_45105 , \9830_b0 , \9831_b0 );
not ( \9831_b0 , w_45109 );
and ( w_45109 , w_45108 , \9831_b1 );
or ( \9836_b1 , \9833_b1 , w_45112 );
or ( \9836_b0 , \9833_b0 , w_45111 );
not ( w_45111 , w_45113 );
and ( w_45113 , w_45112 , w_45110 );
or ( w_45110 , \9834_b1 , w_45114 );
or ( w_45111 , \9834_b0 , \9835_b0 );
not ( \9835_b0 , w_45115 );
and ( w_45115 , w_45114 , \9835_b1 );
or ( \9844_b1 , \9841_b1 , w_45118 );
or ( \9844_b0 , \9841_b0 , w_45117 );
not ( w_45117 , w_45119 );
and ( w_45119 , w_45118 , w_45116 );
or ( w_45116 , \9842_b1 , w_45120 );
or ( w_45117 , \9842_b0 , \9843_b0 );
not ( \9843_b0 , w_45121 );
and ( w_45121 , w_45120 , \9843_b1 );
or ( \9848_b1 , \9845_b1 , w_45124 );
or ( \9848_b0 , \9845_b0 , w_45123 );
not ( w_45123 , w_45125 );
and ( w_45125 , w_45124 , w_45122 );
or ( w_45122 , \9846_b1 , w_45126 );
or ( w_45123 , \9846_b0 , \9847_b0 );
not ( \9847_b0 , w_45127 );
and ( w_45127 , w_45126 , \9847_b1 );
or ( \9880_b1 , \9877_b1 , w_45130 );
or ( \9880_b0 , \9877_b0 , w_45129 );
not ( w_45129 , w_45131 );
and ( w_45131 , w_45130 , w_45128 );
or ( w_45128 , \9878_b1 , w_45132 );
or ( w_45129 , \9878_b0 , \9879_b0 );
not ( \9879_b0 , w_45133 );
and ( w_45133 , w_45132 , \9879_b1 );
or ( \9884_b1 , \9881_b1 , w_45136 );
or ( \9884_b0 , \9881_b0 , w_45135 );
not ( w_45135 , w_45137 );
and ( w_45137 , w_45136 , w_45134 );
or ( w_45134 , \9882_b1 , w_45138 );
or ( w_45135 , \9882_b0 , \9883_b0 );
not ( \9883_b0 , w_45139 );
and ( w_45139 , w_45138 , \9883_b1 );
or ( \9892_b1 , \9889_b1 , w_45142 );
or ( \9892_b0 , \9889_b0 , w_45141 );
not ( w_45141 , w_45143 );
and ( w_45143 , w_45142 , w_45140 );
or ( w_45140 , \9890_b1 , w_45144 );
or ( w_45141 , \9890_b0 , \9891_b0 );
not ( \9891_b0 , w_45145 );
and ( w_45145 , w_45144 , \9891_b1 );
or ( \9896_b1 , \9893_b1 , w_45148 );
or ( \9896_b0 , \9893_b0 , w_45147 );
not ( w_45147 , w_45149 );
and ( w_45149 , w_45148 , w_45146 );
or ( w_45146 , \9894_b1 , w_45150 );
or ( w_45147 , \9894_b0 , \9895_b0 );
not ( \9895_b0 , w_45151 );
and ( w_45151 , w_45150 , \9895_b1 );
or ( \9901_b1 , \9898_b1 , w_45154 );
or ( \9901_b0 , \9898_b0 , w_45153 );
not ( w_45153 , w_45155 );
and ( w_45155 , w_45154 , w_45152 );
or ( w_45152 , \9899_b1 , w_45156 );
or ( w_45153 , \9899_b0 , \9900_b0 );
not ( \9900_b0 , w_45157 );
and ( w_45157 , w_45156 , \9900_b1 );
or ( \9907_b1 , \9904_b1 , w_45160 );
or ( \9907_b0 , \9904_b0 , w_45159 );
not ( w_45159 , w_45161 );
and ( w_45161 , w_45160 , w_45158 );
or ( w_45158 , \9905_b1 , w_45162 );
or ( w_45159 , \9905_b0 , \9906_b0 );
not ( \9906_b0 , w_45163 );
and ( w_45163 , w_45162 , \9906_b1 );
or ( \9967_b1 , \9964_b1 , w_45166 );
or ( \9967_b0 , \9964_b0 , w_45165 );
not ( w_45165 , w_45167 );
and ( w_45167 , w_45166 , w_45164 );
or ( w_45164 , \9965_b1 , w_45168 );
or ( w_45165 , \9965_b0 , \9966_b0 );
not ( \9966_b0 , w_45169 );
and ( w_45169 , w_45168 , \9966_b1 );
or ( \9971_b1 , \9968_b1 , w_45172 );
or ( \9971_b0 , \9968_b0 , w_45171 );
not ( w_45171 , w_45173 );
and ( w_45173 , w_45172 , w_45170 );
or ( w_45170 , \9969_b1 , w_45174 );
or ( w_45171 , \9969_b0 , \9970_b0 );
not ( \9970_b0 , w_45175 );
and ( w_45175 , w_45174 , \9970_b1 );
or ( \9976_b1 , \9973_b1 , w_45178 );
or ( \9976_b0 , \9973_b0 , w_45177 );
not ( w_45177 , w_45179 );
and ( w_45179 , w_45178 , w_45176 );
or ( w_45176 , \9974_b1 , w_45180 );
or ( w_45177 , \9974_b0 , \9975_b0 );
not ( \9975_b0 , w_45181 );
and ( w_45181 , w_45180 , \9975_b1 );
or ( \9984_b1 , \9981_b1 , w_45184 );
or ( \9984_b0 , \9981_b0 , w_45183 );
not ( w_45183 , w_45185 );
and ( w_45185 , w_45184 , w_45182 );
or ( w_45182 , \9982_b1 , w_45186 );
or ( w_45183 , \9982_b0 , \9983_b0 );
not ( \9983_b0 , w_45187 );
and ( w_45187 , w_45186 , \9983_b1 );
or ( \9990_b1 , \9987_b1 , w_45190 );
or ( \9990_b0 , \9987_b0 , w_45189 );
not ( w_45189 , w_45191 );
and ( w_45191 , w_45190 , w_45188 );
or ( w_45188 , \9988_b1 , w_45192 );
or ( w_45189 , \9988_b0 , \9989_b0 );
not ( \9989_b0 , w_45193 );
and ( w_45193 , w_45192 , \9989_b1 );
or ( \9994_b1 , \9991_b1 , w_45196 );
or ( \9994_b0 , \9991_b0 , w_45195 );
not ( w_45195 , w_45197 );
and ( w_45197 , w_45196 , w_45194 );
or ( w_45194 , \9992_b1 , w_45198 );
or ( w_45195 , \9992_b0 , \9993_b0 );
not ( \9993_b0 , w_45199 );
and ( w_45199 , w_45198 , \9993_b1 );
or ( \9998_b1 , \9995_b1 , w_45202 );
or ( \9998_b0 , \9995_b0 , w_45201 );
not ( w_45201 , w_45203 );
and ( w_45203 , w_45202 , w_45200 );
or ( w_45200 , \9996_b1 , w_45204 );
or ( w_45201 , \9996_b0 , \9997_b0 );
not ( \9997_b0 , w_45205 );
and ( w_45205 , w_45204 , \9997_b1 );
or ( \10003_b1 , \10000_b1 , w_45208 );
or ( \10003_b0 , \10000_b0 , w_45207 );
not ( w_45207 , w_45209 );
and ( w_45209 , w_45208 , w_45206 );
or ( w_45206 , \10001_b1 , w_45210 );
or ( w_45207 , \10001_b0 , \10002_b0 );
not ( \10002_b0 , w_45211 );
and ( w_45211 , w_45210 , \10002_b1 );
or ( \10009_b1 , \10006_b1 , w_45214 );
or ( \10009_b0 , \10006_b0 , w_45213 );
not ( w_45213 , w_45215 );
and ( w_45215 , w_45214 , w_45212 );
or ( w_45212 , \10007_b1 , w_45216 );
or ( w_45213 , \10007_b0 , \10008_b0 );
not ( \10008_b0 , w_45217 );
and ( w_45217 , w_45216 , \10008_b1 );
or ( \10013_b1 , \10010_b1 , w_45220 );
or ( \10013_b0 , \10010_b0 , w_45219 );
not ( w_45219 , w_45221 );
and ( w_45221 , w_45220 , w_45218 );
or ( w_45218 , \10011_b1 , w_45222 );
or ( w_45219 , \10011_b0 , \10012_b0 );
not ( \10012_b0 , w_45223 );
and ( w_45223 , w_45222 , \10012_b1 );
or ( \10018_b1 , \10015_b1 , w_45226 );
or ( \10018_b0 , \10015_b0 , w_45225 );
not ( w_45225 , w_45227 );
and ( w_45227 , w_45226 , w_45224 );
or ( w_45224 , \10016_b1 , w_45228 );
or ( w_45225 , \10016_b0 , \10017_b0 );
not ( \10017_b0 , w_45229 );
and ( w_45229 , w_45228 , \10017_b1 );
or ( \10022_b1 , \10019_b1 , w_45232 );
or ( \10022_b0 , \10019_b0 , w_45231 );
not ( w_45231 , w_45233 );
and ( w_45233 , w_45232 , w_45230 );
or ( w_45230 , \10020_b1 , w_45234 );
or ( w_45231 , \10020_b0 , \10021_b0 );
not ( \10021_b0 , w_45235 );
and ( w_45235 , w_45234 , \10021_b1 );
or ( \10027_b1 , \10024_b1 , w_45238 );
or ( \10027_b0 , \10024_b0 , w_45237 );
not ( w_45237 , w_45239 );
and ( w_45239 , w_45238 , w_45236 );
or ( w_45236 , \10025_b1 , w_45240 );
or ( w_45237 , \10025_b0 , \10026_b0 );
not ( \10026_b0 , w_45241 );
and ( w_45241 , w_45240 , \10026_b1 );
or ( \10032_b1 , \10029_b1 , w_45244 );
or ( \10032_b0 , \10029_b0 , w_45243 );
not ( w_45243 , w_45245 );
and ( w_45245 , w_45244 , w_45242 );
or ( w_45242 , \10030_b1 , w_45246 );
or ( w_45243 , \10030_b0 , \10031_b0 );
not ( \10031_b0 , w_45247 );
and ( w_45247 , w_45246 , \10031_b1 );
or ( \10036_b1 , \10033_b1 , w_45250 );
or ( \10036_b0 , \10033_b0 , w_45249 );
not ( w_45249 , w_45251 );
and ( w_45251 , w_45250 , w_45248 );
or ( w_45248 , \10034_b1 , w_45252 );
or ( w_45249 , \10034_b0 , \10035_b0 );
not ( \10035_b0 , w_45253 );
and ( w_45253 , w_45252 , \10035_b1 );
or ( \10041_b1 , \10038_b1 , w_45256 );
or ( \10041_b0 , \10038_b0 , w_45255 );
not ( w_45255 , w_45257 );
and ( w_45257 , w_45256 , w_45254 );
or ( w_45254 , \10039_b1 , w_45258 );
or ( w_45255 , \10039_b0 , \10040_b0 );
not ( \10040_b0 , w_45259 );
and ( w_45259 , w_45258 , \10040_b1 );
or ( \10047_b1 , \10044_b1 , w_45262 );
or ( \10047_b0 , \10044_b0 , w_45261 );
not ( w_45261 , w_45263 );
and ( w_45263 , w_45262 , w_45260 );
or ( w_45260 , \10045_b1 , w_45264 );
or ( w_45261 , \10045_b0 , \10046_b0 );
not ( \10046_b0 , w_45265 );
and ( w_45265 , w_45264 , \10046_b1 );
or ( \10134_b1 , \10131_b1 , w_45268 );
or ( \10134_b0 , \10131_b0 , w_45267 );
not ( w_45267 , w_45269 );
and ( w_45269 , w_45268 , w_45266 );
or ( w_45266 , \10132_b1 , w_45270 );
or ( w_45267 , \10132_b0 , \10133_b0 );
not ( \10133_b0 , w_45271 );
and ( w_45271 , w_45270 , \10133_b1 );
or ( \10138_b1 , \10135_b1 , w_45274 );
or ( \10138_b0 , \10135_b0 , w_45273 );
not ( w_45273 , w_45275 );
and ( w_45275 , w_45274 , w_45272 );
or ( w_45272 , \10136_b1 , w_45276 );
or ( w_45273 , \10136_b0 , \10137_b0 );
not ( \10137_b0 , w_45277 );
and ( w_45277 , w_45276 , \10137_b1 );
or ( \10148_b1 , \10145_b1 , w_45280 );
or ( \10148_b0 , \10145_b0 , w_45279 );
not ( w_45279 , w_45281 );
and ( w_45281 , w_45280 , w_45278 );
or ( w_45278 , \10146_b1 , w_45282 );
or ( w_45279 , \10146_b0 , \10147_b0 );
not ( \10147_b0 , w_45283 );
and ( w_45283 , w_45282 , \10147_b1 );
or ( \10153_b1 , \10150_b1 , w_45286 );
or ( \10153_b0 , \10150_b0 , w_45285 );
not ( w_45285 , w_45287 );
and ( w_45287 , w_45286 , w_45284 );
or ( w_45284 , \10151_b1 , w_45288 );
or ( w_45285 , \10151_b0 , \10152_b0 );
not ( \10152_b0 , w_45289 );
and ( w_45289 , w_45288 , \10152_b1 );
or ( \10157_b1 , \10154_b1 , w_45292 );
or ( \10157_b0 , \10154_b0 , w_45291 );
not ( w_45291 , w_45293 );
and ( w_45293 , w_45292 , w_45290 );
or ( w_45290 , \10155_b1 , w_45294 );
or ( w_45291 , \10155_b0 , \10156_b0 );
not ( \10156_b0 , w_45295 );
and ( w_45295 , w_45294 , \10156_b1 );
or ( \10161_b1 , \10158_b1 , w_45298 );
or ( \10161_b0 , \10158_b0 , w_45297 );
not ( w_45297 , w_45299 );
and ( w_45299 , w_45298 , w_45296 );
or ( w_45296 , \10159_b1 , w_45300 );
or ( w_45297 , \10159_b0 , \10160_b0 );
not ( \10160_b0 , w_45301 );
and ( w_45301 , w_45300 , \10160_b1 );
or ( \10169_b1 , \10166_b1 , w_45304 );
or ( \10169_b0 , \10166_b0 , w_45303 );
not ( w_45303 , w_45305 );
and ( w_45305 , w_45304 , w_45302 );
or ( w_45302 , \10167_b1 , w_45306 );
or ( w_45303 , \10167_b0 , \10168_b0 );
not ( \10168_b0 , w_45307 );
and ( w_45307 , w_45306 , \10168_b1 );
or ( \10173_b1 , \10170_b1 , w_45310 );
or ( \10173_b0 , \10170_b0 , w_45309 );
not ( w_45309 , w_45311 );
and ( w_45311 , w_45310 , w_45308 );
or ( w_45308 , \10171_b1 , w_45312 );
or ( w_45309 , \10171_b0 , \10172_b0 );
not ( \10172_b0 , w_45313 );
and ( w_45313 , w_45312 , \10172_b1 );
or ( \10205_b1 , \10202_b1 , w_45316 );
or ( \10205_b0 , \10202_b0 , w_45315 );
not ( w_45315 , w_45317 );
and ( w_45317 , w_45316 , w_45314 );
or ( w_45314 , \10203_b1 , w_45318 );
or ( w_45315 , \10203_b0 , \10204_b0 );
not ( \10204_b0 , w_45319 );
and ( w_45319 , w_45318 , \10204_b1 );
or ( \10209_b1 , \10206_b1 , w_45322 );
or ( \10209_b0 , \10206_b0 , w_45321 );
not ( w_45321 , w_45323 );
and ( w_45323 , w_45322 , w_45320 );
or ( w_45320 , \10207_b1 , w_45324 );
or ( w_45321 , \10207_b0 , \10208_b0 );
not ( \10208_b0 , w_45325 );
and ( w_45325 , w_45324 , \10208_b1 );
or ( \10217_b1 , \10214_b1 , w_45328 );
or ( \10217_b0 , \10214_b0 , w_45327 );
not ( w_45327 , w_45329 );
and ( w_45329 , w_45328 , w_45326 );
or ( w_45326 , \10215_b1 , w_45330 );
or ( w_45327 , \10215_b0 , \10216_b0 );
not ( \10216_b0 , w_45331 );
and ( w_45331 , w_45330 , \10216_b1 );
or ( \10221_b1 , \10218_b1 , w_45334 );
or ( \10221_b0 , \10218_b0 , w_45333 );
not ( w_45333 , w_45335 );
and ( w_45335 , w_45334 , w_45332 );
or ( w_45332 , \10219_b1 , w_45336 );
or ( w_45333 , \10219_b0 , \10220_b0 );
not ( \10220_b0 , w_45337 );
and ( w_45337 , w_45336 , \10220_b1 );
or ( \10226_b1 , \10223_b1 , w_45340 );
or ( \10226_b0 , \10223_b0 , w_45339 );
not ( w_45339 , w_45341 );
and ( w_45341 , w_45340 , w_45338 );
or ( w_45338 , \10224_b1 , w_45342 );
or ( w_45339 , \10224_b0 , \10225_b0 );
not ( \10225_b0 , w_45343 );
and ( w_45343 , w_45342 , \10225_b1 );
or ( \10232_b1 , \10229_b1 , w_45346 );
or ( \10232_b0 , \10229_b0 , w_45345 );
not ( w_45345 , w_45347 );
and ( w_45347 , w_45346 , w_45344 );
or ( w_45344 , \10230_b1 , w_45348 );
or ( w_45345 , \10230_b0 , \10231_b0 );
not ( \10231_b0 , w_45349 );
and ( w_45349 , w_45348 , \10231_b1 );
or ( \10292_b1 , \10289_b1 , w_45352 );
or ( \10292_b0 , \10289_b0 , w_45351 );
not ( w_45351 , w_45353 );
and ( w_45353 , w_45352 , w_45350 );
or ( w_45350 , \10290_b1 , w_45354 );
or ( w_45351 , \10290_b0 , \10291_b0 );
not ( \10291_b0 , w_45355 );
and ( w_45355 , w_45354 , \10291_b1 );
or ( \10296_b1 , \10293_b1 , w_45358 );
or ( \10296_b0 , \10293_b0 , w_45357 );
not ( w_45357 , w_45359 );
and ( w_45359 , w_45358 , w_45356 );
or ( w_45356 , \10294_b1 , w_45360 );
or ( w_45357 , \10294_b0 , \10295_b0 );
not ( \10295_b0 , w_45361 );
and ( w_45361 , w_45360 , \10295_b1 );
or ( \10301_b1 , \10298_b1 , w_45364 );
or ( \10301_b0 , \10298_b0 , w_45363 );
not ( w_45363 , w_45365 );
and ( w_45365 , w_45364 , w_45362 );
or ( w_45362 , \10299_b1 , w_45366 );
or ( w_45363 , \10299_b0 , \10300_b0 );
not ( \10300_b0 , w_45367 );
and ( w_45367 , w_45366 , \10300_b1 );
or ( \10309_b1 , \10306_b1 , w_45370 );
or ( \10309_b0 , \10306_b0 , w_45369 );
not ( w_45369 , w_45371 );
and ( w_45371 , w_45370 , w_45368 );
or ( w_45368 , \10307_b1 , w_45372 );
or ( w_45369 , \10307_b0 , \10308_b0 );
not ( \10308_b0 , w_45373 );
and ( w_45373 , w_45372 , \10308_b1 );
or ( \10318_b1 , \10315_b1 , w_45376 );
or ( \10318_b0 , \10315_b0 , w_45375 );
not ( w_45375 , w_45377 );
and ( w_45377 , w_45376 , w_45374 );
or ( w_45374 , \10316_b1 , w_45378 );
or ( w_45375 , \10316_b0 , \10317_b0 );
not ( \10317_b0 , w_45379 );
and ( w_45379 , w_45378 , \10317_b1 );
or ( \10322_b1 , \10319_b1 , w_45382 );
or ( \10322_b0 , \10319_b0 , w_45381 );
not ( w_45381 , w_45383 );
and ( w_45383 , w_45382 , w_45380 );
or ( w_45380 , \10320_b1 , w_45384 );
or ( w_45381 , \10320_b0 , \10321_b0 );
not ( \10321_b0 , w_45385 );
and ( w_45385 , w_45384 , \10321_b1 );
or ( \10326_b1 , \10323_b1 , w_45388 );
or ( \10326_b0 , \10323_b0 , w_45387 );
not ( w_45387 , w_45389 );
and ( w_45389 , w_45388 , w_45386 );
or ( w_45386 , \10324_b1 , w_45390 );
or ( w_45387 , \10324_b0 , \10325_b0 );
not ( \10325_b0 , w_45391 );
and ( w_45391 , w_45390 , \10325_b1 );
or ( \10331_b1 , \10328_b1 , w_45394 );
or ( \10331_b0 , \10328_b0 , w_45393 );
not ( w_45393 , w_45395 );
and ( w_45395 , w_45394 , w_45392 );
or ( w_45392 , \10329_b1 , w_45396 );
or ( w_45393 , \10329_b0 , \10330_b0 );
not ( \10330_b0 , w_45397 );
and ( w_45397 , w_45396 , \10330_b1 );
or ( \10337_b1 , \10334_b1 , w_45400 );
or ( \10337_b0 , \10334_b0 , w_45399 );
not ( w_45399 , w_45401 );
and ( w_45401 , w_45400 , w_45398 );
or ( w_45398 , \10335_b1 , w_45402 );
or ( w_45399 , \10335_b0 , \10336_b0 );
not ( \10336_b0 , w_45403 );
and ( w_45403 , w_45402 , \10336_b1 );
or ( \10341_b1 , \10338_b1 , w_45406 );
or ( \10341_b0 , \10338_b0 , w_45405 );
not ( w_45405 , w_45407 );
and ( w_45407 , w_45406 , w_45404 );
or ( w_45404 , \10339_b1 , w_45408 );
or ( w_45405 , \10339_b0 , \10340_b0 );
not ( \10340_b0 , w_45409 );
and ( w_45409 , w_45408 , \10340_b1 );
or ( \10346_b1 , \10343_b1 , w_45412 );
or ( \10346_b0 , \10343_b0 , w_45411 );
not ( w_45411 , w_45413 );
and ( w_45413 , w_45412 , w_45410 );
or ( w_45410 , \10344_b1 , w_45414 );
or ( w_45411 , \10344_b0 , \10345_b0 );
not ( \10345_b0 , w_45415 );
and ( w_45415 , w_45414 , \10345_b1 );
or ( \10350_b1 , \10347_b1 , w_45418 );
or ( \10350_b0 , \10347_b0 , w_45417 );
not ( w_45417 , w_45419 );
and ( w_45419 , w_45418 , w_45416 );
or ( w_45416 , \10348_b1 , w_45420 );
or ( w_45417 , \10348_b0 , \10349_b0 );
not ( \10349_b0 , w_45421 );
and ( w_45421 , w_45420 , \10349_b1 );
or ( \10355_b1 , \10352_b1 , w_45424 );
or ( \10355_b0 , \10352_b0 , w_45423 );
not ( w_45423 , w_45425 );
and ( w_45425 , w_45424 , w_45422 );
or ( w_45422 , \10353_b1 , w_45426 );
or ( w_45423 , \10353_b0 , \10354_b0 );
not ( \10354_b0 , w_45427 );
and ( w_45427 , w_45426 , \10354_b1 );
or ( \10360_b1 , \10357_b1 , w_45430 );
or ( \10360_b0 , \10357_b0 , w_45429 );
not ( w_45429 , w_45431 );
and ( w_45431 , w_45430 , w_45428 );
or ( w_45428 , \10358_b1 , w_45432 );
or ( w_45429 , \10358_b0 , \10359_b0 );
not ( \10359_b0 , w_45433 );
and ( w_45433 , w_45432 , \10359_b1 );
or ( \10364_b1 , \10361_b1 , w_45436 );
or ( \10364_b0 , \10361_b0 , w_45435 );
not ( w_45435 , w_45437 );
and ( w_45437 , w_45436 , w_45434 );
or ( w_45434 , \10362_b1 , w_45438 );
or ( w_45435 , \10362_b0 , \10363_b0 );
not ( \10363_b0 , w_45439 );
and ( w_45439 , w_45438 , \10363_b1 );
or ( \10369_b1 , \10366_b1 , w_45442 );
or ( \10369_b0 , \10366_b0 , w_45441 );
not ( w_45441 , w_45443 );
and ( w_45443 , w_45442 , w_45440 );
or ( w_45440 , \10367_b1 , w_45444 );
or ( w_45441 , \10367_b0 , \10368_b0 );
not ( \10368_b0 , w_45445 );
and ( w_45445 , w_45444 , \10368_b1 );
or ( \10375_b1 , \10372_b1 , w_45448 );
or ( \10375_b0 , \10372_b0 , w_45447 );
not ( w_45447 , w_45449 );
and ( w_45449 , w_45448 , w_45446 );
or ( w_45446 , \10373_b1 , w_45450 );
or ( w_45447 , \10373_b0 , \10374_b0 );
not ( \10374_b0 , w_45451 );
and ( w_45451 , w_45450 , \10374_b1 );
or ( \10462_b1 , \10459_b1 , w_45454 );
or ( \10462_b0 , \10459_b0 , w_45453 );
not ( w_45453 , w_45455 );
and ( w_45455 , w_45454 , w_45452 );
or ( w_45452 , \10460_b1 , w_45456 );
or ( w_45453 , \10460_b0 , \10461_b0 );
not ( \10461_b0 , w_45457 );
and ( w_45457 , w_45456 , \10461_b1 );
or ( \10466_b1 , \10463_b1 , w_45460 );
or ( \10466_b0 , \10463_b0 , w_45459 );
not ( w_45459 , w_45461 );
and ( w_45461 , w_45460 , w_45458 );
or ( w_45458 , \10464_b1 , w_45462 );
or ( w_45459 , \10464_b0 , \10465_b0 );
not ( \10465_b0 , w_45463 );
and ( w_45463 , w_45462 , \10465_b1 );
or ( \10476_b1 , \10473_b1 , w_45466 );
or ( \10476_b0 , \10473_b0 , w_45465 );
not ( w_45465 , w_45467 );
and ( w_45467 , w_45466 , w_45464 );
or ( w_45464 , \10474_b1 , w_45468 );
or ( w_45465 , \10474_b0 , \10475_b0 );
not ( \10475_b0 , w_45469 );
and ( w_45469 , w_45468 , \10475_b1 );
or ( \10481_b1 , \10478_b1 , w_45472 );
or ( \10481_b0 , \10478_b0 , w_45471 );
not ( w_45471 , w_45473 );
and ( w_45473 , w_45472 , w_45470 );
or ( w_45470 , \10479_b1 , w_45474 );
or ( w_45471 , \10479_b0 , \10480_b0 );
not ( \10480_b0 , w_45475 );
and ( w_45475 , w_45474 , \10480_b1 );
or ( \10485_b1 , \10482_b1 , w_45478 );
or ( \10485_b0 , \10482_b0 , w_45477 );
not ( w_45477 , w_45479 );
and ( w_45479 , w_45478 , w_45476 );
or ( w_45476 , \10483_b1 , w_45480 );
or ( w_45477 , \10483_b0 , \10484_b0 );
not ( \10484_b0 , w_45481 );
and ( w_45481 , w_45480 , \10484_b1 );
or ( \10489_b1 , \10486_b1 , w_45484 );
or ( \10489_b0 , \10486_b0 , w_45483 );
not ( w_45483 , w_45485 );
and ( w_45485 , w_45484 , w_45482 );
or ( w_45482 , \10487_b1 , w_45486 );
or ( w_45483 , \10487_b0 , \10488_b0 );
not ( \10488_b0 , w_45487 );
and ( w_45487 , w_45486 , \10488_b1 );
or ( \10497_b1 , \10494_b1 , w_45490 );
or ( \10497_b0 , \10494_b0 , w_45489 );
not ( w_45489 , w_45491 );
and ( w_45491 , w_45490 , w_45488 );
or ( w_45488 , \10495_b1 , w_45492 );
or ( w_45489 , \10495_b0 , \10496_b0 );
not ( \10496_b0 , w_45493 );
and ( w_45493 , w_45492 , \10496_b1 );
or ( \10501_b1 , \10498_b1 , w_45496 );
or ( \10501_b0 , \10498_b0 , w_45495 );
not ( w_45495 , w_45497 );
and ( w_45497 , w_45496 , w_45494 );
or ( w_45494 , \10499_b1 , w_45498 );
or ( w_45495 , \10499_b0 , \10500_b0 );
not ( \10500_b0 , w_45499 );
and ( w_45499 , w_45498 , \10500_b1 );
or ( \10533_b1 , \10530_b1 , w_45502 );
or ( \10533_b0 , \10530_b0 , w_45501 );
not ( w_45501 , w_45503 );
and ( w_45503 , w_45502 , w_45500 );
or ( w_45500 , \10531_b1 , w_45504 );
or ( w_45501 , \10531_b0 , \10532_b0 );
not ( \10532_b0 , w_45505 );
and ( w_45505 , w_45504 , \10532_b1 );
or ( \10537_b1 , \10534_b1 , w_45508 );
or ( \10537_b0 , \10534_b0 , w_45507 );
not ( w_45507 , w_45509 );
and ( w_45509 , w_45508 , w_45506 );
or ( w_45506 , \10535_b1 , w_45510 );
or ( w_45507 , \10535_b0 , \10536_b0 );
not ( \10536_b0 , w_45511 );
and ( w_45511 , w_45510 , \10536_b1 );
or ( \10545_b1 , \10542_b1 , w_45514 );
or ( \10545_b0 , \10542_b0 , w_45513 );
not ( w_45513 , w_45515 );
and ( w_45515 , w_45514 , w_45512 );
or ( w_45512 , \10543_b1 , w_45516 );
or ( w_45513 , \10543_b0 , \10544_b0 );
not ( \10544_b0 , w_45517 );
and ( w_45517 , w_45516 , \10544_b1 );
or ( \10549_b1 , \10546_b1 , w_45520 );
or ( \10549_b0 , \10546_b0 , w_45519 );
not ( w_45519 , w_45521 );
and ( w_45521 , w_45520 , w_45518 );
or ( w_45518 , \10547_b1 , w_45522 );
or ( w_45519 , \10547_b0 , \10548_b0 );
not ( \10548_b0 , w_45523 );
and ( w_45523 , w_45522 , \10548_b1 );
or ( \10554_b1 , \10551_b1 , w_45526 );
or ( \10554_b0 , \10551_b0 , w_45525 );
not ( w_45525 , w_45527 );
and ( w_45527 , w_45526 , w_45524 );
or ( w_45524 , \10552_b1 , w_45528 );
or ( w_45525 , \10552_b0 , \10553_b0 );
not ( \10553_b0 , w_45529 );
and ( w_45529 , w_45528 , \10553_b1 );
or ( \10560_b1 , \10557_b1 , w_45532 );
or ( \10560_b0 , \10557_b0 , w_45531 );
not ( w_45531 , w_45533 );
and ( w_45533 , w_45532 , w_45530 );
or ( w_45530 , \10558_b1 , w_45534 );
or ( w_45531 , \10558_b0 , \10559_b0 );
not ( \10559_b0 , w_45535 );
and ( w_45535 , w_45534 , \10559_b1 );
or ( \10620_b1 , \10617_b1 , w_45538 );
or ( \10620_b0 , \10617_b0 , w_45537 );
not ( w_45537 , w_45539 );
and ( w_45539 , w_45538 , w_45536 );
or ( w_45536 , \10618_b1 , w_45540 );
or ( w_45537 , \10618_b0 , \10619_b0 );
not ( \10619_b0 , w_45541 );
and ( w_45541 , w_45540 , \10619_b1 );
or ( \10624_b1 , \10621_b1 , w_45544 );
or ( \10624_b0 , \10621_b0 , w_45543 );
not ( w_45543 , w_45545 );
and ( w_45545 , w_45544 , w_45542 );
or ( w_45542 , \10622_b1 , w_45546 );
or ( w_45543 , \10622_b0 , \10623_b0 );
not ( \10623_b0 , w_45547 );
and ( w_45547 , w_45546 , \10623_b1 );
or ( \10629_b1 , \10626_b1 , w_45550 );
or ( \10629_b0 , \10626_b0 , w_45549 );
not ( w_45549 , w_45551 );
and ( w_45551 , w_45550 , w_45548 );
or ( w_45548 , \10627_b1 , w_45552 );
or ( w_45549 , \10627_b0 , \10628_b0 );
not ( \10628_b0 , w_45553 );
and ( w_45553 , w_45552 , \10628_b1 );
or ( \10637_b1 , \10634_b1 , w_45556 );
or ( \10637_b0 , \10634_b0 , w_45555 );
not ( w_45555 , w_45557 );
and ( w_45557 , w_45556 , w_45554 );
or ( w_45554 , \10635_b1 , w_45558 );
or ( w_45555 , \10635_b0 , \10636_b0 );
not ( \10636_b0 , w_45559 );
and ( w_45559 , w_45558 , \10636_b1 );
or ( \10643_b1 , \10640_b1 , w_45562 );
or ( \10643_b0 , \10640_b0 , w_45561 );
not ( w_45561 , w_45563 );
and ( w_45563 , w_45562 , w_45560 );
or ( w_45560 , \10641_b1 , w_45564 );
or ( w_45561 , \10641_b0 , \10642_b0 );
not ( \10642_b0 , w_45565 );
and ( w_45565 , w_45564 , \10642_b1 );
or ( \10647_b1 , \10644_b1 , w_45568 );
or ( \10647_b0 , \10644_b0 , w_45567 );
not ( w_45567 , w_45569 );
and ( w_45569 , w_45568 , w_45566 );
or ( w_45566 , \10645_b1 , w_45570 );
or ( w_45567 , \10645_b0 , \10646_b0 );
not ( \10646_b0 , w_45571 );
and ( w_45571 , w_45570 , \10646_b1 );
or ( \10651_b1 , \10648_b1 , w_45574 );
or ( \10651_b0 , \10648_b0 , w_45573 );
not ( w_45573 , w_45575 );
and ( w_45575 , w_45574 , w_45572 );
or ( w_45572 , \10649_b1 , w_45576 );
or ( w_45573 , \10649_b0 , \10650_b0 );
not ( \10650_b0 , w_45577 );
and ( w_45577 , w_45576 , \10650_b1 );
or ( \10656_b1 , \10653_b1 , w_45580 );
or ( \10656_b0 , \10653_b0 , w_45579 );
not ( w_45579 , w_45581 );
and ( w_45581 , w_45580 , w_45578 );
or ( w_45578 , \10654_b1 , w_45582 );
or ( w_45579 , \10654_b0 , \10655_b0 );
not ( \10655_b0 , w_45583 );
and ( w_45583 , w_45582 , \10655_b1 );
or ( \10662_b1 , \10659_b1 , w_45586 );
or ( \10662_b0 , \10659_b0 , w_45585 );
not ( w_45585 , w_45587 );
and ( w_45587 , w_45586 , w_45584 );
or ( w_45584 , \10660_b1 , w_45588 );
or ( w_45585 , \10660_b0 , \10661_b0 );
not ( \10661_b0 , w_45589 );
and ( w_45589 , w_45588 , \10661_b1 );
or ( \10666_b1 , \10663_b1 , w_45592 );
or ( \10666_b0 , \10663_b0 , w_45591 );
not ( w_45591 , w_45593 );
and ( w_45593 , w_45592 , w_45590 );
or ( w_45590 , \10664_b1 , w_45594 );
or ( w_45591 , \10664_b0 , \10665_b0 );
not ( \10665_b0 , w_45595 );
and ( w_45595 , w_45594 , \10665_b1 );
or ( \10671_b1 , \10668_b1 , w_45598 );
or ( \10671_b0 , \10668_b0 , w_45597 );
not ( w_45597 , w_45599 );
and ( w_45599 , w_45598 , w_45596 );
or ( w_45596 , \10669_b1 , w_45600 );
or ( w_45597 , \10669_b0 , \10670_b0 );
not ( \10670_b0 , w_45601 );
and ( w_45601 , w_45600 , \10670_b1 );
or ( \10675_b1 , \10672_b1 , w_45604 );
or ( \10675_b0 , \10672_b0 , w_45603 );
not ( w_45603 , w_45605 );
and ( w_45605 , w_45604 , w_45602 );
or ( w_45602 , \10673_b1 , w_45606 );
or ( w_45603 , \10673_b0 , \10674_b0 );
not ( \10674_b0 , w_45607 );
and ( w_45607 , w_45606 , \10674_b1 );
or ( \10680_b1 , \10677_b1 , w_45610 );
or ( \10680_b0 , \10677_b0 , w_45609 );
not ( w_45609 , w_45611 );
and ( w_45611 , w_45610 , w_45608 );
or ( w_45608 , \10678_b1 , w_45612 );
or ( w_45609 , \10678_b0 , \10679_b0 );
not ( \10679_b0 , w_45613 );
and ( w_45613 , w_45612 , \10679_b1 );
or ( \10685_b1 , \10682_b1 , w_45616 );
or ( \10685_b0 , \10682_b0 , w_45615 );
not ( w_45615 , w_45617 );
and ( w_45617 , w_45616 , w_45614 );
or ( w_45614 , \10683_b1 , w_45618 );
or ( w_45615 , \10683_b0 , \10684_b0 );
not ( \10684_b0 , w_45619 );
and ( w_45619 , w_45618 , \10684_b1 );
or ( \10689_b1 , \10686_b1 , w_45622 );
or ( \10689_b0 , \10686_b0 , w_45621 );
not ( w_45621 , w_45623 );
and ( w_45623 , w_45622 , w_45620 );
or ( w_45620 , \10687_b1 , w_45624 );
or ( w_45621 , \10687_b0 , \10688_b0 );
not ( \10688_b0 , w_45625 );
and ( w_45625 , w_45624 , \10688_b1 );
or ( \10694_b1 , \10691_b1 , w_45628 );
or ( \10694_b0 , \10691_b0 , w_45627 );
not ( w_45627 , w_45629 );
and ( w_45629 , w_45628 , w_45626 );
or ( w_45626 , \10692_b1 , w_45630 );
or ( w_45627 , \10692_b0 , \10693_b0 );
not ( \10693_b0 , w_45631 );
and ( w_45631 , w_45630 , \10693_b1 );
or ( \10700_b1 , \10697_b1 , w_45634 );
or ( \10700_b0 , \10697_b0 , w_45633 );
not ( w_45633 , w_45635 );
and ( w_45635 , w_45634 , w_45632 );
or ( w_45632 , \10698_b1 , w_45636 );
or ( w_45633 , \10698_b0 , \10699_b0 );
not ( \10699_b0 , w_45637 );
and ( w_45637 , w_45636 , \10699_b1 );
or ( \10787_b1 , \10784_b1 , w_45640 );
or ( \10787_b0 , \10784_b0 , w_45639 );
not ( w_45639 , w_45641 );
and ( w_45641 , w_45640 , w_45638 );
or ( w_45638 , \10785_b1 , w_45642 );
or ( w_45639 , \10785_b0 , \10786_b0 );
not ( \10786_b0 , w_45643 );
and ( w_45643 , w_45642 , \10786_b1 );
or ( \10791_b1 , \10788_b1 , w_45646 );
or ( \10791_b0 , \10788_b0 , w_45645 );
not ( w_45645 , w_45647 );
and ( w_45647 , w_45646 , w_45644 );
or ( w_45644 , \10789_b1 , w_45648 );
or ( w_45645 , \10789_b0 , \10790_b0 );
not ( \10790_b0 , w_45649 );
and ( w_45649 , w_45648 , \10790_b1 );
or ( \10801_b1 , \10798_b1 , w_45652 );
or ( \10801_b0 , \10798_b0 , w_45651 );
not ( w_45651 , w_45653 );
and ( w_45653 , w_45652 , w_45650 );
or ( w_45650 , \10799_b1 , w_45654 );
or ( w_45651 , \10799_b0 , \10800_b0 );
not ( \10800_b0 , w_45655 );
and ( w_45655 , w_45654 , \10800_b1 );
or ( \10806_b1 , \10803_b1 , w_45658 );
or ( \10806_b0 , \10803_b0 , w_45657 );
not ( w_45657 , w_45659 );
and ( w_45659 , w_45658 , w_45656 );
or ( w_45656 , \10804_b1 , w_45660 );
or ( w_45657 , \10804_b0 , \10805_b0 );
not ( \10805_b0 , w_45661 );
and ( w_45661 , w_45660 , \10805_b1 );
or ( \10810_b1 , \10807_b1 , w_45664 );
or ( \10810_b0 , \10807_b0 , w_45663 );
not ( w_45663 , w_45665 );
and ( w_45665 , w_45664 , w_45662 );
or ( w_45662 , \10808_b1 , w_45666 );
or ( w_45663 , \10808_b0 , \10809_b0 );
not ( \10809_b0 , w_45667 );
and ( w_45667 , w_45666 , \10809_b1 );
or ( \10814_b1 , \10811_b1 , w_45670 );
or ( \10814_b0 , \10811_b0 , w_45669 );
not ( w_45669 , w_45671 );
and ( w_45671 , w_45670 , w_45668 );
or ( w_45668 , \10812_b1 , w_45672 );
or ( w_45669 , \10812_b0 , \10813_b0 );
not ( \10813_b0 , w_45673 );
and ( w_45673 , w_45672 , \10813_b1 );
or ( \10822_b1 , \10819_b1 , w_45676 );
or ( \10822_b0 , \10819_b0 , w_45675 );
not ( w_45675 , w_45677 );
and ( w_45677 , w_45676 , w_45674 );
or ( w_45674 , \10820_b1 , w_45678 );
or ( w_45675 , \10820_b0 , \10821_b0 );
not ( \10821_b0 , w_45679 );
and ( w_45679 , w_45678 , \10821_b1 );
or ( \10826_b1 , \10823_b1 , w_45682 );
or ( \10826_b0 , \10823_b0 , w_45681 );
not ( w_45681 , w_45683 );
and ( w_45683 , w_45682 , w_45680 );
or ( w_45680 , \10824_b1 , w_45684 );
or ( w_45681 , \10824_b0 , \10825_b0 );
not ( \10825_b0 , w_45685 );
and ( w_45685 , w_45684 , \10825_b1 );
or ( \10858_b1 , \10855_b1 , w_45688 );
or ( \10858_b0 , \10855_b0 , w_45687 );
not ( w_45687 , w_45689 );
and ( w_45689 , w_45688 , w_45686 );
or ( w_45686 , \10856_b1 , w_45690 );
or ( w_45687 , \10856_b0 , \10857_b0 );
not ( \10857_b0 , w_45691 );
and ( w_45691 , w_45690 , \10857_b1 );
or ( \10862_b1 , \10859_b1 , w_45694 );
or ( \10862_b0 , \10859_b0 , w_45693 );
not ( w_45693 , w_45695 );
and ( w_45695 , w_45694 , w_45692 );
or ( w_45692 , \10860_b1 , w_45696 );
or ( w_45693 , \10860_b0 , \10861_b0 );
not ( \10861_b0 , w_45697 );
and ( w_45697 , w_45696 , \10861_b1 );
or ( \10870_b1 , \10867_b1 , w_45700 );
or ( \10870_b0 , \10867_b0 , w_45699 );
not ( w_45699 , w_45701 );
and ( w_45701 , w_45700 , w_45698 );
or ( w_45698 , \10868_b1 , w_45702 );
or ( w_45699 , \10868_b0 , \10869_b0 );
not ( \10869_b0 , w_45703 );
and ( w_45703 , w_45702 , \10869_b1 );
or ( \10874_b1 , \10871_b1 , w_45706 );
or ( \10874_b0 , \10871_b0 , w_45705 );
not ( w_45705 , w_45707 );
and ( w_45707 , w_45706 , w_45704 );
or ( w_45704 , \10872_b1 , w_45708 );
or ( w_45705 , \10872_b0 , \10873_b0 );
not ( \10873_b0 , w_45709 );
and ( w_45709 , w_45708 , \10873_b1 );
or ( \10879_b1 , \10876_b1 , w_45712 );
or ( \10879_b0 , \10876_b0 , w_45711 );
not ( w_45711 , w_45713 );
and ( w_45713 , w_45712 , w_45710 );
or ( w_45710 , \10877_b1 , w_45714 );
or ( w_45711 , \10877_b0 , \10878_b0 );
not ( \10878_b0 , w_45715 );
and ( w_45715 , w_45714 , \10878_b1 );
or ( \10885_b1 , \10882_b1 , w_45718 );
or ( \10885_b0 , \10882_b0 , w_45717 );
not ( w_45717 , w_45719 );
and ( w_45719 , w_45718 , w_45716 );
or ( w_45716 , \10883_b1 , w_45720 );
or ( w_45717 , \10883_b0 , \10884_b0 );
not ( \10884_b0 , w_45721 );
and ( w_45721 , w_45720 , \10884_b1 );
or ( \10945_b1 , \10942_b1 , w_45724 );
or ( \10945_b0 , \10942_b0 , w_45723 );
not ( w_45723 , w_45725 );
and ( w_45725 , w_45724 , w_45722 );
or ( w_45722 , \10943_b1 , w_45726 );
or ( w_45723 , \10943_b0 , \10944_b0 );
not ( \10944_b0 , w_45727 );
and ( w_45727 , w_45726 , \10944_b1 );
or ( \10949_b1 , \10946_b1 , w_45730 );
or ( \10949_b0 , \10946_b0 , w_45729 );
not ( w_45729 , w_45731 );
and ( w_45731 , w_45730 , w_45728 );
or ( w_45728 , \10947_b1 , w_45732 );
or ( w_45729 , \10947_b0 , \10948_b0 );
not ( \10948_b0 , w_45733 );
and ( w_45733 , w_45732 , \10948_b1 );
or ( \10954_b1 , \10951_b1 , w_45736 );
or ( \10954_b0 , \10951_b0 , w_45735 );
not ( w_45735 , w_45737 );
and ( w_45737 , w_45736 , w_45734 );
or ( w_45734 , \10952_b1 , w_45738 );
or ( w_45735 , \10952_b0 , \10953_b0 );
not ( \10953_b0 , w_45739 );
and ( w_45739 , w_45738 , \10953_b1 );
or ( \10962_b1 , \10959_b1 , w_45742 );
or ( \10962_b0 , \10959_b0 , w_45741 );
not ( w_45741 , w_45743 );
and ( w_45743 , w_45742 , w_45740 );
or ( w_45740 , \10960_b1 , w_45744 );
or ( w_45741 , \10960_b0 , \10961_b0 );
not ( \10961_b0 , w_45745 );
and ( w_45745 , w_45744 , \10961_b1 );
or ( \10969_b1 , \10966_b1 , w_45748 );
or ( \10969_b0 , \10966_b0 , w_45747 );
not ( w_45747 , w_45749 );
and ( w_45749 , w_45748 , w_45746 );
or ( w_45746 , \10967_b1 , w_45750 );
or ( w_45747 , \10967_b0 , \10968_b0 );
not ( \10968_b0 , w_45751 );
and ( w_45751 , w_45750 , \10968_b1 );
or ( \10973_b1 , \10970_b1 , w_45754 );
or ( \10973_b0 , \10970_b0 , w_45753 );
not ( w_45753 , w_45755 );
and ( w_45755 , w_45754 , w_45752 );
or ( w_45752 , \10971_b1 , w_45756 );
or ( w_45753 , \10971_b0 , \10972_b0 );
not ( \10972_b0 , w_45757 );
and ( w_45757 , w_45756 , \10972_b1 );
or ( \10977_b1 , \10974_b1 , w_45760 );
or ( \10977_b0 , \10974_b0 , w_45759 );
not ( w_45759 , w_45761 );
and ( w_45761 , w_45760 , w_45758 );
or ( w_45758 , \10975_b1 , w_45762 );
or ( w_45759 , \10975_b0 , \10976_b0 );
not ( \10976_b0 , w_45763 );
and ( w_45763 , w_45762 , \10976_b1 );
or ( \10982_b1 , \10979_b1 , w_45766 );
or ( \10982_b0 , \10979_b0 , w_45765 );
not ( w_45765 , w_45767 );
and ( w_45767 , w_45766 , w_45764 );
or ( w_45764 , \10980_b1 , w_45768 );
or ( w_45765 , \10980_b0 , \10981_b0 );
not ( \10981_b0 , w_45769 );
and ( w_45769 , w_45768 , \10981_b1 );
or ( \10988_b1 , \10985_b1 , w_45772 );
or ( \10988_b0 , \10985_b0 , w_45771 );
not ( w_45771 , w_45773 );
and ( w_45773 , w_45772 , w_45770 );
or ( w_45770 , \10986_b1 , w_45774 );
or ( w_45771 , \10986_b0 , \10987_b0 );
not ( \10987_b0 , w_45775 );
and ( w_45775 , w_45774 , \10987_b1 );
or ( \10992_b1 , \10989_b1 , w_45778 );
or ( \10992_b0 , \10989_b0 , w_45777 );
not ( w_45777 , w_45779 );
and ( w_45779 , w_45778 , w_45776 );
or ( w_45776 , \10990_b1 , w_45780 );
or ( w_45777 , \10990_b0 , \10991_b0 );
not ( \10991_b0 , w_45781 );
and ( w_45781 , w_45780 , \10991_b1 );
or ( \10997_b1 , \10994_b1 , w_45784 );
or ( \10997_b0 , \10994_b0 , w_45783 );
not ( w_45783 , w_45785 );
and ( w_45785 , w_45784 , w_45782 );
or ( w_45782 , \10995_b1 , w_45786 );
or ( w_45783 , \10995_b0 , \10996_b0 );
not ( \10996_b0 , w_45787 );
and ( w_45787 , w_45786 , \10996_b1 );
or ( \11001_b1 , \10998_b1 , w_45790 );
or ( \11001_b0 , \10998_b0 , w_45789 );
not ( w_45789 , w_45791 );
and ( w_45791 , w_45790 , w_45788 );
or ( w_45788 , \10999_b1 , w_45792 );
or ( w_45789 , \10999_b0 , \11000_b0 );
not ( \11000_b0 , w_45793 );
and ( w_45793 , w_45792 , \11000_b1 );
or ( \11006_b1 , \11003_b1 , w_45796 );
or ( \11006_b0 , \11003_b0 , w_45795 );
not ( w_45795 , w_45797 );
and ( w_45797 , w_45796 , w_45794 );
or ( w_45794 , \11004_b1 , w_45798 );
or ( w_45795 , \11004_b0 , \11005_b0 );
not ( \11005_b0 , w_45799 );
and ( w_45799 , w_45798 , \11005_b1 );
or ( \11011_b1 , \11008_b1 , w_45802 );
or ( \11011_b0 , \11008_b0 , w_45801 );
not ( w_45801 , w_45803 );
and ( w_45803 , w_45802 , w_45800 );
or ( w_45800 , \11009_b1 , w_45804 );
or ( w_45801 , \11009_b0 , \11010_b0 );
not ( \11010_b0 , w_45805 );
and ( w_45805 , w_45804 , \11010_b1 );
or ( \11015_b1 , \11012_b1 , w_45808 );
or ( \11015_b0 , \11012_b0 , w_45807 );
not ( w_45807 , w_45809 );
and ( w_45809 , w_45808 , w_45806 );
or ( w_45806 , \11013_b1 , w_45810 );
or ( w_45807 , \11013_b0 , \11014_b0 );
not ( \11014_b0 , w_45811 );
and ( w_45811 , w_45810 , \11014_b1 );
or ( \11020_b1 , \11017_b1 , w_45814 );
or ( \11020_b0 , \11017_b0 , w_45813 );
not ( w_45813 , w_45815 );
and ( w_45815 , w_45814 , w_45812 );
or ( w_45812 , \11018_b1 , w_45816 );
or ( w_45813 , \11018_b0 , \11019_b0 );
not ( \11019_b0 , w_45817 );
and ( w_45817 , w_45816 , \11019_b1 );
or ( \11026_b1 , \11023_b1 , w_45820 );
or ( \11026_b0 , \11023_b0 , w_45819 );
not ( w_45819 , w_45821 );
and ( w_45821 , w_45820 , w_45818 );
or ( w_45818 , \11024_b1 , w_45822 );
or ( w_45819 , \11024_b0 , \11025_b0 );
not ( \11025_b0 , w_45823 );
and ( w_45823 , w_45822 , \11025_b1 );
or ( \11113_b1 , \11110_b1 , w_45826 );
or ( \11113_b0 , \11110_b0 , w_45825 );
not ( w_45825 , w_45827 );
and ( w_45827 , w_45826 , w_45824 );
or ( w_45824 , \11111_b1 , w_45828 );
or ( w_45825 , \11111_b0 , \11112_b0 );
not ( \11112_b0 , w_45829 );
and ( w_45829 , w_45828 , \11112_b1 );
or ( \11117_b1 , \11114_b1 , w_45832 );
or ( \11117_b0 , \11114_b0 , w_45831 );
not ( w_45831 , w_45833 );
and ( w_45833 , w_45832 , w_45830 );
or ( w_45830 , \11115_b1 , w_45834 );
or ( w_45831 , \11115_b0 , \11116_b0 );
not ( \11116_b0 , w_45835 );
and ( w_45835 , w_45834 , \11116_b1 );
or ( \11127_b1 , \11124_b1 , w_45838 );
or ( \11127_b0 , \11124_b0 , w_45837 );
not ( w_45837 , w_45839 );
and ( w_45839 , w_45838 , w_45836 );
or ( w_45836 , \11125_b1 , w_45840 );
or ( w_45837 , \11125_b0 , \11126_b0 );
not ( \11126_b0 , w_45841 );
and ( w_45841 , w_45840 , \11126_b1 );
or ( \11132_b1 , \11129_b1 , w_45844 );
or ( \11132_b0 , \11129_b0 , w_45843 );
not ( w_45843 , w_45845 );
and ( w_45845 , w_45844 , w_45842 );
or ( w_45842 , \11130_b1 , w_45846 );
or ( w_45843 , \11130_b0 , \11131_b0 );
not ( \11131_b0 , w_45847 );
and ( w_45847 , w_45846 , \11131_b1 );
or ( \11136_b1 , \11133_b1 , w_45850 );
or ( \11136_b0 , \11133_b0 , w_45849 );
not ( w_45849 , w_45851 );
and ( w_45851 , w_45850 , w_45848 );
or ( w_45848 , \11134_b1 , w_45852 );
or ( w_45849 , \11134_b0 , \11135_b0 );
not ( \11135_b0 , w_45853 );
and ( w_45853 , w_45852 , \11135_b1 );
or ( \11140_b1 , \11137_b1 , w_45856 );
or ( \11140_b0 , \11137_b0 , w_45855 );
not ( w_45855 , w_45857 );
and ( w_45857 , w_45856 , w_45854 );
or ( w_45854 , \11138_b1 , w_45858 );
or ( w_45855 , \11138_b0 , \11139_b0 );
not ( \11139_b0 , w_45859 );
and ( w_45859 , w_45858 , \11139_b1 );
or ( \11148_b1 , \11145_b1 , w_45862 );
or ( \11148_b0 , \11145_b0 , w_45861 );
not ( w_45861 , w_45863 );
and ( w_45863 , w_45862 , w_45860 );
or ( w_45860 , \11146_b1 , w_45864 );
or ( w_45861 , \11146_b0 , \11147_b0 );
not ( \11147_b0 , w_45865 );
and ( w_45865 , w_45864 , \11147_b1 );
or ( \11152_b1 , \11149_b1 , w_45868 );
or ( \11152_b0 , \11149_b0 , w_45867 );
not ( w_45867 , w_45869 );
and ( w_45869 , w_45868 , w_45866 );
or ( w_45866 , \11150_b1 , w_45870 );
or ( w_45867 , \11150_b0 , \11151_b0 );
not ( \11151_b0 , w_45871 );
and ( w_45871 , w_45870 , \11151_b1 );
or ( \11184_b1 , \11181_b1 , w_45874 );
or ( \11184_b0 , \11181_b0 , w_45873 );
not ( w_45873 , w_45875 );
and ( w_45875 , w_45874 , w_45872 );
or ( w_45872 , \11182_b1 , w_45876 );
or ( w_45873 , \11182_b0 , \11183_b0 );
not ( \11183_b0 , w_45877 );
and ( w_45877 , w_45876 , \11183_b1 );
or ( \11188_b1 , \11185_b1 , w_45880 );
or ( \11188_b0 , \11185_b0 , w_45879 );
not ( w_45879 , w_45881 );
and ( w_45881 , w_45880 , w_45878 );
or ( w_45878 , \11186_b1 , w_45882 );
or ( w_45879 , \11186_b0 , \11187_b0 );
not ( \11187_b0 , w_45883 );
and ( w_45883 , w_45882 , \11187_b1 );
or ( \11196_b1 , \11193_b1 , w_45886 );
or ( \11196_b0 , \11193_b0 , w_45885 );
not ( w_45885 , w_45887 );
and ( w_45887 , w_45886 , w_45884 );
or ( w_45884 , \11194_b1 , w_45888 );
or ( w_45885 , \11194_b0 , \11195_b0 );
not ( \11195_b0 , w_45889 );
and ( w_45889 , w_45888 , \11195_b1 );
or ( \11200_b1 , \11197_b1 , w_45892 );
or ( \11200_b0 , \11197_b0 , w_45891 );
not ( w_45891 , w_45893 );
and ( w_45893 , w_45892 , w_45890 );
or ( w_45890 , \11198_b1 , w_45894 );
or ( w_45891 , \11198_b0 , \11199_b0 );
not ( \11199_b0 , w_45895 );
and ( w_45895 , w_45894 , \11199_b1 );
or ( \11205_b1 , \11202_b1 , w_45898 );
or ( \11205_b0 , \11202_b0 , w_45897 );
not ( w_45897 , w_45899 );
and ( w_45899 , w_45898 , w_45896 );
or ( w_45896 , \11203_b1 , w_45900 );
or ( w_45897 , \11203_b0 , \11204_b0 );
not ( \11204_b0 , w_45901 );
and ( w_45901 , w_45900 , \11204_b1 );
or ( \11211_b1 , \11208_b1 , w_45904 );
or ( \11211_b0 , \11208_b0 , w_45903 );
not ( w_45903 , w_45905 );
and ( w_45905 , w_45904 , w_45902 );
or ( w_45902 , \11209_b1 , w_45906 );
or ( w_45903 , \11209_b0 , \11210_b0 );
not ( \11210_b0 , w_45907 );
and ( w_45907 , w_45906 , \11210_b1 );
or ( \11271_b1 , \11268_b1 , w_45910 );
or ( \11271_b0 , \11268_b0 , w_45909 );
not ( w_45909 , w_45911 );
and ( w_45911 , w_45910 , w_45908 );
or ( w_45908 , \11269_b1 , w_45912 );
or ( w_45909 , \11269_b0 , \11270_b0 );
not ( \11270_b0 , w_45913 );
and ( w_45913 , w_45912 , \11270_b1 );
or ( \11275_b1 , \11272_b1 , w_45916 );
or ( \11275_b0 , \11272_b0 , w_45915 );
not ( w_45915 , w_45917 );
and ( w_45917 , w_45916 , w_45914 );
or ( w_45914 , \11273_b1 , w_45918 );
or ( w_45915 , \11273_b0 , \11274_b0 );
not ( \11274_b0 , w_45919 );
and ( w_45919 , w_45918 , \11274_b1 );
or ( \11280_b1 , \11277_b1 , w_45922 );
or ( \11280_b0 , \11277_b0 , w_45921 );
not ( w_45921 , w_45923 );
and ( w_45923 , w_45922 , w_45920 );
or ( w_45920 , \11278_b1 , w_45924 );
or ( w_45921 , \11278_b0 , \11279_b0 );
not ( \11279_b0 , w_45925 );
and ( w_45925 , w_45924 , \11279_b1 );
or ( \11288_b1 , \11285_b1 , w_45928 );
or ( \11288_b0 , \11285_b0 , w_45927 );
not ( w_45927 , w_45929 );
and ( w_45929 , w_45928 , w_45926 );
or ( w_45926 , \11286_b1 , w_45930 );
or ( w_45927 , \11286_b0 , \11287_b0 );
not ( \11287_b0 , w_45931 );
and ( w_45931 , w_45930 , \11287_b1 );
or ( \11294_b1 , \11291_b1 , w_45934 );
or ( \11294_b0 , \11291_b0 , w_45933 );
not ( w_45933 , w_45935 );
and ( w_45935 , w_45934 , w_45932 );
or ( w_45932 , \11292_b1 , w_45936 );
or ( w_45933 , \11292_b0 , \11293_b0 );
not ( \11293_b0 , w_45937 );
and ( w_45937 , w_45936 , \11293_b1 );
or ( \11298_b1 , \11295_b1 , w_45940 );
or ( \11298_b0 , \11295_b0 , w_45939 );
not ( w_45939 , w_45941 );
and ( w_45941 , w_45940 , w_45938 );
or ( w_45938 , \11296_b1 , w_45942 );
or ( w_45939 , \11296_b0 , \11297_b0 );
not ( \11297_b0 , w_45943 );
and ( w_45943 , w_45942 , \11297_b1 );
or ( \11302_b1 , \11299_b1 , w_45946 );
or ( \11302_b0 , \11299_b0 , w_45945 );
not ( w_45945 , w_45947 );
and ( w_45947 , w_45946 , w_45944 );
or ( w_45944 , \11300_b1 , w_45948 );
or ( w_45945 , \11300_b0 , \11301_b0 );
not ( \11301_b0 , w_45949 );
and ( w_45949 , w_45948 , \11301_b1 );
or ( \11307_b1 , \11304_b1 , w_45952 );
or ( \11307_b0 , \11304_b0 , w_45951 );
not ( w_45951 , w_45953 );
and ( w_45953 , w_45952 , w_45950 );
or ( w_45950 , \11305_b1 , w_45954 );
or ( w_45951 , \11305_b0 , \11306_b0 );
not ( \11306_b0 , w_45955 );
and ( w_45955 , w_45954 , \11306_b1 );
or ( \11313_b1 , \11310_b1 , w_45958 );
or ( \11313_b0 , \11310_b0 , w_45957 );
not ( w_45957 , w_45959 );
and ( w_45959 , w_45958 , w_45956 );
or ( w_45956 , \11311_b1 , w_45960 );
or ( w_45957 , \11311_b0 , \11312_b0 );
not ( \11312_b0 , w_45961 );
and ( w_45961 , w_45960 , \11312_b1 );
or ( \11317_b1 , \11314_b1 , w_45964 );
or ( \11317_b0 , \11314_b0 , w_45963 );
not ( w_45963 , w_45965 );
and ( w_45965 , w_45964 , w_45962 );
or ( w_45962 , \11315_b1 , w_45966 );
or ( w_45963 , \11315_b0 , \11316_b0 );
not ( \11316_b0 , w_45967 );
and ( w_45967 , w_45966 , \11316_b1 );
or ( \11322_b1 , \11319_b1 , w_45970 );
or ( \11322_b0 , \11319_b0 , w_45969 );
not ( w_45969 , w_45971 );
and ( w_45971 , w_45970 , w_45968 );
or ( w_45968 , \11320_b1 , w_45972 );
or ( w_45969 , \11320_b0 , \11321_b0 );
not ( \11321_b0 , w_45973 );
and ( w_45973 , w_45972 , \11321_b1 );
or ( \11326_b1 , \11323_b1 , w_45976 );
or ( \11326_b0 , \11323_b0 , w_45975 );
not ( w_45975 , w_45977 );
and ( w_45977 , w_45976 , w_45974 );
or ( w_45974 , \11324_b1 , w_45978 );
or ( w_45975 , \11324_b0 , \11325_b0 );
not ( \11325_b0 , w_45979 );
and ( w_45979 , w_45978 , \11325_b1 );
or ( \11331_b1 , \11328_b1 , w_45982 );
or ( \11331_b0 , \11328_b0 , w_45981 );
not ( w_45981 , w_45983 );
and ( w_45983 , w_45982 , w_45980 );
or ( w_45980 , \11329_b1 , w_45984 );
or ( w_45981 , \11329_b0 , \11330_b0 );
not ( \11330_b0 , w_45985 );
and ( w_45985 , w_45984 , \11330_b1 );
or ( \11336_b1 , \11333_b1 , w_45988 );
or ( \11336_b0 , \11333_b0 , w_45987 );
not ( w_45987 , w_45989 );
and ( w_45989 , w_45988 , w_45986 );
or ( w_45986 , \11334_b1 , w_45990 );
or ( w_45987 , \11334_b0 , \11335_b0 );
not ( \11335_b0 , w_45991 );
and ( w_45991 , w_45990 , \11335_b1 );
or ( \11340_b1 , \11337_b1 , w_45994 );
or ( \11340_b0 , \11337_b0 , w_45993 );
not ( w_45993 , w_45995 );
and ( w_45995 , w_45994 , w_45992 );
or ( w_45992 , \11338_b1 , w_45996 );
or ( w_45993 , \11338_b0 , \11339_b0 );
not ( \11339_b0 , w_45997 );
and ( w_45997 , w_45996 , \11339_b1 );
or ( \11345_b1 , \11342_b1 , w_46000 );
or ( \11345_b0 , \11342_b0 , w_45999 );
not ( w_45999 , w_46001 );
and ( w_46001 , w_46000 , w_45998 );
or ( w_45998 , \11343_b1 , w_46002 );
or ( w_45999 , \11343_b0 , \11344_b0 );
not ( \11344_b0 , w_46003 );
and ( w_46003 , w_46002 , \11344_b1 );
or ( \11351_b1 , \11348_b1 , w_46006 );
or ( \11351_b0 , \11348_b0 , w_46005 );
not ( w_46005 , w_46007 );
and ( w_46007 , w_46006 , w_46004 );
or ( w_46004 , \11349_b1 , w_46008 );
or ( w_46005 , \11349_b0 , \11350_b0 );
not ( \11350_b0 , w_46009 );
and ( w_46009 , w_46008 , \11350_b1 );
or ( \11438_b1 , \11435_b1 , w_46012 );
or ( \11438_b0 , \11435_b0 , w_46011 );
not ( w_46011 , w_46013 );
and ( w_46013 , w_46012 , w_46010 );
or ( w_46010 , \11436_b1 , w_46014 );
or ( w_46011 , \11436_b0 , \11437_b0 );
not ( \11437_b0 , w_46015 );
and ( w_46015 , w_46014 , \11437_b1 );
or ( \11442_b1 , \11439_b1 , w_46018 );
or ( \11442_b0 , \11439_b0 , w_46017 );
not ( w_46017 , w_46019 );
and ( w_46019 , w_46018 , w_46016 );
or ( w_46016 , \11440_b1 , w_46020 );
or ( w_46017 , \11440_b0 , \11441_b0 );
not ( \11441_b0 , w_46021 );
and ( w_46021 , w_46020 , \11441_b1 );
or ( \11452_b1 , \11449_b1 , w_46024 );
or ( \11452_b0 , \11449_b0 , w_46023 );
not ( w_46023 , w_46025 );
and ( w_46025 , w_46024 , w_46022 );
or ( w_46022 , \11450_b1 , w_46026 );
or ( w_46023 , \11450_b0 , \11451_b0 );
not ( \11451_b0 , w_46027 );
and ( w_46027 , w_46026 , \11451_b1 );
or ( \11457_b1 , \11454_b1 , w_46030 );
or ( \11457_b0 , \11454_b0 , w_46029 );
not ( w_46029 , w_46031 );
and ( w_46031 , w_46030 , w_46028 );
or ( w_46028 , \11455_b1 , w_46032 );
or ( w_46029 , \11455_b0 , \11456_b0 );
not ( \11456_b0 , w_46033 );
and ( w_46033 , w_46032 , \11456_b1 );
or ( \11461_b1 , \11458_b1 , w_46036 );
or ( \11461_b0 , \11458_b0 , w_46035 );
not ( w_46035 , w_46037 );
and ( w_46037 , w_46036 , w_46034 );
or ( w_46034 , \11459_b1 , w_46038 );
or ( w_46035 , \11459_b0 , \11460_b0 );
not ( \11460_b0 , w_46039 );
and ( w_46039 , w_46038 , \11460_b1 );
or ( \11465_b1 , \11462_b1 , w_46042 );
or ( \11465_b0 , \11462_b0 , w_46041 );
not ( w_46041 , w_46043 );
and ( w_46043 , w_46042 , w_46040 );
or ( w_46040 , \11463_b1 , w_46044 );
or ( w_46041 , \11463_b0 , \11464_b0 );
not ( \11464_b0 , w_46045 );
and ( w_46045 , w_46044 , \11464_b1 );
or ( \11473_b1 , \11470_b1 , w_46048 );
or ( \11473_b0 , \11470_b0 , w_46047 );
not ( w_46047 , w_46049 );
and ( w_46049 , w_46048 , w_46046 );
or ( w_46046 , \11471_b1 , w_46050 );
or ( w_46047 , \11471_b0 , \11472_b0 );
not ( \11472_b0 , w_46051 );
and ( w_46051 , w_46050 , \11472_b1 );
or ( \11477_b1 , \11474_b1 , w_46054 );
or ( \11477_b0 , \11474_b0 , w_46053 );
not ( w_46053 , w_46055 );
and ( w_46055 , w_46054 , w_46052 );
or ( w_46052 , \11475_b1 , w_46056 );
or ( w_46053 , \11475_b0 , \11476_b0 );
not ( \11476_b0 , w_46057 );
and ( w_46057 , w_46056 , \11476_b1 );
or ( \11509_b1 , \11506_b1 , w_46060 );
or ( \11509_b0 , \11506_b0 , w_46059 );
not ( w_46059 , w_46061 );
and ( w_46061 , w_46060 , w_46058 );
or ( w_46058 , \11507_b1 , w_46062 );
or ( w_46059 , \11507_b0 , \11508_b0 );
not ( \11508_b0 , w_46063 );
and ( w_46063 , w_46062 , \11508_b1 );
or ( \11513_b1 , \11510_b1 , w_46066 );
or ( \11513_b0 , \11510_b0 , w_46065 );
not ( w_46065 , w_46067 );
and ( w_46067 , w_46066 , w_46064 );
or ( w_46064 , \11511_b1 , w_46068 );
or ( w_46065 , \11511_b0 , \11512_b0 );
not ( \11512_b0 , w_46069 );
and ( w_46069 , w_46068 , \11512_b1 );
or ( \11521_b1 , \11518_b1 , w_46072 );
or ( \11521_b0 , \11518_b0 , w_46071 );
not ( w_46071 , w_46073 );
and ( w_46073 , w_46072 , w_46070 );
or ( w_46070 , \11519_b1 , w_46074 );
or ( w_46071 , \11519_b0 , \11520_b0 );
not ( \11520_b0 , w_46075 );
and ( w_46075 , w_46074 , \11520_b1 );
or ( \11525_b1 , \11522_b1 , w_46078 );
or ( \11525_b0 , \11522_b0 , w_46077 );
not ( w_46077 , w_46079 );
and ( w_46079 , w_46078 , w_46076 );
or ( w_46076 , \11523_b1 , w_46080 );
or ( w_46077 , \11523_b0 , \11524_b0 );
not ( \11524_b0 , w_46081 );
and ( w_46081 , w_46080 , \11524_b1 );
or ( \11530_b1 , \11527_b1 , w_46084 );
or ( \11530_b0 , \11527_b0 , w_46083 );
not ( w_46083 , w_46085 );
and ( w_46085 , w_46084 , w_46082 );
or ( w_46082 , \11528_b1 , w_46086 );
or ( w_46083 , \11528_b0 , \11529_b0 );
not ( \11529_b0 , w_46087 );
and ( w_46087 , w_46086 , \11529_b1 );
or ( \11536_b1 , \11533_b1 , w_46090 );
or ( \11536_b0 , \11533_b0 , w_46089 );
not ( w_46089 , w_46091 );
and ( w_46091 , w_46090 , w_46088 );
or ( w_46088 , \11534_b1 , w_46092 );
or ( w_46089 , \11534_b0 , \11535_b0 );
not ( \11535_b0 , w_46093 );
and ( w_46093 , w_46092 , \11535_b1 );
or ( \11596_b1 , \11593_b1 , w_46096 );
or ( \11596_b0 , \11593_b0 , w_46095 );
not ( w_46095 , w_46097 );
and ( w_46097 , w_46096 , w_46094 );
or ( w_46094 , \11594_b1 , w_46098 );
or ( w_46095 , \11594_b0 , \11595_b0 );
not ( \11595_b0 , w_46099 );
and ( w_46099 , w_46098 , \11595_b1 );
or ( \11600_b1 , \11597_b1 , w_46102 );
or ( \11600_b0 , \11597_b0 , w_46101 );
not ( w_46101 , w_46103 );
and ( w_46103 , w_46102 , w_46100 );
or ( w_46100 , \11598_b1 , w_46104 );
or ( w_46101 , \11598_b0 , \11599_b0 );
not ( \11599_b0 , w_46105 );
and ( w_46105 , w_46104 , \11599_b1 );
or ( \11605_b1 , \11602_b1 , w_46108 );
or ( \11605_b0 , \11602_b0 , w_46107 );
not ( w_46107 , w_46109 );
and ( w_46109 , w_46108 , w_46106 );
or ( w_46106 , \11603_b1 , w_46110 );
or ( w_46107 , \11603_b0 , \11604_b0 );
not ( \11604_b0 , w_46111 );
and ( w_46111 , w_46110 , \11604_b1 );
or ( \11613_b1 , \11610_b1 , w_46114 );
or ( \11613_b0 , \11610_b0 , w_46113 );
not ( w_46113 , w_46115 );
and ( w_46115 , w_46114 , w_46112 );
or ( w_46112 , \11611_b1 , w_46116 );
or ( w_46113 , \11611_b0 , \11612_b0 );
not ( \11612_b0 , w_46117 );
and ( w_46117 , w_46116 , \11612_b1 );
or ( \11621_b1 , \11618_b1 , w_46120 );
or ( \11621_b0 , \11618_b0 , w_46119 );
not ( w_46119 , w_46121 );
and ( w_46121 , w_46120 , w_46118 );
or ( w_46118 , \11619_b1 , w_46122 );
or ( w_46119 , \11619_b0 , \11620_b0 );
not ( \11620_b0 , w_46123 );
and ( w_46123 , w_46122 , \11620_b1 );
or ( \11625_b1 , \11622_b1 , w_46126 );
or ( \11625_b0 , \11622_b0 , w_46125 );
not ( w_46125 , w_46127 );
and ( w_46127 , w_46126 , w_46124 );
or ( w_46124 , \11623_b1 , w_46128 );
or ( w_46125 , \11623_b0 , \11624_b0 );
not ( \11624_b0 , w_46129 );
and ( w_46129 , w_46128 , \11624_b1 );
or ( \11629_b1 , \11626_b1 , w_46132 );
or ( \11629_b0 , \11626_b0 , w_46131 );
not ( w_46131 , w_46133 );
and ( w_46133 , w_46132 , w_46130 );
or ( w_46130 , \11627_b1 , w_46134 );
or ( w_46131 , \11627_b0 , \11628_b0 );
not ( \11628_b0 , w_46135 );
and ( w_46135 , w_46134 , \11628_b1 );
or ( \11634_b1 , \11631_b1 , w_46138 );
or ( \11634_b0 , \11631_b0 , w_46137 );
not ( w_46137 , w_46139 );
and ( w_46139 , w_46138 , w_46136 );
or ( w_46136 , \11632_b1 , w_46140 );
or ( w_46137 , \11632_b0 , \11633_b0 );
not ( \11633_b0 , w_46141 );
and ( w_46141 , w_46140 , \11633_b1 );
or ( \11640_b1 , \11637_b1 , w_46144 );
or ( \11640_b0 , \11637_b0 , w_46143 );
not ( w_46143 , w_46145 );
and ( w_46145 , w_46144 , w_46142 );
or ( w_46142 , \11638_b1 , w_46146 );
or ( w_46143 , \11638_b0 , \11639_b0 );
not ( \11639_b0 , w_46147 );
and ( w_46147 , w_46146 , \11639_b1 );
or ( \11644_b1 , \11641_b1 , w_46150 );
or ( \11644_b0 , \11641_b0 , w_46149 );
not ( w_46149 , w_46151 );
and ( w_46151 , w_46150 , w_46148 );
or ( w_46148 , \11642_b1 , w_46152 );
or ( w_46149 , \11642_b0 , \11643_b0 );
not ( \11643_b0 , w_46153 );
and ( w_46153 , w_46152 , \11643_b1 );
or ( \11649_b1 , \11646_b1 , w_46156 );
or ( \11649_b0 , \11646_b0 , w_46155 );
not ( w_46155 , w_46157 );
and ( w_46157 , w_46156 , w_46154 );
or ( w_46154 , \11647_b1 , w_46158 );
or ( w_46155 , \11647_b0 , \11648_b0 );
not ( \11648_b0 , w_46159 );
and ( w_46159 , w_46158 , \11648_b1 );
or ( \11653_b1 , \11650_b1 , w_46162 );
or ( \11653_b0 , \11650_b0 , w_46161 );
not ( w_46161 , w_46163 );
and ( w_46163 , w_46162 , w_46160 );
or ( w_46160 , \11651_b1 , w_46164 );
or ( w_46161 , \11651_b0 , \11652_b0 );
not ( \11652_b0 , w_46165 );
and ( w_46165 , w_46164 , \11652_b1 );
or ( \11658_b1 , \11655_b1 , w_46168 );
or ( \11658_b0 , \11655_b0 , w_46167 );
not ( w_46167 , w_46169 );
and ( w_46169 , w_46168 , w_46166 );
or ( w_46166 , \11656_b1 , w_46170 );
or ( w_46167 , \11656_b0 , \11657_b0 );
not ( \11657_b0 , w_46171 );
and ( w_46171 , w_46170 , \11657_b1 );
or ( \11663_b1 , \11660_b1 , w_46174 );
or ( \11663_b0 , \11660_b0 , w_46173 );
not ( w_46173 , w_46175 );
and ( w_46175 , w_46174 , w_46172 );
or ( w_46172 , \11661_b1 , w_46176 );
or ( w_46173 , \11661_b0 , \11662_b0 );
not ( \11662_b0 , w_46177 );
and ( w_46177 , w_46176 , \11662_b1 );
or ( \11667_b1 , \11664_b1 , w_46180 );
or ( \11667_b0 , \11664_b0 , w_46179 );
not ( w_46179 , w_46181 );
and ( w_46181 , w_46180 , w_46178 );
or ( w_46178 , \11665_b1 , w_46182 );
or ( w_46179 , \11665_b0 , \11666_b0 );
not ( \11666_b0 , w_46183 );
and ( w_46183 , w_46182 , \11666_b1 );
or ( \11672_b1 , \11669_b1 , w_46186 );
or ( \11672_b0 , \11669_b0 , w_46185 );
not ( w_46185 , w_46187 );
and ( w_46187 , w_46186 , w_46184 );
or ( w_46184 , \11670_b1 , w_46188 );
or ( w_46185 , \11670_b0 , \11671_b0 );
not ( \11671_b0 , w_46189 );
and ( w_46189 , w_46188 , \11671_b1 );
or ( \11678_b1 , \11675_b1 , w_46192 );
or ( \11678_b0 , \11675_b0 , w_46191 );
not ( w_46191 , w_46193 );
and ( w_46193 , w_46192 , w_46190 );
or ( w_46190 , \11676_b1 , w_46194 );
or ( w_46191 , \11676_b0 , \11677_b0 );
not ( \11677_b0 , w_46195 );
and ( w_46195 , w_46194 , \11677_b1 );
or ( \11765_b1 , \11762_b1 , w_46198 );
or ( \11765_b0 , \11762_b0 , w_46197 );
not ( w_46197 , w_46199 );
and ( w_46199 , w_46198 , w_46196 );
or ( w_46196 , \11763_b1 , w_46200 );
or ( w_46197 , \11763_b0 , \11764_b0 );
not ( \11764_b0 , w_46201 );
and ( w_46201 , w_46200 , \11764_b1 );
or ( \11769_b1 , \11766_b1 , w_46204 );
or ( \11769_b0 , \11766_b0 , w_46203 );
not ( w_46203 , w_46205 );
and ( w_46205 , w_46204 , w_46202 );
or ( w_46202 , \11767_b1 , w_46206 );
or ( w_46203 , \11767_b0 , \11768_b0 );
not ( \11768_b0 , w_46207 );
and ( w_46207 , w_46206 , \11768_b1 );
or ( \11779_b1 , \11776_b1 , w_46210 );
or ( \11779_b0 , \11776_b0 , w_46209 );
not ( w_46209 , w_46211 );
and ( w_46211 , w_46210 , w_46208 );
or ( w_46208 , \11777_b1 , w_46212 );
or ( w_46209 , \11777_b0 , \11778_b0 );
not ( \11778_b0 , w_46213 );
and ( w_46213 , w_46212 , \11778_b1 );
or ( \11784_b1 , \11781_b1 , w_46216 );
or ( \11784_b0 , \11781_b0 , w_46215 );
not ( w_46215 , w_46217 );
and ( w_46217 , w_46216 , w_46214 );
or ( w_46214 , \11782_b1 , w_46218 );
or ( w_46215 , \11782_b0 , \11783_b0 );
not ( \11783_b0 , w_46219 );
and ( w_46219 , w_46218 , \11783_b1 );
or ( \11788_b1 , \11785_b1 , w_46222 );
or ( \11788_b0 , \11785_b0 , w_46221 );
not ( w_46221 , w_46223 );
and ( w_46223 , w_46222 , w_46220 );
or ( w_46220 , \11786_b1 , w_46224 );
or ( w_46221 , \11786_b0 , \11787_b0 );
not ( \11787_b0 , w_46225 );
and ( w_46225 , w_46224 , \11787_b1 );
or ( \11792_b1 , \11789_b1 , w_46228 );
or ( \11792_b0 , \11789_b0 , w_46227 );
not ( w_46227 , w_46229 );
and ( w_46229 , w_46228 , w_46226 );
or ( w_46226 , \11790_b1 , w_46230 );
or ( w_46227 , \11790_b0 , \11791_b0 );
not ( \11791_b0 , w_46231 );
and ( w_46231 , w_46230 , \11791_b1 );
or ( \11800_b1 , \11797_b1 , w_46234 );
or ( \11800_b0 , \11797_b0 , w_46233 );
not ( w_46233 , w_46235 );
and ( w_46235 , w_46234 , w_46232 );
or ( w_46232 , \11798_b1 , w_46236 );
or ( w_46233 , \11798_b0 , \11799_b0 );
not ( \11799_b0 , w_46237 );
and ( w_46237 , w_46236 , \11799_b1 );
or ( \11804_b1 , \11801_b1 , w_46240 );
or ( \11804_b0 , \11801_b0 , w_46239 );
not ( w_46239 , w_46241 );
and ( w_46241 , w_46240 , w_46238 );
or ( w_46238 , \11802_b1 , w_46242 );
or ( w_46239 , \11802_b0 , \11803_b0 );
not ( \11803_b0 , w_46243 );
and ( w_46243 , w_46242 , \11803_b1 );
or ( \11836_b1 , \11833_b1 , w_46246 );
or ( \11836_b0 , \11833_b0 , w_46245 );
not ( w_46245 , w_46247 );
and ( w_46247 , w_46246 , w_46244 );
or ( w_46244 , \11834_b1 , w_46248 );
or ( w_46245 , \11834_b0 , \11835_b0 );
not ( \11835_b0 , w_46249 );
and ( w_46249 , w_46248 , \11835_b1 );
or ( \11840_b1 , \11837_b1 , w_46252 );
or ( \11840_b0 , \11837_b0 , w_46251 );
not ( w_46251 , w_46253 );
and ( w_46253 , w_46252 , w_46250 );
or ( w_46250 , \11838_b1 , w_46254 );
or ( w_46251 , \11838_b0 , \11839_b0 );
not ( \11839_b0 , w_46255 );
and ( w_46255 , w_46254 , \11839_b1 );
or ( \11848_b1 , \11845_b1 , w_46258 );
or ( \11848_b0 , \11845_b0 , w_46257 );
not ( w_46257 , w_46259 );
and ( w_46259 , w_46258 , w_46256 );
or ( w_46256 , \11846_b1 , w_46260 );
or ( w_46257 , \11846_b0 , \11847_b0 );
not ( \11847_b0 , w_46261 );
and ( w_46261 , w_46260 , \11847_b1 );
or ( \11852_b1 , \11849_b1 , w_46264 );
or ( \11852_b0 , \11849_b0 , w_46263 );
not ( w_46263 , w_46265 );
and ( w_46265 , w_46264 , w_46262 );
or ( w_46262 , \11850_b1 , w_46266 );
or ( w_46263 , \11850_b0 , \11851_b0 );
not ( \11851_b0 , w_46267 );
and ( w_46267 , w_46266 , \11851_b1 );
or ( \11857_b1 , \11854_b1 , w_46270 );
or ( \11857_b0 , \11854_b0 , w_46269 );
not ( w_46269 , w_46271 );
and ( w_46271 , w_46270 , w_46268 );
or ( w_46268 , \11855_b1 , w_46272 );
or ( w_46269 , \11855_b0 , \11856_b0 );
not ( \11856_b0 , w_46273 );
and ( w_46273 , w_46272 , \11856_b1 );
or ( \11863_b1 , \11860_b1 , w_46276 );
or ( \11863_b0 , \11860_b0 , w_46275 );
not ( w_46275 , w_46277 );
and ( w_46277 , w_46276 , w_46274 );
or ( w_46274 , \11861_b1 , w_46278 );
or ( w_46275 , \11861_b0 , \11862_b0 );
not ( \11862_b0 , w_46279 );
and ( w_46279 , w_46278 , \11862_b1 );
or ( \11923_b1 , \11920_b1 , w_46282 );
or ( \11923_b0 , \11920_b0 , w_46281 );
not ( w_46281 , w_46283 );
and ( w_46283 , w_46282 , w_46280 );
or ( w_46280 , \11921_b1 , w_46284 );
or ( w_46281 , \11921_b0 , \11922_b0 );
not ( \11922_b0 , w_46285 );
and ( w_46285 , w_46284 , \11922_b1 );
or ( \11927_b1 , \11924_b1 , w_46288 );
or ( \11927_b0 , \11924_b0 , w_46287 );
not ( w_46287 , w_46289 );
and ( w_46289 , w_46288 , w_46286 );
or ( w_46286 , \11925_b1 , w_46290 );
or ( w_46287 , \11925_b0 , \11926_b0 );
not ( \11926_b0 , w_46291 );
and ( w_46291 , w_46290 , \11926_b1 );
or ( \11932_b1 , \11929_b1 , w_46294 );
or ( \11932_b0 , \11929_b0 , w_46293 );
not ( w_46293 , w_46295 );
and ( w_46295 , w_46294 , w_46292 );
or ( w_46292 , \11930_b1 , w_46296 );
or ( w_46293 , \11930_b0 , \11931_b0 );
not ( \11931_b0 , w_46297 );
and ( w_46297 , w_46296 , \11931_b1 );
or ( \11940_b1 , \11937_b1 , w_46300 );
or ( \11940_b0 , \11937_b0 , w_46299 );
not ( w_46299 , w_46301 );
and ( w_46301 , w_46300 , w_46298 );
or ( w_46298 , \11938_b1 , w_46302 );
or ( w_46299 , \11938_b0 , \11939_b0 );
not ( \11939_b0 , w_46303 );
and ( w_46303 , w_46302 , \11939_b1 );
or ( \11946_b1 , \11943_b1 , w_46306 );
or ( \11946_b0 , \11943_b0 , w_46305 );
not ( w_46305 , w_46307 );
and ( w_46307 , w_46306 , w_46304 );
or ( w_46304 , \11944_b1 , w_46308 );
or ( w_46305 , \11944_b0 , \11945_b0 );
not ( \11945_b0 , w_46309 );
and ( w_46309 , w_46308 , \11945_b1 );
or ( \11950_b1 , \11947_b1 , w_46312 );
or ( \11950_b0 , \11947_b0 , w_46311 );
not ( w_46311 , w_46313 );
and ( w_46313 , w_46312 , w_46310 );
or ( w_46310 , \11948_b1 , w_46314 );
or ( w_46311 , \11948_b0 , \11949_b0 );
not ( \11949_b0 , w_46315 );
and ( w_46315 , w_46314 , \11949_b1 );
or ( \11954_b1 , \11951_b1 , w_46318 );
or ( \11954_b0 , \11951_b0 , w_46317 );
not ( w_46317 , w_46319 );
and ( w_46319 , w_46318 , w_46316 );
or ( w_46316 , \11952_b1 , w_46320 );
or ( w_46317 , \11952_b0 , \11953_b0 );
not ( \11953_b0 , w_46321 );
and ( w_46321 , w_46320 , \11953_b1 );
or ( \11959_b1 , \11956_b1 , w_46324 );
or ( \11959_b0 , \11956_b0 , w_46323 );
not ( w_46323 , w_46325 );
and ( w_46325 , w_46324 , w_46322 );
or ( w_46322 , \11957_b1 , w_46326 );
or ( w_46323 , \11957_b0 , \11958_b0 );
not ( \11958_b0 , w_46327 );
and ( w_46327 , w_46326 , \11958_b1 );
or ( \11965_b1 , \11962_b1 , w_46330 );
or ( \11965_b0 , \11962_b0 , w_46329 );
not ( w_46329 , w_46331 );
and ( w_46331 , w_46330 , w_46328 );
or ( w_46328 , \11963_b1 , w_46332 );
or ( w_46329 , \11963_b0 , \11964_b0 );
not ( \11964_b0 , w_46333 );
and ( w_46333 , w_46332 , \11964_b1 );
or ( \11969_b1 , \11966_b1 , w_46336 );
or ( \11969_b0 , \11966_b0 , w_46335 );
not ( w_46335 , w_46337 );
and ( w_46337 , w_46336 , w_46334 );
or ( w_46334 , \11967_b1 , w_46338 );
or ( w_46335 , \11967_b0 , \11968_b0 );
not ( \11968_b0 , w_46339 );
and ( w_46339 , w_46338 , \11968_b1 );
or ( \11974_b1 , \11971_b1 , w_46342 );
or ( \11974_b0 , \11971_b0 , w_46341 );
not ( w_46341 , w_46343 );
and ( w_46343 , w_46342 , w_46340 );
or ( w_46340 , \11972_b1 , w_46344 );
or ( w_46341 , \11972_b0 , \11973_b0 );
not ( \11973_b0 , w_46345 );
and ( w_46345 , w_46344 , \11973_b1 );
or ( \11978_b1 , \11975_b1 , w_46348 );
or ( \11978_b0 , \11975_b0 , w_46347 );
not ( w_46347 , w_46349 );
and ( w_46349 , w_46348 , w_46346 );
or ( w_46346 , \11976_b1 , w_46350 );
or ( w_46347 , \11976_b0 , \11977_b0 );
not ( \11977_b0 , w_46351 );
and ( w_46351 , w_46350 , \11977_b1 );
or ( \11983_b1 , \11980_b1 , w_46354 );
or ( \11983_b0 , \11980_b0 , w_46353 );
not ( w_46353 , w_46355 );
and ( w_46355 , w_46354 , w_46352 );
or ( w_46352 , \11981_b1 , w_46356 );
or ( w_46353 , \11981_b0 , \11982_b0 );
not ( \11982_b0 , w_46357 );
and ( w_46357 , w_46356 , \11982_b1 );
or ( \11988_b1 , \11985_b1 , w_46360 );
or ( \11988_b0 , \11985_b0 , w_46359 );
not ( w_46359 , w_46361 );
and ( w_46361 , w_46360 , w_46358 );
or ( w_46358 , \11986_b1 , w_46362 );
or ( w_46359 , \11986_b0 , \11987_b0 );
not ( \11987_b0 , w_46363 );
and ( w_46363 , w_46362 , \11987_b1 );
or ( \11992_b1 , \11989_b1 , w_46366 );
or ( \11992_b0 , \11989_b0 , w_46365 );
not ( w_46365 , w_46367 );
and ( w_46367 , w_46366 , w_46364 );
or ( w_46364 , \11990_b1 , w_46368 );
or ( w_46365 , \11990_b0 , \11991_b0 );
not ( \11991_b0 , w_46369 );
and ( w_46369 , w_46368 , \11991_b1 );
or ( \11997_b1 , \11994_b1 , w_46372 );
or ( \11997_b0 , \11994_b0 , w_46371 );
not ( w_46371 , w_46373 );
and ( w_46373 , w_46372 , w_46370 );
or ( w_46370 , \11995_b1 , w_46374 );
or ( w_46371 , \11995_b0 , \11996_b0 );
not ( \11996_b0 , w_46375 );
and ( w_46375 , w_46374 , \11996_b1 );
or ( \12003_b1 , \12000_b1 , w_46378 );
or ( \12003_b0 , \12000_b0 , w_46377 );
not ( w_46377 , w_46379 );
and ( w_46379 , w_46378 , w_46376 );
or ( w_46376 , \12001_b1 , w_46380 );
or ( w_46377 , \12001_b0 , \12002_b0 );
not ( \12002_b0 , w_46381 );
and ( w_46381 , w_46380 , \12002_b1 );
or ( \12025_b1 , \12022_b1 , w_46384 );
or ( \12025_b0 , \12022_b0 , w_46383 );
not ( w_46383 , w_46385 );
and ( w_46385 , w_46384 , w_46382 );
or ( w_46382 , \12023_b1 , w_46386 );
or ( w_46383 , \12023_b0 , \12024_b0 );
not ( \12024_b0 , w_46387 );
and ( w_46387 , w_46386 , \12024_b1 );
or ( \12029_b1 , \12026_b1 , w_46390 );
or ( \12029_b0 , \12026_b0 , w_46389 );
not ( w_46389 , w_46391 );
and ( w_46391 , w_46390 , w_46388 );
or ( w_46388 , \12027_b1 , w_46392 );
or ( w_46389 , \12027_b0 , \12028_b0 );
not ( \12028_b0 , w_46393 );
and ( w_46393 , w_46392 , \12028_b1 );
or ( \12039_b1 , \12036_b1 , w_46396 );
or ( \12039_b0 , \12036_b0 , w_46395 );
not ( w_46395 , w_46397 );
and ( w_46397 , w_46396 , w_46394 );
or ( w_46394 , \12037_b1 , w_46398 );
or ( w_46395 , \12037_b0 , \12038_b0 );
not ( \12038_b0 , w_46399 );
and ( w_46399 , w_46398 , \12038_b1 );
or ( \12044_b1 , \12041_b1 , w_46402 );
or ( \12044_b0 , \12041_b0 , w_46401 );
not ( w_46401 , w_46403 );
and ( w_46403 , w_46402 , w_46400 );
or ( w_46400 , \12042_b1 , w_46404 );
or ( w_46401 , \12042_b0 , \12043_b0 );
not ( \12043_b0 , w_46405 );
and ( w_46405 , w_46404 , \12043_b1 );
or ( \12048_b1 , \12045_b1 , w_46408 );
or ( \12048_b0 , \12045_b0 , w_46407 );
not ( w_46407 , w_46409 );
and ( w_46409 , w_46408 , w_46406 );
or ( w_46406 , \12046_b1 , w_46410 );
or ( w_46407 , \12046_b0 , \12047_b0 );
not ( \12047_b0 , w_46411 );
and ( w_46411 , w_46410 , \12047_b1 );
or ( \12052_b1 , \12049_b1 , w_46414 );
or ( \12052_b0 , \12049_b0 , w_46413 );
not ( w_46413 , w_46415 );
and ( w_46415 , w_46414 , w_46412 );
or ( w_46412 , \12050_b1 , w_46416 );
or ( w_46413 , \12050_b0 , \12051_b0 );
not ( \12051_b0 , w_46417 );
and ( w_46417 , w_46416 , \12051_b1 );
or ( \12060_b1 , \12057_b1 , w_46420 );
or ( \12060_b0 , \12057_b0 , w_46419 );
not ( w_46419 , w_46421 );
and ( w_46421 , w_46420 , w_46418 );
or ( w_46418 , \12058_b1 , w_46422 );
or ( w_46419 , \12058_b0 , \12059_b0 );
not ( \12059_b0 , w_46423 );
and ( w_46423 , w_46422 , \12059_b1 );
or ( \12064_b1 , \12061_b1 , w_46426 );
or ( \12064_b0 , \12061_b0 , w_46425 );
not ( w_46425 , w_46427 );
and ( w_46427 , w_46426 , w_46424 );
or ( w_46424 , \12062_b1 , w_46428 );
or ( w_46425 , \12062_b0 , \12063_b0 );
not ( \12063_b0 , w_46429 );
and ( w_46429 , w_46428 , \12063_b1 );
or ( \12076_b1 , \12073_b1 , w_46432 );
or ( \12076_b0 , \12073_b0 , w_46431 );
not ( w_46431 , w_46433 );
and ( w_46433 , w_46432 , w_46430 );
or ( w_46430 , \12074_b1 , w_46434 );
or ( w_46431 , \12074_b0 , \12075_b0 );
not ( \12075_b0 , w_46435 );
and ( w_46435 , w_46434 , \12075_b1 );
or ( \12087_b1 , \12084_b1 , w_46438 );
or ( \12087_b0 , \12084_b0 , w_46437 );
not ( w_46437 , w_46439 );
and ( w_46439 , w_46438 , w_46436 );
or ( w_46436 , \12085_b1 , w_46440 );
or ( w_46437 , \12085_b0 , \12086_b0 );
not ( \12086_b0 , w_46441 );
and ( w_46441 , w_46440 , \12086_b1 );
or ( \12091_b1 , \12088_b1 , w_46444 );
or ( \12091_b0 , \12088_b0 , w_46443 );
not ( w_46443 , w_46445 );
and ( w_46445 , w_46444 , w_46442 );
or ( w_46442 , \12089_b1 , w_46446 );
or ( w_46443 , \12089_b0 , \12090_b0 );
not ( \12090_b0 , w_46447 );
and ( w_46447 , w_46446 , \12090_b1 );
or ( \12096_b1 , \12093_b1 , w_46450 );
or ( \12096_b0 , \12093_b0 , w_46449 );
not ( w_46449 , w_46451 );
and ( w_46451 , w_46450 , w_46448 );
or ( w_46448 , \12094_b1 , w_46452 );
or ( w_46449 , \12094_b0 , \12095_b0 );
not ( \12095_b0 , w_46453 );
and ( w_46453 , w_46452 , \12095_b1 );
or ( \12104_b1 , \12101_b1 , w_46456 );
or ( \12104_b0 , \12101_b0 , w_46455 );
not ( w_46455 , w_46457 );
and ( w_46457 , w_46456 , w_46454 );
or ( w_46454 , \12102_b1 , w_46458 );
or ( w_46455 , \12102_b0 , \12103_b0 );
not ( \12103_b0 , w_46459 );
and ( w_46459 , w_46458 , \12103_b1 );
or ( \12111_b1 , \12108_b1 , w_46462 );
or ( \12111_b0 , \12108_b0 , w_46461 );
not ( w_46461 , w_46463 );
and ( w_46463 , w_46462 , w_46460 );
or ( w_46460 , \12109_b1 , w_46464 );
or ( w_46461 , \12109_b0 , \12110_b0 );
not ( \12110_b0 , w_46465 );
and ( w_46465 , w_46464 , \12110_b1 );
or ( \12115_b1 , \12112_b1 , w_46468 );
or ( \12115_b0 , \12112_b0 , w_46467 );
not ( w_46467 , w_46469 );
and ( w_46469 , w_46468 , w_46466 );
or ( w_46466 , \12113_b1 , w_46470 );
or ( w_46467 , \12113_b0 , \12114_b0 );
not ( \12114_b0 , w_46471 );
and ( w_46471 , w_46470 , \12114_b1 );
or ( \12119_b1 , \12116_b1 , w_46474 );
or ( \12119_b0 , \12116_b0 , w_46473 );
not ( w_46473 , w_46475 );
and ( w_46475 , w_46474 , w_46472 );
or ( w_46472 , \12117_b1 , w_46476 );
or ( w_46473 , \12117_b0 , \12118_b0 );
not ( \12118_b0 , w_46477 );
and ( w_46477 , w_46476 , \12118_b1 );
or ( \12124_b1 , \12121_b1 , w_46480 );
or ( \12124_b0 , \12121_b0 , w_46479 );
not ( w_46479 , w_46481 );
and ( w_46481 , w_46480 , w_46478 );
or ( w_46478 , \12122_b1 , w_46482 );
or ( w_46479 , \12122_b0 , \12123_b0 );
not ( \12123_b0 , w_46483 );
and ( w_46483 , w_46482 , \12123_b1 );
or ( \12130_b1 , \12127_b1 , w_46486 );
or ( \12130_b0 , \12127_b0 , w_46485 );
not ( w_46485 , w_46487 );
and ( w_46487 , w_46486 , w_46484 );
or ( w_46484 , \12128_b1 , w_46488 );
or ( w_46485 , \12128_b0 , \12129_b0 );
not ( \12129_b0 , w_46489 );
and ( w_46489 , w_46488 , \12129_b1 );
or ( \12134_b1 , \12131_b1 , w_46492 );
or ( \12134_b0 , \12131_b0 , w_46491 );
not ( w_46491 , w_46493 );
and ( w_46493 , w_46492 , w_46490 );
or ( w_46490 , \12132_b1 , w_46494 );
or ( w_46491 , \12132_b0 , \12133_b0 );
not ( \12133_b0 , w_46495 );
and ( w_46495 , w_46494 , \12133_b1 );
or ( \12148_b1 , \12145_b1 , w_46498 );
or ( \12148_b0 , \12145_b0 , w_46497 );
not ( w_46497 , w_46499 );
and ( w_46499 , w_46498 , w_46496 );
or ( w_46496 , \12146_b1 , w_46500 );
or ( w_46497 , \12146_b0 , \12147_b0 );
not ( \12147_b0 , w_46501 );
and ( w_46501 , w_46500 , \12147_b1 );
or ( \12153_b1 , \12150_b1 , w_46504 );
or ( \12153_b0 , \12150_b0 , w_46503 );
not ( w_46503 , w_46505 );
and ( w_46505 , w_46504 , w_46502 );
or ( w_46502 , \12151_b1 , w_46506 );
or ( w_46503 , \12151_b0 , \12152_b0 );
not ( \12152_b0 , w_46507 );
and ( w_46507 , w_46506 , \12152_b1 );
or ( \12160_b1 , \12157_b1 , w_46510 );
or ( \12160_b0 , \12157_b0 , w_46509 );
not ( w_46509 , w_46511 );
and ( w_46511 , w_46510 , w_46508 );
or ( w_46508 , \12158_b1 , w_46512 );
or ( w_46509 , \12158_b0 , \12159_b0 );
not ( \12159_b0 , w_46513 );
and ( w_46513 , w_46512 , \12159_b1 );
or ( \12164_b1 , \12161_b1 , w_46516 );
or ( \12164_b0 , \12161_b0 , w_46515 );
not ( w_46515 , w_46517 );
and ( w_46517 , w_46516 , w_46514 );
or ( w_46514 , \12162_b1 , w_46518 );
or ( w_46515 , \12162_b0 , \12163_b0 );
not ( \12163_b0 , w_46519 );
and ( w_46519 , w_46518 , \12163_b1 );
or ( \12173_b1 , \12170_b1 , w_46522 );
or ( \12173_b0 , \12170_b0 , w_46521 );
not ( w_46521 , w_46523 );
and ( w_46523 , w_46522 , w_46520 );
or ( w_46520 , \12171_b1 , w_46524 );
or ( w_46521 , \12171_b0 , \12172_b0 );
not ( \12172_b0 , w_46525 );
and ( w_46525 , w_46524 , \12172_b1 );
or ( \12179_b1 , \12176_b1 , w_46528 );
or ( \12179_b0 , \12176_b0 , w_46527 );
not ( w_46527 , w_46529 );
and ( w_46529 , w_46528 , w_46526 );
or ( w_46526 , \12177_b1 , w_46530 );
or ( w_46527 , \12177_b0 , \12178_b0 );
not ( \12178_b0 , w_46531 );
and ( w_46531 , w_46530 , \12178_b1 );
or ( \12189_b1 , \12186_b1 , w_46534 );
or ( \12189_b0 , \12186_b0 , w_46533 );
not ( w_46533 , w_46535 );
and ( w_46535 , w_46534 , w_46532 );
or ( w_46532 , \12187_b1 , w_46536 );
or ( w_46533 , \12187_b0 , \12188_b0 );
not ( \12188_b0 , w_46537 );
and ( w_46537 , w_46536 , \12188_b1 );
or ( \12196_b1 , \12193_b1 , w_46540 );
or ( \12196_b0 , \12193_b0 , w_46539 );
not ( w_46539 , w_46541 );
and ( w_46541 , w_46540 , w_46538 );
or ( w_46538 , \12194_b1 , w_46542 );
or ( w_46539 , \12194_b0 , \12195_b0 );
not ( \12195_b0 , w_46543 );
and ( w_46543 , w_46542 , \12195_b1 );
or ( \12214_b1 , \12207_b1 , w_46546 );
or ( \12214_b0 , \12207_b0 , w_46545 );
not ( w_46545 , w_46547 );
and ( w_46547 , w_46546 , w_46544 );
or ( w_46544 , \12212_b1 , w_46548 );
or ( w_46545 , \12212_b0 , \12213_b0 );
not ( \12213_b0 , w_46549 );
and ( w_46549 , w_46548 , \12213_b1 );
or ( \12230_b1 , \12223_b1 , w_46552 );
or ( \12230_b0 , \12223_b0 , w_46551 );
not ( w_46551 , w_46553 );
and ( w_46553 , w_46552 , w_46550 );
or ( w_46550 , \12228_b1 , w_46554 );
or ( w_46551 , \12228_b0 , \12229_b0 );
not ( \12229_b0 , w_46555 );
and ( w_46555 , w_46554 , \12229_b1 );
or ( \12238_b1 , \12231_b1 , w_46558 );
or ( \12238_b0 , \12231_b0 , w_46557 );
not ( w_46557 , w_46559 );
and ( w_46559 , w_46558 , w_46556 );
or ( w_46556 , \12236_b1 , w_46560 );
or ( w_46557 , \12236_b0 , \12237_b0 );
not ( \12237_b0 , w_46561 );
and ( w_46561 , w_46560 , \12237_b1 );
or ( \12280_b1 , \12273_b1 , w_46564 );
or ( \12280_b0 , \12273_b0 , w_46563 );
not ( w_46563 , w_46565 );
and ( w_46565 , w_46564 , w_46562 );
or ( w_46562 , \12278_b1 , w_46566 );
or ( w_46563 , \12278_b0 , \12279_b0 );
not ( \12279_b0 , w_46567 );
and ( w_46567 , w_46566 , \12279_b1 );
or ( \12296_b1 , \12289_b1 , w_46570 );
or ( \12296_b0 , \12289_b0 , w_46569 );
not ( w_46569 , w_46571 );
and ( w_46571 , w_46570 , w_46568 );
or ( w_46568 , \12294_b1 , w_46572 );
or ( w_46569 , \12294_b0 , \12295_b0 );
not ( \12295_b0 , w_46573 );
and ( w_46573 , w_46572 , \12295_b1 );
or ( \12313_b1 , \12264_b1 , w_46576 );
or ( \12313_b0 , \12264_b0 , w_46575 );
not ( w_46575 , w_46577 );
and ( w_46577 , w_46576 , w_46574 );
or ( w_46574 , \12311_b1 , w_46578 );
or ( w_46575 , \12311_b0 , \12312_b0 );
not ( \12312_b0 , w_46579 );
and ( w_46579 , w_46578 , \12312_b1 );
or ( \12317_b1 , \12314_b1 , w_46582 );
or ( \12317_b0 , \12314_b0 , w_46581 );
not ( w_46581 , w_46583 );
and ( w_46583 , w_46582 , w_46580 );
or ( w_46580 , \12315_b1 , w_46584 );
or ( w_46581 , \12315_b0 , \12316_b0 );
not ( \12316_b0 , w_46585 );
and ( w_46585 , w_46584 , \12316_b1 );
or ( \12321_b1 , \12318_b1 , w_46588 );
or ( \12321_b0 , \12318_b0 , w_46587 );
not ( w_46587 , w_46589 );
and ( w_46589 , w_46588 , w_46586 );
or ( w_46586 , \12319_b1 , w_46590 );
or ( w_46587 , \12319_b0 , \12320_b0 );
not ( \12320_b0 , w_46591 );
and ( w_46591 , w_46590 , \12320_b1 );
or ( \12326_b1 , \12323_b1 , w_46594 );
or ( \12326_b0 , \12323_b0 , w_46593 );
not ( w_46593 , w_46595 );
and ( w_46595 , w_46594 , w_46592 );
or ( w_46592 , \12324_b1 , w_46596 );
or ( w_46593 , \12324_b0 , \12325_b0 );
not ( \12325_b0 , w_46597 );
and ( w_46597 , w_46596 , \12325_b1 );
or ( \12332_b1 , \12329_b1 , w_46600 );
or ( \12332_b0 , \12329_b0 , w_46599 );
not ( w_46599 , w_46601 );
and ( w_46601 , w_46600 , w_46598 );
or ( w_46598 , \12330_b1 , w_46602 );
or ( w_46599 , \12330_b0 , \12331_b0 );
not ( \12331_b0 , w_46603 );
and ( w_46603 , w_46602 , \12331_b1 );
or ( \12391_b1 , \12384_b1 , w_46606 );
or ( \12391_b0 , \12384_b0 , w_46605 );
not ( w_46605 , w_46607 );
and ( w_46607 , w_46606 , w_46604 );
or ( w_46604 , \12389_b1 , w_46608 );
or ( w_46605 , \12389_b0 , \12390_b0 );
not ( \12390_b0 , w_46609 );
and ( w_46609 , w_46608 , \12390_b1 );
or ( \12407_b1 , \12400_b1 , w_46612 );
or ( \12407_b0 , \12400_b0 , w_46611 );
not ( w_46611 , w_46613 );
and ( w_46613 , w_46612 , w_46610 );
or ( w_46610 , \12405_b1 , w_46614 );
or ( w_46611 , \12405_b0 , \12406_b0 );
not ( \12406_b0 , w_46615 );
and ( w_46615 , w_46614 , \12406_b1 );
or ( \12415_b1 , \12408_b1 , w_46618 );
or ( \12415_b0 , \12408_b0 , w_46617 );
not ( w_46617 , w_46619 );
and ( w_46619 , w_46618 , w_46616 );
or ( w_46616 , \12413_b1 , w_46620 );
or ( w_46617 , \12413_b0 , \12414_b0 );
not ( \12414_b0 , w_46621 );
and ( w_46621 , w_46620 , \12414_b1 );
or ( \12425_b1 , \12420_b1 , w_46624 );
or ( \12425_b0 , \12420_b0 , w_46623 );
not ( w_46623 , w_46625 );
and ( w_46625 , w_46624 , w_46622 );
or ( w_46622 , \12423_b1 , w_46626 );
or ( w_46623 , \12423_b0 , \12424_b0 );
not ( \12424_b0 , w_46627 );
and ( w_46627 , w_46626 , \12424_b1 );
or ( \12431_b1 , \12426_b1 , w_46630 );
or ( \12431_b0 , \12426_b0 , w_46629 );
not ( w_46629 , w_46631 );
and ( w_46631 , w_46630 , w_46628 );
or ( w_46628 , \12429_b1 , w_46632 );
or ( w_46629 , \12429_b0 , \12430_b0 );
not ( \12430_b0 , w_46633 );
and ( w_46633 , w_46632 , \12430_b1 );
or ( \12442_b1 , \12437_b1 , w_46636 );
or ( \12442_b0 , \12437_b0 , w_46635 );
not ( w_46635 , w_46637 );
and ( w_46637 , w_46636 , w_46634 );
or ( w_46634 , \12440_b1 , w_46638 );
or ( w_46635 , \12440_b0 , \12441_b0 );
not ( \12441_b0 , w_46639 );
and ( w_46639 , w_46638 , \12441_b1 );
or ( \12447_b1 , \12444_b1 , w_46642 );
or ( \12447_b0 , \12444_b0 , w_46641 );
not ( w_46641 , w_46643 );
and ( w_46643 , w_46642 , w_46640 );
or ( w_46640 , \12445_b1 , w_46644 );
or ( w_46641 , \12445_b0 , \12446_b0 );
not ( \12446_b0 , w_46645 );
and ( w_46645 , w_46644 , \12446_b1 );
or ( \12483_b1 , \12480_b1 , w_46648 );
or ( \12483_b0 , \12480_b0 , w_46647 );
not ( w_46647 , w_46649 );
and ( w_46649 , w_46648 , w_46646 );
or ( w_46646 , \12481_b1 , w_46650 );
or ( w_46647 , \12481_b0 , \12482_b0 );
not ( \12482_b0 , w_46651 );
and ( w_46651 , w_46650 , \12482_b1 );
or ( \12487_b1 , \12484_b1 , w_46654 );
or ( \12487_b0 , \12484_b0 , w_46653 );
not ( w_46653 , w_46655 );
and ( w_46655 , w_46654 , w_46652 );
or ( w_46652 , \12485_b1 , w_46656 );
or ( w_46653 , \12485_b0 , \12486_b0 );
not ( \12486_b0 , w_46657 );
and ( w_46657 , w_46656 , \12486_b1 );
or ( \12496_b1 , \12493_b1 , w_46660 );
or ( \12496_b0 , \12493_b0 , w_46659 );
not ( w_46659 , w_46661 );
and ( w_46661 , w_46660 , w_46658 );
or ( w_46658 , \12494_b1 , w_46662 );
or ( w_46659 , \12494_b0 , \12495_b0 );
not ( \12495_b0 , w_46663 );
and ( w_46663 , w_46662 , \12495_b1 );
or ( \12500_b1 , \12497_b1 , w_46666 );
or ( \12500_b0 , \12497_b0 , w_46665 );
not ( w_46665 , w_46667 );
and ( w_46667 , w_46666 , w_46664 );
or ( w_46664 , \12498_b1 , w_46668 );
or ( w_46665 , \12498_b0 , \12499_b0 );
not ( \12499_b0 , w_46669 );
and ( w_46669 , w_46668 , \12499_b1 );
or ( \12517_b1 , \12514_b1 , w_46672 );
or ( \12517_b0 , \12514_b0 , w_46671 );
not ( w_46671 , w_46673 );
and ( w_46673 , w_46672 , w_46670 );
or ( w_46670 , \12515_b1 , w_46674 );
or ( w_46671 , \12515_b0 , \12516_b0 );
not ( \12516_b0 , w_46675 );
and ( w_46675 , w_46674 , \12516_b1 );
or ( \12523_b1 , \12520_b1 , w_46678 );
or ( \12523_b0 , \12520_b0 , w_46677 );
not ( w_46677 , w_46679 );
and ( w_46679 , w_46678 , w_46676 );
or ( w_46676 , \12521_b1 , w_46680 );
or ( w_46677 , \12521_b0 , \12522_b0 );
not ( \12522_b0 , w_46681 );
and ( w_46681 , w_46680 , \12522_b1 );
or ( \12527_b1 , \12524_b1 , w_46684 );
or ( \12527_b0 , \12524_b0 , w_46683 );
not ( w_46683 , w_46685 );
and ( w_46685 , w_46684 , w_46682 );
or ( w_46682 , \12525_b1 , w_46686 );
or ( w_46683 , \12525_b0 , \12526_b0 );
not ( \12526_b0 , w_46687 );
and ( w_46687 , w_46686 , \12526_b1 );
or ( \12577_b1 , \12574_b1 , w_46690 );
or ( \12577_b0 , \12574_b0 , w_46689 );
not ( w_46689 , w_46691 );
and ( w_46691 , w_46690 , w_46688 );
or ( w_46688 , \12575_b1 , w_46692 );
or ( w_46689 , \12575_b0 , \12576_b0 );
not ( \12576_b0 , w_46693 );
and ( w_46693 , w_46692 , \12576_b1 );
or ( \12583_b1 , \12580_b1 , w_46696 );
or ( \12583_b0 , \12580_b0 , w_46695 );
not ( w_46695 , w_46697 );
and ( w_46697 , w_46696 , w_46694 );
or ( w_46694 , \12581_b1 , w_46698 );
or ( w_46695 , \12581_b0 , \12582_b0 );
not ( \12582_b0 , w_46699 );
and ( w_46699 , w_46698 , \12582_b1 );
or ( \12587_b1 , \12584_b1 , w_46702 );
or ( \12587_b0 , \12584_b0 , w_46701 );
not ( w_46701 , w_46703 );
and ( w_46703 , w_46702 , w_46700 );
or ( w_46700 , \12585_b1 , w_46704 );
or ( w_46701 , \12585_b0 , \12586_b0 );
not ( \12586_b0 , w_46705 );
and ( w_46705 , w_46704 , \12586_b1 );
or ( \12592_b1 , \12589_b1 , w_46708 );
or ( \12592_b0 , \12589_b0 , w_46707 );
not ( w_46707 , w_46709 );
and ( w_46709 , w_46708 , w_46706 );
or ( w_46706 , \12590_b1 , w_46710 );
or ( w_46707 , \12590_b0 , \12591_b0 );
not ( \12591_b0 , w_46711 );
and ( w_46711 , w_46710 , \12591_b1 );
or ( \12599_b1 , \12596_b1 , w_46714 );
or ( \12599_b0 , \12596_b0 , w_46713 );
not ( w_46713 , w_46715 );
and ( w_46715 , w_46714 , w_46712 );
or ( w_46712 , \12597_b1 , w_46716 );
or ( w_46713 , \12597_b0 , \12598_b0 );
not ( \12598_b0 , w_46717 );
and ( w_46717 , w_46716 , \12598_b1 );
or ( \12604_b1 , \12601_b1 , w_46720 );
or ( \12604_b0 , \12601_b0 , w_46719 );
not ( w_46719 , w_46721 );
and ( w_46721 , w_46720 , w_46718 );
or ( w_46718 , \12602_b1 , w_46722 );
or ( w_46719 , \12602_b0 , \12603_b0 );
not ( \12603_b0 , w_46723 );
and ( w_46723 , w_46722 , \12603_b1 );
or ( \12608_b1 , \12605_b1 , w_46726 );
or ( \12608_b0 , \12605_b0 , w_46725 );
not ( w_46725 , w_46727 );
and ( w_46727 , w_46726 , w_46724 );
or ( w_46724 , \12606_b1 , w_46728 );
or ( w_46725 , \12606_b0 , \12607_b0 );
not ( \12607_b0 , w_46729 );
and ( w_46729 , w_46728 , \12607_b1 );
or ( \12645_b1 , \12642_b1 , w_46732 );
or ( \12645_b0 , \12642_b0 , w_46731 );
not ( w_46731 , w_46733 );
and ( w_46733 , w_46732 , w_46730 );
or ( w_46730 , \12643_b1 , w_46734 );
or ( w_46731 , \12643_b0 , \12644_b0 );
not ( \12644_b0 , w_46735 );
and ( w_46735 , w_46734 , \12644_b1 );
or ( \12649_b1 , \12646_b1 , w_46738 );
or ( \12649_b0 , \12646_b0 , w_46737 );
not ( w_46737 , w_46739 );
and ( w_46739 , w_46738 , w_46736 );
or ( w_46736 , \12647_b1 , w_46740 );
or ( w_46737 , \12647_b0 , \12648_b0 );
not ( \12648_b0 , w_46741 );
and ( w_46741 , w_46740 , \12648_b1 );
or ( \12654_b1 , \12651_b1 , w_46744 );
or ( \12654_b0 , \12651_b0 , w_46743 );
not ( w_46743 , w_46745 );
and ( w_46745 , w_46744 , w_46742 );
or ( w_46742 , \12652_b1 , w_46746 );
or ( w_46743 , \12652_b0 , \12653_b0 );
not ( \12653_b0 , w_46747 );
and ( w_46747 , w_46746 , \12653_b1 );
or ( \12661_b1 , \12658_b1 , w_46750 );
or ( \12661_b0 , \12658_b0 , w_46749 );
not ( w_46749 , w_46751 );
and ( w_46751 , w_46750 , w_46748 );
or ( w_46748 , \12659_b1 , w_46752 );
or ( w_46749 , \12659_b0 , \12660_b0 );
not ( \12660_b0 , w_46753 );
and ( w_46753 , w_46752 , \12660_b1 );
or ( \12665_b1 , \12662_b1 , w_46756 );
or ( \12665_b0 , \12662_b0 , w_46755 );
not ( w_46755 , w_46757 );
and ( w_46757 , w_46756 , w_46754 );
or ( w_46754 , \12663_b1 , w_46758 );
or ( w_46755 , \12663_b0 , \12664_b0 );
not ( \12664_b0 , w_46759 );
and ( w_46759 , w_46758 , \12664_b1 );
or ( \12691_b1 , \12688_b1 , w_46762 );
or ( \12691_b0 , \12688_b0 , w_46761 );
not ( w_46761 , w_46763 );
and ( w_46763 , w_46762 , w_46760 );
or ( w_46760 , \12689_b1 , w_46764 );
or ( w_46761 , \12689_b0 , \12690_b0 );
not ( \12690_b0 , w_46765 );
and ( w_46765 , w_46764 , \12690_b1 );
or ( \12695_b1 , \12692_b1 , w_46768 );
or ( \12695_b0 , \12692_b0 , w_46767 );
not ( w_46767 , w_46769 );
and ( w_46769 , w_46768 , w_46766 );
or ( w_46766 , \12693_b1 , w_46770 );
or ( w_46767 , \12693_b0 , \12694_b0 );
not ( \12694_b0 , w_46771 );
and ( w_46771 , w_46770 , \12694_b1 );
or ( \12699_b1 , \12696_b1 , w_46774 );
or ( \12699_b0 , \12696_b0 , w_46773 );
not ( w_46773 , w_46775 );
and ( w_46775 , w_46774 , w_46772 );
or ( w_46772 , \12697_b1 , w_46776 );
or ( w_46773 , \12697_b0 , \12698_b0 );
not ( \12698_b0 , w_46777 );
and ( w_46777 , w_46776 , \12698_b1 );
or ( \12704_b1 , \12701_b1 , w_46780 );
or ( \12704_b0 , \12701_b0 , w_46779 );
not ( w_46779 , w_46781 );
and ( w_46781 , w_46780 , w_46778 );
or ( w_46778 , \12702_b1 , w_46782 );
or ( w_46779 , \12702_b0 , \12703_b0 );
not ( \12703_b0 , w_46783 );
and ( w_46783 , w_46782 , \12703_b1 );
or ( \12709_b1 , \12706_b1 , w_46786 );
or ( \12709_b0 , \12706_b0 , w_46785 );
not ( w_46785 , w_46787 );
and ( w_46787 , w_46786 , w_46784 );
or ( w_46784 , \12707_b1 , w_46788 );
or ( w_46785 , \12707_b0 , \12708_b0 );
not ( \12708_b0 , w_46789 );
and ( w_46789 , w_46788 , \12708_b1 );
or ( \12713_b1 , \12710_b1 , w_46792 );
or ( \12713_b0 , \12710_b0 , w_46791 );
not ( w_46791 , w_46793 );
and ( w_46793 , w_46792 , w_46790 );
or ( w_46790 , \12711_b1 , w_46794 );
or ( w_46791 , \12711_b0 , \12712_b0 );
not ( \12712_b0 , w_46795 );
and ( w_46795 , w_46794 , \12712_b1 );
or ( \12735_b1 , \12732_b1 , w_46798 );
or ( \12735_b0 , \12732_b0 , w_46797 );
not ( w_46797 , w_46799 );
and ( w_46799 , w_46798 , w_46796 );
or ( w_46796 , \12733_b1 , w_46800 );
or ( w_46797 , \12733_b0 , \12734_b0 );
not ( \12734_b0 , w_46801 );
and ( w_46801 , w_46800 , \12734_b1 );
or ( \12739_b1 , \12736_b1 , w_46804 );
or ( \12739_b0 , \12736_b0 , w_46803 );
not ( w_46803 , w_46805 );
and ( w_46805 , w_46804 , w_46802 );
or ( w_46802 , \12737_b1 , w_46806 );
or ( w_46803 , \12737_b0 , \12738_b0 );
not ( \12738_b0 , w_46807 );
and ( w_46807 , w_46806 , \12738_b1 );
or ( \12782_b1 , \12779_b1 , w_46810 );
or ( \12782_b0 , \12779_b0 , w_46809 );
not ( w_46809 , w_46811 );
and ( w_46811 , w_46810 , w_46808 );
or ( w_46808 , \12780_b1 , w_46812 );
or ( w_46809 , \12780_b0 , \12781_b0 );
not ( \12781_b0 , w_46813 );
and ( w_46813 , w_46812 , \12781_b1 );
or ( \12788_b1 , \12785_b1 , w_46816 );
or ( \12788_b0 , \12785_b0 , w_46815 );
not ( w_46815 , w_46817 );
and ( w_46817 , w_46816 , w_46814 );
or ( w_46814 , \12786_b1 , w_46818 );
or ( w_46815 , \12786_b0 , \12787_b0 );
not ( \12787_b0 , w_46819 );
and ( w_46819 , w_46818 , \12787_b1 );
or ( \12834_b1 , \12831_b1 , w_46822 );
or ( \12834_b0 , \12831_b0 , w_46821 );
not ( w_46821 , w_46823 );
and ( w_46823 , w_46822 , w_46820 );
or ( w_46820 , \12832_b1 , w_46824 );
or ( w_46821 , \12832_b0 , \12833_b0 );
not ( \12833_b0 , w_46825 );
and ( w_46825 , w_46824 , \12833_b1 );
or ( \12838_b1 , \12835_b1 , w_46828 );
or ( \12838_b0 , \12835_b0 , w_46827 );
not ( w_46827 , w_46829 );
and ( w_46829 , w_46828 , w_46826 );
or ( w_46826 , \12836_b1 , w_46830 );
or ( w_46827 , \12836_b0 , \12837_b0 );
not ( \12837_b0 , w_46831 );
and ( w_46831 , w_46830 , \12837_b1 );
or ( \12843_b1 , \12840_b1 , w_46834 );
or ( \12843_b0 , \12840_b0 , w_46833 );
not ( w_46833 , w_46835 );
and ( w_46835 , w_46834 , w_46832 );
or ( w_46832 , \12841_b1 , w_46836 );
or ( w_46833 , \12841_b0 , \12842_b0 );
not ( \12842_b0 , w_46837 );
and ( w_46837 , w_46836 , \12842_b1 );
or ( \12850_b1 , \12847_b1 , w_46840 );
or ( \12850_b0 , \12847_b0 , w_46839 );
not ( w_46839 , w_46841 );
and ( w_46841 , w_46840 , w_46838 );
or ( w_46838 , \12848_b1 , w_46842 );
or ( w_46839 , \12848_b0 , \12849_b0 );
not ( \12849_b0 , w_46843 );
and ( w_46843 , w_46842 , \12849_b1 );
or ( \12854_b1 , \12851_b1 , w_46846 );
or ( \12854_b0 , \12851_b0 , w_46845 );
not ( w_46845 , w_46847 );
and ( w_46847 , w_46846 , w_46844 );
or ( w_46844 , \12852_b1 , w_46848 );
or ( w_46845 , \12852_b0 , \12853_b0 );
not ( \12853_b0 , w_46849 );
and ( w_46849 , w_46848 , \12853_b1 );
or ( \12872_b1 , \12869_b1 , w_46852 );
or ( \12872_b0 , \12869_b0 , w_46851 );
not ( w_46851 , w_46853 );
and ( w_46853 , w_46852 , w_46850 );
or ( w_46850 , \12870_b1 , w_46854 );
or ( w_46851 , \12870_b0 , \12871_b0 );
not ( \12871_b0 , w_46855 );
and ( w_46855 , w_46854 , \12871_b1 );
or ( \12878_b1 , \12875_b1 , w_46858 );
or ( \12878_b0 , \12875_b0 , w_46857 );
not ( w_46857 , w_46859 );
and ( w_46859 , w_46858 , w_46856 );
or ( w_46856 , \12876_b1 , w_46860 );
or ( w_46857 , \12876_b0 , \12877_b0 );
not ( \12877_b0 , w_46861 );
and ( w_46861 , w_46860 , \12877_b1 );
or ( \12882_b1 , \12879_b1 , w_46864 );
or ( \12882_b0 , \12879_b0 , w_46863 );
not ( w_46863 , w_46865 );
and ( w_46865 , w_46864 , w_46862 );
or ( w_46862 , \12880_b1 , w_46866 );
or ( w_46863 , \12880_b0 , \12881_b0 );
not ( \12881_b0 , w_46867 );
and ( w_46867 , w_46866 , \12881_b1 );
or ( \12886_b1 , \12883_b1 , w_46870 );
or ( \12886_b0 , \12883_b0 , w_46869 );
not ( w_46869 , w_46871 );
and ( w_46871 , w_46870 , w_46868 );
or ( w_46868 , \12884_b1 , w_46872 );
or ( w_46869 , \12884_b0 , \12885_b0 );
not ( \12885_b0 , w_46873 );
and ( w_46873 , w_46872 , \12885_b1 );
or ( \12891_b1 , \12888_b1 , w_46876 );
or ( \12891_b0 , \12888_b0 , w_46875 );
not ( w_46875 , w_46877 );
and ( w_46877 , w_46876 , w_46874 );
or ( w_46874 , \12889_b1 , w_46878 );
or ( w_46875 , \12889_b0 , \12890_b0 );
not ( \12890_b0 , w_46879 );
and ( w_46879 , w_46878 , \12890_b1 );
or ( \12896_b1 , \12893_b1 , w_46882 );
or ( \12896_b0 , \12893_b0 , w_46881 );
not ( w_46881 , w_46883 );
and ( w_46883 , w_46882 , w_46880 );
or ( w_46880 , \12894_b1 , w_46884 );
or ( w_46881 , \12894_b0 , \12895_b0 );
not ( \12895_b0 , w_46885 );
and ( w_46885 , w_46884 , \12895_b1 );
or ( \12900_b1 , \12897_b1 , w_46888 );
or ( \12900_b0 , \12897_b0 , w_46887 );
not ( w_46887 , w_46889 );
and ( w_46889 , w_46888 , w_46886 );
or ( w_46886 , \12898_b1 , w_46890 );
or ( w_46887 , \12898_b0 , \12899_b0 );
not ( \12899_b0 , w_46891 );
and ( w_46891 , w_46890 , \12899_b1 );
or ( \12952_b1 , \12949_b1 , w_46894 );
or ( \12952_b0 , \12949_b0 , w_46893 );
not ( w_46893 , w_46895 );
and ( w_46895 , w_46894 , w_46892 );
or ( w_46892 , \12950_b1 , w_46896 );
or ( w_46893 , \12950_b0 , \12951_b0 );
not ( \12951_b0 , w_46897 );
and ( w_46897 , w_46896 , \12951_b1 );
or ( \12958_b1 , \12955_b1 , w_46900 );
or ( \12958_b0 , \12955_b0 , w_46899 );
not ( w_46899 , w_46901 );
and ( w_46901 , w_46900 , w_46898 );
or ( w_46898 , \12956_b1 , w_46902 );
or ( w_46899 , \12956_b0 , \12957_b0 );
not ( \12957_b0 , w_46903 );
and ( w_46903 , w_46902 , \12957_b1 );
or ( \12974_b1 , \12971_b1 , w_46906 );
or ( \12974_b0 , \12971_b0 , w_46905 );
not ( w_46905 , w_46907 );
and ( w_46907 , w_46906 , w_46904 );
or ( w_46904 , \12972_b1 , w_46908 );
or ( w_46905 , \12972_b0 , \12973_b0 );
not ( \12973_b0 , w_46909 );
and ( w_46909 , w_46908 , \12973_b1 );
or ( \12979_b1 , \12976_b1 , w_46912 );
or ( \12979_b0 , \12976_b0 , w_46911 );
not ( w_46911 , w_46913 );
and ( w_46913 , w_46912 , w_46910 );
or ( w_46910 , \12977_b1 , w_46914 );
or ( w_46911 , \12977_b0 , \12978_b0 );
not ( \12978_b0 , w_46915 );
and ( w_46915 , w_46914 , \12978_b1 );
or ( \12985_b1 , \12982_b1 , w_46918 );
or ( \12985_b0 , \12982_b0 , w_46917 );
not ( w_46917 , w_46919 );
and ( w_46919 , w_46918 , w_46916 );
or ( w_46916 , \12983_b1 , w_46920 );
or ( w_46917 , \12983_b0 , \12984_b0 );
not ( \12984_b0 , w_46921 );
and ( w_46921 , w_46920 , \12984_b1 );
or ( \13047_b1 , \13044_b1 , w_46924 );
or ( \13047_b0 , \13044_b0 , w_46923 );
not ( w_46923 , w_46925 );
and ( w_46925 , w_46924 , w_46922 );
or ( w_46922 , \13045_b1 , w_46926 );
or ( w_46923 , \13045_b0 , \13046_b0 );
not ( \13046_b0 , w_46927 );
and ( w_46927 , w_46926 , \13046_b1 );
or ( \13051_b1 , \13048_b1 , w_46930 );
or ( \13051_b0 , \13048_b0 , w_46929 );
not ( w_46929 , w_46931 );
and ( w_46931 , w_46930 , w_46928 );
or ( w_46928 , \13049_b1 , w_46932 );
or ( w_46929 , \13049_b0 , \13050_b0 );
not ( \13050_b0 , w_46933 );
and ( w_46933 , w_46932 , \13050_b1 );
or ( \13056_b1 , \13053_b1 , w_46936 );
or ( \13056_b0 , \13053_b0 , w_46935 );
not ( w_46935 , w_46937 );
and ( w_46937 , w_46936 , w_46934 );
or ( w_46934 , \13054_b1 , w_46938 );
or ( w_46935 , \13054_b0 , \13055_b0 );
not ( \13055_b0 , w_46939 );
and ( w_46939 , w_46938 , \13055_b1 );
or ( \13063_b1 , \13060_b1 , w_46942 );
or ( \13063_b0 , \13060_b0 , w_46941 );
not ( w_46941 , w_46943 );
and ( w_46943 , w_46942 , w_46940 );
or ( w_46940 , \13061_b1 , w_46944 );
or ( w_46941 , \13061_b0 , \13062_b0 );
not ( \13062_b0 , w_46945 );
and ( w_46945 , w_46944 , \13062_b1 );
or ( \13067_b1 , \13064_b1 , w_46948 );
or ( \13067_b0 , \13064_b0 , w_46947 );
not ( w_46947 , w_46949 );
and ( w_46949 , w_46948 , w_46946 );
or ( w_46946 , \13065_b1 , w_46950 );
or ( w_46947 , \13065_b0 , \13066_b0 );
not ( \13066_b0 , w_46951 );
and ( w_46951 , w_46950 , \13066_b1 );
or ( \13072_b1 , \13069_b1 , w_46954 );
or ( \13072_b0 , \13069_b0 , w_46953 );
not ( w_46953 , w_46955 );
and ( w_46955 , w_46954 , w_46952 );
or ( w_46952 , \13070_b1 , w_46956 );
or ( w_46953 , \13070_b0 , \13071_b0 );
not ( \13071_b0 , w_46957 );
and ( w_46957 , w_46956 , \13071_b1 );
or ( \13079_b1 , \13076_b1 , w_46960 );
or ( \13079_b0 , \13076_b0 , w_46959 );
not ( w_46959 , w_46961 );
and ( w_46961 , w_46960 , w_46958 );
or ( w_46958 , \13077_b1 , w_46962 );
or ( w_46959 , \13077_b0 , \13078_b0 );
not ( \13078_b0 , w_46963 );
and ( w_46963 , w_46962 , \13078_b1 );
or ( \13087_b1 , \13084_b1 , w_46966 );
or ( \13087_b0 , \13084_b0 , w_46965 );
not ( w_46965 , w_46967 );
and ( w_46967 , w_46966 , w_46964 );
or ( w_46964 , \13085_b1 , w_46968 );
or ( w_46965 , \13085_b0 , \13086_b0 );
not ( \13086_b0 , w_46969 );
and ( w_46969 , w_46968 , \13086_b1 );
or ( \13091_b1 , \13088_b1 , w_46972 );
or ( \13091_b0 , \13088_b0 , w_46971 );
not ( w_46971 , w_46973 );
and ( w_46973 , w_46972 , w_46970 );
or ( w_46970 , \13089_b1 , w_46974 );
or ( w_46971 , \13089_b0 , \13090_b0 );
not ( \13090_b0 , w_46975 );
and ( w_46975 , w_46974 , \13090_b1 );
or ( \13095_b1 , \13092_b1 , w_46978 );
or ( \13095_b0 , \13092_b0 , w_46977 );
not ( w_46977 , w_46979 );
and ( w_46979 , w_46978 , w_46976 );
or ( w_46976 , \13093_b1 , w_46980 );
or ( w_46977 , \13093_b0 , \13094_b0 );
not ( \13094_b0 , w_46981 );
and ( w_46981 , w_46980 , \13094_b1 );
or ( \13103_b1 , \13100_b1 , w_46984 );
or ( \13103_b0 , \13100_b0 , w_46983 );
not ( w_46983 , w_46985 );
and ( w_46985 , w_46984 , w_46982 );
or ( w_46982 , \13101_b1 , w_46986 );
or ( w_46983 , \13101_b0 , \13102_b0 );
not ( \13102_b0 , w_46987 );
and ( w_46987 , w_46986 , \13102_b1 );
or ( \13107_b1 , \13104_b1 , w_46990 );
or ( \13107_b0 , \13104_b0 , w_46989 );
not ( w_46989 , w_46991 );
and ( w_46991 , w_46990 , w_46988 );
or ( w_46988 , \13105_b1 , w_46992 );
or ( w_46989 , \13105_b0 , \13106_b0 );
not ( \13106_b0 , w_46993 );
and ( w_46993 , w_46992 , \13106_b1 );
or ( \13141_b1 , \13138_b1 , w_46996 );
or ( \13141_b0 , \13138_b0 , w_46995 );
not ( w_46995 , w_46997 );
and ( w_46997 , w_46996 , w_46994 );
or ( w_46994 , \13139_b1 , w_46998 );
or ( w_46995 , \13139_b0 , \13140_b0 );
not ( \13140_b0 , w_46999 );
and ( w_46999 , w_46998 , \13140_b1 );
or ( \13176_b1 , \13173_b1 , w_47002 );
or ( \13176_b0 , \13173_b0 , w_47001 );
not ( w_47001 , w_47003 );
and ( w_47003 , w_47002 , w_47000 );
or ( w_47000 , \13174_b1 , w_47004 );
or ( w_47001 , \13174_b0 , \13175_b0 );
not ( \13175_b0 , w_47005 );
and ( w_47005 , w_47004 , \13175_b1 );
or ( \13180_b1 , \13177_b1 , w_47008 );
or ( \13180_b0 , \13177_b0 , w_47007 );
not ( w_47007 , w_47009 );
and ( w_47009 , w_47008 , w_47006 );
or ( w_47006 , \13178_b1 , w_47010 );
or ( w_47007 , \13178_b0 , \13179_b0 );
not ( \13179_b0 , w_47011 );
and ( w_47011 , w_47010 , \13179_b1 );
or ( \13185_b1 , \13182_b1 , w_47014 );
or ( \13185_b0 , \13182_b0 , w_47013 );
not ( w_47013 , w_47015 );
and ( w_47015 , w_47014 , w_47012 );
or ( w_47012 , \13183_b1 , w_47016 );
or ( w_47013 , \13183_b0 , \13184_b0 );
not ( \13184_b0 , w_47017 );
and ( w_47017 , w_47016 , \13184_b1 );
or ( \13193_b1 , \13190_b1 , w_47020 );
or ( \13193_b0 , \13190_b0 , w_47019 );
not ( w_47019 , w_47021 );
and ( w_47021 , w_47020 , w_47018 );
or ( w_47018 , \13191_b1 , w_47022 );
or ( w_47019 , \13191_b0 , \13192_b0 );
not ( \13192_b0 , w_47023 );
and ( w_47023 , w_47022 , \13192_b1 );
or ( \13198_b1 , \13195_b1 , w_47026 );
or ( \13198_b0 , \13195_b0 , w_47025 );
not ( w_47025 , w_47027 );
and ( w_47027 , w_47026 , w_47024 );
or ( w_47024 , \13196_b1 , w_47028 );
or ( w_47025 , \13196_b0 , \13197_b0 );
not ( \13197_b0 , w_47029 );
and ( w_47029 , w_47028 , \13197_b1 );
or ( \13202_b1 , \13199_b1 , w_47032 );
or ( \13202_b0 , \13199_b0 , w_47031 );
not ( w_47031 , w_47033 );
and ( w_47033 , w_47032 , w_47030 );
or ( w_47030 , \13200_b1 , w_47034 );
or ( w_47031 , \13200_b0 , \13201_b0 );
not ( \13201_b0 , w_47035 );
and ( w_47035 , w_47034 , \13201_b1 );
or ( \13206_b1 , \13203_b1 , w_47038 );
or ( \13206_b0 , \13203_b0 , w_47037 );
not ( w_47037 , w_47039 );
and ( w_47039 , w_47038 , w_47036 );
or ( w_47036 , \13204_b1 , w_47040 );
or ( w_47037 , \13204_b0 , \13205_b0 );
not ( \13205_b0 , w_47041 );
and ( w_47041 , w_47040 , \13205_b1 );
or ( \13214_b1 , \13211_b1 , w_47044 );
or ( \13214_b0 , \13211_b0 , w_47043 );
not ( w_47043 , w_47045 );
and ( w_47045 , w_47044 , w_47042 );
or ( w_47042 , \13212_b1 , w_47046 );
or ( w_47043 , \13212_b0 , \13213_b0 );
not ( \13213_b0 , w_47047 );
and ( w_47047 , w_47046 , \13213_b1 );
or ( \13218_b1 , \13215_b1 , w_47050 );
or ( \13218_b0 , \13215_b0 , w_47049 );
not ( w_47049 , w_47051 );
and ( w_47051 , w_47050 , w_47048 );
or ( w_47048 , \13216_b1 , w_47052 );
or ( w_47049 , \13216_b0 , \13217_b0 );
not ( \13217_b0 , w_47053 );
and ( w_47053 , w_47052 , \13217_b1 );
or ( \13263_b1 , \13260_b1 , w_47056 );
or ( \13263_b0 , \13260_b0 , w_47055 );
not ( w_47055 , w_47057 );
and ( w_47057 , w_47056 , w_47054 );
or ( w_47054 , \13261_b1 , w_47058 );
or ( w_47055 , \13261_b0 , \13262_b0 );
not ( \13262_b0 , w_47059 );
and ( w_47059 , w_47058 , \13262_b1 );
or ( \13291_b1 , \13288_b1 , w_47062 );
or ( \13291_b0 , \13288_b0 , w_47061 );
not ( w_47061 , w_47063 );
and ( w_47063 , w_47062 , w_47060 );
or ( w_47060 , \13289_b1 , w_47064 );
or ( w_47061 , \13289_b0 , \13290_b0 );
not ( \13290_b0 , w_47065 );
and ( w_47065 , w_47064 , \13290_b1 );
or ( \13295_b1 , \13292_b1 , w_47068 );
or ( \13295_b0 , \13292_b0 , w_47067 );
not ( w_47067 , w_47069 );
and ( w_47069 , w_47068 , w_47066 );
or ( w_47066 , \13293_b1 , w_47070 );
or ( w_47067 , \13293_b0 , \13294_b0 );
not ( \13294_b0 , w_47071 );
and ( w_47071 , w_47070 , \13294_b1 );
or ( \13300_b1 , \13297_b1 , w_47074 );
or ( \13300_b0 , \13297_b0 , w_47073 );
not ( w_47073 , w_47075 );
and ( w_47075 , w_47074 , w_47072 );
or ( w_47072 , \13298_b1 , w_47076 );
or ( w_47073 , \13298_b0 , \13299_b0 );
not ( \13299_b0 , w_47077 );
and ( w_47077 , w_47076 , \13299_b1 );
or ( \13308_b1 , \13305_b1 , w_47080 );
or ( \13308_b0 , \13305_b0 , w_47079 );
not ( w_47079 , w_47081 );
and ( w_47081 , w_47080 , w_47078 );
or ( w_47078 , \13306_b1 , w_47082 );
or ( w_47079 , \13306_b0 , \13307_b0 );
not ( \13307_b0 , w_47083 );
and ( w_47083 , w_47082 , \13307_b1 );
or ( \13314_b1 , \13311_b1 , w_47086 );
or ( \13314_b0 , \13311_b0 , w_47085 );
not ( w_47085 , w_47087 );
and ( w_47087 , w_47086 , w_47084 );
or ( w_47084 , \13312_b1 , w_47088 );
or ( w_47085 , \13312_b0 , \13313_b0 );
not ( \13313_b0 , w_47089 );
and ( w_47089 , w_47088 , \13313_b1 );
or ( \13329_b1 , \13326_b1 , w_47092 );
or ( \13329_b0 , \13326_b0 , w_47091 );
not ( w_47091 , w_47093 );
and ( w_47093 , w_47092 , w_47090 );
or ( w_47090 , \13327_b1 , w_47094 );
or ( w_47091 , \13327_b0 , \13328_b0 );
not ( \13328_b0 , w_47095 );
and ( w_47095 , w_47094 , \13328_b1 );
or ( \13341_b1 , \13338_b1 , w_47098 );
or ( \13341_b0 , \13338_b0 , w_47097 );
not ( w_47097 , w_47099 );
and ( w_47099 , w_47098 , w_47096 );
or ( w_47096 , \13339_b1 , w_47100 );
or ( w_47097 , \13339_b0 , \13340_b0 );
not ( \13340_b0 , w_47101 );
and ( w_47101 , w_47100 , \13340_b1 );
or ( \13345_b1 , \13342_b1 , w_47104 );
or ( \13345_b0 , \13342_b0 , w_47103 );
not ( w_47103 , w_47105 );
and ( w_47105 , w_47104 , w_47102 );
or ( w_47102 , \13343_b1 , w_47106 );
or ( w_47103 , \13343_b0 , \13344_b0 );
not ( \13344_b0 , w_47107 );
and ( w_47107 , w_47106 , \13344_b1 );
or ( \13350_b1 , \13347_b1 , w_47110 );
or ( \13350_b0 , \13347_b0 , w_47109 );
not ( w_47109 , w_47111 );
and ( w_47111 , w_47110 , w_47108 );
or ( w_47108 , \13348_b1 , w_47112 );
or ( w_47109 , \13348_b0 , \13349_b0 );
not ( \13349_b0 , w_47113 );
and ( w_47113 , w_47112 , \13349_b1 );
or ( \13357_b1 , \13354_b1 , w_47116 );
or ( \13357_b0 , \13354_b0 , w_47115 );
not ( w_47115 , w_47117 );
and ( w_47117 , w_47116 , w_47114 );
or ( w_47114 , \13355_b1 , w_47118 );
or ( w_47115 , \13355_b0 , \13356_b0 );
not ( \13356_b0 , w_47119 );
and ( w_47119 , w_47118 , \13356_b1 );
or ( \13361_b1 , \13358_b1 , w_47122 );
or ( \13361_b0 , \13358_b0 , w_47121 );
not ( w_47121 , w_47123 );
and ( w_47123 , w_47122 , w_47120 );
or ( w_47120 , \13359_b1 , w_47124 );
or ( w_47121 , \13359_b0 , \13360_b0 );
not ( \13360_b0 , w_47125 );
and ( w_47125 , w_47124 , \13360_b1 );
or ( \13366_b1 , \13363_b1 , w_47128 );
or ( \13366_b0 , \13363_b0 , w_47127 );
not ( w_47127 , w_47129 );
and ( w_47129 , w_47128 , w_47126 );
or ( w_47126 , \13364_b1 , w_47130 );
or ( w_47127 , \13364_b0 , \13365_b0 );
not ( \13365_b0 , w_47131 );
and ( w_47131 , w_47130 , \13365_b1 );
or ( \13370_b1 , \13367_b1 , w_47134 );
or ( \13370_b0 , \13367_b0 , w_47133 );
not ( w_47133 , w_47135 );
and ( w_47135 , w_47134 , w_47132 );
or ( w_47132 , \13368_b1 , w_47136 );
or ( w_47133 , \13368_b0 , \13369_b0 );
not ( \13369_b0 , w_47137 );
and ( w_47137 , w_47136 , \13369_b1 );
or ( \13375_b1 , \13372_b1 , w_47140 );
or ( \13375_b0 , \13372_b0 , w_47139 );
not ( w_47139 , w_47141 );
and ( w_47141 , w_47140 , w_47138 );
or ( w_47138 , \13373_b1 , w_47142 );
or ( w_47139 , \13373_b0 , \13374_b0 );
not ( \13374_b0 , w_47143 );
and ( w_47143 , w_47142 , \13374_b1 );
or ( \13382_b1 , \13379_b1 , w_47146 );
or ( \13382_b0 , \13379_b0 , w_47145 );
not ( w_47145 , w_47147 );
and ( w_47147 , w_47146 , w_47144 );
or ( w_47144 , \13380_b1 , w_47148 );
or ( w_47145 , \13380_b0 , \13381_b0 );
not ( \13381_b0 , w_47149 );
and ( w_47149 , w_47148 , \13381_b1 );
or ( \13387_b1 , \13384_b1 , w_47152 );
or ( \13387_b0 , \13384_b0 , w_47151 );
not ( w_47151 , w_47153 );
and ( w_47153 , w_47152 , w_47150 );
or ( w_47150 , \13385_b1 , w_47154 );
or ( w_47151 , \13385_b0 , \13386_b0 );
not ( \13386_b0 , w_47155 );
and ( w_47155 , w_47154 , \13386_b1 );
or ( \13391_b1 , \13388_b1 , w_47158 );
or ( \13391_b0 , \13388_b0 , w_47157 );
not ( w_47157 , w_47159 );
and ( w_47159 , w_47158 , w_47156 );
or ( w_47156 , \13389_b1 , w_47160 );
or ( w_47157 , \13389_b0 , \13390_b0 );
not ( \13390_b0 , w_47161 );
and ( w_47161 , w_47160 , \13390_b1 );
or ( \13405_b1 , \13402_b1 , w_47164 );
or ( \13405_b0 , \13402_b0 , w_47163 );
not ( w_47163 , w_47165 );
and ( w_47165 , w_47164 , w_47162 );
or ( w_47162 , \13403_b1 , w_47166 );
or ( w_47163 , \13403_b0 , \13404_b0 );
not ( \13404_b0 , w_47167 );
and ( w_47167 , w_47166 , \13404_b1 );
or ( \13411_b1 , \13408_b1 , w_47170 );
or ( \13411_b0 , \13408_b0 , w_47169 );
not ( w_47169 , w_47171 );
and ( w_47171 , w_47170 , w_47168 );
or ( w_47168 , \13409_b1 , w_47172 );
or ( w_47169 , \13409_b0 , \13410_b0 );
not ( \13410_b0 , w_47173 );
and ( w_47173 , w_47172 , \13410_b1 );
or ( \13415_b1 , \13412_b1 , w_47176 );
or ( \13415_b0 , \13412_b0 , w_47175 );
not ( w_47175 , w_47177 );
and ( w_47177 , w_47176 , w_47174 );
or ( w_47174 , \13413_b1 , w_47178 );
or ( w_47175 , \13413_b0 , \13414_b0 );
not ( \13414_b0 , w_47179 );
and ( w_47179 , w_47178 , \13414_b1 );
or ( \13420_b1 , \13417_b1 , w_47182 );
or ( \13420_b0 , \13417_b0 , w_47181 );
not ( w_47181 , w_47183 );
and ( w_47183 , w_47182 , w_47180 );
or ( w_47180 , \13418_b1 , w_47184 );
or ( w_47181 , \13418_b0 , \13419_b0 );
not ( \13419_b0 , w_47185 );
and ( w_47185 , w_47184 , \13419_b1 );
or ( \13427_b1 , \13424_b1 , w_47188 );
or ( \13427_b0 , \13424_b0 , w_47187 );
not ( w_47187 , w_47189 );
and ( w_47189 , w_47188 , w_47186 );
or ( w_47186 , \13425_b1 , w_47190 );
or ( w_47187 , \13425_b0 , \13426_b0 );
not ( \13426_b0 , w_47191 );
and ( w_47191 , w_47190 , \13426_b1 );
or ( \13434_b1 , \13431_b1 , w_47194 );
or ( \13434_b0 , \13431_b0 , w_47193 );
not ( w_47193 , w_47195 );
and ( w_47195 , w_47194 , w_47192 );
or ( w_47192 , \13432_b1 , w_47196 );
or ( w_47193 , \13432_b0 , \13433_b0 );
not ( \13433_b0 , w_47197 );
and ( w_47197 , w_47196 , \13433_b1 );
or ( \13438_b1 , \13435_b1 , w_47200 );
or ( \13438_b0 , \13435_b0 , w_47199 );
not ( w_47199 , w_47201 );
and ( w_47201 , w_47200 , w_47198 );
or ( w_47198 , \13436_b1 , w_47202 );
or ( w_47199 , \13436_b0 , \13437_b0 );
not ( \13437_b0 , w_47203 );
and ( w_47203 , w_47202 , \13437_b1 );
or ( \13451_b1 , \13448_b1 , w_47206 );
or ( \13451_b0 , \13448_b0 , w_47205 );
not ( w_47205 , w_47207 );
and ( w_47207 , w_47206 , w_47204 );
or ( w_47204 , \13449_b1 , w_47208 );
or ( w_47205 , \13449_b0 , \13450_b0 );
not ( \13450_b0 , w_47209 );
and ( w_47209 , w_47208 , \13450_b1 );
or ( \13455_b1 , \13452_b1 , w_47212 );
or ( \13455_b0 , \13452_b0 , w_47211 );
not ( w_47211 , w_47213 );
and ( w_47213 , w_47212 , w_47210 );
or ( w_47210 , \13453_b1 , w_47214 );
or ( w_47211 , \13453_b0 , \13454_b0 );
not ( \13454_b0 , w_47215 );
and ( w_47215 , w_47214 , \13454_b1 );
or ( \13467_b1 , \13464_b1 , w_47218 );
or ( \13467_b0 , \13464_b0 , w_47217 );
not ( w_47217 , w_47219 );
and ( w_47219 , w_47218 , w_47216 );
or ( w_47216 , \13465_b1 , w_47220 );
or ( w_47217 , \13465_b0 , \13466_b0 );
not ( \13466_b0 , w_47221 );
and ( w_47221 , w_47220 , \13466_b1 );
or ( \13477_b1 , \13474_b1 , w_47224 );
or ( \13477_b0 , \13474_b0 , w_47223 );
not ( w_47223 , w_47225 );
and ( w_47225 , w_47224 , w_47222 );
or ( w_47222 , \13475_b1 , w_47226 );
or ( w_47223 , \13475_b0 , \13476_b0 );
not ( \13476_b0 , w_47227 );
and ( w_47227 , w_47226 , \13476_b1 );
or ( \13481_b1 , \13478_b1 , w_47230 );
or ( \13481_b0 , \13478_b0 , w_47229 );
not ( w_47229 , w_47231 );
and ( w_47231 , w_47230 , w_47228 );
or ( w_47228 , \13479_b1 , w_47232 );
or ( w_47229 , \13479_b0 , \13480_b0 );
not ( \13480_b0 , w_47233 );
and ( w_47233 , w_47232 , \13480_b1 );
or ( \13493_b1 , \13490_b1 , w_47236 );
or ( \13493_b0 , \13490_b0 , w_47235 );
not ( w_47235 , w_47237 );
and ( w_47237 , w_47236 , w_47234 );
or ( w_47234 , \13491_b1 , w_47238 );
or ( w_47235 , \13491_b0 , \13492_b0 );
not ( \13492_b0 , w_47239 );
and ( w_47239 , w_47238 , \13492_b1 );
or ( \13502_b1 , \13499_b1 , w_47242 );
or ( \13502_b0 , \13499_b0 , w_47241 );
not ( w_47241 , w_47243 );
and ( w_47243 , w_47242 , w_47240 );
or ( w_47240 , \13500_b1 , w_47244 );
or ( w_47241 , \13500_b0 , \13501_b0 );
not ( \13501_b0 , w_47245 );
and ( w_47245 , w_47244 , \13501_b1 );
or ( \13509_b1 , \13506_b1 , w_47248 );
or ( \13509_b0 , \13506_b0 , w_47247 );
not ( w_47247 , w_47249 );
and ( w_47249 , w_47248 , w_47246 );
or ( w_47246 , \13507_b1 , w_47250 );
or ( w_47247 , \13507_b0 , \13508_b0 );
not ( \13508_b0 , w_47251 );
and ( w_47251 , w_47250 , \13508_b1 );
or ( \13540_b1 , \13533_b1 , w_47254 );
or ( \13540_b0 , \13533_b0 , w_47253 );
not ( w_47253 , w_47255 );
and ( w_47255 , w_47254 , w_47252 );
or ( w_47252 , \13538_b1 , w_47256 );
or ( w_47253 , \13538_b0 , \13539_b0 );
not ( \13539_b0 , w_47257 );
and ( w_47257 , w_47256 , \13539_b1 );
or ( \13570_b1 , \13563_b1 , w_47260 );
or ( \13570_b0 , \13563_b0 , w_47259 );
not ( w_47259 , w_47261 );
and ( w_47261 , w_47260 , w_47258 );
or ( w_47258 , \13568_b1 , w_47262 );
or ( w_47259 , \13568_b0 , \13569_b0 );
not ( \13569_b0 , w_47263 );
and ( w_47263 , w_47262 , \13569_b1 );
or ( \13577_b1 , \13572_b1 , w_47266 );
or ( \13577_b0 , \13572_b0 , w_47265 );
not ( w_47265 , w_47267 );
and ( w_47267 , w_47266 , w_47264 );
or ( w_47264 , \13575_b1 , w_47268 );
or ( w_47265 , \13575_b0 , \13576_b0 );
not ( \13576_b0 , w_47269 );
and ( w_47269 , w_47268 , \13576_b1 );
or ( \13582_b1 , \13579_b1 , w_47272 );
or ( \13582_b0 , \13579_b0 , w_47271 );
not ( w_47271 , w_47273 );
and ( w_47273 , w_47272 , w_47270 );
or ( w_47270 , \13580_b1 , w_47274 );
or ( w_47271 , \13580_b0 , \13581_b0 );
not ( \13581_b0 , w_47275 );
and ( w_47275 , w_47274 , \13581_b1 );
or ( \13586_b1 , \13583_b1 , w_47278 );
or ( \13586_b0 , \13583_b0 , w_47277 );
not ( w_47277 , w_47279 );
and ( w_47279 , w_47278 , w_47276 );
or ( w_47276 , \13584_b1 , w_47280 );
or ( w_47277 , \13584_b0 , \13585_b0 );
not ( \13585_b0 , w_47281 );
and ( w_47281 , w_47280 , \13585_b1 );
or ( \13618_b1 , \13615_b1 , w_47284 );
or ( \13618_b0 , \13615_b0 , w_47283 );
not ( w_47283 , w_47285 );
and ( w_47285 , w_47284 , w_47282 );
or ( w_47282 , \13616_b1 , w_47286 );
or ( w_47283 , \13616_b0 , \13617_b0 );
not ( \13617_b0 , w_47287 );
and ( w_47287 , w_47286 , \13617_b1 );
or ( \13642_b1 , \13639_b1 , w_47290 );
or ( \13642_b0 , \13639_b0 , w_47289 );
not ( w_47289 , w_47291 );
and ( w_47291 , w_47290 , w_47288 );
or ( w_47288 , \13640_b1 , w_47292 );
or ( w_47289 , \13640_b0 , \13641_b0 );
not ( \13641_b0 , w_47293 );
and ( w_47293 , w_47292 , \13641_b1 );
or ( \13646_b1 , \13643_b1 , w_47296 );
or ( \13646_b0 , \13643_b0 , w_47295 );
not ( w_47295 , w_47297 );
and ( w_47297 , w_47296 , w_47294 );
or ( w_47294 , \13644_b1 , w_47298 );
or ( w_47295 , \13644_b0 , \13645_b0 );
not ( \13645_b0 , w_47299 );
and ( w_47299 , w_47298 , \13645_b1 );
or ( \13659_b1 , \13656_b1 , w_47302 );
or ( \13659_b0 , \13656_b0 , w_47301 );
not ( w_47301 , w_47303 );
and ( w_47303 , w_47302 , w_47300 );
or ( w_47300 , \13657_b1 , w_47304 );
or ( w_47301 , \13657_b0 , \13658_b0 );
not ( \13658_b0 , w_47305 );
and ( w_47305 , w_47304 , \13658_b1 );
or ( \13681_b1 , \13678_b1 , w_47308 );
or ( \13681_b0 , \13678_b0 , w_47307 );
not ( w_47307 , w_47309 );
and ( w_47309 , w_47308 , w_47306 );
or ( w_47306 , \13679_b1 , w_47310 );
or ( w_47307 , \13679_b0 , \13680_b0 );
not ( \13680_b0 , w_47311 );
and ( w_47311 , w_47310 , \13680_b1 );
or ( \13699_b1 , \13696_b1 , w_47314 );
or ( \13699_b0 , \13696_b0 , w_47313 );
not ( w_47313 , w_47315 );
and ( w_47315 , w_47314 , w_47312 );
or ( w_47312 , \13697_b1 , w_47316 );
or ( w_47313 , \13697_b0 , \13698_b0 );
not ( \13698_b0 , w_47317 );
and ( w_47317 , w_47316 , \13698_b1 );
or ( \13706_b1 , \13703_b1 , w_47320 );
or ( \13706_b0 , \13703_b0 , w_47319 );
not ( w_47319 , w_47321 );
and ( w_47321 , w_47320 , w_47318 );
or ( w_47318 , \13704_b1 , w_47322 );
or ( w_47319 , \13704_b0 , \13705_b0 );
not ( \13705_b0 , w_47323 );
and ( w_47323 , w_47322 , \13705_b1 );
or ( \13710_b1 , \13707_b1 , w_47326 );
or ( \13710_b0 , \13707_b0 , w_47325 );
not ( w_47325 , w_47327 );
and ( w_47327 , w_47326 , w_47324 );
or ( w_47324 , \13708_b1 , w_47328 );
or ( w_47325 , \13708_b0 , \13709_b0 );
not ( \13709_b0 , w_47329 );
and ( w_47329 , w_47328 , \13709_b1 );
or ( \13717_b1 , \13714_b1 , w_47332 );
or ( \13717_b0 , \13714_b0 , w_47331 );
not ( w_47331 , w_47333 );
and ( w_47333 , w_47332 , w_47330 );
or ( w_47330 , \13715_b1 , w_47334 );
or ( w_47331 , \13715_b0 , \13716_b0 );
not ( \13716_b0 , w_47335 );
and ( w_47335 , w_47334 , \13716_b1 );
or ( \13721_b1 , \13718_b1 , w_47338 );
or ( \13721_b0 , \13718_b0 , w_47337 );
not ( w_47337 , w_47339 );
and ( w_47339 , w_47338 , w_47336 );
or ( w_47336 , \13719_b1 , w_47340 );
or ( w_47337 , \13719_b0 , \13720_b0 );
not ( \13720_b0 , w_47341 );
and ( w_47341 , w_47340 , \13720_b1 );
or ( \13733_b1 , \13730_b1 , w_47344 );
or ( \13733_b0 , \13730_b0 , w_47343 );
not ( w_47343 , w_47345 );
and ( w_47345 , w_47344 , w_47342 );
or ( w_47342 , \13731_b1 , w_47346 );
or ( w_47343 , \13731_b0 , \13732_b0 );
not ( \13732_b0 , w_47347 );
and ( w_47347 , w_47346 , \13732_b1 );
or ( \13737_b1 , \13734_b1 , w_47350 );
or ( \13737_b0 , \13734_b0 , w_47349 );
not ( w_47349 , w_47351 );
and ( w_47351 , w_47350 , w_47348 );
or ( w_47348 , \13735_b1 , w_47352 );
or ( w_47349 , \13735_b0 , \13736_b0 );
not ( \13736_b0 , w_47353 );
and ( w_47353 , w_47352 , \13736_b1 );
or ( \13751_b1 , \13748_b1 , w_47356 );
or ( \13751_b0 , \13748_b0 , w_47355 );
not ( w_47355 , w_47357 );
and ( w_47357 , w_47356 , w_47354 );
or ( w_47354 , \13749_b1 , w_47358 );
or ( w_47355 , \13749_b0 , \13750_b0 );
not ( \13750_b0 , w_47359 );
and ( w_47359 , w_47358 , \13750_b1 );
or ( \13764_b1 , \13761_b1 , w_47362 );
or ( \13764_b0 , \13761_b0 , w_47361 );
not ( w_47361 , w_47363 );
and ( w_47363 , w_47362 , w_47360 );
or ( w_47360 , \13762_b1 , w_47364 );
or ( w_47361 , \13762_b0 , \13763_b0 );
not ( \13763_b0 , w_47365 );
and ( w_47365 , w_47364 , \13763_b1 );
or ( \13803_b1 , \13800_b1 , w_47368 );
or ( \13803_b0 , \13800_b0 , w_47367 );
not ( w_47367 , w_47369 );
and ( w_47369 , w_47368 , w_47366 );
or ( w_47366 , \13801_b1 , w_47370 );
or ( w_47367 , \13801_b0 , \13802_b0 );
not ( \13802_b0 , w_47371 );
and ( w_47371 , w_47370 , \13802_b1 );
endmodule

