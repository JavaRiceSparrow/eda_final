// ...
module top(\A[0][9]_b1 ,\A[0][9]_b0 ,\A[0][8]_b1 ,\A[0][8]_b0 ,\A[0][7]_b1 ,\A[0][7]_b0 ,\A[0][6]_b1 ,\A[0][6]_b0 ,\A[0][5]_b1 ,
		\A[0][5]_b0 ,\A[0][4]_b1 ,\A[0][4]_b0 ,\A[0][3]_b1 ,\A[0][3]_b0 ,\A[0][2]_b1 ,\A[0][2]_b0 ,\A[0][1]_b1 ,\A[0][1]_b0 ,
		\A[0][0]_b1 ,\A[0][0]_b0 ,\A[1][9]_b1 ,\A[1][9]_b0 ,\A[1][8]_b1 ,\A[1][8]_b0 ,\A[1][7]_b1 ,\A[1][7]_b0 ,\A[1][6]_b1 ,
		\A[1][6]_b0 ,\A[1][5]_b1 ,\A[1][5]_b0 ,\A[1][4]_b1 ,\A[1][4]_b0 ,\A[1][3]_b1 ,\A[1][3]_b0 ,\A[1][2]_b1 ,\A[1][2]_b0 ,
		\A[1][1]_b1 ,\A[1][1]_b0 ,\A[1][0]_b1 ,\A[1][0]_b0 ,\A[2][9]_b1 ,\A[2][9]_b0 ,\A[2][8]_b1 ,\A[2][8]_b0 ,\A[2][7]_b1 ,
		\A[2][7]_b0 ,\A[2][6]_b1 ,\A[2][6]_b0 ,\A[2][5]_b1 ,\A[2][5]_b0 ,\A[2][4]_b1 ,\A[2][4]_b0 ,\A[2][3]_b1 ,\A[2][3]_b0 ,
		\A[2][2]_b1 ,\A[2][2]_b0 ,\A[2][1]_b1 ,\A[2][1]_b0 ,\A[2][0]_b1 ,\A[2][0]_b0 ,\B[9]_b1 ,\B[9]_b0 ,\B[8]_b1 ,
		\B[8]_b0 ,\B[7]_b1 ,\B[7]_b0 ,\B[6]_b1 ,\B[6]_b0 ,\B[5]_b1 ,\B[5]_b0 ,\B[4]_b1 ,\B[4]_b0 ,
		\B[3]_b1 ,\B[3]_b0 ,\B[2]_b1 ,\B[2]_b0 ,\B[1]_b1 ,\B[1]_b0 ,\B[0]_b1 ,\B[0]_b0 ,\I[7]_b1 ,
		\I[7]_b0 ,\I[6]_b1 ,\I[6]_b0 ,\I[5]_b1 ,\I[5]_b0 ,\I[4]_b1 ,\I[4]_b0 ,\I[3]_b1 ,\I[3]_b0 ,
		\I[2]_b1 ,\I[2]_b0 ,\I[1]_b1 ,\I[1]_b0 ,\I[0]_b1 ,\I[0]_b0 ,\O[19]_b1 ,\O[19]_b0 ,\O[18]_b1 ,
		\O[18]_b0 ,\O[17]_b1 ,\O[17]_b0 ,\O[16]_b1 ,\O[16]_b0 ,\O[15]_b1 ,\O[15]_b0 ,\O[14]_b1 ,\O[14]_b0 ,
		\O[13]_b1 ,\O[13]_b0 ,\O[12]_b1 ,\O[12]_b0 ,\O[11]_b1 ,\O[11]_b0 ,\O[10]_b1 ,\O[10]_b0 ,\O[9]_b1 ,
		\O[9]_b0 ,\O[8]_b1 ,\O[8]_b0 ,\O[7]_b1 ,\O[7]_b0 ,\O[6]_b1 ,\O[6]_b0 ,\O[5]_b1 ,\O[5]_b0 ,
		\O[4]_b1 ,\O[4]_b0 ,\O[3]_b1 ,\O[3]_b0 ,\O[2]_b1 ,\O[2]_b0 ,\O[1]_b1 ,\O[1]_b0 ,\O[0]_b1 ,
		\O[0]_b0 );
input \A[0][9]_b1 ,\A[0][9]_b0 ,\A[0][8]_b1 ,\A[0][8]_b0 ,\A[0][7]_b1 ,\A[0][7]_b0 ,\A[0][6]_b1 ,\A[0][6]_b0 ,\A[0][5]_b1 ,
		\A[0][5]_b0 ,\A[0][4]_b1 ,\A[0][4]_b0 ,\A[0][3]_b1 ,\A[0][3]_b0 ,\A[0][2]_b1 ,\A[0][2]_b0 ,\A[0][1]_b1 ,\A[0][1]_b0 ,
		\A[0][0]_b1 ,\A[0][0]_b0 ,\A[1][9]_b1 ,\A[1][9]_b0 ,\A[1][8]_b1 ,\A[1][8]_b0 ,\A[1][7]_b1 ,\A[1][7]_b0 ,\A[1][6]_b1 ,
		\A[1][6]_b0 ,\A[1][5]_b1 ,\A[1][5]_b0 ,\A[1][4]_b1 ,\A[1][4]_b0 ,\A[1][3]_b1 ,\A[1][3]_b0 ,\A[1][2]_b1 ,\A[1][2]_b0 ,
		\A[1][1]_b1 ,\A[1][1]_b0 ,\A[1][0]_b1 ,\A[1][0]_b0 ,\A[2][9]_b1 ,\A[2][9]_b0 ,\A[2][8]_b1 ,\A[2][8]_b0 ,\A[2][7]_b1 ,
		\A[2][7]_b0 ,\A[2][6]_b1 ,\A[2][6]_b0 ,\A[2][5]_b1 ,\A[2][5]_b0 ,\A[2][4]_b1 ,\A[2][4]_b0 ,\A[2][3]_b1 ,\A[2][3]_b0 ,
		\A[2][2]_b1 ,\A[2][2]_b0 ,\A[2][1]_b1 ,\A[2][1]_b0 ,\A[2][0]_b1 ,\A[2][0]_b0 ,\B[9]_b1 ,\B[9]_b0 ,\B[8]_b1 ,
		\B[8]_b0 ,\B[7]_b1 ,\B[7]_b0 ,\B[6]_b1 ,\B[6]_b0 ,\B[5]_b1 ,\B[5]_b0 ,\B[4]_b1 ,\B[4]_b0 ,
		\B[3]_b1 ,\B[3]_b0 ,\B[2]_b1 ,\B[2]_b0 ,\B[1]_b1 ,\B[1]_b0 ,\B[0]_b1 ,\B[0]_b0 ,\I[7]_b1 ,
		\I[7]_b0 ,\I[6]_b1 ,\I[6]_b0 ,\I[5]_b1 ,\I[5]_b0 ,\I[4]_b1 ,\I[4]_b0 ,\I[3]_b1 ,\I[3]_b0 ,
		\I[2]_b1 ,\I[2]_b0 ,\I[1]_b1 ,\I[1]_b0 ,\I[0]_b1 ,\I[0]_b0 ;
output \O[19]_b1 ,\O[19]_b0 ,\O[18]_b1 ,\O[18]_b0 ,\O[17]_b1 ,\O[17]_b0 ,\O[16]_b1 ,\O[16]_b0 ,\O[15]_b1 ,
		\O[15]_b0 ,\O[14]_b1 ,\O[14]_b0 ,\O[13]_b1 ,\O[13]_b0 ,\O[12]_b1 ,\O[12]_b0 ,\O[11]_b1 ,\O[11]_b0 ,
		\O[10]_b1 ,\O[10]_b0 ,\O[9]_b1 ,\O[9]_b0 ,\O[8]_b1 ,\O[8]_b0 ,\O[7]_b1 ,\O[7]_b0 ,\O[6]_b1 ,
		\O[6]_b0 ,\O[5]_b1 ,\O[5]_b0 ,\O[4]_b1 ,\O[4]_b0 ,\O[3]_b1 ,\O[3]_b0 ,\O[2]_b1 ,\O[2]_b0 ,
		\O[1]_b1 ,\O[1]_b0 ,\O[0]_b1 ,\O[0]_b0 ;

wire \69_ZERO_b1 , \69_ZERO_b0 , \70_b1 , \70_b0 , \71_ONE_b1 , \71_ONE_b0 , \72_b1 , \72_b0 , \73_b1 , \73_b0 , 
		\74_b1 , \74_b0 , \75_b1 , \75_b0 , \76_b1 , \76_b0 , \77_b1 , \77_b0 , \78_b1 , \78_b0 , 
		\79_b1 , \79_b0 , \80_b1 , \80_b0 , \81_b1 , \81_b0 , \82_b1 , \82_b0 , \83_b1 , \83_b0 , 
		\84_b1 , \84_b0 , \85_b1 , \85_b0 , \86_b1 , \86_b0 , \87_b1 , \87_b0 , \88_b1 , \88_b0 , 
		\89_b1 , \89_b0 , \90_b1 , \90_b0 , \91_b1 , \91_b0 , \92_b1 , \92_b0 , \93_b1 , \93_b0 , 
		\94_b1 , \94_b0 , \95_b1 , \95_b0 , \96_b1 , \96_b0 , \97_b1 , \97_b0 , \98_b1 , \98_b0 , 
		\99_b1 , \99_b0 , \100_b1 , \100_b0 , \101_b1 , \101_b0 , \102_b1 , \102_b0 , \103_b1 , \103_b0 , 
		\104_b1 , \104_b0 , \105_b1 , \105_b0 , \106_b1 , \106_b0 , \107_b1 , \107_b0 , \108_b1 , \108_b0 , 
		\109_b1 , \109_b0 , \110_b1 , \110_b0 , \111_b1 , \111_b0 , \112_b1 , \112_b0 , \113_b1 , \113_b0 , 
		\114_b1 , \114_b0 , \115_b1 , \115_b0 , \116_b1 , \116_b0 , \117_b1 , \117_b0 , \118_b1 , \118_b0 , 
		\119_b1 , \119_b0 , \120_b1 , \120_b0 , \121_b1 , \121_b0 , \122_b1 , \122_b0 , \123_b1 , \123_b0 , 
		\124_b1 , \124_b0 , \125_b1 , \125_b0 , \126_b1 , \126_b0 , \127_b1 , \127_b0 , \128_b1 , \128_b0 , 
		\129_b1 , \129_b0 , \130_b1 , \130_b0 , \131_b1 , \131_b0 , \132_b1 , \132_b0 , \133_b1 , \133_b0 , 
		\134_b1 , \134_b0 , \135_b1 , \135_b0 , \136_b1 , \136_b0 , \137_b1 , \137_b0 , \138_b1 , \138_b0 , 
		\139_b1 , \139_b0 , \140_b1 , \140_b0 , \141_b1 , \141_b0 , \142_b1 , \142_b0 , \143_b1 , \143_b0 , 
		\144_b1 , \144_b0 , \145_b1 , \145_b0 , \146_b1 , \146_b0 , \147_b1 , \147_b0 , \148_b1 , \148_b0 , 
		\149_b1 , \149_b0 , \150_b1 , \150_b0 , \151_b1 , \151_b0 , \152_b1 , \152_b0 , \153_b1 , \153_b0 , 
		\154_b1 , \154_b0 , \155_b1 , \155_b0 , \156_b1 , \156_b0 , \157_b1 , \157_b0 , \158_b1 , \158_b0 , 
		\159_b1 , \159_b0 , \160_b1 , \160_b0 , \161_b1 , \161_b0 , \162_b1 , \162_b0 , \163_b1 , \163_b0 , 
		\164_b1 , \164_b0 , \165_b1 , \165_b0 , \166_b1 , \166_b0 , \167_b1 , \167_b0 , \168_b1 , \168_b0 , 
		\169_b1 , \169_b0 , \170_b1 , \170_b0 , \171_b1 , \171_b0 , \172_b1 , \172_b0 , \173_b1 , \173_b0 , 
		\174_b1 , \174_b0 , \175_b1 , \175_b0 , \176_b1 , \176_b0 , \177_b1 , \177_b0 , \178_b1 , \178_b0 , 
		\179_b1 , \179_b0 , \180_b1 , \180_b0 , \181_b1 , \181_b0 , \182_b1 , \182_b0 , \183_b1 , \183_b0 , 
		\184_b1 , \184_b0 , \185_b1 , \185_b0 , \186_b1 , \186_b0 , \187_b1 , \187_b0 , \188_b1 , \188_b0 , 
		\189_b1 , \189_b0 , \190_b1 , \190_b0 , \191_b1 , \191_b0 , \192_b1 , \192_b0 , \193_b1 , \193_b0 , 
		\194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , \197_b1 , \197_b0 , \198_b1 , \198_b0 , 
		\199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , \202_b1 , \202_b0 , \203_b1 , \203_b0 , 
		\204_b1 , \204_b0 , \205_b1 , \205_b0 , \206_b1 , \206_b0 , \207_b1 , \207_b0 , \208_b1 , \208_b0 , 
		\209_b1 , \209_b0 , \210_b1 , \210_b0 , \211_b1 , \211_b0 , \212_b1 , \212_b0 , \213_b1 , \213_b0 , 
		\214_b1 , \214_b0 , \215_b1 , \215_b0 , \216_b1 , \216_b0 , \217_b1 , \217_b0 , \218_b1 , \218_b0 , 
		\219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , \222_b1 , \222_b0 , \223_b1 , \223_b0 , 
		\224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , \227_b1 , \227_b0 , \228_b1 , \228_b0 , 
		\229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , \232_b1 , \232_b0 , \233_b1 , \233_b0 , 
		\234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , \237_b1 , \237_b0 , \238_b1 , \238_b0 , 
		\239_b1 , \239_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , \242_b1 , \242_b0 , \243_b1 , \243_b0 , 
		\244_b1 , \244_b0 , \245_b1 , \245_b0 , \246_b1 , \246_b0 , \247_b1 , \247_b0 , \248_b1 , \248_b0 , 
		\249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , \252_b1 , \252_b0 , \253_b1 , \253_b0 , 
		\254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , \257_b1 , \257_b0 , \258_b1 , \258_b0 , 
		\259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , \262_b1 , \262_b0 , \263_b1 , \263_b0 , 
		\264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , \267_b1 , \267_b0 , \268_b1 , \268_b0 , 
		\269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , \272_b1 , \272_b0 , \273_b1 , \273_b0 , 
		\274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_b1 , \276_b0 , \277_b1 , \277_b0 , \278_b1 , \278_b0 , 
		\279_b1 , \279_b0 , \280_b1 , \280_b0 , \281_b1 , \281_b0 , \282_b1 , \282_b0 , \283_b1 , \283_b0 , 
		\284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , \287_b1 , \287_b0 , \288_b1 , \288_b0 , 
		\289_b1 , \289_b0 , \290_b1 , \290_b0 , \291_b1 , \291_b0 , \292_b1 , \292_b0 , \293_b1 , \293_b0 , 
		\294_b1 , \294_b0 , \295_b1 , \295_b0 , \296_b1 , \296_b0 , \297_b1 , \297_b0 , \298_b1 , \298_b0 , 
		\299_b1 , \299_b0 , \300_b1 , \300_b0 , \301_b1 , \301_b0 , \302_b1 , \302_b0 , \303_b1 , \303_b0 , 
		\304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , \307_b1 , \307_b0 , \308_b1 , \308_b0 , 
		\309_b1 , \309_b0 , \310_b1 , \310_b0 , \311_b1 , \311_b0 , \312_b1 , \312_b0 , \313_b1 , \313_b0 , 
		\314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_b1 , \316_b0 , \317_b1 , \317_b0 , \318_b1 , \318_b0 , 
		\319_b1 , \319_b0 , \320_b1 , \320_b0 , \321_b1 , \321_b0 , \322_b1 , \322_b0 , \323_b1 , \323_b0 , 
		\324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , \327_b1 , \327_b0 , \328_b1 , \328_b0 , 
		\329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_b1 , \331_b0 , \332_b1 , \332_b0 , \333_b1 , \333_b0 , 
		\334_b1 , \334_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , \337_b1 , \337_b0 , \338_b1 , \338_b0 , 
		\339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_b1 , \341_b0 , \342_b1 , \342_b0 , \343_b1 , \343_b0 , 
		\344_b1 , \344_b0 , \345_b1 , \345_b0 , \346_b1 , \346_b0 , \347_b1 , \347_b0 , \348_b1 , \348_b0 , 
		\349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , \352_b1 , \352_b0 , \353_b1 , \353_b0 , 
		\354_b1 , \354_b0 , \355_b1 , \355_b0 , \356_b1 , \356_b0 , \357_b1 , \357_b0 , \358_b1 , \358_b0 , 
		\359_b1 , \359_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , \362_b1 , \362_b0 , \363_b1 , \363_b0 , 
		\364_b1 , \364_b0 , \365_b1 , \365_b0 , \366_b1 , \366_b0 , \367_b1 , \367_b0 , \368_b1 , \368_b0 , 
		\369_b1 , \369_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , \372_b1 , \372_b0 , \373_b1 , \373_b0 , 
		\374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , \377_b1 , \377_b0 , \378_b1 , \378_b0 , 
		\379_b1 , \379_b0 , \380_b1 , \380_b0 , \381_b1 , \381_b0 , \382_b1 , \382_b0 , \383_b1 , \383_b0 , 
		\384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , \387_b1 , \387_b0 , \388_b1 , \388_b0 , 
		\389_b1 , \389_b0 , \390_b1 , \390_b0 , \391_b1 , \391_b0 , \392_b1 , \392_b0 , \393_b1 , \393_b0 , 
		\394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , \397_b1 , \397_b0 , \398_b1 , \398_b0 , 
		\399_b1 , \399_b0 , \400_b1 , \400_b0 , \401_b1 , \401_b0 , \402_b1 , \402_b0 , \403_b1 , \403_b0 , 
		\404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , \407_b1 , \407_b0 , \408_b1 , \408_b0 , 
		\409_b1 , \409_b0 , \410_b1 , \410_b0 , \411_b1 , \411_b0 , \412_b1 , \412_b0 , \413_b1 , \413_b0 , 
		\414_b1 , \414_b0 , \415_b1 , \415_b0 , \416_b1 , \416_b0 , \417_b1 , \417_b0 , \418_b1 , \418_b0 , 
		\419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , \422_b1 , \422_b0 , \423_b1 , \423_b0 , 
		\424_b1 , \424_b0 , \425_b1 , \425_b0 , \426_b1 , \426_b0 , \427_b1 , \427_b0 , \428_b1 , \428_b0 , 
		\429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , \432_b1 , \432_b0 , \433_b1 , \433_b0 , 
		\434_b1 , \434_b0 , \435_b1 , \435_b0 , \436_b1 , \436_b0 , \437_b1 , \437_b0 , \438_b1 , \438_b0 , 
		\439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , \442_b1 , \442_b0 , \443_b1 , \443_b0 , 
		\444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_b1 , \446_b0 , \447_b1 , \447_b0 , \448_b1 , \448_b0 , 
		\449_b1 , \449_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , \452_b1 , \452_b0 , \453_b1 , \453_b0 , 
		\454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_b1 , \456_b0 , \457_b1 , \457_b0 , \458_b1 , \458_b0 , 
		\459_b1 , \459_b0 , \460_b1 , \460_b0 , \461_b1 , \461_b0 , \462_b1 , \462_b0 , \463_b1 , \463_b0 , 
		\464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , \467_b1 , \467_b0 , \468_b1 , \468_b0 , 
		\469_b1 , \469_b0 , \470_b1 , \470_b0 , \471_b1 , \471_b0 , \472_b1 , \472_b0 , \473_b1 , \473_b0 , 
		\474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , \477_b1 , \477_b0 , \478_b1 , \478_b0 , 
		\479_b1 , \479_b0 , \480_b1 , \480_b0 , \481_b1 , \481_b0 , \482_b1 , \482_b0 , \483_b1 , \483_b0 , 
		\484_b1 , \484_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , \487_b1 , \487_b0 , \488_b1 , \488_b0 , 
		\489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , \492_b1 , \492_b0 , \493_b1 , \493_b0 , 
		\494_b1 , \494_b0 , \495_b1 , \495_b0 , \496_b1 , \496_b0 , \497_b1 , \497_b0 , \498_b1 , \498_b0 , 
		\499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , \502_b1 , \502_b0 , \503_b1 , \503_b0 , 
		\504_b1 , \504_b0 , \505_b1 , \505_b0 , \506_b1 , \506_b0 , \507_b1 , \507_b0 , \508_b1 , \508_b0 , 
		\509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , \512_b1 , \512_b0 , \513_b1 , \513_b0 , 
		\514_b1 , \514_b0 , \515_b1 , \515_b0 , \516_b1 , \516_b0 , \517_b1 , \517_b0 , \518_b1 , \518_b0 , 
		\519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , \522_b1 , \522_b0 , \523_b1 , \523_b0 , 
		\524_b1 , \524_b0 , \525_b1 , \525_b0 , \526_b1 , \526_b0 , \527_b1 , \527_b0 , \528_b1 , \528_b0 , 
		\529_b1 , \529_b0 , \530_b1 , \530_b0 , \531_b1 , \531_b0 , \532_b1 , \532_b0 , \533_b1 , \533_b0 , 
		\534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_b1 , \536_b0 , \537_b1 , \537_b0 , \538_b1 , \538_b0 , 
		\539_b1 , \539_b0 , \540_b1 , \540_b0 , \541_b1 , \541_b0 , \542_b1 , \542_b0 , \543_b1 , \543_b0 , 
		\544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , \547_b1 , \547_b0 , \548_b1 , \548_b0 , 
		\549_b1 , \549_b0 , \550_b1 , \550_b0 , \551_b1 , \551_b0 , \552_b1 , \552_b0 , \553_b1 , \553_b0 , 
		\554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , \557_b1 , \557_b0 , \558_b1 , \558_b0 , 
		\559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_b1 , \561_b0 , \562_b1 , \562_b0 , \563_b1 , \563_b0 , 
		\564_b1 , \564_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , \567_b1 , \567_b0 , \568_b1 , \568_b0 , 
		\569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_b1 , \571_b0 , \572_b1 , \572_b0 , \573_b1 , \573_b0 , 
		\574_b1 , \574_b0 , \575_b1 , \575_b0 , \576_b1 , \576_b0 , \577_b1 , \577_b0 , \578_b1 , \578_b0 , 
		\579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , \582_b1 , \582_b0 , \583_b1 , \583_b0 , 
		\584_b1 , \584_b0 , \585_b1 , \585_b0 , \586_b1 , \586_b0 , \587_b1 , \587_b0 , \588_b1 , \588_b0 , 
		\589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , \592_b1 , \592_b0 , \593_b1 , \593_b0 , 
		\594_b1 , \594_b0 , \595_b1 , \595_b0 , \596_b1 , \596_b0 , \597_b1 , \597_b0 , \598_b1 , \598_b0 , 
		\599_b1 , \599_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , \602_b1 , \602_b0 , \603_b1 , \603_b0 , 
		\604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_b1 , \606_b0 , \607_b1 , \607_b0 , \608_b1 , \608_b0 , 
		\609_b1 , \609_b0 , \610_b1 , \610_b0 , \611_b1 , \611_b0 , \612_b1 , \612_b0 , \613_b1 , \613_b0 , 
		\614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , \617_b1 , \617_b0 , \618_b1 , \618_b0 , 
		\619_b1 , \619_b0 , \620_b1 , \620_b0 , \621_b1 , \621_b0 , \622_b1 , \622_b0 , \623_b1 , \623_b0 , 
		\624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , \627_b1 , \627_b0 , \628_b1 , \628_b0 , 
		\629_b1 , \629_b0 , \630_b1 , \630_b0 , \631_b1 , \631_b0 , \632_b1 , \632_b0 , \633_b1 , \633_b0 , 
		\634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , \637_b1 , \637_b0 , \638_b1 , \638_b0 , 
		\639_b1 , \639_b0 , \640_b1 , \640_b0 , \641_b1 , \641_b0 , \642_b1 , \642_b0 , \643_b1 , \643_b0 , 
		\644_b1 , \644_b0 , \645_b1 , \645_b0 , \646_b1 , \646_b0 , \647_b1 , \647_b0 , \648_b1 , \648_b0 , 
		\649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , \652_b1 , \652_b0 , \653_b1 , \653_b0 , 
		\654_b1 , \654_b0 , \655_b1 , \655_b0 , \656_b1 , \656_b0 , \657_b1 , \657_b0 , \658_b1 , \658_b0 , 
		\659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , \662_b1 , \662_b0 , \663_b1 , \663_b0 , 
		\664_b1 , \664_b0 , \665_b1 , \665_b0 , \666_b1 , \666_b0 , \667_b1 , \667_b0 , \668_b1 , \668_b0 , 
		\669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , \672_b1 , \672_b0 , \673_b1 , \673_b0 , 
		\674_b1 , \674_b0 , \675_b1 , \675_b0 , \676_b1 , \676_b0 , \677_b1 , \677_b0 , \678_b1 , \678_b0 , 
		\679_b1 , \679_b0 , \680_b1 , \680_b0 , \681_b1 , \681_b0 , \682_b1 , \682_b0 , \683_b1 , \683_b0 , 
		\684_b1 , \684_b0 , \685_b1 , \685_b0 , \686_b1 , \686_b0 , \687_b1 , \687_b0 , \688_b1 , \688_b0 , 
		\689_b1 , \689_b0 , \690_b1 , \690_b0 , \691_b1 , \691_b0 , \692_b1 , \692_b0 , \693_b1 , \693_b0 , 
		\694_b1 , \694_b0 , \695_b1 , \695_b0 , \696_b1 , \696_b0 , \697_b1 , \697_b0 , \698_b1 , \698_b0 , 
		\699_b1 , \699_b0 , \700_b1 , \700_b0 , \701_b1 , \701_b0 , \702_b1 , \702_b0 , \703_b1 , \703_b0 , 
		\704_b1 , \704_b0 , \705_b1 , \705_b0 , \706_b1 , \706_b0 , \707_b1 , \707_b0 , \708_b1 , \708_b0 , 
		\709_b1 , \709_b0 , \710_b1 , \710_b0 , \711_b1 , \711_b0 , \712_b1 , \712_b0 , \713_b1 , \713_b0 , 
		\714_b1 , \714_b0 , \715_b1 , \715_b0 , \716_b1 , \716_b0 , \717_b1 , \717_b0 , \718_b1 , \718_b0 , 
		\719_b1 , \719_b0 , \720_b1 , \720_b0 , \721_b1 , \721_b0 , \722_b1 , \722_b0 , \723_b1 , \723_b0 , 
		\724_b1 , \724_b0 , \725_b1 , \725_b0 , \726_b1 , \726_b0 , \727_b1 , \727_b0 , \728_b1 , \728_b0 , 
		\729_b1 , \729_b0 , \730_b1 , \730_b0 , \731_b1 , \731_b0 , \732_b1 , \732_b0 , \733_b1 , \733_b0 , 
		\734_b1 , \734_b0 , \735_b1 , \735_b0 , \736_b1 , \736_b0 , \737_b1 , \737_b0 , \738_b1 , \738_b0 , 
		\739_b1 , \739_b0 , \740_b1 , \740_b0 , \741_b1 , \741_b0 , \742_b1 , \742_b0 , \743_b1 , \743_b0 , 
		\744_b1 , \744_b0 , \745_b1 , \745_b0 , \746_b1 , \746_b0 , \747_b1 , \747_b0 , \748_b1 , \748_b0 , 
		\749_b1 , \749_b0 , \750_b1 , \750_b0 , \751_b1 , \751_b0 , \752_b1 , \752_b0 , \753_b1 , \753_b0 , 
		\754_b1 , \754_b0 , \755_b1 , \755_b0 , \756_b1 , \756_b0 , \757_b1 , \757_b0 , \758_b1 , \758_b0 , 
		\759_b1 , \759_b0 , \760_b1 , \760_b0 , \761_b1 , \761_b0 , \762_b1 , \762_b0 , \763_b1 , \763_b0 , 
		\764_b1 , \764_b0 , \765_b1 , \765_b0 , \766_b1 , \766_b0 , \767_b1 , \767_b0 , \768_b1 , \768_b0 , 
		\769_b1 , \769_b0 , \770_b1 , \770_b0 , \771_b1 , \771_b0 , \772_b1 , \772_b0 , \773_b1 , \773_b0 , 
		\774_b1 , \774_b0 , \775_b1 , \775_b0 , \776_b1 , \776_b0 , \777_b1 , \777_b0 , \778_b1 , \778_b0 , 
		\779_b1 , \779_b0 , \780_b1 , \780_b0 , \781_b1 , \781_b0 , \782_b1 , \782_b0 , \783_b1 , \783_b0 , 
		\784_b1 , \784_b0 , \785_b1 , \785_b0 , \786_b1 , \786_b0 , \787_b1 , \787_b0 , \788_b1 , \788_b0 , 
		\789_b1 , \789_b0 , \790_b1 , \790_b0 , \791_b1 , \791_b0 , \792_b1 , \792_b0 , \793_b1 , \793_b0 , 
		\794_b1 , \794_b0 , \795_b1 , \795_b0 , \796_b1 , \796_b0 , \797_b1 , \797_b0 , \798_b1 , \798_b0 , 
		\799_b1 , \799_b0 , \800_b1 , \800_b0 , \801_b1 , \801_b0 , \802_b1 , \802_b0 , \803_b1 , \803_b0 , 
		\804_b1 , \804_b0 , \805_b1 , \805_b0 , \806_b1 , \806_b0 , \807_b1 , \807_b0 , \808_b1 , \808_b0 , 
		\809_b1 , \809_b0 , \810_b1 , \810_b0 , \811_b1 , \811_b0 , \812_b1 , \812_b0 , \813_b1 , \813_b0 , 
		\814_b1 , \814_b0 , \815_b1 , \815_b0 , \816_b1 , \816_b0 , \817_b1 , \817_b0 , \818_b1 , \818_b0 , 
		\819_b1 , \819_b0 , \820_b1 , \820_b0 , \821_b1 , \821_b0 , \822_b1 , \822_b0 , \823_b1 , \823_b0 , 
		\824_b1 , \824_b0 , \825_b1 , \825_b0 , \826_b1 , \826_b0 , \827_b1 , \827_b0 , \828_b1 , \828_b0 , 
		\829_b1 , \829_b0 , \830_b1 , \830_b0 , \831_b1 , \831_b0 , \832_b1 , \832_b0 , \833_b1 , \833_b0 , 
		\834_b1 , \834_b0 , \835_b1 , \835_b0 , \836_b1 , \836_b0 , \837_b1 , \837_b0 , \838_b1 , \838_b0 , 
		\839_b1 , \839_b0 , \840_b1 , \840_b0 , \841_b1 , \841_b0 , \842_b1 , \842_b0 , \843_b1 , \843_b0 , 
		\844_b1 , \844_b0 , \845_b1 , \845_b0 , \846_b1 , \846_b0 , \847_b1 , \847_b0 , \848_b1 , \848_b0 , 
		\849_b1 , \849_b0 , \850_b1 , \850_b0 , \851_b1 , \851_b0 , \852_b1 , \852_b0 , \853_b1 , \853_b0 , 
		\854_b1 , \854_b0 , \855_b1 , \855_b0 , \856_b1 , \856_b0 , \857_b1 , \857_b0 , \858_b1 , \858_b0 , 
		\859_b1 , \859_b0 , \860_b1 , \860_b0 , \861_b1 , \861_b0 , \862_b1 , \862_b0 , \863_b1 , \863_b0 , 
		\864_b1 , \864_b0 , \865_b1 , \865_b0 , \866_b1 , \866_b0 , \867_b1 , \867_b0 , \868_b1 , \868_b0 , 
		\869_b1 , \869_b0 , \870_b1 , \870_b0 , \871_b1 , \871_b0 , \872_b1 , \872_b0 , \873_b1 , \873_b0 , 
		\874_b1 , \874_b0 , \875_b1 , \875_b0 , \876_b1 , \876_b0 , \877_b1 , \877_b0 , \878_b1 , \878_b0 , 
		\879_b1 , \879_b0 , \880_b1 , \880_b0 , \881_b1 , \881_b0 , \882_b1 , \882_b0 , \883_b1 , \883_b0 , 
		\884_b1 , \884_b0 , \885_b1 , \885_b0 , \886_b1 , \886_b0 , \887_b1 , \887_b0 , \888_b1 , \888_b0 , 
		\889_b1 , \889_b0 , \890_b1 , \890_b0 , \891_b1 , \891_b0 , \892_b1 , \892_b0 , \893_b1 , \893_b0 , 
		\894_b1 , \894_b0 , \895_b1 , \895_b0 , \896_b1 , \896_b0 , \897_b1 , \897_b0 , \898_b1 , \898_b0 , 
		\899_b1 , \899_b0 , \900_b1 , \900_b0 , \901_b1 , \901_b0 , \902_b1 , \902_b0 , \903_b1 , \903_b0 , 
		\904_b1 , \904_b0 , \905_b1 , \905_b0 , \906_b1 , \906_b0 , \907_b1 , \907_b0 , \908_b1 , \908_b0 , 
		\909_b1 , \909_b0 , \910_b1 , \910_b0 , \911_b1 , \911_b0 , \912_b1 , \912_b0 , \913_b1 , \913_b0 , 
		\914_b1 , \914_b0 , \915_b1 , \915_b0 , \916_b1 , \916_b0 , \917_b1 , \917_b0 , \918_b1 , \918_b0 , 
		\919_b1 , \919_b0 , \920_b1 , \920_b0 , \921_b1 , \921_b0 , \922_b1 , \922_b0 , \923_b1 , \923_b0 , 
		\924_b1 , \924_b0 , \925_b1 , \925_b0 , \926_b1 , \926_b0 , \927_b1 , \927_b0 , \928_b1 , \928_b0 , 
		\929_b1 , \929_b0 , \930_b1 , \930_b0 , \931_b1 , \931_b0 , \932_b1 , \932_b0 , \933_b1 , \933_b0 , 
		\934_b1 , \934_b0 , \935_b1 , \935_b0 , \936_b1 , \936_b0 , \937_b1 , \937_b0 , \938_b1 , \938_b0 , 
		\939_b1 , \939_b0 , \940_b1 , \940_b0 , \941_b1 , \941_b0 , \942_b1 , \942_b0 , \943_b1 , \943_b0 , 
		\944_b1 , \944_b0 , \945_b1 , \945_b0 , \946_b1 , \946_b0 , \947_b1 , \947_b0 , \948_b1 , \948_b0 , 
		\949_b1 , \949_b0 , \950_b1 , \950_b0 , \951_b1 , \951_b0 , \952_b1 , \952_b0 , \953_b1 , \953_b0 , 
		\954_b1 , \954_b0 , \955_b1 , \955_b0 , \956_b1 , \956_b0 , \957_b1 , \957_b0 , \958_b1 , \958_b0 , 
		\959_b1 , \959_b0 , \960_b1 , \960_b0 , \961_b1 , \961_b0 , \962_b1 , \962_b0 , \963_b1 , \963_b0 , 
		\964_b1 , \964_b0 , \965_b1 , \965_b0 , \966_b1 , \966_b0 , \967_b1 , \967_b0 , \968_b1 , \968_b0 , 
		\969_b1 , \969_b0 , \970_b1 , \970_b0 , \971_b1 , \971_b0 , \972_b1 , \972_b0 , \973_b1 , \973_b0 , 
		\974_b1 , \974_b0 , \975_b1 , \975_b0 , \976_b1 , \976_b0 , \977_b1 , \977_b0 , \978_b1 , \978_b0 , 
		\979_b1 , \979_b0 , \980_b1 , \980_b0 , \981_b1 , \981_b0 , \982_b1 , \982_b0 , \983_b1 , \983_b0 , 
		\984_b1 , \984_b0 , \985_b1 , \985_b0 , \986_b1 , \986_b0 , \987_b1 , \987_b0 , \988_b1 , \988_b0 , 
		\989_b1 , \989_b0 , \990_b1 , \990_b0 , \991_b1 , \991_b0 , \992_b1 , \992_b0 , \993_b1 , \993_b0 , 
		\994_b1 , \994_b0 , \995_b1 , \995_b0 , \996_b1 , \996_b0 , \997_b1 , \997_b0 , \998_b1 , \998_b0 , 
		\999_b1 , \999_b0 , \1000_b1 , \1000_b0 , \1001_b1 , \1001_b0 , \1002_b1 , \1002_b0 , \1003_b1 , \1003_b0 , 
		\1004_b1 , \1004_b0 , \1005_b1 , \1005_b0 , \1006_b1 , \1006_b0 , \1007_b1 , \1007_b0 , \1008_b1 , \1008_b0 , 
		\1009_b1 , \1009_b0 , \1010_b1 , \1010_b0 , \1011_b1 , \1011_b0 , \1012_b1 , \1012_b0 , \1013_b1 , \1013_b0 , 
		\1014_b1 , \1014_b0 , \1015_b1 , \1015_b0 , \1016_b1 , \1016_b0 , \1017_b1 , \1017_b0 , \1018_b1 , \1018_b0 , 
		\1019_b1 , \1019_b0 , \1020_b1 , \1020_b0 , \1021_b1 , \1021_b0 , \1022_b1 , \1022_b0 , \1023_b1 , \1023_b0 , 
		\1024_b1 , \1024_b0 , \1025_b1 , \1025_b0 , \1026_b1 , \1026_b0 , \1027_b1 , \1027_b0 , \1028_b1 , \1028_b0 , 
		\1029_b1 , \1029_b0 , \1030_b1 , \1030_b0 , \1031_b1 , \1031_b0 , \1032_b1 , \1032_b0 , \1033_b1 , \1033_b0 , 
		\1034_b1 , \1034_b0 , \1035_b1 , \1035_b0 , \1036_b1 , \1036_b0 , \1037_b1 , \1037_b0 , \1038_b1 , \1038_b0 , 
		\1039_b1 , \1039_b0 , \1040_b1 , \1040_b0 , \1041_b1 , \1041_b0 , \1042_b1 , \1042_b0 , \1043_b1 , \1043_b0 , 
		\1044_b1 , \1044_b0 , \1045_b1 , \1045_b0 , \1046_b1 , \1046_b0 , \1047_b1 , \1047_b0 , \1048_b1 , \1048_b0 , 
		\1049_b1 , \1049_b0 , \1050_b1 , \1050_b0 , \1051_b1 , \1051_b0 , \1052_b1 , \1052_b0 , \1053_b1 , \1053_b0 , 
		\1054_b1 , \1054_b0 , \1055_b1 , \1055_b0 , \1056_b1 , \1056_b0 , \1057_b1 , \1057_b0 , \1058_b1 , \1058_b0 , 
		\1059_b1 , \1059_b0 , \1060_b1 , \1060_b0 , \1061_b1 , \1061_b0 , \1062_b1 , \1062_b0 , \1063_b1 , \1063_b0 , 
		\1064_b1 , \1064_b0 , \1065_b1 , \1065_b0 , \1066_b1 , \1066_b0 , \1067_b1 , \1067_b0 , \1068_b1 , \1068_b0 , 
		\1069_b1 , \1069_b0 , \1070_b1 , \1070_b0 , \1071_b1 , \1071_b0 , \1072_b1 , \1072_b0 , \1073_b1 , \1073_b0 , 
		\1074_b1 , \1074_b0 , \1075_b1 , \1075_b0 , w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , 
		w_6 , w_7 , w_8 , w_9 , w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , 
		w_16 , w_17 , w_18 , w_19 , w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , 
		w_26 , w_27 , w_28 , w_29 , w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , 
		w_36 , w_37 , w_38 , w_39 , w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , 
		w_46 , w_47 , w_48 , w_49 , w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , 
		w_56 , w_57 , w_58 , w_59 , w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , 
		w_66 , w_67 , w_68 , w_69 , w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , 
		w_76 , w_77 , w_78 , w_79 , w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , 
		w_86 , w_87 , w_88 , w_89 , w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , 
		w_96 , w_97 , w_98 , w_99 , w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , 
		w_106 , w_107 , w_108 , w_109 , w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , 
		w_116 , w_117 , w_118 , w_119 , w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , 
		w_126 , w_127 , w_128 , w_129 , w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , 
		w_136 , w_137 , w_138 , w_139 , w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , 
		w_146 , w_147 , w_148 , w_149 , w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , 
		w_156 , w_157 , w_158 , w_159 , w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , 
		w_166 , w_167 , w_168 , w_169 , w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , 
		w_176 , w_177 , w_178 , w_179 , w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , 
		w_186 , w_187 , w_188 , w_189 , w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , 
		w_196 , w_197 , w_198 , w_199 , w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , 
		w_206 , w_207 , w_208 , w_209 , w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , 
		w_216 , w_217 , w_218 , w_219 , w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , 
		w_226 , w_227 , w_228 , w_229 , w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , 
		w_236 , w_237 , w_238 , w_239 , w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , 
		w_246 , w_247 , w_248 , w_249 , w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , 
		w_256 , w_257 , w_258 , w_259 , w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , 
		w_266 , w_267 , w_268 , w_269 , w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , 
		w_276 , w_277 , w_278 , w_279 , w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , 
		w_286 , w_287 , w_288 , w_289 , w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , 
		w_296 , w_297 , w_298 , w_299 , w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , 
		w_306 , w_307 , w_308 , w_309 , w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , 
		w_316 , w_317 , w_318 , w_319 , w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , 
		w_326 , w_327 , w_328 , w_329 , w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , 
		w_336 , w_337 , w_338 , w_339 , w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , 
		w_346 , w_347 , w_348 , w_349 , w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , 
		w_356 , w_357 , w_358 , w_359 , w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , 
		w_366 , w_367 , w_368 , w_369 , w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , 
		w_376 , w_377 , w_378 , w_379 , w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , 
		w_386 , w_387 , w_388 , w_389 , w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , 
		w_396 , w_397 , w_398 , w_399 , w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , 
		w_406 , w_407 , w_408 , w_409 , w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , 
		w_416 , w_417 , w_418 , w_419 , w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , 
		w_426 , w_427 , w_428 , w_429 , w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , 
		w_436 , w_437 , w_438 , w_439 , w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , 
		w_446 , w_447 , w_448 , w_449 , w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , 
		w_456 , w_457 , w_458 , w_459 , w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , 
		w_466 , w_467 , w_468 , w_469 , w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , 
		w_476 , w_477 , w_478 , w_479 , w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , 
		w_486 , w_487 , w_488 , w_489 , w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , 
		w_496 , w_497 , w_498 , w_499 , w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , 
		w_506 , w_507 , w_508 , w_509 , w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , 
		w_516 , w_517 , w_518 , w_519 , w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , 
		w_526 , w_527 , w_528 , w_529 , w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , 
		w_536 , w_537 , w_538 , w_539 , w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , 
		w_546 , w_547 , w_548 , w_549 , w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , 
		w_556 , w_557 , w_558 , w_559 , w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , 
		w_566 , w_567 , w_568 , w_569 , w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , 
		w_576 , w_577 , w_578 , w_579 , w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , 
		w_586 , w_587 , w_588 , w_589 , w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , 
		w_596 , w_597 , w_598 , w_599 , w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , 
		w_606 , w_607 , w_608 , w_609 , w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , 
		w_616 , w_617 , w_618 , w_619 , w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , 
		w_626 , w_627 , w_628 , w_629 , w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , 
		w_636 , w_637 , w_638 , w_639 , w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , 
		w_646 , w_647 , w_648 , w_649 , w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , 
		w_656 , w_657 , w_658 , w_659 , w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , 
		w_666 , w_667 , w_668 , w_669 , w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , 
		w_676 , w_677 , w_678 , w_679 , w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , 
		w_686 , w_687 , w_688 , w_689 , w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , 
		w_696 , w_697 , w_698 , w_699 , w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , 
		w_706 , w_707 , w_708 , w_709 , w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , 
		w_716 , w_717 , w_718 , w_719 , w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , 
		w_726 , w_727 , w_728 , w_729 , w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , 
		w_736 , w_737 , w_738 , w_739 , w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , 
		w_746 , w_747 , w_748 , w_749 , w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , 
		w_756 , w_757 , w_758 , w_759 , w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , 
		w_766 , w_767 , w_768 , w_769 , w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , 
		w_776 , w_777 , w_778 , w_779 , w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , 
		w_786 , w_787 , w_788 , w_789 , w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , 
		w_796 , w_797 , w_798 , w_799 , w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , 
		w_806 , w_807 , w_808 , w_809 , w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , 
		w_816 , w_817 , w_818 , w_819 , w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , 
		w_826 , w_827 , w_828 , w_829 , w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , 
		w_836 , w_837 , w_838 , w_839 , w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , 
		w_846 , w_847 , w_848 , w_849 , w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , 
		w_856 , w_857 , w_858 , w_859 , w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , 
		w_866 , w_867 , w_868 , w_869 , w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , 
		w_876 , w_877 , w_878 , w_879 , w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , 
		w_886 , w_887 , w_888 , w_889 , w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , 
		w_896 , w_897 , w_898 , w_899 , w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , 
		w_906 , w_907 , w_908 , w_909 , w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , 
		w_916 , w_917 , w_918 , w_919 , w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , 
		w_926 , w_927 , w_928 , w_929 , w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , 
		w_936 , w_937 , w_938 , w_939 , w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , 
		w_946 , w_947 , w_948 , w_949 , w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , 
		w_956 , w_957 , w_958 , w_959 , w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , 
		w_966 , w_967 , w_968 , w_969 , w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , 
		w_976 , w_977 , w_978 , w_979 , w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , 
		w_986 , w_987 , w_988 , w_989 , w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , 
		w_996 , w_997 , w_998 , w_999 , w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , 
		w_1006 , w_1007 , w_1008 , w_1009 , w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , 
		w_1016 , w_1017 , w_1018 , w_1019 , w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , 
		w_1026 , w_1027 , w_1028 , w_1029 , w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , 
		w_1036 , w_1037 , w_1038 , w_1039 , w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , 
		w_1046 , w_1047 , w_1048 , w_1049 , w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , 
		w_1056 , w_1057 , w_1058 , w_1059 , w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , 
		w_1066 , w_1067 , w_1068 , w_1069 , w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , 
		w_1076 , w_1077 , w_1078 , w_1079 , w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , 
		w_1086 , w_1087 , w_1088 , w_1089 , w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , 
		w_1096 , w_1097 , w_1098 , w_1099 , w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , 
		w_1106 , w_1107 , w_1108 , w_1109 , w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , 
		w_1116 , w_1117 , w_1118 , w_1119 , w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , 
		w_1126 , w_1127 , w_1128 , w_1129 , w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , 
		w_1136 , w_1137 , w_1138 , w_1139 , w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , 
		w_1146 , w_1147 , w_1148 , w_1149 , w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , 
		w_1156 , w_1157 , w_1158 , w_1159 , w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , 
		w_1166 , w_1167 , w_1168 , w_1169 , w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , 
		w_1176 , w_1177 , w_1178 , w_1179 , w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , 
		w_1186 , w_1187 , w_1188 , w_1189 , w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , 
		w_1196 , w_1197 , w_1198 , w_1199 , w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , 
		w_1206 , w_1207 , w_1208 , w_1209 , w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , 
		w_1216 , w_1217 , w_1218 , w_1219 , w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , 
		w_1226 , w_1227 , w_1228 , w_1229 , w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , 
		w_1236 , w_1237 , w_1238 , w_1239 , w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , 
		w_1246 , w_1247 , w_1248 , w_1249 , w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , 
		w_1256 , w_1257 , w_1258 , w_1259 , w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , 
		w_1266 , w_1267 , w_1268 , w_1269 , w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , 
		w_1276 , w_1277 , w_1278 , w_1279 , w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , 
		w_1286 , w_1287 , w_1288 , w_1289 , w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , 
		w_1296 , w_1297 , w_1298 , w_1299 , w_1300 , w_1301 , w_1302 , w_1303 , w_1304 , w_1305 , 
		w_1306 , w_1307 , w_1308 , w_1309 , w_1310 , w_1311 , w_1312 , w_1313 , w_1314 , w_1315 , 
		w_1316 , w_1317 , w_1318 , w_1319 , w_1320 , w_1321 , w_1322 , w_1323 , w_1324 , w_1325 , 
		w_1326 , w_1327 , w_1328 , w_1329 , w_1330 , w_1331 , w_1332 , w_1333 , w_1334 , w_1335 , 
		w_1336 , w_1337 , w_1338 , w_1339 , w_1340 , w_1341 , w_1342 , w_1343 , w_1344 , w_1345 , 
		w_1346 , w_1347 , w_1348 , w_1349 , w_1350 , w_1351 , w_1352 , w_1353 , w_1354 , w_1355 , 
		w_1356 , w_1357 , w_1358 , w_1359 , w_1360 , w_1361 , w_1362 , w_1363 , w_1364 , w_1365 , 
		w_1366 , w_1367 , w_1368 , w_1369 , w_1370 , w_1371 , w_1372 , w_1373 , w_1374 , w_1375 , 
		w_1376 , w_1377 , w_1378 , w_1379 , w_1380 , w_1381 , w_1382 , w_1383 , w_1384 , w_1385 , 
		w_1386 , w_1387 , w_1388 , w_1389 , w_1390 , w_1391 , w_1392 , w_1393 , w_1394 , w_1395 , 
		w_1396 , w_1397 , w_1398 , w_1399 , w_1400 , w_1401 , w_1402 , w_1403 , w_1404 , w_1405 , 
		w_1406 , w_1407 , w_1408 , w_1409 , w_1410 , w_1411 , w_1412 , w_1413 , w_1414 , w_1415 , 
		w_1416 , w_1417 , w_1418 , w_1419 , w_1420 , w_1421 , w_1422 , w_1423 , w_1424 , w_1425 , 
		w_1426 , w_1427 , w_1428 , w_1429 , w_1430 , w_1431 , w_1432 , w_1433 , w_1434 , w_1435 , 
		w_1436 , w_1437 , w_1438 , w_1439 , w_1440 , w_1441 , w_1442 , w_1443 , w_1444 , w_1445 , 
		w_1446 , w_1447 , w_1448 , w_1449 , w_1450 , w_1451 , w_1452 , w_1453 , w_1454 , w_1455 , 
		w_1456 , w_1457 , w_1458 , w_1459 , w_1460 , w_1461 , w_1462 , w_1463 , w_1464 , w_1465 , 
		w_1466 , w_1467 , w_1468 , w_1469 , w_1470 , w_1471 , w_1472 , w_1473 , w_1474 , w_1475 , 
		w_1476 , w_1477 , w_1478 , w_1479 , w_1480 , w_1481 , w_1482 , w_1483 , w_1484 , w_1485 , 
		w_1486 , w_1487 , w_1488 , w_1489 , w_1490 , w_1491 , w_1492 , w_1493 , w_1494 , w_1495 , 
		w_1496 , w_1497 , w_1498 , w_1499 , w_1500 , w_1501 , w_1502 , w_1503 , w_1504 , w_1505 , 
		w_1506 , w_1507 , w_1508 , w_1509 , w_1510 , w_1511 , w_1512 , w_1513 , w_1514 , w_1515 , 
		w_1516 , w_1517 , w_1518 , w_1519 , w_1520 , w_1521 , w_1522 , w_1523 , w_1524 , w_1525 , 
		w_1526 , w_1527 , w_1528 , w_1529 , w_1530 , w_1531 , w_1532 , w_1533 , w_1534 , w_1535 , 
		w_1536 , w_1537 , w_1538 , w_1539 , w_1540 , w_1541 , w_1542 , w_1543 , w_1544 , w_1545 , 
		w_1546 , w_1547 , w_1548 , w_1549 , w_1550 , w_1551 , w_1552 , w_1553 , w_1554 , w_1555 , 
		w_1556 , w_1557 , w_1558 , w_1559 , w_1560 , w_1561 , w_1562 , w_1563 , w_1564 , w_1565 , 
		w_1566 , w_1567 , w_1568 , w_1569 , w_1570 , w_1571 , w_1572 , w_1573 , w_1574 , w_1575 , 
		w_1576 , w_1577 , w_1578 , w_1579 , w_1580 , w_1581 , w_1582 , w_1583 , w_1584 , w_1585 , 
		w_1586 , w_1587 , w_1588 , w_1589 , w_1590 , w_1591 , w_1592 , w_1593 , w_1594 , w_1595 , 
		w_1596 , w_1597 , w_1598 , w_1599 , w_1600 , w_1601 , w_1602 , w_1603 , w_1604 , w_1605 , 
		w_1606 , w_1607 , w_1608 , w_1609 , w_1610 , w_1611 , w_1612 , w_1613 , w_1614 , w_1615 , 
		w_1616 , w_1617 , w_1618 , w_1619 , w_1620 , w_1621 , w_1622 , w_1623 , w_1624 , w_1625 , 
		w_1626 , w_1627 , w_1628 , w_1629 , w_1630 , w_1631 , w_1632 , w_1633 , w_1634 , w_1635 , 
		w_1636 , w_1637 , w_1638 , w_1639 , w_1640 , w_1641 , w_1642 , w_1643 , w_1644 , w_1645 , 
		w_1646 , w_1647 , w_1648 , w_1649 , w_1650 , w_1651 , w_1652 , w_1653 , w_1654 , w_1655 , 
		w_1656 , w_1657 , w_1658 , w_1659 , w_1660 , w_1661 , w_1662 , w_1663 , w_1664 , w_1665 , 
		w_1666 , w_1667 , w_1668 , w_1669 , w_1670 , w_1671 , w_1672 , w_1673 , w_1674 , w_1675 , 
		w_1676 , w_1677 , w_1678 , w_1679 , w_1680 , w_1681 , w_1682 , w_1683 , w_1684 , w_1685 , 
		w_1686 , w_1687 , w_1688 , w_1689 , w_1690 , w_1691 , w_1692 , w_1693 , w_1694 , w_1695 , 
		w_1696 , w_1697 , w_1698 , w_1699 , w_1700 , w_1701 , w_1702 , w_1703 , w_1704 , w_1705 , 
		w_1706 , w_1707 , w_1708 , w_1709 , w_1710 , w_1711 , w_1712 , w_1713 , w_1714 , w_1715 , 
		w_1716 , w_1717 , w_1718 , w_1719 , w_1720 , w_1721 , w_1722 , w_1723 , w_1724 , w_1725 , 
		w_1726 , w_1727 , w_1728 , w_1729 , w_1730 , w_1731 , w_1732 , w_1733 , w_1734 , w_1735 , 
		w_1736 , w_1737 , w_1738 , w_1739 , w_1740 , w_1741 , w_1742 , w_1743 , w_1744 , w_1745 , 
		w_1746 , w_1747 , w_1748 , w_1749 , w_1750 , w_1751 , w_1752 , w_1753 , w_1754 , w_1755 , 
		w_1756 , w_1757 , w_1758 , w_1759 , w_1760 , w_1761 , w_1762 , w_1763 , w_1764 , w_1765 , 
		w_1766 , w_1767 , w_1768 , w_1769 , w_1770 , w_1771 , w_1772 , w_1773 , w_1774 , w_1775 , 
		w_1776 , w_1777 , w_1778 , w_1779 , w_1780 , w_1781 , w_1782 , w_1783 , w_1784 , w_1785 , 
		w_1786 , w_1787 , w_1788 , w_1789 , w_1790 , w_1791 , w_1792 , w_1793 , w_1794 , w_1795 , 
		w_1796 , w_1797 , w_1798 , w_1799 , w_1800 , w_1801 , w_1802 , w_1803 , w_1804 , w_1805 , 
		w_1806 , w_1807 , w_1808 , w_1809 , w_1810 , w_1811 , w_1812 , w_1813 , w_1814 , w_1815 , 
		w_1816 , w_1817 , w_1818 , w_1819 , w_1820 , w_1821 , w_1822 , w_1823 , w_1824 , w_1825 , 
		w_1826 , w_1827 , w_1828 , w_1829 , w_1830 , w_1831 , w_1832 , w_1833 , w_1834 , w_1835 , 
		w_1836 , w_1837 , w_1838 , w_1839 , w_1840 , w_1841 , w_1842 , w_1843 , w_1844 , w_1845 , 
		w_1846 , w_1847 , w_1848 , w_1849 , w_1850 , w_1851 , w_1852 , w_1853 , w_1854 , w_1855 , 
		w_1856 , w_1857 , w_1858 , w_1859 , w_1860 , w_1861 , w_1862 , w_1863 , w_1864 , w_1865 , 
		w_1866 , w_1867 , w_1868 , w_1869 , w_1870 , w_1871 , w_1872 , w_1873 , w_1874 , w_1875 , 
		w_1876 , w_1877 , w_1878 , w_1879 , w_1880 , w_1881 , w_1882 , w_1883 , w_1884 , w_1885 , 
		w_1886 , w_1887 , w_1888 , w_1889 , w_1890 , w_1891 , w_1892 , w_1893 , w_1894 , w_1895 , 
		w_1896 , w_1897 , w_1898 , w_1899 , w_1900 , w_1901 , w_1902 , w_1903 , w_1904 , w_1905 , 
		w_1906 , w_1907 , w_1908 , w_1909 , w_1910 , w_1911 , w_1912 , w_1913 , w_1914 , w_1915 , 
		w_1916 , w_1917 , w_1918 , w_1919 , w_1920 , w_1921 , w_1922 , w_1923 , w_1924 , w_1925 , 
		w_1926 , w_1927 , w_1928 , w_1929 , w_1930 , w_1931 , w_1932 , w_1933 , w_1934 , w_1935 , 
		w_1936 , w_1937 , w_1938 , w_1939 , w_1940 , w_1941 , w_1942 , w_1943 , w_1944 , w_1945 , 
		w_1946 , w_1947 , w_1948 , w_1949 , w_1950 , w_1951 , w_1952 , w_1953 , w_1954 , w_1955 , 
		w_1956 , w_1957 , w_1958 , w_1959 , w_1960 , w_1961 , w_1962 , w_1963 , w_1964 , w_1965 , 
		w_1966 , w_1967 , w_1968 , w_1969 , w_1970 , w_1971 , w_1972 , w_1973 , w_1974 , w_1975 , 
		w_1976 , w_1977 , w_1978 , w_1979 , w_1980 , w_1981 , w_1982 , w_1983 , w_1984 , w_1985 , 
		w_1986 , w_1987 , w_1988 , w_1989 , w_1990 , w_1991 , w_1992 , w_1993 , w_1994 , w_1995 , 
		w_1996 , w_1997 , w_1998 , w_1999 , w_2000 , w_2001 , w_2002 , w_2003 , w_2004 , w_2005 , 
		w_2006 , w_2007 , w_2008 , w_2009 , w_2010 , w_2011 , w_2012 , w_2013 , w_2014 , w_2015 , 
		w_2016 , w_2017 , w_2018 , w_2019 , w_2020 , w_2021 , w_2022 , w_2023 , w_2024 , w_2025 , 
		w_2026 , w_2027 , w_2028 , w_2029 , w_2030 , w_2031 , w_2032 , w_2033 , w_2034 , w_2035 , 
		w_2036 , w_2037 , w_2038 , w_2039 , w_2040 , w_2041 , w_2042 , w_2043 , w_2044 , w_2045 , 
		w_2046 , w_2047 , w_2048 , w_2049 , w_2050 , w_2051 , w_2052 , w_2053 , w_2054 , w_2055 , 
		w_2056 , w_2057 , w_2058 , w_2059 , w_2060 , w_2061 , w_2062 , w_2063 , w_2064 , w_2065 , 
		w_2066 , w_2067 , w_2068 , w_2069 , w_2070 , w_2071 , w_2072 , w_2073 , w_2074 , w_2075 , 
		w_2076 , w_2077 , w_2078 , w_2079 , w_2080 , w_2081 , w_2082 , w_2083 , w_2084 , w_2085 , 
		w_2086 , w_2087 , w_2088 , w_2089 , w_2090 , w_2091 , w_2092 , w_2093 , w_2094 , w_2095 , 
		w_2096 , w_2097 , w_2098 , w_2099 , w_2100 , w_2101 , w_2102 , w_2103 , w_2104 , w_2105 , 
		w_2106 , w_2107 , w_2108 , w_2109 , w_2110 , w_2111 , w_2112 , w_2113 , w_2114 , w_2115 , 
		w_2116 , w_2117 , w_2118 , w_2119 , w_2120 , w_2121 , w_2122 , w_2123 , w_2124 , w_2125 , 
		w_2126 , w_2127 , w_2128 , w_2129 , w_2130 , w_2131 , w_2132 , w_2133 , w_2134 , w_2135 , 
		w_2136 , w_2137 , w_2138 , w_2139 , w_2140 , w_2141 , w_2142 , w_2143 , w_2144 , w_2145 , 
		w_2146 , w_2147 , w_2148 , w_2149 , w_2150 , w_2151 , w_2152 , w_2153 , w_2154 , w_2155 , 
		w_2156 , w_2157 , w_2158 , w_2159 , w_2160 , w_2161 , w_2162 , w_2163 , w_2164 , w_2165 , 
		w_2166 , w_2167 , w_2168 , w_2169 , w_2170 , w_2171 , w_2172 , w_2173 , w_2174 , w_2175 , 
		w_2176 , w_2177 , w_2178 , w_2179 , w_2180 , w_2181 , w_2182 , w_2183 , w_2184 , w_2185 , 
		w_2186 , w_2187 , w_2188 , w_2189 , w_2190 , w_2191 , w_2192 , w_2193 , w_2194 , w_2195 , 
		w_2196 , w_2197 , w_2198 , w_2199 , w_2200 , w_2201 , w_2202 , w_2203 , w_2204 , w_2205 , 
		w_2206 , w_2207 , w_2208 , w_2209 , w_2210 , w_2211 , w_2212 , w_2213 , w_2214 , w_2215 , 
		w_2216 , w_2217 , w_2218 , w_2219 , w_2220 , w_2221 , w_2222 , w_2223 , w_2224 , w_2225 , 
		w_2226 , w_2227 , w_2228 , w_2229 , w_2230 , w_2231 , w_2232 , w_2233 , w_2234 , w_2235 , 
		w_2236 , w_2237 , w_2238 , w_2239 , w_2240 , w_2241 , w_2242 , w_2243 , w_2244 , w_2245 , 
		w_2246 , w_2247 , w_2248 , w_2249 , w_2250 , w_2251 , w_2252 , w_2253 , w_2254 , w_2255 , 
		w_2256 , w_2257 , w_2258 , w_2259 , w_2260 , w_2261 , w_2262 , w_2263 , w_2264 , w_2265 , 
		w_2266 , w_2267 , w_2268 , w_2269 , w_2270 , w_2271 , w_2272 , w_2273 , w_2274 , w_2275 , 
		w_2276 , w_2277 , w_2278 , w_2279 , w_2280 , w_2281 , w_2282 , w_2283 , w_2284 , w_2285 , 
		w_2286 , w_2287 , w_2288 , w_2289 , w_2290 , w_2291 , w_2292 , w_2293 , w_2294 , w_2295 , 
		w_2296 , w_2297 , w_2298 , w_2299 , w_2300 , w_2301 , w_2302 , w_2303 , w_2304 , w_2305 , 
		w_2306 , w_2307 , w_2308 , w_2309 , w_2310 , w_2311 , w_2312 , w_2313 , w_2314 , w_2315 , 
		w_2316 , w_2317 , w_2318 , w_2319 , w_2320 , w_2321 , w_2322 , w_2323 , w_2324 , w_2325 , 
		w_2326 , w_2327 , w_2328 , w_2329 , w_2330 , w_2331 , w_2332 , w_2333 , w_2334 , w_2335 , 
		w_2336 , w_2337 , w_2338 , w_2339 , w_2340 , w_2341 , w_2342 , w_2343 , w_2344 , w_2345 , 
		w_2346 , w_2347 , w_2348 , w_2349 , w_2350 , w_2351 , w_2352 , w_2353 , w_2354 , w_2355 , 
		w_2356 , w_2357 , w_2358 , w_2359 , w_2360 , w_2361 , w_2362 , w_2363 , w_2364 , w_2365 , 
		w_2366 , w_2367 , w_2368 , w_2369 , w_2370 , w_2371 , w_2372 , w_2373 , w_2374 , w_2375 , 
		w_2376 , w_2377 , w_2378 , w_2379 , w_2380 , w_2381 , w_2382 , w_2383 , w_2384 , w_2385 , 
		w_2386 , w_2387 , w_2388 , w_2389 , w_2390 , w_2391 , w_2392 , w_2393 , w_2394 , w_2395 , 
		w_2396 , w_2397 , w_2398 , w_2399 , w_2400 , w_2401 , w_2402 , w_2403 , w_2404 , w_2405 , 
		w_2406 , w_2407 , w_2408 , w_2409 , w_2410 , w_2411 , w_2412 , w_2413 , w_2414 , w_2415 , 
		w_2416 , w_2417 , w_2418 , w_2419 , w_2420 , w_2421 , w_2422 , w_2423 , w_2424 , w_2425 , 
		w_2426 , w_2427 , w_2428 , w_2429 , w_2430 , w_2431 , w_2432 , w_2433 , w_2434 , w_2435 , 
		w_2436 , w_2437 , w_2438 , w_2439 , w_2440 , w_2441 , w_2442 , w_2443 , w_2444 , w_2445 , 
		w_2446 , w_2447 , w_2448 , w_2449 , w_2450 , w_2451 , w_2452 , w_2453 , w_2454 , w_2455 , 
		w_2456 , w_2457 , w_2458 , w_2459 , w_2460 , w_2461 , w_2462 , w_2463 , w_2464 , w_2465 , 
		w_2466 , w_2467 , w_2468 , w_2469 , w_2470 , w_2471 , w_2472 , w_2473 , w_2474 , w_2475 , 
		w_2476 , w_2477 , w_2478 , w_2479 , w_2480 , w_2481 , w_2482 , w_2483 , w_2484 , w_2485 , 
		w_2486 , w_2487 , w_2488 , w_2489 , w_2490 , w_2491 , w_2492 , w_2493 , w_2494 , w_2495 , 
		w_2496 , w_2497 , w_2498 , w_2499 , w_2500 , w_2501 , w_2502 , w_2503 , w_2504 , w_2505 , 
		w_2506 , w_2507 , w_2508 , w_2509 , w_2510 , w_2511 , w_2512 , w_2513 , w_2514 , w_2515 , 
		w_2516 , w_2517 , w_2518 , w_2519 , w_2520 , w_2521 , w_2522 , w_2523 , w_2524 , w_2525 , 
		w_2526 , w_2527 , w_2528 , w_2529 , w_2530 , w_2531 , w_2532 , w_2533 , w_2534 , w_2535 , 
		w_2536 , w_2537 , w_2538 , w_2539 , w_2540 , w_2541 , w_2542 , w_2543 , w_2544 , w_2545 , 
		w_2546 , w_2547 , w_2548 , w_2549 , w_2550 , w_2551 , w_2552 , w_2553 , w_2554 , w_2555 , 
		w_2556 , w_2557 , w_2558 , w_2559 , w_2560 , w_2561 , w_2562 , w_2563 , w_2564 , w_2565 , 
		w_2566 , w_2567 , w_2568 , w_2569 , w_2570 , w_2571 , w_2572 , w_2573 , w_2574 , w_2575 , 
		w_2576 , w_2577 , w_2578 , w_2579 , w_2580 , w_2581 , w_2582 , w_2583 , w_2584 , w_2585 , 
		w_2586 , w_2587 , w_2588 , w_2589 , w_2590 , w_2591 , w_2592 , w_2593 , w_2594 , w_2595 , 
		w_2596 , w_2597 , w_2598 , w_2599 , w_2600 , w_2601 , w_2602 , w_2603 , w_2604 , w_2605 , 
		w_2606 , w_2607 , w_2608 , w_2609 , w_2610 , w_2611 , w_2612 , w_2613 , w_2614 , w_2615 , 
		w_2616 , w_2617 , w_2618 , w_2619 , w_2620 , w_2621 , w_2622 , w_2623 , w_2624 , w_2625 , 
		w_2626 , w_2627 , w_2628 , w_2629 , w_2630 , w_2631 , w_2632 , w_2633 , w_2634 , w_2635 , 
		w_2636 , w_2637 , w_2638 , w_2639 , w_2640 , w_2641 , w_2642 , w_2643 , w_2644 , w_2645 , 
		w_2646 , w_2647 , w_2648 , w_2649 , w_2650 , w_2651 , w_2652 , w_2653 , w_2654 , w_2655 , 
		w_2656 , w_2657 , w_2658 , w_2659 , w_2660 , w_2661 , w_2662 , w_2663 , w_2664 , w_2665 , 
		w_2666 , w_2667 , w_2668 , w_2669 , w_2670 , w_2671 , w_2672 , w_2673 , w_2674 , w_2675 , 
		w_2676 , w_2677 , w_2678 , w_2679 , w_2680 , w_2681 , w_2682 , w_2683 , w_2684 , w_2685 , 
		w_2686 , w_2687 , w_2688 , w_2689 , w_2690 , w_2691 , w_2692 , w_2693 , w_2694 , w_2695 , 
		w_2696 , w_2697 , w_2698 , w_2699 , w_2700 , w_2701 , w_2702 , w_2703 , w_2704 , w_2705 , 
		w_2706 , w_2707 , w_2708 , w_2709 , w_2710 , w_2711 , w_2712 , w_2713 , w_2714 , w_2715 , 
		w_2716 , w_2717 , w_2718 , w_2719 , w_2720 , w_2721 , w_2722 , w_2723 , w_2724 , w_2725 , 
		w_2726 , w_2727 , w_2728 , w_2729 , w_2730 , w_2731 , w_2732 , w_2733 , w_2734 , w_2735 , 
		w_2736 , w_2737 , w_2738 , w_2739 , w_2740 , w_2741 , w_2742 , w_2743 , w_2744 , w_2745 , 
		w_2746 , w_2747 , w_2748 , w_2749 , w_2750 , w_2751 , w_2752 , w_2753 , w_2754 , w_2755 , 
		w_2756 , w_2757 , w_2758 , w_2759 , w_2760 , w_2761 , w_2762 , w_2763 , w_2764 , w_2765 , 
		w_2766 , w_2767 , w_2768 , w_2769 , w_2770 , w_2771 , w_2772 , w_2773 , w_2774 , w_2775 , 
		w_2776 , w_2777 , w_2778 , w_2779 , w_2780 , w_2781 , w_2782 , w_2783 , w_2784 , w_2785 , 
		w_2786 , w_2787 , w_2788 , w_2789 , w_2790 , w_2791 , w_2792 , w_2793 , w_2794 , w_2795 , 
		w_2796 , w_2797 , w_2798 , w_2799 , w_2800 , w_2801 , w_2802 , w_2803 , w_2804 , w_2805 , 
		w_2806 , w_2807 , w_2808 , w_2809 , w_2810 , w_2811 , w_2812 , w_2813 , w_2814 , w_2815 , 
		w_2816 , w_2817 , w_2818 , w_2819 , w_2820 , w_2821 , w_2822 , w_2823 , w_2824 , w_2825 , 
		w_2826 , w_2827 , w_2828 , w_2829 , w_2830 , w_2831 , w_2832 , w_2833 , w_2834 , w_2835 , 
		w_2836 , w_2837 , w_2838 , w_2839 , w_2840 , w_2841 , w_2842 , w_2843 , w_2844 , w_2845 , 
		w_2846 , w_2847 , w_2848 , w_2849 , w_2850 , w_2851 , w_2852 , w_2853 , w_2854 , w_2855 , 
		w_2856 , w_2857 , w_2858 , w_2859 , w_2860 , w_2861 , w_2862 , w_2863 , w_2864 , w_2865 , 
		w_2866 , w_2867 , w_2868 , w_2869 , w_2870 , w_2871 , w_2872 , w_2873 , w_2874 , w_2875 , 
		w_2876 , w_2877 , w_2878 , w_2879 , w_2880 , w_2881 , w_2882 , w_2883 , w_2884 , w_2885 , 
		w_2886 , w_2887 , w_2888 , w_2889 , w_2890 , w_2891 , w_2892 , w_2893 , w_2894 , w_2895 , 
		w_2896 , w_2897 , w_2898 , w_2899 , w_2900 , w_2901 , w_2902 , w_2903 , w_2904 , w_2905 , 
		w_2906 , w_2907 , w_2908 , w_2909 , w_2910 , w_2911 , w_2912 , w_2913 , w_2914 , w_2915 , 
		w_2916 , w_2917 , w_2918 , w_2919 , w_2920 , w_2921 , w_2922 , w_2923 , w_2924 , w_2925 , 
		w_2926 , w_2927 , w_2928 , w_2929 , w_2930 , w_2931 , w_2932 , w_2933 , w_2934 , w_2935 , 
		w_2936 , w_2937 , w_2938 , w_2939 , w_2940 , w_2941 , w_2942 , w_2943 , w_2944 , w_2945 , 
		w_2946 , w_2947 , w_2948 , w_2949 , w_2950 , w_2951 , w_2952 , w_2953 , w_2954 , w_2955 , 
		w_2956 , w_2957 , w_2958 , w_2959 , w_2960 , w_2961 , w_2962 , w_2963 , w_2964 , w_2965 , 
		w_2966 , w_2967 , w_2968 , w_2969 , w_2970 , w_2971 , w_2972 , w_2973 , w_2974 , w_2975 , 
		w_2976 , w_2977 , w_2978 , w_2979 , w_2980 , w_2981 , w_2982 , w_2983 , w_2984 , w_2985 , 
		w_2986 , w_2987 , w_2988 , w_2989 , w_2990 , w_2991 , w_2992 , w_2993 , w_2994 , w_2995 , 
		w_2996 , w_2997 , w_2998 , w_2999 , w_3000 , w_3001 , w_3002 , w_3003 , w_3004 , w_3005 , 
		w_3006 , w_3007 , w_3008 , w_3009 , w_3010 , w_3011 , w_3012 , w_3013 , w_3014 , w_3015 , 
		w_3016 , w_3017 , w_3018 , w_3019 , w_3020 , w_3021 , w_3022 , w_3023 , w_3024 , w_3025 , 
		w_3026 , w_3027 , w_3028 , w_3029 , w_3030 , w_3031 , w_3032 , w_3033 , w_3034 , w_3035 , 
		w_3036 , w_3037 , w_3038 , w_3039 , w_3040 , w_3041 , w_3042 , w_3043 , w_3044 , w_3045 , 
		w_3046 , w_3047 , w_3048 , w_3049 , w_3050 , w_3051 , w_3052 , w_3053 , w_3054 , w_3055 , 
		w_3056 , w_3057 , w_3058 , w_3059 , w_3060 , w_3061 , w_3062 , w_3063 , w_3064 , w_3065 , 
		w_3066 , w_3067 , w_3068 , w_3069 , w_3070 , w_3071 , w_3072 , w_3073 , w_3074 , w_3075 , 
		w_3076 , w_3077 , w_3078 , w_3079 , w_3080 , w_3081 , w_3082 , w_3083 , w_3084 , w_3085 , 
		w_3086 , w_3087 , w_3088 , w_3089 , w_3090 , w_3091 , w_3092 , w_3093 , w_3094 , w_3095 , 
		w_3096 , w_3097 , w_3098 , w_3099 , w_3100 , w_3101 , w_3102 , w_3103 , w_3104 , w_3105 , 
		w_3106 , w_3107 , w_3108 , w_3109 , w_3110 , w_3111 , w_3112 , w_3113 , w_3114 , w_3115 , 
		w_3116 , w_3117 , w_3118 , w_3119 , w_3120 , w_3121 , w_3122 , w_3123 , w_3124 , w_3125 , 
		w_3126 , w_3127 , w_3128 , w_3129 , w_3130 , w_3131 , w_3132 , w_3133 , w_3134 , w_3135 , 
		w_3136 , w_3137 , w_3138 , w_3139 , w_3140 , w_3141 , w_3142 , w_3143 , w_3144 , w_3145 , 
		w_3146 , w_3147 , w_3148 , w_3149 , w_3150 , w_3151 , w_3152 , w_3153 , w_3154 , w_3155 , 
		w_3156 , w_3157 , w_3158 , w_3159 , w_3160 , w_3161 , w_3162 , w_3163 , w_3164 , w_3165 , 
		w_3166 , w_3167 , w_3168 , w_3169 , w_3170 , w_3171 , w_3172 , w_3173 , w_3174 , w_3175 , 
		w_3176 , w_3177 , w_3178 , w_3179 , w_3180 , w_3181 , w_3182 , w_3183 , w_3184 , w_3185 , 
		w_3186 , w_3187 , w_3188 , w_3189 , w_3190 , w_3191 , w_3192 , w_3193 , w_3194 , w_3195 , 
		w_3196 , w_3197 , w_3198 , w_3199 , w_3200 , w_3201 , w_3202 , w_3203 , w_3204 , w_3205 , 
		w_3206 , w_3207 , w_3208 , w_3209 , w_3210 , w_3211 , w_3212 , w_3213 , w_3214 , w_3215 , 
		w_3216 , w_3217 , w_3218 , w_3219 , w_3220 , w_3221 , w_3222 , w_3223 , w_3224 , w_3225 , 
		w_3226 , w_3227 , w_3228 , w_3229 , w_3230 , w_3231 , w_3232 , w_3233 , w_3234 , w_3235 , 
		w_3236 , w_3237 , w_3238 , w_3239 , w_3240 , w_3241 , w_3242 , w_3243 , w_3244 , w_3245 , 
		w_3246 , w_3247 , w_3248 , w_3249 , w_3250 , w_3251 , w_3252 , w_3253 , w_3254 , w_3255 , 
		w_3256 , w_3257 , w_3258 , w_3259 , w_3260 , w_3261 , w_3262 , w_3263 , w_3264 , w_3265 , 
		w_3266 , w_3267 , w_3268 , w_3269 , w_3270 , w_3271 , w_3272 , w_3273 , w_3274 , w_3275 , 
		w_3276 , w_3277 , w_3278 , w_3279 , w_3280 , w_3281 , w_3282 , w_3283 , w_3284 , w_3285 , 
		w_3286 , w_3287 , w_3288 , w_3289 ;
buf ( \O[19]_b1 , \943_b1 );
buf ( \O[19]_b0 , \943_b0 );
buf ( \O[18]_b1 , \949_b1 );
buf ( \O[18]_b0 , \949_b0 );
buf ( \O[17]_b1 , \969_b1 );
buf ( \O[17]_b0 , \969_b0 );
buf ( \O[16]_b1 , \1073_b1 );
buf ( \O[16]_b0 , \1073_b0 );
buf ( \O[15]_b1 , \985_b1 );
buf ( \O[15]_b0 , \985_b0 );
buf ( \O[14]_b1 , \1074_b1 );
buf ( \O[14]_b0 , \1074_b0 );
buf ( \O[13]_b1 , \997_b1 );
buf ( \O[13]_b0 , \997_b0 );
buf ( \O[12]_b1 , \1075_b1 );
buf ( \O[12]_b0 , \1075_b0 );
buf ( \O[11]_b1 , \1010_b1 );
buf ( \O[11]_b0 , \1010_b0 );
buf ( \O[10]_b1 , \1017_b1 );
buf ( \O[10]_b0 , \1017_b0 );
buf ( \O[9]_b1 , \1024_b1 );
buf ( \O[9]_b0 , \1024_b0 );
buf ( \O[8]_b1 , \1030_b1 );
buf ( \O[8]_b0 , \1030_b0 );
buf ( \O[7]_b1 , \1039_b1 );
buf ( \O[7]_b0 , \1039_b0 );
buf ( \O[6]_b1 , \1047_b1 );
buf ( \O[6]_b0 , \1047_b0 );
buf ( \O[5]_b1 , \1053_b1 );
buf ( \O[5]_b0 , \1053_b0 );
buf ( \O[4]_b1 , \1059_b1 );
buf ( \O[4]_b0 , \1059_b0 );
buf ( \O[3]_b1 , \1065_b1 );
buf ( \O[3]_b0 , \1065_b0 );
buf ( \O[2]_b1 , \1067_b1 );
buf ( \O[2]_b0 , \1067_b0 );
buf ( \O[1]_b1 , \1071_b1 );
buf ( \O[1]_b0 , \1071_b0 );
buf ( \O[0]_b1 , \1072_b1 );
buf ( \O[0]_b0 , \1072_b0 );
buf ( \72_b1 , \A[0][5]_b1 );
not ( \72_b1 , w_0 );
not ( \72_b0 , w_1 );
and ( w_0 , w_1 , \A[0][5]_b0 );
or ( \73_b1 , \I[1]_b1 , w_3 );
not ( w_3 , w_4 );
and ( \73_b0 , \I[1]_b0 , w_5 );
and ( w_4 ,  , w_5 );
buf ( w_3 , \I[0]_b1 );
not ( w_3 , w_6 );
not (  , w_7 );
and ( w_6 , w_7 , \I[0]_b0 );
buf ( \74_b1 , \73_b1 );
not ( \74_b1 , w_8 );
not ( \74_b0 , w_9 );
and ( w_8 , w_9 , \73_b0 );
or ( \75_b1 , \72_b1 , w_10 );
or ( \75_b0 , \72_b0 , \74_b0 );
not ( \74_b0 , w_11 );
and ( w_11 , w_10 , \74_b1 );
or ( \76_b1 , \A[1][5]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_12 );
and ( \76_b0 , \A[1][5]_b0 , w_13 );
and ( w_12 , w_13 , \I[0]_b0 );
or ( \77_b1 , \A[2][5]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_14 );
and ( \77_b0 , \A[2][5]_b0 , w_15 );
and ( w_14 , w_15 , \I[1]_b0 );
or ( \78_b1 , \76_b1 , w_17 );
not ( w_17 , w_18 );
and ( \78_b0 , \76_b0 , w_19 );
and ( w_18 ,  , w_19 );
buf ( w_17 , \77_b1 );
not ( w_17 , w_20 );
not (  , w_21 );
and ( w_20 , w_21 , \77_b0 );
or ( \79_b1 , \75_b1 , w_23 );
not ( w_23 , w_24 );
and ( \79_b0 , \75_b0 , w_25 );
and ( w_24 ,  , w_25 );
buf ( w_23 , \78_b1 );
not ( w_23 , w_26 );
not (  , w_27 );
and ( w_26 , w_27 , \78_b0 );
buf ( \80_b1 , \79_b1 );
buf ( \80_b0 , \79_b0 );
or ( \81_b1 , \80_b1 , w_29 );
not ( w_29 , w_30 );
and ( \81_b0 , \80_b0 , w_31 );
and ( w_30 ,  , w_31 );
buf ( w_29 , \B[9]_b1 );
not ( w_29 , w_32 );
not (  , w_33 );
and ( w_32 , w_33 , \B[9]_b0 );
buf ( \82_b1 , \A[0][7]_b1 );
not ( \82_b1 , w_34 );
not ( \82_b0 , w_35 );
and ( w_34 , w_35 , \A[0][7]_b0 );
or ( \84_b1 , \A[2][7]_b1 , w_37 );
not ( w_37 , w_38 );
and ( \84_b0 , \A[2][7]_b0 , w_39 );
and ( w_38 ,  , w_39 );
buf ( w_37 , \I[1]_b1 );
not ( w_37 , w_40 );
not (  , w_41 );
and ( w_40 , w_41 , \I[1]_b0 );
or ( \85_b1 , \A[1][7]_b1 , w_43 );
not ( w_43 , w_44 );
and ( \85_b0 , \A[1][7]_b0 , w_45 );
and ( w_44 ,  , w_45 );
buf ( w_43 , \I[0]_b1 );
not ( w_43 , w_46 );
not (  , w_47 );
and ( w_46 , w_47 , \I[0]_b0 );
or ( \86_b1 , \84_b1 , w_49 );
not ( w_49 , w_50 );
and ( \86_b0 , \84_b0 , w_51 );
and ( w_50 ,  , w_51 );
buf ( w_49 , \85_b1 );
not ( w_49 , w_52 );
not (  , w_53 );
and ( w_52 , w_53 , \85_b0 );
or ( \87_b1 , \83_b1 , w_55 );
not ( w_55 , w_56 );
and ( \87_b0 , \83_b0 , w_57 );
and ( w_56 ,  , w_57 );
buf ( w_55 , \86_b1 );
not ( w_55 , w_58 );
not (  , w_59 );
and ( w_58 , w_59 , \86_b0 );
buf ( \88_b1 , \87_b1 );
not ( \88_b1 , w_60 );
not ( \88_b0 , w_61 );
and ( w_60 , w_61 , \87_b0 );
or ( \89_b1 , \88_b1 , w_63 );
not ( w_63 , w_64 );
and ( \89_b0 , \88_b0 , w_65 );
and ( w_64 ,  , w_65 );
buf ( w_63 , \B[7]_b1 );
not ( w_63 , w_66 );
not (  , w_67 );
and ( w_66 , w_67 , \B[7]_b0 );
or ( \90_b1 , \81_b1 , \89_b1 );
xor ( \90_b0 , \81_b0 , w_68 );
not ( w_68 , w_69 );
and ( w_69 , \89_b1 , \89_b0 );
or ( \91_b1 , \80_b1 , w_71 );
not ( w_71 , w_72 );
and ( \91_b0 , \80_b0 , w_73 );
and ( w_72 ,  , w_73 );
buf ( w_71 , \B[8]_b1 );
not ( w_71 , w_74 );
not (  , w_75 );
and ( w_74 , w_75 , \B[8]_b0 );
or ( \92_b1 , \I[1]_b1 , w_77 );
not ( w_77 , w_78 );
and ( \92_b0 , \I[1]_b0 , w_79 );
and ( w_78 ,  , w_79 );
buf ( w_77 , \I[0]_b1 );
not ( w_77 , w_80 );
not (  , w_81 );
and ( w_80 , w_81 , \I[0]_b0 );
buf ( \93_b1 , \92_b1 );
not ( \93_b1 , w_82 );
not ( \93_b0 , w_83 );
and ( w_82 , w_83 , \92_b0 );
buf ( \94_b1 , \A[0][4]_b1 );
not ( \94_b1 , w_84 );
not ( \94_b0 , w_85 );
and ( w_84 , w_85 , \A[0][4]_b0 );
or ( \95_b1 , \93_b1 , w_86 );
or ( \95_b0 , \93_b0 , \94_b0 );
not ( \94_b0 , w_87 );
and ( w_87 , w_86 , \94_b1 );
or ( \96_b1 , \A[1][4]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_88 );
and ( \96_b0 , \A[1][4]_b0 , w_89 );
and ( w_88 , w_89 , \I[0]_b0 );
or ( \97_b1 , \A[2][4]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_90 );
and ( \97_b0 , \A[2][4]_b0 , w_91 );
and ( w_90 , w_91 , \I[1]_b0 );
or ( \98_b1 , \96_b1 , w_93 );
not ( w_93 , w_94 );
and ( \98_b0 , \96_b0 , w_95 );
and ( w_94 ,  , w_95 );
buf ( w_93 , \97_b1 );
not ( w_93 , w_96 );
not (  , w_97 );
and ( w_96 , w_97 , \97_b0 );
or ( \99_b1 , \95_b1 , w_99 );
not ( w_99 , w_100 );
and ( \99_b0 , \95_b0 , w_101 );
and ( w_100 ,  , w_101 );
buf ( w_99 , \98_b1 );
not ( w_99 , w_102 );
not (  , w_103 );
and ( w_102 , w_103 , \98_b0 );
buf ( \100_b1 , \99_b1 );
buf ( \100_b0 , \99_b0 );
or ( \101_b1 , \100_b1 , w_105 );
not ( w_105 , w_106 );
and ( \101_b0 , \100_b0 , w_107 );
and ( w_106 ,  , w_107 );
buf ( w_105 , \B[9]_b1 );
not ( w_105 , w_108 );
not (  , w_109 );
and ( w_108 , w_109 , \B[9]_b0 );
or ( \102_b1 , \91_b1 , \101_b1 );
xor ( \102_b0 , \91_b0 , w_110 );
not ( w_110 , w_111 );
and ( w_111 , \101_b1 , \101_b0 );
or ( \103_b1 , \88_b1 , w_113 );
not ( w_113 , w_114 );
and ( \103_b0 , \88_b0 , w_115 );
and ( w_114 ,  , w_115 );
buf ( w_113 , \B[6]_b1 );
not ( w_113 , w_116 );
not (  , w_117 );
and ( w_116 , w_117 , \B[6]_b0 );
or ( \104_b1 , \102_b1 , \103_b1 );
not ( \103_b1 , w_118 );
and ( \104_b0 , \102_b0 , w_119 );
and ( w_118 , w_119 , \103_b0 );
or ( \105_b1 , \91_b1 , \101_b1 );
not ( \101_b1 , w_120 );
and ( \105_b0 , \91_b0 , w_121 );
and ( w_120 , w_121 , \101_b0 );
or ( \106_b1 , \104_b1 , w_122 );
or ( \106_b0 , \104_b0 , \105_b0 );
not ( \105_b0 , w_123 );
and ( w_123 , w_122 , \105_b1 );
or ( \107_b1 , \90_b1 , \106_b1 );
not ( \106_b1 , w_124 );
and ( \107_b0 , \90_b0 , w_125 );
and ( w_124 , w_125 , \106_b0 );
or ( \108_b1 , \81_b1 , \89_b1 );
not ( \89_b1 , w_126 );
and ( \108_b0 , \81_b0 , w_127 );
and ( w_126 , w_127 , \89_b0 );
or ( \109_b1 , \107_b1 , w_128 );
or ( \109_b0 , \107_b0 , \108_b0 );
not ( \108_b0 , w_129 );
and ( w_129 , w_128 , \108_b1 );
or ( \110_b1 , \88_b1 , w_131 );
not ( w_131 , w_132 );
and ( \110_b0 , \88_b0 , w_133 );
and ( w_132 ,  , w_133 );
buf ( w_131 , \B[8]_b1 );
not ( w_131 , w_134 );
not (  , w_135 );
and ( w_134 , w_135 , \B[8]_b0 );
or ( \111_b1 , \I[1]_b1 , w_137 );
not ( w_137 , w_138 );
and ( \111_b0 , \I[1]_b0 , w_139 );
and ( w_138 ,  , w_139 );
buf ( w_137 , \I[0]_b1 );
not ( w_137 , w_140 );
not (  , w_141 );
and ( w_140 , w_141 , \I[0]_b0 );
buf ( \112_b1 , \111_b1 );
not ( \112_b1 , w_142 );
not ( \112_b0 , w_143 );
and ( w_142 , w_143 , \111_b0 );
buf ( \113_b1 , \A[0][6]_b1 );
not ( \113_b1 , w_144 );
not ( \113_b0 , w_145 );
and ( w_144 , w_145 , \A[0][6]_b0 );
or ( \114_b1 , \112_b1 , w_146 );
or ( \114_b0 , \112_b0 , \113_b0 );
not ( \113_b0 , w_147 );
and ( w_147 , w_146 , \113_b1 );
or ( \115_b1 , \A[1][6]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_148 );
and ( \115_b0 , \A[1][6]_b0 , w_149 );
and ( w_148 , w_149 , \I[0]_b0 );
or ( \116_b1 , \A[2][6]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_150 );
and ( \116_b0 , \A[2][6]_b0 , w_151 );
and ( w_150 , w_151 , \I[1]_b0 );
or ( \117_b1 , \115_b1 , w_153 );
not ( w_153 , w_154 );
and ( \117_b0 , \115_b0 , w_155 );
and ( w_154 ,  , w_155 );
buf ( w_153 , \116_b1 );
not ( w_153 , w_156 );
not (  , w_157 );
and ( w_156 , w_157 , \116_b0 );
or ( \118_b1 , \114_b1 , w_159 );
not ( w_159 , w_160 );
and ( \118_b0 , \114_b0 , w_161 );
and ( w_160 ,  , w_161 );
buf ( w_159 , \117_b1 );
not ( w_159 , w_162 );
not (  , w_163 );
and ( w_162 , w_163 , \117_b0 );
buf ( \119_b1 , \118_b1 );
buf ( \119_b0 , \118_b0 );
or ( \120_b1 , \119_b1 , w_165 );
not ( w_165 , w_166 );
and ( \120_b0 , \119_b0 , w_167 );
and ( w_166 ,  , w_167 );
buf ( w_165 , \B[8]_b1 );
not ( w_165 , w_168 );
not (  , w_169 );
and ( w_168 , w_169 , \B[8]_b0 );
or ( \121_b1 , \I[1]_b1 , w_171 );
not ( w_171 , w_172 );
and ( \121_b0 , \I[1]_b0 , w_173 );
and ( w_172 ,  , w_173 );
buf ( w_171 , \I[0]_b1 );
not ( w_171 , w_174 );
not (  , w_175 );
and ( w_174 , w_175 , \I[0]_b0 );
buf ( \122_b1 , \121_b1 );
not ( \122_b1 , w_176 );
not ( \122_b0 , w_177 );
and ( w_176 , w_177 , \121_b0 );
buf ( \123_b1 , \A[0][9]_b1 );
not ( \123_b1 , w_178 );
not ( \123_b0 , w_179 );
and ( w_178 , w_179 , \A[0][9]_b0 );
or ( \124_b1 , \122_b1 , w_180 );
or ( \124_b0 , \122_b0 , \123_b0 );
not ( \123_b0 , w_181 );
and ( w_181 , w_180 , \123_b1 );
or ( \125_b1 , \A[1][9]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_182 );
and ( \125_b0 , \A[1][9]_b0 , w_183 );
and ( w_182 , w_183 , \I[0]_b0 );
or ( \126_b1 , \A[2][9]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_184 );
and ( \126_b0 , \A[2][9]_b0 , w_185 );
and ( w_184 , w_185 , \I[1]_b0 );
or ( \127_b1 , \125_b1 , w_187 );
not ( w_187 , w_188 );
and ( \127_b0 , \125_b0 , w_189 );
and ( w_188 ,  , w_189 );
buf ( w_187 , \126_b1 );
not ( w_187 , w_190 );
not (  , w_191 );
and ( w_190 , w_191 , \126_b0 );
or ( \128_b1 , \124_b1 , w_193 );
not ( w_193 , w_194 );
and ( \128_b0 , \124_b0 , w_195 );
and ( w_194 ,  , w_195 );
buf ( w_193 , \127_b1 );
not ( w_193 , w_196 );
not (  , w_197 );
and ( w_196 , w_197 , \127_b0 );
buf ( \129_b1 , \128_b1 );
buf ( \129_b0 , \128_b0 );
or ( \130_b1 , \129_b1 , w_199 );
not ( w_199 , w_200 );
and ( \130_b0 , \129_b0 , w_201 );
and ( w_200 ,  , w_201 );
buf ( w_199 , \B[5]_b1 );
not ( w_199 , w_202 );
not (  , w_203 );
and ( w_202 , w_203 , \B[5]_b0 );
or ( \131_b1 , \120_b1 , \130_b1 );
xor ( \131_b0 , \120_b0 , w_204 );
not ( w_204 , w_205 );
and ( w_205 , \130_b1 , \130_b0 );
or ( \132_b1 , \I[1]_b1 , w_207 );
not ( w_207 , w_208 );
and ( \132_b0 , \I[1]_b0 , w_209 );
and ( w_208 ,  , w_209 );
buf ( w_207 , \I[0]_b1 );
not ( w_207 , w_210 );
not (  , w_211 );
and ( w_210 , w_211 , \I[0]_b0 );
buf ( \133_b1 , \132_b1 );
not ( \133_b1 , w_212 );
not ( \133_b0 , w_213 );
and ( w_212 , w_213 , \132_b0 );
buf ( \134_b1 , \A[0][8]_b1 );
not ( \134_b1 , w_214 );
not ( \134_b0 , w_215 );
and ( w_214 , w_215 , \A[0][8]_b0 );
or ( \135_b1 , \133_b1 , w_216 );
or ( \135_b0 , \133_b0 , \134_b0 );
not ( \134_b0 , w_217 );
and ( w_217 , w_216 , \134_b1 );
or ( \136_b1 , \A[1][8]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_218 );
and ( \136_b0 , \A[1][8]_b0 , w_219 );
and ( w_218 , w_219 , \I[0]_b0 );
or ( \137_b1 , \A[2][8]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_220 );
and ( \137_b0 , \A[2][8]_b0 , w_221 );
and ( w_220 , w_221 , \I[1]_b0 );
or ( \138_b1 , \136_b1 , w_223 );
not ( w_223 , w_224 );
and ( \138_b0 , \136_b0 , w_225 );
and ( w_224 ,  , w_225 );
buf ( w_223 , \137_b1 );
not ( w_223 , w_226 );
not (  , w_227 );
and ( w_226 , w_227 , \137_b0 );
or ( \139_b1 , \135_b1 , w_229 );
not ( w_229 , w_230 );
and ( \139_b0 , \135_b0 , w_231 );
and ( w_230 ,  , w_231 );
buf ( w_229 , \138_b1 );
not ( w_229 , w_232 );
not (  , w_233 );
and ( w_232 , w_233 , \138_b0 );
buf ( \140_b1 , \139_b1 );
buf ( \140_b0 , \139_b0 );
or ( \141_b1 , \140_b1 , w_235 );
not ( w_235 , w_236 );
and ( \141_b0 , \140_b0 , w_237 );
and ( w_236 ,  , w_237 );
buf ( w_235 , \B[6]_b1 );
not ( w_235 , w_238 );
not (  , w_239 );
and ( w_238 , w_239 , \B[6]_b0 );
or ( \142_b1 , \131_b1 , \141_b1 );
not ( \141_b1 , w_240 );
and ( \142_b0 , \131_b0 , w_241 );
and ( w_240 , w_241 , \141_b0 );
or ( \143_b1 , \120_b1 , \130_b1 );
not ( \130_b1 , w_242 );
and ( \143_b0 , \120_b0 , w_243 );
and ( w_242 , w_243 , \130_b0 );
or ( \144_b1 , \142_b1 , w_244 );
or ( \144_b0 , \142_b0 , \143_b0 );
not ( \143_b0 , w_245 );
and ( w_245 , w_244 , \143_b1 );
or ( \145_b1 , \110_b1 , \144_b1 );
xor ( \145_b0 , \110_b0 , w_246 );
not ( w_246 , w_247 );
and ( w_247 , \144_b1 , \144_b0 );
or ( \146_b1 , \140_b1 , w_249 );
not ( w_249 , w_250 );
and ( \146_b0 , \140_b0 , w_251 );
and ( w_250 ,  , w_251 );
buf ( w_249 , \B[7]_b1 );
not ( w_249 , w_252 );
not (  , w_253 );
and ( w_252 , w_253 , \B[7]_b0 );
or ( \147_b1 , \129_b1 , w_255 );
not ( w_255 , w_256 );
and ( \147_b0 , \129_b0 , w_257 );
and ( w_256 ,  , w_257 );
buf ( w_255 , \B[6]_b1 );
not ( w_255 , w_258 );
not (  , w_259 );
and ( w_258 , w_259 , \B[6]_b0 );
or ( \148_b1 , \146_b1 , \147_b1 );
xor ( \148_b0 , \146_b0 , w_260 );
not ( w_260 , w_261 );
and ( w_261 , \147_b1 , \147_b0 );
or ( \149_b1 , \119_b1 , w_263 );
not ( w_263 , w_264 );
and ( \149_b0 , \119_b0 , w_265 );
and ( w_264 ,  , w_265 );
buf ( w_263 , \B[9]_b1 );
not ( w_263 , w_266 );
not (  , w_267 );
and ( w_266 , w_267 , \B[9]_b0 );
or ( \150_b1 , \148_b1 , \149_b1 );
xor ( \150_b0 , \148_b0 , w_268 );
not ( w_268 , w_269 );
and ( w_269 , \149_b1 , \149_b0 );
or ( \151_b1 , \145_b1 , \150_b1 );
xor ( \151_b0 , \145_b0 , w_270 );
not ( w_270 , w_271 );
and ( w_271 , \150_b1 , \150_b0 );
or ( \152_b1 , \109_b1 , \151_b1 );
xor ( \152_b0 , \109_b0 , w_272 );
not ( w_272 , w_273 );
and ( w_273 , \151_b1 , \151_b0 );
or ( \153_b1 , \81_b1 , \89_b1 );
xor ( \153_b0 , \81_b0 , w_274 );
not ( w_274 , w_275 );
and ( w_275 , \89_b1 , \89_b0 );
or ( \154_b1 , \153_b1 , \106_b1 );
xor ( \154_b0 , \153_b0 , w_276 );
not ( w_276 , w_277 );
and ( w_277 , \106_b1 , \106_b0 );
or ( \155_b1 , \120_b1 , \130_b1 );
xor ( \155_b0 , \120_b0 , w_278 );
not ( w_278 , w_279 );
and ( w_279 , \130_b1 , \130_b0 );
or ( \156_b1 , \155_b1 , \141_b1 );
xor ( \156_b0 , \155_b0 , w_280 );
not ( w_280 , w_281 );
and ( w_281 , \141_b1 , \141_b0 );
or ( \157_b1 , \154_b1 , w_283 );
not ( w_283 , w_284 );
and ( \157_b0 , \154_b0 , w_285 );
and ( w_284 ,  , w_285 );
buf ( w_283 , \156_b1 );
not ( w_283 , w_286 );
not (  , w_287 );
and ( w_286 , w_287 , \156_b0 );
or ( \158_b1 , \140_b1 , w_289 );
not ( w_289 , w_290 );
and ( \158_b0 , \140_b0 , w_291 );
and ( w_290 ,  , w_291 );
buf ( w_289 , \B[5]_b1 );
not ( w_289 , w_292 );
not (  , w_293 );
and ( w_292 , w_293 , \B[5]_b0 );
or ( \159_b1 , \129_b1 , w_295 );
not ( w_295 , w_296 );
and ( \159_b0 , \129_b0 , w_297 );
and ( w_296 ,  , w_297 );
buf ( w_295 , \B[4]_b1 );
not ( w_295 , w_298 );
not (  , w_299 );
and ( w_298 , w_299 , \B[4]_b0 );
or ( \160_b1 , \158_b1 , \159_b1 );
xor ( \160_b0 , \158_b0 , w_300 );
not ( w_300 , w_301 );
and ( w_301 , \159_b1 , \159_b0 );
or ( \161_b1 , \119_b1 , w_303 );
not ( w_303 , w_304 );
and ( \161_b0 , \119_b0 , w_305 );
and ( w_304 ,  , w_305 );
buf ( w_303 , \B[7]_b1 );
not ( w_303 , w_306 );
not (  , w_307 );
and ( w_306 , w_307 , \B[7]_b0 );
or ( \162_b1 , \160_b1 , \161_b1 );
not ( \161_b1 , w_308 );
and ( \162_b0 , \160_b0 , w_309 );
and ( w_308 , w_309 , \161_b0 );
or ( \163_b1 , \158_b1 , \159_b1 );
not ( \159_b1 , w_310 );
and ( \163_b0 , \158_b0 , w_311 );
and ( w_310 , w_311 , \159_b0 );
or ( \164_b1 , \162_b1 , w_312 );
or ( \164_b0 , \162_b0 , \163_b0 );
not ( \163_b0 , w_313 );
and ( w_313 , w_312 , \163_b1 );
buf ( \165_b1 , \164_b1 );
not ( \165_b1 , w_314 );
not ( \165_b0 , w_315 );
and ( w_314 , w_315 , \164_b0 );
or ( \166_b1 , \157_b1 , \165_b1 );
not ( \165_b1 , w_316 );
and ( \166_b0 , \157_b0 , w_317 );
and ( w_316 , w_317 , \165_b0 );
or ( \167_b1 , \154_b1 , w_319 );
not ( w_319 , w_320 );
and ( \167_b0 , \154_b0 , w_321 );
and ( w_320 ,  , w_321 );
buf ( w_319 , \156_b1 );
not ( w_319 , w_322 );
not (  , w_323 );
and ( w_322 , w_323 , \156_b0 );
or ( \168_b1 , \166_b1 , w_325 );
not ( w_325 , w_326 );
and ( \168_b0 , \166_b0 , w_327 );
and ( w_326 ,  , w_327 );
buf ( w_325 , \167_b1 );
not ( w_325 , w_328 );
not (  , w_329 );
and ( w_328 , w_329 , \167_b0 );
or ( \169_b1 , \152_b1 , \168_b1 );
xor ( \169_b0 , \152_b0 , w_330 );
not ( w_330 , w_331 );
and ( w_331 , \168_b1 , \168_b0 );
buf ( \170_b1 , \169_b1 );
not ( \170_b1 , w_332 );
not ( \170_b0 , w_333 );
and ( w_332 , w_333 , \169_b0 );
or ( \171_b1 , \158_b1 , \159_b1 );
xor ( \171_b0 , \158_b0 , w_334 );
not ( w_334 , w_335 );
and ( w_335 , \159_b1 , \159_b0 );
or ( \172_b1 , \171_b1 , \161_b1 );
xor ( \172_b0 , \171_b0 , w_336 );
not ( w_336 , w_337 );
and ( w_337 , \161_b1 , \161_b0 );
or ( \173_b1 , \139_b1 , w_339 );
not ( w_339 , w_340 );
and ( \173_b0 , \139_b0 , w_341 );
and ( w_340 ,  , w_341 );
buf ( w_339 , \B[4]_b1 );
not ( w_339 , w_342 );
not (  , w_343 );
and ( w_342 , w_343 , \B[4]_b0 );
buf ( \174_b1 , \173_b1 );
not ( \174_b1 , w_344 );
not ( \174_b0 , w_345 );
and ( w_344 , w_345 , \173_b0 );
or ( \175_b1 , \129_b1 , w_347 );
not ( w_347 , w_348 );
and ( \175_b0 , \129_b0 , w_349 );
and ( w_348 ,  , w_349 );
buf ( w_347 , \B[3]_b1 );
not ( w_347 , w_350 );
not (  , w_351 );
and ( w_350 , w_351 , \B[3]_b0 );
buf ( \176_b1 , \175_b1 );
not ( \176_b1 , w_352 );
not ( \176_b0 , w_353 );
and ( w_352 , w_353 , \175_b0 );
or ( \177_b1 , \174_b1 , w_354 );
or ( \177_b0 , \174_b0 , \176_b0 );
not ( \176_b0 , w_355 );
and ( w_355 , w_354 , \176_b1 );
or ( \178_b1 , \119_b1 , \B[6]_b1 );
not ( \B[6]_b1 , w_356 );
and ( \178_b0 , \119_b0 , w_357 );
and ( w_356 , w_357 , \B[6]_b0 );
or ( \179_b1 , \177_b1 , w_359 );
not ( w_359 , w_360 );
and ( \179_b0 , \177_b0 , w_361 );
and ( w_360 ,  , w_361 );
buf ( w_359 , \178_b1 );
not ( w_359 , w_362 );
not (  , w_363 );
and ( w_362 , w_363 , \178_b0 );
buf ( \180_b1 , \175_b1 );
not ( \180_b1 , w_364 );
not ( \180_b0 , w_365 );
and ( w_364 , w_365 , \175_b0 );
buf ( \181_b1 , \173_b1 );
not ( \181_b1 , w_366 );
not ( \181_b0 , w_367 );
and ( w_366 , w_367 , \173_b0 );
or ( \182_b1 , \180_b1 , w_369 );
not ( w_369 , w_370 );
and ( \182_b0 , \180_b0 , w_371 );
and ( w_370 ,  , w_371 );
buf ( w_369 , \181_b1 );
not ( w_369 , w_372 );
not (  , w_373 );
and ( w_372 , w_373 , \181_b0 );
or ( \183_b1 , \179_b1 , w_375 );
not ( w_375 , w_376 );
and ( \183_b0 , \179_b0 , w_377 );
and ( w_376 ,  , w_377 );
buf ( w_375 , \182_b1 );
not ( w_375 , w_378 );
not (  , w_379 );
and ( w_378 , w_379 , \182_b0 );
buf ( \184_b1 , \183_b1 );
not ( \184_b1 , w_380 );
not ( \184_b0 , w_381 );
and ( w_380 , w_381 , \183_b0 );
or ( \185_b1 , \172_b1 , w_383 );
not ( w_383 , w_384 );
and ( \185_b0 , \172_b0 , w_385 );
and ( w_384 ,  , w_385 );
buf ( w_383 , \184_b1 );
not ( w_383 , w_386 );
not (  , w_387 );
and ( w_386 , w_387 , \184_b0 );
buf ( \186_b1 , \185_b1 );
not ( \186_b1 , w_388 );
not ( \186_b0 , w_389 );
and ( w_388 , w_389 , \185_b0 );
or ( \187_b1 , \80_b1 , w_391 );
not ( w_391 , w_392 );
and ( \187_b0 , \80_b0 , w_393 );
and ( w_392 ,  , w_393 );
buf ( w_391 , \B[7]_b1 );
not ( w_391 , w_394 );
not (  , w_395 );
and ( w_394 , w_395 , \B[7]_b0 );
or ( \188_b1 , \88_b1 , w_397 );
not ( w_397 , w_398 );
and ( \188_b0 , \88_b0 , w_399 );
and ( w_398 ,  , w_399 );
buf ( w_397 , \B[5]_b1 );
not ( w_397 , w_400 );
not (  , w_401 );
and ( w_400 , w_401 , \B[5]_b0 );
or ( \189_b1 , \187_b1 , \188_b1 );
not ( \188_b1 , w_402 );
and ( \189_b0 , \187_b0 , w_403 );
and ( w_402 , w_403 , \188_b0 );
or ( \190_b1 , \100_b1 , w_405 );
not ( w_405 , w_406 );
and ( \190_b0 , \100_b0 , w_407 );
and ( w_406 ,  , w_407 );
buf ( w_405 , \B[8]_b1 );
not ( w_405 , w_408 );
not (  , w_409 );
and ( w_408 , w_409 , \B[8]_b0 );
or ( \191_b1 , \189_b1 , w_410 );
or ( \191_b0 , \189_b0 , \190_b0 );
not ( \190_b0 , w_411 );
and ( w_411 , w_410 , \190_b1 );
or ( \192_b1 , \188_b1 , w_412 );
or ( \192_b0 , \188_b0 , \187_b0 );
not ( \187_b0 , w_413 );
and ( w_413 , w_412 , \187_b1 );
or ( \193_b1 , \191_b1 , w_415 );
not ( w_415 , w_416 );
and ( \193_b0 , \191_b0 , w_417 );
and ( w_416 ,  , w_417 );
buf ( w_415 , \192_b1 );
not ( w_415 , w_418 );
not (  , w_419 );
and ( w_418 , w_419 , \192_b0 );
buf ( \194_b1 , \193_b1 );
not ( \194_b1 , w_420 );
not ( \194_b0 , w_421 );
and ( w_420 , w_421 , \193_b0 );
or ( \195_b1 , \186_b1 , w_422 );
or ( \195_b0 , \186_b0 , \194_b0 );
not ( \194_b0 , w_423 );
and ( w_423 , w_422 , \194_b1 );
or ( \196_b1 , \172_b1 , w_424 );
or ( \196_b0 , \172_b0 , \184_b0 );
not ( \184_b0 , w_425 );
and ( w_425 , w_424 , \184_b1 );
or ( \197_b1 , \195_b1 , w_427 );
not ( w_427 , w_428 );
and ( \197_b0 , \195_b0 , w_429 );
and ( w_428 ,  , w_429 );
buf ( w_427 , \196_b1 );
not ( w_427 , w_430 );
not (  , w_431 );
and ( w_430 , w_431 , \196_b0 );
or ( \198_b1 , \156_b1 , \164_b1 );
not ( \164_b1 , w_432 );
and ( \198_b0 , \156_b0 , w_433 );
and ( w_432 , w_433 , \164_b0 );
buf ( \199_b1 , \156_b1 );
not ( \199_b1 , w_434 );
not ( \199_b0 , w_435 );
and ( w_434 , w_435 , \156_b0 );
or ( \200_b1 , \199_b1 , \165_b1 );
not ( \165_b1 , w_436 );
and ( \200_b0 , \199_b0 , w_437 );
and ( w_436 , w_437 , \165_b0 );
or ( \201_b1 , \198_b1 , w_439 );
not ( w_439 , w_440 );
and ( \201_b0 , \198_b0 , w_441 );
and ( w_440 ,  , w_441 );
buf ( w_439 , \200_b1 );
not ( w_439 , w_442 );
not (  , w_443 );
and ( w_442 , w_443 , \200_b0 );
or ( \202_b1 , \201_b1 , \154_b1 );
not ( \154_b1 , w_444 );
and ( \202_b0 , \201_b0 , w_445 );
and ( w_444 , w_445 , \154_b0 );
buf ( \203_b1 , \201_b1 );
not ( \203_b1 , w_446 );
not ( \203_b0 , w_447 );
and ( w_446 , w_447 , \201_b0 );
buf ( \204_b1 , \154_b1 );
not ( \204_b1 , w_448 );
not ( \204_b0 , w_449 );
and ( w_448 , w_449 , \154_b0 );
or ( \205_b1 , \203_b1 , \204_b1 );
not ( \204_b1 , w_450 );
and ( \205_b0 , \203_b0 , w_451 );
and ( w_450 , w_451 , \204_b0 );
or ( \206_b1 , \202_b1 , w_452 );
or ( \206_b0 , \202_b0 , \205_b0 );
not ( \205_b0 , w_453 );
and ( w_453 , w_452 , \205_b1 );
or ( \207_b1 , \197_b1 , \206_b1 );
xor ( \207_b0 , \197_b0 , w_454 );
not ( w_454 , w_455 );
and ( w_455 , \206_b1 , \206_b0 );
or ( \208_b1 , \91_b1 , \101_b1 );
xor ( \208_b0 , \91_b0 , w_456 );
not ( w_456 , w_457 );
and ( w_457 , \101_b1 , \101_b0 );
or ( \209_b1 , \208_b1 , \103_b1 );
xor ( \209_b0 , \208_b0 , w_458 );
not ( w_458 , w_459 );
and ( w_459 , \103_b1 , \103_b0 );
buf ( \210_b1 , \209_b1 );
not ( \210_b1 , w_460 );
not ( \210_b0 , w_461 );
and ( w_460 , w_461 , \209_b0 );
buf ( \211_b1 , \183_b1 );
not ( \211_b1 , w_462 );
not ( \211_b0 , w_463 );
and ( w_462 , w_463 , \183_b0 );
buf ( \212_b1 , \211_b1 );
not ( \212_b1 , w_464 );
not ( \212_b0 , w_465 );
and ( w_464 , w_465 , \211_b0 );
buf ( \213_b1 , \193_b1 );
not ( \213_b1 , w_466 );
not ( \213_b0 , w_467 );
and ( w_466 , w_467 , \193_b0 );
or ( \214_b1 , \212_b1 , \213_b1 );
not ( \213_b1 , w_468 );
and ( \214_b0 , \212_b0 , w_469 );
and ( w_468 , w_469 , \213_b0 );
or ( \215_b1 , \193_b1 , \184_b1 );
not ( \184_b1 , w_470 );
and ( \215_b0 , \193_b0 , w_471 );
and ( w_470 , w_471 , \184_b0 );
or ( \216_b1 , \214_b1 , w_473 );
not ( w_473 , w_474 );
and ( \216_b0 , \214_b0 , w_475 );
and ( w_474 ,  , w_475 );
buf ( w_473 , \215_b1 );
not ( w_473 , w_476 );
not (  , w_477 );
and ( w_476 , w_477 , \215_b0 );
buf ( \217_b1 , \216_b1 );
not ( \217_b1 , w_478 );
not ( \217_b0 , w_479 );
and ( w_478 , w_479 , \216_b0 );
buf ( \218_b1 , \172_b1 );
not ( \218_b1 , w_480 );
not ( \218_b0 , w_481 );
and ( w_480 , w_481 , \172_b0 );
buf ( \219_b1 , \218_b1 );
not ( \219_b1 , w_482 );
not ( \219_b0 , w_483 );
and ( w_482 , w_483 , \218_b0 );
or ( \220_b1 , \217_b1 , w_484 );
or ( \220_b0 , \217_b0 , \219_b0 );
not ( \219_b0 , w_485 );
and ( w_485 , w_484 , \219_b1 );
buf ( \221_b1 , \216_b1 );
not ( \221_b1 , w_486 );
not ( \221_b0 , w_487 );
and ( w_486 , w_487 , \216_b0 );
or ( \222_b1 , \221_b1 , w_489 );
not ( w_489 , w_490 );
and ( \222_b0 , \221_b0 , w_491 );
and ( w_490 ,  , w_491 );
buf ( w_489 , \172_b1 );
not ( w_489 , w_492 );
not (  , w_493 );
and ( w_492 , w_493 , \172_b0 );
or ( \223_b1 , \220_b1 , w_495 );
not ( w_495 , w_496 );
and ( \223_b0 , \220_b0 , w_497 );
and ( w_496 ,  , w_497 );
buf ( w_495 , \222_b1 );
not ( w_495 , w_498 );
not (  , w_499 );
and ( w_498 , w_499 , \222_b0 );
buf ( \224_b1 , \223_b1 );
not ( \224_b1 , w_500 );
not ( \224_b0 , w_501 );
and ( w_500 , w_501 , \223_b0 );
buf ( \225_b1 , \224_b1 );
not ( \225_b1 , w_502 );
not ( \225_b0 , w_503 );
and ( w_502 , w_503 , \224_b0 );
or ( \226_b1 , \210_b1 , w_504 );
or ( \226_b0 , \210_b0 , \225_b0 );
not ( \225_b0 , w_505 );
and ( w_505 , w_504 , \225_b1 );
buf ( \227_b1 , \A[0][3]_b1 );
not ( \227_b1 , w_506 );
not ( \227_b0 , w_507 );
and ( w_506 , w_507 , \A[0][3]_b0 );
or ( \229_b1 , \A[2][3]_b1 , w_509 );
not ( w_509 , w_510 );
and ( \229_b0 , \A[2][3]_b0 , w_511 );
and ( w_510 ,  , w_511 );
buf ( w_509 , \I[1]_b1 );
not ( w_509 , w_512 );
not (  , w_513 );
and ( w_512 , w_513 , \I[1]_b0 );
or ( \230_b1 , \A[1][3]_b1 , w_515 );
not ( w_515 , w_516 );
and ( \230_b0 , \A[1][3]_b0 , w_517 );
and ( w_516 ,  , w_517 );
buf ( w_515 , \I[0]_b1 );
not ( w_515 , w_518 );
not (  , w_519 );
and ( w_518 , w_519 , \I[0]_b0 );
or ( \231_b1 , \229_b1 , w_521 );
not ( w_521 , w_522 );
and ( \231_b0 , \229_b0 , w_523 );
and ( w_522 ,  , w_523 );
buf ( w_521 , \230_b1 );
not ( w_521 , w_524 );
not (  , w_525 );
and ( w_524 , w_525 , \230_b0 );
or ( \232_b1 , \228_b1 , w_527 );
not ( w_527 , w_528 );
and ( \232_b0 , \228_b0 , w_529 );
and ( w_528 ,  , w_529 );
buf ( w_527 , \231_b1 );
not ( w_527 , w_530 );
not (  , w_531 );
and ( w_530 , w_531 , \231_b0 );
buf ( \233_b1 , \232_b1 );
not ( \233_b1 , w_532 );
not ( \233_b0 , w_533 );
and ( w_532 , w_533 , \232_b0 );
buf ( \234_b1 , \233_b1 );
buf ( \234_b0 , \233_b0 );
or ( \235_b1 , \234_b1 , w_535 );
not ( w_535 , w_536 );
and ( \235_b0 , \234_b0 , w_537 );
and ( w_536 ,  , w_537 );
buf ( w_535 , \B[9]_b1 );
not ( w_535 , w_538 );
not (  , w_539 );
and ( w_538 , w_539 , \B[9]_b0 );
or ( \236_b1 , \139_b1 , w_541 );
not ( w_541 , w_542 );
and ( \236_b0 , \139_b0 , w_543 );
and ( w_542 ,  , w_543 );
buf ( w_541 , \B[3]_b1 );
not ( w_541 , w_544 );
not (  , w_545 );
and ( w_544 , w_545 , \B[3]_b0 );
or ( \237_b1 , \119_b1 , w_547 );
not ( w_547 , w_548 );
and ( \237_b0 , \119_b0 , w_549 );
and ( w_548 ,  , w_549 );
buf ( w_547 , \B[5]_b1 );
not ( w_547 , w_550 );
not (  , w_551 );
and ( w_550 , w_551 , \B[5]_b0 );
or ( \238_b1 , \236_b1 , \237_b1 );
xor ( \238_b0 , \236_b0 , w_552 );
not ( w_552 , w_553 );
and ( w_553 , \237_b1 , \237_b0 );
or ( \239_b1 , \129_b1 , w_555 );
not ( w_555 , w_556 );
and ( \239_b0 , \129_b0 , w_557 );
and ( w_556 ,  , w_557 );
buf ( w_555 , \B[2]_b1 );
not ( w_555 , w_558 );
not (  , w_559 );
and ( w_558 , w_559 , \B[2]_b0 );
or ( \240_b1 , \238_b1 , \239_b1 );
not ( \239_b1 , w_560 );
and ( \240_b0 , \238_b0 , w_561 );
and ( w_560 , w_561 , \239_b0 );
or ( \241_b1 , \236_b1 , \237_b1 );
not ( \237_b1 , w_562 );
and ( \241_b0 , \236_b0 , w_563 );
and ( w_562 , w_563 , \237_b0 );
or ( \242_b1 , \240_b1 , w_564 );
or ( \242_b0 , \240_b0 , \241_b0 );
not ( \241_b0 , w_565 );
and ( w_565 , w_564 , \241_b1 );
or ( \243_b1 , \235_b1 , \242_b1 );
xor ( \243_b0 , \235_b0 , w_566 );
not ( w_566 , w_567 );
and ( w_567 , \242_b1 , \242_b0 );
or ( \244_b1 , \80_b1 , w_569 );
not ( w_569 , w_570 );
and ( \244_b0 , \80_b0 , w_571 );
and ( w_570 ,  , w_571 );
buf ( w_569 , \B[6]_b1 );
not ( w_569 , w_572 );
not (  , w_573 );
and ( w_572 , w_573 , \B[6]_b0 );
or ( \245_b1 , \I[1]_b1 , w_575 );
not ( w_575 , w_576 );
and ( \245_b0 , \I[1]_b0 , w_577 );
and ( w_576 ,  , w_577 );
buf ( w_575 , \I[0]_b1 );
not ( w_575 , w_578 );
not (  , w_579 );
and ( w_578 , w_579 , \I[0]_b0 );
buf ( \246_b1 , \245_b1 );
not ( \246_b1 , w_580 );
not ( \246_b0 , w_581 );
and ( w_580 , w_581 , \245_b0 );
buf ( \247_b1 , \A[0][2]_b1 );
not ( \247_b1 , w_582 );
not ( \247_b0 , w_583 );
and ( w_582 , w_583 , \A[0][2]_b0 );
or ( \248_b1 , \246_b1 , w_584 );
or ( \248_b0 , \246_b0 , \247_b0 );
not ( \247_b0 , w_585 );
and ( w_585 , w_584 , \247_b1 );
or ( \249_b1 , \A[1][2]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_586 );
and ( \249_b0 , \A[1][2]_b0 , w_587 );
and ( w_586 , w_587 , \I[0]_b0 );
or ( \250_b1 , \A[2][2]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_588 );
and ( \250_b0 , \A[2][2]_b0 , w_589 );
and ( w_588 , w_589 , \I[1]_b0 );
or ( \251_b1 , \249_b1 , w_591 );
not ( w_591 , w_592 );
and ( \251_b0 , \249_b0 , w_593 );
and ( w_592 ,  , w_593 );
buf ( w_591 , \250_b1 );
not ( w_591 , w_594 );
not (  , w_595 );
and ( w_594 , w_595 , \250_b0 );
or ( \252_b1 , \248_b1 , w_597 );
not ( w_597 , w_598 );
and ( \252_b0 , \248_b0 , w_599 );
and ( w_598 ,  , w_599 );
buf ( w_597 , \251_b1 );
not ( w_597 , w_600 );
not (  , w_601 );
and ( w_600 , w_601 , \251_b0 );
buf ( \253_b1 , \252_b1 );
buf ( \253_b0 , \252_b0 );
or ( \254_b1 , \253_b1 , w_603 );
not ( w_603 , w_604 );
and ( \254_b0 , \253_b0 , w_605 );
and ( w_604 ,  , w_605 );
buf ( w_603 , \B[9]_b1 );
not ( w_603 , w_606 );
not (  , w_607 );
and ( w_606 , w_607 , \B[9]_b0 );
or ( \255_b1 , \244_b1 , \254_b1 );
xor ( \255_b0 , \244_b0 , w_608 );
not ( w_608 , w_609 );
and ( w_609 , \254_b1 , \254_b0 );
or ( \256_b1 , \88_b1 , w_611 );
not ( w_611 , w_612 );
and ( \256_b0 , \88_b0 , w_613 );
and ( w_612 ,  , w_613 );
buf ( w_611 , \B[4]_b1 );
not ( w_611 , w_614 );
not (  , w_615 );
and ( w_614 , w_615 , \B[4]_b0 );
or ( \257_b1 , \255_b1 , \256_b1 );
not ( \256_b1 , w_616 );
and ( \257_b0 , \255_b0 , w_617 );
and ( w_616 , w_617 , \256_b0 );
or ( \258_b1 , \244_b1 , \254_b1 );
not ( \254_b1 , w_618 );
and ( \258_b0 , \244_b0 , w_619 );
and ( w_618 , w_619 , \254_b0 );
or ( \259_b1 , \257_b1 , w_620 );
or ( \259_b0 , \257_b0 , \258_b0 );
not ( \258_b0 , w_621 );
and ( w_621 , w_620 , \258_b1 );
or ( \260_b1 , \243_b1 , \259_b1 );
not ( \259_b1 , w_622 );
and ( \260_b0 , \243_b0 , w_623 );
and ( w_622 , w_623 , \259_b0 );
or ( \261_b1 , \235_b1 , \242_b1 );
not ( \242_b1 , w_624 );
and ( \261_b0 , \235_b0 , w_625 );
and ( w_624 , w_625 , \242_b0 );
or ( \262_b1 , \260_b1 , w_626 );
or ( \262_b0 , \260_b0 , \261_b0 );
not ( \261_b0 , w_627 );
and ( w_627 , w_626 , \261_b1 );
buf ( \263_b1 , \262_b1 );
not ( \263_b1 , w_628 );
not ( \263_b0 , w_629 );
and ( w_628 , w_629 , \262_b0 );
or ( \264_b1 , \226_b1 , w_631 );
not ( w_631 , w_632 );
and ( \264_b0 , \226_b0 , w_633 );
and ( w_632 ,  , w_633 );
buf ( w_631 , \263_b1 );
not ( w_631 , w_634 );
not (  , w_635 );
and ( w_634 , w_635 , \263_b0 );
buf ( \265_b1 , \209_b1 );
not ( \265_b1 , w_636 );
not ( \265_b0 , w_637 );
and ( w_636 , w_637 , \209_b0 );
or ( \266_b1 , \265_b1 , w_639 );
not ( w_639 , w_640 );
and ( \266_b0 , \265_b0 , w_641 );
and ( w_640 ,  , w_641 );
buf ( w_639 , \223_b1 );
not ( w_639 , w_642 );
not (  , w_643 );
and ( w_642 , w_643 , \223_b0 );
or ( \267_b1 , \264_b1 , w_645 );
not ( w_645 , w_646 );
and ( \267_b0 , \264_b0 , w_647 );
and ( w_646 ,  , w_647 );
buf ( w_645 , \266_b1 );
not ( w_645 , w_648 );
not (  , w_649 );
and ( w_648 , w_649 , \266_b0 );
or ( \268_b1 , \207_b1 , \267_b1 );
not ( \267_b1 , w_650 );
and ( \268_b0 , \207_b0 , w_651 );
and ( w_650 , w_651 , \267_b0 );
or ( \269_b1 , \197_b1 , \206_b1 );
not ( \206_b1 , w_652 );
and ( \269_b0 , \197_b0 , w_653 );
and ( w_652 , w_653 , \206_b0 );
or ( \270_b1 , \268_b1 , w_654 );
or ( \270_b0 , \268_b0 , \269_b0 );
not ( \269_b0 , w_655 );
and ( w_655 , w_654 , \269_b1 );
or ( \271_b1 , \170_b1 , w_657 );
not ( w_657 , w_658 );
and ( \271_b0 , \170_b0 , w_659 );
and ( w_658 ,  , w_659 );
buf ( w_657 , \270_b1 );
not ( w_657 , w_660 );
not (  , w_661 );
and ( w_660 , w_661 , \270_b0 );
buf ( \272_b1 , \271_b1 );
not ( \272_b1 , w_662 );
not ( \272_b0 , w_663 );
and ( w_662 , w_663 , \271_b0 );
buf ( \273_b1 , \272_b1 );
not ( \273_b1 , w_664 );
not ( \273_b0 , w_665 );
and ( w_664 , w_665 , \272_b0 );
buf ( \274_b1 , \270_b1 );
not ( \274_b1 , w_666 );
not ( \274_b0 , w_667 );
and ( w_666 , w_667 , \270_b0 );
or ( \275_b1 , \274_b1 , w_669 );
not ( w_669 , w_670 );
and ( \275_b0 , \274_b0 , w_671 );
and ( w_670 ,  , w_671 );
buf ( w_669 , \169_b1 );
not ( w_669 , w_672 );
not (  , w_673 );
and ( w_672 , w_673 , \169_b0 );
or ( \276_b1 , \273_b1 , w_675 );
not ( w_675 , w_676 );
and ( \276_b0 , \273_b0 , w_677 );
and ( w_676 ,  , w_677 );
buf ( w_675 , \275_b1 );
not ( w_675 , w_678 );
not (  , w_679 );
and ( w_678 , w_679 , \275_b0 );
buf ( \277_b1 , \276_b1 );
not ( \277_b1 , w_680 );
not ( \277_b0 , w_681 );
and ( w_680 , w_681 , \276_b0 );
buf ( \280_b1 , \279_b1 );
not ( \280_b1 , w_682 );
not ( \280_b0 , w_683 );
and ( w_682 , w_683 , \279_b0 );
or ( \281_b1 , \278_b1 , w_684 );
or ( \281_b0 , \278_b0 , \280_b0 );
not ( \280_b0 , w_685 );
and ( w_685 , w_684 , \280_b1 );
and ( \282_b0 , \277_b0 , w_686 );
and ( \282_b0 , 1'b1_b0 , w_687 );
and ( w_700 , w_701 , w_688 );
and ( w_688 , 1'b1_b0 , w_689 );
and ( w_701 , 1'b1_b1 , w_690 );
and ( \282_b1 , \277_b0 , w_691 );
and ( \277_b1 , w_702 , w_692 );
and ( w_701 , 1'b1_b0 , w_693 );
and ( \282_b1 , \282_b0 , w_694 );
and ( w_699 , w_703 , \281_b1 );
or ( w_686 , w_687 , w_695 );
or ( w_695 , w_689 , \281_b0 );
or ( w_690 , w_691 , w_696 );
or ( w_696 , w_692 , w_697 );
or ( w_697 , w_693 , w_698 );
or ( w_698 , w_694 , w_699 );
not ( \277_b1 , w_700 );
not ( \277_b0 , w_701 );
not ( \282_b1 , w_702 );
not ( \281_b0 , w_703 );
buf ( \283_b1 , \A[0][1]_b1 );
not ( \283_b1 , w_704 );
not ( \283_b0 , w_705 );
and ( w_704 , w_705 , \A[0][1]_b0 );
or ( \285_b1 , \A[2][1]_b1 , w_707 );
not ( w_707 , w_708 );
and ( \285_b0 , \A[2][1]_b0 , w_709 );
and ( w_708 ,  , w_709 );
buf ( w_707 , \I[1]_b1 );
not ( w_707 , w_710 );
not (  , w_711 );
and ( w_710 , w_711 , \I[1]_b0 );
or ( \286_b1 , \A[1][1]_b1 , w_713 );
not ( w_713 , w_714 );
and ( \286_b0 , \A[1][1]_b0 , w_715 );
and ( w_714 ,  , w_715 );
buf ( w_713 , \I[0]_b1 );
not ( w_713 , w_716 );
not (  , w_717 );
and ( w_716 , w_717 , \I[0]_b0 );
or ( \287_b1 , \285_b1 , w_719 );
not ( w_719 , w_720 );
and ( \287_b0 , \285_b0 , w_721 );
and ( w_720 ,  , w_721 );
buf ( w_719 , \286_b1 );
not ( w_719 , w_722 );
not (  , w_723 );
and ( w_722 , w_723 , \286_b0 );
or ( \288_b1 , \284_b1 , w_725 );
not ( w_725 , w_726 );
and ( \288_b0 , \284_b0 , w_727 );
and ( w_726 ,  , w_727 );
buf ( w_725 , \287_b1 );
not ( w_725 , w_728 );
not (  , w_729 );
and ( w_728 , w_729 , \287_b0 );
buf ( \289_b1 , \288_b1 );
not ( \289_b1 , w_730 );
not ( \289_b0 , w_731 );
and ( w_730 , w_731 , \288_b0 );
or ( \290_b1 , \I[1]_b1 , w_733 );
not ( w_733 , w_734 );
and ( \290_b0 , \I[1]_b0 , w_735 );
and ( w_734 ,  , w_735 );
buf ( w_733 , \I[0]_b1 );
not ( w_733 , w_736 );
not (  , w_737 );
and ( w_736 , w_737 , \I[0]_b0 );
or ( \291_b1 , \290_b1 , w_739 );
not ( w_739 , w_740 );
and ( \291_b0 , \290_b0 , w_741 );
and ( w_740 ,  , w_741 );
buf ( w_739 , \A[0][0]_b1 );
not ( w_739 , w_742 );
not (  , w_743 );
and ( w_742 , w_743 , \A[0][0]_b0 );
or ( \292_b1 , \A[1][0]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_744 );
and ( \292_b0 , \A[1][0]_b0 , w_745 );
and ( w_744 , w_745 , \I[0]_b0 );
or ( \293_b1 , \A[2][0]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_746 );
and ( \293_b0 , \A[2][0]_b0 , w_747 );
and ( w_746 , w_747 , \I[1]_b0 );
or ( \294_b1 , \292_b1 , w_749 );
not ( w_749 , w_750 );
and ( \294_b0 , \292_b0 , w_751 );
and ( w_750 ,  , w_751 );
buf ( w_749 , \293_b1 );
not ( w_749 , w_752 );
not (  , w_753 );
and ( w_752 , w_753 , \293_b0 );
or ( \295_b1 , \291_b1 , w_755 );
not ( w_755 , w_756 );
and ( \295_b0 , \291_b0 , w_757 );
and ( w_756 ,  , w_757 );
buf ( w_755 , \294_b1 );
not ( w_755 , w_758 );
not (  , w_759 );
and ( w_758 , w_759 , \294_b0 );
buf ( \296_b1 , \295_b1 );
buf ( \296_b0 , \295_b0 );
or ( \297_b1 , \129_b1 , w_761 );
not ( w_761 , w_762 );
and ( \297_b0 , \129_b0 , w_763 );
and ( w_762 ,  , w_763 );
buf ( w_761 , \B[8]_b1 );
not ( w_761 , w_764 );
not (  , w_765 );
and ( w_764 , w_765 , \B[8]_b0 );
or ( \298_b1 , \140_b1 , w_767 );
not ( w_767 , w_768 );
and ( \298_b0 , \140_b0 , w_769 );
and ( w_768 ,  , w_769 );
buf ( w_767 , \B[9]_b1 );
not ( w_767 , w_770 );
not (  , w_771 );
and ( w_770 , w_771 , \B[9]_b0 );
or ( \299_b1 , \297_b1 , \298_b1 );
xor ( \299_b0 , \297_b0 , w_772 );
not ( w_772 , w_773 );
and ( w_773 , \298_b1 , \298_b0 );
or ( \300_b1 , \129_b1 , w_775 );
not ( w_775 , w_776 );
and ( \300_b0 , \129_b0 , w_777 );
and ( w_776 ,  , w_777 );
buf ( w_775 , \B[7]_b1 );
not ( w_775 , w_778 );
not (  , w_779 );
and ( w_778 , w_779 , \B[7]_b0 );
or ( \301_b1 , \88_b1 , w_781 );
not ( w_781 , w_782 );
and ( \301_b0 , \88_b0 , w_783 );
and ( w_782 ,  , w_783 );
buf ( w_781 , \B[9]_b1 );
not ( w_781 , w_784 );
not (  , w_785 );
and ( w_784 , w_785 , \B[9]_b0 );
or ( \302_b1 , \300_b1 , \301_b1 );
xor ( \302_b0 , \300_b0 , w_786 );
not ( w_786 , w_787 );
and ( w_787 , \301_b1 , \301_b0 );
or ( \303_b1 , \140_b1 , w_789 );
not ( w_789 , w_790 );
and ( \303_b0 , \140_b0 , w_791 );
and ( w_790 ,  , w_791 );
buf ( w_789 , \B[8]_b1 );
not ( w_789 , w_792 );
not (  , w_793 );
and ( w_792 , w_793 , \B[8]_b0 );
or ( \304_b1 , \302_b1 , \303_b1 );
not ( \303_b1 , w_794 );
and ( \304_b0 , \302_b0 , w_795 );
and ( w_794 , w_795 , \303_b0 );
or ( \305_b1 , \300_b1 , \301_b1 );
not ( \301_b1 , w_796 );
and ( \305_b0 , \300_b0 , w_797 );
and ( w_796 , w_797 , \301_b0 );
or ( \306_b1 , \304_b1 , w_798 );
or ( \306_b0 , \304_b0 , \305_b0 );
not ( \305_b0 , w_799 );
and ( w_799 , w_798 , \305_b1 );
or ( \307_b1 , \299_b1 , \306_b1 );
not ( \306_b1 , w_800 );
and ( \307_b0 , \299_b0 , w_801 );
and ( w_800 , w_801 , \306_b0 );
or ( \308_b1 , \297_b1 , \298_b1 );
not ( \298_b1 , w_802 );
and ( \308_b0 , \297_b0 , w_803 );
and ( w_802 , w_803 , \298_b0 );
or ( \309_b1 , \307_b1 , w_804 );
or ( \309_b0 , \307_b0 , \308_b0 );
not ( \308_b0 , w_805 );
and ( w_805 , w_804 , \308_b1 );
or ( \310_b1 , \129_b1 , w_807 );
not ( w_807 , w_808 );
and ( \310_b0 , \129_b0 , w_809 );
and ( w_808 ,  , w_809 );
buf ( w_807 , \B[9]_b1 );
not ( w_807 , w_810 );
not (  , w_811 );
and ( w_810 , w_811 , \B[9]_b0 );
or ( \311_b1 , \309_b1 , w_813 );
not ( w_813 , w_814 );
and ( \311_b0 , \309_b0 , w_815 );
and ( w_814 ,  , w_815 );
buf ( w_813 , \310_b1 );
not ( w_813 , w_816 );
not (  , w_817 );
and ( w_816 , w_817 , \310_b0 );
buf ( \312_b1 , \311_b1 );
not ( \312_b1 , w_818 );
not ( \312_b0 , w_819 );
and ( w_818 , w_819 , \311_b0 );
or ( \313_b1 , \187_b1 , \190_b1 );
xor ( \313_b0 , \187_b0 , w_820 );
not ( w_820 , w_821 );
and ( w_821 , \190_b1 , \190_b0 );
or ( \314_b1 , \313_b1 , \188_b1 );
xor ( \314_b0 , \313_b0 , w_822 );
not ( w_822 , w_823 );
and ( w_823 , \188_b1 , \188_b0 );
or ( \315_b1 , \175_b1 , \173_b1 );
xor ( \315_b0 , \175_b0 , w_824 );
not ( w_824 , w_825 );
and ( w_825 , \173_b1 , \173_b0 );
or ( \316_b1 , \315_b1 , w_826 );
xor ( \316_b0 , \315_b0 , w_828 );
not ( w_828 , w_829 );
and ( w_829 , w_826 , w_827 );
buf ( w_826 , \178_b1 );
not ( w_826 , w_830 );
not ( w_827 , w_831 );
and ( w_830 , w_831 , \178_b0 );
or ( \317_b1 , \314_b1 , \316_b1 );
not ( \316_b1 , w_832 );
and ( \317_b0 , \314_b0 , w_833 );
and ( w_832 , w_833 , \316_b0 );
or ( \318_b1 , \233_b1 , w_835 );
not ( w_835 , w_836 );
and ( \318_b0 , \233_b0 , w_837 );
and ( w_836 ,  , w_837 );
buf ( w_835 , \B[8]_b1 );
not ( w_835 , w_838 );
not (  , w_839 );
and ( w_838 , w_839 , \B[8]_b0 );
or ( \319_b1 , \100_b1 , w_841 );
not ( w_841 , w_842 );
and ( \319_b0 , \100_b0 , w_843 );
and ( w_842 ,  , w_843 );
buf ( w_841 , \B[7]_b1 );
not ( w_841 , w_844 );
not (  , w_845 );
and ( w_844 , w_845 , \B[7]_b0 );
or ( \320_b1 , \318_b1 , \319_b1 );
xor ( \320_b0 , \318_b0 , w_846 );
not ( w_846 , w_847 );
and ( w_847 , \319_b1 , \319_b0 );
or ( \321_b1 , \129_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_848 );
and ( \321_b0 , \129_b0 , w_849 );
and ( w_848 , w_849 , \B[1]_b0 );
or ( \322_b1 , \139_b1 , \B[2]_b1 );
not ( \B[2]_b1 , w_850 );
and ( \322_b0 , \139_b0 , w_851 );
and ( w_850 , w_851 , \B[2]_b0 );
or ( \323_b1 , \321_b1 , w_853 );
not ( w_853 , w_854 );
and ( \323_b0 , \321_b0 , w_855 );
and ( w_854 ,  , w_855 );
buf ( w_853 , \322_b1 );
not ( w_853 , w_856 );
not (  , w_857 );
and ( w_856 , w_857 , \322_b0 );
or ( \324_b1 , \320_b1 , \323_b1 );
not ( \323_b1 , w_858 );
and ( \324_b0 , \320_b0 , w_859 );
and ( w_858 , w_859 , \323_b0 );
or ( \325_b1 , \318_b1 , \319_b1 );
not ( \319_b1 , w_860 );
and ( \325_b0 , \318_b0 , w_861 );
and ( w_860 , w_861 , \319_b0 );
or ( \326_b1 , \324_b1 , w_862 );
or ( \326_b0 , \324_b0 , \325_b0 );
not ( \325_b0 , w_863 );
and ( w_863 , w_862 , \325_b1 );
or ( \327_b1 , \317_b1 , w_865 );
not ( w_865 , w_866 );
and ( \327_b0 , \317_b0 , w_867 );
and ( w_866 ,  , w_867 );
buf ( w_865 , \326_b1 );
not ( w_865 , w_868 );
not (  , w_869 );
and ( w_868 , w_869 , \326_b0 );
buf ( \328_b1 , \316_b1 );
not ( \328_b1 , w_870 );
not ( \328_b0 , w_871 );
and ( w_870 , w_871 , \316_b0 );
buf ( \329_b1 , \314_b1 );
not ( \329_b1 , w_872 );
not ( \329_b0 , w_873 );
and ( w_872 , w_873 , \314_b0 );
or ( \330_b1 , \328_b1 , \329_b1 );
not ( \329_b1 , w_874 );
and ( \330_b0 , \328_b0 , w_875 );
and ( w_874 , w_875 , \329_b0 );
or ( \331_b1 , \327_b1 , w_877 );
not ( w_877 , w_878 );
and ( \331_b0 , \327_b0 , w_879 );
and ( w_878 ,  , w_879 );
buf ( w_877 , \330_b1 );
not ( w_877 , w_880 );
not (  , w_881 );
and ( w_880 , w_881 , \330_b0 );
buf ( \332_b1 , \331_b1 );
not ( \332_b1 , w_882 );
not ( \332_b0 , w_883 );
and ( w_882 , w_883 , \331_b0 );
or ( \333_b1 , \209_b1 , \262_b1 );
xor ( \333_b0 , \209_b0 , w_884 );
not ( w_884 , w_885 );
and ( w_885 , \262_b1 , \262_b0 );
or ( \334_b1 , \333_b1 , w_886 );
xor ( \334_b0 , \333_b0 , w_888 );
not ( w_888 , w_889 );
and ( w_889 , w_886 , w_887 );
buf ( w_886 , \223_b1 );
not ( w_886 , w_890 );
not ( w_887 , w_891 );
and ( w_890 , w_891 , \223_b0 );
buf ( \335_b1 , \334_b1 );
not ( \335_b1 , w_892 );
not ( \335_b0 , w_893 );
and ( w_892 , w_893 , \334_b0 );
or ( \336_b1 , \332_b1 , w_894 );
or ( \336_b0 , \332_b0 , \335_b0 );
not ( \335_b0 , w_895 );
and ( w_895 , w_894 , \335_b1 );
or ( \337_b1 , \235_b1 , \242_b1 );
xor ( \337_b0 , \235_b0 , w_896 );
not ( w_896 , w_897 );
and ( w_897 , \242_b1 , \242_b0 );
or ( \338_b1 , \337_b1 , \259_b1 );
xor ( \338_b0 , \337_b0 , w_898 );
not ( w_898 , w_899 );
and ( w_899 , \259_b1 , \259_b0 );
or ( \339_b1 , \236_b1 , \237_b1 );
xor ( \339_b0 , \236_b0 , w_900 );
not ( w_900 , w_901 );
and ( w_901 , \237_b1 , \237_b0 );
or ( \340_b1 , \339_b1 , \239_b1 );
xor ( \340_b0 , \339_b0 , w_902 );
not ( w_902 , w_903 );
and ( w_903 , \239_b1 , \239_b0 );
buf ( \341_b1 , \340_b1 );
not ( \341_b1 , w_904 );
not ( \341_b0 , w_905 );
and ( w_904 , w_905 , \340_b0 );
or ( \342_b1 , \119_b1 , w_907 );
not ( w_907 , w_908 );
and ( \342_b0 , \119_b0 , w_909 );
and ( w_908 ,  , w_909 );
buf ( w_907 , \B[4]_b1 );
not ( w_907 , w_910 );
not (  , w_911 );
and ( w_910 , w_911 , \B[4]_b0 );
buf ( \343_b1 , \342_b1 );
not ( \343_b1 , w_912 );
not ( \343_b0 , w_913 );
and ( w_912 , w_913 , \342_b0 );
or ( \344_b1 , \253_b1 , w_915 );
not ( w_915 , w_916 );
and ( \344_b0 , \253_b0 , w_917 );
and ( w_916 ,  , w_917 );
buf ( w_915 , \B[8]_b1 );
not ( w_915 , w_918 );
not (  , w_919 );
and ( w_918 , w_919 , \B[8]_b0 );
buf ( \345_b1 , \344_b1 );
not ( \345_b1 , w_920 );
not ( \345_b0 , w_921 );
and ( w_920 , w_921 , \344_b0 );
or ( \346_b1 , \343_b1 , w_922 );
or ( \346_b0 , \343_b0 , \345_b0 );
not ( \345_b0 , w_923 );
and ( w_923 , w_922 , \345_b1 );
or ( \347_b1 , \289_b1 , \B[9]_b1 );
not ( \B[9]_b1 , w_924 );
and ( \347_b0 , \289_b0 , w_925 );
and ( w_924 , w_925 , \B[9]_b0 );
or ( \348_b1 , \346_b1 , w_927 );
not ( w_927 , w_928 );
and ( \348_b0 , \346_b0 , w_929 );
and ( w_928 ,  , w_929 );
buf ( w_927 , \347_b1 );
not ( w_927 , w_930 );
not (  , w_931 );
and ( w_930 , w_931 , \347_b0 );
buf ( \349_b1 , \342_b1 );
not ( \349_b1 , w_932 );
not ( \349_b0 , w_933 );
and ( w_932 , w_933 , \342_b0 );
buf ( \350_b1 , \344_b1 );
not ( \350_b1 , w_934 );
not ( \350_b0 , w_935 );
and ( w_934 , w_935 , \344_b0 );
or ( \351_b1 , \349_b1 , w_937 );
not ( w_937 , w_938 );
and ( \351_b0 , \349_b0 , w_939 );
and ( w_938 ,  , w_939 );
buf ( w_937 , \350_b1 );
not ( w_937 , w_940 );
not (  , w_941 );
and ( w_940 , w_941 , \350_b0 );
or ( \352_b1 , \348_b1 , w_943 );
not ( w_943 , w_944 );
and ( \352_b0 , \348_b0 , w_945 );
and ( w_944 ,  , w_945 );
buf ( w_943 , \351_b1 );
not ( w_943 , w_946 );
not (  , w_947 );
and ( w_946 , w_947 , \351_b0 );
or ( \353_b1 , \341_b1 , w_949 );
not ( w_949 , w_950 );
and ( \353_b0 , \341_b0 , w_951 );
and ( w_950 ,  , w_951 );
buf ( w_949 , \352_b1 );
not ( w_949 , w_952 );
not (  , w_953 );
and ( w_952 , w_953 , \352_b0 );
buf ( \354_b1 , \352_b1 );
not ( \354_b1 , w_954 );
not ( \354_b0 , w_955 );
and ( w_954 , w_955 , \352_b0 );
buf ( \355_b1 , \354_b1 );
not ( \355_b1 , w_956 );
not ( \355_b0 , w_957 );
and ( w_956 , w_957 , \354_b0 );
buf ( \356_b1 , \340_b1 );
not ( \356_b1 , w_958 );
not ( \356_b0 , w_959 );
and ( w_958 , w_959 , \340_b0 );
or ( \357_b1 , \355_b1 , w_960 );
or ( \357_b0 , \355_b0 , \356_b0 );
not ( \356_b0 , w_961 );
and ( w_961 , w_960 , \356_b1 );
or ( \358_b1 , \80_b1 , w_963 );
not ( w_963 , w_964 );
and ( \358_b0 , \80_b0 , w_965 );
and ( w_964 ,  , w_965 );
buf ( w_963 , \B[5]_b1 );
not ( w_963 , w_966 );
not (  , w_967 );
and ( w_966 , w_967 , \B[5]_b0 );
buf ( \359_b1 , \358_b1 );
not ( \359_b1 , w_968 );
not ( \359_b0 , w_969 );
and ( w_968 , w_969 , \358_b0 );
or ( \360_b1 , \88_b1 , w_971 );
not ( w_971 , w_972 );
and ( \360_b0 , \88_b0 , w_973 );
and ( w_972 ,  , w_973 );
buf ( w_971 , \B[3]_b1 );
not ( w_971 , w_974 );
not (  , w_975 );
and ( w_974 , w_975 , \B[3]_b0 );
buf ( \361_b1 , \360_b1 );
not ( \361_b1 , w_976 );
not ( \361_b0 , w_977 );
and ( w_976 , w_977 , \360_b0 );
or ( \362_b1 , \359_b1 , w_978 );
or ( \362_b0 , \359_b0 , \361_b0 );
not ( \361_b0 , w_979 );
and ( w_979 , w_978 , \361_b1 );
or ( \363_b1 , \100_b1 , w_981 );
not ( w_981 , w_982 );
and ( \363_b0 , \100_b0 , w_983 );
and ( w_982 ,  , w_983 );
buf ( w_981 , \B[6]_b1 );
not ( w_981 , w_984 );
not (  , w_985 );
and ( w_984 , w_985 , \B[6]_b0 );
buf ( \364_b1 , \363_b1 );
not ( \364_b1 , w_986 );
not ( \364_b0 , w_987 );
and ( w_986 , w_987 , \363_b0 );
or ( \365_b1 , \362_b1 , w_989 );
not ( w_989 , w_990 );
and ( \365_b0 , \362_b0 , w_991 );
and ( w_990 ,  , w_991 );
buf ( w_989 , \364_b1 );
not ( w_989 , w_992 );
not (  , w_993 );
and ( w_992 , w_993 , \364_b0 );
or ( \366_b1 , \360_b1 , w_994 );
or ( \366_b0 , \360_b0 , \358_b0 );
not ( \358_b0 , w_995 );
and ( w_995 , w_994 , \358_b1 );
or ( \367_b1 , \365_b1 , w_997 );
not ( w_997 , w_998 );
and ( \367_b0 , \365_b0 , w_999 );
and ( w_998 ,  , w_999 );
buf ( w_997 , \366_b1 );
not ( w_997 , w_1000 );
not (  , w_1001 );
and ( w_1000 , w_1001 , \366_b0 );
or ( \368_b1 , \357_b1 , w_1003 );
not ( w_1003 , w_1004 );
and ( \368_b0 , \357_b0 , w_1005 );
and ( w_1004 ,  , w_1005 );
buf ( w_1003 , \367_b1 );
not ( w_1003 , w_1006 );
not (  , w_1007 );
and ( w_1006 , w_1007 , \367_b0 );
or ( \369_b1 , \353_b1 , \368_b1 );
not ( \368_b1 , w_1008 );
and ( \369_b0 , \353_b0 , w_1009 );
and ( w_1008 , w_1009 , \368_b0 );
or ( \370_b1 , \338_b1 , \369_b1 );
xor ( \370_b0 , \338_b0 , w_1010 );
not ( w_1010 , w_1011 );
and ( w_1011 , \369_b1 , \369_b0 );
or ( \371_b1 , \244_b1 , \254_b1 );
xor ( \371_b0 , \244_b0 , w_1012 );
not ( w_1012 , w_1013 );
and ( w_1013 , \254_b1 , \254_b0 );
or ( \372_b1 , \371_b1 , \256_b1 );
xor ( \372_b0 , \371_b0 , w_1014 );
not ( w_1014 , w_1015 );
and ( w_1015 , \256_b1 , \256_b0 );
or ( \373_b1 , \318_b1 , \319_b1 );
xor ( \373_b0 , \318_b0 , w_1016 );
not ( w_1016 , w_1017 );
and ( w_1017 , \319_b1 , \319_b0 );
or ( \374_b1 , \373_b1 , \323_b1 );
xor ( \374_b0 , \373_b0 , w_1018 );
not ( w_1018 , w_1019 );
and ( w_1019 , \323_b1 , \323_b0 );
or ( \375_b1 , \372_b1 , \374_b1 );
xor ( \375_b0 , \372_b0 , w_1020 );
not ( w_1020 , w_1021 );
and ( w_1021 , \374_b1 , \374_b0 );
or ( \376_b1 , \234_b1 , w_1023 );
not ( w_1023 , w_1024 );
and ( \376_b0 , \234_b0 , w_1025 );
and ( w_1024 ,  , w_1025 );
buf ( w_1023 , \B[7]_b1 );
not ( w_1023 , w_1026 );
not (  , w_1027 );
and ( w_1026 , w_1027 , \B[7]_b0 );
or ( \377_b1 , \129_b1 , w_1029 );
not ( w_1029 , w_1030 );
and ( \377_b0 , \129_b0 , w_1031 );
and ( w_1030 ,  , w_1031 );
buf ( w_1029 , \B[0]_b1 );
not ( w_1029 , w_1032 );
not (  , w_1033 );
and ( w_1032 , w_1033 , \B[0]_b0 );
buf ( \378_b1 , \377_b1 );
not ( \378_b1 , w_1034 );
not ( \378_b0 , w_1035 );
and ( w_1034 , w_1035 , \377_b0 );
or ( \379_b1 , \139_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1036 );
and ( \379_b0 , \139_b0 , w_1037 );
and ( w_1036 , w_1037 , \B[1]_b0 );
or ( \380_b1 , \378_b1 , w_1039 );
not ( w_1039 , w_1040 );
and ( \380_b0 , \378_b0 , w_1041 );
and ( w_1040 ,  , w_1041 );
buf ( w_1039 , \379_b1 );
not ( w_1039 , w_1042 );
not (  , w_1043 );
and ( w_1042 , w_1043 , \379_b0 );
or ( \381_b1 , \376_b1 , \380_b1 );
xor ( \381_b0 , \376_b0 , w_1044 );
not ( w_1044 , w_1045 );
and ( w_1045 , \380_b1 , \380_b0 );
or ( \382_b1 , \322_b1 , w_1046 );
xor ( \382_b0 , \322_b0 , w_1048 );
not ( w_1048 , w_1049 );
and ( w_1049 , w_1046 , w_1047 );
buf ( w_1046 , \321_b1 );
not ( w_1046 , w_1050 );
not ( w_1047 , w_1051 );
and ( w_1050 , w_1051 , \321_b0 );
or ( \383_b1 , \381_b1 , \382_b1 );
not ( \382_b1 , w_1052 );
and ( \383_b0 , \381_b0 , w_1053 );
and ( w_1052 , w_1053 , \382_b0 );
or ( \384_b1 , \376_b1 , \380_b1 );
not ( \380_b1 , w_1054 );
and ( \384_b0 , \376_b0 , w_1055 );
and ( w_1054 , w_1055 , \380_b0 );
or ( \385_b1 , \383_b1 , w_1056 );
or ( \385_b0 , \383_b0 , \384_b0 );
not ( \384_b0 , w_1057 );
and ( w_1057 , w_1056 , \384_b1 );
or ( \386_b1 , \375_b1 , \385_b1 );
not ( \385_b1 , w_1058 );
and ( \386_b0 , \375_b0 , w_1059 );
and ( w_1058 , w_1059 , \385_b0 );
or ( \387_b1 , \372_b1 , \374_b1 );
not ( \374_b1 , w_1060 );
and ( \387_b0 , \372_b0 , w_1061 );
and ( w_1060 , w_1061 , \374_b0 );
or ( \388_b1 , \386_b1 , w_1062 );
or ( \388_b0 , \386_b0 , \387_b0 );
not ( \387_b0 , w_1063 );
and ( w_1063 , w_1062 , \387_b1 );
or ( \389_b1 , \370_b1 , \388_b1 );
not ( \388_b1 , w_1064 );
and ( \389_b0 , \370_b0 , w_1065 );
and ( w_1064 , w_1065 , \388_b0 );
or ( \390_b1 , \338_b1 , \369_b1 );
not ( \369_b1 , w_1066 );
and ( \390_b0 , \338_b0 , w_1067 );
and ( w_1066 , w_1067 , \369_b0 );
or ( \391_b1 , \389_b1 , w_1068 );
or ( \391_b0 , \389_b0 , \390_b0 );
not ( \390_b0 , w_1069 );
and ( w_1069 , w_1068 , \390_b1 );
buf ( \392_b1 , \391_b1 );
not ( \392_b1 , w_1070 );
not ( \392_b0 , w_1071 );
and ( w_1070 , w_1071 , \391_b0 );
or ( \393_b1 , \336_b1 , w_1073 );
not ( w_1073 , w_1074 );
and ( \393_b0 , \336_b0 , w_1075 );
and ( w_1074 ,  , w_1075 );
buf ( w_1073 , \392_b1 );
not ( w_1073 , w_1076 );
not (  , w_1077 );
and ( w_1076 , w_1077 , \392_b0 );
or ( \394_b1 , \334_b1 , w_1078 );
or ( \394_b0 , \334_b0 , \331_b0 );
not ( \331_b0 , w_1079 );
and ( w_1079 , w_1078 , \331_b1 );
or ( \395_b1 , \393_b1 , w_1081 );
not ( w_1081 , w_1082 );
and ( \395_b0 , \393_b0 , w_1083 );
and ( w_1082 ,  , w_1083 );
buf ( w_1081 , \394_b1 );
not ( w_1081 , w_1084 );
not (  , w_1085 );
and ( w_1084 , w_1085 , \394_b0 );
or ( \396_b1 , \197_b1 , \206_b1 );
xor ( \396_b0 , \197_b0 , w_1086 );
not ( w_1086 , w_1087 );
and ( w_1087 , \206_b1 , \206_b0 );
or ( \397_b1 , \396_b1 , \267_b1 );
xor ( \397_b0 , \396_b0 , w_1088 );
not ( w_1088 , w_1089 );
and ( w_1089 , \267_b1 , \267_b0 );
or ( \398_b1 , \395_b1 , w_1090 );
or ( \398_b0 , \395_b0 , \397_b0 );
not ( \397_b0 , w_1091 );
and ( w_1091 , w_1090 , \397_b1 );
or ( \399_b1 , \398_b1 , w_1093 );
not ( w_1093 , w_1094 );
and ( \399_b0 , \398_b0 , w_1095 );
and ( w_1094 ,  , w_1095 );
buf ( w_1093 , \272_b1 );
not ( w_1093 , w_1096 );
not (  , w_1097 );
and ( w_1096 , w_1097 , \272_b0 );
or ( \400_b1 , \146_b1 , \147_b1 );
xor ( \400_b0 , \146_b0 , w_1098 );
not ( w_1098 , w_1099 );
and ( w_1099 , \147_b1 , \147_b0 );
or ( \401_b1 , \400_b1 , \149_b1 );
not ( \149_b1 , w_1100 );
and ( \401_b0 , \400_b0 , w_1101 );
and ( w_1100 , w_1101 , \149_b0 );
or ( \402_b1 , \146_b1 , \147_b1 );
not ( \147_b1 , w_1102 );
and ( \402_b0 , \146_b0 , w_1103 );
and ( w_1102 , w_1103 , \147_b0 );
or ( \403_b1 , \401_b1 , w_1104 );
or ( \403_b0 , \401_b0 , \402_b0 );
not ( \402_b0 , w_1105 );
and ( w_1105 , w_1104 , \402_b1 );
or ( \404_b1 , \300_b1 , \301_b1 );
xor ( \404_b0 , \300_b0 , w_1106 );
not ( w_1106 , w_1107 );
and ( w_1107 , \301_b1 , \301_b0 );
or ( \405_b1 , \404_b1 , \303_b1 );
xor ( \405_b0 , \404_b0 , w_1108 );
not ( w_1108 , w_1109 );
and ( w_1109 , \303_b1 , \303_b0 );
or ( \406_b1 , \403_b1 , \405_b1 );
xor ( \406_b0 , \403_b0 , w_1110 );
not ( w_1110 , w_1111 );
and ( w_1111 , \405_b1 , \405_b0 );
or ( \407_b1 , \110_b1 , \144_b1 );
xor ( \407_b0 , \110_b0 , w_1112 );
not ( w_1112 , w_1113 );
and ( w_1113 , \144_b1 , \144_b0 );
or ( \408_b1 , \407_b1 , \150_b1 );
not ( \150_b1 , w_1114 );
and ( \408_b0 , \407_b0 , w_1115 );
and ( w_1114 , w_1115 , \150_b0 );
or ( \409_b1 , \110_b1 , \144_b1 );
not ( \144_b1 , w_1116 );
and ( \409_b0 , \110_b0 , w_1117 );
and ( w_1116 , w_1117 , \144_b0 );
or ( \410_b1 , \408_b1 , w_1118 );
or ( \410_b0 , \408_b0 , \409_b0 );
not ( \409_b0 , w_1119 );
and ( w_1119 , w_1118 , \409_b1 );
or ( \411_b1 , \406_b1 , \410_b1 );
not ( \410_b1 , w_1120 );
and ( \411_b0 , \406_b0 , w_1121 );
and ( w_1120 , w_1121 , \410_b0 );
or ( \412_b1 , \403_b1 , \405_b1 );
not ( \405_b1 , w_1122 );
and ( \412_b0 , \403_b0 , w_1123 );
and ( w_1122 , w_1123 , \405_b0 );
or ( \413_b1 , \411_b1 , w_1124 );
or ( \413_b0 , \411_b0 , \412_b0 );
not ( \412_b0 , w_1125 );
and ( w_1125 , w_1124 , \412_b1 );
or ( \414_b1 , \297_b1 , \298_b1 );
xor ( \414_b0 , \297_b0 , w_1126 );
not ( w_1126 , w_1127 );
and ( w_1127 , \298_b1 , \298_b0 );
or ( \415_b1 , \414_b1 , \306_b1 );
xor ( \415_b0 , \414_b0 , w_1128 );
not ( w_1128 , w_1129 );
and ( w_1129 , \306_b1 , \306_b0 );
or ( \416_b1 , \413_b1 , w_1131 );
not ( w_1131 , w_1132 );
and ( \416_b0 , \413_b0 , w_1133 );
and ( w_1132 ,  , w_1133 );
buf ( w_1131 , \415_b1 );
not ( w_1131 , w_1134 );
not (  , w_1135 );
and ( w_1134 , w_1135 , \415_b0 );
or ( \417_b1 , \109_b1 , \151_b1 );
xor ( \417_b0 , \109_b0 , w_1136 );
not ( w_1136 , w_1137 );
and ( w_1137 , \151_b1 , \151_b0 );
or ( \418_b1 , \417_b1 , \168_b1 );
not ( \168_b1 , w_1138 );
and ( \418_b0 , \417_b0 , w_1139 );
and ( w_1138 , w_1139 , \168_b0 );
or ( \419_b1 , \109_b1 , \151_b1 );
not ( \151_b1 , w_1140 );
and ( \419_b0 , \109_b0 , w_1141 );
and ( w_1140 , w_1141 , \151_b0 );
or ( \420_b1 , \418_b1 , w_1142 );
or ( \420_b0 , \418_b0 , \419_b0 );
not ( \419_b0 , w_1143 );
and ( w_1143 , w_1142 , \419_b1 );
or ( \421_b1 , \403_b1 , \405_b1 );
xor ( \421_b0 , \403_b0 , w_1144 );
not ( w_1144 , w_1145 );
and ( w_1145 , \405_b1 , \405_b0 );
or ( \422_b1 , \421_b1 , \410_b1 );
xor ( \422_b0 , \421_b0 , w_1146 );
not ( w_1146 , w_1147 );
and ( w_1147 , \410_b1 , \410_b0 );
or ( \423_b1 , \420_b1 , w_1149 );
not ( w_1149 , w_1150 );
and ( \423_b0 , \420_b0 , w_1151 );
and ( w_1150 ,  , w_1151 );
buf ( w_1149 , \422_b1 );
not ( w_1149 , w_1152 );
not (  , w_1153 );
and ( w_1152 , w_1153 , \422_b0 );
or ( \424_b1 , \416_b1 , w_1155 );
not ( w_1155 , w_1156 );
and ( \424_b0 , \416_b0 , w_1157 );
and ( w_1156 ,  , w_1157 );
buf ( w_1155 , \423_b1 );
not ( w_1155 , w_1158 );
not (  , w_1159 );
and ( w_1158 , w_1159 , \423_b0 );
or ( \425_b1 , \399_b1 , w_1161 );
not ( w_1161 , w_1162 );
and ( \425_b0 , \399_b0 , w_1163 );
and ( w_1162 ,  , w_1163 );
buf ( w_1161 , \424_b1 );
not ( w_1161 , w_1164 );
not (  , w_1165 );
and ( w_1164 , w_1165 , \424_b0 );
buf ( \426_b1 , \425_b1 );
not ( \426_b1 , w_1166 );
not ( \426_b0 , w_1167 );
and ( w_1166 , w_1167 , \425_b0 );
or ( \427_b1 , \338_b1 , \369_b1 );
xor ( \427_b0 , \338_b0 , w_1168 );
not ( w_1168 , w_1169 );
and ( w_1169 , \369_b1 , \369_b0 );
or ( \428_b1 , \427_b1 , \388_b1 );
xor ( \428_b0 , \427_b0 , w_1170 );
not ( w_1170 , w_1171 );
and ( w_1171 , \388_b1 , \388_b0 );
or ( \429_b1 , \328_b1 , \329_b1 );
xor ( \429_b0 , \328_b0 , w_1172 );
not ( w_1172 , w_1173 );
and ( w_1173 , \329_b1 , \329_b0 );
or ( \430_b1 , \429_b1 , \326_b1 );
not ( \326_b1 , w_1174 );
and ( \430_b0 , \429_b0 , w_1175 );
and ( w_1174 , w_1175 , \326_b0 );
buf ( \431_b1 , \429_b1 );
not ( \431_b1 , w_1176 );
not ( \431_b0 , w_1177 );
and ( w_1176 , w_1177 , \429_b0 );
buf ( \432_b1 , \326_b1 );
not ( \432_b1 , w_1178 );
not ( \432_b0 , w_1179 );
and ( w_1178 , w_1179 , \326_b0 );
or ( \433_b1 , \431_b1 , \432_b1 );
not ( \432_b1 , w_1180 );
and ( \433_b0 , \431_b0 , w_1181 );
and ( w_1180 , w_1181 , \432_b0 );
or ( \434_b1 , \430_b1 , w_1182 );
or ( \434_b0 , \430_b0 , \433_b0 );
not ( \433_b0 , w_1183 );
and ( w_1183 , w_1182 , \433_b1 );
or ( \435_b1 , \428_b1 , \434_b1 );
xor ( \435_b0 , \428_b0 , w_1184 );
not ( w_1184 , w_1185 );
and ( w_1185 , \434_b1 , \434_b0 );
buf ( \436_b1 , \367_b1 );
not ( \436_b1 , w_1186 );
not ( \436_b0 , w_1187 );
and ( w_1186 , w_1187 , \367_b0 );
buf ( \437_b1 , \354_b1 );
not ( \437_b1 , w_1188 );
not ( \437_b0 , w_1189 );
and ( w_1188 , w_1189 , \354_b0 );
or ( \438_b1 , \436_b1 , w_1190 );
or ( \438_b0 , \436_b0 , \437_b0 );
not ( \437_b0 , w_1191 );
and ( w_1191 , w_1190 , \437_b1 );
buf ( \439_b1 , \367_b1 );
not ( \439_b1 , w_1192 );
not ( \439_b0 , w_1193 );
and ( w_1192 , w_1193 , \367_b0 );
or ( \440_b1 , \439_b1 , w_1195 );
not ( w_1195 , w_1196 );
and ( \440_b0 , \439_b0 , w_1197 );
and ( w_1196 ,  , w_1197 );
buf ( w_1195 , \352_b1 );
not ( w_1195 , w_1198 );
not (  , w_1199 );
and ( w_1198 , w_1199 , \352_b0 );
or ( \441_b1 , \438_b1 , w_1201 );
not ( w_1201 , w_1202 );
and ( \441_b0 , \438_b0 , w_1203 );
and ( w_1202 ,  , w_1203 );
buf ( w_1201 , \440_b1 );
not ( w_1201 , w_1204 );
not (  , w_1205 );
and ( w_1204 , w_1205 , \440_b0 );
or ( \442_b1 , \441_b1 , \340_b1 );
not ( \340_b1 , w_1206 );
and ( \442_b0 , \441_b0 , w_1207 );
and ( w_1206 , w_1207 , \340_b0 );
buf ( \443_b1 , \441_b1 );
not ( \443_b1 , w_1208 );
not ( \443_b0 , w_1209 );
and ( w_1208 , w_1209 , \441_b0 );
buf ( \444_b1 , \340_b1 );
not ( \444_b1 , w_1210 );
not ( \444_b0 , w_1211 );
and ( w_1210 , w_1211 , \340_b0 );
or ( \445_b1 , \443_b1 , \444_b1 );
not ( \444_b1 , w_1212 );
and ( \445_b0 , \443_b0 , w_1213 );
and ( w_1212 , w_1213 , \444_b0 );
or ( \446_b1 , \442_b1 , w_1215 );
not ( w_1215 , w_1216 );
and ( \446_b0 , \442_b0 , w_1217 );
and ( w_1216 ,  , w_1217 );
buf ( w_1215 , \445_b1 );
not ( w_1215 , w_1218 );
not (  , w_1219 );
and ( w_1218 , w_1219 , \445_b0 );
or ( \447_b1 , \80_b1 , w_1221 );
not ( w_1221 , w_1222 );
and ( \447_b0 , \80_b0 , w_1223 );
and ( w_1222 ,  , w_1223 );
buf ( w_1221 , \B[4]_b1 );
not ( w_1221 , w_1224 );
not (  , w_1225 );
and ( w_1224 , w_1225 , \B[4]_b0 );
or ( \448_b1 , \88_b1 , w_1227 );
not ( w_1227 , w_1228 );
and ( \448_b0 , \88_b0 , w_1229 );
and ( w_1228 ,  , w_1229 );
buf ( w_1227 , \B[2]_b1 );
not ( w_1227 , w_1230 );
not (  , w_1231 );
and ( w_1230 , w_1231 , \B[2]_b0 );
or ( \449_b1 , \447_b1 , \448_b1 );
xor ( \449_b0 , \447_b0 , w_1232 );
not ( w_1232 , w_1233 );
and ( w_1233 , \448_b1 , \448_b0 );
or ( \450_b1 , \B[9]_b1 , w_1235 );
not ( w_1235 , w_1236 );
and ( \450_b0 , \B[9]_b0 , w_1237 );
and ( w_1236 ,  , w_1237 );
buf ( w_1235 , \296_b1 );
not ( w_1235 , w_1238 );
not (  , w_1239 );
and ( w_1238 , w_1239 , \296_b0 );
or ( \451_b1 , \449_b1 , \450_b1 );
not ( \450_b1 , w_1240 );
and ( \451_b0 , \449_b0 , w_1241 );
and ( w_1240 , w_1241 , \450_b0 );
or ( \452_b1 , \447_b1 , \448_b1 );
not ( \448_b1 , w_1242 );
and ( \452_b0 , \447_b0 , w_1243 );
and ( w_1242 , w_1243 , \448_b0 );
or ( \453_b1 , \451_b1 , w_1244 );
or ( \453_b0 , \451_b0 , \452_b0 );
not ( \452_b0 , w_1245 );
and ( w_1245 , w_1244 , \452_b1 );
or ( \454_b1 , \358_b1 , \363_b1 );
xor ( \454_b0 , \358_b0 , w_1246 );
not ( w_1246 , w_1247 );
and ( w_1247 , \363_b1 , \363_b0 );
or ( \455_b1 , \454_b1 , \360_b1 );
xor ( \455_b0 , \454_b0 , w_1248 );
not ( w_1248 , w_1249 );
and ( w_1249 , \360_b1 , \360_b0 );
or ( \456_b1 , \453_b1 , \455_b1 );
xor ( \456_b0 , \453_b0 , w_1250 );
not ( w_1250 , w_1251 );
and ( w_1251 , \455_b1 , \455_b0 );
or ( \457_b1 , \119_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_1252 );
and ( \457_b0 , \119_b0 , w_1253 );
and ( w_1252 , w_1253 , \B[3]_b0 );
or ( \458_b1 , \253_b1 , \B[7]_b1 );
not ( \B[7]_b1 , w_1254 );
and ( \458_b0 , \253_b0 , w_1255 );
and ( w_1254 , w_1255 , \B[7]_b0 );
or ( \459_b1 , \457_b1 , w_1256 );
or ( \459_b0 , \457_b0 , \458_b0 );
not ( \458_b0 , w_1257 );
and ( w_1257 , w_1256 , \458_b1 );
or ( \460_b1 , \289_b1 , w_1259 );
not ( w_1259 , w_1260 );
and ( \460_b0 , \289_b0 , w_1261 );
and ( w_1260 ,  , w_1261 );
buf ( w_1259 , \B[8]_b1 );
not ( w_1259 , w_1262 );
not (  , w_1263 );
and ( w_1262 , w_1263 , \B[8]_b0 );
buf ( \461_b1 , \460_b1 );
not ( \461_b1 , w_1264 );
not ( \461_b0 , w_1265 );
and ( w_1264 , w_1265 , \460_b0 );
or ( \462_b1 , \459_b1 , \461_b1 );
not ( \461_b1 , w_1266 );
and ( \462_b0 , \459_b0 , w_1267 );
and ( w_1266 , w_1267 , \461_b0 );
or ( \463_b1 , \457_b1 , \458_b1 );
not ( \458_b1 , w_1268 );
and ( \463_b0 , \457_b0 , w_1269 );
and ( w_1268 , w_1269 , \458_b0 );
or ( \464_b1 , \462_b1 , w_1271 );
not ( w_1271 , w_1272 );
and ( \464_b0 , \462_b0 , w_1273 );
and ( w_1272 ,  , w_1273 );
buf ( w_1271 , \463_b1 );
not ( w_1271 , w_1274 );
not (  , w_1275 );
and ( w_1274 , w_1275 , \463_b0 );
or ( \465_b1 , \456_b1 , \464_b1 );
not ( \464_b1 , w_1276 );
and ( \465_b0 , \456_b0 , w_1277 );
and ( w_1276 , w_1277 , \464_b0 );
or ( \466_b1 , \453_b1 , \455_b1 );
not ( \455_b1 , w_1278 );
and ( \466_b0 , \453_b0 , w_1279 );
and ( w_1278 , w_1279 , \455_b0 );
or ( \467_b1 , \465_b1 , w_1280 );
or ( \467_b0 , \465_b0 , \466_b0 );
not ( \466_b0 , w_1281 );
and ( w_1281 , w_1280 , \466_b1 );
or ( \468_b1 , \446_b1 , \467_b1 );
xor ( \468_b0 , \446_b0 , w_1282 );
not ( w_1282 , w_1283 );
and ( w_1283 , \467_b1 , \467_b0 );
or ( \469_b1 , \342_b1 , \350_b1 );
xor ( \469_b0 , \342_b0 , w_1284 );
not ( w_1284 , w_1285 );
and ( w_1285 , \350_b1 , \350_b0 );
or ( \470_b1 , \469_b1 , \347_b1 );
xor ( \470_b0 , \469_b0 , w_1286 );
not ( w_1286 , w_1287 );
and ( w_1287 , \347_b1 , \347_b0 );
or ( \471_b1 , \234_b1 , w_1289 );
not ( w_1289 , w_1290 );
and ( \471_b0 , \234_b0 , w_1291 );
and ( w_1290 ,  , w_1291 );
buf ( w_1289 , \B[6]_b1 );
not ( w_1289 , w_1292 );
not (  , w_1293 );
and ( w_1292 , w_1293 , \B[6]_b0 );
or ( \472_b1 , \100_b1 , w_1295 );
not ( w_1295 , w_1296 );
and ( \472_b0 , \100_b0 , w_1297 );
and ( w_1296 ,  , w_1297 );
buf ( w_1295 , \B[5]_b1 );
not ( w_1295 , w_1298 );
not (  , w_1299 );
and ( w_1298 , w_1299 , \B[5]_b0 );
or ( \473_b1 , \471_b1 , \472_b1 );
xor ( \473_b0 , \471_b0 , w_1300 );
not ( w_1300 , w_1301 );
and ( w_1301 , \472_b1 , \472_b0 );
buf ( \474_b1 , \379_b1 );
not ( \474_b1 , w_1302 );
not ( \474_b0 , w_1303 );
and ( w_1302 , w_1303 , \379_b0 );
buf ( \475_b1 , \377_b1 );
not ( \475_b1 , w_1304 );
not ( \475_b0 , w_1305 );
and ( w_1304 , w_1305 , \377_b0 );
or ( \476_b1 , \474_b1 , \475_b1 );
not ( \475_b1 , w_1306 );
and ( \476_b0 , \474_b0 , w_1307 );
and ( w_1306 , w_1307 , \475_b0 );
or ( \477_b1 , \379_b1 , \377_b1 );
not ( \377_b1 , w_1308 );
and ( \477_b0 , \379_b0 , w_1309 );
and ( w_1308 , w_1309 , \377_b0 );
or ( \478_b1 , \476_b1 , w_1311 );
not ( w_1311 , w_1312 );
and ( \478_b0 , \476_b0 , w_1313 );
and ( w_1312 ,  , w_1313 );
buf ( w_1311 , \477_b1 );
not ( w_1311 , w_1314 );
not (  , w_1315 );
and ( w_1314 , w_1315 , \477_b0 );
or ( \479_b1 , \473_b1 , \478_b1 );
not ( \478_b1 , w_1316 );
and ( \479_b0 , \473_b0 , w_1317 );
and ( w_1316 , w_1317 , \478_b0 );
or ( \480_b1 , \471_b1 , \472_b1 );
not ( \472_b1 , w_1318 );
and ( \480_b0 , \471_b0 , w_1319 );
and ( w_1318 , w_1319 , \472_b0 );
or ( \481_b1 , \479_b1 , w_1320 );
or ( \481_b0 , \479_b0 , \480_b0 );
not ( \480_b0 , w_1321 );
and ( w_1321 , w_1320 , \480_b1 );
or ( \482_b1 , \470_b1 , \481_b1 );
xor ( \482_b0 , \470_b0 , w_1322 );
not ( w_1322 , w_1323 );
and ( w_1323 , \481_b1 , \481_b0 );
or ( \483_b1 , \88_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_1324 );
and ( \483_b0 , \88_b0 , w_1325 );
and ( w_1324 , w_1325 , \B[0]_b0 );
or ( \484_b1 , \379_b1 , w_1327 );
not ( w_1327 , w_1328 );
and ( \484_b0 , \379_b0 , w_1329 );
and ( w_1328 ,  , w_1329 );
buf ( w_1327 , \483_b1 );
not ( w_1327 , w_1330 );
not (  , w_1331 );
and ( w_1330 , w_1331 , \483_b0 );
or ( \485_b1 , \233_b1 , w_1333 );
not ( w_1333 , w_1334 );
and ( \485_b0 , \233_b0 , w_1335 );
and ( w_1334 ,  , w_1335 );
buf ( w_1333 , \B[5]_b1 );
not ( w_1333 , w_1336 );
not (  , w_1337 );
and ( w_1336 , w_1337 , \B[5]_b0 );
buf ( \486_b1 , \485_b1 );
not ( \486_b1 , w_1338 );
not ( \486_b0 , w_1339 );
and ( w_1338 , w_1339 , \485_b0 );
or ( \487_b1 , \100_b1 , w_1341 );
not ( w_1341 , w_1342 );
and ( \487_b0 , \100_b0 , w_1343 );
and ( w_1342 ,  , w_1343 );
buf ( w_1341 , \B[4]_b1 );
not ( w_1341 , w_1344 );
not (  , w_1345 );
and ( w_1344 , w_1345 , \B[4]_b0 );
buf ( \488_b1 , \487_b1 );
not ( \488_b1 , w_1346 );
not ( \488_b0 , w_1347 );
and ( w_1346 , w_1347 , \487_b0 );
or ( \489_b1 , \486_b1 , w_1348 );
or ( \489_b0 , \486_b0 , \488_b0 );
not ( \488_b0 , w_1349 );
and ( w_1349 , w_1348 , \488_b1 );
or ( \490_b1 , \119_b1 , \B[2]_b1 );
not ( \B[2]_b1 , w_1350 );
and ( \490_b0 , \119_b0 , w_1351 );
and ( w_1350 , w_1351 , \B[2]_b0 );
or ( \491_b1 , \489_b1 , w_1353 );
not ( w_1353 , w_1354 );
and ( \491_b0 , \489_b0 , w_1355 );
and ( w_1354 ,  , w_1355 );
buf ( w_1353 , \490_b1 );
not ( w_1353 , w_1356 );
not (  , w_1357 );
and ( w_1356 , w_1357 , \490_b0 );
buf ( \492_b1 , \487_b1 );
not ( \492_b1 , w_1358 );
not ( \492_b0 , w_1359 );
and ( w_1358 , w_1359 , \487_b0 );
buf ( \493_b1 , \485_b1 );
not ( \493_b1 , w_1360 );
not ( \493_b0 , w_1361 );
and ( w_1360 , w_1361 , \485_b0 );
or ( \494_b1 , \492_b1 , w_1363 );
not ( w_1363 , w_1364 );
and ( \494_b0 , \492_b0 , w_1365 );
and ( w_1364 ,  , w_1365 );
buf ( w_1363 , \493_b1 );
not ( w_1363 , w_1366 );
not (  , w_1367 );
and ( w_1366 , w_1367 , \493_b0 );
or ( \495_b1 , \491_b1 , w_1369 );
not ( w_1369 , w_1370 );
and ( \495_b0 , \491_b0 , w_1371 );
and ( w_1370 ,  , w_1371 );
buf ( w_1369 , \494_b1 );
not ( w_1369 , w_1372 );
not (  , w_1373 );
and ( w_1372 , w_1373 , \494_b0 );
buf ( \496_b1 , \495_b1 );
not ( \496_b1 , w_1374 );
not ( \496_b0 , w_1375 );
and ( w_1374 , w_1375 , \495_b0 );
or ( \497_b1 , \484_b1 , \496_b1 );
xor ( \497_b0 , \484_b0 , w_1376 );
not ( w_1376 , w_1377 );
and ( w_1377 , \496_b1 , \496_b0 );
or ( \498_b1 , \289_b1 , w_1379 );
not ( w_1379 , w_1380 );
and ( \498_b0 , \289_b0 , w_1381 );
and ( w_1380 ,  , w_1381 );
buf ( w_1379 , \B[7]_b1 );
not ( w_1379 , w_1382 );
not (  , w_1383 );
and ( w_1382 , w_1383 , \B[7]_b0 );
or ( \499_b1 , \80_b1 , w_1385 );
not ( w_1385 , w_1386 );
and ( \499_b0 , \80_b0 , w_1387 );
and ( w_1386 ,  , w_1387 );
buf ( w_1385 , \B[3]_b1 );
not ( w_1385 , w_1388 );
not (  , w_1389 );
and ( w_1388 , w_1389 , \B[3]_b0 );
or ( \500_b1 , \498_b1 , w_1391 );
not ( w_1391 , w_1392 );
and ( \500_b0 , \498_b0 , w_1393 );
and ( w_1392 ,  , w_1393 );
buf ( w_1391 , \499_b1 );
not ( w_1391 , w_1394 );
not (  , w_1395 );
and ( w_1394 , w_1395 , \499_b0 );
or ( \501_b1 , \296_b1 , \B[8]_b1 );
not ( \B[8]_b1 , w_1396 );
and ( \501_b0 , \296_b0 , w_1397 );
and ( w_1396 , w_1397 , \B[8]_b0 );
or ( \502_b1 , \500_b1 , \501_b1 );
not ( \501_b1 , w_1398 );
and ( \502_b0 , \500_b0 , w_1399 );
and ( w_1398 , w_1399 , \501_b0 );
or ( \503_b1 , \498_b1 , w_1401 );
not ( w_1401 , w_1402 );
and ( \503_b0 , \498_b0 , w_1403 );
and ( w_1402 ,  , w_1403 );
buf ( w_1401 , \499_b1 );
not ( w_1401 , w_1404 );
not (  , w_1405 );
and ( w_1404 , w_1405 , \499_b0 );
or ( \504_b1 , \502_b1 , w_1407 );
not ( w_1407 , w_1408 );
and ( \504_b0 , \502_b0 , w_1409 );
and ( w_1408 ,  , w_1409 );
buf ( w_1407 , \503_b1 );
not ( w_1407 , w_1410 );
not (  , w_1411 );
and ( w_1410 , w_1411 , \503_b0 );
or ( \505_b1 , \497_b1 , \504_b1 );
not ( \504_b1 , w_1412 );
and ( \505_b0 , \497_b0 , w_1413 );
and ( w_1412 , w_1413 , \504_b0 );
or ( \506_b1 , \484_b1 , \496_b1 );
not ( \496_b1 , w_1414 );
and ( \506_b0 , \484_b0 , w_1415 );
and ( w_1414 , w_1415 , \496_b0 );
or ( \507_b1 , \505_b1 , w_1416 );
or ( \507_b0 , \505_b0 , \506_b0 );
not ( \506_b0 , w_1417 );
and ( w_1417 , w_1416 , \506_b1 );
or ( \508_b1 , \482_b1 , \507_b1 );
not ( \507_b1 , w_1418 );
and ( \508_b0 , \482_b0 , w_1419 );
and ( w_1418 , w_1419 , \507_b0 );
or ( \509_b1 , \470_b1 , \481_b1 );
not ( \481_b1 , w_1420 );
and ( \509_b0 , \470_b0 , w_1421 );
and ( w_1420 , w_1421 , \481_b0 );
or ( \510_b1 , \508_b1 , w_1422 );
or ( \510_b0 , \508_b0 , \509_b0 );
not ( \509_b0 , w_1423 );
and ( w_1423 , w_1422 , \509_b1 );
or ( \511_b1 , \468_b1 , \510_b1 );
not ( \510_b1 , w_1424 );
and ( \511_b0 , \468_b0 , w_1425 );
and ( w_1424 , w_1425 , \510_b0 );
or ( \512_b1 , \446_b1 , \467_b1 );
not ( \467_b1 , w_1426 );
and ( \512_b0 , \446_b0 , w_1427 );
and ( w_1426 , w_1427 , \467_b0 );
or ( \513_b1 , \511_b1 , w_1428 );
or ( \513_b0 , \511_b0 , \512_b0 );
not ( \512_b0 , w_1429 );
and ( w_1429 , w_1428 , \512_b1 );
or ( \514_b1 , \435_b1 , w_1430 );
xor ( \514_b0 , \435_b0 , w_1432 );
not ( w_1432 , w_1433 );
and ( w_1433 , w_1430 , w_1431 );
buf ( w_1430 , \513_b1 );
not ( w_1430 , w_1434 );
not ( w_1431 , w_1435 );
and ( w_1434 , w_1435 , \513_b0 );
or ( \515_b1 , \372_b1 , \374_b1 );
xor ( \515_b0 , \372_b0 , w_1436 );
not ( w_1436 , w_1437 );
and ( w_1437 , \374_b1 , \374_b0 );
or ( \516_b1 , \515_b1 , \385_b1 );
xor ( \516_b0 , \515_b0 , w_1438 );
not ( w_1438 , w_1439 );
and ( w_1439 , \385_b1 , \385_b0 );
or ( \517_b1 , \376_b1 , \380_b1 );
xor ( \517_b0 , \376_b0 , w_1440 );
not ( w_1440 , w_1441 );
and ( w_1441 , \380_b1 , \380_b0 );
or ( \518_b1 , \517_b1 , \382_b1 );
xor ( \518_b0 , \517_b0 , w_1442 );
not ( w_1442 , w_1443 );
and ( w_1443 , \382_b1 , \382_b0 );
or ( \519_b1 , \453_b1 , \455_b1 );
xor ( \519_b0 , \453_b0 , w_1444 );
not ( w_1444 , w_1445 );
and ( w_1445 , \455_b1 , \455_b0 );
or ( \520_b1 , \519_b1 , \464_b1 );
xor ( \520_b0 , \519_b0 , w_1446 );
not ( w_1446 , w_1447 );
and ( w_1447 , \464_b1 , \464_b0 );
or ( \521_b1 , \518_b1 , \520_b1 );
xor ( \521_b0 , \518_b0 , w_1448 );
not ( w_1448 , w_1449 );
and ( w_1449 , \520_b1 , \520_b0 );
or ( \522_b1 , \457_b1 , \458_b1 );
xor ( \522_b0 , \457_b0 , w_1450 );
not ( w_1450 , w_1451 );
and ( w_1451 , \458_b1 , \458_b0 );
or ( \523_b1 , \522_b1 , \461_b1 );
not ( \461_b1 , w_1452 );
and ( \523_b0 , \522_b0 , w_1453 );
and ( w_1452 , w_1453 , \461_b0 );
buf ( \524_b1 , \522_b1 );
not ( \524_b1 , w_1454 );
not ( \524_b0 , w_1455 );
and ( w_1454 , w_1455 , \522_b0 );
or ( \525_b1 , \524_b1 , \460_b1 );
not ( \460_b1 , w_1456 );
and ( \525_b0 , \524_b0 , w_1457 );
and ( w_1456 , w_1457 , \460_b0 );
or ( \526_b1 , \523_b1 , w_1459 );
not ( w_1459 , w_1460 );
and ( \526_b0 , \523_b0 , w_1461 );
and ( w_1460 ,  , w_1461 );
buf ( w_1459 , \525_b1 );
not ( w_1459 , w_1462 );
not (  , w_1463 );
and ( w_1462 , w_1463 , \525_b0 );
buf ( \527_b1 , \526_b1 );
not ( \527_b1 , w_1464 );
not ( \527_b0 , w_1465 );
and ( w_1464 , w_1465 , \526_b0 );
or ( \528_b1 , \447_b1 , \448_b1 );
xor ( \528_b0 , \447_b0 , w_1466 );
not ( w_1466 , w_1467 );
and ( w_1467 , \448_b1 , \448_b0 );
or ( \529_b1 , \528_b1 , \450_b1 );
xor ( \529_b0 , \528_b0 , w_1468 );
not ( w_1468 , w_1469 );
and ( w_1469 , \450_b1 , \450_b0 );
or ( \530_b1 , \527_b1 , w_1471 );
not ( w_1471 , w_1472 );
and ( \530_b0 , \527_b0 , w_1473 );
and ( w_1472 ,  , w_1473 );
buf ( w_1471 , \529_b1 );
not ( w_1471 , w_1474 );
not (  , w_1475 );
and ( w_1474 , w_1475 , \529_b0 );
or ( \531_b1 , \253_b1 , \B[6]_b1 );
not ( \B[6]_b1 , w_1476 );
and ( \531_b0 , \253_b0 , w_1477 );
and ( w_1476 , w_1477 , \B[6]_b0 );
or ( \532_b1 , \88_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1478 );
and ( \532_b0 , \88_b0 , w_1479 );
and ( w_1478 , w_1479 , \B[1]_b0 );
buf ( \533_b1 , \532_b1 );
not ( \533_b1 , w_1480 );
not ( \533_b0 , w_1481 );
and ( w_1480 , w_1481 , \532_b0 );
or ( \534_b1 , \140_b1 , w_1483 );
not ( w_1483 , w_1484 );
and ( \534_b0 , \140_b0 , w_1485 );
and ( w_1484 ,  , w_1485 );
buf ( w_1483 , \B[0]_b1 );
not ( w_1483 , w_1486 );
not (  , w_1487 );
and ( w_1486 , w_1487 , \B[0]_b0 );
buf ( \535_b1 , \534_b1 );
not ( \535_b1 , w_1488 );
not ( \535_b0 , w_1489 );
and ( w_1488 , w_1489 , \534_b0 );
or ( \536_b1 , \533_b1 , w_1490 );
or ( \536_b0 , \533_b0 , \535_b0 );
not ( \535_b0 , w_1491 );
and ( w_1491 , w_1490 , \535_b1 );
or ( \537_b1 , \532_b1 , w_1492 );
or ( \537_b0 , \532_b0 , \534_b0 );
not ( \534_b0 , w_1493 );
and ( w_1493 , w_1492 , \534_b1 );
or ( \538_b1 , \536_b1 , w_1495 );
not ( w_1495 , w_1496 );
and ( \538_b0 , \536_b0 , w_1497 );
and ( w_1496 ,  , w_1497 );
buf ( w_1495 , \537_b1 );
not ( w_1495 , w_1498 );
not (  , w_1499 );
and ( w_1498 , w_1499 , \537_b0 );
or ( \539_b1 , \531_b1 , \538_b1 );
xor ( \539_b0 , \531_b0 , w_1500 );
not ( w_1500 , w_1501 );
and ( w_1501 , \538_b1 , \538_b0 );
or ( \540_b1 , \119_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1502 );
and ( \540_b0 , \119_b0 , w_1503 );
and ( w_1502 , w_1503 , \B[1]_b0 );
or ( \541_b1 , \483_b1 , \540_b1 );
not ( \540_b1 , w_1504 );
and ( \541_b0 , \483_b0 , w_1505 );
and ( w_1504 , w_1505 , \540_b0 );
or ( \542_b1 , \539_b1 , \541_b1 );
not ( \541_b1 , w_1506 );
and ( \542_b0 , \539_b0 , w_1507 );
and ( w_1506 , w_1507 , \541_b0 );
or ( \543_b1 , \531_b1 , \538_b1 );
not ( \538_b1 , w_1508 );
and ( \543_b0 , \531_b0 , w_1509 );
and ( w_1508 , w_1509 , \538_b0 );
or ( \544_b1 , \542_b1 , w_1510 );
or ( \544_b0 , \542_b0 , \543_b0 );
not ( \543_b0 , w_1511 );
and ( w_1511 , w_1510 , \543_b1 );
or ( \545_b1 , \530_b1 , \544_b1 );
not ( \544_b1 , w_1512 );
and ( \545_b0 , \530_b0 , w_1513 );
and ( w_1512 , w_1513 , \544_b0 );
or ( \546_b1 , \527_b1 , w_1515 );
not ( w_1515 , w_1516 );
and ( \546_b0 , \527_b0 , w_1517 );
and ( w_1516 ,  , w_1517 );
buf ( w_1515 , \529_b1 );
not ( w_1515 , w_1518 );
not (  , w_1519 );
and ( w_1518 , w_1519 , \529_b0 );
or ( \547_b1 , \545_b1 , w_1521 );
not ( w_1521 , w_1522 );
and ( \547_b0 , \545_b0 , w_1523 );
and ( w_1522 ,  , w_1523 );
buf ( w_1521 , \546_b1 );
not ( w_1521 , w_1524 );
not (  , w_1525 );
and ( w_1524 , w_1525 , \546_b0 );
or ( \548_b1 , \521_b1 , \547_b1 );
not ( \547_b1 , w_1526 );
and ( \548_b0 , \521_b0 , w_1527 );
and ( w_1526 , w_1527 , \547_b0 );
or ( \549_b1 , \518_b1 , \520_b1 );
not ( \520_b1 , w_1528 );
and ( \549_b0 , \518_b0 , w_1529 );
and ( w_1528 , w_1529 , \520_b0 );
or ( \550_b1 , \548_b1 , w_1530 );
or ( \550_b0 , \548_b0 , \549_b0 );
not ( \549_b0 , w_1531 );
and ( w_1531 , w_1530 , \549_b1 );
or ( \551_b1 , \516_b1 , \550_b1 );
xor ( \551_b0 , \516_b0 , w_1532 );
not ( w_1532 , w_1533 );
and ( w_1533 , \550_b1 , \550_b0 );
or ( \552_b1 , \446_b1 , \467_b1 );
xor ( \552_b0 , \446_b0 , w_1534 );
not ( w_1534 , w_1535 );
and ( w_1535 , \467_b1 , \467_b0 );
or ( \553_b1 , \552_b1 , \510_b1 );
xor ( \553_b0 , \552_b0 , w_1536 );
not ( w_1536 , w_1537 );
and ( w_1537 , \510_b1 , \510_b0 );
or ( \554_b1 , \551_b1 , \553_b1 );
not ( \553_b1 , w_1538 );
and ( \554_b0 , \551_b0 , w_1539 );
and ( w_1538 , w_1539 , \553_b0 );
or ( \555_b1 , \516_b1 , \550_b1 );
not ( \550_b1 , w_1540 );
and ( \555_b0 , \516_b0 , w_1541 );
and ( w_1540 , w_1541 , \550_b0 );
or ( \556_b1 , \554_b1 , w_1542 );
or ( \556_b0 , \554_b0 , \555_b0 );
not ( \555_b0 , w_1543 );
and ( w_1543 , w_1542 , \555_b1 );
or ( \557_b1 , \514_b1 , w_1545 );
not ( w_1545 , w_1546 );
and ( \557_b0 , \514_b0 , w_1547 );
and ( w_1546 ,  , w_1547 );
buf ( w_1545 , \556_b1 );
not ( w_1545 , w_1548 );
not (  , w_1549 );
and ( w_1548 , w_1549 , \556_b0 );
buf ( \558_b1 , \428_b1 );
not ( \558_b1 , w_1550 );
not ( \558_b0 , w_1551 );
and ( w_1550 , w_1551 , \428_b0 );
buf ( \559_b1 , \434_b1 );
not ( \559_b1 , w_1552 );
not ( \559_b0 , w_1553 );
and ( w_1552 , w_1553 , \434_b0 );
buf ( \560_b1 , \559_b1 );
not ( \560_b1 , w_1554 );
not ( \560_b0 , w_1555 );
and ( w_1554 , w_1555 , \559_b0 );
or ( \561_b1 , \558_b1 , w_1556 );
or ( \561_b0 , \558_b0 , \560_b0 );
not ( \560_b0 , w_1557 );
and ( w_1557 , w_1556 , \560_b1 );
buf ( \562_b1 , \513_b1 );
not ( \562_b1 , w_1558 );
not ( \562_b0 , w_1559 );
and ( w_1558 , w_1559 , \513_b0 );
or ( \563_b1 , \561_b1 , w_1561 );
not ( w_1561 , w_1562 );
and ( \563_b0 , \561_b0 , w_1563 );
and ( w_1562 ,  , w_1563 );
buf ( w_1561 , \562_b1 );
not ( w_1561 , w_1564 );
not (  , w_1565 );
and ( w_1564 , w_1565 , \562_b0 );
buf ( \564_b1 , \428_b1 );
not ( \564_b1 , w_1566 );
not ( \564_b0 , w_1567 );
and ( w_1566 , w_1567 , \428_b0 );
or ( \565_b1 , \564_b1 , w_1569 );
not ( w_1569 , w_1570 );
and ( \565_b0 , \564_b0 , w_1571 );
and ( w_1570 ,  , w_1571 );
buf ( w_1569 , \434_b1 );
not ( w_1569 , w_1572 );
not (  , w_1573 );
and ( w_1572 , w_1573 , \434_b0 );
or ( \566_b1 , \563_b1 , w_1575 );
not ( w_1575 , w_1576 );
and ( \566_b0 , \563_b0 , w_1577 );
and ( w_1576 ,  , w_1577 );
buf ( w_1575 , \565_b1 );
not ( w_1575 , w_1578 );
not (  , w_1579 );
and ( w_1578 , w_1579 , \565_b0 );
buf ( \567_b1 , \566_b1 );
not ( \567_b1 , w_1580 );
not ( \567_b0 , w_1581 );
and ( w_1580 , w_1581 , \566_b0 );
or ( \568_b1 , \331_b1 , \391_b1 );
xor ( \568_b0 , \331_b0 , w_1582 );
not ( w_1582 , w_1583 );
and ( w_1583 , \391_b1 , \391_b0 );
or ( \569_b1 , \568_b1 , \334_b1 );
xor ( \569_b0 , \568_b0 , w_1584 );
not ( w_1584 , w_1585 );
and ( w_1585 , \334_b1 , \334_b0 );
or ( \570_b1 , \567_b1 , w_1587 );
not ( w_1587 , w_1588 );
and ( \570_b0 , \567_b0 , w_1589 );
and ( w_1588 ,  , w_1589 );
buf ( w_1587 , \569_b1 );
not ( w_1587 , w_1590 );
not (  , w_1591 );
and ( w_1590 , w_1591 , \569_b0 );
or ( \571_b1 , \557_b1 , w_1593 );
not ( w_1593 , w_1594 );
and ( \571_b0 , \557_b0 , w_1595 );
and ( w_1594 ,  , w_1595 );
buf ( w_1593 , \570_b1 );
not ( w_1593 , w_1596 );
not (  , w_1597 );
and ( w_1596 , w_1597 , \570_b0 );
or ( \572_b1 , \426_b1 , w_1599 );
not ( w_1599 , w_1600 );
and ( \572_b0 , \426_b0 , w_1601 );
and ( w_1600 ,  , w_1601 );
buf ( w_1599 , \571_b1 );
not ( w_1599 , w_1602 );
not (  , w_1603 );
and ( w_1602 , w_1603 , \571_b0 );
buf ( \573_b1 , \572_b1 );
not ( \573_b1 , w_1604 );
not ( \573_b0 , w_1605 );
and ( w_1604 , w_1605 , \572_b0 );
or ( \574_b1 , \119_b1 , w_1607 );
not ( w_1607 , w_1608 );
and ( \574_b0 , \119_b0 , w_1609 );
and ( w_1608 ,  , w_1609 );
buf ( w_1607 , \B[0]_b1 );
not ( w_1607 , w_1610 );
not (  , w_1611 );
and ( w_1610 , w_1611 , \B[0]_b0 );
buf ( \575_b1 , \574_b1 );
not ( \575_b1 , w_1612 );
not ( \575_b0 , w_1613 );
and ( w_1612 , w_1613 , \574_b0 );
or ( \576_b1 , \80_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1614 );
and ( \576_b0 , \80_b0 , w_1615 );
and ( w_1614 , w_1615 , \B[1]_b0 );
buf ( \577_b1 , \576_b1 );
not ( \577_b1 , w_1616 );
not ( \577_b0 , w_1617 );
and ( w_1616 , w_1617 , \576_b0 );
or ( \578_b1 , \575_b1 , \577_b1 );
not ( \577_b1 , w_1618 );
and ( \578_b0 , \575_b0 , w_1619 );
and ( w_1618 , w_1619 , \577_b0 );
or ( \579_b1 , \574_b1 , \576_b1 );
not ( \576_b1 , w_1620 );
and ( \579_b0 , \574_b0 , w_1621 );
and ( w_1620 , w_1621 , \576_b0 );
or ( \580_b1 , \578_b1 , w_1623 );
not ( w_1623 , w_1624 );
and ( \580_b0 , \578_b0 , w_1625 );
and ( w_1624 ,  , w_1625 );
buf ( w_1623 , \579_b1 );
not ( w_1623 , w_1626 );
not (  , w_1627 );
and ( w_1626 , w_1627 , \579_b0 );
or ( \581_b1 , \289_b1 , w_1629 );
not ( w_1629 , w_1630 );
and ( \581_b0 , \289_b0 , w_1631 );
and ( w_1630 ,  , w_1631 );
buf ( w_1629 , \B[4]_b1 );
not ( w_1629 , w_1632 );
not (  , w_1633 );
and ( w_1632 , w_1633 , \B[4]_b0 );
or ( \582_b1 , \234_b1 , w_1635 );
not ( w_1635 , w_1636 );
and ( \582_b0 , \234_b0 , w_1637 );
and ( w_1636 ,  , w_1637 );
buf ( w_1635 , \B[2]_b1 );
not ( w_1635 , w_1638 );
not (  , w_1639 );
and ( w_1638 , w_1639 , \B[2]_b0 );
or ( \583_b1 , \581_b1 , \582_b1 );
xor ( \583_b0 , \581_b0 , w_1640 );
not ( w_1640 , w_1641 );
and ( w_1641 , \582_b1 , \582_b0 );
or ( \584_b1 , \253_b1 , w_1643 );
not ( w_1643 , w_1644 );
and ( \584_b0 , \253_b0 , w_1645 );
and ( w_1644 ,  , w_1645 );
buf ( w_1643 , \B[3]_b1 );
not ( w_1643 , w_1646 );
not (  , w_1647 );
and ( w_1646 , w_1647 , \B[3]_b0 );
or ( \585_b1 , \583_b1 , \584_b1 );
not ( \584_b1 , w_1648 );
and ( \585_b0 , \583_b0 , w_1649 );
and ( w_1648 , w_1649 , \584_b0 );
or ( \586_b1 , \581_b1 , \582_b1 );
not ( \582_b1 , w_1650 );
and ( \586_b0 , \581_b0 , w_1651 );
and ( w_1650 , w_1651 , \582_b0 );
or ( \587_b1 , \585_b1 , w_1652 );
or ( \587_b0 , \585_b0 , \586_b0 );
not ( \586_b0 , w_1653 );
and ( w_1653 , w_1652 , \586_b1 );
or ( \588_b1 , \580_b1 , \587_b1 );
xor ( \588_b0 , \580_b0 , w_1654 );
not ( w_1654 , w_1655 );
and ( w_1655 , \587_b1 , \587_b0 );
or ( \589_b1 , \253_b1 , w_1657 );
not ( w_1657 , w_1658 );
and ( \589_b0 , \253_b0 , w_1659 );
and ( w_1658 ,  , w_1659 );
buf ( w_1657 , \B[4]_b1 );
not ( w_1657 , w_1660 );
not (  , w_1661 );
and ( w_1660 , w_1661 , \B[4]_b0 );
or ( \590_b1 , \233_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_1662 );
and ( \590_b0 , \233_b0 , w_1663 );
and ( w_1662 , w_1663 , \B[3]_b0 );
or ( \591_b1 , \589_b1 , \590_b1 );
xor ( \591_b0 , \589_b0 , w_1664 );
not ( w_1664 , w_1665 );
and ( w_1665 , \590_b1 , \590_b0 );
or ( \592_b1 , \100_b1 , w_1667 );
not ( w_1667 , w_1668 );
and ( \592_b0 , \100_b0 , w_1669 );
and ( w_1668 ,  , w_1669 );
buf ( w_1667 , \B[2]_b1 );
not ( w_1667 , w_1670 );
not (  , w_1671 );
and ( w_1670 , w_1671 , \B[2]_b0 );
or ( \593_b1 , \591_b1 , w_1672 );
xor ( \593_b0 , \591_b0 , w_1674 );
not ( w_1674 , w_1675 );
and ( w_1675 , w_1672 , w_1673 );
buf ( w_1672 , \592_b1 );
not ( w_1672 , w_1676 );
not ( w_1673 , w_1677 );
and ( w_1676 , w_1677 , \592_b0 );
or ( \594_b1 , \588_b1 , \593_b1 );
not ( \593_b1 , w_1678 );
and ( \594_b0 , \588_b0 , w_1679 );
and ( w_1678 , w_1679 , \593_b0 );
or ( \595_b1 , \580_b1 , \587_b1 );
not ( \587_b1 , w_1680 );
and ( \595_b0 , \580_b0 , w_1681 );
and ( w_1680 , w_1681 , \587_b0 );
or ( \596_b1 , \594_b1 , w_1682 );
or ( \596_b0 , \594_b0 , \595_b0 );
not ( \595_b0 , w_1683 );
and ( w_1683 , w_1682 , \595_b1 );
buf ( \597_b1 , \596_b1 );
not ( \597_b1 , w_1684 );
not ( \597_b0 , w_1685 );
and ( w_1684 , w_1685 , \596_b0 );
buf ( \598_b1 , \576_b1 );
not ( \598_b1 , w_1686 );
not ( \598_b0 , w_1687 );
and ( w_1686 , w_1687 , \576_b0 );
or ( \599_b1 , \598_b1 , w_1689 );
not ( w_1689 , w_1690 );
and ( \599_b0 , \598_b0 , w_1691 );
and ( w_1690 ,  , w_1691 );
buf ( w_1689 , \574_b1 );
not ( w_1689 , w_1692 );
not (  , w_1693 );
and ( w_1692 , w_1693 , \574_b0 );
or ( \600_b1 , \483_b1 , \540_b1 );
xor ( \600_b0 , \483_b0 , w_1694 );
not ( w_1694 , w_1695 );
and ( w_1695 , \540_b1 , \540_b0 );
or ( \601_b1 , \599_b1 , \600_b1 );
xor ( \601_b0 , \599_b0 , w_1696 );
not ( w_1696 , w_1697 );
and ( w_1697 , \600_b1 , \600_b0 );
buf ( \602_b1 , \592_b1 );
not ( \602_b1 , w_1698 );
not ( \602_b0 , w_1699 );
and ( w_1698 , w_1699 , \592_b0 );
buf ( \603_b1 , \589_b1 );
not ( \603_b1 , w_1700 );
not ( \603_b0 , w_1701 );
and ( w_1700 , w_1701 , \589_b0 );
or ( \604_b1 , \602_b1 , w_1702 );
or ( \604_b0 , \602_b0 , \603_b0 );
not ( \603_b0 , w_1703 );
and ( w_1703 , w_1702 , \603_b1 );
or ( \605_b1 , \604_b1 , w_1705 );
not ( w_1705 , w_1706 );
and ( \605_b0 , \604_b0 , w_1707 );
and ( w_1706 ,  , w_1707 );
buf ( w_1705 , \590_b1 );
not ( w_1705 , w_1708 );
not (  , w_1709 );
and ( w_1708 , w_1709 , \590_b0 );
or ( \606_b1 , \589_b1 , w_1710 );
or ( \606_b0 , \589_b0 , \592_b0 );
not ( \592_b0 , w_1711 );
and ( w_1711 , w_1710 , \592_b1 );
or ( \607_b1 , \605_b1 , w_1713 );
not ( w_1713 , w_1714 );
and ( \607_b0 , \605_b0 , w_1715 );
and ( w_1714 ,  , w_1715 );
buf ( w_1713 , \606_b1 );
not ( w_1713 , w_1716 );
not (  , w_1717 );
and ( w_1716 , w_1717 , \606_b0 );
or ( \608_b1 , \601_b1 , \607_b1 );
xor ( \608_b0 , \601_b0 , w_1718 );
not ( w_1718 , w_1719 );
and ( w_1719 , \607_b1 , \607_b0 );
buf ( \609_b1 , \608_b1 );
not ( \609_b1 , w_1720 );
not ( \609_b0 , w_1721 );
and ( w_1720 , w_1721 , \608_b0 );
or ( \610_b1 , \597_b1 , \609_b1 );
not ( \609_b1 , w_1722 );
and ( \610_b0 , \597_b0 , w_1723 );
and ( w_1722 , w_1723 , \609_b0 );
or ( \611_b1 , \596_b1 , \608_b1 );
not ( \608_b1 , w_1724 );
and ( \611_b0 , \596_b0 , w_1725 );
and ( w_1724 , w_1725 , \608_b0 );
or ( \612_b1 , \610_b1 , w_1727 );
not ( w_1727 , w_1728 );
and ( \612_b0 , \610_b0 , w_1729 );
and ( w_1728 ,  , w_1729 );
buf ( w_1727 , \611_b1 );
not ( w_1727 , w_1730 );
not (  , w_1731 );
and ( w_1730 , w_1731 , \611_b0 );
or ( \613_b1 , \80_b1 , w_1733 );
not ( w_1733 , w_1734 );
and ( \613_b0 , \80_b0 , w_1735 );
and ( w_1734 ,  , w_1735 );
buf ( w_1733 , \B[2]_b1 );
not ( w_1733 , w_1736 );
not (  , w_1737 );
and ( w_1736 , w_1737 , \B[2]_b0 );
or ( \614_b1 , \253_b1 , w_1739 );
not ( w_1739 , w_1740 );
and ( \614_b0 , \253_b0 , w_1741 );
and ( w_1740 ,  , w_1741 );
buf ( w_1739 , \B[5]_b1 );
not ( w_1739 , w_1742 );
not (  , w_1743 );
and ( w_1742 , w_1743 , \B[5]_b0 );
or ( \615_b1 , \613_b1 , \614_b1 );
xor ( \615_b0 , \613_b0 , w_1744 );
not ( w_1744 , w_1745 );
and ( w_1745 , \614_b1 , \614_b0 );
or ( \616_b1 , \289_b1 , w_1747 );
not ( w_1747 , w_1748 );
and ( \616_b0 , \289_b0 , w_1749 );
and ( w_1748 ,  , w_1749 );
buf ( w_1747 , \B[6]_b1 );
not ( w_1747 , w_1750 );
not (  , w_1751 );
and ( w_1750 , w_1751 , \B[6]_b0 );
or ( \617_b1 , \615_b1 , \616_b1 );
xor ( \617_b0 , \615_b0 , w_1752 );
not ( w_1752 , w_1753 );
and ( w_1753 , \616_b1 , \616_b0 );
buf ( \618_b1 , \617_b1 );
not ( \618_b1 , w_1754 );
not ( \618_b0 , w_1755 );
and ( w_1754 , w_1755 , \617_b0 );
buf ( \619_b1 , \618_b1 );
not ( \619_b1 , w_1756 );
not ( \619_b0 , w_1757 );
and ( w_1756 , w_1757 , \618_b0 );
or ( \620_b1 , \296_b1 , w_1759 );
not ( w_1759 , w_1760 );
and ( \620_b0 , \296_b0 , w_1761 );
and ( w_1760 ,  , w_1761 );
buf ( w_1759 , \B[7]_b1 );
not ( w_1759 , w_1762 );
not (  , w_1763 );
and ( w_1762 , w_1763 , \B[7]_b0 );
or ( \621_b1 , \100_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_1764 );
and ( \621_b0 , \100_b0 , w_1765 );
and ( w_1764 , w_1765 , \B[3]_b0 );
or ( \622_b1 , \620_b1 , \621_b1 );
xor ( \622_b0 , \620_b0 , w_1766 );
not ( w_1766 , w_1767 );
and ( w_1767 , \621_b1 , \621_b0 );
or ( \623_b1 , \234_b1 , w_1769 );
not ( w_1769 , w_1770 );
and ( \623_b0 , \234_b0 , w_1771 );
and ( w_1770 ,  , w_1771 );
buf ( w_1769 , \B[4]_b1 );
not ( w_1769 , w_1772 );
not (  , w_1773 );
and ( w_1772 , w_1773 , \B[4]_b0 );
or ( \624_b1 , \622_b1 , w_1774 );
xor ( \624_b0 , \622_b0 , w_1776 );
not ( w_1776 , w_1777 );
and ( w_1777 , w_1774 , w_1775 );
buf ( w_1774 , \623_b1 );
not ( w_1774 , w_1778 );
not ( w_1775 , w_1779 );
and ( w_1778 , w_1779 , \623_b0 );
buf ( \625_b1 , \624_b1 );
not ( \625_b1 , w_1780 );
not ( \625_b0 , w_1781 );
and ( w_1780 , w_1781 , \624_b0 );
or ( \626_b1 , \619_b1 , w_1782 );
or ( \626_b0 , \619_b0 , \625_b0 );
not ( \625_b0 , w_1783 );
and ( w_1783 , w_1782 , \625_b1 );
buf ( \627_b1 , \624_b1 );
not ( \627_b1 , w_1784 );
not ( \627_b0 , w_1785 );
and ( w_1784 , w_1785 , \624_b0 );
or ( \628_b1 , \627_b1 , w_1787 );
not ( w_1787 , w_1788 );
and ( \628_b0 , \627_b0 , w_1789 );
and ( w_1788 ,  , w_1789 );
buf ( w_1787 , \617_b1 );
not ( w_1787 , w_1790 );
not (  , w_1791 );
and ( w_1790 , w_1791 , \617_b0 );
or ( \629_b1 , \626_b1 , w_1793 );
not ( w_1793 , w_1794 );
and ( \629_b0 , \626_b0 , w_1795 );
and ( w_1794 ,  , w_1795 );
buf ( w_1793 , \628_b1 );
not ( w_1793 , w_1796 );
not (  , w_1797 );
and ( w_1796 , w_1797 , \628_b0 );
or ( \630_b1 , \296_b1 , \B[6]_b1 );
not ( \B[6]_b1 , w_1798 );
and ( \630_b0 , \296_b0 , w_1799 );
and ( w_1798 , w_1799 , \B[6]_b0 );
buf ( \631_b1 , \630_b1 );
not ( \631_b1 , w_1800 );
not ( \631_b0 , w_1801 );
and ( w_1800 , w_1801 , \630_b0 );
or ( \632_b1 , \289_b1 , w_1803 );
not ( w_1803 , w_1804 );
and ( \632_b0 , \289_b0 , w_1805 );
and ( w_1804 ,  , w_1805 );
buf ( w_1803 , \B[5]_b1 );
not ( w_1803 , w_1806 );
not (  , w_1807 );
and ( w_1806 , w_1807 , \B[5]_b0 );
or ( \633_b1 , \631_b1 , w_1808 );
or ( \633_b0 , \631_b0 , \632_b0 );
not ( \632_b0 , w_1809 );
and ( w_1809 , w_1808 , \632_b1 );
buf ( \634_b1 , \632_b1 );
not ( \634_b1 , w_1810 );
not ( \634_b0 , w_1811 );
and ( w_1810 , w_1811 , \632_b0 );
buf ( \635_b1 , \631_b1 );
not ( \635_b1 , w_1812 );
not ( \635_b0 , w_1813 );
and ( w_1812 , w_1813 , \631_b0 );
or ( \636_b1 , \634_b1 , w_1814 );
or ( \636_b0 , \634_b0 , \635_b0 );
not ( \635_b0 , w_1815 );
and ( w_1815 , w_1814 , \635_b1 );
or ( \637_b1 , \100_b1 , w_1817 );
not ( w_1817 , w_1818 );
and ( \637_b0 , \100_b0 , w_1819 );
and ( w_1818 ,  , w_1819 );
buf ( w_1817 , \B[1]_b1 );
not ( w_1817 , w_1820 );
not (  , w_1821 );
and ( w_1820 , w_1821 , \B[1]_b0 );
buf ( \638_b1 , \637_b1 );
not ( \638_b1 , w_1822 );
not ( \638_b0 , w_1823 );
and ( w_1822 , w_1823 , \637_b0 );
or ( \639_b1 , \80_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_1824 );
and ( \639_b0 , \80_b0 , w_1825 );
and ( w_1824 , w_1825 , \B[0]_b0 );
or ( \640_b1 , \638_b1 , w_1827 );
not ( w_1827 , w_1828 );
and ( \640_b0 , \638_b0 , w_1829 );
and ( w_1828 ,  , w_1829 );
buf ( w_1827 , \639_b1 );
not ( w_1827 , w_1830 );
not (  , w_1831 );
and ( w_1830 , w_1831 , \639_b0 );
buf ( \641_b1 , \640_b1 );
not ( \641_b1 , w_1832 );
not ( \641_b0 , w_1833 );
and ( w_1832 , w_1833 , \640_b0 );
or ( \642_b1 , \636_b1 , w_1835 );
not ( w_1835 , w_1836 );
and ( \642_b0 , \636_b0 , w_1837 );
and ( w_1836 ,  , w_1837 );
buf ( w_1835 , \641_b1 );
not ( w_1835 , w_1838 );
not (  , w_1839 );
and ( w_1838 , w_1839 , \641_b0 );
or ( \643_b1 , \633_b1 , w_1841 );
not ( w_1841 , w_1842 );
and ( \643_b0 , \633_b0 , w_1843 );
and ( w_1842 ,  , w_1843 );
buf ( w_1841 , \642_b1 );
not ( w_1841 , w_1844 );
not (  , w_1845 );
and ( w_1844 , w_1845 , \642_b0 );
buf ( \644_b1 , \643_b1 );
not ( \644_b1 , w_1846 );
not ( \644_b0 , w_1847 );
and ( w_1846 , w_1847 , \643_b0 );
or ( \645_b1 , \629_b1 , \644_b1 );
not ( \644_b1 , w_1848 );
and ( \645_b0 , \629_b0 , w_1849 );
and ( w_1848 , w_1849 , \644_b0 );
buf ( \646_b1 , \629_b1 );
not ( \646_b1 , w_1850 );
not ( \646_b0 , w_1851 );
and ( w_1850 , w_1851 , \629_b0 );
or ( \647_b1 , \646_b1 , \643_b1 );
not ( \643_b1 , w_1852 );
and ( \647_b0 , \646_b0 , w_1853 );
and ( w_1852 , w_1853 , \643_b0 );
or ( \648_b1 , \645_b1 , w_1855 );
not ( w_1855 , w_1856 );
and ( \648_b0 , \645_b0 , w_1857 );
and ( w_1856 ,  , w_1857 );
buf ( w_1855 , \647_b1 );
not ( w_1855 , w_1858 );
not (  , w_1859 );
and ( w_1858 , w_1859 , \647_b0 );
buf ( \649_b1 , \648_b1 );
not ( \649_b1 , w_1860 );
not ( \649_b0 , w_1861 );
and ( w_1860 , w_1861 , \648_b0 );
or ( \650_b1 , \612_b1 , \649_b1 );
not ( \649_b1 , w_1862 );
and ( \650_b0 , \612_b0 , w_1863 );
and ( w_1862 , w_1863 , \649_b0 );
buf ( \651_b1 , \612_b1 );
not ( \651_b1 , w_1864 );
not ( \651_b0 , w_1865 );
and ( w_1864 , w_1865 , \612_b0 );
or ( \652_b1 , \651_b1 , \648_b1 );
not ( \648_b1 , w_1866 );
and ( \652_b0 , \651_b0 , w_1867 );
and ( w_1866 , w_1867 , \648_b0 );
or ( \653_b1 , \650_b1 , w_1869 );
not ( w_1869 , w_1870 );
and ( \653_b0 , \650_b0 , w_1871 );
and ( w_1870 ,  , w_1871 );
buf ( w_1869 , \652_b1 );
not ( w_1869 , w_1872 );
not (  , w_1873 );
and ( w_1872 , w_1873 , \652_b0 );
or ( \654_b1 , \630_b1 , \632_b1 );
xor ( \654_b0 , \630_b0 , w_1874 );
not ( w_1874 , w_1875 );
and ( w_1875 , \632_b1 , \632_b0 );
or ( \655_b1 , \654_b1 , w_1876 );
xor ( \655_b0 , \654_b0 , w_1878 );
not ( w_1878 , w_1879 );
and ( w_1879 , w_1876 , w_1877 );
buf ( w_1876 , \640_b1 );
not ( w_1876 , w_1880 );
not ( w_1877 , w_1881 );
and ( w_1880 , w_1881 , \640_b0 );
or ( \656_b1 , \296_b1 , w_1883 );
not ( w_1883 , w_1884 );
and ( \656_b0 , \296_b0 , w_1885 );
and ( w_1884 ,  , w_1885 );
buf ( w_1883 , \B[5]_b1 );
not ( w_1883 , w_1886 );
not (  , w_1887 );
and ( w_1886 , w_1887 , \B[5]_b0 );
or ( \657_b1 , \100_b1 , w_1889 );
not ( w_1889 , w_1890 );
and ( \657_b0 , \100_b0 , w_1891 );
and ( w_1890 ,  , w_1891 );
buf ( w_1889 , \B[0]_b1 );
not ( w_1889 , w_1892 );
not (  , w_1893 );
and ( w_1892 , w_1893 , \B[0]_b0 );
buf ( \658_b1 , \657_b1 );
not ( \658_b1 , w_1894 );
not ( \658_b0 , w_1895 );
and ( w_1894 , w_1895 , \657_b0 );
or ( \659_b1 , \233_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1896 );
and ( \659_b0 , \233_b0 , w_1897 );
and ( w_1896 , w_1897 , \B[1]_b0 );
or ( \660_b1 , \658_b1 , w_1899 );
not ( w_1899 , w_1900 );
and ( \660_b0 , \658_b0 , w_1901 );
and ( w_1900 ,  , w_1901 );
buf ( w_1899 , \659_b1 );
not ( w_1899 , w_1902 );
not (  , w_1903 );
and ( w_1902 , w_1903 , \659_b0 );
or ( \661_b1 , \656_b1 , \660_b1 );
xor ( \661_b0 , \656_b0 , w_1904 );
not ( w_1904 , w_1905 );
and ( w_1905 , \660_b1 , \660_b0 );
buf ( \662_b1 , \639_b1 );
not ( \662_b1 , w_1906 );
not ( \662_b0 , w_1907 );
and ( w_1906 , w_1907 , \639_b0 );
buf ( \663_b1 , \637_b1 );
not ( \663_b1 , w_1908 );
not ( \663_b0 , w_1909 );
and ( w_1908 , w_1909 , \637_b0 );
or ( \664_b1 , \662_b1 , \663_b1 );
not ( \663_b1 , w_1910 );
and ( \664_b0 , \662_b0 , w_1911 );
and ( w_1910 , w_1911 , \663_b0 );
or ( \665_b1 , \637_b1 , \639_b1 );
not ( \639_b1 , w_1912 );
and ( \665_b0 , \637_b0 , w_1913 );
and ( w_1912 , w_1913 , \639_b0 );
or ( \666_b1 , \664_b1 , w_1915 );
not ( w_1915 , w_1916 );
and ( \666_b0 , \664_b0 , w_1917 );
and ( w_1916 ,  , w_1917 );
buf ( w_1915 , \665_b1 );
not ( w_1915 , w_1918 );
not (  , w_1919 );
and ( w_1918 , w_1919 , \665_b0 );
or ( \667_b1 , \661_b1 , \666_b1 );
not ( \666_b1 , w_1920 );
and ( \667_b0 , \661_b0 , w_1921 );
and ( w_1920 , w_1921 , \666_b0 );
or ( \668_b1 , \656_b1 , \660_b1 );
not ( \660_b1 , w_1922 );
and ( \668_b0 , \656_b0 , w_1923 );
and ( w_1922 , w_1923 , \660_b0 );
or ( \669_b1 , \667_b1 , w_1924 );
or ( \669_b0 , \667_b0 , \668_b0 );
not ( \668_b0 , w_1925 );
and ( w_1925 , w_1924 , \668_b1 );
or ( \670_b1 , \655_b1 , \669_b1 );
xor ( \670_b0 , \655_b0 , w_1926 );
not ( w_1926 , w_1927 );
and ( w_1927 , \669_b1 , \669_b0 );
or ( \671_b1 , \580_b1 , \587_b1 );
xor ( \671_b0 , \580_b0 , w_1928 );
not ( w_1928 , w_1929 );
and ( w_1929 , \587_b1 , \587_b0 );
or ( \672_b1 , \671_b1 , \593_b1 );
xor ( \672_b0 , \671_b0 , w_1930 );
not ( w_1930 , w_1931 );
and ( w_1931 , \593_b1 , \593_b0 );
or ( \673_b1 , \670_b1 , \672_b1 );
not ( \672_b1 , w_1932 );
and ( \673_b0 , \670_b0 , w_1933 );
and ( w_1932 , w_1933 , \672_b0 );
or ( \674_b1 , \655_b1 , \669_b1 );
not ( \669_b1 , w_1934 );
and ( \674_b0 , \655_b0 , w_1935 );
and ( w_1934 , w_1935 , \669_b0 );
or ( \675_b1 , \673_b1 , w_1936 );
or ( \675_b0 , \673_b0 , \674_b0 );
not ( \674_b0 , w_1937 );
and ( w_1937 , w_1936 , \674_b1 );
or ( \676_b1 , \653_b1 , w_1939 );
not ( w_1939 , w_1940 );
and ( \676_b0 , \653_b0 , w_1941 );
and ( w_1940 ,  , w_1941 );
buf ( w_1939 , \675_b1 );
not ( w_1939 , w_1942 );
not (  , w_1943 );
and ( w_1942 , w_1943 , \675_b0 );
buf ( \677_b1 , \676_b1 );
not ( \677_b1 , w_1944 );
not ( \677_b0 , w_1945 );
and ( w_1944 , w_1945 , \676_b0 );
or ( \678_b1 , \655_b1 , \669_b1 );
xor ( \678_b0 , \655_b0 , w_1946 );
not ( w_1946 , w_1947 );
and ( w_1947 , \669_b1 , \669_b0 );
or ( \679_b1 , \678_b1 , \672_b1 );
xor ( \679_b0 , \678_b0 , w_1948 );
not ( w_1948 , w_1949 );
and ( w_1949 , \672_b1 , \672_b0 );
or ( \680_b1 , \296_b1 , w_1951 );
not ( w_1951 , w_1952 );
and ( \680_b0 , \296_b0 , w_1953 );
and ( w_1952 ,  , w_1953 );
buf ( w_1951 , \B[4]_b1 );
not ( w_1951 , w_1954 );
not (  , w_1955 );
and ( w_1954 , w_1955 , \B[4]_b0 );
or ( \681_b1 , \253_b1 , w_1957 );
not ( w_1957 , w_1958 );
and ( \681_b0 , \253_b0 , w_1959 );
and ( w_1958 ,  , w_1959 );
buf ( w_1957 , \B[2]_b1 );
not ( w_1957 , w_1960 );
not (  , w_1961 );
and ( w_1960 , w_1961 , \B[2]_b0 );
or ( \682_b1 , \680_b1 , \681_b1 );
xor ( \682_b0 , \680_b0 , w_1962 );
not ( w_1962 , w_1963 );
and ( w_1963 , \681_b1 , \681_b0 );
or ( \683_b1 , \289_b1 , w_1965 );
not ( w_1965 , w_1966 );
and ( \683_b0 , \289_b0 , w_1967 );
and ( w_1966 ,  , w_1967 );
buf ( w_1965 , \B[3]_b1 );
not ( w_1965 , w_1968 );
not (  , w_1969 );
and ( w_1968 , w_1969 , \B[3]_b0 );
or ( \684_b1 , \682_b1 , \683_b1 );
not ( \683_b1 , w_1970 );
and ( \684_b0 , \682_b0 , w_1971 );
and ( w_1970 , w_1971 , \683_b0 );
or ( \685_b1 , \680_b1 , \681_b1 );
not ( \681_b1 , w_1972 );
and ( \685_b0 , \680_b0 , w_1973 );
and ( w_1972 , w_1973 , \681_b0 );
or ( \686_b1 , \684_b1 , w_1974 );
or ( \686_b0 , \684_b0 , \685_b0 );
not ( \685_b0 , w_1975 );
and ( w_1975 , w_1974 , \685_b1 );
or ( \687_b1 , \581_b1 , \582_b1 );
xor ( \687_b0 , \581_b0 , w_1976 );
not ( w_1976 , w_1977 );
and ( w_1977 , \582_b1 , \582_b0 );
or ( \688_b1 , \687_b1 , \584_b1 );
xor ( \688_b0 , \687_b0 , w_1978 );
not ( w_1978 , w_1979 );
and ( w_1979 , \584_b1 , \584_b0 );
or ( \689_b1 , \686_b1 , \688_b1 );
xor ( \689_b0 , \686_b0 , w_1980 );
not ( w_1980 , w_1981 );
and ( w_1981 , \688_b1 , \688_b0 );
or ( \690_b1 , \656_b1 , \660_b1 );
xor ( \690_b0 , \656_b0 , w_1982 );
not ( w_1982 , w_1983 );
and ( w_1983 , \660_b1 , \660_b0 );
or ( \691_b1 , \690_b1 , \666_b1 );
xor ( \691_b0 , \690_b0 , w_1984 );
not ( w_1984 , w_1985 );
and ( w_1985 , \666_b1 , \666_b0 );
or ( \692_b1 , \689_b1 , \691_b1 );
not ( \691_b1 , w_1986 );
and ( \692_b0 , \689_b0 , w_1987 );
and ( w_1986 , w_1987 , \691_b0 );
or ( \693_b1 , \686_b1 , \688_b1 );
not ( \688_b1 , w_1988 );
and ( \693_b0 , \686_b0 , w_1989 );
and ( w_1988 , w_1989 , \688_b0 );
or ( \694_b1 , \692_b1 , w_1990 );
or ( \694_b0 , \692_b0 , \693_b0 );
not ( \693_b0 , w_1991 );
and ( w_1991 , w_1990 , \693_b1 );
or ( \695_b1 , \679_b1 , w_1993 );
not ( w_1993 , w_1994 );
and ( \695_b0 , \679_b0 , w_1995 );
and ( w_1994 ,  , w_1995 );
buf ( w_1993 , \694_b1 );
not ( w_1993 , w_1996 );
not (  , w_1997 );
and ( w_1996 , w_1997 , \694_b0 );
buf ( \696_b1 , \695_b1 );
not ( \696_b1 , w_1998 );
not ( \696_b0 , w_1999 );
and ( w_1998 , w_1999 , \695_b0 );
or ( \697_b1 , \686_b1 , \688_b1 );
xor ( \697_b0 , \686_b0 , w_2000 );
not ( w_2000 , w_2001 );
and ( w_2001 , \688_b1 , \688_b0 );
or ( \698_b1 , \697_b1 , \691_b1 );
xor ( \698_b0 , \697_b0 , w_2002 );
not ( w_2002 , w_2003 );
and ( w_2003 , \691_b1 , \691_b0 );
or ( \699_b1 , \234_b1 , w_2005 );
not ( w_2005 , w_2006 );
and ( \699_b0 , \234_b0 , w_2007 );
and ( w_2006 ,  , w_2007 );
buf ( w_2005 , \B[0]_b1 );
not ( w_2005 , w_2008 );
not (  , w_2009 );
and ( w_2008 , w_2009 , \B[0]_b0 );
buf ( \700_b1 , \699_b1 );
not ( \700_b1 , w_2010 );
not ( \700_b0 , w_2011 );
and ( w_2010 , w_2011 , \699_b0 );
or ( \701_b1 , \253_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_2012 );
and ( \701_b0 , \253_b0 , w_2013 );
and ( w_2012 , w_2013 , \B[1]_b0 );
or ( \702_b1 , \700_b1 , w_2015 );
not ( w_2015 , w_2016 );
and ( \702_b0 , \700_b0 , w_2017 );
and ( w_2016 ,  , w_2017 );
buf ( w_2015 , \701_b1 );
not ( w_2015 , w_2018 );
not (  , w_2019 );
and ( w_2018 , w_2019 , \701_b0 );
buf ( \703_b1 , \659_b1 );
not ( \703_b1 , w_2020 );
not ( \703_b0 , w_2021 );
and ( w_2020 , w_2021 , \659_b0 );
buf ( \704_b1 , \657_b1 );
not ( \704_b1 , w_2022 );
not ( \704_b0 , w_2023 );
and ( w_2022 , w_2023 , \657_b0 );
or ( \705_b1 , \703_b1 , \704_b1 );
not ( \704_b1 , w_2024 );
and ( \705_b0 , \703_b0 , w_2025 );
and ( w_2024 , w_2025 , \704_b0 );
or ( \706_b1 , \659_b1 , \657_b1 );
not ( \657_b1 , w_2026 );
and ( \706_b0 , \659_b0 , w_2027 );
and ( w_2026 , w_2027 , \657_b0 );
or ( \707_b1 , \705_b1 , w_2029 );
not ( w_2029 , w_2030 );
and ( \707_b0 , \705_b0 , w_2031 );
and ( w_2030 ,  , w_2031 );
buf ( w_2029 , \706_b1 );
not ( w_2029 , w_2032 );
not (  , w_2033 );
and ( w_2032 , w_2033 , \706_b0 );
or ( \708_b1 , \702_b1 , \707_b1 );
xor ( \708_b0 , \702_b0 , w_2034 );
not ( w_2034 , w_2035 );
and ( w_2035 , \707_b1 , \707_b0 );
or ( \709_b1 , \680_b1 , \681_b1 );
xor ( \709_b0 , \680_b0 , w_2036 );
not ( w_2036 , w_2037 );
and ( w_2037 , \681_b1 , \681_b0 );
or ( \710_b1 , \709_b1 , \683_b1 );
xor ( \710_b0 , \709_b0 , w_2038 );
not ( w_2038 , w_2039 );
and ( w_2039 , \683_b1 , \683_b0 );
or ( \711_b1 , \708_b1 , \710_b1 );
not ( \710_b1 , w_2040 );
and ( \711_b0 , \708_b0 , w_2041 );
and ( w_2040 , w_2041 , \710_b0 );
or ( \712_b1 , \702_b1 , \707_b1 );
not ( \707_b1 , w_2042 );
and ( \712_b0 , \702_b0 , w_2043 );
and ( w_2042 , w_2043 , \707_b0 );
or ( \713_b1 , \711_b1 , w_2044 );
or ( \713_b0 , \711_b0 , \712_b0 );
not ( \712_b0 , w_2045 );
and ( w_2045 , w_2044 , \712_b1 );
or ( \714_b1 , \698_b1 , w_2047 );
not ( w_2047 , w_2048 );
and ( \714_b0 , \698_b0 , w_2049 );
and ( w_2048 ,  , w_2049 );
buf ( w_2047 , \713_b1 );
not ( w_2047 , w_2050 );
not (  , w_2051 );
and ( w_2050 , w_2051 , \713_b0 );
buf ( \715_b1 , \714_b1 );
not ( \715_b1 , w_2052 );
not ( \715_b0 , w_2053 );
and ( w_2052 , w_2053 , \714_b0 );
or ( \716_b1 , \702_b1 , \707_b1 );
xor ( \716_b0 , \702_b0 , w_2054 );
not ( w_2054 , w_2055 );
and ( w_2055 , \707_b1 , \707_b0 );
or ( \717_b1 , \716_b1 , \710_b1 );
xor ( \717_b0 , \716_b0 , w_2056 );
not ( w_2056 , w_2057 );
and ( w_2057 , \710_b1 , \710_b0 );
buf ( \718_b1 , \701_b1 );
not ( \718_b1 , w_2058 );
not ( \718_b0 , w_2059 );
and ( w_2058 , w_2059 , \701_b0 );
buf ( \719_b1 , \699_b1 );
not ( \719_b1 , w_2060 );
not ( \719_b0 , w_2061 );
and ( w_2060 , w_2061 , \699_b0 );
or ( \720_b1 , \718_b1 , \719_b1 );
not ( \719_b1 , w_2062 );
and ( \720_b0 , \718_b0 , w_2063 );
and ( w_2062 , w_2063 , \719_b0 );
or ( \721_b1 , \699_b1 , \701_b1 );
not ( \701_b1 , w_2064 );
and ( \721_b0 , \699_b0 , w_2065 );
and ( w_2064 , w_2065 , \701_b0 );
or ( \722_b1 , \720_b1 , w_2067 );
not ( w_2067 , w_2068 );
and ( \722_b0 , \720_b0 , w_2069 );
and ( w_2068 ,  , w_2069 );
buf ( w_2067 , \721_b1 );
not ( w_2067 , w_2070 );
not (  , w_2071 );
and ( w_2070 , w_2071 , \721_b0 );
buf ( \723_b1 , \722_b1 );
not ( \723_b1 , w_2072 );
not ( \723_b0 , w_2073 );
and ( w_2072 , w_2073 , \722_b0 );
or ( \724_b1 , \296_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_2074 );
and ( \724_b0 , \296_b0 , w_2075 );
and ( w_2074 , w_2075 , \B[3]_b0 );
buf ( \725_b1 , \724_b1 );
not ( \725_b1 , w_2076 );
not ( \725_b0 , w_2077 );
and ( w_2076 , w_2077 , \724_b0 );
or ( \726_b1 , \289_b1 , w_2079 );
not ( w_2079 , w_2080 );
and ( \726_b0 , \289_b0 , w_2081 );
and ( w_2080 ,  , w_2081 );
buf ( w_2079 , \B[2]_b1 );
not ( w_2079 , w_2082 );
not (  , w_2083 );
and ( w_2082 , w_2083 , \B[2]_b0 );
or ( \727_b1 , \725_b1 , w_2085 );
not ( w_2085 , w_2086 );
and ( \727_b0 , \725_b0 , w_2087 );
and ( w_2086 ,  , w_2087 );
buf ( w_2085 , \726_b1 );
not ( w_2085 , w_2088 );
not (  , w_2089 );
and ( w_2088 , w_2089 , \726_b0 );
or ( \728_b1 , \723_b1 , w_2091 );
not ( w_2091 , w_2092 );
and ( \728_b0 , \723_b0 , w_2093 );
and ( w_2092 ,  , w_2093 );
buf ( w_2091 , \727_b1 );
not ( w_2091 , w_2094 );
not (  , w_2095 );
and ( w_2094 , w_2095 , \727_b0 );
buf ( \729_b1 , \726_b1 );
not ( \729_b1 , w_2096 );
not ( \729_b0 , w_2097 );
and ( w_2096 , w_2097 , \726_b0 );
or ( \730_b1 , \729_b1 , w_2099 );
not ( w_2099 , w_2100 );
and ( \730_b0 , \729_b0 , w_2101 );
and ( w_2100 ,  , w_2101 );
buf ( w_2099 , \724_b1 );
not ( w_2099 , w_2102 );
not (  , w_2103 );
and ( w_2102 , w_2103 , \724_b0 );
or ( \731_b1 , \728_b1 , \730_b1 );
not ( \730_b1 , w_2104 );
and ( \731_b0 , \728_b0 , w_2105 );
and ( w_2104 , w_2105 , \730_b0 );
or ( \732_b1 , \717_b1 , w_2106 );
or ( \732_b0 , \717_b0 , \731_b0 );
not ( \731_b0 , w_2107 );
and ( w_2107 , w_2106 , \731_b1 );
or ( \733_b1 , \253_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_2108 );
and ( \733_b0 , \253_b0 , w_2109 );
and ( w_2108 , w_2109 , \B[0]_b0 );
or ( \734_b1 , \296_b1 , \B[2]_b1 );
not ( \B[2]_b1 , w_2110 );
and ( \734_b0 , \296_b0 , w_2111 );
and ( w_2110 , w_2111 , \B[2]_b0 );
or ( \735_b1 , \733_b1 , \734_b1 );
not ( \734_b1 , w_2112 );
and ( \735_b0 , \733_b0 , w_2113 );
and ( w_2112 , w_2113 , \734_b0 );
buf ( \736_b1 , \735_b1 );
not ( \736_b1 , w_2114 );
not ( \736_b0 , w_2115 );
and ( w_2114 , w_2115 , \735_b0 );
buf ( \737_b1 , \722_b1 );
not ( \737_b1 , w_2116 );
not ( \737_b0 , w_2117 );
and ( w_2116 , w_2117 , \722_b0 );
buf ( \738_b1 , \726_b1 );
not ( \738_b1 , w_2118 );
not ( \738_b0 , w_2119 );
and ( w_2118 , w_2119 , \726_b0 );
buf ( \739_b1 , \724_b1 );
not ( \739_b1 , w_2120 );
not ( \739_b0 , w_2121 );
and ( w_2120 , w_2121 , \724_b0 );
or ( \740_b1 , \738_b1 , w_2122 );
or ( \740_b0 , \738_b0 , \739_b0 );
not ( \739_b0 , w_2123 );
and ( w_2123 , w_2122 , \739_b1 );
or ( \741_b1 , \724_b1 , w_2124 );
or ( \741_b0 , \724_b0 , \726_b0 );
not ( \726_b0 , w_2125 );
and ( w_2125 , w_2124 , \726_b1 );
or ( \742_b1 , \740_b1 , w_2127 );
not ( w_2127 , w_2128 );
and ( \742_b0 , \740_b0 , w_2129 );
and ( w_2128 ,  , w_2129 );
buf ( w_2127 , \741_b1 );
not ( w_2127 , w_2130 );
not (  , w_2131 );
and ( w_2130 , w_2131 , \741_b0 );
buf ( \743_b1 , \742_b1 );
not ( \743_b1 , w_2132 );
not ( \743_b0 , w_2133 );
and ( w_2132 , w_2133 , \742_b0 );
or ( \744_b1 , \737_b1 , \743_b1 );
not ( \743_b1 , w_2134 );
and ( \744_b0 , \737_b0 , w_2135 );
and ( w_2134 , w_2135 , \743_b0 );
or ( \745_b1 , \742_b1 , \722_b1 );
not ( \722_b1 , w_2136 );
and ( \745_b0 , \742_b0 , w_2137 );
and ( w_2136 , w_2137 , \722_b0 );
or ( \746_b1 , \744_b1 , w_2139 );
not ( w_2139 , w_2140 );
and ( \746_b0 , \744_b0 , w_2141 );
and ( w_2140 ,  , w_2141 );
buf ( w_2139 , \745_b1 );
not ( w_2139 , w_2142 );
not (  , w_2143 );
and ( w_2142 , w_2143 , \745_b0 );
or ( \747_b1 , \736_b1 , w_2145 );
not ( w_2145 , w_2146 );
and ( \747_b0 , \736_b0 , w_2147 );
and ( w_2146 ,  , w_2147 );
buf ( w_2145 , \746_b1 );
not ( w_2145 , w_2148 );
not (  , w_2149 );
and ( w_2148 , w_2149 , \746_b0 );
buf ( \748_b1 , \747_b1 );
not ( \748_b1 , w_2150 );
not ( \748_b0 , w_2151 );
and ( w_2150 , w_2151 , \747_b0 );
or ( \749_b1 , \289_b1 , w_2153 );
not ( w_2153 , w_2154 );
and ( \749_b0 , \289_b0 , w_2155 );
and ( w_2154 ,  , w_2155 );
buf ( w_2153 , \B[1]_b1 );
not ( w_2153 , w_2156 );
not (  , w_2157 );
and ( w_2156 , w_2157 , \B[1]_b0 );
buf ( \750_b1 , \749_b1 );
not ( \750_b1 , w_2158 );
not ( \750_b0 , w_2159 );
and ( w_2158 , w_2159 , \749_b0 );
or ( \751_b1 , \296_b1 , w_2161 );
not ( w_2161 , w_2162 );
and ( \751_b0 , \296_b0 , w_2163 );
and ( w_2162 ,  , w_2163 );
buf ( w_2161 , \B[0]_b1 );
not ( w_2161 , w_2164 );
not (  , w_2165 );
and ( w_2164 , w_2165 , \B[0]_b0 );
or ( \752_b1 , \749_b1 , w_2167 );
not ( w_2167 , w_2168 );
and ( \752_b0 , \749_b0 , w_2169 );
and ( w_2168 ,  , w_2169 );
buf ( w_2167 , \751_b1 );
not ( w_2167 , w_2170 );
not (  , w_2171 );
and ( w_2170 , w_2171 , \751_b0 );
or ( \753_b1 , \750_b1 , \752_b1 );
xor ( \753_b0 , \750_b0 , w_2172 );
not ( w_2172 , w_2173 );
and ( w_2173 , \752_b1 , \752_b0 );
or ( \754_b1 , \733_b1 , \734_b1 );
xor ( \754_b0 , \733_b0 , w_2174 );
not ( w_2174 , w_2175 );
and ( w_2175 , \734_b1 , \734_b0 );
or ( \755_b1 , \753_b1 , \754_b1 );
not ( \754_b1 , w_2176 );
and ( \755_b0 , \753_b0 , w_2177 );
and ( w_2176 , w_2177 , \754_b0 );
or ( \756_b1 , \750_b1 , \752_b1 );
not ( \752_b1 , w_2178 );
and ( \756_b0 , \750_b0 , w_2179 );
and ( w_2178 , w_2179 , \752_b0 );
or ( \757_b1 , \755_b1 , w_2180 );
or ( \757_b0 , \755_b0 , \756_b0 );
not ( \756_b0 , w_2181 );
and ( w_2181 , w_2180 , \756_b1 );
buf ( \758_b1 , \757_b1 );
not ( \758_b1 , w_2182 );
not ( \758_b0 , w_2183 );
and ( w_2182 , w_2183 , \757_b0 );
or ( \759_b1 , \748_b1 , w_2184 );
or ( \759_b0 , \748_b0 , \758_b0 );
not ( \758_b0 , w_2185 );
and ( w_2185 , w_2184 , \758_b1 );
buf ( \760_b1 , \746_b1 );
not ( \760_b1 , w_2186 );
not ( \760_b0 , w_2187 );
and ( w_2186 , w_2187 , \746_b0 );
or ( \761_b1 , \760_b1 , w_2189 );
not ( w_2189 , w_2190 );
and ( \761_b0 , \760_b0 , w_2191 );
and ( w_2190 ,  , w_2191 );
buf ( w_2189 , \735_b1 );
not ( w_2189 , w_2192 );
not (  , w_2193 );
and ( w_2192 , w_2193 , \735_b0 );
or ( \762_b1 , \759_b1 , w_2195 );
not ( w_2195 , w_2196 );
and ( \762_b0 , \759_b0 , w_2197 );
and ( w_2196 ,  , w_2197 );
buf ( w_2195 , \761_b1 );
not ( w_2195 , w_2198 );
not (  , w_2199 );
and ( w_2198 , w_2199 , \761_b0 );
or ( \763_b1 , \717_b1 , w_2201 );
not ( w_2201 , w_2202 );
and ( \763_b0 , \717_b0 , w_2203 );
and ( w_2202 ,  , w_2203 );
buf ( w_2201 , \731_b1 );
not ( w_2201 , w_2204 );
not (  , w_2205 );
and ( w_2204 , w_2205 , \731_b0 );
or ( \764_b1 , \762_b1 , w_2207 );
not ( w_2207 , w_2208 );
and ( \764_b0 , \762_b0 , w_2209 );
and ( w_2208 ,  , w_2209 );
buf ( w_2207 , \763_b1 );
not ( w_2207 , w_2210 );
not (  , w_2211 );
and ( w_2210 , w_2211 , \763_b0 );
or ( \765_b1 , \732_b1 , w_2213 );
not ( w_2213 , w_2214 );
and ( \765_b0 , \732_b0 , w_2215 );
and ( w_2214 ,  , w_2215 );
buf ( w_2213 , \764_b1 );
not ( w_2213 , w_2216 );
not (  , w_2217 );
and ( w_2216 , w_2217 , \764_b0 );
buf ( \766_b1 , \765_b1 );
not ( \766_b1 , w_2218 );
not ( \766_b0 , w_2219 );
and ( w_2218 , w_2219 , \765_b0 );
or ( \767_b1 , \715_b1 , w_2220 );
or ( \767_b0 , \715_b0 , \766_b0 );
not ( \766_b0 , w_2221 );
and ( w_2221 , w_2220 , \766_b1 );
or ( \768_b1 , \698_b1 , w_2222 );
or ( \768_b0 , \698_b0 , \713_b0 );
not ( \713_b0 , w_2223 );
and ( w_2223 , w_2222 , \713_b1 );
or ( \769_b1 , \767_b1 , w_2225 );
not ( w_2225 , w_2226 );
and ( \769_b0 , \767_b0 , w_2227 );
and ( w_2226 ,  , w_2227 );
buf ( w_2225 , \768_b1 );
not ( w_2225 , w_2228 );
not (  , w_2229 );
and ( w_2228 , w_2229 , \768_b0 );
buf ( \770_b1 , \769_b1 );
not ( \770_b1 , w_2230 );
not ( \770_b0 , w_2231 );
and ( w_2230 , w_2231 , \769_b0 );
or ( \771_b1 , \696_b1 , w_2232 );
or ( \771_b0 , \696_b0 , \770_b0 );
not ( \770_b0 , w_2233 );
and ( w_2233 , w_2232 , \770_b1 );
buf ( \772_b1 , \679_b1 );
not ( \772_b1 , w_2234 );
not ( \772_b0 , w_2235 );
and ( w_2234 , w_2235 , \679_b0 );
buf ( \773_b1 , \694_b1 );
not ( \773_b1 , w_2236 );
not ( \773_b0 , w_2237 );
and ( w_2236 , w_2237 , \694_b0 );
or ( \774_b1 , \772_b1 , w_2239 );
not ( w_2239 , w_2240 );
and ( \774_b0 , \772_b0 , w_2241 );
and ( w_2240 ,  , w_2241 );
buf ( w_2239 , \773_b1 );
not ( w_2239 , w_2242 );
not (  , w_2243 );
and ( w_2242 , w_2243 , \773_b0 );
or ( \775_b1 , \771_b1 , w_2245 );
not ( w_2245 , w_2246 );
and ( \775_b0 , \771_b0 , w_2247 );
and ( w_2246 ,  , w_2247 );
buf ( w_2245 , \774_b1 );
not ( w_2245 , w_2248 );
not (  , w_2249 );
and ( w_2248 , w_2249 , \774_b0 );
buf ( \776_b1 , \775_b1 );
not ( \776_b1 , w_2250 );
not ( \776_b0 , w_2251 );
and ( w_2250 , w_2251 , \775_b0 );
or ( \777_b1 , \677_b1 , w_2252 );
or ( \777_b0 , \677_b0 , \776_b0 );
not ( \776_b0 , w_2253 );
and ( w_2253 , w_2252 , \776_b1 );
buf ( \778_b1 , \653_b1 );
not ( \778_b1 , w_2254 );
not ( \778_b0 , w_2255 );
and ( w_2254 , w_2255 , \653_b0 );
buf ( \779_b1 , \675_b1 );
not ( \779_b1 , w_2256 );
not ( \779_b0 , w_2257 );
and ( w_2256 , w_2257 , \675_b0 );
or ( \780_b1 , \778_b1 , w_2259 );
not ( w_2259 , w_2260 );
and ( \780_b0 , \778_b0 , w_2261 );
and ( w_2260 ,  , w_2261 );
buf ( w_2259 , \779_b1 );
not ( w_2259 , w_2262 );
not (  , w_2263 );
and ( w_2262 , w_2263 , \779_b0 );
or ( \781_b1 , \777_b1 , w_2265 );
not ( w_2265 , w_2266 );
and ( \781_b0 , \777_b0 , w_2267 );
and ( w_2266 ,  , w_2267 );
buf ( w_2265 , \780_b1 );
not ( w_2265 , w_2268 );
not (  , w_2269 );
and ( w_2268 , w_2269 , \780_b0 );
buf ( \782_b1 , \617_b1 );
not ( \782_b1 , w_2270 );
not ( \782_b0 , w_2271 );
and ( w_2270 , w_2271 , \617_b0 );
buf ( \783_b1 , \624_b1 );
not ( \783_b1 , w_2272 );
not ( \783_b0 , w_2273 );
and ( w_2272 , w_2273 , \624_b0 );
or ( \784_b1 , \782_b1 , w_2274 );
or ( \784_b0 , \782_b0 , \783_b0 );
not ( \783_b0 , w_2275 );
and ( w_2275 , w_2274 , \783_b1 );
or ( \785_b1 , \784_b1 , w_2277 );
not ( w_2277 , w_2278 );
and ( \785_b0 , \784_b0 , w_2279 );
and ( w_2278 ,  , w_2279 );
buf ( w_2277 , \643_b1 );
not ( w_2277 , w_2280 );
not (  , w_2281 );
and ( w_2280 , w_2281 , \643_b0 );
or ( \786_b1 , \627_b1 , w_2283 );
not ( w_2283 , w_2284 );
and ( \786_b0 , \627_b0 , w_2285 );
and ( w_2284 ,  , w_2285 );
buf ( w_2283 , \618_b1 );
not ( w_2283 , w_2286 );
not (  , w_2287 );
and ( w_2286 , w_2287 , \618_b0 );
or ( \787_b1 , \785_b1 , w_2289 );
not ( w_2289 , w_2290 );
and ( \787_b0 , \785_b0 , w_2291 );
and ( w_2290 ,  , w_2291 );
buf ( w_2289 , \786_b1 );
not ( w_2289 , w_2292 );
not (  , w_2293 );
and ( w_2292 , w_2293 , \786_b0 );
buf ( \788_b1 , \623_b1 );
not ( \788_b1 , w_2294 );
not ( \788_b0 , w_2295 );
and ( w_2294 , w_2295 , \623_b0 );
buf ( \789_b1 , \620_b1 );
not ( \789_b1 , w_2296 );
not ( \789_b0 , w_2297 );
and ( w_2296 , w_2297 , \620_b0 );
or ( \790_b1 , \788_b1 , w_2298 );
or ( \790_b0 , \788_b0 , \789_b0 );
not ( \789_b0 , w_2299 );
and ( w_2299 , w_2298 , \789_b1 );
or ( \791_b1 , \790_b1 , w_2301 );
not ( w_2301 , w_2302 );
and ( \791_b0 , \790_b0 , w_2303 );
and ( w_2302 ,  , w_2303 );
buf ( w_2301 , \621_b1 );
not ( w_2301 , w_2304 );
not (  , w_2305 );
and ( w_2304 , w_2305 , \621_b0 );
or ( \792_b1 , \623_b1 , w_2306 );
or ( \792_b0 , \623_b0 , \620_b0 );
not ( \620_b0 , w_2307 );
and ( w_2307 , w_2306 , \620_b1 );
or ( \793_b1 , \791_b1 , w_2309 );
not ( w_2309 , w_2310 );
and ( \793_b0 , \791_b0 , w_2311 );
and ( w_2310 ,  , w_2311 );
buf ( w_2309 , \792_b1 );
not ( w_2309 , w_2312 );
not (  , w_2313 );
and ( w_2312 , w_2313 , \792_b0 );
buf ( \794_b1 , \614_b1 );
not ( \794_b1 , w_2314 );
not ( \794_b0 , w_2315 );
and ( w_2314 , w_2315 , \614_b0 );
buf ( \795_b1 , \616_b1 );
not ( \795_b1 , w_2316 );
not ( \795_b0 , w_2317 );
and ( w_2316 , w_2317 , \616_b0 );
or ( \796_b1 , \794_b1 , w_2318 );
or ( \796_b0 , \794_b0 , \795_b0 );
not ( \795_b0 , w_2319 );
and ( w_2319 , w_2318 , \795_b1 );
buf ( \797_b1 , \613_b1 );
not ( \797_b1 , w_2320 );
not ( \797_b0 , w_2321 );
and ( w_2320 , w_2321 , \613_b0 );
or ( \798_b1 , \796_b1 , w_2323 );
not ( w_2323 , w_2324 );
and ( \798_b0 , \796_b0 , w_2325 );
and ( w_2324 ,  , w_2325 );
buf ( w_2323 , \797_b1 );
not ( w_2323 , w_2326 );
not (  , w_2327 );
and ( w_2326 , w_2327 , \797_b0 );
or ( \799_b1 , \614_b1 , w_2328 );
or ( \799_b0 , \614_b0 , \616_b0 );
not ( \616_b0 , w_2329 );
and ( w_2329 , w_2328 , \616_b1 );
or ( \800_b1 , \798_b1 , w_2331 );
not ( w_2331 , w_2332 );
and ( \800_b0 , \798_b0 , w_2333 );
and ( w_2332 ,  , w_2333 );
buf ( w_2331 , \799_b1 );
not ( w_2331 , w_2334 );
not (  , w_2335 );
and ( w_2334 , w_2335 , \799_b0 );
or ( \801_b1 , \793_b1 , \800_b1 );
xor ( \801_b0 , \793_b0 , w_2336 );
not ( w_2336 , w_2337 );
and ( w_2337 , \800_b1 , \800_b0 );
or ( \802_b1 , \490_b1 , \487_b1 );
xor ( \802_b0 , \490_b0 , w_2338 );
not ( w_2338 , w_2339 );
and ( w_2339 , \487_b1 , \487_b0 );
buf ( \803_b1 , \485_b1 );
not ( \803_b1 , w_2340 );
not ( \803_b0 , w_2341 );
and ( w_2340 , w_2341 , \485_b0 );
or ( \804_b1 , \802_b1 , \803_b1 );
xor ( \804_b0 , \802_b0 , w_2342 );
not ( w_2342 , w_2343 );
and ( w_2343 , \803_b1 , \803_b0 );
buf ( \805_b1 , \804_b1 );
not ( \805_b1 , w_2344 );
not ( \805_b0 , w_2345 );
and ( w_2344 , w_2345 , \804_b0 );
or ( \806_b1 , \801_b1 , \805_b1 );
not ( \805_b1 , w_2346 );
and ( \806_b0 , \801_b0 , w_2347 );
and ( w_2346 , w_2347 , \805_b0 );
buf ( \807_b1 , \801_b1 );
not ( \807_b1 , w_2348 );
not ( \807_b0 , w_2349 );
and ( w_2348 , w_2349 , \801_b0 );
or ( \808_b1 , \807_b1 , \804_b1 );
not ( \804_b1 , w_2350 );
and ( \808_b0 , \807_b0 , w_2351 );
and ( w_2350 , w_2351 , \804_b0 );
or ( \809_b1 , \806_b1 , w_2353 );
not ( w_2353 , w_2354 );
and ( \809_b0 , \806_b0 , w_2355 );
and ( w_2354 ,  , w_2355 );
buf ( w_2353 , \808_b1 );
not ( w_2353 , w_2356 );
not (  , w_2357 );
and ( w_2356 , w_2357 , \808_b0 );
or ( \810_b1 , \787_b1 , \809_b1 );
xor ( \810_b0 , \787_b0 , w_2358 );
not ( w_2358 , w_2359 );
and ( w_2359 , \809_b1 , \809_b0 );
or ( \811_b1 , \499_b1 , \498_b1 );
xor ( \811_b0 , \499_b0 , w_2360 );
not ( w_2360 , w_2361 );
and ( w_2361 , \498_b1 , \498_b0 );
or ( \812_b1 , \811_b1 , \501_b1 );
xor ( \812_b0 , \811_b0 , w_2362 );
not ( w_2362 , w_2363 );
and ( w_2363 , \501_b1 , \501_b0 );
or ( \813_b1 , \531_b1 , \538_b1 );
xor ( \813_b0 , \531_b0 , w_2364 );
not ( w_2364 , w_2365 );
and ( w_2365 , \538_b1 , \538_b0 );
or ( \814_b1 , \813_b1 , \541_b1 );
xor ( \814_b0 , \813_b0 , w_2366 );
not ( w_2366 , w_2367 );
and ( w_2367 , \541_b1 , \541_b0 );
or ( \815_b1 , \812_b1 , \814_b1 );
xor ( \815_b0 , \812_b0 , w_2368 );
not ( w_2368 , w_2369 );
and ( w_2369 , \814_b1 , \814_b0 );
or ( \816_b1 , \599_b1 , \600_b1 );
xor ( \816_b0 , \599_b0 , w_2370 );
not ( w_2370 , w_2371 );
and ( w_2371 , \600_b1 , \600_b0 );
or ( \817_b1 , \816_b1 , \607_b1 );
not ( \607_b1 , w_2372 );
and ( \817_b0 , \816_b0 , w_2373 );
and ( w_2372 , w_2373 , \607_b0 );
or ( \818_b1 , \599_b1 , \600_b1 );
not ( \600_b1 , w_2374 );
and ( \818_b0 , \599_b0 , w_2375 );
and ( w_2374 , w_2375 , \600_b0 );
or ( \819_b1 , \817_b1 , w_2376 );
or ( \819_b0 , \817_b0 , \818_b0 );
not ( \818_b0 , w_2377 );
and ( w_2377 , w_2376 , \818_b1 );
or ( \820_b1 , \815_b1 , \819_b1 );
xor ( \820_b0 , \815_b0 , w_2378 );
not ( w_2378 , w_2379 );
and ( w_2379 , \819_b1 , \819_b0 );
or ( \821_b1 , \810_b1 , \820_b1 );
xor ( \821_b0 , \810_b0 , w_2380 );
not ( w_2380 , w_2381 );
and ( w_2381 , \820_b1 , \820_b0 );
buf ( \822_b1 , \821_b1 );
not ( \822_b1 , w_2382 );
not ( \822_b0 , w_2383 );
and ( w_2382 , w_2383 , \821_b0 );
buf ( \823_b1 , \608_b1 );
not ( \823_b1 , w_2384 );
not ( \823_b0 , w_2385 );
and ( w_2384 , w_2385 , \608_b0 );
buf ( \824_b1 , \649_b1 );
not ( \824_b1 , w_2386 );
not ( \824_b0 , w_2387 );
and ( w_2386 , w_2387 , \649_b0 );
or ( \825_b1 , \823_b1 , w_2388 );
or ( \825_b0 , \823_b0 , \824_b0 );
not ( \824_b0 , w_2389 );
and ( w_2389 , w_2388 , \824_b1 );
buf ( \826_b1 , \608_b1 );
not ( \826_b1 , w_2390 );
not ( \826_b0 , w_2391 );
and ( w_2390 , w_2391 , \608_b0 );
buf ( \827_b1 , \826_b1 );
not ( \827_b1 , w_2392 );
not ( \827_b0 , w_2393 );
and ( w_2392 , w_2393 , \826_b0 );
buf ( \828_b1 , \648_b1 );
not ( \828_b1 , w_2394 );
not ( \828_b0 , w_2395 );
and ( w_2394 , w_2395 , \648_b0 );
or ( \829_b1 , \827_b1 , w_2396 );
or ( \829_b0 , \827_b0 , \828_b0 );
not ( \828_b0 , w_2397 );
and ( w_2397 , w_2396 , \828_b1 );
buf ( \830_b1 , \596_b1 );
not ( \830_b1 , w_2398 );
not ( \830_b0 , w_2399 );
and ( w_2398 , w_2399 , \596_b0 );
or ( \831_b1 , \829_b1 , w_2401 );
not ( w_2401 , w_2402 );
and ( \831_b0 , \829_b0 , w_2403 );
and ( w_2402 ,  , w_2403 );
buf ( w_2401 , \830_b1 );
not ( w_2401 , w_2404 );
not (  , w_2405 );
and ( w_2404 , w_2405 , \830_b0 );
or ( \832_b1 , \825_b1 , w_2407 );
not ( w_2407 , w_2408 );
and ( \832_b0 , \825_b0 , w_2409 );
and ( w_2408 ,  , w_2409 );
buf ( w_2407 , \831_b1 );
not ( w_2407 , w_2410 );
not (  , w_2411 );
and ( w_2410 , w_2411 , \831_b0 );
buf ( \833_b1 , \832_b1 );
not ( \833_b1 , w_2412 );
not ( \833_b0 , w_2413 );
and ( w_2412 , w_2413 , \832_b0 );
or ( \834_b1 , \822_b1 , w_2415 );
not ( w_2415 , w_2416 );
and ( \834_b0 , \822_b0 , w_2417 );
and ( w_2416 ,  , w_2417 );
buf ( w_2415 , \833_b1 );
not ( w_2415 , w_2418 );
not (  , w_2419 );
and ( w_2418 , w_2419 , \833_b0 );
or ( \835_b1 , \781_b1 , w_2421 );
not ( w_2421 , w_2422 );
and ( \835_b0 , \781_b0 , w_2423 );
and ( w_2422 ,  , w_2423 );
buf ( w_2421 , \834_b1 );
not ( w_2421 , w_2424 );
not (  , w_2425 );
and ( w_2424 , w_2425 , \834_b0 );
or ( \836_b1 , \529_b1 , \526_b1 );
not ( \526_b1 , w_2426 );
and ( \836_b0 , \529_b0 , w_2427 );
and ( w_2426 , w_2427 , \526_b0 );
buf ( \837_b1 , \529_b1 );
not ( \837_b1 , w_2428 );
not ( \837_b0 , w_2429 );
and ( w_2428 , w_2429 , \529_b0 );
or ( \838_b1 , \837_b1 , \527_b1 );
not ( \527_b1 , w_2430 );
and ( \838_b0 , \837_b0 , w_2431 );
and ( w_2430 , w_2431 , \527_b0 );
or ( \839_b1 , \836_b1 , w_2432 );
or ( \839_b0 , \836_b0 , \838_b0 );
not ( \838_b0 , w_2433 );
and ( w_2433 , w_2432 , \838_b1 );
or ( \840_b1 , \839_b1 , \544_b1 );
xor ( \840_b0 , \839_b0 , w_2434 );
not ( w_2434 , w_2435 );
and ( w_2435 , \544_b1 , \544_b0 );
or ( \841_b1 , \812_b1 , \814_b1 );
xor ( \841_b0 , \812_b0 , w_2436 );
not ( w_2436 , w_2437 );
and ( w_2437 , \814_b1 , \814_b0 );
or ( \842_b1 , \841_b1 , \819_b1 );
not ( \819_b1 , w_2438 );
and ( \842_b0 , \841_b0 , w_2439 );
and ( w_2438 , w_2439 , \819_b0 );
or ( \843_b1 , \812_b1 , \814_b1 );
not ( \814_b1 , w_2440 );
and ( \843_b0 , \812_b0 , w_2441 );
and ( w_2440 , w_2441 , \814_b0 );
or ( \844_b1 , \842_b1 , w_2442 );
or ( \844_b0 , \842_b0 , \843_b0 );
not ( \843_b0 , w_2443 );
and ( w_2443 , w_2442 , \843_b1 );
or ( \845_b1 , \840_b1 , \844_b1 );
xor ( \845_b0 , \840_b0 , w_2444 );
not ( w_2444 , w_2445 );
and ( w_2445 , \844_b1 , \844_b0 );
or ( \846_b1 , \471_b1 , \472_b1 );
xor ( \846_b0 , \471_b0 , w_2446 );
not ( w_2446 , w_2447 );
and ( w_2447 , \472_b1 , \472_b0 );
or ( \847_b1 , \846_b1 , \478_b1 );
xor ( \847_b0 , \846_b0 , w_2448 );
not ( w_2448 , w_2449 );
and ( w_2449 , \478_b1 , \478_b0 );
or ( \848_b1 , \484_b1 , \496_b1 );
xor ( \848_b0 , \484_b0 , w_2450 );
not ( w_2450 , w_2451 );
and ( w_2451 , \496_b1 , \496_b0 );
or ( \849_b1 , \848_b1 , \504_b1 );
xor ( \849_b0 , \848_b0 , w_2452 );
not ( w_2452 , w_2453 );
and ( w_2453 , \504_b1 , \504_b0 );
or ( \850_b1 , \847_b1 , \849_b1 );
xor ( \850_b0 , \847_b0 , w_2454 );
not ( w_2454 , w_2455 );
and ( w_2455 , \849_b1 , \849_b0 );
or ( \851_b1 , \793_b1 , w_2456 );
or ( \851_b0 , \793_b0 , \800_b0 );
not ( \800_b0 , w_2457 );
and ( w_2457 , w_2456 , \800_b1 );
or ( \852_b1 , \851_b1 , \805_b1 );
not ( \805_b1 , w_2458 );
and ( \852_b0 , \851_b0 , w_2459 );
and ( w_2458 , w_2459 , \805_b0 );
or ( \853_b1 , \793_b1 , \800_b1 );
not ( \800_b1 , w_2460 );
and ( \853_b0 , \793_b0 , w_2461 );
and ( w_2460 , w_2461 , \800_b0 );
or ( \854_b1 , \852_b1 , w_2463 );
not ( w_2463 , w_2464 );
and ( \854_b0 , \852_b0 , w_2465 );
and ( w_2464 ,  , w_2465 );
buf ( w_2463 , \853_b1 );
not ( w_2463 , w_2466 );
not (  , w_2467 );
and ( w_2466 , w_2467 , \853_b0 );
or ( \855_b1 , \850_b1 , \854_b1 );
xor ( \855_b0 , \850_b0 , w_2468 );
not ( w_2468 , w_2469 );
and ( w_2469 , \854_b1 , \854_b0 );
buf ( \856_b1 , \855_b1 );
not ( \856_b1 , w_2470 );
not ( \856_b0 , w_2471 );
and ( w_2470 , w_2471 , \855_b0 );
or ( \857_b1 , \845_b1 , \856_b1 );
not ( \856_b1 , w_2472 );
and ( \857_b0 , \845_b0 , w_2473 );
and ( w_2472 , w_2473 , \856_b0 );
buf ( \858_b1 , \845_b1 );
not ( \858_b1 , w_2474 );
not ( \858_b0 , w_2475 );
and ( w_2474 , w_2475 , \845_b0 );
or ( \859_b1 , \858_b1 , \855_b1 );
not ( \855_b1 , w_2476 );
and ( \859_b0 , \858_b0 , w_2477 );
and ( w_2476 , w_2477 , \855_b0 );
or ( \860_b1 , \857_b1 , w_2479 );
not ( w_2479 , w_2480 );
and ( \860_b0 , \857_b0 , w_2481 );
and ( w_2480 ,  , w_2481 );
buf ( w_2479 , \859_b1 );
not ( w_2479 , w_2482 );
not (  , w_2483 );
and ( w_2482 , w_2483 , \859_b0 );
or ( \861_b1 , \787_b1 , \809_b1 );
xor ( \861_b0 , \787_b0 , w_2484 );
not ( w_2484 , w_2485 );
and ( w_2485 , \809_b1 , \809_b0 );
or ( \862_b1 , \861_b1 , \820_b1 );
not ( \820_b1 , w_2486 );
and ( \862_b0 , \861_b0 , w_2487 );
and ( w_2486 , w_2487 , \820_b0 );
or ( \863_b1 , \787_b1 , \809_b1 );
not ( \809_b1 , w_2488 );
and ( \863_b0 , \787_b0 , w_2489 );
and ( w_2488 , w_2489 , \809_b0 );
or ( \864_b1 , \862_b1 , w_2490 );
or ( \864_b0 , \862_b0 , \863_b0 );
not ( \863_b0 , w_2491 );
and ( w_2491 , w_2490 , \863_b1 );
or ( \865_b1 , \860_b1 , w_2493 );
not ( w_2493 , w_2494 );
and ( \865_b0 , \860_b0 , w_2495 );
and ( w_2494 ,  , w_2495 );
buf ( w_2493 , \864_b1 );
not ( w_2493 , w_2496 );
not (  , w_2497 );
and ( w_2496 , w_2497 , \864_b0 );
or ( \866_b1 , \821_b1 , w_2499 );
not ( w_2499 , w_2500 );
and ( \866_b0 , \821_b0 , w_2501 );
and ( w_2500 ,  , w_2501 );
buf ( w_2499 , \832_b1 );
not ( w_2499 , w_2502 );
not (  , w_2503 );
and ( w_2502 , w_2503 , \832_b0 );
or ( \867_b1 , \865_b1 , \866_b1 );
not ( \866_b1 , w_2504 );
and ( \867_b0 , \865_b0 , w_2505 );
and ( w_2504 , w_2505 , \866_b0 );
or ( \868_b1 , \835_b1 , w_2507 );
not ( w_2507 , w_2508 );
and ( \868_b0 , \835_b0 , w_2509 );
and ( w_2508 ,  , w_2509 );
buf ( w_2507 , \867_b1 );
not ( w_2507 , w_2510 );
not (  , w_2511 );
and ( w_2510 , w_2511 , \867_b0 );
buf ( \869_b1 , \868_b1 );
not ( \869_b1 , w_2512 );
not ( \869_b0 , w_2513 );
and ( w_2512 , w_2513 , \868_b0 );
or ( \870_b1 , \470_b1 , \481_b1 );
xor ( \870_b0 , \470_b0 , w_2514 );
not ( w_2514 , w_2515 );
and ( w_2515 , \481_b1 , \481_b0 );
or ( \871_b1 , \870_b1 , \507_b1 );
xor ( \871_b0 , \870_b0 , w_2516 );
not ( w_2516 , w_2517 );
and ( w_2517 , \507_b1 , \507_b0 );
buf ( \872_b1 , \871_b1 );
not ( \872_b1 , w_2518 );
not ( \872_b0 , w_2519 );
and ( w_2518 , w_2519 , \871_b0 );
or ( \873_b1 , \847_b1 , \849_b1 );
xor ( \873_b0 , \847_b0 , w_2520 );
not ( w_2520 , w_2521 );
and ( w_2521 , \849_b1 , \849_b0 );
or ( \874_b1 , \873_b1 , \854_b1 );
not ( \854_b1 , w_2522 );
and ( \874_b0 , \873_b0 , w_2523 );
and ( w_2522 , w_2523 , \854_b0 );
or ( \875_b1 , \847_b1 , \849_b1 );
not ( \849_b1 , w_2524 );
and ( \875_b0 , \847_b0 , w_2525 );
and ( w_2524 , w_2525 , \849_b0 );
or ( \876_b1 , \874_b1 , w_2526 );
or ( \876_b0 , \874_b0 , \875_b0 );
not ( \875_b0 , w_2527 );
and ( w_2527 , w_2526 , \875_b1 );
buf ( \877_b1 , \876_b1 );
not ( \877_b1 , w_2528 );
not ( \877_b0 , w_2529 );
and ( w_2528 , w_2529 , \876_b0 );
buf ( \878_b1 , \877_b1 );
not ( \878_b1 , w_2530 );
not ( \878_b0 , w_2531 );
and ( w_2530 , w_2531 , \877_b0 );
or ( \879_b1 , \872_b1 , w_2532 );
or ( \879_b0 , \872_b0 , \878_b0 );
not ( \878_b0 , w_2533 );
and ( w_2533 , w_2532 , \878_b1 );
buf ( \880_b1 , \871_b1 );
not ( \880_b1 , w_2534 );
not ( \880_b0 , w_2535 );
and ( w_2534 , w_2535 , \871_b0 );
or ( \881_b1 , \880_b1 , w_2537 );
not ( w_2537 , w_2538 );
and ( \881_b0 , \880_b0 , w_2539 );
and ( w_2538 ,  , w_2539 );
buf ( w_2537 , \876_b1 );
not ( w_2537 , w_2540 );
not (  , w_2541 );
and ( w_2540 , w_2541 , \876_b0 );
or ( \882_b1 , \879_b1 , w_2543 );
not ( w_2543 , w_2544 );
and ( \882_b0 , \879_b0 , w_2545 );
and ( w_2544 ,  , w_2545 );
buf ( w_2543 , \881_b1 );
not ( w_2543 , w_2546 );
not (  , w_2547 );
and ( w_2546 , w_2547 , \881_b0 );
or ( \883_b1 , \518_b1 , \520_b1 );
xor ( \883_b0 , \518_b0 , w_2548 );
not ( w_2548 , w_2549 );
and ( w_2549 , \520_b1 , \520_b0 );
or ( \884_b1 , \883_b1 , \547_b1 );
xor ( \884_b0 , \883_b0 , w_2550 );
not ( w_2550 , w_2551 );
and ( w_2551 , \547_b1 , \547_b0 );
or ( \885_b1 , \882_b1 , \884_b1 );
xor ( \885_b0 , \882_b0 , w_2552 );
not ( w_2552 , w_2553 );
and ( w_2553 , \884_b1 , \884_b0 );
or ( \886_b1 , \844_b1 , w_2554 );
or ( \886_b0 , \844_b0 , \840_b0 );
not ( \840_b0 , w_2555 );
and ( w_2555 , w_2554 , \840_b1 );
or ( \887_b1 , \856_b1 , \886_b1 );
not ( \886_b1 , w_2556 );
and ( \887_b0 , \856_b0 , w_2557 );
and ( w_2556 , w_2557 , \886_b0 );
or ( \888_b1 , \840_b1 , \844_b1 );
not ( \844_b1 , w_2558 );
and ( \888_b0 , \840_b0 , w_2559 );
and ( w_2558 , w_2559 , \844_b0 );
or ( \889_b1 , \887_b1 , w_2561 );
not ( w_2561 , w_2562 );
and ( \889_b0 , \887_b0 , w_2563 );
and ( w_2562 ,  , w_2563 );
buf ( w_2561 , \888_b1 );
not ( w_2561 , w_2564 );
not (  , w_2565 );
and ( w_2564 , w_2565 , \888_b0 );
or ( \890_b1 , \885_b1 , w_2567 );
not ( w_2567 , w_2568 );
and ( \890_b0 , \885_b0 , w_2569 );
and ( w_2568 ,  , w_2569 );
buf ( w_2567 , \889_b1 );
not ( w_2567 , w_2570 );
not (  , w_2571 );
and ( w_2570 , w_2571 , \889_b0 );
buf ( \891_b1 , \860_b1 );
not ( \891_b1 , w_2572 );
not ( \891_b0 , w_2573 );
and ( w_2572 , w_2573 , \860_b0 );
buf ( \892_b1 , \864_b1 );
not ( \892_b1 , w_2574 );
not ( \892_b0 , w_2575 );
and ( w_2574 , w_2575 , \864_b0 );
or ( \893_b1 , \891_b1 , w_2577 );
not ( w_2577 , w_2578 );
and ( \893_b0 , \891_b0 , w_2579 );
and ( w_2578 ,  , w_2579 );
buf ( w_2577 , \892_b1 );
not ( w_2577 , w_2580 );
not (  , w_2581 );
and ( w_2580 , w_2581 , \892_b0 );
or ( \894_b1 , \890_b1 , w_2583 );
not ( w_2583 , w_2584 );
and ( \894_b0 , \890_b0 , w_2585 );
and ( w_2584 ,  , w_2585 );
buf ( w_2583 , \893_b1 );
not ( w_2583 , w_2586 );
not (  , w_2587 );
and ( w_2586 , w_2587 , \893_b0 );
or ( \895_b1 , \516_b1 , \550_b1 );
xor ( \895_b0 , \516_b0 , w_2588 );
not ( w_2588 , w_2589 );
and ( w_2589 , \550_b1 , \550_b0 );
or ( \896_b1 , \895_b1 , w_2590 );
xor ( \896_b0 , \895_b0 , w_2592 );
not ( w_2592 , w_2593 );
and ( w_2593 , w_2590 , w_2591 );
buf ( w_2590 , \553_b1 );
not ( w_2590 , w_2594 );
not ( w_2591 , w_2595 );
and ( w_2594 , w_2595 , \553_b0 );
buf ( \897_b1 , \871_b1 );
not ( \897_b1 , w_2596 );
not ( \897_b0 , w_2597 );
and ( w_2596 , w_2597 , \871_b0 );
buf ( \898_b1 , \884_b1 );
not ( \898_b1 , w_2598 );
not ( \898_b0 , w_2599 );
and ( w_2598 , w_2599 , \884_b0 );
or ( \899_b1 , \897_b1 , w_2600 );
or ( \899_b0 , \897_b0 , \898_b0 );
not ( \898_b0 , w_2601 );
and ( w_2601 , w_2600 , \898_b1 );
buf ( \900_b1 , \876_b1 );
not ( \900_b1 , w_2602 );
not ( \900_b0 , w_2603 );
and ( w_2602 , w_2603 , \876_b0 );
or ( \901_b1 , \899_b1 , w_2605 );
not ( w_2605 , w_2606 );
and ( \901_b0 , \899_b0 , w_2607 );
and ( w_2606 ,  , w_2607 );
buf ( w_2605 , \900_b1 );
not ( w_2605 , w_2608 );
not (  , w_2609 );
and ( w_2608 , w_2609 , \900_b0 );
buf ( \902_b1 , \871_b1 );
not ( \902_b1 , w_2610 );
not ( \902_b0 , w_2611 );
and ( w_2610 , w_2611 , \871_b0 );
buf ( \903_b1 , \884_b1 );
not ( \903_b1 , w_2612 );
not ( \903_b0 , w_2613 );
and ( w_2612 , w_2613 , \884_b0 );
or ( \904_b1 , \902_b1 , w_2615 );
not ( w_2615 , w_2616 );
and ( \904_b0 , \902_b0 , w_2617 );
and ( w_2616 ,  , w_2617 );
buf ( w_2615 , \903_b1 );
not ( w_2615 , w_2618 );
not (  , w_2619 );
and ( w_2618 , w_2619 , \903_b0 );
or ( \905_b1 , \901_b1 , w_2621 );
not ( w_2621 , w_2622 );
and ( \905_b0 , \901_b0 , w_2623 );
and ( w_2622 ,  , w_2623 );
buf ( w_2621 , \904_b1 );
not ( w_2621 , w_2624 );
not (  , w_2625 );
and ( w_2624 , w_2625 , \904_b0 );
or ( \906_b1 , \896_b1 , w_2627 );
not ( w_2627 , w_2628 );
and ( \906_b0 , \896_b0 , w_2629 );
and ( w_2628 ,  , w_2629 );
buf ( w_2627 , \905_b1 );
not ( w_2627 , w_2630 );
not (  , w_2631 );
and ( w_2630 , w_2631 , \905_b0 );
or ( \907_b1 , \894_b1 , w_2633 );
not ( w_2633 , w_2634 );
and ( \907_b0 , \894_b0 , w_2635 );
and ( w_2634 ,  , w_2635 );
buf ( w_2633 , \906_b1 );
not ( w_2633 , w_2636 );
not (  , w_2637 );
and ( w_2636 , w_2637 , \906_b0 );
buf ( \908_b1 , \907_b1 );
not ( \908_b1 , w_2638 );
not ( \908_b0 , w_2639 );
and ( w_2638 , w_2639 , \907_b0 );
or ( \909_b1 , \869_b1 , w_2640 );
or ( \909_b0 , \869_b0 , \908_b0 );
not ( \908_b0 , w_2641 );
and ( w_2641 , w_2640 , \908_b1 );
or ( \910_b1 , \516_b1 , \550_b1 );
xor ( \910_b0 , \516_b0 , w_2642 );
not ( w_2642 , w_2643 );
and ( w_2643 , \550_b1 , \550_b0 );
or ( \911_b1 , \910_b1 , \553_b1 );
xor ( \911_b0 , \910_b0 , w_2644 );
not ( w_2644 , w_2645 );
and ( w_2645 , \553_b1 , \553_b0 );
buf ( \912_b1 , \905_b1 );
not ( \912_b1 , w_2646 );
not ( \912_b0 , w_2647 );
and ( w_2646 , w_2647 , \905_b0 );
or ( \913_b1 , \911_b1 , w_2649 );
not ( w_2649 , w_2650 );
and ( \913_b0 , \911_b0 , w_2651 );
and ( w_2650 ,  , w_2651 );
buf ( w_2649 , \912_b1 );
not ( w_2649 , w_2652 );
not (  , w_2653 );
and ( w_2652 , w_2653 , \912_b0 );
or ( \914_b1 , \885_b1 , w_2655 );
not ( w_2655 , w_2656 );
and ( \914_b0 , \885_b0 , w_2657 );
and ( w_2656 ,  , w_2657 );
buf ( w_2655 , \889_b1 );
not ( w_2655 , w_2658 );
not (  , w_2659 );
and ( w_2658 , w_2659 , \889_b0 );
or ( \915_b1 , \913_b1 , \914_b1 );
not ( \914_b1 , w_2660 );
and ( \915_b0 , \913_b0 , w_2661 );
and ( w_2660 , w_2661 , \914_b0 );
or ( \916_b1 , \911_b1 , w_2663 );
not ( w_2663 , w_2664 );
and ( \916_b0 , \911_b0 , w_2665 );
and ( w_2664 ,  , w_2665 );
buf ( w_2663 , \912_b1 );
not ( w_2663 , w_2666 );
not (  , w_2667 );
and ( w_2666 , w_2667 , \912_b0 );
or ( \917_b1 , \915_b1 , w_2669 );
not ( w_2669 , w_2670 );
and ( \917_b0 , \915_b0 , w_2671 );
and ( w_2670 ,  , w_2671 );
buf ( w_2669 , \916_b1 );
not ( w_2669 , w_2672 );
not (  , w_2673 );
and ( w_2672 , w_2673 , \916_b0 );
or ( \918_b1 , \909_b1 , w_2675 );
not ( w_2675 , w_2676 );
and ( \918_b0 , \909_b0 , w_2677 );
and ( w_2676 ,  , w_2677 );
buf ( w_2675 , \917_b1 );
not ( w_2675 , w_2678 );
not (  , w_2679 );
and ( w_2678 , w_2679 , \917_b0 );
buf ( \919_b1 , \918_b1 );
not ( \919_b1 , w_2680 );
not ( \919_b0 , w_2681 );
and ( w_2680 , w_2681 , \918_b0 );
or ( \920_b1 , \573_b1 , w_2682 );
or ( \920_b0 , \573_b0 , \919_b0 );
not ( \919_b0 , w_2683 );
and ( w_2683 , w_2682 , \919_b1 );
buf ( \921_b1 , \570_b1 );
not ( \921_b1 , w_2684 );
not ( \921_b0 , w_2685 );
and ( w_2684 , w_2685 , \570_b0 );
or ( \922_b1 , \514_b1 , w_2687 );
not ( w_2687 , w_2688 );
and ( \922_b0 , \514_b0 , w_2689 );
and ( w_2688 ,  , w_2689 );
buf ( w_2687 , \556_b1 );
not ( w_2687 , w_2690 );
not (  , w_2691 );
and ( w_2690 , w_2691 , \556_b0 );
buf ( \923_b1 , \922_b1 );
not ( \923_b1 , w_2692 );
not ( \923_b0 , w_2693 );
and ( w_2692 , w_2693 , \922_b0 );
or ( \924_b1 , \921_b1 , w_2694 );
or ( \924_b0 , \921_b0 , \923_b0 );
not ( \923_b0 , w_2695 );
and ( w_2695 , w_2694 , \923_b1 );
buf ( \925_b1 , \569_b1 );
not ( \925_b1 , w_2696 );
not ( \925_b0 , w_2697 );
and ( w_2696 , w_2697 , \569_b0 );
or ( \926_b1 , \925_b1 , w_2699 );
not ( w_2699 , w_2700 );
and ( \926_b0 , \925_b0 , w_2701 );
and ( w_2700 ,  , w_2701 );
buf ( w_2699 , \566_b1 );
not ( w_2699 , w_2702 );
not (  , w_2703 );
and ( w_2702 , w_2703 , \566_b0 );
or ( \927_b1 , \924_b1 , w_2705 );
not ( w_2705 , w_2706 );
and ( \927_b0 , \924_b0 , w_2707 );
and ( w_2706 ,  , w_2707 );
buf ( w_2705 , \926_b1 );
not ( w_2705 , w_2708 );
not (  , w_2709 );
and ( w_2708 , w_2709 , \926_b0 );
or ( \928_b1 , \927_b1 , w_2711 );
not ( w_2711 , w_2712 );
and ( \928_b0 , \927_b0 , w_2713 );
and ( w_2712 ,  , w_2713 );
buf ( w_2711 , \425_b1 );
not ( w_2711 , w_2714 );
not (  , w_2715 );
and ( w_2714 , w_2715 , \425_b0 );
buf ( \929_b1 , \423_b1 );
not ( \929_b1 , w_2716 );
not ( \929_b0 , w_2717 );
and ( w_2716 , w_2717 , \423_b0 );
or ( \930_b1 , \395_b1 , w_2719 );
not ( w_2719 , w_2720 );
and ( \930_b0 , \395_b0 , w_2721 );
and ( w_2720 ,  , w_2721 );
buf ( w_2719 , \397_b1 );
not ( w_2719 , w_2722 );
not (  , w_2723 );
and ( w_2722 , w_2723 , \397_b0 );
or ( \931_b1 , \930_b1 , w_2725 );
not ( w_2725 , w_2726 );
and ( \931_b0 , \930_b0 , w_2727 );
and ( w_2726 ,  , w_2727 );
buf ( w_2725 , \271_b1 );
not ( w_2725 , w_2728 );
not (  , w_2729 );
and ( w_2728 , w_2729 , \271_b0 );
or ( \932_b1 , \931_b1 , w_2731 );
not ( w_2731 , w_2732 );
and ( \932_b0 , \931_b0 , w_2733 );
and ( w_2732 ,  , w_2733 );
buf ( w_2731 , \275_b1 );
not ( w_2731 , w_2734 );
not (  , w_2735 );
and ( w_2734 , w_2735 , \275_b0 );
or ( \933_b1 , \929_b1 , w_2737 );
not ( w_2737 , w_2738 );
and ( \933_b0 , \929_b0 , w_2739 );
and ( w_2738 ,  , w_2739 );
buf ( w_2737 , \932_b1 );
not ( w_2737 , w_2740 );
not (  , w_2741 );
and ( w_2740 , w_2741 , \932_b0 );
or ( \934_b1 , \420_b1 , w_2743 );
not ( w_2743 , w_2744 );
and ( \934_b0 , \420_b0 , w_2745 );
and ( w_2744 ,  , w_2745 );
buf ( w_2743 , \422_b1 );
not ( w_2743 , w_2746 );
not (  , w_2747 );
and ( w_2746 , w_2747 , \422_b0 );
or ( \935_b1 , \933_b1 , w_2748 );
or ( \935_b0 , \933_b0 , \934_b0 );
not ( \934_b0 , w_2749 );
and ( w_2749 , w_2748 , \934_b1 );
or ( \936_b1 , \935_b1 , w_2751 );
not ( w_2751 , w_2752 );
and ( \936_b0 , \935_b0 , w_2753 );
and ( w_2752 ,  , w_2753 );
buf ( w_2751 , \416_b1 );
not ( w_2751 , w_2754 );
not (  , w_2755 );
and ( w_2754 , w_2755 , \416_b0 );
or ( \937_b1 , \413_b1 , w_2756 );
or ( \937_b0 , \413_b0 , \415_b0 );
not ( \415_b0 , w_2757 );
and ( w_2757 , w_2756 , \415_b1 );
or ( \939_b1 , \920_b1 , w_2759 );
not ( w_2759 , w_2760 );
and ( \939_b0 , \920_b0 , w_2761 );
and ( w_2760 ,  , w_2761 );
buf ( w_2759 , \938_b1 );
not ( w_2759 , w_2762 );
not (  , w_2763 );
and ( w_2762 , w_2763 , \938_b0 );
buf ( \940_b1 , \939_b1 );
not ( \940_b1 , w_2764 );
not ( \940_b0 , w_2765 );
and ( w_2764 , w_2765 , \939_b0 );
or ( \941_b1 , \312_b1 , w_2766 );
or ( \941_b0 , \312_b0 , \940_b0 );
not ( \940_b0 , w_2767 );
and ( w_2767 , w_2766 , \940_b1 );
or ( \942_b1 , \309_b1 , w_2768 );
or ( \942_b0 , \309_b0 , \310_b0 );
not ( \310_b0 , w_2769 );
and ( w_2769 , w_2768 , \310_b1 );
or ( \943_b1 , \941_b1 , w_2771 );
not ( w_2771 , w_2772 );
and ( \943_b0 , \941_b0 , w_2773 );
and ( w_2772 ,  , w_2773 );
buf ( w_2771 , \942_b1 );
not ( w_2771 , w_2774 );
not (  , w_2775 );
and ( w_2774 , w_2775 , \942_b0 );
or ( \944_b1 , \311_b1 , w_2777 );
not ( w_2777 , w_2778 );
and ( \944_b0 , \311_b0 , w_2779 );
and ( w_2778 ,  , w_2779 );
buf ( w_2777 , \942_b1 );
not ( w_2777 , w_2780 );
not (  , w_2781 );
and ( w_2780 , w_2781 , \942_b0 );
buf ( \945_b1 , \944_b1 );
not ( \945_b1 , w_2782 );
not ( \945_b0 , w_2783 );
and ( w_2782 , w_2783 , \944_b0 );
buf ( \946_b1 , \939_b1 );
not ( \946_b1 , w_2784 );
not ( \946_b0 , w_2785 );
and ( w_2784 , w_2785 , \939_b0 );
or ( \947_b1 , \945_b1 , w_2786 );
or ( \947_b0 , \945_b0 , \946_b0 );
not ( \946_b0 , w_2787 );
and ( w_2787 , w_2786 , \946_b1 );
or ( \948_b1 , \944_b1 , w_2788 );
or ( \948_b0 , \944_b0 , \939_b0 );
not ( \939_b0 , w_2789 );
and ( w_2789 , w_2788 , \939_b1 );
or ( \949_b1 , \947_b1 , w_2791 );
not ( w_2791 , w_2792 );
and ( \949_b0 , \947_b0 , w_2793 );
and ( w_2792 ,  , w_2793 );
buf ( w_2791 , \948_b1 );
not ( w_2791 , w_2794 );
not (  , w_2795 );
and ( w_2794 , w_2795 , \948_b0 );
buf ( \950_b1 , \423_b1 );
not ( \950_b1 , w_2796 );
not ( \950_b0 , w_2797 );
and ( w_2796 , w_2797 , \423_b0 );
or ( \951_b1 , \571_b1 , w_2799 );
not ( w_2799 , w_2800 );
and ( \951_b0 , \571_b0 , w_2801 );
and ( w_2800 ,  , w_2801 );
buf ( w_2799 , \399_b1 );
not ( w_2799 , w_2802 );
not (  , w_2803 );
and ( w_2802 , w_2803 , \399_b0 );
buf ( \952_b1 , \951_b1 );
not ( \952_b1 , w_2804 );
not ( \952_b0 , w_2805 );
and ( w_2804 , w_2805 , \951_b0 );
buf ( \953_b1 , \918_b1 );
not ( \953_b1 , w_2806 );
not ( \953_b0 , w_2807 );
and ( w_2806 , w_2807 , \918_b0 );
or ( \954_b1 , \952_b1 , w_2808 );
or ( \954_b0 , \952_b0 , \953_b0 );
not ( \953_b0 , w_2809 );
and ( w_2809 , w_2808 , \953_b1 );
or ( \955_b1 , \398_b1 , \272_b1 );
not ( \272_b1 , w_2810 );
and ( \955_b0 , \398_b0 , w_2811 );
and ( w_2810 , w_2811 , \272_b0 );
or ( \956_b1 , \927_b1 , \955_b1 );
not ( \955_b1 , w_2812 );
and ( \956_b0 , \927_b0 , w_2813 );
and ( w_2812 , w_2813 , \955_b0 );
buf ( \957_b1 , \932_b1 );
not ( \957_b1 , w_2814 );
not ( \957_b0 , w_2815 );
and ( w_2814 , w_2815 , \932_b0 );
or ( \958_b1 , \956_b1 , w_2817 );
not ( w_2817 , w_2818 );
and ( \958_b0 , \956_b0 , w_2819 );
and ( w_2818 ,  , w_2819 );
buf ( w_2817 , \957_b1 );
not ( w_2817 , w_2820 );
not (  , w_2821 );
and ( w_2820 , w_2821 , \957_b0 );
or ( \959_b1 , \954_b1 , w_2823 );
not ( w_2823 , w_2824 );
and ( \959_b0 , \954_b0 , w_2825 );
and ( w_2824 ,  , w_2825 );
buf ( w_2823 , \958_b1 );
not ( w_2823 , w_2826 );
not (  , w_2827 );
and ( w_2826 , w_2827 , \958_b0 );
buf ( \960_b1 , \959_b1 );
not ( \960_b1 , w_2828 );
not ( \960_b0 , w_2829 );
and ( w_2828 , w_2829 , \959_b0 );
or ( \961_b1 , \950_b1 , w_2830 );
or ( \961_b0 , \950_b0 , \960_b0 );
not ( \960_b0 , w_2831 );
and ( w_2831 , w_2830 , \960_b1 );
buf ( \962_b1 , \934_b1 );
not ( \962_b1 , w_2832 );
not ( \962_b0 , w_2833 );
and ( w_2832 , w_2833 , \934_b0 );
or ( \963_b1 , \961_b1 , w_2835 );
not ( w_2835 , w_2836 );
and ( \963_b0 , \961_b0 , w_2837 );
and ( w_2836 ,  , w_2837 );
buf ( w_2835 , \962_b1 );
not ( w_2835 , w_2838 );
not (  , w_2839 );
and ( w_2838 , w_2839 , \962_b0 );
or ( \964_b1 , \416_b1 , w_2841 );
not ( w_2841 , w_2842 );
and ( \964_b0 , \416_b0 , w_2843 );
and ( w_2842 ,  , w_2843 );
buf ( w_2841 , \937_b1 );
not ( w_2841 , w_2844 );
not (  , w_2845 );
and ( w_2844 , w_2845 , \937_b0 );
buf ( \965_b1 , \964_b1 );
not ( \965_b1 , w_2846 );
not ( \965_b0 , w_2847 );
and ( w_2846 , w_2847 , \964_b0 );
or ( \966_b1 , \963_b1 , \965_b1 );
not ( \965_b1 , w_2848 );
and ( \966_b0 , \963_b0 , w_2849 );
and ( w_2848 , w_2849 , \965_b0 );
buf ( \967_b1 , \963_b1 );
not ( \967_b1 , w_2850 );
not ( \967_b0 , w_2851 );
and ( w_2850 , w_2851 , \963_b0 );
or ( \968_b1 , \967_b1 , \964_b1 );
not ( \964_b1 , w_2852 );
and ( \968_b0 , \967_b0 , w_2853 );
and ( w_2852 , w_2853 , \964_b0 );
or ( \969_b1 , \966_b1 , w_2855 );
not ( w_2855 , w_2856 );
and ( \969_b0 , \966_b0 , w_2857 );
and ( w_2856 ,  , w_2857 );
buf ( w_2855 , \968_b1 );
not ( w_2855 , w_2858 );
not (  , w_2859 );
and ( w_2858 , w_2859 , \968_b0 );
buf ( \970_b1 , \398_b1 );
buf ( \970_b0 , \398_b0 );
buf ( \971_b1 , \970_b1 );
not ( \971_b1 , w_2860 );
not ( \971_b0 , w_2861 );
and ( w_2860 , w_2861 , \970_b0 );
buf ( \972_b1 , \571_b1 );
not ( \972_b1 , w_2862 );
not ( \972_b0 , w_2863 );
and ( w_2862 , w_2863 , \571_b0 );
buf ( \973_b1 , \972_b1 );
not ( \973_b1 , w_2864 );
not ( \973_b0 , w_2865 );
and ( w_2864 , w_2865 , \972_b0 );
buf ( \974_b1 , \918_b1 );
not ( \974_b1 , w_2866 );
not ( \974_b0 , w_2867 );
and ( w_2866 , w_2867 , \918_b0 );
or ( \975_b1 , \973_b1 , w_2868 );
or ( \975_b0 , \973_b0 , \974_b0 );
not ( \974_b0 , w_2869 );
and ( w_2869 , w_2868 , \974_b1 );
buf ( \976_b1 , \927_b1 );
not ( \976_b1 , w_2870 );
not ( \976_b0 , w_2871 );
and ( w_2870 , w_2871 , \927_b0 );
or ( \977_b1 , \975_b1 , w_2873 );
not ( w_2873 , w_2874 );
and ( \977_b0 , \975_b0 , w_2875 );
and ( w_2874 ,  , w_2875 );
buf ( w_2873 , \976_b1 );
not ( w_2873 , w_2876 );
not (  , w_2877 );
and ( w_2876 , w_2877 , \976_b0 );
buf ( \978_b1 , \977_b1 );
not ( \978_b1 , w_2878 );
not ( \978_b0 , w_2879 );
and ( w_2878 , w_2879 , \977_b0 );
or ( \979_b1 , \971_b1 , w_2880 );
or ( \979_b0 , \971_b0 , \978_b0 );
not ( \978_b0 , w_2881 );
and ( w_2881 , w_2880 , \978_b1 );
buf ( \980_b1 , \930_b1 );
buf ( \980_b0 , \930_b0 );
or ( \981_b1 , \979_b1 , w_2883 );
not ( w_2883 , w_2884 );
and ( \981_b0 , \979_b0 , w_2885 );
and ( w_2884 ,  , w_2885 );
buf ( w_2883 , \980_b1 );
not ( w_2883 , w_2886 );
not (  , w_2887 );
and ( w_2886 , w_2887 , \980_b0 );
or ( \982_b1 , \981_b1 , \276_b1 );
not ( \276_b1 , w_2888 );
and ( \982_b0 , \981_b0 , w_2889 );
and ( w_2888 , w_2889 , \276_b0 );
buf ( \983_b1 , \981_b1 );
not ( \983_b1 , w_2890 );
not ( \983_b0 , w_2891 );
and ( w_2890 , w_2891 , \981_b0 );
or ( \984_b1 , \983_b1 , \282_b1 );
not ( \282_b1 , w_2892 );
and ( \984_b0 , \983_b0 , w_2893 );
and ( w_2892 , w_2893 , \282_b0 );
or ( \985_b1 , \982_b1 , w_2895 );
not ( w_2895 , w_2896 );
and ( \985_b0 , \982_b0 , w_2897 );
and ( w_2896 ,  , w_2897 );
buf ( w_2895 , \984_b1 );
not ( w_2895 , w_2898 );
not (  , w_2899 );
and ( w_2898 , w_2899 , \984_b0 );
buf ( \986_b1 , \557_b1 );
buf ( \986_b0 , \557_b0 );
buf ( \987_b1 , \986_b1 );
not ( \987_b1 , w_2900 );
not ( \987_b0 , w_2901 );
and ( w_2900 , w_2901 , \986_b0 );
buf ( \988_b1 , \918_b1 );
not ( \988_b1 , w_2902 );
not ( \988_b0 , w_2903 );
and ( w_2902 , w_2903 , \918_b0 );
or ( \989_b1 , \987_b1 , w_2904 );
or ( \989_b0 , \987_b0 , \988_b0 );
not ( \988_b0 , w_2905 );
and ( w_2905 , w_2904 , \988_b1 );
buf ( \990_b1 , \922_b1 );
not ( \990_b1 , w_2906 );
not ( \990_b0 , w_2907 );
and ( w_2906 , w_2907 , \922_b0 );
or ( \991_b1 , \989_b1 , w_2909 );
not ( w_2909 , w_2910 );
and ( \991_b0 , \989_b0 , w_2911 );
and ( w_2910 ,  , w_2911 );
buf ( w_2909 , \990_b1 );
not ( w_2909 , w_2912 );
not (  , w_2913 );
and ( w_2912 , w_2913 , \990_b0 );
or ( \992_b1 , \570_b1 , w_2915 );
not ( w_2915 , w_2916 );
and ( \992_b0 , \570_b0 , w_2917 );
and ( w_2916 ,  , w_2917 );
buf ( w_2915 , \926_b1 );
not ( w_2915 , w_2918 );
not (  , w_2919 );
and ( w_2918 , w_2919 , \926_b0 );
buf ( \993_b1 , \992_b1 );
not ( \993_b1 , w_2920 );
not ( \993_b0 , w_2921 );
and ( w_2920 , w_2921 , \992_b0 );
or ( \994_b1 , \991_b1 , \993_b1 );
not ( \993_b1 , w_2922 );
and ( \994_b0 , \991_b0 , w_2923 );
and ( w_2922 , w_2923 , \993_b0 );
buf ( \995_b1 , \991_b1 );
not ( \995_b1 , w_2924 );
not ( \995_b0 , w_2925 );
and ( w_2924 , w_2925 , \991_b0 );
or ( \996_b1 , \995_b1 , \992_b1 );
not ( \992_b1 , w_2926 );
and ( \996_b0 , \995_b0 , w_2927 );
and ( w_2926 , w_2927 , \992_b0 );
or ( \997_b1 , \994_b1 , w_2929 );
not ( w_2929 , w_2930 );
and ( \997_b0 , \994_b0 , w_2931 );
and ( w_2930 ,  , w_2931 );
buf ( w_2929 , \996_b1 );
not ( w_2929 , w_2932 );
not (  , w_2933 );
and ( w_2932 , w_2933 , \996_b0 );
or ( \998_b1 , \868_b1 , w_2935 );
not ( w_2935 , w_2936 );
and ( \998_b0 , \868_b0 , w_2937 );
and ( w_2936 ,  , w_2937 );
buf ( w_2935 , \893_b1 );
not ( w_2935 , w_2938 );
not (  , w_2939 );
and ( w_2938 , w_2939 , \893_b0 );
buf ( \999_b1 , \998_b1 );
not ( \999_b1 , w_2940 );
not ( \999_b0 , w_2941 );
and ( w_2940 , w_2941 , \998_b0 );
buf ( \1000_b1 , \890_b1 );
buf ( \1000_b0 , \890_b0 );
or ( \1001_b1 , \999_b1 , \1000_b1 );
not ( \1000_b1 , w_2942 );
and ( \1001_b0 , \999_b0 , w_2943 );
and ( w_2942 , w_2943 , \1000_b0 );
buf ( \1002_b1 , \914_b1 );
buf ( \1002_b0 , \914_b0 );
or ( \1003_b1 , \1001_b1 , w_2945 );
not ( w_2945 , w_2946 );
and ( \1003_b0 , \1001_b0 , w_2947 );
and ( w_2946 ,  , w_2947 );
buf ( w_2945 , \1002_b1 );
not ( w_2945 , w_2948 );
not (  , w_2949 );
and ( w_2948 , w_2949 , \1002_b0 );
buf ( \1004_b1 , \916_b1 );
not ( \1004_b1 , w_2950 );
not ( \1004_b0 , w_2951 );
and ( w_2950 , w_2951 , \916_b0 );
or ( \1005_b1 , \1004_b1 , w_2953 );
not ( w_2953 , w_2954 );
and ( \1005_b0 , \1004_b0 , w_2955 );
and ( w_2954 ,  , w_2955 );
buf ( w_2953 , \913_b1 );
not ( w_2953 , w_2956 );
not (  , w_2957 );
and ( w_2956 , w_2957 , \913_b0 );
or ( \1006_b1 , \1003_b1 , \1005_b1 );
not ( \1005_b1 , w_2958 );
and ( \1006_b0 , \1003_b0 , w_2959 );
and ( w_2958 , w_2959 , \1005_b0 );
buf ( \1007_b1 , \1003_b1 );
not ( \1007_b1 , w_2960 );
not ( \1007_b0 , w_2961 );
and ( w_2960 , w_2961 , \1003_b0 );
buf ( \1008_b1 , \1005_b1 );
not ( \1008_b1 , w_2962 );
not ( \1008_b0 , w_2963 );
and ( w_2962 , w_2963 , \1005_b0 );
or ( \1009_b1 , \1007_b1 , \1008_b1 );
not ( \1008_b1 , w_2964 );
and ( \1009_b0 , \1007_b0 , w_2965 );
and ( w_2964 , w_2965 , \1008_b0 );
or ( \1010_b1 , \1006_b1 , w_2967 );
not ( w_2967 , w_2968 );
and ( \1010_b0 , \1006_b0 , w_2969 );
and ( w_2968 ,  , w_2969 );
buf ( w_2967 , \1009_b1 );
not ( w_2967 , w_2970 );
not (  , w_2971 );
and ( w_2970 , w_2971 , \1009_b0 );
buf ( \1011_b1 , \1002_b1 );
not ( \1011_b1 , w_2972 );
not ( \1011_b0 , w_2973 );
and ( w_2972 , w_2973 , \1002_b0 );
or ( \1012_b1 , \1011_b1 , w_2975 );
not ( w_2975 , w_2976 );
and ( \1012_b0 , \1011_b0 , w_2977 );
and ( w_2976 ,  , w_2977 );
buf ( w_2975 , \1000_b1 );
not ( w_2975 , w_2978 );
not (  , w_2979 );
and ( w_2978 , w_2979 , \1000_b0 );
or ( \1013_b1 , \998_b1 , \1012_b1 );
not ( \1012_b1 , w_2980 );
and ( \1013_b0 , \998_b0 , w_2981 );
and ( w_2980 , w_2981 , \1012_b0 );
buf ( \1014_b1 , \998_b1 );
not ( \1014_b1 , w_2982 );
not ( \1014_b0 , w_2983 );
and ( w_2982 , w_2983 , \998_b0 );
buf ( \1015_b1 , \1012_b1 );
not ( \1015_b1 , w_2984 );
not ( \1015_b0 , w_2985 );
and ( w_2984 , w_2985 , \1012_b0 );
or ( \1016_b1 , \1014_b1 , \1015_b1 );
not ( \1015_b1 , w_2986 );
and ( \1016_b0 , \1014_b0 , w_2987 );
and ( w_2986 , w_2987 , \1015_b0 );
or ( \1017_b1 , \1013_b1 , w_2989 );
not ( w_2989 , w_2990 );
and ( \1017_b0 , \1013_b0 , w_2991 );
and ( w_2990 ,  , w_2991 );
buf ( w_2989 , \1016_b1 );
not ( w_2989 , w_2992 );
not (  , w_2993 );
and ( w_2992 , w_2993 , \1016_b0 );
or ( \1018_b1 , \835_b1 , w_2995 );
not ( w_2995 , w_2996 );
and ( \1018_b0 , \835_b0 , w_2997 );
and ( w_2996 ,  , w_2997 );
buf ( w_2995 , \866_b1 );
not ( w_2995 , w_2998 );
not (  , w_2999 );
and ( w_2998 , w_2999 , \866_b0 );
or ( \1019_b1 , \893_b1 , w_3001 );
not ( w_3001 , w_3002 );
and ( \1019_b0 , \893_b0 , w_3003 );
and ( w_3002 ,  , w_3003 );
buf ( w_3001 , \865_b1 );
not ( w_3001 , w_3004 );
not (  , w_3005 );
and ( w_3004 , w_3005 , \865_b0 );
buf ( \1020_b1 , \1019_b1 );
not ( \1020_b1 , w_3006 );
not ( \1020_b0 , w_3007 );
and ( w_3006 , w_3007 , \1019_b0 );
or ( \1021_b1 , \1018_b1 , \1020_b1 );
not ( \1020_b1 , w_3008 );
and ( \1021_b0 , \1018_b0 , w_3009 );
and ( w_3008 , w_3009 , \1020_b0 );
buf ( \1022_b1 , \1018_b1 );
not ( \1022_b1 , w_3010 );
not ( \1022_b0 , w_3011 );
and ( w_3010 , w_3011 , \1018_b0 );
or ( \1023_b1 , \1022_b1 , \1019_b1 );
not ( \1019_b1 , w_3012 );
and ( \1023_b0 , \1022_b0 , w_3013 );
and ( w_3012 , w_3013 , \1019_b0 );
or ( \1024_b1 , \1021_b1 , w_3015 );
not ( w_3015 , w_3016 );
and ( \1024_b0 , \1021_b0 , w_3017 );
and ( w_3016 ,  , w_3017 );
buf ( w_3015 , \1023_b1 );
not ( w_3015 , w_3018 );
not (  , w_3019 );
and ( w_3018 , w_3019 , \1023_b0 );
or ( \1025_b1 , \834_b1 , w_3021 );
not ( w_3021 , w_3022 );
and ( \1025_b0 , \834_b0 , w_3023 );
and ( w_3022 ,  , w_3023 );
buf ( w_3021 , \866_b1 );
not ( w_3021 , w_3024 );
not (  , w_3025 );
and ( w_3024 , w_3025 , \866_b0 );
buf ( \1026_b1 , \1025_b1 );
not ( \1026_b1 , w_3026 );
not ( \1026_b0 , w_3027 );
and ( w_3026 , w_3027 , \1025_b0 );
or ( \1027_b1 , \781_b1 , \1026_b1 );
not ( \1026_b1 , w_3028 );
and ( \1027_b0 , \781_b0 , w_3029 );
and ( w_3028 , w_3029 , \1026_b0 );
buf ( \1028_b1 , \781_b1 );
not ( \1028_b1 , w_3030 );
not ( \1028_b0 , w_3031 );
and ( w_3030 , w_3031 , \781_b0 );
or ( \1029_b1 , \1028_b1 , \1025_b1 );
not ( \1025_b1 , w_3032 );
and ( \1029_b0 , \1028_b0 , w_3033 );
and ( w_3032 , w_3033 , \1025_b0 );
or ( \1030_b1 , \1027_b1 , w_3035 );
not ( w_3035 , w_3036 );
and ( \1030_b0 , \1027_b0 , w_3037 );
and ( w_3036 ,  , w_3037 );
buf ( w_3035 , \1029_b1 );
not ( w_3035 , w_3038 );
not (  , w_3039 );
and ( w_3038 , w_3039 , \1029_b0 );
or ( \1031_b1 , \970_b1 , w_3041 );
not ( w_3041 , w_3042 );
and ( \1031_b0 , \970_b0 , w_3043 );
and ( w_3042 ,  , w_3043 );
buf ( w_3041 , \980_b1 );
not ( w_3041 , w_3044 );
not (  , w_3045 );
and ( w_3044 , w_3045 , \980_b0 );
or ( \1032_b1 , \990_b1 , w_3047 );
not ( w_3047 , w_3048 );
and ( \1032_b0 , \990_b0 , w_3049 );
and ( w_3048 ,  , w_3049 );
buf ( w_3047 , \986_b1 );
not ( w_3047 , w_3050 );
not (  , w_3051 );
and ( w_3050 , w_3051 , \986_b0 );
or ( \1033_b1 , \780_b1 , w_3053 );
not ( w_3053 , w_3054 );
and ( \1033_b0 , \780_b0 , w_3055 );
and ( w_3054 ,  , w_3055 );
buf ( w_3053 , \676_b1 );
not ( w_3053 , w_3056 );
not (  , w_3057 );
and ( w_3056 , w_3057 , \676_b0 );
buf ( \1034_b1 , \1033_b1 );
not ( \1034_b1 , w_3058 );
not ( \1034_b0 , w_3059 );
and ( w_3058 , w_3059 , \1033_b0 );
buf ( \1035_b1 , \775_b1 );
buf ( \1035_b0 , \775_b0 );
buf ( \1036_b1 , \1035_b1 );
not ( \1036_b1 , w_3060 );
not ( \1036_b0 , w_3061 );
and ( w_3060 , w_3061 , \1035_b0 );
or ( \1037_b1 , \1034_b1 , w_3062 );
or ( \1037_b0 , \1034_b0 , \1036_b0 );
not ( \1036_b0 , w_3063 );
and ( w_3063 , w_3062 , \1036_b1 );
or ( \1038_b1 , \1035_b1 , w_3064 );
or ( \1038_b0 , \1035_b0 , \1033_b0 );
not ( \1033_b0 , w_3065 );
and ( w_3065 , w_3064 , \1033_b1 );
or ( \1039_b1 , \1037_b1 , w_3067 );
not ( w_3067 , w_3068 );
and ( \1039_b0 , \1037_b0 , w_3069 );
and ( w_3068 ,  , w_3069 );
buf ( w_3067 , \1038_b1 );
not ( w_3067 , w_3070 );
not (  , w_3071 );
and ( w_3070 , w_3071 , \1038_b0 );
or ( \1040_b1 , \423_b1 , w_3073 );
not ( w_3073 , w_3074 );
and ( \1040_b0 , \423_b0 , w_3075 );
and ( w_3074 ,  , w_3075 );
buf ( w_3073 , \962_b1 );
not ( w_3073 , w_3076 );
not (  , w_3077 );
and ( w_3076 , w_3077 , \962_b0 );
buf ( \1041_b1 , \769_b1 );
buf ( \1041_b0 , \769_b0 );
buf ( \1042_b1 , \1041_b1 );
not ( \1042_b1 , w_3078 );
not ( \1042_b0 , w_3079 );
and ( w_3078 , w_3079 , \1041_b0 );
or ( \1043_b1 , \774_b1 , w_3081 );
not ( w_3081 , w_3082 );
and ( \1043_b0 , \774_b0 , w_3083 );
and ( w_3082 ,  , w_3083 );
buf ( w_3081 , \695_b1 );
not ( w_3081 , w_3084 );
not (  , w_3085 );
and ( w_3084 , w_3085 , \695_b0 );
buf ( \1044_b1 , \1043_b1 );
not ( \1044_b1 , w_3086 );
not ( \1044_b0 , w_3087 );
and ( w_3086 , w_3087 , \1043_b0 );
or ( \1045_b1 , \1042_b1 , w_3088 );
or ( \1045_b0 , \1042_b0 , \1044_b0 );
not ( \1044_b0 , w_3089 );
and ( w_3089 , w_3088 , \1044_b1 );
or ( \1046_b1 , \1041_b1 , w_3090 );
or ( \1046_b0 , \1041_b0 , \1043_b0 );
not ( \1043_b0 , w_3091 );
and ( w_3091 , w_3090 , \1043_b1 );
or ( \1047_b1 , \1045_b1 , w_3093 );
not ( w_3093 , w_3094 );
and ( \1047_b0 , \1045_b0 , w_3095 );
and ( w_3094 ,  , w_3095 );
buf ( w_3093 , \1046_b1 );
not ( w_3093 , w_3096 );
not (  , w_3097 );
and ( w_3096 , w_3097 , \1046_b0 );
or ( \1048_b1 , \768_b1 , \714_b1 );
not ( \714_b1 , w_3098 );
and ( \1048_b0 , \768_b0 , w_3099 );
and ( w_3098 , w_3099 , \714_b0 );
or ( \1049_b1 , \1048_b1 , \765_b1 );
not ( \765_b1 , w_3100 );
and ( \1049_b0 , \1048_b0 , w_3101 );
and ( w_3100 , w_3101 , \765_b0 );
buf ( \1050_b1 , \1048_b1 );
not ( \1050_b1 , w_3102 );
not ( \1050_b0 , w_3103 );
and ( w_3102 , w_3103 , \1048_b0 );
buf ( \1051_b1 , \765_b1 );
not ( \1051_b1 , w_3104 );
not ( \1051_b0 , w_3105 );
and ( w_3104 , w_3105 , \765_b0 );
or ( \1052_b1 , \1050_b1 , \1051_b1 );
not ( \1051_b1 , w_3106 );
and ( \1052_b0 , \1050_b0 , w_3107 );
and ( w_3106 , w_3107 , \1051_b0 );
or ( \1053_b1 , \1049_b1 , w_3109 );
not ( w_3109 , w_3110 );
and ( \1053_b0 , \1049_b0 , w_3111 );
and ( w_3110 ,  , w_3111 );
buf ( w_3109 , \1052_b1 );
not ( w_3109 , w_3112 );
not (  , w_3113 );
and ( w_3112 , w_3113 , \1052_b0 );
or ( \1054_b1 , \732_b1 , w_3115 );
not ( w_3115 , w_3116 );
and ( \1054_b0 , \732_b0 , w_3117 );
and ( w_3116 ,  , w_3117 );
buf ( w_3115 , \763_b1 );
not ( w_3115 , w_3118 );
not (  , w_3119 );
and ( w_3118 , w_3119 , \763_b0 );
buf ( \1055_b1 , \762_b1 );
not ( \1055_b1 , w_3120 );
not ( \1055_b0 , w_3121 );
and ( w_3120 , w_3121 , \762_b0 );
or ( \1056_b1 , \1054_b1 , \1055_b1 );
not ( \1055_b1 , w_3122 );
and ( \1056_b0 , \1054_b0 , w_3123 );
and ( w_3122 , w_3123 , \1055_b0 );
buf ( \1057_b1 , \1054_b1 );
not ( \1057_b1 , w_3124 );
not ( \1057_b0 , w_3125 );
and ( w_3124 , w_3125 , \1054_b0 );
or ( \1058_b1 , \1057_b1 , \762_b1 );
not ( \762_b1 , w_3126 );
and ( \1058_b0 , \1057_b0 , w_3127 );
and ( w_3126 , w_3127 , \762_b0 );
or ( \1059_b1 , \1056_b1 , w_3129 );
not ( w_3129 , w_3130 );
and ( \1059_b0 , \1056_b0 , w_3131 );
and ( w_3130 ,  , w_3131 );
buf ( w_3129 , \1058_b1 );
not ( w_3129 , w_3132 );
not (  , w_3133 );
and ( w_3132 , w_3133 , \1058_b0 );
or ( \1060_b1 , \761_b1 , w_3135 );
not ( w_3135 , w_3136 );
and ( \1060_b0 , \761_b0 , w_3137 );
and ( w_3136 ,  , w_3137 );
buf ( w_3135 , \747_b1 );
not ( w_3135 , w_3138 );
not (  , w_3139 );
and ( w_3138 , w_3139 , \747_b0 );
buf ( \1061_b1 , \1060_b1 );
not ( \1061_b1 , w_3140 );
not ( \1061_b0 , w_3141 );
and ( w_3140 , w_3141 , \1060_b0 );
buf ( \1062_b1 , \757_b1 );
not ( \1062_b1 , w_3142 );
not ( \1062_b0 , w_3143 );
and ( w_3142 , w_3143 , \757_b0 );
or ( \1063_b1 , \1061_b1 , w_3144 );
or ( \1063_b0 , \1061_b0 , \1062_b0 );
not ( \1062_b0 , w_3145 );
and ( w_3145 , w_3144 , \1062_b1 );
or ( \1064_b1 , \757_b1 , w_3146 );
or ( \1064_b0 , \757_b0 , \1060_b0 );
not ( \1060_b0 , w_3147 );
and ( w_3147 , w_3146 , \1060_b1 );
or ( \1065_b1 , \1063_b1 , w_3149 );
not ( w_3149 , w_3150 );
and ( \1065_b0 , \1063_b0 , w_3151 );
and ( w_3150 ,  , w_3151 );
buf ( w_3149 , \1064_b1 );
not ( w_3149 , w_3152 );
not (  , w_3153 );
and ( w_3152 , w_3153 , \1064_b0 );
or ( \1066_b1 , \750_b1 , \752_b1 );
xor ( \1066_b0 , \750_b0 , w_3154 );
not ( w_3154 , w_3155 );
and ( w_3155 , \752_b1 , \752_b0 );
or ( \1067_b1 , \1066_b1 , \754_b1 );
xor ( \1067_b0 , \1066_b0 , w_3156 );
not ( w_3156 , w_3157 );
and ( w_3157 , \754_b1 , \754_b0 );
or ( \1068_b1 , \289_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_3158 );
and ( \1068_b0 , \289_b0 , w_3159 );
and ( w_3158 , w_3159 , \B[0]_b0 );
or ( \1069_b1 , \296_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_3160 );
and ( \1069_b0 , \296_b0 , w_3161 );
and ( w_3160 , w_3161 , \B[1]_b0 );
or ( \1070_b1 , \1068_b1 , w_3163 );
not ( w_3163 , w_3164 );
and ( \1070_b0 , \1068_b0 , w_3165 );
and ( w_3164 ,  , w_3165 );
buf ( w_3163 , \1069_b1 );
not ( w_3163 , w_3166 );
not (  , w_3167 );
and ( w_3166 , w_3167 , \1069_b0 );
or ( \1071_b1 , \752_b1 , w_3169 );
not ( w_3169 , w_3170 );
and ( \1071_b0 , \752_b0 , w_3171 );
and ( w_3170 ,  , w_3171 );
buf ( w_3169 , \1070_b1 );
not ( w_3169 , w_3172 );
not (  , w_3173 );
and ( w_3172 , w_3173 , \1070_b0 );
buf ( \1072_b1 , \751_b1 );
not ( \1072_b1 , w_3174 );
not ( \1072_b0 , w_3175 );
and ( w_3174 , w_3175 , \751_b0 );
or ( \1073_b1 , \959_b1 , w_3176 );
xor ( \1073_b0 , \959_b0 , w_3178 );
not ( w_3178 , w_3179 );
and ( w_3179 , w_3176 , w_3177 );
buf ( w_3176 , \1040_b1 );
not ( w_3176 , w_3180 );
not ( w_3177 , w_3181 );
and ( w_3180 , w_3181 , \1040_b0 );
or ( \1074_b1 , \977_b1 , w_3182 );
xor ( \1074_b0 , \977_b0 , w_3184 );
not ( w_3184 , w_3185 );
and ( w_3185 , w_3182 , w_3183 );
buf ( w_3182 , \1031_b1 );
not ( w_3182 , w_3186 );
not ( w_3183 , w_3187 );
and ( w_3186 , w_3187 , \1031_b0 );
or ( \1075_b1 , \1032_b1 , w_3188 );
xor ( \1075_b0 , \1032_b0 , w_3190 );
not ( w_3190 , w_3191 );
and ( w_3191 , w_3188 , w_3189 );
buf ( w_3188 , \918_b1 );
not ( w_3188 , w_3192 );
not ( w_3189 , w_3193 );
and ( w_3192 , w_3193 , \918_b0 );
or ( \83_b1 , \82_b1 , w_3198 );
or ( \83_b0 , \82_b0 , w_3195 );
not ( w_3195 , w_3199 );
and ( w_3199 , w_3198 , w_3194 );
or ( w_3194 , \I[0]_b1 , w_3200 );
or ( w_3195 , \I[0]_b0 , w_3197 );
not ( w_3197 , w_3201 );
and ( w_3201 , w_3200 , w_3196 );
buf ( w_3196 , \I[1]_b1 );
not ( w_3196 , w_3202 );
not ( w_3197 , w_3203 );
and ( w_3202 , w_3203 , \I[1]_b0 );
or ( \228_b1 , \227_b1 , w_3208 );
or ( \228_b0 , \227_b0 , w_3205 );
not ( w_3205 , w_3209 );
and ( w_3209 , w_3208 , w_3204 );
or ( w_3204 , \I[0]_b1 , w_3210 );
or ( w_3205 , \I[0]_b0 , w_3207 );
not ( w_3207 , w_3211 );
and ( w_3211 , w_3210 , w_3206 );
buf ( w_3206 , \I[1]_b1 );
not ( w_3206 , w_3212 );
not ( w_3207 , w_3213 );
and ( w_3212 , w_3213 , \I[1]_b0 );
or ( \278_b1 , \I[7]_b1 , w_3226 );
or ( \278_b0 , \I[7]_b0 , w_3215 );
not ( w_3215 , w_3227 );
and ( w_3227 , w_3226 , w_3214 );
or ( w_3214 , \I[6]_b1 , w_3228 );
or ( w_3215 , \I[6]_b0 , w_3217 );
not ( w_3217 , w_3229 );
and ( w_3229 , w_3228 , w_3216 );
or ( w_3216 , \I[5]_b1 , w_3230 );
or ( w_3217 , \I[5]_b0 , w_3219 );
not ( w_3219 , w_3231 );
and ( w_3231 , w_3230 , w_3218 );
or ( w_3218 , \I[4]_b1 , w_3232 );
or ( w_3219 , \I[4]_b0 , w_3221 );
not ( w_3221 , w_3233 );
and ( w_3233 , w_3232 , w_3220 );
or ( w_3220 , \I[3]_b1 , w_3234 );
or ( w_3221 , \I[3]_b0 , w_3223 );
not ( w_3223 , w_3235 );
and ( w_3235 , w_3234 , w_3222 );
or ( w_3222 , \I[2]_b1 , w_3236 );
or ( w_3223 , \I[2]_b0 , w_3225 );
not ( w_3225 , w_3237 );
and ( w_3237 , w_3236 , w_3224 );
or ( w_3224 , \I[1]_b1 , w_3238 );
or ( w_3225 , \I[1]_b0 , \I[0]_b0 );
not ( \I[0]_b0 , w_3239 );
and ( w_3239 , w_3238 , \I[0]_b1 );
or ( \279_b1 , \B[9]_b1 , w_3240 );
not ( w_3240 , w_3256 );
and ( \279_b0 , \B[9]_b0 , w_3257 );
and ( w_3256 , w_3257 , w_3241 );
or ( w_3240 , \B[8]_b1 , w_3242 );
not ( w_3242 , w_3258 );
and ( w_3241 , \B[8]_b0 , w_3259 );
and ( w_3258 , w_3259 , w_3243 );
or ( w_3242 , \B[7]_b1 , w_3244 );
not ( w_3244 , w_3260 );
and ( w_3243 , \B[7]_b0 , w_3261 );
and ( w_3260 , w_3261 , w_3245 );
or ( w_3244 , \B[6]_b1 , w_3246 );
not ( w_3246 , w_3262 );
and ( w_3245 , \B[6]_b0 , w_3263 );
and ( w_3262 , w_3263 , w_3247 );
or ( w_3246 , \B[5]_b1 , w_3248 );
not ( w_3248 , w_3264 );
and ( w_3247 , \B[5]_b0 , w_3265 );
and ( w_3264 , w_3265 , w_3249 );
or ( w_3248 , \B[4]_b1 , w_3250 );
not ( w_3250 , w_3266 );
and ( w_3249 , \B[4]_b0 , w_3267 );
and ( w_3266 , w_3267 , w_3251 );
or ( w_3250 , \B[3]_b1 , w_3252 );
not ( w_3252 , w_3268 );
and ( w_3251 , \B[3]_b0 , w_3269 );
and ( w_3268 , w_3269 , w_3253 );
or ( w_3252 , \B[2]_b1 , w_3254 );
not ( w_3254 , w_3270 );
and ( w_3253 , \B[2]_b0 , w_3271 );
and ( w_3270 , w_3271 , w_3255 );
or ( w_3254 , \B[1]_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_3272 );
and ( w_3255 , \B[1]_b0 , w_3273 );
and ( w_3272 , w_3273 , \B[0]_b0 );
or ( \284_b1 , \283_b1 , w_3278 );
or ( \284_b0 , \283_b0 , w_3275 );
not ( w_3275 , w_3279 );
and ( w_3279 , w_3278 , w_3274 );
or ( w_3274 , \I[0]_b1 , w_3280 );
or ( w_3275 , \I[0]_b0 , w_3277 );
not ( w_3277 , w_3281 );
and ( w_3281 , w_3280 , w_3276 );
buf ( w_3276 , \I[1]_b1 );
not ( w_3276 , w_3282 );
not ( w_3277 , w_3283 );
and ( w_3282 , w_3283 , \I[1]_b0 );
or ( \938_b1 , \928_b1 , w_3284 );
not ( w_3284 , w_3286 );
and ( \938_b0 , \928_b0 , w_3287 );
and ( w_3286 , w_3287 , w_3285 );
or ( w_3284 , \936_b1 , \937_b1 );
not ( \937_b1 , w_3288 );
and ( w_3285 , \936_b0 , w_3289 );
and ( w_3288 , w_3289 , \937_b0 );
endmodule

