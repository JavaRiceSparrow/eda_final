// ...
module top(\A[2][9]_b1 ,\A[2][9]_b0 ,\A[2][8]_b1 ,\A[2][8]_b0 ,\A[2][7]_b1 ,\A[2][7]_b0 ,\A[2][6]_b1 ,\A[2][6]_b0 ,\A[2][5]_b1 ,
		\A[2][5]_b0 ,\A[2][4]_b1 ,\A[2][4]_b0 ,\A[2][3]_b1 ,\A[2][3]_b0 ,\A[2][2]_b1 ,\A[2][2]_b0 ,\A[2][1]_b1 ,\A[2][1]_b0 ,
		\A[2][0]_b1 ,\A[2][0]_b0 ,\A[1][9]_b1 ,\A[1][9]_b0 ,\A[1][8]_b1 ,\A[1][8]_b0 ,\A[1][7]_b1 ,\A[1][7]_b0 ,\A[1][6]_b1 ,
		\A[1][6]_b0 ,\A[1][5]_b1 ,\A[1][5]_b0 ,\A[1][4]_b1 ,\A[1][4]_b0 ,\A[1][3]_b1 ,\A[1][3]_b0 ,\A[1][2]_b1 ,\A[1][2]_b0 ,
		\A[1][1]_b1 ,\A[1][1]_b0 ,\A[1][0]_b1 ,\A[1][0]_b0 ,\A[0][9]_b1 ,\A[0][9]_b0 ,\A[0][8]_b1 ,\A[0][8]_b0 ,\A[0][7]_b1 ,
		\A[0][7]_b0 ,\A[0][6]_b1 ,\A[0][6]_b0 ,\A[0][5]_b1 ,\A[0][5]_b0 ,\A[0][4]_b1 ,\A[0][4]_b0 ,\A[0][3]_b1 ,\A[0][3]_b0 ,
		\A[0][2]_b1 ,\A[0][2]_b0 ,\A[0][1]_b1 ,\A[0][1]_b0 ,\A[0][0]_b1 ,\A[0][0]_b0 ,\B[9]_b1 ,\B[9]_b0 ,\B[8]_b1 ,
		\B[8]_b0 ,\B[7]_b1 ,\B[7]_b0 ,\B[6]_b1 ,\B[6]_b0 ,\B[5]_b1 ,\B[5]_b0 ,\B[4]_b1 ,\B[4]_b0 ,
		\B[3]_b1 ,\B[3]_b0 ,\B[2]_b1 ,\B[2]_b0 ,\B[1]_b1 ,\B[1]_b0 ,\B[0]_b1 ,\B[0]_b0 ,\I[7]_b1 ,
		\I[7]_b0 ,\I[6]_b1 ,\I[6]_b0 ,\I[5]_b1 ,\I[5]_b0 ,\I[4]_b1 ,\I[4]_b0 ,\I[3]_b1 ,\I[3]_b0 ,
		\I[2]_b1 ,\I[2]_b0 ,\I[1]_b1 ,\I[1]_b0 ,\I[0]_b1 ,\I[0]_b0 ,\O[19]_b1 ,\O[19]_b0 ,\O[18]_b1 ,
		\O[18]_b0 ,\O[17]_b1 ,\O[17]_b0 ,\O[16]_b1 ,\O[16]_b0 ,\O[15]_b1 ,\O[15]_b0 ,\O[14]_b1 ,\O[14]_b0 ,
		\O[13]_b1 ,\O[13]_b0 ,\O[12]_b1 ,\O[12]_b0 ,\O[11]_b1 ,\O[11]_b0 ,\O[10]_b1 ,\O[10]_b0 ,\O[9]_b1 ,
		\O[9]_b0 ,\O[8]_b1 ,\O[8]_b0 ,\O[7]_b1 ,\O[7]_b0 ,\O[6]_b1 ,\O[6]_b0 ,\O[5]_b1 ,\O[5]_b0 ,
		\O[4]_b1 ,\O[4]_b0 ,\O[3]_b1 ,\O[3]_b0 ,\O[2]_b1 ,\O[2]_b0 ,\O[1]_b1 ,\O[1]_b0 ,\O[0]_b1 ,
		\O[0]_b0 );
input \A[2][9]_b1 ,\A[2][9]_b0 ,\A[2][8]_b1 ,\A[2][8]_b0 ,\A[2][7]_b1 ,\A[2][7]_b0 ,\A[2][6]_b1 ,\A[2][6]_b0 ,\A[2][5]_b1 ,
		\A[2][5]_b0 ,\A[2][4]_b1 ,\A[2][4]_b0 ,\A[2][3]_b1 ,\A[2][3]_b0 ,\A[2][2]_b1 ,\A[2][2]_b0 ,\A[2][1]_b1 ,\A[2][1]_b0 ,
		\A[2][0]_b1 ,\A[2][0]_b0 ,\A[1][9]_b1 ,\A[1][9]_b0 ,\A[1][8]_b1 ,\A[1][8]_b0 ,\A[1][7]_b1 ,\A[1][7]_b0 ,\A[1][6]_b1 ,
		\A[1][6]_b0 ,\A[1][5]_b1 ,\A[1][5]_b0 ,\A[1][4]_b1 ,\A[1][4]_b0 ,\A[1][3]_b1 ,\A[1][3]_b0 ,\A[1][2]_b1 ,\A[1][2]_b0 ,
		\A[1][1]_b1 ,\A[1][1]_b0 ,\A[1][0]_b1 ,\A[1][0]_b0 ,\A[0][9]_b1 ,\A[0][9]_b0 ,\A[0][8]_b1 ,\A[0][8]_b0 ,\A[0][7]_b1 ,
		\A[0][7]_b0 ,\A[0][6]_b1 ,\A[0][6]_b0 ,\A[0][5]_b1 ,\A[0][5]_b0 ,\A[0][4]_b1 ,\A[0][4]_b0 ,\A[0][3]_b1 ,\A[0][3]_b0 ,
		\A[0][2]_b1 ,\A[0][2]_b0 ,\A[0][1]_b1 ,\A[0][1]_b0 ,\A[0][0]_b1 ,\A[0][0]_b0 ,\B[9]_b1 ,\B[9]_b0 ,\B[8]_b1 ,
		\B[8]_b0 ,\B[7]_b1 ,\B[7]_b0 ,\B[6]_b1 ,\B[6]_b0 ,\B[5]_b1 ,\B[5]_b0 ,\B[4]_b1 ,\B[4]_b0 ,
		\B[3]_b1 ,\B[3]_b0 ,\B[2]_b1 ,\B[2]_b0 ,\B[1]_b1 ,\B[1]_b0 ,\B[0]_b1 ,\B[0]_b0 ,\I[7]_b1 ,
		\I[7]_b0 ,\I[6]_b1 ,\I[6]_b0 ,\I[5]_b1 ,\I[5]_b0 ,\I[4]_b1 ,\I[4]_b0 ,\I[3]_b1 ,\I[3]_b0 ,
		\I[2]_b1 ,\I[2]_b0 ,\I[1]_b1 ,\I[1]_b0 ,\I[0]_b1 ,\I[0]_b0 ;
output \O[19]_b1 ,\O[19]_b0 ,\O[18]_b1 ,\O[18]_b0 ,\O[17]_b1 ,\O[17]_b0 ,\O[16]_b1 ,\O[16]_b0 ,\O[15]_b1 ,
		\O[15]_b0 ,\O[14]_b1 ,\O[14]_b0 ,\O[13]_b1 ,\O[13]_b0 ,\O[12]_b1 ,\O[12]_b0 ,\O[11]_b1 ,\O[11]_b0 ,
		\O[10]_b1 ,\O[10]_b0 ,\O[9]_b1 ,\O[9]_b0 ,\O[8]_b1 ,\O[8]_b0 ,\O[7]_b1 ,\O[7]_b0 ,\O[6]_b1 ,
		\O[6]_b0 ,\O[5]_b1 ,\O[5]_b0 ,\O[4]_b1 ,\O[4]_b0 ,\O[3]_b1 ,\O[3]_b0 ,\O[2]_b1 ,\O[2]_b0 ,
		\O[1]_b1 ,\O[1]_b0 ,\O[0]_b1 ,\O[0]_b0 ;

wire \69_ZERO_b1 , \69_ZERO_b0 , \70_ZERO_b1 , \70_ZERO_b0 , \71_ZERO_b1 , \71_ZERO_b0 , \72_ZERO_b1 , \72_ZERO_b0 , \73_ZERO_b1 , \73_ZERO_b0 , 
		\74_ZERO_b1 , \74_ZERO_b0 , \75_ZERO_b1 , \75_ZERO_b0 , \76_b1 , \76_b0 , \77_b1 , \77_b0 , \78_b1 , \78_b0 , 
		\79_b1 , \79_b0 , \80_b1 , \80_b0 , \81_b1 , \81_b0 , \82_b1 , \82_b0 , \83_b1 , \83_b0 , 
		\84_b1 , \84_b0 , \85_b1 , \85_b0 , \86_ONE_b1 , \86_ONE_b0 , \87_ONE_b1 , \87_ONE_b0 , \88_b1 , \88_b0 , 
		\89_b1 , \89_b0 , \90_b1 , \90_b0 , \91_b1 , \91_b0 , \92_b1 , \92_b0 , \93_b1 , \93_b0 , 
		\94_b1 , \94_b0 , \95_b1 , \95_b0 , \96_b1 , \96_b0 , \97_b1 , \97_b0 , \98_b1 , \98_b0 , 
		\99_b1 , \99_b0 , \100_b1 , \100_b0 , \101_b1 , \101_b0 , \102_b1 , \102_b0 , \103_b1 , \103_b0 , 
		\104_b1 , \104_b0 , \105_b1 , \105_b0 , \106_b1 , \106_b0 , \107_b1 , \107_b0 , \108_b1 , \108_b0 , 
		\109_A[9]_b1 , \109_A[9]_b0 , \110_b1 , \110_b0 , \111_b1 , \111_b0 , \112_b1 , \112_b0 , \113_b1 , \113_b0 , 
		\114_b1 , \114_b0 , \115_A[8]_b1 , \115_A[8]_b0 , \116_b1 , \116_b0 , \117_b1 , \117_b0 , \118_b1 , \118_b0 , 
		\119_b1 , \119_b0 , \120_b1 , \120_b0 , \121_A[7]_b1 , \121_A[7]_b0 , \122_b1 , \122_b0 , \123_b1 , \123_b0 , 
		\124_b1 , \124_b0 , \125_b1 , \125_b0 , \126_b1 , \126_b0 , \127_A[6]_b1 , \127_A[6]_b0 , \128_b1 , \128_b0 , 
		\129_b1 , \129_b0 , \130_b1 , \130_b0 , \131_b1 , \131_b0 , \132_b1 , \132_b0 , \133_A[5]_b1 , \133_A[5]_b0 , 
		\134_b1 , \134_b0 , \135_b1 , \135_b0 , \136_b1 , \136_b0 , \137_b1 , \137_b0 , \138_b1 , \138_b0 , 
		\139_A[4]_b1 , \139_A[4]_b0 , \140_b1 , \140_b0 , \141_b1 , \141_b0 , \142_b1 , \142_b0 , \143_b1 , \143_b0 , 
		\144_b1 , \144_b0 , \145_A[3]_b1 , \145_A[3]_b0 , \146_b1 , \146_b0 , \147_b1 , \147_b0 , \148_b1 , \148_b0 , 
		\149_b1 , \149_b0 , \150_b1 , \150_b0 , \151_A[2]_b1 , \151_A[2]_b0 , \152_b1 , \152_b0 , \153_b1 , \153_b0 , 
		\154_b1 , \154_b0 , \155_b1 , \155_b0 , \156_b1 , \156_b0 , \157_A[1]_b1 , \157_A[1]_b0 , \158_b1 , \158_b0 , 
		\159_b1 , \159_b0 , \160_b1 , \160_b0 , \161_b1 , \161_b0 , \162_b1 , \162_b0 , \163_A[0]_b1 , \163_A[0]_b0 , 
		\164_B[9]_b1 , \164_B[9]_b0 , \165_B[8]_b1 , \165_B[8]_b0 , \166_B[7]_b1 , \166_B[7]_b0 , \167_B[6]_b1 , \167_B[6]_b0 , \168_B[5]_b1 , \168_B[5]_b0 , 
		\169_B[4]_b1 , \169_B[4]_b0 , \170_B[3]_b1 , \170_B[3]_b0 , \171_B[2]_b1 , \171_B[2]_b0 , \172_B[1]_b1 , \172_B[1]_b0 , \173_B[0]_b1 , \173_B[0]_b0 , 
		\174_b1 , \174_b0 , \175_b1 , \175_b0 , \176_b1 , \176_b0 , \177_b1 , \177_b0 , \178_b1 , \178_b0 , 
		\179_b1 , \179_b0 , \180_b1 , \180_b0 , \181_b1 , \181_b0 , \182_b1 , \182_b0 , \183_b1 , \183_b0 , 
		\184_b1 , \184_b0 , \185_b1 , \185_b0 , \186_b1 , \186_b0 , \187_b1 , \187_b0 , \188_b1 , \188_b0 , 
		\189_b1 , \189_b0 , \190_b1 , \190_b0 , \191_b1 , \191_b0 , \192_b1 , \192_b0 , \193_b1 , \193_b0 , 
		\194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , \197_b1 , \197_b0 , \198_b1 , \198_b0 , 
		\199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , \202_b1 , \202_b0 , \203_b1 , \203_b0 , 
		\204_b1 , \204_b0 , \205_b1 , \205_b0 , \206_b1 , \206_b0 , \207_b1 , \207_b0 , \208_b1 , \208_b0 , 
		\209_b1 , \209_b0 , \210_b1 , \210_b0 , \211_b1 , \211_b0 , \212_b1 , \212_b0 , \213_b1 , \213_b0 , 
		\214_b1 , \214_b0 , \215_b1 , \215_b0 , \216_b1 , \216_b0 , \217_b1 , \217_b0 , \218_b1 , \218_b0 , 
		\219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , \222_b1 , \222_b0 , \223_b1 , \223_b0 , 
		\224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , \227_b1 , \227_b0 , \228_b1 , \228_b0 , 
		\229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , \232_b1 , \232_b0 , \233_b1 , \233_b0 , 
		\234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , \237_b1 , \237_b0 , \238_b1 , \238_b0 , 
		\239_b1 , \239_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , \242_b1 , \242_b0 , \243_b1 , \243_b0 , 
		\244_b1 , \244_b0 , \245_b1 , \245_b0 , \246_b1 , \246_b0 , \247_b1 , \247_b0 , \248_b1 , \248_b0 , 
		\249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , \252_b1 , \252_b0 , \253_b1 , \253_b0 , 
		\254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , \257_b1 , \257_b0 , \258_b1 , \258_b0 , 
		\259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , \262_b1 , \262_b0 , \263_b1 , \263_b0 , 
		\264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , \267_b1 , \267_b0 , \268_b1 , \268_b0 , 
		\269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , \272_b1 , \272_b0 , \273_b1 , \273_b0 , 
		\274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_b1 , \276_b0 , \277_b1 , \277_b0 , \278_b1 , \278_b0 , 
		\279_b1 , \279_b0 , \280_b1 , \280_b0 , \281_b1 , \281_b0 , \282_b1 , \282_b0 , \283_b1 , \283_b0 , 
		\284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , \287_b1 , \287_b0 , \288_b1 , \288_b0 , 
		\289_b1 , \289_b0 , \290_b1 , \290_b0 , \291_b1 , \291_b0 , \292_b1 , \292_b0 , \293_b1 , \293_b0 , 
		\294_b1 , \294_b0 , \295_b1 , \295_b0 , \296_b1 , \296_b0 , \297_b1 , \297_b0 , \298_b1 , \298_b0 , 
		\299_b1 , \299_b0 , \300_b1 , \300_b0 , \301_b1 , \301_b0 , \302_b1 , \302_b0 , \303_b1 , \303_b0 , 
		\304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , \307_b1 , \307_b0 , \308_b1 , \308_b0 , 
		\309_b1 , \309_b0 , \310_b1 , \310_b0 , \311_b1 , \311_b0 , \312_b1 , \312_b0 , \313_b1 , \313_b0 , 
		\314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_b1 , \316_b0 , \317_b1 , \317_b0 , \318_b1 , \318_b0 , 
		\319_b1 , \319_b0 , \320_b1 , \320_b0 , \321_b1 , \321_b0 , \322_b1 , \322_b0 , \323_b1 , \323_b0 , 
		\324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , \327_b1 , \327_b0 , \328_b1 , \328_b0 , 
		\329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_b1 , \331_b0 , \332_b1 , \332_b0 , \333_b1 , \333_b0 , 
		\334_b1 , \334_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , \337_b1 , \337_b0 , \338_b1 , \338_b0 , 
		\339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_b1 , \341_b0 , \342_b1 , \342_b0 , \343_b1 , \343_b0 , 
		\344_b1 , \344_b0 , \345_b1 , \345_b0 , \346_b1 , \346_b0 , \347_b1 , \347_b0 , \348_b1 , \348_b0 , 
		\349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , \352_b1 , \352_b0 , \353_b1 , \353_b0 , 
		\354_b1 , \354_b0 , \355_b1 , \355_b0 , \356_b1 , \356_b0 , \357_b1 , \357_b0 , \358_b1 , \358_b0 , 
		\359_b1 , \359_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , \362_b1 , \362_b0 , \363_b1 , \363_b0 , 
		\364_b1 , \364_b0 , \365_b1 , \365_b0 , \366_b1 , \366_b0 , \367_b1 , \367_b0 , \368_b1 , \368_b0 , 
		\369_b1 , \369_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , \372_b1 , \372_b0 , \373_b1 , \373_b0 , 
		\374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , \377_b1 , \377_b0 , \378_b1 , \378_b0 , 
		\379_b1 , \379_b0 , \380_b1 , \380_b0 , \381_b1 , \381_b0 , \382_b1 , \382_b0 , \383_b1 , \383_b0 , 
		\384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , \387_b1 , \387_b0 , \388_b1 , \388_b0 , 
		\389_b1 , \389_b0 , \390_b1 , \390_b0 , \391_b1 , \391_b0 , \392_b1 , \392_b0 , \393_b1 , \393_b0 , 
		\394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , \397_b1 , \397_b0 , \398_b1 , \398_b0 , 
		\399_b1 , \399_b0 , \400_b1 , \400_b0 , \401_b1 , \401_b0 , \402_b1 , \402_b0 , \403_b1 , \403_b0 , 
		\404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , \407_b1 , \407_b0 , \408_b1 , \408_b0 , 
		\409_b1 , \409_b0 , \410_b1 , \410_b0 , \411_b1 , \411_b0 , \412_b1 , \412_b0 , \413_b1 , \413_b0 , 
		\414_b1 , \414_b0 , \415_b1 , \415_b0 , \416_b1 , \416_b0 , \417_b1 , \417_b0 , \418_b1 , \418_b0 , 
		\419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , \422_b1 , \422_b0 , \423_b1 , \423_b0 , 
		\424_b1 , \424_b0 , \425_b1 , \425_b0 , \426_b1 , \426_b0 , \427_b1 , \427_b0 , \428_b1 , \428_b0 , 
		\429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , \432_b1 , \432_b0 , \433_b1 , \433_b0 , 
		\434_b1 , \434_b0 , \435_b1 , \435_b0 , \436_b1 , \436_b0 , \437_b1 , \437_b0 , \438_b1 , \438_b0 , 
		\439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , \442_b1 , \442_b0 , \443_b1 , \443_b0 , 
		\444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_b1 , \446_b0 , \447_b1 , \447_b0 , \448_b1 , \448_b0 , 
		\449_b1 , \449_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , \452_b1 , \452_b0 , \453_b1 , \453_b0 , 
		\454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_b1 , \456_b0 , \457_b1 , \457_b0 , \458_b1 , \458_b0 , 
		\459_b1 , \459_b0 , \460_b1 , \460_b0 , \461_b1 , \461_b0 , \462_b1 , \462_b0 , \463_b1 , \463_b0 , 
		\464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , \467_b1 , \467_b0 , \468_b1 , \468_b0 , 
		\469_b1 , \469_b0 , \470_b1 , \470_b0 , \471_b1 , \471_b0 , \472_b1 , \472_b0 , \473_b1 , \473_b0 , 
		\474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , \477_b1 , \477_b0 , \478_b1 , \478_b0 , 
		\479_b1 , \479_b0 , \480_b1 , \480_b0 , \481_b1 , \481_b0 , \482_b1 , \482_b0 , \483_b1 , \483_b0 , 
		\484_b1 , \484_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , \487_b1 , \487_b0 , \488_b1 , \488_b0 , 
		\489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , \492_b1 , \492_b0 , \493_b1 , \493_b0 , 
		\494_b1 , \494_b0 , \495_b1 , \495_b0 , \496_b1 , \496_b0 , \497_b1 , \497_b0 , \498_b1 , \498_b0 , 
		\499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , \502_b1 , \502_b0 , \503_b1 , \503_b0 , 
		\504_b1 , \504_b0 , \505_b1 , \505_b0 , \506_b1 , \506_b0 , \507_b1 , \507_b0 , \508_b1 , \508_b0 , 
		\509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , \512_b1 , \512_b0 , \513_b1 , \513_b0 , 
		\514_b1 , \514_b0 , \515_b1 , \515_b0 , \516_b1 , \516_b0 , \517_b1 , \517_b0 , \518_b1 , \518_b0 , 
		\519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , \522_b1 , \522_b0 , \523_b1 , \523_b0 , 
		\524_b1 , \524_b0 , \525_b1 , \525_b0 , \526_b1 , \526_b0 , \527_b1 , \527_b0 , \528_b1 , \528_b0 , 
		\529_b1 , \529_b0 , \530_b1 , \530_b0 , \531_b1 , \531_b0 , \532_b1 , \532_b0 , \533_b1 , \533_b0 , 
		\534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_b1 , \536_b0 , \537_b1 , \537_b0 , \538_b1 , \538_b0 , 
		\539_b1 , \539_b0 , \540_b1 , \540_b0 , \541_b1 , \541_b0 , \542_b1 , \542_b0 , \543_b1 , \543_b0 , 
		\544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , \547_b1 , \547_b0 , \548_b1 , \548_b0 , 
		\549_b1 , \549_b0 , \550_b1 , \550_b0 , \551_b1 , \551_b0 , \552_b1 , \552_b0 , \553_b1 , \553_b0 , 
		\554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , \557_b1 , \557_b0 , \558_b1 , \558_b0 , 
		\559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_b1 , \561_b0 , \562_b1 , \562_b0 , \563_b1 , \563_b0 , 
		\564_b1 , \564_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , \567_b1 , \567_b0 , \568_b1 , \568_b0 , 
		\569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_b1 , \571_b0 , \572_b1 , \572_b0 , \573_b1 , \573_b0 , 
		\574_b1 , \574_b0 , \575_b1 , \575_b0 , \576_b1 , \576_b0 , \577_b1 , \577_b0 , \578_b1 , \578_b0 , 
		\579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , \582_b1 , \582_b0 , \583_b1 , \583_b0 , 
		\584_b1 , \584_b0 , \585_b1 , \585_b0 , \586_b1 , \586_b0 , \587_b1 , \587_b0 , \588_b1 , \588_b0 , 
		\589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , \592_b1 , \592_b0 , \593_b1 , \593_b0 , 
		\594_b1 , \594_b0 , \595_b1 , \595_b0 , \596_b1 , \596_b0 , \597_b1 , \597_b0 , \598_b1 , \598_b0 , 
		\599_b1 , \599_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , \602_b1 , \602_b0 , \603_b1 , \603_b0 , 
		\604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_b1 , \606_b0 , \607_b1 , \607_b0 , \608_b1 , \608_b0 , 
		\609_b1 , \609_b0 , \610_b1 , \610_b0 , \611_b1 , \611_b0 , \612_b1 , \612_b0 , \613_b1 , \613_b0 , 
		\614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , \617_b1 , \617_b0 , \618_b1 , \618_b0 , 
		\619_b1 , \619_b0 , \620_b1 , \620_b0 , \621_b1 , \621_b0 , \622_b1 , \622_b0 , \623_b1 , \623_b0 , 
		\624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , \627_b1 , \627_b0 , \628_b1 , \628_b0 , 
		\629_b1 , \629_b0 , \630_b1 , \630_b0 , \631_b1 , \631_b0 , \632_b1 , \632_b0 , \633_b1 , \633_b0 , 
		\634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , \637_b1 , \637_b0 , \638_b1 , \638_b0 , 
		\639_b1 , \639_b0 , \640_b1 , \640_b0 , \641_b1 , \641_b0 , \642_b1 , \642_b0 , \643_b1 , \643_b0 , 
		\644_b1 , \644_b0 , \645_b1 , \645_b0 , \646_b1 , \646_b0 , \647_b1 , \647_b0 , \648_b1 , \648_b0 , 
		\649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , \652_b1 , \652_b0 , \653_b1 , \653_b0 , 
		\654_b1 , \654_b0 , \655_b1 , \655_b0 , \656_b1 , \656_b0 , \657_b1 , \657_b0 , \658_b1 , \658_b0 , 
		\659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , \662_b1 , \662_b0 , \663_b1 , \663_b0 , 
		\664_b1 , \664_b0 , \665_b1 , \665_b0 , \666_b1 , \666_b0 , \667_b1 , \667_b0 , \668_b1 , \668_b0 , 
		\669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , \672_b1 , \672_b0 , \673_b1 , \673_b0 , 
		\674_b1 , \674_b0 , \675_Z[19]_b1 , \675_Z[19]_b0 , \676_b1 , \676_b0 , \677_Z[18]_b1 , \677_Z[18]_b0 , \678_b1 , \678_b0 , 
		\679_Z[17]_b1 , \679_Z[17]_b0 , \680_b1 , \680_b0 , \681_Z[16]_b1 , \681_Z[16]_b0 , \682_b1 , \682_b0 , \683_Z[15]_b1 , \683_Z[15]_b0 , 
		\684_b1 , \684_b0 , \685_Z[14]_b1 , \685_Z[14]_b0 , \686_b1 , \686_b0 , \687_Z[13]_b1 , \687_Z[13]_b0 , \688_b1 , \688_b0 , 
		\689_Z[12]_b1 , \689_Z[12]_b0 , \690_b1 , \690_b0 , \691_Z[11]_b1 , \691_Z[11]_b0 , \692_b1 , \692_b0 , \693_Z[10]_b1 , \693_Z[10]_b0 , 
		\694_b1 , \694_b0 , \695_Z[9]_b1 , \695_Z[9]_b0 , \696_b1 , \696_b0 , \697_Z[8]_b1 , \697_Z[8]_b0 , \698_b1 , \698_b0 , 
		\699_Z[7]_b1 , \699_Z[7]_b0 , \700_b1 , \700_b0 , \701_Z[6]_b1 , \701_Z[6]_b0 , \702_b1 , \702_b0 , \703_Z[5]_b1 , \703_Z[5]_b0 , 
		\704_b1 , \704_b0 , \705_Z[4]_b1 , \705_Z[4]_b0 , \706_b1 , \706_b0 , \707_Z[3]_b1 , \707_Z[3]_b0 , \708_b1 , \708_b0 , 
		\709_Z[2]_b1 , \709_Z[2]_b0 , \710_b1 , \710_b0 , \711_Z[1]_b1 , \711_Z[1]_b0 , \712_b1 , \712_b0 , \713_Z[0]_b1 , \713_Z[0]_b0 , 
		w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , w_6 , w_7 , w_8 , w_9 , 
		w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , w_16 , w_17 , w_18 , w_19 , 
		w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , w_26 , w_27 , w_28 , w_29 , 
		w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , w_36 , w_37 , w_38 , w_39 , 
		w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , w_46 , w_47 , w_48 , w_49 , 
		w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , w_56 , w_57 , w_58 , w_59 , 
		w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , w_66 , w_67 , w_68 , w_69 , 
		w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , w_76 , w_77 , w_78 , w_79 , 
		w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , w_86 , w_87 , w_88 , w_89 , 
		w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , w_96 , w_97 , w_98 , w_99 , 
		w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , w_106 , w_107 , w_108 , w_109 , 
		w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , w_116 , w_117 , w_118 , w_119 , 
		w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , w_126 , w_127 , w_128 , w_129 , 
		w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , w_136 , w_137 , w_138 , w_139 , 
		w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , w_146 , w_147 , w_148 , w_149 , 
		w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , w_156 , w_157 , w_158 , w_159 , 
		w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , w_166 , w_167 , w_168 , w_169 , 
		w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , w_176 , w_177 , w_178 , w_179 , 
		w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , w_186 , w_187 , w_188 , w_189 , 
		w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , w_196 , w_197 , w_198 , w_199 , 
		w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , w_206 , w_207 , w_208 , w_209 , 
		w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , w_216 , w_217 , w_218 , w_219 , 
		w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , w_226 , w_227 , w_228 , w_229 , 
		w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , w_236 , w_237 , w_238 , w_239 , 
		w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , w_246 , w_247 , w_248 , w_249 , 
		w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , w_256 , w_257 , w_258 , w_259 , 
		w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , w_266 , w_267 , w_268 , w_269 , 
		w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , w_276 , w_277 , w_278 , w_279 , 
		w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , w_286 , w_287 , w_288 , w_289 , 
		w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , w_296 , w_297 , w_298 , w_299 , 
		w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , w_306 , w_307 , w_308 , w_309 , 
		w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , w_316 , w_317 , w_318 , w_319 , 
		w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , w_326 , w_327 , w_328 , w_329 , 
		w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , w_336 , w_337 , w_338 , w_339 , 
		w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , w_346 , w_347 , w_348 , w_349 , 
		w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , w_356 , w_357 , w_358 , w_359 , 
		w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , w_366 , w_367 , w_368 , w_369 , 
		w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , w_376 , w_377 , w_378 , w_379 , 
		w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , w_386 , w_387 , w_388 , w_389 , 
		w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , w_396 , w_397 , w_398 , w_399 , 
		w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , w_406 , w_407 , w_408 , w_409 , 
		w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , w_416 , w_417 , w_418 , w_419 , 
		w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , w_426 , w_427 , w_428 , w_429 , 
		w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , w_436 , w_437 , w_438 , w_439 , 
		w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , w_446 , w_447 , w_448 , w_449 , 
		w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , w_456 , w_457 , w_458 , w_459 , 
		w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , w_466 , w_467 , w_468 , w_469 , 
		w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , w_476 , w_477 , w_478 , w_479 , 
		w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , w_486 , w_487 , w_488 , w_489 , 
		w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , w_496 , w_497 , w_498 , w_499 , 
		w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , w_506 , w_507 , w_508 , w_509 , 
		w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , w_516 , w_517 , w_518 , w_519 , 
		w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , w_526 , w_527 , w_528 , w_529 , 
		w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , w_536 , w_537 , w_538 , w_539 , 
		w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , w_546 , w_547 , w_548 , w_549 , 
		w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , w_556 , w_557 , w_558 , w_559 , 
		w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , w_566 , w_567 , w_568 , w_569 , 
		w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , w_576 , w_577 , w_578 , w_579 , 
		w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , w_586 , w_587 , w_588 , w_589 , 
		w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , w_596 , w_597 , w_598 , w_599 , 
		w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , w_606 , w_607 , w_608 , w_609 , 
		w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , w_616 , w_617 , w_618 , w_619 , 
		w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , w_626 , w_627 , w_628 , w_629 , 
		w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , w_636 , w_637 , w_638 , w_639 , 
		w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , w_646 , w_647 , w_648 , w_649 , 
		w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , w_656 , w_657 , w_658 , w_659 , 
		w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , w_666 , w_667 , w_668 , w_669 , 
		w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , w_676 , w_677 , w_678 , w_679 , 
		w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , w_686 , w_687 , w_688 , w_689 , 
		w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , w_696 , w_697 , w_698 , w_699 , 
		w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , w_706 , w_707 , w_708 , w_709 , 
		w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , w_716 , w_717 , w_718 , w_719 , 
		w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , w_726 , w_727 , w_728 , w_729 , 
		w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , w_736 , w_737 , w_738 , w_739 , 
		w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , w_746 , w_747 , w_748 , w_749 , 
		w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , w_756 , w_757 , w_758 , w_759 , 
		w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , w_766 , w_767 , w_768 , w_769 , 
		w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , w_776 , w_777 , w_778 , w_779 , 
		w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , w_786 , w_787 , w_788 , w_789 , 
		w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , w_796 , w_797 , w_798 , w_799 , 
		w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , w_806 , w_807 , w_808 , w_809 , 
		w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , w_816 , w_817 , w_818 , w_819 , 
		w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , w_826 , w_827 , w_828 , w_829 , 
		w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , w_836 , w_837 , w_838 , w_839 , 
		w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , w_846 , w_847 , w_848 , w_849 , 
		w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , w_856 , w_857 , w_858 , w_859 , 
		w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , w_866 , w_867 , w_868 , w_869 , 
		w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , w_876 , w_877 , w_878 , w_879 , 
		w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , w_886 , w_887 , w_888 , w_889 , 
		w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , w_896 , w_897 , w_898 , w_899 , 
		w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , w_906 , w_907 , w_908 , w_909 , 
		w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , w_916 , w_917 , w_918 , w_919 , 
		w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , w_926 , w_927 , w_928 , w_929 , 
		w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , w_936 , w_937 , w_938 , w_939 , 
		w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , w_946 , w_947 , w_948 , w_949 , 
		w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , w_956 , w_957 , w_958 , w_959 , 
		w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , w_966 , w_967 , w_968 , w_969 , 
		w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , w_976 , w_977 , w_978 , w_979 , 
		w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , w_986 , w_987 , w_988 , w_989 , 
		w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , w_996 , w_997 , w_998 , w_999 , 
		w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , w_1006 , w_1007 , w_1008 , w_1009 , 
		w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , w_1016 , w_1017 , w_1018 , w_1019 , 
		w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , w_1026 , w_1027 , w_1028 , w_1029 , 
		w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , w_1036 , w_1037 , w_1038 , w_1039 , 
		w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , w_1046 , w_1047 , w_1048 , w_1049 , 
		w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , w_1056 , w_1057 , w_1058 , w_1059 , 
		w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , w_1066 , w_1067 , w_1068 , w_1069 , 
		w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , w_1076 , w_1077 , w_1078 , w_1079 , 
		w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , w_1086 , w_1087 , w_1088 , w_1089 , 
		w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , w_1096 , w_1097 , w_1098 , w_1099 , 
		w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , w_1106 , w_1107 , w_1108 , w_1109 , 
		w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , w_1116 , w_1117 , w_1118 , w_1119 , 
		w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , w_1126 , w_1127 , w_1128 , w_1129 , 
		w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , w_1136 , w_1137 , w_1138 , w_1139 , 
		w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , w_1146 , w_1147 , w_1148 , w_1149 , 
		w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , w_1156 , w_1157 , w_1158 , w_1159 , 
		w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , w_1166 , w_1167 , w_1168 , w_1169 , 
		w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , w_1176 , w_1177 , w_1178 , w_1179 , 
		w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , w_1186 , w_1187 , w_1188 , w_1189 , 
		w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , w_1196 , w_1197 , w_1198 , w_1199 , 
		w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , w_1206 , w_1207 , w_1208 , w_1209 , 
		w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , w_1216 , w_1217 , w_1218 , w_1219 , 
		w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , w_1226 , w_1227 , w_1228 , w_1229 , 
		w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , w_1236 , w_1237 , w_1238 , w_1239 , 
		w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , w_1246 , w_1247 , w_1248 , w_1249 , 
		w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , w_1256 , w_1257 , w_1258 , w_1259 , 
		w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , w_1266 , w_1267 , w_1268 , w_1269 , 
		w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , w_1276 , w_1277 , w_1278 , w_1279 , 
		w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , w_1286 , w_1287 , w_1288 , w_1289 , 
		w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , w_1296 , w_1297 ;
buf ( \O[19]_b1 , \675_Z[19]_b1 );
buf ( \O[19]_b0 , \675_Z[19]_b0 );
buf ( \O[18]_b1 , \677_Z[18]_b1 );
buf ( \O[18]_b0 , \677_Z[18]_b0 );
buf ( \O[17]_b1 , \679_Z[17]_b1 );
buf ( \O[17]_b0 , \679_Z[17]_b0 );
buf ( \O[16]_b1 , \681_Z[16]_b1 );
buf ( \O[16]_b0 , \681_Z[16]_b0 );
buf ( \O[15]_b1 , \683_Z[15]_b1 );
buf ( \O[15]_b0 , \683_Z[15]_b0 );
buf ( \O[14]_b1 , \685_Z[14]_b1 );
buf ( \O[14]_b0 , \685_Z[14]_b0 );
buf ( \O[13]_b1 , \687_Z[13]_b1 );
buf ( \O[13]_b0 , \687_Z[13]_b0 );
buf ( \O[12]_b1 , \689_Z[12]_b1 );
buf ( \O[12]_b0 , \689_Z[12]_b0 );
buf ( \O[11]_b1 , \691_Z[11]_b1 );
buf ( \O[11]_b0 , \691_Z[11]_b0 );
buf ( \O[10]_b1 , \693_Z[10]_b1 );
buf ( \O[10]_b0 , \693_Z[10]_b0 );
buf ( \O[9]_b1 , \695_Z[9]_b1 );
buf ( \O[9]_b0 , \695_Z[9]_b0 );
buf ( \O[8]_b1 , \697_Z[8]_b1 );
buf ( \O[8]_b0 , \697_Z[8]_b0 );
buf ( \O[7]_b1 , \699_Z[7]_b1 );
buf ( \O[7]_b0 , \699_Z[7]_b0 );
buf ( \O[6]_b1 , \701_Z[6]_b1 );
buf ( \O[6]_b0 , \701_Z[6]_b0 );
buf ( \O[5]_b1 , \703_Z[5]_b1 );
buf ( \O[5]_b0 , \703_Z[5]_b0 );
buf ( \O[4]_b1 , \705_Z[4]_b1 );
buf ( \O[4]_b0 , \705_Z[4]_b0 );
buf ( \O[3]_b1 , \707_Z[3]_b1 );
buf ( \O[3]_b0 , \707_Z[3]_b0 );
buf ( \O[2]_b1 , \709_Z[2]_b1 );
buf ( \O[2]_b0 , \709_Z[2]_b0 );
buf ( \O[1]_b1 , \711_Z[1]_b1 );
buf ( \O[1]_b0 , \711_Z[1]_b0 );
buf ( \O[0]_b1 , \713_Z[0]_b1 );
buf ( \O[0]_b0 , \713_Z[0]_b0 );
buf ( \88_b1 , \I[1]_b1 );
not ( \88_b1 , w_0 );
not ( \88_b0 , w_1 );
and ( w_0 , w_1 , \I[1]_b0 );
or ( \90_b1 , \A[2][9]_b1 , \89_b1 );
not ( \89_b1 , w_2 );
and ( \90_b0 , \A[2][9]_b0 , w_3 );
and ( w_2 , w_3 , \89_b0 );
buf ( \91_b1 , \I[0]_b1 );
not ( \91_b1 , w_4 );
not ( \91_b0 , w_5 );
and ( w_4 , w_5 , \I[0]_b0 );
or ( \93_b1 , \A[1][9]_b1 , \92_b1 );
not ( \92_b1 , w_6 );
and ( \93_b0 , \A[1][9]_b0 , w_7 );
and ( w_6 , w_7 , \92_b0 );
or ( \95_b1 , \A[0][9]_b1 , \94_b1 );
not ( \94_b1 , w_8 );
and ( \95_b0 , \A[0][9]_b0 , w_9 );
and ( w_8 , w_9 , \94_b0 );
buf ( \97_b1 , \I[2]_b1 );
buf ( \97_b0 , \I[2]_b0 );
buf ( \98_b1 , \I[3]_b1 );
buf ( \98_b0 , \I[3]_b0 );
buf ( \99_b1 , \I[4]_b1 );
buf ( \99_b0 , \I[4]_b0 );
buf ( \100_b1 , \I[5]_b1 );
buf ( \100_b0 , \I[5]_b0 );
buf ( \101_b1 , \I[6]_b1 );
buf ( \101_b0 , \I[6]_b0 );
buf ( \102_b1 , \I[7]_b1 );
buf ( \102_b0 , \I[7]_b0 );
buf ( \103_b1 , \I[1]_b1 );
buf ( \103_b0 , \I[1]_b0 );
buf ( \104_b1 , \I[0]_b1 );
buf ( \104_b0 , \I[0]_b0 );
or ( \105_b1 , \103_b1 , \104_b1 );
not ( \104_b1 , w_10 );
and ( \105_b0 , \103_b0 , w_11 );
and ( w_10 , w_11 , \104_b0 );
buf ( \107_b1 , \106_b1 );
buf ( \107_b0 , \106_b0 );
and ( \108_b1 , \96_b1 , w_12 );
xor ( w_12 , \96_b0 , \107_b1 );
not ( \107_b1 , w_13 );
and ( \108_b0 , w_13 , \107_b0 );
buf ( \109_A[9]_b1 , \108_b1 );
buf ( \109_A[9]_b0 , \108_b0 );
or ( \110_b1 , \A[2][8]_b1 , \89_b1 );
not ( \89_b1 , w_14 );
and ( \110_b0 , \A[2][8]_b0 , w_15 );
and ( w_14 , w_15 , \89_b0 );
or ( \111_b1 , \A[1][8]_b1 , \92_b1 );
not ( \92_b1 , w_16 );
and ( \111_b0 , \A[1][8]_b0 , w_17 );
and ( w_16 , w_17 , \92_b0 );
or ( \112_b1 , \A[0][8]_b1 , \94_b1 );
not ( \94_b1 , w_18 );
and ( \112_b0 , \A[0][8]_b0 , w_19 );
and ( w_18 , w_19 , \94_b0 );
and ( \114_b1 , \113_b1 , w_20 );
xor ( w_20 , \113_b0 , \107_b1 );
not ( \107_b1 , w_21 );
and ( \114_b0 , w_21 , \107_b0 );
buf ( \115_A[8]_b1 , \114_b1 );
buf ( \115_A[8]_b0 , \114_b0 );
or ( \116_b1 , \A[2][7]_b1 , \89_b1 );
not ( \89_b1 , w_22 );
and ( \116_b0 , \A[2][7]_b0 , w_23 );
and ( w_22 , w_23 , \89_b0 );
or ( \117_b1 , \A[1][7]_b1 , \92_b1 );
not ( \92_b1 , w_24 );
and ( \117_b0 , \A[1][7]_b0 , w_25 );
and ( w_24 , w_25 , \92_b0 );
or ( \118_b1 , \A[0][7]_b1 , \94_b1 );
not ( \94_b1 , w_26 );
and ( \118_b0 , \A[0][7]_b0 , w_27 );
and ( w_26 , w_27 , \94_b0 );
and ( \120_b1 , \119_b1 , w_28 );
xor ( w_28 , \119_b0 , \107_b1 );
not ( \107_b1 , w_29 );
and ( \120_b0 , w_29 , \107_b0 );
buf ( \121_A[7]_b1 , \120_b1 );
buf ( \121_A[7]_b0 , \120_b0 );
or ( \122_b1 , \A[2][6]_b1 , \89_b1 );
not ( \89_b1 , w_30 );
and ( \122_b0 , \A[2][6]_b0 , w_31 );
and ( w_30 , w_31 , \89_b0 );
or ( \123_b1 , \A[1][6]_b1 , \92_b1 );
not ( \92_b1 , w_32 );
and ( \123_b0 , \A[1][6]_b0 , w_33 );
and ( w_32 , w_33 , \92_b0 );
or ( \124_b1 , \A[0][6]_b1 , \94_b1 );
not ( \94_b1 , w_34 );
and ( \124_b0 , \A[0][6]_b0 , w_35 );
and ( w_34 , w_35 , \94_b0 );
and ( \126_b1 , \125_b1 , w_36 );
xor ( w_36 , \125_b0 , \107_b1 );
not ( \107_b1 , w_37 );
and ( \126_b0 , w_37 , \107_b0 );
buf ( \127_A[6]_b1 , \126_b1 );
buf ( \127_A[6]_b0 , \126_b0 );
or ( \128_b1 , \A[2][5]_b1 , \89_b1 );
not ( \89_b1 , w_38 );
and ( \128_b0 , \A[2][5]_b0 , w_39 );
and ( w_38 , w_39 , \89_b0 );
or ( \129_b1 , \A[1][5]_b1 , \92_b1 );
not ( \92_b1 , w_40 );
and ( \129_b0 , \A[1][5]_b0 , w_41 );
and ( w_40 , w_41 , \92_b0 );
or ( \130_b1 , \A[0][5]_b1 , \94_b1 );
not ( \94_b1 , w_42 );
and ( \130_b0 , \A[0][5]_b0 , w_43 );
and ( w_42 , w_43 , \94_b0 );
and ( \132_b1 , \131_b1 , w_44 );
xor ( w_44 , \131_b0 , \107_b1 );
not ( \107_b1 , w_45 );
and ( \132_b0 , w_45 , \107_b0 );
buf ( \133_A[5]_b1 , \132_b1 );
buf ( \133_A[5]_b0 , \132_b0 );
or ( \134_b1 , \A[2][4]_b1 , \89_b1 );
not ( \89_b1 , w_46 );
and ( \134_b0 , \A[2][4]_b0 , w_47 );
and ( w_46 , w_47 , \89_b0 );
or ( \135_b1 , \A[1][4]_b1 , \92_b1 );
not ( \92_b1 , w_48 );
and ( \135_b0 , \A[1][4]_b0 , w_49 );
and ( w_48 , w_49 , \92_b0 );
or ( \136_b1 , \A[0][4]_b1 , \94_b1 );
not ( \94_b1 , w_50 );
and ( \136_b0 , \A[0][4]_b0 , w_51 );
and ( w_50 , w_51 , \94_b0 );
and ( \138_b1 , \137_b1 , w_52 );
xor ( w_52 , \137_b0 , \107_b1 );
not ( \107_b1 , w_53 );
and ( \138_b0 , w_53 , \107_b0 );
buf ( \139_A[4]_b1 , \138_b1 );
buf ( \139_A[4]_b0 , \138_b0 );
or ( \140_b1 , \A[2][3]_b1 , \89_b1 );
not ( \89_b1 , w_54 );
and ( \140_b0 , \A[2][3]_b0 , w_55 );
and ( w_54 , w_55 , \89_b0 );
or ( \141_b1 , \A[1][3]_b1 , \92_b1 );
not ( \92_b1 , w_56 );
and ( \141_b0 , \A[1][3]_b0 , w_57 );
and ( w_56 , w_57 , \92_b0 );
or ( \142_b1 , \A[0][3]_b1 , \94_b1 );
not ( \94_b1 , w_58 );
and ( \142_b0 , \A[0][3]_b0 , w_59 );
and ( w_58 , w_59 , \94_b0 );
and ( \144_b1 , \143_b1 , w_60 );
xor ( w_60 , \143_b0 , \107_b1 );
not ( \107_b1 , w_61 );
and ( \144_b0 , w_61 , \107_b0 );
buf ( \145_A[3]_b1 , \144_b1 );
buf ( \145_A[3]_b0 , \144_b0 );
or ( \146_b1 , \A[2][2]_b1 , \89_b1 );
not ( \89_b1 , w_62 );
and ( \146_b0 , \A[2][2]_b0 , w_63 );
and ( w_62 , w_63 , \89_b0 );
or ( \147_b1 , \A[1][2]_b1 , \92_b1 );
not ( \92_b1 , w_64 );
and ( \147_b0 , \A[1][2]_b0 , w_65 );
and ( w_64 , w_65 , \92_b0 );
or ( \148_b1 , \A[0][2]_b1 , \94_b1 );
not ( \94_b1 , w_66 );
and ( \148_b0 , \A[0][2]_b0 , w_67 );
and ( w_66 , w_67 , \94_b0 );
and ( \150_b1 , \149_b1 , w_68 );
xor ( w_68 , \149_b0 , \107_b1 );
not ( \107_b1 , w_69 );
and ( \150_b0 , w_69 , \107_b0 );
buf ( \151_A[2]_b1 , \150_b1 );
buf ( \151_A[2]_b0 , \150_b0 );
or ( \152_b1 , \A[2][1]_b1 , \89_b1 );
not ( \89_b1 , w_70 );
and ( \152_b0 , \A[2][1]_b0 , w_71 );
and ( w_70 , w_71 , \89_b0 );
or ( \153_b1 , \A[1][1]_b1 , \92_b1 );
not ( \92_b1 , w_72 );
and ( \153_b0 , \A[1][1]_b0 , w_73 );
and ( w_72 , w_73 , \92_b0 );
or ( \154_b1 , \A[0][1]_b1 , \94_b1 );
not ( \94_b1 , w_74 );
and ( \154_b0 , \A[0][1]_b0 , w_75 );
and ( w_74 , w_75 , \94_b0 );
and ( \156_b1 , \155_b1 , w_76 );
xor ( w_76 , \155_b0 , \107_b1 );
not ( \107_b1 , w_77 );
and ( \156_b0 , w_77 , \107_b0 );
buf ( \157_A[1]_b1 , \156_b1 );
buf ( \157_A[1]_b0 , \156_b0 );
or ( \158_b1 , \A[2][0]_b1 , \89_b1 );
not ( \89_b1 , w_78 );
and ( \158_b0 , \A[2][0]_b0 , w_79 );
and ( w_78 , w_79 , \89_b0 );
or ( \159_b1 , \A[1][0]_b1 , \92_b1 );
not ( \92_b1 , w_80 );
and ( \159_b0 , \A[1][0]_b0 , w_81 );
and ( w_80 , w_81 , \92_b0 );
or ( \160_b1 , \A[0][0]_b1 , \94_b1 );
not ( \94_b1 , w_82 );
and ( \160_b0 , \A[0][0]_b0 , w_83 );
and ( w_82 , w_83 , \94_b0 );
and ( \162_b1 , \161_b1 , w_84 );
xor ( w_84 , \161_b0 , \107_b1 );
not ( \107_b1 , w_85 );
and ( \162_b0 , w_85 , \107_b0 );
buf ( \163_A[0]_b1 , \162_b1 );
buf ( \163_A[0]_b0 , \162_b0 );
buf ( \164_B[9]_b1 , \B[9]_b1 );
buf ( \164_B[9]_b0 , \B[9]_b0 );
buf ( \165_B[8]_b1 , \B[8]_b1 );
buf ( \165_B[8]_b0 , \B[8]_b0 );
buf ( \166_B[7]_b1 , \B[7]_b1 );
buf ( \166_B[7]_b0 , \B[7]_b0 );
buf ( \167_B[6]_b1 , \B[6]_b1 );
buf ( \167_B[6]_b0 , \B[6]_b0 );
buf ( \168_B[5]_b1 , \B[5]_b1 );
buf ( \168_B[5]_b0 , \B[5]_b0 );
buf ( \169_B[4]_b1 , \B[4]_b1 );
buf ( \169_B[4]_b0 , \B[4]_b0 );
buf ( \170_B[3]_b1 , \B[3]_b1 );
buf ( \170_B[3]_b0 , \B[3]_b0 );
buf ( \171_B[2]_b1 , \B[2]_b1 );
buf ( \171_B[2]_b0 , \B[2]_b0 );
buf ( \172_B[1]_b1 , \B[1]_b1 );
buf ( \172_B[1]_b0 , \B[1]_b0 );
buf ( \173_B[0]_b1 , \B[0]_b1 );
buf ( \173_B[0]_b0 , \B[0]_b0 );
or ( \174_b1 , \109_A[9]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_86 );
and ( \174_b0 , \109_A[9]_b0 , w_87 );
and ( w_86 , w_87 , \172_B[1]_b0 );
or ( \175_b1 , \109_A[9]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_88 );
and ( \175_b0 , \109_A[9]_b0 , w_89 );
and ( w_88 , w_89 , \173_B[0]_b0 );
or ( \176_b1 , \115_A[8]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_90 );
and ( \176_b0 , \115_A[8]_b0 , w_91 );
and ( w_90 , w_91 , \172_B[1]_b0 );
or ( \177_b1 , \175_b1 , \176_b1 );
not ( \176_b1 , w_92 );
and ( \177_b0 , \175_b0 , w_93 );
and ( w_92 , w_93 , \176_b0 );
or ( \178_b1 , \175_b1 , \176_b1 );
xor ( \178_b0 , \175_b0 , w_94 );
not ( w_94 , w_95 );
and ( w_95 , \176_b1 , \176_b0 );
or ( \179_b1 , \115_A[8]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_96 );
and ( \179_b0 , \115_A[8]_b0 , w_97 );
and ( w_96 , w_97 , \173_B[0]_b0 );
or ( \180_b1 , \121_A[7]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_98 );
and ( \180_b0 , \121_A[7]_b0 , w_99 );
and ( w_98 , w_99 , \172_B[1]_b0 );
or ( \181_b1 , \179_b1 , \180_b1 );
not ( \180_b1 , w_100 );
and ( \181_b0 , \179_b0 , w_101 );
and ( w_100 , w_101 , \180_b0 );
or ( \182_b1 , \179_b1 , \180_b1 );
xor ( \182_b0 , \179_b0 , w_102 );
not ( w_102 , w_103 );
and ( w_103 , \180_b1 , \180_b0 );
or ( \183_b1 , \121_A[7]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_104 );
and ( \183_b0 , \121_A[7]_b0 , w_105 );
and ( w_104 , w_105 , \173_B[0]_b0 );
or ( \184_b1 , \127_A[6]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_106 );
and ( \184_b0 , \127_A[6]_b0 , w_107 );
and ( w_106 , w_107 , \172_B[1]_b0 );
or ( \185_b1 , \183_b1 , \184_b1 );
not ( \184_b1 , w_108 );
and ( \185_b0 , \183_b0 , w_109 );
and ( w_108 , w_109 , \184_b0 );
or ( \186_b1 , \183_b1 , \184_b1 );
xor ( \186_b0 , \183_b0 , w_110 );
not ( w_110 , w_111 );
and ( w_111 , \184_b1 , \184_b0 );
or ( \187_b1 , \127_A[6]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_112 );
and ( \187_b0 , \127_A[6]_b0 , w_113 );
and ( w_112 , w_113 , \173_B[0]_b0 );
or ( \188_b1 , \133_A[5]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_114 );
and ( \188_b0 , \133_A[5]_b0 , w_115 );
and ( w_114 , w_115 , \172_B[1]_b0 );
or ( \189_b1 , \187_b1 , \188_b1 );
not ( \188_b1 , w_116 );
and ( \189_b0 , \187_b0 , w_117 );
and ( w_116 , w_117 , \188_b0 );
or ( \190_b1 , \187_b1 , \188_b1 );
xor ( \190_b0 , \187_b0 , w_118 );
not ( w_118 , w_119 );
and ( w_119 , \188_b1 , \188_b0 );
or ( \191_b1 , \133_A[5]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_120 );
and ( \191_b0 , \133_A[5]_b0 , w_121 );
and ( w_120 , w_121 , \173_B[0]_b0 );
or ( \192_b1 , \139_A[4]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_122 );
and ( \192_b0 , \139_A[4]_b0 , w_123 );
and ( w_122 , w_123 , \172_B[1]_b0 );
or ( \193_b1 , \191_b1 , \192_b1 );
not ( \192_b1 , w_124 );
and ( \193_b0 , \191_b0 , w_125 );
and ( w_124 , w_125 , \192_b0 );
or ( \194_b1 , \191_b1 , \192_b1 );
xor ( \194_b0 , \191_b0 , w_126 );
not ( w_126 , w_127 );
and ( w_127 , \192_b1 , \192_b0 );
or ( \195_b1 , \139_A[4]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_128 );
and ( \195_b0 , \139_A[4]_b0 , w_129 );
and ( w_128 , w_129 , \173_B[0]_b0 );
or ( \196_b1 , \145_A[3]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_130 );
and ( \196_b0 , \145_A[3]_b0 , w_131 );
and ( w_130 , w_131 , \172_B[1]_b0 );
or ( \197_b1 , \195_b1 , \196_b1 );
not ( \196_b1 , w_132 );
and ( \197_b0 , \195_b0 , w_133 );
and ( w_132 , w_133 , \196_b0 );
or ( \198_b1 , \195_b1 , \196_b1 );
xor ( \198_b0 , \195_b0 , w_134 );
not ( w_134 , w_135 );
and ( w_135 , \196_b1 , \196_b0 );
or ( \199_b1 , \145_A[3]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_136 );
and ( \199_b0 , \145_A[3]_b0 , w_137 );
and ( w_136 , w_137 , \173_B[0]_b0 );
or ( \200_b1 , \151_A[2]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_138 );
and ( \200_b0 , \151_A[2]_b0 , w_139 );
and ( w_138 , w_139 , \172_B[1]_b0 );
or ( \201_b1 , \199_b1 , \200_b1 );
not ( \200_b1 , w_140 );
and ( \201_b0 , \199_b0 , w_141 );
and ( w_140 , w_141 , \200_b0 );
or ( \202_b1 , \199_b1 , \200_b1 );
xor ( \202_b0 , \199_b0 , w_142 );
not ( w_142 , w_143 );
and ( w_143 , \200_b1 , \200_b0 );
or ( \203_b1 , \151_A[2]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_144 );
and ( \203_b0 , \151_A[2]_b0 , w_145 );
and ( w_144 , w_145 , \173_B[0]_b0 );
or ( \204_b1 , \157_A[1]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_146 );
and ( \204_b0 , \157_A[1]_b0 , w_147 );
and ( w_146 , w_147 , \172_B[1]_b0 );
or ( \205_b1 , \203_b1 , \204_b1 );
not ( \204_b1 , w_148 );
and ( \205_b0 , \203_b0 , w_149 );
and ( w_148 , w_149 , \204_b0 );
or ( \206_b1 , \203_b1 , \204_b1 );
xor ( \206_b0 , \203_b0 , w_150 );
not ( w_150 , w_151 );
and ( w_151 , \204_b1 , \204_b0 );
or ( \207_b1 , \157_A[1]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_152 );
and ( \207_b0 , \157_A[1]_b0 , w_153 );
and ( w_152 , w_153 , \173_B[0]_b0 );
or ( \208_b1 , \163_A[0]_b1 , \172_B[1]_b1 );
not ( \172_B[1]_b1 , w_154 );
and ( \208_b0 , \163_A[0]_b0 , w_155 );
and ( w_154 , w_155 , \172_B[1]_b0 );
or ( \209_b1 , \207_b1 , \208_b1 );
not ( \208_b1 , w_156 );
and ( \209_b0 , \207_b0 , w_157 );
and ( w_156 , w_157 , \208_b0 );
or ( \210_b1 , \206_b1 , \209_b1 );
not ( \209_b1 , w_158 );
and ( \210_b0 , \206_b0 , w_159 );
and ( w_158 , w_159 , \209_b0 );
or ( \211_b1 , \205_b1 , w_160 );
or ( \211_b0 , \205_b0 , \210_b0 );
not ( \210_b0 , w_161 );
and ( w_161 , w_160 , \210_b1 );
or ( \212_b1 , \202_b1 , \211_b1 );
not ( \211_b1 , w_162 );
and ( \212_b0 , \202_b0 , w_163 );
and ( w_162 , w_163 , \211_b0 );
or ( \213_b1 , \201_b1 , w_164 );
or ( \213_b0 , \201_b0 , \212_b0 );
not ( \212_b0 , w_165 );
and ( w_165 , w_164 , \212_b1 );
or ( \214_b1 , \198_b1 , \213_b1 );
not ( \213_b1 , w_166 );
and ( \214_b0 , \198_b0 , w_167 );
and ( w_166 , w_167 , \213_b0 );
or ( \215_b1 , \197_b1 , w_168 );
or ( \215_b0 , \197_b0 , \214_b0 );
not ( \214_b0 , w_169 );
and ( w_169 , w_168 , \214_b1 );
or ( \216_b1 , \194_b1 , \215_b1 );
not ( \215_b1 , w_170 );
and ( \216_b0 , \194_b0 , w_171 );
and ( w_170 , w_171 , \215_b0 );
or ( \217_b1 , \193_b1 , w_172 );
or ( \217_b0 , \193_b0 , \216_b0 );
not ( \216_b0 , w_173 );
and ( w_173 , w_172 , \216_b1 );
or ( \218_b1 , \190_b1 , \217_b1 );
not ( \217_b1 , w_174 );
and ( \218_b0 , \190_b0 , w_175 );
and ( w_174 , w_175 , \217_b0 );
or ( \219_b1 , \189_b1 , w_176 );
or ( \219_b0 , \189_b0 , \218_b0 );
not ( \218_b0 , w_177 );
and ( w_177 , w_176 , \218_b1 );
or ( \220_b1 , \186_b1 , \219_b1 );
not ( \219_b1 , w_178 );
and ( \220_b0 , \186_b0 , w_179 );
and ( w_178 , w_179 , \219_b0 );
or ( \221_b1 , \185_b1 , w_180 );
or ( \221_b0 , \185_b0 , \220_b0 );
not ( \220_b0 , w_181 );
and ( w_181 , w_180 , \220_b1 );
or ( \222_b1 , \182_b1 , \221_b1 );
not ( \221_b1 , w_182 );
and ( \222_b0 , \182_b0 , w_183 );
and ( w_182 , w_183 , \221_b0 );
or ( \223_b1 , \181_b1 , w_184 );
or ( \223_b0 , \181_b0 , \222_b0 );
not ( \222_b0 , w_185 );
and ( w_185 , w_184 , \222_b1 );
or ( \224_b1 , \178_b1 , \223_b1 );
not ( \223_b1 , w_186 );
and ( \224_b0 , \178_b0 , w_187 );
and ( w_186 , w_187 , \223_b0 );
or ( \225_b1 , \177_b1 , w_188 );
or ( \225_b0 , \177_b0 , \224_b0 );
not ( \224_b0 , w_189 );
and ( w_189 , w_188 , \224_b1 );
or ( \226_b1 , \174_b1 , \225_b1 );
not ( \225_b1 , w_190 );
and ( \226_b0 , \174_b0 , w_191 );
and ( w_190 , w_191 , \225_b0 );
or ( \227_b1 , \109_A[9]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_192 );
and ( \227_b0 , \109_A[9]_b0 , w_193 );
and ( w_192 , w_193 , \171_B[2]_b0 );
or ( \228_b1 , \226_b1 , \227_b1 );
not ( \227_b1 , w_194 );
and ( \228_b0 , \226_b0 , w_195 );
and ( w_194 , w_195 , \227_b0 );
or ( \229_b1 , \226_b1 , \227_b1 );
xor ( \229_b0 , \226_b0 , w_196 );
not ( w_196 , w_197 );
and ( w_197 , \227_b1 , \227_b0 );
or ( \230_b1 , \174_b1 , \225_b1 );
xor ( \230_b0 , \174_b0 , w_198 );
not ( w_198 , w_199 );
and ( w_199 , \225_b1 , \225_b0 );
or ( \231_b1 , \115_A[8]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_200 );
and ( \231_b0 , \115_A[8]_b0 , w_201 );
and ( w_200 , w_201 , \171_B[2]_b0 );
or ( \232_b1 , \230_b1 , \231_b1 );
not ( \231_b1 , w_202 );
and ( \232_b0 , \230_b0 , w_203 );
and ( w_202 , w_203 , \231_b0 );
or ( \233_b1 , \230_b1 , \231_b1 );
xor ( \233_b0 , \230_b0 , w_204 );
not ( w_204 , w_205 );
and ( w_205 , \231_b1 , \231_b0 );
or ( \234_b1 , \178_b1 , \223_b1 );
xor ( \234_b0 , \178_b0 , w_206 );
not ( w_206 , w_207 );
and ( w_207 , \223_b1 , \223_b0 );
or ( \235_b1 , \121_A[7]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_208 );
and ( \235_b0 , \121_A[7]_b0 , w_209 );
and ( w_208 , w_209 , \171_B[2]_b0 );
or ( \236_b1 , \234_b1 , \235_b1 );
not ( \235_b1 , w_210 );
and ( \236_b0 , \234_b0 , w_211 );
and ( w_210 , w_211 , \235_b0 );
or ( \237_b1 , \234_b1 , \235_b1 );
xor ( \237_b0 , \234_b0 , w_212 );
not ( w_212 , w_213 );
and ( w_213 , \235_b1 , \235_b0 );
or ( \238_b1 , \182_b1 , \221_b1 );
xor ( \238_b0 , \182_b0 , w_214 );
not ( w_214 , w_215 );
and ( w_215 , \221_b1 , \221_b0 );
or ( \239_b1 , \127_A[6]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_216 );
and ( \239_b0 , \127_A[6]_b0 , w_217 );
and ( w_216 , w_217 , \171_B[2]_b0 );
or ( \240_b1 , \238_b1 , \239_b1 );
not ( \239_b1 , w_218 );
and ( \240_b0 , \238_b0 , w_219 );
and ( w_218 , w_219 , \239_b0 );
or ( \241_b1 , \238_b1 , \239_b1 );
xor ( \241_b0 , \238_b0 , w_220 );
not ( w_220 , w_221 );
and ( w_221 , \239_b1 , \239_b0 );
or ( \242_b1 , \186_b1 , \219_b1 );
xor ( \242_b0 , \186_b0 , w_222 );
not ( w_222 , w_223 );
and ( w_223 , \219_b1 , \219_b0 );
or ( \243_b1 , \133_A[5]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_224 );
and ( \243_b0 , \133_A[5]_b0 , w_225 );
and ( w_224 , w_225 , \171_B[2]_b0 );
or ( \244_b1 , \242_b1 , \243_b1 );
not ( \243_b1 , w_226 );
and ( \244_b0 , \242_b0 , w_227 );
and ( w_226 , w_227 , \243_b0 );
or ( \245_b1 , \242_b1 , \243_b1 );
xor ( \245_b0 , \242_b0 , w_228 );
not ( w_228 , w_229 );
and ( w_229 , \243_b1 , \243_b0 );
or ( \246_b1 , \190_b1 , \217_b1 );
xor ( \246_b0 , \190_b0 , w_230 );
not ( w_230 , w_231 );
and ( w_231 , \217_b1 , \217_b0 );
or ( \247_b1 , \139_A[4]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_232 );
and ( \247_b0 , \139_A[4]_b0 , w_233 );
and ( w_232 , w_233 , \171_B[2]_b0 );
or ( \248_b1 , \246_b1 , \247_b1 );
not ( \247_b1 , w_234 );
and ( \248_b0 , \246_b0 , w_235 );
and ( w_234 , w_235 , \247_b0 );
or ( \249_b1 , \246_b1 , \247_b1 );
xor ( \249_b0 , \246_b0 , w_236 );
not ( w_236 , w_237 );
and ( w_237 , \247_b1 , \247_b0 );
or ( \250_b1 , \194_b1 , \215_b1 );
xor ( \250_b0 , \194_b0 , w_238 );
not ( w_238 , w_239 );
and ( w_239 , \215_b1 , \215_b0 );
or ( \251_b1 , \145_A[3]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_240 );
and ( \251_b0 , \145_A[3]_b0 , w_241 );
and ( w_240 , w_241 , \171_B[2]_b0 );
or ( \252_b1 , \250_b1 , \251_b1 );
not ( \251_b1 , w_242 );
and ( \252_b0 , \250_b0 , w_243 );
and ( w_242 , w_243 , \251_b0 );
or ( \253_b1 , \250_b1 , \251_b1 );
xor ( \253_b0 , \250_b0 , w_244 );
not ( w_244 , w_245 );
and ( w_245 , \251_b1 , \251_b0 );
or ( \254_b1 , \198_b1 , \213_b1 );
xor ( \254_b0 , \198_b0 , w_246 );
not ( w_246 , w_247 );
and ( w_247 , \213_b1 , \213_b0 );
or ( \255_b1 , \151_A[2]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_248 );
and ( \255_b0 , \151_A[2]_b0 , w_249 );
and ( w_248 , w_249 , \171_B[2]_b0 );
or ( \256_b1 , \254_b1 , \255_b1 );
not ( \255_b1 , w_250 );
and ( \256_b0 , \254_b0 , w_251 );
and ( w_250 , w_251 , \255_b0 );
or ( \257_b1 , \254_b1 , \255_b1 );
xor ( \257_b0 , \254_b0 , w_252 );
not ( w_252 , w_253 );
and ( w_253 , \255_b1 , \255_b0 );
or ( \258_b1 , \202_b1 , \211_b1 );
xor ( \258_b0 , \202_b0 , w_254 );
not ( w_254 , w_255 );
and ( w_255 , \211_b1 , \211_b0 );
or ( \259_b1 , \157_A[1]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_256 );
and ( \259_b0 , \157_A[1]_b0 , w_257 );
and ( w_256 , w_257 , \171_B[2]_b0 );
or ( \260_b1 , \258_b1 , \259_b1 );
not ( \259_b1 , w_258 );
and ( \260_b0 , \258_b0 , w_259 );
and ( w_258 , w_259 , \259_b0 );
or ( \261_b1 , \258_b1 , \259_b1 );
xor ( \261_b0 , \258_b0 , w_260 );
not ( w_260 , w_261 );
and ( w_261 , \259_b1 , \259_b0 );
or ( \262_b1 , \206_b1 , \209_b1 );
xor ( \262_b0 , \206_b0 , w_262 );
not ( w_262 , w_263 );
and ( w_263 , \209_b1 , \209_b0 );
or ( \263_b1 , \163_A[0]_b1 , \171_B[2]_b1 );
not ( \171_B[2]_b1 , w_264 );
and ( \263_b0 , \163_A[0]_b0 , w_265 );
and ( w_264 , w_265 , \171_B[2]_b0 );
or ( \264_b1 , \262_b1 , \263_b1 );
not ( \263_b1 , w_266 );
and ( \264_b0 , \262_b0 , w_267 );
and ( w_266 , w_267 , \263_b0 );
or ( \265_b1 , \261_b1 , \264_b1 );
not ( \264_b1 , w_268 );
and ( \265_b0 , \261_b0 , w_269 );
and ( w_268 , w_269 , \264_b0 );
or ( \266_b1 , \260_b1 , w_270 );
or ( \266_b0 , \260_b0 , \265_b0 );
not ( \265_b0 , w_271 );
and ( w_271 , w_270 , \265_b1 );
or ( \267_b1 , \257_b1 , \266_b1 );
not ( \266_b1 , w_272 );
and ( \267_b0 , \257_b0 , w_273 );
and ( w_272 , w_273 , \266_b0 );
or ( \268_b1 , \256_b1 , w_274 );
or ( \268_b0 , \256_b0 , \267_b0 );
not ( \267_b0 , w_275 );
and ( w_275 , w_274 , \267_b1 );
or ( \269_b1 , \253_b1 , \268_b1 );
not ( \268_b1 , w_276 );
and ( \269_b0 , \253_b0 , w_277 );
and ( w_276 , w_277 , \268_b0 );
or ( \270_b1 , \252_b1 , w_278 );
or ( \270_b0 , \252_b0 , \269_b0 );
not ( \269_b0 , w_279 );
and ( w_279 , w_278 , \269_b1 );
or ( \271_b1 , \249_b1 , \270_b1 );
not ( \270_b1 , w_280 );
and ( \271_b0 , \249_b0 , w_281 );
and ( w_280 , w_281 , \270_b0 );
or ( \272_b1 , \248_b1 , w_282 );
or ( \272_b0 , \248_b0 , \271_b0 );
not ( \271_b0 , w_283 );
and ( w_283 , w_282 , \271_b1 );
or ( \273_b1 , \245_b1 , \272_b1 );
not ( \272_b1 , w_284 );
and ( \273_b0 , \245_b0 , w_285 );
and ( w_284 , w_285 , \272_b0 );
or ( \274_b1 , \244_b1 , w_286 );
or ( \274_b0 , \244_b0 , \273_b0 );
not ( \273_b0 , w_287 );
and ( w_287 , w_286 , \273_b1 );
or ( \275_b1 , \241_b1 , \274_b1 );
not ( \274_b1 , w_288 );
and ( \275_b0 , \241_b0 , w_289 );
and ( w_288 , w_289 , \274_b0 );
or ( \276_b1 , \240_b1 , w_290 );
or ( \276_b0 , \240_b0 , \275_b0 );
not ( \275_b0 , w_291 );
and ( w_291 , w_290 , \275_b1 );
or ( \277_b1 , \237_b1 , \276_b1 );
not ( \276_b1 , w_292 );
and ( \277_b0 , \237_b0 , w_293 );
and ( w_292 , w_293 , \276_b0 );
or ( \278_b1 , \236_b1 , w_294 );
or ( \278_b0 , \236_b0 , \277_b0 );
not ( \277_b0 , w_295 );
and ( w_295 , w_294 , \277_b1 );
or ( \279_b1 , \233_b1 , \278_b1 );
not ( \278_b1 , w_296 );
and ( \279_b0 , \233_b0 , w_297 );
and ( w_296 , w_297 , \278_b0 );
or ( \280_b1 , \232_b1 , w_298 );
or ( \280_b0 , \232_b0 , \279_b0 );
not ( \279_b0 , w_299 );
and ( w_299 , w_298 , \279_b1 );
or ( \281_b1 , \229_b1 , \280_b1 );
not ( \280_b1 , w_300 );
and ( \281_b0 , \229_b0 , w_301 );
and ( w_300 , w_301 , \280_b0 );
or ( \282_b1 , \228_b1 , w_302 );
or ( \282_b0 , \228_b0 , \281_b0 );
not ( \281_b0 , w_303 );
and ( w_303 , w_302 , \281_b1 );
or ( \283_b1 , \109_A[9]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_304 );
and ( \283_b0 , \109_A[9]_b0 , w_305 );
and ( w_304 , w_305 , \170_B[3]_b0 );
or ( \284_b1 , \282_b1 , \283_b1 );
not ( \283_b1 , w_306 );
and ( \284_b0 , \282_b0 , w_307 );
and ( w_306 , w_307 , \283_b0 );
or ( \285_b1 , \282_b1 , \283_b1 );
xor ( \285_b0 , \282_b0 , w_308 );
not ( w_308 , w_309 );
and ( w_309 , \283_b1 , \283_b0 );
or ( \286_b1 , \229_b1 , \280_b1 );
xor ( \286_b0 , \229_b0 , w_310 );
not ( w_310 , w_311 );
and ( w_311 , \280_b1 , \280_b0 );
or ( \287_b1 , \115_A[8]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_312 );
and ( \287_b0 , \115_A[8]_b0 , w_313 );
and ( w_312 , w_313 , \170_B[3]_b0 );
or ( \288_b1 , \286_b1 , \287_b1 );
not ( \287_b1 , w_314 );
and ( \288_b0 , \286_b0 , w_315 );
and ( w_314 , w_315 , \287_b0 );
or ( \289_b1 , \286_b1 , \287_b1 );
xor ( \289_b0 , \286_b0 , w_316 );
not ( w_316 , w_317 );
and ( w_317 , \287_b1 , \287_b0 );
or ( \290_b1 , \233_b1 , \278_b1 );
xor ( \290_b0 , \233_b0 , w_318 );
not ( w_318 , w_319 );
and ( w_319 , \278_b1 , \278_b0 );
or ( \291_b1 , \121_A[7]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_320 );
and ( \291_b0 , \121_A[7]_b0 , w_321 );
and ( w_320 , w_321 , \170_B[3]_b0 );
or ( \292_b1 , \290_b1 , \291_b1 );
not ( \291_b1 , w_322 );
and ( \292_b0 , \290_b0 , w_323 );
and ( w_322 , w_323 , \291_b0 );
or ( \293_b1 , \290_b1 , \291_b1 );
xor ( \293_b0 , \290_b0 , w_324 );
not ( w_324 , w_325 );
and ( w_325 , \291_b1 , \291_b0 );
or ( \294_b1 , \237_b1 , \276_b1 );
xor ( \294_b0 , \237_b0 , w_326 );
not ( w_326 , w_327 );
and ( w_327 , \276_b1 , \276_b0 );
or ( \295_b1 , \127_A[6]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_328 );
and ( \295_b0 , \127_A[6]_b0 , w_329 );
and ( w_328 , w_329 , \170_B[3]_b0 );
or ( \296_b1 , \294_b1 , \295_b1 );
not ( \295_b1 , w_330 );
and ( \296_b0 , \294_b0 , w_331 );
and ( w_330 , w_331 , \295_b0 );
or ( \297_b1 , \294_b1 , \295_b1 );
xor ( \297_b0 , \294_b0 , w_332 );
not ( w_332 , w_333 );
and ( w_333 , \295_b1 , \295_b0 );
or ( \298_b1 , \241_b1 , \274_b1 );
xor ( \298_b0 , \241_b0 , w_334 );
not ( w_334 , w_335 );
and ( w_335 , \274_b1 , \274_b0 );
or ( \299_b1 , \133_A[5]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_336 );
and ( \299_b0 , \133_A[5]_b0 , w_337 );
and ( w_336 , w_337 , \170_B[3]_b0 );
or ( \300_b1 , \298_b1 , \299_b1 );
not ( \299_b1 , w_338 );
and ( \300_b0 , \298_b0 , w_339 );
and ( w_338 , w_339 , \299_b0 );
or ( \301_b1 , \298_b1 , \299_b1 );
xor ( \301_b0 , \298_b0 , w_340 );
not ( w_340 , w_341 );
and ( w_341 , \299_b1 , \299_b0 );
or ( \302_b1 , \245_b1 , \272_b1 );
xor ( \302_b0 , \245_b0 , w_342 );
not ( w_342 , w_343 );
and ( w_343 , \272_b1 , \272_b0 );
or ( \303_b1 , \139_A[4]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_344 );
and ( \303_b0 , \139_A[4]_b0 , w_345 );
and ( w_344 , w_345 , \170_B[3]_b0 );
or ( \304_b1 , \302_b1 , \303_b1 );
not ( \303_b1 , w_346 );
and ( \304_b0 , \302_b0 , w_347 );
and ( w_346 , w_347 , \303_b0 );
or ( \305_b1 , \302_b1 , \303_b1 );
xor ( \305_b0 , \302_b0 , w_348 );
not ( w_348 , w_349 );
and ( w_349 , \303_b1 , \303_b0 );
or ( \306_b1 , \249_b1 , \270_b1 );
xor ( \306_b0 , \249_b0 , w_350 );
not ( w_350 , w_351 );
and ( w_351 , \270_b1 , \270_b0 );
or ( \307_b1 , \145_A[3]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_352 );
and ( \307_b0 , \145_A[3]_b0 , w_353 );
and ( w_352 , w_353 , \170_B[3]_b0 );
or ( \308_b1 , \306_b1 , \307_b1 );
not ( \307_b1 , w_354 );
and ( \308_b0 , \306_b0 , w_355 );
and ( w_354 , w_355 , \307_b0 );
or ( \309_b1 , \306_b1 , \307_b1 );
xor ( \309_b0 , \306_b0 , w_356 );
not ( w_356 , w_357 );
and ( w_357 , \307_b1 , \307_b0 );
or ( \310_b1 , \253_b1 , \268_b1 );
xor ( \310_b0 , \253_b0 , w_358 );
not ( w_358 , w_359 );
and ( w_359 , \268_b1 , \268_b0 );
or ( \311_b1 , \151_A[2]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_360 );
and ( \311_b0 , \151_A[2]_b0 , w_361 );
and ( w_360 , w_361 , \170_B[3]_b0 );
or ( \312_b1 , \310_b1 , \311_b1 );
not ( \311_b1 , w_362 );
and ( \312_b0 , \310_b0 , w_363 );
and ( w_362 , w_363 , \311_b0 );
or ( \313_b1 , \310_b1 , \311_b1 );
xor ( \313_b0 , \310_b0 , w_364 );
not ( w_364 , w_365 );
and ( w_365 , \311_b1 , \311_b0 );
or ( \314_b1 , \257_b1 , \266_b1 );
xor ( \314_b0 , \257_b0 , w_366 );
not ( w_366 , w_367 );
and ( w_367 , \266_b1 , \266_b0 );
or ( \315_b1 , \157_A[1]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_368 );
and ( \315_b0 , \157_A[1]_b0 , w_369 );
and ( w_368 , w_369 , \170_B[3]_b0 );
or ( \316_b1 , \314_b1 , \315_b1 );
not ( \315_b1 , w_370 );
and ( \316_b0 , \314_b0 , w_371 );
and ( w_370 , w_371 , \315_b0 );
or ( \317_b1 , \314_b1 , \315_b1 );
xor ( \317_b0 , \314_b0 , w_372 );
not ( w_372 , w_373 );
and ( w_373 , \315_b1 , \315_b0 );
or ( \318_b1 , \261_b1 , \264_b1 );
xor ( \318_b0 , \261_b0 , w_374 );
not ( w_374 , w_375 );
and ( w_375 , \264_b1 , \264_b0 );
or ( \319_b1 , \163_A[0]_b1 , \170_B[3]_b1 );
not ( \170_B[3]_b1 , w_376 );
and ( \319_b0 , \163_A[0]_b0 , w_377 );
and ( w_376 , w_377 , \170_B[3]_b0 );
or ( \320_b1 , \318_b1 , \319_b1 );
not ( \319_b1 , w_378 );
and ( \320_b0 , \318_b0 , w_379 );
and ( w_378 , w_379 , \319_b0 );
or ( \321_b1 , \317_b1 , \320_b1 );
not ( \320_b1 , w_380 );
and ( \321_b0 , \317_b0 , w_381 );
and ( w_380 , w_381 , \320_b0 );
or ( \322_b1 , \316_b1 , w_382 );
or ( \322_b0 , \316_b0 , \321_b0 );
not ( \321_b0 , w_383 );
and ( w_383 , w_382 , \321_b1 );
or ( \323_b1 , \313_b1 , \322_b1 );
not ( \322_b1 , w_384 );
and ( \323_b0 , \313_b0 , w_385 );
and ( w_384 , w_385 , \322_b0 );
or ( \324_b1 , \312_b1 , w_386 );
or ( \324_b0 , \312_b0 , \323_b0 );
not ( \323_b0 , w_387 );
and ( w_387 , w_386 , \323_b1 );
or ( \325_b1 , \309_b1 , \324_b1 );
not ( \324_b1 , w_388 );
and ( \325_b0 , \309_b0 , w_389 );
and ( w_388 , w_389 , \324_b0 );
or ( \326_b1 , \308_b1 , w_390 );
or ( \326_b0 , \308_b0 , \325_b0 );
not ( \325_b0 , w_391 );
and ( w_391 , w_390 , \325_b1 );
or ( \327_b1 , \305_b1 , \326_b1 );
not ( \326_b1 , w_392 );
and ( \327_b0 , \305_b0 , w_393 );
and ( w_392 , w_393 , \326_b0 );
or ( \328_b1 , \304_b1 , w_394 );
or ( \328_b0 , \304_b0 , \327_b0 );
not ( \327_b0 , w_395 );
and ( w_395 , w_394 , \327_b1 );
or ( \329_b1 , \301_b1 , \328_b1 );
not ( \328_b1 , w_396 );
and ( \329_b0 , \301_b0 , w_397 );
and ( w_396 , w_397 , \328_b0 );
or ( \330_b1 , \300_b1 , w_398 );
or ( \330_b0 , \300_b0 , \329_b0 );
not ( \329_b0 , w_399 );
and ( w_399 , w_398 , \329_b1 );
or ( \331_b1 , \297_b1 , \330_b1 );
not ( \330_b1 , w_400 );
and ( \331_b0 , \297_b0 , w_401 );
and ( w_400 , w_401 , \330_b0 );
or ( \332_b1 , \296_b1 , w_402 );
or ( \332_b0 , \296_b0 , \331_b0 );
not ( \331_b0 , w_403 );
and ( w_403 , w_402 , \331_b1 );
or ( \333_b1 , \293_b1 , \332_b1 );
not ( \332_b1 , w_404 );
and ( \333_b0 , \293_b0 , w_405 );
and ( w_404 , w_405 , \332_b0 );
or ( \334_b1 , \292_b1 , w_406 );
or ( \334_b0 , \292_b0 , \333_b0 );
not ( \333_b0 , w_407 );
and ( w_407 , w_406 , \333_b1 );
or ( \335_b1 , \289_b1 , \334_b1 );
not ( \334_b1 , w_408 );
and ( \335_b0 , \289_b0 , w_409 );
and ( w_408 , w_409 , \334_b0 );
or ( \336_b1 , \288_b1 , w_410 );
or ( \336_b0 , \288_b0 , \335_b0 );
not ( \335_b0 , w_411 );
and ( w_411 , w_410 , \335_b1 );
or ( \337_b1 , \285_b1 , \336_b1 );
not ( \336_b1 , w_412 );
and ( \337_b0 , \285_b0 , w_413 );
and ( w_412 , w_413 , \336_b0 );
or ( \338_b1 , \284_b1 , w_414 );
or ( \338_b0 , \284_b0 , \337_b0 );
not ( \337_b0 , w_415 );
and ( w_415 , w_414 , \337_b1 );
or ( \339_b1 , \109_A[9]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_416 );
and ( \339_b0 , \109_A[9]_b0 , w_417 );
and ( w_416 , w_417 , \169_B[4]_b0 );
or ( \340_b1 , \338_b1 , \339_b1 );
not ( \339_b1 , w_418 );
and ( \340_b0 , \338_b0 , w_419 );
and ( w_418 , w_419 , \339_b0 );
or ( \341_b1 , \338_b1 , \339_b1 );
xor ( \341_b0 , \338_b0 , w_420 );
not ( w_420 , w_421 );
and ( w_421 , \339_b1 , \339_b0 );
or ( \342_b1 , \285_b1 , \336_b1 );
xor ( \342_b0 , \285_b0 , w_422 );
not ( w_422 , w_423 );
and ( w_423 , \336_b1 , \336_b0 );
or ( \343_b1 , \115_A[8]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_424 );
and ( \343_b0 , \115_A[8]_b0 , w_425 );
and ( w_424 , w_425 , \169_B[4]_b0 );
or ( \344_b1 , \342_b1 , \343_b1 );
not ( \343_b1 , w_426 );
and ( \344_b0 , \342_b0 , w_427 );
and ( w_426 , w_427 , \343_b0 );
or ( \345_b1 , \342_b1 , \343_b1 );
xor ( \345_b0 , \342_b0 , w_428 );
not ( w_428 , w_429 );
and ( w_429 , \343_b1 , \343_b0 );
or ( \346_b1 , \289_b1 , \334_b1 );
xor ( \346_b0 , \289_b0 , w_430 );
not ( w_430 , w_431 );
and ( w_431 , \334_b1 , \334_b0 );
or ( \347_b1 , \121_A[7]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_432 );
and ( \347_b0 , \121_A[7]_b0 , w_433 );
and ( w_432 , w_433 , \169_B[4]_b0 );
or ( \348_b1 , \346_b1 , \347_b1 );
not ( \347_b1 , w_434 );
and ( \348_b0 , \346_b0 , w_435 );
and ( w_434 , w_435 , \347_b0 );
or ( \349_b1 , \346_b1 , \347_b1 );
xor ( \349_b0 , \346_b0 , w_436 );
not ( w_436 , w_437 );
and ( w_437 , \347_b1 , \347_b0 );
or ( \350_b1 , \293_b1 , \332_b1 );
xor ( \350_b0 , \293_b0 , w_438 );
not ( w_438 , w_439 );
and ( w_439 , \332_b1 , \332_b0 );
or ( \351_b1 , \127_A[6]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_440 );
and ( \351_b0 , \127_A[6]_b0 , w_441 );
and ( w_440 , w_441 , \169_B[4]_b0 );
or ( \352_b1 , \350_b1 , \351_b1 );
not ( \351_b1 , w_442 );
and ( \352_b0 , \350_b0 , w_443 );
and ( w_442 , w_443 , \351_b0 );
or ( \353_b1 , \350_b1 , \351_b1 );
xor ( \353_b0 , \350_b0 , w_444 );
not ( w_444 , w_445 );
and ( w_445 , \351_b1 , \351_b0 );
or ( \354_b1 , \297_b1 , \330_b1 );
xor ( \354_b0 , \297_b0 , w_446 );
not ( w_446 , w_447 );
and ( w_447 , \330_b1 , \330_b0 );
or ( \355_b1 , \133_A[5]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_448 );
and ( \355_b0 , \133_A[5]_b0 , w_449 );
and ( w_448 , w_449 , \169_B[4]_b0 );
or ( \356_b1 , \354_b1 , \355_b1 );
not ( \355_b1 , w_450 );
and ( \356_b0 , \354_b0 , w_451 );
and ( w_450 , w_451 , \355_b0 );
or ( \357_b1 , \354_b1 , \355_b1 );
xor ( \357_b0 , \354_b0 , w_452 );
not ( w_452 , w_453 );
and ( w_453 , \355_b1 , \355_b0 );
or ( \358_b1 , \301_b1 , \328_b1 );
xor ( \358_b0 , \301_b0 , w_454 );
not ( w_454 , w_455 );
and ( w_455 , \328_b1 , \328_b0 );
or ( \359_b1 , \139_A[4]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_456 );
and ( \359_b0 , \139_A[4]_b0 , w_457 );
and ( w_456 , w_457 , \169_B[4]_b0 );
or ( \360_b1 , \358_b1 , \359_b1 );
not ( \359_b1 , w_458 );
and ( \360_b0 , \358_b0 , w_459 );
and ( w_458 , w_459 , \359_b0 );
or ( \361_b1 , \358_b1 , \359_b1 );
xor ( \361_b0 , \358_b0 , w_460 );
not ( w_460 , w_461 );
and ( w_461 , \359_b1 , \359_b0 );
or ( \362_b1 , \305_b1 , \326_b1 );
xor ( \362_b0 , \305_b0 , w_462 );
not ( w_462 , w_463 );
and ( w_463 , \326_b1 , \326_b0 );
or ( \363_b1 , \145_A[3]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_464 );
and ( \363_b0 , \145_A[3]_b0 , w_465 );
and ( w_464 , w_465 , \169_B[4]_b0 );
or ( \364_b1 , \362_b1 , \363_b1 );
not ( \363_b1 , w_466 );
and ( \364_b0 , \362_b0 , w_467 );
and ( w_466 , w_467 , \363_b0 );
or ( \365_b1 , \362_b1 , \363_b1 );
xor ( \365_b0 , \362_b0 , w_468 );
not ( w_468 , w_469 );
and ( w_469 , \363_b1 , \363_b0 );
or ( \366_b1 , \309_b1 , \324_b1 );
xor ( \366_b0 , \309_b0 , w_470 );
not ( w_470 , w_471 );
and ( w_471 , \324_b1 , \324_b0 );
or ( \367_b1 , \151_A[2]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_472 );
and ( \367_b0 , \151_A[2]_b0 , w_473 );
and ( w_472 , w_473 , \169_B[4]_b0 );
or ( \368_b1 , \366_b1 , \367_b1 );
not ( \367_b1 , w_474 );
and ( \368_b0 , \366_b0 , w_475 );
and ( w_474 , w_475 , \367_b0 );
or ( \369_b1 , \366_b1 , \367_b1 );
xor ( \369_b0 , \366_b0 , w_476 );
not ( w_476 , w_477 );
and ( w_477 , \367_b1 , \367_b0 );
or ( \370_b1 , \313_b1 , \322_b1 );
xor ( \370_b0 , \313_b0 , w_478 );
not ( w_478 , w_479 );
and ( w_479 , \322_b1 , \322_b0 );
or ( \371_b1 , \157_A[1]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_480 );
and ( \371_b0 , \157_A[1]_b0 , w_481 );
and ( w_480 , w_481 , \169_B[4]_b0 );
or ( \372_b1 , \370_b1 , \371_b1 );
not ( \371_b1 , w_482 );
and ( \372_b0 , \370_b0 , w_483 );
and ( w_482 , w_483 , \371_b0 );
or ( \373_b1 , \370_b1 , \371_b1 );
xor ( \373_b0 , \370_b0 , w_484 );
not ( w_484 , w_485 );
and ( w_485 , \371_b1 , \371_b0 );
or ( \374_b1 , \317_b1 , \320_b1 );
xor ( \374_b0 , \317_b0 , w_486 );
not ( w_486 , w_487 );
and ( w_487 , \320_b1 , \320_b0 );
or ( \375_b1 , \163_A[0]_b1 , \169_B[4]_b1 );
not ( \169_B[4]_b1 , w_488 );
and ( \375_b0 , \163_A[0]_b0 , w_489 );
and ( w_488 , w_489 , \169_B[4]_b0 );
or ( \376_b1 , \374_b1 , \375_b1 );
not ( \375_b1 , w_490 );
and ( \376_b0 , \374_b0 , w_491 );
and ( w_490 , w_491 , \375_b0 );
or ( \377_b1 , \373_b1 , \376_b1 );
not ( \376_b1 , w_492 );
and ( \377_b0 , \373_b0 , w_493 );
and ( w_492 , w_493 , \376_b0 );
or ( \378_b1 , \372_b1 , w_494 );
or ( \378_b0 , \372_b0 , \377_b0 );
not ( \377_b0 , w_495 );
and ( w_495 , w_494 , \377_b1 );
or ( \379_b1 , \369_b1 , \378_b1 );
not ( \378_b1 , w_496 );
and ( \379_b0 , \369_b0 , w_497 );
and ( w_496 , w_497 , \378_b0 );
or ( \380_b1 , \368_b1 , w_498 );
or ( \380_b0 , \368_b0 , \379_b0 );
not ( \379_b0 , w_499 );
and ( w_499 , w_498 , \379_b1 );
or ( \381_b1 , \365_b1 , \380_b1 );
not ( \380_b1 , w_500 );
and ( \381_b0 , \365_b0 , w_501 );
and ( w_500 , w_501 , \380_b0 );
or ( \382_b1 , \364_b1 , w_502 );
or ( \382_b0 , \364_b0 , \381_b0 );
not ( \381_b0 , w_503 );
and ( w_503 , w_502 , \381_b1 );
or ( \383_b1 , \361_b1 , \382_b1 );
not ( \382_b1 , w_504 );
and ( \383_b0 , \361_b0 , w_505 );
and ( w_504 , w_505 , \382_b0 );
or ( \384_b1 , \360_b1 , w_506 );
or ( \384_b0 , \360_b0 , \383_b0 );
not ( \383_b0 , w_507 );
and ( w_507 , w_506 , \383_b1 );
or ( \385_b1 , \357_b1 , \384_b1 );
not ( \384_b1 , w_508 );
and ( \385_b0 , \357_b0 , w_509 );
and ( w_508 , w_509 , \384_b0 );
or ( \386_b1 , \356_b1 , w_510 );
or ( \386_b0 , \356_b0 , \385_b0 );
not ( \385_b0 , w_511 );
and ( w_511 , w_510 , \385_b1 );
or ( \387_b1 , \353_b1 , \386_b1 );
not ( \386_b1 , w_512 );
and ( \387_b0 , \353_b0 , w_513 );
and ( w_512 , w_513 , \386_b0 );
or ( \388_b1 , \352_b1 , w_514 );
or ( \388_b0 , \352_b0 , \387_b0 );
not ( \387_b0 , w_515 );
and ( w_515 , w_514 , \387_b1 );
or ( \389_b1 , \349_b1 , \388_b1 );
not ( \388_b1 , w_516 );
and ( \389_b0 , \349_b0 , w_517 );
and ( w_516 , w_517 , \388_b0 );
or ( \390_b1 , \348_b1 , w_518 );
or ( \390_b0 , \348_b0 , \389_b0 );
not ( \389_b0 , w_519 );
and ( w_519 , w_518 , \389_b1 );
or ( \391_b1 , \345_b1 , \390_b1 );
not ( \390_b1 , w_520 );
and ( \391_b0 , \345_b0 , w_521 );
and ( w_520 , w_521 , \390_b0 );
or ( \392_b1 , \344_b1 , w_522 );
or ( \392_b0 , \344_b0 , \391_b0 );
not ( \391_b0 , w_523 );
and ( w_523 , w_522 , \391_b1 );
or ( \393_b1 , \341_b1 , \392_b1 );
not ( \392_b1 , w_524 );
and ( \393_b0 , \341_b0 , w_525 );
and ( w_524 , w_525 , \392_b0 );
or ( \394_b1 , \340_b1 , w_526 );
or ( \394_b0 , \340_b0 , \393_b0 );
not ( \393_b0 , w_527 );
and ( w_527 , w_526 , \393_b1 );
or ( \395_b1 , \109_A[9]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_528 );
and ( \395_b0 , \109_A[9]_b0 , w_529 );
and ( w_528 , w_529 , \168_B[5]_b0 );
or ( \396_b1 , \394_b1 , \395_b1 );
not ( \395_b1 , w_530 );
and ( \396_b0 , \394_b0 , w_531 );
and ( w_530 , w_531 , \395_b0 );
or ( \397_b1 , \394_b1 , \395_b1 );
xor ( \397_b0 , \394_b0 , w_532 );
not ( w_532 , w_533 );
and ( w_533 , \395_b1 , \395_b0 );
or ( \398_b1 , \341_b1 , \392_b1 );
xor ( \398_b0 , \341_b0 , w_534 );
not ( w_534 , w_535 );
and ( w_535 , \392_b1 , \392_b0 );
or ( \399_b1 , \115_A[8]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_536 );
and ( \399_b0 , \115_A[8]_b0 , w_537 );
and ( w_536 , w_537 , \168_B[5]_b0 );
or ( \400_b1 , \398_b1 , \399_b1 );
not ( \399_b1 , w_538 );
and ( \400_b0 , \398_b0 , w_539 );
and ( w_538 , w_539 , \399_b0 );
or ( \401_b1 , \398_b1 , \399_b1 );
xor ( \401_b0 , \398_b0 , w_540 );
not ( w_540 , w_541 );
and ( w_541 , \399_b1 , \399_b0 );
or ( \402_b1 , \345_b1 , \390_b1 );
xor ( \402_b0 , \345_b0 , w_542 );
not ( w_542 , w_543 );
and ( w_543 , \390_b1 , \390_b0 );
or ( \403_b1 , \121_A[7]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_544 );
and ( \403_b0 , \121_A[7]_b0 , w_545 );
and ( w_544 , w_545 , \168_B[5]_b0 );
or ( \404_b1 , \402_b1 , \403_b1 );
not ( \403_b1 , w_546 );
and ( \404_b0 , \402_b0 , w_547 );
and ( w_546 , w_547 , \403_b0 );
or ( \405_b1 , \402_b1 , \403_b1 );
xor ( \405_b0 , \402_b0 , w_548 );
not ( w_548 , w_549 );
and ( w_549 , \403_b1 , \403_b0 );
or ( \406_b1 , \349_b1 , \388_b1 );
xor ( \406_b0 , \349_b0 , w_550 );
not ( w_550 , w_551 );
and ( w_551 , \388_b1 , \388_b0 );
or ( \407_b1 , \127_A[6]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_552 );
and ( \407_b0 , \127_A[6]_b0 , w_553 );
and ( w_552 , w_553 , \168_B[5]_b0 );
or ( \408_b1 , \406_b1 , \407_b1 );
not ( \407_b1 , w_554 );
and ( \408_b0 , \406_b0 , w_555 );
and ( w_554 , w_555 , \407_b0 );
or ( \409_b1 , \406_b1 , \407_b1 );
xor ( \409_b0 , \406_b0 , w_556 );
not ( w_556 , w_557 );
and ( w_557 , \407_b1 , \407_b0 );
or ( \410_b1 , \353_b1 , \386_b1 );
xor ( \410_b0 , \353_b0 , w_558 );
not ( w_558 , w_559 );
and ( w_559 , \386_b1 , \386_b0 );
or ( \411_b1 , \133_A[5]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_560 );
and ( \411_b0 , \133_A[5]_b0 , w_561 );
and ( w_560 , w_561 , \168_B[5]_b0 );
or ( \412_b1 , \410_b1 , \411_b1 );
not ( \411_b1 , w_562 );
and ( \412_b0 , \410_b0 , w_563 );
and ( w_562 , w_563 , \411_b0 );
or ( \413_b1 , \410_b1 , \411_b1 );
xor ( \413_b0 , \410_b0 , w_564 );
not ( w_564 , w_565 );
and ( w_565 , \411_b1 , \411_b0 );
or ( \414_b1 , \357_b1 , \384_b1 );
xor ( \414_b0 , \357_b0 , w_566 );
not ( w_566 , w_567 );
and ( w_567 , \384_b1 , \384_b0 );
or ( \415_b1 , \139_A[4]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_568 );
and ( \415_b0 , \139_A[4]_b0 , w_569 );
and ( w_568 , w_569 , \168_B[5]_b0 );
or ( \416_b1 , \414_b1 , \415_b1 );
not ( \415_b1 , w_570 );
and ( \416_b0 , \414_b0 , w_571 );
and ( w_570 , w_571 , \415_b0 );
or ( \417_b1 , \414_b1 , \415_b1 );
xor ( \417_b0 , \414_b0 , w_572 );
not ( w_572 , w_573 );
and ( w_573 , \415_b1 , \415_b0 );
or ( \418_b1 , \361_b1 , \382_b1 );
xor ( \418_b0 , \361_b0 , w_574 );
not ( w_574 , w_575 );
and ( w_575 , \382_b1 , \382_b0 );
or ( \419_b1 , \145_A[3]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_576 );
and ( \419_b0 , \145_A[3]_b0 , w_577 );
and ( w_576 , w_577 , \168_B[5]_b0 );
or ( \420_b1 , \418_b1 , \419_b1 );
not ( \419_b1 , w_578 );
and ( \420_b0 , \418_b0 , w_579 );
and ( w_578 , w_579 , \419_b0 );
or ( \421_b1 , \418_b1 , \419_b1 );
xor ( \421_b0 , \418_b0 , w_580 );
not ( w_580 , w_581 );
and ( w_581 , \419_b1 , \419_b0 );
or ( \422_b1 , \365_b1 , \380_b1 );
xor ( \422_b0 , \365_b0 , w_582 );
not ( w_582 , w_583 );
and ( w_583 , \380_b1 , \380_b0 );
or ( \423_b1 , \151_A[2]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_584 );
and ( \423_b0 , \151_A[2]_b0 , w_585 );
and ( w_584 , w_585 , \168_B[5]_b0 );
or ( \424_b1 , \422_b1 , \423_b1 );
not ( \423_b1 , w_586 );
and ( \424_b0 , \422_b0 , w_587 );
and ( w_586 , w_587 , \423_b0 );
or ( \425_b1 , \422_b1 , \423_b1 );
xor ( \425_b0 , \422_b0 , w_588 );
not ( w_588 , w_589 );
and ( w_589 , \423_b1 , \423_b0 );
or ( \426_b1 , \369_b1 , \378_b1 );
xor ( \426_b0 , \369_b0 , w_590 );
not ( w_590 , w_591 );
and ( w_591 , \378_b1 , \378_b0 );
or ( \427_b1 , \157_A[1]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_592 );
and ( \427_b0 , \157_A[1]_b0 , w_593 );
and ( w_592 , w_593 , \168_B[5]_b0 );
or ( \428_b1 , \426_b1 , \427_b1 );
not ( \427_b1 , w_594 );
and ( \428_b0 , \426_b0 , w_595 );
and ( w_594 , w_595 , \427_b0 );
or ( \429_b1 , \426_b1 , \427_b1 );
xor ( \429_b0 , \426_b0 , w_596 );
not ( w_596 , w_597 );
and ( w_597 , \427_b1 , \427_b0 );
or ( \430_b1 , \373_b1 , \376_b1 );
xor ( \430_b0 , \373_b0 , w_598 );
not ( w_598 , w_599 );
and ( w_599 , \376_b1 , \376_b0 );
or ( \431_b1 , \163_A[0]_b1 , \168_B[5]_b1 );
not ( \168_B[5]_b1 , w_600 );
and ( \431_b0 , \163_A[0]_b0 , w_601 );
and ( w_600 , w_601 , \168_B[5]_b0 );
or ( \432_b1 , \430_b1 , \431_b1 );
not ( \431_b1 , w_602 );
and ( \432_b0 , \430_b0 , w_603 );
and ( w_602 , w_603 , \431_b0 );
or ( \433_b1 , \429_b1 , \432_b1 );
not ( \432_b1 , w_604 );
and ( \433_b0 , \429_b0 , w_605 );
and ( w_604 , w_605 , \432_b0 );
or ( \434_b1 , \428_b1 , w_606 );
or ( \434_b0 , \428_b0 , \433_b0 );
not ( \433_b0 , w_607 );
and ( w_607 , w_606 , \433_b1 );
or ( \435_b1 , \425_b1 , \434_b1 );
not ( \434_b1 , w_608 );
and ( \435_b0 , \425_b0 , w_609 );
and ( w_608 , w_609 , \434_b0 );
or ( \436_b1 , \424_b1 , w_610 );
or ( \436_b0 , \424_b0 , \435_b0 );
not ( \435_b0 , w_611 );
and ( w_611 , w_610 , \435_b1 );
or ( \437_b1 , \421_b1 , \436_b1 );
not ( \436_b1 , w_612 );
and ( \437_b0 , \421_b0 , w_613 );
and ( w_612 , w_613 , \436_b0 );
or ( \438_b1 , \420_b1 , w_614 );
or ( \438_b0 , \420_b0 , \437_b0 );
not ( \437_b0 , w_615 );
and ( w_615 , w_614 , \437_b1 );
or ( \439_b1 , \417_b1 , \438_b1 );
not ( \438_b1 , w_616 );
and ( \439_b0 , \417_b0 , w_617 );
and ( w_616 , w_617 , \438_b0 );
or ( \440_b1 , \416_b1 , w_618 );
or ( \440_b0 , \416_b0 , \439_b0 );
not ( \439_b0 , w_619 );
and ( w_619 , w_618 , \439_b1 );
or ( \441_b1 , \413_b1 , \440_b1 );
not ( \440_b1 , w_620 );
and ( \441_b0 , \413_b0 , w_621 );
and ( w_620 , w_621 , \440_b0 );
or ( \442_b1 , \412_b1 , w_622 );
or ( \442_b0 , \412_b0 , \441_b0 );
not ( \441_b0 , w_623 );
and ( w_623 , w_622 , \441_b1 );
or ( \443_b1 , \409_b1 , \442_b1 );
not ( \442_b1 , w_624 );
and ( \443_b0 , \409_b0 , w_625 );
and ( w_624 , w_625 , \442_b0 );
or ( \444_b1 , \408_b1 , w_626 );
or ( \444_b0 , \408_b0 , \443_b0 );
not ( \443_b0 , w_627 );
and ( w_627 , w_626 , \443_b1 );
or ( \445_b1 , \405_b1 , \444_b1 );
not ( \444_b1 , w_628 );
and ( \445_b0 , \405_b0 , w_629 );
and ( w_628 , w_629 , \444_b0 );
or ( \446_b1 , \404_b1 , w_630 );
or ( \446_b0 , \404_b0 , \445_b0 );
not ( \445_b0 , w_631 );
and ( w_631 , w_630 , \445_b1 );
or ( \447_b1 , \401_b1 , \446_b1 );
not ( \446_b1 , w_632 );
and ( \447_b0 , \401_b0 , w_633 );
and ( w_632 , w_633 , \446_b0 );
or ( \448_b1 , \400_b1 , w_634 );
or ( \448_b0 , \400_b0 , \447_b0 );
not ( \447_b0 , w_635 );
and ( w_635 , w_634 , \447_b1 );
or ( \449_b1 , \397_b1 , \448_b1 );
not ( \448_b1 , w_636 );
and ( \449_b0 , \397_b0 , w_637 );
and ( w_636 , w_637 , \448_b0 );
or ( \450_b1 , \396_b1 , w_638 );
or ( \450_b0 , \396_b0 , \449_b0 );
not ( \449_b0 , w_639 );
and ( w_639 , w_638 , \449_b1 );
or ( \451_b1 , \109_A[9]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_640 );
and ( \451_b0 , \109_A[9]_b0 , w_641 );
and ( w_640 , w_641 , \167_B[6]_b0 );
or ( \452_b1 , \450_b1 , \451_b1 );
not ( \451_b1 , w_642 );
and ( \452_b0 , \450_b0 , w_643 );
and ( w_642 , w_643 , \451_b0 );
or ( \453_b1 , \450_b1 , \451_b1 );
xor ( \453_b0 , \450_b0 , w_644 );
not ( w_644 , w_645 );
and ( w_645 , \451_b1 , \451_b0 );
or ( \454_b1 , \397_b1 , \448_b1 );
xor ( \454_b0 , \397_b0 , w_646 );
not ( w_646 , w_647 );
and ( w_647 , \448_b1 , \448_b0 );
or ( \455_b1 , \115_A[8]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_648 );
and ( \455_b0 , \115_A[8]_b0 , w_649 );
and ( w_648 , w_649 , \167_B[6]_b0 );
or ( \456_b1 , \454_b1 , \455_b1 );
not ( \455_b1 , w_650 );
and ( \456_b0 , \454_b0 , w_651 );
and ( w_650 , w_651 , \455_b0 );
or ( \457_b1 , \454_b1 , \455_b1 );
xor ( \457_b0 , \454_b0 , w_652 );
not ( w_652 , w_653 );
and ( w_653 , \455_b1 , \455_b0 );
or ( \458_b1 , \401_b1 , \446_b1 );
xor ( \458_b0 , \401_b0 , w_654 );
not ( w_654 , w_655 );
and ( w_655 , \446_b1 , \446_b0 );
or ( \459_b1 , \121_A[7]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_656 );
and ( \459_b0 , \121_A[7]_b0 , w_657 );
and ( w_656 , w_657 , \167_B[6]_b0 );
or ( \460_b1 , \458_b1 , \459_b1 );
not ( \459_b1 , w_658 );
and ( \460_b0 , \458_b0 , w_659 );
and ( w_658 , w_659 , \459_b0 );
or ( \461_b1 , \458_b1 , \459_b1 );
xor ( \461_b0 , \458_b0 , w_660 );
not ( w_660 , w_661 );
and ( w_661 , \459_b1 , \459_b0 );
or ( \462_b1 , \405_b1 , \444_b1 );
xor ( \462_b0 , \405_b0 , w_662 );
not ( w_662 , w_663 );
and ( w_663 , \444_b1 , \444_b0 );
or ( \463_b1 , \127_A[6]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_664 );
and ( \463_b0 , \127_A[6]_b0 , w_665 );
and ( w_664 , w_665 , \167_B[6]_b0 );
or ( \464_b1 , \462_b1 , \463_b1 );
not ( \463_b1 , w_666 );
and ( \464_b0 , \462_b0 , w_667 );
and ( w_666 , w_667 , \463_b0 );
or ( \465_b1 , \462_b1 , \463_b1 );
xor ( \465_b0 , \462_b0 , w_668 );
not ( w_668 , w_669 );
and ( w_669 , \463_b1 , \463_b0 );
or ( \466_b1 , \409_b1 , \442_b1 );
xor ( \466_b0 , \409_b0 , w_670 );
not ( w_670 , w_671 );
and ( w_671 , \442_b1 , \442_b0 );
or ( \467_b1 , \133_A[5]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_672 );
and ( \467_b0 , \133_A[5]_b0 , w_673 );
and ( w_672 , w_673 , \167_B[6]_b0 );
or ( \468_b1 , \466_b1 , \467_b1 );
not ( \467_b1 , w_674 );
and ( \468_b0 , \466_b0 , w_675 );
and ( w_674 , w_675 , \467_b0 );
or ( \469_b1 , \466_b1 , \467_b1 );
xor ( \469_b0 , \466_b0 , w_676 );
not ( w_676 , w_677 );
and ( w_677 , \467_b1 , \467_b0 );
or ( \470_b1 , \413_b1 , \440_b1 );
xor ( \470_b0 , \413_b0 , w_678 );
not ( w_678 , w_679 );
and ( w_679 , \440_b1 , \440_b0 );
or ( \471_b1 , \139_A[4]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_680 );
and ( \471_b0 , \139_A[4]_b0 , w_681 );
and ( w_680 , w_681 , \167_B[6]_b0 );
or ( \472_b1 , \470_b1 , \471_b1 );
not ( \471_b1 , w_682 );
and ( \472_b0 , \470_b0 , w_683 );
and ( w_682 , w_683 , \471_b0 );
or ( \473_b1 , \470_b1 , \471_b1 );
xor ( \473_b0 , \470_b0 , w_684 );
not ( w_684 , w_685 );
and ( w_685 , \471_b1 , \471_b0 );
or ( \474_b1 , \417_b1 , \438_b1 );
xor ( \474_b0 , \417_b0 , w_686 );
not ( w_686 , w_687 );
and ( w_687 , \438_b1 , \438_b0 );
or ( \475_b1 , \145_A[3]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_688 );
and ( \475_b0 , \145_A[3]_b0 , w_689 );
and ( w_688 , w_689 , \167_B[6]_b0 );
or ( \476_b1 , \474_b1 , \475_b1 );
not ( \475_b1 , w_690 );
and ( \476_b0 , \474_b0 , w_691 );
and ( w_690 , w_691 , \475_b0 );
or ( \477_b1 , \474_b1 , \475_b1 );
xor ( \477_b0 , \474_b0 , w_692 );
not ( w_692 , w_693 );
and ( w_693 , \475_b1 , \475_b0 );
or ( \478_b1 , \421_b1 , \436_b1 );
xor ( \478_b0 , \421_b0 , w_694 );
not ( w_694 , w_695 );
and ( w_695 , \436_b1 , \436_b0 );
or ( \479_b1 , \151_A[2]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_696 );
and ( \479_b0 , \151_A[2]_b0 , w_697 );
and ( w_696 , w_697 , \167_B[6]_b0 );
or ( \480_b1 , \478_b1 , \479_b1 );
not ( \479_b1 , w_698 );
and ( \480_b0 , \478_b0 , w_699 );
and ( w_698 , w_699 , \479_b0 );
or ( \481_b1 , \478_b1 , \479_b1 );
xor ( \481_b0 , \478_b0 , w_700 );
not ( w_700 , w_701 );
and ( w_701 , \479_b1 , \479_b0 );
or ( \482_b1 , \425_b1 , \434_b1 );
xor ( \482_b0 , \425_b0 , w_702 );
not ( w_702 , w_703 );
and ( w_703 , \434_b1 , \434_b0 );
or ( \483_b1 , \157_A[1]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_704 );
and ( \483_b0 , \157_A[1]_b0 , w_705 );
and ( w_704 , w_705 , \167_B[6]_b0 );
or ( \484_b1 , \482_b1 , \483_b1 );
not ( \483_b1 , w_706 );
and ( \484_b0 , \482_b0 , w_707 );
and ( w_706 , w_707 , \483_b0 );
or ( \485_b1 , \482_b1 , \483_b1 );
xor ( \485_b0 , \482_b0 , w_708 );
not ( w_708 , w_709 );
and ( w_709 , \483_b1 , \483_b0 );
or ( \486_b1 , \429_b1 , \432_b1 );
xor ( \486_b0 , \429_b0 , w_710 );
not ( w_710 , w_711 );
and ( w_711 , \432_b1 , \432_b0 );
or ( \487_b1 , \163_A[0]_b1 , \167_B[6]_b1 );
not ( \167_B[6]_b1 , w_712 );
and ( \487_b0 , \163_A[0]_b0 , w_713 );
and ( w_712 , w_713 , \167_B[6]_b0 );
or ( \488_b1 , \486_b1 , \487_b1 );
not ( \487_b1 , w_714 );
and ( \488_b0 , \486_b0 , w_715 );
and ( w_714 , w_715 , \487_b0 );
or ( \489_b1 , \485_b1 , \488_b1 );
not ( \488_b1 , w_716 );
and ( \489_b0 , \485_b0 , w_717 );
and ( w_716 , w_717 , \488_b0 );
or ( \490_b1 , \484_b1 , w_718 );
or ( \490_b0 , \484_b0 , \489_b0 );
not ( \489_b0 , w_719 );
and ( w_719 , w_718 , \489_b1 );
or ( \491_b1 , \481_b1 , \490_b1 );
not ( \490_b1 , w_720 );
and ( \491_b0 , \481_b0 , w_721 );
and ( w_720 , w_721 , \490_b0 );
or ( \492_b1 , \480_b1 , w_722 );
or ( \492_b0 , \480_b0 , \491_b0 );
not ( \491_b0 , w_723 );
and ( w_723 , w_722 , \491_b1 );
or ( \493_b1 , \477_b1 , \492_b1 );
not ( \492_b1 , w_724 );
and ( \493_b0 , \477_b0 , w_725 );
and ( w_724 , w_725 , \492_b0 );
or ( \494_b1 , \476_b1 , w_726 );
or ( \494_b0 , \476_b0 , \493_b0 );
not ( \493_b0 , w_727 );
and ( w_727 , w_726 , \493_b1 );
or ( \495_b1 , \473_b1 , \494_b1 );
not ( \494_b1 , w_728 );
and ( \495_b0 , \473_b0 , w_729 );
and ( w_728 , w_729 , \494_b0 );
or ( \496_b1 , \472_b1 , w_730 );
or ( \496_b0 , \472_b0 , \495_b0 );
not ( \495_b0 , w_731 );
and ( w_731 , w_730 , \495_b1 );
or ( \497_b1 , \469_b1 , \496_b1 );
not ( \496_b1 , w_732 );
and ( \497_b0 , \469_b0 , w_733 );
and ( w_732 , w_733 , \496_b0 );
or ( \498_b1 , \468_b1 , w_734 );
or ( \498_b0 , \468_b0 , \497_b0 );
not ( \497_b0 , w_735 );
and ( w_735 , w_734 , \497_b1 );
or ( \499_b1 , \465_b1 , \498_b1 );
not ( \498_b1 , w_736 );
and ( \499_b0 , \465_b0 , w_737 );
and ( w_736 , w_737 , \498_b0 );
or ( \500_b1 , \464_b1 , w_738 );
or ( \500_b0 , \464_b0 , \499_b0 );
not ( \499_b0 , w_739 );
and ( w_739 , w_738 , \499_b1 );
or ( \501_b1 , \461_b1 , \500_b1 );
not ( \500_b1 , w_740 );
and ( \501_b0 , \461_b0 , w_741 );
and ( w_740 , w_741 , \500_b0 );
or ( \502_b1 , \460_b1 , w_742 );
or ( \502_b0 , \460_b0 , \501_b0 );
not ( \501_b0 , w_743 );
and ( w_743 , w_742 , \501_b1 );
or ( \503_b1 , \457_b1 , \502_b1 );
not ( \502_b1 , w_744 );
and ( \503_b0 , \457_b0 , w_745 );
and ( w_744 , w_745 , \502_b0 );
or ( \504_b1 , \456_b1 , w_746 );
or ( \504_b0 , \456_b0 , \503_b0 );
not ( \503_b0 , w_747 );
and ( w_747 , w_746 , \503_b1 );
or ( \505_b1 , \453_b1 , \504_b1 );
not ( \504_b1 , w_748 );
and ( \505_b0 , \453_b0 , w_749 );
and ( w_748 , w_749 , \504_b0 );
or ( \506_b1 , \452_b1 , w_750 );
or ( \506_b0 , \452_b0 , \505_b0 );
not ( \505_b0 , w_751 );
and ( w_751 , w_750 , \505_b1 );
or ( \507_b1 , \109_A[9]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_752 );
and ( \507_b0 , \109_A[9]_b0 , w_753 );
and ( w_752 , w_753 , \166_B[7]_b0 );
or ( \508_b1 , \506_b1 , \507_b1 );
not ( \507_b1 , w_754 );
and ( \508_b0 , \506_b0 , w_755 );
and ( w_754 , w_755 , \507_b0 );
or ( \509_b1 , \506_b1 , \507_b1 );
xor ( \509_b0 , \506_b0 , w_756 );
not ( w_756 , w_757 );
and ( w_757 , \507_b1 , \507_b0 );
or ( \510_b1 , \453_b1 , \504_b1 );
xor ( \510_b0 , \453_b0 , w_758 );
not ( w_758 , w_759 );
and ( w_759 , \504_b1 , \504_b0 );
or ( \511_b1 , \115_A[8]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_760 );
and ( \511_b0 , \115_A[8]_b0 , w_761 );
and ( w_760 , w_761 , \166_B[7]_b0 );
or ( \512_b1 , \510_b1 , \511_b1 );
not ( \511_b1 , w_762 );
and ( \512_b0 , \510_b0 , w_763 );
and ( w_762 , w_763 , \511_b0 );
or ( \513_b1 , \510_b1 , \511_b1 );
xor ( \513_b0 , \510_b0 , w_764 );
not ( w_764 , w_765 );
and ( w_765 , \511_b1 , \511_b0 );
or ( \514_b1 , \457_b1 , \502_b1 );
xor ( \514_b0 , \457_b0 , w_766 );
not ( w_766 , w_767 );
and ( w_767 , \502_b1 , \502_b0 );
or ( \515_b1 , \121_A[7]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_768 );
and ( \515_b0 , \121_A[7]_b0 , w_769 );
and ( w_768 , w_769 , \166_B[7]_b0 );
or ( \516_b1 , \514_b1 , \515_b1 );
not ( \515_b1 , w_770 );
and ( \516_b0 , \514_b0 , w_771 );
and ( w_770 , w_771 , \515_b0 );
or ( \517_b1 , \514_b1 , \515_b1 );
xor ( \517_b0 , \514_b0 , w_772 );
not ( w_772 , w_773 );
and ( w_773 , \515_b1 , \515_b0 );
or ( \518_b1 , \461_b1 , \500_b1 );
xor ( \518_b0 , \461_b0 , w_774 );
not ( w_774 , w_775 );
and ( w_775 , \500_b1 , \500_b0 );
or ( \519_b1 , \127_A[6]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_776 );
and ( \519_b0 , \127_A[6]_b0 , w_777 );
and ( w_776 , w_777 , \166_B[7]_b0 );
or ( \520_b1 , \518_b1 , \519_b1 );
not ( \519_b1 , w_778 );
and ( \520_b0 , \518_b0 , w_779 );
and ( w_778 , w_779 , \519_b0 );
or ( \521_b1 , \518_b1 , \519_b1 );
xor ( \521_b0 , \518_b0 , w_780 );
not ( w_780 , w_781 );
and ( w_781 , \519_b1 , \519_b0 );
or ( \522_b1 , \465_b1 , \498_b1 );
xor ( \522_b0 , \465_b0 , w_782 );
not ( w_782 , w_783 );
and ( w_783 , \498_b1 , \498_b0 );
or ( \523_b1 , \133_A[5]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_784 );
and ( \523_b0 , \133_A[5]_b0 , w_785 );
and ( w_784 , w_785 , \166_B[7]_b0 );
or ( \524_b1 , \522_b1 , \523_b1 );
not ( \523_b1 , w_786 );
and ( \524_b0 , \522_b0 , w_787 );
and ( w_786 , w_787 , \523_b0 );
or ( \525_b1 , \522_b1 , \523_b1 );
xor ( \525_b0 , \522_b0 , w_788 );
not ( w_788 , w_789 );
and ( w_789 , \523_b1 , \523_b0 );
or ( \526_b1 , \469_b1 , \496_b1 );
xor ( \526_b0 , \469_b0 , w_790 );
not ( w_790 , w_791 );
and ( w_791 , \496_b1 , \496_b0 );
or ( \527_b1 , \139_A[4]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_792 );
and ( \527_b0 , \139_A[4]_b0 , w_793 );
and ( w_792 , w_793 , \166_B[7]_b0 );
or ( \528_b1 , \526_b1 , \527_b1 );
not ( \527_b1 , w_794 );
and ( \528_b0 , \526_b0 , w_795 );
and ( w_794 , w_795 , \527_b0 );
or ( \529_b1 , \526_b1 , \527_b1 );
xor ( \529_b0 , \526_b0 , w_796 );
not ( w_796 , w_797 );
and ( w_797 , \527_b1 , \527_b0 );
or ( \530_b1 , \473_b1 , \494_b1 );
xor ( \530_b0 , \473_b0 , w_798 );
not ( w_798 , w_799 );
and ( w_799 , \494_b1 , \494_b0 );
or ( \531_b1 , \145_A[3]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_800 );
and ( \531_b0 , \145_A[3]_b0 , w_801 );
and ( w_800 , w_801 , \166_B[7]_b0 );
or ( \532_b1 , \530_b1 , \531_b1 );
not ( \531_b1 , w_802 );
and ( \532_b0 , \530_b0 , w_803 );
and ( w_802 , w_803 , \531_b0 );
or ( \533_b1 , \530_b1 , \531_b1 );
xor ( \533_b0 , \530_b0 , w_804 );
not ( w_804 , w_805 );
and ( w_805 , \531_b1 , \531_b0 );
or ( \534_b1 , \477_b1 , \492_b1 );
xor ( \534_b0 , \477_b0 , w_806 );
not ( w_806 , w_807 );
and ( w_807 , \492_b1 , \492_b0 );
or ( \535_b1 , \151_A[2]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_808 );
and ( \535_b0 , \151_A[2]_b0 , w_809 );
and ( w_808 , w_809 , \166_B[7]_b0 );
or ( \536_b1 , \534_b1 , \535_b1 );
not ( \535_b1 , w_810 );
and ( \536_b0 , \534_b0 , w_811 );
and ( w_810 , w_811 , \535_b0 );
or ( \537_b1 , \534_b1 , \535_b1 );
xor ( \537_b0 , \534_b0 , w_812 );
not ( w_812 , w_813 );
and ( w_813 , \535_b1 , \535_b0 );
or ( \538_b1 , \481_b1 , \490_b1 );
xor ( \538_b0 , \481_b0 , w_814 );
not ( w_814 , w_815 );
and ( w_815 , \490_b1 , \490_b0 );
or ( \539_b1 , \157_A[1]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_816 );
and ( \539_b0 , \157_A[1]_b0 , w_817 );
and ( w_816 , w_817 , \166_B[7]_b0 );
or ( \540_b1 , \538_b1 , \539_b1 );
not ( \539_b1 , w_818 );
and ( \540_b0 , \538_b0 , w_819 );
and ( w_818 , w_819 , \539_b0 );
or ( \541_b1 , \538_b1 , \539_b1 );
xor ( \541_b0 , \538_b0 , w_820 );
not ( w_820 , w_821 );
and ( w_821 , \539_b1 , \539_b0 );
or ( \542_b1 , \485_b1 , \488_b1 );
xor ( \542_b0 , \485_b0 , w_822 );
not ( w_822 , w_823 );
and ( w_823 , \488_b1 , \488_b0 );
or ( \543_b1 , \163_A[0]_b1 , \166_B[7]_b1 );
not ( \166_B[7]_b1 , w_824 );
and ( \543_b0 , \163_A[0]_b0 , w_825 );
and ( w_824 , w_825 , \166_B[7]_b0 );
or ( \544_b1 , \542_b1 , \543_b1 );
not ( \543_b1 , w_826 );
and ( \544_b0 , \542_b0 , w_827 );
and ( w_826 , w_827 , \543_b0 );
or ( \545_b1 , \541_b1 , \544_b1 );
not ( \544_b1 , w_828 );
and ( \545_b0 , \541_b0 , w_829 );
and ( w_828 , w_829 , \544_b0 );
or ( \546_b1 , \540_b1 , w_830 );
or ( \546_b0 , \540_b0 , \545_b0 );
not ( \545_b0 , w_831 );
and ( w_831 , w_830 , \545_b1 );
or ( \547_b1 , \537_b1 , \546_b1 );
not ( \546_b1 , w_832 );
and ( \547_b0 , \537_b0 , w_833 );
and ( w_832 , w_833 , \546_b0 );
or ( \548_b1 , \536_b1 , w_834 );
or ( \548_b0 , \536_b0 , \547_b0 );
not ( \547_b0 , w_835 );
and ( w_835 , w_834 , \547_b1 );
or ( \549_b1 , \533_b1 , \548_b1 );
not ( \548_b1 , w_836 );
and ( \549_b0 , \533_b0 , w_837 );
and ( w_836 , w_837 , \548_b0 );
or ( \550_b1 , \532_b1 , w_838 );
or ( \550_b0 , \532_b0 , \549_b0 );
not ( \549_b0 , w_839 );
and ( w_839 , w_838 , \549_b1 );
or ( \551_b1 , \529_b1 , \550_b1 );
not ( \550_b1 , w_840 );
and ( \551_b0 , \529_b0 , w_841 );
and ( w_840 , w_841 , \550_b0 );
or ( \552_b1 , \528_b1 , w_842 );
or ( \552_b0 , \528_b0 , \551_b0 );
not ( \551_b0 , w_843 );
and ( w_843 , w_842 , \551_b1 );
or ( \553_b1 , \525_b1 , \552_b1 );
not ( \552_b1 , w_844 );
and ( \553_b0 , \525_b0 , w_845 );
and ( w_844 , w_845 , \552_b0 );
or ( \554_b1 , \524_b1 , w_846 );
or ( \554_b0 , \524_b0 , \553_b0 );
not ( \553_b0 , w_847 );
and ( w_847 , w_846 , \553_b1 );
or ( \555_b1 , \521_b1 , \554_b1 );
not ( \554_b1 , w_848 );
and ( \555_b0 , \521_b0 , w_849 );
and ( w_848 , w_849 , \554_b0 );
or ( \556_b1 , \520_b1 , w_850 );
or ( \556_b0 , \520_b0 , \555_b0 );
not ( \555_b0 , w_851 );
and ( w_851 , w_850 , \555_b1 );
or ( \557_b1 , \517_b1 , \556_b1 );
not ( \556_b1 , w_852 );
and ( \557_b0 , \517_b0 , w_853 );
and ( w_852 , w_853 , \556_b0 );
or ( \558_b1 , \516_b1 , w_854 );
or ( \558_b0 , \516_b0 , \557_b0 );
not ( \557_b0 , w_855 );
and ( w_855 , w_854 , \557_b1 );
or ( \559_b1 , \513_b1 , \558_b1 );
not ( \558_b1 , w_856 );
and ( \559_b0 , \513_b0 , w_857 );
and ( w_856 , w_857 , \558_b0 );
or ( \560_b1 , \512_b1 , w_858 );
or ( \560_b0 , \512_b0 , \559_b0 );
not ( \559_b0 , w_859 );
and ( w_859 , w_858 , \559_b1 );
or ( \561_b1 , \509_b1 , \560_b1 );
not ( \560_b1 , w_860 );
and ( \561_b0 , \509_b0 , w_861 );
and ( w_860 , w_861 , \560_b0 );
or ( \562_b1 , \508_b1 , w_862 );
or ( \562_b0 , \508_b0 , \561_b0 );
not ( \561_b0 , w_863 );
and ( w_863 , w_862 , \561_b1 );
or ( \563_b1 , \109_A[9]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_864 );
and ( \563_b0 , \109_A[9]_b0 , w_865 );
and ( w_864 , w_865 , \165_B[8]_b0 );
or ( \564_b1 , \562_b1 , \563_b1 );
not ( \563_b1 , w_866 );
and ( \564_b0 , \562_b0 , w_867 );
and ( w_866 , w_867 , \563_b0 );
or ( \565_b1 , \562_b1 , \563_b1 );
xor ( \565_b0 , \562_b0 , w_868 );
not ( w_868 , w_869 );
and ( w_869 , \563_b1 , \563_b0 );
or ( \566_b1 , \509_b1 , \560_b1 );
xor ( \566_b0 , \509_b0 , w_870 );
not ( w_870 , w_871 );
and ( w_871 , \560_b1 , \560_b0 );
or ( \567_b1 , \115_A[8]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_872 );
and ( \567_b0 , \115_A[8]_b0 , w_873 );
and ( w_872 , w_873 , \165_B[8]_b0 );
or ( \568_b1 , \566_b1 , \567_b1 );
not ( \567_b1 , w_874 );
and ( \568_b0 , \566_b0 , w_875 );
and ( w_874 , w_875 , \567_b0 );
or ( \569_b1 , \566_b1 , \567_b1 );
xor ( \569_b0 , \566_b0 , w_876 );
not ( w_876 , w_877 );
and ( w_877 , \567_b1 , \567_b0 );
or ( \570_b1 , \513_b1 , \558_b1 );
xor ( \570_b0 , \513_b0 , w_878 );
not ( w_878 , w_879 );
and ( w_879 , \558_b1 , \558_b0 );
or ( \571_b1 , \121_A[7]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_880 );
and ( \571_b0 , \121_A[7]_b0 , w_881 );
and ( w_880 , w_881 , \165_B[8]_b0 );
or ( \572_b1 , \570_b1 , \571_b1 );
not ( \571_b1 , w_882 );
and ( \572_b0 , \570_b0 , w_883 );
and ( w_882 , w_883 , \571_b0 );
or ( \573_b1 , \570_b1 , \571_b1 );
xor ( \573_b0 , \570_b0 , w_884 );
not ( w_884 , w_885 );
and ( w_885 , \571_b1 , \571_b0 );
or ( \574_b1 , \517_b1 , \556_b1 );
xor ( \574_b0 , \517_b0 , w_886 );
not ( w_886 , w_887 );
and ( w_887 , \556_b1 , \556_b0 );
or ( \575_b1 , \127_A[6]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_888 );
and ( \575_b0 , \127_A[6]_b0 , w_889 );
and ( w_888 , w_889 , \165_B[8]_b0 );
or ( \576_b1 , \574_b1 , \575_b1 );
not ( \575_b1 , w_890 );
and ( \576_b0 , \574_b0 , w_891 );
and ( w_890 , w_891 , \575_b0 );
or ( \577_b1 , \574_b1 , \575_b1 );
xor ( \577_b0 , \574_b0 , w_892 );
not ( w_892 , w_893 );
and ( w_893 , \575_b1 , \575_b0 );
or ( \578_b1 , \521_b1 , \554_b1 );
xor ( \578_b0 , \521_b0 , w_894 );
not ( w_894 , w_895 );
and ( w_895 , \554_b1 , \554_b0 );
or ( \579_b1 , \133_A[5]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_896 );
and ( \579_b0 , \133_A[5]_b0 , w_897 );
and ( w_896 , w_897 , \165_B[8]_b0 );
or ( \580_b1 , \578_b1 , \579_b1 );
not ( \579_b1 , w_898 );
and ( \580_b0 , \578_b0 , w_899 );
and ( w_898 , w_899 , \579_b0 );
or ( \581_b1 , \578_b1 , \579_b1 );
xor ( \581_b0 , \578_b0 , w_900 );
not ( w_900 , w_901 );
and ( w_901 , \579_b1 , \579_b0 );
or ( \582_b1 , \525_b1 , \552_b1 );
xor ( \582_b0 , \525_b0 , w_902 );
not ( w_902 , w_903 );
and ( w_903 , \552_b1 , \552_b0 );
or ( \583_b1 , \139_A[4]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_904 );
and ( \583_b0 , \139_A[4]_b0 , w_905 );
and ( w_904 , w_905 , \165_B[8]_b0 );
or ( \584_b1 , \582_b1 , \583_b1 );
not ( \583_b1 , w_906 );
and ( \584_b0 , \582_b0 , w_907 );
and ( w_906 , w_907 , \583_b0 );
or ( \585_b1 , \582_b1 , \583_b1 );
xor ( \585_b0 , \582_b0 , w_908 );
not ( w_908 , w_909 );
and ( w_909 , \583_b1 , \583_b0 );
or ( \586_b1 , \529_b1 , \550_b1 );
xor ( \586_b0 , \529_b0 , w_910 );
not ( w_910 , w_911 );
and ( w_911 , \550_b1 , \550_b0 );
or ( \587_b1 , \145_A[3]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_912 );
and ( \587_b0 , \145_A[3]_b0 , w_913 );
and ( w_912 , w_913 , \165_B[8]_b0 );
or ( \588_b1 , \586_b1 , \587_b1 );
not ( \587_b1 , w_914 );
and ( \588_b0 , \586_b0 , w_915 );
and ( w_914 , w_915 , \587_b0 );
or ( \589_b1 , \586_b1 , \587_b1 );
xor ( \589_b0 , \586_b0 , w_916 );
not ( w_916 , w_917 );
and ( w_917 , \587_b1 , \587_b0 );
or ( \590_b1 , \533_b1 , \548_b1 );
xor ( \590_b0 , \533_b0 , w_918 );
not ( w_918 , w_919 );
and ( w_919 , \548_b1 , \548_b0 );
or ( \591_b1 , \151_A[2]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_920 );
and ( \591_b0 , \151_A[2]_b0 , w_921 );
and ( w_920 , w_921 , \165_B[8]_b0 );
or ( \592_b1 , \590_b1 , \591_b1 );
not ( \591_b1 , w_922 );
and ( \592_b0 , \590_b0 , w_923 );
and ( w_922 , w_923 , \591_b0 );
or ( \593_b1 , \590_b1 , \591_b1 );
xor ( \593_b0 , \590_b0 , w_924 );
not ( w_924 , w_925 );
and ( w_925 , \591_b1 , \591_b0 );
or ( \594_b1 , \537_b1 , \546_b1 );
xor ( \594_b0 , \537_b0 , w_926 );
not ( w_926 , w_927 );
and ( w_927 , \546_b1 , \546_b0 );
or ( \595_b1 , \157_A[1]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_928 );
and ( \595_b0 , \157_A[1]_b0 , w_929 );
and ( w_928 , w_929 , \165_B[8]_b0 );
or ( \596_b1 , \594_b1 , \595_b1 );
not ( \595_b1 , w_930 );
and ( \596_b0 , \594_b0 , w_931 );
and ( w_930 , w_931 , \595_b0 );
or ( \597_b1 , \594_b1 , \595_b1 );
xor ( \597_b0 , \594_b0 , w_932 );
not ( w_932 , w_933 );
and ( w_933 , \595_b1 , \595_b0 );
or ( \598_b1 , \541_b1 , \544_b1 );
xor ( \598_b0 , \541_b0 , w_934 );
not ( w_934 , w_935 );
and ( w_935 , \544_b1 , \544_b0 );
or ( \599_b1 , \163_A[0]_b1 , \165_B[8]_b1 );
not ( \165_B[8]_b1 , w_936 );
and ( \599_b0 , \163_A[0]_b0 , w_937 );
and ( w_936 , w_937 , \165_B[8]_b0 );
or ( \600_b1 , \598_b1 , \599_b1 );
not ( \599_b1 , w_938 );
and ( \600_b0 , \598_b0 , w_939 );
and ( w_938 , w_939 , \599_b0 );
or ( \601_b1 , \597_b1 , \600_b1 );
not ( \600_b1 , w_940 );
and ( \601_b0 , \597_b0 , w_941 );
and ( w_940 , w_941 , \600_b0 );
or ( \602_b1 , \596_b1 , w_942 );
or ( \602_b0 , \596_b0 , \601_b0 );
not ( \601_b0 , w_943 );
and ( w_943 , w_942 , \601_b1 );
or ( \603_b1 , \593_b1 , \602_b1 );
not ( \602_b1 , w_944 );
and ( \603_b0 , \593_b0 , w_945 );
and ( w_944 , w_945 , \602_b0 );
or ( \604_b1 , \592_b1 , w_946 );
or ( \604_b0 , \592_b0 , \603_b0 );
not ( \603_b0 , w_947 );
and ( w_947 , w_946 , \603_b1 );
or ( \605_b1 , \589_b1 , \604_b1 );
not ( \604_b1 , w_948 );
and ( \605_b0 , \589_b0 , w_949 );
and ( w_948 , w_949 , \604_b0 );
or ( \606_b1 , \588_b1 , w_950 );
or ( \606_b0 , \588_b0 , \605_b0 );
not ( \605_b0 , w_951 );
and ( w_951 , w_950 , \605_b1 );
or ( \607_b1 , \585_b1 , \606_b1 );
not ( \606_b1 , w_952 );
and ( \607_b0 , \585_b0 , w_953 );
and ( w_952 , w_953 , \606_b0 );
or ( \608_b1 , \584_b1 , w_954 );
or ( \608_b0 , \584_b0 , \607_b0 );
not ( \607_b0 , w_955 );
and ( w_955 , w_954 , \607_b1 );
or ( \609_b1 , \581_b1 , \608_b1 );
not ( \608_b1 , w_956 );
and ( \609_b0 , \581_b0 , w_957 );
and ( w_956 , w_957 , \608_b0 );
or ( \610_b1 , \580_b1 , w_958 );
or ( \610_b0 , \580_b0 , \609_b0 );
not ( \609_b0 , w_959 );
and ( w_959 , w_958 , \609_b1 );
or ( \611_b1 , \577_b1 , \610_b1 );
not ( \610_b1 , w_960 );
and ( \611_b0 , \577_b0 , w_961 );
and ( w_960 , w_961 , \610_b0 );
or ( \612_b1 , \576_b1 , w_962 );
or ( \612_b0 , \576_b0 , \611_b0 );
not ( \611_b0 , w_963 );
and ( w_963 , w_962 , \611_b1 );
or ( \613_b1 , \573_b1 , \612_b1 );
not ( \612_b1 , w_964 );
and ( \613_b0 , \573_b0 , w_965 );
and ( w_964 , w_965 , \612_b0 );
or ( \614_b1 , \572_b1 , w_966 );
or ( \614_b0 , \572_b0 , \613_b0 );
not ( \613_b0 , w_967 );
and ( w_967 , w_966 , \613_b1 );
or ( \615_b1 , \569_b1 , \614_b1 );
not ( \614_b1 , w_968 );
and ( \615_b0 , \569_b0 , w_969 );
and ( w_968 , w_969 , \614_b0 );
or ( \616_b1 , \568_b1 , w_970 );
or ( \616_b0 , \568_b0 , \615_b0 );
not ( \615_b0 , w_971 );
and ( w_971 , w_970 , \615_b1 );
or ( \617_b1 , \565_b1 , \616_b1 );
not ( \616_b1 , w_972 );
and ( \617_b0 , \565_b0 , w_973 );
and ( w_972 , w_973 , \616_b0 );
or ( \618_b1 , \564_b1 , w_974 );
or ( \618_b0 , \564_b0 , \617_b0 );
not ( \617_b0 , w_975 );
and ( w_975 , w_974 , \617_b1 );
or ( \619_b1 , \109_A[9]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_976 );
and ( \619_b0 , \109_A[9]_b0 , w_977 );
and ( w_976 , w_977 , \164_B[9]_b0 );
or ( \620_b1 , \618_b1 , \619_b1 );
not ( \619_b1 , w_978 );
and ( \620_b0 , \618_b0 , w_979 );
and ( w_978 , w_979 , \619_b0 );
or ( \621_b1 , \618_b1 , \619_b1 );
xor ( \621_b0 , \618_b0 , w_980 );
not ( w_980 , w_981 );
and ( w_981 , \619_b1 , \619_b0 );
or ( \622_b1 , \565_b1 , \616_b1 );
xor ( \622_b0 , \565_b0 , w_982 );
not ( w_982 , w_983 );
and ( w_983 , \616_b1 , \616_b0 );
or ( \623_b1 , \115_A[8]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_984 );
and ( \623_b0 , \115_A[8]_b0 , w_985 );
and ( w_984 , w_985 , \164_B[9]_b0 );
or ( \624_b1 , \622_b1 , \623_b1 );
not ( \623_b1 , w_986 );
and ( \624_b0 , \622_b0 , w_987 );
and ( w_986 , w_987 , \623_b0 );
or ( \625_b1 , \622_b1 , \623_b1 );
xor ( \625_b0 , \622_b0 , w_988 );
not ( w_988 , w_989 );
and ( w_989 , \623_b1 , \623_b0 );
or ( \626_b1 , \569_b1 , \614_b1 );
xor ( \626_b0 , \569_b0 , w_990 );
not ( w_990 , w_991 );
and ( w_991 , \614_b1 , \614_b0 );
or ( \627_b1 , \121_A[7]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_992 );
and ( \627_b0 , \121_A[7]_b0 , w_993 );
and ( w_992 , w_993 , \164_B[9]_b0 );
or ( \628_b1 , \626_b1 , \627_b1 );
not ( \627_b1 , w_994 );
and ( \628_b0 , \626_b0 , w_995 );
and ( w_994 , w_995 , \627_b0 );
or ( \629_b1 , \626_b1 , \627_b1 );
xor ( \629_b0 , \626_b0 , w_996 );
not ( w_996 , w_997 );
and ( w_997 , \627_b1 , \627_b0 );
or ( \630_b1 , \573_b1 , \612_b1 );
xor ( \630_b0 , \573_b0 , w_998 );
not ( w_998 , w_999 );
and ( w_999 , \612_b1 , \612_b0 );
or ( \631_b1 , \127_A[6]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1000 );
and ( \631_b0 , \127_A[6]_b0 , w_1001 );
and ( w_1000 , w_1001 , \164_B[9]_b0 );
or ( \632_b1 , \630_b1 , \631_b1 );
not ( \631_b1 , w_1002 );
and ( \632_b0 , \630_b0 , w_1003 );
and ( w_1002 , w_1003 , \631_b0 );
or ( \633_b1 , \630_b1 , \631_b1 );
xor ( \633_b0 , \630_b0 , w_1004 );
not ( w_1004 , w_1005 );
and ( w_1005 , \631_b1 , \631_b0 );
or ( \634_b1 , \577_b1 , \610_b1 );
xor ( \634_b0 , \577_b0 , w_1006 );
not ( w_1006 , w_1007 );
and ( w_1007 , \610_b1 , \610_b0 );
or ( \635_b1 , \133_A[5]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1008 );
and ( \635_b0 , \133_A[5]_b0 , w_1009 );
and ( w_1008 , w_1009 , \164_B[9]_b0 );
or ( \636_b1 , \634_b1 , \635_b1 );
not ( \635_b1 , w_1010 );
and ( \636_b0 , \634_b0 , w_1011 );
and ( w_1010 , w_1011 , \635_b0 );
or ( \637_b1 , \634_b1 , \635_b1 );
xor ( \637_b0 , \634_b0 , w_1012 );
not ( w_1012 , w_1013 );
and ( w_1013 , \635_b1 , \635_b0 );
or ( \638_b1 , \581_b1 , \608_b1 );
xor ( \638_b0 , \581_b0 , w_1014 );
not ( w_1014 , w_1015 );
and ( w_1015 , \608_b1 , \608_b0 );
or ( \639_b1 , \139_A[4]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1016 );
and ( \639_b0 , \139_A[4]_b0 , w_1017 );
and ( w_1016 , w_1017 , \164_B[9]_b0 );
or ( \640_b1 , \638_b1 , \639_b1 );
not ( \639_b1 , w_1018 );
and ( \640_b0 , \638_b0 , w_1019 );
and ( w_1018 , w_1019 , \639_b0 );
or ( \641_b1 , \638_b1 , \639_b1 );
xor ( \641_b0 , \638_b0 , w_1020 );
not ( w_1020 , w_1021 );
and ( w_1021 , \639_b1 , \639_b0 );
or ( \642_b1 , \585_b1 , \606_b1 );
xor ( \642_b0 , \585_b0 , w_1022 );
not ( w_1022 , w_1023 );
and ( w_1023 , \606_b1 , \606_b0 );
or ( \643_b1 , \145_A[3]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1024 );
and ( \643_b0 , \145_A[3]_b0 , w_1025 );
and ( w_1024 , w_1025 , \164_B[9]_b0 );
or ( \644_b1 , \642_b1 , \643_b1 );
not ( \643_b1 , w_1026 );
and ( \644_b0 , \642_b0 , w_1027 );
and ( w_1026 , w_1027 , \643_b0 );
or ( \645_b1 , \642_b1 , \643_b1 );
xor ( \645_b0 , \642_b0 , w_1028 );
not ( w_1028 , w_1029 );
and ( w_1029 , \643_b1 , \643_b0 );
or ( \646_b1 , \589_b1 , \604_b1 );
xor ( \646_b0 , \589_b0 , w_1030 );
not ( w_1030 , w_1031 );
and ( w_1031 , \604_b1 , \604_b0 );
or ( \647_b1 , \151_A[2]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1032 );
and ( \647_b0 , \151_A[2]_b0 , w_1033 );
and ( w_1032 , w_1033 , \164_B[9]_b0 );
or ( \648_b1 , \646_b1 , \647_b1 );
not ( \647_b1 , w_1034 );
and ( \648_b0 , \646_b0 , w_1035 );
and ( w_1034 , w_1035 , \647_b0 );
or ( \649_b1 , \646_b1 , \647_b1 );
xor ( \649_b0 , \646_b0 , w_1036 );
not ( w_1036 , w_1037 );
and ( w_1037 , \647_b1 , \647_b0 );
or ( \650_b1 , \593_b1 , \602_b1 );
xor ( \650_b0 , \593_b0 , w_1038 );
not ( w_1038 , w_1039 );
and ( w_1039 , \602_b1 , \602_b0 );
or ( \651_b1 , \157_A[1]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1040 );
and ( \651_b0 , \157_A[1]_b0 , w_1041 );
and ( w_1040 , w_1041 , \164_B[9]_b0 );
or ( \652_b1 , \650_b1 , \651_b1 );
not ( \651_b1 , w_1042 );
and ( \652_b0 , \650_b0 , w_1043 );
and ( w_1042 , w_1043 , \651_b0 );
or ( \653_b1 , \650_b1 , \651_b1 );
xor ( \653_b0 , \650_b0 , w_1044 );
not ( w_1044 , w_1045 );
and ( w_1045 , \651_b1 , \651_b0 );
or ( \654_b1 , \597_b1 , \600_b1 );
xor ( \654_b0 , \597_b0 , w_1046 );
not ( w_1046 , w_1047 );
and ( w_1047 , \600_b1 , \600_b0 );
or ( \655_b1 , \163_A[0]_b1 , \164_B[9]_b1 );
not ( \164_B[9]_b1 , w_1048 );
and ( \655_b0 , \163_A[0]_b0 , w_1049 );
and ( w_1048 , w_1049 , \164_B[9]_b0 );
or ( \656_b1 , \654_b1 , \655_b1 );
not ( \655_b1 , w_1050 );
and ( \656_b0 , \654_b0 , w_1051 );
and ( w_1050 , w_1051 , \655_b0 );
or ( \657_b1 , \653_b1 , \656_b1 );
not ( \656_b1 , w_1052 );
and ( \657_b0 , \653_b0 , w_1053 );
and ( w_1052 , w_1053 , \656_b0 );
or ( \658_b1 , \652_b1 , w_1054 );
or ( \658_b0 , \652_b0 , \657_b0 );
not ( \657_b0 , w_1055 );
and ( w_1055 , w_1054 , \657_b1 );
or ( \659_b1 , \649_b1 , \658_b1 );
not ( \658_b1 , w_1056 );
and ( \659_b0 , \649_b0 , w_1057 );
and ( w_1056 , w_1057 , \658_b0 );
or ( \660_b1 , \648_b1 , w_1058 );
or ( \660_b0 , \648_b0 , \659_b0 );
not ( \659_b0 , w_1059 );
and ( w_1059 , w_1058 , \659_b1 );
or ( \661_b1 , \645_b1 , \660_b1 );
not ( \660_b1 , w_1060 );
and ( \661_b0 , \645_b0 , w_1061 );
and ( w_1060 , w_1061 , \660_b0 );
or ( \662_b1 , \644_b1 , w_1062 );
or ( \662_b0 , \644_b0 , \661_b0 );
not ( \661_b0 , w_1063 );
and ( w_1063 , w_1062 , \661_b1 );
or ( \663_b1 , \641_b1 , \662_b1 );
not ( \662_b1 , w_1064 );
and ( \663_b0 , \641_b0 , w_1065 );
and ( w_1064 , w_1065 , \662_b0 );
or ( \664_b1 , \640_b1 , w_1066 );
or ( \664_b0 , \640_b0 , \663_b0 );
not ( \663_b0 , w_1067 );
and ( w_1067 , w_1066 , \663_b1 );
or ( \665_b1 , \637_b1 , \664_b1 );
not ( \664_b1 , w_1068 );
and ( \665_b0 , \637_b0 , w_1069 );
and ( w_1068 , w_1069 , \664_b0 );
or ( \666_b1 , \636_b1 , w_1070 );
or ( \666_b0 , \636_b0 , \665_b0 );
not ( \665_b0 , w_1071 );
and ( w_1071 , w_1070 , \665_b1 );
or ( \667_b1 , \633_b1 , \666_b1 );
not ( \666_b1 , w_1072 );
and ( \667_b0 , \633_b0 , w_1073 );
and ( w_1072 , w_1073 , \666_b0 );
or ( \668_b1 , \632_b1 , w_1074 );
or ( \668_b0 , \632_b0 , \667_b0 );
not ( \667_b0 , w_1075 );
and ( w_1075 , w_1074 , \667_b1 );
or ( \669_b1 , \629_b1 , \668_b1 );
not ( \668_b1 , w_1076 );
and ( \669_b0 , \629_b0 , w_1077 );
and ( w_1076 , w_1077 , \668_b0 );
or ( \670_b1 , \628_b1 , w_1078 );
or ( \670_b0 , \628_b0 , \669_b0 );
not ( \669_b0 , w_1079 );
and ( w_1079 , w_1078 , \669_b1 );
or ( \671_b1 , \625_b1 , \670_b1 );
not ( \670_b1 , w_1080 );
and ( \671_b0 , \625_b0 , w_1081 );
and ( w_1080 , w_1081 , \670_b0 );
or ( \672_b1 , \624_b1 , w_1082 );
or ( \672_b0 , \624_b0 , \671_b0 );
not ( \671_b0 , w_1083 );
and ( w_1083 , w_1082 , \671_b1 );
or ( \673_b1 , \621_b1 , \672_b1 );
not ( \672_b1 , w_1084 );
and ( \673_b0 , \621_b0 , w_1085 );
and ( w_1084 , w_1085 , \672_b0 );
or ( \674_b1 , \620_b1 , w_1086 );
or ( \674_b0 , \620_b0 , \673_b0 );
not ( \673_b0 , w_1087 );
and ( w_1087 , w_1086 , \673_b1 );
buf ( \675_Z[19]_b1 , \674_b1 );
buf ( \675_Z[19]_b0 , \674_b0 );
or ( \676_b1 , \621_b1 , \672_b1 );
xor ( \676_b0 , \621_b0 , w_1088 );
not ( w_1088 , w_1089 );
and ( w_1089 , \672_b1 , \672_b0 );
buf ( \677_Z[18]_b1 , \676_b1 );
buf ( \677_Z[18]_b0 , \676_b0 );
or ( \678_b1 , \625_b1 , \670_b1 );
xor ( \678_b0 , \625_b0 , w_1090 );
not ( w_1090 , w_1091 );
and ( w_1091 , \670_b1 , \670_b0 );
buf ( \679_Z[17]_b1 , \678_b1 );
buf ( \679_Z[17]_b0 , \678_b0 );
or ( \680_b1 , \629_b1 , \668_b1 );
xor ( \680_b0 , \629_b0 , w_1092 );
not ( w_1092 , w_1093 );
and ( w_1093 , \668_b1 , \668_b0 );
buf ( \681_Z[16]_b1 , \680_b1 );
buf ( \681_Z[16]_b0 , \680_b0 );
or ( \682_b1 , \633_b1 , \666_b1 );
xor ( \682_b0 , \633_b0 , w_1094 );
not ( w_1094 , w_1095 );
and ( w_1095 , \666_b1 , \666_b0 );
buf ( \683_Z[15]_b1 , \682_b1 );
buf ( \683_Z[15]_b0 , \682_b0 );
or ( \684_b1 , \637_b1 , \664_b1 );
xor ( \684_b0 , \637_b0 , w_1096 );
not ( w_1096 , w_1097 );
and ( w_1097 , \664_b1 , \664_b0 );
buf ( \685_Z[14]_b1 , \684_b1 );
buf ( \685_Z[14]_b0 , \684_b0 );
or ( \686_b1 , \641_b1 , \662_b1 );
xor ( \686_b0 , \641_b0 , w_1098 );
not ( w_1098 , w_1099 );
and ( w_1099 , \662_b1 , \662_b0 );
buf ( \687_Z[13]_b1 , \686_b1 );
buf ( \687_Z[13]_b0 , \686_b0 );
or ( \688_b1 , \645_b1 , \660_b1 );
xor ( \688_b0 , \645_b0 , w_1100 );
not ( w_1100 , w_1101 );
and ( w_1101 , \660_b1 , \660_b0 );
buf ( \689_Z[12]_b1 , \688_b1 );
buf ( \689_Z[12]_b0 , \688_b0 );
or ( \690_b1 , \649_b1 , \658_b1 );
xor ( \690_b0 , \649_b0 , w_1102 );
not ( w_1102 , w_1103 );
and ( w_1103 , \658_b1 , \658_b0 );
buf ( \691_Z[11]_b1 , \690_b1 );
buf ( \691_Z[11]_b0 , \690_b0 );
or ( \692_b1 , \653_b1 , \656_b1 );
xor ( \692_b0 , \653_b0 , w_1104 );
not ( w_1104 , w_1105 );
and ( w_1105 , \656_b1 , \656_b0 );
buf ( \693_Z[10]_b1 , \692_b1 );
buf ( \693_Z[10]_b0 , \692_b0 );
or ( \694_b1 , \654_b1 , \655_b1 );
xor ( \694_b0 , \654_b0 , w_1106 );
not ( w_1106 , w_1107 );
and ( w_1107 , \655_b1 , \655_b0 );
buf ( \695_Z[9]_b1 , \694_b1 );
buf ( \695_Z[9]_b0 , \694_b0 );
or ( \696_b1 , \598_b1 , \599_b1 );
xor ( \696_b0 , \598_b0 , w_1108 );
not ( w_1108 , w_1109 );
and ( w_1109 , \599_b1 , \599_b0 );
buf ( \697_Z[8]_b1 , \696_b1 );
buf ( \697_Z[8]_b0 , \696_b0 );
or ( \698_b1 , \542_b1 , \543_b1 );
xor ( \698_b0 , \542_b0 , w_1110 );
not ( w_1110 , w_1111 );
and ( w_1111 , \543_b1 , \543_b0 );
buf ( \699_Z[7]_b1 , \698_b1 );
buf ( \699_Z[7]_b0 , \698_b0 );
or ( \700_b1 , \486_b1 , \487_b1 );
xor ( \700_b0 , \486_b0 , w_1112 );
not ( w_1112 , w_1113 );
and ( w_1113 , \487_b1 , \487_b0 );
buf ( \701_Z[6]_b1 , \700_b1 );
buf ( \701_Z[6]_b0 , \700_b0 );
or ( \702_b1 , \430_b1 , \431_b1 );
xor ( \702_b0 , \430_b0 , w_1114 );
not ( w_1114 , w_1115 );
and ( w_1115 , \431_b1 , \431_b0 );
buf ( \703_Z[5]_b1 , \702_b1 );
buf ( \703_Z[5]_b0 , \702_b0 );
or ( \704_b1 , \374_b1 , \375_b1 );
xor ( \704_b0 , \374_b0 , w_1116 );
not ( w_1116 , w_1117 );
and ( w_1117 , \375_b1 , \375_b0 );
buf ( \705_Z[4]_b1 , \704_b1 );
buf ( \705_Z[4]_b0 , \704_b0 );
or ( \706_b1 , \318_b1 , \319_b1 );
xor ( \706_b0 , \318_b0 , w_1118 );
not ( w_1118 , w_1119 );
and ( w_1119 , \319_b1 , \319_b0 );
buf ( \707_Z[3]_b1 , \706_b1 );
buf ( \707_Z[3]_b0 , \706_b0 );
or ( \708_b1 , \262_b1 , \263_b1 );
xor ( \708_b0 , \262_b0 , w_1120 );
not ( w_1120 , w_1121 );
and ( w_1121 , \263_b1 , \263_b0 );
buf ( \709_Z[2]_b1 , \708_b1 );
buf ( \709_Z[2]_b0 , \708_b0 );
or ( \710_b1 , \207_b1 , \208_b1 );
xor ( \710_b0 , \207_b0 , w_1122 );
not ( w_1122 , w_1123 );
and ( w_1123 , \208_b1 , \208_b0 );
buf ( \711_Z[1]_b1 , \710_b1 );
buf ( \711_Z[1]_b0 , \710_b0 );
or ( \712_b1 , \163_A[0]_b1 , \173_B[0]_b1 );
not ( \173_B[0]_b1 , w_1124 );
and ( \712_b0 , \163_A[0]_b0 , w_1125 );
and ( w_1124 , w_1125 , \173_B[0]_b0 );
buf ( \713_Z[0]_b1 , \712_b1 );
buf ( \713_Z[0]_b0 , \712_b0 );
or ( \89_b1 , \I[0]_b1 , w_1140 );
or ( \89_b0 , \I[0]_b0 , w_1127 );
not ( w_1127 , w_1141 );
and ( w_1141 , w_1140 , w_1126 );
or ( w_1126 , \88_b1 , w_1142 );
or ( w_1127 , \88_b0 , w_1129 );
not ( w_1129 , w_1143 );
and ( w_1143 , w_1142 , w_1128 );
or ( w_1128 , \I[2]_b1 , w_1144 );
or ( w_1129 , \I[2]_b0 , w_1131 );
not ( w_1131 , w_1145 );
and ( w_1145 , w_1144 , w_1130 );
or ( w_1130 , \I[3]_b1 , w_1146 );
or ( w_1131 , \I[3]_b0 , w_1133 );
not ( w_1133 , w_1147 );
and ( w_1147 , w_1146 , w_1132 );
or ( w_1132 , \I[4]_b1 , w_1148 );
or ( w_1133 , \I[4]_b0 , w_1135 );
not ( w_1135 , w_1149 );
and ( w_1149 , w_1148 , w_1134 );
or ( w_1134 , \I[5]_b1 , w_1150 );
or ( w_1135 , \I[5]_b0 , w_1137 );
not ( w_1137 , w_1151 );
and ( w_1151 , w_1150 , w_1136 );
or ( w_1136 , \I[6]_b1 , w_1152 );
or ( w_1137 , \I[6]_b0 , w_1139 );
not ( w_1139 , w_1153 );
and ( w_1153 , w_1152 , w_1138 );
buf ( w_1138 , \I[7]_b1 );
not ( w_1138 , w_1154 );
not ( w_1139 , w_1155 );
and ( w_1154 , w_1155 , \I[7]_b0 );
or ( \92_b1 , \91_b1 , w_1170 );
or ( \92_b0 , \91_b0 , w_1157 );
not ( w_1157 , w_1171 );
and ( w_1171 , w_1170 , w_1156 );
or ( w_1156 , \I[1]_b1 , w_1172 );
or ( w_1157 , \I[1]_b0 , w_1159 );
not ( w_1159 , w_1173 );
and ( w_1173 , w_1172 , w_1158 );
or ( w_1158 , \I[2]_b1 , w_1174 );
or ( w_1159 , \I[2]_b0 , w_1161 );
not ( w_1161 , w_1175 );
and ( w_1175 , w_1174 , w_1160 );
or ( w_1160 , \I[3]_b1 , w_1176 );
or ( w_1161 , \I[3]_b0 , w_1163 );
not ( w_1163 , w_1177 );
and ( w_1177 , w_1176 , w_1162 );
or ( w_1162 , \I[4]_b1 , w_1178 );
or ( w_1163 , \I[4]_b0 , w_1165 );
not ( w_1165 , w_1179 );
and ( w_1179 , w_1178 , w_1164 );
or ( w_1164 , \I[5]_b1 , w_1180 );
or ( w_1165 , \I[5]_b0 , w_1167 );
not ( w_1167 , w_1181 );
and ( w_1181 , w_1180 , w_1166 );
or ( w_1166 , \I[6]_b1 , w_1182 );
or ( w_1167 , \I[6]_b0 , w_1169 );
not ( w_1169 , w_1183 );
and ( w_1183 , w_1182 , w_1168 );
buf ( w_1168 , \I[7]_b1 );
not ( w_1168 , w_1184 );
not ( w_1169 , w_1185 );
and ( w_1184 , w_1185 , \I[7]_b0 );
or ( \94_b1 , \I[0]_b1 , w_1200 );
or ( \94_b0 , \I[0]_b0 , w_1187 );
not ( w_1187 , w_1201 );
and ( w_1201 , w_1200 , w_1186 );
or ( w_1186 , \I[1]_b1 , w_1202 );
or ( w_1187 , \I[1]_b0 , w_1189 );
not ( w_1189 , w_1203 );
and ( w_1203 , w_1202 , w_1188 );
or ( w_1188 , \I[2]_b1 , w_1204 );
or ( w_1189 , \I[2]_b0 , w_1191 );
not ( w_1191 , w_1205 );
and ( w_1205 , w_1204 , w_1190 );
or ( w_1190 , \I[3]_b1 , w_1206 );
or ( w_1191 , \I[3]_b0 , w_1193 );
not ( w_1193 , w_1207 );
and ( w_1207 , w_1206 , w_1192 );
or ( w_1192 , \I[4]_b1 , w_1208 );
or ( w_1193 , \I[4]_b0 , w_1195 );
not ( w_1195 , w_1209 );
and ( w_1209 , w_1208 , w_1194 );
or ( w_1194 , \I[5]_b1 , w_1210 );
or ( w_1195 , \I[5]_b0 , w_1197 );
not ( w_1197 , w_1211 );
and ( w_1211 , w_1210 , w_1196 );
or ( w_1196 , \I[6]_b1 , w_1212 );
or ( w_1197 , \I[6]_b0 , w_1199 );
not ( w_1199 , w_1213 );
and ( w_1213 , w_1212 , w_1198 );
buf ( w_1198 , \I[7]_b1 );
not ( w_1198 , w_1214 );
not ( w_1199 , w_1215 );
and ( w_1214 , w_1215 , \I[7]_b0 );
or ( \96_b1 , \90_b1 , w_1218 );
or ( \96_b0 , \90_b0 , w_1217 );
not ( w_1217 , w_1219 );
and ( w_1219 , w_1218 , w_1216 );
or ( w_1216 , \93_b1 , w_1220 );
or ( w_1217 , \93_b0 , \95_b0 );
not ( \95_b0 , w_1221 );
and ( w_1221 , w_1220 , \95_b1 );
or ( \106_b1 , \97_b1 , w_1232 );
or ( \106_b0 , \97_b0 , w_1223 );
not ( w_1223 , w_1233 );
and ( w_1233 , w_1232 , w_1222 );
or ( w_1222 , \98_b1 , w_1234 );
or ( w_1223 , \98_b0 , w_1225 );
not ( w_1225 , w_1235 );
and ( w_1235 , w_1234 , w_1224 );
or ( w_1224 , \99_b1 , w_1236 );
or ( w_1225 , \99_b0 , w_1227 );
not ( w_1227 , w_1237 );
and ( w_1237 , w_1236 , w_1226 );
or ( w_1226 , \100_b1 , w_1238 );
or ( w_1227 , \100_b0 , w_1229 );
not ( w_1229 , w_1239 );
and ( w_1239 , w_1238 , w_1228 );
or ( w_1228 , \101_b1 , w_1240 );
or ( w_1229 , \101_b0 , w_1231 );
not ( w_1231 , w_1241 );
and ( w_1241 , w_1240 , w_1230 );
or ( w_1230 , \102_b1 , w_1242 );
or ( w_1231 , \102_b0 , \105_b0 );
not ( \105_b0 , w_1243 );
and ( w_1243 , w_1242 , \105_b1 );
or ( \113_b1 , \110_b1 , w_1246 );
or ( \113_b0 , \110_b0 , w_1245 );
not ( w_1245 , w_1247 );
and ( w_1247 , w_1246 , w_1244 );
or ( w_1244 , \111_b1 , w_1248 );
or ( w_1245 , \111_b0 , \112_b0 );
not ( \112_b0 , w_1249 );
and ( w_1249 , w_1248 , \112_b1 );
or ( \119_b1 , \116_b1 , w_1252 );
or ( \119_b0 , \116_b0 , w_1251 );
not ( w_1251 , w_1253 );
and ( w_1253 , w_1252 , w_1250 );
or ( w_1250 , \117_b1 , w_1254 );
or ( w_1251 , \117_b0 , \118_b0 );
not ( \118_b0 , w_1255 );
and ( w_1255 , w_1254 , \118_b1 );
or ( \125_b1 , \122_b1 , w_1258 );
or ( \125_b0 , \122_b0 , w_1257 );
not ( w_1257 , w_1259 );
and ( w_1259 , w_1258 , w_1256 );
or ( w_1256 , \123_b1 , w_1260 );
or ( w_1257 , \123_b0 , \124_b0 );
not ( \124_b0 , w_1261 );
and ( w_1261 , w_1260 , \124_b1 );
or ( \131_b1 , \128_b1 , w_1264 );
or ( \131_b0 , \128_b0 , w_1263 );
not ( w_1263 , w_1265 );
and ( w_1265 , w_1264 , w_1262 );
or ( w_1262 , \129_b1 , w_1266 );
or ( w_1263 , \129_b0 , \130_b0 );
not ( \130_b0 , w_1267 );
and ( w_1267 , w_1266 , \130_b1 );
or ( \137_b1 , \134_b1 , w_1270 );
or ( \137_b0 , \134_b0 , w_1269 );
not ( w_1269 , w_1271 );
and ( w_1271 , w_1270 , w_1268 );
or ( w_1268 , \135_b1 , w_1272 );
or ( w_1269 , \135_b0 , \136_b0 );
not ( \136_b0 , w_1273 );
and ( w_1273 , w_1272 , \136_b1 );
or ( \143_b1 , \140_b1 , w_1276 );
or ( \143_b0 , \140_b0 , w_1275 );
not ( w_1275 , w_1277 );
and ( w_1277 , w_1276 , w_1274 );
or ( w_1274 , \141_b1 , w_1278 );
or ( w_1275 , \141_b0 , \142_b0 );
not ( \142_b0 , w_1279 );
and ( w_1279 , w_1278 , \142_b1 );
or ( \149_b1 , \146_b1 , w_1282 );
or ( \149_b0 , \146_b0 , w_1281 );
not ( w_1281 , w_1283 );
and ( w_1283 , w_1282 , w_1280 );
or ( w_1280 , \147_b1 , w_1284 );
or ( w_1281 , \147_b0 , \148_b0 );
not ( \148_b0 , w_1285 );
and ( w_1285 , w_1284 , \148_b1 );
or ( \155_b1 , \152_b1 , w_1288 );
or ( \155_b0 , \152_b0 , w_1287 );
not ( w_1287 , w_1289 );
and ( w_1289 , w_1288 , w_1286 );
or ( w_1286 , \153_b1 , w_1290 );
or ( w_1287 , \153_b0 , \154_b0 );
not ( \154_b0 , w_1291 );
and ( w_1291 , w_1290 , \154_b1 );
or ( \161_b1 , \158_b1 , w_1294 );
or ( \161_b0 , \158_b0 , w_1293 );
not ( w_1293 , w_1295 );
and ( w_1295 , w_1294 , w_1292 );
or ( w_1292 , \159_b1 , w_1296 );
or ( w_1293 , \159_b0 , \160_b0 );
not ( \160_b0 , w_1297 );
and ( w_1297 , w_1296 , \160_b1 );
endmodule

