// ...
module top(\a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,
		\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,
		\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,
		\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,\a[0]_b1 ,\a[0]_b0 ,\b[15]_b1 ,\b[15]_b0 ,\b[14]_b1 ,\b[14]_b0 ,
		\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,\b[10]_b0 ,\b[9]_b1 ,
		\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,\b[5]_b1 ,\b[5]_b0 ,
		\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,\b[1]_b0 ,\b[0]_b1 ,
		\b[0]_b0 ,\c[15]_b1 ,\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,
		\c[11]_b1 ,\c[11]_b0 ,\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,
		\c[7]_b0 ,\c[6]_b1 ,\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,
		\c[2]_b1 ,\c[2]_b0 ,\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,
		\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,
		\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,
		\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,
		\d[0]_b1 ,\d[0]_b0 ,\o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,
		\o[28]_b0 ,\o[27]_b1 ,\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,
		\o[23]_b1 ,\o[23]_b0 ,\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,
		\o[19]_b0 ,\o[18]_b1 ,\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,
		\o[14]_b1 ,\o[14]_b0 ,\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,
		\o[10]_b0 ,\o[9]_b1 ,\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,
		\o[5]_b1 ,\o[5]_b0 ,\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,
		\o[1]_b0 ,\o[0]_b1 ,\o[0]_b0 );
input \a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,
		\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,
		\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,
		\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,\a[0]_b1 ,\a[0]_b0 ,\b[15]_b1 ,\b[15]_b0 ,\b[14]_b1 ,\b[14]_b0 ,
		\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,\b[10]_b0 ,\b[9]_b1 ,
		\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,\b[5]_b1 ,\b[5]_b0 ,
		\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,\b[1]_b0 ,\b[0]_b1 ,
		\b[0]_b0 ,\c[15]_b1 ,\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,
		\c[11]_b1 ,\c[11]_b0 ,\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,
		\c[7]_b0 ,\c[6]_b1 ,\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,
		\c[2]_b1 ,\c[2]_b0 ,\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,
		\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,
		\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,
		\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,
		\d[0]_b1 ,\d[0]_b0 ;
output \o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,\o[28]_b0 ,\o[27]_b1 ,
		\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,\o[23]_b1 ,\o[23]_b0 ,
		\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,\o[19]_b0 ,\o[18]_b1 ,
		\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,\o[14]_b1 ,\o[14]_b0 ,
		\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,\o[10]_b0 ,\o[9]_b1 ,
		\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,\o[5]_b1 ,\o[5]_b0 ,
		\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,\o[1]_b0 ,\o[0]_b1 ,
		\o[0]_b0 ;

wire \97_ZERO_b1 , \97_ZERO_b0 , \98_ONE_b1 , \98_ONE_b0 , \99_b1 , \99_b0 , \100_b1 , \100_b0 , \101_b1 , \101_b0 , 
		\102_b1 , \102_b0 , \103_b1 , \103_b0 , \104_b1 , \104_b0 , \105_b1 , \105_b0 , \106_b1 , \106_b0 , 
		\107_b1 , \107_b0 , \108_b1 , \108_b0 , \109_b1 , \109_b0 , \110_b1 , \110_b0 , \111_b1 , \111_b0 , 
		\112_b1 , \112_b0 , \113_b1 , \113_b0 , \114_b1 , \114_b0 , \115_b1 , \115_b0 , \116_b1 , \116_b0 , 
		\117_b1 , \117_b0 , \118_b1 , \118_b0 , \119_b1 , \119_b0 , \120_b1 , \120_b0 , \121_b1 , \121_b0 , 
		\122_b1 , \122_b0 , \123_b1 , \123_b0 , \124_b1 , \124_b0 , \125_b1 , \125_b0 , \126_b1 , \126_b0 , 
		\127_b1 , \127_b0 , \128_b1 , \128_b0 , \129_b1 , \129_b0 , \130_b1 , \130_b0 , \131_b1 , \131_b0 , 
		\132_b1 , \132_b0 , \133_b1 , \133_b0 , \134_b1 , \134_b0 , \135_b1 , \135_b0 , \136_b1 , \136_b0 , 
		\137_b1 , \137_b0 , \138_b1 , \138_b0 , \139_b1 , \139_b0 , \140_b1 , \140_b0 , \141_b1 , \141_b0 , 
		\142_b1 , \142_b0 , \143_b1 , \143_b0 , \144_b1 , \144_b0 , \145_b1 , \145_b0 , \146_b1 , \146_b0 , 
		\147_b1 , \147_b0 , \148_b1 , \148_b0 , \149_b1 , \149_b0 , \150_b1 , \150_b0 , \151_b1 , \151_b0 , 
		\152_b1 , \152_b0 , \153_b1 , \153_b0 , \154_b1 , \154_b0 , \155_b1 , \155_b0 , \156_b1 , \156_b0 , 
		\157_b1 , \157_b0 , \158_b1 , \158_b0 , \159_b1 , \159_b0 , \160_b1 , \160_b0 , \161_b1 , \161_b0 , 
		\162_b1 , \162_b0 , \163_b1 , \163_b0 , \164_b1 , \164_b0 , \165_b1 , \165_b0 , \166_b1 , \166_b0 , 
		\167_b1 , \167_b0 , \168_b1 , \168_b0 , \169_b1 , \169_b0 , \170_b1 , \170_b0 , \171_b1 , \171_b0 , 
		\172_b1 , \172_b0 , \173_b1 , \173_b0 , \174_b1 , \174_b0 , \175_b1 , \175_b0 , \176_b1 , \176_b0 , 
		\177_b1 , \177_b0 , \178_b1 , \178_b0 , \179_b1 , \179_b0 , \180_b1 , \180_b0 , \181_b1 , \181_b0 , 
		\182_b1 , \182_b0 , \183_b1 , \183_b0 , \184_b1 , \184_b0 , \185_b1 , \185_b0 , \186_b1 , \186_b0 , 
		\187_b1 , \187_b0 , \188_b1 , \188_b0 , \189_b1 , \189_b0 , \190_b1 , \190_b0 , \191_b1 , \191_b0 , 
		\192_b1 , \192_b0 , \193_b1 , \193_b0 , \194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , 
		\197_b1 , \197_b0 , \198_b1 , \198_b0 , \199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , 
		\202_b1 , \202_b0 , \203_b1 , \203_b0 , \204_b1 , \204_b0 , \205_b1 , \205_b0 , \206_b1 , \206_b0 , 
		\207_b1 , \207_b0 , \208_b1 , \208_b0 , \209_b1 , \209_b0 , \210_b1 , \210_b0 , \211_b1 , \211_b0 , 
		\212_b1 , \212_b0 , \213_b1 , \213_b0 , \214_b1 , \214_b0 , \215_b1 , \215_b0 , \216_b1 , \216_b0 , 
		\217_b1 , \217_b0 , \218_b1 , \218_b0 , \219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , 
		\222_b1 , \222_b0 , \223_b1 , \223_b0 , \224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , 
		\227_b1 , \227_b0 , \228_b1 , \228_b0 , \229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , 
		\232_b1 , \232_b0 , \233_b1 , \233_b0 , \234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , 
		\237_b1 , \237_b0 , \238_b1 , \238_b0 , \239_b1 , \239_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , 
		\242_b1 , \242_b0 , \243_b1 , \243_b0 , \244_b1 , \244_b0 , \245_b1 , \245_b0 , \246_b1 , \246_b0 , 
		\247_b1 , \247_b0 , \248_b1 , \248_b0 , \249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , 
		\252_b1 , \252_b0 , \253_b1 , \253_b0 , \254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , 
		\257_b1 , \257_b0 , \258_b1 , \258_b0 , \259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , 
		\262_b1 , \262_b0 , \263_b1 , \263_b0 , \264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , 
		\267_b1 , \267_b0 , \268_b1 , \268_b0 , \269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , 
		\272_b1 , \272_b0 , \273_b1 , \273_b0 , \274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_b1 , \276_b0 , 
		\277_b1 , \277_b0 , \278_b1 , \278_b0 , \279_b1 , \279_b0 , \280_b1 , \280_b0 , \281_b1 , \281_b0 , 
		\282_b1 , \282_b0 , \283_b1 , \283_b0 , \284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , 
		\287_b1 , \287_b0 , \288_b1 , \288_b0 , \289_b1 , \289_b0 , \290_b1 , \290_b0 , \291_b1 , \291_b0 , 
		\292_b1 , \292_b0 , \293_b1 , \293_b0 , \294_b1 , \294_b0 , \295_b1 , \295_b0 , \296_b1 , \296_b0 , 
		\297_b1 , \297_b0 , \298_b1 , \298_b0 , \299_b1 , \299_b0 , \300_b1 , \300_b0 , \301_b1 , \301_b0 , 
		\302_b1 , \302_b0 , \303_b1 , \303_b0 , \304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , 
		\307_b1 , \307_b0 , \308_b1 , \308_b0 , \309_b1 , \309_b0 , \310_b1 , \310_b0 , \311_b1 , \311_b0 , 
		\312_b1 , \312_b0 , \313_b1 , \313_b0 , \314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_b1 , \316_b0 , 
		\317_b1 , \317_b0 , \318_b1 , \318_b0 , \319_b1 , \319_b0 , \320_b1 , \320_b0 , \321_b1 , \321_b0 , 
		\322_b1 , \322_b0 , \323_b1 , \323_b0 , \324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , 
		\327_b1 , \327_b0 , \328_b1 , \328_b0 , \329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_b1 , \331_b0 , 
		\332_b1 , \332_b0 , \333_b1 , \333_b0 , \334_b1 , \334_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , 
		\337_b1 , \337_b0 , \338_b1 , \338_b0 , \339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_b1 , \341_b0 , 
		\342_b1 , \342_b0 , \343_b1 , \343_b0 , \344_b1 , \344_b0 , \345_b1 , \345_b0 , \346_b1 , \346_b0 , 
		\347_b1 , \347_b0 , \348_b1 , \348_b0 , \349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , 
		\352_b1 , \352_b0 , \353_b1 , \353_b0 , \354_b1 , \354_b0 , \355_b1 , \355_b0 , \356_b1 , \356_b0 , 
		\357_b1 , \357_b0 , \358_b1 , \358_b0 , \359_b1 , \359_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , 
		\362_b1 , \362_b0 , \363_b1 , \363_b0 , \364_b1 , \364_b0 , \365_b1 , \365_b0 , \366_b1 , \366_b0 , 
		\367_b1 , \367_b0 , \368_b1 , \368_b0 , \369_b1 , \369_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , 
		\372_b1 , \372_b0 , \373_b1 , \373_b0 , \374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , 
		\377_b1 , \377_b0 , \378_b1 , \378_b0 , \379_b1 , \379_b0 , \380_b1 , \380_b0 , \381_b1 , \381_b0 , 
		\382_b1 , \382_b0 , \383_b1 , \383_b0 , \384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , 
		\387_b1 , \387_b0 , \388_b1 , \388_b0 , \389_b1 , \389_b0 , \390_b1 , \390_b0 , \391_b1 , \391_b0 , 
		\392_b1 , \392_b0 , \393_b1 , \393_b0 , \394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , 
		\397_b1 , \397_b0 , \398_b1 , \398_b0 , \399_b1 , \399_b0 , \400_b1 , \400_b0 , \401_b1 , \401_b0 , 
		\402_b1 , \402_b0 , \403_b1 , \403_b0 , \404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , 
		\407_b1 , \407_b0 , \408_b1 , \408_b0 , \409_b1 , \409_b0 , \410_b1 , \410_b0 , \411_b1 , \411_b0 , 
		\412_b1 , \412_b0 , \413_b1 , \413_b0 , \414_b1 , \414_b0 , \415_b1 , \415_b0 , \416_b1 , \416_b0 , 
		\417_b1 , \417_b0 , \418_b1 , \418_b0 , \419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , 
		\422_b1 , \422_b0 , \423_b1 , \423_b0 , \424_b1 , \424_b0 , \425_b1 , \425_b0 , \426_b1 , \426_b0 , 
		\427_b1 , \427_b0 , \428_b1 , \428_b0 , \429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , 
		\432_b1 , \432_b0 , \433_b1 , \433_b0 , \434_b1 , \434_b0 , \435_b1 , \435_b0 , \436_b1 , \436_b0 , 
		\437_b1 , \437_b0 , \438_b1 , \438_b0 , \439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , 
		\442_b1 , \442_b0 , \443_b1 , \443_b0 , \444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_b1 , \446_b0 , 
		\447_b1 , \447_b0 , \448_b1 , \448_b0 , \449_b1 , \449_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , 
		\452_b1 , \452_b0 , \453_b1 , \453_b0 , \454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_b1 , \456_b0 , 
		\457_b1 , \457_b0 , \458_b1 , \458_b0 , \459_b1 , \459_b0 , \460_b1 , \460_b0 , \461_b1 , \461_b0 , 
		\462_b1 , \462_b0 , \463_b1 , \463_b0 , \464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , 
		\467_b1 , \467_b0 , \468_b1 , \468_b0 , \469_b1 , \469_b0 , \470_b1 , \470_b0 , \471_b1 , \471_b0 , 
		\472_b1 , \472_b0 , \473_b1 , \473_b0 , \474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , 
		\477_b1 , \477_b0 , \478_b1 , \478_b0 , \479_b1 , \479_b0 , \480_b1 , \480_b0 , \481_b1 , \481_b0 , 
		\482_b1 , \482_b0 , \483_b1 , \483_b0 , \484_b1 , \484_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , 
		\487_b1 , \487_b0 , \488_b1 , \488_b0 , \489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , 
		\492_b1 , \492_b0 , \493_b1 , \493_b0 , \494_b1 , \494_b0 , \495_b1 , \495_b0 , \496_b1 , \496_b0 , 
		\497_b1 , \497_b0 , \498_b1 , \498_b0 , \499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , 
		\502_b1 , \502_b0 , \503_b1 , \503_b0 , \504_b1 , \504_b0 , \505_b1 , \505_b0 , \506_b1 , \506_b0 , 
		\507_b1 , \507_b0 , \508_b1 , \508_b0 , \509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , 
		\512_b1 , \512_b0 , \513_b1 , \513_b0 , \514_b1 , \514_b0 , \515_b1 , \515_b0 , \516_b1 , \516_b0 , 
		\517_b1 , \517_b0 , \518_b1 , \518_b0 , \519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , 
		\522_b1 , \522_b0 , \523_b1 , \523_b0 , \524_b1 , \524_b0 , \525_b1 , \525_b0 , \526_b1 , \526_b0 , 
		\527_b1 , \527_b0 , \528_b1 , \528_b0 , \529_b1 , \529_b0 , \530_b1 , \530_b0 , \531_b1 , \531_b0 , 
		\532_b1 , \532_b0 , \533_b1 , \533_b0 , \534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_b1 , \536_b0 , 
		\537_b1 , \537_b0 , \538_b1 , \538_b0 , \539_b1 , \539_b0 , \540_b1 , \540_b0 , \541_b1 , \541_b0 , 
		\542_b1 , \542_b0 , \543_b1 , \543_b0 , \544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , 
		\547_b1 , \547_b0 , \548_b1 , \548_b0 , \549_b1 , \549_b0 , \550_b1 , \550_b0 , \551_b1 , \551_b0 , 
		\552_b1 , \552_b0 , \553_b1 , \553_b0 , \554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , 
		\557_b1 , \557_b0 , \558_b1 , \558_b0 , \559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_b1 , \561_b0 , 
		\562_b1 , \562_b0 , \563_b1 , \563_b0 , \564_b1 , \564_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , 
		\567_b1 , \567_b0 , \568_b1 , \568_b0 , \569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_b1 , \571_b0 , 
		\572_b1 , \572_b0 , \573_b1 , \573_b0 , \574_b1 , \574_b0 , \575_b1 , \575_b0 , \576_b1 , \576_b0 , 
		\577_b1 , \577_b0 , \578_b1 , \578_b0 , \579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , 
		\582_b1 , \582_b0 , \583_b1 , \583_b0 , \584_b1 , \584_b0 , \585_b1 , \585_b0 , \586_b1 , \586_b0 , 
		\587_b1 , \587_b0 , \588_b1 , \588_b0 , \589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , 
		\592_b1 , \592_b0 , \593_b1 , \593_b0 , \594_b1 , \594_b0 , \595_b1 , \595_b0 , \596_b1 , \596_b0 , 
		\597_b1 , \597_b0 , \598_b1 , \598_b0 , \599_b1 , \599_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , 
		\602_b1 , \602_b0 , \603_b1 , \603_b0 , \604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_b1 , \606_b0 , 
		\607_b1 , \607_b0 , \608_b1 , \608_b0 , \609_b1 , \609_b0 , \610_b1 , \610_b0 , \611_b1 , \611_b0 , 
		\612_b1 , \612_b0 , \613_b1 , \613_b0 , \614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , 
		\617_b1 , \617_b0 , \618_b1 , \618_b0 , \619_b1 , \619_b0 , \620_b1 , \620_b0 , \621_b1 , \621_b0 , 
		\622_b1 , \622_b0 , \623_b1 , \623_b0 , \624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , 
		\627_b1 , \627_b0 , \628_b1 , \628_b0 , \629_b1 , \629_b0 , \630_b1 , \630_b0 , \631_b1 , \631_b0 , 
		\632_b1 , \632_b0 , \633_b1 , \633_b0 , \634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , 
		\637_b1 , \637_b0 , \638_b1 , \638_b0 , \639_b1 , \639_b0 , \640_b1 , \640_b0 , \641_b1 , \641_b0 , 
		\642_b1 , \642_b0 , \643_b1 , \643_b0 , \644_b1 , \644_b0 , \645_b1 , \645_b0 , \646_b1 , \646_b0 , 
		\647_b1 , \647_b0 , \648_b1 , \648_b0 , \649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , 
		\652_b1 , \652_b0 , \653_b1 , \653_b0 , \654_b1 , \654_b0 , \655_b1 , \655_b0 , \656_b1 , \656_b0 , 
		\657_b1 , \657_b0 , \658_b1 , \658_b0 , \659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , 
		\662_b1 , \662_b0 , \663_b1 , \663_b0 , \664_b1 , \664_b0 , \665_b1 , \665_b0 , \666_b1 , \666_b0 , 
		\667_b1 , \667_b0 , \668_b1 , \668_b0 , \669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , 
		\672_b1 , \672_b0 , \673_b1 , \673_b0 , \674_b1 , \674_b0 , \675_b1 , \675_b0 , \676_b1 , \676_b0 , 
		\677_b1 , \677_b0 , \678_b1 , \678_b0 , \679_b1 , \679_b0 , \680_b1 , \680_b0 , \681_b1 , \681_b0 , 
		\682_b1 , \682_b0 , \683_b1 , \683_b0 , \684_b1 , \684_b0 , \685_b1 , \685_b0 , \686_b1 , \686_b0 , 
		\687_b1 , \687_b0 , \688_b1 , \688_b0 , \689_b1 , \689_b0 , \690_b1 , \690_b0 , \691_b1 , \691_b0 , 
		\692_b1 , \692_b0 , \693_b1 , \693_b0 , \694_b1 , \694_b0 , \695_b1 , \695_b0 , \696_b1 , \696_b0 , 
		\697_b1 , \697_b0 , \698_b1 , \698_b0 , \699_b1 , \699_b0 , \700_b1 , \700_b0 , \701_b1 , \701_b0 , 
		\702_b1 , \702_b0 , \703_b1 , \703_b0 , \704_b1 , \704_b0 , \705_b1 , \705_b0 , \706_b1 , \706_b0 , 
		\707_b1 , \707_b0 , \708_b1 , \708_b0 , \709_b1 , \709_b0 , \710_b1 , \710_b0 , \711_b1 , \711_b0 , 
		\712_b1 , \712_b0 , \713_b1 , \713_b0 , \714_b1 , \714_b0 , \715_b1 , \715_b0 , \716_b1 , \716_b0 , 
		\717_b1 , \717_b0 , \718_b1 , \718_b0 , \719_b1 , \719_b0 , \720_b1 , \720_b0 , \721_b1 , \721_b0 , 
		\722_b1 , \722_b0 , \723_b1 , \723_b0 , \724_b1 , \724_b0 , \725_b1 , \725_b0 , \726_b1 , \726_b0 , 
		\727_b1 , \727_b0 , \728_b1 , \728_b0 , \729_b1 , \729_b0 , \730_b1 , \730_b0 , \731_b1 , \731_b0 , 
		\732_b1 , \732_b0 , \733_b1 , \733_b0 , \734_b1 , \734_b0 , \735_b1 , \735_b0 , \736_b1 , \736_b0 , 
		\737_b1 , \737_b0 , \738_b1 , \738_b0 , \739_b1 , \739_b0 , \740_b1 , \740_b0 , \741_b1 , \741_b0 , 
		\742_b1 , \742_b0 , \743_b1 , \743_b0 , \744_b1 , \744_b0 , \745_b1 , \745_b0 , \746_b1 , \746_b0 , 
		\747_b1 , \747_b0 , \748_b1 , \748_b0 , \749_b1 , \749_b0 , \750_b1 , \750_b0 , \751_b1 , \751_b0 , 
		\752_b1 , \752_b0 , \753_b1 , \753_b0 , \754_b1 , \754_b0 , \755_b1 , \755_b0 , \756_b1 , \756_b0 , 
		\757_b1 , \757_b0 , \758_b1 , \758_b0 , \759_b1 , \759_b0 , \760_b1 , \760_b0 , \761_b1 , \761_b0 , 
		\762_b1 , \762_b0 , \763_b1 , \763_b0 , \764_b1 , \764_b0 , \765_b1 , \765_b0 , \766_b1 , \766_b0 , 
		\767_b1 , \767_b0 , \768_b1 , \768_b0 , \769_b1 , \769_b0 , \770_b1 , \770_b0 , \771_b1 , \771_b0 , 
		\772_b1 , \772_b0 , \773_b1 , \773_b0 , \774_b1 , \774_b0 , \775_b1 , \775_b0 , \776_b1 , \776_b0 , 
		\777_b1 , \777_b0 , \778_b1 , \778_b0 , \779_b1 , \779_b0 , \780_b1 , \780_b0 , \781_b1 , \781_b0 , 
		\782_b1 , \782_b0 , \783_b1 , \783_b0 , \784_b1 , \784_b0 , \785_b1 , \785_b0 , \786_b1 , \786_b0 , 
		\787_b1 , \787_b0 , \788_b1 , \788_b0 , \789_b1 , \789_b0 , \790_b1 , \790_b0 , \791_b1 , \791_b0 , 
		\792_b1 , \792_b0 , \793_b1 , \793_b0 , \794_b1 , \794_b0 , \795_b1 , \795_b0 , \796_b1 , \796_b0 , 
		\797_b1 , \797_b0 , \798_b1 , \798_b0 , \799_b1 , \799_b0 , \800_b1 , \800_b0 , \801_b1 , \801_b0 , 
		\802_b1 , \802_b0 , \803_b1 , \803_b0 , \804_b1 , \804_b0 , \805_b1 , \805_b0 , \806_b1 , \806_b0 , 
		\807_b1 , \807_b0 , \808_b1 , \808_b0 , \809_b1 , \809_b0 , \810_b1 , \810_b0 , \811_b1 , \811_b0 , 
		\812_b1 , \812_b0 , \813_b1 , \813_b0 , \814_b1 , \814_b0 , \815_b1 , \815_b0 , \816_b1 , \816_b0 , 
		\817_b1 , \817_b0 , \818_b1 , \818_b0 , \819_b1 , \819_b0 , \820_b1 , \820_b0 , \821_b1 , \821_b0 , 
		\822_b1 , \822_b0 , \823_b1 , \823_b0 , \824_b1 , \824_b0 , \825_b1 , \825_b0 , \826_b1 , \826_b0 , 
		\827_b1 , \827_b0 , \828_b1 , \828_b0 , \829_b1 , \829_b0 , \830_b1 , \830_b0 , \831_b1 , \831_b0 , 
		\832_b1 , \832_b0 , \833_b1 , \833_b0 , \834_b1 , \834_b0 , \835_b1 , \835_b0 , \836_b1 , \836_b0 , 
		\837_b1 , \837_b0 , \838_b1 , \838_b0 , \839_b1 , \839_b0 , \840_b1 , \840_b0 , \841_b1 , \841_b0 , 
		\842_b1 , \842_b0 , \843_b1 , \843_b0 , \844_b1 , \844_b0 , \845_b1 , \845_b0 , \846_b1 , \846_b0 , 
		\847_b1 , \847_b0 , \848_b1 , \848_b0 , \849_b1 , \849_b0 , \850_b1 , \850_b0 , \851_b1 , \851_b0 , 
		\852_b1 , \852_b0 , \853_b1 , \853_b0 , \854_b1 , \854_b0 , \855_b1 , \855_b0 , \856_b1 , \856_b0 , 
		\857_b1 , \857_b0 , \858_b1 , \858_b0 , \859_b1 , \859_b0 , \860_b1 , \860_b0 , \861_b1 , \861_b0 , 
		\862_b1 , \862_b0 , \863_b1 , \863_b0 , \864_b1 , \864_b0 , \865_b1 , \865_b0 , \866_b1 , \866_b0 , 
		\867_b1 , \867_b0 , \868_b1 , \868_b0 , \869_b1 , \869_b0 , \870_b1 , \870_b0 , \871_b1 , \871_b0 , 
		\872_b1 , \872_b0 , \873_b1 , \873_b0 , \874_b1 , \874_b0 , \875_b1 , \875_b0 , \876_b1 , \876_b0 , 
		\877_b1 , \877_b0 , \878_b1 , \878_b0 , \879_b1 , \879_b0 , \880_b1 , \880_b0 , \881_b1 , \881_b0 , 
		\882_b1 , \882_b0 , \883_b1 , \883_b0 , \884_b1 , \884_b0 , \885_b1 , \885_b0 , \886_b1 , \886_b0 , 
		\887_b1 , \887_b0 , \888_b1 , \888_b0 , \889_b1 , \889_b0 , \890_b1 , \890_b0 , \891_b1 , \891_b0 , 
		\892_b1 , \892_b0 , \893_b1 , \893_b0 , \894_b1 , \894_b0 , \895_b1 , \895_b0 , \896_b1 , \896_b0 , 
		\897_b1 , \897_b0 , \898_b1 , \898_b0 , \899_b1 , \899_b0 , \900_b1 , \900_b0 , \901_b1 , \901_b0 , 
		\902_b1 , \902_b0 , \903_b1 , \903_b0 , \904_b1 , \904_b0 , \905_b1 , \905_b0 , \906_b1 , \906_b0 , 
		\907_b1 , \907_b0 , \908_b1 , \908_b0 , \909_b1 , \909_b0 , \910_b1 , \910_b0 , \911_b1 , \911_b0 , 
		\912_b1 , \912_b0 , \913_b1 , \913_b0 , \914_b1 , \914_b0 , \915_b1 , \915_b0 , \916_b1 , \916_b0 , 
		\917_b1 , \917_b0 , \918_b1 , \918_b0 , \919_b1 , \919_b0 , \920_b1 , \920_b0 , \921_b1 , \921_b0 , 
		\922_b1 , \922_b0 , \923_b1 , \923_b0 , \924_b1 , \924_b0 , \925_b1 , \925_b0 , \926_b1 , \926_b0 , 
		\927_b1 , \927_b0 , \928_b1 , \928_b0 , \929_b1 , \929_b0 , \930_b1 , \930_b0 , \931_b1 , \931_b0 , 
		\932_b1 , \932_b0 , \933_b1 , \933_b0 , \934_b1 , \934_b0 , \935_b1 , \935_b0 , \936_b1 , \936_b0 , 
		\937_b1 , \937_b0 , \938_b1 , \938_b0 , \939_b1 , \939_b0 , \940_b1 , \940_b0 , \941_b1 , \941_b0 , 
		\942_b1 , \942_b0 , \943_b1 , \943_b0 , \944_b1 , \944_b0 , \945_b1 , \945_b0 , \946_b1 , \946_b0 , 
		\947_b1 , \947_b0 , \948_b1 , \948_b0 , \949_b1 , \949_b0 , \950_b1 , \950_b0 , \951_b1 , \951_b0 , 
		\952_b1 , \952_b0 , \953_b1 , \953_b0 , \954_b1 , \954_b0 , \955_b1 , \955_b0 , \956_b1 , \956_b0 , 
		\957_b1 , \957_b0 , \958_b1 , \958_b0 , \959_b1 , \959_b0 , \960_b1 , \960_b0 , \961_b1 , \961_b0 , 
		\962_b1 , \962_b0 , \963_b1 , \963_b0 , \964_b1 , \964_b0 , \965_b1 , \965_b0 , \966_b1 , \966_b0 , 
		\967_b1 , \967_b0 , \968_b1 , \968_b0 , \969_b1 , \969_b0 , \970_b1 , \970_b0 , \971_b1 , \971_b0 , 
		\972_b1 , \972_b0 , \973_b1 , \973_b0 , \974_b1 , \974_b0 , \975_b1 , \975_b0 , \976_b1 , \976_b0 , 
		\977_b1 , \977_b0 , \978_b1 , \978_b0 , \979_b1 , \979_b0 , \980_b1 , \980_b0 , \981_b1 , \981_b0 , 
		\982_b1 , \982_b0 , \983_b1 , \983_b0 , \984_b1 , \984_b0 , \985_b1 , \985_b0 , \986_b1 , \986_b0 , 
		\987_b1 , \987_b0 , \988_b1 , \988_b0 , \989_b1 , \989_b0 , \990_b1 , \990_b0 , \991_b1 , \991_b0 , 
		\992_b1 , \992_b0 , \993_b1 , \993_b0 , \994_b1 , \994_b0 , \995_b1 , \995_b0 , \996_b1 , \996_b0 , 
		\997_b1 , \997_b0 , \998_b1 , \998_b0 , \999_b1 , \999_b0 , \1000_b1 , \1000_b0 , \1001_b1 , \1001_b0 , 
		\1002_b1 , \1002_b0 , \1003_b1 , \1003_b0 , \1004_b1 , \1004_b0 , \1005_b1 , \1005_b0 , \1006_b1 , \1006_b0 , 
		\1007_b1 , \1007_b0 , \1008_b1 , \1008_b0 , \1009_b1 , \1009_b0 , \1010_b1 , \1010_b0 , \1011_b1 , \1011_b0 , 
		\1012_b1 , \1012_b0 , \1013_b1 , \1013_b0 , \1014_b1 , \1014_b0 , \1015_b1 , \1015_b0 , \1016_b1 , \1016_b0 , 
		\1017_b1 , \1017_b0 , \1018_b1 , \1018_b0 , \1019_b1 , \1019_b0 , \1020_b1 , \1020_b0 , \1021_b1 , \1021_b0 , 
		\1022_b1 , \1022_b0 , \1023_b1 , \1023_b0 , \1024_b1 , \1024_b0 , \1025_b1 , \1025_b0 , \1026_b1 , \1026_b0 , 
		\1027_b1 , \1027_b0 , \1028_b1 , \1028_b0 , \1029_b1 , \1029_b0 , \1030_b1 , \1030_b0 , \1031_b1 , \1031_b0 , 
		\1032_b1 , \1032_b0 , \1033_b1 , \1033_b0 , \1034_b1 , \1034_b0 , \1035_b1 , \1035_b0 , \1036_b1 , \1036_b0 , 
		\1037_b1 , \1037_b0 , \1038_b1 , \1038_b0 , \1039_b1 , \1039_b0 , \1040_b1 , \1040_b0 , \1041_b1 , \1041_b0 , 
		\1042_b1 , \1042_b0 , \1043_b1 , \1043_b0 , \1044_b1 , \1044_b0 , \1045_b1 , \1045_b0 , \1046_b1 , \1046_b0 , 
		\1047_b1 , \1047_b0 , \1048_b1 , \1048_b0 , \1049_b1 , \1049_b0 , \1050_b1 , \1050_b0 , \1051_b1 , \1051_b0 , 
		\1052_b1 , \1052_b0 , \1053_b1 , \1053_b0 , \1054_b1 , \1054_b0 , \1055_b1 , \1055_b0 , \1056_b1 , \1056_b0 , 
		\1057_b1 , \1057_b0 , \1058_b1 , \1058_b0 , \1059_b1 , \1059_b0 , \1060_b1 , \1060_b0 , \1061_b1 , \1061_b0 , 
		\1062_b1 , \1062_b0 , \1063_b1 , \1063_b0 , \1064_b1 , \1064_b0 , \1065_b1 , \1065_b0 , \1066_b1 , \1066_b0 , 
		\1067_b1 , \1067_b0 , \1068_b1 , \1068_b0 , \1069_b1 , \1069_b0 , \1070_b1 , \1070_b0 , \1071_b1 , \1071_b0 , 
		\1072_b1 , \1072_b0 , \1073_b1 , \1073_b0 , \1074_b1 , \1074_b0 , \1075_b1 , \1075_b0 , \1076_b1 , \1076_b0 , 
		\1077_b1 , \1077_b0 , \1078_b1 , \1078_b0 , \1079_b1 , \1079_b0 , \1080_b1 , \1080_b0 , \1081_b1 , \1081_b0 , 
		\1082_b1 , \1082_b0 , \1083_b1 , \1083_b0 , \1084_b1 , \1084_b0 , \1085_b1 , \1085_b0 , \1086_b1 , \1086_b0 , 
		\1087_b1 , \1087_b0 , \1088_b1 , \1088_b0 , \1089_b1 , \1089_b0 , \1090_b1 , \1090_b0 , \1091_b1 , \1091_b0 , 
		\1092_b1 , \1092_b0 , \1093_b1 , \1093_b0 , \1094_b1 , \1094_b0 , \1095_b1 , \1095_b0 , \1096_b1 , \1096_b0 , 
		\1097_b1 , \1097_b0 , \1098_b1 , \1098_b0 , \1099_b1 , \1099_b0 , \1100_b1 , \1100_b0 , \1101_b1 , \1101_b0 , 
		\1102_b1 , \1102_b0 , \1103_b1 , \1103_b0 , \1104_b1 , \1104_b0 , \1105_b1 , \1105_b0 , \1106_b1 , \1106_b0 , 
		\1107_b1 , \1107_b0 , \1108_b1 , \1108_b0 , \1109_b1 , \1109_b0 , \1110_b1 , \1110_b0 , \1111_b1 , \1111_b0 , 
		\1112_b1 , \1112_b0 , \1113_b1 , \1113_b0 , \1114_b1 , \1114_b0 , \1115_b1 , \1115_b0 , \1116_b1 , \1116_b0 , 
		\1117_b1 , \1117_b0 , \1118_b1 , \1118_b0 , \1119_b1 , \1119_b0 , \1120_b1 , \1120_b0 , \1121_b1 , \1121_b0 , 
		\1122_b1 , \1122_b0 , \1123_b1 , \1123_b0 , \1124_b1 , \1124_b0 , \1125_b1 , \1125_b0 , \1126_b1 , \1126_b0 , 
		\1127_b1 , \1127_b0 , \1128_b1 , \1128_b0 , \1129_b1 , \1129_b0 , \1130_b1 , \1130_b0 , \1131_b1 , \1131_b0 , 
		\1132_b1 , \1132_b0 , \1133_b1 , \1133_b0 , \1134_b1 , \1134_b0 , \1135_b1 , \1135_b0 , \1136_b1 , \1136_b0 , 
		\1137_b1 , \1137_b0 , \1138_b1 , \1138_b0 , \1139_b1 , \1139_b0 , \1140_b1 , \1140_b0 , \1141_b1 , \1141_b0 , 
		\1142_b1 , \1142_b0 , \1143_b1 , \1143_b0 , \1144_b1 , \1144_b0 , \1145_b1 , \1145_b0 , \1146_b1 , \1146_b0 , 
		\1147_b1 , \1147_b0 , \1148_b1 , \1148_b0 , \1149_b1 , \1149_b0 , \1150_b1 , \1150_b0 , \1151_b1 , \1151_b0 , 
		\1152_b1 , \1152_b0 , \1153_b1 , \1153_b0 , \1154_b1 , \1154_b0 , \1155_b1 , \1155_b0 , \1156_b1 , \1156_b0 , 
		\1157_b1 , \1157_b0 , \1158_b1 , \1158_b0 , \1159_b1 , \1159_b0 , \1160_b1 , \1160_b0 , \1161_b1 , \1161_b0 , 
		\1162_b1 , \1162_b0 , \1163_b1 , \1163_b0 , \1164_b1 , \1164_b0 , \1165_b1 , \1165_b0 , \1166_b1 , \1166_b0 , 
		\1167_b1 , \1167_b0 , \1168_b1 , \1168_b0 , \1169_b1 , \1169_b0 , \1170_b1 , \1170_b0 , \1171_b1 , \1171_b0 , 
		\1172_b1 , \1172_b0 , \1173_b1 , \1173_b0 , \1174_b1 , \1174_b0 , \1175_b1 , \1175_b0 , \1176_b1 , \1176_b0 , 
		\1177_b1 , \1177_b0 , \1178_b1 , \1178_b0 , \1179_b1 , \1179_b0 , \1180_b1 , \1180_b0 , \1181_b1 , \1181_b0 , 
		\1182_b1 , \1182_b0 , \1183_b1 , \1183_b0 , \1184_b1 , \1184_b0 , \1185_b1 , \1185_b0 , \1186_b1 , \1186_b0 , 
		\1187_b1 , \1187_b0 , \1188_b1 , \1188_b0 , \1189_b1 , \1189_b0 , \1190_b1 , \1190_b0 , \1191_b1 , \1191_b0 , 
		\1192_b1 , \1192_b0 , \1193_b1 , \1193_b0 , \1194_b1 , \1194_b0 , \1195_b1 , \1195_b0 , \1196_b1 , \1196_b0 , 
		\1197_b1 , \1197_b0 , \1198_b1 , \1198_b0 , \1199_b1 , \1199_b0 , \1200_b1 , \1200_b0 , \1201_b1 , \1201_b0 , 
		\1202_b1 , \1202_b0 , \1203_b1 , \1203_b0 , \1204_b1 , \1204_b0 , \1205_b1 , \1205_b0 , \1206_b1 , \1206_b0 , 
		\1207_b1 , \1207_b0 , \1208_b1 , \1208_b0 , \1209_b1 , \1209_b0 , \1210_b1 , \1210_b0 , \1211_b1 , \1211_b0 , 
		\1212_b1 , \1212_b0 , \1213_b1 , \1213_b0 , \1214_b1 , \1214_b0 , \1215_b1 , \1215_b0 , \1216_b1 , \1216_b0 , 
		\1217_b1 , \1217_b0 , \1218_b1 , \1218_b0 , \1219_b1 , \1219_b0 , \1220_b1 , \1220_b0 , \1221_b1 , \1221_b0 , 
		\1222_b1 , \1222_b0 , \1223_b1 , \1223_b0 , \1224_b1 , \1224_b0 , \1225_b1 , \1225_b0 , \1226_b1 , \1226_b0 , 
		\1227_b1 , \1227_b0 , \1228_b1 , \1228_b0 , \1229_b1 , \1229_b0 , \1230_b1 , \1230_b0 , \1231_b1 , \1231_b0 , 
		\1232_b1 , \1232_b0 , \1233_b1 , \1233_b0 , \1234_b1 , \1234_b0 , \1235_b1 , \1235_b0 , \1236_b1 , \1236_b0 , 
		\1237_b1 , \1237_b0 , \1238_b1 , \1238_b0 , \1239_b1 , \1239_b0 , \1240_b1 , \1240_b0 , \1241_b1 , \1241_b0 , 
		\1242_b1 , \1242_b0 , \1243_b1 , \1243_b0 , \1244_b1 , \1244_b0 , \1245_b1 , \1245_b0 , \1246_b1 , \1246_b0 , 
		\1247_b1 , \1247_b0 , \1248_b1 , \1248_b0 , \1249_b1 , \1249_b0 , \1250_b1 , \1250_b0 , \1251_b1 , \1251_b0 , 
		\1252_b1 , \1252_b0 , \1253_b1 , \1253_b0 , \1254_b1 , \1254_b0 , \1255_b1 , \1255_b0 , \1256_b1 , \1256_b0 , 
		\1257_b1 , \1257_b0 , \1258_b1 , \1258_b0 , \1259_b1 , \1259_b0 , \1260_b1 , \1260_b0 , \1261_b1 , \1261_b0 , 
		\1262_b1 , \1262_b0 , \1263_b1 , \1263_b0 , \1264_b1 , \1264_b0 , \1265_b1 , \1265_b0 , \1266_b1 , \1266_b0 , 
		\1267_b1 , \1267_b0 , \1268_b1 , \1268_b0 , \1269_b1 , \1269_b0 , \1270_b1 , \1270_b0 , \1271_b1 , \1271_b0 , 
		\1272_b1 , \1272_b0 , \1273_b1 , \1273_b0 , \1274_b1 , \1274_b0 , \1275_b1 , \1275_b0 , \1276_b1 , \1276_b0 , 
		\1277_b1 , \1277_b0 , \1278_b1 , \1278_b0 , \1279_b1 , \1279_b0 , \1280_b1 , \1280_b0 , \1281_b1 , \1281_b0 , 
		\1282_b1 , \1282_b0 , \1283_b1 , \1283_b0 , \1284_b1 , \1284_b0 , \1285_b1 , \1285_b0 , \1286_b1 , \1286_b0 , 
		\1287_b1 , \1287_b0 , \1288_b1 , \1288_b0 , \1289_b1 , \1289_b0 , \1290_b1 , \1290_b0 , \1291_b1 , \1291_b0 , 
		\1292_b1 , \1292_b0 , \1293_b1 , \1293_b0 , \1294_b1 , \1294_b0 , \1295_b1 , \1295_b0 , \1296_b1 , \1296_b0 , 
		\1297_b1 , \1297_b0 , \1298_b1 , \1298_b0 , \1299_b1 , \1299_b0 , \1300_b1 , \1300_b0 , \1301_b1 , \1301_b0 , 
		\1302_b1 , \1302_b0 , \1303_b1 , \1303_b0 , \1304_b1 , \1304_b0 , \1305_b1 , \1305_b0 , \1306_b1 , \1306_b0 , 
		\1307_b1 , \1307_b0 , \1308_b1 , \1308_b0 , \1309_b1 , \1309_b0 , \1310_b1 , \1310_b0 , \1311_b1 , \1311_b0 , 
		\1312_b1 , \1312_b0 , \1313_b1 , \1313_b0 , \1314_b1 , \1314_b0 , \1315_b1 , \1315_b0 , \1316_b1 , \1316_b0 , 
		\1317_b1 , \1317_b0 , \1318_b1 , \1318_b0 , \1319_b1 , \1319_b0 , \1320_b1 , \1320_b0 , \1321_b1 , \1321_b0 , 
		\1322_b1 , \1322_b0 , \1323_b1 , \1323_b0 , \1324_b1 , \1324_b0 , \1325_b1 , \1325_b0 , \1326_b1 , \1326_b0 , 
		\1327_b1 , \1327_b0 , \1328_b1 , \1328_b0 , \1329_b1 , \1329_b0 , \1330_b1 , \1330_b0 , \1331_b1 , \1331_b0 , 
		\1332_b1 , \1332_b0 , \1333_b1 , \1333_b0 , \1334_b1 , \1334_b0 , \1335_b1 , \1335_b0 , \1336_b1 , \1336_b0 , 
		\1337_b1 , \1337_b0 , \1338_b1 , \1338_b0 , \1339_b1 , \1339_b0 , \1340_b1 , \1340_b0 , \1341_b1 , \1341_b0 , 
		\1342_b1 , \1342_b0 , \1343_b1 , \1343_b0 , \1344_b1 , \1344_b0 , \1345_b1 , \1345_b0 , \1346_b1 , \1346_b0 , 
		\1347_b1 , \1347_b0 , \1348_b1 , \1348_b0 , \1349_b1 , \1349_b0 , \1350_b1 , \1350_b0 , \1351_b1 , \1351_b0 , 
		\1352_b1 , \1352_b0 , \1353_b1 , \1353_b0 , \1354_b1 , \1354_b0 , \1355_b1 , \1355_b0 , \1356_b1 , \1356_b0 , 
		\1357_b1 , \1357_b0 , \1358_b1 , \1358_b0 , \1359_b1 , \1359_b0 , \1360_b1 , \1360_b0 , \1361_b1 , \1361_b0 , 
		\1362_b1 , \1362_b0 , \1363_b1 , \1363_b0 , \1364_b1 , \1364_b0 , \1365_b1 , \1365_b0 , \1366_b1 , \1366_b0 , 
		\1367_b1 , \1367_b0 , \1368_b1 , \1368_b0 , \1369_b1 , \1369_b0 , \1370_b1 , \1370_b0 , \1371_b1 , \1371_b0 , 
		\1372_b1 , \1372_b0 , \1373_b1 , \1373_b0 , \1374_b1 , \1374_b0 , \1375_b1 , \1375_b0 , \1376_b1 , \1376_b0 , 
		\1377_b1 , \1377_b0 , \1378_b1 , \1378_b0 , \1379_b1 , \1379_b0 , \1380_b1 , \1380_b0 , \1381_b1 , \1381_b0 , 
		\1382_b1 , \1382_b0 , \1383_b1 , \1383_b0 , \1384_b1 , \1384_b0 , \1385_b1 , \1385_b0 , \1386_b1 , \1386_b0 , 
		\1387_b1 , \1387_b0 , \1388_b1 , \1388_b0 , \1389_b1 , \1389_b0 , \1390_b1 , \1390_b0 , \1391_b1 , \1391_b0 , 
		\1392_b1 , \1392_b0 , \1393_b1 , \1393_b0 , \1394_b1 , \1394_b0 , \1395_b1 , \1395_b0 , \1396_b1 , \1396_b0 , 
		\1397_b1 , \1397_b0 , \1398_b1 , \1398_b0 , \1399_b1 , \1399_b0 , \1400_b1 , \1400_b0 , \1401_b1 , \1401_b0 , 
		\1402_b1 , \1402_b0 , \1403_b1 , \1403_b0 , \1404_b1 , \1404_b0 , \1405_b1 , \1405_b0 , \1406_b1 , \1406_b0 , 
		\1407_b1 , \1407_b0 , \1408_b1 , \1408_b0 , \1409_b1 , \1409_b0 , \1410_b1 , \1410_b0 , \1411_b1 , \1411_b0 , 
		\1412_b1 , \1412_b0 , \1413_b1 , \1413_b0 , \1414_b1 , \1414_b0 , \1415_b1 , \1415_b0 , \1416_b1 , \1416_b0 , 
		\1417_b1 , \1417_b0 , \1418_b1 , \1418_b0 , \1419_b1 , \1419_b0 , \1420_b1 , \1420_b0 , \1421_b1 , \1421_b0 , 
		\1422_b1 , \1422_b0 , \1423_b1 , \1423_b0 , \1424_b1 , \1424_b0 , \1425_b1 , \1425_b0 , \1426_b1 , \1426_b0 , 
		\1427_b1 , \1427_b0 , \1428_b1 , \1428_b0 , \1429_b1 , \1429_b0 , \1430_b1 , \1430_b0 , \1431_b1 , \1431_b0 , 
		\1432_b1 , \1432_b0 , \1433_b1 , \1433_b0 , \1434_b1 , \1434_b0 , \1435_b1 , \1435_b0 , \1436_b1 , \1436_b0 , 
		\1437_b1 , \1437_b0 , \1438_b1 , \1438_b0 , \1439_b1 , \1439_b0 , \1440_b1 , \1440_b0 , \1441_b1 , \1441_b0 , 
		\1442_b1 , \1442_b0 , \1443_b1 , \1443_b0 , \1444_b1 , \1444_b0 , \1445_b1 , \1445_b0 , \1446_b1 , \1446_b0 , 
		\1447_b1 , \1447_b0 , \1448_b1 , \1448_b0 , \1449_b1 , \1449_b0 , \1450_b1 , \1450_b0 , \1451_b1 , \1451_b0 , 
		\1452_b1 , \1452_b0 , \1453_b1 , \1453_b0 , \1454_b1 , \1454_b0 , \1455_b1 , \1455_b0 , \1456_b1 , \1456_b0 , 
		\1457_b1 , \1457_b0 , \1458_b1 , \1458_b0 , \1459_b1 , \1459_b0 , \1460_b1 , \1460_b0 , \1461_b1 , \1461_b0 , 
		\1462_b1 , \1462_b0 , \1463_b1 , \1463_b0 , \1464_b1 , \1464_b0 , \1465_b1 , \1465_b0 , \1466_b1 , \1466_b0 , 
		\1467_b1 , \1467_b0 , \1468_b1 , \1468_b0 , \1469_b1 , \1469_b0 , \1470_b1 , \1470_b0 , \1471_b1 , \1471_b0 , 
		\1472_b1 , \1472_b0 , \1473_b1 , \1473_b0 , \1474_b1 , \1474_b0 , \1475_b1 , \1475_b0 , \1476_b1 , \1476_b0 , 
		\1477_b1 , \1477_b0 , \1478_b1 , \1478_b0 , \1479_b1 , \1479_b0 , \1480_b1 , \1480_b0 , \1481_b1 , \1481_b0 , 
		\1482_b1 , \1482_b0 , \1483_b1 , \1483_b0 , \1484_b1 , \1484_b0 , \1485_b1 , \1485_b0 , \1486_b1 , \1486_b0 , 
		\1487_b1 , \1487_b0 , \1488_b1 , \1488_b0 , \1489_b1 , \1489_b0 , \1490_b1 , \1490_b0 , \1491_b1 , \1491_b0 , 
		\1492_b1 , \1492_b0 , \1493_b1 , \1493_b0 , \1494_b1 , \1494_b0 , \1495_b1 , \1495_b0 , \1496_b1 , \1496_b0 , 
		\1497_b1 , \1497_b0 , \1498_b1 , \1498_b0 , \1499_b1 , \1499_b0 , \1500_b1 , \1500_b0 , \1501_b1 , \1501_b0 , 
		\1502_b1 , \1502_b0 , \1503_b1 , \1503_b0 , \1504_b1 , \1504_b0 , \1505_b1 , \1505_b0 , \1506_b1 , \1506_b0 , 
		\1507_b1 , \1507_b0 , \1508_b1 , \1508_b0 , \1509_b1 , \1509_b0 , \1510_b1 , \1510_b0 , \1511_b1 , \1511_b0 , 
		\1512_b1 , \1512_b0 , \1513_b1 , \1513_b0 , \1514_b1 , \1514_b0 , \1515_b1 , \1515_b0 , \1516_b1 , \1516_b0 , 
		\1517_b1 , \1517_b0 , \1518_b1 , \1518_b0 , \1519_b1 , \1519_b0 , \1520_b1 , \1520_b0 , \1521_b1 , \1521_b0 , 
		\1522_b1 , \1522_b0 , \1523_b1 , \1523_b0 , \1524_b1 , \1524_b0 , \1525_b1 , \1525_b0 , \1526_b1 , \1526_b0 , 
		\1527_b1 , \1527_b0 , \1528_b1 , \1528_b0 , \1529_b1 , \1529_b0 , \1530_b1 , \1530_b0 , \1531_b1 , \1531_b0 , 
		\1532_b1 , \1532_b0 , \1533_b1 , \1533_b0 , \1534_b1 , \1534_b0 , \1535_b1 , \1535_b0 , \1536_b1 , \1536_b0 , 
		\1537_b1 , \1537_b0 , \1538_b1 , \1538_b0 , \1539_b1 , \1539_b0 , \1540_b1 , \1540_b0 , \1541_b1 , \1541_b0 , 
		\1542_b1 , \1542_b0 , \1543_b1 , \1543_b0 , \1544_b1 , \1544_b0 , \1545_b1 , \1545_b0 , \1546_b1 , \1546_b0 , 
		\1547_b1 , \1547_b0 , \1548_b1 , \1548_b0 , \1549_b1 , \1549_b0 , \1550_b1 , \1550_b0 , \1551_b1 , \1551_b0 , 
		\1552_b1 , \1552_b0 , \1553_b1 , \1553_b0 , \1554_b1 , \1554_b0 , \1555_b1 , \1555_b0 , \1556_b1 , \1556_b0 , 
		\1557_b1 , \1557_b0 , \1558_b1 , \1558_b0 , \1559_b1 , \1559_b0 , \1560_b1 , \1560_b0 , \1561_b1 , \1561_b0 , 
		\1562_b1 , \1562_b0 , \1563_b1 , \1563_b0 , \1564_b1 , \1564_b0 , \1565_b1 , \1565_b0 , \1566_b1 , \1566_b0 , 
		\1567_b1 , \1567_b0 , \1568_b1 , \1568_b0 , \1569_b1 , \1569_b0 , \1570_b1 , \1570_b0 , \1571_b1 , \1571_b0 , 
		\1572_b1 , \1572_b0 , \1573_b1 , \1573_b0 , \1574_b1 , \1574_b0 , \1575_b1 , \1575_b0 , \1576_b1 , \1576_b0 , 
		\1577_b1 , \1577_b0 , \1578_b1 , \1578_b0 , \1579_b1 , \1579_b0 , \1580_b1 , \1580_b0 , \1581_b1 , \1581_b0 , 
		\1582_b1 , \1582_b0 , \1583_b1 , \1583_b0 , \1584_b1 , \1584_b0 , \1585_b1 , \1585_b0 , \1586_b1 , \1586_b0 , 
		\1587_b1 , \1587_b0 , \1588_b1 , \1588_b0 , \1589_b1 , \1589_b0 , \1590_b1 , \1590_b0 , \1591_b1 , \1591_b0 , 
		\1592_b1 , \1592_b0 , \1593_b1 , \1593_b0 , \1594_b1 , \1594_b0 , \1595_b1 , \1595_b0 , \1596_b1 , \1596_b0 , 
		\1597_b1 , \1597_b0 , \1598_b1 , \1598_b0 , \1599_b1 , \1599_b0 , \1600_b1 , \1600_b0 , \1601_b1 , \1601_b0 , 
		\1602_b1 , \1602_b0 , \1603_b1 , \1603_b0 , \1604_b1 , \1604_b0 , \1605_b1 , \1605_b0 , \1606_b1 , \1606_b0 , 
		\1607_b1 , \1607_b0 , \1608_b1 , \1608_b0 , \1609_b1 , \1609_b0 , \1610_b1 , \1610_b0 , \1611_b1 , \1611_b0 , 
		\1612_b1 , \1612_b0 , \1613_b1 , \1613_b0 , \1614_b1 , \1614_b0 , \1615_b1 , \1615_b0 , \1616_b1 , \1616_b0 , 
		\1617_b1 , \1617_b0 , \1618_b1 , \1618_b0 , \1619_b1 , \1619_b0 , \1620_b1 , \1620_b0 , \1621_b1 , \1621_b0 , 
		\1622_b1 , \1622_b0 , \1623_b1 , \1623_b0 , \1624_b1 , \1624_b0 , \1625_b1 , \1625_b0 , \1626_b1 , \1626_b0 , 
		\1627_b1 , \1627_b0 , \1628_b1 , \1628_b0 , \1629_b1 , \1629_b0 , \1630_b1 , \1630_b0 , \1631_b1 , \1631_b0 , 
		\1632_b1 , \1632_b0 , \1633_b1 , \1633_b0 , \1634_b1 , \1634_b0 , \1635_b1 , \1635_b0 , \1636_b1 , \1636_b0 , 
		\1637_b1 , \1637_b0 , \1638_b1 , \1638_b0 , \1639_b1 , \1639_b0 , \1640_b1 , \1640_b0 , \1641_b1 , \1641_b0 , 
		\1642_b1 , \1642_b0 , \1643_b1 , \1643_b0 , \1644_b1 , \1644_b0 , \1645_b1 , \1645_b0 , \1646_b1 , \1646_b0 , 
		\1647_b1 , \1647_b0 , \1648_b1 , \1648_b0 , \1649_b1 , \1649_b0 , \1650_b1 , \1650_b0 , \1651_b1 , \1651_b0 , 
		\1652_b1 , \1652_b0 , \1653_b1 , \1653_b0 , \1654_b1 , \1654_b0 , \1655_b1 , \1655_b0 , \1656_b1 , \1656_b0 , 
		\1657_b1 , \1657_b0 , \1658_b1 , \1658_b0 , \1659_b1 , \1659_b0 , \1660_b1 , \1660_b0 , \1661_b1 , \1661_b0 , 
		\1662_b1 , \1662_b0 , \1663_b1 , \1663_b0 , \1664_b1 , \1664_b0 , \1665_b1 , \1665_b0 , \1666_b1 , \1666_b0 , 
		\1667_b1 , \1667_b0 , \1668_b1 , \1668_b0 , \1669_b1 , \1669_b0 , \1670_b1 , \1670_b0 , \1671_b1 , \1671_b0 , 
		\1672_b1 , \1672_b0 , \1673_b1 , \1673_b0 , \1674_b1 , \1674_b0 , \1675_b1 , \1675_b0 , \1676_b1 , \1676_b0 , 
		\1677_b1 , \1677_b0 , \1678_b1 , \1678_b0 , \1679_b1 , \1679_b0 , \1680_b1 , \1680_b0 , \1681_b1 , \1681_b0 , 
		\1682_b1 , \1682_b0 , \1683_b1 , \1683_b0 , \1684_b1 , \1684_b0 , \1685_b1 , \1685_b0 , \1686_b1 , \1686_b0 , 
		\1687_b1 , \1687_b0 , \1688_b1 , \1688_b0 , \1689_b1 , \1689_b0 , \1690_b1 , \1690_b0 , \1691_b1 , \1691_b0 , 
		\1692_b1 , \1692_b0 , \1693_b1 , \1693_b0 , \1694_b1 , \1694_b0 , \1695_b1 , \1695_b0 , \1696_b1 , \1696_b0 , 
		\1697_b1 , \1697_b0 , \1698_b1 , \1698_b0 , \1699_b1 , \1699_b0 , \1700_b1 , \1700_b0 , \1701_b1 , \1701_b0 , 
		\1702_b1 , \1702_b0 , \1703_b1 , \1703_b0 , \1704_b1 , \1704_b0 , \1705_b1 , \1705_b0 , \1706_b1 , \1706_b0 , 
		\1707_b1 , \1707_b0 , \1708_b1 , \1708_b0 , \1709_b1 , \1709_b0 , \1710_b1 , \1710_b0 , \1711_b1 , \1711_b0 , 
		\1712_b1 , \1712_b0 , \1713_b1 , \1713_b0 , \1714_b1 , \1714_b0 , \1715_b1 , \1715_b0 , \1716_b1 , \1716_b0 , 
		\1717_b1 , \1717_b0 , \1718_b1 , \1718_b0 , \1719_b1 , \1719_b0 , \1720_b1 , \1720_b0 , \1721_b1 , \1721_b0 , 
		\1722_b1 , \1722_b0 , \1723_b1 , \1723_b0 , \1724_b1 , \1724_b0 , \1725_b1 , \1725_b0 , \1726_b1 , \1726_b0 , 
		\1727_b1 , \1727_b0 , \1728_b1 , \1728_b0 , \1729_b1 , \1729_b0 , \1730_b1 , \1730_b0 , \1731_b1 , \1731_b0 , 
		\1732_b1 , \1732_b0 , \1733_b1 , \1733_b0 , \1734_b1 , \1734_b0 , \1735_b1 , \1735_b0 , \1736_b1 , \1736_b0 , 
		\1737_b1 , \1737_b0 , \1738_b1 , \1738_b0 , \1739_b1 , \1739_b0 , \1740_b1 , \1740_b0 , \1741_b1 , \1741_b0 , 
		\1742_b1 , \1742_b0 , \1743_b1 , \1743_b0 , \1744_b1 , \1744_b0 , \1745_b1 , \1745_b0 , \1746_b1 , \1746_b0 , 
		\1747_b1 , \1747_b0 , \1748_b1 , \1748_b0 , \1749_b1 , \1749_b0 , \1750_b1 , \1750_b0 , \1751_b1 , \1751_b0 , 
		\1752_b1 , \1752_b0 , \1753_b1 , \1753_b0 , \1754_b1 , \1754_b0 , \1755_b1 , \1755_b0 , \1756_b1 , \1756_b0 , 
		\1757_b1 , \1757_b0 , \1758_b1 , \1758_b0 , \1759_b1 , \1759_b0 , \1760_b1 , \1760_b0 , \1761_b1 , \1761_b0 , 
		\1762_b1 , \1762_b0 , \1763_b1 , \1763_b0 , \1764_b1 , \1764_b0 , \1765_b1 , \1765_b0 , \1766_b1 , \1766_b0 , 
		\1767_b1 , \1767_b0 , \1768_b1 , \1768_b0 , \1769_b1 , \1769_b0 , \1770_b1 , \1770_b0 , \1771_b1 , \1771_b0 , 
		\1772_b1 , \1772_b0 , \1773_b1 , \1773_b0 , \1774_b1 , \1774_b0 , \1775_b1 , \1775_b0 , \1776_b1 , \1776_b0 , 
		\1777_b1 , \1777_b0 , \1778_b1 , \1778_b0 , \1779_b1 , \1779_b0 , \1780_b1 , \1780_b0 , \1781_b1 , \1781_b0 , 
		\1782_b1 , \1782_b0 , \1783_b1 , \1783_b0 , \1784_b1 , \1784_b0 , \1785_b1 , \1785_b0 , \1786_b1 , \1786_b0 , 
		\1787_b1 , \1787_b0 , \1788_b1 , \1788_b0 , \1789_b1 , \1789_b0 , \1790_b1 , \1790_b0 , \1791_b1 , \1791_b0 , 
		\1792_b1 , \1792_b0 , \1793_b1 , \1793_b0 , \1794_b1 , \1794_b0 , \1795_b1 , \1795_b0 , \1796_b1 , \1796_b0 , 
		\1797_b1 , \1797_b0 , \1798_b1 , \1798_b0 , \1799_b1 , \1799_b0 , \1800_b1 , \1800_b0 , \1801_b1 , \1801_b0 , 
		\1802_b1 , \1802_b0 , \1803_b1 , \1803_b0 , \1804_b1 , \1804_b0 , \1805_b1 , \1805_b0 , \1806_b1 , \1806_b0 , 
		\1807_b1 , \1807_b0 , \1808_b1 , \1808_b0 , \1809_b1 , \1809_b0 , \1810_b1 , \1810_b0 , \1811_b1 , \1811_b0 , 
		\1812_b1 , \1812_b0 , \1813_b1 , \1813_b0 , \1814_b1 , \1814_b0 , \1815_b1 , \1815_b0 , \1816_b1 , \1816_b0 , 
		\1817_b1 , \1817_b0 , \1818_b1 , \1818_b0 , \1819_b1 , \1819_b0 , \1820_b1 , \1820_b0 , \1821_b1 , \1821_b0 , 
		\1822_b1 , \1822_b0 , \1823_b1 , \1823_b0 , \1824_b1 , \1824_b0 , \1825_b1 , \1825_b0 , \1826_b1 , \1826_b0 , 
		\1827_b1 , \1827_b0 , \1828_b1 , \1828_b0 , \1829_b1 , \1829_b0 , \1830_b1 , \1830_b0 , \1831_b1 , \1831_b0 , 
		\1832_b1 , \1832_b0 , \1833_b1 , \1833_b0 , \1834_b1 , \1834_b0 , \1835_b1 , \1835_b0 , \1836_b1 , \1836_b0 , 
		\1837_b1 , \1837_b0 , \1838_b1 , \1838_b0 , \1839_b1 , \1839_b0 , \1840_b1 , \1840_b0 , \1841_b1 , \1841_b0 , 
		\1842_b1 , \1842_b0 , \1843_b1 , \1843_b0 , \1844_b1 , \1844_b0 , \1845_b1 , \1845_b0 , \1846_b1 , \1846_b0 , 
		\1847_b1 , \1847_b0 , \1848_b1 , \1848_b0 , \1849_b1 , \1849_b0 , \1850_b1 , \1850_b0 , \1851_b1 , \1851_b0 , 
		\1852_b1 , \1852_b0 , \1853_b1 , \1853_b0 , \1854_b1 , \1854_b0 , \1855_b1 , \1855_b0 , \1856_b1 , \1856_b0 , 
		\1857_b1 , \1857_b0 , \1858_b1 , \1858_b0 , \1859_b1 , \1859_b0 , \1860_b1 , \1860_b0 , \1861_b1 , \1861_b0 , 
		\1862_b1 , \1862_b0 , \1863_b1 , \1863_b0 , \1864_b1 , \1864_b0 , \1865_b1 , \1865_b0 , \1866_b1 , \1866_b0 , 
		\1867_b1 , \1867_b0 , \1868_b1 , \1868_b0 , \1869_b1 , \1869_b0 , \1870_b1 , \1870_b0 , \1871_b1 , \1871_b0 , 
		\1872_b1 , \1872_b0 , \1873_b1 , \1873_b0 , \1874_b1 , \1874_b0 , \1875_b1 , \1875_b0 , \1876_b1 , \1876_b0 , 
		\1877_b1 , \1877_b0 , \1878_b1 , \1878_b0 , \1879_b1 , \1879_b0 , \1880_b1 , \1880_b0 , \1881_b1 , \1881_b0 , 
		\1882_b1 , \1882_b0 , \1883_b1 , \1883_b0 , \1884_b1 , \1884_b0 , \1885_b1 , \1885_b0 , \1886_b1 , \1886_b0 , 
		\1887_b1 , \1887_b0 , \1888_b1 , \1888_b0 , \1889_b1 , \1889_b0 , \1890_b1 , \1890_b0 , \1891_b1 , \1891_b0 , 
		\1892_b1 , \1892_b0 , \1893_b1 , \1893_b0 , \1894_b1 , \1894_b0 , \1895_b1 , \1895_b0 , \1896_b1 , \1896_b0 , 
		\1897_b1 , \1897_b0 , \1898_b1 , \1898_b0 , \1899_b1 , \1899_b0 , \1900_b1 , \1900_b0 , \1901_b1 , \1901_b0 , 
		\1902_b1 , \1902_b0 , \1903_b1 , \1903_b0 , \1904_b1 , \1904_b0 , \1905_b1 , \1905_b0 , \1906_b1 , \1906_b0 , 
		\1907_b1 , \1907_b0 , \1908_b1 , \1908_b0 , \1909_b1 , \1909_b0 , \1910_b1 , \1910_b0 , \1911_b1 , \1911_b0 , 
		\1912_b1 , \1912_b0 , \1913_b1 , \1913_b0 , \1914_b1 , \1914_b0 , \1915_b1 , \1915_b0 , \1916_b1 , \1916_b0 , 
		\1917_b1 , \1917_b0 , \1918_b1 , \1918_b0 , \1919_b1 , \1919_b0 , \1920_b1 , \1920_b0 , \1921_b1 , \1921_b0 , 
		\1922_b1 , \1922_b0 , \1923_b1 , \1923_b0 , \1924_b1 , \1924_b0 , \1925_b1 , \1925_b0 , \1926_b1 , \1926_b0 , 
		\1927_b1 , \1927_b0 , \1928_b1 , \1928_b0 , \1929_b1 , \1929_b0 , \1930_b1 , \1930_b0 , \1931_b1 , \1931_b0 , 
		\1932_b1 , \1932_b0 , \1933_b1 , \1933_b0 , \1934_b1 , \1934_b0 , \1935_b1 , \1935_b0 , \1936_b1 , \1936_b0 , 
		\1937_b1 , \1937_b0 , \1938_b1 , \1938_b0 , \1939_b1 , \1939_b0 , \1940_b1 , \1940_b0 , \1941_b1 , \1941_b0 , 
		\1942_b1 , \1942_b0 , \1943_b1 , \1943_b0 , \1944_b1 , \1944_b0 , \1945_b1 , \1945_b0 , \1946_b1 , \1946_b0 , 
		\1947_b1 , \1947_b0 , \1948_b1 , \1948_b0 , \1949_b1 , \1949_b0 , \1950_b1 , \1950_b0 , \1951_b1 , \1951_b0 , 
		\1952_b1 , \1952_b0 , \1953_b1 , \1953_b0 , \1954_b1 , \1954_b0 , \1955_b1 , \1955_b0 , \1956_b1 , \1956_b0 , 
		\1957_b1 , \1957_b0 , \1958_b1 , \1958_b0 , \1959_b1 , \1959_b0 , \1960_b1 , \1960_b0 , \1961_b1 , \1961_b0 , 
		\1962_b1 , \1962_b0 , \1963_b1 , \1963_b0 , \1964_b1 , \1964_b0 , \1965_b1 , \1965_b0 , \1966_b1 , \1966_b0 , 
		\1967_b1 , \1967_b0 , \1968_b1 , \1968_b0 , \1969_b1 , \1969_b0 , \1970_b1 , \1970_b0 , \1971_b1 , \1971_b0 , 
		\1972_b1 , \1972_b0 , \1973_b1 , \1973_b0 , \1974_b1 , \1974_b0 , \1975_b1 , \1975_b0 , \1976_b1 , \1976_b0 , 
		\1977_b1 , \1977_b0 , \1978_b1 , \1978_b0 , \1979_b1 , \1979_b0 , \1980_b1 , \1980_b0 , \1981_b1 , \1981_b0 , 
		\1982_b1 , \1982_b0 , \1983_b1 , \1983_b0 , \1984_b1 , \1984_b0 , \1985_b1 , \1985_b0 , \1986_b1 , \1986_b0 , 
		\1987_b1 , \1987_b0 , \1988_b1 , \1988_b0 , \1989_b1 , \1989_b0 , \1990_b1 , \1990_b0 , \1991_b1 , \1991_b0 , 
		\1992_b1 , \1992_b0 , \1993_b1 , \1993_b0 , \1994_b1 , \1994_b0 , \1995_b1 , \1995_b0 , \1996_b1 , \1996_b0 , 
		\1997_b1 , \1997_b0 , \1998_b1 , \1998_b0 , \1999_b1 , \1999_b0 , \2000_b1 , \2000_b0 , \2001_b1 , \2001_b0 , 
		\2002_b1 , \2002_b0 , \2003_b1 , \2003_b0 , \2004_b1 , \2004_b0 , \2005_b1 , \2005_b0 , \2006_b1 , \2006_b0 , 
		\2007_b1 , \2007_b0 , \2008_b1 , \2008_b0 , \2009_b1 , \2009_b0 , \2010_b1 , \2010_b0 , \2011_b1 , \2011_b0 , 
		\2012_b1 , \2012_b0 , \2013_b1 , \2013_b0 , \2014_b1 , \2014_b0 , \2015_b1 , \2015_b0 , \2016_b1 , \2016_b0 , 
		\2017_b1 , \2017_b0 , \2018_b1 , \2018_b0 , \2019_b1 , \2019_b0 , \2020_b1 , \2020_b0 , \2021_b1 , \2021_b0 , 
		\2022_b1 , \2022_b0 , \2023_b1 , \2023_b0 , \2024_b1 , \2024_b0 , \2025_b1 , \2025_b0 , \2026_b1 , \2026_b0 , 
		\2027_b1 , \2027_b0 , \2028_b1 , \2028_b0 , \2029_b1 , \2029_b0 , \2030_b1 , \2030_b0 , \2031_b1 , \2031_b0 , 
		\2032_b1 , \2032_b0 , \2033_b1 , \2033_b0 , \2034_b1 , \2034_b0 , \2035_b1 , \2035_b0 , \2036_b1 , \2036_b0 , 
		\2037_b1 , \2037_b0 , \2038_b1 , \2038_b0 , \2039_b1 , \2039_b0 , \2040_b1 , \2040_b0 , \2041_b1 , \2041_b0 , 
		\2042_b1 , \2042_b0 , \2043_b1 , \2043_b0 , \2044_b1 , \2044_b0 , \2045_b1 , \2045_b0 , \2046_b1 , \2046_b0 , 
		\2047_b1 , \2047_b0 , \2048_b1 , \2048_b0 , \2049_b1 , \2049_b0 , \2050_b1 , \2050_b0 , \2051_b1 , \2051_b0 , 
		\2052_b1 , \2052_b0 , \2053_b1 , \2053_b0 , \2054_b1 , \2054_b0 , \2055_b1 , \2055_b0 , \2056_b1 , \2056_b0 , 
		\2057_b1 , \2057_b0 , \2058_b1 , \2058_b0 , \2059_b1 , \2059_b0 , \2060_b1 , \2060_b0 , \2061_b1 , \2061_b0 , 
		\2062_b1 , \2062_b0 , \2063_b1 , \2063_b0 , \2064_b1 , \2064_b0 , \2065_b1 , \2065_b0 , \2066_b1 , \2066_b0 , 
		\2067_b1 , \2067_b0 , \2068_b1 , \2068_b0 , \2069_b1 , \2069_b0 , \2070_b1 , \2070_b0 , \2071_b1 , \2071_b0 , 
		\2072_b1 , \2072_b0 , \2073_b1 , \2073_b0 , \2074_b1 , \2074_b0 , \2075_b1 , \2075_b0 , \2076_b1 , \2076_b0 , 
		\2077_b1 , \2077_b0 , \2078_b1 , \2078_b0 , \2079_b1 , \2079_b0 , \2080_b1 , \2080_b0 , \2081_b1 , \2081_b0 , 
		\2082_b1 , \2082_b0 , \2083_b1 , \2083_b0 , \2084_b1 , \2084_b0 , \2085_b1 , \2085_b0 , \2086_b1 , \2086_b0 , 
		\2087_b1 , \2087_b0 , \2088_b1 , \2088_b0 , \2089_b1 , \2089_b0 , \2090_b1 , \2090_b0 , \2091_b1 , \2091_b0 , 
		\2092_b1 , \2092_b0 , \2093_b1 , \2093_b0 , \2094_b1 , \2094_b0 , \2095_b1 , \2095_b0 , \2096_b1 , \2096_b0 , 
		\2097_b1 , \2097_b0 , \2098_b1 , \2098_b0 , \2099_b1 , \2099_b0 , \2100_b1 , \2100_b0 , \2101_b1 , \2101_b0 , 
		\2102_b1 , \2102_b0 , \2103_b1 , \2103_b0 , \2104_b1 , \2104_b0 , \2105_b1 , \2105_b0 , \2106_b1 , \2106_b0 , 
		\2107_b1 , \2107_b0 , \2108_b1 , \2108_b0 , \2109_b1 , \2109_b0 , \2110_b1 , \2110_b0 , \2111_b1 , \2111_b0 , 
		\2112_b1 , \2112_b0 , \2113_b1 , \2113_b0 , \2114_b1 , \2114_b0 , \2115_b1 , \2115_b0 , \2116_b1 , \2116_b0 , 
		\2117_b1 , \2117_b0 , \2118_b1 , \2118_b0 , \2119_b1 , \2119_b0 , \2120_b1 , \2120_b0 , \2121_b1 , \2121_b0 , 
		\2122_b1 , \2122_b0 , \2123_b1 , \2123_b0 , \2124_b1 , \2124_b0 , \2125_b1 , \2125_b0 , \2126_b1 , \2126_b0 , 
		\2127_b1 , \2127_b0 , \2128_b1 , \2128_b0 , \2129_b1 , \2129_b0 , \2130_b1 , \2130_b0 , \2131_b1 , \2131_b0 , 
		\2132_b1 , \2132_b0 , \2133_b1 , \2133_b0 , \2134_b1 , \2134_b0 , \2135_b1 , \2135_b0 , \2136_b1 , \2136_b0 , 
		\2137_b1 , \2137_b0 , \2138_b1 , \2138_b0 , \2139_b1 , \2139_b0 , \2140_b1 , \2140_b0 , \2141_b1 , \2141_b0 , 
		\2142_b1 , \2142_b0 , \2143_b1 , \2143_b0 , \2144_b1 , \2144_b0 , \2145_b1 , \2145_b0 , \2146_b1 , \2146_b0 , 
		\2147_b1 , \2147_b0 , \2148_b1 , \2148_b0 , \2149_b1 , \2149_b0 , \2150_b1 , \2150_b0 , \2151_b1 , \2151_b0 , 
		\2152_b1 , \2152_b0 , \2153_b1 , \2153_b0 , \2154_b1 , \2154_b0 , \2155_b1 , \2155_b0 , \2156_b1 , \2156_b0 , 
		\2157_b1 , \2157_b0 , \2158_b1 , \2158_b0 , \2159_b1 , \2159_b0 , \2160_b1 , \2160_b0 , \2161_b1 , \2161_b0 , 
		\2162_b1 , \2162_b0 , \2163_b1 , \2163_b0 , \2164_b1 , \2164_b0 , \2165_b1 , \2165_b0 , \2166_b1 , \2166_b0 , 
		\2167_b1 , \2167_b0 , \2168_b1 , \2168_b0 , \2169_b1 , \2169_b0 , \2170_b1 , \2170_b0 , \2171_b1 , \2171_b0 , 
		\2172_b1 , \2172_b0 , \2173_b1 , \2173_b0 , \2174_b1 , \2174_b0 , \2175_b1 , \2175_b0 , \2176_b1 , \2176_b0 , 
		\2177_b1 , \2177_b0 , \2178_b1 , \2178_b0 , \2179_b1 , \2179_b0 , \2180_b1 , \2180_b0 , \2181_b1 , \2181_b0 , 
		\2182_b1 , \2182_b0 , \2183_b1 , \2183_b0 , \2184_b1 , \2184_b0 , \2185_b1 , \2185_b0 , \2186_b1 , \2186_b0 , 
		\2187_b1 , \2187_b0 , \2188_b1 , \2188_b0 , \2189_b1 , \2189_b0 , \2190_b1 , \2190_b0 , \2191_b1 , \2191_b0 , 
		\2192_b1 , \2192_b0 , \2193_b1 , \2193_b0 , \2194_b1 , \2194_b0 , \2195_b1 , \2195_b0 , \2196_b1 , \2196_b0 , 
		\2197_b1 , \2197_b0 , \2198_b1 , \2198_b0 , \2199_b1 , \2199_b0 , \2200_b1 , \2200_b0 , \2201_b1 , \2201_b0 , 
		\2202_b1 , \2202_b0 , \2203_b1 , \2203_b0 , \2204_b1 , \2204_b0 , \2205_b1 , \2205_b0 , \2206_b1 , \2206_b0 , 
		\2207_b1 , \2207_b0 , \2208_b1 , \2208_b0 , \2209_b1 , \2209_b0 , \2210_b1 , \2210_b0 , \2211_b1 , \2211_b0 , 
		\2212_b1 , \2212_b0 , \2213_b1 , \2213_b0 , \2214_b1 , \2214_b0 , \2215_b1 , \2215_b0 , \2216_b1 , \2216_b0 , 
		\2217_b1 , \2217_b0 , \2218_b1 , \2218_b0 , \2219_b1 , \2219_b0 , \2220_b1 , \2220_b0 , \2221_b1 , \2221_b0 , 
		\2222_b1 , \2222_b0 , \2223_b1 , \2223_b0 , \2224_b1 , \2224_b0 , \2225_b1 , \2225_b0 , \2226_b1 , \2226_b0 , 
		\2227_b1 , \2227_b0 , \2228_b1 , \2228_b0 , \2229_b1 , \2229_b0 , \2230_b1 , \2230_b0 , \2231_b1 , \2231_b0 , 
		\2232_b1 , \2232_b0 , \2233_b1 , \2233_b0 , \2234_b1 , \2234_b0 , \2235_b1 , \2235_b0 , \2236_b1 , \2236_b0 , 
		\2237_b1 , \2237_b0 , \2238_b1 , \2238_b0 , \2239_b1 , \2239_b0 , \2240_b1 , \2240_b0 , \2241_b1 , \2241_b0 , 
		\2242_b1 , \2242_b0 , \2243_b1 , \2243_b0 , \2244_b1 , \2244_b0 , \2245_b1 , \2245_b0 , \2246_b1 , \2246_b0 , 
		\2247_b1 , \2247_b0 , \2248_b1 , \2248_b0 , \2249_b1 , \2249_b0 , \2250_b1 , \2250_b0 , \2251_b1 , \2251_b0 , 
		\2252_b1 , \2252_b0 , \2253_b1 , \2253_b0 , \2254_b1 , \2254_b0 , \2255_b1 , \2255_b0 , \2256_b1 , \2256_b0 , 
		\2257_b1 , \2257_b0 , \2258_b1 , \2258_b0 , \2259_b1 , \2259_b0 , \2260_b1 , \2260_b0 , \2261_b1 , \2261_b0 , 
		\2262_b1 , \2262_b0 , \2263_b1 , \2263_b0 , \2264_b1 , \2264_b0 , \2265_b1 , \2265_b0 , \2266_b1 , \2266_b0 , 
		\2267_b1 , \2267_b0 , \2268_b1 , \2268_b0 , \2269_b1 , \2269_b0 , \2270_b1 , \2270_b0 , \2271_b1 , \2271_b0 , 
		\2272_b1 , \2272_b0 , \2273_b1 , \2273_b0 , \2274_b1 , \2274_b0 , \2275_b1 , \2275_b0 , \2276_b1 , \2276_b0 , 
		\2277_b1 , \2277_b0 , \2278_b1 , \2278_b0 , \2279_b1 , \2279_b0 , \2280_b1 , \2280_b0 , \2281_b1 , \2281_b0 , 
		\2282_b1 , \2282_b0 , \2283_b1 , \2283_b0 , \2284_b1 , \2284_b0 , \2285_b1 , \2285_b0 , \2286_b1 , \2286_b0 , 
		\2287_b1 , \2287_b0 , \2288_b1 , \2288_b0 , \2289_b1 , \2289_b0 , \2290_b1 , \2290_b0 , \2291_b1 , \2291_b0 , 
		\2292_b1 , \2292_b0 , \2293_b1 , \2293_b0 , \2294_b1 , \2294_b0 , \2295_b1 , \2295_b0 , \2296_b1 , \2296_b0 , 
		\2297_b1 , \2297_b0 , \2298_b1 , \2298_b0 , \2299_b1 , \2299_b0 , \2300_b1 , \2300_b0 , \2301_b1 , \2301_b0 , 
		\2302_b1 , \2302_b0 , \2303_b1 , \2303_b0 , \2304_b1 , \2304_b0 , \2305_b1 , \2305_b0 , \2306_b1 , \2306_b0 , 
		\2307_b1 , \2307_b0 , \2308_b1 , \2308_b0 , \2309_b1 , \2309_b0 , \2310_b1 , \2310_b0 , \2311_b1 , \2311_b0 , 
		\2312_b1 , \2312_b0 , \2313_b1 , \2313_b0 , \2314_b1 , \2314_b0 , \2315_b1 , \2315_b0 , \2316_b1 , \2316_b0 , 
		\2317_b1 , \2317_b0 , \2318_b1 , \2318_b0 , \2319_b1 , \2319_b0 , \2320_b1 , \2320_b0 , \2321_b1 , \2321_b0 , 
		\2322_b1 , \2322_b0 , \2323_b1 , \2323_b0 , \2324_b1 , \2324_b0 , \2325_b1 , \2325_b0 , \2326_b1 , \2326_b0 , 
		\2327_b1 , \2327_b0 , \2328_b1 , \2328_b0 , \2329_b1 , \2329_b0 , \2330_b1 , \2330_b0 , \2331_b1 , \2331_b0 , 
		\2332_b1 , \2332_b0 , \2333_b1 , \2333_b0 , \2334_b1 , \2334_b0 , \2335_b1 , \2335_b0 , \2336_b1 , \2336_b0 , 
		\2337_b1 , \2337_b0 , \2338_b1 , \2338_b0 , \2339_b1 , \2339_b0 , \2340_b1 , \2340_b0 , \2341_b1 , \2341_b0 , 
		\2342_b1 , \2342_b0 , \2343_b1 , \2343_b0 , \2344_b1 , \2344_b0 , \2345_b1 , \2345_b0 , \2346_b1 , \2346_b0 , 
		\2347_b1 , \2347_b0 , \2348_b1 , \2348_b0 , \2349_b1 , \2349_b0 , \2350_b1 , \2350_b0 , \2351_b1 , \2351_b0 , 
		\2352_b1 , \2352_b0 , \2353_b1 , \2353_b0 , \2354_b1 , \2354_b0 , \2355_b1 , \2355_b0 , \2356_b1 , \2356_b0 , 
		\2357_b1 , \2357_b0 , \2358_b1 , \2358_b0 , \2359_b1 , \2359_b0 , \2360_b1 , \2360_b0 , \2361_b1 , \2361_b0 , 
		\2362_b1 , \2362_b0 , \2363_b1 , \2363_b0 , \2364_b1 , \2364_b0 , \2365_b1 , \2365_b0 , \2366_b1 , \2366_b0 , 
		\2367_b1 , \2367_b0 , \2368_b1 , \2368_b0 , \2369_b1 , \2369_b0 , \2370_b1 , \2370_b0 , \2371_b1 , \2371_b0 , 
		\2372_b1 , \2372_b0 , \2373_b1 , \2373_b0 , \2374_b1 , \2374_b0 , \2375_b1 , \2375_b0 , \2376_b1 , \2376_b0 , 
		\2377_b1 , \2377_b0 , \2378_b1 , \2378_b0 , \2379_b1 , \2379_b0 , \2380_b1 , \2380_b0 , \2381_b1 , \2381_b0 , 
		\2382_b1 , \2382_b0 , \2383_b1 , \2383_b0 , \2384_b1 , \2384_b0 , \2385_b1 , \2385_b0 , \2386_b1 , \2386_b0 , 
		\2387_b1 , \2387_b0 , \2388_b1 , \2388_b0 , \2389_b1 , \2389_b0 , \2390_b1 , \2390_b0 , \2391_b1 , \2391_b0 , 
		\2392_b1 , \2392_b0 , \2393_b1 , \2393_b0 , \2394_b1 , \2394_b0 , \2395_b1 , \2395_b0 , \2396_b1 , \2396_b0 , 
		\2397_b1 , \2397_b0 , \2398_b1 , \2398_b0 , \2399_b1 , \2399_b0 , \2400_b1 , \2400_b0 , \2401_b1 , \2401_b0 , 
		\2402_b1 , \2402_b0 , \2403_b1 , \2403_b0 , \2404_b1 , \2404_b0 , \2405_b1 , \2405_b0 , \2406_b1 , \2406_b0 , 
		\2407_b1 , \2407_b0 , \2408_b1 , \2408_b0 , \2409_b1 , \2409_b0 , \2410_b1 , \2410_b0 , \2411_b1 , \2411_b0 , 
		\2412_b1 , \2412_b0 , \2413_b1 , \2413_b0 , \2414_b1 , \2414_b0 , \2415_b1 , \2415_b0 , \2416_b1 , \2416_b0 , 
		\2417_b1 , \2417_b0 , \2418_b1 , \2418_b0 , \2419_b1 , \2419_b0 , \2420_b1 , \2420_b0 , \2421_b1 , \2421_b0 , 
		\2422_b1 , \2422_b0 , \2423_b1 , \2423_b0 , \2424_b1 , \2424_b0 , \2425_b1 , \2425_b0 , \2426_b1 , \2426_b0 , 
		\2427_b1 , \2427_b0 , \2428_b1 , \2428_b0 , \2429_b1 , \2429_b0 , \2430_b1 , \2430_b0 , \2431_b1 , \2431_b0 , 
		\2432_b1 , \2432_b0 , \2433_b1 , \2433_b0 , \2434_b1 , \2434_b0 , \2435_b1 , \2435_b0 , \2436_b1 , \2436_b0 , 
		\2437_b1 , \2437_b0 , \2438_b1 , \2438_b0 , \2439_b1 , \2439_b0 , \2440_b1 , \2440_b0 , \2441_b1 , \2441_b0 , 
		\2442_b1 , \2442_b0 , \2443_b1 , \2443_b0 , \2444_b1 , \2444_b0 , \2445_b1 , \2445_b0 , \2446_b1 , \2446_b0 , 
		\2447_b1 , \2447_b0 , \2448_b1 , \2448_b0 , \2449_b1 , \2449_b0 , \2450_b1 , \2450_b0 , \2451_b1 , \2451_b0 , 
		\2452_b1 , \2452_b0 , \2453_b1 , \2453_b0 , \2454_b1 , \2454_b0 , \2455_b1 , \2455_b0 , \2456_b1 , \2456_b0 , 
		\2457_b1 , \2457_b0 , \2458_b1 , \2458_b0 , \2459_b1 , \2459_b0 , \2460_b1 , \2460_b0 , \2461_b1 , \2461_b0 , 
		\2462_b1 , \2462_b0 , \2463_b1 , \2463_b0 , \2464_b1 , \2464_b0 , \2465_b1 , \2465_b0 , \2466_b1 , \2466_b0 , 
		\2467_b1 , \2467_b0 , \2468_b1 , \2468_b0 , \2469_b1 , \2469_b0 , \2470_b1 , \2470_b0 , \2471_b1 , \2471_b0 , 
		\2472_b1 , \2472_b0 , \2473_b1 , \2473_b0 , \2474_b1 , \2474_b0 , \2475_b1 , \2475_b0 , \2476_b1 , \2476_b0 , 
		\2477_b1 , \2477_b0 , \2478_b1 , \2478_b0 , \2479_b1 , \2479_b0 , \2480_b1 , \2480_b0 , \2481_b1 , \2481_b0 , 
		\2482_b1 , \2482_b0 , \2483_b1 , \2483_b0 , \2484_b1 , \2484_b0 , \2485_b1 , \2485_b0 , \2486_b1 , \2486_b0 , 
		\2487_b1 , \2487_b0 , \2488_b1 , \2488_b0 , \2489_b1 , \2489_b0 , \2490_b1 , \2490_b0 , \2491_b1 , \2491_b0 , 
		\2492_b1 , \2492_b0 , \2493_b1 , \2493_b0 , \2494_b1 , \2494_b0 , \2495_b1 , \2495_b0 , \2496_b1 , \2496_b0 , 
		\2497_b1 , \2497_b0 , \2498_b1 , \2498_b0 , \2499_b1 , \2499_b0 , \2500_b1 , \2500_b0 , \2501_b1 , \2501_b0 , 
		\2502_b1 , \2502_b0 , \2503_b1 , \2503_b0 , \2504_b1 , \2504_b0 , \2505_b1 , \2505_b0 , \2506_b1 , \2506_b0 , 
		\2507_b1 , \2507_b0 , \2508_b1 , \2508_b0 , \2509_b1 , \2509_b0 , \2510_b1 , \2510_b0 , \2511_b1 , \2511_b0 , 
		\2512_b1 , \2512_b0 , \2513_b1 , \2513_b0 , \2514_b1 , \2514_b0 , \2515_b1 , \2515_b0 , \2516_b1 , \2516_b0 , 
		\2517_b1 , \2517_b0 , \2518_b1 , \2518_b0 , \2519_b1 , \2519_b0 , \2520_b1 , \2520_b0 , \2521_b1 , \2521_b0 , 
		\2522_b1 , \2522_b0 , \2523_b1 , \2523_b0 , \2524_b1 , \2524_b0 , \2525_b1 , \2525_b0 , \2526_b1 , \2526_b0 , 
		\2527_b1 , \2527_b0 , \2528_b1 , \2528_b0 , \2529_b1 , \2529_b0 , \2530_b1 , \2530_b0 , \2531_b1 , \2531_b0 , 
		\2532_b1 , \2532_b0 , \2533_b1 , \2533_b0 , \2534_b1 , \2534_b0 , \2535_b1 , \2535_b0 , \2536_b1 , \2536_b0 , 
		\2537_b1 , \2537_b0 , \2538_b1 , \2538_b0 , \2539_b1 , \2539_b0 , \2540_b1 , \2540_b0 , \2541_b1 , \2541_b0 , 
		\2542_b1 , \2542_b0 , \2543_b1 , \2543_b0 , \2544_b1 , \2544_b0 , \2545_b1 , \2545_b0 , \2546_b1 , \2546_b0 , 
		\2547_b1 , \2547_b0 , \2548_b1 , \2548_b0 , \2549_b1 , \2549_b0 , \2550_b1 , \2550_b0 , \2551_b1 , \2551_b0 , 
		\2552_b1 , \2552_b0 , \2553_b1 , \2553_b0 , \2554_b1 , \2554_b0 , \2555_b1 , \2555_b0 , \2556_b1 , \2556_b0 , 
		\2557_b1 , \2557_b0 , \2558_b1 , \2558_b0 , \2559_b1 , \2559_b0 , \2560_b1 , \2560_b0 , \2561_b1 , \2561_b0 , 
		\2562_b1 , \2562_b0 , \2563_b1 , \2563_b0 , \2564_b1 , \2564_b0 , \2565_b1 , \2565_b0 , \2566_b1 , \2566_b0 , 
		\2567_b1 , \2567_b0 , \2568_b1 , \2568_b0 , \2569_b1 , \2569_b0 , \2570_b1 , \2570_b0 , \2571_b1 , \2571_b0 , 
		\2572_b1 , \2572_b0 , \2573_b1 , \2573_b0 , \2574_b1 , \2574_b0 , \2575_b1 , \2575_b0 , \2576_b1 , \2576_b0 , 
		\2577_b1 , \2577_b0 , \2578_b1 , \2578_b0 , \2579_b1 , \2579_b0 , \2580_b1 , \2580_b0 , \2581_b1 , \2581_b0 , 
		\2582_b1 , \2582_b0 , \2583_b1 , \2583_b0 , \2584_b1 , \2584_b0 , \2585_b1 , \2585_b0 , \2586_b1 , \2586_b0 , 
		\2587_b1 , \2587_b0 , \2588_b1 , \2588_b0 , \2589_b1 , \2589_b0 , \2590_b1 , \2590_b0 , \2591_b1 , \2591_b0 , 
		\2592_b1 , \2592_b0 , \2593_b1 , \2593_b0 , \2594_b1 , \2594_b0 , \2595_b1 , \2595_b0 , \2596_b1 , \2596_b0 , 
		\2597_b1 , \2597_b0 , \2598_b1 , \2598_b0 , \2599_b1 , \2599_b0 , \2600_b1 , \2600_b0 , \2601_b1 , \2601_b0 , 
		\2602_b1 , \2602_b0 , \2603_b1 , \2603_b0 , \2604_b1 , \2604_b0 , \2605_b1 , \2605_b0 , \2606_b1 , \2606_b0 , 
		\2607_b1 , \2607_b0 , \2608_b1 , \2608_b0 , \2609_b1 , \2609_b0 , \2610_b1 , \2610_b0 , \2611_b1 , \2611_b0 , 
		\2612_b1 , \2612_b0 , \2613_b1 , \2613_b0 , \2614_b1 , \2614_b0 , \2615_b1 , \2615_b0 , \2616_b1 , \2616_b0 , 
		\2617_b1 , \2617_b0 , \2618_b1 , \2618_b0 , \2619_b1 , \2619_b0 , \2620_b1 , \2620_b0 , \2621_b1 , \2621_b0 , 
		\2622_b1 , \2622_b0 , \2623_b1 , \2623_b0 , \2624_b1 , \2624_b0 , \2625_b1 , \2625_b0 , \2626_b1 , \2626_b0 , 
		\2627_b1 , \2627_b0 , \2628_b1 , \2628_b0 , \2629_b1 , \2629_b0 , \2630_b1 , \2630_b0 , \2631_b1 , \2631_b0 , 
		\2632_b1 , \2632_b0 , \2633_b1 , \2633_b0 , \2634_b1 , \2634_b0 , \2635_b1 , \2635_b0 , \2636_b1 , \2636_b0 , 
		\2637_b1 , \2637_b0 , \2638_b1 , \2638_b0 , \2639_b1 , \2639_b0 , \2640_b1 , \2640_b0 , \2641_b1 , \2641_b0 , 
		\2642_b1 , \2642_b0 , \2643_b1 , \2643_b0 , \2644_b1 , \2644_b0 , \2645_b1 , \2645_b0 , \2646_b1 , \2646_b0 , 
		\2647_b1 , \2647_b0 , \2648_b1 , \2648_b0 , \2649_b1 , \2649_b0 , \2650_b1 , \2650_b0 , \2651_b1 , \2651_b0 , 
		\2652_b1 , \2652_b0 , \2653_b1 , \2653_b0 , \2654_b1 , \2654_b0 , \2655_b1 , \2655_b0 , \2656_b1 , \2656_b0 , 
		\2657_b1 , \2657_b0 , \2658_b1 , \2658_b0 , \2659_b1 , \2659_b0 , \2660_b1 , \2660_b0 , \2661_b1 , \2661_b0 , 
		\2662_b1 , \2662_b0 , \2663_b1 , \2663_b0 , \2664_b1 , \2664_b0 , \2665_b1 , \2665_b0 , \2666_b1 , \2666_b0 , 
		\2667_b1 , \2667_b0 , \2668_b1 , \2668_b0 , \2669_b1 , \2669_b0 , \2670_b1 , \2670_b0 , \2671_b1 , \2671_b0 , 
		\2672_b1 , \2672_b0 , \2673_b1 , \2673_b0 , \2674_b1 , \2674_b0 , \2675_b1 , \2675_b0 , \2676_b1 , \2676_b0 , 
		\2677_b1 , \2677_b0 , \2678_b1 , \2678_b0 , \2679_b1 , \2679_b0 , \2680_b1 , \2680_b0 , \2681_b1 , \2681_b0 , 
		\2682_b1 , \2682_b0 , \2683_b1 , \2683_b0 , \2684_b1 , \2684_b0 , \2685_b1 , \2685_b0 , \2686_b1 , \2686_b0 , 
		\2687_b1 , \2687_b0 , \2688_b1 , \2688_b0 , \2689_b1 , \2689_b0 , \2690_b1 , \2690_b0 , \2691_b1 , \2691_b0 , 
		\2692_b1 , \2692_b0 , \2693_b1 , \2693_b0 , \2694_b1 , \2694_b0 , \2695_b1 , \2695_b0 , \2696_b1 , \2696_b0 , 
		\2697_b1 , \2697_b0 , \2698_b1 , \2698_b0 , \2699_b1 , \2699_b0 , \2700_b1 , \2700_b0 , \2701_b1 , \2701_b0 , 
		\2702_b1 , \2702_b0 , \2703_b1 , \2703_b0 , \2704_b1 , \2704_b0 , \2705_b1 , \2705_b0 , \2706_b1 , \2706_b0 , 
		\2707_b1 , \2707_b0 , \2708_b1 , \2708_b0 , \2709_b1 , \2709_b0 , \2710_b1 , \2710_b0 , \2711_b1 , \2711_b0 , 
		\2712_b1 , \2712_b0 , \2713_b1 , \2713_b0 , \2714_b1 , \2714_b0 , \2715_b1 , \2715_b0 , \2716_b1 , \2716_b0 , 
		\2717_b1 , \2717_b0 , \2718_b1 , \2718_b0 , \2719_b1 , \2719_b0 , \2720_b1 , \2720_b0 , \2721_b1 , \2721_b0 , 
		\2722_b1 , \2722_b0 , \2723_b1 , \2723_b0 , \2724_b1 , \2724_b0 , \2725_b1 , \2725_b0 , \2726_b1 , \2726_b0 , 
		\2727_b1 , \2727_b0 , \2728_b1 , \2728_b0 , \2729_b1 , \2729_b0 , \2730_b1 , \2730_b0 , \2731_b1 , \2731_b0 , 
		\2732_b1 , \2732_b0 , \2733_b1 , \2733_b0 , \2734_b1 , \2734_b0 , \2735_b1 , \2735_b0 , \2736_b1 , \2736_b0 , 
		\2737_b1 , \2737_b0 , \2738_b1 , \2738_b0 , \2739_b1 , \2739_b0 , \2740_b1 , \2740_b0 , \2741_b1 , \2741_b0 , 
		\2742_b1 , \2742_b0 , \2743_b1 , \2743_b0 , \2744_b1 , \2744_b0 , \2745_b1 , \2745_b0 , \2746_b1 , \2746_b0 , 
		\2747_b1 , \2747_b0 , \2748_b1 , \2748_b0 , \2749_b1 , \2749_b0 , \2750_b1 , \2750_b0 , \2751_b1 , \2751_b0 , 
		\2752_b1 , \2752_b0 , \2753_b1 , \2753_b0 , \2754_b1 , \2754_b0 , \2755_b1 , \2755_b0 , \2756_b1 , \2756_b0 , 
		\2757_b1 , \2757_b0 , \2758_b1 , \2758_b0 , \2759_b1 , \2759_b0 , \2760_b1 , \2760_b0 , \2761_b1 , \2761_b0 , 
		\2762_b1 , \2762_b0 , \2763_b1 , \2763_b0 , \2764_b1 , \2764_b0 , \2765_b1 , \2765_b0 , \2766_b1 , \2766_b0 , 
		\2767_b1 , \2767_b0 , \2768_b1 , \2768_b0 , \2769_b1 , \2769_b0 , \2770_b1 , \2770_b0 , \2771_b1 , \2771_b0 , 
		\2772_b1 , \2772_b0 , \2773_b1 , \2773_b0 , \2774_b1 , \2774_b0 , \2775_b1 , \2775_b0 , \2776_b1 , \2776_b0 , 
		\2777_b1 , \2777_b0 , \2778_b1 , \2778_b0 , \2779_b1 , \2779_b0 , \2780_b1 , \2780_b0 , \2781_b1 , \2781_b0 , 
		\2782_b1 , \2782_b0 , \2783_b1 , \2783_b0 , \2784_b1 , \2784_b0 , \2785_b1 , \2785_b0 , \2786_b1 , \2786_b0 , 
		\2787_b1 , \2787_b0 , \2788_b1 , \2788_b0 , \2789_b1 , \2789_b0 , \2790_b1 , \2790_b0 , \2791_b1 , \2791_b0 , 
		\2792_b1 , \2792_b0 , \2793_b1 , \2793_b0 , \2794_b1 , \2794_b0 , \2795_b1 , \2795_b0 , \2796_b1 , \2796_b0 , 
		\2797_b1 , \2797_b0 , \2798_b1 , \2798_b0 , \2799_b1 , \2799_b0 , \2800_b1 , \2800_b0 , \2801_b1 , \2801_b0 , 
		\2802_b1 , \2802_b0 , \2803_b1 , \2803_b0 , \2804_b1 , \2804_b0 , \2805_b1 , \2805_b0 , \2806_b1 , \2806_b0 , 
		\2807_b1 , \2807_b0 , \2808_b1 , \2808_b0 , \2809_b1 , \2809_b0 , \2810_b1 , \2810_b0 , \2811_b1 , \2811_b0 , 
		\2812_b1 , \2812_b0 , \2813_b1 , \2813_b0 , \2814_b1 , \2814_b0 , \2815_b1 , \2815_b0 , \2816_b1 , \2816_b0 , 
		\2817_b1 , \2817_b0 , \2818_b1 , \2818_b0 , \2819_b1 , \2819_b0 , \2820_b1 , \2820_b0 , \2821_b1 , \2821_b0 , 
		\2822_b1 , \2822_b0 , \2823_b1 , \2823_b0 , \2824_b1 , \2824_b0 , \2825_b1 , \2825_b0 , \2826_b1 , \2826_b0 , 
		\2827_b1 , \2827_b0 , \2828_b1 , \2828_b0 , \2829_b1 , \2829_b0 , \2830_b1 , \2830_b0 , \2831_b1 , \2831_b0 , 
		\2832_b1 , \2832_b0 , \2833_b1 , \2833_b0 , \2834_b1 , \2834_b0 , \2835_b1 , \2835_b0 , \2836_b1 , \2836_b0 , 
		\2837_b1 , \2837_b0 , \2838_b1 , \2838_b0 , \2839_b1 , \2839_b0 , \2840_b1 , \2840_b0 , \2841_b1 , \2841_b0 , 
		\2842_b1 , \2842_b0 , \2843_b1 , \2843_b0 , \2844_b1 , \2844_b0 , \2845_b1 , \2845_b0 , \2846_b1 , \2846_b0 , 
		\2847_b1 , \2847_b0 , \2848_b1 , \2848_b0 , \2849_b1 , \2849_b0 , \2850_b1 , \2850_b0 , \2851_b1 , \2851_b0 , 
		\2852_b1 , \2852_b0 , \2853_b1 , \2853_b0 , \2854_b1 , \2854_b0 , \2855_b1 , \2855_b0 , \2856_b1 , \2856_b0 , 
		\2857_b1 , \2857_b0 , \2858_b1 , \2858_b0 , \2859_b1 , \2859_b0 , \2860_b1 , \2860_b0 , \2861_b1 , \2861_b0 , 
		\2862_b1 , \2862_b0 , \2863_b1 , \2863_b0 , \2864_b1 , \2864_b0 , \2865_b1 , \2865_b0 , \2866_b1 , \2866_b0 , 
		\2867_b1 , \2867_b0 , \2868_b1 , \2868_b0 , \2869_b1 , \2869_b0 , \2870_b1 , \2870_b0 , \2871_b1 , \2871_b0 , 
		\2872_b1 , \2872_b0 , \2873_b1 , \2873_b0 , \2874_b1 , \2874_b0 , \2875_b1 , \2875_b0 , \2876_b1 , \2876_b0 , 
		\2877_b1 , \2877_b0 , \2878_b1 , \2878_b0 , \2879_b1 , \2879_b0 , \2880_b1 , \2880_b0 , \2881_b1 , \2881_b0 , 
		\2882_b1 , \2882_b0 , \2883_b1 , \2883_b0 , \2884_b1 , \2884_b0 , \2885_b1 , \2885_b0 , \2886_b1 , \2886_b0 , 
		\2887_b1 , \2887_b0 , \2888_b1 , \2888_b0 , \2889_b1 , \2889_b0 , \2890_b1 , \2890_b0 , \2891_b1 , \2891_b0 , 
		\2892_b1 , \2892_b0 , \2893_b1 , \2893_b0 , \2894_b1 , \2894_b0 , \2895_b1 , \2895_b0 , \2896_b1 , \2896_b0 , 
		\2897_b1 , \2897_b0 , \2898_b1 , \2898_b0 , \2899_b1 , \2899_b0 , \2900_b1 , \2900_b0 , \2901_b1 , \2901_b0 , 
		\2902_b1 , \2902_b0 , \2903_b1 , \2903_b0 , \2904_b1 , \2904_b0 , \2905_b1 , \2905_b0 , \2906_b1 , \2906_b0 , 
		\2907_b1 , \2907_b0 , \2908_b1 , \2908_b0 , \2909_b1 , \2909_b0 , \2910_b1 , \2910_b0 , \2911_b1 , \2911_b0 , 
		\2912_b1 , \2912_b0 , \2913_b1 , \2913_b0 , \2914_b1 , \2914_b0 , \2915_b1 , \2915_b0 , \2916_b1 , \2916_b0 , 
		\2917_b1 , \2917_b0 , \2918_b1 , \2918_b0 , \2919_b1 , \2919_b0 , \2920_b1 , \2920_b0 , \2921_b1 , \2921_b0 , 
		\2922_b1 , \2922_b0 , \2923_b1 , \2923_b0 , \2924_b1 , \2924_b0 , \2925_b1 , \2925_b0 , \2926_b1 , \2926_b0 , 
		\2927_b1 , \2927_b0 , \2928_b1 , \2928_b0 , \2929_b1 , \2929_b0 , \2930_b1 , \2930_b0 , \2931_b1 , \2931_b0 , 
		\2932_b1 , \2932_b0 , \2933_b1 , \2933_b0 , \2934_b1 , \2934_b0 , \2935_b1 , \2935_b0 , \2936_b1 , \2936_b0 , 
		\2937_b1 , \2937_b0 , \2938_b1 , \2938_b0 , \2939_b1 , \2939_b0 , \2940_b1 , \2940_b0 , \2941_b1 , \2941_b0 , 
		\2942_b1 , \2942_b0 , \2943_b1 , \2943_b0 , \2944_b1 , \2944_b0 , \2945_b1 , \2945_b0 , \2946_b1 , \2946_b0 , 
		\2947_b1 , \2947_b0 , \2948_b1 , \2948_b0 , \2949_b1 , \2949_b0 , \2950_b1 , \2950_b0 , \2951_b1 , \2951_b0 , 
		\2952_b1 , \2952_b0 , \2953_b1 , \2953_b0 , \2954_b1 , \2954_b0 , \2955_b1 , \2955_b0 , \2956_b1 , \2956_b0 , 
		\2957_b1 , \2957_b0 , \2958_b1 , \2958_b0 , \2959_b1 , \2959_b0 , \2960_b1 , \2960_b0 , \2961_b1 , \2961_b0 , 
		\2962_b1 , \2962_b0 , \2963_b1 , \2963_b0 , \2964_b1 , \2964_b0 , \2965_b1 , \2965_b0 , \2966_b1 , \2966_b0 , 
		\2967_b1 , \2967_b0 , \2968_b1 , \2968_b0 , \2969_b1 , \2969_b0 , \2970_b1 , \2970_b0 , \2971_b1 , \2971_b0 , 
		\2972_b1 , \2972_b0 , \2973_b1 , \2973_b0 , \2974_b1 , \2974_b0 , \2975_b1 , \2975_b0 , \2976_b1 , \2976_b0 , 
		\2977_b1 , \2977_b0 , \2978_b1 , \2978_b0 , \2979_b1 , \2979_b0 , \2980_b1 , \2980_b0 , \2981_b1 , \2981_b0 , 
		\2982_b1 , \2982_b0 , \2983_b1 , \2983_b0 , \2984_b1 , \2984_b0 , \2985_b1 , \2985_b0 , \2986_b1 , \2986_b0 , 
		\2987_b1 , \2987_b0 , \2988_b1 , \2988_b0 , \2989_b1 , \2989_b0 , \2990_b1 , \2990_b0 , \2991_b1 , \2991_b0 , 
		\2992_b1 , \2992_b0 , \2993_b1 , \2993_b0 , \2994_b1 , \2994_b0 , \2995_b1 , \2995_b0 , \2996_b1 , \2996_b0 , 
		\2997_b1 , \2997_b0 , \2998_b1 , \2998_b0 , \2999_b1 , \2999_b0 , \3000_b1 , \3000_b0 , \3001_b1 , \3001_b0 , 
		\3002_b1 , \3002_b0 , \3003_b1 , \3003_b0 , \3004_b1 , \3004_b0 , \3005_b1 , \3005_b0 , \3006_b1 , \3006_b0 , 
		\3007_b1 , \3007_b0 , \3008_b1 , \3008_b0 , \3009_b1 , \3009_b0 , \3010_b1 , \3010_b0 , \3011_b1 , \3011_b0 , 
		\3012_b1 , \3012_b0 , \3013_b1 , \3013_b0 , \3014_b1 , \3014_b0 , \3015_b1 , \3015_b0 , \3016_b1 , \3016_b0 , 
		\3017_b1 , \3017_b0 , \3018_b1 , \3018_b0 , \3019_b1 , \3019_b0 , \3020_b1 , \3020_b0 , \3021_b1 , \3021_b0 , 
		\3022_b1 , \3022_b0 , \3023_b1 , \3023_b0 , \3024_b1 , \3024_b0 , \3025_b1 , \3025_b0 , \3026_b1 , \3026_b0 , 
		\3027_b1 , \3027_b0 , \3028_b1 , \3028_b0 , \3029_b1 , \3029_b0 , \3030_b1 , \3030_b0 , \3031_b1 , \3031_b0 , 
		\3032_b1 , \3032_b0 , \3033_b1 , \3033_b0 , \3034_b1 , \3034_b0 , \3035_b1 , \3035_b0 , \3036_b1 , \3036_b0 , 
		\3037_b1 , \3037_b0 , \3038_b1 , \3038_b0 , \3039_b1 , \3039_b0 , \3040_b1 , \3040_b0 , \3041_b1 , \3041_b0 , 
		\3042_b1 , \3042_b0 , \3043_b1 , \3043_b0 , \3044_b1 , \3044_b0 , \3045_b1 , \3045_b0 , \3046_b1 , \3046_b0 , 
		\3047_b1 , \3047_b0 , \3048_b1 , \3048_b0 , \3049_b1 , \3049_b0 , \3050_b1 , \3050_b0 , \3051_b1 , \3051_b0 , 
		\3052_b1 , \3052_b0 , \3053_b1 , \3053_b0 , \3054_b1 , \3054_b0 , \3055_b1 , \3055_b0 , \3056_b1 , \3056_b0 , 
		\3057_b1 , \3057_b0 , \3058_b1 , \3058_b0 , \3059_b1 , \3059_b0 , \3060_b1 , \3060_b0 , \3061_b1 , \3061_b0 , 
		\3062_b1 , \3062_b0 , \3063_b1 , \3063_b0 , \3064_b1 , \3064_b0 , \3065_b1 , \3065_b0 , \3066_b1 , \3066_b0 , 
		\3067_b1 , \3067_b0 , \3068_b1 , \3068_b0 , \3069_b1 , \3069_b0 , \3070_b1 , \3070_b0 , \3071_b1 , \3071_b0 , 
		\3072_b1 , \3072_b0 , \3073_b1 , \3073_b0 , \3074_b1 , \3074_b0 , \3075_b1 , \3075_b0 , \3076_b1 , \3076_b0 , 
		\3077_b1 , \3077_b0 , \3078_b1 , \3078_b0 , \3079_b1 , \3079_b0 , \3080_b1 , \3080_b0 , \3081_b1 , \3081_b0 , 
		\3082_b1 , \3082_b0 , \3083_b1 , \3083_b0 , \3084_b1 , \3084_b0 , \3085_b1 , \3085_b0 , \3086_b1 , \3086_b0 , 
		\3087_b1 , \3087_b0 , \3088_b1 , \3088_b0 , \3089_b1 , \3089_b0 , \3090_b1 , \3090_b0 , \3091_b1 , \3091_b0 , 
		\3092_b1 , \3092_b0 , \3093_b1 , \3093_b0 , \3094_b1 , \3094_b0 , \3095_b1 , \3095_b0 , \3096_b1 , \3096_b0 , 
		\3097_b1 , \3097_b0 , \3098_b1 , \3098_b0 , \3099_b1 , \3099_b0 , \3100_b1 , \3100_b0 , \3101_b1 , \3101_b0 , 
		\3102_b1 , \3102_b0 , \3103_b1 , \3103_b0 , \3104_b1 , \3104_b0 , \3105_b1 , \3105_b0 , \3106_b1 , \3106_b0 , 
		\3107_b1 , \3107_b0 , \3108_b1 , \3108_b0 , \3109_b1 , \3109_b0 , \3110_b1 , \3110_b0 , \3111_b1 , \3111_b0 , 
		\3112_b1 , \3112_b0 , \3113_b1 , \3113_b0 , \3114_b1 , \3114_b0 , \3115_b1 , \3115_b0 , \3116_b1 , \3116_b0 , 
		\3117_b1 , \3117_b0 , \3118_b1 , \3118_b0 , \3119_b1 , \3119_b0 , \3120_b1 , \3120_b0 , \3121_b1 , \3121_b0 , 
		\3122_b1 , \3122_b0 , \3123_b1 , \3123_b0 , \3124_b1 , \3124_b0 , \3125_b1 , \3125_b0 , \3126_b1 , \3126_b0 , 
		\3127_b1 , \3127_b0 , \3128_b1 , \3128_b0 , \3129_b1 , \3129_b0 , \3130_b1 , \3130_b0 , \3131_b1 , \3131_b0 , 
		\3132_b1 , \3132_b0 , \3133_b1 , \3133_b0 , \3134_b1 , \3134_b0 , \3135_b1 , \3135_b0 , \3136_b1 , \3136_b0 , 
		\3137_b1 , \3137_b0 , \3138_b1 , \3138_b0 , \3139_b1 , \3139_b0 , \3140_b1 , \3140_b0 , \3141_b1 , \3141_b0 , 
		\3142_b1 , \3142_b0 , \3143_b1 , \3143_b0 , \3144_b1 , \3144_b0 , \3145_b1 , \3145_b0 , \3146_b1 , \3146_b0 , 
		\3147_b1 , \3147_b0 , \3148_b1 , \3148_b0 , \3149_b1 , \3149_b0 , \3150_b1 , \3150_b0 , \3151_b1 , \3151_b0 , 
		\3152_b1 , \3152_b0 , \3153_b1 , \3153_b0 , \3154_b1 , \3154_b0 , \3155_b1 , \3155_b0 , \3156_b1 , \3156_b0 , 
		\3157_b1 , \3157_b0 , \3158_b1 , \3158_b0 , \3159_b1 , \3159_b0 , \3160_b1 , \3160_b0 , \3161_b1 , \3161_b0 , 
		\3162_b1 , \3162_b0 , \3163_b1 , \3163_b0 , \3164_b1 , \3164_b0 , \3165_b1 , \3165_b0 , \3166_b1 , \3166_b0 , 
		\3167_b1 , \3167_b0 , \3168_b1 , \3168_b0 , \3169_b1 , \3169_b0 , \3170_b1 , \3170_b0 , \3171_b1 , \3171_b0 , 
		\3172_b1 , \3172_b0 , \3173_b1 , \3173_b0 , \3174_b1 , \3174_b0 , \3175_b1 , \3175_b0 , \3176_b1 , \3176_b0 , 
		\3177_b1 , \3177_b0 , \3178_b1 , \3178_b0 , \3179_b1 , \3179_b0 , \3180_b1 , \3180_b0 , \3181_b1 , \3181_b0 , 
		\3182_b1 , \3182_b0 , \3183_b1 , \3183_b0 , \3184_b1 , \3184_b0 , \3185_b1 , \3185_b0 , \3186_b1 , \3186_b0 , 
		\3187_b1 , \3187_b0 , \3188_b1 , \3188_b0 , \3189_b1 , \3189_b0 , \3190_b1 , \3190_b0 , \3191_b1 , \3191_b0 , 
		\3192_b1 , \3192_b0 , \3193_b1 , \3193_b0 , \3194_b1 , \3194_b0 , \3195_b1 , \3195_b0 , \3196_b1 , \3196_b0 , 
		\3197_b1 , \3197_b0 , \3198_b1 , \3198_b0 , \3199_b1 , \3199_b0 , \3200_b1 , \3200_b0 , \3201_b1 , \3201_b0 , 
		\3202_b1 , \3202_b0 , \3203_b1 , \3203_b0 , \3204_b1 , \3204_b0 , \3205_b1 , \3205_b0 , \3206_b1 , \3206_b0 , 
		\3207_b1 , \3207_b0 , \3208_b1 , \3208_b0 , \3209_b1 , \3209_b0 , \3210_b1 , \3210_b0 , \3211_b1 , \3211_b0 , 
		\3212_b1 , \3212_b0 , \3213_b1 , \3213_b0 , \3214_b1 , \3214_b0 , \3215_b1 , \3215_b0 , \3216_b1 , \3216_b0 , 
		\3217_b1 , \3217_b0 , \3218_b1 , \3218_b0 , \3219_b1 , \3219_b0 , \3220_b1 , \3220_b0 , \3221_b1 , \3221_b0 , 
		\3222_b1 , \3222_b0 , \3223_b1 , \3223_b0 , \3224_b1 , \3224_b0 , \3225_b1 , \3225_b0 , \3226_b1 , \3226_b0 , 
		\3227_b1 , \3227_b0 , \3228_b1 , \3228_b0 , \3229_b1 , \3229_b0 , \3230_b1 , \3230_b0 , \3231_b1 , \3231_b0 , 
		\3232_b1 , \3232_b0 , \3233_b1 , \3233_b0 , \3234_b1 , \3234_b0 , \3235_b1 , \3235_b0 , \3236_b1 , \3236_b0 , 
		\3237_b1 , \3237_b0 , \3238_b1 , \3238_b0 , \3239_b1 , \3239_b0 , \3240_b1 , \3240_b0 , \3241_b1 , \3241_b0 , 
		\3242_b1 , \3242_b0 , \3243_b1 , \3243_b0 , \3244_b1 , \3244_b0 , \3245_b1 , \3245_b0 , \3246_b1 , \3246_b0 , 
		\3247_b1 , \3247_b0 , \3248_b1 , \3248_b0 , \3249_b1 , \3249_b0 , \3250_b1 , \3250_b0 , \3251_b1 , \3251_b0 , 
		\3252_b1 , \3252_b0 , \3253_b1 , \3253_b0 , \3254_b1 , \3254_b0 , \3255_b1 , \3255_b0 , \3256_b1 , \3256_b0 , 
		\3257_b1 , \3257_b0 , \3258_b1 , \3258_b0 , \3259_b1 , \3259_b0 , \3260_b1 , \3260_b0 , \3261_b1 , \3261_b0 , 
		\3262_b1 , \3262_b0 , \3263_b1 , \3263_b0 , \3264_b1 , \3264_b0 , \3265_b1 , \3265_b0 , \3266_b1 , \3266_b0 , 
		\3267_b1 , \3267_b0 , \3268_b1 , \3268_b0 , \3269_b1 , \3269_b0 , \3270_b1 , \3270_b0 , \3271_b1 , \3271_b0 , 
		\3272_b1 , \3272_b0 , \3273_b1 , \3273_b0 , \3274_b1 , \3274_b0 , \3275_b1 , \3275_b0 , \3276_b1 , \3276_b0 , 
		\3277_b1 , \3277_b0 , \3278_b1 , \3278_b0 , \3279_b1 , \3279_b0 , \3280_b1 , \3280_b0 , \3281_b1 , \3281_b0 , 
		\3282_b1 , \3282_b0 , \3283_b1 , \3283_b0 , \3284_b1 , \3284_b0 , \3285_b1 , \3285_b0 , \3286_b1 , \3286_b0 , 
		\3287_b1 , \3287_b0 , \3288_b1 , \3288_b0 , \3289_b1 , \3289_b0 , \3290_b1 , \3290_b0 , \3291_b1 , \3291_b0 , 
		\3292_b1 , \3292_b0 , \3293_b1 , \3293_b0 , \3294_b1 , \3294_b0 , \3295_b1 , \3295_b0 , \3296_b1 , \3296_b0 , 
		\3297_b1 , \3297_b0 , \3298_b1 , \3298_b0 , \3299_b1 , \3299_b0 , \3300_b1 , \3300_b0 , \3301_b1 , \3301_b0 , 
		\3302_b1 , \3302_b0 , \3303_b1 , \3303_b0 , \3304_b1 , \3304_b0 , \3305_b1 , \3305_b0 , \3306_b1 , \3306_b0 , 
		\3307_b1 , \3307_b0 , \3308_b1 , \3308_b0 , \3309_b1 , \3309_b0 , \3310_b1 , \3310_b0 , \3311_b1 , \3311_b0 , 
		\3312_b1 , \3312_b0 , \3313_b1 , \3313_b0 , \3314_b1 , \3314_b0 , \3315_b1 , \3315_b0 , \3316_b1 , \3316_b0 , 
		\3317_b1 , \3317_b0 , \3318_b1 , \3318_b0 , \3319_b1 , \3319_b0 , \3320_b1 , \3320_b0 , \3321_b1 , \3321_b0 , 
		\3322_b1 , \3322_b0 , \3323_b1 , \3323_b0 , \3324_b1 , \3324_b0 , \3325_b1 , \3325_b0 , \3326_b1 , \3326_b0 , 
		\3327_b1 , \3327_b0 , \3328_b1 , \3328_b0 , \3329_b1 , \3329_b0 , \3330_b1 , \3330_b0 , \3331_b1 , \3331_b0 , 
		\3332_b1 , \3332_b0 , \3333_b1 , \3333_b0 , \3334_b1 , \3334_b0 , \3335_b1 , \3335_b0 , \3336_b1 , \3336_b0 , 
		\3337_b1 , \3337_b0 , \3338_b1 , \3338_b0 , \3339_b1 , \3339_b0 , \3340_b1 , \3340_b0 , \3341_b1 , \3341_b0 , 
		\3342_b1 , \3342_b0 , \3343_b1 , \3343_b0 , \3344_b1 , \3344_b0 , \3345_b1 , \3345_b0 , \3346_b1 , \3346_b0 , 
		\3347_b1 , \3347_b0 , \3348_b1 , \3348_b0 , \3349_b1 , \3349_b0 , \3350_b1 , \3350_b0 , \3351_b1 , \3351_b0 , 
		\3352_b1 , \3352_b0 , \3353_b1 , \3353_b0 , \3354_b1 , \3354_b0 , \3355_b1 , \3355_b0 , \3356_b1 , \3356_b0 , 
		\3357_b1 , \3357_b0 , \3358_b1 , \3358_b0 , \3359_b1 , \3359_b0 , \3360_b1 , \3360_b0 , \3361_b1 , \3361_b0 , 
		\3362_b1 , \3362_b0 , \3363_b1 , \3363_b0 , \3364_b1 , \3364_b0 , \3365_b1 , \3365_b0 , \3366_b1 , \3366_b0 , 
		\3367_b1 , \3367_b0 , \3368_b1 , \3368_b0 , \3369_b1 , \3369_b0 , \3370_b1 , \3370_b0 , \3371_b1 , \3371_b0 , 
		\3372_b1 , \3372_b0 , \3373_b1 , \3373_b0 , \3374_b1 , \3374_b0 , \3375_b1 , \3375_b0 , \3376_b1 , \3376_b0 , 
		\3377_b1 , \3377_b0 , \3378_b1 , \3378_b0 , \3379_b1 , \3379_b0 , \3380_b1 , \3380_b0 , \3381_b1 , \3381_b0 , 
		\3382_b1 , \3382_b0 , \3383_b1 , \3383_b0 , \3384_b1 , \3384_b0 , \3385_b1 , \3385_b0 , \3386_b1 , \3386_b0 , 
		\3387_b1 , \3387_b0 , \3388_b1 , \3388_b0 , \3389_b1 , \3389_b0 , \3390_b1 , \3390_b0 , \3391_b1 , \3391_b0 , 
		\3392_b1 , \3392_b0 , \3393_b1 , \3393_b0 , \3394_b1 , \3394_b0 , \3395_b1 , \3395_b0 , \3396_b1 , \3396_b0 , 
		\3397_b1 , \3397_b0 , \3398_b1 , \3398_b0 , \3399_b1 , \3399_b0 , \3400_b1 , \3400_b0 , \3401_b1 , \3401_b0 , 
		\3402_b1 , \3402_b0 , \3403_b1 , \3403_b0 , \3404_b1 , \3404_b0 , \3405_b1 , \3405_b0 , \3406_b1 , \3406_b0 , 
		\3407_b1 , \3407_b0 , \3408_b1 , \3408_b0 , \3409_b1 , \3409_b0 , \3410_b1 , \3410_b0 , \3411_b1 , \3411_b0 , 
		\3412_b1 , \3412_b0 , \3413_b1 , \3413_b0 , \3414_b1 , \3414_b0 , \3415_b1 , \3415_b0 , \3416_b1 , \3416_b0 , 
		\3417_b1 , \3417_b0 , \3418_b1 , \3418_b0 , \3419_b1 , \3419_b0 , \3420_b1 , \3420_b0 , \3421_b1 , \3421_b0 , 
		\3422_b1 , \3422_b0 , \3423_b1 , \3423_b0 , \3424_b1 , \3424_b0 , \3425_b1 , \3425_b0 , \3426_b1 , \3426_b0 , 
		\3427_b1 , \3427_b0 , \3428_b1 , \3428_b0 , \3429_b1 , \3429_b0 , \3430_b1 , \3430_b0 , \3431_b1 , \3431_b0 , 
		\3432_b1 , \3432_b0 , \3433_b1 , \3433_b0 , \3434_b1 , \3434_b0 , \3435_b1 , \3435_b0 , \3436_b1 , \3436_b0 , 
		\3437_b1 , \3437_b0 , \3438_b1 , \3438_b0 , \3439_b1 , \3439_b0 , \3440_b1 , \3440_b0 , \3441_b1 , \3441_b0 , 
		\3442_b1 , \3442_b0 , \3443_b1 , \3443_b0 , \3444_b1 , \3444_b0 , \3445_b1 , \3445_b0 , \3446_b1 , \3446_b0 , 
		\3447_b1 , \3447_b0 , \3448_b1 , \3448_b0 , \3449_b1 , \3449_b0 , \3450_b1 , \3450_b0 , \3451_b1 , \3451_b0 , 
		\3452_b1 , \3452_b0 , \3453_b1 , \3453_b0 , \3454_b1 , \3454_b0 , \3455_b1 , \3455_b0 , \3456_b1 , \3456_b0 , 
		\3457_b1 , \3457_b0 , \3458_b1 , \3458_b0 , \3459_b1 , \3459_b0 , \3460_b1 , \3460_b0 , \3461_b1 , \3461_b0 , 
		\3462_b1 , \3462_b0 , \3463_b1 , \3463_b0 , \3464_b1 , \3464_b0 , \3465_b1 , \3465_b0 , \3466_b1 , \3466_b0 , 
		\3467_b1 , \3467_b0 , \3468_b1 , \3468_b0 , \3469_b1 , \3469_b0 , \3470_b1 , \3470_b0 , \3471_b1 , \3471_b0 , 
		\3472_b1 , \3472_b0 , \3473_b1 , \3473_b0 , \3474_b1 , \3474_b0 , \3475_b1 , \3475_b0 , \3476_b1 , \3476_b0 , 
		\3477_b1 , \3477_b0 , \3478_b1 , \3478_b0 , \3479_b1 , \3479_b0 , \3480_b1 , \3480_b0 , \3481_b1 , \3481_b0 , 
		\3482_b1 , \3482_b0 , \3483_b1 , \3483_b0 , \3484_b1 , \3484_b0 , \3485_b1 , \3485_b0 , \3486_b1 , \3486_b0 , 
		\3487_b1 , \3487_b0 , \3488_b1 , \3488_b0 , \3489_b1 , \3489_b0 , \3490_b1 , \3490_b0 , \3491_b1 , \3491_b0 , 
		\3492_b1 , \3492_b0 , \3493_b1 , \3493_b0 , \3494_b1 , \3494_b0 , \3495_b1 , \3495_b0 , \3496_b1 , \3496_b0 , 
		\3497_b1 , \3497_b0 , \3498_b1 , \3498_b0 , \3499_b1 , \3499_b0 , \3500_b1 , \3500_b0 , \3501_b1 , \3501_b0 , 
		\3502_b1 , \3502_b0 , \3503_b1 , \3503_b0 , \3504_b1 , \3504_b0 , \3505_b1 , \3505_b0 , \3506_b1 , \3506_b0 , 
		\3507_b1 , \3507_b0 , \3508_b1 , \3508_b0 , \3509_b1 , \3509_b0 , \3510_b1 , \3510_b0 , \3511_b1 , \3511_b0 , 
		\3512_b1 , \3512_b0 , \3513_b1 , \3513_b0 , \3514_b1 , \3514_b0 , \3515_b1 , \3515_b0 , \3516_b1 , \3516_b0 , 
		\3517_b1 , \3517_b0 , \3518_b1 , \3518_b0 , \3519_b1 , \3519_b0 , \3520_b1 , \3520_b0 , \3521_b1 , \3521_b0 , 
		\3522_b1 , \3522_b0 , \3523_b1 , \3523_b0 , \3524_b1 , \3524_b0 , \3525_b1 , \3525_b0 , \3526_b1 , \3526_b0 , 
		\3527_b1 , \3527_b0 , \3528_b1 , \3528_b0 , \3529_b1 , \3529_b0 , \3530_b1 , \3530_b0 , \3531_b1 , \3531_b0 , 
		\3532_b1 , \3532_b0 , \3533_b1 , \3533_b0 , \3534_b1 , \3534_b0 , \3535_b1 , \3535_b0 , \3536_b1 , \3536_b0 , 
		\3537_b1 , \3537_b0 , \3538_b1 , \3538_b0 , \3539_b1 , \3539_b0 , \3540_b1 , \3540_b0 , \3541_b1 , \3541_b0 , 
		\3542_b1 , \3542_b0 , \3543_b1 , \3543_b0 , \3544_b1 , \3544_b0 , \3545_b1 , \3545_b0 , \3546_b1 , \3546_b0 , 
		\3547_b1 , \3547_b0 , \3548_b1 , \3548_b0 , \3549_b1 , \3549_b0 , \3550_b1 , \3550_b0 , \3551_b1 , \3551_b0 , 
		\3552_b1 , \3552_b0 , \3553_b1 , \3553_b0 , \3554_b1 , \3554_b0 , \3555_b1 , \3555_b0 , \3556_b1 , \3556_b0 , 
		\3557_b1 , \3557_b0 , \3558_b1 , \3558_b0 , \3559_b1 , \3559_b0 , \3560_b1 , \3560_b0 , \3561_b1 , \3561_b0 , 
		\3562_b1 , \3562_b0 , \3563_b1 , \3563_b0 , \3564_b1 , \3564_b0 , \3565_b1 , \3565_b0 , \3566_b1 , \3566_b0 , 
		\3567_b1 , \3567_b0 , \3568_b1 , \3568_b0 , \3569_b1 , \3569_b0 , \3570_b1 , \3570_b0 , \3571_b1 , \3571_b0 , 
		\3572_b1 , \3572_b0 , \3573_b1 , \3573_b0 , \3574_b1 , \3574_b0 , \3575_b1 , \3575_b0 , \3576_b1 , \3576_b0 , 
		\3577_b1 , \3577_b0 , \3578_b1 , \3578_b0 , \3579_b1 , \3579_b0 , \3580_b1 , \3580_b0 , \3581_b1 , \3581_b0 , 
		\3582_b1 , \3582_b0 , \3583_b1 , \3583_b0 , \3584_b1 , \3584_b0 , \3585_b1 , \3585_b0 , \3586_b1 , \3586_b0 , 
		\3587_b1 , \3587_b0 , \3588_b1 , \3588_b0 , \3589_b1 , \3589_b0 , \3590_b1 , \3590_b0 , \3591_b1 , \3591_b0 , 
		\3592_b1 , \3592_b0 , \3593_b1 , \3593_b0 , \3594_b1 , \3594_b0 , \3595_b1 , \3595_b0 , \3596_b1 , \3596_b0 , 
		\3597_b1 , \3597_b0 , \3598_b1 , \3598_b0 , \3599_b1 , \3599_b0 , \3600_b1 , \3600_b0 , \3601_b1 , \3601_b0 , 
		\3602_b1 , \3602_b0 , \3603_b1 , \3603_b0 , \3604_b1 , \3604_b0 , \3605_b1 , \3605_b0 , \3606_b1 , \3606_b0 , 
		\3607_b1 , \3607_b0 , \3608_b1 , \3608_b0 , \3609_b1 , \3609_b0 , \3610_b1 , \3610_b0 , \3611_b1 , \3611_b0 , 
		\3612_b1 , \3612_b0 , \3613_b1 , \3613_b0 , \3614_b1 , \3614_b0 , \3615_b1 , \3615_b0 , \3616_b1 , \3616_b0 , 
		\3617_b1 , \3617_b0 , \3618_b1 , \3618_b0 , \3619_b1 , \3619_b0 , \3620_b1 , \3620_b0 , \3621_b1 , \3621_b0 , 
		\3622_b1 , \3622_b0 , \3623_b1 , \3623_b0 , \3624_b1 , \3624_b0 , \3625_b1 , \3625_b0 , \3626_b1 , \3626_b0 , 
		\3627_b1 , \3627_b0 , \3628_b1 , \3628_b0 , \3629_b1 , \3629_b0 , \3630_b1 , \3630_b0 , \3631_b1 , \3631_b0 , 
		\3632_b1 , \3632_b0 , \3633_b1 , \3633_b0 , \3634_b1 , \3634_b0 , \3635_b1 , \3635_b0 , \3636_b1 , \3636_b0 , 
		\3637_b1 , \3637_b0 , \3638_b1 , \3638_b0 , \3639_b1 , \3639_b0 , \3640_b1 , \3640_b0 , \3641_b1 , \3641_b0 , 
		\3642_b1 , \3642_b0 , \3643_b1 , \3643_b0 , \3644_b1 , \3644_b0 , \3645_b1 , \3645_b0 , \3646_b1 , \3646_b0 , 
		\3647_b1 , \3647_b0 , \3648_b1 , \3648_b0 , \3649_b1 , \3649_b0 , \3650_b1 , \3650_b0 , \3651_b1 , \3651_b0 , 
		\3652_b1 , \3652_b0 , \3653_b1 , \3653_b0 , \3654_b1 , \3654_b0 , \3655_b1 , \3655_b0 , \3656_b1 , \3656_b0 , 
		\3657_b1 , \3657_b0 , \3658_b1 , \3658_b0 , \3659_b1 , \3659_b0 , \3660_b1 , \3660_b0 , \3661_b1 , \3661_b0 , 
		\3662_b1 , \3662_b0 , \3663_b1 , \3663_b0 , \3664_b1 , \3664_b0 , \3665_b1 , \3665_b0 , \3666_b1 , \3666_b0 , 
		\3667_b1 , \3667_b0 , \3668_b1 , \3668_b0 , \3669_b1 , \3669_b0 , \3670_b1 , \3670_b0 , \3671_b1 , \3671_b0 , 
		\3672_b1 , \3672_b0 , \3673_b1 , \3673_b0 , \3674_b1 , \3674_b0 , \3675_b1 , \3675_b0 , \3676_b1 , \3676_b0 , 
		\3677_b1 , \3677_b0 , \3678_b1 , \3678_b0 , \3679_b1 , \3679_b0 , \3680_b1 , \3680_b0 , \3681_b1 , \3681_b0 , 
		\3682_b1 , \3682_b0 , \3683_b1 , \3683_b0 , \3684_b1 , \3684_b0 , \3685_b1 , \3685_b0 , \3686_b1 , \3686_b0 , 
		\3687_b1 , \3687_b0 , \3688_b1 , \3688_b0 , \3689_b1 , \3689_b0 , \3690_b1 , \3690_b0 , \3691_b1 , \3691_b0 , 
		\3692_b1 , \3692_b0 , \3693_b1 , \3693_b0 , \3694_b1 , \3694_b0 , \3695_b1 , \3695_b0 , \3696_b1 , \3696_b0 , 
		\3697_b1 , \3697_b0 , \3698_b1 , \3698_b0 , \3699_b1 , \3699_b0 , \3700_b1 , \3700_b0 , \3701_b1 , \3701_b0 , 
		\3702_b1 , \3702_b0 , \3703_b1 , \3703_b0 , \3704_b1 , \3704_b0 , \3705_b1 , \3705_b0 , \3706_b1 , \3706_b0 , 
		\3707_b1 , \3707_b0 , \3708_b1 , \3708_b0 , \3709_b1 , \3709_b0 , \3710_b1 , \3710_b0 , \3711_b1 , \3711_b0 , 
		\3712_b1 , \3712_b0 , \3713_b1 , \3713_b0 , \3714_b1 , \3714_b0 , \3715_b1 , \3715_b0 , \3716_b1 , \3716_b0 , 
		\3717_b1 , \3717_b0 , \3718_b1 , \3718_b0 , \3719_b1 , \3719_b0 , \3720_b1 , \3720_b0 , \3721_b1 , \3721_b0 , 
		\3722_b1 , \3722_b0 , \3723_b1 , \3723_b0 , \3724_b1 , \3724_b0 , \3725_b1 , \3725_b0 , \3726_b1 , \3726_b0 , 
		\3727_b1 , \3727_b0 , \3728_b1 , \3728_b0 , \3729_b1 , \3729_b0 , \3730_b1 , \3730_b0 , \3731_b1 , \3731_b0 , 
		\3732_b1 , \3732_b0 , \3733_b1 , \3733_b0 , \3734_b1 , \3734_b0 , \3735_b1 , \3735_b0 , \3736_b1 , \3736_b0 , 
		\3737_b1 , \3737_b0 , \3738_b1 , \3738_b0 , \3739_b1 , \3739_b0 , \3740_b1 , \3740_b0 , \3741_b1 , \3741_b0 , 
		\3742_b1 , \3742_b0 , \3743_b1 , \3743_b0 , \3744_b1 , \3744_b0 , \3745_b1 , \3745_b0 , \3746_b1 , \3746_b0 , 
		\3747_b1 , \3747_b0 , \3748_b1 , \3748_b0 , \3749_b1 , \3749_b0 , \3750_b1 , \3750_b0 , \3751_b1 , \3751_b0 , 
		\3752_b1 , \3752_b0 , \3753_b1 , \3753_b0 , \3754_b1 , \3754_b0 , \3755_b1 , \3755_b0 , \3756_b1 , \3756_b0 , 
		\3757_b1 , \3757_b0 , \3758_b1 , \3758_b0 , \3759_b1 , \3759_b0 , \3760_b1 , \3760_b0 , \3761_b1 , \3761_b0 , 
		\3762_b1 , \3762_b0 , \3763_b1 , \3763_b0 , \3764_b1 , \3764_b0 , \3765_b1 , \3765_b0 , \3766_b1 , \3766_b0 , 
		\3767_b1 , \3767_b0 , \3768_b1 , \3768_b0 , \3769_b1 , \3769_b0 , \3770_b1 , \3770_b0 , \3771_b1 , \3771_b0 , 
		\3772_b1 , \3772_b0 , \3773_b1 , \3773_b0 , \3774_b1 , \3774_b0 , \3775_b1 , \3775_b0 , \3776_b1 , \3776_b0 , 
		\3777_b1 , \3777_b0 , \3778_b1 , \3778_b0 , \3779_b1 , \3779_b0 , \3780_b1 , \3780_b0 , \3781_b1 , \3781_b0 , 
		\3782_b1 , \3782_b0 , \3783_b1 , \3783_b0 , \3784_b1 , \3784_b0 , \3785_b1 , \3785_b0 , \3786_b1 , \3786_b0 , 
		\3787_b1 , \3787_b0 , \3788_b1 , \3788_b0 , \3789_b1 , \3789_b0 , \3790_b1 , \3790_b0 , \3791_b1 , \3791_b0 , 
		\3792_b1 , \3792_b0 , \3793_b1 , \3793_b0 , \3794_b1 , \3794_b0 , \3795_b1 , \3795_b0 , \3796_b1 , \3796_b0 , 
		\3797_b1 , \3797_b0 , \3798_b1 , \3798_b0 , \3799_b1 , \3799_b0 , \3800_b1 , \3800_b0 , \3801_b1 , \3801_b0 , 
		\3802_b1 , \3802_b0 , \3803_b1 , \3803_b0 , \3804_b1 , \3804_b0 , \3805_b1 , \3805_b0 , \3806_b1 , \3806_b0 , 
		\3807_b1 , \3807_b0 , \3808_b1 , \3808_b0 , \3809_b1 , \3809_b0 , \3810_b1 , \3810_b0 , \3811_b1 , \3811_b0 , 
		\3812_b1 , \3812_b0 , \3813_b1 , \3813_b0 , \3814_b1 , \3814_b0 , \3815_b1 , \3815_b0 , \3816_b1 , \3816_b0 , 
		\3817_b1 , \3817_b0 , \3818_b1 , \3818_b0 , \3819_b1 , \3819_b0 , \3820_b1 , \3820_b0 , \3821_b1 , \3821_b0 , 
		\3822_b1 , \3822_b0 , \3823_b1 , \3823_b0 , \3824_b1 , \3824_b0 , \3825_b1 , \3825_b0 , \3826_b1 , \3826_b0 , 
		\3827_b1 , \3827_b0 , \3828_b1 , \3828_b0 , \3829_b1 , \3829_b0 , \3830_b1 , \3830_b0 , \3831_b1 , \3831_b0 , 
		\3832_b1 , \3832_b0 , \3833_b1 , \3833_b0 , \3834_b1 , \3834_b0 , \3835_b1 , \3835_b0 , \3836_b1 , \3836_b0 , 
		\3837_b1 , \3837_b0 , \3838_b1 , \3838_b0 , \3839_b1 , \3839_b0 , \3840_b1 , \3840_b0 , \3841_b1 , \3841_b0 , 
		\3842_b1 , \3842_b0 , \3843_b1 , \3843_b0 , \3844_b1 , \3844_b0 , \3845_b1 , \3845_b0 , \3846_b1 , \3846_b0 , 
		\3847_b1 , \3847_b0 , \3848_b1 , \3848_b0 , \3849_b1 , \3849_b0 , \3850_b1 , \3850_b0 , \3851_b1 , \3851_b0 , 
		\3852_b1 , \3852_b0 , \3853_b1 , \3853_b0 , \3854_b1 , \3854_b0 , \3855_b1 , \3855_b0 , \3856_b1 , \3856_b0 , 
		\3857_b1 , \3857_b0 , \3858_b1 , \3858_b0 , \3859_b1 , \3859_b0 , \3860_b1 , \3860_b0 , \3861_b1 , \3861_b0 , 
		\3862_b1 , \3862_b0 , \3863_b1 , \3863_b0 , \3864_b1 , \3864_b0 , \3865_b1 , \3865_b0 , \3866_b1 , \3866_b0 , 
		\3867_b1 , \3867_b0 , \3868_b1 , \3868_b0 , \3869_b1 , \3869_b0 , \3870_b1 , \3870_b0 , \3871_b1 , \3871_b0 , 
		\3872_b1 , \3872_b0 , \3873_b1 , \3873_b0 , \3874_b1 , \3874_b0 , \3875_b1 , \3875_b0 , \3876_b1 , \3876_b0 , 
		\3877_b1 , \3877_b0 , \3878_b1 , \3878_b0 , \3879_b1 , \3879_b0 , \3880_b1 , \3880_b0 , \3881_b1 , \3881_b0 , 
		\3882_b1 , \3882_b0 , \3883_b1 , \3883_b0 , \3884_b1 , \3884_b0 , \3885_b1 , \3885_b0 , \3886_b1 , \3886_b0 , 
		\3887_b1 , \3887_b0 , \3888_b1 , \3888_b0 , \3889_b1 , \3889_b0 , \3890_b1 , \3890_b0 , \3891_b1 , \3891_b0 , 
		\3892_b1 , \3892_b0 , \3893_b1 , \3893_b0 , \3894_b1 , \3894_b0 , \3895_b1 , \3895_b0 , \3896_b1 , \3896_b0 , 
		\3897_b1 , \3897_b0 , \3898_b1 , \3898_b0 , \3899_b1 , \3899_b0 , \3900_b1 , \3900_b0 , \3901_b1 , \3901_b0 , 
		\3902_b1 , \3902_b0 , \3903_b1 , \3903_b0 , \3904_b1 , \3904_b0 , \3905_b1 , \3905_b0 , \3906_b1 , \3906_b0 , 
		\3907_b1 , \3907_b0 , \3908_b1 , \3908_b0 , \3909_b1 , \3909_b0 , \3910_b1 , \3910_b0 , \3911_b1 , \3911_b0 , 
		\3912_b1 , \3912_b0 , \3913_b1 , \3913_b0 , \3914_b1 , \3914_b0 , \3915_b1 , \3915_b0 , \3916_b1 , \3916_b0 , 
		\3917_b1 , \3917_b0 , \3918_b1 , \3918_b0 , \3919_b1 , \3919_b0 , \3920_b1 , \3920_b0 , \3921_b1 , \3921_b0 , 
		\3922_b1 , \3922_b0 , \3923_b1 , \3923_b0 , \3924_b1 , \3924_b0 , \3925_b1 , \3925_b0 , \3926_b1 , \3926_b0 , 
		\3927_b1 , \3927_b0 , \3928_b1 , \3928_b0 , \3929_b1 , \3929_b0 , \3930_b1 , \3930_b0 , \3931_b1 , \3931_b0 , 
		\3932_b1 , \3932_b0 , \3933_b1 , \3933_b0 , \3934_b1 , \3934_b0 , \3935_b1 , \3935_b0 , \3936_b1 , \3936_b0 , 
		\3937_b1 , \3937_b0 , \3938_b1 , \3938_b0 , \3939_b1 , \3939_b0 , \3940_b1 , \3940_b0 , \3941_b1 , \3941_b0 , 
		\3942_b1 , \3942_b0 , \3943_b1 , \3943_b0 , \3944_b1 , \3944_b0 , \3945_b1 , \3945_b0 , \3946_b1 , \3946_b0 , 
		\3947_b1 , \3947_b0 , \3948_b1 , \3948_b0 , \3949_b1 , \3949_b0 , \3950_b1 , \3950_b0 , \3951_b1 , \3951_b0 , 
		\3952_b1 , \3952_b0 , \3953_b1 , \3953_b0 , \3954_b1 , \3954_b0 , \3955_b1 , \3955_b0 , \3956_b1 , \3956_b0 , 
		\3957_b1 , \3957_b0 , \3958_b1 , \3958_b0 , \3959_b1 , \3959_b0 , \3960_b1 , \3960_b0 , \3961_b1 , \3961_b0 , 
		\3962_b1 , \3962_b0 , \3963_b1 , \3963_b0 , \3964_b1 , \3964_b0 , \3965_b1 , \3965_b0 , \3966_b1 , \3966_b0 , 
		\3967_b1 , \3967_b0 , \3968_b1 , \3968_b0 , \3969_b1 , \3969_b0 , \3970_b1 , \3970_b0 , \3971_b1 , \3971_b0 , 
		\3972_b1 , \3972_b0 , \3973_b1 , \3973_b0 , \3974_b1 , \3974_b0 , \3975_b1 , \3975_b0 , \3976_b1 , \3976_b0 , 
		\3977_b1 , \3977_b0 , \3978_b1 , \3978_b0 , \3979_b1 , \3979_b0 , \3980_b1 , \3980_b0 , \3981_b1 , \3981_b0 , 
		\3982_b1 , \3982_b0 , \3983_b1 , \3983_b0 , \3984_b1 , \3984_b0 , \3985_b1 , \3985_b0 , \3986_b1 , \3986_b0 , 
		\3987_b1 , \3987_b0 , \3988_b1 , \3988_b0 , \3989_b1 , \3989_b0 , \3990_b1 , \3990_b0 , \3991_b1 , \3991_b0 , 
		\3992_b1 , \3992_b0 , \3993_b1 , \3993_b0 , \3994_b1 , \3994_b0 , \3995_b1 , \3995_b0 , \3996_b1 , \3996_b0 , 
		\3997_b1 , \3997_b0 , \3998_b1 , \3998_b0 , \3999_b1 , \3999_b0 , \4000_b1 , \4000_b0 , \4001_b1 , \4001_b0 , 
		\4002_b1 , \4002_b0 , \4003_b1 , \4003_b0 , \4004_b1 , \4004_b0 , \4005_b1 , \4005_b0 , \4006_b1 , \4006_b0 , 
		\4007_b1 , \4007_b0 , \4008_b1 , \4008_b0 , \4009_b1 , \4009_b0 , \4010_b1 , \4010_b0 , \4011_b1 , \4011_b0 , 
		\4012_b1 , \4012_b0 , \4013_b1 , \4013_b0 , \4014_b1 , \4014_b0 , \4015_b1 , \4015_b0 , \4016_b1 , \4016_b0 , 
		\4017_b1 , \4017_b0 , \4018_b1 , \4018_b0 , \4019_b1 , \4019_b0 , \4020_b1 , \4020_b0 , \4021_b1 , \4021_b0 , 
		\4022_b1 , \4022_b0 , \4023_b1 , \4023_b0 , \4024_b1 , \4024_b0 , \4025_b1 , \4025_b0 , \4026_b1 , \4026_b0 , 
		\4027_b1 , \4027_b0 , \4028_b1 , \4028_b0 , \4029_b1 , \4029_b0 , \4030_b1 , \4030_b0 , \4031_b1 , \4031_b0 , 
		\4032_b1 , \4032_b0 , \4033_b1 , \4033_b0 , \4034_b1 , \4034_b0 , \4035_b1 , \4035_b0 , \4036_b1 , \4036_b0 , 
		\4037_b1 , \4037_b0 , \4038_b1 , \4038_b0 , \4039_b1 , \4039_b0 , \4040_b1 , \4040_b0 , \4041_b1 , \4041_b0 , 
		\4042_b1 , \4042_b0 , \4043_b1 , \4043_b0 , \4044_b1 , \4044_b0 , \4045_b1 , \4045_b0 , \4046_b1 , \4046_b0 , 
		\4047_b1 , \4047_b0 , \4048_b1 , \4048_b0 , \4049_b1 , \4049_b0 , \4050_b1 , \4050_b0 , \4051_b1 , \4051_b0 , 
		\4052_b1 , \4052_b0 , \4053_b1 , \4053_b0 , \4054_b1 , \4054_b0 , \4055_b1 , \4055_b0 , \4056_b1 , \4056_b0 , 
		\4057_b1 , \4057_b0 , \4058_b1 , \4058_b0 , \4059_b1 , \4059_b0 , \4060_b1 , \4060_b0 , \4061_b1 , \4061_b0 , 
		\4062_b1 , \4062_b0 , \4063_b1 , \4063_b0 , \4064_b1 , \4064_b0 , \4065_b1 , \4065_b0 , \4066_b1 , \4066_b0 , 
		\4067_b1 , \4067_b0 , \4068_b1 , \4068_b0 , \4069_b1 , \4069_b0 , \4070_b1 , \4070_b0 , \4071_b1 , \4071_b0 , 
		\4072_b1 , \4072_b0 , \4073_b1 , \4073_b0 , \4074_b1 , \4074_b0 , \4075_b1 , \4075_b0 , \4076_b1 , \4076_b0 , 
		\4077_b1 , \4077_b0 , \4078_b1 , \4078_b0 , \4079_b1 , \4079_b0 , \4080_b1 , \4080_b0 , \4081_b1 , \4081_b0 , 
		\4082_b1 , \4082_b0 , \4083_b1 , \4083_b0 , \4084_b1 , \4084_b0 , \4085_b1 , \4085_b0 , \4086_b1 , \4086_b0 , 
		\4087_b1 , \4087_b0 , \4088_b1 , \4088_b0 , \4089_b1 , \4089_b0 , \4090_b1 , \4090_b0 , \4091_b1 , \4091_b0 , 
		\4092_b1 , \4092_b0 , \4093_b1 , \4093_b0 , \4094_b1 , \4094_b0 , \4095_b1 , \4095_b0 , \4096_b1 , \4096_b0 , 
		\4097_b1 , \4097_b0 , \4098_b1 , \4098_b0 , \4099_b1 , \4099_b0 , \4100_b1 , \4100_b0 , \4101_b1 , \4101_b0 , 
		\4102_b1 , \4102_b0 , \4103_b1 , \4103_b0 , \4104_b1 , \4104_b0 , \4105_b1 , \4105_b0 , \4106_b1 , \4106_b0 , 
		\4107_b1 , \4107_b0 , \4108_b1 , \4108_b0 , \4109_b1 , \4109_b0 , \4110_b1 , \4110_b0 , \4111_b1 , \4111_b0 , 
		\4112_b1 , \4112_b0 , \4113_b1 , \4113_b0 , \4114_b1 , \4114_b0 , \4115_b1 , \4115_b0 , \4116_b1 , \4116_b0 , 
		\4117_b1 , \4117_b0 , \4118_b1 , \4118_b0 , \4119_b1 , \4119_b0 , \4120_b1 , \4120_b0 , \4121_b1 , \4121_b0 , 
		\4122_b1 , \4122_b0 , \4123_b1 , \4123_b0 , \4124_b1 , \4124_b0 , \4125_b1 , \4125_b0 , \4126_b1 , \4126_b0 , 
		\4127_b1 , \4127_b0 , \4128_b1 , \4128_b0 , \4129_b1 , \4129_b0 , \4130_b1 , \4130_b0 , \4131_b1 , \4131_b0 , 
		\4132_b1 , \4132_b0 , \4133_b1 , \4133_b0 , \4134_b1 , \4134_b0 , \4135_b1 , \4135_b0 , \4136_b1 , \4136_b0 , 
		\4137_b1 , \4137_b0 , \4138_b1 , \4138_b0 , \4139_b1 , \4139_b0 , \4140_b1 , \4140_b0 , \4141_b1 , \4141_b0 , 
		\4142_b1 , \4142_b0 , \4143_b1 , \4143_b0 , \4144_b1 , \4144_b0 , \4145_b1 , \4145_b0 , \4146_b1 , \4146_b0 , 
		\4147_b1 , \4147_b0 , \4148_b1 , \4148_b0 , \4149_b1 , \4149_b0 , \4150_b1 , \4150_b0 , \4151_b1 , \4151_b0 , 
		\4152_b1 , \4152_b0 , \4153_b1 , \4153_b0 , \4154_b1 , \4154_b0 , \4155_b1 , \4155_b0 , \4156_b1 , \4156_b0 , 
		\4157_b1 , \4157_b0 , \4158_b1 , \4158_b0 , \4159_b1 , \4159_b0 , \4160_b1 , \4160_b0 , \4161_b1 , \4161_b0 , 
		\4162_b1 , \4162_b0 , \4163_b1 , \4163_b0 , \4164_b1 , \4164_b0 , \4165_b1 , \4165_b0 , \4166_b1 , \4166_b0 , 
		\4167_b1 , \4167_b0 , \4168_b1 , \4168_b0 , \4169_b1 , \4169_b0 , \4170_b1 , \4170_b0 , \4171_b1 , \4171_b0 , 
		\4172_b1 , \4172_b0 , \4173_b1 , \4173_b0 , \4174_b1 , \4174_b0 , \4175_b1 , \4175_b0 , \4176_b1 , \4176_b0 , 
		\4177_b1 , \4177_b0 , \4178_b1 , \4178_b0 , \4179_b1 , \4179_b0 , \4180_b1 , \4180_b0 , \4181_b1 , \4181_b0 , 
		\4182_b1 , \4182_b0 , \4183_b1 , \4183_b0 , \4184_b1 , \4184_b0 , \4185_b1 , \4185_b0 , \4186_b1 , \4186_b0 , 
		\4187_b1 , \4187_b0 , \4188_b1 , \4188_b0 , \4189_b1 , \4189_b0 , \4190_b1 , \4190_b0 , \4191_b1 , \4191_b0 , 
		\4192_b1 , \4192_b0 , \4193_b1 , \4193_b0 , \4194_b1 , \4194_b0 , \4195_b1 , \4195_b0 , \4196_b1 , \4196_b0 , 
		\4197_b1 , \4197_b0 , \4198_b1 , \4198_b0 , \4199_b1 , \4199_b0 , \4200_b1 , \4200_b0 , \4201_b1 , \4201_b0 , 
		\4202_b1 , \4202_b0 , \4203_b1 , \4203_b0 , \4204_b1 , \4204_b0 , \4205_b1 , \4205_b0 , \4206_b1 , \4206_b0 , 
		\4207_b1 , \4207_b0 , \4208_b1 , \4208_b0 , \4209_b1 , \4209_b0 , \4210_b1 , \4210_b0 , \4211_b1 , \4211_b0 , 
		\4212_b1 , \4212_b0 , \4213_b1 , \4213_b0 , \4214_b1 , \4214_b0 , \4215_b1 , \4215_b0 , \4216_b1 , \4216_b0 , 
		\4217_b1 , \4217_b0 , \4218_b1 , \4218_b0 , \4219_b1 , \4219_b0 , \4220_b1 , \4220_b0 , \4221_b1 , \4221_b0 , 
		\4222_b1 , \4222_b0 , \4223_b1 , \4223_b0 , \4224_b1 , \4224_b0 , \4225_b1 , \4225_b0 , \4226_b1 , \4226_b0 , 
		\4227_b1 , \4227_b0 , \4228_b1 , \4228_b0 , \4229_b1 , \4229_b0 , \4230_b1 , \4230_b0 , \4231_b1 , \4231_b0 , 
		\4232_b1 , \4232_b0 , \4233_b1 , \4233_b0 , \4234_b1 , \4234_b0 , \4235_b1 , \4235_b0 , \4236_b1 , \4236_b0 , 
		\4237_b1 , \4237_b0 , \4238_b1 , \4238_b0 , \4239_b1 , \4239_b0 , \4240_b1 , \4240_b0 , \4241_b1 , \4241_b0 , 
		\4242_b1 , \4242_b0 , \4243_b1 , \4243_b0 , \4244_b1 , \4244_b0 , \4245_b1 , \4245_b0 , \4246_b1 , \4246_b0 , 
		\4247_b1 , \4247_b0 , \4248_b1 , \4248_b0 , \4249_b1 , \4249_b0 , \4250_b1 , \4250_b0 , \4251_b1 , \4251_b0 , 
		\4252_b1 , \4252_b0 , \4253_b1 , \4253_b0 , \4254_b1 , \4254_b0 , \4255_b1 , \4255_b0 , \4256_b1 , \4256_b0 , 
		\4257_b1 , \4257_b0 , \4258_b1 , \4258_b0 , \4259_b1 , \4259_b0 , \4260_b1 , \4260_b0 , \4261_b1 , \4261_b0 , 
		\4262_b1 , \4262_b0 , \4263_b1 , \4263_b0 , \4264_b1 , \4264_b0 , \4265_b1 , \4265_b0 , \4266_b1 , \4266_b0 , 
		\4267_b1 , \4267_b0 , \4268_b1 , \4268_b0 , \4269_b1 , \4269_b0 , \4270_b1 , \4270_b0 , \4271_b1 , \4271_b0 , 
		\4272_b1 , \4272_b0 , \4273_b1 , \4273_b0 , \4274_b1 , \4274_b0 , \4275_b1 , \4275_b0 , \4276_b1 , \4276_b0 , 
		\4277_b1 , \4277_b0 , \4278_b1 , \4278_b0 , \4279_b1 , \4279_b0 , \4280_b1 , \4280_b0 , \4281_b1 , \4281_b0 , 
		\4282_b1 , \4282_b0 , \4283_b1 , \4283_b0 , \4284_b1 , \4284_b0 , \4285_b1 , \4285_b0 , \4286_b1 , \4286_b0 , 
		\4287_b1 , \4287_b0 , \4288_b1 , \4288_b0 , \4289_b1 , \4289_b0 , \4290_b1 , \4290_b0 , \4291_b1 , \4291_b0 , 
		\4292_b1 , \4292_b0 , \4293_b1 , \4293_b0 , \4294_b1 , \4294_b0 , \4295_b1 , \4295_b0 , \4296_b1 , \4296_b0 , 
		\4297_b1 , \4297_b0 , \4298_b1 , \4298_b0 , \4299_b1 , \4299_b0 , \4300_b1 , \4300_b0 , \4301_b1 , \4301_b0 , 
		\4302_b1 , \4302_b0 , \4303_b1 , \4303_b0 , \4304_b1 , \4304_b0 , \4305_b1 , \4305_b0 , \4306_b1 , \4306_b0 , 
		\4307_b1 , \4307_b0 , \4308_b1 , \4308_b0 , \4309_b1 , \4309_b0 , \4310_b1 , \4310_b0 , \4311_b1 , \4311_b0 , 
		\4312_b1 , \4312_b0 , \4313_b1 , \4313_b0 , \4314_b1 , \4314_b0 , \4315_b1 , \4315_b0 , \4316_b1 , \4316_b0 , 
		\4317_b1 , \4317_b0 , \4318_b1 , \4318_b0 , \4319_b1 , \4319_b0 , \4320_b1 , \4320_b0 , \4321_b1 , \4321_b0 , 
		\4322_b1 , \4322_b0 , \4323_b1 , \4323_b0 , \4324_b1 , \4324_b0 , \4325_b1 , \4325_b0 , \4326_b1 , \4326_b0 , 
		\4327_b1 , \4327_b0 , \4328_b1 , \4328_b0 , \4329_b1 , \4329_b0 , \4330_b1 , \4330_b0 , \4331_b1 , \4331_b0 , 
		\4332_b1 , \4332_b0 , \4333_b1 , \4333_b0 , \4334_b1 , \4334_b0 , \4335_b1 , \4335_b0 , \4336_b1 , \4336_b0 , 
		\4337_b1 , \4337_b0 , \4338_b1 , \4338_b0 , \4339_b1 , \4339_b0 , \4340_b1 , \4340_b0 , \4341_b1 , \4341_b0 , 
		\4342_b1 , \4342_b0 , \4343_b1 , \4343_b0 , \4344_b1 , \4344_b0 , \4345_b1 , \4345_b0 , \4346_b1 , \4346_b0 , 
		\4347_b1 , \4347_b0 , \4348_b1 , \4348_b0 , \4349_b1 , \4349_b0 , \4350_b1 , \4350_b0 , \4351_b1 , \4351_b0 , 
		\4352_b1 , \4352_b0 , \4353_b1 , \4353_b0 , \4354_b1 , \4354_b0 , \4355_b1 , \4355_b0 , \4356_b1 , \4356_b0 , 
		\4357_b1 , \4357_b0 , \4358_b1 , \4358_b0 , \4359_b1 , \4359_b0 , \4360_b1 , \4360_b0 , \4361_b1 , \4361_b0 , 
		\4362_b1 , \4362_b0 , \4363_b1 , \4363_b0 , \4364_b1 , \4364_b0 , \4365_b1 , \4365_b0 , \4366_b1 , \4366_b0 , 
		\4367_b1 , \4367_b0 , \4368_b1 , \4368_b0 , \4369_b1 , \4369_b0 , \4370_b1 , \4370_b0 , \4371_b1 , \4371_b0 , 
		\4372_b1 , \4372_b0 , \4373_b1 , \4373_b0 , \4374_b1 , \4374_b0 , \4375_b1 , \4375_b0 , \4376_b1 , \4376_b0 , 
		\4377_b1 , \4377_b0 , \4378_b1 , \4378_b0 , \4379_b1 , \4379_b0 , \4380_b1 , \4380_b0 , \4381_b1 , \4381_b0 , 
		\4382_b1 , \4382_b0 , \4383_b1 , \4383_b0 , \4384_b1 , \4384_b0 , \4385_b1 , \4385_b0 , \4386_b1 , \4386_b0 , 
		\4387_b1 , \4387_b0 , \4388_b1 , \4388_b0 , \4389_b1 , \4389_b0 , \4390_b1 , \4390_b0 , \4391_b1 , \4391_b0 , 
		\4392_b1 , \4392_b0 , \4393_b1 , \4393_b0 , \4394_b1 , \4394_b0 , \4395_b1 , \4395_b0 , \4396_b1 , \4396_b0 , 
		\4397_b1 , \4397_b0 , \4398_b1 , \4398_b0 , \4399_b1 , \4399_b0 , \4400_b1 , \4400_b0 , \4401_b1 , \4401_b0 , 
		\4402_b1 , \4402_b0 , \4403_b1 , \4403_b0 , \4404_b1 , \4404_b0 , \4405_b1 , \4405_b0 , \4406_b1 , \4406_b0 , 
		\4407_b1 , \4407_b0 , \4408_b1 , \4408_b0 , \4409_b1 , \4409_b0 , \4410_b1 , \4410_b0 , \4411_b1 , \4411_b0 , 
		\4412_b1 , \4412_b0 , \4413_b1 , \4413_b0 , \4414_b1 , \4414_b0 , \4415_b1 , \4415_b0 , \4416_b1 , \4416_b0 , 
		\4417_b1 , \4417_b0 , \4418_b1 , \4418_b0 , \4419_b1 , \4419_b0 , \4420_b1 , \4420_b0 , \4421_b1 , \4421_b0 , 
		\4422_b1 , \4422_b0 , \4423_b1 , \4423_b0 , \4424_b1 , \4424_b0 , \4425_b1 , \4425_b0 , \4426_b1 , \4426_b0 , 
		\4427_b1 , \4427_b0 , \4428_b1 , \4428_b0 , \4429_b1 , \4429_b0 , \4430_b1 , \4430_b0 , \4431_b1 , \4431_b0 , 
		\4432_b1 , \4432_b0 , \4433_b1 , \4433_b0 , \4434_b1 , \4434_b0 , \4435_b1 , \4435_b0 , \4436_b1 , \4436_b0 , 
		\4437_b1 , \4437_b0 , \4438_b1 , \4438_b0 , \4439_b1 , \4439_b0 , \4440_b1 , \4440_b0 , \4441_b1 , \4441_b0 , 
		\4442_b1 , \4442_b0 , \4443_b1 , \4443_b0 , \4444_b1 , \4444_b0 , \4445_b1 , \4445_b0 , \4446_b1 , \4446_b0 , 
		\4447_b1 , \4447_b0 , \4448_b1 , \4448_b0 , \4449_b1 , \4449_b0 , \4450_b1 , \4450_b0 , \4451_b1 , \4451_b0 , 
		\4452_b1 , \4452_b0 , \4453_b1 , \4453_b0 , \4454_b1 , \4454_b0 , \4455_b1 , \4455_b0 , \4456_b1 , \4456_b0 , 
		\4457_b1 , \4457_b0 , \4458_b1 , \4458_b0 , \4459_b1 , \4459_b0 , \4460_b1 , \4460_b0 , \4461_b1 , \4461_b0 , 
		\4462_b1 , \4462_b0 , \4463_b1 , \4463_b0 , \4464_b1 , \4464_b0 , \4465_b1 , \4465_b0 , \4466_b1 , \4466_b0 , 
		\4467_b1 , \4467_b0 , \4468_b1 , \4468_b0 , \4469_b1 , \4469_b0 , \4470_b1 , \4470_b0 , \4471_b1 , \4471_b0 , 
		\4472_b1 , \4472_b0 , \4473_b1 , \4473_b0 , \4474_b1 , \4474_b0 , \4475_b1 , \4475_b0 , \4476_b1 , \4476_b0 , 
		\4477_b1 , \4477_b0 , \4478_b1 , \4478_b0 , \4479_b1 , \4479_b0 , \4480_b1 , \4480_b0 , \4481_b1 , \4481_b0 , 
		\4482_b1 , \4482_b0 , \4483_b1 , \4483_b0 , \4484_b1 , \4484_b0 , \4485_b1 , \4485_b0 , \4486_b1 , \4486_b0 , 
		\4487_b1 , \4487_b0 , \4488_b1 , \4488_b0 , \4489_b1 , \4489_b0 , \4490_b1 , \4490_b0 , \4491_b1 , \4491_b0 , 
		\4492_b1 , \4492_b0 , \4493_b1 , \4493_b0 , \4494_b1 , \4494_b0 , \4495_b1 , \4495_b0 , \4496_b1 , \4496_b0 , 
		\4497_b1 , \4497_b0 , \4498_b1 , \4498_b0 , \4499_b1 , \4499_b0 , \4500_b1 , \4500_b0 , \4501_b1 , \4501_b0 , 
		\4502_b1 , \4502_b0 , \4503_b1 , \4503_b0 , \4504_b1 , \4504_b0 , \4505_b1 , \4505_b0 , \4506_b1 , \4506_b0 , 
		\4507_b1 , \4507_b0 , \4508_b1 , \4508_b0 , \4509_b1 , \4509_b0 , \4510_b1 , \4510_b0 , \4511_b1 , \4511_b0 , 
		\4512_b1 , \4512_b0 , \4513_b1 , \4513_b0 , \4514_b1 , \4514_b0 , \4515_b1 , \4515_b0 , \4516_b1 , \4516_b0 , 
		\4517_b1 , \4517_b0 , \4518_b1 , \4518_b0 , \4519_b1 , \4519_b0 , \4520_b1 , \4520_b0 , \4521_b1 , \4521_b0 , 
		\4522_b1 , \4522_b0 , \4523_b1 , \4523_b0 , \4524_b1 , \4524_b0 , \4525_b1 , \4525_b0 , \4526_b1 , \4526_b0 , 
		\4527_b1 , \4527_b0 , \4528_b1 , \4528_b0 , \4529_b1 , \4529_b0 , \4530_b1 , \4530_b0 , \4531_b1 , \4531_b0 , 
		\4532_b1 , \4532_b0 , \4533_b1 , \4533_b0 , \4534_b1 , \4534_b0 , \4535_b1 , \4535_b0 , \4536_b1 , \4536_b0 , 
		\4537_b1 , \4537_b0 , \4538_b1 , \4538_b0 , \4539_b1 , \4539_b0 , \4540_b1 , \4540_b0 , \4541_b1 , \4541_b0 , 
		\4542_b1 , \4542_b0 , \4543_b1 , \4543_b0 , \4544_b1 , \4544_b0 , \4545_b1 , \4545_b0 , \4546_b1 , \4546_b0 , 
		\4547_b1 , \4547_b0 , \4548_b1 , \4548_b0 , \4549_b1 , \4549_b0 , \4550_b1 , \4550_b0 , \4551_b1 , \4551_b0 , 
		\4552_b1 , \4552_b0 , \4553_b1 , \4553_b0 , \4554_b1 , \4554_b0 , \4555_b1 , \4555_b0 , \4556_b1 , \4556_b0 , 
		\4557_b1 , \4557_b0 , \4558_b1 , \4558_b0 , \4559_b1 , \4559_b0 , \4560_b1 , \4560_b0 , \4561_b1 , \4561_b0 , 
		\4562_b1 , \4562_b0 , \4563_b1 , \4563_b0 , \4564_b1 , \4564_b0 , \4565_b1 , \4565_b0 , \4566_b1 , \4566_b0 , 
		\4567_b1 , \4567_b0 , \4568_b1 , \4568_b0 , \4569_b1 , \4569_b0 , \4570_b1 , \4570_b0 , \4571_b1 , \4571_b0 , 
		\4572_b1 , \4572_b0 , \4573_b1 , \4573_b0 , \4574_b1 , \4574_b0 , \4575_b1 , \4575_b0 , \4576_b1 , \4576_b0 , 
		\4577_b1 , \4577_b0 , \4578_b1 , \4578_b0 , \4579_b1 , \4579_b0 , \4580_b1 , \4580_b0 , \4581_b1 , \4581_b0 , 
		\4582_b1 , \4582_b0 , \4583_b1 , \4583_b0 , \4584_b1 , \4584_b0 , \4585_b1 , \4585_b0 , \4586_b1 , \4586_b0 , 
		\4587_b1 , \4587_b0 , \4588_b1 , \4588_b0 , \4589_b1 , \4589_b0 , \4590_b1 , \4590_b0 , \4591_b1 , \4591_b0 , 
		\4592_b1 , \4592_b0 , \4593_b1 , \4593_b0 , \4594_b1 , \4594_b0 , \4595_b1 , \4595_b0 , \4596_b1 , \4596_b0 , 
		\4597_b1 , \4597_b0 , \4598_b1 , \4598_b0 , \4599_b1 , \4599_b0 , \4600_b1 , \4600_b0 , \4601_b1 , \4601_b0 , 
		\4602_b1 , \4602_b0 , \4603_b1 , \4603_b0 , \4604_b1 , \4604_b0 , \4605_b1 , \4605_b0 , \4606_b1 , \4606_b0 , 
		\4607_b1 , \4607_b0 , \4608_b1 , \4608_b0 , \4609_b1 , \4609_b0 , \4610_b1 , \4610_b0 , \4611_b1 , \4611_b0 , 
		\4612_b1 , \4612_b0 , \4613_b1 , \4613_b0 , \4614_b1 , \4614_b0 , \4615_b1 , \4615_b0 , \4616_b1 , \4616_b0 , 
		\4617_b1 , \4617_b0 , \4618_b1 , \4618_b0 , \4619_b1 , \4619_b0 , \4620_b1 , \4620_b0 , \4621_b1 , \4621_b0 , 
		\4622_b1 , \4622_b0 , \4623_b1 , \4623_b0 , \4624_b1 , \4624_b0 , \4625_b1 , \4625_b0 , \4626_b1 , \4626_b0 , 
		\4627_b1 , \4627_b0 , \4628_b1 , \4628_b0 , \4629_b1 , \4629_b0 , \4630_b1 , \4630_b0 , \4631_b1 , \4631_b0 , 
		\4632_b1 , \4632_b0 , \4633_b1 , \4633_b0 , \4634_b1 , \4634_b0 , \4635_b1 , \4635_b0 , \4636_b1 , \4636_b0 , 
		\4637_b1 , \4637_b0 , \4638_b1 , \4638_b0 , \4639_b1 , \4639_b0 , \4640_b1 , \4640_b0 , \4641_b1 , \4641_b0 , 
		\4642_b1 , \4642_b0 , \4643_b1 , \4643_b0 , \4644_b1 , \4644_b0 , \4645_b1 , \4645_b0 , \4646_b1 , \4646_b0 , 
		\4647_b1 , \4647_b0 , \4648_b1 , \4648_b0 , \4649_b1 , \4649_b0 , \4650_b1 , \4650_b0 , \4651_b1 , \4651_b0 , 
		\4652_b1 , \4652_b0 , \4653_b1 , \4653_b0 , \4654_b1 , \4654_b0 , \4655_b1 , \4655_b0 , \4656_b1 , \4656_b0 , 
		\4657_b1 , \4657_b0 , \4658_b1 , \4658_b0 , \4659_b1 , \4659_b0 , \4660_b1 , \4660_b0 , \4661_b1 , \4661_b0 , 
		\4662_b1 , \4662_b0 , \4663_b1 , \4663_b0 , \4664_b1 , \4664_b0 , \4665_b1 , \4665_b0 , \4666_b1 , \4666_b0 , 
		\4667_b1 , \4667_b0 , \4668_b1 , \4668_b0 , \4669_b1 , \4669_b0 , \4670_b1 , \4670_b0 , \4671_b1 , \4671_b0 , 
		\4672_b1 , \4672_b0 , \4673_b1 , \4673_b0 , \4674_b1 , \4674_b0 , \4675_b1 , \4675_b0 , \4676_b1 , \4676_b0 , 
		\4677_b1 , \4677_b0 , \4678_b1 , \4678_b0 , \4679_b1 , \4679_b0 , \4680_b1 , \4680_b0 , \4681_b1 , \4681_b0 , 
		\4682_b1 , \4682_b0 , \4683_b1 , \4683_b0 , \4684_b1 , \4684_b0 , \4685_b1 , \4685_b0 , \4686_b1 , \4686_b0 , 
		\4687_b1 , \4687_b0 , \4688_b1 , \4688_b0 , \4689_b1 , \4689_b0 , \4690_b1 , \4690_b0 , \4691_b1 , \4691_b0 , 
		\4692_b1 , \4692_b0 , \4693_b1 , \4693_b0 , \4694_b1 , \4694_b0 , \4695_b1 , \4695_b0 , \4696_b1 , \4696_b0 , 
		\4697_b1 , \4697_b0 , \4698_b1 , \4698_b0 , \4699_b1 , \4699_b0 , \4700_b1 , \4700_b0 , \4701_b1 , \4701_b0 , 
		\4702_b1 , \4702_b0 , \4703_b1 , \4703_b0 , \4704_b1 , \4704_b0 , \4705_b1 , \4705_b0 , \4706_b1 , \4706_b0 , 
		\4707_b1 , \4707_b0 , \4708_b1 , \4708_b0 , \4709_b1 , \4709_b0 , \4710_b1 , \4710_b0 , \4711_b1 , \4711_b0 , 
		\4712_b1 , \4712_b0 , \4713_b1 , \4713_b0 , \4714_b1 , \4714_b0 , \4715_b1 , \4715_b0 , \4716_b1 , \4716_b0 , 
		\4717_b1 , \4717_b0 , \4718_b1 , \4718_b0 , \4719_b1 , \4719_b0 , \4720_b1 , \4720_b0 , \4721_b1 , \4721_b0 , 
		\4722_b1 , \4722_b0 , \4723_b1 , \4723_b0 , \4724_b1 , \4724_b0 , \4725_b1 , \4725_b0 , \4726_b1 , \4726_b0 , 
		\4727_b1 , \4727_b0 , \4728_b1 , \4728_b0 , \4729_b1 , \4729_b0 , \4730_b1 , \4730_b0 , \4731_b1 , \4731_b0 , 
		\4732_b1 , \4732_b0 , \4733_b1 , \4733_b0 , \4734_b1 , \4734_b0 , \4735_b1 , \4735_b0 , \4736_b1 , \4736_b0 , 
		\4737_b1 , \4737_b0 , \4738_b1 , \4738_b0 , \4739_b1 , \4739_b0 , \4740_b1 , \4740_b0 , \4741_b1 , \4741_b0 , 
		\4742_b1 , \4742_b0 , \4743_b1 , \4743_b0 , \4744_b1 , \4744_b0 , \4745_b1 , \4745_b0 , \4746_b1 , \4746_b0 , 
		\4747_b1 , \4747_b0 , \4748_b1 , \4748_b0 , \4749_b1 , \4749_b0 , \4750_b1 , \4750_b0 , \4751_b1 , \4751_b0 , 
		\4752_b1 , \4752_b0 , \4753_b1 , \4753_b0 , \4754_b1 , \4754_b0 , \4755_b1 , \4755_b0 , \4756_b1 , \4756_b0 , 
		\4757_b1 , \4757_b0 , \4758_b1 , \4758_b0 , \4759_b1 , \4759_b0 , \4760_b1 , \4760_b0 , \4761_b1 , \4761_b0 , 
		\4762_b1 , \4762_b0 , \4763_b1 , \4763_b0 , \4764_b1 , \4764_b0 , \4765_b1 , \4765_b0 , \4766_b1 , \4766_b0 , 
		\4767_b1 , \4767_b0 , \4768_b1 , \4768_b0 , \4769_b1 , \4769_b0 , \4770_b1 , \4770_b0 , \4771_b1 , \4771_b0 , 
		\4772_b1 , \4772_b0 , \4773_b1 , \4773_b0 , \4774_b1 , \4774_b0 , \4775_b1 , \4775_b0 , \4776_b1 , \4776_b0 , 
		\4777_b1 , \4777_b0 , \4778_b1 , \4778_b0 , \4779_b1 , \4779_b0 , \4780_b1 , \4780_b0 , \4781_b1 , \4781_b0 , 
		\4782_b1 , \4782_b0 , \4783_b1 , \4783_b0 , \4784_b1 , \4784_b0 , \4785_b1 , \4785_b0 , \4786_b1 , \4786_b0 , 
		\4787_b1 , \4787_b0 , \4788_b1 , \4788_b0 , \4789_b1 , \4789_b0 , \4790_b1 , \4790_b0 , \4791_b1 , \4791_b0 , 
		\4792_b1 , \4792_b0 , \4793_b1 , \4793_b0 , \4794_b1 , \4794_b0 , \4795_b1 , \4795_b0 , \4796_b1 , \4796_b0 , 
		\4797_b1 , \4797_b0 , \4798_b1 , \4798_b0 , \4799_b1 , \4799_b0 , \4800_b1 , \4800_b0 , \4801_b1 , \4801_b0 , 
		\4802_b1 , \4802_b0 , \4803_b1 , \4803_b0 , \4804_b1 , \4804_b0 , \4805_b1 , \4805_b0 , \4806_b1 , \4806_b0 , 
		\4807_b1 , \4807_b0 , \4808_b1 , \4808_b0 , \4809_b1 , \4809_b0 , \4810_b1 , \4810_b0 , \4811_b1 , \4811_b0 , 
		\4812_b1 , \4812_b0 , \4813_b1 , \4813_b0 , \4814_b1 , \4814_b0 , \4815_b1 , \4815_b0 , \4816_b1 , \4816_b0 , 
		\4817_b1 , \4817_b0 , \4818_b1 , \4818_b0 , \4819_b1 , \4819_b0 , \4820_b1 , \4820_b0 , \4821_b1 , \4821_b0 , 
		\4822_b1 , \4822_b0 , \4823_b1 , \4823_b0 , \4824_b1 , \4824_b0 , \4825_b1 , \4825_b0 , \4826_b1 , \4826_b0 , 
		\4827_b1 , \4827_b0 , \4828_b1 , \4828_b0 , \4829_b1 , \4829_b0 , \4830_b1 , \4830_b0 , \4831_b1 , \4831_b0 , 
		\4832_b1 , \4832_b0 , \4833_b1 , \4833_b0 , \4834_b1 , \4834_b0 , \4835_b1 , \4835_b0 , \4836_b1 , \4836_b0 , 
		\4837_b1 , \4837_b0 , \4838_b1 , \4838_b0 , \4839_b1 , \4839_b0 , \4840_b1 , \4840_b0 , \4841_b1 , \4841_b0 , 
		\4842_b1 , \4842_b0 , \4843_b1 , \4843_b0 , \4844_b1 , \4844_b0 , \4845_b1 , \4845_b0 , \4846_b1 , \4846_b0 , 
		\4847_b1 , \4847_b0 , \4848_b1 , \4848_b0 , \4849_b1 , \4849_b0 , \4850_b1 , \4850_b0 , \4851_b1 , \4851_b0 , 
		\4852_b1 , \4852_b0 , \4853_b1 , \4853_b0 , \4854_b1 , \4854_b0 , \4855_b1 , \4855_b0 , \4856_b1 , \4856_b0 , 
		\4857_b1 , \4857_b0 , \4858_b1 , \4858_b0 , \4859_b1 , \4859_b0 , \4860_b1 , \4860_b0 , \4861_b1 , \4861_b0 , 
		\4862_b1 , \4862_b0 , \4863_b1 , \4863_b0 , \4864_b1 , \4864_b0 , \4865_b1 , \4865_b0 , \4866_b1 , \4866_b0 , 
		\4867_b1 , \4867_b0 , \4868_b1 , \4868_b0 , \4869_b1 , \4869_b0 , \4870_b1 , \4870_b0 , \4871_b1 , \4871_b0 , 
		\4872_b1 , \4872_b0 , \4873_b1 , \4873_b0 , \4874_b1 , \4874_b0 , \4875_b1 , \4875_b0 , \4876_b1 , \4876_b0 , 
		\4877_b1 , \4877_b0 , \4878_b1 , \4878_b0 , \4879_b1 , \4879_b0 , \4880_b1 , \4880_b0 , \4881_b1 , \4881_b0 , 
		\4882_b1 , \4882_b0 , \4883_b1 , \4883_b0 , \4884_b1 , \4884_b0 , \4885_b1 , \4885_b0 , \4886_b1 , \4886_b0 , 
		\4887_b1 , \4887_b0 , \4888_b1 , \4888_b0 , \4889_b1 , \4889_b0 , \4890_b1 , \4890_b0 , \4891_b1 , \4891_b0 , 
		\4892_b1 , \4892_b0 , \4893_b1 , \4893_b0 , \4894_b1 , \4894_b0 , \4895_b1 , \4895_b0 , \4896_b1 , \4896_b0 , 
		\4897_b1 , \4897_b0 , \4898_b1 , \4898_b0 , \4899_b1 , \4899_b0 , \4900_b1 , \4900_b0 , \4901_b1 , \4901_b0 , 
		\4902_b1 , \4902_b0 , \4903_b1 , \4903_b0 , \4904_b1 , \4904_b0 , \4905_b1 , \4905_b0 , \4906_b1 , \4906_b0 , 
		\4907_b1 , \4907_b0 , \4908_b1 , \4908_b0 , \4909_b1 , \4909_b0 , \4910_b1 , \4910_b0 , \4911_b1 , \4911_b0 , 
		\4912_b1 , \4912_b0 , \4913_b1 , \4913_b0 , \4914_b1 , \4914_b0 , \4915_b1 , \4915_b0 , \4916_b1 , \4916_b0 , 
		\4917_b1 , \4917_b0 , \4918_b1 , \4918_b0 , \4919_b1 , \4919_b0 , \4920_b1 , \4920_b0 , \4921_b1 , \4921_b0 , 
		\4922_b1 , \4922_b0 , \4923_b1 , \4923_b0 , \4924_b1 , \4924_b0 , \4925_b1 , \4925_b0 , \4926_b1 , \4926_b0 , 
		\4927_b1 , \4927_b0 , \4928_b1 , \4928_b0 , \4929_b1 , \4929_b0 , \4930_b1 , \4930_b0 , \4931_b1 , \4931_b0 , 
		\4932_b1 , \4932_b0 , \4933_b1 , \4933_b0 , \4934_b1 , \4934_b0 , \4935_b1 , \4935_b0 , \4936_b1 , \4936_b0 , 
		\4937_b1 , \4937_b0 , \4938_b1 , \4938_b0 , \4939_b1 , \4939_b0 , \4940_b1 , \4940_b0 , \4941_b1 , \4941_b0 , 
		\4942_b1 , \4942_b0 , \4943_b1 , \4943_b0 , \4944_b1 , \4944_b0 , \4945_b1 , \4945_b0 , \4946_b1 , \4946_b0 , 
		\4947_b1 , \4947_b0 , \4948_b1 , \4948_b0 , \4949_b1 , \4949_b0 , \4950_b1 , \4950_b0 , \4951_b1 , \4951_b0 , 
		\4952_b1 , \4952_b0 , \4953_b1 , \4953_b0 , \4954_b1 , \4954_b0 , \4955_b1 , \4955_b0 , \4956_b1 , \4956_b0 , 
		\4957_b1 , \4957_b0 , \4958_b1 , \4958_b0 , \4959_b1 , \4959_b0 , \4960_b1 , \4960_b0 , \4961_b1 , \4961_b0 , 
		\4962_b1 , \4962_b0 , \4963_b1 , \4963_b0 , \4964_b1 , \4964_b0 , \4965_b1 , \4965_b0 , \4966_b1 , \4966_b0 , 
		\4967_b1 , \4967_b0 , \4968_b1 , \4968_b0 , \4969_b1 , \4969_b0 , \4970_b1 , \4970_b0 , \4971_b1 , \4971_b0 , 
		\4972_b1 , \4972_b0 , \4973_b1 , \4973_b0 , \4974_b1 , \4974_b0 , \4975_b1 , \4975_b0 , \4976_b1 , \4976_b0 , 
		\4977_b1 , \4977_b0 , \4978_b1 , \4978_b0 , \4979_b1 , \4979_b0 , \4980_b1 , \4980_b0 , \4981_b1 , \4981_b0 , 
		\4982_b1 , \4982_b0 , \4983_b1 , \4983_b0 , \4984_b1 , \4984_b0 , \4985_b1 , \4985_b0 , \4986_b1 , \4986_b0 , 
		\4987_b1 , \4987_b0 , \4988_b1 , \4988_b0 , \4989_b1 , \4989_b0 , \4990_b1 , \4990_b0 , \4991_b1 , \4991_b0 , 
		\4992_b1 , \4992_b0 , \4993_b1 , \4993_b0 , \4994_b1 , \4994_b0 , \4995_b1 , \4995_b0 , \4996_b1 , \4996_b0 , 
		\4997_b1 , \4997_b0 , \4998_b1 , \4998_b0 , \4999_b1 , \4999_b0 , \5000_b1 , \5000_b0 , \5001_b1 , \5001_b0 , 
		\5002_b1 , \5002_b0 , \5003_b1 , \5003_b0 , \5004_b1 , \5004_b0 , \5005_b1 , \5005_b0 , \5006_b1 , \5006_b0 , 
		\5007_b1 , \5007_b0 , \5008_b1 , \5008_b0 , \5009_b1 , \5009_b0 , \5010_b1 , \5010_b0 , \5011_b1 , \5011_b0 , 
		\5012_b1 , \5012_b0 , \5013_b1 , \5013_b0 , \5014_b1 , \5014_b0 , \5015_b1 , \5015_b0 , \5016_b1 , \5016_b0 , 
		\5017_b1 , \5017_b0 , \5018_b1 , \5018_b0 , \5019_b1 , \5019_b0 , \5020_b1 , \5020_b0 , \5021_b1 , \5021_b0 , 
		\5022_b1 , \5022_b0 , \5023_b1 , \5023_b0 , \5024_b1 , \5024_b0 , \5025_b1 , \5025_b0 , \5026_b1 , \5026_b0 , 
		\5027_b1 , \5027_b0 , \5028_b1 , \5028_b0 , \5029_b1 , \5029_b0 , \5030_b1 , \5030_b0 , \5031_b1 , \5031_b0 , 
		\5032_b1 , \5032_b0 , \5033_b1 , \5033_b0 , \5034_b1 , \5034_b0 , \5035_b1 , \5035_b0 , \5036_b1 , \5036_b0 , 
		\5037_b1 , \5037_b0 , \5038_b1 , \5038_b0 , \5039_b1 , \5039_b0 , \5040_b1 , \5040_b0 , \5041_b1 , \5041_b0 , 
		\5042_b1 , \5042_b0 , \5043_b1 , \5043_b0 , \5044_b1 , \5044_b0 , \5045_b1 , \5045_b0 , \5046_b1 , \5046_b0 , 
		\5047_b1 , \5047_b0 , \5048_b1 , \5048_b0 , \5049_b1 , \5049_b0 , \5050_b1 , \5050_b0 , \5051_b1 , \5051_b0 , 
		\5052_b1 , \5052_b0 , \5053_b1 , \5053_b0 , \5054_b1 , \5054_b0 , \5055_b1 , \5055_b0 , \5056_b1 , \5056_b0 , 
		\5057_b1 , \5057_b0 , \5058_b1 , \5058_b0 , \5059_b1 , \5059_b0 , \5060_b1 , \5060_b0 , \5061_b1 , \5061_b0 , 
		\5062_b1 , \5062_b0 , \5063_b1 , \5063_b0 , \5064_b1 , \5064_b0 , \5065_b1 , \5065_b0 , \5066_b1 , \5066_b0 , 
		\5067_b1 , \5067_b0 , \5068_b1 , \5068_b0 , \5069_b1 , \5069_b0 , \5070_b1 , \5070_b0 , \5071_b1 , \5071_b0 , 
		\5072_b1 , \5072_b0 , \5073_b1 , \5073_b0 , \5074_b1 , \5074_b0 , \5075_b1 , \5075_b0 , \5076_b1 , \5076_b0 , 
		\5077_b1 , \5077_b0 , \5078_b1 , \5078_b0 , \5079_b1 , \5079_b0 , \5080_b1 , \5080_b0 , \5081_b1 , \5081_b0 , 
		\5082_b1 , \5082_b0 , \5083_b1 , \5083_b0 , \5084_b1 , \5084_b0 , \5085_b1 , \5085_b0 , \5086_b1 , \5086_b0 , 
		\5087_b1 , \5087_b0 , \5088_b1 , \5088_b0 , \5089_b1 , \5089_b0 , \5090_b1 , \5090_b0 , \5091_b1 , \5091_b0 , 
		\5092_b1 , \5092_b0 , \5093_b1 , \5093_b0 , \5094_b1 , \5094_b0 , \5095_b1 , \5095_b0 , \5096_b1 , \5096_b0 , 
		\5097_b1 , \5097_b0 , \5098_b1 , \5098_b0 , \5099_b1 , \5099_b0 , \5100_b1 , \5100_b0 , \5101_b1 , \5101_b0 , 
		\5102_b1 , \5102_b0 , \5103_b1 , \5103_b0 , \5104_b1 , \5104_b0 , \5105_b1 , \5105_b0 , \5106_b1 , \5106_b0 , 
		\5107_b1 , \5107_b0 , \5108_b1 , \5108_b0 , \5109_b1 , \5109_b0 , \5110_b1 , \5110_b0 , \5111_b1 , \5111_b0 , 
		\5112_b1 , \5112_b0 , \5113_b1 , \5113_b0 , \5114_b1 , \5114_b0 , \5115_b1 , \5115_b0 , \5116_b1 , \5116_b0 , 
		\5117_b1 , \5117_b0 , \5118_b1 , \5118_b0 , \5119_b1 , \5119_b0 , \5120_b1 , \5120_b0 , \5121_b1 , \5121_b0 , 
		\5122_b1 , \5122_b0 , \5123_b1 , \5123_b0 , \5124_b1 , \5124_b0 , \5125_b1 , \5125_b0 , \5126_b1 , \5126_b0 , 
		\5127_b1 , \5127_b0 , \5128_b1 , \5128_b0 , \5129_b1 , \5129_b0 , \5130_b1 , \5130_b0 , \5131_b1 , \5131_b0 , 
		\5132_b1 , \5132_b0 , \5133_b1 , \5133_b0 , \5134_b1 , \5134_b0 , \5135_b1 , \5135_b0 , \5136_b1 , \5136_b0 , 
		\5137_b1 , \5137_b0 , \5138_b1 , \5138_b0 , \5139_b1 , \5139_b0 , \5140_b1 , \5140_b0 , \5141_b1 , \5141_b0 , 
		\5142_b1 , \5142_b0 , \5143_b1 , \5143_b0 , \5144_b1 , \5144_b0 , \5145_b1 , \5145_b0 , \5146_b1 , \5146_b0 , 
		\5147_b1 , \5147_b0 , \5148_b1 , \5148_b0 , \5149_b1 , \5149_b0 , \5150_b1 , \5150_b0 , \5151_b1 , \5151_b0 , 
		\5152_b1 , \5152_b0 , \5153_b1 , \5153_b0 , \5154_b1 , \5154_b0 , \5155_b1 , \5155_b0 , \5156_b1 , \5156_b0 , 
		\5157_b1 , \5157_b0 , \5158_b1 , \5158_b0 , \5159_b1 , \5159_b0 , \5160_b1 , \5160_b0 , \5161_b1 , \5161_b0 , 
		\5162_b1 , \5162_b0 , \5163_b1 , \5163_b0 , \5164_b1 , \5164_b0 , \5165_b1 , \5165_b0 , \5166_b1 , \5166_b0 , 
		\5167_b1 , \5167_b0 , \5168_b1 , \5168_b0 , \5169_b1 , \5169_b0 , \5170_b1 , \5170_b0 , \5171_b1 , \5171_b0 , 
		\5172_b1 , \5172_b0 , \5173_b1 , \5173_b0 , \5174_b1 , \5174_b0 , \5175_b1 , \5175_b0 , \5176_b1 , \5176_b0 , 
		\5177_b1 , \5177_b0 , \5178_b1 , \5178_b0 , \5179_b1 , \5179_b0 , \5180_b1 , \5180_b0 , \5181_b1 , \5181_b0 , 
		\5182_b1 , \5182_b0 , \5183_b1 , \5183_b0 , \5184_b1 , \5184_b0 , \5185_b1 , \5185_b0 , \5186_b1 , \5186_b0 , 
		\5187_b1 , \5187_b0 , \5188_b1 , \5188_b0 , \5189_b1 , \5189_b0 , \5190_b1 , \5190_b0 , \5191_b1 , \5191_b0 , 
		\5192_b1 , \5192_b0 , \5193_b1 , \5193_b0 , \5194_b1 , \5194_b0 , \5195_b1 , \5195_b0 , \5196_b1 , \5196_b0 , 
		\5197_b1 , \5197_b0 , \5198_b1 , \5198_b0 , \5199_b1 , \5199_b0 , \5200_b1 , \5200_b0 , \5201_b1 , \5201_b0 , 
		\5202_b1 , \5202_b0 , \5203_b1 , \5203_b0 , \5204_b1 , \5204_b0 , \5205_b1 , \5205_b0 , \5206_b1 , \5206_b0 , 
		\5207_b1 , \5207_b0 , \5208_b1 , \5208_b0 , \5209_b1 , \5209_b0 , \5210_b1 , \5210_b0 , \5211_b1 , \5211_b0 , 
		\5212_b1 , \5212_b0 , \5213_b1 , \5213_b0 , \5214_b1 , \5214_b0 , \5215_b1 , \5215_b0 , \5216_b1 , \5216_b0 , 
		\5217_b1 , \5217_b0 , \5218_b1 , \5218_b0 , \5219_b1 , \5219_b0 , \5220_b1 , \5220_b0 , \5221_b1 , \5221_b0 , 
		\5222_b1 , \5222_b0 , \5223_b1 , \5223_b0 , \5224_b1 , \5224_b0 , \5225_b1 , \5225_b0 , \5226_b1 , \5226_b0 , 
		\5227_b1 , \5227_b0 , \5228_b1 , \5228_b0 , \5229_b1 , \5229_b0 , \5230_b1 , \5230_b0 , \5231_b1 , \5231_b0 , 
		\5232_b1 , \5232_b0 , \5233_b1 , \5233_b0 , \5234_b1 , \5234_b0 , \5235_b1 , \5235_b0 , \5236_b1 , \5236_b0 , 
		\5237_b1 , \5237_b0 , \5238_b1 , \5238_b0 , \5239_b1 , \5239_b0 , \5240_b1 , \5240_b0 , \5241_b1 , \5241_b0 , 
		\5242_b1 , \5242_b0 , \5243_b1 , \5243_b0 , \5244_b1 , \5244_b0 , \5245_b1 , \5245_b0 , \5246_b1 , \5246_b0 , 
		\5247_b1 , \5247_b0 , \5248_b1 , \5248_b0 , \5249_b1 , \5249_b0 , \5250_b1 , \5250_b0 , \5251_b1 , \5251_b0 , 
		\5252_b1 , \5252_b0 , \5253_b1 , \5253_b0 , \5254_b1 , \5254_b0 , \5255_b1 , \5255_b0 , \5256_b1 , \5256_b0 , 
		\5257_b1 , \5257_b0 , \5258_b1 , \5258_b0 , \5259_b1 , \5259_b0 , \5260_b1 , \5260_b0 , \5261_b1 , \5261_b0 , 
		\5262_b1 , \5262_b0 , \5263_b1 , \5263_b0 , \5264_b1 , \5264_b0 , \5265_b1 , \5265_b0 , \5266_b1 , \5266_b0 , 
		\5267_b1 , \5267_b0 , \5268_b1 , \5268_b0 , \5269_b1 , \5269_b0 , \5270_b1 , \5270_b0 , \5271_b1 , \5271_b0 , 
		\5272_b1 , \5272_b0 , \5273_b1 , \5273_b0 , \5274_b1 , \5274_b0 , \5275_b1 , \5275_b0 , \5276_b1 , \5276_b0 , 
		\5277_b1 , \5277_b0 , \5278_b1 , \5278_b0 , \5279_b1 , \5279_b0 , \5280_b1 , \5280_b0 , \5281_b1 , \5281_b0 , 
		\5282_b1 , \5282_b0 , \5283_b1 , \5283_b0 , \5284_b1 , \5284_b0 , \5285_b1 , \5285_b0 , \5286_b1 , \5286_b0 , 
		\5287_b1 , \5287_b0 , \5288_b1 , \5288_b0 , \5289_b1 , \5289_b0 , \5290_b1 , \5290_b0 , \5291_b1 , \5291_b0 , 
		\5292_b1 , \5292_b0 , \5293_b1 , \5293_b0 , \5294_b1 , \5294_b0 , \5295_b1 , \5295_b0 , \5296_b1 , \5296_b0 , 
		\5297_b1 , \5297_b0 , \5298_b1 , \5298_b0 , \5299_b1 , \5299_b0 , \5300_b1 , \5300_b0 , \5301_b1 , \5301_b0 , 
		\5302_b1 , \5302_b0 , \5303_b1 , \5303_b0 , \5304_b1 , \5304_b0 , \5305_b1 , \5305_b0 , \5306_b1 , \5306_b0 , 
		\5307_b1 , \5307_b0 , \5308_b1 , \5308_b0 , \5309_b1 , \5309_b0 , \5310_b1 , \5310_b0 , \5311_b1 , \5311_b0 , 
		\5312_b1 , \5312_b0 , \5313_b1 , \5313_b0 , \5314_b1 , \5314_b0 , \5315_b1 , \5315_b0 , \5316_b1 , \5316_b0 , 
		\5317_b1 , \5317_b0 , \5318_b1 , \5318_b0 , \5319_b1 , \5319_b0 , \5320_b1 , \5320_b0 , \5321_b1 , \5321_b0 , 
		\5322_b1 , \5322_b0 , \5323_b1 , \5323_b0 , \5324_b1 , \5324_b0 , \5325_b1 , \5325_b0 , \5326_b1 , \5326_b0 , 
		\5327_b1 , \5327_b0 , \5328_b1 , \5328_b0 , \5329_b1 , \5329_b0 , \5330_b1 , \5330_b0 , \5331_b1 , \5331_b0 , 
		\5332_b1 , \5332_b0 , \5333_b1 , \5333_b0 , \5334_b1 , \5334_b0 , \5335_b1 , \5335_b0 , \5336_b1 , \5336_b0 , 
		\5337_b1 , \5337_b0 , \5338_b1 , \5338_b0 , \5339_b1 , \5339_b0 , \5340_b1 , \5340_b0 , \5341_b1 , \5341_b0 , 
		\5342_b1 , \5342_b0 , \5343_b1 , \5343_b0 , \5344_b1 , \5344_b0 , \5345_b1 , \5345_b0 , \5346_b1 , \5346_b0 , 
		\5347_b1 , \5347_b0 , \5348_b1 , \5348_b0 , \5349_b1 , \5349_b0 , \5350_b1 , \5350_b0 , \5351_b1 , \5351_b0 , 
		\5352_b1 , \5352_b0 , \5353_b1 , \5353_b0 , \5354_b1 , \5354_b0 , \5355_b1 , \5355_b0 , \5356_b1 , \5356_b0 , 
		\5357_b1 , \5357_b0 , \5358_b1 , \5358_b0 , \5359_b1 , \5359_b0 , \5360_b1 , \5360_b0 , \5361_b1 , \5361_b0 , 
		\5362_b1 , \5362_b0 , \5363_b1 , \5363_b0 , \5364_b1 , \5364_b0 , \5365_b1 , \5365_b0 , \5366_b1 , \5366_b0 , 
		\5367_b1 , \5367_b0 , \5368_b1 , \5368_b0 , \5369_b1 , \5369_b0 , \5370_b1 , \5370_b0 , \5371_b1 , \5371_b0 , 
		\5372_b1 , \5372_b0 , \5373_b1 , \5373_b0 , \5374_b1 , \5374_b0 , \5375_b1 , \5375_b0 , \5376_b1 , \5376_b0 , 
		\5377_b1 , \5377_b0 , \5378_b1 , \5378_b0 , \5379_b1 , \5379_b0 , \5380_b1 , \5380_b0 , \5381_b1 , \5381_b0 , 
		\5382_b1 , \5382_b0 , \5383_b1 , \5383_b0 , \5384_b1 , \5384_b0 , \5385_b1 , \5385_b0 , \5386_b1 , \5386_b0 , 
		\5387_b1 , \5387_b0 , \5388_b1 , \5388_b0 , \5389_b1 , \5389_b0 , \5390_b1 , \5390_b0 , \5391_b1 , \5391_b0 , 
		\5392_b1 , \5392_b0 , \5393_b1 , \5393_b0 , \5394_b1 , \5394_b0 , \5395_b1 , \5395_b0 , \5396_b1 , \5396_b0 , 
		\5397_b1 , \5397_b0 , \5398_b1 , \5398_b0 , \5399_b1 , \5399_b0 , \5400_b1 , \5400_b0 , \5401_b1 , \5401_b0 , 
		\5402_b1 , \5402_b0 , \5403_b1 , \5403_b0 , \5404_b1 , \5404_b0 , \5405_b1 , \5405_b0 , \5406_b1 , \5406_b0 , 
		\5407_b1 , \5407_b0 , \5408_b1 , \5408_b0 , \5409_b1 , \5409_b0 , \5410_b1 , \5410_b0 , \5411_b1 , \5411_b0 , 
		\5412_b1 , \5412_b0 , \5413_b1 , \5413_b0 , \5414_b1 , \5414_b0 , \5415_b1 , \5415_b0 , \5416_b1 , \5416_b0 , 
		\5417_b1 , \5417_b0 , \5418_b1 , \5418_b0 , \5419_b1 , \5419_b0 , \5420_b1 , \5420_b0 , \5421_b1 , \5421_b0 , 
		\5422_b1 , \5422_b0 , \5423_b1 , \5423_b0 , \5424_b1 , \5424_b0 , \5425_b1 , \5425_b0 , \5426_b1 , \5426_b0 , 
		\5427_b1 , \5427_b0 , \5428_b1 , \5428_b0 , \5429_b1 , \5429_b0 , \5430_b1 , \5430_b0 , \5431_b1 , \5431_b0 , 
		\5432_b1 , \5432_b0 , \5433_b1 , \5433_b0 , \5434_b1 , \5434_b0 , \5435_b1 , \5435_b0 , \5436_b1 , \5436_b0 , 
		\5437_b1 , \5437_b0 , \5438_b1 , \5438_b0 , \5439_b1 , \5439_b0 , \5440_b1 , \5440_b0 , \5441_b1 , \5441_b0 , 
		\5442_b1 , \5442_b0 , \5443_b1 , \5443_b0 , \5444_b1 , \5444_b0 , \5445_b1 , \5445_b0 , \5446_b1 , \5446_b0 , 
		\5447_b1 , \5447_b0 , \5448_b1 , \5448_b0 , \5449_b1 , \5449_b0 , \5450_b1 , \5450_b0 , \5451_b1 , \5451_b0 , 
		\5452_b1 , \5452_b0 , \5453_b1 , \5453_b0 , \5454_b1 , \5454_b0 , \5455_b1 , \5455_b0 , \5456_b1 , \5456_b0 , 
		\5457_b1 , \5457_b0 , \5458_b1 , \5458_b0 , \5459_b1 , \5459_b0 , \5460_b1 , \5460_b0 , \5461_b1 , \5461_b0 , 
		\5462_b1 , \5462_b0 , \5463_b1 , \5463_b0 , \5464_b1 , \5464_b0 , \5465_b1 , \5465_b0 , \5466_b1 , \5466_b0 , 
		\5467_b1 , \5467_b0 , \5468_b1 , \5468_b0 , \5469_b1 , \5469_b0 , \5470_b1 , \5470_b0 , \5471_b1 , \5471_b0 , 
		\5472_b1 , \5472_b0 , \5473_b1 , \5473_b0 , \5474_b1 , \5474_b0 , \5475_b1 , \5475_b0 , \5476_b1 , \5476_b0 , 
		\5477_b1 , \5477_b0 , \5478_b1 , \5478_b0 , \5479_b1 , \5479_b0 , \5480_b1 , \5480_b0 , \5481_b1 , \5481_b0 , 
		\5482_b1 , \5482_b0 , \5483_b1 , \5483_b0 , \5484_b1 , \5484_b0 , \5485_b1 , \5485_b0 , \5486_b1 , \5486_b0 , 
		\5487_b1 , \5487_b0 , \5488_b1 , \5488_b0 , \5489_b1 , \5489_b0 , \5490_b1 , \5490_b0 , \5491_b1 , \5491_b0 , 
		\5492_b1 , \5492_b0 , \5493_b1 , \5493_b0 , \5494_b1 , \5494_b0 , \5495_b1 , \5495_b0 , \5496_b1 , \5496_b0 , 
		\5497_b1 , \5497_b0 , \5498_b1 , \5498_b0 , \5499_b1 , \5499_b0 , \5500_b1 , \5500_b0 , \5501_b1 , \5501_b0 , 
		\5502_b1 , \5502_b0 , \5503_b1 , \5503_b0 , \5504_b1 , \5504_b0 , \5505_b1 , \5505_b0 , \5506_b1 , \5506_b0 , 
		\5507_b1 , \5507_b0 , \5508_b1 , \5508_b0 , \5509_b1 , \5509_b0 , \5510_b1 , \5510_b0 , \5511_b1 , \5511_b0 , 
		\5512_b1 , \5512_b0 , \5513_b1 , \5513_b0 , \5514_b1 , \5514_b0 , \5515_b1 , \5515_b0 , \5516_b1 , \5516_b0 , 
		\5517_b1 , \5517_b0 , \5518_b1 , \5518_b0 , \5519_b1 , \5519_b0 , \5520_b1 , \5520_b0 , \5521_b1 , \5521_b0 , 
		\5522_b1 , \5522_b0 , \5523_b1 , \5523_b0 , \5524_b1 , \5524_b0 , \5525_b1 , \5525_b0 , \5526_b1 , \5526_b0 , 
		\5527_b1 , \5527_b0 , \5528_b1 , \5528_b0 , \5529_b1 , \5529_b0 , \5530_b1 , \5530_b0 , \5531_b1 , \5531_b0 , 
		\5532_b1 , \5532_b0 , \5533_b1 , \5533_b0 , \5534_b1 , \5534_b0 , \5535_b1 , \5535_b0 , \5536_b1 , \5536_b0 , 
		\5537_b1 , \5537_b0 , \5538_b1 , \5538_b0 , \5539_b1 , \5539_b0 , \5540_b1 , \5540_b0 , \5541_b1 , \5541_b0 , 
		\5542_b1 , \5542_b0 , \5543_b1 , \5543_b0 , \5544_b1 , \5544_b0 , \5545_b1 , \5545_b0 , \5546_b1 , \5546_b0 , 
		\5547_b1 , \5547_b0 , \5548_b1 , \5548_b0 , \5549_b1 , \5549_b0 , \5550_b1 , \5550_b0 , \5551_b1 , \5551_b0 , 
		\5552_b1 , \5552_b0 , \5553_b1 , \5553_b0 , \5554_b1 , \5554_b0 , \5555_b1 , \5555_b0 , \5556_b1 , \5556_b0 , 
		\5557_b1 , \5557_b0 , \5558_b1 , \5558_b0 , \5559_b1 , \5559_b0 , \5560_b1 , \5560_b0 , \5561_b1 , \5561_b0 , 
		\5562_b1 , \5562_b0 , \5563_b1 , \5563_b0 , \5564_b1 , \5564_b0 , \5565_b1 , \5565_b0 , \5566_b1 , \5566_b0 , 
		\5567_b1 , \5567_b0 , \5568_b1 , \5568_b0 , \5569_b1 , \5569_b0 , \5570_b1 , \5570_b0 , \5571_b1 , \5571_b0 , 
		\5572_b1 , \5572_b0 , \5573_b1 , \5573_b0 , \5574_b1 , \5574_b0 , \5575_b1 , \5575_b0 , \5576_b1 , \5576_b0 , 
		\5577_b1 , \5577_b0 , \5578_b1 , \5578_b0 , \5579_b1 , \5579_b0 , \5580_b1 , \5580_b0 , \5581_b1 , \5581_b0 , 
		\5582_b1 , \5582_b0 , \5583_b1 , \5583_b0 , \5584_b1 , \5584_b0 , \5585_b1 , \5585_b0 , \5586_b1 , \5586_b0 , 
		\5587_b1 , \5587_b0 , \5588_b1 , \5588_b0 , \5589_b1 , \5589_b0 , \5590_b1 , \5590_b0 , \5591_b1 , \5591_b0 , 
		\5592_b1 , \5592_b0 , \5593_b1 , \5593_b0 , \5594_b1 , \5594_b0 , \5595_b1 , \5595_b0 , \5596_b1 , \5596_b0 , 
		\5597_b1 , \5597_b0 , \5598_b1 , \5598_b0 , \5599_b1 , \5599_b0 , \5600_b1 , \5600_b0 , \5601_b1 , \5601_b0 , 
		\5602_b1 , \5602_b0 , \5603_b1 , \5603_b0 , \5604_b1 , \5604_b0 , \5605_b1 , \5605_b0 , \5606_b1 , \5606_b0 , 
		\5607_b1 , \5607_b0 , \5608_b1 , \5608_b0 , \5609_b1 , \5609_b0 , \5610_b1 , \5610_b0 , \5611_b1 , \5611_b0 , 
		\5612_b1 , \5612_b0 , \5613_b1 , \5613_b0 , \5614_b1 , \5614_b0 , \5615_b1 , \5615_b0 , \5616_b1 , \5616_b0 , 
		\5617_b1 , \5617_b0 , \5618_b1 , \5618_b0 , \5619_b1 , \5619_b0 , \5620_b1 , \5620_b0 , \5621_b1 , \5621_b0 , 
		\5622_b1 , \5622_b0 , \5623_b1 , \5623_b0 , \5624_b1 , \5624_b0 , \5625_b1 , \5625_b0 , \5626_b1 , \5626_b0 , 
		\5627_b1 , \5627_b0 , \5628_b1 , \5628_b0 , \5629_b1 , \5629_b0 , \5630_b1 , \5630_b0 , \5631_b1 , \5631_b0 , 
		\5632_b1 , \5632_b0 , \5633_b1 , \5633_b0 , \5634_b1 , \5634_b0 , \5635_b1 , \5635_b0 , \5636_b1 , \5636_b0 , 
		\5637_b1 , \5637_b0 , \5638_b1 , \5638_b0 , \5639_b1 , \5639_b0 , \5640_b1 , \5640_b0 , \5641_b1 , \5641_b0 , 
		\5642_b1 , \5642_b0 , \5643_b1 , \5643_b0 , \5644_b1 , \5644_b0 , \5645_b1 , \5645_b0 , \5646_b1 , \5646_b0 , 
		\5647_b1 , \5647_b0 , \5648_b1 , \5648_b0 , \5649_b1 , \5649_b0 , \5650_b1 , \5650_b0 , \5651_b1 , \5651_b0 , 
		\5652_b1 , \5652_b0 , \5653_b1 , \5653_b0 , \5654_b1 , \5654_b0 , \5655_b1 , \5655_b0 , \5656_b1 , \5656_b0 , 
		\5657_b1 , \5657_b0 , \5658_b1 , \5658_b0 , \5659_b1 , \5659_b0 , \5660_b1 , \5660_b0 , \5661_b1 , \5661_b0 , 
		\5662_b1 , \5662_b0 , \5663_b1 , \5663_b0 , \5664_b1 , \5664_b0 , \5665_b1 , \5665_b0 , \5666_b1 , \5666_b0 , 
		\5667_b1 , \5667_b0 , \5668_b1 , \5668_b0 , \5669_b1 , \5669_b0 , \5670_b1 , \5670_b0 , \5671_b1 , \5671_b0 , 
		\5672_b1 , \5672_b0 , \5673_b1 , \5673_b0 , \5674_b1 , \5674_b0 , \5675_b1 , \5675_b0 , \5676_b1 , \5676_b0 , 
		\5677_b1 , \5677_b0 , \5678_b1 , \5678_b0 , \5679_b1 , \5679_b0 , \5680_b1 , \5680_b0 , \5681_b1 , \5681_b0 , 
		\5682_b1 , \5682_b0 , \5683_b1 , \5683_b0 , \5684_b1 , \5684_b0 , \5685_b1 , \5685_b0 , \5686_b1 , \5686_b0 , 
		\5687_b1 , \5687_b0 , \5688_b1 , \5688_b0 , \5689_b1 , \5689_b0 , \5690_b1 , \5690_b0 , \5691_b1 , \5691_b0 , 
		\5692_b1 , \5692_b0 , \5693_b1 , \5693_b0 , \5694_b1 , \5694_b0 , \5695_b1 , \5695_b0 , \5696_b1 , \5696_b0 , 
		\5697_b1 , \5697_b0 , \5698_b1 , \5698_b0 , \5699_b1 , \5699_b0 , \5700_b1 , \5700_b0 , \5701_b1 , \5701_b0 , 
		\5702_b1 , \5702_b0 , \5703_b1 , \5703_b0 , \5704_b1 , \5704_b0 , \5705_b1 , \5705_b0 , \5706_b1 , \5706_b0 , 
		\5707_b1 , \5707_b0 , \5708_b1 , \5708_b0 , \5709_b1 , \5709_b0 , \5710_b1 , \5710_b0 , \5711_b1 , \5711_b0 , 
		\5712_b1 , \5712_b0 , \5713_b1 , \5713_b0 , \5714_b1 , \5714_b0 , \5715_b1 , \5715_b0 , \5716_b1 , \5716_b0 , 
		\5717_b1 , \5717_b0 , \5718_b1 , \5718_b0 , \5719_b1 , \5719_b0 , \5720_b1 , \5720_b0 , \5721_b1 , \5721_b0 , 
		\5722_b1 , \5722_b0 , \5723_b1 , \5723_b0 , \5724_b1 , \5724_b0 , \5725_b1 , \5725_b0 , \5726_b1 , \5726_b0 , 
		\5727_b1 , \5727_b0 , \5728_b1 , \5728_b0 , \5729_b1 , \5729_b0 , \5730_b1 , \5730_b0 , \5731_b1 , \5731_b0 , 
		\5732_b1 , \5732_b0 , \5733_b1 , \5733_b0 , \5734_b1 , \5734_b0 , \5735_b1 , \5735_b0 , \5736_b1 , \5736_b0 , 
		\5737_b1 , \5737_b0 , \5738_b1 , \5738_b0 , \5739_b1 , \5739_b0 , \5740_b1 , \5740_b0 , \5741_b1 , \5741_b0 , 
		\5742_b1 , \5742_b0 , \5743_b1 , \5743_b0 , \5744_b1 , \5744_b0 , \5745_b1 , \5745_b0 , \5746_b1 , \5746_b0 , 
		\5747_b1 , \5747_b0 , \5748_b1 , \5748_b0 , \5749_b1 , \5749_b0 , \5750_b1 , \5750_b0 , \5751_b1 , \5751_b0 , 
		\5752_b1 , \5752_b0 , \5753_b1 , \5753_b0 , \5754_b1 , \5754_b0 , \5755_b1 , \5755_b0 , \5756_b1 , \5756_b0 , 
		\5757_b1 , \5757_b0 , \5758_b1 , \5758_b0 , \5759_b1 , \5759_b0 , \5760_b1 , \5760_b0 , \5761_b1 , \5761_b0 , 
		\5762_b1 , \5762_b0 , \5763_b1 , \5763_b0 , \5764_b1 , \5764_b0 , \5765_b1 , \5765_b0 , \5766_b1 , \5766_b0 , 
		\5767_b1 , \5767_b0 , \5768_b1 , \5768_b0 , \5769_b1 , \5769_b0 , \5770_b1 , \5770_b0 , \5771_b1 , \5771_b0 , 
		\5772_b1 , \5772_b0 , \5773_b1 , \5773_b0 , \5774_b1 , \5774_b0 , \5775_b1 , \5775_b0 , \5776_b1 , \5776_b0 , 
		\5777_b1 , \5777_b0 , \5778_b1 , \5778_b0 , \5779_b1 , \5779_b0 , \5780_b1 , \5780_b0 , \5781_b1 , \5781_b0 , 
		\5782_b1 , \5782_b0 , \5783_b1 , \5783_b0 , \5784_b1 , \5784_b0 , \5785_b1 , \5785_b0 , \5786_b1 , \5786_b0 , 
		\5787_b1 , \5787_b0 , \5788_b1 , \5788_b0 , \5789_b1 , \5789_b0 , \5790_b1 , \5790_b0 , \5791_b1 , \5791_b0 , 
		\5792_b1 , \5792_b0 , \5793_b1 , \5793_b0 , \5794_b1 , \5794_b0 , \5795_b1 , \5795_b0 , \5796_b1 , \5796_b0 , 
		\5797_b1 , \5797_b0 , \5798_b1 , \5798_b0 , \5799_b1 , \5799_b0 , \5800_b1 , \5800_b0 , \5801_b1 , \5801_b0 , 
		\5802_b1 , \5802_b0 , \5803_b1 , \5803_b0 , \5804_b1 , \5804_b0 , \5805_b1 , \5805_b0 , \5806_b1 , \5806_b0 , 
		\5807_b1 , \5807_b0 , \5808_b1 , \5808_b0 , \5809_b1 , \5809_b0 , \5810_b1 , \5810_b0 , \5811_b1 , \5811_b0 , 
		\5812_b1 , \5812_b0 , \5813_b1 , \5813_b0 , \5814_b1 , \5814_b0 , \5815_b1 , \5815_b0 , \5816_b1 , \5816_b0 , 
		\5817_b1 , \5817_b0 , \5818_b1 , \5818_b0 , \5819_b1 , \5819_b0 , \5820_b1 , \5820_b0 , \5821_b1 , \5821_b0 , 
		\5822_b1 , \5822_b0 , \5823_b1 , \5823_b0 , \5824_b1 , \5824_b0 , \5825_b1 , \5825_b0 , \5826_b1 , \5826_b0 , 
		\5827_b1 , \5827_b0 , \5828_b1 , \5828_b0 , \5829_b1 , \5829_b0 , \5830_b1 , \5830_b0 , \5831_b1 , \5831_b0 , 
		\5832_b1 , \5832_b0 , \5833_b1 , \5833_b0 , \5834_b1 , \5834_b0 , \5835_b1 , \5835_b0 , \5836_b1 , \5836_b0 , 
		\5837_b1 , \5837_b0 , \5838_b1 , \5838_b0 , \5839_b1 , \5839_b0 , \5840_b1 , \5840_b0 , \5841_b1 , \5841_b0 , 
		\5842_b1 , \5842_b0 , \5843_b1 , \5843_b0 , \5844_b1 , \5844_b0 , \5845_b1 , \5845_b0 , \5846_b1 , \5846_b0 , 
		\5847_b1 , \5847_b0 , \5848_b1 , \5848_b0 , \5849_b1 , \5849_b0 , \5850_b1 , \5850_b0 , \5851_b1 , \5851_b0 , 
		\5852_b1 , \5852_b0 , \5853_b1 , \5853_b0 , \5854_b1 , \5854_b0 , \5855_b1 , \5855_b0 , \5856_b1 , \5856_b0 , 
		\5857_b1 , \5857_b0 , \5858_b1 , \5858_b0 , \5859_b1 , \5859_b0 , \5860_b1 , \5860_b0 , \5861_b1 , \5861_b0 , 
		\5862_b1 , \5862_b0 , \5863_b1 , \5863_b0 , \5864_b1 , \5864_b0 , \5865_b1 , \5865_b0 , \5866_b1 , \5866_b0 , 
		\5867_b1 , \5867_b0 , \5868_b1 , \5868_b0 , \5869_b1 , \5869_b0 , \5870_b1 , \5870_b0 , \5871_b1 , \5871_b0 , 
		\5872_b1 , \5872_b0 , \5873_b1 , \5873_b0 , \5874_b1 , \5874_b0 , \5875_b1 , \5875_b0 , \5876_b1 , \5876_b0 , 
		\5877_b1 , \5877_b0 , \5878_b1 , \5878_b0 , \5879_b1 , \5879_b0 , \5880_b1 , \5880_b0 , \5881_b1 , \5881_b0 , 
		\5882_b1 , \5882_b0 , \5883_b1 , \5883_b0 , \5884_b1 , \5884_b0 , \5885_b1 , \5885_b0 , \5886_b1 , \5886_b0 , 
		\5887_b1 , \5887_b0 , \5888_b1 , \5888_b0 , \5889_b1 , \5889_b0 , \5890_b1 , \5890_b0 , \5891_b1 , \5891_b0 , 
		\5892_b1 , \5892_b0 , \5893_b1 , \5893_b0 , \5894_b1 , \5894_b0 , \5895_b1 , \5895_b0 , \5896_b1 , \5896_b0 , 
		\5897_b1 , \5897_b0 , \5898_b1 , \5898_b0 , \5899_b1 , \5899_b0 , \5900_b1 , \5900_b0 , \5901_b1 , \5901_b0 , 
		\5902_b1 , \5902_b0 , \5903_b1 , \5903_b0 , \5904_b1 , \5904_b0 , \5905_b1 , \5905_b0 , \5906_b1 , \5906_b0 , 
		\5907_b1 , \5907_b0 , \5908_b1 , \5908_b0 , \5909_b1 , \5909_b0 , \5910_b1 , \5910_b0 , \5911_b1 , \5911_b0 , 
		\5912_b1 , \5912_b0 , \5913_b1 , \5913_b0 , \5914_b1 , \5914_b0 , \5915_b1 , \5915_b0 , \5916_b1 , \5916_b0 , 
		\5917_b1 , \5917_b0 , \5918_b1 , \5918_b0 , \5919_b1 , \5919_b0 , \5920_b1 , \5920_b0 , \5921_b1 , \5921_b0 , 
		\5922_b1 , \5922_b0 , \5923_b1 , \5923_b0 , \5924_b1 , \5924_b0 , \5925_b1 , \5925_b0 , \5926_b1 , \5926_b0 , 
		\5927_b1 , \5927_b0 , \5928_b1 , \5928_b0 , \5929_b1 , \5929_b0 , \5930_b1 , \5930_b0 , \5931_b1 , \5931_b0 , 
		\5932_b1 , \5932_b0 , \5933_b1 , \5933_b0 , \5934_b1 , \5934_b0 , \5935_b1 , \5935_b0 , \5936_b1 , \5936_b0 , 
		\5937_b1 , \5937_b0 , \5938_b1 , \5938_b0 , \5939_b1 , \5939_b0 , \5940_b1 , \5940_b0 , \5941_b1 , \5941_b0 , 
		\5942_b1 , \5942_b0 , \5943_b1 , \5943_b0 , \5944_b1 , \5944_b0 , \5945_b1 , \5945_b0 , \5946_b1 , \5946_b0 , 
		\5947_b1 , \5947_b0 , \5948_b1 , \5948_b0 , \5949_b1 , \5949_b0 , \5950_b1 , \5950_b0 , \5951_b1 , \5951_b0 , 
		\5952_b1 , \5952_b0 , \5953_b1 , \5953_b0 , \5954_b1 , \5954_b0 , \5955_b1 , \5955_b0 , \5956_b1 , \5956_b0 , 
		\5957_b1 , \5957_b0 , \5958_b1 , \5958_b0 , \5959_b1 , \5959_b0 , \5960_b1 , \5960_b0 , \5961_b1 , \5961_b0 , 
		\5962_b1 , \5962_b0 , \5963_b1 , \5963_b0 , \5964_b1 , \5964_b0 , \5965_b1 , \5965_b0 , \5966_b1 , \5966_b0 , 
		\5967_b1 , \5967_b0 , \5968_b1 , \5968_b0 , \5969_b1 , \5969_b0 , \5970_b1 , \5970_b0 , \5971_b1 , \5971_b0 , 
		\5972_b1 , \5972_b0 , \5973_b1 , \5973_b0 , \5974_b1 , \5974_b0 , \5975_b1 , \5975_b0 , \5976_b1 , \5976_b0 , 
		\5977_b1 , \5977_b0 , \5978_b1 , \5978_b0 , \5979_b1 , \5979_b0 , \5980_b1 , \5980_b0 , \5981_b1 , \5981_b0 , 
		\5982_b1 , \5982_b0 , \5983_b1 , \5983_b0 , \5984_b1 , \5984_b0 , \5985_b1 , \5985_b0 , \5986_b1 , \5986_b0 , 
		\5987_b1 , \5987_b0 , \5988_b1 , \5988_b0 , \5989_b1 , \5989_b0 , \5990_b1 , \5990_b0 , \5991_b1 , \5991_b0 , 
		\5992_b1 , \5992_b0 , \5993_b1 , \5993_b0 , \5994_b1 , \5994_b0 , \5995_b1 , \5995_b0 , \5996_b1 , \5996_b0 , 
		\5997_b1 , \5997_b0 , \5998_b1 , \5998_b0 , \5999_b1 , \5999_b0 , \6000_b1 , \6000_b0 , \6001_b1 , \6001_b0 , 
		\6002_b1 , \6002_b0 , \6003_b1 , \6003_b0 , \6004_b1 , \6004_b0 , \6005_b1 , \6005_b0 , \6006_b1 , \6006_b0 , 
		\6007_b1 , \6007_b0 , \6008_b1 , \6008_b0 , \6009_b1 , \6009_b0 , \6010_b1 , \6010_b0 , \6011_b1 , \6011_b0 , 
		\6012_b1 , \6012_b0 , \6013_b1 , \6013_b0 , \6014_b1 , \6014_b0 , \6015_b1 , \6015_b0 , \6016_b1 , \6016_b0 , 
		\6017_b1 , \6017_b0 , \6018_b1 , \6018_b0 , \6019_b1 , \6019_b0 , \6020_b1 , \6020_b0 , \6021_b1 , \6021_b0 , 
		\6022_b1 , \6022_b0 , \6023_b1 , \6023_b0 , \6024_b1 , \6024_b0 , \6025_b1 , \6025_b0 , \6026_b1 , \6026_b0 , 
		\6027_b1 , \6027_b0 , \6028_b1 , \6028_b0 , \6029_b1 , \6029_b0 , \6030_b1 , \6030_b0 , \6031_b1 , \6031_b0 , 
		\6032_b1 , \6032_b0 , \6033_b1 , \6033_b0 , \6034_b1 , \6034_b0 , \6035_b1 , \6035_b0 , \6036_b1 , \6036_b0 , 
		\6037_b1 , \6037_b0 , \6038_b1 , \6038_b0 , \6039_b1 , \6039_b0 , \6040_b1 , \6040_b0 , \6041_b1 , \6041_b0 , 
		\6042_b1 , \6042_b0 , \6043_b1 , \6043_b0 , \6044_b1 , \6044_b0 , \6045_b1 , \6045_b0 , \6046_b1 , \6046_b0 , 
		\6047_b1 , \6047_b0 , \6048_b1 , \6048_b0 , \6049_b1 , \6049_b0 , \6050_b1 , \6050_b0 , \6051_b1 , \6051_b0 , 
		\6052_b1 , \6052_b0 , \6053_b1 , \6053_b0 , \6054_b1 , \6054_b0 , \6055_b1 , \6055_b0 , \6056_b1 , \6056_b0 , 
		\6057_b1 , \6057_b0 , \6058_b1 , \6058_b0 , \6059_b1 , \6059_b0 , \6060_b1 , \6060_b0 , \6061_b1 , \6061_b0 , 
		\6062_b1 , \6062_b0 , \6063_b1 , \6063_b0 , \6064_b1 , \6064_b0 , \6065_b1 , \6065_b0 , \6066_b1 , \6066_b0 , 
		\6067_b1 , \6067_b0 , \6068_b1 , \6068_b0 , \6069_b1 , \6069_b0 , \6070_b1 , \6070_b0 , \6071_b1 , \6071_b0 , 
		\6072_b1 , \6072_b0 , \6073_b1 , \6073_b0 , \6074_b1 , \6074_b0 , \6075_b1 , \6075_b0 , \6076_b1 , \6076_b0 , 
		\6077_b1 , \6077_b0 , \6078_b1 , \6078_b0 , \6079_b1 , \6079_b0 , \6080_b1 , \6080_b0 , \6081_b1 , \6081_b0 , 
		\6082_b1 , \6082_b0 , \6083_b1 , \6083_b0 , \6084_b1 , \6084_b0 , \6085_b1 , \6085_b0 , \6086_b1 , \6086_b0 , 
		\6087_b1 , \6087_b0 , \6088_b1 , \6088_b0 , \6089_b1 , \6089_b0 , \6090_b1 , \6090_b0 , \6091_b1 , \6091_b0 , 
		\6092_b1 , \6092_b0 , \6093_b1 , \6093_b0 , \6094_b1 , \6094_b0 , \6095_b1 , \6095_b0 , \6096_b1 , \6096_b0 , 
		\6097_b1 , \6097_b0 , \6098_b1 , \6098_b0 , \6099_b1 , \6099_b0 , \6100_b1 , \6100_b0 , \6101_b1 , \6101_b0 , 
		\6102_b1 , \6102_b0 , \6103_b1 , \6103_b0 , \6104_b1 , \6104_b0 , \6105_b1 , \6105_b0 , \6106_b1 , \6106_b0 , 
		\6107_b1 , \6107_b0 , \6108_b1 , \6108_b0 , \6109_b1 , \6109_b0 , \6110_b1 , \6110_b0 , \6111_b1 , \6111_b0 , 
		\6112_b1 , \6112_b0 , \6113_b1 , \6113_b0 , \6114_b1 , \6114_b0 , \6115_b1 , \6115_b0 , \6116_b1 , \6116_b0 , 
		\6117_b1 , \6117_b0 , \6118_b1 , \6118_b0 , \6119_b1 , \6119_b0 , \6120_b1 , \6120_b0 , \6121_b1 , \6121_b0 , 
		\6122_b1 , \6122_b0 , \6123_b1 , \6123_b0 , \6124_b1 , \6124_b0 , \6125_b1 , \6125_b0 , \6126_b1 , \6126_b0 , 
		\6127_b1 , \6127_b0 , \6128_b1 , \6128_b0 , \6129_b1 , \6129_b0 , \6130_b1 , \6130_b0 , \6131_b1 , \6131_b0 , 
		\6132_b1 , \6132_b0 , \6133_b1 , \6133_b0 , \6134_b1 , \6134_b0 , \6135_b1 , \6135_b0 , \6136_b1 , \6136_b0 , 
		\6137_b1 , \6137_b0 , \6138_b1 , \6138_b0 , \6139_b1 , \6139_b0 , \6140_b1 , \6140_b0 , \6141_b1 , \6141_b0 , 
		\6142_b1 , \6142_b0 , \6143_b1 , \6143_b0 , \6144_b1 , \6144_b0 , \6145_b1 , \6145_b0 , \6146_b1 , \6146_b0 , 
		\6147_b1 , \6147_b0 , \6148_b1 , \6148_b0 , \6149_b1 , \6149_b0 , \6150_b1 , \6150_b0 , \6151_b1 , \6151_b0 , 
		\6152_b1 , \6152_b0 , \6153_b1 , \6153_b0 , \6154_b1 , \6154_b0 , \6155_b1 , \6155_b0 , \6156_b1 , \6156_b0 , 
		\6157_b1 , \6157_b0 , \6158_b1 , \6158_b0 , \6159_b1 , \6159_b0 , \6160_b1 , \6160_b0 , \6161_b1 , \6161_b0 , 
		\6162_b1 , \6162_b0 , \6163_b1 , \6163_b0 , \6164_b1 , \6164_b0 , \6165_b1 , \6165_b0 , \6166_b1 , \6166_b0 , 
		\6167_b1 , \6167_b0 , \6168_b1 , \6168_b0 , \6169_b1 , \6169_b0 , \6170_b1 , \6170_b0 , \6171_b1 , \6171_b0 , 
		\6172_b1 , \6172_b0 , \6173_b1 , \6173_b0 , \6174_b1 , \6174_b0 , \6175_b1 , \6175_b0 , \6176_b1 , \6176_b0 , 
		\6177_b1 , \6177_b0 , \6178_b1 , \6178_b0 , \6179_b1 , \6179_b0 , \6180_b1 , \6180_b0 , \6181_b1 , \6181_b0 , 
		\6182_b1 , \6182_b0 , \6183_b1 , \6183_b0 , \6184_b1 , \6184_b0 , \6185_b1 , \6185_b0 , \6186_b1 , \6186_b0 , 
		\6187_b1 , \6187_b0 , \6188_b1 , \6188_b0 , \6189_b1 , \6189_b0 , \6190_b1 , \6190_b0 , \6191_b1 , \6191_b0 , 
		\6192_b1 , \6192_b0 , \6193_b1 , \6193_b0 , \6194_b1 , \6194_b0 , \6195_b1 , \6195_b0 , \6196_b1 , \6196_b0 , 
		\6197_b1 , \6197_b0 , \6198_b1 , \6198_b0 , \6199_b1 , \6199_b0 , \6200_b1 , \6200_b0 , \6201_b1 , \6201_b0 , 
		\6202_b1 , \6202_b0 , \6203_b1 , \6203_b0 , \6204_b1 , \6204_b0 , \6205_b1 , \6205_b0 , \6206_b1 , \6206_b0 , 
		\6207_b1 , \6207_b0 , \6208_b1 , \6208_b0 , \6209_b1 , \6209_b0 , \6210_b1 , \6210_b0 , \6211_b1 , \6211_b0 , 
		\6212_b1 , \6212_b0 , \6213_b1 , \6213_b0 , \6214_b1 , \6214_b0 , \6215_b1 , \6215_b0 , \6216_b1 , \6216_b0 , 
		\6217_b1 , \6217_b0 , \6218_b1 , \6218_b0 , \6219_b1 , \6219_b0 , \6220_b1 , \6220_b0 , \6221_b1 , \6221_b0 , 
		\6222_b1 , \6222_b0 , \6223_b1 , \6223_b0 , \6224_b1 , \6224_b0 , \6225_b1 , \6225_b0 , \6226_b1 , \6226_b0 , 
		\6227_b1 , \6227_b0 , \6228_b1 , \6228_b0 , \6229_b1 , \6229_b0 , \6230_b1 , \6230_b0 , \6231_b1 , \6231_b0 , 
		\6232_b1 , \6232_b0 , \6233_b1 , \6233_b0 , \6234_b1 , \6234_b0 , \6235_b1 , \6235_b0 , \6236_b1 , \6236_b0 , 
		\6237_b1 , \6237_b0 , \6238_b1 , \6238_b0 , \6239_b1 , \6239_b0 , \6240_b1 , \6240_b0 , \6241_b1 , \6241_b0 , 
		\6242_b1 , \6242_b0 , \6243_b1 , \6243_b0 , \6244_b1 , \6244_b0 , \6245_b1 , \6245_b0 , \6246_b1 , \6246_b0 , 
		\6247_b1 , \6247_b0 , \6248_b1 , \6248_b0 , \6249_b1 , \6249_b0 , \6250_b1 , \6250_b0 , \6251_b1 , \6251_b0 , 
		\6252_b1 , \6252_b0 , \6253_b1 , \6253_b0 , \6254_b1 , \6254_b0 , \6255_b1 , \6255_b0 , \6256_b1 , \6256_b0 , 
		\6257_b1 , \6257_b0 , \6258_b1 , \6258_b0 , \6259_b1 , \6259_b0 , \6260_b1 , \6260_b0 , \6261_b1 , \6261_b0 , 
		\6262_b1 , \6262_b0 , \6263_b1 , \6263_b0 , \6264_b1 , \6264_b0 , \6265_b1 , \6265_b0 , \6266_b1 , \6266_b0 , 
		\6267_b1 , \6267_b0 , \6268_b1 , \6268_b0 , \6269_b1 , \6269_b0 , \6270_b1 , \6270_b0 , \6271_b1 , \6271_b0 , 
		\6272_b1 , \6272_b0 , \6273_b1 , \6273_b0 , \6274_b1 , \6274_b0 , \6275_b1 , \6275_b0 , \6276_b1 , \6276_b0 , 
		\6277_b1 , \6277_b0 , \6278_b1 , \6278_b0 , \6279_b1 , \6279_b0 , \6280_b1 , \6280_b0 , \6281_b1 , \6281_b0 , 
		\6282_b1 , \6282_b0 , \6283_b1 , \6283_b0 , \6284_b1 , \6284_b0 , \6285_b1 , \6285_b0 , \6286_b1 , \6286_b0 , 
		\6287_b1 , \6287_b0 , \6288_b1 , \6288_b0 , \6289_b1 , \6289_b0 , \6290_b1 , \6290_b0 , \6291_b1 , \6291_b0 , 
		\6292_b1 , \6292_b0 , \6293_b1 , \6293_b0 , \6294_b1 , \6294_b0 , \6295_b1 , \6295_b0 , \6296_b1 , \6296_b0 , 
		\6297_b1 , \6297_b0 , \6298_b1 , \6298_b0 , \6299_b1 , \6299_b0 , \6300_b1 , \6300_b0 , \6301_b1 , \6301_b0 , 
		\6302_b1 , \6302_b0 , \6303_b1 , \6303_b0 , \6304_b1 , \6304_b0 , \6305_b1 , \6305_b0 , \6306_b1 , \6306_b0 , 
		\6307_b1 , \6307_b0 , \6308_b1 , \6308_b0 , \6309_b1 , \6309_b0 , \6310_b1 , \6310_b0 , \6311_b1 , \6311_b0 , 
		\6312_b1 , \6312_b0 , \6313_b1 , \6313_b0 , \6314_b1 , \6314_b0 , \6315_b1 , \6315_b0 , \6316_b1 , \6316_b0 , 
		\6317_b1 , \6317_b0 , \6318_b1 , \6318_b0 , \6319_b1 , \6319_b0 , \6320_b1 , \6320_b0 , \6321_b1 , \6321_b0 , 
		\6322_b1 , \6322_b0 , \6323_b1 , \6323_b0 , \6324_b1 , \6324_b0 , \6325_b1 , \6325_b0 , \6326_b1 , \6326_b0 , 
		\6327_b1 , \6327_b0 , \6328_b1 , \6328_b0 , \6329_b1 , \6329_b0 , \6330_b1 , \6330_b0 , \6331_b1 , \6331_b0 , 
		\6332_b1 , \6332_b0 , \6333_b1 , \6333_b0 , \6334_b1 , \6334_b0 , \6335_b1 , \6335_b0 , \6336_b1 , \6336_b0 , 
		\6337_b1 , \6337_b0 , \6338_b1 , \6338_b0 , \6339_b1 , \6339_b0 , \6340_b1 , \6340_b0 , \6341_b1 , \6341_b0 , 
		\6342_b1 , \6342_b0 , \6343_b1 , \6343_b0 , \6344_b1 , \6344_b0 , \6345_b1 , \6345_b0 , \6346_b1 , \6346_b0 , 
		\6347_b1 , \6347_b0 , \6348_b1 , \6348_b0 , \6349_b1 , \6349_b0 , \6350_b1 , \6350_b0 , \6351_b1 , \6351_b0 , 
		\6352_b1 , \6352_b0 , \6353_b1 , \6353_b0 , \6354_b1 , \6354_b0 , \6355_b1 , \6355_b0 , \6356_b1 , \6356_b0 , 
		\6357_b1 , \6357_b0 , \6358_b1 , \6358_b0 , \6359_b1 , \6359_b0 , \6360_b1 , \6360_b0 , \6361_b1 , \6361_b0 , 
		\6362_b1 , \6362_b0 , \6363_b1 , \6363_b0 , \6364_b1 , \6364_b0 , \6365_b1 , \6365_b0 , \6366_b1 , \6366_b0 , 
		\6367_b1 , \6367_b0 , \6368_b1 , \6368_b0 , \6369_b1 , \6369_b0 , \6370_b1 , \6370_b0 , \6371_b1 , \6371_b0 , 
		\6372_b1 , \6372_b0 , \6373_b1 , \6373_b0 , \6374_b1 , \6374_b0 , \6375_b1 , \6375_b0 , \6376_b1 , \6376_b0 , 
		\6377_b1 , \6377_b0 , \6378_b1 , \6378_b0 , \6379_b1 , \6379_b0 , \6380_b1 , \6380_b0 , \6381_b1 , \6381_b0 , 
		\6382_b1 , \6382_b0 , \6383_b1 , \6383_b0 , \6384_b1 , \6384_b0 , \6385_b1 , \6385_b0 , \6386_b1 , \6386_b0 , 
		\6387_b1 , \6387_b0 , \6388_b1 , \6388_b0 , \6389_b1 , \6389_b0 , \6390_b1 , \6390_b0 , \6391_b1 , \6391_b0 , 
		\6392_b1 , \6392_b0 , \6393_b1 , \6393_b0 , \6394_b1 , \6394_b0 , \6395_b1 , \6395_b0 , \6396_b1 , \6396_b0 , 
		\6397_b1 , \6397_b0 , \6398_b1 , \6398_b0 , \6399_b1 , \6399_b0 , \6400_b1 , \6400_b0 , \6401_b1 , \6401_b0 , 
		\6402_b1 , \6402_b0 , \6403_b1 , \6403_b0 , \6404_b1 , \6404_b0 , \6405_b1 , \6405_b0 , \6406_b1 , \6406_b0 , 
		\6407_b1 , \6407_b0 , \6408_b1 , \6408_b0 , \6409_b1 , \6409_b0 , \6410_b1 , \6410_b0 , \6411_b1 , \6411_b0 , 
		\6412_b1 , \6412_b0 , \6413_b1 , \6413_b0 , \6414_b1 , \6414_b0 , \6415_b1 , \6415_b0 , \6416_b1 , \6416_b0 , 
		\6417_b1 , \6417_b0 , \6418_b1 , \6418_b0 , \6419_b1 , \6419_b0 , \6420_b1 , \6420_b0 , \6421_b1 , \6421_b0 , 
		\6422_b1 , \6422_b0 , \6423_b1 , \6423_b0 , \6424_b1 , \6424_b0 , \6425_b1 , \6425_b0 , \6426_b1 , \6426_b0 , 
		\6427_b1 , \6427_b0 , \6428_b1 , \6428_b0 , \6429_b1 , \6429_b0 , \6430_b1 , \6430_b0 , \6431_b1 , \6431_b0 , 
		\6432_b1 , \6432_b0 , \6433_b1 , \6433_b0 , \6434_b1 , \6434_b0 , \6435_b1 , \6435_b0 , \6436_b1 , \6436_b0 , 
		\6437_b1 , \6437_b0 , \6438_b1 , \6438_b0 , \6439_b1 , \6439_b0 , \6440_b1 , \6440_b0 , \6441_b1 , \6441_b0 , 
		\6442_b1 , \6442_b0 , \6443_b1 , \6443_b0 , \6444_b1 , \6444_b0 , \6445_b1 , \6445_b0 , \6446_b1 , \6446_b0 , 
		\6447_b1 , \6447_b0 , \6448_b1 , \6448_b0 , \6449_b1 , \6449_b0 , \6450_b1 , \6450_b0 , \6451_b1 , \6451_b0 , 
		\6452_b1 , \6452_b0 , \6453_b1 , \6453_b0 , \6454_b1 , \6454_b0 , \6455_b1 , \6455_b0 , \6456_b1 , \6456_b0 , 
		\6457_b1 , \6457_b0 , \6458_b1 , \6458_b0 , \6459_b1 , \6459_b0 , \6460_b1 , \6460_b0 , \6461_b1 , \6461_b0 , 
		\6462_b1 , \6462_b0 , \6463_b1 , \6463_b0 , \6464_b1 , \6464_b0 , \6465_b1 , \6465_b0 , \6466_b1 , \6466_b0 , 
		\6467_b1 , \6467_b0 , \6468_b1 , \6468_b0 , \6469_b1 , \6469_b0 , \6470_b1 , \6470_b0 , \6471_b1 , \6471_b0 , 
		\6472_b1 , \6472_b0 , \6473_b1 , \6473_b0 , \6474_b1 , \6474_b0 , \6475_b1 , \6475_b0 , \6476_b1 , \6476_b0 , 
		\6477_b1 , \6477_b0 , \6478_b1 , \6478_b0 , \6479_b1 , \6479_b0 , \6480_b1 , \6480_b0 , \6481_b1 , \6481_b0 , 
		\6482_b1 , \6482_b0 , \6483_b1 , \6483_b0 , \6484_b1 , \6484_b0 , \6485_b1 , \6485_b0 , \6486_b1 , \6486_b0 , 
		\6487_b1 , \6487_b0 , \6488_b1 , \6488_b0 , \6489_b1 , \6489_b0 , \6490_b1 , \6490_b0 , \6491_b1 , \6491_b0 , 
		\6492_b1 , \6492_b0 , \6493_b1 , \6493_b0 , \6494_b1 , \6494_b0 , \6495_b1 , \6495_b0 , \6496_b1 , \6496_b0 , 
		\6497_b1 , \6497_b0 , \6498_b1 , \6498_b0 , \6499_b1 , \6499_b0 , \6500_b1 , \6500_b0 , \6501_b1 , \6501_b0 , 
		\6502_b1 , \6502_b0 , \6503_b1 , \6503_b0 , \6504_b1 , \6504_b0 , \6505_b1 , \6505_b0 , \6506_b1 , \6506_b0 , 
		\6507_b1 , \6507_b0 , \6508_b1 , \6508_b0 , \6509_b1 , \6509_b0 , \6510_b1 , \6510_b0 , \6511_b1 , \6511_b0 , 
		\6512_b1 , \6512_b0 , \6513_b1 , \6513_b0 , \6514_b1 , \6514_b0 , \6515_b1 , \6515_b0 , \6516_b1 , \6516_b0 , 
		\6517_b1 , \6517_b0 , \6518_b1 , \6518_b0 , \6519_b1 , \6519_b0 , \6520_b1 , \6520_b0 , \6521_b1 , \6521_b0 , 
		\6522_b1 , \6522_b0 , \6523_b1 , \6523_b0 , \6524_b1 , \6524_b0 , \6525_b1 , \6525_b0 , \6526_b1 , \6526_b0 , 
		\6527_b1 , \6527_b0 , \6528_b1 , \6528_b0 , \6529_b1 , \6529_b0 , \6530_b1 , \6530_b0 , \6531_b1 , \6531_b0 , 
		\6532_b1 , \6532_b0 , \6533_b1 , \6533_b0 , \6534_b1 , \6534_b0 , \6535_b1 , \6535_b0 , \6536_b1 , \6536_b0 , 
		\6537_b1 , \6537_b0 , \6538_b1 , \6538_b0 , \6539_b1 , \6539_b0 , \6540_b1 , \6540_b0 , \6541_b1 , \6541_b0 , 
		\6542_b1 , \6542_b0 , \6543_b1 , \6543_b0 , \6544_b1 , \6544_b0 , \6545_b1 , \6545_b0 , \6546_b1 , \6546_b0 , 
		\6547_b1 , \6547_b0 , \6548_b1 , \6548_b0 , \6549_b1 , \6549_b0 , \6550_b1 , \6550_b0 , \6551_b1 , \6551_b0 , 
		\6552_b1 , \6552_b0 , \6553_b1 , \6553_b0 , \6554_b1 , \6554_b0 , \6555_b1 , \6555_b0 , \6556_b1 , \6556_b0 , 
		\6557_b1 , \6557_b0 , \6558_b1 , \6558_b0 , \6559_b1 , \6559_b0 , \6560_b1 , \6560_b0 , \6561_b1 , \6561_b0 , 
		\6562_b1 , \6562_b0 , \6563_b1 , \6563_b0 , \6564_b1 , \6564_b0 , \6565_b1 , \6565_b0 , \6566_b1 , \6566_b0 , 
		\6567_b1 , \6567_b0 , \6568_b1 , \6568_b0 , \6569_b1 , \6569_b0 , \6570_b1 , \6570_b0 , \6571_b1 , \6571_b0 , 
		\6572_b1 , \6572_b0 , \6573_b1 , \6573_b0 , \6574_b1 , \6574_b0 , \6575_b1 , \6575_b0 , \6576_b1 , \6576_b0 , 
		\6577_b1 , \6577_b0 , \6578_b1 , \6578_b0 , \6579_b1 , \6579_b0 , \6580_b1 , \6580_b0 , \6581_b1 , \6581_b0 , 
		\6582_b1 , \6582_b0 , \6583_b1 , \6583_b0 , \6584_b1 , \6584_b0 , \6585_b1 , \6585_b0 , \6586_b1 , \6586_b0 , 
		\6587_b1 , \6587_b0 , \6588_b1 , \6588_b0 , \6589_b1 , \6589_b0 , \6590_b1 , \6590_b0 , \6591_b1 , \6591_b0 , 
		\6592_b1 , \6592_b0 , \6593_b1 , \6593_b0 , \6594_b1 , \6594_b0 , \6595_b1 , \6595_b0 , \6596_b1 , \6596_b0 , 
		\6597_b1 , \6597_b0 , \6598_b1 , \6598_b0 , \6599_b1 , \6599_b0 , \6600_b1 , \6600_b0 , \6601_b1 , \6601_b0 , 
		\6602_b1 , \6602_b0 , \6603_b1 , \6603_b0 , \6604_b1 , \6604_b0 , \6605_b1 , \6605_b0 , \6606_b1 , \6606_b0 , 
		\6607_b1 , \6607_b0 , \6608_b1 , \6608_b0 , \6609_b1 , \6609_b0 , \6610_b1 , \6610_b0 , \6611_b1 , \6611_b0 , 
		\6612_b1 , \6612_b0 , \6613_b1 , \6613_b0 , \6614_b1 , \6614_b0 , \6615_b1 , \6615_b0 , \6616_b1 , \6616_b0 , 
		\6617_b1 , \6617_b0 , \6618_b1 , \6618_b0 , \6619_b1 , \6619_b0 , \6620_b1 , \6620_b0 , \6621_b1 , \6621_b0 , 
		\6622_b1 , \6622_b0 , \6623_b1 , \6623_b0 , \6624_b1 , \6624_b0 , \6625_b1 , \6625_b0 , \6626_b1 , \6626_b0 , 
		\6627_b1 , \6627_b0 , \6628_b1 , \6628_b0 , \6629_b1 , \6629_b0 , \6630_b1 , \6630_b0 , \6631_b1 , \6631_b0 , 
		\6632_b1 , \6632_b0 , \6633_b1 , \6633_b0 , \6634_b1 , \6634_b0 , \6635_b1 , \6635_b0 , \6636_b1 , \6636_b0 , 
		\6637_b1 , \6637_b0 , \6638_b1 , \6638_b0 , \6639_b1 , \6639_b0 , \6640_b1 , \6640_b0 , \6641_b1 , \6641_b0 , 
		\6642_b1 , \6642_b0 , \6643_b1 , \6643_b0 , \6644_b1 , \6644_b0 , \6645_b1 , \6645_b0 , \6646_b1 , \6646_b0 , 
		\6647_b1 , \6647_b0 , \6648_b1 , \6648_b0 , \6649_b1 , \6649_b0 , \6650_b1 , \6650_b0 , \6651_b1 , \6651_b0 , 
		\6652_b1 , \6652_b0 , \6653_b1 , \6653_b0 , \6654_b1 , \6654_b0 , \6655_b1 , \6655_b0 , \6656_b1 , \6656_b0 , 
		\6657_b1 , \6657_b0 , \6658_b1 , \6658_b0 , \6659_b1 , \6659_b0 , \6660_b1 , \6660_b0 , \6661_b1 , \6661_b0 , 
		\6662_b1 , \6662_b0 , \6663_b1 , \6663_b0 , \6664_b1 , \6664_b0 , \6665_b1 , \6665_b0 , \6666_b1 , \6666_b0 , 
		\6667_b1 , \6667_b0 , \6668_b1 , \6668_b0 , \6669_b1 , \6669_b0 , \6670_b1 , \6670_b0 , \6671_b1 , \6671_b0 , 
		\6672_b1 , \6672_b0 , \6673_b1 , \6673_b0 , \6674_b1 , \6674_b0 , \6675_b1 , \6675_b0 , \6676_b1 , \6676_b0 , 
		\6677_b1 , \6677_b0 , \6678_b1 , \6678_b0 , \6679_b1 , \6679_b0 , \6680_b1 , \6680_b0 , \6681_b1 , \6681_b0 , 
		\6682_b1 , \6682_b0 , \6683_b1 , \6683_b0 , \6684_b1 , \6684_b0 , \6685_b1 , \6685_b0 , \6686_b1 , \6686_b0 , 
		\6687_b1 , \6687_b0 , \6688_b1 , \6688_b0 , \6689_b1 , \6689_b0 , \6690_b1 , \6690_b0 , \6691_b1 , \6691_b0 , 
		\6692_b1 , \6692_b0 , \6693_b1 , \6693_b0 , \6694_b1 , \6694_b0 , \6695_b1 , \6695_b0 , \6696_b1 , \6696_b0 , 
		\6697_b1 , \6697_b0 , \6698_b1 , \6698_b0 , \6699_b1 , \6699_b0 , \6700_b1 , \6700_b0 , \6701_b1 , \6701_b0 , 
		\6702_b1 , \6702_b0 , \6703_b1 , \6703_b0 , \6704_b1 , \6704_b0 , \6705_b1 , \6705_b0 , \6706_b1 , \6706_b0 , 
		\6707_b1 , \6707_b0 , \6708_b1 , \6708_b0 , \6709_b1 , \6709_b0 , \6710_b1 , \6710_b0 , \6711_b1 , \6711_b0 , 
		\6712_b1 , \6712_b0 , \6713_b1 , \6713_b0 , \6714_b1 , \6714_b0 , \6715_b1 , \6715_b0 , \6716_b1 , \6716_b0 , 
		\6717_b1 , \6717_b0 , \6718_b1 , \6718_b0 , \6719_b1 , \6719_b0 , \6720_b1 , \6720_b0 , \6721_b1 , \6721_b0 , 
		\6722_b1 , \6722_b0 , \6723_b1 , \6723_b0 , \6724_b1 , \6724_b0 , \6725_b1 , \6725_b0 , \6726_b1 , \6726_b0 , 
		\6727_b1 , \6727_b0 , \6728_b1 , \6728_b0 , \6729_b1 , \6729_b0 , \6730_b1 , \6730_b0 , \6731_b1 , \6731_b0 , 
		\6732_b1 , \6732_b0 , \6733_b1 , \6733_b0 , \6734_b1 , \6734_b0 , \6735_b1 , \6735_b0 , \6736_b1 , \6736_b0 , 
		\6737_b1 , \6737_b0 , \6738_b1 , \6738_b0 , \6739_b1 , \6739_b0 , \6740_b1 , \6740_b0 , \6741_b1 , \6741_b0 , 
		\6742_b1 , \6742_b0 , \6743_b1 , \6743_b0 , \6744_b1 , \6744_b0 , \6745_b1 , \6745_b0 , \6746_b1 , \6746_b0 , 
		\6747_b1 , \6747_b0 , \6748_b1 , \6748_b0 , \6749_b1 , \6749_b0 , \6750_b1 , \6750_b0 , \6751_b1 , \6751_b0 , 
		\6752_b1 , \6752_b0 , \6753_b1 , \6753_b0 , \6754_b1 , \6754_b0 , \6755_b1 , \6755_b0 , \6756_b1 , \6756_b0 , 
		\6757_b1 , \6757_b0 , \6758_b1 , \6758_b0 , \6759_b1 , \6759_b0 , \6760_b1 , \6760_b0 , \6761_b1 , \6761_b0 , 
		\6762_b1 , \6762_b0 , \6763_b1 , \6763_b0 , \6764_b1 , \6764_b0 , \6765_b1 , \6765_b0 , \6766_b1 , \6766_b0 , 
		\6767_b1 , \6767_b0 , \6768_b1 , \6768_b0 , \6769_b1 , \6769_b0 , \6770_b1 , \6770_b0 , \6771_b1 , \6771_b0 , 
		\6772_b1 , \6772_b0 , \6773_b1 , \6773_b0 , \6774_b1 , \6774_b0 , \6775_b1 , \6775_b0 , \6776_b1 , \6776_b0 , 
		\6777_b1 , \6777_b0 , \6778_b1 , \6778_b0 , \6779_b1 , \6779_b0 , \6780_b1 , \6780_b0 , \6781_b1 , \6781_b0 , 
		\6782_b1 , \6782_b0 , \6783_b1 , \6783_b0 , \6784_b1 , \6784_b0 , \6785_b1 , \6785_b0 , \6786_b1 , \6786_b0 , 
		\6787_b1 , \6787_b0 , \6788_b1 , \6788_b0 , \6789_b1 , \6789_b0 , \6790_b1 , \6790_b0 , \6791_b1 , \6791_b0 , 
		\6792_b1 , \6792_b0 , \6793_b1 , \6793_b0 , \6794_b1 , \6794_b0 , \6795_b1 , \6795_b0 , \6796_b1 , \6796_b0 , 
		\6797_b1 , \6797_b0 , \6798_b1 , \6798_b0 , \6799_b1 , \6799_b0 , \6800_b1 , \6800_b0 , \6801_b1 , \6801_b0 , 
		\6802_b1 , \6802_b0 , \6803_b1 , \6803_b0 , \6804_b1 , \6804_b0 , \6805_b1 , \6805_b0 , \6806_b1 , \6806_b0 , 
		\6807_b1 , \6807_b0 , \6808_b1 , \6808_b0 , \6809_b1 , \6809_b0 , \6810_b1 , \6810_b0 , \6811_b1 , \6811_b0 , 
		\6812_b1 , \6812_b0 , \6813_b1 , \6813_b0 , \6814_b1 , \6814_b0 , \6815_b1 , \6815_b0 , \6816_b1 , \6816_b0 , 
		\6817_b1 , \6817_b0 , \6818_b1 , \6818_b0 , \6819_b1 , \6819_b0 , \6820_b1 , \6820_b0 , \6821_b1 , \6821_b0 , 
		\6822_b1 , \6822_b0 , \6823_b1 , \6823_b0 , \6824_b1 , \6824_b0 , \6825_b1 , \6825_b0 , \6826_b1 , \6826_b0 , 
		\6827_b1 , \6827_b0 , \6828_b1 , \6828_b0 , \6829_b1 , \6829_b0 , \6830_b1 , \6830_b0 , \6831_b1 , \6831_b0 , 
		\6832_b1 , \6832_b0 , \6833_b1 , \6833_b0 , \6834_b1 , \6834_b0 , \6835_b1 , \6835_b0 , \6836_b1 , \6836_b0 , 
		\6837_b1 , \6837_b0 , \6838_b1 , \6838_b0 , \6839_b1 , \6839_b0 , \6840_b1 , \6840_b0 , \6841_b1 , \6841_b0 , 
		\6842_b1 , \6842_b0 , \6843_b1 , \6843_b0 , \6844_b1 , \6844_b0 , \6845_b1 , \6845_b0 , \6846_b1 , \6846_b0 , 
		\6847_b1 , \6847_b0 , \6848_b1 , \6848_b0 , \6849_b1 , \6849_b0 , \6850_b1 , \6850_b0 , \6851_b1 , \6851_b0 , 
		\6852_b1 , \6852_b0 , \6853_b1 , \6853_b0 , \6854_b1 , \6854_b0 , \6855_b1 , \6855_b0 , \6856_b1 , \6856_b0 , 
		\6857_b1 , \6857_b0 , \6858_b1 , \6858_b0 , \6859_b1 , \6859_b0 , \6860_b1 , \6860_b0 , \6861_b1 , \6861_b0 , 
		\6862_b1 , \6862_b0 , \6863_b1 , \6863_b0 , \6864_b1 , \6864_b0 , \6865_b1 , \6865_b0 , \6866_b1 , \6866_b0 , 
		\6867_b1 , \6867_b0 , \6868_b1 , \6868_b0 , \6869_b1 , \6869_b0 , \6870_b1 , \6870_b0 , \6871_b1 , \6871_b0 , 
		\6872_b1 , \6872_b0 , \6873_b1 , \6873_b0 , \6874_b1 , \6874_b0 , \6875_b1 , \6875_b0 , \6876_b1 , \6876_b0 , 
		\6877_b1 , \6877_b0 , \6878_b1 , \6878_b0 , \6879_b1 , \6879_b0 , \6880_b1 , \6880_b0 , \6881_b1 , \6881_b0 , 
		\6882_b1 , \6882_b0 , \6883_b1 , \6883_b0 , \6884_b1 , \6884_b0 , \6885_b1 , \6885_b0 , \6886_b1 , \6886_b0 , 
		\6887_b1 , \6887_b0 , \6888_b1 , \6888_b0 , \6889_b1 , \6889_b0 , \6890_b1 , \6890_b0 , \6891_b1 , \6891_b0 , 
		\6892_b1 , \6892_b0 , \6893_b1 , \6893_b0 , \6894_b1 , \6894_b0 , \6895_b1 , \6895_b0 , \6896_b1 , \6896_b0 , 
		\6897_b1 , \6897_b0 , \6898_b1 , \6898_b0 , \6899_b1 , \6899_b0 , \6900_b1 , \6900_b0 , \6901_b1 , \6901_b0 , 
		\6902_b1 , \6902_b0 , \6903_b1 , \6903_b0 , \6904_b1 , \6904_b0 , \6905_b1 , \6905_b0 , \6906_b1 , \6906_b0 , 
		\6907_b1 , \6907_b0 , \6908_b1 , \6908_b0 , \6909_b1 , \6909_b0 , \6910_b1 , \6910_b0 , \6911_b1 , \6911_b0 , 
		\6912_b1 , \6912_b0 , \6913_b1 , \6913_b0 , \6914_b1 , \6914_b0 , \6915_b1 , \6915_b0 , \6916_b1 , \6916_b0 , 
		\6917_b1 , \6917_b0 , \6918_b1 , \6918_b0 , \6919_b1 , \6919_b0 , \6920_b1 , \6920_b0 , \6921_b1 , \6921_b0 , 
		\6922_b1 , \6922_b0 , \6923_b1 , \6923_b0 , \6924_b1 , \6924_b0 , \6925_b1 , \6925_b0 , \6926_b1 , \6926_b0 , 
		\6927_b1 , \6927_b0 , \6928_b1 , \6928_b0 , \6929_b1 , \6929_b0 , \6930_b1 , \6930_b0 , \6931_b1 , \6931_b0 , 
		\6932_b1 , \6932_b0 , \6933_b1 , \6933_b0 , \6934_b1 , \6934_b0 , \6935_b1 , \6935_b0 , \6936_b1 , \6936_b0 , 
		\6937_b1 , \6937_b0 , \6938_b1 , \6938_b0 , \6939_b1 , \6939_b0 , \6940_b1 , \6940_b0 , \6941_b1 , \6941_b0 , 
		\6942_b1 , \6942_b0 , \6943_b1 , \6943_b0 , \6944_b1 , \6944_b0 , \6945_b1 , \6945_b0 , \6946_b1 , \6946_b0 , 
		\6947_b1 , \6947_b0 , \6948_b1 , \6948_b0 , \6949_b1 , \6949_b0 , \6950_b1 , \6950_b0 , \6951_b1 , \6951_b0 , 
		\6952_b1 , \6952_b0 , \6953_b1 , \6953_b0 , \6954_b1 , \6954_b0 , \6955_b1 , \6955_b0 , \6956_b1 , \6956_b0 , 
		\6957_b1 , \6957_b0 , \6958_b1 , \6958_b0 , \6959_b1 , \6959_b0 , \6960_b1 , \6960_b0 , \6961_b1 , \6961_b0 , 
		\6962_b1 , \6962_b0 , \6963_b1 , \6963_b0 , \6964_b1 , \6964_b0 , \6965_b1 , \6965_b0 , \6966_b1 , \6966_b0 , 
		\6967_b1 , \6967_b0 , \6968_b1 , \6968_b0 , \6969_b1 , \6969_b0 , \6970_b1 , \6970_b0 , \6971_b1 , \6971_b0 , 
		\6972_b1 , \6972_b0 , \6973_b1 , \6973_b0 , \6974_b1 , \6974_b0 , \6975_b1 , \6975_b0 , \6976_b1 , \6976_b0 , 
		\6977_b1 , \6977_b0 , \6978_b1 , \6978_b0 , \6979_b1 , \6979_b0 , \6980_b1 , \6980_b0 , \6981_b1 , \6981_b0 , 
		\6982_b1 , \6982_b0 , \6983_b1 , \6983_b0 , \6984_b1 , \6984_b0 , \6985_b1 , \6985_b0 , \6986_b1 , \6986_b0 , 
		\6987_b1 , \6987_b0 , \6988_b1 , \6988_b0 , \6989_b1 , \6989_b0 , \6990_b1 , \6990_b0 , \6991_b1 , \6991_b0 , 
		\6992_b1 , \6992_b0 , \6993_b1 , \6993_b0 , \6994_b1 , \6994_b0 , \6995_b1 , \6995_b0 , \6996_b1 , \6996_b0 , 
		\6997_b1 , \6997_b0 , \6998_b1 , \6998_b0 , \6999_b1 , \6999_b0 , \7000_b1 , \7000_b0 , \7001_b1 , \7001_b0 , 
		\7002_b1 , \7002_b0 , \7003_b1 , \7003_b0 , \7004_b1 , \7004_b0 , \7005_b1 , \7005_b0 , \7006_b1 , \7006_b0 , 
		\7007_b1 , \7007_b0 , \7008_b1 , \7008_b0 , \7009_b1 , \7009_b0 , \7010_b1 , \7010_b0 , \7011_b1 , \7011_b0 , 
		\7012_b1 , \7012_b0 , \7013_b1 , \7013_b0 , \7014_b1 , \7014_b0 , \7015_b1 , \7015_b0 , \7016_b1 , \7016_b0 , 
		\7017_b1 , \7017_b0 , \7018_b1 , \7018_b0 , \7019_b1 , \7019_b0 , \7020_b1 , \7020_b0 , \7021_b1 , \7021_b0 , 
		\7022_b1 , \7022_b0 , \7023_b1 , \7023_b0 , \7024_b1 , \7024_b0 , \7025_b1 , \7025_b0 , \7026_b1 , \7026_b0 , 
		\7027_b1 , \7027_b0 , \7028_b1 , \7028_b0 , \7029_b1 , \7029_b0 , \7030_b1 , \7030_b0 , \7031_b1 , \7031_b0 , 
		\7032_b1 , \7032_b0 , \7033_b1 , \7033_b0 , \7034_b1 , \7034_b0 , \7035_b1 , \7035_b0 , \7036_b1 , \7036_b0 , 
		\7037_b1 , \7037_b0 , \7038_b1 , \7038_b0 , \7039_b1 , \7039_b0 , \7040_b1 , \7040_b0 , \7041_b1 , \7041_b0 , 
		\7042_b1 , \7042_b0 , \7043_b1 , \7043_b0 , \7044_b1 , \7044_b0 , \7045_b1 , \7045_b0 , \7046_b1 , \7046_b0 , 
		\7047_b1 , \7047_b0 , \7048_b1 , \7048_b0 , \7049_b1 , \7049_b0 , \7050_b1 , \7050_b0 , \7051_b1 , \7051_b0 , 
		\7052_b1 , \7052_b0 , \7053_b1 , \7053_b0 , \7054_b1 , \7054_b0 , \7055_b1 , \7055_b0 , \7056_b1 , \7056_b0 , 
		\7057_b1 , \7057_b0 , \7058_b1 , \7058_b0 , \7059_b1 , \7059_b0 , \7060_b1 , \7060_b0 , \7061_b1 , \7061_b0 , 
		\7062_b1 , \7062_b0 , \7063_b1 , \7063_b0 , \7064_b1 , \7064_b0 , \7065_b1 , \7065_b0 , \7066_b1 , \7066_b0 , 
		\7067_b1 , \7067_b0 , \7068_b1 , \7068_b0 , \7069_b1 , \7069_b0 , \7070_b1 , \7070_b0 , \7071_b1 , \7071_b0 , 
		\7072_b1 , \7072_b0 , \7073_b1 , \7073_b0 , \7074_b1 , \7074_b0 , \7075_b1 , \7075_b0 , \7076_b1 , \7076_b0 , 
		\7077_b1 , \7077_b0 , \7078_b1 , \7078_b0 , \7079_b1 , \7079_b0 , \7080_b1 , \7080_b0 , \7081_b1 , \7081_b0 , 
		\7082_b1 , \7082_b0 , \7083_b1 , \7083_b0 , \7084_b1 , \7084_b0 , \7085_b1 , \7085_b0 , \7086_b1 , \7086_b0 , 
		\7087_b1 , \7087_b0 , \7088_b1 , \7088_b0 , \7089_b1 , \7089_b0 , \7090_b1 , \7090_b0 , \7091_b1 , \7091_b0 , 
		\7092_b1 , \7092_b0 , \7093_b1 , \7093_b0 , \7094_b1 , \7094_b0 , \7095_b1 , \7095_b0 , \7096_b1 , \7096_b0 , 
		\7097_b1 , \7097_b0 , \7098_b1 , \7098_b0 , \7099_b1 , \7099_b0 , \7100_b1 , \7100_b0 , \7101_b1 , \7101_b0 , 
		\7102_b1 , \7102_b0 , \7103_b1 , \7103_b0 , \7104_b1 , \7104_b0 , \7105_b1 , \7105_b0 , \7106_b1 , \7106_b0 , 
		\7107_b1 , \7107_b0 , \7108_b1 , \7108_b0 , \7109_b1 , \7109_b0 , \7110_b1 , \7110_b0 , \7111_b1 , \7111_b0 , 
		\7112_b1 , \7112_b0 , \7113_b1 , \7113_b0 , \7114_b1 , \7114_b0 , \7115_b1 , \7115_b0 , \7116_b1 , \7116_b0 , 
		\7117_b1 , \7117_b0 , \7118_b1 , \7118_b0 , \7119_b1 , \7119_b0 , \7120_b1 , \7120_b0 , \7121_b1 , \7121_b0 , 
		\7122_b1 , \7122_b0 , \7123_b1 , \7123_b0 , \7124_b1 , \7124_b0 , \7125_b1 , \7125_b0 , \7126_b1 , \7126_b0 , 
		\7127_b1 , \7127_b0 , \7128_b1 , \7128_b0 , \7129_b1 , \7129_b0 , \7130_b1 , \7130_b0 , \7131_b1 , \7131_b0 , 
		\7132_b1 , \7132_b0 , \7133_b1 , \7133_b0 , \7134_b1 , \7134_b0 , \7135_b1 , \7135_b0 , \7136_b1 , \7136_b0 , 
		\7137_b1 , \7137_b0 , \7138_b1 , \7138_b0 , \7139_b1 , \7139_b0 , \7140_b1 , \7140_b0 , \7141_b1 , \7141_b0 , 
		\7142_b1 , \7142_b0 , \7143_b1 , \7143_b0 , \7144_b1 , \7144_b0 , \7145_b1 , \7145_b0 , \7146_b1 , \7146_b0 , 
		\7147_b1 , \7147_b0 , \7148_b1 , \7148_b0 , \7149_b1 , \7149_b0 , \7150_b1 , \7150_b0 , \7151_b1 , \7151_b0 , 
		\7152_b1 , \7152_b0 , \7153_b1 , \7153_b0 , \7154_b1 , \7154_b0 , \7155_b1 , \7155_b0 , \7156_b1 , \7156_b0 , 
		\7157_b1 , \7157_b0 , \7158_b1 , \7158_b0 , \7159_b1 , \7159_b0 , \7160_b1 , \7160_b0 , \7161_b1 , \7161_b0 , 
		\7162_b1 , \7162_b0 , \7163_b1 , \7163_b0 , \7164_b1 , \7164_b0 , \7165_b1 , \7165_b0 , \7166_b1 , \7166_b0 , 
		\7167_b1 , \7167_b0 , \7168_b1 , \7168_b0 , \7169_b1 , \7169_b0 , \7170_b1 , \7170_b0 , \7171_b1 , \7171_b0 , 
		\7172_b1 , \7172_b0 , \7173_b1 , \7173_b0 , \7174_b1 , \7174_b0 , \7175_b1 , \7175_b0 , \7176_b1 , \7176_b0 , 
		\7177_b1 , \7177_b0 , \7178_b1 , \7178_b0 , \7179_b1 , \7179_b0 , \7180_b1 , \7180_b0 , \7181_b1 , \7181_b0 , 
		\7182_b1 , \7182_b0 , \7183_b1 , \7183_b0 , \7184_b1 , \7184_b0 , \7185_b1 , \7185_b0 , \7186_b1 , \7186_b0 , 
		\7187_b1 , \7187_b0 , \7188_b1 , \7188_b0 , \7189_b1 , \7189_b0 , \7190_b1 , \7190_b0 , \7191_b1 , \7191_b0 , 
		\7192_b1 , \7192_b0 , \7193_b1 , \7193_b0 , \7194_b1 , \7194_b0 , \7195_b1 , \7195_b0 , \7196_b1 , \7196_b0 , 
		\7197_b1 , \7197_b0 , \7198_b1 , \7198_b0 , \7199_b1 , \7199_b0 , \7200_b1 , \7200_b0 , \7201_b1 , \7201_b0 , 
		\7202_b1 , \7202_b0 , \7203_b1 , \7203_b0 , \7204_b1 , \7204_b0 , \7205_b1 , \7205_b0 , \7206_b1 , \7206_b0 , 
		\7207_b1 , \7207_b0 , \7208_b1 , \7208_b0 , \7209_b1 , \7209_b0 , \7210_b1 , \7210_b0 , \7211_b1 , \7211_b0 , 
		\7212_b1 , \7212_b0 , \7213_b1 , \7213_b0 , \7214_b1 , \7214_b0 , \7215_b1 , \7215_b0 , \7216_b1 , \7216_b0 , 
		\7217_b1 , \7217_b0 , \7218_b1 , \7218_b0 , \7219_b1 , \7219_b0 , \7220_b1 , \7220_b0 , \7221_b1 , \7221_b0 , 
		\7222_b1 , \7222_b0 , \7223_b1 , \7223_b0 , \7224_b1 , \7224_b0 , \7225_b1 , \7225_b0 , \7226_b1 , \7226_b0 , 
		\7227_b1 , \7227_b0 , \7228_b1 , \7228_b0 , \7229_b1 , \7229_b0 , \7230_b1 , \7230_b0 , \7231_b1 , \7231_b0 , 
		\7232_b1 , \7232_b0 , \7233_b1 , \7233_b0 , \7234_b1 , \7234_b0 , \7235_b1 , \7235_b0 , \7236_b1 , \7236_b0 , 
		\7237_b1 , \7237_b0 , \7238_b1 , \7238_b0 , \7239_b1 , \7239_b0 , \7240_b1 , \7240_b0 , \7241_b1 , \7241_b0 , 
		\7242_b1 , \7242_b0 , \7243_b1 , \7243_b0 , \7244_b1 , \7244_b0 , \7245_b1 , \7245_b0 , \7246_b1 , \7246_b0 , 
		\7247_b1 , \7247_b0 , \7248_b1 , \7248_b0 , \7249_b1 , \7249_b0 , \7250_b1 , \7250_b0 , \7251_b1 , \7251_b0 , 
		\7252_b1 , \7252_b0 , \7253_b1 , \7253_b0 , \7254_b1 , \7254_b0 , \7255_b1 , \7255_b0 , \7256_b1 , \7256_b0 , 
		\7257_b1 , \7257_b0 , \7258_b1 , \7258_b0 , \7259_b1 , \7259_b0 , \7260_b1 , \7260_b0 , \7261_b1 , \7261_b0 , 
		\7262_b1 , \7262_b0 , \7263_b1 , \7263_b0 , \7264_b1 , \7264_b0 , \7265_b1 , \7265_b0 , \7266_b1 , \7266_b0 , 
		\7267_b1 , \7267_b0 , \7268_b1 , \7268_b0 , \7269_b1 , \7269_b0 , \7270_b1 , \7270_b0 , \7271_b1 , \7271_b0 , 
		\7272_b1 , \7272_b0 , \7273_b1 , \7273_b0 , \7274_b1 , \7274_b0 , \7275_b1 , \7275_b0 , \7276_b1 , \7276_b0 , 
		\7277_b1 , \7277_b0 , \7278_b1 , \7278_b0 , \7279_b1 , \7279_b0 , \7280_b1 , \7280_b0 , \7281_b1 , \7281_b0 , 
		\7282_b1 , \7282_b0 , \7283_b1 , \7283_b0 , \7284_b1 , \7284_b0 , \7285_b1 , \7285_b0 , \7286_b1 , \7286_b0 , 
		\7287_b1 , \7287_b0 , \7288_b1 , \7288_b0 , \7289_b1 , \7289_b0 , \7290_b1 , \7290_b0 , \7291_b1 , \7291_b0 , 
		\7292_b1 , \7292_b0 , \7293_b1 , \7293_b0 , \7294_b1 , \7294_b0 , \7295_b1 , \7295_b0 , \7296_b1 , \7296_b0 , 
		\7297_b1 , \7297_b0 , \7298_b1 , \7298_b0 , \7299_b1 , \7299_b0 , \7300_b1 , \7300_b0 , \7301_b1 , \7301_b0 , 
		\7302_b1 , \7302_b0 , \7303_b1 , \7303_b0 , \7304_b1 , \7304_b0 , \7305_b1 , \7305_b0 , \7306_b1 , \7306_b0 , 
		\7307_b1 , \7307_b0 , \7308_b1 , \7308_b0 , \7309_b1 , \7309_b0 , \7310_b1 , \7310_b0 , \7311_b1 , \7311_b0 , 
		\7312_b1 , \7312_b0 , \7313_b1 , \7313_b0 , \7314_b1 , \7314_b0 , \7315_b1 , \7315_b0 , \7316_b1 , \7316_b0 , 
		\7317_b1 , \7317_b0 , \7318_b1 , \7318_b0 , \7319_b1 , \7319_b0 , \7320_b1 , \7320_b0 , \7321_b1 , \7321_b0 , 
		\7322_b1 , \7322_b0 , \7323_b1 , \7323_b0 , \7324_b1 , \7324_b0 , \7325_b1 , \7325_b0 , \7326_b1 , \7326_b0 , 
		\7327_b1 , \7327_b0 , \7328_b1 , \7328_b0 , \7329_b1 , \7329_b0 , \7330_b1 , \7330_b0 , \7331_b1 , \7331_b0 , 
		\7332_b1 , \7332_b0 , \7333_b1 , \7333_b0 , \7334_b1 , \7334_b0 , \7335_b1 , \7335_b0 , \7336_b1 , \7336_b0 , 
		\7337_b1 , \7337_b0 , \7338_b1 , \7338_b0 , \7339_b1 , \7339_b0 , \7340_b1 , \7340_b0 , \7341_b1 , \7341_b0 , 
		\7342_b1 , \7342_b0 , \7343_b1 , \7343_b0 , \7344_b1 , \7344_b0 , \7345_b1 , \7345_b0 , \7346_b1 , \7346_b0 , 
		\7347_b1 , \7347_b0 , \7348_b1 , \7348_b0 , \7349_b1 , \7349_b0 , \7350_b1 , \7350_b0 , \7351_b1 , \7351_b0 , 
		\7352_b1 , \7352_b0 , \7353_b1 , \7353_b0 , \7354_b1 , \7354_b0 , \7355_b1 , \7355_b0 , \7356_b1 , \7356_b0 , 
		\7357_b1 , \7357_b0 , \7358_b1 , \7358_b0 , \7359_b1 , \7359_b0 , \7360_b1 , \7360_b0 , \7361_b1 , \7361_b0 , 
		\7362_b1 , \7362_b0 , \7363_b1 , \7363_b0 , \7364_b1 , \7364_b0 , \7365_b1 , \7365_b0 , \7366_b1 , \7366_b0 , 
		\7367_b1 , \7367_b0 , \7368_b1 , \7368_b0 , \7369_b1 , \7369_b0 , \7370_b1 , \7370_b0 , \7371_b1 , \7371_b0 , 
		\7372_b1 , \7372_b0 , \7373_b1 , \7373_b0 , \7374_b1 , \7374_b0 , \7375_b1 , \7375_b0 , \7376_b1 , \7376_b0 , 
		\7377_b1 , \7377_b0 , \7378_b1 , \7378_b0 , \7379_b1 , \7379_b0 , \7380_b1 , \7380_b0 , \7381_b1 , \7381_b0 , 
		\7382_b1 , \7382_b0 , \7383_b1 , \7383_b0 , \7384_b1 , \7384_b0 , \7385_b1 , \7385_b0 , \7386_b1 , \7386_b0 , 
		\7387_b1 , \7387_b0 , \7388_b1 , \7388_b0 , \7389_b1 , \7389_b0 , \7390_b1 , \7390_b0 , \7391_b1 , \7391_b0 , 
		\7392_b1 , \7392_b0 , \7393_b1 , \7393_b0 , \7394_b1 , \7394_b0 , \7395_b1 , \7395_b0 , \7396_b1 , \7396_b0 , 
		\7397_b1 , \7397_b0 , \7398_b1 , \7398_b0 , \7399_b1 , \7399_b0 , \7400_b1 , \7400_b0 , \7401_b1 , \7401_b0 , 
		\7402_b1 , \7402_b0 , \7403_b1 , \7403_b0 , \7404_b1 , \7404_b0 , \7405_b1 , \7405_b0 , \7406_b1 , \7406_b0 , 
		\7407_b1 , \7407_b0 , \7408_b1 , \7408_b0 , \7409_b1 , \7409_b0 , \7410_b1 , \7410_b0 , \7411_b1 , \7411_b0 , 
		\7412_b1 , \7412_b0 , \7413_b1 , \7413_b0 , \7414_b1 , \7414_b0 , \7415_b1 , \7415_b0 , \7416_b1 , \7416_b0 , 
		\7417_b1 , \7417_b0 , \7418_b1 , \7418_b0 , \7419_b1 , \7419_b0 , \7420_b1 , \7420_b0 , \7421_b1 , \7421_b0 , 
		\7422_b1 , \7422_b0 , \7423_b1 , \7423_b0 , \7424_b1 , \7424_b0 , \7425_b1 , \7425_b0 , \7426_b1 , \7426_b0 , 
		\7427_b1 , \7427_b0 , \7428_b1 , \7428_b0 , \7429_b1 , \7429_b0 , \7430_b1 , \7430_b0 , \7431_b1 , \7431_b0 , 
		\7432_b1 , \7432_b0 , \7433_b1 , \7433_b0 , \7434_b1 , \7434_b0 , \7435_b1 , \7435_b0 , \7436_b1 , \7436_b0 , 
		\7437_b1 , \7437_b0 , \7438_b1 , \7438_b0 , \7439_b1 , \7439_b0 , \7440_b1 , \7440_b0 , \7441_b1 , \7441_b0 , 
		\7442_b1 , \7442_b0 , \7443_b1 , \7443_b0 , \7444_b1 , \7444_b0 , \7445_b1 , \7445_b0 , \7446_b1 , \7446_b0 , 
		\7447_b1 , \7447_b0 , \7448_b1 , \7448_b0 , \7449_b1 , \7449_b0 , \7450_b1 , \7450_b0 , \7451_b1 , \7451_b0 , 
		\7452_b1 , \7452_b0 , \7453_b1 , \7453_b0 , \7454_b1 , \7454_b0 , \7455_b1 , \7455_b0 , \7456_b1 , \7456_b0 , 
		\7457_b1 , \7457_b0 , \7458_b1 , \7458_b0 , \7459_b1 , \7459_b0 , \7460_b1 , \7460_b0 , \7461_b1 , \7461_b0 , 
		\7462_b1 , \7462_b0 , \7463_b1 , \7463_b0 , \7464_b1 , \7464_b0 , \7465_b1 , \7465_b0 , \7466_b1 , \7466_b0 , 
		\7467_b1 , \7467_b0 , \7468_b1 , \7468_b0 , \7469_b1 , \7469_b0 , \7470_b1 , \7470_b0 , \7471_b1 , \7471_b0 , 
		\7472_b1 , \7472_b0 , \7473_b1 , \7473_b0 , \7474_b1 , \7474_b0 , \7475_b1 , \7475_b0 , \7476_b1 , \7476_b0 , 
		\7477_b1 , \7477_b0 , \7478_b1 , \7478_b0 , \7479_b1 , \7479_b0 , \7480_b1 , \7480_b0 , \7481_b1 , \7481_b0 , 
		\7482_b1 , \7482_b0 , \7483_b1 , \7483_b0 , \7484_b1 , \7484_b0 , \7485_b1 , \7485_b0 , \7486_b1 , \7486_b0 , 
		\7487_b1 , \7487_b0 , \7488_b1 , \7488_b0 , \7489_b1 , \7489_b0 , \7490_b1 , \7490_b0 , \7491_b1 , \7491_b0 , 
		\7492_b1 , \7492_b0 , \7493_b1 , \7493_b0 , \7494_b1 , \7494_b0 , \7495_b1 , \7495_b0 , \7496_b1 , \7496_b0 , 
		\7497_b1 , \7497_b0 , \7498_b1 , \7498_b0 , \7499_b1 , \7499_b0 , \7500_b1 , \7500_b0 , \7501_b1 , \7501_b0 , 
		\7502_b1 , \7502_b0 , \7503_b1 , \7503_b0 , \7504_b1 , \7504_b0 , \7505_b1 , \7505_b0 , \7506_b1 , \7506_b0 , 
		\7507_b1 , \7507_b0 , \7508_b1 , \7508_b0 , w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , 
		w_6 , w_7 , w_8 , w_9 , w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , 
		w_16 , w_17 , w_18 , w_19 , w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , 
		w_26 , w_27 , w_28 , w_29 , w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , 
		w_36 , w_37 , w_38 , w_39 , w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , 
		w_46 , w_47 , w_48 , w_49 , w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , 
		w_56 , w_57 , w_58 , w_59 , w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , 
		w_66 , w_67 , w_68 , w_69 , w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , 
		w_76 , w_77 , w_78 , w_79 , w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , 
		w_86 , w_87 , w_88 , w_89 , w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , 
		w_96 , w_97 , w_98 , w_99 , w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , 
		w_106 , w_107 , w_108 , w_109 , w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , 
		w_116 , w_117 , w_118 , w_119 , w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , 
		w_126 , w_127 , w_128 , w_129 , w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , 
		w_136 , w_137 , w_138 , w_139 , w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , 
		w_146 , w_147 , w_148 , w_149 , w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , 
		w_156 , w_157 , w_158 , w_159 , w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , 
		w_166 , w_167 , w_168 , w_169 , w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , 
		w_176 , w_177 , w_178 , w_179 , w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , 
		w_186 , w_187 , w_188 , w_189 , w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , 
		w_196 , w_197 , w_198 , w_199 , w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , 
		w_206 , w_207 , w_208 , w_209 , w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , 
		w_216 , w_217 , w_218 , w_219 , w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , 
		w_226 , w_227 , w_228 , w_229 , w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , 
		w_236 , w_237 , w_238 , w_239 , w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , 
		w_246 , w_247 , w_248 , w_249 , w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , 
		w_256 , w_257 , w_258 , w_259 , w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , 
		w_266 , w_267 , w_268 , w_269 , w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , 
		w_276 , w_277 , w_278 , w_279 , w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , 
		w_286 , w_287 , w_288 , w_289 , w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , 
		w_296 , w_297 , w_298 , w_299 , w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , 
		w_306 , w_307 , w_308 , w_309 , w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , 
		w_316 , w_317 , w_318 , w_319 , w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , 
		w_326 , w_327 , w_328 , w_329 , w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , 
		w_336 , w_337 , w_338 , w_339 , w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , 
		w_346 , w_347 , w_348 , w_349 , w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , 
		w_356 , w_357 , w_358 , w_359 , w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , 
		w_366 , w_367 , w_368 , w_369 , w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , 
		w_376 , w_377 , w_378 , w_379 , w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , 
		w_386 , w_387 , w_388 , w_389 , w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , 
		w_396 , w_397 , w_398 , w_399 , w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , 
		w_406 , w_407 , w_408 , w_409 , w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , 
		w_416 , w_417 , w_418 , w_419 , w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , 
		w_426 , w_427 , w_428 , w_429 , w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , 
		w_436 , w_437 , w_438 , w_439 , w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , 
		w_446 , w_447 , w_448 , w_449 , w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , 
		w_456 , w_457 , w_458 , w_459 , w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , 
		w_466 , w_467 , w_468 , w_469 , w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , 
		w_476 , w_477 , w_478 , w_479 , w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , 
		w_486 , w_487 , w_488 , w_489 , w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , 
		w_496 , w_497 , w_498 , w_499 , w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , 
		w_506 , w_507 , w_508 , w_509 , w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , 
		w_516 , w_517 , w_518 , w_519 , w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , 
		w_526 , w_527 , w_528 , w_529 , w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , 
		w_536 , w_537 , w_538 , w_539 , w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , 
		w_546 , w_547 , w_548 , w_549 , w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , 
		w_556 , w_557 , w_558 , w_559 , w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , 
		w_566 , w_567 , w_568 , w_569 , w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , 
		w_576 , w_577 , w_578 , w_579 , w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , 
		w_586 , w_587 , w_588 , w_589 , w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , 
		w_596 , w_597 , w_598 , w_599 , w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , 
		w_606 , w_607 , w_608 , w_609 , w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , 
		w_616 , w_617 , w_618 , w_619 , w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , 
		w_626 , w_627 , w_628 , w_629 , w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , 
		w_636 , w_637 , w_638 , w_639 , w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , 
		w_646 , w_647 , w_648 , w_649 , w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , 
		w_656 , w_657 , w_658 , w_659 , w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , 
		w_666 , w_667 , w_668 , w_669 , w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , 
		w_676 , w_677 , w_678 , w_679 , w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , 
		w_686 , w_687 , w_688 , w_689 , w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , 
		w_696 , w_697 , w_698 , w_699 , w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , 
		w_706 , w_707 , w_708 , w_709 , w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , 
		w_716 , w_717 , w_718 , w_719 , w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , 
		w_726 , w_727 , w_728 , w_729 , w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , 
		w_736 , w_737 , w_738 , w_739 , w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , 
		w_746 , w_747 , w_748 , w_749 , w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , 
		w_756 , w_757 , w_758 , w_759 , w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , 
		w_766 , w_767 , w_768 , w_769 , w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , 
		w_776 , w_777 , w_778 , w_779 , w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , 
		w_786 , w_787 , w_788 , w_789 , w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , 
		w_796 , w_797 , w_798 , w_799 , w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , 
		w_806 , w_807 , w_808 , w_809 , w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , 
		w_816 , w_817 , w_818 , w_819 , w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , 
		w_826 , w_827 , w_828 , w_829 , w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , 
		w_836 , w_837 , w_838 , w_839 , w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , 
		w_846 , w_847 , w_848 , w_849 , w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , 
		w_856 , w_857 , w_858 , w_859 , w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , 
		w_866 , w_867 , w_868 , w_869 , w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , 
		w_876 , w_877 , w_878 , w_879 , w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , 
		w_886 , w_887 , w_888 , w_889 , w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , 
		w_896 , w_897 , w_898 , w_899 , w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , 
		w_906 , w_907 , w_908 , w_909 , w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , 
		w_916 , w_917 , w_918 , w_919 , w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , 
		w_926 , w_927 , w_928 , w_929 , w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , 
		w_936 , w_937 , w_938 , w_939 , w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , 
		w_946 , w_947 , w_948 , w_949 , w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , 
		w_956 , w_957 , w_958 , w_959 , w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , 
		w_966 , w_967 , w_968 , w_969 , w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , 
		w_976 , w_977 , w_978 , w_979 , w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , 
		w_986 , w_987 , w_988 , w_989 , w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , 
		w_996 , w_997 , w_998 , w_999 , w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , 
		w_1006 , w_1007 , w_1008 , w_1009 , w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , 
		w_1016 , w_1017 , w_1018 , w_1019 , w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , 
		w_1026 , w_1027 , w_1028 , w_1029 , w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , 
		w_1036 , w_1037 , w_1038 , w_1039 , w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , 
		w_1046 , w_1047 , w_1048 , w_1049 , w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , 
		w_1056 , w_1057 , w_1058 , w_1059 , w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , 
		w_1066 , w_1067 , w_1068 , w_1069 , w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , 
		w_1076 , w_1077 , w_1078 , w_1079 , w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , 
		w_1086 , w_1087 , w_1088 , w_1089 , w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , 
		w_1096 , w_1097 , w_1098 , w_1099 , w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , 
		w_1106 , w_1107 , w_1108 , w_1109 , w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , 
		w_1116 , w_1117 , w_1118 , w_1119 , w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , 
		w_1126 , w_1127 , w_1128 , w_1129 , w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , 
		w_1136 , w_1137 , w_1138 , w_1139 , w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , 
		w_1146 , w_1147 , w_1148 , w_1149 , w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , 
		w_1156 , w_1157 , w_1158 , w_1159 , w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , 
		w_1166 , w_1167 , w_1168 , w_1169 , w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , 
		w_1176 , w_1177 , w_1178 , w_1179 , w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , 
		w_1186 , w_1187 , w_1188 , w_1189 , w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , 
		w_1196 , w_1197 , w_1198 , w_1199 , w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , 
		w_1206 , w_1207 , w_1208 , w_1209 , w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , 
		w_1216 , w_1217 , w_1218 , w_1219 , w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , 
		w_1226 , w_1227 , w_1228 , w_1229 , w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , 
		w_1236 , w_1237 , w_1238 , w_1239 , w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , 
		w_1246 , w_1247 , w_1248 , w_1249 , w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , 
		w_1256 , w_1257 , w_1258 , w_1259 , w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , 
		w_1266 , w_1267 , w_1268 , w_1269 , w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , 
		w_1276 , w_1277 , w_1278 , w_1279 , w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , 
		w_1286 , w_1287 , w_1288 , w_1289 , w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , 
		w_1296 , w_1297 , w_1298 , w_1299 , w_1300 , w_1301 , w_1302 , w_1303 , w_1304 , w_1305 , 
		w_1306 , w_1307 , w_1308 , w_1309 , w_1310 , w_1311 , w_1312 , w_1313 , w_1314 , w_1315 , 
		w_1316 , w_1317 , w_1318 , w_1319 , w_1320 , w_1321 , w_1322 , w_1323 , w_1324 , w_1325 , 
		w_1326 , w_1327 , w_1328 , w_1329 , w_1330 , w_1331 , w_1332 , w_1333 , w_1334 , w_1335 , 
		w_1336 , w_1337 , w_1338 , w_1339 , w_1340 , w_1341 , w_1342 , w_1343 , w_1344 , w_1345 , 
		w_1346 , w_1347 , w_1348 , w_1349 , w_1350 , w_1351 , w_1352 , w_1353 , w_1354 , w_1355 , 
		w_1356 , w_1357 , w_1358 , w_1359 , w_1360 , w_1361 , w_1362 , w_1363 , w_1364 , w_1365 , 
		w_1366 , w_1367 , w_1368 , w_1369 , w_1370 , w_1371 , w_1372 , w_1373 , w_1374 , w_1375 , 
		w_1376 , w_1377 , w_1378 , w_1379 , w_1380 , w_1381 , w_1382 , w_1383 , w_1384 , w_1385 , 
		w_1386 , w_1387 , w_1388 , w_1389 , w_1390 , w_1391 , w_1392 , w_1393 , w_1394 , w_1395 , 
		w_1396 , w_1397 , w_1398 , w_1399 , w_1400 , w_1401 , w_1402 , w_1403 , w_1404 , w_1405 , 
		w_1406 , w_1407 , w_1408 , w_1409 , w_1410 , w_1411 , w_1412 , w_1413 , w_1414 , w_1415 , 
		w_1416 , w_1417 , w_1418 , w_1419 , w_1420 , w_1421 , w_1422 , w_1423 , w_1424 , w_1425 , 
		w_1426 , w_1427 , w_1428 , w_1429 , w_1430 , w_1431 , w_1432 , w_1433 , w_1434 , w_1435 , 
		w_1436 , w_1437 , w_1438 , w_1439 , w_1440 , w_1441 , w_1442 , w_1443 , w_1444 , w_1445 , 
		w_1446 , w_1447 , w_1448 , w_1449 , w_1450 , w_1451 , w_1452 , w_1453 , w_1454 , w_1455 , 
		w_1456 , w_1457 , w_1458 , w_1459 , w_1460 , w_1461 , w_1462 , w_1463 , w_1464 , w_1465 , 
		w_1466 , w_1467 , w_1468 , w_1469 , w_1470 , w_1471 , w_1472 , w_1473 , w_1474 , w_1475 , 
		w_1476 , w_1477 , w_1478 , w_1479 , w_1480 , w_1481 , w_1482 , w_1483 , w_1484 , w_1485 , 
		w_1486 , w_1487 , w_1488 , w_1489 , w_1490 , w_1491 , w_1492 , w_1493 , w_1494 , w_1495 , 
		w_1496 , w_1497 , w_1498 , w_1499 , w_1500 , w_1501 , w_1502 , w_1503 , w_1504 , w_1505 , 
		w_1506 , w_1507 , w_1508 , w_1509 , w_1510 , w_1511 , w_1512 , w_1513 , w_1514 , w_1515 , 
		w_1516 , w_1517 , w_1518 , w_1519 , w_1520 , w_1521 , w_1522 , w_1523 , w_1524 , w_1525 , 
		w_1526 , w_1527 , w_1528 , w_1529 , w_1530 , w_1531 , w_1532 , w_1533 , w_1534 , w_1535 , 
		w_1536 , w_1537 , w_1538 , w_1539 , w_1540 , w_1541 , w_1542 , w_1543 , w_1544 , w_1545 , 
		w_1546 , w_1547 , w_1548 , w_1549 , w_1550 , w_1551 , w_1552 , w_1553 , w_1554 , w_1555 , 
		w_1556 , w_1557 , w_1558 , w_1559 , w_1560 , w_1561 , w_1562 , w_1563 , w_1564 , w_1565 , 
		w_1566 , w_1567 , w_1568 , w_1569 , w_1570 , w_1571 , w_1572 , w_1573 , w_1574 , w_1575 , 
		w_1576 , w_1577 , w_1578 , w_1579 , w_1580 , w_1581 , w_1582 , w_1583 , w_1584 , w_1585 , 
		w_1586 , w_1587 , w_1588 , w_1589 , w_1590 , w_1591 , w_1592 , w_1593 , w_1594 , w_1595 , 
		w_1596 , w_1597 , w_1598 , w_1599 , w_1600 , w_1601 , w_1602 , w_1603 , w_1604 , w_1605 , 
		w_1606 , w_1607 , w_1608 , w_1609 , w_1610 , w_1611 , w_1612 , w_1613 , w_1614 , w_1615 , 
		w_1616 , w_1617 , w_1618 , w_1619 , w_1620 , w_1621 , w_1622 , w_1623 , w_1624 , w_1625 , 
		w_1626 , w_1627 , w_1628 , w_1629 , w_1630 , w_1631 , w_1632 , w_1633 , w_1634 , w_1635 , 
		w_1636 , w_1637 , w_1638 , w_1639 , w_1640 , w_1641 , w_1642 , w_1643 , w_1644 , w_1645 , 
		w_1646 , w_1647 , w_1648 , w_1649 , w_1650 , w_1651 , w_1652 , w_1653 , w_1654 , w_1655 , 
		w_1656 , w_1657 , w_1658 , w_1659 , w_1660 , w_1661 , w_1662 , w_1663 , w_1664 , w_1665 , 
		w_1666 , w_1667 , w_1668 , w_1669 , w_1670 , w_1671 , w_1672 , w_1673 , w_1674 , w_1675 , 
		w_1676 , w_1677 , w_1678 , w_1679 , w_1680 , w_1681 , w_1682 , w_1683 , w_1684 , w_1685 , 
		w_1686 , w_1687 , w_1688 , w_1689 , w_1690 , w_1691 , w_1692 , w_1693 , w_1694 , w_1695 , 
		w_1696 , w_1697 , w_1698 , w_1699 , w_1700 , w_1701 , w_1702 , w_1703 , w_1704 , w_1705 , 
		w_1706 , w_1707 , w_1708 , w_1709 , w_1710 , w_1711 , w_1712 , w_1713 , w_1714 , w_1715 , 
		w_1716 , w_1717 , w_1718 , w_1719 , w_1720 , w_1721 , w_1722 , w_1723 , w_1724 , w_1725 , 
		w_1726 , w_1727 , w_1728 , w_1729 , w_1730 , w_1731 , w_1732 , w_1733 , w_1734 , w_1735 , 
		w_1736 , w_1737 , w_1738 , w_1739 , w_1740 , w_1741 , w_1742 , w_1743 , w_1744 , w_1745 , 
		w_1746 , w_1747 , w_1748 , w_1749 , w_1750 , w_1751 , w_1752 , w_1753 , w_1754 , w_1755 , 
		w_1756 , w_1757 , w_1758 , w_1759 , w_1760 , w_1761 , w_1762 , w_1763 , w_1764 , w_1765 , 
		w_1766 , w_1767 , w_1768 , w_1769 , w_1770 , w_1771 , w_1772 , w_1773 , w_1774 , w_1775 , 
		w_1776 , w_1777 , w_1778 , w_1779 , w_1780 , w_1781 , w_1782 , w_1783 , w_1784 , w_1785 , 
		w_1786 , w_1787 , w_1788 , w_1789 , w_1790 , w_1791 , w_1792 , w_1793 , w_1794 , w_1795 , 
		w_1796 , w_1797 , w_1798 , w_1799 , w_1800 , w_1801 , w_1802 , w_1803 , w_1804 , w_1805 , 
		w_1806 , w_1807 , w_1808 , w_1809 , w_1810 , w_1811 , w_1812 , w_1813 , w_1814 , w_1815 , 
		w_1816 , w_1817 , w_1818 , w_1819 , w_1820 , w_1821 , w_1822 , w_1823 , w_1824 , w_1825 , 
		w_1826 , w_1827 , w_1828 , w_1829 , w_1830 , w_1831 , w_1832 , w_1833 , w_1834 , w_1835 , 
		w_1836 , w_1837 , w_1838 , w_1839 , w_1840 , w_1841 , w_1842 , w_1843 , w_1844 , w_1845 , 
		w_1846 , w_1847 , w_1848 , w_1849 , w_1850 , w_1851 , w_1852 , w_1853 , w_1854 , w_1855 , 
		w_1856 , w_1857 , w_1858 , w_1859 , w_1860 , w_1861 , w_1862 , w_1863 , w_1864 , w_1865 , 
		w_1866 , w_1867 , w_1868 , w_1869 , w_1870 , w_1871 , w_1872 , w_1873 , w_1874 , w_1875 , 
		w_1876 , w_1877 , w_1878 , w_1879 , w_1880 , w_1881 , w_1882 , w_1883 , w_1884 , w_1885 , 
		w_1886 , w_1887 , w_1888 , w_1889 , w_1890 , w_1891 , w_1892 , w_1893 , w_1894 , w_1895 , 
		w_1896 , w_1897 , w_1898 , w_1899 , w_1900 , w_1901 , w_1902 , w_1903 , w_1904 , w_1905 , 
		w_1906 , w_1907 , w_1908 , w_1909 , w_1910 , w_1911 , w_1912 , w_1913 , w_1914 , w_1915 , 
		w_1916 , w_1917 , w_1918 , w_1919 , w_1920 , w_1921 , w_1922 , w_1923 , w_1924 , w_1925 , 
		w_1926 , w_1927 , w_1928 , w_1929 , w_1930 , w_1931 , w_1932 , w_1933 , w_1934 , w_1935 , 
		w_1936 , w_1937 , w_1938 , w_1939 , w_1940 , w_1941 , w_1942 , w_1943 , w_1944 , w_1945 , 
		w_1946 , w_1947 , w_1948 , w_1949 , w_1950 , w_1951 , w_1952 , w_1953 , w_1954 , w_1955 , 
		w_1956 , w_1957 , w_1958 , w_1959 , w_1960 , w_1961 , w_1962 , w_1963 , w_1964 , w_1965 , 
		w_1966 , w_1967 , w_1968 , w_1969 , w_1970 , w_1971 , w_1972 , w_1973 , w_1974 , w_1975 , 
		w_1976 , w_1977 , w_1978 , w_1979 , w_1980 , w_1981 , w_1982 , w_1983 , w_1984 , w_1985 , 
		w_1986 , w_1987 , w_1988 , w_1989 , w_1990 , w_1991 , w_1992 , w_1993 , w_1994 , w_1995 , 
		w_1996 , w_1997 , w_1998 , w_1999 , w_2000 , w_2001 , w_2002 , w_2003 , w_2004 , w_2005 , 
		w_2006 , w_2007 , w_2008 , w_2009 , w_2010 , w_2011 , w_2012 , w_2013 , w_2014 , w_2015 , 
		w_2016 , w_2017 , w_2018 , w_2019 , w_2020 , w_2021 , w_2022 , w_2023 , w_2024 , w_2025 , 
		w_2026 , w_2027 , w_2028 , w_2029 , w_2030 , w_2031 , w_2032 , w_2033 , w_2034 , w_2035 , 
		w_2036 , w_2037 , w_2038 , w_2039 , w_2040 , w_2041 , w_2042 , w_2043 , w_2044 , w_2045 , 
		w_2046 , w_2047 , w_2048 , w_2049 , w_2050 , w_2051 , w_2052 , w_2053 , w_2054 , w_2055 , 
		w_2056 , w_2057 , w_2058 , w_2059 , w_2060 , w_2061 , w_2062 , w_2063 , w_2064 , w_2065 , 
		w_2066 , w_2067 , w_2068 , w_2069 , w_2070 , w_2071 , w_2072 , w_2073 , w_2074 , w_2075 , 
		w_2076 , w_2077 , w_2078 , w_2079 , w_2080 , w_2081 , w_2082 , w_2083 , w_2084 , w_2085 , 
		w_2086 , w_2087 , w_2088 , w_2089 , w_2090 , w_2091 , w_2092 , w_2093 , w_2094 , w_2095 , 
		w_2096 , w_2097 , w_2098 , w_2099 , w_2100 , w_2101 , w_2102 , w_2103 , w_2104 , w_2105 , 
		w_2106 , w_2107 , w_2108 , w_2109 , w_2110 , w_2111 , w_2112 , w_2113 , w_2114 , w_2115 , 
		w_2116 , w_2117 , w_2118 , w_2119 , w_2120 , w_2121 , w_2122 , w_2123 , w_2124 , w_2125 , 
		w_2126 , w_2127 , w_2128 , w_2129 , w_2130 , w_2131 , w_2132 , w_2133 , w_2134 , w_2135 , 
		w_2136 , w_2137 , w_2138 , w_2139 , w_2140 , w_2141 , w_2142 , w_2143 , w_2144 , w_2145 , 
		w_2146 , w_2147 , w_2148 , w_2149 , w_2150 , w_2151 , w_2152 , w_2153 , w_2154 , w_2155 , 
		w_2156 , w_2157 , w_2158 , w_2159 , w_2160 , w_2161 , w_2162 , w_2163 , w_2164 , w_2165 , 
		w_2166 , w_2167 , w_2168 , w_2169 , w_2170 , w_2171 , w_2172 , w_2173 , w_2174 , w_2175 , 
		w_2176 , w_2177 , w_2178 , w_2179 , w_2180 , w_2181 , w_2182 , w_2183 , w_2184 , w_2185 , 
		w_2186 , w_2187 , w_2188 , w_2189 , w_2190 , w_2191 , w_2192 , w_2193 , w_2194 , w_2195 , 
		w_2196 , w_2197 , w_2198 , w_2199 , w_2200 , w_2201 , w_2202 , w_2203 , w_2204 , w_2205 , 
		w_2206 , w_2207 , w_2208 , w_2209 , w_2210 , w_2211 , w_2212 , w_2213 , w_2214 , w_2215 , 
		w_2216 , w_2217 , w_2218 , w_2219 , w_2220 , w_2221 , w_2222 , w_2223 , w_2224 , w_2225 , 
		w_2226 , w_2227 , w_2228 , w_2229 , w_2230 , w_2231 , w_2232 , w_2233 , w_2234 , w_2235 , 
		w_2236 , w_2237 , w_2238 , w_2239 , w_2240 , w_2241 , w_2242 , w_2243 , w_2244 , w_2245 , 
		w_2246 , w_2247 , w_2248 , w_2249 , w_2250 , w_2251 , w_2252 , w_2253 , w_2254 , w_2255 , 
		w_2256 , w_2257 , w_2258 , w_2259 , w_2260 , w_2261 , w_2262 , w_2263 , w_2264 , w_2265 , 
		w_2266 , w_2267 , w_2268 , w_2269 , w_2270 , w_2271 , w_2272 , w_2273 , w_2274 , w_2275 , 
		w_2276 , w_2277 , w_2278 , w_2279 , w_2280 , w_2281 , w_2282 , w_2283 , w_2284 , w_2285 , 
		w_2286 , w_2287 , w_2288 , w_2289 , w_2290 , w_2291 , w_2292 , w_2293 , w_2294 , w_2295 , 
		w_2296 , w_2297 , w_2298 , w_2299 , w_2300 , w_2301 , w_2302 , w_2303 , w_2304 , w_2305 , 
		w_2306 , w_2307 , w_2308 , w_2309 , w_2310 , w_2311 , w_2312 , w_2313 , w_2314 , w_2315 , 
		w_2316 , w_2317 , w_2318 , w_2319 , w_2320 , w_2321 , w_2322 , w_2323 , w_2324 , w_2325 , 
		w_2326 , w_2327 , w_2328 , w_2329 , w_2330 , w_2331 , w_2332 , w_2333 , w_2334 , w_2335 , 
		w_2336 , w_2337 , w_2338 , w_2339 , w_2340 , w_2341 , w_2342 , w_2343 , w_2344 , w_2345 , 
		w_2346 , w_2347 , w_2348 , w_2349 , w_2350 , w_2351 , w_2352 , w_2353 , w_2354 , w_2355 , 
		w_2356 , w_2357 , w_2358 , w_2359 , w_2360 , w_2361 , w_2362 , w_2363 , w_2364 , w_2365 , 
		w_2366 , w_2367 , w_2368 , w_2369 , w_2370 , w_2371 , w_2372 , w_2373 , w_2374 , w_2375 , 
		w_2376 , w_2377 , w_2378 , w_2379 , w_2380 , w_2381 , w_2382 , w_2383 , w_2384 , w_2385 , 
		w_2386 , w_2387 , w_2388 , w_2389 , w_2390 , w_2391 , w_2392 , w_2393 , w_2394 , w_2395 , 
		w_2396 , w_2397 , w_2398 , w_2399 , w_2400 , w_2401 , w_2402 , w_2403 , w_2404 , w_2405 , 
		w_2406 , w_2407 , w_2408 , w_2409 , w_2410 , w_2411 , w_2412 , w_2413 , w_2414 , w_2415 , 
		w_2416 , w_2417 , w_2418 , w_2419 , w_2420 , w_2421 , w_2422 , w_2423 , w_2424 , w_2425 , 
		w_2426 , w_2427 , w_2428 , w_2429 , w_2430 , w_2431 , w_2432 , w_2433 , w_2434 , w_2435 , 
		w_2436 , w_2437 , w_2438 , w_2439 , w_2440 , w_2441 , w_2442 , w_2443 , w_2444 , w_2445 , 
		w_2446 , w_2447 , w_2448 , w_2449 , w_2450 , w_2451 , w_2452 , w_2453 , w_2454 , w_2455 , 
		w_2456 , w_2457 , w_2458 , w_2459 , w_2460 , w_2461 , w_2462 , w_2463 , w_2464 , w_2465 , 
		w_2466 , w_2467 , w_2468 , w_2469 , w_2470 , w_2471 , w_2472 , w_2473 , w_2474 , w_2475 , 
		w_2476 , w_2477 , w_2478 , w_2479 , w_2480 , w_2481 , w_2482 , w_2483 , w_2484 , w_2485 , 
		w_2486 , w_2487 , w_2488 , w_2489 , w_2490 , w_2491 , w_2492 , w_2493 , w_2494 , w_2495 , 
		w_2496 , w_2497 , w_2498 , w_2499 , w_2500 , w_2501 , w_2502 , w_2503 , w_2504 , w_2505 , 
		w_2506 , w_2507 , w_2508 , w_2509 , w_2510 , w_2511 , w_2512 , w_2513 , w_2514 , w_2515 , 
		w_2516 , w_2517 , w_2518 , w_2519 , w_2520 , w_2521 , w_2522 , w_2523 , w_2524 , w_2525 , 
		w_2526 , w_2527 , w_2528 , w_2529 , w_2530 , w_2531 , w_2532 , w_2533 , w_2534 , w_2535 , 
		w_2536 , w_2537 , w_2538 , w_2539 , w_2540 , w_2541 , w_2542 , w_2543 , w_2544 , w_2545 , 
		w_2546 , w_2547 , w_2548 , w_2549 , w_2550 , w_2551 , w_2552 , w_2553 , w_2554 , w_2555 , 
		w_2556 , w_2557 , w_2558 , w_2559 , w_2560 , w_2561 , w_2562 , w_2563 , w_2564 , w_2565 , 
		w_2566 , w_2567 , w_2568 , w_2569 , w_2570 , w_2571 , w_2572 , w_2573 , w_2574 , w_2575 , 
		w_2576 , w_2577 , w_2578 , w_2579 , w_2580 , w_2581 , w_2582 , w_2583 , w_2584 , w_2585 , 
		w_2586 , w_2587 , w_2588 , w_2589 , w_2590 , w_2591 , w_2592 , w_2593 , w_2594 , w_2595 , 
		w_2596 , w_2597 , w_2598 , w_2599 , w_2600 , w_2601 , w_2602 , w_2603 , w_2604 , w_2605 , 
		w_2606 , w_2607 , w_2608 , w_2609 , w_2610 , w_2611 , w_2612 , w_2613 , w_2614 , w_2615 , 
		w_2616 , w_2617 , w_2618 , w_2619 , w_2620 , w_2621 , w_2622 , w_2623 , w_2624 , w_2625 , 
		w_2626 , w_2627 , w_2628 , w_2629 , w_2630 , w_2631 , w_2632 , w_2633 , w_2634 , w_2635 , 
		w_2636 , w_2637 , w_2638 , w_2639 , w_2640 , w_2641 , w_2642 , w_2643 , w_2644 , w_2645 , 
		w_2646 , w_2647 , w_2648 , w_2649 , w_2650 , w_2651 , w_2652 , w_2653 , w_2654 , w_2655 , 
		w_2656 , w_2657 , w_2658 , w_2659 , w_2660 , w_2661 , w_2662 , w_2663 , w_2664 , w_2665 , 
		w_2666 , w_2667 , w_2668 , w_2669 , w_2670 , w_2671 , w_2672 , w_2673 , w_2674 , w_2675 , 
		w_2676 , w_2677 , w_2678 , w_2679 , w_2680 , w_2681 , w_2682 , w_2683 , w_2684 , w_2685 , 
		w_2686 , w_2687 , w_2688 , w_2689 , w_2690 , w_2691 , w_2692 , w_2693 , w_2694 , w_2695 , 
		w_2696 , w_2697 , w_2698 , w_2699 , w_2700 , w_2701 , w_2702 , w_2703 , w_2704 , w_2705 , 
		w_2706 , w_2707 , w_2708 , w_2709 , w_2710 , w_2711 , w_2712 , w_2713 , w_2714 , w_2715 , 
		w_2716 , w_2717 , w_2718 , w_2719 , w_2720 , w_2721 , w_2722 , w_2723 , w_2724 , w_2725 , 
		w_2726 , w_2727 , w_2728 , w_2729 , w_2730 , w_2731 , w_2732 , w_2733 , w_2734 , w_2735 , 
		w_2736 , w_2737 , w_2738 , w_2739 , w_2740 , w_2741 , w_2742 , w_2743 , w_2744 , w_2745 , 
		w_2746 , w_2747 , w_2748 , w_2749 , w_2750 , w_2751 , w_2752 , w_2753 , w_2754 , w_2755 , 
		w_2756 , w_2757 , w_2758 , w_2759 , w_2760 , w_2761 , w_2762 , w_2763 , w_2764 , w_2765 , 
		w_2766 , w_2767 , w_2768 , w_2769 , w_2770 , w_2771 , w_2772 , w_2773 , w_2774 , w_2775 , 
		w_2776 , w_2777 , w_2778 , w_2779 , w_2780 , w_2781 , w_2782 , w_2783 , w_2784 , w_2785 , 
		w_2786 , w_2787 , w_2788 , w_2789 , w_2790 , w_2791 , w_2792 , w_2793 , w_2794 , w_2795 , 
		w_2796 , w_2797 , w_2798 , w_2799 , w_2800 , w_2801 , w_2802 , w_2803 , w_2804 , w_2805 , 
		w_2806 , w_2807 , w_2808 , w_2809 , w_2810 , w_2811 , w_2812 , w_2813 , w_2814 , w_2815 , 
		w_2816 , w_2817 , w_2818 , w_2819 , w_2820 , w_2821 , w_2822 , w_2823 , w_2824 , w_2825 , 
		w_2826 , w_2827 , w_2828 , w_2829 , w_2830 , w_2831 , w_2832 , w_2833 , w_2834 , w_2835 , 
		w_2836 , w_2837 , w_2838 , w_2839 , w_2840 , w_2841 , w_2842 , w_2843 , w_2844 , w_2845 , 
		w_2846 , w_2847 , w_2848 , w_2849 , w_2850 , w_2851 , w_2852 , w_2853 , w_2854 , w_2855 , 
		w_2856 , w_2857 , w_2858 , w_2859 , w_2860 , w_2861 , w_2862 , w_2863 , w_2864 , w_2865 , 
		w_2866 , w_2867 , w_2868 , w_2869 , w_2870 , w_2871 , w_2872 , w_2873 , w_2874 , w_2875 , 
		w_2876 , w_2877 , w_2878 , w_2879 , w_2880 , w_2881 , w_2882 , w_2883 , w_2884 , w_2885 , 
		w_2886 , w_2887 , w_2888 , w_2889 , w_2890 , w_2891 , w_2892 , w_2893 , w_2894 , w_2895 , 
		w_2896 , w_2897 , w_2898 , w_2899 , w_2900 , w_2901 , w_2902 , w_2903 , w_2904 , w_2905 , 
		w_2906 , w_2907 , w_2908 , w_2909 , w_2910 , w_2911 , w_2912 , w_2913 , w_2914 , w_2915 , 
		w_2916 , w_2917 , w_2918 , w_2919 , w_2920 , w_2921 , w_2922 , w_2923 , w_2924 , w_2925 , 
		w_2926 , w_2927 , w_2928 , w_2929 , w_2930 , w_2931 , w_2932 , w_2933 , w_2934 , w_2935 , 
		w_2936 , w_2937 , w_2938 , w_2939 , w_2940 , w_2941 , w_2942 , w_2943 , w_2944 , w_2945 , 
		w_2946 , w_2947 , w_2948 , w_2949 , w_2950 , w_2951 , w_2952 , w_2953 , w_2954 , w_2955 , 
		w_2956 , w_2957 , w_2958 , w_2959 , w_2960 , w_2961 , w_2962 , w_2963 , w_2964 , w_2965 , 
		w_2966 , w_2967 , w_2968 , w_2969 , w_2970 , w_2971 , w_2972 , w_2973 , w_2974 , w_2975 , 
		w_2976 , w_2977 , w_2978 , w_2979 , w_2980 , w_2981 , w_2982 , w_2983 , w_2984 , w_2985 , 
		w_2986 , w_2987 , w_2988 , w_2989 , w_2990 , w_2991 , w_2992 , w_2993 , w_2994 , w_2995 , 
		w_2996 , w_2997 , w_2998 , w_2999 , w_3000 , w_3001 , w_3002 , w_3003 , w_3004 , w_3005 , 
		w_3006 , w_3007 , w_3008 , w_3009 , w_3010 , w_3011 , w_3012 , w_3013 , w_3014 , w_3015 , 
		w_3016 , w_3017 , w_3018 , w_3019 , w_3020 , w_3021 , w_3022 , w_3023 , w_3024 , w_3025 , 
		w_3026 , w_3027 , w_3028 , w_3029 , w_3030 , w_3031 , w_3032 , w_3033 , w_3034 , w_3035 , 
		w_3036 , w_3037 , w_3038 , w_3039 , w_3040 , w_3041 , w_3042 , w_3043 , w_3044 , w_3045 , 
		w_3046 , w_3047 , w_3048 , w_3049 , w_3050 , w_3051 , w_3052 , w_3053 , w_3054 , w_3055 , 
		w_3056 , w_3057 , w_3058 , w_3059 , w_3060 , w_3061 , w_3062 , w_3063 , w_3064 , w_3065 , 
		w_3066 , w_3067 , w_3068 , w_3069 , w_3070 , w_3071 , w_3072 , w_3073 , w_3074 , w_3075 , 
		w_3076 , w_3077 , w_3078 , w_3079 , w_3080 , w_3081 , w_3082 , w_3083 , w_3084 , w_3085 , 
		w_3086 , w_3087 , w_3088 , w_3089 , w_3090 , w_3091 , w_3092 , w_3093 , w_3094 , w_3095 , 
		w_3096 , w_3097 , w_3098 , w_3099 , w_3100 , w_3101 , w_3102 , w_3103 , w_3104 , w_3105 , 
		w_3106 , w_3107 , w_3108 , w_3109 , w_3110 , w_3111 , w_3112 , w_3113 , w_3114 , w_3115 , 
		w_3116 , w_3117 , w_3118 , w_3119 , w_3120 , w_3121 , w_3122 , w_3123 , w_3124 , w_3125 , 
		w_3126 , w_3127 , w_3128 , w_3129 , w_3130 , w_3131 , w_3132 , w_3133 , w_3134 , w_3135 , 
		w_3136 , w_3137 , w_3138 , w_3139 , w_3140 , w_3141 , w_3142 , w_3143 , w_3144 , w_3145 , 
		w_3146 , w_3147 , w_3148 , w_3149 , w_3150 , w_3151 , w_3152 , w_3153 , w_3154 , w_3155 , 
		w_3156 , w_3157 , w_3158 , w_3159 , w_3160 , w_3161 , w_3162 , w_3163 , w_3164 , w_3165 , 
		w_3166 , w_3167 , w_3168 , w_3169 , w_3170 , w_3171 , w_3172 , w_3173 , w_3174 , w_3175 , 
		w_3176 , w_3177 , w_3178 , w_3179 , w_3180 , w_3181 , w_3182 , w_3183 , w_3184 , w_3185 , 
		w_3186 , w_3187 , w_3188 , w_3189 , w_3190 , w_3191 , w_3192 , w_3193 , w_3194 , w_3195 , 
		w_3196 , w_3197 , w_3198 , w_3199 , w_3200 , w_3201 , w_3202 , w_3203 , w_3204 , w_3205 , 
		w_3206 , w_3207 , w_3208 , w_3209 , w_3210 , w_3211 , w_3212 , w_3213 , w_3214 , w_3215 , 
		w_3216 , w_3217 , w_3218 , w_3219 , w_3220 , w_3221 , w_3222 , w_3223 , w_3224 , w_3225 , 
		w_3226 , w_3227 , w_3228 , w_3229 , w_3230 , w_3231 , w_3232 , w_3233 , w_3234 , w_3235 , 
		w_3236 , w_3237 , w_3238 , w_3239 , w_3240 , w_3241 , w_3242 , w_3243 , w_3244 , w_3245 , 
		w_3246 , w_3247 , w_3248 , w_3249 , w_3250 , w_3251 , w_3252 , w_3253 , w_3254 , w_3255 , 
		w_3256 , w_3257 , w_3258 , w_3259 , w_3260 , w_3261 , w_3262 , w_3263 , w_3264 , w_3265 , 
		w_3266 , w_3267 , w_3268 , w_3269 , w_3270 , w_3271 , w_3272 , w_3273 , w_3274 , w_3275 , 
		w_3276 , w_3277 , w_3278 , w_3279 , w_3280 , w_3281 , w_3282 , w_3283 , w_3284 , w_3285 , 
		w_3286 , w_3287 , w_3288 , w_3289 , w_3290 , w_3291 , w_3292 , w_3293 , w_3294 , w_3295 , 
		w_3296 , w_3297 , w_3298 , w_3299 , w_3300 , w_3301 , w_3302 , w_3303 , w_3304 , w_3305 , 
		w_3306 , w_3307 , w_3308 , w_3309 , w_3310 , w_3311 , w_3312 , w_3313 , w_3314 , w_3315 , 
		w_3316 , w_3317 , w_3318 , w_3319 , w_3320 , w_3321 , w_3322 , w_3323 , w_3324 , w_3325 , 
		w_3326 , w_3327 , w_3328 , w_3329 , w_3330 , w_3331 , w_3332 , w_3333 , w_3334 , w_3335 , 
		w_3336 , w_3337 , w_3338 , w_3339 , w_3340 , w_3341 , w_3342 , w_3343 , w_3344 , w_3345 , 
		w_3346 , w_3347 , w_3348 , w_3349 , w_3350 , w_3351 , w_3352 , w_3353 , w_3354 , w_3355 , 
		w_3356 , w_3357 , w_3358 , w_3359 , w_3360 , w_3361 , w_3362 , w_3363 , w_3364 , w_3365 , 
		w_3366 , w_3367 , w_3368 , w_3369 , w_3370 , w_3371 , w_3372 , w_3373 , w_3374 , w_3375 , 
		w_3376 , w_3377 , w_3378 , w_3379 , w_3380 , w_3381 , w_3382 , w_3383 , w_3384 , w_3385 , 
		w_3386 , w_3387 , w_3388 , w_3389 , w_3390 , w_3391 , w_3392 , w_3393 , w_3394 , w_3395 , 
		w_3396 , w_3397 , w_3398 , w_3399 , w_3400 , w_3401 , w_3402 , w_3403 , w_3404 , w_3405 , 
		w_3406 , w_3407 , w_3408 , w_3409 , w_3410 , w_3411 , w_3412 , w_3413 , w_3414 , w_3415 , 
		w_3416 , w_3417 , w_3418 , w_3419 , w_3420 , w_3421 , w_3422 , w_3423 , w_3424 , w_3425 , 
		w_3426 , w_3427 , w_3428 , w_3429 , w_3430 , w_3431 , w_3432 , w_3433 , w_3434 , w_3435 , 
		w_3436 , w_3437 , w_3438 , w_3439 , w_3440 , w_3441 , w_3442 , w_3443 , w_3444 , w_3445 , 
		w_3446 , w_3447 , w_3448 , w_3449 , w_3450 , w_3451 , w_3452 , w_3453 , w_3454 , w_3455 , 
		w_3456 , w_3457 , w_3458 , w_3459 , w_3460 , w_3461 , w_3462 , w_3463 , w_3464 , w_3465 , 
		w_3466 , w_3467 , w_3468 , w_3469 , w_3470 , w_3471 , w_3472 , w_3473 , w_3474 , w_3475 , 
		w_3476 , w_3477 , w_3478 , w_3479 , w_3480 , w_3481 , w_3482 , w_3483 , w_3484 , w_3485 , 
		w_3486 , w_3487 , w_3488 , w_3489 , w_3490 , w_3491 , w_3492 , w_3493 , w_3494 , w_3495 , 
		w_3496 , w_3497 , w_3498 , w_3499 , w_3500 , w_3501 , w_3502 , w_3503 , w_3504 , w_3505 , 
		w_3506 , w_3507 , w_3508 , w_3509 , w_3510 , w_3511 , w_3512 , w_3513 , w_3514 , w_3515 , 
		w_3516 , w_3517 , w_3518 , w_3519 , w_3520 , w_3521 , w_3522 , w_3523 , w_3524 , w_3525 , 
		w_3526 , w_3527 , w_3528 , w_3529 , w_3530 , w_3531 , w_3532 , w_3533 , w_3534 , w_3535 , 
		w_3536 , w_3537 , w_3538 , w_3539 , w_3540 , w_3541 , w_3542 , w_3543 , w_3544 , w_3545 , 
		w_3546 , w_3547 , w_3548 , w_3549 , w_3550 , w_3551 , w_3552 , w_3553 , w_3554 , w_3555 , 
		w_3556 , w_3557 , w_3558 , w_3559 , w_3560 , w_3561 , w_3562 , w_3563 , w_3564 , w_3565 , 
		w_3566 , w_3567 , w_3568 , w_3569 , w_3570 , w_3571 , w_3572 , w_3573 , w_3574 , w_3575 , 
		w_3576 , w_3577 , w_3578 , w_3579 , w_3580 , w_3581 , w_3582 , w_3583 , w_3584 , w_3585 , 
		w_3586 , w_3587 , w_3588 , w_3589 , w_3590 , w_3591 , w_3592 , w_3593 , w_3594 , w_3595 , 
		w_3596 , w_3597 , w_3598 , w_3599 , w_3600 , w_3601 , w_3602 , w_3603 , w_3604 , w_3605 , 
		w_3606 , w_3607 , w_3608 , w_3609 , w_3610 , w_3611 , w_3612 , w_3613 , w_3614 , w_3615 , 
		w_3616 , w_3617 , w_3618 , w_3619 , w_3620 , w_3621 , w_3622 , w_3623 , w_3624 , w_3625 , 
		w_3626 , w_3627 , w_3628 , w_3629 , w_3630 , w_3631 , w_3632 , w_3633 , w_3634 , w_3635 , 
		w_3636 , w_3637 , w_3638 , w_3639 , w_3640 , w_3641 , w_3642 , w_3643 , w_3644 , w_3645 , 
		w_3646 , w_3647 , w_3648 , w_3649 , w_3650 , w_3651 , w_3652 , w_3653 , w_3654 , w_3655 , 
		w_3656 , w_3657 , w_3658 , w_3659 , w_3660 , w_3661 , w_3662 , w_3663 , w_3664 , w_3665 , 
		w_3666 , w_3667 , w_3668 , w_3669 , w_3670 , w_3671 , w_3672 , w_3673 , w_3674 , w_3675 , 
		w_3676 , w_3677 , w_3678 , w_3679 , w_3680 , w_3681 , w_3682 , w_3683 , w_3684 , w_3685 , 
		w_3686 , w_3687 , w_3688 , w_3689 , w_3690 , w_3691 , w_3692 , w_3693 , w_3694 , w_3695 , 
		w_3696 , w_3697 , w_3698 , w_3699 , w_3700 , w_3701 , w_3702 , w_3703 , w_3704 , w_3705 , 
		w_3706 , w_3707 , w_3708 , w_3709 , w_3710 , w_3711 , w_3712 , w_3713 , w_3714 , w_3715 , 
		w_3716 , w_3717 , w_3718 , w_3719 , w_3720 , w_3721 , w_3722 , w_3723 , w_3724 , w_3725 , 
		w_3726 , w_3727 , w_3728 , w_3729 , w_3730 , w_3731 , w_3732 , w_3733 , w_3734 , w_3735 , 
		w_3736 , w_3737 , w_3738 , w_3739 , w_3740 , w_3741 , w_3742 , w_3743 , w_3744 , w_3745 , 
		w_3746 , w_3747 , w_3748 , w_3749 , w_3750 , w_3751 , w_3752 , w_3753 , w_3754 , w_3755 , 
		w_3756 , w_3757 , w_3758 , w_3759 , w_3760 , w_3761 , w_3762 , w_3763 , w_3764 , w_3765 , 
		w_3766 , w_3767 , w_3768 , w_3769 , w_3770 , w_3771 , w_3772 , w_3773 , w_3774 , w_3775 , 
		w_3776 , w_3777 , w_3778 , w_3779 , w_3780 , w_3781 , w_3782 , w_3783 , w_3784 , w_3785 , 
		w_3786 , w_3787 , w_3788 , w_3789 , w_3790 , w_3791 , w_3792 , w_3793 , w_3794 , w_3795 , 
		w_3796 , w_3797 , w_3798 , w_3799 , w_3800 , w_3801 , w_3802 , w_3803 , w_3804 , w_3805 , 
		w_3806 , w_3807 , w_3808 , w_3809 , w_3810 , w_3811 , w_3812 , w_3813 , w_3814 , w_3815 , 
		w_3816 , w_3817 , w_3818 , w_3819 , w_3820 , w_3821 , w_3822 , w_3823 , w_3824 , w_3825 , 
		w_3826 , w_3827 , w_3828 , w_3829 , w_3830 , w_3831 , w_3832 , w_3833 , w_3834 , w_3835 , 
		w_3836 , w_3837 , w_3838 , w_3839 , w_3840 , w_3841 , w_3842 , w_3843 , w_3844 , w_3845 , 
		w_3846 , w_3847 , w_3848 , w_3849 , w_3850 , w_3851 , w_3852 , w_3853 , w_3854 , w_3855 , 
		w_3856 , w_3857 , w_3858 , w_3859 , w_3860 , w_3861 , w_3862 , w_3863 , w_3864 , w_3865 , 
		w_3866 , w_3867 , w_3868 , w_3869 , w_3870 , w_3871 , w_3872 , w_3873 , w_3874 , w_3875 , 
		w_3876 , w_3877 , w_3878 , w_3879 , w_3880 , w_3881 , w_3882 , w_3883 , w_3884 , w_3885 , 
		w_3886 , w_3887 , w_3888 , w_3889 , w_3890 , w_3891 , w_3892 , w_3893 , w_3894 , w_3895 , 
		w_3896 , w_3897 , w_3898 , w_3899 , w_3900 , w_3901 , w_3902 , w_3903 , w_3904 , w_3905 , 
		w_3906 , w_3907 , w_3908 , w_3909 , w_3910 , w_3911 , w_3912 , w_3913 , w_3914 , w_3915 , 
		w_3916 , w_3917 , w_3918 , w_3919 , w_3920 , w_3921 , w_3922 , w_3923 , w_3924 , w_3925 , 
		w_3926 , w_3927 , w_3928 , w_3929 , w_3930 , w_3931 , w_3932 , w_3933 , w_3934 , w_3935 , 
		w_3936 , w_3937 , w_3938 , w_3939 , w_3940 , w_3941 , w_3942 , w_3943 , w_3944 , w_3945 , 
		w_3946 , w_3947 , w_3948 , w_3949 , w_3950 , w_3951 , w_3952 , w_3953 , w_3954 , w_3955 , 
		w_3956 , w_3957 , w_3958 , w_3959 , w_3960 , w_3961 , w_3962 , w_3963 , w_3964 , w_3965 , 
		w_3966 , w_3967 , w_3968 , w_3969 , w_3970 , w_3971 , w_3972 , w_3973 , w_3974 , w_3975 , 
		w_3976 , w_3977 , w_3978 , w_3979 , w_3980 , w_3981 , w_3982 , w_3983 , w_3984 , w_3985 , 
		w_3986 , w_3987 , w_3988 , w_3989 , w_3990 , w_3991 , w_3992 , w_3993 , w_3994 , w_3995 , 
		w_3996 , w_3997 , w_3998 , w_3999 , w_4000 , w_4001 , w_4002 , w_4003 , w_4004 , w_4005 , 
		w_4006 , w_4007 , w_4008 , w_4009 , w_4010 , w_4011 , w_4012 , w_4013 , w_4014 , w_4015 , 
		w_4016 , w_4017 , w_4018 , w_4019 , w_4020 , w_4021 , w_4022 , w_4023 , w_4024 , w_4025 , 
		w_4026 , w_4027 , w_4028 , w_4029 , w_4030 , w_4031 , w_4032 , w_4033 , w_4034 , w_4035 , 
		w_4036 , w_4037 , w_4038 , w_4039 , w_4040 , w_4041 , w_4042 , w_4043 , w_4044 , w_4045 , 
		w_4046 , w_4047 , w_4048 , w_4049 , w_4050 , w_4051 , w_4052 , w_4053 , w_4054 , w_4055 , 
		w_4056 , w_4057 , w_4058 , w_4059 , w_4060 , w_4061 , w_4062 , w_4063 , w_4064 , w_4065 , 
		w_4066 , w_4067 , w_4068 , w_4069 , w_4070 , w_4071 , w_4072 , w_4073 , w_4074 , w_4075 , 
		w_4076 , w_4077 , w_4078 , w_4079 , w_4080 , w_4081 , w_4082 , w_4083 , w_4084 , w_4085 , 
		w_4086 , w_4087 , w_4088 , w_4089 , w_4090 , w_4091 , w_4092 , w_4093 , w_4094 , w_4095 , 
		w_4096 , w_4097 , w_4098 , w_4099 , w_4100 , w_4101 , w_4102 , w_4103 , w_4104 , w_4105 , 
		w_4106 , w_4107 , w_4108 , w_4109 , w_4110 , w_4111 , w_4112 , w_4113 , w_4114 , w_4115 , 
		w_4116 , w_4117 , w_4118 , w_4119 , w_4120 , w_4121 , w_4122 , w_4123 , w_4124 , w_4125 , 
		w_4126 , w_4127 , w_4128 , w_4129 , w_4130 , w_4131 , w_4132 , w_4133 , w_4134 , w_4135 , 
		w_4136 , w_4137 , w_4138 , w_4139 , w_4140 , w_4141 , w_4142 , w_4143 , w_4144 , w_4145 , 
		w_4146 , w_4147 , w_4148 , w_4149 , w_4150 , w_4151 , w_4152 , w_4153 , w_4154 , w_4155 , 
		w_4156 , w_4157 , w_4158 , w_4159 , w_4160 , w_4161 , w_4162 , w_4163 , w_4164 , w_4165 , 
		w_4166 , w_4167 , w_4168 , w_4169 , w_4170 , w_4171 , w_4172 , w_4173 , w_4174 , w_4175 , 
		w_4176 , w_4177 , w_4178 , w_4179 , w_4180 , w_4181 , w_4182 , w_4183 , w_4184 , w_4185 , 
		w_4186 , w_4187 , w_4188 , w_4189 , w_4190 , w_4191 , w_4192 , w_4193 , w_4194 , w_4195 , 
		w_4196 , w_4197 , w_4198 , w_4199 , w_4200 , w_4201 , w_4202 , w_4203 , w_4204 , w_4205 , 
		w_4206 , w_4207 , w_4208 , w_4209 , w_4210 , w_4211 , w_4212 , w_4213 , w_4214 , w_4215 , 
		w_4216 , w_4217 , w_4218 , w_4219 , w_4220 , w_4221 , w_4222 , w_4223 , w_4224 , w_4225 , 
		w_4226 , w_4227 , w_4228 , w_4229 , w_4230 , w_4231 , w_4232 , w_4233 , w_4234 , w_4235 , 
		w_4236 , w_4237 , w_4238 , w_4239 , w_4240 , w_4241 , w_4242 , w_4243 , w_4244 , w_4245 , 
		w_4246 , w_4247 , w_4248 , w_4249 , w_4250 , w_4251 , w_4252 , w_4253 , w_4254 , w_4255 , 
		w_4256 , w_4257 , w_4258 , w_4259 , w_4260 , w_4261 , w_4262 , w_4263 , w_4264 , w_4265 , 
		w_4266 , w_4267 , w_4268 , w_4269 , w_4270 , w_4271 , w_4272 , w_4273 , w_4274 , w_4275 , 
		w_4276 , w_4277 , w_4278 , w_4279 , w_4280 , w_4281 , w_4282 , w_4283 , w_4284 , w_4285 , 
		w_4286 , w_4287 , w_4288 , w_4289 , w_4290 , w_4291 , w_4292 , w_4293 , w_4294 , w_4295 , 
		w_4296 , w_4297 , w_4298 , w_4299 , w_4300 , w_4301 , w_4302 , w_4303 , w_4304 , w_4305 , 
		w_4306 , w_4307 , w_4308 , w_4309 , w_4310 , w_4311 , w_4312 , w_4313 , w_4314 , w_4315 , 
		w_4316 , w_4317 , w_4318 , w_4319 , w_4320 , w_4321 , w_4322 , w_4323 , w_4324 , w_4325 , 
		w_4326 , w_4327 , w_4328 , w_4329 , w_4330 , w_4331 , w_4332 , w_4333 , w_4334 , w_4335 , 
		w_4336 , w_4337 , w_4338 , w_4339 , w_4340 , w_4341 , w_4342 , w_4343 , w_4344 , w_4345 , 
		w_4346 , w_4347 , w_4348 , w_4349 , w_4350 , w_4351 , w_4352 , w_4353 , w_4354 , w_4355 , 
		w_4356 , w_4357 , w_4358 , w_4359 , w_4360 , w_4361 , w_4362 , w_4363 , w_4364 , w_4365 , 
		w_4366 , w_4367 , w_4368 , w_4369 , w_4370 , w_4371 , w_4372 , w_4373 , w_4374 , w_4375 , 
		w_4376 , w_4377 , w_4378 , w_4379 , w_4380 , w_4381 , w_4382 , w_4383 , w_4384 , w_4385 , 
		w_4386 , w_4387 , w_4388 , w_4389 , w_4390 , w_4391 , w_4392 , w_4393 , w_4394 , w_4395 , 
		w_4396 , w_4397 , w_4398 , w_4399 , w_4400 , w_4401 , w_4402 , w_4403 , w_4404 , w_4405 , 
		w_4406 , w_4407 , w_4408 , w_4409 , w_4410 , w_4411 , w_4412 , w_4413 , w_4414 , w_4415 , 
		w_4416 , w_4417 , w_4418 , w_4419 , w_4420 , w_4421 , w_4422 , w_4423 , w_4424 , w_4425 , 
		w_4426 , w_4427 , w_4428 , w_4429 , w_4430 , w_4431 , w_4432 , w_4433 , w_4434 , w_4435 , 
		w_4436 , w_4437 , w_4438 , w_4439 , w_4440 , w_4441 , w_4442 , w_4443 , w_4444 , w_4445 , 
		w_4446 , w_4447 , w_4448 , w_4449 , w_4450 , w_4451 , w_4452 , w_4453 , w_4454 , w_4455 , 
		w_4456 , w_4457 , w_4458 , w_4459 , w_4460 , w_4461 , w_4462 , w_4463 , w_4464 , w_4465 , 
		w_4466 , w_4467 , w_4468 , w_4469 , w_4470 , w_4471 , w_4472 , w_4473 , w_4474 , w_4475 , 
		w_4476 , w_4477 , w_4478 , w_4479 , w_4480 , w_4481 , w_4482 , w_4483 , w_4484 , w_4485 , 
		w_4486 , w_4487 , w_4488 , w_4489 , w_4490 , w_4491 , w_4492 , w_4493 , w_4494 , w_4495 , 
		w_4496 , w_4497 , w_4498 , w_4499 , w_4500 , w_4501 , w_4502 , w_4503 , w_4504 , w_4505 , 
		w_4506 , w_4507 , w_4508 , w_4509 , w_4510 , w_4511 , w_4512 , w_4513 , w_4514 , w_4515 , 
		w_4516 , w_4517 , w_4518 , w_4519 , w_4520 , w_4521 , w_4522 , w_4523 , w_4524 , w_4525 , 
		w_4526 , w_4527 , w_4528 , w_4529 , w_4530 , w_4531 , w_4532 , w_4533 , w_4534 , w_4535 , 
		w_4536 , w_4537 , w_4538 , w_4539 , w_4540 , w_4541 , w_4542 , w_4543 , w_4544 , w_4545 , 
		w_4546 , w_4547 , w_4548 , w_4549 , w_4550 , w_4551 , w_4552 , w_4553 , w_4554 , w_4555 , 
		w_4556 , w_4557 , w_4558 , w_4559 , w_4560 , w_4561 , w_4562 , w_4563 , w_4564 , w_4565 , 
		w_4566 , w_4567 , w_4568 , w_4569 , w_4570 , w_4571 , w_4572 , w_4573 , w_4574 , w_4575 , 
		w_4576 , w_4577 , w_4578 , w_4579 , w_4580 , w_4581 , w_4582 , w_4583 , w_4584 , w_4585 , 
		w_4586 , w_4587 , w_4588 , w_4589 , w_4590 , w_4591 , w_4592 , w_4593 , w_4594 , w_4595 , 
		w_4596 , w_4597 , w_4598 , w_4599 , w_4600 , w_4601 , w_4602 , w_4603 , w_4604 , w_4605 , 
		w_4606 , w_4607 , w_4608 , w_4609 , w_4610 , w_4611 , w_4612 , w_4613 , w_4614 , w_4615 , 
		w_4616 , w_4617 , w_4618 , w_4619 , w_4620 , w_4621 , w_4622 , w_4623 , w_4624 , w_4625 , 
		w_4626 , w_4627 , w_4628 , w_4629 , w_4630 , w_4631 , w_4632 , w_4633 , w_4634 , w_4635 , 
		w_4636 , w_4637 , w_4638 , w_4639 , w_4640 , w_4641 , w_4642 , w_4643 , w_4644 , w_4645 , 
		w_4646 , w_4647 , w_4648 , w_4649 , w_4650 , w_4651 , w_4652 , w_4653 , w_4654 , w_4655 , 
		w_4656 , w_4657 , w_4658 , w_4659 , w_4660 , w_4661 , w_4662 , w_4663 , w_4664 , w_4665 , 
		w_4666 , w_4667 , w_4668 , w_4669 , w_4670 , w_4671 , w_4672 , w_4673 , w_4674 , w_4675 , 
		w_4676 , w_4677 , w_4678 , w_4679 , w_4680 , w_4681 , w_4682 , w_4683 , w_4684 , w_4685 , 
		w_4686 , w_4687 , w_4688 , w_4689 , w_4690 , w_4691 , w_4692 , w_4693 , w_4694 , w_4695 , 
		w_4696 , w_4697 , w_4698 , w_4699 , w_4700 , w_4701 , w_4702 , w_4703 , w_4704 , w_4705 , 
		w_4706 , w_4707 , w_4708 , w_4709 , w_4710 , w_4711 , w_4712 , w_4713 , w_4714 , w_4715 , 
		w_4716 , w_4717 , w_4718 , w_4719 , w_4720 , w_4721 , w_4722 , w_4723 , w_4724 , w_4725 , 
		w_4726 , w_4727 , w_4728 , w_4729 , w_4730 , w_4731 , w_4732 , w_4733 , w_4734 , w_4735 , 
		w_4736 , w_4737 , w_4738 , w_4739 , w_4740 , w_4741 , w_4742 , w_4743 , w_4744 , w_4745 , 
		w_4746 , w_4747 , w_4748 , w_4749 , w_4750 , w_4751 , w_4752 , w_4753 , w_4754 , w_4755 , 
		w_4756 , w_4757 , w_4758 , w_4759 , w_4760 , w_4761 , w_4762 , w_4763 , w_4764 , w_4765 , 
		w_4766 , w_4767 , w_4768 , w_4769 , w_4770 , w_4771 , w_4772 , w_4773 , w_4774 , w_4775 , 
		w_4776 , w_4777 , w_4778 , w_4779 , w_4780 , w_4781 , w_4782 , w_4783 , w_4784 , w_4785 , 
		w_4786 , w_4787 , w_4788 , w_4789 , w_4790 , w_4791 , w_4792 , w_4793 , w_4794 , w_4795 , 
		w_4796 , w_4797 , w_4798 , w_4799 , w_4800 , w_4801 , w_4802 , w_4803 , w_4804 , w_4805 , 
		w_4806 , w_4807 , w_4808 , w_4809 , w_4810 , w_4811 , w_4812 , w_4813 , w_4814 , w_4815 , 
		w_4816 , w_4817 , w_4818 , w_4819 , w_4820 , w_4821 , w_4822 , w_4823 , w_4824 , w_4825 , 
		w_4826 , w_4827 , w_4828 , w_4829 , w_4830 , w_4831 , w_4832 , w_4833 , w_4834 , w_4835 , 
		w_4836 , w_4837 , w_4838 , w_4839 , w_4840 , w_4841 , w_4842 , w_4843 , w_4844 , w_4845 , 
		w_4846 , w_4847 , w_4848 , w_4849 , w_4850 , w_4851 , w_4852 , w_4853 , w_4854 , w_4855 , 
		w_4856 , w_4857 , w_4858 , w_4859 , w_4860 , w_4861 , w_4862 , w_4863 , w_4864 , w_4865 , 
		w_4866 , w_4867 , w_4868 , w_4869 , w_4870 , w_4871 , w_4872 , w_4873 , w_4874 , w_4875 , 
		w_4876 , w_4877 , w_4878 , w_4879 , w_4880 , w_4881 , w_4882 , w_4883 , w_4884 , w_4885 , 
		w_4886 , w_4887 , w_4888 , w_4889 , w_4890 , w_4891 , w_4892 , w_4893 , w_4894 , w_4895 , 
		w_4896 , w_4897 , w_4898 , w_4899 , w_4900 , w_4901 , w_4902 , w_4903 , w_4904 , w_4905 , 
		w_4906 , w_4907 , w_4908 , w_4909 , w_4910 , w_4911 , w_4912 , w_4913 , w_4914 , w_4915 , 
		w_4916 , w_4917 , w_4918 , w_4919 , w_4920 , w_4921 , w_4922 , w_4923 , w_4924 , w_4925 , 
		w_4926 , w_4927 , w_4928 , w_4929 , w_4930 , w_4931 , w_4932 , w_4933 , w_4934 , w_4935 , 
		w_4936 , w_4937 , w_4938 , w_4939 , w_4940 , w_4941 , w_4942 , w_4943 , w_4944 , w_4945 , 
		w_4946 , w_4947 , w_4948 , w_4949 , w_4950 , w_4951 , w_4952 , w_4953 , w_4954 , w_4955 , 
		w_4956 , w_4957 , w_4958 , w_4959 , w_4960 , w_4961 , w_4962 , w_4963 , w_4964 , w_4965 , 
		w_4966 , w_4967 , w_4968 , w_4969 , w_4970 , w_4971 , w_4972 , w_4973 , w_4974 , w_4975 , 
		w_4976 , w_4977 , w_4978 , w_4979 , w_4980 , w_4981 , w_4982 , w_4983 , w_4984 , w_4985 , 
		w_4986 , w_4987 , w_4988 , w_4989 , w_4990 , w_4991 , w_4992 , w_4993 , w_4994 , w_4995 , 
		w_4996 , w_4997 , w_4998 , w_4999 , w_5000 , w_5001 , w_5002 , w_5003 , w_5004 , w_5005 , 
		w_5006 , w_5007 , w_5008 , w_5009 , w_5010 , w_5011 , w_5012 , w_5013 , w_5014 , w_5015 , 
		w_5016 , w_5017 , w_5018 , w_5019 , w_5020 , w_5021 , w_5022 , w_5023 , w_5024 , w_5025 , 
		w_5026 , w_5027 , w_5028 , w_5029 , w_5030 , w_5031 , w_5032 , w_5033 , w_5034 , w_5035 , 
		w_5036 , w_5037 , w_5038 , w_5039 , w_5040 , w_5041 , w_5042 , w_5043 , w_5044 , w_5045 , 
		w_5046 , w_5047 , w_5048 , w_5049 , w_5050 , w_5051 , w_5052 , w_5053 , w_5054 , w_5055 , 
		w_5056 , w_5057 , w_5058 , w_5059 , w_5060 , w_5061 , w_5062 , w_5063 , w_5064 , w_5065 , 
		w_5066 , w_5067 , w_5068 , w_5069 , w_5070 , w_5071 , w_5072 , w_5073 , w_5074 , w_5075 , 
		w_5076 , w_5077 , w_5078 , w_5079 , w_5080 , w_5081 , w_5082 , w_5083 , w_5084 , w_5085 , 
		w_5086 , w_5087 , w_5088 , w_5089 , w_5090 , w_5091 , w_5092 , w_5093 , w_5094 , w_5095 , 
		w_5096 , w_5097 , w_5098 , w_5099 , w_5100 , w_5101 , w_5102 , w_5103 , w_5104 , w_5105 , 
		w_5106 , w_5107 , w_5108 , w_5109 , w_5110 , w_5111 , w_5112 , w_5113 , w_5114 , w_5115 , 
		w_5116 , w_5117 , w_5118 , w_5119 , w_5120 , w_5121 , w_5122 , w_5123 , w_5124 , w_5125 , 
		w_5126 , w_5127 , w_5128 , w_5129 , w_5130 , w_5131 , w_5132 , w_5133 , w_5134 , w_5135 , 
		w_5136 , w_5137 , w_5138 , w_5139 , w_5140 , w_5141 , w_5142 , w_5143 , w_5144 , w_5145 , 
		w_5146 , w_5147 , w_5148 , w_5149 , w_5150 , w_5151 , w_5152 , w_5153 , w_5154 , w_5155 , 
		w_5156 , w_5157 , w_5158 , w_5159 , w_5160 , w_5161 , w_5162 , w_5163 , w_5164 , w_5165 , 
		w_5166 , w_5167 , w_5168 , w_5169 , w_5170 , w_5171 , w_5172 , w_5173 , w_5174 , w_5175 , 
		w_5176 , w_5177 , w_5178 , w_5179 , w_5180 , w_5181 , w_5182 , w_5183 , w_5184 , w_5185 , 
		w_5186 , w_5187 , w_5188 , w_5189 , w_5190 , w_5191 , w_5192 , w_5193 , w_5194 , w_5195 , 
		w_5196 , w_5197 , w_5198 , w_5199 , w_5200 , w_5201 , w_5202 , w_5203 , w_5204 , w_5205 , 
		w_5206 , w_5207 , w_5208 , w_5209 , w_5210 , w_5211 , w_5212 , w_5213 , w_5214 , w_5215 , 
		w_5216 , w_5217 , w_5218 , w_5219 , w_5220 , w_5221 , w_5222 , w_5223 , w_5224 , w_5225 , 
		w_5226 , w_5227 , w_5228 , w_5229 , w_5230 , w_5231 , w_5232 , w_5233 , w_5234 , w_5235 , 
		w_5236 , w_5237 , w_5238 , w_5239 , w_5240 , w_5241 , w_5242 , w_5243 , w_5244 , w_5245 , 
		w_5246 , w_5247 , w_5248 , w_5249 , w_5250 , w_5251 , w_5252 , w_5253 , w_5254 , w_5255 , 
		w_5256 , w_5257 , w_5258 , w_5259 , w_5260 , w_5261 , w_5262 , w_5263 , w_5264 , w_5265 , 
		w_5266 , w_5267 , w_5268 , w_5269 , w_5270 , w_5271 , w_5272 , w_5273 , w_5274 , w_5275 , 
		w_5276 , w_5277 , w_5278 , w_5279 , w_5280 , w_5281 , w_5282 , w_5283 , w_5284 , w_5285 , 
		w_5286 , w_5287 , w_5288 , w_5289 , w_5290 , w_5291 , w_5292 , w_5293 , w_5294 , w_5295 , 
		w_5296 , w_5297 , w_5298 , w_5299 , w_5300 , w_5301 , w_5302 , w_5303 , w_5304 , w_5305 , 
		w_5306 , w_5307 , w_5308 , w_5309 , w_5310 , w_5311 , w_5312 , w_5313 , w_5314 , w_5315 , 
		w_5316 , w_5317 , w_5318 , w_5319 , w_5320 , w_5321 , w_5322 , w_5323 , w_5324 , w_5325 , 
		w_5326 , w_5327 , w_5328 , w_5329 , w_5330 , w_5331 , w_5332 , w_5333 , w_5334 , w_5335 , 
		w_5336 , w_5337 , w_5338 , w_5339 , w_5340 , w_5341 , w_5342 , w_5343 , w_5344 , w_5345 , 
		w_5346 , w_5347 , w_5348 , w_5349 , w_5350 , w_5351 , w_5352 , w_5353 , w_5354 , w_5355 , 
		w_5356 , w_5357 , w_5358 , w_5359 , w_5360 , w_5361 , w_5362 , w_5363 , w_5364 , w_5365 , 
		w_5366 , w_5367 , w_5368 , w_5369 , w_5370 , w_5371 , w_5372 , w_5373 , w_5374 , w_5375 , 
		w_5376 , w_5377 , w_5378 , w_5379 , w_5380 , w_5381 , w_5382 , w_5383 , w_5384 , w_5385 , 
		w_5386 , w_5387 , w_5388 , w_5389 , w_5390 , w_5391 , w_5392 , w_5393 , w_5394 , w_5395 , 
		w_5396 , w_5397 , w_5398 , w_5399 , w_5400 , w_5401 , w_5402 , w_5403 , w_5404 , w_5405 , 
		w_5406 , w_5407 , w_5408 , w_5409 , w_5410 , w_5411 , w_5412 , w_5413 , w_5414 , w_5415 , 
		w_5416 , w_5417 , w_5418 , w_5419 , w_5420 , w_5421 , w_5422 , w_5423 , w_5424 , w_5425 , 
		w_5426 , w_5427 , w_5428 , w_5429 , w_5430 , w_5431 , w_5432 , w_5433 , w_5434 , w_5435 , 
		w_5436 , w_5437 , w_5438 , w_5439 , w_5440 , w_5441 , w_5442 , w_5443 , w_5444 , w_5445 , 
		w_5446 , w_5447 , w_5448 , w_5449 , w_5450 , w_5451 , w_5452 , w_5453 , w_5454 , w_5455 , 
		w_5456 , w_5457 , w_5458 , w_5459 , w_5460 , w_5461 , w_5462 , w_5463 , w_5464 , w_5465 , 
		w_5466 , w_5467 , w_5468 , w_5469 , w_5470 , w_5471 , w_5472 , w_5473 , w_5474 , w_5475 , 
		w_5476 , w_5477 , w_5478 , w_5479 , w_5480 , w_5481 , w_5482 , w_5483 , w_5484 , w_5485 , 
		w_5486 , w_5487 , w_5488 , w_5489 , w_5490 , w_5491 , w_5492 , w_5493 , w_5494 , w_5495 , 
		w_5496 , w_5497 , w_5498 , w_5499 , w_5500 , w_5501 , w_5502 , w_5503 , w_5504 , w_5505 , 
		w_5506 , w_5507 , w_5508 , w_5509 , w_5510 , w_5511 , w_5512 , w_5513 , w_5514 , w_5515 , 
		w_5516 , w_5517 , w_5518 , w_5519 , w_5520 , w_5521 , w_5522 , w_5523 , w_5524 , w_5525 , 
		w_5526 , w_5527 , w_5528 , w_5529 , w_5530 , w_5531 , w_5532 , w_5533 , w_5534 , w_5535 , 
		w_5536 , w_5537 , w_5538 , w_5539 , w_5540 , w_5541 , w_5542 , w_5543 , w_5544 , w_5545 , 
		w_5546 , w_5547 , w_5548 , w_5549 , w_5550 , w_5551 , w_5552 , w_5553 , w_5554 , w_5555 , 
		w_5556 , w_5557 , w_5558 , w_5559 , w_5560 , w_5561 , w_5562 , w_5563 , w_5564 , w_5565 , 
		w_5566 , w_5567 , w_5568 , w_5569 , w_5570 , w_5571 , w_5572 , w_5573 , w_5574 , w_5575 , 
		w_5576 , w_5577 , w_5578 , w_5579 , w_5580 , w_5581 , w_5582 , w_5583 , w_5584 , w_5585 , 
		w_5586 , w_5587 , w_5588 , w_5589 , w_5590 , w_5591 , w_5592 , w_5593 , w_5594 , w_5595 , 
		w_5596 , w_5597 , w_5598 , w_5599 , w_5600 , w_5601 , w_5602 , w_5603 , w_5604 , w_5605 , 
		w_5606 , w_5607 , w_5608 , w_5609 , w_5610 , w_5611 , w_5612 , w_5613 , w_5614 , w_5615 , 
		w_5616 , w_5617 , w_5618 , w_5619 , w_5620 , w_5621 , w_5622 , w_5623 , w_5624 , w_5625 , 
		w_5626 , w_5627 , w_5628 , w_5629 , w_5630 , w_5631 , w_5632 , w_5633 , w_5634 , w_5635 , 
		w_5636 , w_5637 , w_5638 , w_5639 , w_5640 , w_5641 , w_5642 , w_5643 , w_5644 , w_5645 , 
		w_5646 , w_5647 , w_5648 , w_5649 , w_5650 , w_5651 , w_5652 , w_5653 , w_5654 , w_5655 , 
		w_5656 , w_5657 , w_5658 , w_5659 , w_5660 , w_5661 , w_5662 , w_5663 , w_5664 , w_5665 , 
		w_5666 , w_5667 , w_5668 , w_5669 , w_5670 , w_5671 , w_5672 , w_5673 , w_5674 , w_5675 , 
		w_5676 , w_5677 , w_5678 , w_5679 , w_5680 , w_5681 , w_5682 , w_5683 , w_5684 , w_5685 , 
		w_5686 , w_5687 , w_5688 , w_5689 , w_5690 , w_5691 , w_5692 , w_5693 , w_5694 , w_5695 , 
		w_5696 , w_5697 , w_5698 , w_5699 , w_5700 , w_5701 , w_5702 , w_5703 , w_5704 , w_5705 , 
		w_5706 , w_5707 , w_5708 , w_5709 , w_5710 , w_5711 , w_5712 , w_5713 , w_5714 , w_5715 , 
		w_5716 , w_5717 , w_5718 , w_5719 , w_5720 , w_5721 , w_5722 , w_5723 , w_5724 , w_5725 , 
		w_5726 , w_5727 , w_5728 , w_5729 , w_5730 , w_5731 , w_5732 , w_5733 , w_5734 , w_5735 , 
		w_5736 , w_5737 , w_5738 , w_5739 , w_5740 , w_5741 , w_5742 , w_5743 , w_5744 , w_5745 , 
		w_5746 , w_5747 , w_5748 , w_5749 , w_5750 , w_5751 , w_5752 , w_5753 , w_5754 , w_5755 , 
		w_5756 , w_5757 , w_5758 , w_5759 , w_5760 , w_5761 , w_5762 , w_5763 , w_5764 , w_5765 , 
		w_5766 , w_5767 , w_5768 , w_5769 , w_5770 , w_5771 , w_5772 , w_5773 , w_5774 , w_5775 , 
		w_5776 , w_5777 , w_5778 , w_5779 , w_5780 , w_5781 , w_5782 , w_5783 , w_5784 , w_5785 , 
		w_5786 , w_5787 , w_5788 , w_5789 , w_5790 , w_5791 , w_5792 , w_5793 , w_5794 , w_5795 , 
		w_5796 , w_5797 , w_5798 , w_5799 , w_5800 , w_5801 , w_5802 , w_5803 , w_5804 , w_5805 , 
		w_5806 , w_5807 , w_5808 , w_5809 , w_5810 , w_5811 , w_5812 , w_5813 , w_5814 , w_5815 , 
		w_5816 , w_5817 , w_5818 , w_5819 , w_5820 , w_5821 , w_5822 , w_5823 , w_5824 , w_5825 , 
		w_5826 , w_5827 , w_5828 , w_5829 , w_5830 , w_5831 , w_5832 , w_5833 , w_5834 , w_5835 , 
		w_5836 , w_5837 , w_5838 , w_5839 , w_5840 , w_5841 , w_5842 , w_5843 , w_5844 , w_5845 , 
		w_5846 , w_5847 , w_5848 , w_5849 , w_5850 , w_5851 , w_5852 , w_5853 , w_5854 , w_5855 , 
		w_5856 , w_5857 , w_5858 , w_5859 , w_5860 , w_5861 , w_5862 , w_5863 , w_5864 , w_5865 , 
		w_5866 , w_5867 , w_5868 , w_5869 , w_5870 , w_5871 , w_5872 , w_5873 , w_5874 , w_5875 , 
		w_5876 , w_5877 , w_5878 , w_5879 , w_5880 , w_5881 , w_5882 , w_5883 , w_5884 , w_5885 , 
		w_5886 , w_5887 , w_5888 , w_5889 , w_5890 , w_5891 , w_5892 , w_5893 , w_5894 , w_5895 , 
		w_5896 , w_5897 , w_5898 , w_5899 , w_5900 , w_5901 , w_5902 , w_5903 , w_5904 , w_5905 , 
		w_5906 , w_5907 , w_5908 , w_5909 , w_5910 , w_5911 , w_5912 , w_5913 , w_5914 , w_5915 , 
		w_5916 , w_5917 , w_5918 , w_5919 , w_5920 , w_5921 , w_5922 , w_5923 , w_5924 , w_5925 , 
		w_5926 , w_5927 , w_5928 , w_5929 , w_5930 , w_5931 , w_5932 , w_5933 , w_5934 , w_5935 , 
		w_5936 , w_5937 , w_5938 , w_5939 , w_5940 , w_5941 , w_5942 , w_5943 , w_5944 , w_5945 , 
		w_5946 , w_5947 , w_5948 , w_5949 , w_5950 , w_5951 , w_5952 , w_5953 , w_5954 , w_5955 , 
		w_5956 , w_5957 , w_5958 , w_5959 , w_5960 , w_5961 , w_5962 , w_5963 , w_5964 , w_5965 , 
		w_5966 , w_5967 , w_5968 , w_5969 , w_5970 , w_5971 , w_5972 , w_5973 , w_5974 , w_5975 , 
		w_5976 , w_5977 , w_5978 , w_5979 , w_5980 , w_5981 , w_5982 , w_5983 , w_5984 , w_5985 , 
		w_5986 , w_5987 , w_5988 , w_5989 , w_5990 , w_5991 , w_5992 , w_5993 , w_5994 , w_5995 , 
		w_5996 , w_5997 , w_5998 , w_5999 , w_6000 , w_6001 , w_6002 , w_6003 , w_6004 , w_6005 , 
		w_6006 , w_6007 , w_6008 , w_6009 , w_6010 , w_6011 , w_6012 , w_6013 , w_6014 , w_6015 , 
		w_6016 , w_6017 , w_6018 , w_6019 , w_6020 , w_6021 , w_6022 , w_6023 , w_6024 , w_6025 , 
		w_6026 , w_6027 , w_6028 , w_6029 , w_6030 , w_6031 , w_6032 , w_6033 , w_6034 , w_6035 , 
		w_6036 , w_6037 , w_6038 , w_6039 , w_6040 , w_6041 , w_6042 , w_6043 , w_6044 , w_6045 , 
		w_6046 , w_6047 , w_6048 , w_6049 , w_6050 , w_6051 , w_6052 , w_6053 , w_6054 , w_6055 , 
		w_6056 , w_6057 , w_6058 , w_6059 , w_6060 , w_6061 , w_6062 , w_6063 , w_6064 , w_6065 , 
		w_6066 , w_6067 , w_6068 , w_6069 , w_6070 , w_6071 , w_6072 , w_6073 , w_6074 , w_6075 , 
		w_6076 , w_6077 , w_6078 , w_6079 , w_6080 , w_6081 , w_6082 , w_6083 , w_6084 , w_6085 , 
		w_6086 , w_6087 , w_6088 , w_6089 , w_6090 , w_6091 , w_6092 , w_6093 , w_6094 , w_6095 , 
		w_6096 , w_6097 , w_6098 , w_6099 , w_6100 , w_6101 , w_6102 , w_6103 , w_6104 , w_6105 , 
		w_6106 , w_6107 , w_6108 , w_6109 , w_6110 , w_6111 , w_6112 , w_6113 , w_6114 , w_6115 , 
		w_6116 , w_6117 , w_6118 , w_6119 , w_6120 , w_6121 , w_6122 , w_6123 , w_6124 , w_6125 , 
		w_6126 , w_6127 , w_6128 , w_6129 , w_6130 , w_6131 , w_6132 , w_6133 , w_6134 , w_6135 , 
		w_6136 , w_6137 , w_6138 , w_6139 , w_6140 , w_6141 , w_6142 , w_6143 , w_6144 , w_6145 , 
		w_6146 , w_6147 , w_6148 , w_6149 , w_6150 , w_6151 , w_6152 , w_6153 , w_6154 , w_6155 , 
		w_6156 , w_6157 , w_6158 , w_6159 , w_6160 , w_6161 , w_6162 , w_6163 , w_6164 , w_6165 , 
		w_6166 , w_6167 , w_6168 , w_6169 , w_6170 , w_6171 , w_6172 , w_6173 , w_6174 , w_6175 , 
		w_6176 , w_6177 , w_6178 , w_6179 , w_6180 , w_6181 , w_6182 , w_6183 , w_6184 , w_6185 , 
		w_6186 , w_6187 , w_6188 , w_6189 , w_6190 , w_6191 , w_6192 , w_6193 , w_6194 , w_6195 , 
		w_6196 , w_6197 , w_6198 , w_6199 , w_6200 , w_6201 , w_6202 , w_6203 , w_6204 , w_6205 , 
		w_6206 , w_6207 , w_6208 , w_6209 , w_6210 , w_6211 , w_6212 , w_6213 , w_6214 , w_6215 , 
		w_6216 , w_6217 , w_6218 , w_6219 , w_6220 , w_6221 , w_6222 , w_6223 , w_6224 , w_6225 , 
		w_6226 , w_6227 , w_6228 , w_6229 , w_6230 , w_6231 , w_6232 , w_6233 , w_6234 , w_6235 , 
		w_6236 , w_6237 , w_6238 , w_6239 , w_6240 , w_6241 , w_6242 , w_6243 , w_6244 , w_6245 , 
		w_6246 , w_6247 , w_6248 , w_6249 , w_6250 , w_6251 , w_6252 , w_6253 , w_6254 , w_6255 , 
		w_6256 , w_6257 , w_6258 , w_6259 , w_6260 , w_6261 , w_6262 , w_6263 , w_6264 , w_6265 , 
		w_6266 , w_6267 , w_6268 , w_6269 , w_6270 , w_6271 , w_6272 , w_6273 , w_6274 , w_6275 , 
		w_6276 , w_6277 , w_6278 , w_6279 , w_6280 , w_6281 , w_6282 , w_6283 , w_6284 , w_6285 , 
		w_6286 , w_6287 , w_6288 , w_6289 , w_6290 , w_6291 , w_6292 , w_6293 , w_6294 , w_6295 , 
		w_6296 , w_6297 , w_6298 , w_6299 , w_6300 , w_6301 , w_6302 , w_6303 , w_6304 , w_6305 , 
		w_6306 , w_6307 , w_6308 , w_6309 , w_6310 , w_6311 , w_6312 , w_6313 , w_6314 , w_6315 , 
		w_6316 , w_6317 , w_6318 , w_6319 , w_6320 , w_6321 , w_6322 , w_6323 , w_6324 , w_6325 , 
		w_6326 , w_6327 , w_6328 , w_6329 , w_6330 , w_6331 , w_6332 , w_6333 , w_6334 , w_6335 , 
		w_6336 , w_6337 , w_6338 , w_6339 , w_6340 , w_6341 , w_6342 , w_6343 , w_6344 , w_6345 , 
		w_6346 , w_6347 , w_6348 , w_6349 , w_6350 , w_6351 , w_6352 , w_6353 , w_6354 , w_6355 , 
		w_6356 , w_6357 , w_6358 , w_6359 , w_6360 , w_6361 , w_6362 , w_6363 , w_6364 , w_6365 , 
		w_6366 , w_6367 , w_6368 , w_6369 , w_6370 , w_6371 , w_6372 , w_6373 , w_6374 , w_6375 , 
		w_6376 , w_6377 , w_6378 , w_6379 , w_6380 , w_6381 , w_6382 , w_6383 , w_6384 , w_6385 , 
		w_6386 , w_6387 , w_6388 , w_6389 , w_6390 , w_6391 , w_6392 , w_6393 , w_6394 , w_6395 , 
		w_6396 , w_6397 , w_6398 , w_6399 , w_6400 , w_6401 , w_6402 , w_6403 , w_6404 , w_6405 , 
		w_6406 , w_6407 , w_6408 , w_6409 , w_6410 , w_6411 , w_6412 , w_6413 , w_6414 , w_6415 , 
		w_6416 , w_6417 , w_6418 , w_6419 , w_6420 , w_6421 , w_6422 , w_6423 , w_6424 , w_6425 , 
		w_6426 , w_6427 , w_6428 , w_6429 , w_6430 , w_6431 , w_6432 , w_6433 , w_6434 , w_6435 , 
		w_6436 , w_6437 , w_6438 , w_6439 , w_6440 , w_6441 , w_6442 , w_6443 , w_6444 , w_6445 , 
		w_6446 , w_6447 , w_6448 , w_6449 , w_6450 , w_6451 , w_6452 , w_6453 , w_6454 , w_6455 , 
		w_6456 , w_6457 , w_6458 , w_6459 , w_6460 , w_6461 , w_6462 , w_6463 , w_6464 , w_6465 , 
		w_6466 , w_6467 , w_6468 , w_6469 , w_6470 , w_6471 , w_6472 , w_6473 , w_6474 , w_6475 , 
		w_6476 , w_6477 , w_6478 , w_6479 , w_6480 , w_6481 , w_6482 , w_6483 , w_6484 , w_6485 , 
		w_6486 , w_6487 , w_6488 , w_6489 , w_6490 , w_6491 , w_6492 , w_6493 , w_6494 , w_6495 , 
		w_6496 , w_6497 , w_6498 , w_6499 , w_6500 , w_6501 , w_6502 , w_6503 , w_6504 , w_6505 , 
		w_6506 , w_6507 , w_6508 , w_6509 , w_6510 , w_6511 , w_6512 , w_6513 , w_6514 , w_6515 , 
		w_6516 , w_6517 , w_6518 , w_6519 , w_6520 , w_6521 , w_6522 , w_6523 , w_6524 , w_6525 , 
		w_6526 , w_6527 , w_6528 , w_6529 , w_6530 , w_6531 , w_6532 , w_6533 , w_6534 , w_6535 , 
		w_6536 , w_6537 , w_6538 , w_6539 , w_6540 , w_6541 , w_6542 , w_6543 , w_6544 , w_6545 , 
		w_6546 , w_6547 , w_6548 , w_6549 , w_6550 , w_6551 , w_6552 , w_6553 , w_6554 , w_6555 , 
		w_6556 , w_6557 , w_6558 , w_6559 , w_6560 , w_6561 , w_6562 , w_6563 , w_6564 , w_6565 , 
		w_6566 , w_6567 , w_6568 , w_6569 , w_6570 , w_6571 , w_6572 , w_6573 , w_6574 , w_6575 , 
		w_6576 , w_6577 , w_6578 , w_6579 , w_6580 , w_6581 , w_6582 , w_6583 , w_6584 , w_6585 , 
		w_6586 , w_6587 , w_6588 , w_6589 , w_6590 , w_6591 , w_6592 , w_6593 , w_6594 , w_6595 , 
		w_6596 , w_6597 , w_6598 , w_6599 , w_6600 , w_6601 , w_6602 , w_6603 , w_6604 , w_6605 , 
		w_6606 , w_6607 , w_6608 , w_6609 , w_6610 , w_6611 , w_6612 , w_6613 , w_6614 , w_6615 , 
		w_6616 , w_6617 , w_6618 , w_6619 , w_6620 , w_6621 , w_6622 , w_6623 , w_6624 , w_6625 , 
		w_6626 , w_6627 , w_6628 , w_6629 , w_6630 , w_6631 , w_6632 , w_6633 , w_6634 , w_6635 , 
		w_6636 , w_6637 , w_6638 , w_6639 , w_6640 , w_6641 , w_6642 , w_6643 , w_6644 , w_6645 , 
		w_6646 , w_6647 , w_6648 , w_6649 , w_6650 , w_6651 , w_6652 , w_6653 , w_6654 , w_6655 , 
		w_6656 , w_6657 , w_6658 , w_6659 , w_6660 , w_6661 , w_6662 , w_6663 , w_6664 , w_6665 , 
		w_6666 , w_6667 , w_6668 , w_6669 , w_6670 , w_6671 , w_6672 , w_6673 , w_6674 , w_6675 , 
		w_6676 , w_6677 , w_6678 , w_6679 , w_6680 , w_6681 , w_6682 , w_6683 , w_6684 , w_6685 , 
		w_6686 , w_6687 , w_6688 , w_6689 , w_6690 , w_6691 , w_6692 , w_6693 , w_6694 , w_6695 , 
		w_6696 , w_6697 , w_6698 , w_6699 , w_6700 , w_6701 , w_6702 , w_6703 , w_6704 , w_6705 , 
		w_6706 , w_6707 , w_6708 , w_6709 , w_6710 , w_6711 , w_6712 , w_6713 , w_6714 , w_6715 , 
		w_6716 , w_6717 , w_6718 , w_6719 , w_6720 , w_6721 , w_6722 , w_6723 , w_6724 , w_6725 , 
		w_6726 , w_6727 , w_6728 , w_6729 , w_6730 , w_6731 , w_6732 , w_6733 , w_6734 , w_6735 , 
		w_6736 , w_6737 , w_6738 , w_6739 , w_6740 , w_6741 , w_6742 , w_6743 , w_6744 , w_6745 , 
		w_6746 , w_6747 , w_6748 , w_6749 , w_6750 , w_6751 , w_6752 , w_6753 , w_6754 , w_6755 , 
		w_6756 , w_6757 , w_6758 , w_6759 , w_6760 , w_6761 , w_6762 , w_6763 , w_6764 , w_6765 , 
		w_6766 , w_6767 , w_6768 , w_6769 , w_6770 , w_6771 , w_6772 , w_6773 , w_6774 , w_6775 , 
		w_6776 , w_6777 , w_6778 , w_6779 , w_6780 , w_6781 , w_6782 , w_6783 , w_6784 , w_6785 , 
		w_6786 , w_6787 , w_6788 , w_6789 , w_6790 , w_6791 , w_6792 , w_6793 , w_6794 , w_6795 , 
		w_6796 , w_6797 , w_6798 , w_6799 , w_6800 , w_6801 , w_6802 , w_6803 , w_6804 , w_6805 , 
		w_6806 , w_6807 , w_6808 , w_6809 , w_6810 , w_6811 , w_6812 , w_6813 , w_6814 , w_6815 , 
		w_6816 , w_6817 , w_6818 , w_6819 , w_6820 , w_6821 , w_6822 , w_6823 , w_6824 , w_6825 , 
		w_6826 , w_6827 , w_6828 , w_6829 , w_6830 , w_6831 , w_6832 , w_6833 , w_6834 , w_6835 , 
		w_6836 , w_6837 , w_6838 , w_6839 , w_6840 , w_6841 , w_6842 , w_6843 , w_6844 , w_6845 , 
		w_6846 , w_6847 , w_6848 , w_6849 , w_6850 , w_6851 , w_6852 , w_6853 , w_6854 , w_6855 , 
		w_6856 , w_6857 , w_6858 , w_6859 , w_6860 , w_6861 , w_6862 , w_6863 , w_6864 , w_6865 , 
		w_6866 , w_6867 , w_6868 , w_6869 , w_6870 , w_6871 , w_6872 , w_6873 , w_6874 , w_6875 , 
		w_6876 , w_6877 , w_6878 , w_6879 , w_6880 , w_6881 , w_6882 , w_6883 , w_6884 , w_6885 , 
		w_6886 , w_6887 , w_6888 , w_6889 , w_6890 , w_6891 , w_6892 , w_6893 , w_6894 , w_6895 , 
		w_6896 , w_6897 , w_6898 , w_6899 , w_6900 , w_6901 , w_6902 , w_6903 , w_6904 , w_6905 , 
		w_6906 , w_6907 , w_6908 , w_6909 , w_6910 , w_6911 , w_6912 , w_6913 , w_6914 , w_6915 , 
		w_6916 , w_6917 , w_6918 , w_6919 , w_6920 , w_6921 , w_6922 , w_6923 , w_6924 , w_6925 , 
		w_6926 , w_6927 , w_6928 , w_6929 , w_6930 , w_6931 , w_6932 , w_6933 , w_6934 , w_6935 , 
		w_6936 , w_6937 , w_6938 , w_6939 , w_6940 , w_6941 , w_6942 , w_6943 , w_6944 , w_6945 , 
		w_6946 , w_6947 , w_6948 , w_6949 , w_6950 , w_6951 , w_6952 , w_6953 , w_6954 , w_6955 , 
		w_6956 , w_6957 , w_6958 , w_6959 , w_6960 , w_6961 , w_6962 , w_6963 , w_6964 , w_6965 , 
		w_6966 , w_6967 , w_6968 , w_6969 , w_6970 , w_6971 , w_6972 , w_6973 , w_6974 , w_6975 , 
		w_6976 , w_6977 , w_6978 , w_6979 , w_6980 , w_6981 , w_6982 , w_6983 , w_6984 , w_6985 , 
		w_6986 , w_6987 , w_6988 , w_6989 , w_6990 , w_6991 , w_6992 , w_6993 , w_6994 , w_6995 , 
		w_6996 , w_6997 , w_6998 , w_6999 , w_7000 , w_7001 , w_7002 , w_7003 , w_7004 , w_7005 , 
		w_7006 , w_7007 , w_7008 , w_7009 , w_7010 , w_7011 , w_7012 , w_7013 , w_7014 , w_7015 , 
		w_7016 , w_7017 , w_7018 , w_7019 , w_7020 , w_7021 , w_7022 , w_7023 , w_7024 , w_7025 , 
		w_7026 , w_7027 , w_7028 , w_7029 , w_7030 , w_7031 , w_7032 , w_7033 , w_7034 , w_7035 , 
		w_7036 , w_7037 , w_7038 , w_7039 , w_7040 , w_7041 , w_7042 , w_7043 , w_7044 , w_7045 , 
		w_7046 , w_7047 , w_7048 , w_7049 , w_7050 , w_7051 , w_7052 , w_7053 , w_7054 , w_7055 , 
		w_7056 , w_7057 , w_7058 , w_7059 , w_7060 , w_7061 , w_7062 , w_7063 , w_7064 , w_7065 , 
		w_7066 , w_7067 , w_7068 , w_7069 , w_7070 , w_7071 , w_7072 , w_7073 , w_7074 , w_7075 , 
		w_7076 , w_7077 , w_7078 , w_7079 , w_7080 , w_7081 , w_7082 , w_7083 , w_7084 , w_7085 , 
		w_7086 , w_7087 , w_7088 , w_7089 , w_7090 , w_7091 , w_7092 , w_7093 , w_7094 , w_7095 , 
		w_7096 , w_7097 , w_7098 , w_7099 , w_7100 , w_7101 , w_7102 , w_7103 , w_7104 , w_7105 , 
		w_7106 , w_7107 , w_7108 , w_7109 , w_7110 , w_7111 , w_7112 , w_7113 , w_7114 , w_7115 , 
		w_7116 , w_7117 , w_7118 , w_7119 , w_7120 , w_7121 , w_7122 , w_7123 , w_7124 , w_7125 , 
		w_7126 , w_7127 , w_7128 , w_7129 , w_7130 , w_7131 , w_7132 , w_7133 , w_7134 , w_7135 , 
		w_7136 , w_7137 , w_7138 , w_7139 , w_7140 , w_7141 , w_7142 , w_7143 , w_7144 , w_7145 , 
		w_7146 , w_7147 , w_7148 , w_7149 , w_7150 , w_7151 , w_7152 , w_7153 , w_7154 , w_7155 , 
		w_7156 , w_7157 , w_7158 , w_7159 , w_7160 , w_7161 , w_7162 , w_7163 , w_7164 , w_7165 , 
		w_7166 , w_7167 , w_7168 , w_7169 , w_7170 , w_7171 , w_7172 , w_7173 , w_7174 , w_7175 , 
		w_7176 , w_7177 , w_7178 , w_7179 , w_7180 , w_7181 , w_7182 , w_7183 , w_7184 , w_7185 , 
		w_7186 , w_7187 , w_7188 , w_7189 , w_7190 , w_7191 , w_7192 , w_7193 , w_7194 , w_7195 , 
		w_7196 , w_7197 , w_7198 , w_7199 , w_7200 , w_7201 , w_7202 , w_7203 , w_7204 , w_7205 , 
		w_7206 , w_7207 , w_7208 , w_7209 , w_7210 , w_7211 , w_7212 , w_7213 , w_7214 , w_7215 , 
		w_7216 , w_7217 , w_7218 , w_7219 , w_7220 , w_7221 , w_7222 , w_7223 , w_7224 , w_7225 , 
		w_7226 , w_7227 , w_7228 , w_7229 , w_7230 , w_7231 , w_7232 , w_7233 , w_7234 , w_7235 , 
		w_7236 , w_7237 , w_7238 , w_7239 , w_7240 , w_7241 , w_7242 , w_7243 , w_7244 , w_7245 , 
		w_7246 , w_7247 , w_7248 , w_7249 , w_7250 , w_7251 , w_7252 , w_7253 , w_7254 , w_7255 , 
		w_7256 , w_7257 , w_7258 , w_7259 , w_7260 , w_7261 , w_7262 , w_7263 , w_7264 , w_7265 , 
		w_7266 , w_7267 , w_7268 , w_7269 , w_7270 , w_7271 , w_7272 , w_7273 , w_7274 , w_7275 , 
		w_7276 , w_7277 , w_7278 , w_7279 , w_7280 , w_7281 , w_7282 , w_7283 , w_7284 , w_7285 , 
		w_7286 , w_7287 , w_7288 , w_7289 , w_7290 , w_7291 , w_7292 , w_7293 , w_7294 , w_7295 , 
		w_7296 , w_7297 , w_7298 , w_7299 , w_7300 , w_7301 , w_7302 , w_7303 , w_7304 , w_7305 , 
		w_7306 , w_7307 , w_7308 , w_7309 , w_7310 , w_7311 , w_7312 , w_7313 , w_7314 , w_7315 , 
		w_7316 , w_7317 , w_7318 , w_7319 , w_7320 , w_7321 , w_7322 , w_7323 , w_7324 , w_7325 , 
		w_7326 , w_7327 , w_7328 , w_7329 , w_7330 , w_7331 , w_7332 , w_7333 , w_7334 , w_7335 , 
		w_7336 , w_7337 , w_7338 , w_7339 , w_7340 , w_7341 , w_7342 , w_7343 , w_7344 , w_7345 , 
		w_7346 , w_7347 , w_7348 , w_7349 , w_7350 , w_7351 , w_7352 , w_7353 , w_7354 , w_7355 , 
		w_7356 , w_7357 , w_7358 , w_7359 , w_7360 , w_7361 , w_7362 , w_7363 , w_7364 , w_7365 , 
		w_7366 , w_7367 , w_7368 , w_7369 , w_7370 , w_7371 , w_7372 , w_7373 , w_7374 , w_7375 , 
		w_7376 , w_7377 , w_7378 , w_7379 , w_7380 , w_7381 , w_7382 , w_7383 , w_7384 , w_7385 , 
		w_7386 , w_7387 , w_7388 , w_7389 , w_7390 , w_7391 , w_7392 , w_7393 , w_7394 , w_7395 , 
		w_7396 , w_7397 , w_7398 , w_7399 , w_7400 , w_7401 , w_7402 , w_7403 , w_7404 , w_7405 , 
		w_7406 , w_7407 , w_7408 , w_7409 , w_7410 , w_7411 , w_7412 , w_7413 , w_7414 , w_7415 , 
		w_7416 , w_7417 , w_7418 , w_7419 , w_7420 , w_7421 , w_7422 , w_7423 , w_7424 , w_7425 , 
		w_7426 , w_7427 , w_7428 , w_7429 , w_7430 , w_7431 , w_7432 , w_7433 , w_7434 , w_7435 , 
		w_7436 , w_7437 , w_7438 , w_7439 , w_7440 , w_7441 , w_7442 , w_7443 , w_7444 , w_7445 , 
		w_7446 , w_7447 , w_7448 , w_7449 , w_7450 , w_7451 , w_7452 , w_7453 , w_7454 , w_7455 , 
		w_7456 , w_7457 , w_7458 , w_7459 , w_7460 , w_7461 , w_7462 , w_7463 , w_7464 , w_7465 , 
		w_7466 , w_7467 , w_7468 , w_7469 , w_7470 , w_7471 , w_7472 , w_7473 , w_7474 , w_7475 , 
		w_7476 , w_7477 , w_7478 , w_7479 , w_7480 , w_7481 , w_7482 , w_7483 , w_7484 , w_7485 , 
		w_7486 , w_7487 , w_7488 , w_7489 , w_7490 , w_7491 , w_7492 , w_7493 , w_7494 , w_7495 , 
		w_7496 , w_7497 , w_7498 , w_7499 , w_7500 , w_7501 , w_7502 , w_7503 , w_7504 , w_7505 , 
		w_7506 , w_7507 , w_7508 , w_7509 , w_7510 , w_7511 , w_7512 , w_7513 , w_7514 , w_7515 , 
		w_7516 , w_7517 , w_7518 , w_7519 , w_7520 , w_7521 , w_7522 , w_7523 , w_7524 , w_7525 , 
		w_7526 , w_7527 , w_7528 , w_7529 , w_7530 , w_7531 , w_7532 , w_7533 , w_7534 , w_7535 , 
		w_7536 , w_7537 , w_7538 , w_7539 , w_7540 , w_7541 , w_7542 , w_7543 , w_7544 , w_7545 , 
		w_7546 , w_7547 , w_7548 , w_7549 , w_7550 , w_7551 , w_7552 , w_7553 , w_7554 , w_7555 , 
		w_7556 , w_7557 , w_7558 , w_7559 , w_7560 , w_7561 , w_7562 , w_7563 , w_7564 , w_7565 , 
		w_7566 , w_7567 , w_7568 , w_7569 , w_7570 , w_7571 , w_7572 , w_7573 , w_7574 , w_7575 , 
		w_7576 , w_7577 , w_7578 , w_7579 , w_7580 , w_7581 , w_7582 , w_7583 , w_7584 , w_7585 , 
		w_7586 , w_7587 , w_7588 , w_7589 , w_7590 , w_7591 , w_7592 , w_7593 , w_7594 , w_7595 , 
		w_7596 , w_7597 , w_7598 , w_7599 , w_7600 , w_7601 , w_7602 , w_7603 , w_7604 , w_7605 , 
		w_7606 , w_7607 , w_7608 , w_7609 , w_7610 , w_7611 , w_7612 , w_7613 , w_7614 , w_7615 , 
		w_7616 , w_7617 , w_7618 , w_7619 , w_7620 , w_7621 , w_7622 , w_7623 , w_7624 , w_7625 , 
		w_7626 , w_7627 , w_7628 , w_7629 , w_7630 , w_7631 , w_7632 , w_7633 , w_7634 , w_7635 , 
		w_7636 , w_7637 , w_7638 , w_7639 , w_7640 , w_7641 , w_7642 , w_7643 , w_7644 , w_7645 , 
		w_7646 , w_7647 , w_7648 , w_7649 , w_7650 , w_7651 , w_7652 , w_7653 , w_7654 , w_7655 , 
		w_7656 , w_7657 , w_7658 , w_7659 , w_7660 , w_7661 , w_7662 , w_7663 , w_7664 , w_7665 , 
		w_7666 , w_7667 , w_7668 , w_7669 , w_7670 , w_7671 , w_7672 , w_7673 , w_7674 , w_7675 , 
		w_7676 , w_7677 , w_7678 , w_7679 , w_7680 , w_7681 , w_7682 , w_7683 , w_7684 , w_7685 , 
		w_7686 , w_7687 , w_7688 , w_7689 , w_7690 , w_7691 , w_7692 , w_7693 , w_7694 , w_7695 , 
		w_7696 , w_7697 , w_7698 , w_7699 , w_7700 , w_7701 , w_7702 , w_7703 , w_7704 , w_7705 , 
		w_7706 , w_7707 , w_7708 , w_7709 , w_7710 , w_7711 , w_7712 , w_7713 , w_7714 , w_7715 , 
		w_7716 , w_7717 , w_7718 , w_7719 , w_7720 , w_7721 , w_7722 , w_7723 , w_7724 , w_7725 , 
		w_7726 , w_7727 , w_7728 , w_7729 , w_7730 , w_7731 , w_7732 , w_7733 , w_7734 , w_7735 , 
		w_7736 , w_7737 , w_7738 , w_7739 , w_7740 , w_7741 , w_7742 , w_7743 , w_7744 , w_7745 , 
		w_7746 , w_7747 , w_7748 , w_7749 , w_7750 , w_7751 , w_7752 , w_7753 , w_7754 , w_7755 , 
		w_7756 , w_7757 , w_7758 , w_7759 , w_7760 , w_7761 , w_7762 , w_7763 , w_7764 , w_7765 , 
		w_7766 , w_7767 , w_7768 , w_7769 , w_7770 , w_7771 , w_7772 , w_7773 , w_7774 , w_7775 , 
		w_7776 , w_7777 , w_7778 , w_7779 , w_7780 , w_7781 , w_7782 , w_7783 , w_7784 , w_7785 , 
		w_7786 , w_7787 , w_7788 , w_7789 , w_7790 , w_7791 , w_7792 , w_7793 , w_7794 , w_7795 , 
		w_7796 , w_7797 , w_7798 , w_7799 , w_7800 , w_7801 , w_7802 , w_7803 , w_7804 , w_7805 , 
		w_7806 , w_7807 , w_7808 , w_7809 , w_7810 , w_7811 , w_7812 , w_7813 , w_7814 , w_7815 , 
		w_7816 , w_7817 , w_7818 , w_7819 , w_7820 , w_7821 , w_7822 , w_7823 , w_7824 , w_7825 , 
		w_7826 , w_7827 , w_7828 , w_7829 , w_7830 , w_7831 , w_7832 , w_7833 , w_7834 , w_7835 , 
		w_7836 , w_7837 , w_7838 , w_7839 , w_7840 , w_7841 , w_7842 , w_7843 , w_7844 , w_7845 , 
		w_7846 , w_7847 , w_7848 , w_7849 , w_7850 , w_7851 , w_7852 , w_7853 , w_7854 , w_7855 , 
		w_7856 , w_7857 , w_7858 , w_7859 , w_7860 , w_7861 , w_7862 , w_7863 , w_7864 , w_7865 , 
		w_7866 , w_7867 , w_7868 , w_7869 , w_7870 , w_7871 , w_7872 , w_7873 , w_7874 , w_7875 , 
		w_7876 , w_7877 , w_7878 , w_7879 , w_7880 , w_7881 , w_7882 , w_7883 , w_7884 , w_7885 , 
		w_7886 , w_7887 , w_7888 , w_7889 , w_7890 , w_7891 , w_7892 , w_7893 , w_7894 , w_7895 , 
		w_7896 , w_7897 , w_7898 , w_7899 , w_7900 , w_7901 , w_7902 , w_7903 , w_7904 , w_7905 , 
		w_7906 , w_7907 , w_7908 , w_7909 , w_7910 , w_7911 , w_7912 , w_7913 , w_7914 , w_7915 , 
		w_7916 , w_7917 , w_7918 , w_7919 , w_7920 , w_7921 , w_7922 , w_7923 , w_7924 , w_7925 , 
		w_7926 , w_7927 , w_7928 , w_7929 , w_7930 , w_7931 , w_7932 , w_7933 , w_7934 , w_7935 , 
		w_7936 , w_7937 , w_7938 , w_7939 , w_7940 , w_7941 , w_7942 , w_7943 , w_7944 , w_7945 , 
		w_7946 , w_7947 , w_7948 , w_7949 , w_7950 , w_7951 , w_7952 , w_7953 , w_7954 , w_7955 , 
		w_7956 , w_7957 , w_7958 , w_7959 , w_7960 , w_7961 , w_7962 , w_7963 , w_7964 , w_7965 , 
		w_7966 , w_7967 , w_7968 , w_7969 , w_7970 , w_7971 , w_7972 , w_7973 , w_7974 , w_7975 , 
		w_7976 , w_7977 , w_7978 , w_7979 , w_7980 , w_7981 , w_7982 , w_7983 , w_7984 , w_7985 , 
		w_7986 , w_7987 , w_7988 , w_7989 , w_7990 , w_7991 , w_7992 , w_7993 , w_7994 , w_7995 , 
		w_7996 , w_7997 , w_7998 , w_7999 , w_8000 , w_8001 , w_8002 , w_8003 , w_8004 , w_8005 , 
		w_8006 , w_8007 , w_8008 , w_8009 , w_8010 , w_8011 , w_8012 , w_8013 , w_8014 , w_8015 , 
		w_8016 , w_8017 , w_8018 , w_8019 , w_8020 , w_8021 , w_8022 , w_8023 , w_8024 , w_8025 , 
		w_8026 , w_8027 , w_8028 , w_8029 , w_8030 , w_8031 , w_8032 , w_8033 , w_8034 , w_8035 , 
		w_8036 , w_8037 , w_8038 , w_8039 , w_8040 , w_8041 , w_8042 , w_8043 , w_8044 , w_8045 , 
		w_8046 , w_8047 , w_8048 , w_8049 , w_8050 , w_8051 , w_8052 , w_8053 , w_8054 , w_8055 , 
		w_8056 , w_8057 , w_8058 , w_8059 , w_8060 , w_8061 , w_8062 , w_8063 , w_8064 , w_8065 , 
		w_8066 , w_8067 , w_8068 , w_8069 , w_8070 , w_8071 , w_8072 , w_8073 , w_8074 , w_8075 , 
		w_8076 , w_8077 , w_8078 , w_8079 , w_8080 , w_8081 , w_8082 , w_8083 , w_8084 , w_8085 , 
		w_8086 , w_8087 , w_8088 , w_8089 , w_8090 , w_8091 , w_8092 , w_8093 , w_8094 , w_8095 , 
		w_8096 , w_8097 , w_8098 , w_8099 , w_8100 , w_8101 , w_8102 , w_8103 , w_8104 , w_8105 , 
		w_8106 , w_8107 , w_8108 , w_8109 , w_8110 , w_8111 , w_8112 , w_8113 , w_8114 , w_8115 , 
		w_8116 , w_8117 , w_8118 , w_8119 , w_8120 , w_8121 , w_8122 , w_8123 , w_8124 , w_8125 , 
		w_8126 , w_8127 , w_8128 , w_8129 , w_8130 , w_8131 , w_8132 , w_8133 , w_8134 , w_8135 , 
		w_8136 , w_8137 , w_8138 , w_8139 , w_8140 , w_8141 , w_8142 , w_8143 , w_8144 , w_8145 , 
		w_8146 , w_8147 , w_8148 , w_8149 , w_8150 , w_8151 , w_8152 , w_8153 , w_8154 , w_8155 , 
		w_8156 , w_8157 , w_8158 , w_8159 , w_8160 , w_8161 , w_8162 , w_8163 , w_8164 , w_8165 , 
		w_8166 , w_8167 , w_8168 , w_8169 , w_8170 , w_8171 , w_8172 , w_8173 , w_8174 , w_8175 , 
		w_8176 , w_8177 , w_8178 , w_8179 , w_8180 , w_8181 , w_8182 , w_8183 , w_8184 , w_8185 , 
		w_8186 , w_8187 , w_8188 , w_8189 , w_8190 , w_8191 , w_8192 , w_8193 , w_8194 , w_8195 , 
		w_8196 , w_8197 , w_8198 , w_8199 , w_8200 , w_8201 , w_8202 , w_8203 , w_8204 , w_8205 , 
		w_8206 , w_8207 , w_8208 , w_8209 , w_8210 , w_8211 , w_8212 , w_8213 , w_8214 , w_8215 , 
		w_8216 , w_8217 , w_8218 , w_8219 , w_8220 , w_8221 , w_8222 , w_8223 , w_8224 , w_8225 , 
		w_8226 , w_8227 , w_8228 , w_8229 , w_8230 , w_8231 , w_8232 , w_8233 , w_8234 , w_8235 , 
		w_8236 , w_8237 , w_8238 , w_8239 , w_8240 , w_8241 , w_8242 , w_8243 , w_8244 , w_8245 , 
		w_8246 , w_8247 , w_8248 , w_8249 , w_8250 , w_8251 , w_8252 , w_8253 , w_8254 , w_8255 , 
		w_8256 , w_8257 , w_8258 , w_8259 , w_8260 , w_8261 , w_8262 , w_8263 , w_8264 , w_8265 , 
		w_8266 , w_8267 , w_8268 , w_8269 , w_8270 , w_8271 , w_8272 , w_8273 , w_8274 , w_8275 , 
		w_8276 , w_8277 , w_8278 , w_8279 , w_8280 , w_8281 , w_8282 , w_8283 , w_8284 , w_8285 , 
		w_8286 , w_8287 , w_8288 , w_8289 , w_8290 , w_8291 , w_8292 , w_8293 , w_8294 , w_8295 , 
		w_8296 , w_8297 , w_8298 , w_8299 , w_8300 , w_8301 , w_8302 , w_8303 , w_8304 , w_8305 , 
		w_8306 , w_8307 , w_8308 , w_8309 , w_8310 , w_8311 , w_8312 , w_8313 , w_8314 , w_8315 , 
		w_8316 , w_8317 , w_8318 , w_8319 , w_8320 , w_8321 , w_8322 , w_8323 , w_8324 , w_8325 , 
		w_8326 , w_8327 , w_8328 , w_8329 , w_8330 , w_8331 , w_8332 , w_8333 , w_8334 , w_8335 , 
		w_8336 , w_8337 , w_8338 , w_8339 , w_8340 , w_8341 , w_8342 , w_8343 , w_8344 , w_8345 , 
		w_8346 , w_8347 , w_8348 , w_8349 , w_8350 , w_8351 , w_8352 , w_8353 , w_8354 , w_8355 , 
		w_8356 , w_8357 , w_8358 , w_8359 , w_8360 , w_8361 , w_8362 , w_8363 , w_8364 , w_8365 , 
		w_8366 , w_8367 , w_8368 , w_8369 , w_8370 , w_8371 , w_8372 , w_8373 , w_8374 , w_8375 , 
		w_8376 , w_8377 , w_8378 , w_8379 , w_8380 , w_8381 , w_8382 , w_8383 , w_8384 , w_8385 , 
		w_8386 , w_8387 , w_8388 , w_8389 , w_8390 , w_8391 , w_8392 , w_8393 , w_8394 , w_8395 , 
		w_8396 , w_8397 , w_8398 , w_8399 , w_8400 , w_8401 , w_8402 , w_8403 , w_8404 , w_8405 , 
		w_8406 , w_8407 , w_8408 , w_8409 , w_8410 , w_8411 , w_8412 , w_8413 , w_8414 , w_8415 , 
		w_8416 , w_8417 , w_8418 , w_8419 , w_8420 , w_8421 , w_8422 , w_8423 , w_8424 , w_8425 , 
		w_8426 , w_8427 , w_8428 , w_8429 , w_8430 , w_8431 , w_8432 , w_8433 , w_8434 , w_8435 , 
		w_8436 , w_8437 , w_8438 , w_8439 , w_8440 , w_8441 , w_8442 , w_8443 , w_8444 , w_8445 , 
		w_8446 , w_8447 , w_8448 , w_8449 , w_8450 , w_8451 , w_8452 , w_8453 , w_8454 , w_8455 , 
		w_8456 , w_8457 , w_8458 , w_8459 , w_8460 , w_8461 , w_8462 , w_8463 , w_8464 , w_8465 , 
		w_8466 , w_8467 , w_8468 , w_8469 , w_8470 , w_8471 , w_8472 , w_8473 , w_8474 , w_8475 , 
		w_8476 , w_8477 , w_8478 , w_8479 , w_8480 , w_8481 , w_8482 , w_8483 , w_8484 , w_8485 , 
		w_8486 , w_8487 , w_8488 , w_8489 , w_8490 , w_8491 , w_8492 , w_8493 , w_8494 , w_8495 , 
		w_8496 , w_8497 , w_8498 , w_8499 , w_8500 , w_8501 , w_8502 , w_8503 , w_8504 , w_8505 , 
		w_8506 , w_8507 , w_8508 , w_8509 , w_8510 , w_8511 , w_8512 , w_8513 , w_8514 , w_8515 , 
		w_8516 , w_8517 , w_8518 , w_8519 , w_8520 , w_8521 , w_8522 , w_8523 , w_8524 , w_8525 , 
		w_8526 , w_8527 , w_8528 , w_8529 , w_8530 , w_8531 , w_8532 , w_8533 , w_8534 , w_8535 , 
		w_8536 , w_8537 , w_8538 , w_8539 , w_8540 , w_8541 , w_8542 , w_8543 , w_8544 , w_8545 , 
		w_8546 , w_8547 , w_8548 , w_8549 , w_8550 , w_8551 , w_8552 , w_8553 , w_8554 , w_8555 , 
		w_8556 , w_8557 , w_8558 , w_8559 , w_8560 , w_8561 , w_8562 , w_8563 , w_8564 , w_8565 , 
		w_8566 , w_8567 , w_8568 , w_8569 , w_8570 , w_8571 , w_8572 , w_8573 , w_8574 , w_8575 , 
		w_8576 , w_8577 , w_8578 , w_8579 , w_8580 , w_8581 , w_8582 , w_8583 , w_8584 , w_8585 , 
		w_8586 , w_8587 , w_8588 , w_8589 , w_8590 , w_8591 , w_8592 , w_8593 , w_8594 , w_8595 , 
		w_8596 , w_8597 , w_8598 , w_8599 , w_8600 , w_8601 , w_8602 , w_8603 , w_8604 , w_8605 , 
		w_8606 , w_8607 , w_8608 , w_8609 , w_8610 , w_8611 , w_8612 , w_8613 , w_8614 , w_8615 , 
		w_8616 , w_8617 , w_8618 , w_8619 , w_8620 , w_8621 , w_8622 , w_8623 , w_8624 , w_8625 , 
		w_8626 , w_8627 , w_8628 , w_8629 , w_8630 , w_8631 , w_8632 , w_8633 , w_8634 , w_8635 , 
		w_8636 , w_8637 , w_8638 , w_8639 , w_8640 , w_8641 , w_8642 , w_8643 , w_8644 , w_8645 , 
		w_8646 , w_8647 , w_8648 , w_8649 , w_8650 , w_8651 , w_8652 , w_8653 , w_8654 , w_8655 , 
		w_8656 , w_8657 , w_8658 , w_8659 , w_8660 , w_8661 , w_8662 , w_8663 , w_8664 , w_8665 , 
		w_8666 , w_8667 , w_8668 , w_8669 , w_8670 , w_8671 , w_8672 , w_8673 , w_8674 , w_8675 , 
		w_8676 , w_8677 , w_8678 , w_8679 , w_8680 , w_8681 , w_8682 , w_8683 , w_8684 , w_8685 , 
		w_8686 , w_8687 , w_8688 , w_8689 , w_8690 , w_8691 , w_8692 , w_8693 , w_8694 , w_8695 , 
		w_8696 , w_8697 , w_8698 , w_8699 , w_8700 , w_8701 , w_8702 , w_8703 , w_8704 , w_8705 , 
		w_8706 , w_8707 , w_8708 , w_8709 , w_8710 , w_8711 , w_8712 , w_8713 , w_8714 , w_8715 , 
		w_8716 , w_8717 , w_8718 , w_8719 , w_8720 , w_8721 , w_8722 , w_8723 , w_8724 , w_8725 , 
		w_8726 , w_8727 , w_8728 , w_8729 , w_8730 , w_8731 , w_8732 , w_8733 , w_8734 , w_8735 , 
		w_8736 , w_8737 , w_8738 , w_8739 , w_8740 , w_8741 , w_8742 , w_8743 , w_8744 , w_8745 , 
		w_8746 , w_8747 , w_8748 , w_8749 , w_8750 , w_8751 , w_8752 , w_8753 , w_8754 , w_8755 , 
		w_8756 , w_8757 , w_8758 , w_8759 , w_8760 , w_8761 , w_8762 , w_8763 , w_8764 , w_8765 , 
		w_8766 , w_8767 , w_8768 , w_8769 , w_8770 , w_8771 , w_8772 , w_8773 , w_8774 , w_8775 , 
		w_8776 , w_8777 , w_8778 , w_8779 , w_8780 , w_8781 , w_8782 , w_8783 , w_8784 , w_8785 , 
		w_8786 , w_8787 , w_8788 , w_8789 , w_8790 , w_8791 , w_8792 , w_8793 , w_8794 , w_8795 , 
		w_8796 , w_8797 , w_8798 , w_8799 , w_8800 , w_8801 , w_8802 , w_8803 , w_8804 , w_8805 , 
		w_8806 , w_8807 , w_8808 , w_8809 , w_8810 , w_8811 , w_8812 , w_8813 , w_8814 , w_8815 , 
		w_8816 , w_8817 , w_8818 , w_8819 , w_8820 , w_8821 , w_8822 , w_8823 , w_8824 , w_8825 , 
		w_8826 , w_8827 , w_8828 , w_8829 , w_8830 , w_8831 , w_8832 , w_8833 , w_8834 , w_8835 , 
		w_8836 , w_8837 , w_8838 , w_8839 , w_8840 , w_8841 , w_8842 , w_8843 , w_8844 , w_8845 , 
		w_8846 , w_8847 , w_8848 , w_8849 , w_8850 , w_8851 , w_8852 , w_8853 , w_8854 , w_8855 , 
		w_8856 , w_8857 , w_8858 , w_8859 , w_8860 , w_8861 , w_8862 , w_8863 , w_8864 , w_8865 , 
		w_8866 , w_8867 , w_8868 , w_8869 , w_8870 , w_8871 , w_8872 , w_8873 , w_8874 , w_8875 , 
		w_8876 , w_8877 , w_8878 , w_8879 , w_8880 , w_8881 , w_8882 , w_8883 , w_8884 , w_8885 , 
		w_8886 , w_8887 , w_8888 , w_8889 , w_8890 , w_8891 , w_8892 , w_8893 , w_8894 , w_8895 , 
		w_8896 , w_8897 , w_8898 , w_8899 , w_8900 , w_8901 , w_8902 , w_8903 , w_8904 , w_8905 , 
		w_8906 , w_8907 , w_8908 , w_8909 , w_8910 , w_8911 , w_8912 , w_8913 , w_8914 , w_8915 , 
		w_8916 , w_8917 , w_8918 , w_8919 , w_8920 , w_8921 , w_8922 , w_8923 , w_8924 , w_8925 , 
		w_8926 , w_8927 , w_8928 , w_8929 , w_8930 , w_8931 , w_8932 , w_8933 , w_8934 , w_8935 , 
		w_8936 , w_8937 , w_8938 , w_8939 , w_8940 , w_8941 , w_8942 , w_8943 , w_8944 , w_8945 , 
		w_8946 , w_8947 , w_8948 , w_8949 , w_8950 , w_8951 , w_8952 , w_8953 , w_8954 , w_8955 , 
		w_8956 , w_8957 , w_8958 , w_8959 , w_8960 , w_8961 , w_8962 , w_8963 , w_8964 , w_8965 , 
		w_8966 , w_8967 , w_8968 , w_8969 , w_8970 , w_8971 , w_8972 , w_8973 , w_8974 , w_8975 , 
		w_8976 , w_8977 , w_8978 , w_8979 , w_8980 , w_8981 , w_8982 , w_8983 , w_8984 , w_8985 , 
		w_8986 , w_8987 , w_8988 , w_8989 , w_8990 , w_8991 , w_8992 , w_8993 , w_8994 , w_8995 , 
		w_8996 , w_8997 , w_8998 , w_8999 , w_9000 , w_9001 , w_9002 , w_9003 , w_9004 , w_9005 , 
		w_9006 , w_9007 , w_9008 , w_9009 , w_9010 , w_9011 , w_9012 , w_9013 , w_9014 , w_9015 , 
		w_9016 , w_9017 , w_9018 , w_9019 , w_9020 , w_9021 , w_9022 , w_9023 , w_9024 , w_9025 , 
		w_9026 , w_9027 , w_9028 , w_9029 , w_9030 , w_9031 , w_9032 , w_9033 , w_9034 , w_9035 , 
		w_9036 , w_9037 , w_9038 , w_9039 , w_9040 , w_9041 , w_9042 , w_9043 , w_9044 , w_9045 , 
		w_9046 , w_9047 , w_9048 , w_9049 , w_9050 , w_9051 , w_9052 , w_9053 , w_9054 , w_9055 , 
		w_9056 , w_9057 , w_9058 , w_9059 , w_9060 , w_9061 , w_9062 , w_9063 , w_9064 , w_9065 , 
		w_9066 , w_9067 , w_9068 , w_9069 , w_9070 , w_9071 , w_9072 , w_9073 , w_9074 , w_9075 , 
		w_9076 , w_9077 , w_9078 , w_9079 , w_9080 , w_9081 , w_9082 , w_9083 , w_9084 , w_9085 , 
		w_9086 , w_9087 , w_9088 , w_9089 , w_9090 , w_9091 , w_9092 , w_9093 , w_9094 , w_9095 , 
		w_9096 , w_9097 , w_9098 , w_9099 , w_9100 , w_9101 , w_9102 , w_9103 , w_9104 , w_9105 , 
		w_9106 , w_9107 , w_9108 , w_9109 , w_9110 , w_9111 , w_9112 , w_9113 , w_9114 , w_9115 , 
		w_9116 , w_9117 , w_9118 , w_9119 , w_9120 , w_9121 , w_9122 , w_9123 , w_9124 , w_9125 , 
		w_9126 , w_9127 , w_9128 , w_9129 , w_9130 , w_9131 , w_9132 , w_9133 , w_9134 , w_9135 , 
		w_9136 , w_9137 , w_9138 , w_9139 , w_9140 , w_9141 , w_9142 , w_9143 , w_9144 , w_9145 , 
		w_9146 , w_9147 , w_9148 , w_9149 , w_9150 , w_9151 , w_9152 , w_9153 , w_9154 , w_9155 , 
		w_9156 , w_9157 , w_9158 , w_9159 , w_9160 , w_9161 , w_9162 , w_9163 , w_9164 , w_9165 , 
		w_9166 , w_9167 , w_9168 , w_9169 , w_9170 , w_9171 , w_9172 , w_9173 , w_9174 , w_9175 , 
		w_9176 , w_9177 , w_9178 , w_9179 , w_9180 , w_9181 , w_9182 , w_9183 , w_9184 , w_9185 , 
		w_9186 , w_9187 , w_9188 , w_9189 , w_9190 , w_9191 , w_9192 , w_9193 , w_9194 , w_9195 , 
		w_9196 , w_9197 , w_9198 , w_9199 , w_9200 , w_9201 , w_9202 , w_9203 , w_9204 , w_9205 , 
		w_9206 , w_9207 , w_9208 , w_9209 , w_9210 , w_9211 , w_9212 , w_9213 , w_9214 , w_9215 , 
		w_9216 , w_9217 , w_9218 , w_9219 , w_9220 , w_9221 , w_9222 , w_9223 , w_9224 , w_9225 , 
		w_9226 , w_9227 , w_9228 , w_9229 , w_9230 , w_9231 , w_9232 , w_9233 , w_9234 , w_9235 , 
		w_9236 , w_9237 , w_9238 , w_9239 , w_9240 , w_9241 , w_9242 , w_9243 , w_9244 , w_9245 , 
		w_9246 , w_9247 , w_9248 , w_9249 , w_9250 , w_9251 , w_9252 , w_9253 , w_9254 , w_9255 , 
		w_9256 , w_9257 , w_9258 , w_9259 , w_9260 , w_9261 , w_9262 , w_9263 , w_9264 , w_9265 , 
		w_9266 , w_9267 , w_9268 , w_9269 , w_9270 , w_9271 , w_9272 , w_9273 , w_9274 , w_9275 , 
		w_9276 , w_9277 , w_9278 , w_9279 , w_9280 , w_9281 , w_9282 , w_9283 , w_9284 , w_9285 , 
		w_9286 , w_9287 , w_9288 , w_9289 , w_9290 , w_9291 , w_9292 , w_9293 , w_9294 , w_9295 , 
		w_9296 , w_9297 , w_9298 , w_9299 , w_9300 , w_9301 , w_9302 , w_9303 , w_9304 , w_9305 , 
		w_9306 , w_9307 , w_9308 , w_9309 , w_9310 , w_9311 , w_9312 , w_9313 , w_9314 , w_9315 , 
		w_9316 , w_9317 , w_9318 , w_9319 , w_9320 , w_9321 , w_9322 , w_9323 , w_9324 , w_9325 , 
		w_9326 , w_9327 , w_9328 , w_9329 , w_9330 , w_9331 , w_9332 , w_9333 , w_9334 , w_9335 , 
		w_9336 , w_9337 , w_9338 , w_9339 , w_9340 , w_9341 , w_9342 , w_9343 , w_9344 , w_9345 , 
		w_9346 , w_9347 , w_9348 , w_9349 , w_9350 , w_9351 , w_9352 , w_9353 , w_9354 , w_9355 , 
		w_9356 , w_9357 , w_9358 , w_9359 , w_9360 , w_9361 , w_9362 , w_9363 , w_9364 , w_9365 , 
		w_9366 , w_9367 , w_9368 , w_9369 , w_9370 , w_9371 , w_9372 , w_9373 , w_9374 , w_9375 , 
		w_9376 , w_9377 , w_9378 , w_9379 , w_9380 , w_9381 , w_9382 , w_9383 , w_9384 , w_9385 , 
		w_9386 , w_9387 , w_9388 , w_9389 , w_9390 , w_9391 , w_9392 , w_9393 , w_9394 , w_9395 , 
		w_9396 , w_9397 , w_9398 , w_9399 , w_9400 , w_9401 , w_9402 , w_9403 , w_9404 , w_9405 , 
		w_9406 , w_9407 , w_9408 , w_9409 , w_9410 , w_9411 , w_9412 , w_9413 , w_9414 , w_9415 , 
		w_9416 , w_9417 , w_9418 , w_9419 , w_9420 , w_9421 , w_9422 , w_9423 , w_9424 , w_9425 , 
		w_9426 , w_9427 , w_9428 , w_9429 , w_9430 , w_9431 , w_9432 , w_9433 , w_9434 , w_9435 , 
		w_9436 , w_9437 , w_9438 , w_9439 , w_9440 , w_9441 , w_9442 , w_9443 , w_9444 , w_9445 , 
		w_9446 , w_9447 , w_9448 , w_9449 , w_9450 , w_9451 , w_9452 , w_9453 , w_9454 , w_9455 , 
		w_9456 , w_9457 , w_9458 , w_9459 , w_9460 , w_9461 , w_9462 , w_9463 , w_9464 , w_9465 , 
		w_9466 , w_9467 , w_9468 , w_9469 , w_9470 , w_9471 , w_9472 , w_9473 , w_9474 , w_9475 , 
		w_9476 , w_9477 , w_9478 , w_9479 , w_9480 , w_9481 , w_9482 , w_9483 , w_9484 , w_9485 , 
		w_9486 , w_9487 , w_9488 , w_9489 , w_9490 , w_9491 , w_9492 , w_9493 , w_9494 , w_9495 , 
		w_9496 , w_9497 , w_9498 , w_9499 , w_9500 , w_9501 , w_9502 , w_9503 , w_9504 , w_9505 , 
		w_9506 , w_9507 , w_9508 , w_9509 , w_9510 , w_9511 , w_9512 , w_9513 , w_9514 , w_9515 , 
		w_9516 , w_9517 , w_9518 , w_9519 , w_9520 , w_9521 , w_9522 , w_9523 , w_9524 , w_9525 , 
		w_9526 , w_9527 , w_9528 , w_9529 , w_9530 , w_9531 , w_9532 , w_9533 , w_9534 , w_9535 , 
		w_9536 , w_9537 , w_9538 , w_9539 , w_9540 , w_9541 , w_9542 , w_9543 , w_9544 , w_9545 , 
		w_9546 , w_9547 , w_9548 , w_9549 , w_9550 , w_9551 , w_9552 , w_9553 , w_9554 , w_9555 , 
		w_9556 , w_9557 , w_9558 , w_9559 , w_9560 , w_9561 , w_9562 , w_9563 , w_9564 , w_9565 , 
		w_9566 , w_9567 , w_9568 , w_9569 , w_9570 , w_9571 , w_9572 , w_9573 , w_9574 , w_9575 , 
		w_9576 , w_9577 , w_9578 , w_9579 , w_9580 , w_9581 , w_9582 , w_9583 , w_9584 , w_9585 , 
		w_9586 , w_9587 , w_9588 , w_9589 , w_9590 , w_9591 , w_9592 , w_9593 , w_9594 , w_9595 , 
		w_9596 , w_9597 , w_9598 , w_9599 , w_9600 , w_9601 , w_9602 , w_9603 , w_9604 , w_9605 , 
		w_9606 , w_9607 , w_9608 , w_9609 , w_9610 , w_9611 , w_9612 , w_9613 , w_9614 , w_9615 , 
		w_9616 , w_9617 , w_9618 , w_9619 , w_9620 , w_9621 , w_9622 , w_9623 , w_9624 , w_9625 , 
		w_9626 , w_9627 , w_9628 , w_9629 , w_9630 , w_9631 , w_9632 , w_9633 , w_9634 , w_9635 , 
		w_9636 , w_9637 , w_9638 , w_9639 , w_9640 , w_9641 , w_9642 , w_9643 , w_9644 , w_9645 , 
		w_9646 , w_9647 , w_9648 , w_9649 , w_9650 , w_9651 , w_9652 , w_9653 , w_9654 , w_9655 , 
		w_9656 , w_9657 , w_9658 , w_9659 , w_9660 , w_9661 , w_9662 , w_9663 , w_9664 , w_9665 , 
		w_9666 , w_9667 , w_9668 , w_9669 , w_9670 , w_9671 , w_9672 , w_9673 , w_9674 , w_9675 , 
		w_9676 , w_9677 , w_9678 , w_9679 , w_9680 , w_9681 , w_9682 , w_9683 , w_9684 , w_9685 , 
		w_9686 , w_9687 , w_9688 , w_9689 , w_9690 , w_9691 , w_9692 , w_9693 , w_9694 , w_9695 , 
		w_9696 , w_9697 , w_9698 , w_9699 , w_9700 , w_9701 , w_9702 , w_9703 , w_9704 , w_9705 , 
		w_9706 , w_9707 , w_9708 , w_9709 , w_9710 , w_9711 , w_9712 , w_9713 , w_9714 , w_9715 , 
		w_9716 , w_9717 , w_9718 , w_9719 , w_9720 , w_9721 , w_9722 , w_9723 , w_9724 , w_9725 , 
		w_9726 , w_9727 , w_9728 , w_9729 , w_9730 , w_9731 , w_9732 , w_9733 , w_9734 , w_9735 , 
		w_9736 , w_9737 , w_9738 , w_9739 , w_9740 , w_9741 , w_9742 , w_9743 , w_9744 , w_9745 , 
		w_9746 , w_9747 , w_9748 , w_9749 , w_9750 , w_9751 , w_9752 , w_9753 , w_9754 , w_9755 , 
		w_9756 , w_9757 , w_9758 , w_9759 , w_9760 , w_9761 , w_9762 , w_9763 , w_9764 , w_9765 , 
		w_9766 , w_9767 , w_9768 , w_9769 , w_9770 , w_9771 , w_9772 , w_9773 , w_9774 , w_9775 , 
		w_9776 , w_9777 , w_9778 , w_9779 , w_9780 , w_9781 , w_9782 , w_9783 , w_9784 , w_9785 , 
		w_9786 , w_9787 , w_9788 , w_9789 , w_9790 , w_9791 , w_9792 , w_9793 , w_9794 , w_9795 , 
		w_9796 , w_9797 , w_9798 , w_9799 , w_9800 , w_9801 , w_9802 , w_9803 , w_9804 , w_9805 , 
		w_9806 , w_9807 , w_9808 , w_9809 , w_9810 , w_9811 , w_9812 , w_9813 , w_9814 , w_9815 , 
		w_9816 , w_9817 , w_9818 , w_9819 , w_9820 , w_9821 , w_9822 , w_9823 , w_9824 , w_9825 , 
		w_9826 , w_9827 , w_9828 , w_9829 , w_9830 , w_9831 , w_9832 , w_9833 , w_9834 , w_9835 , 
		w_9836 , w_9837 , w_9838 , w_9839 , w_9840 , w_9841 , w_9842 , w_9843 , w_9844 , w_9845 , 
		w_9846 , w_9847 , w_9848 , w_9849 , w_9850 , w_9851 , w_9852 , w_9853 , w_9854 , w_9855 , 
		w_9856 , w_9857 , w_9858 , w_9859 , w_9860 , w_9861 , w_9862 , w_9863 , w_9864 , w_9865 , 
		w_9866 , w_9867 , w_9868 , w_9869 , w_9870 , w_9871 , w_9872 , w_9873 , w_9874 , w_9875 , 
		w_9876 , w_9877 , w_9878 , w_9879 , w_9880 , w_9881 , w_9882 , w_9883 , w_9884 , w_9885 , 
		w_9886 , w_9887 , w_9888 , w_9889 , w_9890 , w_9891 , w_9892 , w_9893 , w_9894 , w_9895 , 
		w_9896 , w_9897 , w_9898 , w_9899 , w_9900 , w_9901 , w_9902 , w_9903 , w_9904 , w_9905 , 
		w_9906 , w_9907 , w_9908 , w_9909 , w_9910 , w_9911 , w_9912 , w_9913 , w_9914 , w_9915 , 
		w_9916 , w_9917 , w_9918 , w_9919 , w_9920 , w_9921 , w_9922 , w_9923 , w_9924 , w_9925 , 
		w_9926 , w_9927 , w_9928 , w_9929 , w_9930 , w_9931 , w_9932 , w_9933 , w_9934 , w_9935 , 
		w_9936 , w_9937 , w_9938 , w_9939 , w_9940 , w_9941 , w_9942 , w_9943 , w_9944 , w_9945 , 
		w_9946 , w_9947 , w_9948 , w_9949 , w_9950 , w_9951 , w_9952 , w_9953 , w_9954 , w_9955 , 
		w_9956 , w_9957 , w_9958 , w_9959 , w_9960 , w_9961 , w_9962 , w_9963 , w_9964 , w_9965 , 
		w_9966 , w_9967 , w_9968 , w_9969 , w_9970 , w_9971 , w_9972 , w_9973 , w_9974 , w_9975 , 
		w_9976 , w_9977 , w_9978 , w_9979 , w_9980 , w_9981 , w_9982 , w_9983 , w_9984 , w_9985 , 
		w_9986 , w_9987 , w_9988 , w_9989 , w_9990 , w_9991 , w_9992 , w_9993 , w_9994 , w_9995 , 
		w_9996 , w_9997 , w_9998 , w_9999 , w_10000 , w_10001 , w_10002 , w_10003 , w_10004 , w_10005 , 
		w_10006 , w_10007 , w_10008 , w_10009 , w_10010 , w_10011 , w_10012 , w_10013 , w_10014 , w_10015 , 
		w_10016 , w_10017 , w_10018 , w_10019 , w_10020 , w_10021 , w_10022 , w_10023 , w_10024 , w_10025 , 
		w_10026 , w_10027 , w_10028 , w_10029 , w_10030 , w_10031 , w_10032 , w_10033 , w_10034 , w_10035 , 
		w_10036 , w_10037 , w_10038 , w_10039 , w_10040 , w_10041 , w_10042 , w_10043 , w_10044 , w_10045 , 
		w_10046 , w_10047 , w_10048 , w_10049 , w_10050 , w_10051 , w_10052 , w_10053 , w_10054 , w_10055 , 
		w_10056 , w_10057 , w_10058 , w_10059 , w_10060 , w_10061 , w_10062 , w_10063 , w_10064 , w_10065 , 
		w_10066 , w_10067 , w_10068 , w_10069 , w_10070 , w_10071 , w_10072 , w_10073 , w_10074 , w_10075 , 
		w_10076 , w_10077 , w_10078 , w_10079 , w_10080 , w_10081 , w_10082 , w_10083 , w_10084 , w_10085 , 
		w_10086 , w_10087 , w_10088 , w_10089 , w_10090 , w_10091 , w_10092 , w_10093 , w_10094 , w_10095 , 
		w_10096 , w_10097 , w_10098 , w_10099 , w_10100 , w_10101 , w_10102 , w_10103 , w_10104 , w_10105 , 
		w_10106 , w_10107 , w_10108 , w_10109 , w_10110 , w_10111 , w_10112 , w_10113 , w_10114 , w_10115 , 
		w_10116 , w_10117 , w_10118 , w_10119 , w_10120 , w_10121 , w_10122 , w_10123 , w_10124 , w_10125 , 
		w_10126 , w_10127 , w_10128 , w_10129 , w_10130 , w_10131 , w_10132 , w_10133 , w_10134 , w_10135 , 
		w_10136 , w_10137 , w_10138 , w_10139 , w_10140 , w_10141 , w_10142 , w_10143 , w_10144 , w_10145 , 
		w_10146 , w_10147 , w_10148 , w_10149 , w_10150 , w_10151 , w_10152 , w_10153 , w_10154 , w_10155 , 
		w_10156 , w_10157 , w_10158 , w_10159 , w_10160 , w_10161 , w_10162 , w_10163 , w_10164 , w_10165 , 
		w_10166 , w_10167 , w_10168 , w_10169 , w_10170 , w_10171 , w_10172 , w_10173 , w_10174 , w_10175 , 
		w_10176 , w_10177 , w_10178 , w_10179 , w_10180 , w_10181 , w_10182 , w_10183 , w_10184 , w_10185 , 
		w_10186 , w_10187 , w_10188 , w_10189 , w_10190 , w_10191 , w_10192 , w_10193 , w_10194 , w_10195 , 
		w_10196 , w_10197 , w_10198 , w_10199 , w_10200 , w_10201 , w_10202 , w_10203 , w_10204 , w_10205 , 
		w_10206 , w_10207 , w_10208 , w_10209 , w_10210 , w_10211 , w_10212 , w_10213 , w_10214 , w_10215 , 
		w_10216 , w_10217 , w_10218 , w_10219 , w_10220 , w_10221 , w_10222 , w_10223 , w_10224 , w_10225 , 
		w_10226 , w_10227 , w_10228 , w_10229 , w_10230 , w_10231 , w_10232 , w_10233 , w_10234 , w_10235 , 
		w_10236 , w_10237 , w_10238 , w_10239 , w_10240 , w_10241 , w_10242 , w_10243 , w_10244 , w_10245 , 
		w_10246 , w_10247 , w_10248 , w_10249 , w_10250 , w_10251 , w_10252 , w_10253 , w_10254 , w_10255 , 
		w_10256 , w_10257 , w_10258 , w_10259 , w_10260 , w_10261 , w_10262 , w_10263 , w_10264 , w_10265 , 
		w_10266 , w_10267 , w_10268 , w_10269 , w_10270 , w_10271 , w_10272 , w_10273 , w_10274 , w_10275 , 
		w_10276 , w_10277 , w_10278 , w_10279 , w_10280 , w_10281 , w_10282 , w_10283 , w_10284 , w_10285 , 
		w_10286 , w_10287 , w_10288 , w_10289 , w_10290 , w_10291 , w_10292 , w_10293 , w_10294 , w_10295 , 
		w_10296 , w_10297 , w_10298 , w_10299 , w_10300 , w_10301 , w_10302 , w_10303 , w_10304 , w_10305 , 
		w_10306 , w_10307 , w_10308 , w_10309 , w_10310 , w_10311 , w_10312 , w_10313 , w_10314 , w_10315 , 
		w_10316 , w_10317 , w_10318 , w_10319 , w_10320 , w_10321 , w_10322 , w_10323 , w_10324 , w_10325 , 
		w_10326 , w_10327 , w_10328 , w_10329 , w_10330 , w_10331 , w_10332 , w_10333 , w_10334 , w_10335 , 
		w_10336 , w_10337 , w_10338 , w_10339 , w_10340 , w_10341 , w_10342 , w_10343 , w_10344 , w_10345 , 
		w_10346 , w_10347 , w_10348 , w_10349 , w_10350 , w_10351 , w_10352 , w_10353 , w_10354 , w_10355 , 
		w_10356 , w_10357 , w_10358 , w_10359 , w_10360 , w_10361 , w_10362 , w_10363 , w_10364 , w_10365 , 
		w_10366 , w_10367 , w_10368 , w_10369 , w_10370 , w_10371 , w_10372 , w_10373 , w_10374 , w_10375 , 
		w_10376 , w_10377 , w_10378 , w_10379 , w_10380 , w_10381 , w_10382 , w_10383 , w_10384 , w_10385 , 
		w_10386 , w_10387 , w_10388 , w_10389 , w_10390 , w_10391 , w_10392 , w_10393 , w_10394 , w_10395 , 
		w_10396 , w_10397 , w_10398 , w_10399 , w_10400 , w_10401 , w_10402 , w_10403 , w_10404 , w_10405 , 
		w_10406 , w_10407 , w_10408 , w_10409 , w_10410 , w_10411 , w_10412 , w_10413 , w_10414 , w_10415 , 
		w_10416 , w_10417 , w_10418 , w_10419 , w_10420 , w_10421 , w_10422 , w_10423 , w_10424 , w_10425 , 
		w_10426 , w_10427 , w_10428 , w_10429 , w_10430 , w_10431 , w_10432 , w_10433 , w_10434 , w_10435 , 
		w_10436 , w_10437 , w_10438 , w_10439 , w_10440 , w_10441 , w_10442 , w_10443 , w_10444 , w_10445 , 
		w_10446 , w_10447 , w_10448 , w_10449 , w_10450 , w_10451 , w_10452 , w_10453 , w_10454 , w_10455 , 
		w_10456 , w_10457 , w_10458 , w_10459 , w_10460 , w_10461 , w_10462 , w_10463 , w_10464 , w_10465 , 
		w_10466 , w_10467 , w_10468 , w_10469 , w_10470 , w_10471 , w_10472 , w_10473 , w_10474 , w_10475 , 
		w_10476 , w_10477 , w_10478 , w_10479 , w_10480 , w_10481 , w_10482 , w_10483 , w_10484 , w_10485 , 
		w_10486 , w_10487 , w_10488 , w_10489 , w_10490 , w_10491 , w_10492 , w_10493 , w_10494 , w_10495 , 
		w_10496 , w_10497 , w_10498 , w_10499 , w_10500 , w_10501 , w_10502 , w_10503 , w_10504 , w_10505 , 
		w_10506 , w_10507 , w_10508 , w_10509 , w_10510 , w_10511 , w_10512 , w_10513 , w_10514 , w_10515 , 
		w_10516 , w_10517 , w_10518 , w_10519 , w_10520 , w_10521 , w_10522 , w_10523 , w_10524 , w_10525 , 
		w_10526 , w_10527 , w_10528 , w_10529 , w_10530 , w_10531 , w_10532 , w_10533 , w_10534 , w_10535 , 
		w_10536 , w_10537 , w_10538 , w_10539 , w_10540 , w_10541 , w_10542 , w_10543 , w_10544 , w_10545 , 
		w_10546 , w_10547 , w_10548 , w_10549 , w_10550 , w_10551 , w_10552 , w_10553 , w_10554 , w_10555 , 
		w_10556 , w_10557 , w_10558 , w_10559 , w_10560 , w_10561 , w_10562 , w_10563 , w_10564 , w_10565 , 
		w_10566 , w_10567 , w_10568 , w_10569 , w_10570 , w_10571 , w_10572 , w_10573 , w_10574 , w_10575 , 
		w_10576 , w_10577 , w_10578 , w_10579 , w_10580 , w_10581 , w_10582 , w_10583 , w_10584 , w_10585 , 
		w_10586 , w_10587 , w_10588 , w_10589 , w_10590 , w_10591 , w_10592 , w_10593 , w_10594 , w_10595 , 
		w_10596 , w_10597 , w_10598 , w_10599 , w_10600 , w_10601 , w_10602 , w_10603 , w_10604 , w_10605 , 
		w_10606 , w_10607 , w_10608 , w_10609 , w_10610 , w_10611 , w_10612 , w_10613 , w_10614 , w_10615 , 
		w_10616 , w_10617 , w_10618 , w_10619 , w_10620 , w_10621 , w_10622 , w_10623 , w_10624 , w_10625 , 
		w_10626 , w_10627 , w_10628 , w_10629 , w_10630 , w_10631 , w_10632 , w_10633 , w_10634 , w_10635 , 
		w_10636 , w_10637 , w_10638 , w_10639 , w_10640 , w_10641 , w_10642 , w_10643 , w_10644 , w_10645 , 
		w_10646 , w_10647 , w_10648 , w_10649 , w_10650 , w_10651 , w_10652 , w_10653 , w_10654 , w_10655 , 
		w_10656 , w_10657 , w_10658 , w_10659 , w_10660 , w_10661 , w_10662 , w_10663 , w_10664 , w_10665 , 
		w_10666 , w_10667 , w_10668 , w_10669 , w_10670 , w_10671 , w_10672 , w_10673 , w_10674 , w_10675 , 
		w_10676 , w_10677 , w_10678 , w_10679 , w_10680 , w_10681 , w_10682 , w_10683 , w_10684 , w_10685 , 
		w_10686 , w_10687 , w_10688 , w_10689 , w_10690 , w_10691 , w_10692 , w_10693 , w_10694 , w_10695 , 
		w_10696 , w_10697 , w_10698 , w_10699 , w_10700 , w_10701 , w_10702 , w_10703 , w_10704 , w_10705 , 
		w_10706 , w_10707 , w_10708 , w_10709 , w_10710 , w_10711 , w_10712 , w_10713 , w_10714 , w_10715 , 
		w_10716 , w_10717 , w_10718 , w_10719 , w_10720 , w_10721 , w_10722 , w_10723 , w_10724 , w_10725 , 
		w_10726 , w_10727 , w_10728 , w_10729 , w_10730 , w_10731 , w_10732 , w_10733 , w_10734 , w_10735 , 
		w_10736 , w_10737 , w_10738 , w_10739 , w_10740 , w_10741 , w_10742 , w_10743 , w_10744 , w_10745 , 
		w_10746 , w_10747 , w_10748 , w_10749 , w_10750 , w_10751 , w_10752 , w_10753 , w_10754 , w_10755 , 
		w_10756 , w_10757 , w_10758 , w_10759 , w_10760 , w_10761 , w_10762 , w_10763 , w_10764 , w_10765 , 
		w_10766 , w_10767 , w_10768 , w_10769 , w_10770 , w_10771 , w_10772 , w_10773 , w_10774 , w_10775 , 
		w_10776 , w_10777 , w_10778 , w_10779 , w_10780 , w_10781 , w_10782 , w_10783 , w_10784 , w_10785 , 
		w_10786 , w_10787 , w_10788 , w_10789 , w_10790 , w_10791 , w_10792 , w_10793 , w_10794 , w_10795 , 
		w_10796 , w_10797 , w_10798 , w_10799 , w_10800 , w_10801 , w_10802 , w_10803 , w_10804 , w_10805 , 
		w_10806 , w_10807 , w_10808 , w_10809 , w_10810 , w_10811 , w_10812 , w_10813 , w_10814 , w_10815 , 
		w_10816 , w_10817 , w_10818 , w_10819 , w_10820 , w_10821 , w_10822 , w_10823 , w_10824 , w_10825 , 
		w_10826 , w_10827 , w_10828 , w_10829 , w_10830 , w_10831 , w_10832 , w_10833 , w_10834 , w_10835 , 
		w_10836 , w_10837 , w_10838 , w_10839 , w_10840 , w_10841 , w_10842 , w_10843 , w_10844 , w_10845 , 
		w_10846 , w_10847 , w_10848 , w_10849 , w_10850 , w_10851 , w_10852 , w_10853 , w_10854 , w_10855 , 
		w_10856 , w_10857 , w_10858 , w_10859 , w_10860 , w_10861 , w_10862 , w_10863 , w_10864 , w_10865 , 
		w_10866 , w_10867 , w_10868 , w_10869 , w_10870 , w_10871 , w_10872 , w_10873 , w_10874 , w_10875 , 
		w_10876 , w_10877 , w_10878 , w_10879 , w_10880 , w_10881 , w_10882 , w_10883 , w_10884 , w_10885 , 
		w_10886 , w_10887 , w_10888 , w_10889 , w_10890 , w_10891 , w_10892 , w_10893 , w_10894 , w_10895 , 
		w_10896 , w_10897 , w_10898 , w_10899 , w_10900 , w_10901 , w_10902 , w_10903 , w_10904 , w_10905 , 
		w_10906 , w_10907 , w_10908 , w_10909 , w_10910 , w_10911 , w_10912 , w_10913 , w_10914 , w_10915 , 
		w_10916 , w_10917 , w_10918 , w_10919 , w_10920 , w_10921 , w_10922 , w_10923 , w_10924 , w_10925 , 
		w_10926 , w_10927 , w_10928 , w_10929 , w_10930 , w_10931 , w_10932 , w_10933 , w_10934 , w_10935 , 
		w_10936 , w_10937 , w_10938 , w_10939 , w_10940 , w_10941 , w_10942 , w_10943 , w_10944 , w_10945 , 
		w_10946 , w_10947 , w_10948 , w_10949 , w_10950 , w_10951 , w_10952 , w_10953 , w_10954 , w_10955 , 
		w_10956 , w_10957 , w_10958 , w_10959 , w_10960 , w_10961 , w_10962 , w_10963 , w_10964 , w_10965 , 
		w_10966 , w_10967 , w_10968 , w_10969 , w_10970 , w_10971 , w_10972 , w_10973 , w_10974 , w_10975 , 
		w_10976 , w_10977 , w_10978 , w_10979 , w_10980 , w_10981 , w_10982 , w_10983 , w_10984 , w_10985 , 
		w_10986 , w_10987 , w_10988 , w_10989 , w_10990 , w_10991 , w_10992 , w_10993 , w_10994 , w_10995 , 
		w_10996 , w_10997 , w_10998 , w_10999 , w_11000 , w_11001 , w_11002 , w_11003 , w_11004 , w_11005 , 
		w_11006 , w_11007 , w_11008 , w_11009 , w_11010 , w_11011 , w_11012 , w_11013 , w_11014 , w_11015 , 
		w_11016 , w_11017 , w_11018 , w_11019 , w_11020 , w_11021 , w_11022 , w_11023 , w_11024 , w_11025 , 
		w_11026 , w_11027 , w_11028 , w_11029 , w_11030 , w_11031 , w_11032 , w_11033 , w_11034 , w_11035 , 
		w_11036 , w_11037 , w_11038 , w_11039 , w_11040 , w_11041 , w_11042 , w_11043 , w_11044 , w_11045 , 
		w_11046 , w_11047 , w_11048 , w_11049 , w_11050 , w_11051 , w_11052 , w_11053 , w_11054 , w_11055 , 
		w_11056 , w_11057 , w_11058 , w_11059 , w_11060 , w_11061 , w_11062 , w_11063 , w_11064 , w_11065 , 
		w_11066 , w_11067 , w_11068 , w_11069 , w_11070 , w_11071 , w_11072 , w_11073 , w_11074 , w_11075 , 
		w_11076 , w_11077 , w_11078 , w_11079 , w_11080 , w_11081 , w_11082 , w_11083 , w_11084 , w_11085 , 
		w_11086 , w_11087 , w_11088 , w_11089 , w_11090 , w_11091 , w_11092 , w_11093 , w_11094 , w_11095 , 
		w_11096 , w_11097 , w_11098 , w_11099 , w_11100 , w_11101 , w_11102 , w_11103 , w_11104 , w_11105 , 
		w_11106 , w_11107 , w_11108 , w_11109 , w_11110 , w_11111 , w_11112 , w_11113 , w_11114 , w_11115 , 
		w_11116 , w_11117 , w_11118 , w_11119 , w_11120 , w_11121 , w_11122 , w_11123 , w_11124 , w_11125 , 
		w_11126 , w_11127 , w_11128 , w_11129 , w_11130 , w_11131 , w_11132 , w_11133 , w_11134 , w_11135 , 
		w_11136 , w_11137 , w_11138 , w_11139 , w_11140 , w_11141 , w_11142 , w_11143 , w_11144 , w_11145 , 
		w_11146 , w_11147 , w_11148 , w_11149 , w_11150 , w_11151 , w_11152 , w_11153 , w_11154 , w_11155 , 
		w_11156 , w_11157 , w_11158 , w_11159 , w_11160 , w_11161 , w_11162 , w_11163 , w_11164 , w_11165 , 
		w_11166 , w_11167 , w_11168 , w_11169 , w_11170 , w_11171 , w_11172 , w_11173 , w_11174 , w_11175 , 
		w_11176 , w_11177 , w_11178 , w_11179 , w_11180 , w_11181 , w_11182 , w_11183 , w_11184 , w_11185 , 
		w_11186 , w_11187 , w_11188 , w_11189 , w_11190 , w_11191 , w_11192 , w_11193 , w_11194 , w_11195 , 
		w_11196 , w_11197 , w_11198 , w_11199 , w_11200 , w_11201 , w_11202 , w_11203 , w_11204 , w_11205 , 
		w_11206 , w_11207 , w_11208 , w_11209 , w_11210 , w_11211 , w_11212 , w_11213 , w_11214 , w_11215 , 
		w_11216 , w_11217 , w_11218 , w_11219 , w_11220 , w_11221 , w_11222 , w_11223 , w_11224 , w_11225 , 
		w_11226 , w_11227 , w_11228 , w_11229 , w_11230 , w_11231 , w_11232 , w_11233 , w_11234 , w_11235 , 
		w_11236 , w_11237 , w_11238 , w_11239 , w_11240 , w_11241 , w_11242 , w_11243 , w_11244 , w_11245 , 
		w_11246 , w_11247 , w_11248 , w_11249 , w_11250 , w_11251 , w_11252 , w_11253 , w_11254 , w_11255 , 
		w_11256 , w_11257 , w_11258 , w_11259 , w_11260 , w_11261 , w_11262 , w_11263 , w_11264 , w_11265 , 
		w_11266 , w_11267 , w_11268 , w_11269 , w_11270 , w_11271 , w_11272 , w_11273 , w_11274 , w_11275 , 
		w_11276 , w_11277 , w_11278 , w_11279 , w_11280 , w_11281 , w_11282 , w_11283 , w_11284 , w_11285 , 
		w_11286 , w_11287 , w_11288 , w_11289 , w_11290 , w_11291 , w_11292 , w_11293 , w_11294 , w_11295 , 
		w_11296 , w_11297 , w_11298 , w_11299 , w_11300 , w_11301 , w_11302 , w_11303 , w_11304 , w_11305 , 
		w_11306 , w_11307 , w_11308 , w_11309 , w_11310 , w_11311 , w_11312 , w_11313 , w_11314 , w_11315 , 
		w_11316 , w_11317 , w_11318 , w_11319 , w_11320 , w_11321 , w_11322 , w_11323 , w_11324 , w_11325 , 
		w_11326 , w_11327 , w_11328 , w_11329 , w_11330 , w_11331 , w_11332 , w_11333 , w_11334 , w_11335 , 
		w_11336 , w_11337 , w_11338 , w_11339 , w_11340 , w_11341 , w_11342 , w_11343 , w_11344 , w_11345 , 
		w_11346 , w_11347 , w_11348 , w_11349 , w_11350 , w_11351 , w_11352 , w_11353 , w_11354 , w_11355 , 
		w_11356 , w_11357 , w_11358 , w_11359 , w_11360 , w_11361 , w_11362 , w_11363 , w_11364 , w_11365 , 
		w_11366 , w_11367 , w_11368 , w_11369 , w_11370 , w_11371 , w_11372 , w_11373 , w_11374 , w_11375 , 
		w_11376 , w_11377 , w_11378 , w_11379 , w_11380 , w_11381 , w_11382 , w_11383 , w_11384 , w_11385 , 
		w_11386 , w_11387 , w_11388 , w_11389 , w_11390 , w_11391 , w_11392 , w_11393 , w_11394 , w_11395 , 
		w_11396 , w_11397 , w_11398 , w_11399 , w_11400 , w_11401 , w_11402 , w_11403 , w_11404 , w_11405 , 
		w_11406 , w_11407 , w_11408 , w_11409 , w_11410 , w_11411 , w_11412 , w_11413 , w_11414 , w_11415 , 
		w_11416 , w_11417 , w_11418 , w_11419 , w_11420 , w_11421 , w_11422 , w_11423 , w_11424 , w_11425 , 
		w_11426 , w_11427 , w_11428 , w_11429 , w_11430 , w_11431 , w_11432 , w_11433 , w_11434 , w_11435 , 
		w_11436 , w_11437 , w_11438 , w_11439 , w_11440 , w_11441 , w_11442 , w_11443 , w_11444 , w_11445 , 
		w_11446 , w_11447 , w_11448 , w_11449 , w_11450 , w_11451 , w_11452 , w_11453 , w_11454 , w_11455 , 
		w_11456 , w_11457 , w_11458 , w_11459 , w_11460 , w_11461 , w_11462 , w_11463 , w_11464 , w_11465 , 
		w_11466 , w_11467 , w_11468 , w_11469 , w_11470 , w_11471 , w_11472 , w_11473 , w_11474 , w_11475 , 
		w_11476 , w_11477 , w_11478 , w_11479 , w_11480 , w_11481 , w_11482 , w_11483 , w_11484 , w_11485 , 
		w_11486 , w_11487 , w_11488 , w_11489 , w_11490 , w_11491 , w_11492 , w_11493 , w_11494 , w_11495 , 
		w_11496 , w_11497 , w_11498 , w_11499 , w_11500 , w_11501 , w_11502 , w_11503 , w_11504 , w_11505 , 
		w_11506 , w_11507 , w_11508 , w_11509 , w_11510 , w_11511 , w_11512 , w_11513 , w_11514 , w_11515 , 
		w_11516 , w_11517 , w_11518 , w_11519 , w_11520 , w_11521 , w_11522 , w_11523 , w_11524 , w_11525 , 
		w_11526 , w_11527 , w_11528 , w_11529 , w_11530 , w_11531 , w_11532 , w_11533 , w_11534 , w_11535 , 
		w_11536 , w_11537 , w_11538 , w_11539 , w_11540 , w_11541 , w_11542 , w_11543 , w_11544 , w_11545 , 
		w_11546 , w_11547 , w_11548 , w_11549 , w_11550 , w_11551 , w_11552 , w_11553 , w_11554 , w_11555 , 
		w_11556 , w_11557 , w_11558 , w_11559 , w_11560 , w_11561 , w_11562 , w_11563 , w_11564 , w_11565 , 
		w_11566 , w_11567 , w_11568 , w_11569 , w_11570 , w_11571 , w_11572 , w_11573 , w_11574 , w_11575 , 
		w_11576 , w_11577 , w_11578 , w_11579 , w_11580 , w_11581 , w_11582 , w_11583 , w_11584 , w_11585 , 
		w_11586 , w_11587 , w_11588 , w_11589 , w_11590 , w_11591 , w_11592 , w_11593 , w_11594 , w_11595 , 
		w_11596 , w_11597 , w_11598 , w_11599 , w_11600 , w_11601 , w_11602 , w_11603 , w_11604 , w_11605 , 
		w_11606 , w_11607 , w_11608 , w_11609 , w_11610 , w_11611 , w_11612 , w_11613 , w_11614 , w_11615 , 
		w_11616 , w_11617 , w_11618 , w_11619 , w_11620 , w_11621 , w_11622 , w_11623 , w_11624 , w_11625 , 
		w_11626 , w_11627 , w_11628 , w_11629 , w_11630 , w_11631 , w_11632 , w_11633 , w_11634 , w_11635 , 
		w_11636 , w_11637 , w_11638 , w_11639 , w_11640 , w_11641 , w_11642 , w_11643 , w_11644 , w_11645 , 
		w_11646 , w_11647 , w_11648 , w_11649 , w_11650 , w_11651 , w_11652 , w_11653 , w_11654 , w_11655 , 
		w_11656 , w_11657 , w_11658 , w_11659 , w_11660 , w_11661 , w_11662 , w_11663 , w_11664 , w_11665 , 
		w_11666 , w_11667 , w_11668 , w_11669 , w_11670 , w_11671 , w_11672 , w_11673 , w_11674 , w_11675 , 
		w_11676 , w_11677 , w_11678 , w_11679 , w_11680 , w_11681 , w_11682 , w_11683 , w_11684 , w_11685 , 
		w_11686 , w_11687 , w_11688 , w_11689 , w_11690 , w_11691 , w_11692 , w_11693 , w_11694 , w_11695 , 
		w_11696 , w_11697 , w_11698 , w_11699 , w_11700 , w_11701 , w_11702 , w_11703 , w_11704 , w_11705 , 
		w_11706 , w_11707 , w_11708 , w_11709 , w_11710 , w_11711 , w_11712 , w_11713 , w_11714 , w_11715 , 
		w_11716 , w_11717 , w_11718 , w_11719 , w_11720 , w_11721 , w_11722 , w_11723 , w_11724 , w_11725 , 
		w_11726 , w_11727 , w_11728 , w_11729 , w_11730 , w_11731 , w_11732 , w_11733 , w_11734 , w_11735 , 
		w_11736 , w_11737 , w_11738 , w_11739 , w_11740 , w_11741 , w_11742 , w_11743 , w_11744 , w_11745 , 
		w_11746 , w_11747 , w_11748 , w_11749 , w_11750 , w_11751 , w_11752 , w_11753 , w_11754 , w_11755 , 
		w_11756 , w_11757 , w_11758 , w_11759 , w_11760 , w_11761 , w_11762 , w_11763 , w_11764 , w_11765 , 
		w_11766 , w_11767 , w_11768 , w_11769 , w_11770 , w_11771 , w_11772 , w_11773 , w_11774 , w_11775 , 
		w_11776 , w_11777 , w_11778 , w_11779 , w_11780 , w_11781 , w_11782 , w_11783 , w_11784 , w_11785 , 
		w_11786 , w_11787 , w_11788 , w_11789 , w_11790 , w_11791 , w_11792 , w_11793 , w_11794 , w_11795 , 
		w_11796 , w_11797 , w_11798 , w_11799 , w_11800 , w_11801 , w_11802 , w_11803 , w_11804 , w_11805 , 
		w_11806 , w_11807 , w_11808 , w_11809 , w_11810 , w_11811 , w_11812 , w_11813 , w_11814 , w_11815 , 
		w_11816 , w_11817 , w_11818 , w_11819 , w_11820 , w_11821 , w_11822 , w_11823 , w_11824 , w_11825 , 
		w_11826 , w_11827 , w_11828 , w_11829 , w_11830 , w_11831 , w_11832 , w_11833 , w_11834 , w_11835 , 
		w_11836 , w_11837 , w_11838 , w_11839 , w_11840 , w_11841 , w_11842 , w_11843 , w_11844 , w_11845 , 
		w_11846 , w_11847 , w_11848 , w_11849 , w_11850 , w_11851 , w_11852 , w_11853 , w_11854 , w_11855 , 
		w_11856 , w_11857 , w_11858 , w_11859 , w_11860 , w_11861 , w_11862 , w_11863 , w_11864 , w_11865 , 
		w_11866 , w_11867 , w_11868 , w_11869 , w_11870 , w_11871 , w_11872 , w_11873 , w_11874 , w_11875 , 
		w_11876 , w_11877 , w_11878 , w_11879 , w_11880 , w_11881 , w_11882 , w_11883 , w_11884 , w_11885 , 
		w_11886 , w_11887 , w_11888 , w_11889 , w_11890 , w_11891 , w_11892 , w_11893 , w_11894 , w_11895 , 
		w_11896 , w_11897 , w_11898 , w_11899 , w_11900 , w_11901 , w_11902 , w_11903 , w_11904 , w_11905 , 
		w_11906 , w_11907 , w_11908 , w_11909 , w_11910 , w_11911 , w_11912 , w_11913 , w_11914 , w_11915 , 
		w_11916 , w_11917 , w_11918 , w_11919 , w_11920 , w_11921 , w_11922 , w_11923 , w_11924 , w_11925 , 
		w_11926 , w_11927 , w_11928 , w_11929 , w_11930 , w_11931 , w_11932 , w_11933 , w_11934 , w_11935 , 
		w_11936 , w_11937 , w_11938 , w_11939 , w_11940 , w_11941 , w_11942 , w_11943 , w_11944 , w_11945 , 
		w_11946 , w_11947 , w_11948 , w_11949 , w_11950 , w_11951 , w_11952 , w_11953 , w_11954 , w_11955 , 
		w_11956 , w_11957 , w_11958 , w_11959 , w_11960 , w_11961 , w_11962 , w_11963 , w_11964 , w_11965 , 
		w_11966 , w_11967 , w_11968 , w_11969 , w_11970 , w_11971 , w_11972 , w_11973 , w_11974 , w_11975 , 
		w_11976 , w_11977 , w_11978 , w_11979 , w_11980 , w_11981 , w_11982 , w_11983 , w_11984 , w_11985 , 
		w_11986 , w_11987 , w_11988 , w_11989 , w_11990 , w_11991 , w_11992 , w_11993 , w_11994 , w_11995 , 
		w_11996 , w_11997 , w_11998 , w_11999 , w_12000 , w_12001 , w_12002 , w_12003 , w_12004 , w_12005 , 
		w_12006 , w_12007 , w_12008 , w_12009 , w_12010 , w_12011 , w_12012 , w_12013 , w_12014 , w_12015 , 
		w_12016 , w_12017 , w_12018 , w_12019 , w_12020 , w_12021 , w_12022 , w_12023 , w_12024 , w_12025 , 
		w_12026 , w_12027 , w_12028 , w_12029 , w_12030 , w_12031 , w_12032 , w_12033 , w_12034 , w_12035 , 
		w_12036 , w_12037 , w_12038 , w_12039 , w_12040 , w_12041 , w_12042 , w_12043 , w_12044 , w_12045 , 
		w_12046 , w_12047 , w_12048 , w_12049 , w_12050 , w_12051 , w_12052 , w_12053 , w_12054 , w_12055 , 
		w_12056 , w_12057 , w_12058 , w_12059 , w_12060 , w_12061 , w_12062 , w_12063 , w_12064 , w_12065 , 
		w_12066 , w_12067 , w_12068 , w_12069 , w_12070 , w_12071 , w_12072 , w_12073 , w_12074 , w_12075 , 
		w_12076 , w_12077 , w_12078 , w_12079 , w_12080 , w_12081 , w_12082 , w_12083 , w_12084 , w_12085 , 
		w_12086 , w_12087 , w_12088 , w_12089 , w_12090 , w_12091 , w_12092 , w_12093 , w_12094 , w_12095 , 
		w_12096 , w_12097 , w_12098 , w_12099 , w_12100 , w_12101 , w_12102 , w_12103 , w_12104 , w_12105 , 
		w_12106 , w_12107 , w_12108 , w_12109 , w_12110 , w_12111 , w_12112 , w_12113 , w_12114 , w_12115 , 
		w_12116 , w_12117 , w_12118 , w_12119 , w_12120 , w_12121 , w_12122 , w_12123 , w_12124 , w_12125 , 
		w_12126 , w_12127 , w_12128 , w_12129 , w_12130 , w_12131 , w_12132 , w_12133 , w_12134 , w_12135 , 
		w_12136 , w_12137 , w_12138 , w_12139 , w_12140 , w_12141 , w_12142 , w_12143 , w_12144 , w_12145 , 
		w_12146 , w_12147 , w_12148 , w_12149 , w_12150 , w_12151 , w_12152 , w_12153 , w_12154 , w_12155 , 
		w_12156 , w_12157 , w_12158 , w_12159 , w_12160 , w_12161 , w_12162 , w_12163 , w_12164 , w_12165 , 
		w_12166 , w_12167 , w_12168 , w_12169 , w_12170 , w_12171 , w_12172 , w_12173 , w_12174 , w_12175 , 
		w_12176 , w_12177 , w_12178 , w_12179 , w_12180 , w_12181 , w_12182 , w_12183 , w_12184 , w_12185 , 
		w_12186 , w_12187 , w_12188 , w_12189 , w_12190 , w_12191 , w_12192 , w_12193 , w_12194 , w_12195 , 
		w_12196 , w_12197 , w_12198 , w_12199 , w_12200 , w_12201 , w_12202 , w_12203 , w_12204 , w_12205 , 
		w_12206 , w_12207 , w_12208 , w_12209 , w_12210 , w_12211 , w_12212 , w_12213 , w_12214 , w_12215 , 
		w_12216 , w_12217 , w_12218 , w_12219 , w_12220 , w_12221 , w_12222 , w_12223 , w_12224 , w_12225 , 
		w_12226 , w_12227 , w_12228 , w_12229 , w_12230 , w_12231 , w_12232 , w_12233 , w_12234 , w_12235 , 
		w_12236 , w_12237 , w_12238 , w_12239 , w_12240 , w_12241 , w_12242 , w_12243 , w_12244 , w_12245 , 
		w_12246 , w_12247 , w_12248 , w_12249 , w_12250 , w_12251 , w_12252 , w_12253 , w_12254 , w_12255 , 
		w_12256 , w_12257 , w_12258 , w_12259 , w_12260 , w_12261 , w_12262 , w_12263 , w_12264 , w_12265 , 
		w_12266 , w_12267 , w_12268 , w_12269 , w_12270 , w_12271 , w_12272 , w_12273 , w_12274 , w_12275 , 
		w_12276 , w_12277 , w_12278 , w_12279 , w_12280 , w_12281 , w_12282 , w_12283 , w_12284 , w_12285 , 
		w_12286 , w_12287 , w_12288 , w_12289 , w_12290 , w_12291 , w_12292 , w_12293 , w_12294 , w_12295 , 
		w_12296 , w_12297 , w_12298 , w_12299 , w_12300 , w_12301 , w_12302 , w_12303 , w_12304 , w_12305 , 
		w_12306 , w_12307 , w_12308 , w_12309 , w_12310 , w_12311 , w_12312 , w_12313 , w_12314 , w_12315 , 
		w_12316 , w_12317 , w_12318 , w_12319 , w_12320 , w_12321 , w_12322 , w_12323 , w_12324 , w_12325 , 
		w_12326 , w_12327 , w_12328 , w_12329 , w_12330 , w_12331 , w_12332 , w_12333 , w_12334 , w_12335 , 
		w_12336 , w_12337 , w_12338 , w_12339 , w_12340 , w_12341 , w_12342 , w_12343 , w_12344 , w_12345 , 
		w_12346 , w_12347 , w_12348 , w_12349 , w_12350 , w_12351 , w_12352 , w_12353 , w_12354 , w_12355 , 
		w_12356 , w_12357 , w_12358 , w_12359 , w_12360 , w_12361 , w_12362 , w_12363 , w_12364 , w_12365 , 
		w_12366 , w_12367 , w_12368 , w_12369 , w_12370 , w_12371 , w_12372 , w_12373 , w_12374 , w_12375 , 
		w_12376 , w_12377 , w_12378 , w_12379 , w_12380 , w_12381 , w_12382 , w_12383 , w_12384 , w_12385 , 
		w_12386 , w_12387 , w_12388 , w_12389 , w_12390 , w_12391 , w_12392 , w_12393 , w_12394 , w_12395 , 
		w_12396 , w_12397 , w_12398 , w_12399 , w_12400 , w_12401 , w_12402 , w_12403 , w_12404 , w_12405 , 
		w_12406 , w_12407 , w_12408 , w_12409 , w_12410 , w_12411 , w_12412 , w_12413 , w_12414 , w_12415 , 
		w_12416 , w_12417 , w_12418 , w_12419 , w_12420 , w_12421 , w_12422 , w_12423 , w_12424 , w_12425 , 
		w_12426 , w_12427 , w_12428 , w_12429 , w_12430 , w_12431 , w_12432 , w_12433 , w_12434 , w_12435 , 
		w_12436 , w_12437 , w_12438 , w_12439 , w_12440 , w_12441 , w_12442 , w_12443 , w_12444 , w_12445 , 
		w_12446 , w_12447 , w_12448 , w_12449 , w_12450 , w_12451 , w_12452 , w_12453 , w_12454 , w_12455 , 
		w_12456 , w_12457 , w_12458 , w_12459 , w_12460 , w_12461 , w_12462 , w_12463 , w_12464 , w_12465 , 
		w_12466 , w_12467 , w_12468 , w_12469 , w_12470 , w_12471 , w_12472 , w_12473 , w_12474 , w_12475 , 
		w_12476 , w_12477 , w_12478 , w_12479 , w_12480 , w_12481 , w_12482 , w_12483 , w_12484 , w_12485 , 
		w_12486 , w_12487 , w_12488 , w_12489 , w_12490 , w_12491 , w_12492 , w_12493 , w_12494 , w_12495 , 
		w_12496 , w_12497 , w_12498 , w_12499 , w_12500 , w_12501 , w_12502 , w_12503 , w_12504 , w_12505 , 
		w_12506 , w_12507 , w_12508 , w_12509 , w_12510 , w_12511 , w_12512 , w_12513 , w_12514 , w_12515 , 
		w_12516 , w_12517 , w_12518 , w_12519 , w_12520 , w_12521 , w_12522 , w_12523 , w_12524 , w_12525 , 
		w_12526 , w_12527 , w_12528 , w_12529 , w_12530 , w_12531 , w_12532 , w_12533 , w_12534 , w_12535 , 
		w_12536 , w_12537 , w_12538 , w_12539 , w_12540 , w_12541 , w_12542 , w_12543 , w_12544 , w_12545 , 
		w_12546 , w_12547 , w_12548 , w_12549 , w_12550 , w_12551 , w_12552 , w_12553 , w_12554 , w_12555 , 
		w_12556 , w_12557 , w_12558 , w_12559 , w_12560 , w_12561 , w_12562 , w_12563 , w_12564 , w_12565 , 
		w_12566 , w_12567 , w_12568 , w_12569 , w_12570 , w_12571 , w_12572 , w_12573 , w_12574 , w_12575 , 
		w_12576 , w_12577 , w_12578 , w_12579 , w_12580 , w_12581 , w_12582 , w_12583 , w_12584 , w_12585 , 
		w_12586 , w_12587 , w_12588 , w_12589 , w_12590 , w_12591 , w_12592 , w_12593 , w_12594 , w_12595 , 
		w_12596 , w_12597 , w_12598 , w_12599 , w_12600 , w_12601 , w_12602 , w_12603 , w_12604 , w_12605 , 
		w_12606 , w_12607 , w_12608 , w_12609 , w_12610 , w_12611 , w_12612 , w_12613 , w_12614 , w_12615 , 
		w_12616 , w_12617 , w_12618 , w_12619 , w_12620 , w_12621 , w_12622 , w_12623 , w_12624 , w_12625 , 
		w_12626 , w_12627 , w_12628 , w_12629 , w_12630 , w_12631 , w_12632 , w_12633 , w_12634 , w_12635 , 
		w_12636 , w_12637 , w_12638 , w_12639 , w_12640 , w_12641 , w_12642 , w_12643 , w_12644 , w_12645 , 
		w_12646 , w_12647 , w_12648 , w_12649 , w_12650 , w_12651 , w_12652 , w_12653 , w_12654 , w_12655 , 
		w_12656 , w_12657 , w_12658 , w_12659 , w_12660 , w_12661 , w_12662 , w_12663 , w_12664 , w_12665 , 
		w_12666 , w_12667 , w_12668 , w_12669 , w_12670 , w_12671 , w_12672 , w_12673 , w_12674 , w_12675 , 
		w_12676 , w_12677 , w_12678 , w_12679 , w_12680 , w_12681 , w_12682 , w_12683 , w_12684 , w_12685 , 
		w_12686 , w_12687 , w_12688 , w_12689 , w_12690 , w_12691 , w_12692 , w_12693 , w_12694 , w_12695 , 
		w_12696 , w_12697 , w_12698 , w_12699 , w_12700 , w_12701 , w_12702 , w_12703 , w_12704 , w_12705 , 
		w_12706 , w_12707 , w_12708 , w_12709 , w_12710 , w_12711 , w_12712 , w_12713 , w_12714 , w_12715 , 
		w_12716 , w_12717 , w_12718 , w_12719 , w_12720 , w_12721 , w_12722 , w_12723 , w_12724 , w_12725 , 
		w_12726 , w_12727 , w_12728 , w_12729 , w_12730 , w_12731 , w_12732 , w_12733 , w_12734 , w_12735 , 
		w_12736 , w_12737 , w_12738 , w_12739 , w_12740 , w_12741 , w_12742 , w_12743 , w_12744 , w_12745 , 
		w_12746 , w_12747 , w_12748 , w_12749 , w_12750 , w_12751 , w_12752 , w_12753 , w_12754 , w_12755 , 
		w_12756 , w_12757 , w_12758 , w_12759 , w_12760 , w_12761 , w_12762 , w_12763 , w_12764 , w_12765 , 
		w_12766 , w_12767 , w_12768 , w_12769 , w_12770 , w_12771 , w_12772 , w_12773 , w_12774 , w_12775 , 
		w_12776 , w_12777 , w_12778 , w_12779 , w_12780 , w_12781 , w_12782 , w_12783 , w_12784 , w_12785 , 
		w_12786 , w_12787 , w_12788 , w_12789 , w_12790 , w_12791 , w_12792 , w_12793 , w_12794 , w_12795 , 
		w_12796 , w_12797 , w_12798 , w_12799 , w_12800 , w_12801 , w_12802 , w_12803 , w_12804 , w_12805 , 
		w_12806 , w_12807 , w_12808 , w_12809 , w_12810 , w_12811 , w_12812 , w_12813 , w_12814 , w_12815 , 
		w_12816 , w_12817 , w_12818 , w_12819 , w_12820 , w_12821 , w_12822 , w_12823 , w_12824 , w_12825 , 
		w_12826 , w_12827 , w_12828 , w_12829 , w_12830 , w_12831 , w_12832 , w_12833 , w_12834 , w_12835 , 
		w_12836 , w_12837 , w_12838 , w_12839 , w_12840 , w_12841 , w_12842 , w_12843 , w_12844 , w_12845 , 
		w_12846 , w_12847 , w_12848 , w_12849 , w_12850 , w_12851 , w_12852 , w_12853 , w_12854 , w_12855 , 
		w_12856 , w_12857 , w_12858 , w_12859 , w_12860 , w_12861 , w_12862 , w_12863 , w_12864 , w_12865 , 
		w_12866 , w_12867 , w_12868 , w_12869 , w_12870 , w_12871 , w_12872 , w_12873 , w_12874 , w_12875 , 
		w_12876 , w_12877 , w_12878 , w_12879 , w_12880 , w_12881 , w_12882 , w_12883 , w_12884 , w_12885 , 
		w_12886 , w_12887 , w_12888 , w_12889 , w_12890 , w_12891 , w_12892 , w_12893 , w_12894 , w_12895 , 
		w_12896 , w_12897 , w_12898 , w_12899 , w_12900 , w_12901 , w_12902 , w_12903 , w_12904 , w_12905 , 
		w_12906 , w_12907 , w_12908 , w_12909 , w_12910 , w_12911 , w_12912 , w_12913 , w_12914 , w_12915 , 
		w_12916 , w_12917 , w_12918 , w_12919 , w_12920 , w_12921 , w_12922 , w_12923 , w_12924 , w_12925 , 
		w_12926 , w_12927 , w_12928 , w_12929 , w_12930 , w_12931 , w_12932 , w_12933 , w_12934 , w_12935 , 
		w_12936 , w_12937 , w_12938 , w_12939 , w_12940 , w_12941 , w_12942 , w_12943 , w_12944 , w_12945 , 
		w_12946 , w_12947 , w_12948 , w_12949 , w_12950 , w_12951 , w_12952 , w_12953 , w_12954 , w_12955 , 
		w_12956 , w_12957 , w_12958 , w_12959 , w_12960 , w_12961 , w_12962 , w_12963 , w_12964 , w_12965 , 
		w_12966 , w_12967 , w_12968 , w_12969 , w_12970 , w_12971 , w_12972 , w_12973 , w_12974 , w_12975 , 
		w_12976 , w_12977 , w_12978 , w_12979 , w_12980 , w_12981 , w_12982 , w_12983 , w_12984 , w_12985 , 
		w_12986 , w_12987 , w_12988 , w_12989 , w_12990 , w_12991 , w_12992 , w_12993 , w_12994 , w_12995 , 
		w_12996 , w_12997 , w_12998 , w_12999 , w_13000 , w_13001 , w_13002 , w_13003 , w_13004 , w_13005 , 
		w_13006 , w_13007 , w_13008 , w_13009 , w_13010 , w_13011 , w_13012 , w_13013 , w_13014 , w_13015 , 
		w_13016 , w_13017 , w_13018 , w_13019 , w_13020 , w_13021 , w_13022 , w_13023 , w_13024 , w_13025 , 
		w_13026 , w_13027 , w_13028 , w_13029 , w_13030 , w_13031 , w_13032 , w_13033 , w_13034 , w_13035 , 
		w_13036 , w_13037 , w_13038 , w_13039 , w_13040 , w_13041 , w_13042 , w_13043 , w_13044 , w_13045 , 
		w_13046 , w_13047 , w_13048 , w_13049 , w_13050 , w_13051 , w_13052 , w_13053 , w_13054 , w_13055 , 
		w_13056 , w_13057 , w_13058 , w_13059 , w_13060 , w_13061 , w_13062 , w_13063 , w_13064 , w_13065 , 
		w_13066 , w_13067 , w_13068 , w_13069 , w_13070 , w_13071 , w_13072 , w_13073 , w_13074 , w_13075 , 
		w_13076 , w_13077 , w_13078 , w_13079 , w_13080 , w_13081 , w_13082 , w_13083 , w_13084 , w_13085 , 
		w_13086 , w_13087 , w_13088 , w_13089 , w_13090 , w_13091 , w_13092 , w_13093 , w_13094 , w_13095 , 
		w_13096 , w_13097 , w_13098 , w_13099 , w_13100 , w_13101 , w_13102 , w_13103 , w_13104 , w_13105 , 
		w_13106 , w_13107 , w_13108 , w_13109 , w_13110 , w_13111 , w_13112 , w_13113 , w_13114 , w_13115 , 
		w_13116 , w_13117 , w_13118 , w_13119 , w_13120 , w_13121 , w_13122 , w_13123 , w_13124 , w_13125 , 
		w_13126 , w_13127 , w_13128 , w_13129 , w_13130 , w_13131 , w_13132 , w_13133 , w_13134 , w_13135 , 
		w_13136 , w_13137 , w_13138 , w_13139 , w_13140 , w_13141 , w_13142 , w_13143 , w_13144 , w_13145 , 
		w_13146 , w_13147 , w_13148 , w_13149 , w_13150 , w_13151 , w_13152 , w_13153 , w_13154 , w_13155 , 
		w_13156 , w_13157 , w_13158 , w_13159 , w_13160 , w_13161 , w_13162 , w_13163 , w_13164 , w_13165 , 
		w_13166 , w_13167 , w_13168 , w_13169 , w_13170 , w_13171 , w_13172 , w_13173 , w_13174 , w_13175 , 
		w_13176 , w_13177 , w_13178 , w_13179 , w_13180 , w_13181 , w_13182 , w_13183 , w_13184 , w_13185 , 
		w_13186 , w_13187 , w_13188 , w_13189 , w_13190 , w_13191 , w_13192 , w_13193 , w_13194 , w_13195 , 
		w_13196 , w_13197 , w_13198 , w_13199 , w_13200 , w_13201 , w_13202 , w_13203 , w_13204 , w_13205 , 
		w_13206 , w_13207 , w_13208 , w_13209 , w_13210 , w_13211 , w_13212 , w_13213 , w_13214 , w_13215 , 
		w_13216 , w_13217 , w_13218 , w_13219 , w_13220 , w_13221 , w_13222 , w_13223 , w_13224 , w_13225 , 
		w_13226 , w_13227 , w_13228 , w_13229 , w_13230 , w_13231 , w_13232 , w_13233 , w_13234 , w_13235 , 
		w_13236 , w_13237 , w_13238 , w_13239 , w_13240 , w_13241 , w_13242 , w_13243 , w_13244 , w_13245 , 
		w_13246 , w_13247 , w_13248 , w_13249 , w_13250 , w_13251 , w_13252 , w_13253 , w_13254 , w_13255 , 
		w_13256 , w_13257 , w_13258 , w_13259 , w_13260 , w_13261 , w_13262 , w_13263 , w_13264 , w_13265 , 
		w_13266 , w_13267 , w_13268 , w_13269 , w_13270 , w_13271 , w_13272 , w_13273 , w_13274 , w_13275 , 
		w_13276 , w_13277 , w_13278 , w_13279 , w_13280 , w_13281 , w_13282 , w_13283 , w_13284 , w_13285 , 
		w_13286 , w_13287 , w_13288 , w_13289 , w_13290 , w_13291 , w_13292 , w_13293 , w_13294 , w_13295 , 
		w_13296 , w_13297 , w_13298 , w_13299 , w_13300 , w_13301 , w_13302 , w_13303 , w_13304 , w_13305 , 
		w_13306 , w_13307 , w_13308 , w_13309 , w_13310 , w_13311 , w_13312 , w_13313 , w_13314 , w_13315 , 
		w_13316 , w_13317 , w_13318 , w_13319 , w_13320 , w_13321 , w_13322 , w_13323 , w_13324 , w_13325 , 
		w_13326 , w_13327 , w_13328 , w_13329 , w_13330 , w_13331 , w_13332 , w_13333 , w_13334 , w_13335 , 
		w_13336 , w_13337 , w_13338 , w_13339 , w_13340 , w_13341 , w_13342 , w_13343 , w_13344 , w_13345 , 
		w_13346 , w_13347 , w_13348 , w_13349 , w_13350 , w_13351 , w_13352 , w_13353 , w_13354 , w_13355 , 
		w_13356 , w_13357 , w_13358 , w_13359 , w_13360 , w_13361 , w_13362 , w_13363 , w_13364 , w_13365 , 
		w_13366 , w_13367 , w_13368 , w_13369 , w_13370 , w_13371 , w_13372 , w_13373 , w_13374 , w_13375 , 
		w_13376 , w_13377 , w_13378 , w_13379 , w_13380 , w_13381 , w_13382 , w_13383 , w_13384 , w_13385 , 
		w_13386 , w_13387 , w_13388 , w_13389 , w_13390 , w_13391 , w_13392 , w_13393 , w_13394 , w_13395 , 
		w_13396 , w_13397 , w_13398 , w_13399 , w_13400 , w_13401 , w_13402 , w_13403 , w_13404 , w_13405 , 
		w_13406 , w_13407 , w_13408 , w_13409 , w_13410 , w_13411 , w_13412 , w_13413 , w_13414 , w_13415 , 
		w_13416 , w_13417 , w_13418 , w_13419 , w_13420 , w_13421 , w_13422 , w_13423 , w_13424 , w_13425 , 
		w_13426 , w_13427 , w_13428 , w_13429 , w_13430 , w_13431 , w_13432 , w_13433 , w_13434 , w_13435 , 
		w_13436 , w_13437 , w_13438 , w_13439 , w_13440 , w_13441 , w_13442 , w_13443 , w_13444 , w_13445 , 
		w_13446 , w_13447 , w_13448 , w_13449 , w_13450 , w_13451 , w_13452 , w_13453 , w_13454 , w_13455 , 
		w_13456 , w_13457 , w_13458 , w_13459 , w_13460 , w_13461 , w_13462 , w_13463 , w_13464 , w_13465 , 
		w_13466 , w_13467 , w_13468 , w_13469 , w_13470 , w_13471 , w_13472 , w_13473 , w_13474 , w_13475 , 
		w_13476 , w_13477 , w_13478 , w_13479 , w_13480 , w_13481 , w_13482 , w_13483 , w_13484 , w_13485 , 
		w_13486 , w_13487 , w_13488 , w_13489 , w_13490 , w_13491 , w_13492 , w_13493 , w_13494 , w_13495 , 
		w_13496 , w_13497 , w_13498 , w_13499 , w_13500 , w_13501 , w_13502 , w_13503 , w_13504 , w_13505 , 
		w_13506 , w_13507 , w_13508 , w_13509 , w_13510 , w_13511 , w_13512 , w_13513 , w_13514 , w_13515 , 
		w_13516 , w_13517 , w_13518 , w_13519 , w_13520 , w_13521 , w_13522 , w_13523 , w_13524 , w_13525 , 
		w_13526 , w_13527 , w_13528 , w_13529 , w_13530 , w_13531 , w_13532 , w_13533 , w_13534 , w_13535 , 
		w_13536 , w_13537 , w_13538 , w_13539 , w_13540 , w_13541 , w_13542 , w_13543 , w_13544 , w_13545 , 
		w_13546 , w_13547 , w_13548 , w_13549 , w_13550 , w_13551 , w_13552 , w_13553 , w_13554 , w_13555 , 
		w_13556 , w_13557 , w_13558 , w_13559 , w_13560 , w_13561 , w_13562 , w_13563 , w_13564 , w_13565 , 
		w_13566 , w_13567 , w_13568 , w_13569 , w_13570 , w_13571 , w_13572 , w_13573 , w_13574 , w_13575 , 
		w_13576 , w_13577 , w_13578 , w_13579 , w_13580 , w_13581 , w_13582 , w_13583 , w_13584 , w_13585 , 
		w_13586 , w_13587 , w_13588 , w_13589 , w_13590 , w_13591 , w_13592 , w_13593 , w_13594 , w_13595 , 
		w_13596 , w_13597 , w_13598 , w_13599 , w_13600 , w_13601 , w_13602 , w_13603 , w_13604 , w_13605 , 
		w_13606 , w_13607 , w_13608 , w_13609 , w_13610 , w_13611 , w_13612 , w_13613 , w_13614 , w_13615 , 
		w_13616 , w_13617 , w_13618 , w_13619 , w_13620 , w_13621 , w_13622 , w_13623 , w_13624 , w_13625 , 
		w_13626 , w_13627 , w_13628 , w_13629 , w_13630 , w_13631 , w_13632 , w_13633 , w_13634 , w_13635 , 
		w_13636 , w_13637 , w_13638 , w_13639 , w_13640 , w_13641 , w_13642 , w_13643 , w_13644 , w_13645 , 
		w_13646 , w_13647 , w_13648 , w_13649 , w_13650 , w_13651 , w_13652 , w_13653 , w_13654 , w_13655 , 
		w_13656 , w_13657 , w_13658 , w_13659 , w_13660 , w_13661 , w_13662 , w_13663 , w_13664 , w_13665 , 
		w_13666 , w_13667 , w_13668 , w_13669 , w_13670 , w_13671 , w_13672 , w_13673 , w_13674 , w_13675 , 
		w_13676 , w_13677 , w_13678 , w_13679 , w_13680 , w_13681 , w_13682 , w_13683 , w_13684 , w_13685 , 
		w_13686 , w_13687 , w_13688 , w_13689 , w_13690 , w_13691 , w_13692 , w_13693 , w_13694 , w_13695 , 
		w_13696 , w_13697 , w_13698 , w_13699 , w_13700 , w_13701 , w_13702 , w_13703 , w_13704 , w_13705 , 
		w_13706 , w_13707 , w_13708 , w_13709 , w_13710 , w_13711 , w_13712 , w_13713 , w_13714 , w_13715 , 
		w_13716 , w_13717 , w_13718 , w_13719 , w_13720 , w_13721 , w_13722 , w_13723 , w_13724 , w_13725 , 
		w_13726 , w_13727 , w_13728 , w_13729 , w_13730 , w_13731 , w_13732 , w_13733 , w_13734 , w_13735 , 
		w_13736 , w_13737 , w_13738 , w_13739 , w_13740 , w_13741 , w_13742 , w_13743 , w_13744 , w_13745 , 
		w_13746 , w_13747 , w_13748 , w_13749 , w_13750 , w_13751 , w_13752 , w_13753 , w_13754 , w_13755 , 
		w_13756 , w_13757 , w_13758 , w_13759 , w_13760 , w_13761 , w_13762 , w_13763 , w_13764 , w_13765 , 
		w_13766 , w_13767 , w_13768 , w_13769 , w_13770 , w_13771 , w_13772 , w_13773 , w_13774 , w_13775 , 
		w_13776 , w_13777 , w_13778 , w_13779 , w_13780 , w_13781 , w_13782 , w_13783 , w_13784 , w_13785 , 
		w_13786 , w_13787 , w_13788 , w_13789 , w_13790 , w_13791 , w_13792 , w_13793 , w_13794 , w_13795 , 
		w_13796 , w_13797 , w_13798 , w_13799 , w_13800 , w_13801 , w_13802 , w_13803 , w_13804 , w_13805 , 
		w_13806 , w_13807 , w_13808 , w_13809 , w_13810 , w_13811 , w_13812 , w_13813 , w_13814 , w_13815 , 
		w_13816 , w_13817 , w_13818 , w_13819 , w_13820 , w_13821 , w_13822 , w_13823 , w_13824 , w_13825 , 
		w_13826 , w_13827 , w_13828 , w_13829 , w_13830 , w_13831 , w_13832 , w_13833 , w_13834 , w_13835 , 
		w_13836 , w_13837 , w_13838 , w_13839 , w_13840 , w_13841 , w_13842 , w_13843 , w_13844 , w_13845 , 
		w_13846 , w_13847 , w_13848 , w_13849 , w_13850 , w_13851 , w_13852 , w_13853 , w_13854 , w_13855 , 
		w_13856 , w_13857 , w_13858 , w_13859 , w_13860 , w_13861 , w_13862 , w_13863 , w_13864 , w_13865 , 
		w_13866 , w_13867 , w_13868 , w_13869 , w_13870 , w_13871 , w_13872 , w_13873 , w_13874 , w_13875 , 
		w_13876 , w_13877 , w_13878 , w_13879 , w_13880 , w_13881 , w_13882 , w_13883 , w_13884 , w_13885 , 
		w_13886 , w_13887 , w_13888 , w_13889 , w_13890 , w_13891 , w_13892 , w_13893 , w_13894 , w_13895 , 
		w_13896 , w_13897 , w_13898 , w_13899 , w_13900 , w_13901 , w_13902 , w_13903 , w_13904 , w_13905 , 
		w_13906 , w_13907 , w_13908 , w_13909 , w_13910 , w_13911 , w_13912 , w_13913 , w_13914 , w_13915 , 
		w_13916 , w_13917 , w_13918 , w_13919 , w_13920 , w_13921 , w_13922 , w_13923 , w_13924 , w_13925 , 
		w_13926 , w_13927 , w_13928 , w_13929 , w_13930 , w_13931 , w_13932 , w_13933 , w_13934 , w_13935 , 
		w_13936 , w_13937 , w_13938 , w_13939 , w_13940 , w_13941 , w_13942 , w_13943 , w_13944 , w_13945 , 
		w_13946 , w_13947 , w_13948 , w_13949 , w_13950 , w_13951 , w_13952 , w_13953 , w_13954 , w_13955 , 
		w_13956 , w_13957 , w_13958 , w_13959 , w_13960 , w_13961 , w_13962 , w_13963 , w_13964 , w_13965 , 
		w_13966 , w_13967 , w_13968 , w_13969 , w_13970 , w_13971 , w_13972 , w_13973 , w_13974 , w_13975 , 
		w_13976 , w_13977 , w_13978 , w_13979 , w_13980 , w_13981 , w_13982 , w_13983 , w_13984 , w_13985 , 
		w_13986 , w_13987 , w_13988 , w_13989 , w_13990 , w_13991 , w_13992 , w_13993 , w_13994 , w_13995 , 
		w_13996 , w_13997 , w_13998 , w_13999 , w_14000 , w_14001 , w_14002 , w_14003 , w_14004 , w_14005 , 
		w_14006 , w_14007 , w_14008 , w_14009 , w_14010 , w_14011 , w_14012 , w_14013 , w_14014 , w_14015 , 
		w_14016 , w_14017 , w_14018 , w_14019 , w_14020 , w_14021 , w_14022 , w_14023 , w_14024 , w_14025 , 
		w_14026 , w_14027 , w_14028 , w_14029 , w_14030 , w_14031 , w_14032 , w_14033 , w_14034 , w_14035 , 
		w_14036 , w_14037 , w_14038 , w_14039 , w_14040 , w_14041 , w_14042 , w_14043 , w_14044 , w_14045 , 
		w_14046 , w_14047 , w_14048 , w_14049 , w_14050 , w_14051 , w_14052 , w_14053 , w_14054 , w_14055 , 
		w_14056 , w_14057 , w_14058 , w_14059 , w_14060 , w_14061 , w_14062 , w_14063 , w_14064 , w_14065 , 
		w_14066 , w_14067 , w_14068 , w_14069 , w_14070 , w_14071 , w_14072 , w_14073 , w_14074 , w_14075 , 
		w_14076 , w_14077 , w_14078 , w_14079 , w_14080 , w_14081 , w_14082 , w_14083 , w_14084 , w_14085 , 
		w_14086 , w_14087 , w_14088 , w_14089 , w_14090 , w_14091 , w_14092 , w_14093 , w_14094 , w_14095 , 
		w_14096 , w_14097 , w_14098 , w_14099 , w_14100 , w_14101 , w_14102 , w_14103 , w_14104 , w_14105 , 
		w_14106 , w_14107 , w_14108 , w_14109 , w_14110 , w_14111 , w_14112 , w_14113 , w_14114 , w_14115 , 
		w_14116 , w_14117 , w_14118 , w_14119 , w_14120 , w_14121 , w_14122 , w_14123 , w_14124 , w_14125 , 
		w_14126 , w_14127 , w_14128 , w_14129 , w_14130 , w_14131 , w_14132 , w_14133 , w_14134 , w_14135 , 
		w_14136 , w_14137 , w_14138 , w_14139 , w_14140 , w_14141 , w_14142 , w_14143 , w_14144 , w_14145 , 
		w_14146 , w_14147 , w_14148 , w_14149 , w_14150 , w_14151 , w_14152 , w_14153 , w_14154 , w_14155 , 
		w_14156 , w_14157 , w_14158 , w_14159 , w_14160 , w_14161 , w_14162 , w_14163 , w_14164 , w_14165 , 
		w_14166 , w_14167 , w_14168 , w_14169 , w_14170 , w_14171 , w_14172 , w_14173 , w_14174 , w_14175 , 
		w_14176 , w_14177 , w_14178 , w_14179 , w_14180 , w_14181 , w_14182 , w_14183 , w_14184 , w_14185 , 
		w_14186 , w_14187 , w_14188 , w_14189 , w_14190 , w_14191 , w_14192 , w_14193 , w_14194 , w_14195 , 
		w_14196 , w_14197 , w_14198 , w_14199 , w_14200 , w_14201 , w_14202 , w_14203 , w_14204 , w_14205 , 
		w_14206 , w_14207 , w_14208 , w_14209 , w_14210 , w_14211 , w_14212 , w_14213 , w_14214 , w_14215 , 
		w_14216 , w_14217 , w_14218 , w_14219 , w_14220 , w_14221 , w_14222 , w_14223 , w_14224 , w_14225 , 
		w_14226 , w_14227 , w_14228 , w_14229 , w_14230 , w_14231 , w_14232 , w_14233 , w_14234 , w_14235 , 
		w_14236 , w_14237 , w_14238 , w_14239 , w_14240 , w_14241 , w_14242 , w_14243 , w_14244 , w_14245 , 
		w_14246 , w_14247 , w_14248 , w_14249 , w_14250 , w_14251 , w_14252 , w_14253 , w_14254 , w_14255 , 
		w_14256 , w_14257 , w_14258 , w_14259 , w_14260 , w_14261 , w_14262 , w_14263 , w_14264 , w_14265 , 
		w_14266 , w_14267 , w_14268 , w_14269 , w_14270 , w_14271 , w_14272 , w_14273 , w_14274 , w_14275 , 
		w_14276 , w_14277 , w_14278 , w_14279 , w_14280 , w_14281 , w_14282 , w_14283 , w_14284 , w_14285 , 
		w_14286 , w_14287 , w_14288 , w_14289 , w_14290 , w_14291 , w_14292 , w_14293 , w_14294 , w_14295 , 
		w_14296 , w_14297 , w_14298 , w_14299 , w_14300 , w_14301 , w_14302 , w_14303 , w_14304 , w_14305 , 
		w_14306 , w_14307 , w_14308 , w_14309 , w_14310 , w_14311 , w_14312 , w_14313 , w_14314 , w_14315 , 
		w_14316 , w_14317 , w_14318 , w_14319 , w_14320 , w_14321 , w_14322 , w_14323 , w_14324 , w_14325 , 
		w_14326 , w_14327 , w_14328 , w_14329 , w_14330 , w_14331 , w_14332 , w_14333 , w_14334 , w_14335 , 
		w_14336 , w_14337 , w_14338 , w_14339 , w_14340 , w_14341 , w_14342 , w_14343 , w_14344 , w_14345 , 
		w_14346 , w_14347 , w_14348 , w_14349 , w_14350 , w_14351 , w_14352 , w_14353 , w_14354 , w_14355 , 
		w_14356 , w_14357 , w_14358 , w_14359 , w_14360 , w_14361 , w_14362 , w_14363 , w_14364 , w_14365 , 
		w_14366 , w_14367 , w_14368 , w_14369 , w_14370 , w_14371 , w_14372 , w_14373 , w_14374 , w_14375 , 
		w_14376 , w_14377 , w_14378 , w_14379 , w_14380 , w_14381 , w_14382 , w_14383 , w_14384 , w_14385 , 
		w_14386 , w_14387 , w_14388 , w_14389 , w_14390 , w_14391 , w_14392 , w_14393 , w_14394 , w_14395 , 
		w_14396 , w_14397 , w_14398 , w_14399 , w_14400 , w_14401 , w_14402 , w_14403 , w_14404 , w_14405 , 
		w_14406 , w_14407 , w_14408 , w_14409 , w_14410 , w_14411 , w_14412 , w_14413 , w_14414 , w_14415 , 
		w_14416 , w_14417 , w_14418 , w_14419 , w_14420 , w_14421 , w_14422 , w_14423 , w_14424 , w_14425 , 
		w_14426 , w_14427 , w_14428 , w_14429 , w_14430 , w_14431 , w_14432 , w_14433 , w_14434 , w_14435 , 
		w_14436 , w_14437 , w_14438 , w_14439 , w_14440 , w_14441 , w_14442 , w_14443 , w_14444 , w_14445 , 
		w_14446 , w_14447 , w_14448 , w_14449 , w_14450 , w_14451 , w_14452 , w_14453 , w_14454 , w_14455 , 
		w_14456 , w_14457 , w_14458 , w_14459 , w_14460 , w_14461 , w_14462 , w_14463 , w_14464 , w_14465 , 
		w_14466 , w_14467 , w_14468 , w_14469 , w_14470 , w_14471 , w_14472 , w_14473 , w_14474 , w_14475 , 
		w_14476 , w_14477 , w_14478 , w_14479 , w_14480 , w_14481 , w_14482 , w_14483 , w_14484 , w_14485 , 
		w_14486 , w_14487 , w_14488 , w_14489 , w_14490 , w_14491 , w_14492 , w_14493 , w_14494 , w_14495 , 
		w_14496 , w_14497 , w_14498 , w_14499 , w_14500 , w_14501 , w_14502 , w_14503 , w_14504 , w_14505 , 
		w_14506 , w_14507 , w_14508 , w_14509 , w_14510 , w_14511 , w_14512 , w_14513 , w_14514 , w_14515 , 
		w_14516 , w_14517 , w_14518 , w_14519 , w_14520 , w_14521 , w_14522 , w_14523 , w_14524 , w_14525 , 
		w_14526 , w_14527 , w_14528 , w_14529 , w_14530 , w_14531 , w_14532 , w_14533 , w_14534 , w_14535 , 
		w_14536 , w_14537 , w_14538 , w_14539 , w_14540 , w_14541 , w_14542 , w_14543 , w_14544 , w_14545 , 
		w_14546 , w_14547 , w_14548 , w_14549 , w_14550 , w_14551 , w_14552 , w_14553 , w_14554 , w_14555 , 
		w_14556 , w_14557 , w_14558 , w_14559 , w_14560 , w_14561 , w_14562 , w_14563 , w_14564 , w_14565 , 
		w_14566 , w_14567 , w_14568 , w_14569 , w_14570 , w_14571 , w_14572 , w_14573 , w_14574 , w_14575 , 
		w_14576 , w_14577 , w_14578 , w_14579 , w_14580 , w_14581 , w_14582 , w_14583 , w_14584 , w_14585 , 
		w_14586 , w_14587 , w_14588 , w_14589 , w_14590 , w_14591 , w_14592 , w_14593 , w_14594 , w_14595 , 
		w_14596 , w_14597 , w_14598 , w_14599 , w_14600 , w_14601 , w_14602 , w_14603 , w_14604 , w_14605 , 
		w_14606 , w_14607 , w_14608 , w_14609 , w_14610 , w_14611 , w_14612 , w_14613 , w_14614 , w_14615 , 
		w_14616 , w_14617 , w_14618 , w_14619 , w_14620 , w_14621 , w_14622 , w_14623 , w_14624 , w_14625 , 
		w_14626 , w_14627 , w_14628 , w_14629 , w_14630 , w_14631 , w_14632 , w_14633 , w_14634 , w_14635 , 
		w_14636 , w_14637 , w_14638 , w_14639 , w_14640 , w_14641 , w_14642 , w_14643 , w_14644 , w_14645 , 
		w_14646 , w_14647 , w_14648 , w_14649 , w_14650 , w_14651 , w_14652 , w_14653 , w_14654 , w_14655 , 
		w_14656 , w_14657 , w_14658 , w_14659 , w_14660 , w_14661 , w_14662 , w_14663 , w_14664 , w_14665 , 
		w_14666 , w_14667 , w_14668 , w_14669 , w_14670 , w_14671 , w_14672 , w_14673 , w_14674 , w_14675 , 
		w_14676 , w_14677 , w_14678 , w_14679 , w_14680 , w_14681 , w_14682 , w_14683 , w_14684 , w_14685 , 
		w_14686 , w_14687 , w_14688 , w_14689 , w_14690 , w_14691 , w_14692 , w_14693 , w_14694 , w_14695 , 
		w_14696 , w_14697 , w_14698 , w_14699 , w_14700 , w_14701 , w_14702 , w_14703 , w_14704 , w_14705 , 
		w_14706 , w_14707 , w_14708 , w_14709 , w_14710 , w_14711 , w_14712 , w_14713 , w_14714 , w_14715 , 
		w_14716 , w_14717 , w_14718 , w_14719 , w_14720 , w_14721 , w_14722 , w_14723 , w_14724 , w_14725 , 
		w_14726 , w_14727 , w_14728 , w_14729 , w_14730 , w_14731 , w_14732 , w_14733 , w_14734 , w_14735 , 
		w_14736 , w_14737 , w_14738 , w_14739 , w_14740 , w_14741 , w_14742 , w_14743 , w_14744 , w_14745 , 
		w_14746 , w_14747 , w_14748 , w_14749 , w_14750 , w_14751 , w_14752 , w_14753 , w_14754 , w_14755 , 
		w_14756 , w_14757 , w_14758 , w_14759 , w_14760 , w_14761 , w_14762 , w_14763 , w_14764 , w_14765 , 
		w_14766 , w_14767 , w_14768 , w_14769 , w_14770 , w_14771 , w_14772 , w_14773 , w_14774 , w_14775 , 
		w_14776 , w_14777 , w_14778 , w_14779 , w_14780 , w_14781 , w_14782 , w_14783 , w_14784 , w_14785 , 
		w_14786 , w_14787 , w_14788 , w_14789 , w_14790 , w_14791 , w_14792 , w_14793 , w_14794 , w_14795 , 
		w_14796 , w_14797 , w_14798 , w_14799 , w_14800 , w_14801 , w_14802 , w_14803 , w_14804 , w_14805 , 
		w_14806 , w_14807 , w_14808 , w_14809 , w_14810 , w_14811 , w_14812 , w_14813 , w_14814 , w_14815 , 
		w_14816 , w_14817 , w_14818 , w_14819 , w_14820 , w_14821 , w_14822 , w_14823 , w_14824 , w_14825 , 
		w_14826 , w_14827 , w_14828 , w_14829 , w_14830 , w_14831 , w_14832 , w_14833 , w_14834 , w_14835 , 
		w_14836 , w_14837 , w_14838 , w_14839 , w_14840 , w_14841 , w_14842 , w_14843 , w_14844 , w_14845 , 
		w_14846 , w_14847 , w_14848 , w_14849 , w_14850 , w_14851 , w_14852 , w_14853 , w_14854 , w_14855 , 
		w_14856 , w_14857 , w_14858 , w_14859 , w_14860 , w_14861 , w_14862 , w_14863 , w_14864 , w_14865 , 
		w_14866 , w_14867 , w_14868 , w_14869 , w_14870 , w_14871 , w_14872 , w_14873 , w_14874 , w_14875 , 
		w_14876 , w_14877 , w_14878 , w_14879 , w_14880 , w_14881 , w_14882 , w_14883 , w_14884 , w_14885 , 
		w_14886 , w_14887 , w_14888 , w_14889 , w_14890 , w_14891 , w_14892 , w_14893 , w_14894 , w_14895 , 
		w_14896 , w_14897 , w_14898 , w_14899 , w_14900 , w_14901 , w_14902 , w_14903 , w_14904 , w_14905 , 
		w_14906 , w_14907 , w_14908 , w_14909 , w_14910 , w_14911 , w_14912 , w_14913 , w_14914 , w_14915 , 
		w_14916 , w_14917 , w_14918 , w_14919 , w_14920 , w_14921 , w_14922 , w_14923 , w_14924 , w_14925 , 
		w_14926 , w_14927 , w_14928 , w_14929 , w_14930 , w_14931 , w_14932 , w_14933 , w_14934 , w_14935 , 
		w_14936 , w_14937 , w_14938 , w_14939 , w_14940 , w_14941 , w_14942 , w_14943 , w_14944 , w_14945 , 
		w_14946 , w_14947 , w_14948 , w_14949 , w_14950 , w_14951 , w_14952 , w_14953 , w_14954 , w_14955 , 
		w_14956 , w_14957 , w_14958 , w_14959 , w_14960 , w_14961 , w_14962 , w_14963 , w_14964 , w_14965 , 
		w_14966 , w_14967 , w_14968 , w_14969 , w_14970 , w_14971 , w_14972 , w_14973 , w_14974 , w_14975 , 
		w_14976 , w_14977 , w_14978 , w_14979 , w_14980 , w_14981 , w_14982 , w_14983 , w_14984 , w_14985 , 
		w_14986 , w_14987 , w_14988 , w_14989 , w_14990 , w_14991 , w_14992 , w_14993 , w_14994 , w_14995 , 
		w_14996 , w_14997 , w_14998 , w_14999 , w_15000 , w_15001 , w_15002 , w_15003 , w_15004 , w_15005 , 
		w_15006 , w_15007 , w_15008 , w_15009 , w_15010 , w_15011 , w_15012 , w_15013 , w_15014 , w_15015 , 
		w_15016 , w_15017 , w_15018 , w_15019 , w_15020 , w_15021 , w_15022 , w_15023 , w_15024 , w_15025 , 
		w_15026 , w_15027 , w_15028 , w_15029 , w_15030 , w_15031 , w_15032 , w_15033 , w_15034 , w_15035 , 
		w_15036 , w_15037 , w_15038 , w_15039 , w_15040 , w_15041 , w_15042 , w_15043 , w_15044 , w_15045 , 
		w_15046 , w_15047 , w_15048 , w_15049 , w_15050 , w_15051 , w_15052 , w_15053 , w_15054 , w_15055 , 
		w_15056 , w_15057 , w_15058 , w_15059 , w_15060 , w_15061 , w_15062 , w_15063 , w_15064 , w_15065 , 
		w_15066 , w_15067 , w_15068 , w_15069 , w_15070 , w_15071 , w_15072 , w_15073 , w_15074 , w_15075 , 
		w_15076 , w_15077 , w_15078 , w_15079 , w_15080 , w_15081 , w_15082 , w_15083 , w_15084 , w_15085 , 
		w_15086 , w_15087 , w_15088 , w_15089 , w_15090 , w_15091 , w_15092 , w_15093 , w_15094 , w_15095 , 
		w_15096 , w_15097 , w_15098 , w_15099 , w_15100 , w_15101 , w_15102 , w_15103 , w_15104 , w_15105 , 
		w_15106 , w_15107 , w_15108 , w_15109 , w_15110 , w_15111 , w_15112 , w_15113 , w_15114 , w_15115 , 
		w_15116 , w_15117 , w_15118 , w_15119 , w_15120 , w_15121 , w_15122 , w_15123 , w_15124 , w_15125 , 
		w_15126 , w_15127 , w_15128 , w_15129 , w_15130 , w_15131 , w_15132 , w_15133 , w_15134 , w_15135 , 
		w_15136 , w_15137 , w_15138 , w_15139 , w_15140 , w_15141 , w_15142 , w_15143 , w_15144 , w_15145 , 
		w_15146 , w_15147 , w_15148 , w_15149 , w_15150 , w_15151 , w_15152 , w_15153 , w_15154 , w_15155 , 
		w_15156 , w_15157 , w_15158 , w_15159 , w_15160 , w_15161 , w_15162 , w_15163 , w_15164 , w_15165 , 
		w_15166 , w_15167 , w_15168 , w_15169 , w_15170 , w_15171 , w_15172 , w_15173 , w_15174 , w_15175 , 
		w_15176 , w_15177 , w_15178 , w_15179 , w_15180 , w_15181 , w_15182 , w_15183 , w_15184 , w_15185 , 
		w_15186 , w_15187 , w_15188 , w_15189 , w_15190 , w_15191 , w_15192 , w_15193 , w_15194 , w_15195 , 
		w_15196 , w_15197 , w_15198 , w_15199 , w_15200 , w_15201 , w_15202 , w_15203 , w_15204 , w_15205 , 
		w_15206 , w_15207 , w_15208 , w_15209 , w_15210 , w_15211 , w_15212 , w_15213 , w_15214 , w_15215 , 
		w_15216 , w_15217 , w_15218 , w_15219 , w_15220 , w_15221 , w_15222 , w_15223 , w_15224 , w_15225 , 
		w_15226 , w_15227 , w_15228 , w_15229 , w_15230 , w_15231 , w_15232 , w_15233 , w_15234 , w_15235 , 
		w_15236 , w_15237 , w_15238 , w_15239 , w_15240 , w_15241 , w_15242 , w_15243 , w_15244 , w_15245 , 
		w_15246 , w_15247 , w_15248 , w_15249 , w_15250 , w_15251 , w_15252 , w_15253 , w_15254 , w_15255 , 
		w_15256 , w_15257 , w_15258 , w_15259 , w_15260 , w_15261 , w_15262 , w_15263 , w_15264 , w_15265 , 
		w_15266 , w_15267 , w_15268 , w_15269 , w_15270 , w_15271 , w_15272 , w_15273 , w_15274 , w_15275 , 
		w_15276 , w_15277 , w_15278 , w_15279 , w_15280 , w_15281 , w_15282 , w_15283 , w_15284 , w_15285 , 
		w_15286 , w_15287 , w_15288 , w_15289 , w_15290 , w_15291 , w_15292 , w_15293 , w_15294 , w_15295 , 
		w_15296 , w_15297 , w_15298 , w_15299 , w_15300 , w_15301 , w_15302 , w_15303 , w_15304 , w_15305 , 
		w_15306 , w_15307 , w_15308 , w_15309 , w_15310 , w_15311 , w_15312 , w_15313 , w_15314 , w_15315 , 
		w_15316 , w_15317 , w_15318 , w_15319 , w_15320 , w_15321 , w_15322 , w_15323 , w_15324 , w_15325 , 
		w_15326 , w_15327 , w_15328 , w_15329 , w_15330 , w_15331 , w_15332 , w_15333 , w_15334 , w_15335 , 
		w_15336 , w_15337 , w_15338 , w_15339 , w_15340 , w_15341 , w_15342 , w_15343 , w_15344 , w_15345 , 
		w_15346 , w_15347 , w_15348 , w_15349 , w_15350 , w_15351 , w_15352 , w_15353 , w_15354 , w_15355 , 
		w_15356 , w_15357 , w_15358 , w_15359 , w_15360 , w_15361 , w_15362 , w_15363 , w_15364 , w_15365 , 
		w_15366 , w_15367 , w_15368 , w_15369 , w_15370 , w_15371 , w_15372 , w_15373 , w_15374 , w_15375 , 
		w_15376 , w_15377 , w_15378 , w_15379 , w_15380 , w_15381 , w_15382 , w_15383 , w_15384 , w_15385 , 
		w_15386 , w_15387 , w_15388 , w_15389 , w_15390 , w_15391 , w_15392 , w_15393 , w_15394 , w_15395 , 
		w_15396 , w_15397 , w_15398 , w_15399 , w_15400 , w_15401 , w_15402 , w_15403 , w_15404 , w_15405 , 
		w_15406 , w_15407 , w_15408 , w_15409 , w_15410 , w_15411 , w_15412 , w_15413 , w_15414 , w_15415 , 
		w_15416 , w_15417 , w_15418 , w_15419 , w_15420 , w_15421 , w_15422 , w_15423 , w_15424 , w_15425 , 
		w_15426 , w_15427 , w_15428 , w_15429 , w_15430 , w_15431 , w_15432 , w_15433 , w_15434 , w_15435 , 
		w_15436 , w_15437 , w_15438 , w_15439 , w_15440 , w_15441 , w_15442 , w_15443 , w_15444 , w_15445 , 
		w_15446 , w_15447 , w_15448 , w_15449 , w_15450 , w_15451 , w_15452 , w_15453 , w_15454 , w_15455 , 
		w_15456 , w_15457 , w_15458 , w_15459 , w_15460 , w_15461 , w_15462 , w_15463 , w_15464 , w_15465 , 
		w_15466 , w_15467 , w_15468 , w_15469 , w_15470 , w_15471 , w_15472 , w_15473 , w_15474 , w_15475 , 
		w_15476 , w_15477 , w_15478 , w_15479 , w_15480 , w_15481 , w_15482 , w_15483 , w_15484 , w_15485 , 
		w_15486 , w_15487 , w_15488 , w_15489 , w_15490 , w_15491 , w_15492 , w_15493 , w_15494 , w_15495 , 
		w_15496 , w_15497 , w_15498 , w_15499 , w_15500 , w_15501 , w_15502 , w_15503 , w_15504 , w_15505 , 
		w_15506 , w_15507 , w_15508 , w_15509 , w_15510 , w_15511 , w_15512 , w_15513 , w_15514 , w_15515 , 
		w_15516 , w_15517 , w_15518 , w_15519 , w_15520 , w_15521 , w_15522 , w_15523 , w_15524 , w_15525 , 
		w_15526 , w_15527 , w_15528 , w_15529 , w_15530 , w_15531 , w_15532 , w_15533 , w_15534 , w_15535 , 
		w_15536 , w_15537 , w_15538 , w_15539 , w_15540 , w_15541 , w_15542 , w_15543 , w_15544 , w_15545 , 
		w_15546 , w_15547 , w_15548 , w_15549 , w_15550 , w_15551 , w_15552 , w_15553 , w_15554 , w_15555 , 
		w_15556 , w_15557 , w_15558 , w_15559 , w_15560 , w_15561 , w_15562 , w_15563 , w_15564 , w_15565 , 
		w_15566 , w_15567 , w_15568 , w_15569 , w_15570 , w_15571 , w_15572 , w_15573 , w_15574 , w_15575 , 
		w_15576 , w_15577 , w_15578 , w_15579 , w_15580 , w_15581 , w_15582 , w_15583 , w_15584 , w_15585 , 
		w_15586 , w_15587 , w_15588 , w_15589 , w_15590 , w_15591 , w_15592 , w_15593 , w_15594 , w_15595 , 
		w_15596 , w_15597 , w_15598 , w_15599 , w_15600 , w_15601 , w_15602 , w_15603 , w_15604 , w_15605 , 
		w_15606 , w_15607 , w_15608 , w_15609 , w_15610 , w_15611 , w_15612 , w_15613 , w_15614 , w_15615 , 
		w_15616 , w_15617 , w_15618 , w_15619 , w_15620 , w_15621 , w_15622 , w_15623 , w_15624 , w_15625 , 
		w_15626 , w_15627 , w_15628 , w_15629 , w_15630 , w_15631 , w_15632 , w_15633 , w_15634 , w_15635 , 
		w_15636 , w_15637 , w_15638 , w_15639 , w_15640 , w_15641 , w_15642 , w_15643 , w_15644 , w_15645 , 
		w_15646 , w_15647 , w_15648 , w_15649 , w_15650 , w_15651 , w_15652 , w_15653 , w_15654 , w_15655 , 
		w_15656 , w_15657 , w_15658 , w_15659 , w_15660 , w_15661 , w_15662 , w_15663 , w_15664 , w_15665 , 
		w_15666 , w_15667 , w_15668 , w_15669 , w_15670 , w_15671 , w_15672 , w_15673 , w_15674 , w_15675 , 
		w_15676 , w_15677 , w_15678 , w_15679 , w_15680 , w_15681 , w_15682 , w_15683 , w_15684 , w_15685 , 
		w_15686 , w_15687 , w_15688 , w_15689 , w_15690 , w_15691 , w_15692 , w_15693 , w_15694 , w_15695 , 
		w_15696 , w_15697 , w_15698 , w_15699 , w_15700 , w_15701 , w_15702 , w_15703 , w_15704 , w_15705 , 
		w_15706 , w_15707 , w_15708 , w_15709 , w_15710 , w_15711 , w_15712 , w_15713 , w_15714 , w_15715 , 
		w_15716 , w_15717 , w_15718 , w_15719 , w_15720 , w_15721 , w_15722 , w_15723 , w_15724 , w_15725 , 
		w_15726 , w_15727 , w_15728 , w_15729 , w_15730 , w_15731 , w_15732 , w_15733 , w_15734 , w_15735 , 
		w_15736 , w_15737 , w_15738 , w_15739 , w_15740 , w_15741 , w_15742 , w_15743 , w_15744 , w_15745 , 
		w_15746 , w_15747 , w_15748 , w_15749 , w_15750 , w_15751 , w_15752 , w_15753 , w_15754 , w_15755 , 
		w_15756 , w_15757 , w_15758 , w_15759 , w_15760 , w_15761 , w_15762 , w_15763 , w_15764 , w_15765 , 
		w_15766 , w_15767 , w_15768 , w_15769 , w_15770 , w_15771 , w_15772 , w_15773 , w_15774 , w_15775 , 
		w_15776 , w_15777 , w_15778 , w_15779 , w_15780 , w_15781 , w_15782 , w_15783 , w_15784 , w_15785 , 
		w_15786 , w_15787 , w_15788 , w_15789 , w_15790 , w_15791 , w_15792 , w_15793 , w_15794 , w_15795 , 
		w_15796 , w_15797 , w_15798 , w_15799 , w_15800 , w_15801 , w_15802 , w_15803 , w_15804 , w_15805 , 
		w_15806 , w_15807 , w_15808 , w_15809 , w_15810 , w_15811 , w_15812 , w_15813 , w_15814 , w_15815 , 
		w_15816 , w_15817 , w_15818 , w_15819 , w_15820 , w_15821 , w_15822 , w_15823 , w_15824 , w_15825 , 
		w_15826 , w_15827 , w_15828 , w_15829 , w_15830 , w_15831 , w_15832 , w_15833 , w_15834 , w_15835 , 
		w_15836 , w_15837 , w_15838 , w_15839 , w_15840 , w_15841 , w_15842 , w_15843 , w_15844 , w_15845 , 
		w_15846 , w_15847 , w_15848 , w_15849 , w_15850 , w_15851 , w_15852 , w_15853 , w_15854 , w_15855 , 
		w_15856 , w_15857 , w_15858 , w_15859 , w_15860 , w_15861 , w_15862 , w_15863 , w_15864 , w_15865 , 
		w_15866 , w_15867 , w_15868 , w_15869 , w_15870 , w_15871 , w_15872 , w_15873 , w_15874 , w_15875 , 
		w_15876 , w_15877 , w_15878 , w_15879 , w_15880 , w_15881 , w_15882 , w_15883 , w_15884 , w_15885 , 
		w_15886 , w_15887 , w_15888 , w_15889 , w_15890 , w_15891 , w_15892 , w_15893 , w_15894 , w_15895 , 
		w_15896 , w_15897 , w_15898 , w_15899 , w_15900 , w_15901 , w_15902 , w_15903 , w_15904 , w_15905 , 
		w_15906 , w_15907 , w_15908 , w_15909 , w_15910 , w_15911 , w_15912 , w_15913 , w_15914 , w_15915 , 
		w_15916 , w_15917 , w_15918 , w_15919 , w_15920 , w_15921 , w_15922 , w_15923 , w_15924 , w_15925 , 
		w_15926 , w_15927 , w_15928 , w_15929 , w_15930 , w_15931 , w_15932 , w_15933 , w_15934 , w_15935 , 
		w_15936 , w_15937 , w_15938 , w_15939 , w_15940 , w_15941 , w_15942 , w_15943 , w_15944 , w_15945 , 
		w_15946 , w_15947 , w_15948 , w_15949 , w_15950 , w_15951 , w_15952 , w_15953 , w_15954 , w_15955 , 
		w_15956 , w_15957 , w_15958 , w_15959 , w_15960 , w_15961 , w_15962 , w_15963 , w_15964 , w_15965 , 
		w_15966 , w_15967 , w_15968 , w_15969 , w_15970 , w_15971 , w_15972 , w_15973 , w_15974 , w_15975 , 
		w_15976 , w_15977 , w_15978 , w_15979 , w_15980 , w_15981 , w_15982 , w_15983 , w_15984 , w_15985 , 
		w_15986 , w_15987 , w_15988 , w_15989 , w_15990 , w_15991 , w_15992 , w_15993 , w_15994 , w_15995 , 
		w_15996 , w_15997 , w_15998 , w_15999 , w_16000 , w_16001 , w_16002 , w_16003 , w_16004 , w_16005 , 
		w_16006 , w_16007 , w_16008 , w_16009 , w_16010 , w_16011 , w_16012 , w_16013 , w_16014 , w_16015 , 
		w_16016 , w_16017 , w_16018 , w_16019 , w_16020 , w_16021 , w_16022 , w_16023 , w_16024 , w_16025 , 
		w_16026 , w_16027 , w_16028 , w_16029 , w_16030 , w_16031 , w_16032 , w_16033 , w_16034 , w_16035 , 
		w_16036 , w_16037 , w_16038 , w_16039 , w_16040 , w_16041 , w_16042 , w_16043 , w_16044 , w_16045 , 
		w_16046 , w_16047 , w_16048 , w_16049 , w_16050 , w_16051 , w_16052 , w_16053 , w_16054 , w_16055 , 
		w_16056 , w_16057 , w_16058 , w_16059 , w_16060 , w_16061 , w_16062 , w_16063 , w_16064 , w_16065 , 
		w_16066 , w_16067 , w_16068 , w_16069 , w_16070 , w_16071 , w_16072 , w_16073 , w_16074 , w_16075 , 
		w_16076 , w_16077 , w_16078 , w_16079 , w_16080 , w_16081 , w_16082 , w_16083 , w_16084 , w_16085 , 
		w_16086 , w_16087 , w_16088 , w_16089 , w_16090 , w_16091 , w_16092 , w_16093 , w_16094 , w_16095 , 
		w_16096 , w_16097 , w_16098 , w_16099 , w_16100 , w_16101 , w_16102 , w_16103 , w_16104 , w_16105 , 
		w_16106 , w_16107 , w_16108 , w_16109 , w_16110 , w_16111 , w_16112 , w_16113 , w_16114 , w_16115 , 
		w_16116 , w_16117 , w_16118 , w_16119 , w_16120 , w_16121 , w_16122 , w_16123 , w_16124 , w_16125 , 
		w_16126 , w_16127 , w_16128 , w_16129 , w_16130 , w_16131 , w_16132 , w_16133 , w_16134 , w_16135 , 
		w_16136 , w_16137 , w_16138 , w_16139 , w_16140 , w_16141 , w_16142 , w_16143 , w_16144 , w_16145 , 
		w_16146 , w_16147 , w_16148 , w_16149 , w_16150 , w_16151 , w_16152 , w_16153 , w_16154 , w_16155 , 
		w_16156 , w_16157 , w_16158 , w_16159 , w_16160 , w_16161 , w_16162 , w_16163 , w_16164 , w_16165 , 
		w_16166 , w_16167 , w_16168 , w_16169 , w_16170 , w_16171 , w_16172 , w_16173 , w_16174 , w_16175 , 
		w_16176 , w_16177 , w_16178 , w_16179 , w_16180 , w_16181 , w_16182 , w_16183 , w_16184 , w_16185 , 
		w_16186 , w_16187 , w_16188 , w_16189 , w_16190 , w_16191 , w_16192 , w_16193 , w_16194 , w_16195 , 
		w_16196 , w_16197 , w_16198 , w_16199 , w_16200 , w_16201 , w_16202 , w_16203 , w_16204 , w_16205 , 
		w_16206 , w_16207 , w_16208 , w_16209 , w_16210 , w_16211 , w_16212 , w_16213 , w_16214 , w_16215 , 
		w_16216 , w_16217 , w_16218 , w_16219 , w_16220 , w_16221 , w_16222 , w_16223 , w_16224 , w_16225 , 
		w_16226 , w_16227 , w_16228 , w_16229 , w_16230 , w_16231 , w_16232 , w_16233 , w_16234 , w_16235 , 
		w_16236 , w_16237 , w_16238 , w_16239 , w_16240 , w_16241 , w_16242 , w_16243 , w_16244 , w_16245 , 
		w_16246 , w_16247 , w_16248 , w_16249 , w_16250 , w_16251 , w_16252 , w_16253 , w_16254 , w_16255 , 
		w_16256 , w_16257 , w_16258 , w_16259 , w_16260 , w_16261 , w_16262 , w_16263 , w_16264 , w_16265 , 
		w_16266 , w_16267 , w_16268 , w_16269 , w_16270 , w_16271 , w_16272 , w_16273 , w_16274 , w_16275 , 
		w_16276 , w_16277 , w_16278 , w_16279 , w_16280 , w_16281 , w_16282 , w_16283 , w_16284 , w_16285 , 
		w_16286 , w_16287 , w_16288 , w_16289 , w_16290 , w_16291 , w_16292 , w_16293 , w_16294 , w_16295 , 
		w_16296 , w_16297 , w_16298 , w_16299 , w_16300 , w_16301 , w_16302 , w_16303 , w_16304 , w_16305 , 
		w_16306 , w_16307 , w_16308 , w_16309 , w_16310 , w_16311 , w_16312 , w_16313 , w_16314 , w_16315 , 
		w_16316 , w_16317 , w_16318 , w_16319 , w_16320 , w_16321 , w_16322 , w_16323 , w_16324 , w_16325 , 
		w_16326 , w_16327 , w_16328 , w_16329 , w_16330 , w_16331 , w_16332 , w_16333 , w_16334 , w_16335 , 
		w_16336 , w_16337 , w_16338 , w_16339 , w_16340 , w_16341 , w_16342 , w_16343 , w_16344 , w_16345 , 
		w_16346 , w_16347 , w_16348 , w_16349 , w_16350 , w_16351 , w_16352 , w_16353 , w_16354 , w_16355 , 
		w_16356 , w_16357 , w_16358 , w_16359 , w_16360 , w_16361 , w_16362 , w_16363 , w_16364 , w_16365 , 
		w_16366 , w_16367 , w_16368 , w_16369 , w_16370 , w_16371 , w_16372 , w_16373 , w_16374 , w_16375 , 
		w_16376 , w_16377 , w_16378 , w_16379 , w_16380 , w_16381 , w_16382 , w_16383 , w_16384 , w_16385 , 
		w_16386 , w_16387 , w_16388 , w_16389 , w_16390 , w_16391 , w_16392 , w_16393 , w_16394 , w_16395 , 
		w_16396 , w_16397 , w_16398 , w_16399 , w_16400 , w_16401 , w_16402 , w_16403 , w_16404 , w_16405 , 
		w_16406 , w_16407 , w_16408 , w_16409 , w_16410 , w_16411 , w_16412 , w_16413 , w_16414 , w_16415 , 
		w_16416 , w_16417 , w_16418 , w_16419 , w_16420 , w_16421 , w_16422 , w_16423 , w_16424 , w_16425 , 
		w_16426 , w_16427 , w_16428 , w_16429 , w_16430 , w_16431 , w_16432 , w_16433 , w_16434 , w_16435 , 
		w_16436 , w_16437 , w_16438 , w_16439 , w_16440 , w_16441 , w_16442 , w_16443 , w_16444 , w_16445 , 
		w_16446 , w_16447 , w_16448 , w_16449 , w_16450 , w_16451 , w_16452 , w_16453 , w_16454 , w_16455 , 
		w_16456 , w_16457 , w_16458 , w_16459 , w_16460 , w_16461 , w_16462 , w_16463 , w_16464 , w_16465 , 
		w_16466 , w_16467 , w_16468 , w_16469 , w_16470 , w_16471 , w_16472 , w_16473 , w_16474 , w_16475 , 
		w_16476 , w_16477 , w_16478 , w_16479 , w_16480 , w_16481 , w_16482 , w_16483 , w_16484 , w_16485 , 
		w_16486 , w_16487 , w_16488 , w_16489 , w_16490 , w_16491 , w_16492 , w_16493 , w_16494 , w_16495 , 
		w_16496 , w_16497 , w_16498 , w_16499 , w_16500 , w_16501 , w_16502 , w_16503 , w_16504 , w_16505 , 
		w_16506 , w_16507 , w_16508 , w_16509 , w_16510 , w_16511 , w_16512 , w_16513 , w_16514 , w_16515 , 
		w_16516 , w_16517 , w_16518 , w_16519 , w_16520 , w_16521 , w_16522 , w_16523 , w_16524 , w_16525 , 
		w_16526 , w_16527 , w_16528 , w_16529 , w_16530 , w_16531 , w_16532 , w_16533 , w_16534 , w_16535 , 
		w_16536 , w_16537 , w_16538 , w_16539 , w_16540 , w_16541 , w_16542 , w_16543 , w_16544 , w_16545 , 
		w_16546 , w_16547 , w_16548 , w_16549 , w_16550 , w_16551 , w_16552 , w_16553 , w_16554 , w_16555 , 
		w_16556 , w_16557 , w_16558 , w_16559 , w_16560 , w_16561 , w_16562 , w_16563 , w_16564 , w_16565 , 
		w_16566 , w_16567 , w_16568 , w_16569 , w_16570 , w_16571 , w_16572 , w_16573 , w_16574 , w_16575 , 
		w_16576 , w_16577 , w_16578 , w_16579 , w_16580 , w_16581 , w_16582 , w_16583 , w_16584 , w_16585 , 
		w_16586 , w_16587 , w_16588 , w_16589 , w_16590 , w_16591 , w_16592 , w_16593 , w_16594 , w_16595 , 
		w_16596 , w_16597 , w_16598 , w_16599 , w_16600 , w_16601 , w_16602 , w_16603 , w_16604 , w_16605 , 
		w_16606 , w_16607 , w_16608 , w_16609 , w_16610 , w_16611 , w_16612 , w_16613 , w_16614 , w_16615 , 
		w_16616 , w_16617 , w_16618 , w_16619 , w_16620 , w_16621 , w_16622 , w_16623 , w_16624 , w_16625 , 
		w_16626 , w_16627 , w_16628 , w_16629 , w_16630 , w_16631 , w_16632 , w_16633 , w_16634 , w_16635 , 
		w_16636 , w_16637 , w_16638 , w_16639 , w_16640 , w_16641 , w_16642 , w_16643 , w_16644 , w_16645 , 
		w_16646 , w_16647 , w_16648 , w_16649 , w_16650 , w_16651 , w_16652 , w_16653 , w_16654 , w_16655 , 
		w_16656 , w_16657 , w_16658 , w_16659 , w_16660 , w_16661 , w_16662 , w_16663 , w_16664 , w_16665 , 
		w_16666 , w_16667 , w_16668 , w_16669 , w_16670 , w_16671 , w_16672 , w_16673 , w_16674 , w_16675 , 
		w_16676 , w_16677 , w_16678 , w_16679 , w_16680 , w_16681 , w_16682 , w_16683 , w_16684 , w_16685 , 
		w_16686 , w_16687 , w_16688 , w_16689 , w_16690 , w_16691 , w_16692 , w_16693 , w_16694 , w_16695 , 
		w_16696 , w_16697 , w_16698 , w_16699 , w_16700 , w_16701 , w_16702 , w_16703 , w_16704 , w_16705 , 
		w_16706 , w_16707 , w_16708 , w_16709 , w_16710 , w_16711 , w_16712 , w_16713 , w_16714 , w_16715 , 
		w_16716 , w_16717 , w_16718 , w_16719 , w_16720 , w_16721 , w_16722 , w_16723 , w_16724 , w_16725 , 
		w_16726 , w_16727 , w_16728 , w_16729 , w_16730 , w_16731 , w_16732 , w_16733 , w_16734 , w_16735 , 
		w_16736 , w_16737 , w_16738 , w_16739 , w_16740 , w_16741 , w_16742 , w_16743 , w_16744 , w_16745 , 
		w_16746 , w_16747 , w_16748 , w_16749 , w_16750 , w_16751 , w_16752 , w_16753 , w_16754 , w_16755 , 
		w_16756 , w_16757 , w_16758 , w_16759 , w_16760 , w_16761 , w_16762 , w_16763 , w_16764 , w_16765 , 
		w_16766 , w_16767 , w_16768 , w_16769 , w_16770 , w_16771 , w_16772 , w_16773 , w_16774 , w_16775 , 
		w_16776 , w_16777 , w_16778 , w_16779 , w_16780 , w_16781 , w_16782 , w_16783 , w_16784 , w_16785 , 
		w_16786 , w_16787 , w_16788 , w_16789 , w_16790 , w_16791 , w_16792 , w_16793 , w_16794 , w_16795 , 
		w_16796 , w_16797 , w_16798 , w_16799 , w_16800 , w_16801 , w_16802 , w_16803 , w_16804 , w_16805 , 
		w_16806 , w_16807 , w_16808 , w_16809 , w_16810 , w_16811 , w_16812 , w_16813 , w_16814 , w_16815 , 
		w_16816 , w_16817 , w_16818 , w_16819 , w_16820 , w_16821 , w_16822 , w_16823 , w_16824 , w_16825 , 
		w_16826 , w_16827 , w_16828 , w_16829 , w_16830 , w_16831 , w_16832 , w_16833 , w_16834 , w_16835 , 
		w_16836 , w_16837 , w_16838 , w_16839 , w_16840 , w_16841 , w_16842 , w_16843 , w_16844 , w_16845 , 
		w_16846 , w_16847 , w_16848 , w_16849 , w_16850 , w_16851 , w_16852 , w_16853 , w_16854 , w_16855 , 
		w_16856 , w_16857 , w_16858 , w_16859 , w_16860 , w_16861 , w_16862 , w_16863 , w_16864 , w_16865 , 
		w_16866 , w_16867 , w_16868 , w_16869 , w_16870 , w_16871 , w_16872 , w_16873 , w_16874 , w_16875 , 
		w_16876 , w_16877 , w_16878 , w_16879 , w_16880 , w_16881 , w_16882 , w_16883 , w_16884 , w_16885 , 
		w_16886 , w_16887 , w_16888 , w_16889 , w_16890 , w_16891 , w_16892 , w_16893 , w_16894 , w_16895 , 
		w_16896 , w_16897 , w_16898 , w_16899 , w_16900 , w_16901 , w_16902 , w_16903 , w_16904 , w_16905 , 
		w_16906 , w_16907 , w_16908 , w_16909 , w_16910 , w_16911 , w_16912 , w_16913 , w_16914 , w_16915 , 
		w_16916 , w_16917 , w_16918 , w_16919 , w_16920 , w_16921 , w_16922 , w_16923 , w_16924 , w_16925 , 
		w_16926 , w_16927 , w_16928 , w_16929 , w_16930 , w_16931 , w_16932 , w_16933 , w_16934 , w_16935 , 
		w_16936 , w_16937 , w_16938 , w_16939 , w_16940 , w_16941 , w_16942 , w_16943 , w_16944 , w_16945 , 
		w_16946 , w_16947 , w_16948 , w_16949 , w_16950 , w_16951 , w_16952 , w_16953 , w_16954 , w_16955 , 
		w_16956 , w_16957 , w_16958 , w_16959 , w_16960 , w_16961 , w_16962 , w_16963 , w_16964 , w_16965 , 
		w_16966 , w_16967 , w_16968 , w_16969 , w_16970 , w_16971 , w_16972 , w_16973 , w_16974 , w_16975 , 
		w_16976 , w_16977 , w_16978 , w_16979 , w_16980 , w_16981 , w_16982 , w_16983 , w_16984 , w_16985 , 
		w_16986 , w_16987 , w_16988 , w_16989 , w_16990 , w_16991 , w_16992 , w_16993 , w_16994 , w_16995 , 
		w_16996 , w_16997 , w_16998 , w_16999 , w_17000 , w_17001 , w_17002 , w_17003 , w_17004 , w_17005 , 
		w_17006 , w_17007 , w_17008 , w_17009 , w_17010 , w_17011 , w_17012 , w_17013 , w_17014 , w_17015 , 
		w_17016 , w_17017 , w_17018 , w_17019 , w_17020 , w_17021 , w_17022 , w_17023 , w_17024 , w_17025 , 
		w_17026 , w_17027 , w_17028 , w_17029 , w_17030 , w_17031 , w_17032 , w_17033 , w_17034 , w_17035 , 
		w_17036 , w_17037 , w_17038 , w_17039 , w_17040 , w_17041 , w_17042 , w_17043 , w_17044 , w_17045 , 
		w_17046 , w_17047 , w_17048 , w_17049 , w_17050 , w_17051 , w_17052 , w_17053 , w_17054 , w_17055 , 
		w_17056 , w_17057 , w_17058 , w_17059 , w_17060 , w_17061 , w_17062 , w_17063 , w_17064 , w_17065 , 
		w_17066 , w_17067 , w_17068 , w_17069 , w_17070 , w_17071 , w_17072 , w_17073 , w_17074 , w_17075 , 
		w_17076 , w_17077 , w_17078 , w_17079 , w_17080 , w_17081 , w_17082 , w_17083 , w_17084 , w_17085 , 
		w_17086 , w_17087 , w_17088 , w_17089 , w_17090 , w_17091 , w_17092 , w_17093 , w_17094 , w_17095 , 
		w_17096 , w_17097 , w_17098 , w_17099 , w_17100 , w_17101 , w_17102 , w_17103 , w_17104 , w_17105 , 
		w_17106 , w_17107 , w_17108 , w_17109 , w_17110 , w_17111 , w_17112 , w_17113 , w_17114 , w_17115 , 
		w_17116 , w_17117 , w_17118 , w_17119 , w_17120 , w_17121 , w_17122 , w_17123 , w_17124 , w_17125 , 
		w_17126 , w_17127 , w_17128 , w_17129 , w_17130 , w_17131 , w_17132 , w_17133 , w_17134 , w_17135 , 
		w_17136 , w_17137 , w_17138 , w_17139 , w_17140 , w_17141 , w_17142 , w_17143 , w_17144 , w_17145 , 
		w_17146 , w_17147 , w_17148 , w_17149 , w_17150 , w_17151 , w_17152 , w_17153 , w_17154 , w_17155 , 
		w_17156 , w_17157 , w_17158 , w_17159 , w_17160 , w_17161 , w_17162 , w_17163 , w_17164 , w_17165 , 
		w_17166 , w_17167 , w_17168 , w_17169 , w_17170 , w_17171 , w_17172 , w_17173 , w_17174 , w_17175 , 
		w_17176 , w_17177 , w_17178 , w_17179 , w_17180 , w_17181 , w_17182 , w_17183 , w_17184 , w_17185 , 
		w_17186 , w_17187 , w_17188 , w_17189 , w_17190 , w_17191 , w_17192 , w_17193 , w_17194 , w_17195 , 
		w_17196 , w_17197 , w_17198 , w_17199 , w_17200 , w_17201 , w_17202 , w_17203 , w_17204 , w_17205 , 
		w_17206 , w_17207 , w_17208 , w_17209 , w_17210 , w_17211 , w_17212 , w_17213 , w_17214 , w_17215 , 
		w_17216 , w_17217 , w_17218 , w_17219 , w_17220 , w_17221 , w_17222 , w_17223 , w_17224 , w_17225 , 
		w_17226 , w_17227 , w_17228 , w_17229 , w_17230 , w_17231 , w_17232 , w_17233 , w_17234 , w_17235 , 
		w_17236 , w_17237 , w_17238 , w_17239 , w_17240 , w_17241 , w_17242 , w_17243 , w_17244 , w_17245 , 
		w_17246 , w_17247 , w_17248 , w_17249 , w_17250 , w_17251 , w_17252 , w_17253 , w_17254 , w_17255 , 
		w_17256 , w_17257 , w_17258 , w_17259 , w_17260 , w_17261 , w_17262 , w_17263 , w_17264 , w_17265 , 
		w_17266 , w_17267 , w_17268 , w_17269 , w_17270 , w_17271 , w_17272 , w_17273 , w_17274 , w_17275 , 
		w_17276 , w_17277 , w_17278 , w_17279 , w_17280 , w_17281 , w_17282 , w_17283 , w_17284 , w_17285 , 
		w_17286 , w_17287 , w_17288 , w_17289 , w_17290 , w_17291 , w_17292 , w_17293 , w_17294 , w_17295 , 
		w_17296 , w_17297 , w_17298 , w_17299 , w_17300 , w_17301 , w_17302 , w_17303 , w_17304 , w_17305 , 
		w_17306 , w_17307 , w_17308 , w_17309 , w_17310 , w_17311 , w_17312 , w_17313 , w_17314 , w_17315 , 
		w_17316 , w_17317 , w_17318 , w_17319 , w_17320 , w_17321 , w_17322 , w_17323 , w_17324 , w_17325 , 
		w_17326 , w_17327 , w_17328 , w_17329 , w_17330 , w_17331 , w_17332 , w_17333 , w_17334 , w_17335 , 
		w_17336 , w_17337 , w_17338 , w_17339 , w_17340 , w_17341 , w_17342 , w_17343 , w_17344 , w_17345 , 
		w_17346 , w_17347 , w_17348 , w_17349 , w_17350 , w_17351 , w_17352 , w_17353 , w_17354 , w_17355 , 
		w_17356 , w_17357 , w_17358 , w_17359 , w_17360 , w_17361 , w_17362 , w_17363 , w_17364 , w_17365 , 
		w_17366 , w_17367 , w_17368 , w_17369 , w_17370 , w_17371 , w_17372 , w_17373 , w_17374 , w_17375 , 
		w_17376 , w_17377 , w_17378 , w_17379 , w_17380 , w_17381 , w_17382 , w_17383 , w_17384 , w_17385 , 
		w_17386 , w_17387 , w_17388 , w_17389 , w_17390 , w_17391 , w_17392 , w_17393 , w_17394 , w_17395 , 
		w_17396 , w_17397 , w_17398 , w_17399 , w_17400 , w_17401 , w_17402 , w_17403 , w_17404 , w_17405 , 
		w_17406 , w_17407 , w_17408 , w_17409 , w_17410 , w_17411 , w_17412 , w_17413 , w_17414 , w_17415 , 
		w_17416 , w_17417 , w_17418 , w_17419 , w_17420 , w_17421 , w_17422 , w_17423 , w_17424 , w_17425 , 
		w_17426 , w_17427 , w_17428 , w_17429 , w_17430 , w_17431 , w_17432 , w_17433 , w_17434 , w_17435 , 
		w_17436 , w_17437 , w_17438 , w_17439 , w_17440 , w_17441 , w_17442 , w_17443 , w_17444 , w_17445 , 
		w_17446 , w_17447 , w_17448 , w_17449 , w_17450 , w_17451 , w_17452 , w_17453 , w_17454 , w_17455 , 
		w_17456 , w_17457 , w_17458 , w_17459 , w_17460 , w_17461 , w_17462 , w_17463 , w_17464 , w_17465 , 
		w_17466 , w_17467 , w_17468 , w_17469 , w_17470 , w_17471 , w_17472 , w_17473 , w_17474 , w_17475 , 
		w_17476 , w_17477 , w_17478 , w_17479 , w_17480 , w_17481 , w_17482 , w_17483 , w_17484 , w_17485 , 
		w_17486 , w_17487 , w_17488 , w_17489 , w_17490 , w_17491 , w_17492 , w_17493 , w_17494 , w_17495 , 
		w_17496 , w_17497 , w_17498 , w_17499 , w_17500 , w_17501 , w_17502 , w_17503 , w_17504 , w_17505 , 
		w_17506 , w_17507 , w_17508 , w_17509 , w_17510 , w_17511 , w_17512 , w_17513 , w_17514 , w_17515 , 
		w_17516 , w_17517 , w_17518 , w_17519 , w_17520 , w_17521 , w_17522 , w_17523 , w_17524 , w_17525 , 
		w_17526 , w_17527 , w_17528 , w_17529 , w_17530 , w_17531 , w_17532 , w_17533 , w_17534 , w_17535 , 
		w_17536 , w_17537 , w_17538 , w_17539 , w_17540 , w_17541 , w_17542 , w_17543 , w_17544 , w_17545 , 
		w_17546 , w_17547 , w_17548 , w_17549 , w_17550 , w_17551 , w_17552 , w_17553 , w_17554 , w_17555 , 
		w_17556 , w_17557 , w_17558 , w_17559 , w_17560 , w_17561 , w_17562 , w_17563 , w_17564 , w_17565 , 
		w_17566 , w_17567 , w_17568 , w_17569 , w_17570 , w_17571 , w_17572 , w_17573 , w_17574 , w_17575 , 
		w_17576 , w_17577 , w_17578 , w_17579 , w_17580 , w_17581 , w_17582 , w_17583 , w_17584 , w_17585 , 
		w_17586 , w_17587 , w_17588 , w_17589 , w_17590 , w_17591 , w_17592 , w_17593 , w_17594 , w_17595 , 
		w_17596 , w_17597 , w_17598 , w_17599 , w_17600 , w_17601 , w_17602 , w_17603 , w_17604 , w_17605 , 
		w_17606 , w_17607 , w_17608 , w_17609 , w_17610 , w_17611 , w_17612 , w_17613 , w_17614 , w_17615 , 
		w_17616 , w_17617 , w_17618 , w_17619 , w_17620 , w_17621 , w_17622 , w_17623 , w_17624 , w_17625 , 
		w_17626 , w_17627 , w_17628 , w_17629 , w_17630 , w_17631 , w_17632 , w_17633 , w_17634 , w_17635 , 
		w_17636 , w_17637 , w_17638 , w_17639 , w_17640 , w_17641 , w_17642 , w_17643 , w_17644 , w_17645 , 
		w_17646 , w_17647 , w_17648 , w_17649 , w_17650 , w_17651 , w_17652 , w_17653 , w_17654 , w_17655 , 
		w_17656 , w_17657 , w_17658 , w_17659 , w_17660 , w_17661 , w_17662 , w_17663 , w_17664 , w_17665 , 
		w_17666 , w_17667 , w_17668 , w_17669 , w_17670 , w_17671 , w_17672 , w_17673 , w_17674 , w_17675 , 
		w_17676 , w_17677 , w_17678 , w_17679 , w_17680 , w_17681 , w_17682 , w_17683 , w_17684 , w_17685 , 
		w_17686 , w_17687 , w_17688 , w_17689 , w_17690 , w_17691 , w_17692 , w_17693 , w_17694 , w_17695 , 
		w_17696 , w_17697 , w_17698 , w_17699 , w_17700 , w_17701 , w_17702 , w_17703 , w_17704 , w_17705 , 
		w_17706 , w_17707 , w_17708 , w_17709 , w_17710 , w_17711 , w_17712 , w_17713 , w_17714 , w_17715 , 
		w_17716 , w_17717 , w_17718 , w_17719 , w_17720 , w_17721 , w_17722 , w_17723 , w_17724 , w_17725 , 
		w_17726 , w_17727 , w_17728 , w_17729 , w_17730 , w_17731 , w_17732 , w_17733 , w_17734 , w_17735 , 
		w_17736 , w_17737 , w_17738 , w_17739 , w_17740 , w_17741 , w_17742 , w_17743 , w_17744 , w_17745 , 
		w_17746 , w_17747 , w_17748 , w_17749 , w_17750 , w_17751 , w_17752 , w_17753 , w_17754 , w_17755 , 
		w_17756 , w_17757 , w_17758 , w_17759 , w_17760 , w_17761 , w_17762 , w_17763 , w_17764 , w_17765 , 
		w_17766 , w_17767 , w_17768 , w_17769 , w_17770 , w_17771 , w_17772 , w_17773 , w_17774 , w_17775 , 
		w_17776 , w_17777 , w_17778 , w_17779 , w_17780 , w_17781 , w_17782 , w_17783 , w_17784 , w_17785 , 
		w_17786 , w_17787 , w_17788 , w_17789 , w_17790 , w_17791 , w_17792 , w_17793 , w_17794 , w_17795 , 
		w_17796 , w_17797 , w_17798 , w_17799 , w_17800 , w_17801 , w_17802 , w_17803 , w_17804 , w_17805 , 
		w_17806 , w_17807 , w_17808 , w_17809 , w_17810 , w_17811 , w_17812 , w_17813 , w_17814 , w_17815 , 
		w_17816 , w_17817 , w_17818 , w_17819 , w_17820 , w_17821 , w_17822 , w_17823 , w_17824 , w_17825 , 
		w_17826 , w_17827 , w_17828 , w_17829 , w_17830 , w_17831 , w_17832 , w_17833 , w_17834 , w_17835 , 
		w_17836 , w_17837 , w_17838 , w_17839 , w_17840 , w_17841 , w_17842 , w_17843 , w_17844 , w_17845 , 
		w_17846 , w_17847 , w_17848 , w_17849 , w_17850 , w_17851 , w_17852 , w_17853 , w_17854 , w_17855 , 
		w_17856 , w_17857 , w_17858 , w_17859 , w_17860 , w_17861 , w_17862 , w_17863 , w_17864 , w_17865 , 
		w_17866 , w_17867 , w_17868 , w_17869 , w_17870 , w_17871 , w_17872 , w_17873 , w_17874 , w_17875 , 
		w_17876 , w_17877 , w_17878 , w_17879 , w_17880 , w_17881 , w_17882 , w_17883 , w_17884 , w_17885 , 
		w_17886 , w_17887 , w_17888 , w_17889 , w_17890 , w_17891 , w_17892 , w_17893 , w_17894 , w_17895 , 
		w_17896 , w_17897 , w_17898 , w_17899 , w_17900 , w_17901 , w_17902 , w_17903 , w_17904 , w_17905 , 
		w_17906 , w_17907 , w_17908 , w_17909 , w_17910 , w_17911 , w_17912 , w_17913 , w_17914 , w_17915 , 
		w_17916 , w_17917 , w_17918 , w_17919 , w_17920 , w_17921 , w_17922 , w_17923 , w_17924 , w_17925 , 
		w_17926 , w_17927 , w_17928 , w_17929 , w_17930 , w_17931 , w_17932 , w_17933 , w_17934 , w_17935 , 
		w_17936 , w_17937 , w_17938 , w_17939 , w_17940 , w_17941 , w_17942 , w_17943 , w_17944 , w_17945 , 
		w_17946 , w_17947 , w_17948 , w_17949 , w_17950 , w_17951 , w_17952 , w_17953 , w_17954 , w_17955 , 
		w_17956 , w_17957 , w_17958 , w_17959 , w_17960 , w_17961 , w_17962 , w_17963 , w_17964 , w_17965 , 
		w_17966 , w_17967 , w_17968 , w_17969 , w_17970 , w_17971 , w_17972 , w_17973 , w_17974 , w_17975 , 
		w_17976 , w_17977 , w_17978 , w_17979 , w_17980 , w_17981 , w_17982 , w_17983 , w_17984 , w_17985 , 
		w_17986 , w_17987 , w_17988 , w_17989 , w_17990 , w_17991 , w_17992 , w_17993 , w_17994 , w_17995 , 
		w_17996 , w_17997 , w_17998 , w_17999 , w_18000 , w_18001 , w_18002 , w_18003 , w_18004 , w_18005 , 
		w_18006 , w_18007 , w_18008 , w_18009 , w_18010 , w_18011 , w_18012 , w_18013 , w_18014 , w_18015 , 
		w_18016 , w_18017 , w_18018 , w_18019 , w_18020 , w_18021 , w_18022 , w_18023 , w_18024 , w_18025 , 
		w_18026 , w_18027 , w_18028 , w_18029 , w_18030 , w_18031 , w_18032 , w_18033 , w_18034 , w_18035 , 
		w_18036 , w_18037 , w_18038 , w_18039 , w_18040 , w_18041 , w_18042 , w_18043 , w_18044 , w_18045 , 
		w_18046 , w_18047 , w_18048 , w_18049 , w_18050 , w_18051 , w_18052 , w_18053 , w_18054 , w_18055 , 
		w_18056 , w_18057 , w_18058 , w_18059 , w_18060 , w_18061 , w_18062 , w_18063 , w_18064 , w_18065 , 
		w_18066 , w_18067 , w_18068 , w_18069 , w_18070 , w_18071 , w_18072 , w_18073 , w_18074 , w_18075 , 
		w_18076 , w_18077 , w_18078 , w_18079 , w_18080 , w_18081 , w_18082 , w_18083 , w_18084 , w_18085 , 
		w_18086 , w_18087 , w_18088 , w_18089 , w_18090 , w_18091 , w_18092 , w_18093 , w_18094 , w_18095 , 
		w_18096 , w_18097 , w_18098 , w_18099 , w_18100 , w_18101 , w_18102 , w_18103 , w_18104 , w_18105 , 
		w_18106 , w_18107 , w_18108 , w_18109 , w_18110 , w_18111 , w_18112 , w_18113 , w_18114 , w_18115 , 
		w_18116 , w_18117 , w_18118 , w_18119 , w_18120 , w_18121 , w_18122 , w_18123 , w_18124 , w_18125 , 
		w_18126 , w_18127 , w_18128 , w_18129 , w_18130 , w_18131 , w_18132 , w_18133 , w_18134 , w_18135 , 
		w_18136 , w_18137 , w_18138 , w_18139 , w_18140 , w_18141 , w_18142 , w_18143 , w_18144 , w_18145 , 
		w_18146 , w_18147 , w_18148 , w_18149 , w_18150 , w_18151 , w_18152 , w_18153 , w_18154 , w_18155 , 
		w_18156 , w_18157 , w_18158 , w_18159 , w_18160 , w_18161 , w_18162 , w_18163 , w_18164 , w_18165 , 
		w_18166 , w_18167 , w_18168 , w_18169 , w_18170 , w_18171 , w_18172 , w_18173 , w_18174 , w_18175 , 
		w_18176 , w_18177 , w_18178 , w_18179 , w_18180 , w_18181 , w_18182 , w_18183 , w_18184 , w_18185 , 
		w_18186 , w_18187 , w_18188 , w_18189 , w_18190 , w_18191 , w_18192 , w_18193 , w_18194 , w_18195 , 
		w_18196 , w_18197 , w_18198 , w_18199 , w_18200 , w_18201 , w_18202 , w_18203 , w_18204 , w_18205 , 
		w_18206 , w_18207 , w_18208 , w_18209 , w_18210 , w_18211 , w_18212 , w_18213 , w_18214 , w_18215 , 
		w_18216 , w_18217 , w_18218 , w_18219 , w_18220 , w_18221 , w_18222 , w_18223 , w_18224 , w_18225 , 
		w_18226 , w_18227 , w_18228 , w_18229 , w_18230 , w_18231 , w_18232 , w_18233 , w_18234 , w_18235 , 
		w_18236 , w_18237 , w_18238 , w_18239 , w_18240 , w_18241 , w_18242 , w_18243 , w_18244 , w_18245 , 
		w_18246 , w_18247 , w_18248 , w_18249 , w_18250 , w_18251 , w_18252 , w_18253 , w_18254 , w_18255 , 
		w_18256 , w_18257 , w_18258 , w_18259 , w_18260 , w_18261 , w_18262 , w_18263 , w_18264 , w_18265 , 
		w_18266 , w_18267 , w_18268 , w_18269 , w_18270 , w_18271 , w_18272 , w_18273 , w_18274 , w_18275 , 
		w_18276 , w_18277 , w_18278 , w_18279 , w_18280 , w_18281 , w_18282 , w_18283 , w_18284 , w_18285 , 
		w_18286 , w_18287 , w_18288 , w_18289 , w_18290 , w_18291 , w_18292 , w_18293 , w_18294 , w_18295 , 
		w_18296 , w_18297 , w_18298 , w_18299 , w_18300 , w_18301 , w_18302 , w_18303 , w_18304 , w_18305 , 
		w_18306 , w_18307 , w_18308 , w_18309 , w_18310 , w_18311 , w_18312 , w_18313 , w_18314 , w_18315 , 
		w_18316 , w_18317 , w_18318 , w_18319 , w_18320 , w_18321 , w_18322 , w_18323 , w_18324 , w_18325 , 
		w_18326 , w_18327 , w_18328 , w_18329 , w_18330 , w_18331 , w_18332 , w_18333 , w_18334 , w_18335 , 
		w_18336 , w_18337 , w_18338 , w_18339 , w_18340 , w_18341 , w_18342 , w_18343 , w_18344 , w_18345 , 
		w_18346 , w_18347 , w_18348 , w_18349 , w_18350 , w_18351 , w_18352 , w_18353 , w_18354 , w_18355 , 
		w_18356 , w_18357 , w_18358 , w_18359 , w_18360 , w_18361 , w_18362 , w_18363 , w_18364 , w_18365 , 
		w_18366 , w_18367 , w_18368 , w_18369 , w_18370 , w_18371 , w_18372 , w_18373 , w_18374 , w_18375 , 
		w_18376 , w_18377 , w_18378 , w_18379 , w_18380 , w_18381 , w_18382 , w_18383 , w_18384 , w_18385 , 
		w_18386 , w_18387 , w_18388 , w_18389 , w_18390 , w_18391 , w_18392 , w_18393 , w_18394 , w_18395 , 
		w_18396 , w_18397 , w_18398 , w_18399 , w_18400 , w_18401 , w_18402 , w_18403 , w_18404 , w_18405 , 
		w_18406 , w_18407 , w_18408 , w_18409 , w_18410 , w_18411 , w_18412 , w_18413 , w_18414 , w_18415 , 
		w_18416 , w_18417 , w_18418 , w_18419 , w_18420 , w_18421 , w_18422 , w_18423 , w_18424 , w_18425 , 
		w_18426 , w_18427 , w_18428 , w_18429 , w_18430 , w_18431 , w_18432 , w_18433 , w_18434 , w_18435 , 
		w_18436 , w_18437 , w_18438 , w_18439 , w_18440 , w_18441 , w_18442 , w_18443 , w_18444 , w_18445 , 
		w_18446 , w_18447 , w_18448 , w_18449 , w_18450 , w_18451 , w_18452 , w_18453 , w_18454 , w_18455 , 
		w_18456 , w_18457 , w_18458 , w_18459 , w_18460 , w_18461 , w_18462 , w_18463 , w_18464 , w_18465 , 
		w_18466 , w_18467 , w_18468 , w_18469 , w_18470 , w_18471 , w_18472 , w_18473 , w_18474 , w_18475 , 
		w_18476 , w_18477 , w_18478 , w_18479 , w_18480 , w_18481 , w_18482 , w_18483 , w_18484 , w_18485 , 
		w_18486 , w_18487 , w_18488 , w_18489 , w_18490 , w_18491 , w_18492 , w_18493 , w_18494 , w_18495 , 
		w_18496 , w_18497 , w_18498 , w_18499 , w_18500 , w_18501 , w_18502 , w_18503 , w_18504 , w_18505 , 
		w_18506 , w_18507 , w_18508 , w_18509 , w_18510 , w_18511 , w_18512 , w_18513 , w_18514 , w_18515 , 
		w_18516 , w_18517 , w_18518 , w_18519 , w_18520 , w_18521 , w_18522 , w_18523 , w_18524 , w_18525 , 
		w_18526 , w_18527 , w_18528 , w_18529 , w_18530 , w_18531 , w_18532 , w_18533 , w_18534 , w_18535 , 
		w_18536 , w_18537 , w_18538 , w_18539 , w_18540 , w_18541 , w_18542 , w_18543 , w_18544 , w_18545 , 
		w_18546 , w_18547 , w_18548 , w_18549 , w_18550 , w_18551 , w_18552 , w_18553 , w_18554 , w_18555 , 
		w_18556 , w_18557 , w_18558 , w_18559 , w_18560 , w_18561 , w_18562 , w_18563 , w_18564 , w_18565 , 
		w_18566 , w_18567 , w_18568 , w_18569 , w_18570 , w_18571 , w_18572 , w_18573 , w_18574 , w_18575 , 
		w_18576 , w_18577 , w_18578 , w_18579 , w_18580 , w_18581 , w_18582 , w_18583 , w_18584 , w_18585 , 
		w_18586 , w_18587 , w_18588 , w_18589 , w_18590 , w_18591 , w_18592 , w_18593 , w_18594 , w_18595 , 
		w_18596 , w_18597 , w_18598 , w_18599 , w_18600 , w_18601 , w_18602 , w_18603 , w_18604 , w_18605 , 
		w_18606 , w_18607 , w_18608 , w_18609 , w_18610 , w_18611 , w_18612 , w_18613 , w_18614 , w_18615 , 
		w_18616 , w_18617 , w_18618 , w_18619 , w_18620 , w_18621 , w_18622 , w_18623 , w_18624 , w_18625 , 
		w_18626 , w_18627 , w_18628 , w_18629 , w_18630 , w_18631 , w_18632 , w_18633 , w_18634 , w_18635 , 
		w_18636 , w_18637 , w_18638 , w_18639 , w_18640 , w_18641 , w_18642 , w_18643 , w_18644 , w_18645 , 
		w_18646 , w_18647 , w_18648 , w_18649 , w_18650 , w_18651 , w_18652 , w_18653 , w_18654 , w_18655 , 
		w_18656 , w_18657 , w_18658 , w_18659 , w_18660 , w_18661 , w_18662 , w_18663 , w_18664 , w_18665 , 
		w_18666 , w_18667 , w_18668 , w_18669 , w_18670 , w_18671 , w_18672 , w_18673 , w_18674 , w_18675 , 
		w_18676 , w_18677 , w_18678 , w_18679 , w_18680 , w_18681 , w_18682 , w_18683 , w_18684 , w_18685 , 
		w_18686 , w_18687 , w_18688 , w_18689 , w_18690 , w_18691 , w_18692 , w_18693 , w_18694 , w_18695 , 
		w_18696 , w_18697 , w_18698 , w_18699 , w_18700 , w_18701 , w_18702 , w_18703 , w_18704 , w_18705 , 
		w_18706 , w_18707 , w_18708 , w_18709 , w_18710 , w_18711 , w_18712 , w_18713 , w_18714 , w_18715 , 
		w_18716 , w_18717 , w_18718 , w_18719 , w_18720 , w_18721 , w_18722 , w_18723 , w_18724 , w_18725 , 
		w_18726 , w_18727 , w_18728 , w_18729 , w_18730 , w_18731 , w_18732 , w_18733 , w_18734 , w_18735 , 
		w_18736 , w_18737 , w_18738 , w_18739 , w_18740 , w_18741 , w_18742 , w_18743 , w_18744 , w_18745 , 
		w_18746 , w_18747 , w_18748 , w_18749 , w_18750 , w_18751 , w_18752 , w_18753 , w_18754 , w_18755 , 
		w_18756 , w_18757 , w_18758 , w_18759 , w_18760 , w_18761 , w_18762 , w_18763 , w_18764 , w_18765 , 
		w_18766 , w_18767 , w_18768 , w_18769 , w_18770 , w_18771 , w_18772 , w_18773 , w_18774 , w_18775 , 
		w_18776 , w_18777 , w_18778 , w_18779 , w_18780 , w_18781 , w_18782 , w_18783 , w_18784 , w_18785 , 
		w_18786 , w_18787 , w_18788 , w_18789 , w_18790 , w_18791 , w_18792 , w_18793 , w_18794 , w_18795 , 
		w_18796 , w_18797 , w_18798 , w_18799 , w_18800 , w_18801 , w_18802 , w_18803 , w_18804 , w_18805 , 
		w_18806 , w_18807 , w_18808 , w_18809 , w_18810 , w_18811 , w_18812 , w_18813 , w_18814 , w_18815 , 
		w_18816 , w_18817 , w_18818 , w_18819 , w_18820 , w_18821 , w_18822 , w_18823 , w_18824 , w_18825 , 
		w_18826 , w_18827 , w_18828 , w_18829 , w_18830 , w_18831 , w_18832 , w_18833 , w_18834 , w_18835 , 
		w_18836 , w_18837 , w_18838 , w_18839 , w_18840 , w_18841 , w_18842 , w_18843 , w_18844 , w_18845 , 
		w_18846 , w_18847 , w_18848 , w_18849 , w_18850 , w_18851 , w_18852 , w_18853 , w_18854 , w_18855 , 
		w_18856 , w_18857 , w_18858 , w_18859 , w_18860 , w_18861 , w_18862 , w_18863 , w_18864 , w_18865 , 
		w_18866 , w_18867 , w_18868 , w_18869 , w_18870 , w_18871 , w_18872 , w_18873 , w_18874 , w_18875 , 
		w_18876 , w_18877 , w_18878 , w_18879 , w_18880 , w_18881 , w_18882 , w_18883 , w_18884 , w_18885 , 
		w_18886 , w_18887 , w_18888 , w_18889 , w_18890 , w_18891 , w_18892 , w_18893 , w_18894 , w_18895 , 
		w_18896 , w_18897 , w_18898 , w_18899 , w_18900 , w_18901 , w_18902 , w_18903 , w_18904 , w_18905 , 
		w_18906 , w_18907 , w_18908 , w_18909 , w_18910 , w_18911 , w_18912 , w_18913 , w_18914 , w_18915 , 
		w_18916 , w_18917 , w_18918 , w_18919 , w_18920 , w_18921 , w_18922 , w_18923 , w_18924 , w_18925 , 
		w_18926 , w_18927 , w_18928 , w_18929 , w_18930 , w_18931 , w_18932 , w_18933 , w_18934 , w_18935 , 
		w_18936 , w_18937 , w_18938 , w_18939 , w_18940 , w_18941 , w_18942 , w_18943 , w_18944 , w_18945 , 
		w_18946 , w_18947 , w_18948 , w_18949 , w_18950 , w_18951 , w_18952 , w_18953 , w_18954 , w_18955 , 
		w_18956 , w_18957 , w_18958 , w_18959 , w_18960 , w_18961 , w_18962 , w_18963 , w_18964 , w_18965 , 
		w_18966 , w_18967 , w_18968 , w_18969 , w_18970 , w_18971 , w_18972 , w_18973 , w_18974 , w_18975 , 
		w_18976 , w_18977 , w_18978 , w_18979 , w_18980 , w_18981 , w_18982 , w_18983 , w_18984 , w_18985 , 
		w_18986 , w_18987 , w_18988 , w_18989 , w_18990 , w_18991 , w_18992 , w_18993 , w_18994 , w_18995 , 
		w_18996 , w_18997 , w_18998 , w_18999 , w_19000 , w_19001 , w_19002 , w_19003 , w_19004 , w_19005 , 
		w_19006 , w_19007 , w_19008 , w_19009 , w_19010 , w_19011 , w_19012 , w_19013 , w_19014 , w_19015 , 
		w_19016 , w_19017 , w_19018 , w_19019 , w_19020 , w_19021 , w_19022 , w_19023 , w_19024 , w_19025 , 
		w_19026 , w_19027 , w_19028 , w_19029 , w_19030 , w_19031 , w_19032 , w_19033 , w_19034 , w_19035 , 
		w_19036 , w_19037 , w_19038 , w_19039 , w_19040 , w_19041 , w_19042 , w_19043 , w_19044 , w_19045 , 
		w_19046 , w_19047 , w_19048 , w_19049 , w_19050 , w_19051 , w_19052 , w_19053 , w_19054 , w_19055 , 
		w_19056 , w_19057 , w_19058 , w_19059 , w_19060 , w_19061 , w_19062 , w_19063 , w_19064 , w_19065 , 
		w_19066 , w_19067 , w_19068 , w_19069 , w_19070 , w_19071 , w_19072 , w_19073 , w_19074 , w_19075 , 
		w_19076 , w_19077 , w_19078 , w_19079 , w_19080 , w_19081 , w_19082 , w_19083 , w_19084 , w_19085 , 
		w_19086 , w_19087 , w_19088 , w_19089 , w_19090 , w_19091 , w_19092 , w_19093 , w_19094 , w_19095 , 
		w_19096 , w_19097 , w_19098 , w_19099 , w_19100 , w_19101 , w_19102 , w_19103 , w_19104 , w_19105 , 
		w_19106 , w_19107 , w_19108 , w_19109 , w_19110 , w_19111 , w_19112 , w_19113 , w_19114 , w_19115 , 
		w_19116 , w_19117 , w_19118 , w_19119 , w_19120 , w_19121 , w_19122 , w_19123 , w_19124 , w_19125 , 
		w_19126 , w_19127 , w_19128 , w_19129 , w_19130 , w_19131 , w_19132 , w_19133 , w_19134 , w_19135 , 
		w_19136 , w_19137 , w_19138 , w_19139 , w_19140 , w_19141 , w_19142 , w_19143 , w_19144 , w_19145 , 
		w_19146 , w_19147 , w_19148 , w_19149 , w_19150 , w_19151 , w_19152 , w_19153 , w_19154 , w_19155 , 
		w_19156 , w_19157 , w_19158 , w_19159 , w_19160 , w_19161 , w_19162 , w_19163 , w_19164 , w_19165 , 
		w_19166 , w_19167 , w_19168 , w_19169 , w_19170 , w_19171 , w_19172 , w_19173 , w_19174 , w_19175 , 
		w_19176 , w_19177 , w_19178 , w_19179 , w_19180 , w_19181 , w_19182 , w_19183 , w_19184 , w_19185 , 
		w_19186 , w_19187 , w_19188 , w_19189 , w_19190 , w_19191 , w_19192 , w_19193 , w_19194 , w_19195 , 
		w_19196 , w_19197 , w_19198 , w_19199 , w_19200 , w_19201 , w_19202 , w_19203 , w_19204 , w_19205 , 
		w_19206 , w_19207 , w_19208 , w_19209 , w_19210 , w_19211 , w_19212 , w_19213 , w_19214 , w_19215 , 
		w_19216 , w_19217 , w_19218 , w_19219 , w_19220 , w_19221 , w_19222 , w_19223 , w_19224 , w_19225 , 
		w_19226 , w_19227 , w_19228 , w_19229 , w_19230 , w_19231 , w_19232 , w_19233 , w_19234 , w_19235 , 
		w_19236 , w_19237 , w_19238 , w_19239 , w_19240 , w_19241 , w_19242 , w_19243 , w_19244 , w_19245 , 
		w_19246 , w_19247 , w_19248 , w_19249 , w_19250 , w_19251 , w_19252 , w_19253 , w_19254 , w_19255 , 
		w_19256 , w_19257 , w_19258 , w_19259 , w_19260 , w_19261 , w_19262 , w_19263 , w_19264 , w_19265 , 
		w_19266 , w_19267 , w_19268 , w_19269 , w_19270 , w_19271 , w_19272 , w_19273 , w_19274 , w_19275 , 
		w_19276 , w_19277 , w_19278 , w_19279 , w_19280 , w_19281 , w_19282 , w_19283 , w_19284 , w_19285 , 
		w_19286 , w_19287 , w_19288 , w_19289 , w_19290 , w_19291 , w_19292 , w_19293 , w_19294 , w_19295 , 
		w_19296 , w_19297 , w_19298 , w_19299 , w_19300 , w_19301 , w_19302 , w_19303 , w_19304 , w_19305 , 
		w_19306 , w_19307 , w_19308 , w_19309 , w_19310 , w_19311 , w_19312 , w_19313 , w_19314 , w_19315 , 
		w_19316 , w_19317 , w_19318 , w_19319 , w_19320 , w_19321 , w_19322 , w_19323 , w_19324 , w_19325 , 
		w_19326 , w_19327 , w_19328 , w_19329 , w_19330 , w_19331 , w_19332 , w_19333 , w_19334 , w_19335 , 
		w_19336 , w_19337 , w_19338 , w_19339 , w_19340 , w_19341 , w_19342 , w_19343 , w_19344 , w_19345 , 
		w_19346 , w_19347 , w_19348 , w_19349 , w_19350 , w_19351 , w_19352 , w_19353 , w_19354 , w_19355 , 
		w_19356 , w_19357 , w_19358 , w_19359 , w_19360 , w_19361 , w_19362 , w_19363 , w_19364 , w_19365 , 
		w_19366 , w_19367 , w_19368 , w_19369 , w_19370 , w_19371 , w_19372 , w_19373 , w_19374 , w_19375 , 
		w_19376 , w_19377 , w_19378 , w_19379 , w_19380 , w_19381 , w_19382 , w_19383 , w_19384 , w_19385 , 
		w_19386 , w_19387 , w_19388 , w_19389 , w_19390 , w_19391 , w_19392 , w_19393 , w_19394 , w_19395 , 
		w_19396 , w_19397 , w_19398 , w_19399 , w_19400 , w_19401 , w_19402 , w_19403 , w_19404 , w_19405 , 
		w_19406 , w_19407 , w_19408 , w_19409 , w_19410 , w_19411 , w_19412 , w_19413 , w_19414 , w_19415 , 
		w_19416 , w_19417 , w_19418 , w_19419 , w_19420 , w_19421 , w_19422 , w_19423 , w_19424 , w_19425 , 
		w_19426 , w_19427 , w_19428 , w_19429 , w_19430 , w_19431 , w_19432 , w_19433 , w_19434 , w_19435 , 
		w_19436 , w_19437 , w_19438 , w_19439 , w_19440 , w_19441 , w_19442 , w_19443 , w_19444 , w_19445 , 
		w_19446 , w_19447 , w_19448 , w_19449 , w_19450 , w_19451 , w_19452 , w_19453 , w_19454 , w_19455 , 
		w_19456 , w_19457 , w_19458 , w_19459 , w_19460 , w_19461 , w_19462 , w_19463 , w_19464 , w_19465 , 
		w_19466 , w_19467 , w_19468 , w_19469 , w_19470 , w_19471 , w_19472 , w_19473 , w_19474 , w_19475 , 
		w_19476 , w_19477 , w_19478 , w_19479 , w_19480 , w_19481 , w_19482 , w_19483 , w_19484 , w_19485 , 
		w_19486 , w_19487 , w_19488 , w_19489 , w_19490 , w_19491 , w_19492 , w_19493 , w_19494 , w_19495 , 
		w_19496 , w_19497 , w_19498 , w_19499 , w_19500 , w_19501 , w_19502 , w_19503 , w_19504 , w_19505 , 
		w_19506 , w_19507 , w_19508 , w_19509 , w_19510 , w_19511 , w_19512 , w_19513 , w_19514 , w_19515 , 
		w_19516 , w_19517 , w_19518 , w_19519 , w_19520 , w_19521 , w_19522 , w_19523 , w_19524 , w_19525 , 
		w_19526 , w_19527 , w_19528 , w_19529 , w_19530 , w_19531 , w_19532 , w_19533 , w_19534 , w_19535 , 
		w_19536 , w_19537 , w_19538 , w_19539 , w_19540 , w_19541 , w_19542 , w_19543 , w_19544 , w_19545 , 
		w_19546 , w_19547 , w_19548 , w_19549 , w_19550 , w_19551 , w_19552 , w_19553 , w_19554 , w_19555 , 
		w_19556 , w_19557 , w_19558 , w_19559 , w_19560 , w_19561 , w_19562 , w_19563 , w_19564 , w_19565 , 
		w_19566 , w_19567 , w_19568 , w_19569 , w_19570 , w_19571 , w_19572 , w_19573 , w_19574 , w_19575 , 
		w_19576 , w_19577 , w_19578 , w_19579 , w_19580 , w_19581 , w_19582 , w_19583 , w_19584 , w_19585 , 
		w_19586 , w_19587 , w_19588 , w_19589 , w_19590 , w_19591 , w_19592 , w_19593 , w_19594 , w_19595 , 
		w_19596 , w_19597 , w_19598 , w_19599 , w_19600 , w_19601 , w_19602 , w_19603 , w_19604 , w_19605 , 
		w_19606 , w_19607 , w_19608 , w_19609 , w_19610 , w_19611 , w_19612 , w_19613 , w_19614 , w_19615 , 
		w_19616 , w_19617 , w_19618 , w_19619 , w_19620 , w_19621 , w_19622 , w_19623 , w_19624 , w_19625 , 
		w_19626 , w_19627 , w_19628 , w_19629 , w_19630 , w_19631 , w_19632 , w_19633 , w_19634 , w_19635 , 
		w_19636 , w_19637 , w_19638 , w_19639 , w_19640 , w_19641 , w_19642 , w_19643 , w_19644 , w_19645 , 
		w_19646 , w_19647 , w_19648 , w_19649 , w_19650 , w_19651 , w_19652 , w_19653 , w_19654 , w_19655 , 
		w_19656 , w_19657 , w_19658 , w_19659 , w_19660 , w_19661 , w_19662 , w_19663 , w_19664 , w_19665 , 
		w_19666 , w_19667 , w_19668 , w_19669 , w_19670 , w_19671 , w_19672 , w_19673 , w_19674 , w_19675 , 
		w_19676 , w_19677 , w_19678 , w_19679 , w_19680 , w_19681 , w_19682 , w_19683 , w_19684 , w_19685 , 
		w_19686 , w_19687 , w_19688 , w_19689 , w_19690 , w_19691 , w_19692 , w_19693 , w_19694 , w_19695 , 
		w_19696 , w_19697 , w_19698 , w_19699 , w_19700 , w_19701 , w_19702 , w_19703 , w_19704 , w_19705 , 
		w_19706 , w_19707 , w_19708 , w_19709 , w_19710 , w_19711 , w_19712 , w_19713 , w_19714 , w_19715 , 
		w_19716 , w_19717 , w_19718 , w_19719 , w_19720 , w_19721 , w_19722 , w_19723 , w_19724 , w_19725 , 
		w_19726 , w_19727 , w_19728 , w_19729 , w_19730 , w_19731 , w_19732 , w_19733 , w_19734 , w_19735 , 
		w_19736 , w_19737 , w_19738 , w_19739 , w_19740 , w_19741 , w_19742 , w_19743 , w_19744 , w_19745 , 
		w_19746 , w_19747 , w_19748 , w_19749 , w_19750 , w_19751 , w_19752 , w_19753 , w_19754 , w_19755 , 
		w_19756 , w_19757 , w_19758 , w_19759 , w_19760 , w_19761 , w_19762 , w_19763 , w_19764 , w_19765 , 
		w_19766 , w_19767 , w_19768 , w_19769 , w_19770 , w_19771 , w_19772 , w_19773 , w_19774 , w_19775 , 
		w_19776 , w_19777 , w_19778 , w_19779 , w_19780 , w_19781 , w_19782 , w_19783 , w_19784 , w_19785 , 
		w_19786 , w_19787 , w_19788 , w_19789 , w_19790 , w_19791 , w_19792 , w_19793 , w_19794 , w_19795 , 
		w_19796 , w_19797 , w_19798 , w_19799 , w_19800 , w_19801 , w_19802 , w_19803 , w_19804 , w_19805 , 
		w_19806 , w_19807 , w_19808 , w_19809 , w_19810 , w_19811 , w_19812 , w_19813 , w_19814 , w_19815 , 
		w_19816 , w_19817 , w_19818 , w_19819 , w_19820 , w_19821 , w_19822 , w_19823 , w_19824 , w_19825 , 
		w_19826 , w_19827 , w_19828 , w_19829 , w_19830 , w_19831 , w_19832 , w_19833 , w_19834 , w_19835 , 
		w_19836 , w_19837 , w_19838 , w_19839 , w_19840 , w_19841 , w_19842 , w_19843 , w_19844 , w_19845 , 
		w_19846 , w_19847 , w_19848 , w_19849 , w_19850 , w_19851 , w_19852 , w_19853 , w_19854 , w_19855 , 
		w_19856 , w_19857 , w_19858 , w_19859 , w_19860 , w_19861 , w_19862 , w_19863 , w_19864 , w_19865 , 
		w_19866 , w_19867 , w_19868 , w_19869 , w_19870 , w_19871 , w_19872 , w_19873 , w_19874 , w_19875 , 
		w_19876 , w_19877 , w_19878 , w_19879 , w_19880 , w_19881 , w_19882 , w_19883 , w_19884 , w_19885 , 
		w_19886 , w_19887 , w_19888 , w_19889 , w_19890 , w_19891 , w_19892 , w_19893 , w_19894 , w_19895 , 
		w_19896 , w_19897 , w_19898 , w_19899 , w_19900 , w_19901 , w_19902 , w_19903 , w_19904 , w_19905 , 
		w_19906 , w_19907 , w_19908 , w_19909 , w_19910 , w_19911 , w_19912 , w_19913 , w_19914 , w_19915 , 
		w_19916 , w_19917 , w_19918 , w_19919 , w_19920 , w_19921 , w_19922 , w_19923 , w_19924 , w_19925 , 
		w_19926 , w_19927 , w_19928 , w_19929 , w_19930 , w_19931 , w_19932 , w_19933 , w_19934 , w_19935 , 
		w_19936 , w_19937 , w_19938 , w_19939 , w_19940 , w_19941 , w_19942 , w_19943 , w_19944 , w_19945 , 
		w_19946 , w_19947 , w_19948 , w_19949 , w_19950 , w_19951 , w_19952 , w_19953 , w_19954 , w_19955 , 
		w_19956 , w_19957 , w_19958 , w_19959 , w_19960 , w_19961 , w_19962 , w_19963 , w_19964 , w_19965 , 
		w_19966 , w_19967 , w_19968 , w_19969 , w_19970 , w_19971 , w_19972 , w_19973 , w_19974 , w_19975 , 
		w_19976 , w_19977 , w_19978 , w_19979 , w_19980 , w_19981 , w_19982 , w_19983 , w_19984 , w_19985 , 
		w_19986 , w_19987 , w_19988 , w_19989 , w_19990 , w_19991 , w_19992 , w_19993 , w_19994 , w_19995 , 
		w_19996 , w_19997 , w_19998 , w_19999 , w_20000 , w_20001 , w_20002 , w_20003 , w_20004 , w_20005 , 
		w_20006 , w_20007 , w_20008 , w_20009 , w_20010 , w_20011 , w_20012 , w_20013 , w_20014 , w_20015 , 
		w_20016 , w_20017 , w_20018 , w_20019 , w_20020 , w_20021 , w_20022 , w_20023 , w_20024 , w_20025 , 
		w_20026 , w_20027 , w_20028 , w_20029 , w_20030 , w_20031 , w_20032 , w_20033 , w_20034 , w_20035 , 
		w_20036 , w_20037 , w_20038 , w_20039 , w_20040 , w_20041 , w_20042 , w_20043 , w_20044 , w_20045 , 
		w_20046 , w_20047 , w_20048 , w_20049 , w_20050 , w_20051 , w_20052 , w_20053 , w_20054 , w_20055 , 
		w_20056 , w_20057 , w_20058 , w_20059 , w_20060 , w_20061 , w_20062 , w_20063 , w_20064 , w_20065 , 
		w_20066 , w_20067 , w_20068 , w_20069 , w_20070 , w_20071 , w_20072 , w_20073 , w_20074 , w_20075 , 
		w_20076 , w_20077 , w_20078 , w_20079 , w_20080 , w_20081 , w_20082 , w_20083 , w_20084 , w_20085 , 
		w_20086 , w_20087 , w_20088 , w_20089 , w_20090 , w_20091 , w_20092 , w_20093 , w_20094 , w_20095 , 
		w_20096 , w_20097 , w_20098 , w_20099 , w_20100 , w_20101 , w_20102 , w_20103 , w_20104 , w_20105 , 
		w_20106 , w_20107 , w_20108 , w_20109 , w_20110 , w_20111 , w_20112 , w_20113 , w_20114 , w_20115 , 
		w_20116 , w_20117 , w_20118 , w_20119 , w_20120 , w_20121 , w_20122 , w_20123 , w_20124 , w_20125 , 
		w_20126 , w_20127 , w_20128 , w_20129 , w_20130 , w_20131 , w_20132 , w_20133 , w_20134 , w_20135 , 
		w_20136 , w_20137 , w_20138 , w_20139 , w_20140 , w_20141 , w_20142 , w_20143 , w_20144 , w_20145 , 
		w_20146 , w_20147 , w_20148 , w_20149 , w_20150 , w_20151 , w_20152 , w_20153 , w_20154 , w_20155 , 
		w_20156 , w_20157 , w_20158 , w_20159 , w_20160 , w_20161 , w_20162 , w_20163 , w_20164 , w_20165 , 
		w_20166 , w_20167 , w_20168 , w_20169 , w_20170 , w_20171 , w_20172 , w_20173 , w_20174 , w_20175 , 
		w_20176 , w_20177 , w_20178 , w_20179 , w_20180 , w_20181 , w_20182 , w_20183 , w_20184 , w_20185 , 
		w_20186 , w_20187 , w_20188 , w_20189 , w_20190 , w_20191 , w_20192 , w_20193 , w_20194 , w_20195 , 
		w_20196 , w_20197 , w_20198 , w_20199 , w_20200 , w_20201 , w_20202 , w_20203 , w_20204 , w_20205 , 
		w_20206 , w_20207 , w_20208 , w_20209 , w_20210 , w_20211 , w_20212 , w_20213 , w_20214 , w_20215 , 
		w_20216 , w_20217 , w_20218 , w_20219 , w_20220 , w_20221 , w_20222 , w_20223 , w_20224 , w_20225 , 
		w_20226 , w_20227 , w_20228 , w_20229 , w_20230 , w_20231 , w_20232 , w_20233 , w_20234 , w_20235 , 
		w_20236 , w_20237 , w_20238 , w_20239 , w_20240 , w_20241 , w_20242 , w_20243 , w_20244 , w_20245 , 
		w_20246 , w_20247 , w_20248 , w_20249 , w_20250 , w_20251 , w_20252 , w_20253 , w_20254 , w_20255 , 
		w_20256 , w_20257 , w_20258 , w_20259 , w_20260 , w_20261 , w_20262 , w_20263 , w_20264 , w_20265 , 
		w_20266 , w_20267 , w_20268 , w_20269 , w_20270 , w_20271 , w_20272 , w_20273 , w_20274 , w_20275 , 
		w_20276 , w_20277 , w_20278 , w_20279 , w_20280 , w_20281 , w_20282 , w_20283 , w_20284 , w_20285 , 
		w_20286 , w_20287 , w_20288 , w_20289 , w_20290 , w_20291 , w_20292 , w_20293 , w_20294 , w_20295 , 
		w_20296 , w_20297 , w_20298 , w_20299 , w_20300 , w_20301 , w_20302 , w_20303 , w_20304 , w_20305 , 
		w_20306 , w_20307 , w_20308 , w_20309 , w_20310 , w_20311 , w_20312 , w_20313 , w_20314 , w_20315 , 
		w_20316 , w_20317 , w_20318 , w_20319 , w_20320 , w_20321 , w_20322 , w_20323 , w_20324 , w_20325 , 
		w_20326 , w_20327 , w_20328 , w_20329 , w_20330 , w_20331 , w_20332 , w_20333 , w_20334 , w_20335 , 
		w_20336 , w_20337 , w_20338 , w_20339 , w_20340 , w_20341 , w_20342 , w_20343 , w_20344 , w_20345 , 
		w_20346 , w_20347 , w_20348 , w_20349 , w_20350 , w_20351 , w_20352 , w_20353 , w_20354 , w_20355 , 
		w_20356 , w_20357 , w_20358 , w_20359 , w_20360 , w_20361 , w_20362 , w_20363 , w_20364 , w_20365 , 
		w_20366 , w_20367 , w_20368 , w_20369 , w_20370 , w_20371 , w_20372 , w_20373 , w_20374 , w_20375 , 
		w_20376 , w_20377 , w_20378 , w_20379 , w_20380 , w_20381 , w_20382 , w_20383 , w_20384 , w_20385 , 
		w_20386 , w_20387 , w_20388 , w_20389 , w_20390 , w_20391 , w_20392 , w_20393 , w_20394 , w_20395 , 
		w_20396 , w_20397 , w_20398 , w_20399 , w_20400 , w_20401 , w_20402 , w_20403 , w_20404 , w_20405 , 
		w_20406 , w_20407 , w_20408 , w_20409 , w_20410 , w_20411 , w_20412 , w_20413 , w_20414 , w_20415 , 
		w_20416 , w_20417 , w_20418 , w_20419 , w_20420 , w_20421 , w_20422 , w_20423 , w_20424 , w_20425 , 
		w_20426 , w_20427 , w_20428 , w_20429 , w_20430 , w_20431 , w_20432 , w_20433 , w_20434 , w_20435 , 
		w_20436 , w_20437 , w_20438 , w_20439 , w_20440 , w_20441 , w_20442 , w_20443 , w_20444 , w_20445 , 
		w_20446 , w_20447 , w_20448 , w_20449 , w_20450 , w_20451 , w_20452 , w_20453 , w_20454 , w_20455 , 
		w_20456 , w_20457 , w_20458 , w_20459 , w_20460 , w_20461 , w_20462 , w_20463 , w_20464 , w_20465 , 
		w_20466 , w_20467 , w_20468 , w_20469 , w_20470 , w_20471 , w_20472 , w_20473 , w_20474 , w_20475 , 
		w_20476 , w_20477 , w_20478 , w_20479 , w_20480 , w_20481 , w_20482 , w_20483 , w_20484 , w_20485 , 
		w_20486 , w_20487 , w_20488 , w_20489 , w_20490 , w_20491 , w_20492 , w_20493 , w_20494 , w_20495 , 
		w_20496 , w_20497 , w_20498 , w_20499 , w_20500 , w_20501 , w_20502 , w_20503 , w_20504 , w_20505 , 
		w_20506 , w_20507 , w_20508 , w_20509 , w_20510 , w_20511 , w_20512 , w_20513 , w_20514 , w_20515 , 
		w_20516 , w_20517 , w_20518 , w_20519 , w_20520 , w_20521 , w_20522 , w_20523 , w_20524 , w_20525 , 
		w_20526 , w_20527 , w_20528 , w_20529 , w_20530 , w_20531 , w_20532 , w_20533 , w_20534 , w_20535 , 
		w_20536 , w_20537 , w_20538 , w_20539 , w_20540 , w_20541 , w_20542 , w_20543 , w_20544 , w_20545 , 
		w_20546 , w_20547 , w_20548 , w_20549 , w_20550 , w_20551 , w_20552 , w_20553 , w_20554 , w_20555 , 
		w_20556 , w_20557 , w_20558 , w_20559 , w_20560 , w_20561 , w_20562 , w_20563 , w_20564 , w_20565 , 
		w_20566 , w_20567 , w_20568 , w_20569 , w_20570 , w_20571 , w_20572 , w_20573 , w_20574 , w_20575 , 
		w_20576 , w_20577 , w_20578 , w_20579 , w_20580 , w_20581 , w_20582 , w_20583 , w_20584 , w_20585 , 
		w_20586 , w_20587 , w_20588 , w_20589 , w_20590 , w_20591 , w_20592 , w_20593 , w_20594 , w_20595 , 
		w_20596 , w_20597 , w_20598 , w_20599 , w_20600 , w_20601 , w_20602 , w_20603 , w_20604 , w_20605 , 
		w_20606 , w_20607 , w_20608 , w_20609 , w_20610 , w_20611 , w_20612 , w_20613 , w_20614 , w_20615 , 
		w_20616 , w_20617 , w_20618 , w_20619 , w_20620 , w_20621 , w_20622 , w_20623 , w_20624 , w_20625 , 
		w_20626 , w_20627 , w_20628 , w_20629 , w_20630 , w_20631 , w_20632 , w_20633 , w_20634 , w_20635 , 
		w_20636 , w_20637 , w_20638 , w_20639 , w_20640 , w_20641 , w_20642 , w_20643 , w_20644 , w_20645 , 
		w_20646 , w_20647 , w_20648 , w_20649 , w_20650 , w_20651 , w_20652 , w_20653 , w_20654 , w_20655 , 
		w_20656 , w_20657 , w_20658 , w_20659 , w_20660 , w_20661 , w_20662 , w_20663 , w_20664 , w_20665 , 
		w_20666 , w_20667 , w_20668 , w_20669 , w_20670 , w_20671 , w_20672 , w_20673 , w_20674 , w_20675 , 
		w_20676 , w_20677 , w_20678 , w_20679 , w_20680 , w_20681 , w_20682 , w_20683 , w_20684 , w_20685 , 
		w_20686 , w_20687 , w_20688 , w_20689 , w_20690 , w_20691 , w_20692 , w_20693 , w_20694 , w_20695 , 
		w_20696 , w_20697 , w_20698 , w_20699 , w_20700 , w_20701 , w_20702 , w_20703 , w_20704 , w_20705 , 
		w_20706 , w_20707 , w_20708 , w_20709 , w_20710 , w_20711 , w_20712 , w_20713 , w_20714 , w_20715 , 
		w_20716 , w_20717 , w_20718 , w_20719 , w_20720 , w_20721 , w_20722 , w_20723 , w_20724 , w_20725 , 
		w_20726 , w_20727 , w_20728 , w_20729 , w_20730 , w_20731 , w_20732 , w_20733 , w_20734 , w_20735 , 
		w_20736 , w_20737 , w_20738 , w_20739 , w_20740 , w_20741 , w_20742 , w_20743 , w_20744 , w_20745 , 
		w_20746 , w_20747 , w_20748 , w_20749 , w_20750 , w_20751 , w_20752 , w_20753 , w_20754 , w_20755 , 
		w_20756 , w_20757 , w_20758 , w_20759 , w_20760 , w_20761 , w_20762 , w_20763 , w_20764 , w_20765 , 
		w_20766 , w_20767 , w_20768 , w_20769 , w_20770 , w_20771 , w_20772 , w_20773 , w_20774 , w_20775 , 
		w_20776 , w_20777 , w_20778 , w_20779 , w_20780 , w_20781 , w_20782 , w_20783 , w_20784 , w_20785 , 
		w_20786 , w_20787 , w_20788 , w_20789 , w_20790 , w_20791 , w_20792 , w_20793 , w_20794 , w_20795 , 
		w_20796 , w_20797 , w_20798 , w_20799 , w_20800 , w_20801 , w_20802 , w_20803 , w_20804 , w_20805 , 
		w_20806 , w_20807 , w_20808 , w_20809 , w_20810 , w_20811 , w_20812 , w_20813 , w_20814 , w_20815 , 
		w_20816 , w_20817 , w_20818 , w_20819 , w_20820 , w_20821 , w_20822 , w_20823 , w_20824 , w_20825 , 
		w_20826 , w_20827 , w_20828 , w_20829 , w_20830 , w_20831 , w_20832 , w_20833 , w_20834 , w_20835 , 
		w_20836 , w_20837 , w_20838 , w_20839 , w_20840 , w_20841 , w_20842 , w_20843 , w_20844 , w_20845 , 
		w_20846 , w_20847 , w_20848 , w_20849 , w_20850 , w_20851 , w_20852 , w_20853 , w_20854 , w_20855 , 
		w_20856 , w_20857 , w_20858 , w_20859 , w_20860 , w_20861 , w_20862 , w_20863 , w_20864 , w_20865 , 
		w_20866 , w_20867 , w_20868 , w_20869 , w_20870 , w_20871 , w_20872 , w_20873 , w_20874 , w_20875 , 
		w_20876 , w_20877 , w_20878 , w_20879 , w_20880 , w_20881 , w_20882 , w_20883 , w_20884 , w_20885 , 
		w_20886 , w_20887 , w_20888 , w_20889 , w_20890 , w_20891 , w_20892 , w_20893 , w_20894 , w_20895 , 
		w_20896 , w_20897 , w_20898 , w_20899 , w_20900 , w_20901 , w_20902 , w_20903 , w_20904 , w_20905 , 
		w_20906 , w_20907 , w_20908 , w_20909 , w_20910 , w_20911 , w_20912 , w_20913 , w_20914 , w_20915 , 
		w_20916 , w_20917 , w_20918 , w_20919 , w_20920 , w_20921 , w_20922 , w_20923 , w_20924 , w_20925 , 
		w_20926 , w_20927 , w_20928 , w_20929 , w_20930 , w_20931 , w_20932 , w_20933 , w_20934 , w_20935 , 
		w_20936 , w_20937 , w_20938 , w_20939 , w_20940 , w_20941 , w_20942 , w_20943 , w_20944 , w_20945 , 
		w_20946 , w_20947 , w_20948 , w_20949 , w_20950 , w_20951 , w_20952 , w_20953 , w_20954 , w_20955 , 
		w_20956 , w_20957 , w_20958 , w_20959 , w_20960 , w_20961 , w_20962 , w_20963 , w_20964 , w_20965 , 
		w_20966 , w_20967 , w_20968 , w_20969 , w_20970 , w_20971 , w_20972 , w_20973 , w_20974 , w_20975 , 
		w_20976 , w_20977 , w_20978 , w_20979 , w_20980 , w_20981 , w_20982 , w_20983 , w_20984 , w_20985 , 
		w_20986 , w_20987 , w_20988 , w_20989 , w_20990 , w_20991 , w_20992 , w_20993 , w_20994 , w_20995 , 
		w_20996 , w_20997 , w_20998 , w_20999 , w_21000 , w_21001 , w_21002 , w_21003 , w_21004 , w_21005 , 
		w_21006 , w_21007 , w_21008 , w_21009 , w_21010 , w_21011 , w_21012 , w_21013 , w_21014 , w_21015 , 
		w_21016 , w_21017 , w_21018 , w_21019 , w_21020 , w_21021 , w_21022 , w_21023 , w_21024 , w_21025 , 
		w_21026 , w_21027 , w_21028 , w_21029 , w_21030 , w_21031 , w_21032 , w_21033 , w_21034 , w_21035 , 
		w_21036 , w_21037 , w_21038 , w_21039 , w_21040 , w_21041 , w_21042 , w_21043 , w_21044 , w_21045 , 
		w_21046 , w_21047 , w_21048 , w_21049 , w_21050 , w_21051 , w_21052 , w_21053 , w_21054 , w_21055 , 
		w_21056 , w_21057 , w_21058 , w_21059 , w_21060 , w_21061 , w_21062 , w_21063 , w_21064 , w_21065 , 
		w_21066 , w_21067 , w_21068 , w_21069 , w_21070 , w_21071 , w_21072 , w_21073 , w_21074 , w_21075 , 
		w_21076 , w_21077 , w_21078 , w_21079 , w_21080 , w_21081 , w_21082 , w_21083 , w_21084 , w_21085 , 
		w_21086 , w_21087 , w_21088 , w_21089 , w_21090 , w_21091 , w_21092 , w_21093 , w_21094 , w_21095 , 
		w_21096 , w_21097 , w_21098 , w_21099 , w_21100 , w_21101 , w_21102 , w_21103 , w_21104 , w_21105 , 
		w_21106 , w_21107 , w_21108 , w_21109 , w_21110 , w_21111 , w_21112 , w_21113 , w_21114 , w_21115 , 
		w_21116 , w_21117 , w_21118 , w_21119 , w_21120 , w_21121 , w_21122 , w_21123 , w_21124 , w_21125 , 
		w_21126 , w_21127 , w_21128 , w_21129 , w_21130 , w_21131 , w_21132 , w_21133 , w_21134 , w_21135 , 
		w_21136 , w_21137 , w_21138 , w_21139 , w_21140 , w_21141 , w_21142 , w_21143 , w_21144 , w_21145 , 
		w_21146 , w_21147 , w_21148 , w_21149 , w_21150 , w_21151 , w_21152 , w_21153 , w_21154 , w_21155 , 
		w_21156 , w_21157 , w_21158 , w_21159 , w_21160 , w_21161 , w_21162 , w_21163 , w_21164 , w_21165 , 
		w_21166 , w_21167 , w_21168 , w_21169 , w_21170 , w_21171 , w_21172 , w_21173 , w_21174 , w_21175 , 
		w_21176 , w_21177 , w_21178 , w_21179 , w_21180 , w_21181 , w_21182 , w_21183 , w_21184 , w_21185 , 
		w_21186 , w_21187 , w_21188 , w_21189 , w_21190 , w_21191 , w_21192 , w_21193 , w_21194 , w_21195 , 
		w_21196 , w_21197 , w_21198 , w_21199 , w_21200 , w_21201 , w_21202 , w_21203 , w_21204 , w_21205 , 
		w_21206 , w_21207 , w_21208 , w_21209 , w_21210 , w_21211 , w_21212 , w_21213 , w_21214 , w_21215 , 
		w_21216 , w_21217 , w_21218 , w_21219 , w_21220 , w_21221 , w_21222 , w_21223 , w_21224 , w_21225 , 
		w_21226 , w_21227 , w_21228 , w_21229 , w_21230 , w_21231 , w_21232 , w_21233 , w_21234 , w_21235 , 
		w_21236 , w_21237 , w_21238 , w_21239 , w_21240 , w_21241 , w_21242 , w_21243 , w_21244 , w_21245 , 
		w_21246 , w_21247 , w_21248 , w_21249 , w_21250 , w_21251 , w_21252 , w_21253 , w_21254 , w_21255 , 
		w_21256 , w_21257 , w_21258 , w_21259 , w_21260 , w_21261 , w_21262 , w_21263 , w_21264 , w_21265 , 
		w_21266 , w_21267 , w_21268 , w_21269 , w_21270 , w_21271 , w_21272 , w_21273 , w_21274 , w_21275 , 
		w_21276 , w_21277 , w_21278 , w_21279 , w_21280 , w_21281 , w_21282 , w_21283 , w_21284 , w_21285 , 
		w_21286 , w_21287 , w_21288 , w_21289 , w_21290 , w_21291 , w_21292 , w_21293 , w_21294 , w_21295 , 
		w_21296 , w_21297 , w_21298 , w_21299 , w_21300 , w_21301 , w_21302 , w_21303 , w_21304 , w_21305 , 
		w_21306 , w_21307 , w_21308 , w_21309 , w_21310 , w_21311 , w_21312 , w_21313 , w_21314 , w_21315 , 
		w_21316 , w_21317 , w_21318 , w_21319 , w_21320 , w_21321 , w_21322 , w_21323 , w_21324 , w_21325 , 
		w_21326 , w_21327 , w_21328 , w_21329 , w_21330 , w_21331 , w_21332 , w_21333 , w_21334 , w_21335 , 
		w_21336 , w_21337 , w_21338 , w_21339 , w_21340 , w_21341 , w_21342 , w_21343 , w_21344 , w_21345 , 
		w_21346 , w_21347 , w_21348 , w_21349 , w_21350 , w_21351 , w_21352 , w_21353 , w_21354 , w_21355 , 
		w_21356 , w_21357 , w_21358 , w_21359 , w_21360 , w_21361 , w_21362 , w_21363 , w_21364 , w_21365 , 
		w_21366 , w_21367 , w_21368 , w_21369 , w_21370 , w_21371 , w_21372 , w_21373 , w_21374 , w_21375 , 
		w_21376 , w_21377 , w_21378 , w_21379 , w_21380 , w_21381 , w_21382 , w_21383 , w_21384 , w_21385 , 
		w_21386 , w_21387 , w_21388 , w_21389 , w_21390 , w_21391 , w_21392 , w_21393 , w_21394 , w_21395 , 
		w_21396 , w_21397 , w_21398 , w_21399 , w_21400 , w_21401 , w_21402 , w_21403 , w_21404 , w_21405 , 
		w_21406 , w_21407 , w_21408 , w_21409 , w_21410 , w_21411 , w_21412 , w_21413 , w_21414 , w_21415 , 
		w_21416 , w_21417 , w_21418 , w_21419 , w_21420 , w_21421 , w_21422 , w_21423 , w_21424 , w_21425 , 
		w_21426 , w_21427 , w_21428 , w_21429 , w_21430 , w_21431 , w_21432 , w_21433 , w_21434 , w_21435 , 
		w_21436 , w_21437 , w_21438 , w_21439 , w_21440 , w_21441 , w_21442 , w_21443 , w_21444 , w_21445 , 
		w_21446 , w_21447 , w_21448 , w_21449 , w_21450 , w_21451 , w_21452 , w_21453 , w_21454 , w_21455 , 
		w_21456 , w_21457 , w_21458 , w_21459 , w_21460 , w_21461 , w_21462 , w_21463 , w_21464 , w_21465 , 
		w_21466 , w_21467 , w_21468 , w_21469 , w_21470 , w_21471 , w_21472 , w_21473 , w_21474 , w_21475 , 
		w_21476 , w_21477 , w_21478 , w_21479 , w_21480 , w_21481 , w_21482 , w_21483 , w_21484 , w_21485 , 
		w_21486 , w_21487 , w_21488 , w_21489 , w_21490 , w_21491 , w_21492 , w_21493 , w_21494 , w_21495 , 
		w_21496 , w_21497 , w_21498 , w_21499 , w_21500 , w_21501 , w_21502 , w_21503 , w_21504 , w_21505 , 
		w_21506 , w_21507 , w_21508 , w_21509 , w_21510 , w_21511 , w_21512 , w_21513 , w_21514 , w_21515 , 
		w_21516 , w_21517 , w_21518 , w_21519 , w_21520 , w_21521 , w_21522 , w_21523 , w_21524 , w_21525 , 
		w_21526 , w_21527 , w_21528 , w_21529 , w_21530 , w_21531 , w_21532 , w_21533 , w_21534 , w_21535 , 
		w_21536 , w_21537 , w_21538 , w_21539 , w_21540 , w_21541 , w_21542 , w_21543 , w_21544 , w_21545 , 
		w_21546 , w_21547 , w_21548 , w_21549 , w_21550 , w_21551 , w_21552 , w_21553 , w_21554 , w_21555 , 
		w_21556 , w_21557 , w_21558 , w_21559 , w_21560 , w_21561 , w_21562 , w_21563 , w_21564 , w_21565 , 
		w_21566 , w_21567 , w_21568 , w_21569 , w_21570 , w_21571 , w_21572 , w_21573 , w_21574 , w_21575 , 
		w_21576 , w_21577 , w_21578 , w_21579 , w_21580 , w_21581 , w_21582 , w_21583 , w_21584 , w_21585 , 
		w_21586 , w_21587 , w_21588 , w_21589 , w_21590 , w_21591 , w_21592 , w_21593 , w_21594 , w_21595 , 
		w_21596 , w_21597 , w_21598 , w_21599 , w_21600 , w_21601 , w_21602 , w_21603 , w_21604 , w_21605 , 
		w_21606 , w_21607 , w_21608 , w_21609 , w_21610 , w_21611 , w_21612 , w_21613 , w_21614 , w_21615 , 
		w_21616 , w_21617 , w_21618 , w_21619 , w_21620 , w_21621 , w_21622 , w_21623 , w_21624 , w_21625 , 
		w_21626 , w_21627 , w_21628 , w_21629 , w_21630 , w_21631 , w_21632 , w_21633 , w_21634 , w_21635 , 
		w_21636 , w_21637 , w_21638 , w_21639 , w_21640 , w_21641 , w_21642 , w_21643 , w_21644 , w_21645 , 
		w_21646 , w_21647 , w_21648 , w_21649 , w_21650 , w_21651 , w_21652 , w_21653 , w_21654 , w_21655 , 
		w_21656 , w_21657 , w_21658 , w_21659 , w_21660 , w_21661 , w_21662 , w_21663 , w_21664 , w_21665 , 
		w_21666 , w_21667 , w_21668 , w_21669 , w_21670 , w_21671 , w_21672 , w_21673 , w_21674 , w_21675 , 
		w_21676 , w_21677 , w_21678 , w_21679 , w_21680 , w_21681 , w_21682 , w_21683 , w_21684 , w_21685 , 
		w_21686 , w_21687 , w_21688 , w_21689 , w_21690 , w_21691 , w_21692 , w_21693 , w_21694 , w_21695 , 
		w_21696 , w_21697 , w_21698 , w_21699 , w_21700 , w_21701 , w_21702 , w_21703 , w_21704 , w_21705 , 
		w_21706 , w_21707 , w_21708 , w_21709 , w_21710 , w_21711 , w_21712 , w_21713 , w_21714 , w_21715 , 
		w_21716 , w_21717 , w_21718 , w_21719 , w_21720 , w_21721 , w_21722 , w_21723 , w_21724 , w_21725 , 
		w_21726 , w_21727 , w_21728 , w_21729 , w_21730 , w_21731 , w_21732 , w_21733 , w_21734 , w_21735 , 
		w_21736 , w_21737 , w_21738 , w_21739 , w_21740 , w_21741 , w_21742 , w_21743 , w_21744 , w_21745 , 
		w_21746 , w_21747 , w_21748 , w_21749 , w_21750 , w_21751 , w_21752 , w_21753 , w_21754 , w_21755 , 
		w_21756 , w_21757 , w_21758 , w_21759 , w_21760 , w_21761 , w_21762 , w_21763 , w_21764 , w_21765 , 
		w_21766 , w_21767 , w_21768 , w_21769 , w_21770 , w_21771 , w_21772 , w_21773 , w_21774 , w_21775 , 
		w_21776 , w_21777 , w_21778 , w_21779 , w_21780 , w_21781 , w_21782 , w_21783 , w_21784 , w_21785 , 
		w_21786 , w_21787 , w_21788 , w_21789 , w_21790 , w_21791 , w_21792 , w_21793 , w_21794 , w_21795 , 
		w_21796 , w_21797 , w_21798 , w_21799 , w_21800 , w_21801 , w_21802 , w_21803 , w_21804 , w_21805 , 
		w_21806 , w_21807 , w_21808 , w_21809 , w_21810 , w_21811 , w_21812 , w_21813 , w_21814 , w_21815 , 
		w_21816 , w_21817 , w_21818 , w_21819 , w_21820 , w_21821 , w_21822 , w_21823 , w_21824 , w_21825 , 
		w_21826 , w_21827 , w_21828 , w_21829 , w_21830 , w_21831 , w_21832 , w_21833 , w_21834 , w_21835 , 
		w_21836 , w_21837 , w_21838 , w_21839 , w_21840 , w_21841 , w_21842 , w_21843 , w_21844 , w_21845 , 
		w_21846 , w_21847 , w_21848 , w_21849 , w_21850 , w_21851 , w_21852 , w_21853 , w_21854 , w_21855 , 
		w_21856 , w_21857 , w_21858 , w_21859 , w_21860 , w_21861 , w_21862 , w_21863 , w_21864 , w_21865 , 
		w_21866 , w_21867 , w_21868 , w_21869 , w_21870 , w_21871 , w_21872 , w_21873 , w_21874 , w_21875 , 
		w_21876 , w_21877 , w_21878 , w_21879 , w_21880 , w_21881 , w_21882 , w_21883 , w_21884 , w_21885 , 
		w_21886 , w_21887 , w_21888 , w_21889 , w_21890 , w_21891 , w_21892 , w_21893 , w_21894 , w_21895 , 
		w_21896 , w_21897 , w_21898 , w_21899 , w_21900 , w_21901 , w_21902 , w_21903 , w_21904 , w_21905 , 
		w_21906 , w_21907 , w_21908 , w_21909 , w_21910 , w_21911 , w_21912 , w_21913 , w_21914 , w_21915 , 
		w_21916 , w_21917 , w_21918 , w_21919 , w_21920 , w_21921 , w_21922 , w_21923 , w_21924 , w_21925 , 
		w_21926 , w_21927 , w_21928 , w_21929 , w_21930 , w_21931 , w_21932 , w_21933 , w_21934 , w_21935 , 
		w_21936 , w_21937 , w_21938 , w_21939 , w_21940 , w_21941 , w_21942 , w_21943 , w_21944 , w_21945 , 
		w_21946 , w_21947 , w_21948 , w_21949 , w_21950 , w_21951 , w_21952 , w_21953 , w_21954 , w_21955 , 
		w_21956 , w_21957 , w_21958 , w_21959 , w_21960 , w_21961 , w_21962 , w_21963 , w_21964 , w_21965 , 
		w_21966 , w_21967 , w_21968 , w_21969 , w_21970 , w_21971 , w_21972 , w_21973 , w_21974 , w_21975 , 
		w_21976 , w_21977 , w_21978 , w_21979 , w_21980 , w_21981 , w_21982 , w_21983 , w_21984 , w_21985 , 
		w_21986 , w_21987 , w_21988 , w_21989 , w_21990 , w_21991 , w_21992 , w_21993 , w_21994 , w_21995 , 
		w_21996 , w_21997 , w_21998 , w_21999 , w_22000 , w_22001 , w_22002 , w_22003 , w_22004 , w_22005 , 
		w_22006 , w_22007 , w_22008 , w_22009 , w_22010 , w_22011 , w_22012 , w_22013 , w_22014 , w_22015 , 
		w_22016 , w_22017 , w_22018 , w_22019 , w_22020 , w_22021 , w_22022 , w_22023 , w_22024 , w_22025 , 
		w_22026 , w_22027 , w_22028 , w_22029 , w_22030 , w_22031 , w_22032 , w_22033 , w_22034 , w_22035 , 
		w_22036 , w_22037 , w_22038 , w_22039 , w_22040 , w_22041 , w_22042 , w_22043 , w_22044 , w_22045 , 
		w_22046 , w_22047 , w_22048 , w_22049 , w_22050 , w_22051 , w_22052 , w_22053 , w_22054 , w_22055 , 
		w_22056 , w_22057 , w_22058 , w_22059 , w_22060 , w_22061 , w_22062 , w_22063 , w_22064 , w_22065 , 
		w_22066 , w_22067 , w_22068 , w_22069 , w_22070 , w_22071 , w_22072 , w_22073 , w_22074 , w_22075 , 
		w_22076 , w_22077 , w_22078 , w_22079 , w_22080 , w_22081 , w_22082 , w_22083 , w_22084 , w_22085 , 
		w_22086 , w_22087 , w_22088 , w_22089 , w_22090 , w_22091 , w_22092 , w_22093 , w_22094 , w_22095 , 
		w_22096 , w_22097 , w_22098 , w_22099 , w_22100 , w_22101 , w_22102 , w_22103 , w_22104 , w_22105 , 
		w_22106 , w_22107 , w_22108 , w_22109 , w_22110 , w_22111 , w_22112 , w_22113 , w_22114 , w_22115 , 
		w_22116 , w_22117 , w_22118 , w_22119 , w_22120 , w_22121 , w_22122 , w_22123 , w_22124 , w_22125 , 
		w_22126 , w_22127 , w_22128 , w_22129 , w_22130 , w_22131 , w_22132 , w_22133 , w_22134 , w_22135 , 
		w_22136 , w_22137 , w_22138 , w_22139 , w_22140 , w_22141 , w_22142 , w_22143 , w_22144 , w_22145 , 
		w_22146 , w_22147 , w_22148 , w_22149 , w_22150 , w_22151 , w_22152 , w_22153 , w_22154 , w_22155 , 
		w_22156 , w_22157 , w_22158 , w_22159 , w_22160 , w_22161 , w_22162 , w_22163 , w_22164 , w_22165 , 
		w_22166 , w_22167 , w_22168 , w_22169 , w_22170 , w_22171 , w_22172 , w_22173 , w_22174 , w_22175 , 
		w_22176 , w_22177 , w_22178 , w_22179 , w_22180 , w_22181 , w_22182 , w_22183 , w_22184 , w_22185 , 
		w_22186 , w_22187 , w_22188 , w_22189 , w_22190 , w_22191 , w_22192 , w_22193 , w_22194 , w_22195 , 
		w_22196 , w_22197 , w_22198 , w_22199 , w_22200 , w_22201 , w_22202 , w_22203 , w_22204 , w_22205 , 
		w_22206 , w_22207 , w_22208 , w_22209 , w_22210 , w_22211 , w_22212 , w_22213 , w_22214 , w_22215 , 
		w_22216 , w_22217 , w_22218 , w_22219 , w_22220 , w_22221 , w_22222 , w_22223 , w_22224 , w_22225 , 
		w_22226 , w_22227 , w_22228 , w_22229 , w_22230 , w_22231 , w_22232 , w_22233 , w_22234 , w_22235 , 
		w_22236 , w_22237 , w_22238 , w_22239 , w_22240 , w_22241 , w_22242 , w_22243 , w_22244 , w_22245 , 
		w_22246 , w_22247 , w_22248 , w_22249 , w_22250 , w_22251 , w_22252 , w_22253 , w_22254 , w_22255 , 
		w_22256 , w_22257 , w_22258 , w_22259 , w_22260 , w_22261 , w_22262 , w_22263 , w_22264 , w_22265 , 
		w_22266 , w_22267 , w_22268 , w_22269 , w_22270 , w_22271 , w_22272 , w_22273 , w_22274 , w_22275 , 
		w_22276 , w_22277 , w_22278 , w_22279 , w_22280 , w_22281 , w_22282 , w_22283 , w_22284 , w_22285 , 
		w_22286 , w_22287 , w_22288 , w_22289 , w_22290 , w_22291 , w_22292 , w_22293 , w_22294 , w_22295 , 
		w_22296 , w_22297 , w_22298 , w_22299 , w_22300 , w_22301 , w_22302 , w_22303 , w_22304 , w_22305 , 
		w_22306 , w_22307 , w_22308 , w_22309 , w_22310 , w_22311 , w_22312 , w_22313 , w_22314 , w_22315 , 
		w_22316 , w_22317 , w_22318 , w_22319 , w_22320 , w_22321 , w_22322 , w_22323 , w_22324 , w_22325 , 
		w_22326 , w_22327 , w_22328 , w_22329 , w_22330 , w_22331 , w_22332 , w_22333 , w_22334 , w_22335 , 
		w_22336 , w_22337 , w_22338 , w_22339 , w_22340 , w_22341 , w_22342 , w_22343 , w_22344 , w_22345 , 
		w_22346 , w_22347 , w_22348 , w_22349 , w_22350 , w_22351 , w_22352 , w_22353 , w_22354 , w_22355 , 
		w_22356 , w_22357 , w_22358 , w_22359 , w_22360 , w_22361 , w_22362 , w_22363 , w_22364 , w_22365 , 
		w_22366 , w_22367 , w_22368 , w_22369 , w_22370 , w_22371 , w_22372 , w_22373 , w_22374 , w_22375 , 
		w_22376 , w_22377 , w_22378 , w_22379 , w_22380 , w_22381 , w_22382 , w_22383 , w_22384 , w_22385 , 
		w_22386 , w_22387 , w_22388 , w_22389 , w_22390 , w_22391 , w_22392 , w_22393 , w_22394 , w_22395 , 
		w_22396 , w_22397 , w_22398 , w_22399 , w_22400 , w_22401 , w_22402 , w_22403 , w_22404 , w_22405 , 
		w_22406 , w_22407 , w_22408 , w_22409 , w_22410 , w_22411 , w_22412 , w_22413 , w_22414 , w_22415 , 
		w_22416 , w_22417 , w_22418 , w_22419 , w_22420 , w_22421 , w_22422 , w_22423 , w_22424 , w_22425 , 
		w_22426 , w_22427 , w_22428 , w_22429 , w_22430 , w_22431 , w_22432 , w_22433 , w_22434 , w_22435 , 
		w_22436 , w_22437 , w_22438 , w_22439 , w_22440 , w_22441 , w_22442 , w_22443 , w_22444 , w_22445 , 
		w_22446 , w_22447 , w_22448 , w_22449 , w_22450 , w_22451 , w_22452 , w_22453 , w_22454 , w_22455 , 
		w_22456 , w_22457 , w_22458 , w_22459 , w_22460 , w_22461 , w_22462 , w_22463 , w_22464 , w_22465 , 
		w_22466 , w_22467 , w_22468 , w_22469 , w_22470 , w_22471 , w_22472 , w_22473 , w_22474 , w_22475 , 
		w_22476 , w_22477 , w_22478 , w_22479 , w_22480 , w_22481 , w_22482 , w_22483 , w_22484 , w_22485 , 
		w_22486 , w_22487 , w_22488 , w_22489 , w_22490 , w_22491 , w_22492 , w_22493 , w_22494 , w_22495 , 
		w_22496 , w_22497 , w_22498 , w_22499 , w_22500 , w_22501 , w_22502 , w_22503 , w_22504 , w_22505 , 
		w_22506 , w_22507 , w_22508 , w_22509 , w_22510 , w_22511 , w_22512 , w_22513 , w_22514 , w_22515 , 
		w_22516 , w_22517 , w_22518 , w_22519 , w_22520 , w_22521 , w_22522 , w_22523 , w_22524 , w_22525 , 
		w_22526 , w_22527 , w_22528 , w_22529 , w_22530 , w_22531 , w_22532 , w_22533 , w_22534 , w_22535 , 
		w_22536 , w_22537 , w_22538 , w_22539 , w_22540 , w_22541 , w_22542 , w_22543 , w_22544 , w_22545 , 
		w_22546 , w_22547 , w_22548 , w_22549 , w_22550 , w_22551 , w_22552 , w_22553 , w_22554 , w_22555 , 
		w_22556 , w_22557 , w_22558 , w_22559 , w_22560 , w_22561 , w_22562 , w_22563 , w_22564 , w_22565 , 
		w_22566 , w_22567 , w_22568 , w_22569 , w_22570 , w_22571 , w_22572 , w_22573 , w_22574 , w_22575 , 
		w_22576 , w_22577 , w_22578 , w_22579 , w_22580 , w_22581 , w_22582 , w_22583 , w_22584 , w_22585 , 
		w_22586 , w_22587 , w_22588 , w_22589 , w_22590 , w_22591 , w_22592 , w_22593 , w_22594 , w_22595 , 
		w_22596 , w_22597 , w_22598 , w_22599 , w_22600 , w_22601 , w_22602 , w_22603 , w_22604 , w_22605 , 
		w_22606 , w_22607 , w_22608 , w_22609 , w_22610 , w_22611 , w_22612 , w_22613 , w_22614 , w_22615 , 
		w_22616 , w_22617 , w_22618 , w_22619 , w_22620 , w_22621 , w_22622 , w_22623 , w_22624 , w_22625 , 
		w_22626 , w_22627 , w_22628 , w_22629 , w_22630 , w_22631 , w_22632 , w_22633 , w_22634 , w_22635 , 
		w_22636 , w_22637 , w_22638 , w_22639 , w_22640 , w_22641 , w_22642 , w_22643 , w_22644 , w_22645 , 
		w_22646 , w_22647 , w_22648 , w_22649 , w_22650 , w_22651 , w_22652 , w_22653 , w_22654 , w_22655 , 
		w_22656 , w_22657 , w_22658 , w_22659 , w_22660 , w_22661 , w_22662 , w_22663 , w_22664 , w_22665 , 
		w_22666 , w_22667 , w_22668 , w_22669 , w_22670 , w_22671 , w_22672 , w_22673 , w_22674 , w_22675 , 
		w_22676 , w_22677 , w_22678 , w_22679 , w_22680 , w_22681 , w_22682 , w_22683 , w_22684 , w_22685 , 
		w_22686 , w_22687 , w_22688 , w_22689 , w_22690 , w_22691 , w_22692 , w_22693 , w_22694 , w_22695 , 
		w_22696 , w_22697 , w_22698 , w_22699 , w_22700 , w_22701 , w_22702 , w_22703 , w_22704 , w_22705 , 
		w_22706 , w_22707 , w_22708 , w_22709 , w_22710 , w_22711 , w_22712 , w_22713 , w_22714 , w_22715 , 
		w_22716 , w_22717 , w_22718 , w_22719 , w_22720 , w_22721 , w_22722 , w_22723 , w_22724 , w_22725 , 
		w_22726 , w_22727 , w_22728 , w_22729 , w_22730 , w_22731 , w_22732 , w_22733 , w_22734 , w_22735 , 
		w_22736 , w_22737 , w_22738 , w_22739 , w_22740 , w_22741 , w_22742 , w_22743 , w_22744 , w_22745 , 
		w_22746 , w_22747 , w_22748 , w_22749 , w_22750 , w_22751 , w_22752 , w_22753 , w_22754 , w_22755 , 
		w_22756 , w_22757 , w_22758 , w_22759 , w_22760 , w_22761 , w_22762 , w_22763 , w_22764 , w_22765 , 
		w_22766 , w_22767 , w_22768 , w_22769 , w_22770 , w_22771 , w_22772 , w_22773 , w_22774 , w_22775 , 
		w_22776 , w_22777 , w_22778 , w_22779 , w_22780 , w_22781 , w_22782 , w_22783 , w_22784 , w_22785 , 
		w_22786 , w_22787 , w_22788 , w_22789 , w_22790 , w_22791 , w_22792 , w_22793 , w_22794 , w_22795 , 
		w_22796 , w_22797 , w_22798 , w_22799 , w_22800 , w_22801 , w_22802 , w_22803 , w_22804 , w_22805 , 
		w_22806 , w_22807 , w_22808 , w_22809 , w_22810 , w_22811 , w_22812 , w_22813 , w_22814 , w_22815 , 
		w_22816 , w_22817 , w_22818 , w_22819 , w_22820 , w_22821 , w_22822 , w_22823 , w_22824 , w_22825 , 
		w_22826 , w_22827 , w_22828 , w_22829 , w_22830 , w_22831 , w_22832 , w_22833 , w_22834 , w_22835 , 
		w_22836 , w_22837 , w_22838 , w_22839 , w_22840 , w_22841 , w_22842 , w_22843 , w_22844 , w_22845 , 
		w_22846 , w_22847 , w_22848 , w_22849 , w_22850 , w_22851 , w_22852 , w_22853 , w_22854 , w_22855 , 
		w_22856 , w_22857 , w_22858 , w_22859 , w_22860 , w_22861 , w_22862 , w_22863 , w_22864 , w_22865 , 
		w_22866 , w_22867 , w_22868 , w_22869 , w_22870 , w_22871 , w_22872 , w_22873 , w_22874 , w_22875 , 
		w_22876 , w_22877 , w_22878 , w_22879 , w_22880 , w_22881 , w_22882 , w_22883 , w_22884 , w_22885 , 
		w_22886 , w_22887 , w_22888 , w_22889 , w_22890 , w_22891 , w_22892 , w_22893 , w_22894 , w_22895 , 
		w_22896 , w_22897 , w_22898 , w_22899 , w_22900 , w_22901 , w_22902 , w_22903 , w_22904 , w_22905 , 
		w_22906 , w_22907 , w_22908 , w_22909 , w_22910 , w_22911 , w_22912 , w_22913 , w_22914 , w_22915 , 
		w_22916 , w_22917 , w_22918 , w_22919 , w_22920 , w_22921 , w_22922 , w_22923 , w_22924 , w_22925 , 
		w_22926 , w_22927 , w_22928 , w_22929 , w_22930 , w_22931 , w_22932 , w_22933 , w_22934 , w_22935 , 
		w_22936 , w_22937 , w_22938 , w_22939 , w_22940 , w_22941 , w_22942 , w_22943 , w_22944 , w_22945 , 
		w_22946 , w_22947 , w_22948 , w_22949 , w_22950 , w_22951 , w_22952 , w_22953 , w_22954 , w_22955 , 
		w_22956 , w_22957 , w_22958 , w_22959 , w_22960 , w_22961 , w_22962 , w_22963 , w_22964 , w_22965 , 
		w_22966 , w_22967 , w_22968 , w_22969 , w_22970 , w_22971 , w_22972 , w_22973 , w_22974 , w_22975 , 
		w_22976 , w_22977 , w_22978 , w_22979 , w_22980 , w_22981 , w_22982 , w_22983 , w_22984 , w_22985 , 
		w_22986 , w_22987 , w_22988 , w_22989 , w_22990 , w_22991 , w_22992 , w_22993 , w_22994 , w_22995 , 
		w_22996 , w_22997 , w_22998 , w_22999 , w_23000 , w_23001 , w_23002 , w_23003 , w_23004 , w_23005 , 
		w_23006 , w_23007 , w_23008 , w_23009 , w_23010 , w_23011 , w_23012 , w_23013 , w_23014 , w_23015 , 
		w_23016 , w_23017 , w_23018 , w_23019 , w_23020 , w_23021 , w_23022 , w_23023 , w_23024 , w_23025 , 
		w_23026 , w_23027 , w_23028 , w_23029 , w_23030 , w_23031 , w_23032 , w_23033 , w_23034 , w_23035 , 
		w_23036 , w_23037 , w_23038 , w_23039 , w_23040 , w_23041 , w_23042 , w_23043 , w_23044 , w_23045 , 
		w_23046 , w_23047 , w_23048 , w_23049 , w_23050 , w_23051 , w_23052 , w_23053 , w_23054 , w_23055 , 
		w_23056 , w_23057 , w_23058 , w_23059 , w_23060 , w_23061 , w_23062 , w_23063 , w_23064 , w_23065 , 
		w_23066 , w_23067 , w_23068 , w_23069 , w_23070 , w_23071 , w_23072 , w_23073 , w_23074 , w_23075 , 
		w_23076 , w_23077 , w_23078 , w_23079 , w_23080 , w_23081 , w_23082 , w_23083 , w_23084 , w_23085 , 
		w_23086 , w_23087 , w_23088 , w_23089 , w_23090 , w_23091 , w_23092 , w_23093 , w_23094 , w_23095 , 
		w_23096 , w_23097 , w_23098 , w_23099 , w_23100 , w_23101 , w_23102 , w_23103 , w_23104 , w_23105 , 
		w_23106 , w_23107 , w_23108 , w_23109 , w_23110 , w_23111 , w_23112 , w_23113 , w_23114 , w_23115 , 
		w_23116 , w_23117 , w_23118 , w_23119 , w_23120 , w_23121 , w_23122 , w_23123 , w_23124 , w_23125 , 
		w_23126 , w_23127 , w_23128 , w_23129 , w_23130 , w_23131 , w_23132 , w_23133 , w_23134 , w_23135 , 
		w_23136 , w_23137 , w_23138 , w_23139 , w_23140 , w_23141 , w_23142 , w_23143 , w_23144 , w_23145 , 
		w_23146 , w_23147 , w_23148 , w_23149 , w_23150 , w_23151 , w_23152 , w_23153 , w_23154 , w_23155 , 
		w_23156 , w_23157 , w_23158 , w_23159 , w_23160 , w_23161 , w_23162 , w_23163 , w_23164 , w_23165 , 
		w_23166 , w_23167 , w_23168 , w_23169 , w_23170 , w_23171 , w_23172 , w_23173 , w_23174 , w_23175 , 
		w_23176 , w_23177 , w_23178 , w_23179 , w_23180 , w_23181 , w_23182 , w_23183 , w_23184 , w_23185 , 
		w_23186 , w_23187 , w_23188 , w_23189 , w_23190 , w_23191 , w_23192 , w_23193 , w_23194 , w_23195 , 
		w_23196 , w_23197 , w_23198 , w_23199 , w_23200 , w_23201 , w_23202 , w_23203 , w_23204 , w_23205 , 
		w_23206 , w_23207 , w_23208 , w_23209 , w_23210 , w_23211 , w_23212 , w_23213 , w_23214 , w_23215 , 
		w_23216 , w_23217 , w_23218 , w_23219 , w_23220 , w_23221 , w_23222 , w_23223 , w_23224 , w_23225 , 
		w_23226 , w_23227 , w_23228 , w_23229 , w_23230 , w_23231 , w_23232 , w_23233 , w_23234 , w_23235 , 
		w_23236 , w_23237 , w_23238 , w_23239 , w_23240 , w_23241 , w_23242 , w_23243 , w_23244 , w_23245 , 
		w_23246 , w_23247 , w_23248 , w_23249 , w_23250 , w_23251 , w_23252 , w_23253 , w_23254 , w_23255 , 
		w_23256 , w_23257 , w_23258 , w_23259 , w_23260 , w_23261 , w_23262 , w_23263 , w_23264 , w_23265 , 
		w_23266 , w_23267 , w_23268 , w_23269 , w_23270 , w_23271 , w_23272 , w_23273 , w_23274 , w_23275 , 
		w_23276 , w_23277 , w_23278 , w_23279 , w_23280 , w_23281 , w_23282 , w_23283 , w_23284 , w_23285 , 
		w_23286 , w_23287 , w_23288 , w_23289 , w_23290 , w_23291 , w_23292 , w_23293 , w_23294 , w_23295 , 
		w_23296 , w_23297 , w_23298 , w_23299 , w_23300 , w_23301 , w_23302 , w_23303 , w_23304 , w_23305 , 
		w_23306 , w_23307 , w_23308 , w_23309 , w_23310 , w_23311 , w_23312 , w_23313 , w_23314 , w_23315 , 
		w_23316 , w_23317 , w_23318 , w_23319 , w_23320 , w_23321 , w_23322 , w_23323 , w_23324 , w_23325 , 
		w_23326 , w_23327 , w_23328 , w_23329 , w_23330 , w_23331 , w_23332 , w_23333 , w_23334 , w_23335 , 
		w_23336 , w_23337 , w_23338 , w_23339 , w_23340 , w_23341 , w_23342 , w_23343 , w_23344 , w_23345 , 
		w_23346 , w_23347 , w_23348 , w_23349 , w_23350 , w_23351 , w_23352 , w_23353 , w_23354 , w_23355 , 
		w_23356 , w_23357 , w_23358 , w_23359 , w_23360 , w_23361 , w_23362 , w_23363 , w_23364 , w_23365 , 
		w_23366 , w_23367 , w_23368 , w_23369 , w_23370 , w_23371 , w_23372 , w_23373 , w_23374 , w_23375 , 
		w_23376 , w_23377 , w_23378 , w_23379 , w_23380 , w_23381 , w_23382 , w_23383 , w_23384 , w_23385 , 
		w_23386 , w_23387 , w_23388 , w_23389 , w_23390 , w_23391 , w_23392 , w_23393 , w_23394 , w_23395 , 
		w_23396 , w_23397 , w_23398 , w_23399 , w_23400 , w_23401 , w_23402 , w_23403 , w_23404 , w_23405 , 
		w_23406 , w_23407 , w_23408 , w_23409 , w_23410 , w_23411 , w_23412 , w_23413 , w_23414 , w_23415 , 
		w_23416 , w_23417 , w_23418 , w_23419 , w_23420 , w_23421 , w_23422 , w_23423 , w_23424 , w_23425 , 
		w_23426 , w_23427 , w_23428 , w_23429 , w_23430 , w_23431 , w_23432 , w_23433 , w_23434 , w_23435 , 
		w_23436 , w_23437 , w_23438 , w_23439 , w_23440 , w_23441 , w_23442 , w_23443 , w_23444 , w_23445 , 
		w_23446 , w_23447 , w_23448 , w_23449 , w_23450 , w_23451 , w_23452 , w_23453 , w_23454 , w_23455 , 
		w_23456 , w_23457 , w_23458 , w_23459 , w_23460 , w_23461 , w_23462 , w_23463 , w_23464 , w_23465 , 
		w_23466 , w_23467 , w_23468 , w_23469 , w_23470 , w_23471 , w_23472 , w_23473 , w_23474 , w_23475 , 
		w_23476 , w_23477 , w_23478 , w_23479 , w_23480 , w_23481 , w_23482 , w_23483 , w_23484 , w_23485 , 
		w_23486 , w_23487 , w_23488 , w_23489 , w_23490 , w_23491 , w_23492 , w_23493 , w_23494 , w_23495 , 
		w_23496 , w_23497 , w_23498 , w_23499 , w_23500 , w_23501 , w_23502 , w_23503 , w_23504 , w_23505 , 
		w_23506 , w_23507 , w_23508 , w_23509 , w_23510 , w_23511 , w_23512 , w_23513 , w_23514 , w_23515 , 
		w_23516 , w_23517 , w_23518 , w_23519 , w_23520 , w_23521 , w_23522 , w_23523 , w_23524 , w_23525 , 
		w_23526 , w_23527 , w_23528 , w_23529 , w_23530 , w_23531 , w_23532 , w_23533 , w_23534 , w_23535 , 
		w_23536 , w_23537 , w_23538 , w_23539 , w_23540 , w_23541 , w_23542 , w_23543 , w_23544 , w_23545 , 
		w_23546 , w_23547 , w_23548 , w_23549 , w_23550 , w_23551 , w_23552 , w_23553 , w_23554 , w_23555 , 
		w_23556 , w_23557 , w_23558 , w_23559 , w_23560 , w_23561 , w_23562 , w_23563 , w_23564 , w_23565 , 
		w_23566 , w_23567 , w_23568 , w_23569 , w_23570 , w_23571 , w_23572 , w_23573 , w_23574 , w_23575 , 
		w_23576 , w_23577 , w_23578 , w_23579 , w_23580 , w_23581 , w_23582 , w_23583 , w_23584 , w_23585 , 
		w_23586 , w_23587 , w_23588 , w_23589 , w_23590 , w_23591 , w_23592 , w_23593 , w_23594 , w_23595 , 
		w_23596 , w_23597 , w_23598 , w_23599 , w_23600 , w_23601 , w_23602 , w_23603 , w_23604 , w_23605 , 
		w_23606 , w_23607 , w_23608 , w_23609 , w_23610 , w_23611 , w_23612 , w_23613 , w_23614 , w_23615 , 
		w_23616 , w_23617 , w_23618 , w_23619 , w_23620 , w_23621 , w_23622 , w_23623 , w_23624 , w_23625 , 
		w_23626 , w_23627 , w_23628 , w_23629 , w_23630 , w_23631 , w_23632 , w_23633 , w_23634 , w_23635 , 
		w_23636 , w_23637 , w_23638 , w_23639 , w_23640 , w_23641 , w_23642 , w_23643 , w_23644 , w_23645 , 
		w_23646 , w_23647 , w_23648 , w_23649 , w_23650 , w_23651 , w_23652 , w_23653 , w_23654 , w_23655 , 
		w_23656 , w_23657 , w_23658 , w_23659 , w_23660 , w_23661 , w_23662 , w_23663 , w_23664 , w_23665 , 
		w_23666 , w_23667 , w_23668 , w_23669 , w_23670 , w_23671 , w_23672 , w_23673 , w_23674 , w_23675 , 
		w_23676 , w_23677 , w_23678 , w_23679 , w_23680 , w_23681 , w_23682 , w_23683 , w_23684 , w_23685 , 
		w_23686 , w_23687 , w_23688 , w_23689 , w_23690 , w_23691 , w_23692 , w_23693 , w_23694 , w_23695 , 
		w_23696 , w_23697 , w_23698 , w_23699 , w_23700 , w_23701 , w_23702 , w_23703 , w_23704 , w_23705 , 
		w_23706 , w_23707 , w_23708 , w_23709 , w_23710 , w_23711 , w_23712 , w_23713 , w_23714 , w_23715 , 
		w_23716 , w_23717 , w_23718 , w_23719 , w_23720 , w_23721 , w_23722 , w_23723 , w_23724 , w_23725 , 
		w_23726 , w_23727 , w_23728 , w_23729 , w_23730 , w_23731 , w_23732 , w_23733 , w_23734 , w_23735 , 
		w_23736 , w_23737 , w_23738 , w_23739 , w_23740 , w_23741 , w_23742 , w_23743 , w_23744 , w_23745 , 
		w_23746 , w_23747 , w_23748 , w_23749 , w_23750 , w_23751 , w_23752 , w_23753 , w_23754 , w_23755 , 
		w_23756 , w_23757 , w_23758 , w_23759 , w_23760 , w_23761 , w_23762 , w_23763 , w_23764 , w_23765 , 
		w_23766 , w_23767 , w_23768 , w_23769 , w_23770 , w_23771 , w_23772 , w_23773 , w_23774 , w_23775 , 
		w_23776 , w_23777 , w_23778 , w_23779 , w_23780 , w_23781 , w_23782 , w_23783 , w_23784 , w_23785 , 
		w_23786 , w_23787 , w_23788 , w_23789 , w_23790 , w_23791 , w_23792 , w_23793 , w_23794 , w_23795 , 
		w_23796 , w_23797 , w_23798 , w_23799 , w_23800 , w_23801 , w_23802 , w_23803 , w_23804 , w_23805 , 
		w_23806 , w_23807 , w_23808 , w_23809 , w_23810 , w_23811 , w_23812 , w_23813 , w_23814 , w_23815 , 
		w_23816 , w_23817 , w_23818 , w_23819 , w_23820 , w_23821 , w_23822 , w_23823 , w_23824 , w_23825 , 
		w_23826 , w_23827 , w_23828 , w_23829 , w_23830 , w_23831 , w_23832 , w_23833 , w_23834 , w_23835 , 
		w_23836 , w_23837 , w_23838 , w_23839 , w_23840 , w_23841 , w_23842 , w_23843 , w_23844 , w_23845 , 
		w_23846 , w_23847 , w_23848 , w_23849 , w_23850 , w_23851 , w_23852 , w_23853 , w_23854 , w_23855 , 
		w_23856 , w_23857 , w_23858 , w_23859 , w_23860 , w_23861 , w_23862 , w_23863 , w_23864 , w_23865 , 
		w_23866 , w_23867 , w_23868 , w_23869 , w_23870 , w_23871 , w_23872 , w_23873 , w_23874 , w_23875 , 
		w_23876 , w_23877 , w_23878 , w_23879 , w_23880 , w_23881 , w_23882 , w_23883 , w_23884 , w_23885 , 
		w_23886 , w_23887 , w_23888 , w_23889 , w_23890 , w_23891 , w_23892 , w_23893 , w_23894 , w_23895 , 
		w_23896 , w_23897 , w_23898 , w_23899 , w_23900 , w_23901 , w_23902 , w_23903 , w_23904 , w_23905 , 
		w_23906 , w_23907 , w_23908 , w_23909 , w_23910 , w_23911 , w_23912 , w_23913 , w_23914 , w_23915 , 
		w_23916 , w_23917 , w_23918 , w_23919 , w_23920 , w_23921 , w_23922 , w_23923 , w_23924 , w_23925 , 
		w_23926 , w_23927 , w_23928 , w_23929 , w_23930 , w_23931 , w_23932 , w_23933 , w_23934 , w_23935 , 
		w_23936 , w_23937 , w_23938 , w_23939 , w_23940 , w_23941 , w_23942 , w_23943 , w_23944 , w_23945 , 
		w_23946 , w_23947 , w_23948 , w_23949 , w_23950 , w_23951 , w_23952 , w_23953 , w_23954 , w_23955 , 
		w_23956 , w_23957 , w_23958 , w_23959 , w_23960 , w_23961 , w_23962 , w_23963 , w_23964 , w_23965 , 
		w_23966 , w_23967 , w_23968 , w_23969 , w_23970 , w_23971 , w_23972 , w_23973 , w_23974 , w_23975 , 
		w_23976 , w_23977 , w_23978 , w_23979 , w_23980 , w_23981 , w_23982 , w_23983 , w_23984 , w_23985 , 
		w_23986 , w_23987 , w_23988 , w_23989 , w_23990 , w_23991 , w_23992 , w_23993 , w_23994 , w_23995 , 
		w_23996 , w_23997 , w_23998 , w_23999 , w_24000 , w_24001 , w_24002 , w_24003 , w_24004 , w_24005 , 
		w_24006 , w_24007 , w_24008 , w_24009 , w_24010 , w_24011 , w_24012 , w_24013 , w_24014 , w_24015 , 
		w_24016 , w_24017 , w_24018 , w_24019 , w_24020 , w_24021 , w_24022 , w_24023 , w_24024 , w_24025 , 
		w_24026 , w_24027 , w_24028 , w_24029 , w_24030 , w_24031 , w_24032 , w_24033 , w_24034 , w_24035 , 
		w_24036 , w_24037 , w_24038 , w_24039 , w_24040 , w_24041 , w_24042 , w_24043 , w_24044 , w_24045 , 
		w_24046 , w_24047 , w_24048 , w_24049 , w_24050 , w_24051 , w_24052 , w_24053 , w_24054 , w_24055 , 
		w_24056 , w_24057 , w_24058 , w_24059 , w_24060 , w_24061 , w_24062 , w_24063 , w_24064 , w_24065 , 
		w_24066 , w_24067 , w_24068 , w_24069 , w_24070 , w_24071 , w_24072 , w_24073 , w_24074 , w_24075 , 
		w_24076 , w_24077 , w_24078 , w_24079 , w_24080 , w_24081 , w_24082 , w_24083 , w_24084 , w_24085 , 
		w_24086 , w_24087 , w_24088 , w_24089 , w_24090 , w_24091 , w_24092 , w_24093 , w_24094 , w_24095 , 
		w_24096 , w_24097 , w_24098 , w_24099 , w_24100 , w_24101 , w_24102 , w_24103 , w_24104 , w_24105 , 
		w_24106 , w_24107 , w_24108 , w_24109 , w_24110 , w_24111 , w_24112 , w_24113 , w_24114 , w_24115 , 
		w_24116 , w_24117 , w_24118 , w_24119 , w_24120 , w_24121 , w_24122 , w_24123 , w_24124 , w_24125 , 
		w_24126 , w_24127 , w_24128 , w_24129 , w_24130 , w_24131 , w_24132 , w_24133 , w_24134 , w_24135 , 
		w_24136 , w_24137 , w_24138 , w_24139 , w_24140 , w_24141 , w_24142 , w_24143 , w_24144 , w_24145 , 
		w_24146 , w_24147 , w_24148 , w_24149 , w_24150 , w_24151 , w_24152 , w_24153 , w_24154 , w_24155 , 
		w_24156 , w_24157 , w_24158 , w_24159 , w_24160 , w_24161 , w_24162 , w_24163 , w_24164 , w_24165 , 
		w_24166 , w_24167 , w_24168 , w_24169 , w_24170 , w_24171 , w_24172 , w_24173 , w_24174 , w_24175 , 
		w_24176 , w_24177 , w_24178 , w_24179 , w_24180 , w_24181 , w_24182 , w_24183 , w_24184 , w_24185 , 
		w_24186 , w_24187 , w_24188 , w_24189 , w_24190 , w_24191 , w_24192 , w_24193 , w_24194 , w_24195 , 
		w_24196 , w_24197 , w_24198 , w_24199 , w_24200 , w_24201 , w_24202 , w_24203 , w_24204 , w_24205 , 
		w_24206 , w_24207 , w_24208 , w_24209 , w_24210 , w_24211 , w_24212 , w_24213 , w_24214 , w_24215 , 
		w_24216 , w_24217 , w_24218 , w_24219 , w_24220 , w_24221 , w_24222 , w_24223 , w_24224 , w_24225 , 
		w_24226 , w_24227 , w_24228 , w_24229 , w_24230 , w_24231 , w_24232 , w_24233 , w_24234 , w_24235 , 
		w_24236 , w_24237 , w_24238 , w_24239 , w_24240 , w_24241 , w_24242 , w_24243 , w_24244 , w_24245 , 
		w_24246 , w_24247 , w_24248 , w_24249 , w_24250 , w_24251 , w_24252 , w_24253 , w_24254 , w_24255 , 
		w_24256 , w_24257 , w_24258 , w_24259 , w_24260 , w_24261 , w_24262 , w_24263 , w_24264 , w_24265 , 
		w_24266 , w_24267 , w_24268 , w_24269 , w_24270 , w_24271 , w_24272 , w_24273 , w_24274 , w_24275 , 
		w_24276 , w_24277 , w_24278 , w_24279 , w_24280 , w_24281 , w_24282 , w_24283 , w_24284 , w_24285 , 
		w_24286 , w_24287 , w_24288 , w_24289 , w_24290 , w_24291 , w_24292 , w_24293 , w_24294 , w_24295 , 
		w_24296 , w_24297 , w_24298 , w_24299 , w_24300 , w_24301 , w_24302 , w_24303 , w_24304 , w_24305 , 
		w_24306 , w_24307 , w_24308 , w_24309 , w_24310 , w_24311 , w_24312 , w_24313 , w_24314 , w_24315 , 
		w_24316 , w_24317 , w_24318 , w_24319 , w_24320 , w_24321 , w_24322 , w_24323 , w_24324 , w_24325 , 
		w_24326 , w_24327 , w_24328 , w_24329 , w_24330 , w_24331 , w_24332 , w_24333 , w_24334 , w_24335 , 
		w_24336 , w_24337 , w_24338 , w_24339 , w_24340 , w_24341 , w_24342 , w_24343 , w_24344 , w_24345 , 
		w_24346 , w_24347 , w_24348 , w_24349 , w_24350 , w_24351 , w_24352 , w_24353 , w_24354 , w_24355 , 
		w_24356 , w_24357 , w_24358 , w_24359 , w_24360 , w_24361 , w_24362 , w_24363 , w_24364 , w_24365 , 
		w_24366 , w_24367 , w_24368 , w_24369 , w_24370 , w_24371 , w_24372 , w_24373 , w_24374 , w_24375 , 
		w_24376 , w_24377 , w_24378 , w_24379 , w_24380 , w_24381 , w_24382 , w_24383 , w_24384 , w_24385 , 
		w_24386 , w_24387 , w_24388 , w_24389 , w_24390 , w_24391 , w_24392 , w_24393 , w_24394 , w_24395 , 
		w_24396 , w_24397 , w_24398 , w_24399 , w_24400 , w_24401 , w_24402 , w_24403 , w_24404 , w_24405 , 
		w_24406 , w_24407 , w_24408 , w_24409 , w_24410 , w_24411 , w_24412 , w_24413 , w_24414 , w_24415 , 
		w_24416 , w_24417 , w_24418 , w_24419 , w_24420 , w_24421 , w_24422 , w_24423 , w_24424 , w_24425 , 
		w_24426 , w_24427 , w_24428 , w_24429 , w_24430 , w_24431 , w_24432 , w_24433 , w_24434 , w_24435 , 
		w_24436 , w_24437 , w_24438 , w_24439 , w_24440 , w_24441 , w_24442 , w_24443 , w_24444 , w_24445 , 
		w_24446 , w_24447 , w_24448 , w_24449 , w_24450 , w_24451 , w_24452 , w_24453 , w_24454 , w_24455 , 
		w_24456 , w_24457 , w_24458 , w_24459 , w_24460 , w_24461 , w_24462 , w_24463 , w_24464 , w_24465 , 
		w_24466 , w_24467 , w_24468 , w_24469 , w_24470 , w_24471 , w_24472 , w_24473 , w_24474 , w_24475 , 
		w_24476 , w_24477 , w_24478 , w_24479 , w_24480 , w_24481 , w_24482 , w_24483 , w_24484 , w_24485 , 
		w_24486 , w_24487 , w_24488 , w_24489 , w_24490 , w_24491 , w_24492 , w_24493 , w_24494 , w_24495 , 
		w_24496 , w_24497 , w_24498 , w_24499 , w_24500 , w_24501 , w_24502 , w_24503 , w_24504 , w_24505 , 
		w_24506 , w_24507 , w_24508 , w_24509 , w_24510 , w_24511 , w_24512 , w_24513 , w_24514 , w_24515 , 
		w_24516 , w_24517 , w_24518 , w_24519 , w_24520 , w_24521 , w_24522 , w_24523 , w_24524 , w_24525 , 
		w_24526 , w_24527 , w_24528 , w_24529 , w_24530 , w_24531 , w_24532 , w_24533 , w_24534 , w_24535 , 
		w_24536 , w_24537 , w_24538 , w_24539 , w_24540 , w_24541 , w_24542 , w_24543 , w_24544 , w_24545 , 
		w_24546 , w_24547 , w_24548 , w_24549 , w_24550 , w_24551 , w_24552 , w_24553 , w_24554 , w_24555 , 
		w_24556 , w_24557 , w_24558 , w_24559 , w_24560 , w_24561 , w_24562 , w_24563 , w_24564 , w_24565 , 
		w_24566 , w_24567 , w_24568 , w_24569 , w_24570 , w_24571 , w_24572 , w_24573 , w_24574 , w_24575 , 
		w_24576 , w_24577 , w_24578 , w_24579 , w_24580 , w_24581 , w_24582 , w_24583 , w_24584 , w_24585 , 
		w_24586 , w_24587 , w_24588 , w_24589 , w_24590 , w_24591 , w_24592 , w_24593 , w_24594 , w_24595 , 
		w_24596 , w_24597 , w_24598 , w_24599 , w_24600 , w_24601 , w_24602 , w_24603 , w_24604 , w_24605 , 
		w_24606 , w_24607 , w_24608 , w_24609 , w_24610 , w_24611 , w_24612 , w_24613 , w_24614 , w_24615 , 
		w_24616 , w_24617 , w_24618 , w_24619 , w_24620 , w_24621 , w_24622 , w_24623 , w_24624 , w_24625 , 
		w_24626 , w_24627 , w_24628 , w_24629 , w_24630 , w_24631 , w_24632 , w_24633 , w_24634 , w_24635 , 
		w_24636 , w_24637 , w_24638 , w_24639 , w_24640 , w_24641 , w_24642 , w_24643 , w_24644 , w_24645 , 
		w_24646 , w_24647 , w_24648 , w_24649 , w_24650 , w_24651 , w_24652 , w_24653 , w_24654 , w_24655 , 
		w_24656 , w_24657 , w_24658 , w_24659 , w_24660 , w_24661 , w_24662 , w_24663 , w_24664 , w_24665 , 
		w_24666 , w_24667 , w_24668 , w_24669 , w_24670 , w_24671 , w_24672 , w_24673 , w_24674 , w_24675 , 
		w_24676 , w_24677 , w_24678 , w_24679 , w_24680 , w_24681 , w_24682 , w_24683 , w_24684 , w_24685 , 
		w_24686 , w_24687 , w_24688 , w_24689 , w_24690 , w_24691 , w_24692 , w_24693 , w_24694 , w_24695 , 
		w_24696 , w_24697 , w_24698 , w_24699 , w_24700 , w_24701 , w_24702 , w_24703 , w_24704 , w_24705 , 
		w_24706 , w_24707 , w_24708 , w_24709 , w_24710 , w_24711 , w_24712 , w_24713 , w_24714 , w_24715 , 
		w_24716 , w_24717 , w_24718 , w_24719 , w_24720 , w_24721 , w_24722 , w_24723 , w_24724 , w_24725 , 
		w_24726 , w_24727 , w_24728 , w_24729 , w_24730 , w_24731 , w_24732 , w_24733 , w_24734 , w_24735 , 
		w_24736 , w_24737 , w_24738 , w_24739 , w_24740 , w_24741 , w_24742 , w_24743 , w_24744 , w_24745 , 
		w_24746 , w_24747 , w_24748 , w_24749 , w_24750 , w_24751 , w_24752 , w_24753 , w_24754 , w_24755 , 
		w_24756 , w_24757 , w_24758 , w_24759 , w_24760 , w_24761 , w_24762 , w_24763 , w_24764 , w_24765 , 
		w_24766 , w_24767 , w_24768 , w_24769 , w_24770 , w_24771 , w_24772 , w_24773 , w_24774 , w_24775 , 
		w_24776 , w_24777 , w_24778 , w_24779 , w_24780 , w_24781 , w_24782 , w_24783 , w_24784 , w_24785 , 
		w_24786 , w_24787 , w_24788 , w_24789 , w_24790 , w_24791 , w_24792 , w_24793 , w_24794 , w_24795 , 
		w_24796 , w_24797 , w_24798 , w_24799 , w_24800 , w_24801 , w_24802 , w_24803 , w_24804 , w_24805 , 
		w_24806 , w_24807 , w_24808 , w_24809 , w_24810 , w_24811 , w_24812 , w_24813 , w_24814 , w_24815 , 
		w_24816 , w_24817 , w_24818 , w_24819 , w_24820 , w_24821 , w_24822 , w_24823 , w_24824 , w_24825 , 
		w_24826 , w_24827 , w_24828 , w_24829 , w_24830 , w_24831 , w_24832 , w_24833 , w_24834 , w_24835 , 
		w_24836 , w_24837 , w_24838 , w_24839 , w_24840 , w_24841 , w_24842 , w_24843 , w_24844 , w_24845 , 
		w_24846 , w_24847 , w_24848 , w_24849 , w_24850 , w_24851 , w_24852 , w_24853 , w_24854 , w_24855 , 
		w_24856 , w_24857 , w_24858 , w_24859 , w_24860 , w_24861 , w_24862 , w_24863 , w_24864 , w_24865 , 
		w_24866 , w_24867 , w_24868 , w_24869 , w_24870 , w_24871 , w_24872 , w_24873 , w_24874 , w_24875 , 
		w_24876 , w_24877 , w_24878 , w_24879 , w_24880 , w_24881 , w_24882 , w_24883 , w_24884 , w_24885 , 
		w_24886 , w_24887 , w_24888 , w_24889 , w_24890 , w_24891 , w_24892 , w_24893 , w_24894 , w_24895 , 
		w_24896 , w_24897 , w_24898 , w_24899 , w_24900 , w_24901 , w_24902 , w_24903 , w_24904 , w_24905 , 
		w_24906 , w_24907 , w_24908 , w_24909 , w_24910 , w_24911 , w_24912 , w_24913 , w_24914 , w_24915 , 
		w_24916 , w_24917 , w_24918 , w_24919 , w_24920 , w_24921 , w_24922 , w_24923 , w_24924 , w_24925 , 
		w_24926 , w_24927 ;
buf ( \o[31]_b1 , \7238_b1 );
buf ( \o[31]_b0 , \7238_b0 );
buf ( \o[30]_b1 , \7251_b1 );
buf ( \o[30]_b0 , \7251_b0 );
buf ( \o[29]_b1 , \7262_b1 );
buf ( \o[29]_b0 , \7262_b0 );
buf ( \o[28]_b1 , \7274_b1 );
buf ( \o[28]_b0 , \7274_b0 );
buf ( \o[27]_b1 , \7288_b1 );
buf ( \o[27]_b0 , \7288_b0 );
buf ( \o[26]_b1 , \7300_b1 );
buf ( \o[26]_b0 , \7300_b0 );
buf ( \o[25]_b1 , \7311_b1 );
buf ( \o[25]_b0 , \7311_b0 );
buf ( \o[24]_b1 , \7343_b1 );
buf ( \o[24]_b0 , \7343_b0 );
buf ( \o[23]_b1 , \7337_b1 );
buf ( \o[23]_b0 , \7337_b0 );
buf ( \o[22]_b1 , \7508_b1 );
buf ( \o[22]_b0 , \7508_b0 );
buf ( \o[21]_b1 , \7354_b1 );
buf ( \o[21]_b0 , \7354_b0 );
buf ( \o[20]_b1 , \7360_b1 );
buf ( \o[20]_b0 , \7360_b0 );
buf ( \o[19]_b1 , \7375_b1 );
buf ( \o[19]_b0 , \7375_b0 );
buf ( \o[18]_b1 , \7381_b1 );
buf ( \o[18]_b0 , \7381_b0 );
buf ( \o[17]_b1 , \7392_b1 );
buf ( \o[17]_b0 , \7392_b0 );
buf ( \o[16]_b1 , \7398_b1 );
buf ( \o[16]_b0 , \7398_b0 );
buf ( \o[15]_b1 , \7418_b1 );
buf ( \o[15]_b0 , \7418_b0 );
buf ( \o[14]_b1 , \7426_b1 );
buf ( \o[14]_b0 , \7426_b0 );
buf ( \o[13]_b1 , \7436_b1 );
buf ( \o[13]_b0 , \7436_b0 );
buf ( \o[12]_b1 , \7458_b1 );
buf ( \o[12]_b0 , \7458_b0 );
buf ( \o[11]_b1 , \7452_b1 );
buf ( \o[11]_b0 , \7452_b0 );
buf ( \o[10]_b1 , \7464_b1 );
buf ( \o[10]_b0 , \7464_b0 );
buf ( \o[9]_b1 , \7474_b1 );
buf ( \o[9]_b0 , \7474_b0 );
buf ( \o[8]_b1 , \7480_b1 );
buf ( \o[8]_b0 , \7480_b0 );
buf ( \o[7]_b1 , \7482_b1 );
buf ( \o[7]_b0 , \7482_b0 );
buf ( \o[6]_b1 , \7507_b1 );
buf ( \o[6]_b0 , \7507_b0 );
buf ( \o[5]_b1 , \7488_b1 );
buf ( \o[5]_b0 , \7488_b0 );
buf ( \o[4]_b1 , \7495_b1 );
buf ( \o[4]_b0 , \7495_b0 );
buf ( \o[3]_b1 , \7497_b1 );
buf ( \o[3]_b0 , \7497_b0 );
buf ( \o[2]_b1 , \7502_b1 );
buf ( \o[2]_b0 , \7502_b0 );
buf ( \o[1]_b1 , \7505_b1 );
buf ( \o[1]_b0 , \7505_b0 );
buf ( \o[0]_b1 , \7506_b1 );
buf ( \o[0]_b0 , \7506_b0 );
buf ( \99_b1 , \d[15]_b1 );
not ( \99_b1 , w_0 );
not ( \99_b0 , w_1 );
and ( w_0 , w_1 , \d[15]_b0 );
or ( \100_b1 , \b[3]_b1 , \a[2]_b1 );
xor ( \100_b0 , \b[3]_b0 , w_2 );
not ( w_2 , w_3 );
and ( w_3 , \a[2]_b1 , \a[2]_b0 );
buf ( \101_b1 , \100_b1 );
not ( \101_b1 , w_4 );
not ( \101_b0 , w_5 );
and ( w_4 , w_5 , \100_b0 );
or ( \102_b1 , \b[3]_b1 , w_6 );
xor ( \102_b0 , \b[3]_b0 , w_8 );
not ( w_8 , w_9 );
and ( w_9 , w_6 , w_7 );
buf ( w_6 , \b[2]_b1 );
not ( w_6 , w_10 );
not ( w_7 , w_11 );
and ( w_10 , w_11 , \b[2]_b0 );
or ( \103_b1 , \b[2]_b1 , \b[1]_b1 );
xor ( \103_b0 , \b[2]_b0 , w_12 );
not ( w_12 , w_13 );
and ( w_13 , \b[1]_b1 , \b[1]_b0 );
or ( \104_b1 , \102_b1 , w_15 );
not ( w_15 , w_16 );
and ( \104_b0 , \102_b0 , w_17 );
and ( w_16 ,  , w_17 );
buf ( w_15 , \103_b1 );
not ( w_15 , w_18 );
not (  , w_19 );
and ( w_18 , w_19 , \103_b0 );
buf ( \105_b1 , \104_b1 );
not ( \105_b1 , w_20 );
not ( \105_b0 , w_21 );
and ( w_20 , w_21 , \104_b0 );
or ( \106_b1 , \101_b1 , w_22 );
or ( \106_b0 , \101_b0 , \105_b0 );
not ( \105_b0 , w_23 );
and ( w_23 , w_22 , \105_b1 );
or ( \107_b1 , \b[3]_b1 , \a[3]_b1 );
xor ( \107_b0 , \b[3]_b0 , w_24 );
not ( w_24 , w_25 );
and ( w_25 , \a[3]_b1 , \a[3]_b0 );
or ( \108_b1 , \103_b1 , w_27 );
not ( w_27 , w_28 );
and ( \108_b0 , \103_b0 , w_29 );
and ( w_28 ,  , w_29 );
buf ( w_27 , \107_b1 );
not ( w_27 , w_30 );
not (  , w_31 );
and ( w_30 , w_31 , \107_b0 );
or ( \109_b1 , \106_b1 , w_33 );
not ( w_33 , w_34 );
and ( \109_b0 , \106_b0 , w_35 );
and ( w_34 ,  , w_35 );
buf ( w_33 , \108_b1 );
not ( w_33 , w_36 );
not (  , w_37 );
and ( w_36 , w_37 , \108_b0 );
or ( \110_b1 , \a[0]_b1 , w_38 );
or ( \110_b0 , \a[0]_b0 , \b[4]_b0 );
not ( \b[4]_b0 , w_39 );
and ( w_39 , w_38 , \b[4]_b1 );
or ( \111_b1 , \110_b1 , w_41 );
not ( w_41 , w_42 );
and ( \111_b0 , \110_b0 , w_43 );
and ( w_42 ,  , w_43 );
buf ( w_41 , \b[3]_b1 );
not ( w_41 , w_44 );
not (  , w_45 );
and ( w_44 , w_45 , \b[3]_b0 );
or ( \112_b1 , \a[0]_b1 , w_47 );
not ( w_47 , w_48 );
and ( \112_b0 , \a[0]_b0 , w_49 );
and ( w_48 ,  , w_49 );
buf ( w_47 , \b[4]_b1 );
not ( w_47 , w_50 );
not (  , w_51 );
and ( w_50 , w_51 , \b[4]_b0 );
buf ( \114_b1 , \113_b1 );
not ( \114_b1 , w_52 );
not ( \114_b0 , w_53 );
and ( w_52 , w_53 , \113_b0 );
or ( \115_b1 , \109_b1 , \114_b1 );
not ( \114_b1 , w_54 );
and ( \115_b0 , \109_b0 , w_55 );
and ( w_54 , w_55 , \114_b0 );
buf ( \116_b1 , \115_b1 );
not ( \116_b1 , w_56 );
not ( \116_b0 , w_57 );
and ( w_56 , w_57 , \115_b0 );
or ( \117_b1 , \a[5]_b1 , \b[1]_b1 );
xor ( \117_b0 , \a[5]_b0 , w_58 );
not ( w_58 , w_59 );
and ( w_59 , \b[1]_b1 , \b[1]_b0 );
buf ( \118_b1 , \117_b1 );
not ( \118_b1 , w_60 );
not ( \118_b0 , w_61 );
and ( w_60 , w_61 , \117_b0 );
buf ( \119_b1 , \b[1]_b1 );
not ( \119_b1 , w_62 );
not ( \119_b0 , w_63 );
and ( w_62 , w_63 , \b[1]_b0 );
or ( \120_b1 , \119_b1 , w_65 );
not ( w_65 , w_66 );
and ( \120_b0 , \119_b0 , w_67 );
and ( w_66 ,  , w_67 );
buf ( w_65 , \b[0]_b1 );
not ( w_65 , w_68 );
not (  , w_69 );
and ( w_68 , w_69 , \b[0]_b0 );
buf ( \121_b1 , \120_b1 );
not ( \121_b1 , w_70 );
not ( \121_b0 , w_71 );
and ( w_70 , w_71 , \120_b0 );
or ( \122_b1 , \118_b1 , w_72 );
or ( \122_b0 , \118_b0 , \121_b0 );
not ( \121_b0 , w_73 );
and ( w_73 , w_72 , \121_b1 );
or ( \123_b1 , \a[6]_b1 , \b[1]_b1 );
xor ( \123_b0 , \a[6]_b0 , w_74 );
not ( w_74 , w_75 );
and ( w_75 , \b[1]_b1 , \b[1]_b0 );
or ( \124_b1 , \123_b1 , w_77 );
not ( w_77 , w_78 );
and ( \124_b0 , \123_b0 , w_79 );
and ( w_78 ,  , w_79 );
buf ( w_77 , \b[0]_b1 );
not ( w_77 , w_80 );
not (  , w_81 );
and ( w_80 , w_81 , \b[0]_b0 );
or ( \125_b1 , \122_b1 , w_83 );
not ( w_83 , w_84 );
and ( \125_b0 , \122_b0 , w_85 );
and ( w_84 ,  , w_85 );
buf ( w_83 , \124_b1 );
not ( w_83 , w_86 );
not (  , w_87 );
and ( w_86 , w_87 , \124_b0 );
buf ( \126_b1 , \125_b1 );
not ( \126_b1 , w_88 );
not ( \126_b0 , w_89 );
and ( w_88 , w_89 , \125_b0 );
or ( \127_b1 , \116_b1 , w_91 );
not ( w_91 , w_92 );
and ( \127_b0 , \116_b0 , w_93 );
and ( w_92 ,  , w_93 );
buf ( w_91 , \126_b1 );
not ( w_91 , w_94 );
not (  , w_95 );
and ( w_94 , w_95 , \126_b0 );
buf ( \128_b1 , \127_b1 );
not ( \128_b1 , w_96 );
not ( \128_b0 , w_97 );
and ( w_96 , w_97 , \127_b0 );
or ( \129_b1 , \b[6]_b1 , \b[5]_b1 );
xor ( \129_b0 , \b[6]_b0 , w_98 );
not ( w_98 , w_99 );
and ( w_99 , \b[5]_b1 , \b[5]_b0 );
or ( \130_b1 , \129_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_100 );
and ( \130_b0 , \129_b0 , w_101 );
and ( w_100 , w_101 , \a[0]_b0 );
or ( \131_b1 , \a[1]_b1 , \b[5]_b1 );
xor ( \131_b0 , \a[1]_b0 , w_102 );
not ( w_102 , w_103 );
and ( w_103 , \b[5]_b1 , \b[5]_b0 );
buf ( \132_b1 , \131_b1 );
not ( \132_b1 , w_104 );
not ( \132_b0 , w_105 );
and ( w_104 , w_105 , \131_b0 );
or ( \133_b1 , \b[5]_b1 , \b[4]_b1 );
xor ( \133_b0 , \b[5]_b0 , w_106 );
not ( w_106 , w_107 );
and ( w_107 , \b[4]_b1 , \b[4]_b0 );
buf ( \134_b1 , \133_b1 );
not ( \134_b1 , w_108 );
not ( \134_b0 , w_109 );
and ( w_108 , w_109 , \133_b0 );
or ( \135_b1 , \b[4]_b1 , \b[3]_b1 );
xor ( \135_b0 , \b[4]_b0 , w_110 );
not ( w_110 , w_111 );
and ( w_111 , \b[3]_b1 , \b[3]_b0 );
or ( \136_b1 , \134_b1 , w_113 );
not ( w_113 , w_114 );
and ( \136_b0 , \134_b0 , w_115 );
and ( w_114 ,  , w_115 );
buf ( w_113 , \135_b1 );
not ( w_113 , w_116 );
not (  , w_117 );
and ( w_116 , w_117 , \135_b0 );
buf ( \137_b1 , \136_b1 );
not ( \137_b1 , w_118 );
not ( \137_b0 , w_119 );
and ( w_118 , w_119 , \136_b0 );
or ( \138_b1 , \132_b1 , w_120 );
or ( \138_b0 , \132_b0 , \137_b0 );
not ( \137_b0 , w_121 );
and ( w_121 , w_120 , \137_b1 );
or ( \139_b1 , \b[4]_b1 , \b[3]_b1 );
xor ( \139_b0 , \b[4]_b0 , w_122 );
not ( w_122 , w_123 );
and ( w_123 , \b[3]_b1 , \b[3]_b0 );
or ( \140_b1 , \a[2]_b1 , \b[5]_b1 );
xor ( \140_b0 , \a[2]_b0 , w_124 );
not ( w_124 , w_125 );
and ( w_125 , \b[5]_b1 , \b[5]_b0 );
or ( \141_b1 , \139_b1 , w_127 );
not ( w_127 , w_128 );
and ( \141_b0 , \139_b0 , w_129 );
and ( w_128 ,  , w_129 );
buf ( w_127 , \140_b1 );
not ( w_127 , w_130 );
not (  , w_131 );
and ( w_130 , w_131 , \140_b0 );
or ( \142_b1 , \138_b1 , w_133 );
not ( w_133 , w_134 );
and ( \142_b0 , \138_b0 , w_135 );
and ( w_134 ,  , w_135 );
buf ( w_133 , \141_b1 );
not ( w_133 , w_136 );
not (  , w_137 );
and ( w_136 , w_137 , \141_b0 );
or ( \143_b1 , \130_b1 , \142_b1 );
xor ( \143_b0 , \130_b0 , w_138 );
not ( w_138 , w_139 );
and ( w_139 , \142_b1 , \142_b0 );
buf ( \144_b1 , \107_b1 );
not ( \144_b1 , w_140 );
not ( \144_b0 , w_141 );
and ( w_140 , w_141 , \107_b0 );
buf ( \145_b1 , \104_b1 );
not ( \145_b1 , w_142 );
not ( \145_b0 , w_143 );
and ( w_142 , w_143 , \104_b0 );
or ( \146_b1 , \144_b1 , w_144 );
or ( \146_b0 , \144_b0 , \145_b0 );
not ( \145_b0 , w_145 );
and ( w_145 , w_144 , \145_b1 );
or ( \147_b1 , \b[2]_b1 , \b[1]_b1 );
xor ( \147_b0 , \b[2]_b0 , w_146 );
not ( w_146 , w_147 );
and ( w_147 , \b[1]_b1 , \b[1]_b0 );
or ( \148_b1 , \a[4]_b1 , \b[3]_b1 );
xor ( \148_b0 , \a[4]_b0 , w_148 );
not ( w_148 , w_149 );
and ( w_149 , \b[3]_b1 , \b[3]_b0 );
or ( \149_b1 , \147_b1 , w_151 );
not ( w_151 , w_152 );
and ( \149_b0 , \147_b0 , w_153 );
and ( w_152 ,  , w_153 );
buf ( w_151 , \148_b1 );
not ( w_151 , w_154 );
not (  , w_155 );
and ( w_154 , w_155 , \148_b0 );
or ( \150_b1 , \146_b1 , w_157 );
not ( w_157 , w_158 );
and ( \150_b0 , \146_b0 , w_159 );
and ( w_158 ,  , w_159 );
buf ( w_157 , \149_b1 );
not ( w_157 , w_160 );
not (  , w_161 );
and ( w_160 , w_161 , \149_b0 );
or ( \151_b1 , \143_b1 , \150_b1 );
xor ( \151_b0 , \143_b0 , w_162 );
not ( w_162 , w_163 );
and ( w_163 , \150_b1 , \150_b0 );
buf ( \152_b1 , \151_b1 );
not ( \152_b1 , w_164 );
not ( \152_b0 , w_165 );
and ( w_164 , w_165 , \151_b0 );
or ( \153_b1 , \128_b1 , w_166 );
or ( \153_b0 , \128_b0 , \152_b0 );
not ( \152_b0 , w_167 );
and ( w_167 , w_166 , \152_b1 );
or ( \154_b1 , \115_b1 , w_169 );
not ( w_169 , w_170 );
and ( \154_b0 , \115_b0 , w_171 );
and ( w_170 ,  , w_171 );
buf ( w_169 , \125_b1 );
not ( w_169 , w_172 );
not (  , w_173 );
and ( w_172 , w_173 , \125_b0 );
or ( \155_b1 , \153_b1 , w_175 );
not ( w_175 , w_176 );
and ( \155_b0 , \153_b0 , w_177 );
and ( w_176 ,  , w_177 );
buf ( w_175 , \154_b1 );
not ( w_175 , w_178 );
not (  , w_179 );
and ( w_178 , w_179 , \154_b0 );
or ( \156_b1 , \a[0]_b1 , w_180 );
or ( \156_b0 , \a[0]_b0 , \b[6]_b0 );
not ( \b[6]_b0 , w_181 );
and ( w_181 , w_180 , \b[6]_b1 );
or ( \157_b1 , \156_b1 , w_183 );
not ( w_183 , w_184 );
and ( \157_b0 , \156_b0 , w_185 );
and ( w_184 ,  , w_185 );
buf ( w_183 , \b[5]_b1 );
not ( w_183 , w_186 );
not (  , w_187 );
and ( w_186 , w_187 , \b[5]_b0 );
or ( \158_b1 , \a[0]_b1 , w_189 );
not ( w_189 , w_190 );
and ( \158_b0 , \a[0]_b0 , w_191 );
and ( w_190 ,  , w_191 );
buf ( w_189 , \b[6]_b1 );
not ( w_189 , w_192 );
not (  , w_193 );
and ( w_192 , w_193 , \b[6]_b0 );
buf ( \160_b1 , \159_b1 );
not ( \160_b1 , w_194 );
not ( \160_b0 , w_195 );
and ( w_194 , w_195 , \159_b0 );
buf ( \161_b1 , \148_b1 );
not ( \161_b1 , w_196 );
not ( \161_b0 , w_197 );
and ( w_196 , w_197 , \148_b0 );
buf ( \162_b1 , \104_b1 );
not ( \162_b1 , w_198 );
not ( \162_b0 , w_199 );
and ( w_198 , w_199 , \104_b0 );
or ( \163_b1 , \161_b1 , w_200 );
or ( \163_b0 , \161_b0 , \162_b0 );
not ( \162_b0 , w_201 );
and ( w_201 , w_200 , \162_b1 );
or ( \164_b1 , \b[3]_b1 , \a[5]_b1 );
xor ( \164_b0 , \b[3]_b0 , w_202 );
not ( w_202 , w_203 );
and ( w_203 , \a[5]_b1 , \a[5]_b0 );
or ( \165_b1 , \147_b1 , w_205 );
not ( w_205 , w_206 );
and ( \165_b0 , \147_b0 , w_207 );
and ( w_206 ,  , w_207 );
buf ( w_205 , \164_b1 );
not ( w_205 , w_208 );
not (  , w_209 );
and ( w_208 , w_209 , \164_b0 );
or ( \166_b1 , \163_b1 , w_211 );
not ( w_211 , w_212 );
and ( \166_b0 , \163_b0 , w_213 );
and ( w_212 ,  , w_213 );
buf ( w_211 , \165_b1 );
not ( w_211 , w_214 );
not (  , w_215 );
and ( w_214 , w_215 , \165_b0 );
buf ( \167_b1 , \166_b1 );
not ( \167_b1 , w_216 );
not ( \167_b0 , w_217 );
and ( w_216 , w_217 , \166_b0 );
or ( \168_b1 , \160_b1 , w_218 );
or ( \168_b0 , \160_b0 , \167_b0 );
not ( \167_b0 , w_219 );
and ( w_219 , w_218 , \167_b1 );
or ( \169_b1 , \166_b1 , w_220 );
or ( \169_b0 , \166_b0 , \159_b0 );
not ( \159_b0 , w_221 );
and ( w_221 , w_220 , \159_b1 );
or ( \170_b1 , \168_b1 , w_223 );
not ( w_223 , w_224 );
and ( \170_b0 , \168_b0 , w_225 );
and ( w_224 ,  , w_225 );
buf ( w_223 , \169_b1 );
not ( w_223 , w_226 );
not (  , w_227 );
and ( w_226 , w_227 , \169_b0 );
or ( \171_b1 , \130_b1 , \142_b1 );
xor ( \171_b0 , \130_b0 , w_228 );
not ( w_228 , w_229 );
and ( w_229 , \142_b1 , \142_b0 );
or ( \172_b1 , \171_b1 , \150_b1 );
not ( \150_b1 , w_230 );
and ( \172_b0 , \171_b0 , w_231 );
and ( w_230 , w_231 , \150_b0 );
or ( \173_b1 , \130_b1 , \142_b1 );
not ( \142_b1 , w_232 );
and ( \173_b0 , \130_b0 , w_233 );
and ( w_232 , w_233 , \142_b0 );
or ( \174_b1 , \172_b1 , w_234 );
or ( \174_b0 , \172_b0 , \173_b0 );
not ( \173_b0 , w_235 );
and ( w_235 , w_234 , \173_b1 );
or ( \175_b1 , \170_b1 , \174_b1 );
xor ( \175_b0 , \170_b0 , w_236 );
not ( w_236 , w_237 );
and ( w_237 , \174_b1 , \174_b0 );
buf ( \176_b1 , \123_b1 );
not ( \176_b1 , w_238 );
not ( \176_b0 , w_239 );
and ( w_238 , w_239 , \123_b0 );
buf ( \177_b1 , \120_b1 );
not ( \177_b1 , w_240 );
not ( \177_b0 , w_241 );
and ( w_240 , w_241 , \120_b0 );
or ( \178_b1 , \176_b1 , w_242 );
or ( \178_b0 , \176_b0 , \177_b0 );
not ( \177_b0 , w_243 );
and ( w_243 , w_242 , \177_b1 );
or ( \179_b1 , \a[7]_b1 , \b[1]_b1 );
xor ( \179_b0 , \a[7]_b0 , w_244 );
not ( w_244 , w_245 );
and ( w_245 , \b[1]_b1 , \b[1]_b0 );
or ( \180_b1 , \179_b1 , w_247 );
not ( w_247 , w_248 );
and ( \180_b0 , \179_b0 , w_249 );
and ( w_248 ,  , w_249 );
buf ( w_247 , \b[0]_b1 );
not ( w_247 , w_250 );
not (  , w_251 );
and ( w_250 , w_251 , \b[0]_b0 );
or ( \181_b1 , \178_b1 , w_253 );
not ( w_253 , w_254 );
and ( \181_b0 , \178_b0 , w_255 );
and ( w_254 ,  , w_255 );
buf ( w_253 , \180_b1 );
not ( w_253 , w_256 );
not (  , w_257 );
and ( w_256 , w_257 , \180_b0 );
or ( \182_b1 , \a[0]_b1 , \b[7]_b1 );
xor ( \182_b0 , \a[0]_b0 , w_258 );
not ( w_258 , w_259 );
and ( w_259 , \b[7]_b1 , \b[7]_b0 );
buf ( \183_b1 , \182_b1 );
not ( \183_b1 , w_260 );
not ( \183_b0 , w_261 );
and ( w_260 , w_261 , \182_b0 );
or ( \184_b1 , \b[6]_b1 , \b[5]_b1 );
xor ( \184_b0 , \b[6]_b0 , w_262 );
not ( w_262 , w_263 );
and ( w_263 , \b[5]_b1 , \b[5]_b0 );
or ( \185_b1 , \b[7]_b1 , w_264 );
xor ( \185_b0 , \b[7]_b0 , w_266 );
not ( w_266 , w_267 );
and ( w_267 , w_264 , w_265 );
buf ( w_264 , \b[6]_b1 );
not ( w_264 , w_268 );
not ( w_265 , w_269 );
and ( w_268 , w_269 , \b[6]_b0 );
or ( \186_b1 , \184_b1 , w_271 );
not ( w_271 , w_272 );
and ( \186_b0 , \184_b0 , w_273 );
and ( w_272 ,  , w_273 );
buf ( w_271 , \185_b1 );
not ( w_271 , w_274 );
not (  , w_275 );
and ( w_274 , w_275 , \185_b0 );
buf ( \187_b1 , \186_b1 );
not ( \187_b1 , w_276 );
not ( \187_b0 , w_277 );
and ( w_276 , w_277 , \186_b0 );
or ( \188_b1 , \183_b1 , w_278 );
or ( \188_b0 , \183_b0 , \187_b0 );
not ( \187_b0 , w_279 );
and ( w_279 , w_278 , \187_b1 );
or ( \189_b1 , \b[7]_b1 , \a[1]_b1 );
xor ( \189_b0 , \b[7]_b0 , w_280 );
not ( w_280 , w_281 );
and ( w_281 , \a[1]_b1 , \a[1]_b0 );
or ( \190_b1 , \129_b1 , w_283 );
not ( w_283 , w_284 );
and ( \190_b0 , \129_b0 , w_285 );
and ( w_284 ,  , w_285 );
buf ( w_283 , \189_b1 );
not ( w_283 , w_286 );
not (  , w_287 );
and ( w_286 , w_287 , \189_b0 );
or ( \191_b1 , \188_b1 , w_289 );
not ( w_289 , w_290 );
and ( \191_b0 , \188_b0 , w_291 );
and ( w_290 ,  , w_291 );
buf ( w_289 , \190_b1 );
not ( w_289 , w_292 );
not (  , w_293 );
and ( w_292 , w_293 , \190_b0 );
or ( \192_b1 , \181_b1 , \191_b1 );
xor ( \192_b0 , \181_b0 , w_294 );
not ( w_294 , w_295 );
and ( w_295 , \191_b1 , \191_b0 );
buf ( \193_b1 , \140_b1 );
not ( \193_b1 , w_296 );
not ( \193_b0 , w_297 );
and ( w_296 , w_297 , \140_b0 );
buf ( \194_b1 , \133_b1 );
not ( \194_b1 , w_298 );
not ( \194_b0 , w_299 );
and ( w_298 , w_299 , \133_b0 );
or ( \195_b1 , \194_b1 , w_301 );
not ( w_301 , w_302 );
and ( \195_b0 , \194_b0 , w_303 );
and ( w_302 ,  , w_303 );
buf ( w_301 , \135_b1 );
not ( w_301 , w_304 );
not (  , w_305 );
and ( w_304 , w_305 , \135_b0 );
buf ( \196_b1 , \195_b1 );
not ( \196_b1 , w_306 );
not ( \196_b0 , w_307 );
and ( w_306 , w_307 , \195_b0 );
or ( \197_b1 , \193_b1 , w_308 );
or ( \197_b0 , \193_b0 , \196_b0 );
not ( \196_b0 , w_309 );
and ( w_309 , w_308 , \196_b1 );
or ( \198_b1 , \a[3]_b1 , \b[5]_b1 );
xor ( \198_b0 , \a[3]_b0 , w_310 );
not ( w_310 , w_311 );
and ( w_311 , \b[5]_b1 , \b[5]_b0 );
or ( \199_b1 , \139_b1 , w_313 );
not ( w_313 , w_314 );
and ( \199_b0 , \139_b0 , w_315 );
and ( w_314 ,  , w_315 );
buf ( w_313 , \198_b1 );
not ( w_313 , w_316 );
not (  , w_317 );
and ( w_316 , w_317 , \198_b0 );
or ( \200_b1 , \197_b1 , w_319 );
not ( w_319 , w_320 );
and ( \200_b0 , \197_b0 , w_321 );
and ( w_320 ,  , w_321 );
buf ( w_319 , \199_b1 );
not ( w_319 , w_322 );
not (  , w_323 );
and ( w_322 , w_323 , \199_b0 );
or ( \201_b1 , \192_b1 , \200_b1 );
xor ( \201_b0 , \192_b0 , w_324 );
not ( w_324 , w_325 );
and ( w_325 , \200_b1 , \200_b0 );
or ( \202_b1 , \175_b1 , \201_b1 );
xor ( \202_b0 , \175_b0 , w_326 );
not ( w_326 , w_327 );
and ( w_327 , \201_b1 , \201_b0 );
or ( \203_b1 , \155_b1 , \202_b1 );
xor ( \203_b0 , \155_b0 , w_328 );
not ( w_328 , w_329 );
and ( w_329 , \202_b1 , \202_b0 );
buf ( \204_b1 , \109_b1 );
not ( \204_b1 , w_330 );
not ( \204_b0 , w_331 );
and ( w_330 , w_331 , \109_b0 );
or ( \205_b1 , \204_b1 , w_332 );
xor ( \205_b0 , \204_b0 , w_334 );
not ( w_334 , w_335 );
and ( w_335 , w_332 , w_333 );
buf ( w_332 , \113_b1 );
not ( w_332 , w_336 );
not ( w_333 , w_337 );
and ( w_336 , w_337 , \113_b0 );
buf ( \206_b1 , \117_b1 );
not ( \206_b1 , w_338 );
not ( \206_b0 , w_339 );
and ( w_338 , w_339 , \117_b0 );
buf ( \207_b1 , \206_b1 );
not ( \207_b1 , w_340 );
not ( \207_b0 , w_341 );
and ( w_340 , w_341 , \206_b0 );
buf ( \208_b1 , \b[0]_b1 );
not ( \208_b1 , w_342 );
not ( \208_b0 , w_343 );
and ( w_342 , w_343 , \b[0]_b0 );
buf ( \209_b1 , \208_b1 );
not ( \209_b1 , w_344 );
not ( \209_b0 , w_345 );
and ( w_344 , w_345 , \208_b0 );
or ( \210_b1 , \207_b1 , \209_b1 );
not ( \209_b1 , w_346 );
and ( \210_b0 , \207_b0 , w_347 );
and ( w_346 , w_347 , \209_b0 );
buf ( \211_b1 , \b[1]_b1 );
not ( \211_b1 , w_348 );
not ( \211_b0 , w_349 );
and ( w_348 , w_349 , \b[1]_b0 );
or ( \212_b1 , \211_b1 , w_351 );
not ( w_351 , w_352 );
and ( \212_b0 , \211_b0 , w_353 );
and ( w_352 ,  , w_353 );
buf ( w_351 , \b[0]_b1 );
not ( w_351 , w_354 );
not (  , w_355 );
and ( w_354 , w_355 , \b[0]_b0 );
or ( \213_b1 , \a[4]_b1 , \b[1]_b1 );
xor ( \213_b0 , \a[4]_b0 , w_356 );
not ( w_356 , w_357 );
and ( w_357 , \b[1]_b1 , \b[1]_b0 );
or ( \214_b1 , \212_b1 , \213_b1 );
not ( \213_b1 , w_358 );
and ( \214_b0 , \212_b0 , w_359 );
and ( w_358 , w_359 , \213_b0 );
or ( \215_b1 , \210_b1 , w_361 );
not ( w_361 , w_362 );
and ( \215_b0 , \210_b0 , w_363 );
and ( w_362 ,  , w_363 );
buf ( w_361 , \214_b1 );
not ( w_361 , w_364 );
not (  , w_365 );
and ( w_364 , w_365 , \214_b0 );
or ( \216_b1 , \a[0]_b1 , \b[5]_b1 );
xor ( \216_b0 , \a[0]_b0 , w_366 );
not ( w_366 , w_367 );
and ( w_367 , \b[5]_b1 , \b[5]_b0 );
or ( \217_b1 , \b[4]_b1 , w_369 );
not ( w_369 , w_370 );
and ( \217_b0 , \b[4]_b0 , w_371 );
and ( w_370 ,  , w_371 );
buf ( w_369 , \b[3]_b1 );
not ( w_369 , w_372 );
not (  , w_373 );
and ( w_372 , w_373 , \b[3]_b0 );
or ( \219_b1 , \b[4]_b1 , \b[3]_b1 );
not ( \b[3]_b1 , w_374 );
and ( \219_b0 , \b[4]_b0 , w_375 );
and ( w_374 , w_375 , \b[3]_b0 );
or ( \221_b1 , \135_b1 , w_377 );
not ( w_377 , w_378 );
and ( \221_b0 , \135_b0 , w_379 );
and ( w_378 ,  , w_379 );
buf ( w_377 , \131_b1 );
not ( w_377 , w_380 );
not (  , w_381 );
and ( w_380 , w_381 , \131_b0 );
or ( \223_b1 , \215_b1 , \222_b1 );
not ( \222_b1 , w_382 );
and ( \223_b0 , \215_b0 , w_383 );
and ( w_382 , w_383 , \222_b0 );
or ( \224_b1 , \205_b1 , w_384 );
or ( \224_b0 , \205_b0 , \223_b0 );
not ( \223_b0 , w_385 );
and ( w_385 , w_384 , \223_b1 );
or ( \225_b1 , \222_b1 , w_386 );
or ( \225_b0 , \222_b0 , \215_b0 );
not ( \215_b0 , w_387 );
and ( w_387 , w_386 , \215_b1 );
or ( \226_b1 , \224_b1 , w_389 );
not ( w_389 , w_390 );
and ( \226_b0 , \224_b0 , w_391 );
and ( w_390 ,  , w_391 );
buf ( w_389 , \225_b1 );
not ( w_389 , w_392 );
not (  , w_393 );
and ( w_392 , w_393 , \225_b0 );
buf ( \227_b1 , \226_b1 );
not ( \227_b1 , w_394 );
not ( \227_b0 , w_395 );
and ( w_394 , w_395 , \226_b0 );
buf ( \228_b1 , \151_b1 );
not ( \228_b1 , w_396 );
not ( \228_b0 , w_397 );
and ( w_396 , w_397 , \151_b0 );
or ( \229_b1 , \109_b1 , \114_b1 );
not ( \114_b1 , w_398 );
and ( \229_b0 , \109_b0 , w_399 );
and ( w_398 , w_399 , \114_b0 );
buf ( \230_b1 , \229_b1 );
not ( \230_b1 , w_400 );
not ( \230_b0 , w_401 );
and ( w_400 , w_401 , \229_b0 );
buf ( \231_b1 , \126_b1 );
not ( \231_b1 , w_402 );
not ( \231_b0 , w_403 );
and ( w_402 , w_403 , \126_b0 );
or ( \232_b1 , \230_b1 , \231_b1 );
not ( \231_b1 , w_404 );
and ( \232_b0 , \230_b0 , w_405 );
and ( w_404 , w_405 , \231_b0 );
or ( \233_b1 , \115_b1 , \126_b1 );
not ( \126_b1 , w_406 );
and ( \233_b0 , \115_b0 , w_407 );
and ( w_406 , w_407 , \126_b0 );
or ( \234_b1 , \232_b1 , w_409 );
not ( w_409 , w_410 );
and ( \234_b0 , \232_b0 , w_411 );
and ( w_410 ,  , w_411 );
buf ( w_409 , \233_b1 );
not ( w_409 , w_412 );
not (  , w_413 );
and ( w_412 , w_413 , \233_b0 );
buf ( \235_b1 , \234_b1 );
not ( \235_b1 , w_414 );
not ( \235_b0 , w_415 );
and ( w_414 , w_415 , \234_b0 );
or ( \236_b1 , \228_b1 , \235_b1 );
not ( \235_b1 , w_416 );
and ( \236_b0 , \228_b0 , w_417 );
and ( w_416 , w_417 , \235_b0 );
or ( \237_b1 , \151_b1 , \234_b1 );
not ( \234_b1 , w_418 );
and ( \237_b0 , \151_b0 , w_419 );
and ( w_418 , w_419 , \234_b0 );
or ( \238_b1 , \236_b1 , w_421 );
not ( w_421 , w_422 );
and ( \238_b0 , \236_b0 , w_423 );
and ( w_422 ,  , w_423 );
buf ( w_421 , \237_b1 );
not ( w_421 , w_424 );
not (  , w_425 );
and ( w_424 , w_425 , \237_b0 );
or ( \239_b1 , \227_b1 , w_427 );
not ( w_427 , w_428 );
and ( \239_b0 , \227_b0 , w_429 );
and ( w_428 ,  , w_429 );
buf ( w_427 , \238_b1 );
not ( w_427 , w_430 );
not (  , w_431 );
and ( w_430 , w_431 , \238_b0 );
buf ( \240_b1 , \239_b1 );
not ( \240_b1 , w_432 );
not ( \240_b0 , w_433 );
and ( w_432 , w_433 , \239_b0 );
or ( \241_b1 , \139_b1 , w_435 );
not ( w_435 , w_436 );
and ( \241_b0 , \139_b0 , w_437 );
and ( w_436 ,  , w_437 );
buf ( w_435 , \a[0]_b1 );
not ( w_435 , w_438 );
not (  , w_439 );
and ( w_438 , w_439 , \a[0]_b0 );
buf ( \242_b1 , \241_b1 );
not ( \242_b1 , w_440 );
not ( \242_b0 , w_441 );
and ( w_440 , w_441 , \241_b0 );
or ( \243_b1 , \a[3]_b1 , \b[1]_b1 );
xor ( \243_b0 , \a[3]_b0 , w_442 );
not ( w_442 , w_443 );
and ( w_443 , \b[1]_b1 , \b[1]_b0 );
buf ( \244_b1 , \243_b1 );
not ( \244_b1 , w_444 );
not ( \244_b0 , w_445 );
and ( w_444 , w_445 , \243_b0 );
buf ( \245_b1 , \212_b1 );
not ( \245_b1 , w_446 );
not ( \245_b0 , w_447 );
and ( w_446 , w_447 , \212_b0 );
or ( \246_b1 , \244_b1 , w_448 );
or ( \246_b0 , \244_b0 , \245_b0 );
not ( \245_b0 , w_449 );
and ( w_449 , w_448 , \245_b1 );
or ( \247_b1 , \213_b1 , w_451 );
not ( w_451 , w_452 );
and ( \247_b0 , \213_b0 , w_453 );
and ( w_452 ,  , w_453 );
buf ( w_451 , \b[0]_b1 );
not ( w_451 , w_454 );
not (  , w_455 );
and ( w_454 , w_455 , \b[0]_b0 );
or ( \248_b1 , \246_b1 , w_457 );
not ( w_457 , w_458 );
and ( \248_b0 , \246_b0 , w_459 );
and ( w_458 ,  , w_459 );
buf ( w_457 , \247_b1 );
not ( w_457 , w_460 );
not (  , w_461 );
and ( w_460 , w_461 , \247_b0 );
buf ( \249_b1 , \248_b1 );
not ( \249_b1 , w_462 );
not ( \249_b0 , w_463 );
and ( w_462 , w_463 , \248_b0 );
buf ( \250_b1 , \249_b1 );
not ( \250_b1 , w_464 );
not ( \250_b0 , w_465 );
and ( w_464 , w_465 , \249_b0 );
or ( \251_b1 , \242_b1 , w_466 );
or ( \251_b0 , \242_b0 , \250_b0 );
not ( \250_b0 , w_467 );
and ( w_467 , w_466 , \250_b1 );
or ( \252_b1 , \a[1]_b1 , \b[3]_b1 );
xor ( \252_b0 , \a[1]_b0 , w_468 );
not ( w_468 , w_469 );
and ( w_469 , \b[3]_b1 , \b[3]_b0 );
buf ( \253_b1 , \252_b1 );
not ( \253_b1 , w_470 );
not ( \253_b0 , w_471 );
and ( w_470 , w_471 , \252_b0 );
buf ( \254_b1 , \104_b1 );
not ( \254_b1 , w_472 );
not ( \254_b0 , w_473 );
and ( w_472 , w_473 , \104_b0 );
or ( \255_b1 , \253_b1 , w_474 );
or ( \255_b0 , \253_b0 , \254_b0 );
not ( \254_b0 , w_475 );
and ( w_475 , w_474 , \254_b1 );
or ( \256_b1 , \147_b1 , w_477 );
not ( w_477 , w_478 );
and ( \256_b0 , \147_b0 , w_479 );
and ( w_478 ,  , w_479 );
buf ( w_477 , \100_b1 );
not ( w_477 , w_480 );
not (  , w_481 );
and ( w_480 , w_481 , \100_b0 );
or ( \257_b1 , \255_b1 , w_483 );
not ( w_483 , w_484 );
and ( \257_b0 , \255_b0 , w_485 );
and ( w_484 ,  , w_485 );
buf ( w_483 , \256_b1 );
not ( w_483 , w_486 );
not (  , w_487 );
and ( w_486 , w_487 , \256_b0 );
or ( \258_b1 , \251_b1 , w_489 );
not ( w_489 , w_490 );
and ( \258_b0 , \251_b0 , w_491 );
and ( w_490 ,  , w_491 );
buf ( w_489 , \257_b1 );
not ( w_489 , w_492 );
not (  , w_493 );
and ( w_492 , w_493 , \257_b0 );
buf ( \259_b1 , \241_b1 );
not ( \259_b1 , w_494 );
not ( \259_b0 , w_495 );
and ( w_494 , w_495 , \241_b0 );
or ( \260_b1 , \259_b1 , w_497 );
not ( w_497 , w_498 );
and ( \260_b0 , \259_b0 , w_499 );
and ( w_498 ,  , w_499 );
buf ( w_497 , \248_b1 );
not ( w_497 , w_500 );
not (  , w_501 );
and ( w_500 , w_501 , \248_b0 );
or ( \261_b1 , \258_b1 , w_503 );
not ( w_503 , w_504 );
and ( \261_b0 , \258_b0 , w_505 );
and ( w_504 ,  , w_505 );
buf ( w_503 , \260_b1 );
not ( w_503 , w_506 );
not (  , w_507 );
and ( w_506 , w_507 , \260_b0 );
buf ( \262_b1 , \261_b1 );
not ( \262_b1 , w_508 );
not ( \262_b0 , w_509 );
and ( w_508 , w_509 , \261_b0 );
buf ( \263_b1 , \262_b1 );
not ( \263_b1 , w_510 );
not ( \263_b0 , w_511 );
and ( w_510 , w_511 , \262_b0 );
or ( \264_b1 , \113_b1 , \204_b1 );
xor ( \264_b0 , \113_b0 , w_512 );
not ( w_512 , w_513 );
and ( w_513 , \204_b1 , \204_b0 );
or ( \265_b1 , \215_b1 , \222_b1 );
xor ( \265_b0 , \215_b0 , w_514 );
not ( w_514 , w_515 );
and ( w_515 , \222_b1 , \222_b0 );
or ( \266_b1 , \264_b1 , w_516 );
xor ( \266_b0 , \264_b0 , w_518 );
not ( w_518 , w_519 );
and ( w_519 , w_516 , w_517 );
buf ( w_516 , \265_b1 );
not ( w_516 , w_520 );
not ( w_517 , w_521 );
and ( w_520 , w_521 , \265_b0 );
buf ( \267_b1 , \266_b1 );
not ( \267_b1 , w_522 );
not ( \267_b0 , w_523 );
and ( w_522 , w_523 , \266_b0 );
or ( \268_b1 , \263_b1 , w_524 );
or ( \268_b0 , \263_b0 , \267_b0 );
not ( \267_b0 , w_525 );
and ( w_525 , w_524 , \267_b1 );
or ( \269_b1 , \248_b1 , \241_b1 );
not ( \241_b1 , w_526 );
and ( \269_b0 , \248_b0 , w_527 );
and ( w_526 , w_527 , \241_b0 );
buf ( \270_b1 , \248_b1 );
not ( \270_b1 , w_528 );
not ( \270_b0 , w_529 );
and ( w_528 , w_529 , \248_b0 );
or ( \271_b1 , \139_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_530 );
and ( \271_b0 , \139_b0 , w_531 );
and ( w_530 , w_531 , \a[0]_b0 );
or ( \272_b1 , \270_b1 , \271_b1 );
not ( \271_b1 , w_532 );
and ( \272_b0 , \270_b0 , w_533 );
and ( w_532 , w_533 , \271_b0 );
or ( \273_b1 , \269_b1 , w_535 );
not ( w_535 , w_536 );
and ( \273_b0 , \269_b0 , w_537 );
and ( w_536 ,  , w_537 );
buf ( w_535 , \272_b1 );
not ( w_535 , w_538 );
not (  , w_539 );
and ( w_538 , w_539 , \272_b0 );
or ( \274_b1 , \273_b1 , \257_b1 );
not ( \257_b1 , w_540 );
and ( \274_b0 , \273_b0 , w_541 );
and ( w_540 , w_541 , \257_b0 );
buf ( \275_b1 , \273_b1 );
not ( \275_b1 , w_542 );
not ( \275_b0 , w_543 );
and ( w_542 , w_543 , \273_b0 );
buf ( \276_b1 , \257_b1 );
not ( \276_b1 , w_544 );
not ( \276_b0 , w_545 );
and ( w_544 , w_545 , \257_b0 );
or ( \277_b1 , \275_b1 , \276_b1 );
not ( \276_b1 , w_546 );
and ( \277_b0 , \275_b0 , w_547 );
and ( w_546 , w_547 , \276_b0 );
or ( \278_b1 , \274_b1 , w_549 );
not ( w_549 , w_550 );
and ( \278_b0 , \274_b0 , w_551 );
and ( w_550 ,  , w_551 );
buf ( w_549 , \277_b1 );
not ( w_549 , w_552 );
not (  , w_553 );
and ( w_552 , w_553 , \277_b0 );
or ( \279_b1 , \a[0]_b1 , w_555 );
not ( w_555 , w_556 );
and ( \279_b0 , \a[0]_b0 , w_557 );
and ( w_556 ,  , w_557 );
buf ( w_555 , \b[2]_b1 );
not ( w_555 , w_558 );
not (  , w_559 );
and ( w_558 , w_559 , \b[2]_b0 );
or ( \280_b1 , \a[0]_b1 , w_560 );
or ( \280_b0 , \a[0]_b0 , \b[2]_b0 );
not ( \b[2]_b0 , w_561 );
and ( w_561 , w_560 , \b[2]_b1 );
or ( \281_b1 , \280_b1 , w_563 );
not ( w_563 , w_564 );
and ( \281_b0 , \280_b0 , w_565 );
and ( w_564 ,  , w_565 );
buf ( w_563 , \b[1]_b1 );
not ( w_563 , w_566 );
not (  , w_567 );
and ( w_566 , w_567 , \b[1]_b0 );
buf ( \283_b1 , \282_b1 );
not ( \283_b1 , w_568 );
not ( \283_b0 , w_569 );
and ( w_568 , w_569 , \282_b0 );
or ( \284_b1 , \a[2]_b1 , \b[1]_b1 );
xor ( \284_b0 , \a[2]_b0 , w_570 );
not ( w_570 , w_571 );
and ( w_571 , \b[1]_b1 , \b[1]_b0 );
buf ( \285_b1 , \284_b1 );
not ( \285_b1 , w_572 );
not ( \285_b0 , w_573 );
and ( w_572 , w_573 , \284_b0 );
buf ( \286_b1 , \212_b1 );
not ( \286_b1 , w_574 );
not ( \286_b0 , w_575 );
and ( w_574 , w_575 , \212_b0 );
or ( \287_b1 , \285_b1 , w_576 );
or ( \287_b0 , \285_b0 , \286_b0 );
not ( \286_b0 , w_577 );
and ( w_577 , w_576 , \286_b1 );
or ( \288_b1 , \243_b1 , w_579 );
not ( w_579 , w_580 );
and ( \288_b0 , \243_b0 , w_581 );
and ( w_580 ,  , w_581 );
buf ( w_579 , \b[0]_b1 );
not ( w_579 , w_582 );
not (  , w_583 );
and ( w_582 , w_583 , \b[0]_b0 );
or ( \289_b1 , \287_b1 , w_585 );
not ( w_585 , w_586 );
and ( \289_b0 , \287_b0 , w_587 );
and ( w_586 ,  , w_587 );
buf ( w_585 , \288_b1 );
not ( w_585 , w_588 );
not (  , w_589 );
and ( w_588 , w_589 , \288_b0 );
or ( \290_b1 , \283_b1 , w_591 );
not ( w_591 , w_592 );
and ( \290_b0 , \283_b0 , w_593 );
and ( w_592 ,  , w_593 );
buf ( w_591 , \289_b1 );
not ( w_591 , w_594 );
not (  , w_595 );
and ( w_594 , w_595 , \289_b0 );
or ( \291_b1 , \278_b1 , w_597 );
not ( w_597 , w_598 );
and ( \291_b0 , \278_b0 , w_599 );
and ( w_598 ,  , w_599 );
buf ( w_597 , \290_b1 );
not ( w_597 , w_600 );
not (  , w_601 );
and ( w_600 , w_601 , \290_b0 );
buf ( \292_b1 , \291_b1 );
not ( \292_b1 , w_602 );
not ( \292_b0 , w_603 );
and ( w_602 , w_603 , \291_b0 );
or ( \293_b1 , \b[3]_b1 , \a[0]_b1 );
xor ( \293_b0 , \b[3]_b0 , w_604 );
not ( w_604 , w_605 );
and ( w_605 , \a[0]_b1 , \a[0]_b0 );
buf ( \294_b1 , \293_b1 );
not ( \294_b1 , w_606 );
not ( \294_b0 , w_607 );
and ( w_606 , w_607 , \293_b0 );
or ( \295_b1 , \102_b1 , w_609 );
not ( w_609 , w_610 );
and ( \295_b0 , \102_b0 , w_611 );
and ( w_610 ,  , w_611 );
buf ( w_609 , \103_b1 );
not ( w_609 , w_612 );
not (  , w_613 );
and ( w_612 , w_613 , \103_b0 );
buf ( \296_b1 , \295_b1 );
not ( \296_b1 , w_614 );
not ( \296_b0 , w_615 );
and ( w_614 , w_615 , \295_b0 );
or ( \297_b1 , \294_b1 , w_616 );
or ( \297_b0 , \294_b0 , \296_b0 );
not ( \296_b0 , w_617 );
and ( w_617 , w_616 , \296_b1 );
or ( \298_b1 , \147_b1 , w_619 );
not ( w_619 , w_620 );
and ( \298_b0 , \147_b0 , w_621 );
and ( w_620 ,  , w_621 );
buf ( w_619 , \252_b1 );
not ( w_619 , w_622 );
not (  , w_623 );
and ( w_622 , w_623 , \252_b0 );
or ( \299_b1 , \297_b1 , w_625 );
not ( w_625 , w_626 );
and ( \299_b0 , \297_b0 , w_627 );
and ( w_626 ,  , w_627 );
buf ( w_625 , \298_b1 );
not ( w_625 , w_628 );
not (  , w_629 );
and ( w_628 , w_629 , \298_b0 );
buf ( \300_b1 , \299_b1 );
not ( \300_b1 , w_630 );
not ( \300_b0 , w_631 );
and ( w_630 , w_631 , \299_b0 );
or ( \301_b1 , \289_b1 , \282_b1 );
xor ( \301_b0 , \289_b0 , w_632 );
not ( w_632 , w_633 );
and ( w_633 , \282_b1 , \282_b0 );
or ( \302_b1 , \300_b1 , w_635 );
not ( w_635 , w_636 );
and ( \302_b0 , \300_b0 , w_637 );
and ( w_636 ,  , w_637 );
buf ( w_635 , \301_b1 );
not ( w_635 , w_638 );
not (  , w_639 );
and ( w_638 , w_639 , \301_b0 );
buf ( \303_b1 , \302_b1 );
not ( \303_b1 , w_640 );
not ( \303_b0 , w_641 );
and ( w_640 , w_641 , \302_b0 );
or ( \304_b1 , \147_b1 , w_643 );
not ( w_643 , w_644 );
and ( \304_b0 , \147_b0 , w_645 );
and ( w_644 ,  , w_645 );
buf ( w_643 , \a[0]_b1 );
not ( w_643 , w_646 );
not (  , w_647 );
and ( w_646 , w_647 , \a[0]_b0 );
buf ( \305_b1 , \304_b1 );
not ( \305_b1 , w_648 );
not ( \305_b0 , w_649 );
and ( w_648 , w_649 , \304_b0 );
or ( \306_b1 , \b[1]_b1 , \a[1]_b1 );
xor ( \306_b0 , \b[1]_b0 , w_650 );
not ( w_650 , w_651 );
and ( w_651 , \a[1]_b1 , \a[1]_b0 );
buf ( \307_b1 , \306_b1 );
not ( \307_b1 , w_652 );
not ( \307_b0 , w_653 );
and ( w_652 , w_653 , \306_b0 );
buf ( \308_b1 , \120_b1 );
not ( \308_b1 , w_654 );
not ( \308_b0 , w_655 );
and ( w_654 , w_655 , \120_b0 );
or ( \309_b1 , \307_b1 , w_656 );
or ( \309_b0 , \307_b0 , \308_b0 );
not ( \308_b0 , w_657 );
and ( w_657 , w_656 , \308_b1 );
or ( \310_b1 , \284_b1 , w_659 );
not ( w_659 , w_660 );
and ( \310_b0 , \284_b0 , w_661 );
and ( w_660 ,  , w_661 );
buf ( w_659 , \b[0]_b1 );
not ( w_659 , w_662 );
not (  , w_663 );
and ( w_662 , w_663 , \b[0]_b0 );
or ( \311_b1 , \309_b1 , w_665 );
not ( w_665 , w_666 );
and ( \311_b0 , \309_b0 , w_667 );
and ( w_666 ,  , w_667 );
buf ( w_665 , \310_b1 );
not ( w_665 , w_668 );
not (  , w_669 );
and ( w_668 , w_669 , \310_b0 );
or ( \312_b1 , \305_b1 , w_671 );
not ( w_671 , w_672 );
and ( \312_b0 , \305_b0 , w_673 );
and ( w_672 ,  , w_673 );
buf ( w_671 , \311_b1 );
not ( w_671 , w_674 );
not (  , w_675 );
and ( w_674 , w_675 , \311_b0 );
buf ( \313_b1 , \b[0]_b1 );
not ( \313_b1 , w_676 );
not ( \313_b0 , w_677 );
and ( w_676 , w_677 , \b[0]_b0 );
buf ( \314_b1 , \306_b1 );
not ( \314_b1 , w_678 );
not ( \314_b0 , w_679 );
and ( w_678 , w_679 , \306_b0 );
buf ( \315_b1 , \314_b1 );
not ( \315_b1 , w_680 );
not ( \315_b0 , w_681 );
and ( w_680 , w_681 , \314_b0 );
or ( \316_b1 , \313_b1 , w_682 );
or ( \316_b0 , \313_b0 , \315_b0 );
not ( \315_b0 , w_683 );
and ( w_683 , w_682 , \315_b1 );
or ( \317_b1 , \a[0]_b1 , w_685 );
not ( w_685 , w_686 );
and ( \317_b0 , \a[0]_b0 , w_687 );
and ( w_686 ,  , w_687 );
buf ( w_685 , \b[0]_b1 );
not ( w_685 , w_688 );
not (  , w_689 );
and ( w_688 , w_689 , \b[0]_b0 );
or ( \318_b1 , \317_b1 , w_691 );
not ( w_691 , w_692 );
and ( \318_b0 , \317_b0 , w_693 );
and ( w_692 ,  , w_693 );
buf ( w_691 , \b[1]_b1 );
not ( w_691 , w_694 );
not (  , w_695 );
and ( w_694 , w_695 , \b[1]_b0 );
or ( \319_b1 , \318_b1 , w_697 );
not ( w_697 , w_698 );
and ( \319_b0 , \318_b0 , w_699 );
and ( w_698 ,  , w_699 );
buf ( w_697 , \a[0]_b1 );
not ( w_697 , w_700 );
not (  , w_701 );
and ( w_700 , w_701 , \a[0]_b0 );
or ( \320_b1 , \316_b1 , w_703 );
not ( w_703 , w_704 );
and ( \320_b0 , \316_b0 , w_705 );
and ( w_704 ,  , w_705 );
buf ( w_703 , \319_b1 );
not ( w_703 , w_706 );
not (  , w_707 );
and ( w_706 , w_707 , \319_b0 );
or ( \321_b1 , \312_b1 , w_708 );
or ( \321_b0 , \312_b0 , \320_b0 );
not ( \320_b0 , w_709 );
and ( w_709 , w_708 , \320_b1 );
buf ( \322_b1 , \304_b1 );
not ( \322_b1 , w_710 );
not ( \322_b0 , w_711 );
and ( w_710 , w_711 , \304_b0 );
or ( \323_b1 , \322_b1 , w_713 );
not ( w_713 , w_714 );
and ( \323_b0 , \322_b0 , w_715 );
and ( w_714 ,  , w_715 );
buf ( w_713 , \311_b1 );
not ( w_713 , w_716 );
not (  , w_717 );
and ( w_716 , w_717 , \311_b0 );
or ( \324_b1 , \321_b1 , w_719 );
not ( w_719 , w_720 );
and ( \324_b0 , \321_b0 , w_721 );
and ( w_720 ,  , w_721 );
buf ( w_719 , \323_b1 );
not ( w_719 , w_722 );
not (  , w_723 );
and ( w_722 , w_723 , \323_b0 );
buf ( \325_b1 , \324_b1 );
not ( \325_b1 , w_724 );
not ( \325_b0 , w_725 );
and ( w_724 , w_725 , \324_b0 );
or ( \326_b1 , \303_b1 , w_726 );
or ( \326_b0 , \303_b0 , \325_b0 );
not ( \325_b0 , w_727 );
and ( w_727 , w_726 , \325_b1 );
buf ( \327_b1 , \301_b1 );
not ( \327_b1 , w_728 );
not ( \327_b0 , w_729 );
and ( w_728 , w_729 , \301_b0 );
or ( \328_b1 , \327_b1 , w_731 );
not ( w_731 , w_732 );
and ( \328_b0 , \327_b0 , w_733 );
and ( w_732 ,  , w_733 );
buf ( w_731 , \299_b1 );
not ( w_731 , w_734 );
not (  , w_735 );
and ( w_734 , w_735 , \299_b0 );
or ( \329_b1 , \326_b1 , w_737 );
not ( w_737 , w_738 );
and ( \329_b0 , \326_b0 , w_739 );
and ( w_738 ,  , w_739 );
buf ( w_737 , \328_b1 );
not ( w_737 , w_740 );
not (  , w_741 );
and ( w_740 , w_741 , \328_b0 );
buf ( \330_b1 , \329_b1 );
not ( \330_b1 , w_742 );
not ( \330_b0 , w_743 );
and ( w_742 , w_743 , \329_b0 );
or ( \331_b1 , \292_b1 , w_744 );
or ( \331_b0 , \292_b0 , \330_b0 );
not ( \330_b0 , w_745 );
and ( w_745 , w_744 , \330_b1 );
buf ( \332_b1 , \278_b1 );
not ( \332_b1 , w_746 );
not ( \332_b0 , w_747 );
and ( w_746 , w_747 , \278_b0 );
buf ( \333_b1 , \290_b1 );
not ( \333_b1 , w_748 );
not ( \333_b0 , w_749 );
and ( w_748 , w_749 , \290_b0 );
or ( \334_b1 , \332_b1 , w_751 );
not ( w_751 , w_752 );
and ( \334_b0 , \332_b0 , w_753 );
and ( w_752 ,  , w_753 );
buf ( w_751 , \333_b1 );
not ( w_751 , w_754 );
not (  , w_755 );
and ( w_754 , w_755 , \333_b0 );
or ( \335_b1 , \331_b1 , w_757 );
not ( w_757 , w_758 );
and ( \335_b0 , \331_b0 , w_759 );
and ( w_758 ,  , w_759 );
buf ( w_757 , \334_b1 );
not ( w_757 , w_760 );
not (  , w_761 );
and ( w_760 , w_761 , \334_b0 );
or ( \336_b1 , \268_b1 , w_763 );
not ( w_763 , w_764 );
and ( \336_b0 , \268_b0 , w_765 );
and ( w_764 ,  , w_765 );
buf ( w_763 , \335_b1 );
not ( w_763 , w_766 );
not (  , w_767 );
and ( w_766 , w_767 , \335_b0 );
buf ( \337_b1 , \266_b1 );
not ( \337_b1 , w_768 );
not ( \337_b0 , w_769 );
and ( w_768 , w_769 , \266_b0 );
or ( \338_b1 , \337_b1 , w_771 );
not ( w_771 , w_772 );
and ( \338_b0 , \337_b0 , w_773 );
and ( w_772 ,  , w_773 );
buf ( w_771 , \261_b1 );
not ( w_771 , w_774 );
not (  , w_775 );
and ( w_774 , w_775 , \261_b0 );
or ( \339_b1 , \336_b1 , w_777 );
not ( w_777 , w_778 );
and ( \339_b0 , \336_b0 , w_779 );
and ( w_778 ,  , w_779 );
buf ( w_777 , \338_b1 );
not ( w_777 , w_780 );
not (  , w_781 );
and ( w_780 , w_781 , \338_b0 );
buf ( \340_b1 , \339_b1 );
not ( \340_b1 , w_782 );
not ( \340_b0 , w_783 );
and ( w_782 , w_783 , \339_b0 );
or ( \341_b1 , \240_b1 , w_784 );
or ( \341_b0 , \240_b0 , \340_b0 );
not ( \340_b0 , w_785 );
and ( w_785 , w_784 , \340_b1 );
buf ( \342_b1 , \238_b1 );
not ( \342_b1 , w_786 );
not ( \342_b0 , w_787 );
and ( w_786 , w_787 , \238_b0 );
or ( \343_b1 , \342_b1 , w_789 );
not ( w_789 , w_790 );
and ( \343_b0 , \342_b0 , w_791 );
and ( w_790 ,  , w_791 );
buf ( w_789 , \226_b1 );
not ( w_789 , w_792 );
not (  , w_793 );
and ( w_792 , w_793 , \226_b0 );
or ( \344_b1 , \341_b1 , w_795 );
not ( w_795 , w_796 );
and ( \344_b0 , \341_b0 , w_797 );
and ( w_796 ,  , w_797 );
buf ( w_795 , \343_b1 );
not ( w_795 , w_798 );
not (  , w_799 );
and ( w_798 , w_799 , \343_b0 );
or ( \345_b1 , \203_b1 , \344_b1 );
not ( \344_b1 , w_800 );
and ( \345_b0 , \203_b0 , w_801 );
and ( w_800 , w_801 , \344_b0 );
or ( \346_b1 , \155_b1 , \202_b1 );
not ( \202_b1 , w_802 );
and ( \346_b0 , \155_b0 , w_803 );
and ( w_802 , w_803 , \202_b0 );
or ( \347_b1 , \345_b1 , w_804 );
or ( \347_b0 , \345_b0 , \346_b0 );
not ( \346_b0 , w_805 );
and ( w_805 , w_804 , \346_b1 );
buf ( \348_b1 , \120_b1 );
not ( \348_b1 , w_806 );
not ( \348_b0 , w_807 );
and ( w_806 , w_807 , \120_b0 );
or ( \349_b1 , \a[8]_b1 , \b[1]_b1 );
xor ( \349_b0 , \a[8]_b0 , w_808 );
not ( w_808 , w_809 );
and ( w_809 , \b[1]_b1 , \b[1]_b0 );
buf ( \350_b1 , \349_b1 );
not ( \350_b1 , w_810 );
not ( \350_b0 , w_811 );
and ( w_810 , w_811 , \349_b0 );
or ( \351_b1 , \348_b1 , w_812 );
or ( \351_b0 , \348_b0 , \350_b0 );
not ( \350_b0 , w_813 );
and ( w_813 , w_812 , \350_b1 );
or ( \352_b1 , \a[9]_b1 , \b[1]_b1 );
xor ( \352_b0 , \a[9]_b0 , w_814 );
not ( w_814 , w_815 );
and ( w_815 , \b[1]_b1 , \b[1]_b0 );
or ( \353_b1 , \352_b1 , w_817 );
not ( w_817 , w_818 );
and ( \353_b0 , \352_b0 , w_819 );
and ( w_818 ,  , w_819 );
buf ( w_817 , \b[0]_b1 );
not ( w_817 , w_820 );
not (  , w_821 );
and ( w_820 , w_821 , \b[0]_b0 );
or ( \354_b1 , \351_b1 , w_823 );
not ( w_823 , w_824 );
and ( \354_b0 , \351_b0 , w_825 );
and ( w_824 ,  , w_825 );
buf ( w_823 , \353_b1 );
not ( w_823 , w_826 );
not (  , w_827 );
and ( w_826 , w_827 , \353_b0 );
or ( \355_b1 , \b[7]_b1 , \a[2]_b1 );
xor ( \355_b0 , \b[7]_b0 , w_828 );
not ( w_828 , w_829 );
and ( w_829 , \a[2]_b1 , \a[2]_b0 );
buf ( \356_b1 , \355_b1 );
not ( \356_b1 , w_830 );
not ( \356_b0 , w_831 );
and ( w_830 , w_831 , \355_b0 );
buf ( \357_b1 , \186_b1 );
not ( \357_b1 , w_832 );
not ( \357_b0 , w_833 );
and ( w_832 , w_833 , \186_b0 );
or ( \358_b1 , \356_b1 , w_834 );
or ( \358_b0 , \356_b0 , \357_b0 );
not ( \357_b0 , w_835 );
and ( w_835 , w_834 , \357_b1 );
or ( \359_b1 , \a[3]_b1 , \b[7]_b1 );
xor ( \359_b0 , \a[3]_b0 , w_836 );
not ( w_836 , w_837 );
and ( w_837 , \b[7]_b1 , \b[7]_b0 );
or ( \360_b1 , \359_b1 , w_839 );
not ( w_839 , w_840 );
and ( \360_b0 , \359_b0 , w_841 );
and ( w_840 ,  , w_841 );
buf ( w_839 , \129_b1 );
not ( w_839 , w_842 );
not (  , w_843 );
and ( w_842 , w_843 , \129_b0 );
or ( \361_b1 , \358_b1 , w_845 );
not ( w_845 , w_846 );
and ( \361_b0 , \358_b0 , w_847 );
and ( w_846 ,  , w_847 );
buf ( w_845 , \360_b1 );
not ( w_845 , w_848 );
not (  , w_849 );
and ( w_848 , w_849 , \360_b0 );
or ( \362_b1 , \354_b1 , \361_b1 );
xor ( \362_b0 , \354_b0 , w_850 );
not ( w_850 , w_851 );
and ( w_851 , \361_b1 , \361_b0 );
or ( \363_b1 , \a[6]_b1 , \b[3]_b1 );
xor ( \363_b0 , \a[6]_b0 , w_852 );
not ( w_852 , w_853 );
and ( w_853 , \b[3]_b1 , \b[3]_b0 );
buf ( \364_b1 , \363_b1 );
not ( \364_b1 , w_854 );
not ( \364_b0 , w_855 );
and ( w_854 , w_855 , \363_b0 );
buf ( \365_b1 , \295_b1 );
not ( \365_b1 , w_856 );
not ( \365_b0 , w_857 );
and ( w_856 , w_857 , \295_b0 );
or ( \366_b1 , \364_b1 , w_858 );
or ( \366_b0 , \364_b0 , \365_b0 );
not ( \365_b0 , w_859 );
and ( w_859 , w_858 , \365_b1 );
or ( \367_b1 , \a[7]_b1 , \b[3]_b1 );
xor ( \367_b0 , \a[7]_b0 , w_860 );
not ( w_860 , w_861 );
and ( w_861 , \b[3]_b1 , \b[3]_b0 );
or ( \368_b1 , \147_b1 , w_863 );
not ( w_863 , w_864 );
and ( \368_b0 , \147_b0 , w_865 );
and ( w_864 ,  , w_865 );
buf ( w_863 , \367_b1 );
not ( w_863 , w_866 );
not (  , w_867 );
and ( w_866 , w_867 , \367_b0 );
or ( \369_b1 , \366_b1 , w_869 );
not ( w_869 , w_870 );
and ( \369_b0 , \366_b0 , w_871 );
and ( w_870 ,  , w_871 );
buf ( w_869 , \368_b1 );
not ( w_869 , w_872 );
not (  , w_873 );
and ( w_872 , w_873 , \368_b0 );
or ( \370_b1 , \362_b1 , \369_b1 );
xor ( \370_b0 , \362_b0 , w_874 );
not ( w_874 , w_875 );
and ( w_875 , \369_b1 , \369_b0 );
buf ( \371_b1 , \370_b1 );
not ( \371_b1 , w_876 );
not ( \371_b0 , w_877 );
and ( w_876 , w_877 , \370_b0 );
buf ( \372_b1 , \371_b1 );
not ( \372_b1 , w_878 );
not ( \372_b0 , w_879 );
and ( w_878 , w_879 , \371_b0 );
buf ( \373_b1 , \189_b1 );
not ( \373_b1 , w_880 );
not ( \373_b0 , w_881 );
and ( w_880 , w_881 , \189_b0 );
or ( \374_b1 , \185_b1 , w_883 );
not ( w_883 , w_884 );
and ( \374_b0 , \185_b0 , w_885 );
and ( w_884 ,  , w_885 );
buf ( w_883 , \184_b1 );
not ( w_883 , w_886 );
not (  , w_887 );
and ( w_886 , w_887 , \184_b0 );
buf ( \375_b1 , \374_b1 );
not ( \375_b1 , w_888 );
not ( \375_b0 , w_889 );
and ( w_888 , w_889 , \374_b0 );
or ( \376_b1 , \373_b1 , w_890 );
or ( \376_b0 , \373_b0 , \375_b0 );
not ( \375_b0 , w_891 );
and ( w_891 , w_890 , \375_b1 );
or ( \377_b1 , \129_b1 , w_893 );
not ( w_893 , w_894 );
and ( \377_b0 , \129_b0 , w_895 );
and ( w_894 ,  , w_895 );
buf ( w_893 , \355_b1 );
not ( w_893 , w_896 );
not (  , w_897 );
and ( w_896 , w_897 , \355_b0 );
or ( \378_b1 , \376_b1 , w_899 );
not ( w_899 , w_900 );
and ( \378_b0 , \376_b0 , w_901 );
and ( w_900 ,  , w_901 );
buf ( w_899 , \377_b1 );
not ( w_899 , w_902 );
not (  , w_903 );
and ( w_902 , w_903 , \377_b0 );
buf ( \379_b1 , \198_b1 );
not ( \379_b1 , w_904 );
not ( \379_b0 , w_905 );
and ( w_904 , w_905 , \198_b0 );
buf ( \380_b1 , \195_b1 );
not ( \380_b1 , w_906 );
not ( \380_b0 , w_907 );
and ( w_906 , w_907 , \195_b0 );
or ( \381_b1 , \379_b1 , w_908 );
or ( \381_b0 , \379_b0 , \380_b0 );
not ( \380_b0 , w_909 );
and ( w_909 , w_908 , \380_b1 );
or ( \382_b1 , \a[4]_b1 , \b[5]_b1 );
xor ( \382_b0 , \a[4]_b0 , w_910 );
not ( w_910 , w_911 );
and ( w_911 , \b[5]_b1 , \b[5]_b0 );
or ( \383_b1 , \139_b1 , w_913 );
not ( w_913 , w_914 );
and ( \383_b0 , \139_b0 , w_915 );
and ( w_914 ,  , w_915 );
buf ( w_913 , \382_b1 );
not ( w_913 , w_916 );
not (  , w_917 );
and ( w_916 , w_917 , \382_b0 );
or ( \384_b1 , \381_b1 , w_919 );
not ( w_919 , w_920 );
and ( \384_b0 , \381_b0 , w_921 );
and ( w_920 ,  , w_921 );
buf ( w_919 , \383_b1 );
not ( w_919 , w_922 );
not (  , w_923 );
and ( w_922 , w_923 , \383_b0 );
or ( \385_b1 , \378_b1 , \384_b1 );
xor ( \385_b0 , \378_b0 , w_924 );
not ( w_924 , w_925 );
and ( w_925 , \384_b1 , \384_b0 );
buf ( \386_b1 , \166_b1 );
not ( \386_b1 , w_926 );
not ( \386_b0 , w_927 );
and ( w_926 , w_927 , \166_b0 );
or ( \387_b1 , \386_b1 , w_929 );
not ( w_929 , w_930 );
and ( \387_b0 , \386_b0 , w_931 );
and ( w_930 ,  , w_931 );
buf ( w_929 , \159_b1 );
not ( w_929 , w_932 );
not (  , w_933 );
and ( w_932 , w_933 , \159_b0 );
or ( \388_b1 , \385_b1 , \387_b1 );
not ( \387_b1 , w_934 );
and ( \388_b0 , \385_b0 , w_935 );
and ( w_934 , w_935 , \387_b0 );
or ( \389_b1 , \378_b1 , \384_b1 );
not ( \384_b1 , w_936 );
and ( \389_b0 , \378_b0 , w_937 );
and ( w_936 , w_937 , \384_b0 );
or ( \390_b1 , \388_b1 , w_938 );
or ( \390_b0 , \388_b0 , \389_b0 );
not ( \389_b0 , w_939 );
and ( w_939 , w_938 , \389_b1 );
buf ( \391_b1 , \390_b1 );
not ( \391_b1 , w_940 );
not ( \391_b0 , w_941 );
and ( w_940 , w_941 , \390_b0 );
or ( \392_b1 , \372_b1 , w_942 );
or ( \392_b0 , \372_b0 , \391_b0 );
not ( \391_b0 , w_943 );
and ( w_943 , w_942 , \391_b1 );
buf ( \393_b1 , \370_b1 );
not ( \393_b1 , w_944 );
not ( \393_b0 , w_945 );
and ( w_944 , w_945 , \370_b0 );
or ( \394_b1 , \393_b1 , w_946 );
or ( \394_b0 , \393_b0 , \390_b0 );
not ( \390_b0 , w_947 );
and ( w_947 , w_946 , \390_b1 );
or ( \395_b1 , \392_b1 , w_949 );
not ( w_949 , w_950 );
and ( \395_b0 , \392_b0 , w_951 );
and ( w_950 ,  , w_951 );
buf ( w_949 , \394_b1 );
not ( w_949 , w_952 );
not (  , w_953 );
and ( w_952 , w_953 , \394_b0 );
buf ( \396_b1 , \395_b1 );
not ( \396_b1 , w_954 );
not ( \396_b0 , w_955 );
and ( w_954 , w_955 , \395_b0 );
or ( \397_b1 , \a[0]_b1 , \b[9]_b1 );
xor ( \397_b0 , \a[0]_b0 , w_956 );
not ( w_956 , w_957 );
and ( w_957 , \b[9]_b1 , \b[9]_b0 );
buf ( \398_b1 , \397_b1 );
not ( \398_b1 , w_958 );
not ( \398_b0 , w_959 );
and ( w_958 , w_959 , \397_b0 );
or ( \399_b1 , \b[9]_b1 , w_960 );
xor ( \399_b0 , \b[9]_b0 , w_962 );
not ( w_962 , w_963 );
and ( w_963 , w_960 , w_961 );
buf ( w_960 , \b[8]_b1 );
not ( w_960 , w_964 );
not ( w_961 , w_965 );
and ( w_964 , w_965 , \b[8]_b0 );
or ( \400_b1 , \b[8]_b1 , \b[7]_b1 );
xor ( \400_b0 , \b[8]_b0 , w_966 );
not ( w_966 , w_967 );
and ( w_967 , \b[7]_b1 , \b[7]_b0 );
or ( \401_b1 , \399_b1 , w_969 );
not ( w_969 , w_970 );
and ( \401_b0 , \399_b0 , w_971 );
and ( w_970 ,  , w_971 );
buf ( w_969 , \400_b1 );
not ( w_969 , w_972 );
not (  , w_973 );
and ( w_972 , w_973 , \400_b0 );
buf ( \402_b1 , \401_b1 );
not ( \402_b1 , w_974 );
not ( \402_b0 , w_975 );
and ( w_974 , w_975 , \401_b0 );
or ( \403_b1 , \398_b1 , w_976 );
or ( \403_b0 , \398_b0 , \402_b0 );
not ( \402_b0 , w_977 );
and ( w_977 , w_976 , \402_b1 );
or ( \404_b1 , \a[1]_b1 , \b[9]_b1 );
xor ( \404_b0 , \a[1]_b0 , w_978 );
not ( w_978 , w_979 );
and ( w_979 , \b[9]_b1 , \b[9]_b0 );
or ( \405_b1 , \400_b1 , w_981 );
not ( w_981 , w_982 );
and ( \405_b0 , \400_b0 , w_983 );
and ( w_982 ,  , w_983 );
buf ( w_981 , \404_b1 );
not ( w_981 , w_984 );
not (  , w_985 );
and ( w_984 , w_985 , \404_b0 );
or ( \406_b1 , \403_b1 , w_987 );
not ( w_987 , w_988 );
and ( \406_b0 , \403_b0 , w_989 );
and ( w_988 ,  , w_989 );
buf ( w_987 , \405_b1 );
not ( w_987 , w_990 );
not (  , w_991 );
and ( w_990 , w_991 , \405_b0 );
buf ( \407_b1 , \406_b1 );
not ( \407_b1 , w_992 );
not ( \407_b0 , w_993 );
and ( w_992 , w_993 , \406_b0 );
buf ( \408_b1 , \407_b1 );
not ( \408_b1 , w_994 );
not ( \408_b0 , w_995 );
and ( w_994 , w_995 , \407_b0 );
or ( \409_b1 , \a[0]_b1 , w_996 );
or ( \409_b0 , \a[0]_b0 , \b[8]_b0 );
not ( \b[8]_b0 , w_997 );
and ( w_997 , w_996 , \b[8]_b1 );
or ( \410_b1 , \409_b1 , w_999 );
not ( w_999 , w_1000 );
and ( \410_b0 , \409_b0 , w_1001 );
and ( w_1000 ,  , w_1001 );
buf ( w_999 , \b[7]_b1 );
not ( w_999 , w_1002 );
not (  , w_1003 );
and ( w_1002 , w_1003 , \b[7]_b0 );
or ( \411_b1 , \a[0]_b1 , w_1005 );
not ( w_1005 , w_1006 );
and ( \411_b0 , \a[0]_b0 , w_1007 );
and ( w_1006 ,  , w_1007 );
buf ( w_1005 , \b[8]_b1 );
not ( w_1005 , w_1008 );
not (  , w_1009 );
and ( w_1008 , w_1009 , \b[8]_b0 );
buf ( \413_b1 , \382_b1 );
not ( \413_b1 , w_1010 );
not ( \413_b0 , w_1011 );
and ( w_1010 , w_1011 , \382_b0 );
buf ( \414_b1 , \136_b1 );
not ( \414_b1 , w_1012 );
not ( \414_b0 , w_1013 );
and ( w_1012 , w_1013 , \136_b0 );
or ( \415_b1 , \413_b1 , w_1014 );
or ( \415_b0 , \413_b0 , \414_b0 );
not ( \414_b0 , w_1015 );
and ( w_1015 , w_1014 , \414_b1 );
or ( \416_b1 , \a[5]_b1 , \b[5]_b1 );
xor ( \416_b0 , \a[5]_b0 , w_1016 );
not ( w_1016 , w_1017 );
and ( w_1017 , \b[5]_b1 , \b[5]_b0 );
or ( \417_b1 , \139_b1 , w_1019 );
not ( w_1019 , w_1020 );
and ( \417_b0 , \139_b0 , w_1021 );
and ( w_1020 ,  , w_1021 );
buf ( w_1019 , \416_b1 );
not ( w_1019 , w_1022 );
not (  , w_1023 );
and ( w_1022 , w_1023 , \416_b0 );
or ( \418_b1 , \415_b1 , w_1025 );
not ( w_1025 , w_1026 );
and ( \418_b0 , \415_b0 , w_1027 );
and ( w_1026 ,  , w_1027 );
buf ( w_1025 , \417_b1 );
not ( w_1025 , w_1028 );
not (  , w_1029 );
and ( w_1028 , w_1029 , \417_b0 );
or ( \419_b1 , \412_b1 , \418_b1 );
xor ( \419_b0 , \412_b0 , w_1030 );
not ( w_1030 , w_1031 );
and ( w_1031 , \418_b1 , \418_b0 );
buf ( \420_b1 , \419_b1 );
not ( \420_b1 , w_1032 );
not ( \420_b0 , w_1033 );
and ( w_1032 , w_1033 , \419_b0 );
or ( \421_b1 , \408_b1 , w_1034 );
or ( \421_b0 , \408_b0 , \420_b0 );
not ( \420_b0 , w_1035 );
and ( w_1035 , w_1034 , \420_b1 );
or ( \422_b1 , \419_b1 , w_1036 );
or ( \422_b0 , \419_b0 , \407_b0 );
not ( \407_b0 , w_1037 );
and ( w_1037 , w_1036 , \407_b1 );
or ( \423_b1 , \421_b1 , w_1039 );
not ( w_1039 , w_1040 );
and ( \423_b0 , \421_b0 , w_1041 );
and ( w_1040 ,  , w_1041 );
buf ( w_1039 , \422_b1 );
not ( w_1039 , w_1042 );
not (  , w_1043 );
and ( w_1042 , w_1043 , \422_b0 );
or ( \424_b1 , \400_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_1044 );
and ( \424_b0 , \400_b0 , w_1045 );
and ( w_1044 , w_1045 , \a[0]_b0 );
buf ( \425_b1 , \179_b1 );
not ( \425_b1 , w_1046 );
not ( \425_b0 , w_1047 );
and ( w_1046 , w_1047 , \179_b0 );
buf ( \426_b1 , \120_b1 );
not ( \426_b1 , w_1048 );
not ( \426_b0 , w_1049 );
and ( w_1048 , w_1049 , \120_b0 );
or ( \427_b1 , \425_b1 , w_1050 );
or ( \427_b0 , \425_b0 , \426_b0 );
not ( \426_b0 , w_1051 );
and ( w_1051 , w_1050 , \426_b1 );
or ( \428_b1 , \349_b1 , w_1053 );
not ( w_1053 , w_1054 );
and ( \428_b0 , \349_b0 , w_1055 );
and ( w_1054 ,  , w_1055 );
buf ( w_1053 , \b[0]_b1 );
not ( w_1053 , w_1056 );
not (  , w_1057 );
and ( w_1056 , w_1057 , \b[0]_b0 );
or ( \429_b1 , \427_b1 , w_1059 );
not ( w_1059 , w_1060 );
and ( \429_b0 , \427_b0 , w_1061 );
and ( w_1060 ,  , w_1061 );
buf ( w_1059 , \428_b1 );
not ( w_1059 , w_1062 );
not (  , w_1063 );
and ( w_1062 , w_1063 , \428_b0 );
or ( \430_b1 , \424_b1 , \429_b1 );
xor ( \430_b0 , \424_b0 , w_1064 );
not ( w_1064 , w_1065 );
and ( w_1065 , \429_b1 , \429_b0 );
buf ( \431_b1 , \164_b1 );
not ( \431_b1 , w_1066 );
not ( \431_b0 , w_1067 );
and ( w_1066 , w_1067 , \164_b0 );
buf ( \432_b1 , \295_b1 );
not ( \432_b1 , w_1068 );
not ( \432_b0 , w_1069 );
and ( w_1068 , w_1069 , \295_b0 );
or ( \433_b1 , \431_b1 , w_1070 );
or ( \433_b0 , \431_b0 , \432_b0 );
not ( \432_b0 , w_1071 );
and ( w_1071 , w_1070 , \432_b1 );
or ( \434_b1 , \147_b1 , w_1073 );
not ( w_1073 , w_1074 );
and ( \434_b0 , \147_b0 , w_1075 );
and ( w_1074 ,  , w_1075 );
buf ( w_1073 , \363_b1 );
not ( w_1073 , w_1076 );
not (  , w_1077 );
and ( w_1076 , w_1077 , \363_b0 );
or ( \435_b1 , \433_b1 , w_1079 );
not ( w_1079 , w_1080 );
and ( \435_b0 , \433_b0 , w_1081 );
and ( w_1080 ,  , w_1081 );
buf ( w_1079 , \434_b1 );
not ( w_1079 , w_1082 );
not (  , w_1083 );
and ( w_1082 , w_1083 , \434_b0 );
or ( \436_b1 , \430_b1 , \435_b1 );
not ( \435_b1 , w_1084 );
and ( \436_b0 , \430_b0 , w_1085 );
and ( w_1084 , w_1085 , \435_b0 );
or ( \437_b1 , \424_b1 , \429_b1 );
not ( \429_b1 , w_1086 );
and ( \437_b0 , \424_b0 , w_1087 );
and ( w_1086 , w_1087 , \429_b0 );
or ( \438_b1 , \436_b1 , w_1088 );
or ( \438_b0 , \436_b0 , \437_b0 );
not ( \437_b0 , w_1089 );
and ( w_1089 , w_1088 , \437_b1 );
or ( \439_b1 , \423_b1 , w_1090 );
xor ( \439_b0 , \423_b0 , w_1092 );
not ( w_1092 , w_1093 );
and ( w_1093 , w_1090 , w_1091 );
buf ( w_1090 , \438_b1 );
not ( w_1090 , w_1094 );
not ( w_1091 , w_1095 );
and ( w_1094 , w_1095 , \438_b0 );
buf ( \440_b1 , \439_b1 );
not ( \440_b1 , w_1096 );
not ( \440_b0 , w_1097 );
and ( w_1096 , w_1097 , \439_b0 );
or ( \441_b1 , \396_b1 , \440_b1 );
not ( \440_b1 , w_1098 );
and ( \441_b0 , \396_b0 , w_1099 );
and ( w_1098 , w_1099 , \440_b0 );
or ( \442_b1 , \439_b1 , \395_b1 );
not ( \395_b1 , w_1100 );
and ( \442_b0 , \439_b0 , w_1101 );
and ( w_1100 , w_1101 , \395_b0 );
or ( \443_b1 , \441_b1 , w_1103 );
not ( w_1103 , w_1104 );
and ( \443_b0 , \441_b0 , w_1105 );
and ( w_1104 ,  , w_1105 );
buf ( w_1103 , \442_b1 );
not ( w_1103 , w_1106 );
not (  , w_1107 );
and ( w_1106 , w_1107 , \442_b0 );
or ( \444_b1 , \424_b1 , \429_b1 );
xor ( \444_b0 , \424_b0 , w_1108 );
not ( w_1108 , w_1109 );
and ( w_1109 , \429_b1 , \429_b0 );
or ( \445_b1 , \444_b1 , \435_b1 );
xor ( \445_b0 , \444_b0 , w_1110 );
not ( w_1110 , w_1111 );
and ( w_1111 , \435_b1 , \435_b0 );
buf ( \446_b1 , \445_b1 );
not ( \446_b1 , w_1112 );
not ( \446_b0 , w_1113 );
and ( w_1112 , w_1113 , \445_b0 );
buf ( \447_b1 , \446_b1 );
not ( \447_b1 , w_1114 );
not ( \447_b0 , w_1115 );
and ( w_1114 , w_1115 , \446_b0 );
or ( \448_b1 , \181_b1 , \191_b1 );
xor ( \448_b0 , \181_b0 , w_1116 );
not ( w_1116 , w_1117 );
and ( w_1117 , \191_b1 , \191_b0 );
or ( \449_b1 , \448_b1 , \200_b1 );
not ( \200_b1 , w_1118 );
and ( \449_b0 , \448_b0 , w_1119 );
and ( w_1118 , w_1119 , \200_b0 );
or ( \450_b1 , \181_b1 , \191_b1 );
not ( \191_b1 , w_1120 );
and ( \450_b0 , \181_b0 , w_1121 );
and ( w_1120 , w_1121 , \191_b0 );
or ( \451_b1 , \449_b1 , w_1122 );
or ( \451_b0 , \449_b0 , \450_b0 );
not ( \450_b0 , w_1123 );
and ( w_1123 , w_1122 , \450_b1 );
buf ( \452_b1 , \451_b1 );
not ( \452_b1 , w_1124 );
not ( \452_b0 , w_1125 );
and ( w_1124 , w_1125 , \451_b0 );
buf ( \453_b1 , \452_b1 );
not ( \453_b1 , w_1126 );
not ( \453_b0 , w_1127 );
and ( w_1126 , w_1127 , \452_b0 );
or ( \454_b1 , \447_b1 , w_1128 );
or ( \454_b0 , \447_b0 , \453_b0 );
not ( \453_b0 , w_1129 );
and ( w_1129 , w_1128 , \453_b1 );
or ( \455_b1 , \378_b1 , \384_b1 );
xor ( \455_b0 , \378_b0 , w_1130 );
not ( w_1130 , w_1131 );
and ( w_1131 , \384_b1 , \384_b0 );
or ( \456_b1 , \455_b1 , \387_b1 );
xor ( \456_b0 , \455_b0 , w_1132 );
not ( w_1132 , w_1133 );
and ( w_1133 , \387_b1 , \387_b0 );
or ( \457_b1 , \454_b1 , w_1135 );
not ( w_1135 , w_1136 );
and ( \457_b0 , \454_b0 , w_1137 );
and ( w_1136 ,  , w_1137 );
buf ( w_1135 , \456_b1 );
not ( w_1135 , w_1138 );
not (  , w_1139 );
and ( w_1138 , w_1139 , \456_b0 );
buf ( \458_b1 , \446_b1 );
not ( \458_b1 , w_1140 );
not ( \458_b0 , w_1141 );
and ( w_1140 , w_1141 , \446_b0 );
or ( \459_b1 , \458_b1 , w_1143 );
not ( w_1143 , w_1144 );
and ( \459_b0 , \458_b0 , w_1145 );
and ( w_1144 ,  , w_1145 );
buf ( w_1143 , \451_b1 );
not ( w_1143 , w_1146 );
not (  , w_1147 );
and ( w_1146 , w_1147 , \451_b0 );
or ( \460_b1 , \457_b1 , w_1149 );
not ( w_1149 , w_1150 );
and ( \460_b0 , \457_b0 , w_1151 );
and ( w_1150 ,  , w_1151 );
buf ( w_1149 , \459_b1 );
not ( w_1149 , w_1152 );
not (  , w_1153 );
and ( w_1152 , w_1153 , \459_b0 );
buf ( \461_b1 , \460_b1 );
not ( \461_b1 , w_1154 );
not ( \461_b0 , w_1155 );
and ( w_1154 , w_1155 , \460_b0 );
or ( \462_b1 , \443_b1 , w_1157 );
not ( w_1157 , w_1158 );
and ( \462_b0 , \443_b0 , w_1159 );
and ( w_1158 ,  , w_1159 );
buf ( w_1157 , \461_b1 );
not ( w_1157 , w_1160 );
not (  , w_1161 );
and ( w_1160 , w_1161 , \461_b0 );
or ( \463_b1 , \445_b1 , \452_b1 );
xor ( \463_b0 , \445_b0 , w_1162 );
not ( w_1162 , w_1163 );
and ( w_1163 , \452_b1 , \452_b0 );
or ( \464_b1 , \463_b1 , \456_b1 );
xor ( \464_b0 , \463_b0 , w_1164 );
not ( w_1164 , w_1165 );
and ( w_1165 , \456_b1 , \456_b0 );
or ( \465_b1 , \170_b1 , \174_b1 );
xor ( \465_b0 , \170_b0 , w_1166 );
not ( w_1166 , w_1167 );
and ( w_1167 , \174_b1 , \174_b0 );
or ( \466_b1 , \465_b1 , \201_b1 );
not ( \201_b1 , w_1168 );
and ( \466_b0 , \465_b0 , w_1169 );
and ( w_1168 , w_1169 , \201_b0 );
or ( \467_b1 , \170_b1 , \174_b1 );
not ( \174_b1 , w_1170 );
and ( \467_b0 , \170_b0 , w_1171 );
and ( w_1170 , w_1171 , \174_b0 );
or ( \468_b1 , \466_b1 , w_1172 );
or ( \468_b0 , \466_b0 , \467_b0 );
not ( \467_b0 , w_1173 );
and ( w_1173 , w_1172 , \467_b1 );
buf ( \469_b1 , \468_b1 );
not ( \469_b1 , w_1174 );
not ( \469_b0 , w_1175 );
and ( w_1174 , w_1175 , \468_b0 );
or ( \470_b1 , \464_b1 , w_1177 );
not ( w_1177 , w_1178 );
and ( \470_b0 , \464_b0 , w_1179 );
and ( w_1178 ,  , w_1179 );
buf ( w_1177 , \469_b1 );
not ( w_1177 , w_1180 );
not (  , w_1181 );
and ( w_1180 , w_1181 , \469_b0 );
or ( \471_b1 , \462_b1 , \470_b1 );
not ( \470_b1 , w_1182 );
and ( \471_b0 , \462_b0 , w_1183 );
and ( w_1182 , w_1183 , \470_b0 );
buf ( \472_b1 , \374_b1 );
not ( \472_b1 , w_1184 );
not ( \472_b0 , w_1185 );
and ( w_1184 , w_1185 , \374_b0 );
buf ( \473_b1 , \359_b1 );
not ( \473_b1 , w_1186 );
not ( \473_b0 , w_1187 );
and ( w_1186 , w_1187 , \359_b0 );
or ( \474_b1 , \472_b1 , w_1188 );
or ( \474_b0 , \472_b0 , \473_b0 );
not ( \473_b0 , w_1189 );
and ( w_1189 , w_1188 , \473_b1 );
or ( \475_b1 , \a[4]_b1 , \b[7]_b1 );
xor ( \475_b0 , \a[4]_b0 , w_1190 );
not ( w_1190 , w_1191 );
and ( w_1191 , \b[7]_b1 , \b[7]_b0 );
or ( \476_b1 , \129_b1 , w_1193 );
not ( w_1193 , w_1194 );
and ( \476_b0 , \129_b0 , w_1195 );
and ( w_1194 ,  , w_1195 );
buf ( w_1193 , \475_b1 );
not ( w_1193 , w_1196 );
not (  , w_1197 );
and ( w_1196 , w_1197 , \475_b0 );
or ( \477_b1 , \474_b1 , w_1199 );
not ( w_1199 , w_1200 );
and ( \477_b0 , \474_b0 , w_1201 );
and ( w_1200 ,  , w_1201 );
buf ( w_1199 , \476_b1 );
not ( w_1199 , w_1202 );
not (  , w_1203 );
and ( w_1202 , w_1203 , \476_b0 );
buf ( \478_b1 , \404_b1 );
not ( \478_b1 , w_1204 );
not ( \478_b0 , w_1205 );
and ( w_1204 , w_1205 , \404_b0 );
buf ( \479_b1 , \401_b1 );
not ( \479_b1 , w_1206 );
not ( \479_b0 , w_1207 );
and ( w_1206 , w_1207 , \401_b0 );
or ( \480_b1 , \478_b1 , w_1208 );
or ( \480_b0 , \478_b0 , \479_b0 );
not ( \479_b0 , w_1209 );
and ( w_1209 , w_1208 , \479_b1 );
or ( \481_b1 , \a[2]_b1 , \b[9]_b1 );
xor ( \481_b0 , \a[2]_b0 , w_1210 );
not ( w_1210 , w_1211 );
and ( w_1211 , \b[9]_b1 , \b[9]_b0 );
or ( \482_b1 , \400_b1 , w_1213 );
not ( w_1213 , w_1214 );
and ( \482_b0 , \400_b0 , w_1215 );
and ( w_1214 ,  , w_1215 );
buf ( w_1213 , \481_b1 );
not ( w_1213 , w_1216 );
not (  , w_1217 );
and ( w_1216 , w_1217 , \481_b0 );
or ( \483_b1 , \480_b1 , w_1219 );
not ( w_1219 , w_1220 );
and ( \483_b0 , \480_b0 , w_1221 );
and ( w_1220 ,  , w_1221 );
buf ( w_1219 , \482_b1 );
not ( w_1219 , w_1222 );
not (  , w_1223 );
and ( w_1222 , w_1223 , \482_b0 );
or ( \484_b1 , \477_b1 , \483_b1 );
xor ( \484_b0 , \477_b0 , w_1224 );
not ( w_1224 , w_1225 );
and ( w_1225 , \483_b1 , \483_b0 );
buf ( \485_b1 , \367_b1 );
not ( \485_b1 , w_1226 );
not ( \485_b0 , w_1227 );
and ( w_1226 , w_1227 , \367_b0 );
buf ( \486_b1 , \295_b1 );
buf ( \486_b0 , \295_b0 );
buf ( \487_b1 , \486_b1 );
not ( \487_b1 , w_1228 );
not ( \487_b0 , w_1229 );
and ( w_1228 , w_1229 , \486_b0 );
or ( \488_b1 , \485_b1 , w_1230 );
or ( \488_b0 , \485_b0 , \487_b0 );
not ( \487_b0 , w_1231 );
and ( w_1231 , w_1230 , \487_b1 );
or ( \489_b1 , \a[8]_b1 , \b[3]_b1 );
xor ( \489_b0 , \a[8]_b0 , w_1232 );
not ( w_1232 , w_1233 );
and ( w_1233 , \b[3]_b1 , \b[3]_b0 );
or ( \490_b1 , \147_b1 , w_1235 );
not ( w_1235 , w_1236 );
and ( \490_b0 , \147_b0 , w_1237 );
and ( w_1236 ,  , w_1237 );
buf ( w_1235 , \489_b1 );
not ( w_1235 , w_1238 );
not (  , w_1239 );
and ( w_1238 , w_1239 , \489_b0 );
or ( \491_b1 , \488_b1 , w_1241 );
not ( w_1241 , w_1242 );
and ( \491_b0 , \488_b0 , w_1243 );
and ( w_1242 ,  , w_1243 );
buf ( w_1241 , \490_b1 );
not ( w_1241 , w_1244 );
not (  , w_1245 );
and ( w_1244 , w_1245 , \490_b0 );
or ( \492_b1 , \484_b1 , \491_b1 );
xor ( \492_b0 , \484_b0 , w_1246 );
not ( w_1246 , w_1247 );
and ( w_1247 , \491_b1 , \491_b0 );
buf ( \493_b1 , \406_b1 );
not ( \493_b1 , w_1248 );
not ( \493_b0 , w_1249 );
and ( w_1248 , w_1249 , \406_b0 );
buf ( \494_b1 , \419_b1 );
not ( \494_b1 , w_1250 );
not ( \494_b0 , w_1251 );
and ( w_1250 , w_1251 , \419_b0 );
or ( \495_b1 , \493_b1 , w_1252 );
or ( \495_b0 , \493_b0 , \494_b0 );
not ( \494_b0 , w_1253 );
and ( w_1253 , w_1252 , \494_b1 );
or ( \496_b1 , \419_b1 , w_1254 );
or ( \496_b0 , \419_b0 , \406_b0 );
not ( \406_b0 , w_1255 );
and ( w_1255 , w_1254 , \406_b1 );
or ( \497_b1 , \496_b1 , w_1257 );
not ( w_1257 , w_1258 );
and ( \497_b0 , \496_b0 , w_1259 );
and ( w_1258 ,  , w_1259 );
buf ( w_1257 , \438_b1 );
not ( w_1257 , w_1260 );
not (  , w_1261 );
and ( w_1260 , w_1261 , \438_b0 );
or ( \498_b1 , \495_b1 , w_1263 );
not ( w_1263 , w_1264 );
and ( \498_b0 , \495_b0 , w_1265 );
and ( w_1264 ,  , w_1265 );
buf ( w_1263 , \497_b1 );
not ( w_1263 , w_1266 );
not (  , w_1267 );
and ( w_1266 , w_1267 , \497_b0 );
or ( \499_b1 , \492_b1 , \498_b1 );
xor ( \499_b0 , \492_b0 , w_1268 );
not ( w_1268 , w_1269 );
and ( w_1269 , \498_b1 , \498_b0 );
or ( \500_b1 , \412_b1 , \418_b1 );
not ( \418_b1 , w_1270 );
and ( \500_b0 , \412_b0 , w_1271 );
and ( w_1270 , w_1271 , \418_b0 );
or ( \501_b1 , \354_b1 , \361_b1 );
xor ( \501_b0 , \354_b0 , w_1272 );
not ( w_1272 , w_1273 );
and ( w_1273 , \361_b1 , \361_b0 );
or ( \502_b1 , \501_b1 , \369_b1 );
not ( \369_b1 , w_1274 );
and ( \502_b0 , \501_b0 , w_1275 );
and ( w_1274 , w_1275 , \369_b0 );
or ( \503_b1 , \354_b1 , \361_b1 );
not ( \361_b1 , w_1276 );
and ( \503_b0 , \354_b0 , w_1277 );
and ( w_1276 , w_1277 , \361_b0 );
or ( \504_b1 , \502_b1 , w_1278 );
or ( \504_b0 , \502_b0 , \503_b0 );
not ( \503_b0 , w_1279 );
and ( w_1279 , w_1278 , \503_b1 );
or ( \505_b1 , \500_b1 , \504_b1 );
xor ( \505_b0 , \500_b0 , w_1280 );
not ( w_1280 , w_1281 );
and ( w_1281 , \504_b1 , \504_b0 );
or ( \506_b1 , \b[10]_b1 , \b[9]_b1 );
xor ( \506_b0 , \b[10]_b0 , w_1282 );
not ( w_1282 , w_1283 );
and ( w_1283 , \b[9]_b1 , \b[9]_b0 );
or ( \507_b1 , \506_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_1284 );
and ( \507_b0 , \506_b0 , w_1285 );
and ( w_1284 , w_1285 , \a[0]_b0 );
buf ( \508_b1 , \352_b1 );
not ( \508_b1 , w_1286 );
not ( \508_b0 , w_1287 );
and ( w_1286 , w_1287 , \352_b0 );
buf ( \509_b1 , \120_b1 );
not ( \509_b1 , w_1288 );
not ( \509_b0 , w_1289 );
and ( w_1288 , w_1289 , \120_b0 );
or ( \510_b1 , \508_b1 , w_1290 );
or ( \510_b0 , \508_b0 , \509_b0 );
not ( \509_b0 , w_1291 );
and ( w_1291 , w_1290 , \509_b1 );
or ( \511_b1 , \a[10]_b1 , \b[1]_b1 );
xor ( \511_b0 , \a[10]_b0 , w_1292 );
not ( w_1292 , w_1293 );
and ( w_1293 , \b[1]_b1 , \b[1]_b0 );
or ( \512_b1 , \b[0]_b1 , w_1295 );
not ( w_1295 , w_1296 );
and ( \512_b0 , \b[0]_b0 , w_1297 );
and ( w_1296 ,  , w_1297 );
buf ( w_1295 , \511_b1 );
not ( w_1295 , w_1298 );
not (  , w_1299 );
and ( w_1298 , w_1299 , \511_b0 );
or ( \513_b1 , \510_b1 , w_1301 );
not ( w_1301 , w_1302 );
and ( \513_b0 , \510_b0 , w_1303 );
and ( w_1302 ,  , w_1303 );
buf ( w_1301 , \512_b1 );
not ( w_1301 , w_1304 );
not (  , w_1305 );
and ( w_1304 , w_1305 , \512_b0 );
or ( \514_b1 , \507_b1 , \513_b1 );
xor ( \514_b0 , \507_b0 , w_1306 );
not ( w_1306 , w_1307 );
and ( w_1307 , \513_b1 , \513_b0 );
buf ( \515_b1 , \195_b1 );
not ( \515_b1 , w_1308 );
not ( \515_b0 , w_1309 );
and ( w_1308 , w_1309 , \195_b0 );
buf ( \516_b1 , \416_b1 );
not ( \516_b1 , w_1310 );
not ( \516_b0 , w_1311 );
and ( w_1310 , w_1311 , \416_b0 );
or ( \517_b1 , \515_b1 , w_1312 );
or ( \517_b0 , \515_b0 , \516_b0 );
not ( \516_b0 , w_1313 );
and ( w_1313 , w_1312 , \516_b1 );
or ( \518_b1 , \a[6]_b1 , \b[5]_b1 );
xor ( \518_b0 , \a[6]_b0 , w_1314 );
not ( w_1314 , w_1315 );
and ( w_1315 , \b[5]_b1 , \b[5]_b0 );
or ( \519_b1 , \139_b1 , w_1317 );
not ( w_1317 , w_1318 );
and ( \519_b0 , \139_b0 , w_1319 );
and ( w_1318 ,  , w_1319 );
buf ( w_1317 , \518_b1 );
not ( w_1317 , w_1320 );
not (  , w_1321 );
and ( w_1320 , w_1321 , \518_b0 );
or ( \520_b1 , \517_b1 , w_1323 );
not ( w_1323 , w_1324 );
and ( \520_b0 , \517_b0 , w_1325 );
and ( w_1324 ,  , w_1325 );
buf ( w_1323 , \519_b1 );
not ( w_1323 , w_1326 );
not (  , w_1327 );
and ( w_1326 , w_1327 , \519_b0 );
or ( \521_b1 , \514_b1 , \520_b1 );
xor ( \521_b0 , \514_b0 , w_1328 );
not ( w_1328 , w_1329 );
and ( w_1329 , \520_b1 , \520_b0 );
or ( \522_b1 , \505_b1 , \521_b1 );
xor ( \522_b0 , \505_b0 , w_1330 );
not ( w_1330 , w_1331 );
and ( w_1331 , \521_b1 , \521_b0 );
or ( \523_b1 , \499_b1 , w_1332 );
xor ( \523_b0 , \499_b0 , w_1334 );
not ( w_1334 , w_1335 );
and ( w_1335 , w_1332 , w_1333 );
buf ( w_1332 , \522_b1 );
not ( w_1332 , w_1336 );
not ( w_1333 , w_1337 );
and ( w_1336 , w_1337 , \522_b0 );
buf ( \524_b1 , \393_b1 );
not ( \524_b1 , w_1338 );
not ( \524_b0 , w_1339 );
and ( w_1338 , w_1339 , \393_b0 );
buf ( \525_b1 , \439_b1 );
not ( \525_b1 , w_1340 );
not ( \525_b0 , w_1341 );
and ( w_1340 , w_1341 , \439_b0 );
or ( \526_b1 , \524_b1 , w_1342 );
or ( \526_b0 , \524_b0 , \525_b0 );
not ( \525_b0 , w_1343 );
and ( w_1343 , w_1342 , \525_b1 );
buf ( \527_b1 , \390_b1 );
buf ( \527_b0 , \390_b0 );
or ( \528_b1 , \526_b1 , w_1345 );
not ( w_1345 , w_1346 );
and ( \528_b0 , \526_b0 , w_1347 );
and ( w_1346 ,  , w_1347 );
buf ( w_1345 , \527_b1 );
not ( w_1345 , w_1348 );
not (  , w_1349 );
and ( w_1348 , w_1349 , \527_b0 );
or ( \529_b1 , \439_b1 , w_1350 );
or ( \529_b0 , \439_b0 , \393_b0 );
not ( \393_b0 , w_1351 );
and ( w_1351 , w_1350 , \393_b1 );
or ( \530_b1 , \528_b1 , w_1353 );
not ( w_1353 , w_1354 );
and ( \530_b0 , \528_b0 , w_1355 );
and ( w_1354 ,  , w_1355 );
buf ( w_1353 , \529_b1 );
not ( w_1353 , w_1356 );
not (  , w_1357 );
and ( w_1356 , w_1357 , \529_b0 );
buf ( \531_b1 , \530_b1 );
not ( \531_b1 , w_1358 );
not ( \531_b0 , w_1359 );
and ( w_1358 , w_1359 , \530_b0 );
or ( \532_b1 , \523_b1 , w_1361 );
not ( w_1361 , w_1362 );
and ( \532_b0 , \523_b0 , w_1363 );
and ( w_1362 ,  , w_1363 );
buf ( w_1361 , \531_b1 );
not ( w_1361 , w_1364 );
not (  , w_1365 );
and ( w_1364 , w_1365 , \531_b0 );
buf ( \534_b1 , \460_b1 );
not ( \534_b1 , w_1366 );
not ( \534_b0 , w_1367 );
and ( w_1366 , w_1367 , \460_b0 );
buf ( \535_b1 , \443_b1 );
not ( \535_b1 , w_1368 );
not ( \535_b0 , w_1369 );
and ( w_1368 , w_1369 , \443_b0 );
buf ( \536_b1 , \535_b1 );
not ( \536_b1 , w_1370 );
not ( \536_b0 , w_1371 );
and ( w_1370 , w_1371 , \535_b0 );
or ( \537_b1 , \534_b1 , w_1372 );
or ( \537_b0 , \534_b0 , \536_b0 );
not ( \536_b0 , w_1373 );
and ( w_1373 , w_1372 , \536_b1 );
buf ( \538_b1 , \469_b1 );
not ( \538_b1 , w_1374 );
not ( \538_b0 , w_1375 );
and ( w_1374 , w_1375 , \469_b0 );
buf ( \539_b1 , \464_b1 );
not ( \539_b1 , w_1376 );
not ( \539_b0 , w_1377 );
and ( w_1376 , w_1377 , \464_b0 );
or ( \540_b1 , \538_b1 , w_1379 );
not ( w_1379 , w_1380 );
and ( \540_b0 , \538_b0 , w_1381 );
and ( w_1380 ,  , w_1381 );
buf ( w_1379 , \539_b1 );
not ( w_1379 , w_1382 );
not (  , w_1383 );
and ( w_1382 , w_1383 , \539_b0 );
or ( \541_b1 , \537_b1 , w_1385 );
not ( w_1385 , w_1386 );
and ( \541_b0 , \537_b0 , w_1387 );
and ( w_1386 ,  , w_1387 );
buf ( w_1385 , \540_b1 );
not ( w_1385 , w_1388 );
not (  , w_1389 );
and ( w_1388 , w_1389 , \540_b0 );
buf ( \542_b1 , \462_b1 );
buf ( \542_b0 , \462_b0 );
buf ( \544_b1 , \523_b1 );
not ( \544_b1 , w_1390 );
not ( \544_b0 , w_1391 );
and ( w_1390 , w_1391 , \523_b0 );
buf ( \545_b1 , \531_b1 );
not ( \545_b1 , w_1392 );
not ( \545_b0 , w_1393 );
and ( w_1392 , w_1393 , \531_b0 );
or ( \546_b1 , \544_b1 , w_1395 );
not ( w_1395 , w_1396 );
and ( \546_b0 , \544_b0 , w_1397 );
and ( w_1396 ,  , w_1397 );
buf ( w_1395 , \545_b1 );
not ( w_1395 , w_1398 );
not (  , w_1399 );
and ( w_1398 , w_1399 , \545_b0 );
or ( \548_b1 , \522_b1 , w_1401 );
not ( w_1401 , w_1402 );
and ( \548_b0 , \522_b0 , w_1403 );
and ( w_1402 ,  , w_1403 );
buf ( w_1401 , \492_b1 );
not ( w_1401 , w_1404 );
not (  , w_1405 );
and ( w_1404 , w_1405 , \492_b0 );
or ( \549_b1 , \522_b1 , w_1406 );
or ( \549_b0 , \522_b0 , \492_b0 );
not ( \492_b0 , w_1407 );
and ( w_1407 , w_1406 , \492_b1 );
or ( \550_b1 , \549_b1 , w_1409 );
not ( w_1409 , w_1410 );
and ( \550_b0 , \549_b0 , w_1411 );
and ( w_1410 ,  , w_1411 );
buf ( w_1409 , \498_b1 );
not ( w_1409 , w_1412 );
not (  , w_1413 );
and ( w_1412 , w_1413 , \498_b0 );
or ( \551_b1 , \548_b1 , w_1415 );
not ( w_1415 , w_1416 );
and ( \551_b0 , \548_b0 , w_1417 );
and ( w_1416 ,  , w_1417 );
buf ( w_1415 , \550_b1 );
not ( w_1415 , w_1418 );
not (  , w_1419 );
and ( w_1418 , w_1419 , \550_b0 );
or ( \552_b1 , \507_b1 , \513_b1 );
xor ( \552_b0 , \507_b0 , w_1420 );
not ( w_1420 , w_1421 );
and ( w_1421 , \513_b1 , \513_b0 );
or ( \553_b1 , \552_b1 , \520_b1 );
not ( \520_b1 , w_1422 );
and ( \553_b0 , \552_b0 , w_1423 );
and ( w_1422 , w_1423 , \520_b0 );
or ( \554_b1 , \507_b1 , \513_b1 );
not ( \513_b1 , w_1424 );
and ( \554_b0 , \507_b0 , w_1425 );
and ( w_1424 , w_1425 , \513_b0 );
or ( \555_b1 , \553_b1 , w_1426 );
or ( \555_b0 , \553_b0 , \554_b0 );
not ( \554_b0 , w_1427 );
and ( w_1427 , w_1426 , \554_b1 );
or ( \556_b1 , \b[11]_b1 , \b[10]_b1 );
xor ( \556_b0 , \b[11]_b0 , w_1428 );
not ( w_1428 , w_1429 );
and ( w_1429 , \b[10]_b1 , \b[10]_b0 );
or ( \557_b1 , \a[0]_b1 , \b[11]_b1 );
xor ( \557_b0 , \a[0]_b0 , w_1430 );
not ( w_1430 , w_1431 );
and ( w_1431 , \b[11]_b1 , \b[11]_b0 );
or ( \558_b1 , \556_b1 , w_1433 );
not ( w_1433 , w_1434 );
and ( \558_b0 , \556_b0 , w_1435 );
and ( w_1434 ,  , w_1435 );
buf ( w_1433 , \557_b1 );
not ( w_1433 , w_1436 );
not (  , w_1437 );
and ( w_1436 , w_1437 , \557_b0 );
or ( \559_b1 , \558_b1 , w_1438 );
or ( \559_b0 , \558_b0 , \506_b0 );
not ( \506_b0 , w_1439 );
and ( w_1439 , w_1438 , \506_b1 );
or ( \560_b1 , \a[1]_b1 , \b[11]_b1 );
xor ( \560_b0 , \a[1]_b0 , w_1440 );
not ( w_1440 , w_1441 );
and ( w_1441 , \b[11]_b1 , \b[11]_b0 );
or ( \561_b1 , \506_b1 , w_1443 );
not ( w_1443 , w_1444 );
and ( \561_b0 , \506_b0 , w_1445 );
and ( w_1444 ,  , w_1445 );
buf ( w_1443 , \560_b1 );
not ( w_1443 , w_1446 );
not (  , w_1447 );
and ( w_1446 , w_1447 , \560_b0 );
or ( \562_b1 , \559_b1 , w_1449 );
not ( w_1449 , w_1450 );
and ( \562_b0 , \559_b0 , w_1451 );
and ( w_1450 ,  , w_1451 );
buf ( w_1449 , \561_b1 );
not ( w_1449 , w_1452 );
not (  , w_1453 );
and ( w_1452 , w_1453 , \561_b0 );
or ( \563_b1 , \a[0]_b1 , w_1454 );
or ( \563_b0 , \a[0]_b0 , \b[10]_b0 );
not ( \b[10]_b0 , w_1455 );
and ( w_1455 , w_1454 , \b[10]_b1 );
or ( \564_b1 , \563_b1 , w_1457 );
not ( w_1457 , w_1458 );
and ( \564_b0 , \563_b0 , w_1459 );
and ( w_1458 ,  , w_1459 );
buf ( w_1457 , \b[9]_b1 );
not ( w_1457 , w_1460 );
not (  , w_1461 );
and ( w_1460 , w_1461 , \b[9]_b0 );
or ( \565_b1 , \a[0]_b1 , w_1463 );
not ( w_1463 , w_1464 );
and ( \565_b0 , \a[0]_b0 , w_1465 );
and ( w_1464 ,  , w_1465 );
buf ( w_1463 , \b[10]_b1 );
not ( w_1463 , w_1466 );
not (  , w_1467 );
and ( w_1466 , w_1467 , \b[10]_b0 );
buf ( \567_b1 , \566_b1 );
not ( \567_b1 , w_1468 );
not ( \567_b0 , w_1469 );
and ( w_1468 , w_1469 , \566_b0 );
or ( \568_b1 , \562_b1 , \567_b1 );
not ( \567_b1 , w_1470 );
and ( \568_b0 , \562_b0 , w_1471 );
and ( w_1470 , w_1471 , \567_b0 );
buf ( \569_b1 , \562_b1 );
not ( \569_b1 , w_1472 );
not ( \569_b0 , w_1473 );
and ( w_1472 , w_1473 , \562_b0 );
or ( \570_b1 , \569_b1 , \566_b1 );
not ( \566_b1 , w_1474 );
and ( \570_b0 , \569_b0 , w_1475 );
and ( w_1474 , w_1475 , \566_b0 );
or ( \571_b1 , \568_b1 , w_1477 );
not ( w_1477 , w_1478 );
and ( \571_b0 , \568_b0 , w_1479 );
and ( w_1478 ,  , w_1479 );
buf ( w_1477 , \570_b1 );
not ( w_1477 , w_1480 );
not (  , w_1481 );
and ( w_1480 , w_1481 , \570_b0 );
buf ( \572_b1 , \511_b1 );
not ( \572_b1 , w_1482 );
not ( \572_b0 , w_1483 );
and ( w_1482 , w_1483 , \511_b0 );
buf ( \573_b1 , \120_b1 );
not ( \573_b1 , w_1484 );
not ( \573_b0 , w_1485 );
and ( w_1484 , w_1485 , \120_b0 );
or ( \574_b1 , \572_b1 , w_1486 );
or ( \574_b0 , \572_b0 , \573_b0 );
not ( \573_b0 , w_1487 );
and ( w_1487 , w_1486 , \573_b1 );
or ( \575_b1 , \a[11]_b1 , \b[1]_b1 );
xor ( \575_b0 , \a[11]_b0 , w_1488 );
not ( w_1488 , w_1489 );
and ( w_1489 , \b[1]_b1 , \b[1]_b0 );
or ( \576_b1 , \575_b1 , w_1491 );
not ( w_1491 , w_1492 );
and ( \576_b0 , \575_b0 , w_1493 );
and ( w_1492 ,  , w_1493 );
buf ( w_1491 , \b[0]_b1 );
not ( w_1491 , w_1494 );
not (  , w_1495 );
and ( w_1494 , w_1495 , \b[0]_b0 );
or ( \577_b1 , \574_b1 , w_1497 );
not ( w_1497 , w_1498 );
and ( \577_b0 , \574_b0 , w_1499 );
and ( w_1498 ,  , w_1499 );
buf ( w_1497 , \576_b1 );
not ( w_1497 , w_1500 );
not (  , w_1501 );
and ( w_1500 , w_1501 , \576_b0 );
buf ( \578_b1 , \577_b1 );
not ( \578_b1 , w_1502 );
not ( \578_b0 , w_1503 );
and ( w_1502 , w_1503 , \577_b0 );
or ( \579_b1 , \571_b1 , \578_b1 );
not ( \578_b1 , w_1504 );
and ( \579_b0 , \571_b0 , w_1505 );
and ( w_1504 , w_1505 , \578_b0 );
buf ( \580_b1 , \571_b1 );
not ( \580_b1 , w_1506 );
not ( \580_b0 , w_1507 );
and ( w_1506 , w_1507 , \571_b0 );
or ( \581_b1 , \580_b1 , \577_b1 );
not ( \577_b1 , w_1508 );
and ( \581_b0 , \580_b0 , w_1509 );
and ( w_1508 , w_1509 , \577_b0 );
or ( \582_b1 , \579_b1 , w_1511 );
not ( w_1511 , w_1512 );
and ( \582_b0 , \579_b0 , w_1513 );
and ( w_1512 ,  , w_1513 );
buf ( w_1511 , \581_b1 );
not ( w_1511 , w_1514 );
not (  , w_1515 );
and ( w_1514 , w_1515 , \581_b0 );
or ( \583_b1 , \555_b1 , \582_b1 );
xor ( \583_b0 , \555_b0 , w_1516 );
not ( w_1516 , w_1517 );
and ( w_1517 , \582_b1 , \582_b0 );
or ( \584_b1 , \477_b1 , \483_b1 );
xor ( \584_b0 , \477_b0 , w_1518 );
not ( w_1518 , w_1519 );
and ( w_1519 , \483_b1 , \483_b0 );
or ( \585_b1 , \584_b1 , \491_b1 );
not ( \491_b1 , w_1520 );
and ( \585_b0 , \584_b0 , w_1521 );
and ( w_1520 , w_1521 , \491_b0 );
or ( \586_b1 , \477_b1 , \483_b1 );
not ( \483_b1 , w_1522 );
and ( \586_b0 , \477_b0 , w_1523 );
and ( w_1522 , w_1523 , \483_b0 );
or ( \587_b1 , \585_b1 , w_1524 );
or ( \587_b0 , \585_b0 , \586_b0 );
not ( \586_b0 , w_1525 );
and ( w_1525 , w_1524 , \586_b1 );
or ( \588_b1 , \583_b1 , w_1526 );
xor ( \588_b0 , \583_b0 , w_1528 );
not ( w_1528 , w_1529 );
and ( w_1529 , w_1526 , w_1527 );
buf ( w_1526 , \587_b1 );
not ( w_1526 , w_1530 );
not ( w_1527 , w_1531 );
and ( w_1530 , w_1531 , \587_b0 );
buf ( \589_b1 , \481_b1 );
not ( \589_b1 , w_1532 );
not ( \589_b0 , w_1533 );
and ( w_1532 , w_1533 , \481_b0 );
buf ( \590_b1 , \401_b1 );
not ( \590_b1 , w_1534 );
not ( \590_b0 , w_1535 );
and ( w_1534 , w_1535 , \401_b0 );
or ( \591_b1 , \589_b1 , w_1536 );
or ( \591_b0 , \589_b0 , \590_b0 );
not ( \590_b0 , w_1537 );
and ( w_1537 , w_1536 , \590_b1 );
or ( \592_b1 , \a[3]_b1 , \b[9]_b1 );
xor ( \592_b0 , \a[3]_b0 , w_1538 );
not ( w_1538 , w_1539 );
and ( w_1539 , \b[9]_b1 , \b[9]_b0 );
or ( \593_b1 , \400_b1 , w_1541 );
not ( w_1541 , w_1542 );
and ( \593_b0 , \400_b0 , w_1543 );
and ( w_1542 ,  , w_1543 );
buf ( w_1541 , \592_b1 );
not ( w_1541 , w_1544 );
not (  , w_1545 );
and ( w_1544 , w_1545 , \592_b0 );
or ( \594_b1 , \591_b1 , w_1547 );
not ( w_1547 , w_1548 );
and ( \594_b0 , \591_b0 , w_1549 );
and ( w_1548 ,  , w_1549 );
buf ( w_1547 , \593_b1 );
not ( w_1547 , w_1550 );
not (  , w_1551 );
and ( w_1550 , w_1551 , \593_b0 );
buf ( \595_b1 , \518_b1 );
not ( \595_b1 , w_1552 );
not ( \595_b0 , w_1553 );
and ( w_1552 , w_1553 , \518_b0 );
buf ( \596_b1 , \195_b1 );
not ( \596_b1 , w_1554 );
not ( \596_b0 , w_1555 );
and ( w_1554 , w_1555 , \195_b0 );
or ( \597_b1 , \595_b1 , w_1556 );
or ( \597_b0 , \595_b0 , \596_b0 );
not ( \596_b0 , w_1557 );
and ( w_1557 , w_1556 , \596_b1 );
or ( \598_b1 , \a[7]_b1 , \b[5]_b1 );
xor ( \598_b0 , \a[7]_b0 , w_1558 );
not ( w_1558 , w_1559 );
and ( w_1559 , \b[5]_b1 , \b[5]_b0 );
or ( \599_b1 , \139_b1 , w_1561 );
not ( w_1561 , w_1562 );
and ( \599_b0 , \139_b0 , w_1563 );
and ( w_1562 ,  , w_1563 );
buf ( w_1561 , \598_b1 );
not ( w_1561 , w_1564 );
not (  , w_1565 );
and ( w_1564 , w_1565 , \598_b0 );
or ( \600_b1 , \597_b1 , w_1567 );
not ( w_1567 , w_1568 );
and ( \600_b0 , \597_b0 , w_1569 );
and ( w_1568 ,  , w_1569 );
buf ( w_1567 , \599_b1 );
not ( w_1567 , w_1570 );
not (  , w_1571 );
and ( w_1570 , w_1571 , \599_b0 );
or ( \601_b1 , \594_b1 , w_1572 );
xor ( \601_b0 , \594_b0 , w_1574 );
not ( w_1574 , w_1575 );
and ( w_1575 , w_1572 , w_1573 );
buf ( w_1572 , \600_b1 );
not ( w_1572 , w_1576 );
not ( w_1573 , w_1577 );
and ( w_1576 , w_1577 , \600_b0 );
buf ( \602_b1 , \489_b1 );
not ( \602_b1 , w_1578 );
not ( \602_b0 , w_1579 );
and ( w_1578 , w_1579 , \489_b0 );
buf ( \603_b1 , \486_b1 );
not ( \603_b1 , w_1580 );
not ( \603_b0 , w_1581 );
and ( w_1580 , w_1581 , \486_b0 );
or ( \604_b1 , \602_b1 , w_1582 );
or ( \604_b0 , \602_b0 , \603_b0 );
not ( \603_b0 , w_1583 );
and ( w_1583 , w_1582 , \603_b1 );
buf ( \605_b1 , \b[3]_b1 );
not ( \605_b1 , w_1584 );
not ( \605_b0 , w_1585 );
and ( w_1584 , w_1585 , \b[3]_b0 );
or ( \606_b1 , \605_b1 , w_1587 );
not ( w_1587 , w_1588 );
and ( \606_b0 , \605_b0 , w_1589 );
and ( w_1588 ,  , w_1589 );
buf ( w_1587 , \a[9]_b1 );
not ( w_1587 , w_1590 );
not (  , w_1591 );
and ( w_1590 , w_1591 , \a[9]_b0 );
buf ( \607_b1 , \606_b1 );
not ( \607_b1 , w_1592 );
not ( \607_b0 , w_1593 );
and ( w_1592 , w_1593 , \606_b0 );
buf ( \608_b1 , \a[9]_b1 );
not ( \608_b1 , w_1594 );
not ( \608_b0 , w_1595 );
and ( w_1594 , w_1595 , \a[9]_b0 );
or ( \609_b1 , \608_b1 , w_1597 );
not ( w_1597 , w_1598 );
and ( \609_b0 , \608_b0 , w_1599 );
and ( w_1598 ,  , w_1599 );
buf ( w_1597 , \b[3]_b1 );
not ( w_1597 , w_1600 );
not (  , w_1601 );
and ( w_1600 , w_1601 , \b[3]_b0 );
buf ( \610_b1 , \609_b1 );
not ( \610_b1 , w_1602 );
not ( \610_b0 , w_1603 );
and ( w_1602 , w_1603 , \609_b0 );
or ( \611_b1 , \607_b1 , w_1604 );
or ( \611_b0 , \607_b0 , \610_b0 );
not ( \610_b0 , w_1605 );
and ( w_1605 , w_1604 , \610_b1 );
or ( \612_b1 , \611_b1 , w_1607 );
not ( w_1607 , w_1608 );
and ( \612_b0 , \611_b0 , w_1609 );
and ( w_1608 ,  , w_1609 );
buf ( w_1607 , \147_b1 );
not ( w_1607 , w_1610 );
not (  , w_1611 );
and ( w_1610 , w_1611 , \147_b0 );
or ( \613_b1 , \604_b1 , w_1613 );
not ( w_1613 , w_1614 );
and ( \613_b0 , \604_b0 , w_1615 );
and ( w_1614 ,  , w_1615 );
buf ( w_1613 , \612_b1 );
not ( w_1613 , w_1616 );
not (  , w_1617 );
and ( w_1616 , w_1617 , \612_b0 );
buf ( \614_b1 , \613_b1 );
not ( \614_b1 , w_1618 );
not ( \614_b0 , w_1619 );
and ( w_1618 , w_1619 , \613_b0 );
buf ( \615_b1 , \475_b1 );
not ( \615_b1 , w_1620 );
not ( \615_b0 , w_1621 );
and ( w_1620 , w_1621 , \475_b0 );
buf ( \616_b1 , \374_b1 );
not ( \616_b1 , w_1622 );
not ( \616_b0 , w_1623 );
and ( w_1622 , w_1623 , \374_b0 );
or ( \617_b1 , \615_b1 , w_1624 );
or ( \617_b0 , \615_b0 , \616_b0 );
not ( \616_b0 , w_1625 );
and ( w_1625 , w_1624 , \616_b1 );
or ( \618_b1 , \a[5]_b1 , \b[7]_b1 );
xor ( \618_b0 , \a[5]_b0 , w_1626 );
not ( w_1626 , w_1627 );
and ( w_1627 , \b[7]_b1 , \b[7]_b0 );
or ( \619_b1 , \129_b1 , w_1629 );
not ( w_1629 , w_1630 );
and ( \619_b0 , \129_b0 , w_1631 );
and ( w_1630 ,  , w_1631 );
buf ( w_1629 , \618_b1 );
not ( w_1629 , w_1632 );
not (  , w_1633 );
and ( w_1632 , w_1633 , \618_b0 );
or ( \620_b1 , \617_b1 , w_1635 );
not ( w_1635 , w_1636 );
and ( \620_b0 , \617_b0 , w_1637 );
and ( w_1636 ,  , w_1637 );
buf ( w_1635 , \619_b1 );
not ( w_1635 , w_1638 );
not (  , w_1639 );
and ( w_1638 , w_1639 , \619_b0 );
buf ( \621_b1 , \620_b1 );
not ( \621_b1 , w_1640 );
not ( \621_b0 , w_1641 );
and ( w_1640 , w_1641 , \620_b0 );
buf ( \622_b1 , \621_b1 );
not ( \622_b1 , w_1642 );
not ( \622_b0 , w_1643 );
and ( w_1642 , w_1643 , \621_b0 );
or ( \623_b1 , \614_b1 , \622_b1 );
not ( \622_b1 , w_1644 );
and ( \623_b0 , \614_b0 , w_1645 );
and ( w_1644 , w_1645 , \622_b0 );
or ( \624_b1 , \613_b1 , \621_b1 );
not ( \621_b1 , w_1646 );
and ( \624_b0 , \613_b0 , w_1647 );
and ( w_1646 , w_1647 , \621_b0 );
or ( \625_b1 , \623_b1 , w_1649 );
not ( w_1649 , w_1650 );
and ( \625_b0 , \623_b0 , w_1651 );
and ( w_1650 ,  , w_1651 );
buf ( w_1649 , \624_b1 );
not ( w_1649 , w_1652 );
not (  , w_1653 );
and ( w_1652 , w_1653 , \624_b0 );
buf ( \626_b1 , \625_b1 );
not ( \626_b1 , w_1654 );
not ( \626_b0 , w_1655 );
and ( w_1654 , w_1655 , \625_b0 );
or ( \627_b1 , \601_b1 , \626_b1 );
xor ( \627_b0 , \601_b0 , w_1656 );
not ( w_1656 , w_1657 );
and ( w_1657 , \626_b1 , \626_b0 );
buf ( \628_b1 , \627_b1 );
not ( \628_b1 , w_1658 );
not ( \628_b0 , w_1659 );
and ( w_1658 , w_1659 , \627_b0 );
or ( \629_b1 , \588_b1 , \628_b1 );
not ( \628_b1 , w_1660 );
and ( \629_b0 , \588_b0 , w_1661 );
and ( w_1660 , w_1661 , \628_b0 );
buf ( \630_b1 , \588_b1 );
not ( \630_b1 , w_1662 );
not ( \630_b0 , w_1663 );
and ( w_1662 , w_1663 , \588_b0 );
or ( \631_b1 , \630_b1 , \627_b1 );
not ( \627_b1 , w_1664 );
and ( \631_b0 , \630_b0 , w_1665 );
and ( w_1664 , w_1665 , \627_b0 );
or ( \632_b1 , \629_b1 , w_1667 );
not ( w_1667 , w_1668 );
and ( \632_b0 , \629_b0 , w_1669 );
and ( w_1668 ,  , w_1669 );
buf ( w_1667 , \631_b1 );
not ( w_1667 , w_1670 );
not (  , w_1671 );
and ( w_1670 , w_1671 , \631_b0 );
or ( \633_b1 , \500_b1 , \504_b1 );
xor ( \633_b0 , \500_b0 , w_1672 );
not ( w_1672 , w_1673 );
and ( w_1673 , \504_b1 , \504_b0 );
or ( \634_b1 , \633_b1 , \521_b1 );
not ( \521_b1 , w_1674 );
and ( \634_b0 , \633_b0 , w_1675 );
and ( w_1674 , w_1675 , \521_b0 );
or ( \635_b1 , \500_b1 , \504_b1 );
not ( \504_b1 , w_1676 );
and ( \635_b0 , \500_b0 , w_1677 );
and ( w_1676 , w_1677 , \504_b0 );
or ( \636_b1 , \634_b1 , w_1678 );
or ( \636_b0 , \634_b0 , \635_b0 );
not ( \635_b0 , w_1679 );
and ( w_1679 , w_1678 , \635_b1 );
buf ( \637_b1 , \636_b1 );
not ( \637_b1 , w_1680 );
not ( \637_b0 , w_1681 );
and ( w_1680 , w_1681 , \636_b0 );
or ( \638_b1 , \632_b1 , \637_b1 );
not ( \637_b1 , w_1682 );
and ( \638_b0 , \632_b0 , w_1683 );
and ( w_1682 , w_1683 , \637_b0 );
buf ( \639_b1 , \632_b1 );
not ( \639_b1 , w_1684 );
not ( \639_b0 , w_1685 );
and ( w_1684 , w_1685 , \632_b0 );
or ( \640_b1 , \639_b1 , \636_b1 );
not ( \636_b1 , w_1686 );
and ( \640_b0 , \639_b0 , w_1687 );
and ( w_1686 , w_1687 , \636_b0 );
or ( \641_b1 , \638_b1 , w_1689 );
not ( w_1689 , w_1690 );
and ( \641_b0 , \638_b0 , w_1691 );
and ( w_1690 ,  , w_1691 );
buf ( w_1689 , \640_b1 );
not ( w_1689 , w_1692 );
not (  , w_1693 );
and ( w_1692 , w_1693 , \640_b0 );
or ( \642_b1 , \551_b1 , \641_b1 );
xor ( \642_b0 , \551_b0 , w_1694 );
not ( w_1694 , w_1695 );
and ( w_1695 , \641_b1 , \641_b0 );
buf ( \643_b1 , \642_b1 );
not ( \643_b1 , w_1696 );
not ( \643_b0 , w_1697 );
and ( w_1696 , w_1697 , \642_b0 );
or ( \644_b1 , \547_b1 , \643_b1 );
not ( \643_b1 , w_1698 );
and ( \644_b0 , \547_b0 , w_1699 );
and ( w_1698 , w_1699 , \643_b0 );
buf ( \645_b1 , \547_b1 );
not ( \645_b1 , w_1700 );
not ( \645_b0 , w_1701 );
and ( w_1700 , w_1701 , \547_b0 );
or ( \646_b1 , \645_b1 , \642_b1 );
not ( \642_b1 , w_1702 );
and ( \646_b0 , \645_b0 , w_1703 );
and ( w_1702 , w_1703 , \642_b0 );
or ( \647_b1 , \644_b1 , w_1705 );
not ( w_1705 , w_1706 );
and ( \647_b0 , \644_b0 , w_1707 );
and ( w_1706 ,  , w_1707 );
buf ( w_1705 , \646_b1 );
not ( w_1705 , w_1708 );
not (  , w_1709 );
and ( w_1708 , w_1709 , \646_b0 );
buf ( \648_b1 , \647_b1 );
buf ( \648_b0 , \647_b0 );
buf ( \649_b1 , \648_b1 );
buf ( \649_b0 , \648_b0 );
buf ( \650_b1 , \649_b1 );
not ( \650_b1 , w_1710 );
not ( \650_b0 , w_1711 );
and ( w_1710 , w_1711 , \649_b0 );
or ( \651_b1 , \99_b1 , w_1712 );
or ( \651_b0 , \99_b0 , \650_b0 );
not ( \650_b0 , w_1713 );
and ( w_1713 , w_1712 , \650_b1 );
buf ( \652_b1 , \535_b1 );
not ( \652_b1 , w_1714 );
not ( \652_b0 , w_1715 );
and ( w_1714 , w_1715 , \535_b0 );
or ( \653_b1 , \652_b1 , w_1717 );
not ( w_1717 , w_1718 );
and ( \653_b0 , \652_b0 , w_1719 );
and ( w_1718 ,  , w_1719 );
buf ( w_1717 , \461_b1 );
not ( w_1717 , w_1720 );
not (  , w_1721 );
and ( w_1720 , w_1721 , \461_b0 );
buf ( \654_b1 , \653_b1 );
not ( \654_b1 , w_1722 );
not ( \654_b0 , w_1723 );
and ( w_1722 , w_1723 , \653_b0 );
or ( \655_b1 , \654_b1 , w_1725 );
not ( w_1725 , w_1726 );
and ( \655_b0 , \654_b0 , w_1727 );
and ( w_1726 ,  , w_1727 );
buf ( w_1725 , \542_b1 );
not ( w_1725 , w_1728 );
not (  , w_1729 );
and ( w_1728 , w_1729 , \542_b0 );
buf ( \656_b1 , \655_b1 );
not ( \656_b1 , w_1730 );
not ( \656_b0 , w_1731 );
and ( w_1730 , w_1731 , \655_b0 );
buf ( \657_b1 , \470_b1 );
not ( \657_b1 , w_1732 );
not ( \657_b0 , w_1733 );
and ( w_1732 , w_1733 , \470_b0 );
buf ( \658_b1 , \347_b1 );
not ( \658_b1 , w_1734 );
not ( \658_b0 , w_1735 );
and ( w_1734 , w_1735 , \347_b0 );
or ( \659_b1 , \657_b1 , w_1736 );
or ( \659_b0 , \657_b0 , \658_b0 );
not ( \658_b0 , w_1737 );
and ( w_1737 , w_1736 , \658_b1 );
or ( \660_b1 , \539_b1 , w_1739 );
not ( w_1739 , w_1740 );
and ( \660_b0 , \539_b0 , w_1741 );
and ( w_1740 ,  , w_1741 );
buf ( w_1739 , \468_b1 );
not ( w_1739 , w_1742 );
not (  , w_1743 );
and ( w_1742 , w_1743 , \468_b0 );
buf ( \661_b1 , \660_b1 );
buf ( \661_b0 , \660_b0 );
or ( \662_b1 , \659_b1 , w_1745 );
not ( w_1745 , w_1746 );
and ( \662_b0 , \659_b0 , w_1747 );
and ( w_1746 ,  , w_1747 );
buf ( w_1745 , \661_b1 );
not ( w_1745 , w_1748 );
not (  , w_1749 );
and ( w_1748 , w_1749 , \661_b0 );
buf ( \663_b1 , \662_b1 );
not ( \663_b1 , w_1750 );
not ( \663_b0 , w_1751 );
and ( w_1750 , w_1751 , \662_b0 );
or ( \664_b1 , \656_b1 , w_1752 );
or ( \664_b0 , \656_b0 , \663_b0 );
not ( \663_b0 , w_1753 );
and ( w_1753 , w_1752 , \663_b1 );
or ( \665_b1 , \662_b1 , w_1754 );
or ( \665_b0 , \662_b0 , \655_b0 );
not ( \655_b0 , w_1755 );
and ( w_1755 , w_1754 , \655_b1 );
or ( \666_b1 , \664_b1 , w_1757 );
not ( w_1757 , w_1758 );
and ( \666_b0 , \664_b0 , w_1759 );
and ( w_1758 ,  , w_1759 );
buf ( w_1757 , \665_b1 );
not ( w_1757 , w_1760 );
not (  , w_1761 );
and ( w_1760 , w_1761 , \665_b0 );
buf ( \667_b1 , \666_b1 );
buf ( \667_b0 , \666_b0 );
or ( \668_b1 , \667_b1 , \b[15]_b1 );
not ( \b[15]_b1 , w_1762 );
and ( \668_b0 , \667_b0 , w_1763 );
and ( w_1762 , w_1763 , \b[15]_b0 );
or ( \669_b1 , \a[11]_b1 , w_1765 );
not ( w_1765 , w_1766 );
and ( \669_b0 , \a[11]_b0 , w_1767 );
and ( w_1766 ,  , w_1767 );
buf ( w_1765 , \d[11]_b1 );
not ( w_1765 , w_1768 );
not (  , w_1769 );
and ( w_1768 , w_1769 , \d[11]_b0 );
buf ( \670_b1 , \669_b1 );
not ( \670_b1 , w_1770 );
not ( \670_b0 , w_1771 );
and ( w_1770 , w_1771 , \669_b0 );
or ( \672_b1 , \a[10]_b1 , w_1773 );
not ( w_1773 , w_1774 );
and ( \672_b0 , \a[10]_b0 , w_1775 );
and ( w_1774 ,  , w_1775 );
buf ( w_1773 , \d[10]_b1 );
not ( w_1773 , w_1776 );
not (  , w_1777 );
and ( w_1776 , w_1777 , \d[10]_b0 );
or ( \673_b1 , \a[9]_b1 , w_1779 );
not ( w_1779 , w_1780 );
and ( \673_b0 , \a[9]_b0 , w_1781 );
and ( w_1780 ,  , w_1781 );
buf ( w_1779 , \d[9]_b1 );
not ( w_1779 , w_1782 );
not (  , w_1783 );
and ( w_1782 , w_1783 , \d[9]_b0 );
or ( \674_b1 , \a[3]_b1 , w_1785 );
not ( w_1785 , w_1786 );
and ( \674_b0 , \a[3]_b0 , w_1787 );
and ( w_1786 ,  , w_1787 );
buf ( w_1785 , \d[3]_b1 );
not ( w_1785 , w_1788 );
not (  , w_1789 );
and ( w_1788 , w_1789 , \d[3]_b0 );
or ( \679_b1 , \a[1]_b1 , \d[1]_b1 );
not ( \d[1]_b1 , w_1790 );
and ( \679_b0 , \a[1]_b0 , w_1791 );
and ( w_1790 , w_1791 , \d[1]_b0 );
or ( \680_b1 , \a[1]_b1 , w_1793 );
not ( w_1793 , w_1794 );
and ( \680_b0 , \a[1]_b0 , w_1795 );
and ( w_1794 ,  , w_1795 );
buf ( w_1793 , \d[1]_b1 );
not ( w_1793 , w_1796 );
not (  , w_1797 );
and ( w_1796 , w_1797 , \d[1]_b0 );
or ( \681_b1 , \a[0]_b1 , w_1799 );
not ( w_1799 , w_1800 );
and ( \681_b0 , \a[0]_b0 , w_1801 );
and ( w_1800 ,  , w_1801 );
buf ( w_1799 , \d[0]_b1 );
not ( w_1799 , w_1802 );
not (  , w_1803 );
and ( w_1802 , w_1803 , \d[0]_b0 );
or ( \683_b1 , \a[2]_b1 , w_1805 );
not ( w_1805 , w_1806 );
and ( \683_b0 , \a[2]_b0 , w_1807 );
and ( w_1806 ,  , w_1807 );
buf ( w_1805 , \d[2]_b1 );
not ( w_1805 , w_1808 );
not (  , w_1809 );
and ( w_1808 , w_1809 , \d[2]_b0 );
or ( \684_b1 , \a[0]_b1 , w_1811 );
not ( w_1811 , w_1812 );
and ( \684_b0 , \a[0]_b0 , w_1813 );
and ( w_1812 ,  , w_1813 );
buf ( w_1811 , \d[0]_b1 );
not ( w_1811 , w_1814 );
not (  , w_1815 );
and ( w_1814 , w_1815 , \d[0]_b0 );
or ( \686_b1 , \a[14]_b1 , w_1816 );
or ( \686_b0 , \a[14]_b0 , \d[14]_b0 );
not ( \d[14]_b0 , w_1817 );
and ( w_1817 , w_1816 , \d[14]_b1 );
buf ( \687_b1 , \d[12]_b1 );
not ( \687_b1 , w_1818 );
not ( \687_b0 , w_1819 );
and ( w_1818 , w_1819 , \d[12]_b0 );
buf ( \688_b1 , \a[12]_b1 );
not ( \688_b1 , w_1820 );
not ( \688_b0 , w_1821 );
and ( w_1820 , w_1821 , \a[12]_b0 );
or ( \689_b1 , \687_b1 , w_1823 );
not ( w_1823 , w_1824 );
and ( \689_b0 , \687_b0 , w_1825 );
and ( w_1824 ,  , w_1825 );
buf ( w_1823 , \688_b1 );
not ( w_1823 , w_1826 );
not (  , w_1827 );
and ( w_1826 , w_1827 , \688_b0 );
or ( \692_b1 , \691_b1 , w_1829 );
not ( w_1829 , w_1830 );
and ( \692_b0 , \691_b0 , w_1831 );
and ( w_1830 ,  , w_1831 );
buf ( w_1829 , \d[15]_b1 );
not ( w_1829 , w_1832 );
not (  , w_1833 );
and ( w_1832 , w_1833 , \d[15]_b0 );
buf ( \693_b1 , \692_b1 );
not ( \693_b1 , w_1834 );
not ( \693_b0 , w_1835 );
and ( w_1834 , w_1835 , \692_b0 );
or ( \694_b1 , \660_b1 , w_1837 );
not ( w_1837 , w_1838 );
and ( \694_b0 , \660_b0 , w_1839 );
and ( w_1838 ,  , w_1839 );
buf ( w_1837 , \470_b1 );
not ( w_1837 , w_1840 );
not (  , w_1841 );
and ( w_1840 , w_1841 , \470_b0 );
or ( \695_b1 , \347_b1 , w_1842 );
xor ( \695_b0 , \347_b0 , w_1844 );
not ( w_1844 , w_1845 );
and ( w_1845 , w_1842 , w_1843 );
buf ( w_1842 , \694_b1 );
not ( w_1842 , w_1846 );
not ( w_1843 , w_1847 );
and ( w_1846 , w_1847 , \694_b0 );
buf ( \696_b1 , \695_b1 );
not ( \696_b1 , w_1848 );
not ( \696_b0 , w_1849 );
and ( w_1848 , w_1849 , \695_b0 );
buf ( \697_b1 , \696_b1 );
not ( \697_b1 , w_1850 );
not ( \697_b0 , w_1851 );
and ( w_1850 , w_1851 , \696_b0 );
buf ( \698_b1 , \697_b1 );
not ( \698_b1 , w_1852 );
not ( \698_b0 , w_1853 );
and ( w_1852 , w_1853 , \697_b0 );
or ( \699_b1 , \693_b1 , w_1854 );
or ( \699_b0 , \693_b0 , \698_b0 );
not ( \698_b0 , w_1855 );
and ( w_1855 , w_1854 , \698_b1 );
buf ( \700_b1 , \262_b1 );
not ( \700_b1 , w_1856 );
not ( \700_b0 , w_1857 );
and ( w_1856 , w_1857 , \262_b0 );
buf ( \701_b1 , \266_b1 );
not ( \701_b1 , w_1858 );
not ( \701_b0 , w_1859 );
and ( w_1858 , w_1859 , \266_b0 );
or ( \702_b1 , \700_b1 , w_1860 );
or ( \702_b0 , \700_b0 , \701_b0 );
not ( \701_b0 , w_1861 );
and ( w_1861 , w_1860 , \701_b1 );
or ( \703_b1 , \702_b1 , w_1863 );
not ( w_1863 , w_1864 );
and ( \703_b0 , \702_b0 , w_1865 );
and ( w_1864 ,  , w_1865 );
buf ( w_1863 , \338_b1 );
not ( w_1863 , w_1866 );
not (  , w_1867 );
and ( w_1866 , w_1867 , \338_b0 );
buf ( \704_b1 , \335_b1 );
buf ( \704_b0 , \335_b0 );
or ( \705_b1 , \703_b1 , w_1868 );
xor ( \705_b0 , \703_b0 , w_1870 );
not ( w_1870 , w_1871 );
and ( w_1871 , w_1868 , w_1869 );
buf ( w_1868 , \704_b1 );
not ( w_1868 , w_1872 );
not ( w_1869 , w_1873 );
and ( w_1872 , w_1873 , \704_b0 );
buf ( \706_b1 , \705_b1 );
not ( \706_b1 , w_1874 );
not ( \706_b0 , w_1875 );
and ( w_1874 , w_1875 , \705_b0 );
buf ( \707_b1 , \706_b1 );
not ( \707_b1 , w_1876 );
not ( \707_b0 , w_1877 );
and ( w_1876 , w_1877 , \706_b0 );
buf ( \708_b1 , \b[15]_b1 );
not ( \708_b1 , w_1878 );
not ( \708_b0 , w_1879 );
and ( w_1878 , w_1879 , \b[15]_b0 );
buf ( \709_b1 , \d[15]_b1 );
not ( \709_b1 , w_1880 );
not ( \709_b0 , w_1881 );
and ( w_1880 , w_1881 , \d[15]_b0 );
or ( \710_b1 , \708_b1 , \709_b1 );
not ( \709_b1 , w_1882 );
and ( \710_b0 , \708_b0 , w_1883 );
and ( w_1882 , w_1883 , \709_b0 );
or ( \711_b1 , \b[15]_b1 , \d[15]_b1 );
not ( \d[15]_b1 , w_1884 );
and ( \711_b0 , \b[15]_b0 , w_1885 );
and ( w_1884 , w_1885 , \d[15]_b0 );
or ( \712_b1 , \710_b1 , w_1887 );
not ( w_1887 , w_1888 );
and ( \712_b0 , \710_b0 , w_1889 );
and ( w_1888 ,  , w_1889 );
buf ( w_1887 , \711_b1 );
not ( w_1887 , w_1890 );
not (  , w_1891 );
and ( w_1890 , w_1891 , \711_b0 );
buf ( \713_b1 , \712_b1 );
not ( \713_b1 , w_1892 );
not ( \713_b0 , w_1893 );
and ( w_1892 , w_1893 , \712_b0 );
or ( \714_b1 , \b[0]_b1 , w_1895 );
not ( w_1895 , w_1896 );
and ( \714_b0 , \b[0]_b0 , w_1897 );
and ( w_1896 ,  , w_1897 );
buf ( w_1895 , \d[0]_b1 );
not ( w_1895 , w_1898 );
not (  , w_1899 );
and ( w_1898 , w_1899 , \d[0]_b0 );
or ( \715_b1 , \b[1]_b1 , w_1901 );
not ( w_1901 , w_1902 );
and ( \715_b0 , \b[1]_b0 , w_1903 );
and ( w_1902 ,  , w_1903 );
buf ( w_1901 , \d[1]_b1 );
not ( w_1901 , w_1904 );
not (  , w_1905 );
and ( w_1904 , w_1905 , \d[1]_b0 );
or ( \716_b1 , \714_b1 , w_1907 );
not ( w_1907 , w_1908 );
and ( \716_b0 , \714_b0 , w_1909 );
and ( w_1908 ,  , w_1909 );
buf ( w_1907 , \715_b1 );
not ( w_1907 , w_1910 );
not (  , w_1911 );
and ( w_1910 , w_1911 , \715_b0 );
or ( \717_b1 , \b[1]_b1 , w_1912 );
or ( \717_b0 , \b[1]_b0 , \d[1]_b0 );
not ( \d[1]_b0 , w_1913 );
and ( w_1913 , w_1912 , \d[1]_b1 );
or ( \718_b1 , \b[2]_b1 , w_1915 );
not ( w_1915 , w_1916 );
and ( \718_b0 , \b[2]_b0 , w_1917 );
and ( w_1916 ,  , w_1917 );
buf ( w_1915 , \d[2]_b1 );
not ( w_1915 , w_1918 );
not (  , w_1919 );
and ( w_1918 , w_1919 , \d[2]_b0 );
buf ( \719_b1 , \718_b1 );
not ( \719_b1 , w_1920 );
not ( \719_b0 , w_1921 );
and ( w_1920 , w_1921 , \718_b0 );
or ( \721_b1 , \b[3]_b1 , w_1923 );
not ( w_1923 , w_1924 );
and ( \721_b0 , \b[3]_b0 , w_1925 );
and ( w_1924 ,  , w_1925 );
buf ( w_1923 , \d[3]_b1 );
not ( w_1923 , w_1926 );
not (  , w_1927 );
and ( w_1926 , w_1927 , \d[3]_b0 );
or ( \722_b1 , \b[2]_b1 , w_1929 );
not ( w_1929 , w_1930 );
and ( \722_b0 , \b[2]_b0 , w_1931 );
and ( w_1930 ,  , w_1931 );
buf ( w_1929 , \d[2]_b1 );
not ( w_1929 , w_1932 );
not (  , w_1933 );
and ( w_1932 , w_1933 , \d[2]_b0 );
buf ( \724_b1 , \723_b1 );
not ( \724_b1 , w_1934 );
not ( \724_b0 , w_1935 );
and ( w_1934 , w_1935 , \723_b0 );
or ( \725_b1 , \b[5]_b1 , w_1937 );
not ( w_1937 , w_1938 );
and ( \725_b0 , \b[5]_b0 , w_1939 );
and ( w_1938 ,  , w_1939 );
buf ( w_1937 , \d[5]_b1 );
not ( w_1937 , w_1940 );
not (  , w_1941 );
and ( w_1940 , w_1941 , \d[5]_b0 );
or ( \726_b1 , \b[4]_b1 , w_1943 );
not ( w_1943 , w_1944 );
and ( \726_b0 , \b[4]_b0 , w_1945 );
and ( w_1944 ,  , w_1945 );
buf ( w_1943 , \d[4]_b1 );
not ( w_1943 , w_1946 );
not (  , w_1947 );
and ( w_1946 , w_1947 , \d[4]_b0 );
or ( \727_b1 , \725_b1 , w_1949 );
not ( w_1949 , w_1950 );
and ( \727_b0 , \725_b0 , w_1951 );
and ( w_1950 ,  , w_1951 );
buf ( w_1949 , \726_b1 );
not ( w_1949 , w_1952 );
not (  , w_1953 );
and ( w_1952 , w_1953 , \726_b0 );
or ( \728_b1 , \b[6]_b1 , w_1955 );
not ( w_1955 , w_1956 );
and ( \728_b0 , \b[6]_b0 , w_1957 );
and ( w_1956 ,  , w_1957 );
buf ( w_1955 , \d[6]_b1 );
not ( w_1955 , w_1958 );
not (  , w_1959 );
and ( w_1958 , w_1959 , \d[6]_b0 );
or ( \729_b1 , \b[7]_b1 , w_1961 );
not ( w_1961 , w_1962 );
and ( \729_b0 , \b[7]_b0 , w_1963 );
and ( w_1962 ,  , w_1963 );
buf ( w_1961 , \d[7]_b1 );
not ( w_1961 , w_1964 );
not (  , w_1965 );
and ( w_1964 , w_1965 , \d[7]_b0 );
or ( \730_b1 , \728_b1 , w_1967 );
not ( w_1967 , w_1968 );
and ( \730_b0 , \728_b0 , w_1969 );
and ( w_1968 ,  , w_1969 );
buf ( w_1967 , \729_b1 );
not ( w_1967 , w_1970 );
not (  , w_1971 );
and ( w_1970 , w_1971 , \729_b0 );
or ( \731_b1 , \727_b1 , w_1973 );
not ( w_1973 , w_1974 );
and ( \731_b0 , \727_b0 , w_1975 );
and ( w_1974 ,  , w_1975 );
buf ( w_1973 , \730_b1 );
not ( w_1973 , w_1976 );
not (  , w_1977 );
and ( w_1976 , w_1977 , \730_b0 );
or ( \732_b1 , \b[3]_b1 , w_1979 );
not ( w_1979 , w_1980 );
and ( \732_b0 , \b[3]_b0 , w_1981 );
and ( w_1980 ,  , w_1981 );
buf ( w_1979 , \d[3]_b1 );
not ( w_1979 , w_1982 );
not (  , w_1983 );
and ( w_1982 , w_1983 , \d[3]_b0 );
or ( \733_b1 , \731_b1 , w_1985 );
not ( w_1985 , w_1986 );
and ( \733_b0 , \731_b0 , w_1987 );
and ( w_1986 ,  , w_1987 );
buf ( w_1985 , \732_b1 );
not ( w_1985 , w_1988 );
not (  , w_1989 );
and ( w_1988 , w_1989 , \732_b0 );
buf ( \734_b1 , \733_b1 );
not ( \734_b1 , w_1990 );
not ( \734_b0 , w_1991 );
and ( w_1990 , w_1991 , \733_b0 );
or ( \735_b1 , \724_b1 , w_1992 );
or ( \735_b0 , \724_b0 , \734_b0 );
not ( \734_b0 , w_1993 );
and ( w_1993 , w_1992 , \734_b1 );
or ( \736_b1 , \b[7]_b1 , w_1995 );
not ( w_1995 , w_1996 );
and ( \736_b0 , \b[7]_b0 , w_1997 );
and ( w_1996 ,  , w_1997 );
buf ( w_1995 , \d[7]_b1 );
not ( w_1995 , w_1998 );
not (  , w_1999 );
and ( w_1998 , w_1999 , \d[7]_b0 );
buf ( \737_b1 , \736_b1 );
not ( \737_b1 , w_2000 );
not ( \737_b0 , w_2001 );
and ( w_2000 , w_2001 , \736_b0 );
buf ( \738_b1 , \730_b1 );
not ( \738_b1 , w_2002 );
not ( \738_b0 , w_2003 );
and ( w_2002 , w_2003 , \730_b0 );
buf ( \739_b1 , \738_b1 );
not ( \739_b1 , w_2004 );
not ( \739_b0 , w_2005 );
and ( w_2004 , w_2005 , \738_b0 );
or ( \740_b1 , \737_b1 , w_2006 );
or ( \740_b0 , \737_b0 , \739_b0 );
not ( \739_b0 , w_2007 );
and ( w_2007 , w_2006 , \739_b1 );
or ( \741_b1 , \b[6]_b1 , w_2009 );
not ( w_2009 , w_2010 );
and ( \741_b0 , \b[6]_b0 , w_2011 );
and ( w_2010 ,  , w_2011 );
buf ( w_2009 , \d[6]_b1 );
not ( w_2009 , w_2012 );
not (  , w_2013 );
and ( w_2012 , w_2013 , \d[6]_b0 );
or ( \742_b1 , \b[5]_b1 , w_2015 );
not ( w_2015 , w_2016 );
and ( \742_b0 , \b[5]_b0 , w_2017 );
and ( w_2016 ,  , w_2017 );
buf ( w_2015 , \d[5]_b1 );
not ( w_2015 , w_2018 );
not (  , w_2019 );
and ( w_2018 , w_2019 , \d[5]_b0 );
or ( \743_b1 , \b[4]_b1 , w_2021 );
not ( w_2021 , w_2022 );
and ( \743_b0 , \b[4]_b0 , w_2023 );
and ( w_2022 ,  , w_2023 );
buf ( w_2021 , \d[4]_b1 );
not ( w_2021 , w_2024 );
not (  , w_2025 );
and ( w_2024 , w_2025 , \d[4]_b0 );
or ( \744_b1 , \725_b1 , w_2026 );
or ( \744_b0 , \725_b0 , \743_b0 );
not ( \743_b0 , w_2027 );
and ( w_2027 , w_2026 , \743_b1 );
or ( \746_b1 , \740_b1 , w_2029 );
not ( w_2029 , w_2030 );
and ( \746_b0 , \740_b0 , w_2031 );
and ( w_2030 ,  , w_2031 );
buf ( w_2029 , \745_b1 );
not ( w_2029 , w_2032 );
not (  , w_2033 );
and ( w_2032 , w_2033 , \745_b0 );
or ( \747_b1 , \735_b1 , w_2035 );
not ( w_2035 , w_2036 );
and ( \747_b0 , \735_b0 , w_2037 );
and ( w_2036 ,  , w_2037 );
buf ( w_2035 , \746_b1 );
not ( w_2035 , w_2038 );
not (  , w_2039 );
and ( w_2038 , w_2039 , \746_b0 );
or ( \748_b1 , \b[11]_b1 , w_2041 );
not ( w_2041 , w_2042 );
and ( \748_b0 , \b[11]_b0 , w_2043 );
and ( w_2042 ,  , w_2043 );
buf ( w_2041 , \d[11]_b1 );
not ( w_2041 , w_2044 );
not (  , w_2045 );
and ( w_2044 , w_2045 , \d[11]_b0 );
or ( \749_b1 , \b[10]_b1 , w_2047 );
not ( w_2047 , w_2048 );
and ( \749_b0 , \b[10]_b0 , w_2049 );
and ( w_2048 ,  , w_2049 );
buf ( w_2047 , \d[10]_b1 );
not ( w_2047 , w_2050 );
not (  , w_2051 );
and ( w_2050 , w_2051 , \d[10]_b0 );
or ( \750_b1 , \748_b1 , w_2053 );
not ( w_2053 , w_2054 );
and ( \750_b0 , \748_b0 , w_2055 );
and ( w_2054 ,  , w_2055 );
buf ( w_2053 , \749_b1 );
not ( w_2053 , w_2056 );
not (  , w_2057 );
and ( w_2056 , w_2057 , \749_b0 );
or ( \751_b1 , \b[9]_b1 , w_2059 );
not ( w_2059 , w_2060 );
and ( \751_b0 , \b[9]_b0 , w_2061 );
and ( w_2060 ,  , w_2061 );
buf ( w_2059 , \d[9]_b1 );
not ( w_2059 , w_2062 );
not (  , w_2063 );
and ( w_2062 , w_2063 , \d[9]_b0 );
or ( \752_b1 , \b[8]_b1 , w_2065 );
not ( w_2065 , w_2066 );
and ( \752_b0 , \b[8]_b0 , w_2067 );
and ( w_2066 ,  , w_2067 );
buf ( w_2065 , \d[8]_b1 );
not ( w_2065 , w_2068 );
not (  , w_2069 );
and ( w_2068 , w_2069 , \d[8]_b0 );
or ( \753_b1 , \751_b1 , w_2071 );
not ( w_2071 , w_2072 );
and ( \753_b0 , \751_b0 , w_2073 );
and ( w_2072 ,  , w_2073 );
buf ( w_2071 , \752_b1 );
not ( w_2071 , w_2074 );
not (  , w_2075 );
and ( w_2074 , w_2075 , \752_b0 );
or ( \754_b1 , \750_b1 , \753_b1 );
not ( \753_b1 , w_2076 );
and ( \754_b0 , \750_b0 , w_2077 );
and ( w_2076 , w_2077 , \753_b0 );
or ( \755_b1 , \b[14]_b1 , w_2079 );
not ( w_2079 , w_2080 );
and ( \755_b0 , \b[14]_b0 , w_2081 );
and ( w_2080 ,  , w_2081 );
buf ( w_2079 , \d[14]_b1 );
not ( w_2079 , w_2082 );
not (  , w_2083 );
and ( w_2082 , w_2083 , \d[14]_b0 );
buf ( \756_b1 , \755_b1 );
not ( \756_b1 , w_2084 );
not ( \756_b0 , w_2085 );
and ( w_2084 , w_2085 , \755_b0 );
or ( \757_b1 , \b[13]_b1 , w_2087 );
not ( w_2087 , w_2088 );
and ( \757_b0 , \b[13]_b0 , w_2089 );
and ( w_2088 ,  , w_2089 );
buf ( w_2087 , \d[13]_b1 );
not ( w_2087 , w_2090 );
not (  , w_2091 );
and ( w_2090 , w_2091 , \d[13]_b0 );
or ( \758_b1 , \b[12]_b1 , w_2093 );
not ( w_2093 , w_2094 );
and ( \758_b0 , \b[12]_b0 , w_2095 );
and ( w_2094 ,  , w_2095 );
buf ( w_2093 , \d[12]_b1 );
not ( w_2093 , w_2096 );
not (  , w_2097 );
and ( w_2096 , w_2097 , \d[12]_b0 );
or ( \759_b1 , \757_b1 , w_2099 );
not ( w_2099 , w_2100 );
and ( \759_b0 , \757_b0 , w_2101 );
and ( w_2100 ,  , w_2101 );
buf ( w_2099 , \758_b1 );
not ( w_2099 , w_2102 );
not (  , w_2103 );
and ( w_2102 , w_2103 , \758_b0 );
or ( \760_b1 , \756_b1 , w_2105 );
not ( w_2105 , w_2106 );
and ( \760_b0 , \756_b0 , w_2107 );
and ( w_2106 ,  , w_2107 );
buf ( w_2105 , \759_b1 );
not ( w_2105 , w_2108 );
not (  , w_2109 );
and ( w_2108 , w_2109 , \759_b0 );
buf ( \761_b1 , \760_b1 );
not ( \761_b1 , w_2110 );
not ( \761_b0 , w_2111 );
and ( w_2110 , w_2111 , \760_b0 );
or ( \763_b1 , \b[8]_b1 , w_2113 );
not ( w_2113 , w_2114 );
and ( \763_b0 , \b[8]_b0 , w_2115 );
and ( w_2114 ,  , w_2115 );
buf ( w_2113 , \d[8]_b1 );
not ( w_2113 , w_2116 );
not (  , w_2117 );
and ( w_2116 , w_2117 , \d[8]_b0 );
or ( \764_b1 , \751_b1 , w_2118 );
or ( \764_b0 , \751_b0 , \763_b0 );
not ( \763_b0 , w_2119 );
and ( w_2119 , w_2118 , \763_b1 );
or ( \765_b1 , \b[9]_b1 , w_2121 );
not ( w_2121 , w_2122 );
and ( \765_b0 , \b[9]_b0 , w_2123 );
and ( w_2122 ,  , w_2123 );
buf ( w_2121 , \d[9]_b1 );
not ( w_2121 , w_2124 );
not (  , w_2125 );
and ( w_2124 , w_2125 , \d[9]_b0 );
or ( \766_b1 , \764_b1 , w_2127 );
not ( w_2127 , w_2128 );
and ( \766_b0 , \764_b0 , w_2129 );
and ( w_2128 ,  , w_2129 );
buf ( w_2127 , \765_b1 );
not ( w_2127 , w_2130 );
not (  , w_2131 );
and ( w_2130 , w_2131 , \765_b0 );
buf ( \767_b1 , \766_b1 );
not ( \767_b1 , w_2132 );
not ( \767_b0 , w_2133 );
and ( w_2132 , w_2133 , \766_b0 );
buf ( \768_b1 , \750_b1 );
not ( \768_b1 , w_2134 );
not ( \768_b0 , w_2135 );
and ( w_2134 , w_2135 , \750_b0 );
or ( \769_b1 , \767_b1 , w_2136 );
or ( \769_b0 , \767_b0 , \768_b0 );
not ( \768_b0 , w_2137 );
and ( w_2137 , w_2136 , \768_b1 );
buf ( \770_b1 , \748_b1 );
not ( \770_b1 , w_2138 );
not ( \770_b0 , w_2139 );
and ( w_2138 , w_2139 , \748_b0 );
or ( \771_b1 , \b[10]_b1 , w_2141 );
not ( w_2141 , w_2142 );
and ( \771_b0 , \b[10]_b0 , w_2143 );
and ( w_2142 ,  , w_2143 );
buf ( w_2141 , \d[10]_b1 );
not ( w_2141 , w_2144 );
not (  , w_2145 );
and ( w_2144 , w_2145 , \d[10]_b0 );
buf ( \772_b1 , \771_b1 );
not ( \772_b1 , w_2146 );
not ( \772_b0 , w_2147 );
and ( w_2146 , w_2147 , \771_b0 );
or ( \773_b1 , \770_b1 , \772_b1 );
not ( \772_b1 , w_2148 );
and ( \773_b0 , \770_b0 , w_2149 );
and ( w_2148 , w_2149 , \772_b0 );
or ( \774_b1 , \b[11]_b1 , \d[11]_b1 );
not ( \d[11]_b1 , w_2150 );
and ( \774_b0 , \b[11]_b0 , w_2151 );
and ( w_2150 , w_2151 , \d[11]_b0 );
or ( \775_b1 , \773_b1 , w_2153 );
not ( w_2153 , w_2154 );
and ( \775_b0 , \773_b0 , w_2155 );
and ( w_2154 ,  , w_2155 );
buf ( w_2153 , \774_b1 );
not ( w_2153 , w_2156 );
not (  , w_2157 );
and ( w_2156 , w_2157 , \774_b0 );
or ( \776_b1 , \769_b1 , w_2159 );
not ( w_2159 , w_2160 );
and ( \776_b0 , \769_b0 , w_2161 );
and ( w_2160 ,  , w_2161 );
buf ( w_2159 , \775_b1 );
not ( w_2159 , w_2162 );
not (  , w_2163 );
and ( w_2162 , w_2163 , \775_b0 );
buf ( \777_b1 , \776_b1 );
not ( \777_b1 , w_2164 );
not ( \777_b0 , w_2165 );
and ( w_2164 , w_2165 , \776_b0 );
or ( \778_b1 , \777_b1 , w_2166 );
or ( \778_b0 , \777_b0 , \760_b0 );
not ( \760_b0 , w_2167 );
and ( w_2167 , w_2166 , \760_b1 );
or ( \779_b1 , \b[12]_b1 , w_2169 );
not ( w_2169 , w_2170 );
and ( \779_b0 , \b[12]_b0 , w_2171 );
and ( w_2170 ,  , w_2171 );
buf ( w_2169 , \d[12]_b1 );
not ( w_2169 , w_2172 );
not (  , w_2173 );
and ( w_2172 , w_2173 , \d[12]_b0 );
or ( \780_b1 , \757_b1 , w_2174 );
or ( \780_b0 , \757_b0 , \779_b0 );
not ( \779_b0 , w_2175 );
and ( w_2175 , w_2174 , \779_b1 );
or ( \781_b1 , \b[13]_b1 , w_2177 );
not ( w_2177 , w_2178 );
and ( \781_b0 , \b[13]_b0 , w_2179 );
and ( w_2178 ,  , w_2179 );
buf ( w_2177 , \d[13]_b1 );
not ( w_2177 , w_2180 );
not (  , w_2181 );
and ( w_2180 , w_2181 , \d[13]_b0 );
or ( \782_b1 , \780_b1 , w_2183 );
not ( w_2183 , w_2184 );
and ( \782_b0 , \780_b0 , w_2185 );
and ( w_2184 ,  , w_2185 );
buf ( w_2183 , \781_b1 );
not ( w_2183 , w_2186 );
not (  , w_2187 );
and ( w_2186 , w_2187 , \781_b0 );
buf ( \783_b1 , \782_b1 );
not ( \783_b1 , w_2188 );
not ( \783_b0 , w_2189 );
and ( w_2188 , w_2189 , \782_b0 );
or ( \784_b1 , \755_b1 , w_2190 );
or ( \784_b0 , \755_b0 , \783_b0 );
not ( \783_b0 , w_2191 );
and ( w_2191 , w_2190 , \783_b1 );
or ( \785_b1 , \b[14]_b1 , w_2193 );
not ( w_2193 , w_2194 );
and ( \785_b0 , \b[14]_b0 , w_2195 );
and ( w_2194 ,  , w_2195 );
buf ( w_2193 , \d[14]_b1 );
not ( w_2193 , w_2196 );
not (  , w_2197 );
and ( w_2196 , w_2197 , \d[14]_b0 );
or ( \787_b1 , \762_b1 , w_2199 );
not ( w_2199 , w_2200 );
and ( \787_b0 , \762_b0 , w_2201 );
and ( w_2200 ,  , w_2201 );
buf ( w_2199 , \786_b1 );
not ( w_2199 , w_2202 );
not (  , w_2203 );
and ( w_2202 , w_2203 , \786_b0 );
buf ( \788_b1 , \787_b1 );
not ( \788_b1 , w_2204 );
not ( \788_b0 , w_2205 );
and ( w_2204 , w_2205 , \787_b0 );
or ( \789_b1 , \713_b1 , w_2206 );
or ( \789_b0 , \713_b0 , \788_b0 );
not ( \788_b0 , w_2207 );
and ( w_2207 , w_2206 , \788_b1 );
or ( \790_b1 , \787_b1 , w_2208 );
or ( \790_b0 , \787_b0 , \712_b0 );
not ( \712_b0 , w_2209 );
and ( w_2209 , w_2208 , \712_b1 );
or ( \791_b1 , \789_b1 , w_2211 );
not ( w_2211 , w_2212 );
and ( \791_b0 , \789_b0 , w_2213 );
and ( w_2212 ,  , w_2213 );
buf ( w_2211 , \790_b1 );
not ( w_2211 , w_2214 );
not (  , w_2215 );
and ( w_2214 , w_2215 , \790_b0 );
or ( \792_b1 , \707_b1 , \791_b1 );
not ( \791_b1 , w_2216 );
and ( \792_b0 , \707_b0 , w_2217 );
and ( w_2216 , w_2217 , \791_b0 );
buf ( \793_b1 , \a[15]_b1 );
not ( \793_b1 , w_2218 );
not ( \793_b0 , w_2219 );
and ( w_2218 , w_2219 , \a[15]_b0 );
buf ( \794_b1 , \c[15]_b1 );
not ( \794_b1 , w_2220 );
not ( \794_b0 , w_2221 );
and ( w_2220 , w_2221 , \c[15]_b0 );
or ( \795_b1 , \793_b1 , \794_b1 );
not ( \794_b1 , w_2222 );
and ( \795_b0 , \793_b0 , w_2223 );
and ( w_2222 , w_2223 , \794_b0 );
or ( \796_b1 , \a[15]_b1 , \c[15]_b1 );
not ( \c[15]_b1 , w_2224 );
and ( \796_b0 , \a[15]_b0 , w_2225 );
and ( w_2224 , w_2225 , \c[15]_b0 );
or ( \797_b1 , \795_b1 , w_2227 );
not ( w_2227 , w_2228 );
and ( \797_b0 , \795_b0 , w_2229 );
and ( w_2228 ,  , w_2229 );
buf ( w_2227 , \796_b1 );
not ( w_2227 , w_2230 );
not (  , w_2231 );
and ( w_2230 , w_2231 , \796_b0 );
buf ( \798_b1 , \797_b1 );
not ( \798_b1 , w_2232 );
not ( \798_b0 , w_2233 );
and ( w_2232 , w_2233 , \797_b0 );
or ( \799_b1 , \a[0]_b1 , w_2235 );
not ( w_2235 , w_2236 );
and ( \799_b0 , \a[0]_b0 , w_2237 );
and ( w_2236 ,  , w_2237 );
buf ( w_2235 , \c[0]_b1 );
not ( w_2235 , w_2238 );
not (  , w_2239 );
and ( w_2238 , w_2239 , \c[0]_b0 );
or ( \800_b1 , \a[1]_b1 , w_2241 );
not ( w_2241 , w_2242 );
and ( \800_b0 , \a[1]_b0 , w_2243 );
and ( w_2242 ,  , w_2243 );
buf ( w_2241 , \c[1]_b1 );
not ( w_2241 , w_2244 );
not (  , w_2245 );
and ( w_2244 , w_2245 , \c[1]_b0 );
or ( \801_b1 , \799_b1 , w_2247 );
not ( w_2247 , w_2248 );
and ( \801_b0 , \799_b0 , w_2249 );
and ( w_2248 ,  , w_2249 );
buf ( w_2247 , \800_b1 );
not ( w_2247 , w_2250 );
not (  , w_2251 );
and ( w_2250 , w_2251 , \800_b0 );
or ( \802_b1 , \a[1]_b1 , w_2252 );
or ( \802_b0 , \a[1]_b0 , \c[1]_b0 );
not ( \c[1]_b0 , w_2253 );
and ( w_2253 , w_2252 , \c[1]_b1 );
or ( \803_b1 , \a[2]_b1 , w_2255 );
not ( w_2255 , w_2256 );
and ( \803_b0 , \a[2]_b0 , w_2257 );
and ( w_2256 ,  , w_2257 );
buf ( w_2255 , \c[2]_b1 );
not ( w_2255 , w_2258 );
not (  , w_2259 );
and ( w_2258 , w_2259 , \c[2]_b0 );
buf ( \804_b1 , \803_b1 );
not ( \804_b1 , w_2260 );
not ( \804_b0 , w_2261 );
and ( w_2260 , w_2261 , \803_b0 );
or ( \806_b1 , \a[3]_b1 , w_2263 );
not ( w_2263 , w_2264 );
and ( \806_b0 , \a[3]_b0 , w_2265 );
and ( w_2264 ,  , w_2265 );
buf ( w_2263 , \c[3]_b1 );
not ( w_2263 , w_2266 );
not (  , w_2267 );
and ( w_2266 , w_2267 , \c[3]_b0 );
or ( \807_b1 , \a[2]_b1 , w_2269 );
not ( w_2269 , w_2270 );
and ( \807_b0 , \a[2]_b0 , w_2271 );
and ( w_2270 ,  , w_2271 );
buf ( w_2269 , \c[2]_b1 );
not ( w_2269 , w_2272 );
not (  , w_2273 );
and ( w_2272 , w_2273 , \c[2]_b0 );
buf ( \809_b1 , \808_b1 );
not ( \809_b1 , w_2274 );
not ( \809_b0 , w_2275 );
and ( w_2274 , w_2275 , \808_b0 );
or ( \810_b1 , \a[5]_b1 , w_2277 );
not ( w_2277 , w_2278 );
and ( \810_b0 , \a[5]_b0 , w_2279 );
and ( w_2278 ,  , w_2279 );
buf ( w_2277 , \c[5]_b1 );
not ( w_2277 , w_2280 );
not (  , w_2281 );
and ( w_2280 , w_2281 , \c[5]_b0 );
or ( \811_b1 , \a[4]_b1 , w_2283 );
not ( w_2283 , w_2284 );
and ( \811_b0 , \a[4]_b0 , w_2285 );
and ( w_2284 ,  , w_2285 );
buf ( w_2283 , \c[4]_b1 );
not ( w_2283 , w_2286 );
not (  , w_2287 );
and ( w_2286 , w_2287 , \c[4]_b0 );
or ( \812_b1 , \810_b1 , w_2289 );
not ( w_2289 , w_2290 );
and ( \812_b0 , \810_b0 , w_2291 );
and ( w_2290 ,  , w_2291 );
buf ( w_2289 , \811_b1 );
not ( w_2289 , w_2292 );
not (  , w_2293 );
and ( w_2292 , w_2293 , \811_b0 );
or ( \813_b1 , \a[6]_b1 , w_2295 );
not ( w_2295 , w_2296 );
and ( \813_b0 , \a[6]_b0 , w_2297 );
and ( w_2296 ,  , w_2297 );
buf ( w_2295 , \c[6]_b1 );
not ( w_2295 , w_2298 );
not (  , w_2299 );
and ( w_2298 , w_2299 , \c[6]_b0 );
or ( \814_b1 , \a[7]_b1 , w_2301 );
not ( w_2301 , w_2302 );
and ( \814_b0 , \a[7]_b0 , w_2303 );
and ( w_2302 ,  , w_2303 );
buf ( w_2301 , \c[7]_b1 );
not ( w_2301 , w_2304 );
not (  , w_2305 );
and ( w_2304 , w_2305 , \c[7]_b0 );
or ( \815_b1 , \813_b1 , w_2307 );
not ( w_2307 , w_2308 );
and ( \815_b0 , \813_b0 , w_2309 );
and ( w_2308 ,  , w_2309 );
buf ( w_2307 , \814_b1 );
not ( w_2307 , w_2310 );
not (  , w_2311 );
and ( w_2310 , w_2311 , \814_b0 );
or ( \816_b1 , \812_b1 , w_2313 );
not ( w_2313 , w_2314 );
and ( \816_b0 , \812_b0 , w_2315 );
and ( w_2314 ,  , w_2315 );
buf ( w_2313 , \815_b1 );
not ( w_2313 , w_2316 );
not (  , w_2317 );
and ( w_2316 , w_2317 , \815_b0 );
or ( \817_b1 , \a[3]_b1 , w_2319 );
not ( w_2319 , w_2320 );
and ( \817_b0 , \a[3]_b0 , w_2321 );
and ( w_2320 ,  , w_2321 );
buf ( w_2319 , \c[3]_b1 );
not ( w_2319 , w_2322 );
not (  , w_2323 );
and ( w_2322 , w_2323 , \c[3]_b0 );
or ( \818_b1 , \816_b1 , w_2325 );
not ( w_2325 , w_2326 );
and ( \818_b0 , \816_b0 , w_2327 );
and ( w_2326 ,  , w_2327 );
buf ( w_2325 , \817_b1 );
not ( w_2325 , w_2328 );
not (  , w_2329 );
and ( w_2328 , w_2329 , \817_b0 );
buf ( \819_b1 , \818_b1 );
not ( \819_b1 , w_2330 );
not ( \819_b0 , w_2331 );
and ( w_2330 , w_2331 , \818_b0 );
or ( \820_b1 , \809_b1 , w_2332 );
or ( \820_b0 , \809_b0 , \819_b0 );
not ( \819_b0 , w_2333 );
and ( w_2333 , w_2332 , \819_b1 );
or ( \821_b1 , \a[7]_b1 , w_2335 );
not ( w_2335 , w_2336 );
and ( \821_b0 , \a[7]_b0 , w_2337 );
and ( w_2336 ,  , w_2337 );
buf ( w_2335 , \c[7]_b1 );
not ( w_2335 , w_2338 );
not (  , w_2339 );
and ( w_2338 , w_2339 , \c[7]_b0 );
buf ( \822_b1 , \821_b1 );
not ( \822_b1 , w_2340 );
not ( \822_b0 , w_2341 );
and ( w_2340 , w_2341 , \821_b0 );
buf ( \823_b1 , \815_b1 );
not ( \823_b1 , w_2342 );
not ( \823_b0 , w_2343 );
and ( w_2342 , w_2343 , \815_b0 );
buf ( \824_b1 , \823_b1 );
not ( \824_b1 , w_2344 );
not ( \824_b0 , w_2345 );
and ( w_2344 , w_2345 , \823_b0 );
or ( \825_b1 , \822_b1 , w_2346 );
or ( \825_b0 , \822_b0 , \824_b0 );
not ( \824_b0 , w_2347 );
and ( w_2347 , w_2346 , \824_b1 );
or ( \826_b1 , \a[6]_b1 , w_2349 );
not ( w_2349 , w_2350 );
and ( \826_b0 , \a[6]_b0 , w_2351 );
and ( w_2350 ,  , w_2351 );
buf ( w_2349 , \c[6]_b1 );
not ( w_2349 , w_2352 );
not (  , w_2353 );
and ( w_2352 , w_2353 , \c[6]_b0 );
or ( \827_b1 , \a[5]_b1 , w_2355 );
not ( w_2355 , w_2356 );
and ( \827_b0 , \a[5]_b0 , w_2357 );
and ( w_2356 ,  , w_2357 );
buf ( w_2355 , \c[5]_b1 );
not ( w_2355 , w_2358 );
not (  , w_2359 );
and ( w_2358 , w_2359 , \c[5]_b0 );
or ( \828_b1 , \a[4]_b1 , w_2361 );
not ( w_2361 , w_2362 );
and ( \828_b0 , \a[4]_b0 , w_2363 );
and ( w_2362 ,  , w_2363 );
buf ( w_2361 , \c[4]_b1 );
not ( w_2361 , w_2364 );
not (  , w_2365 );
and ( w_2364 , w_2365 , \c[4]_b0 );
or ( \829_b1 , \810_b1 , w_2366 );
or ( \829_b0 , \810_b0 , \828_b0 );
not ( \828_b0 , w_2367 );
and ( w_2367 , w_2366 , \828_b1 );
or ( \831_b1 , \825_b1 , w_2369 );
not ( w_2369 , w_2370 );
and ( \831_b0 , \825_b0 , w_2371 );
and ( w_2370 ,  , w_2371 );
buf ( w_2369 , \830_b1 );
not ( w_2369 , w_2372 );
not (  , w_2373 );
and ( w_2372 , w_2373 , \830_b0 );
or ( \832_b1 , \820_b1 , w_2375 );
not ( w_2375 , w_2376 );
and ( \832_b0 , \820_b0 , w_2377 );
and ( w_2376 ,  , w_2377 );
buf ( w_2375 , \831_b1 );
not ( w_2375 , w_2378 );
not (  , w_2379 );
and ( w_2378 , w_2379 , \831_b0 );
or ( \833_b1 , \a[11]_b1 , w_2381 );
not ( w_2381 , w_2382 );
and ( \833_b0 , \a[11]_b0 , w_2383 );
and ( w_2382 ,  , w_2383 );
buf ( w_2381 , \c[11]_b1 );
not ( w_2381 , w_2384 );
not (  , w_2385 );
and ( w_2384 , w_2385 , \c[11]_b0 );
or ( \834_b1 , \a[10]_b1 , w_2387 );
not ( w_2387 , w_2388 );
and ( \834_b0 , \a[10]_b0 , w_2389 );
and ( w_2388 ,  , w_2389 );
buf ( w_2387 , \c[10]_b1 );
not ( w_2387 , w_2390 );
not (  , w_2391 );
and ( w_2390 , w_2391 , \c[10]_b0 );
or ( \835_b1 , \833_b1 , w_2393 );
not ( w_2393 , w_2394 );
and ( \835_b0 , \833_b0 , w_2395 );
and ( w_2394 ,  , w_2395 );
buf ( w_2393 , \834_b1 );
not ( w_2393 , w_2396 );
not (  , w_2397 );
and ( w_2396 , w_2397 , \834_b0 );
or ( \836_b1 , \a[9]_b1 , w_2399 );
not ( w_2399 , w_2400 );
and ( \836_b0 , \a[9]_b0 , w_2401 );
and ( w_2400 ,  , w_2401 );
buf ( w_2399 , \c[9]_b1 );
not ( w_2399 , w_2402 );
not (  , w_2403 );
and ( w_2402 , w_2403 , \c[9]_b0 );
or ( \837_b1 , \a[8]_b1 , w_2405 );
not ( w_2405 , w_2406 );
and ( \837_b0 , \a[8]_b0 , w_2407 );
and ( w_2406 ,  , w_2407 );
buf ( w_2405 , \c[8]_b1 );
not ( w_2405 , w_2408 );
not (  , w_2409 );
and ( w_2408 , w_2409 , \c[8]_b0 );
or ( \838_b1 , \836_b1 , w_2411 );
not ( w_2411 , w_2412 );
and ( \838_b0 , \836_b0 , w_2413 );
and ( w_2412 ,  , w_2413 );
buf ( w_2411 , \837_b1 );
not ( w_2411 , w_2414 );
not (  , w_2415 );
and ( w_2414 , w_2415 , \837_b0 );
or ( \839_b1 , \835_b1 , \838_b1 );
not ( \838_b1 , w_2416 );
and ( \839_b0 , \835_b0 , w_2417 );
and ( w_2416 , w_2417 , \838_b0 );
or ( \840_b1 , \a[14]_b1 , w_2419 );
not ( w_2419 , w_2420 );
and ( \840_b0 , \a[14]_b0 , w_2421 );
and ( w_2420 ,  , w_2421 );
buf ( w_2419 , \c[14]_b1 );
not ( w_2419 , w_2422 );
not (  , w_2423 );
and ( w_2422 , w_2423 , \c[14]_b0 );
buf ( \841_b1 , \840_b1 );
not ( \841_b1 , w_2424 );
not ( \841_b0 , w_2425 );
and ( w_2424 , w_2425 , \840_b0 );
or ( \842_b1 , \a[13]_b1 , w_2427 );
not ( w_2427 , w_2428 );
and ( \842_b0 , \a[13]_b0 , w_2429 );
and ( w_2428 ,  , w_2429 );
buf ( w_2427 , \c[13]_b1 );
not ( w_2427 , w_2430 );
not (  , w_2431 );
and ( w_2430 , w_2431 , \c[13]_b0 );
or ( \843_b1 , \a[12]_b1 , w_2433 );
not ( w_2433 , w_2434 );
and ( \843_b0 , \a[12]_b0 , w_2435 );
and ( w_2434 ,  , w_2435 );
buf ( w_2433 , \c[12]_b1 );
not ( w_2433 , w_2436 );
not (  , w_2437 );
and ( w_2436 , w_2437 , \c[12]_b0 );
or ( \844_b1 , \842_b1 , w_2439 );
not ( w_2439 , w_2440 );
and ( \844_b0 , \842_b0 , w_2441 );
and ( w_2440 ,  , w_2441 );
buf ( w_2439 , \843_b1 );
not ( w_2439 , w_2442 );
not (  , w_2443 );
and ( w_2442 , w_2443 , \843_b0 );
or ( \845_b1 , \841_b1 , w_2445 );
not ( w_2445 , w_2446 );
and ( \845_b0 , \841_b0 , w_2447 );
and ( w_2446 ,  , w_2447 );
buf ( w_2445 , \844_b1 );
not ( w_2445 , w_2448 );
not (  , w_2449 );
and ( w_2448 , w_2449 , \844_b0 );
buf ( \846_b1 , \845_b1 );
not ( \846_b1 , w_2450 );
not ( \846_b0 , w_2451 );
and ( w_2450 , w_2451 , \845_b0 );
or ( \848_b1 , \a[8]_b1 , w_2453 );
not ( w_2453 , w_2454 );
and ( \848_b0 , \a[8]_b0 , w_2455 );
and ( w_2454 ,  , w_2455 );
buf ( w_2453 , \c[8]_b1 );
not ( w_2453 , w_2456 );
not (  , w_2457 );
and ( w_2456 , w_2457 , \c[8]_b0 );
or ( \849_b1 , \836_b1 , w_2458 );
or ( \849_b0 , \836_b0 , \848_b0 );
not ( \848_b0 , w_2459 );
and ( w_2459 , w_2458 , \848_b1 );
or ( \850_b1 , \a[9]_b1 , w_2461 );
not ( w_2461 , w_2462 );
and ( \850_b0 , \a[9]_b0 , w_2463 );
and ( w_2462 ,  , w_2463 );
buf ( w_2461 , \c[9]_b1 );
not ( w_2461 , w_2464 );
not (  , w_2465 );
and ( w_2464 , w_2465 , \c[9]_b0 );
or ( \851_b1 , \849_b1 , w_2467 );
not ( w_2467 , w_2468 );
and ( \851_b0 , \849_b0 , w_2469 );
and ( w_2468 ,  , w_2469 );
buf ( w_2467 , \850_b1 );
not ( w_2467 , w_2470 );
not (  , w_2471 );
and ( w_2470 , w_2471 , \850_b0 );
buf ( \852_b1 , \851_b1 );
not ( \852_b1 , w_2472 );
not ( \852_b0 , w_2473 );
and ( w_2472 , w_2473 , \851_b0 );
buf ( \853_b1 , \835_b1 );
not ( \853_b1 , w_2474 );
not ( \853_b0 , w_2475 );
and ( w_2474 , w_2475 , \835_b0 );
or ( \854_b1 , \852_b1 , w_2476 );
or ( \854_b0 , \852_b0 , \853_b0 );
not ( \853_b0 , w_2477 );
and ( w_2477 , w_2476 , \853_b1 );
buf ( \855_b1 , \833_b1 );
not ( \855_b1 , w_2478 );
not ( \855_b0 , w_2479 );
and ( w_2478 , w_2479 , \833_b0 );
or ( \856_b1 , \a[10]_b1 , w_2481 );
not ( w_2481 , w_2482 );
and ( \856_b0 , \a[10]_b0 , w_2483 );
and ( w_2482 ,  , w_2483 );
buf ( w_2481 , \c[10]_b1 );
not ( w_2481 , w_2484 );
not (  , w_2485 );
and ( w_2484 , w_2485 , \c[10]_b0 );
buf ( \857_b1 , \856_b1 );
not ( \857_b1 , w_2486 );
not ( \857_b0 , w_2487 );
and ( w_2486 , w_2487 , \856_b0 );
or ( \858_b1 , \855_b1 , \857_b1 );
not ( \857_b1 , w_2488 );
and ( \858_b0 , \855_b0 , w_2489 );
and ( w_2488 , w_2489 , \857_b0 );
or ( \859_b1 , \a[11]_b1 , \c[11]_b1 );
not ( \c[11]_b1 , w_2490 );
and ( \859_b0 , \a[11]_b0 , w_2491 );
and ( w_2490 , w_2491 , \c[11]_b0 );
or ( \860_b1 , \858_b1 , w_2493 );
not ( w_2493 , w_2494 );
and ( \860_b0 , \858_b0 , w_2495 );
and ( w_2494 ,  , w_2495 );
buf ( w_2493 , \859_b1 );
not ( w_2493 , w_2496 );
not (  , w_2497 );
and ( w_2496 , w_2497 , \859_b0 );
or ( \861_b1 , \854_b1 , w_2499 );
not ( w_2499 , w_2500 );
and ( \861_b0 , \854_b0 , w_2501 );
and ( w_2500 ,  , w_2501 );
buf ( w_2499 , \860_b1 );
not ( w_2499 , w_2502 );
not (  , w_2503 );
and ( w_2502 , w_2503 , \860_b0 );
buf ( \862_b1 , \861_b1 );
not ( \862_b1 , w_2504 );
not ( \862_b0 , w_2505 );
and ( w_2504 , w_2505 , \861_b0 );
or ( \863_b1 , \862_b1 , w_2506 );
or ( \863_b0 , \862_b0 , \845_b0 );
not ( \845_b0 , w_2507 );
and ( w_2507 , w_2506 , \845_b1 );
or ( \864_b1 , \a[12]_b1 , w_2509 );
not ( w_2509 , w_2510 );
and ( \864_b0 , \a[12]_b0 , w_2511 );
and ( w_2510 ,  , w_2511 );
buf ( w_2509 , \c[12]_b1 );
not ( w_2509 , w_2512 );
not (  , w_2513 );
and ( w_2512 , w_2513 , \c[12]_b0 );
or ( \865_b1 , \842_b1 , w_2514 );
or ( \865_b0 , \842_b0 , \864_b0 );
not ( \864_b0 , w_2515 );
and ( w_2515 , w_2514 , \864_b1 );
or ( \866_b1 , \a[13]_b1 , w_2517 );
not ( w_2517 , w_2518 );
and ( \866_b0 , \a[13]_b0 , w_2519 );
and ( w_2518 ,  , w_2519 );
buf ( w_2517 , \c[13]_b1 );
not ( w_2517 , w_2520 );
not (  , w_2521 );
and ( w_2520 , w_2521 , \c[13]_b0 );
or ( \867_b1 , \865_b1 , w_2523 );
not ( w_2523 , w_2524 );
and ( \867_b0 , \865_b0 , w_2525 );
and ( w_2524 ,  , w_2525 );
buf ( w_2523 , \866_b1 );
not ( w_2523 , w_2526 );
not (  , w_2527 );
and ( w_2526 , w_2527 , \866_b0 );
buf ( \868_b1 , \867_b1 );
not ( \868_b1 , w_2528 );
not ( \868_b0 , w_2529 );
and ( w_2528 , w_2529 , \867_b0 );
or ( \869_b1 , \840_b1 , w_2530 );
or ( \869_b0 , \840_b0 , \868_b0 );
not ( \868_b0 , w_2531 );
and ( w_2531 , w_2530 , \868_b1 );
or ( \870_b1 , \a[14]_b1 , w_2533 );
not ( w_2533 , w_2534 );
and ( \870_b0 , \a[14]_b0 , w_2535 );
and ( w_2534 ,  , w_2535 );
buf ( w_2533 , \c[14]_b1 );
not ( w_2533 , w_2536 );
not (  , w_2537 );
and ( w_2536 , w_2537 , \c[14]_b0 );
or ( \872_b1 , \847_b1 , w_2539 );
not ( w_2539 , w_2540 );
and ( \872_b0 , \847_b0 , w_2541 );
and ( w_2540 ,  , w_2541 );
buf ( w_2539 , \871_b1 );
not ( w_2539 , w_2542 );
not (  , w_2543 );
and ( w_2542 , w_2543 , \871_b0 );
buf ( \873_b1 , \872_b1 );
not ( \873_b1 , w_2544 );
not ( \873_b0 , w_2545 );
and ( w_2544 , w_2545 , \872_b0 );
or ( \874_b1 , \798_b1 , w_2546 );
or ( \874_b0 , \798_b0 , \873_b0 );
not ( \873_b0 , w_2547 );
and ( w_2547 , w_2546 , \873_b1 );
or ( \875_b1 , \872_b1 , w_2548 );
or ( \875_b0 , \872_b0 , \797_b0 );
not ( \797_b0 , w_2549 );
and ( w_2549 , w_2548 , \797_b1 );
or ( \876_b1 , \874_b1 , w_2551 );
not ( w_2551 , w_2552 );
and ( \876_b0 , \874_b0 , w_2553 );
and ( w_2552 ,  , w_2553 );
buf ( w_2551 , \875_b1 );
not ( w_2551 , w_2554 );
not (  , w_2555 );
and ( w_2554 , w_2555 , \875_b0 );
buf ( \877_b1 , \876_b1 );
not ( \877_b1 , w_2556 );
not ( \877_b0 , w_2557 );
and ( w_2556 , w_2557 , \876_b0 );
or ( \878_b1 , \334_b1 , w_2559 );
not ( w_2559 , w_2560 );
and ( \878_b0 , \334_b0 , w_2561 );
and ( w_2560 ,  , w_2561 );
buf ( w_2559 , \291_b1 );
not ( w_2559 , w_2562 );
not (  , w_2563 );
and ( w_2562 , w_2563 , \291_b0 );
or ( \879_b1 , \878_b1 , w_2564 );
xor ( \879_b0 , \878_b0 , w_2566 );
not ( w_2566 , w_2567 );
and ( w_2567 , w_2564 , w_2565 );
buf ( w_2564 , \329_b1 );
not ( w_2564 , w_2568 );
not ( w_2565 , w_2569 );
and ( w_2568 , w_2569 , \329_b0 );
buf ( \880_b1 , \879_b1 );
buf ( \880_b0 , \879_b0 );
buf ( \881_b1 , \880_b1 );
not ( \881_b1 , w_2570 );
not ( \881_b0 , w_2571 );
and ( w_2570 , w_2571 , \880_b0 );
or ( \882_b1 , \877_b1 , w_2572 );
or ( \882_b0 , \877_b0 , \881_b0 );
not ( \881_b0 , w_2573 );
and ( w_2573 , w_2572 , \881_b1 );
or ( \883_b1 , \314_b1 , w_2574 );
or ( \883_b0 , \314_b0 , \208_b0 );
not ( \208_b0 , w_2575 );
and ( w_2575 , w_2574 , \208_b1 );
or ( \884_b1 , \883_b1 , w_2577 );
not ( w_2577 , w_2578 );
and ( \884_b0 , \883_b0 , w_2579 );
and ( w_2578 ,  , w_2579 );
buf ( w_2577 , \318_b1 );
not ( w_2577 , w_2580 );
not (  , w_2581 );
and ( w_2580 , w_2581 , \318_b0 );
or ( \885_b1 , \320_b1 , \884_b1 );
not ( \884_b1 , w_2582 );
and ( \885_b0 , \320_b0 , w_2583 );
and ( w_2582 , w_2583 , \884_b0 );
buf ( \886_b1 , \885_b1 );
not ( \886_b1 , w_2584 );
not ( \886_b0 , w_2585 );
and ( w_2584 , w_2585 , \885_b0 );
buf ( \887_b1 , \886_b1 );
not ( \887_b1 , w_2586 );
not ( \887_b0 , w_2587 );
and ( w_2586 , w_2587 , \886_b0 );
buf ( \888_b1 , \b[15]_b1 );
not ( \888_b1 , w_2588 );
not ( \888_b0 , w_2589 );
and ( w_2588 , w_2589 , \b[15]_b0 );
buf ( \889_b1 , \888_b1 );
not ( \889_b1 , w_2590 );
not ( \889_b0 , w_2591 );
and ( w_2590 , w_2591 , \888_b0 );
or ( \890_b1 , \887_b1 , \889_b1 );
not ( \889_b1 , w_2592 );
and ( \890_b0 , \887_b0 , w_2593 );
and ( w_2592 , w_2593 , \889_b0 );
or ( \891_b1 , \328_b1 , w_2595 );
not ( w_2595 , w_2596 );
and ( \891_b0 , \328_b0 , w_2597 );
and ( w_2596 ,  , w_2597 );
buf ( w_2595 , \302_b1 );
not ( w_2595 , w_2598 );
not (  , w_2599 );
and ( w_2598 , w_2599 , \302_b0 );
or ( \892_b1 , \891_b1 , w_2600 );
xor ( \892_b0 , \891_b0 , w_2602 );
not ( w_2602 , w_2603 );
and ( w_2603 , w_2600 , w_2601 );
buf ( w_2600 , \324_b1 );
not ( w_2600 , w_2604 );
not ( w_2601 , w_2605 );
and ( w_2604 , w_2605 , \324_b0 );
buf ( \893_b1 , \892_b1 );
not ( \893_b1 , w_2606 );
not ( \893_b0 , w_2607 );
and ( w_2606 , w_2607 , \892_b0 );
buf ( \894_b1 , \893_b1 );
not ( \894_b1 , w_2608 );
not ( \894_b0 , w_2609 );
and ( w_2608 , w_2609 , \893_b0 );
or ( \895_b1 , \894_b1 , \d[15]_b1 );
not ( \d[15]_b1 , w_2610 );
and ( \895_b0 , \894_b0 , w_2611 );
and ( w_2610 , w_2611 , \d[15]_b0 );
or ( \896_b1 , \890_b1 , w_2613 );
not ( w_2613 , w_2614 );
and ( \896_b0 , \890_b0 , w_2615 );
and ( w_2614 ,  , w_2615 );
buf ( w_2613 , \895_b1 );
not ( w_2613 , w_2616 );
not (  , w_2617 );
and ( w_2616 , w_2617 , \895_b0 );
or ( \897_b1 , \882_b1 , w_2619 );
not ( w_2619 , w_2620 );
and ( \897_b0 , \882_b0 , w_2621 );
and ( w_2620 ,  , w_2621 );
buf ( w_2619 , \896_b1 );
not ( w_2619 , w_2622 );
not (  , w_2623 );
and ( w_2622 , w_2623 , \896_b0 );
or ( \898_b1 , \792_b1 , w_2625 );
not ( w_2625 , w_2626 );
and ( \898_b0 , \792_b0 , w_2627 );
and ( w_2626 ,  , w_2627 );
buf ( w_2625 , \897_b1 );
not ( w_2625 , w_2628 );
not (  , w_2629 );
and ( w_2628 , w_2629 , \897_b0 );
or ( \899_b1 , \699_b1 , w_2631 );
not ( w_2631 , w_2632 );
and ( \899_b0 , \699_b0 , w_2633 );
and ( w_2632 ,  , w_2633 );
buf ( w_2631 , \898_b1 );
not ( w_2631 , w_2634 );
not (  , w_2635 );
and ( w_2634 , w_2635 , \898_b0 );
or ( \900_b1 , \668_b1 , w_2637 );
not ( w_2637 , w_2638 );
and ( \900_b0 , \668_b0 , w_2639 );
and ( w_2638 ,  , w_2639 );
buf ( w_2637 , \899_b1 );
not ( w_2637 , w_2640 );
not (  , w_2641 );
and ( w_2640 , w_2641 , \899_b0 );
or ( \901_b1 , \651_b1 , w_2643 );
not ( w_2643 , w_2644 );
and ( \901_b0 , \651_b0 , w_2645 );
and ( w_2644 ,  , w_2645 );
buf ( w_2643 , \900_b1 );
not ( w_2643 , w_2646 );
not (  , w_2647 );
and ( w_2646 , w_2647 , \900_b0 );
buf ( \902_b1 , \685_b1 );
not ( \902_b1 , w_2648 );
not ( \902_b0 , w_2649 );
and ( w_2648 , w_2649 , \685_b0 );
buf ( \903_b1 , \697_b1 );
buf ( \903_b0 , \697_b0 );
or ( \904_b1 , \902_b1 , \903_b1 );
not ( \903_b1 , w_2650 );
and ( \904_b0 , \902_b0 , w_2651 );
and ( w_2650 , w_2651 , \903_b0 );
buf ( \905_b1 , \312_b1 );
not ( \905_b1 , w_2652 );
not ( \905_b0 , w_2653 );
and ( w_2652 , w_2653 , \312_b0 );
or ( \906_b1 , \905_b1 , w_2655 );
not ( w_2655 , w_2656 );
and ( \906_b0 , \905_b0 , w_2657 );
and ( w_2656 ,  , w_2657 );
buf ( w_2655 , \323_b1 );
not ( w_2655 , w_2658 );
not (  , w_2659 );
and ( w_2658 , w_2659 , \323_b0 );
or ( \907_b1 , \906_b1 , \320_b1 );
xor ( \907_b0 , \906_b0 , w_2660 );
not ( w_2660 , w_2661 );
and ( w_2661 , \320_b1 , \320_b0 );
buf ( \908_b1 , \907_b1 );
not ( \908_b1 , w_2662 );
not ( \908_b0 , w_2663 );
and ( w_2662 , w_2663 , \907_b0 );
buf ( \909_b1 , \908_b1 );
not ( \909_b1 , w_2664 );
not ( \909_b0 , w_2665 );
and ( w_2664 , w_2665 , \908_b0 );
or ( \910_b1 , \904_b1 , w_2667 );
not ( w_2667 , w_2668 );
and ( \910_b0 , \904_b0 , w_2669 );
and ( w_2668 ,  , w_2669 );
buf ( w_2667 , \909_b1 );
not ( w_2667 , w_2670 );
not (  , w_2671 );
and ( w_2670 , w_2671 , \909_b0 );
buf ( \911_b1 , \471_b1 );
not ( \911_b1 , w_2672 );
not ( \911_b0 , w_2673 );
and ( w_2672 , w_2673 , \471_b0 );
buf ( \912_b1 , \347_b1 );
not ( \912_b1 , w_2674 );
not ( \912_b0 , w_2675 );
and ( w_2674 , w_2675 , \347_b0 );
or ( \913_b1 , \911_b1 , w_2676 );
or ( \913_b0 , \911_b0 , \912_b0 );
not ( \912_b0 , w_2677 );
and ( w_2677 , w_2676 , \912_b1 );
or ( \914_b1 , \541_b1 , w_2679 );
not ( w_2679 , w_2680 );
and ( \914_b0 , \541_b0 , w_2681 );
and ( w_2680 ,  , w_2681 );
buf ( w_2679 , \542_b1 );
not ( w_2679 , w_2682 );
not (  , w_2683 );
and ( w_2682 , w_2683 , \542_b0 );
or ( \915_b1 , \913_b1 , w_2685 );
not ( w_2685 , w_2686 );
and ( \915_b0 , \913_b0 , w_2687 );
and ( w_2686 ,  , w_2687 );
buf ( w_2685 , \914_b1 );
not ( w_2685 , w_2688 );
not (  , w_2689 );
and ( w_2688 , w_2689 , \914_b0 );
or ( \916_b1 , \523_b1 , w_2690 );
xor ( \916_b0 , \523_b0 , w_2692 );
not ( w_2692 , w_2693 );
and ( w_2693 , w_2690 , w_2691 );
buf ( w_2690 , \531_b1 );
not ( w_2690 , w_2694 );
not ( w_2691 , w_2695 );
and ( w_2694 , w_2695 , \531_b0 );
buf ( \917_b1 , \916_b1 );
not ( \917_b1 , w_2696 );
not ( \917_b0 , w_2697 );
and ( w_2696 , w_2697 , \916_b0 );
or ( \918_b1 , \915_b1 , \917_b1 );
not ( \917_b1 , w_2698 );
and ( \918_b0 , \915_b0 , w_2699 );
and ( w_2698 , w_2699 , \917_b0 );
buf ( \919_b1 , \915_b1 );
not ( \919_b1 , w_2700 );
not ( \919_b0 , w_2701 );
and ( w_2700 , w_2701 , \915_b0 );
or ( \920_b1 , \919_b1 , \916_b1 );
not ( \916_b1 , w_2702 );
and ( \920_b0 , \919_b0 , w_2703 );
and ( w_2702 , w_2703 , \916_b0 );
or ( \921_b1 , \918_b1 , w_2705 );
not ( w_2705 , w_2706 );
and ( \921_b0 , \918_b0 , w_2707 );
and ( w_2706 ,  , w_2707 );
buf ( w_2705 , \920_b1 );
not ( w_2705 , w_2708 );
not (  , w_2709 );
and ( w_2708 , w_2709 , \920_b0 );
buf ( \922_b1 , \921_b1 );
buf ( \922_b0 , \921_b0 );
or ( \923_b1 , \922_b1 , w_2711 );
not ( w_2711 , w_2712 );
and ( \923_b0 , \922_b0 , w_2713 );
and ( w_2712 ,  , w_2713 );
buf ( w_2711 , \b[15]_b1 );
not ( w_2711 , w_2714 );
not (  , w_2715 );
and ( w_2714 , w_2715 , \b[15]_b0 );
or ( \924_b1 , \910_b1 , \923_b1 );
not ( \923_b1 , w_2716 );
and ( \924_b0 , \910_b0 , w_2717 );
and ( w_2716 , w_2717 , \923_b0 );
buf ( \925_b1 , \c[15]_b1 );
not ( \925_b1 , w_2718 );
not ( \925_b0 , w_2719 );
and ( w_2718 , w_2719 , \c[15]_b0 );
or ( \926_b1 , \924_b1 , w_2721 );
not ( w_2721 , w_2722 );
and ( \926_b0 , \924_b0 , w_2723 );
and ( w_2722 ,  , w_2723 );
buf ( w_2721 , \925_b1 );
not ( w_2721 , w_2724 );
not (  , w_2725 );
and ( w_2724 , w_2725 , \925_b0 );
or ( \927_b1 , \901_b1 , w_2727 );
not ( w_2727 , w_2728 );
and ( \927_b0 , \901_b0 , w_2729 );
and ( w_2728 ,  , w_2729 );
buf ( w_2727 , \926_b1 );
not ( w_2727 , w_2730 );
not (  , w_2731 );
and ( w_2730 , w_2731 , \926_b0 );
or ( \928_b1 , \d[5]_b1 , \a[6]_b1 );
xor ( \928_b0 , \d[5]_b0 , w_2732 );
not ( w_2732 , w_2733 );
and ( w_2733 , \a[6]_b1 , \a[6]_b0 );
buf ( \929_b1 , \928_b1 );
not ( \929_b1 , w_2734 );
not ( \929_b0 , w_2735 );
and ( w_2734 , w_2735 , \928_b0 );
or ( \930_b1 , \d[5]_b1 , \d[4]_b1 );
xor ( \930_b0 , \d[5]_b0 , w_2736 );
not ( w_2736 , w_2737 );
and ( w_2737 , \d[4]_b1 , \d[4]_b0 );
buf ( \931_b1 , \930_b1 );
not ( \931_b1 , w_2738 );
not ( \931_b0 , w_2739 );
and ( w_2738 , w_2739 , \930_b0 );
or ( \932_b1 , \d[4]_b1 , \d[3]_b1 );
xor ( \932_b0 , \d[4]_b0 , w_2740 );
not ( w_2740 , w_2741 );
and ( w_2741 , \d[3]_b1 , \d[3]_b0 );
or ( \933_b1 , \931_b1 , w_2743 );
not ( w_2743 , w_2744 );
and ( \933_b0 , \931_b0 , w_2745 );
and ( w_2744 ,  , w_2745 );
buf ( w_2743 , \932_b1 );
not ( w_2743 , w_2746 );
not (  , w_2747 );
and ( w_2746 , w_2747 , \932_b0 );
buf ( \934_b1 , \933_b1 );
not ( \934_b1 , w_2748 );
not ( \934_b0 , w_2749 );
and ( w_2748 , w_2749 , \933_b0 );
or ( \935_b1 , \929_b1 , w_2750 );
or ( \935_b0 , \929_b0 , \934_b0 );
not ( \934_b0 , w_2751 );
and ( w_2751 , w_2750 , \934_b1 );
buf ( \936_b1 , \932_b1 );
buf ( \936_b0 , \932_b0 );
or ( \937_b1 , \d[5]_b1 , \a[7]_b1 );
xor ( \937_b0 , \d[5]_b0 , w_2752 );
not ( w_2752 , w_2753 );
and ( w_2753 , \a[7]_b1 , \a[7]_b0 );
or ( \938_b1 , \936_b1 , w_2755 );
not ( w_2755 , w_2756 );
and ( \938_b0 , \936_b0 , w_2757 );
and ( w_2756 ,  , w_2757 );
buf ( w_2755 , \937_b1 );
not ( w_2755 , w_2758 );
not (  , w_2759 );
and ( w_2758 , w_2759 , \937_b0 );
or ( \939_b1 , \935_b1 , w_2761 );
not ( w_2761 , w_2762 );
and ( \939_b0 , \935_b0 , w_2763 );
and ( w_2762 ,  , w_2763 );
buf ( w_2761 , \938_b1 );
not ( w_2761 , w_2764 );
not (  , w_2765 );
and ( w_2764 , w_2765 , \938_b0 );
or ( \940_b1 , \a[0]_b1 , \d[11]_b1 );
xor ( \940_b0 , \a[0]_b0 , w_2766 );
not ( w_2766 , w_2767 );
and ( w_2767 , \d[11]_b1 , \d[11]_b0 );
buf ( \941_b1 , \940_b1 );
not ( \941_b1 , w_2768 );
not ( \941_b0 , w_2769 );
and ( w_2768 , w_2769 , \940_b0 );
or ( \942_b1 , \d[11]_b1 , w_2770 );
xor ( \942_b0 , \d[11]_b0 , w_2772 );
not ( w_2772 , w_2773 );
and ( w_2773 , w_2770 , w_2771 );
buf ( w_2770 , \d[10]_b1 );
not ( w_2770 , w_2774 );
not ( w_2771 , w_2775 );
and ( w_2774 , w_2775 , \d[10]_b0 );
or ( \943_b1 , \d[10]_b1 , \d[9]_b1 );
xor ( \943_b0 , \d[10]_b0 , w_2776 );
not ( w_2776 , w_2777 );
and ( w_2777 , \d[9]_b1 , \d[9]_b0 );
or ( \944_b1 , \942_b1 , w_2779 );
not ( w_2779 , w_2780 );
and ( \944_b0 , \942_b0 , w_2781 );
and ( w_2780 ,  , w_2781 );
buf ( w_2779 , \943_b1 );
not ( w_2779 , w_2782 );
not (  , w_2783 );
and ( w_2782 , w_2783 , \943_b0 );
buf ( \945_b1 , \944_b1 );
not ( \945_b1 , w_2784 );
not ( \945_b0 , w_2785 );
and ( w_2784 , w_2785 , \944_b0 );
or ( \946_b1 , \941_b1 , w_2786 );
or ( \946_b0 , \941_b0 , \945_b0 );
not ( \945_b0 , w_2787 );
and ( w_2787 , w_2786 , \945_b1 );
or ( \947_b1 , \d[10]_b1 , \d[9]_b1 );
xor ( \947_b0 , \d[10]_b0 , w_2788 );
not ( w_2788 , w_2789 );
and ( w_2789 , \d[9]_b1 , \d[9]_b0 );
or ( \948_b1 , \a[1]_b1 , \d[11]_b1 );
xor ( \948_b0 , \a[1]_b0 , w_2790 );
not ( w_2790 , w_2791 );
and ( w_2791 , \d[11]_b1 , \d[11]_b0 );
or ( \949_b1 , \947_b1 , w_2793 );
not ( w_2793 , w_2794 );
and ( \949_b0 , \947_b0 , w_2795 );
and ( w_2794 ,  , w_2795 );
buf ( w_2793 , \948_b1 );
not ( w_2793 , w_2796 );
not (  , w_2797 );
and ( w_2796 , w_2797 , \948_b0 );
or ( \950_b1 , \946_b1 , w_2799 );
not ( w_2799 , w_2800 );
and ( \950_b0 , \946_b0 , w_2801 );
and ( w_2800 ,  , w_2801 );
buf ( w_2799 , \949_b1 );
not ( w_2799 , w_2802 );
not (  , w_2803 );
and ( w_2802 , w_2803 , \949_b0 );
buf ( \951_b1 , \950_b1 );
not ( \951_b1 , w_2804 );
not ( \951_b0 , w_2805 );
and ( w_2804 , w_2805 , \950_b0 );
or ( \952_b1 , \939_b1 , \951_b1 );
xor ( \952_b0 , \939_b0 , w_2806 );
not ( w_2806 , w_2807 );
and ( w_2807 , \951_b1 , \951_b0 );
or ( \953_b1 , \a[0]_b1 , w_2808 );
or ( \953_b0 , \a[0]_b0 , \d[10]_b0 );
not ( \d[10]_b0 , w_2809 );
and ( w_2809 , w_2808 , \d[10]_b1 );
or ( \954_b1 , \953_b1 , w_2811 );
not ( w_2811 , w_2812 );
and ( \954_b0 , \953_b0 , w_2813 );
and ( w_2812 ,  , w_2813 );
buf ( w_2811 , \d[9]_b1 );
not ( w_2811 , w_2814 );
not (  , w_2815 );
and ( w_2814 , w_2815 , \d[9]_b0 );
or ( \955_b1 , \a[0]_b1 , w_2817 );
not ( w_2817 , w_2818 );
and ( \955_b0 , \a[0]_b0 , w_2819 );
and ( w_2818 ,  , w_2819 );
buf ( w_2817 , \d[10]_b1 );
not ( w_2817 , w_2820 );
not (  , w_2821 );
and ( w_2820 , w_2821 , \d[10]_b0 );
or ( \957_b1 , \a[8]_b1 , \d[3]_b1 );
xor ( \957_b0 , \a[8]_b0 , w_2822 );
not ( w_2822 , w_2823 );
and ( w_2823 , \d[3]_b1 , \d[3]_b0 );
buf ( \958_b1 , \957_b1 );
not ( \958_b1 , w_2824 );
not ( \958_b0 , w_2825 );
and ( w_2824 , w_2825 , \957_b0 );
or ( \959_b1 , \d[2]_b1 , \d[1]_b1 );
xor ( \959_b0 , \d[2]_b0 , w_2826 );
not ( w_2826 , w_2827 );
and ( w_2827 , \d[1]_b1 , \d[1]_b0 );
buf ( \960_b1 , \959_b1 );
not ( \960_b1 , w_2828 );
not ( \960_b0 , w_2829 );
and ( w_2828 , w_2829 , \959_b0 );
or ( \961_b1 , \d[3]_b1 , \d[2]_b1 );
xor ( \961_b0 , \d[3]_b0 , w_2830 );
not ( w_2830 , w_2831 );
and ( w_2831 , \d[2]_b1 , \d[2]_b0 );
or ( \962_b1 , \960_b1 , \961_b1 );
not ( \961_b1 , w_2832 );
and ( \962_b0 , \960_b0 , w_2833 );
and ( w_2832 , w_2833 , \961_b0 );
buf ( \963_b1 , \962_b1 );
not ( \963_b1 , w_2834 );
not ( \963_b0 , w_2835 );
and ( w_2834 , w_2835 , \962_b0 );
or ( \964_b1 , \958_b1 , w_2836 );
or ( \964_b0 , \958_b0 , \963_b0 );
not ( \963_b0 , w_2837 );
and ( w_2837 , w_2836 , \963_b1 );
buf ( \965_b1 , \959_b1 );
buf ( \965_b0 , \959_b0 );
or ( \966_b1 , \a[9]_b1 , \d[3]_b1 );
xor ( \966_b0 , \a[9]_b0 , w_2838 );
not ( w_2838 , w_2839 );
and ( w_2839 , \d[3]_b1 , \d[3]_b0 );
or ( \967_b1 , \965_b1 , w_2841 );
not ( w_2841 , w_2842 );
and ( \967_b0 , \965_b0 , w_2843 );
and ( w_2842 ,  , w_2843 );
buf ( w_2841 , \966_b1 );
not ( w_2841 , w_2844 );
not (  , w_2845 );
and ( w_2844 , w_2845 , \966_b0 );
or ( \968_b1 , \964_b1 , w_2847 );
not ( w_2847 , w_2848 );
and ( \968_b0 , \964_b0 , w_2849 );
and ( w_2848 ,  , w_2849 );
buf ( w_2847 , \967_b1 );
not ( w_2847 , w_2850 );
not (  , w_2851 );
and ( w_2850 , w_2851 , \967_b0 );
or ( \969_b1 , \956_b1 , \968_b1 );
xor ( \969_b0 , \956_b0 , w_2852 );
not ( w_2852 , w_2853 );
and ( w_2853 , \968_b1 , \968_b0 );
or ( \970_b1 , \952_b1 , w_2854 );
xor ( \970_b0 , \952_b0 , w_2856 );
not ( w_2856 , w_2857 );
and ( w_2857 , w_2854 , w_2855 );
buf ( w_2854 , \969_b1 );
not ( w_2854 , w_2858 );
not ( w_2855 , w_2859 );
and ( w_2858 , w_2859 , \969_b0 );
or ( \971_b1 , \a[0]_b1 , w_2860 );
or ( \971_b0 , \a[0]_b0 , \d[8]_b0 );
not ( \d[8]_b0 , w_2861 );
and ( w_2861 , w_2860 , \d[8]_b1 );
or ( \972_b1 , \971_b1 , w_2863 );
not ( w_2863 , w_2864 );
and ( \972_b0 , \971_b0 , w_2865 );
and ( w_2864 ,  , w_2865 );
buf ( w_2863 , \d[7]_b1 );
not ( w_2863 , w_2866 );
not (  , w_2867 );
and ( w_2866 , w_2867 , \d[7]_b0 );
or ( \973_b1 , \a[0]_b1 , w_2869 );
not ( w_2869 , w_2870 );
and ( \973_b0 , \a[0]_b0 , w_2871 );
and ( w_2870 ,  , w_2871 );
buf ( w_2869 , \d[8]_b1 );
not ( w_2869 , w_2872 );
not (  , w_2873 );
and ( w_2872 , w_2873 , \d[8]_b0 );
buf ( \975_b1 , \974_b1 );
not ( \975_b1 , w_2874 );
not ( \975_b0 , w_2875 );
and ( w_2874 , w_2875 , \974_b0 );
or ( \976_b1 , \a[6]_b1 , \d[3]_b1 );
xor ( \976_b0 , \a[6]_b0 , w_2876 );
not ( w_2876 , w_2877 );
and ( w_2877 , \d[3]_b1 , \d[3]_b0 );
buf ( \977_b1 , \976_b1 );
not ( \977_b1 , w_2878 );
not ( \977_b0 , w_2879 );
and ( w_2878 , w_2879 , \976_b0 );
or ( \978_b1 , \d[3]_b1 , \d[2]_b1 );
xor ( \978_b0 , \d[3]_b0 , w_2880 );
not ( w_2880 , w_2881 );
and ( w_2881 , \d[2]_b1 , \d[2]_b0 );
buf ( \979_b1 , \978_b1 );
not ( \979_b1 , w_2882 );
not ( \979_b0 , w_2883 );
and ( w_2882 , w_2883 , \978_b0 );
or ( \980_b1 , \979_b1 , w_2885 );
not ( w_2885 , w_2886 );
and ( \980_b0 , \979_b0 , w_2887 );
and ( w_2886 ,  , w_2887 );
buf ( w_2885 , \959_b1 );
not ( w_2885 , w_2888 );
not (  , w_2889 );
and ( w_2888 , w_2889 , \959_b0 );
buf ( \981_b1 , \980_b1 );
not ( \981_b1 , w_2890 );
not ( \981_b0 , w_2891 );
and ( w_2890 , w_2891 , \980_b0 );
or ( \982_b1 , \977_b1 , w_2892 );
or ( \982_b0 , \977_b0 , \981_b0 );
not ( \981_b0 , w_2893 );
and ( w_2893 , w_2892 , \981_b1 );
or ( \983_b1 , \a[7]_b1 , \d[3]_b1 );
xor ( \983_b0 , \a[7]_b0 , w_2894 );
not ( w_2894 , w_2895 );
and ( w_2895 , \d[3]_b1 , \d[3]_b0 );
or ( \984_b1 , \965_b1 , w_2897 );
not ( w_2897 , w_2898 );
and ( \984_b0 , \965_b0 , w_2899 );
and ( w_2898 ,  , w_2899 );
buf ( w_2897 , \983_b1 );
not ( w_2897 , w_2900 );
not (  , w_2901 );
and ( w_2900 , w_2901 , \983_b0 );
or ( \985_b1 , \982_b1 , w_2903 );
not ( w_2903 , w_2904 );
and ( \985_b0 , \982_b0 , w_2905 );
and ( w_2904 ,  , w_2905 );
buf ( w_2903 , \984_b1 );
not ( w_2903 , w_2906 );
not (  , w_2907 );
and ( w_2906 , w_2907 , \984_b0 );
or ( \986_b1 , \975_b1 , w_2909 );
not ( w_2909 , w_2910 );
and ( \986_b0 , \975_b0 , w_2911 );
and ( w_2910 ,  , w_2911 );
buf ( w_2909 , \985_b1 );
not ( w_2909 , w_2912 );
not (  , w_2913 );
and ( w_2912 , w_2913 , \985_b0 );
buf ( \987_b1 , \986_b1 );
not ( \987_b1 , w_2914 );
not ( \987_b0 , w_2915 );
and ( w_2914 , w_2915 , \986_b0 );
or ( \988_b1 , \943_b1 , w_2917 );
not ( w_2917 , w_2918 );
and ( \988_b0 , \943_b0 , w_2919 );
and ( w_2918 ,  , w_2919 );
buf ( w_2917 , \a[0]_b1 );
not ( w_2917 , w_2920 );
not (  , w_2921 );
and ( w_2920 , w_2921 , \a[0]_b0 );
buf ( \989_b1 , \988_b1 );
not ( \989_b1 , w_2922 );
not ( \989_b0 , w_2923 );
and ( w_2922 , w_2923 , \988_b0 );
or ( \990_b1 , \983_b1 , w_2925 );
not ( w_2925 , w_2926 );
and ( \990_b0 , \983_b0 , w_2927 );
and ( w_2926 ,  , w_2927 );
buf ( w_2925 , \978_b1 );
not ( w_2925 , w_2928 );
not (  , w_2929 );
and ( w_2928 , w_2929 , \978_b0 );
or ( \991_b1 , \959_b1 , w_2930 );
or ( \991_b0 , \959_b0 , \990_b0 );
not ( \990_b0 , w_2931 );
and ( w_2931 , w_2930 , \990_b1 );
or ( \992_b1 , \959_b1 , w_2933 );
not ( w_2933 , w_2934 );
and ( \992_b0 , \959_b0 , w_2935 );
and ( w_2934 ,  , w_2935 );
buf ( w_2933 , \957_b1 );
not ( w_2933 , w_2936 );
not (  , w_2937 );
and ( w_2936 , w_2937 , \957_b0 );
or ( \993_b1 , \991_b1 , w_2939 );
not ( w_2939 , w_2940 );
and ( \993_b0 , \991_b0 , w_2941 );
and ( w_2940 ,  , w_2941 );
buf ( w_2939 , \992_b1 );
not ( w_2939 , w_2942 );
not (  , w_2943 );
and ( w_2942 , w_2943 , \992_b0 );
or ( \994_b1 , \989_b1 , \993_b1 );
xor ( \994_b0 , \989_b0 , w_2944 );
not ( w_2944 , w_2945 );
and ( w_2945 , \993_b1 , \993_b0 );
or ( \995_b1 , \d[7]_b1 , \a[3]_b1 );
xor ( \995_b0 , \d[7]_b0 , w_2946 );
not ( w_2946 , w_2947 );
and ( w_2947 , \a[3]_b1 , \a[3]_b0 );
buf ( \996_b1 , \995_b1 );
not ( \996_b1 , w_2948 );
not ( \996_b0 , w_2949 );
and ( w_2948 , w_2949 , \995_b0 );
or ( \997_b1 , \d[7]_b1 , w_2950 );
xor ( \997_b0 , \d[7]_b0 , w_2952 );
not ( w_2952 , w_2953 );
and ( w_2953 , w_2950 , w_2951 );
buf ( w_2950 , \d[6]_b1 );
not ( w_2950 , w_2954 );
not ( w_2951 , w_2955 );
and ( w_2954 , w_2955 , \d[6]_b0 );
or ( \998_b1 , \d[6]_b1 , \d[5]_b1 );
xor ( \998_b0 , \d[6]_b0 , w_2956 );
not ( w_2956 , w_2957 );
and ( w_2957 , \d[5]_b1 , \d[5]_b0 );
or ( \999_b1 , \997_b1 , w_2959 );
not ( w_2959 , w_2960 );
and ( \999_b0 , \997_b0 , w_2961 );
and ( w_2960 ,  , w_2961 );
buf ( w_2959 , \998_b1 );
not ( w_2959 , w_2962 );
not (  , w_2963 );
and ( w_2962 , w_2963 , \998_b0 );
buf ( \1000_b1 , \999_b1 );
not ( \1000_b1 , w_2964 );
not ( \1000_b0 , w_2965 );
and ( w_2964 , w_2965 , \999_b0 );
or ( \1001_b1 , \996_b1 , w_2966 );
or ( \1001_b0 , \996_b0 , \1000_b0 );
not ( \1000_b0 , w_2967 );
and ( w_2967 , w_2966 , \1000_b1 );
buf ( \1002_b1 , \998_b1 );
not ( \1002_b1 , w_2968 );
not ( \1002_b0 , w_2969 );
and ( w_2968 , w_2969 , \998_b0 );
buf ( \1003_b1 , \1002_b1 );
not ( \1003_b1 , w_2970 );
not ( \1003_b0 , w_2971 );
and ( w_2970 , w_2971 , \1002_b0 );
or ( \1004_b1 , \d[7]_b1 , \a[4]_b1 );
xor ( \1004_b0 , \d[7]_b0 , w_2972 );
not ( w_2972 , w_2973 );
and ( w_2973 , \a[4]_b1 , \a[4]_b0 );
or ( \1005_b1 , \1003_b1 , w_2975 );
not ( w_2975 , w_2976 );
and ( \1005_b0 , \1003_b0 , w_2977 );
and ( w_2976 ,  , w_2977 );
buf ( w_2975 , \1004_b1 );
not ( w_2975 , w_2978 );
not (  , w_2979 );
and ( w_2978 , w_2979 , \1004_b0 );
or ( \1006_b1 , \1001_b1 , w_2981 );
not ( w_2981 , w_2982 );
and ( \1006_b0 , \1001_b0 , w_2983 );
and ( w_2982 ,  , w_2983 );
buf ( w_2981 , \1005_b1 );
not ( w_2981 , w_2984 );
not (  , w_2985 );
and ( w_2984 , w_2985 , \1005_b0 );
or ( \1007_b1 , \994_b1 , w_2986 );
xor ( \1007_b0 , \994_b0 , w_2988 );
not ( w_2988 , w_2989 );
and ( w_2989 , w_2986 , w_2987 );
buf ( w_2986 , \1006_b1 );
not ( w_2986 , w_2990 );
not ( w_2987 , w_2991 );
and ( w_2990 , w_2991 , \1006_b0 );
buf ( \1008_b1 , \1007_b1 );
not ( \1008_b1 , w_2992 );
not ( \1008_b0 , w_2993 );
and ( w_2992 , w_2993 , \1007_b0 );
or ( \1009_b1 , \987_b1 , w_2994 );
or ( \1009_b0 , \987_b0 , \1008_b0 );
not ( \1008_b0 , w_2995 );
and ( w_2995 , w_2994 , \1008_b1 );
buf ( \1010_b1 , \d[0]_b1 );
not ( \1010_b1 , w_2996 );
not ( \1010_b0 , w_2997 );
and ( w_2996 , w_2997 , \d[0]_b0 );
or ( \1011_b1 , \1010_b1 , w_2999 );
not ( w_2999 , w_3000 );
and ( \1011_b0 , \1010_b0 , w_3001 );
and ( w_3000 ,  , w_3001 );
buf ( w_2999 , \d[1]_b1 );
not ( w_2999 , w_3002 );
not (  , w_3003 );
and ( w_3002 , w_3003 , \d[1]_b0 );
buf ( \1012_b1 , \1011_b1 );
not ( \1012_b1 , w_3004 );
not ( \1012_b0 , w_3005 );
and ( w_3004 , w_3005 , \1011_b0 );
or ( \1013_b1 , \d[1]_b1 , \a[8]_b1 );
xor ( \1013_b0 , \d[1]_b0 , w_3006 );
not ( w_3006 , w_3007 );
and ( w_3007 , \a[8]_b1 , \a[8]_b0 );
or ( \1014_b1 , \1012_b1 , \1013_b1 );
not ( \1013_b1 , w_3008 );
and ( \1014_b0 , \1012_b0 , w_3009 );
and ( w_3008 , w_3009 , \1013_b0 );
or ( \1015_b1 , \d[1]_b1 , \a[9]_b1 );
xor ( \1015_b0 , \d[1]_b0 , w_3010 );
not ( w_3010 , w_3011 );
and ( w_3011 , \a[9]_b1 , \a[9]_b0 );
or ( \1016_b1 , \1015_b1 , \d[0]_b1 );
not ( \d[0]_b1 , w_3012 );
and ( \1016_b0 , \1015_b0 , w_3013 );
and ( w_3012 , w_3013 , \d[0]_b0 );
or ( \1017_b1 , \1014_b1 , w_3015 );
not ( w_3015 , w_3016 );
and ( \1017_b0 , \1014_b0 , w_3017 );
and ( w_3016 ,  , w_3017 );
buf ( w_3015 , \1016_b1 );
not ( w_3015 , w_3018 );
not (  , w_3019 );
and ( w_3018 , w_3019 , \1016_b0 );
buf ( \1018_b1 , \1017_b1 );
not ( \1018_b1 , w_3020 );
not ( \1018_b0 , w_3021 );
and ( w_3020 , w_3021 , \1017_b0 );
buf ( \1019_b1 , \1018_b1 );
not ( \1019_b1 , w_3022 );
not ( \1019_b0 , w_3023 );
and ( w_3022 , w_3023 , \1018_b0 );
or ( \1020_b1 , \d[9]_b1 , \a[0]_b1 );
xor ( \1020_b0 , \d[9]_b0 , w_3024 );
not ( w_3024 , w_3025 );
and ( w_3025 , \a[0]_b1 , \a[0]_b0 );
buf ( \1021_b1 , \1020_b1 );
not ( \1021_b1 , w_3026 );
not ( \1021_b0 , w_3027 );
and ( w_3026 , w_3027 , \1020_b0 );
or ( \1022_b1 , \d[9]_b1 , w_3028 );
or ( \1022_b0 , \d[9]_b0 , \d[8]_b0 );
not ( \d[8]_b0 , w_3029 );
and ( w_3029 , w_3028 , \d[8]_b1 );
buf ( \1023_b1 , \d[7]_b1 );
not ( \1023_b1 , w_3030 );
not ( \1023_b0 , w_3031 );
and ( w_3030 , w_3031 , \d[7]_b0 );
or ( \1024_b1 , \1023_b1 , w_3033 );
not ( w_3033 , w_3034 );
and ( \1024_b0 , \1023_b0 , w_3035 );
and ( w_3034 ,  , w_3035 );
buf ( w_3033 , \d[8]_b1 );
not ( w_3033 , w_3036 );
not (  , w_3037 );
and ( w_3036 , w_3037 , \d[8]_b0 );
or ( \1025_b1 , \d[9]_b1 , w_3039 );
not ( w_3039 , w_3040 );
and ( \1025_b0 , \d[9]_b0 , w_3041 );
and ( w_3040 ,  , w_3041 );
buf ( w_3039 , \d[7]_b1 );
not ( w_3039 , w_3042 );
not (  , w_3043 );
and ( w_3042 , w_3043 , \d[7]_b0 );
buf ( \1027_b1 , \1026_b1 );
not ( \1027_b1 , w_3044 );
not ( \1027_b0 , w_3045 );
and ( w_3044 , w_3045 , \1026_b0 );
or ( \1028_b1 , \1021_b1 , w_3046 );
or ( \1028_b0 , \1021_b0 , \1027_b0 );
not ( \1027_b0 , w_3047 );
and ( w_3047 , w_3046 , \1027_b1 );
or ( \1029_b1 , \d[8]_b1 , \d[7]_b1 );
xor ( \1029_b0 , \d[8]_b0 , w_3048 );
not ( w_3048 , w_3049 );
and ( w_3049 , \d[7]_b1 , \d[7]_b0 );
or ( \1030_b1 , \d[9]_b1 , \a[1]_b1 );
xor ( \1030_b0 , \d[9]_b0 , w_3050 );
not ( w_3050 , w_3051 );
and ( w_3051 , \a[1]_b1 , \a[1]_b0 );
or ( \1031_b1 , \1029_b1 , w_3053 );
not ( w_3053 , w_3054 );
and ( \1031_b0 , \1029_b0 , w_3055 );
and ( w_3054 ,  , w_3055 );
buf ( w_3053 , \1030_b1 );
not ( w_3053 , w_3056 );
not (  , w_3057 );
and ( w_3056 , w_3057 , \1030_b0 );
or ( \1032_b1 , \1028_b1 , w_3059 );
not ( w_3059 , w_3060 );
and ( \1032_b0 , \1028_b0 , w_3061 );
and ( w_3060 ,  , w_3061 );
buf ( w_3059 , \1031_b1 );
not ( w_3059 , w_3062 );
not (  , w_3063 );
and ( w_3062 , w_3063 , \1031_b0 );
buf ( \1033_b1 , \1032_b1 );
not ( \1033_b1 , w_3064 );
not ( \1033_b0 , w_3065 );
and ( w_3064 , w_3065 , \1032_b0 );
or ( \1034_b1 , \1019_b1 , w_3066 );
or ( \1034_b0 , \1019_b0 , \1033_b0 );
not ( \1033_b0 , w_3067 );
and ( w_3067 , w_3066 , \1033_b1 );
or ( \1035_b1 , \1032_b1 , w_3068 );
or ( \1035_b0 , \1032_b0 , \1018_b0 );
not ( \1018_b0 , w_3069 );
and ( w_3069 , w_3068 , \1018_b1 );
or ( \1036_b1 , \d[7]_b1 , \a[2]_b1 );
xor ( \1036_b0 , \d[7]_b0 , w_3070 );
not ( w_3070 , w_3071 );
and ( w_3071 , \a[2]_b1 , \a[2]_b0 );
buf ( \1037_b1 , \1036_b1 );
not ( \1037_b1 , w_3072 );
not ( \1037_b0 , w_3073 );
and ( w_3072 , w_3073 , \1036_b0 );
or ( \1038_b1 , \997_b1 , w_3075 );
not ( w_3075 , w_3076 );
and ( \1038_b0 , \997_b0 , w_3077 );
and ( w_3076 ,  , w_3077 );
buf ( w_3075 , \998_b1 );
not ( w_3075 , w_3078 );
not (  , w_3079 );
and ( w_3078 , w_3079 , \998_b0 );
buf ( \1039_b1 , \1038_b1 );
not ( \1039_b1 , w_3080 );
not ( \1039_b0 , w_3081 );
and ( w_3080 , w_3081 , \1038_b0 );
or ( \1040_b1 , \1037_b1 , w_3082 );
or ( \1040_b0 , \1037_b0 , \1039_b0 );
not ( \1039_b0 , w_3083 );
and ( w_3083 , w_3082 , \1039_b1 );
buf ( \1041_b1 , \1002_b1 );
not ( \1041_b1 , w_3084 );
not ( \1041_b0 , w_3085 );
and ( w_3084 , w_3085 , \1002_b0 );
or ( \1042_b1 , \1041_b1 , w_3087 );
not ( w_3087 , w_3088 );
and ( \1042_b0 , \1041_b0 , w_3089 );
and ( w_3088 ,  , w_3089 );
buf ( w_3087 , \995_b1 );
not ( w_3087 , w_3090 );
not (  , w_3091 );
and ( w_3090 , w_3091 , \995_b0 );
or ( \1043_b1 , \1040_b1 , w_3093 );
not ( w_3093 , w_3094 );
and ( \1043_b0 , \1040_b0 , w_3095 );
and ( w_3094 ,  , w_3095 );
buf ( w_3093 , \1042_b1 );
not ( w_3093 , w_3096 );
not (  , w_3097 );
and ( w_3096 , w_3097 , \1042_b0 );
or ( \1044_b1 , \1035_b1 , w_3099 );
not ( w_3099 , w_3100 );
and ( \1044_b0 , \1035_b0 , w_3101 );
and ( w_3100 ,  , w_3101 );
buf ( w_3099 , \1043_b1 );
not ( w_3099 , w_3102 );
not (  , w_3103 );
and ( w_3102 , w_3103 , \1043_b0 );
or ( \1045_b1 , \1034_b1 , w_3105 );
not ( w_3105 , w_3106 );
and ( \1045_b0 , \1034_b0 , w_3107 );
and ( w_3106 ,  , w_3107 );
buf ( w_3105 , \1044_b1 );
not ( w_3105 , w_3108 );
not (  , w_3109 );
and ( w_3108 , w_3109 , \1044_b0 );
or ( \1046_b1 , \1009_b1 , w_3111 );
not ( w_3111 , w_3112 );
and ( \1046_b0 , \1009_b0 , w_3113 );
and ( w_3112 ,  , w_3113 );
buf ( w_3111 , \1045_b1 );
not ( w_3111 , w_3114 );
not (  , w_3115 );
and ( w_3114 , w_3115 , \1045_b0 );
buf ( \1047_b1 , \986_b1 );
not ( \1047_b1 , w_3116 );
not ( \1047_b0 , w_3117 );
and ( w_3116 , w_3117 , \986_b0 );
buf ( \1048_b1 , \1007_b1 );
not ( \1048_b1 , w_3118 );
not ( \1048_b0 , w_3119 );
and ( w_3118 , w_3119 , \1007_b0 );
or ( \1049_b1 , \1047_b1 , w_3121 );
not ( w_3121 , w_3122 );
and ( \1049_b0 , \1047_b0 , w_3123 );
and ( w_3122 ,  , w_3123 );
buf ( w_3121 , \1048_b1 );
not ( w_3121 , w_3124 );
not (  , w_3125 );
and ( w_3124 , w_3125 , \1048_b0 );
or ( \1050_b1 , \1046_b1 , w_3127 );
not ( w_3127 , w_3128 );
and ( \1050_b0 , \1046_b0 , w_3129 );
and ( w_3128 ,  , w_3129 );
buf ( w_3127 , \1049_b1 );
not ( w_3127 , w_3130 );
not (  , w_3131 );
and ( w_3130 , w_3131 , \1049_b0 );
or ( \1051_b1 , \970_b1 , \1050_b1 );
xor ( \1051_b0 , \970_b0 , w_3132 );
not ( w_3132 , w_3133 );
and ( w_3133 , \1050_b1 , \1050_b0 );
or ( \1052_b1 , \a[2]_b1 , \d[9]_b1 );
xor ( \1052_b0 , \a[2]_b0 , w_3134 );
not ( w_3134 , w_3135 );
and ( w_3135 , \d[9]_b1 , \d[9]_b0 );
buf ( \1053_b1 , \1052_b1 );
not ( \1053_b1 , w_3136 );
not ( \1053_b0 , w_3137 );
and ( w_3136 , w_3137 , \1052_b0 );
buf ( \1054_b1 , \d[7]_b1 );
not ( \1054_b1 , w_3138 );
not ( \1054_b0 , w_3139 );
and ( w_3138 , w_3139 , \d[7]_b0 );
buf ( \1055_b1 , \d[8]_b1 );
not ( \1055_b1 , w_3140 );
not ( \1055_b0 , w_3141 );
and ( w_3140 , w_3141 , \d[8]_b0 );
buf ( \1056_b1 , \1055_b1 );
not ( \1056_b1 , w_3142 );
not ( \1056_b0 , w_3143 );
and ( w_3142 , w_3143 , \1055_b0 );
or ( \1057_b1 , \1054_b1 , w_3144 );
or ( \1057_b0 , \1054_b0 , \1056_b0 );
not ( \1056_b0 , w_3145 );
and ( w_3145 , w_3144 , \1056_b1 );
or ( \1058_b1 , \1057_b1 , w_3147 );
not ( w_3147 , w_3148 );
and ( \1058_b0 , \1057_b0 , w_3149 );
and ( w_3148 ,  , w_3149 );
buf ( w_3147 , \1024_b1 );
not ( w_3147 , w_3150 );
not (  , w_3151 );
and ( w_3150 , w_3151 , \1024_b0 );
buf ( \1059_b1 , \1058_b1 );
not ( \1059_b1 , w_3152 );
not ( \1059_b0 , w_3153 );
and ( w_3152 , w_3153 , \1058_b0 );
or ( \1060_b1 , \1053_b1 , w_3154 );
or ( \1060_b0 , \1053_b0 , \1059_b0 );
not ( \1059_b0 , w_3155 );
and ( w_3155 , w_3154 , \1059_b1 );
or ( \1061_b1 , \1026_b1 , w_3157 );
not ( w_3157 , w_3158 );
and ( \1061_b0 , \1026_b0 , w_3159 );
and ( w_3158 ,  , w_3159 );
buf ( w_3157 , \1030_b1 );
not ( w_3157 , w_3160 );
not (  , w_3161 );
and ( w_3160 , w_3161 , \1030_b0 );
or ( \1062_b1 , \1060_b1 , w_3163 );
not ( w_3163 , w_3164 );
and ( \1062_b0 , \1060_b0 , w_3165 );
and ( w_3164 ,  , w_3165 );
buf ( w_3163 , \1061_b1 );
not ( w_3163 , w_3166 );
not (  , w_3167 );
and ( w_3166 , w_3167 , \1061_b0 );
buf ( \1063_b1 , \1062_b1 );
not ( \1063_b1 , w_3168 );
not ( \1063_b0 , w_3169 );
and ( w_3168 , w_3169 , \1062_b0 );
buf ( \1064_b1 , \1015_b1 );
not ( \1064_b1 , w_3170 );
not ( \1064_b0 , w_3171 );
and ( w_3170 , w_3171 , \1015_b0 );
buf ( \1065_b1 , \1011_b1 );
not ( \1065_b1 , w_3172 );
not ( \1065_b0 , w_3173 );
and ( w_3172 , w_3173 , \1011_b0 );
buf ( \1066_b1 , \1065_b1 );
not ( \1066_b1 , w_3174 );
not ( \1066_b0 , w_3175 );
and ( w_3174 , w_3175 , \1065_b0 );
or ( \1067_b1 , \1064_b1 , w_3176 );
or ( \1067_b0 , \1064_b0 , \1066_b0 );
not ( \1066_b0 , w_3177 );
and ( w_3177 , w_3176 , \1066_b1 );
or ( \1068_b1 , \a[10]_b1 , \d[1]_b1 );
xor ( \1068_b0 , \a[10]_b0 , w_3178 );
not ( w_3178 , w_3179 );
and ( w_3179 , \d[1]_b1 , \d[1]_b0 );
or ( \1069_b1 , \1068_b1 , w_3181 );
not ( w_3181 , w_3182 );
and ( \1069_b0 , \1068_b0 , w_3183 );
and ( w_3182 ,  , w_3183 );
buf ( w_3181 , \d[0]_b1 );
not ( w_3181 , w_3184 );
not (  , w_3185 );
and ( w_3184 , w_3185 , \d[0]_b0 );
or ( \1070_b1 , \1067_b1 , w_3187 );
not ( w_3187 , w_3188 );
and ( \1070_b0 , \1067_b0 , w_3189 );
and ( w_3188 ,  , w_3189 );
buf ( w_3187 , \1069_b1 );
not ( w_3187 , w_3190 );
not (  , w_3191 );
and ( w_3190 , w_3191 , \1069_b0 );
buf ( \1071_b1 , \1070_b1 );
not ( \1071_b1 , w_3192 );
not ( \1071_b0 , w_3193 );
and ( w_3192 , w_3193 , \1070_b0 );
or ( \1072_b1 , \1063_b1 , w_3194 );
or ( \1072_b0 , \1063_b0 , \1071_b0 );
not ( \1071_b0 , w_3195 );
and ( w_3195 , w_3194 , \1071_b1 );
or ( \1073_b1 , \1070_b1 , w_3196 );
or ( \1073_b0 , \1070_b0 , \1062_b0 );
not ( \1062_b0 , w_3197 );
and ( w_3197 , w_3196 , \1062_b1 );
or ( \1074_b1 , \a[5]_b1 , \d[5]_b1 );
xor ( \1074_b0 , \a[5]_b0 , w_3198 );
not ( w_3198 , w_3199 );
and ( w_3199 , \d[5]_b1 , \d[5]_b0 );
buf ( \1075_b1 , \1074_b1 );
not ( \1075_b1 , w_3200 );
not ( \1075_b0 , w_3201 );
and ( w_3200 , w_3201 , \1074_b0 );
buf ( \1076_b1 , \933_b1 );
not ( \1076_b1 , w_3202 );
not ( \1076_b0 , w_3203 );
and ( w_3202 , w_3203 , \933_b0 );
or ( \1077_b1 , \1075_b1 , w_3204 );
or ( \1077_b0 , \1075_b0 , \1076_b0 );
not ( \1076_b0 , w_3205 );
and ( w_3205 , w_3204 , \1076_b1 );
or ( \1078_b1 , \936_b1 , w_3207 );
not ( w_3207 , w_3208 );
and ( \1078_b0 , \936_b0 , w_3209 );
and ( w_3208 ,  , w_3209 );
buf ( w_3207 , \928_b1 );
not ( w_3207 , w_3210 );
not (  , w_3211 );
and ( w_3210 , w_3211 , \928_b0 );
or ( \1079_b1 , \1077_b1 , w_3213 );
not ( w_3213 , w_3214 );
and ( \1079_b0 , \1077_b0 , w_3215 );
and ( w_3214 ,  , w_3215 );
buf ( w_3213 , \1078_b1 );
not ( w_3213 , w_3216 );
not (  , w_3217 );
and ( w_3216 , w_3217 , \1078_b0 );
or ( \1080_b1 , \1073_b1 , w_3219 );
not ( w_3219 , w_3220 );
and ( \1080_b0 , \1073_b0 , w_3221 );
and ( w_3220 ,  , w_3221 );
buf ( w_3219 , \1079_b1 );
not ( w_3219 , w_3222 );
not (  , w_3223 );
and ( w_3222 , w_3223 , \1079_b0 );
or ( \1081_b1 , \1072_b1 , w_3225 );
not ( w_3225 , w_3226 );
and ( \1081_b0 , \1072_b0 , w_3227 );
and ( w_3226 ,  , w_3227 );
buf ( w_3225 , \1080_b1 );
not ( w_3225 , w_3228 );
not (  , w_3229 );
and ( w_3228 , w_3229 , \1080_b0 );
buf ( \1082_b1 , \993_b1 );
not ( \1082_b1 , w_3230 );
not ( \1082_b0 , w_3231 );
and ( w_3230 , w_3231 , \993_b0 );
or ( \1083_b1 , \1082_b1 , w_3233 );
not ( w_3233 , w_3234 );
and ( \1083_b0 , \1082_b0 , w_3235 );
and ( w_3234 ,  , w_3235 );
buf ( w_3233 , \988_b1 );
not ( w_3233 , w_3236 );
not (  , w_3237 );
and ( w_3236 , w_3237 , \988_b0 );
buf ( \1084_b1 , \1083_b1 );
not ( \1084_b1 , w_3238 );
not ( \1084_b0 , w_3239 );
and ( w_3238 , w_3239 , \1083_b0 );
buf ( \1085_b1 , \1006_b1 );
not ( \1085_b1 , w_3240 );
not ( \1085_b0 , w_3241 );
and ( w_3240 , w_3241 , \1006_b0 );
or ( \1086_b1 , \1084_b1 , w_3242 );
or ( \1086_b0 , \1084_b0 , \1085_b0 );
not ( \1085_b0 , w_3243 );
and ( w_3243 , w_3242 , \1085_b1 );
or ( \1087_b1 , \993_b1 , w_3245 );
not ( w_3245 , w_3246 );
and ( \1087_b0 , \993_b0 , w_3247 );
and ( w_3246 ,  , w_3247 );
buf ( w_3245 , \989_b1 );
not ( w_3245 , w_3248 );
not (  , w_3249 );
and ( w_3248 , w_3249 , \989_b0 );
or ( \1088_b1 , \1086_b1 , w_3251 );
not ( w_3251 , w_3252 );
and ( \1088_b0 , \1086_b0 , w_3253 );
and ( w_3252 ,  , w_3253 );
buf ( w_3251 , \1087_b1 );
not ( w_3251 , w_3254 );
not (  , w_3255 );
and ( w_3254 , w_3255 , \1087_b0 );
or ( \1089_b1 , \1081_b1 , \1088_b1 );
xor ( \1089_b0 , \1081_b0 , w_3256 );
not ( w_3256 , w_3257 );
and ( w_3257 , \1088_b1 , \1088_b0 );
buf ( \1090_b1 , \1068_b1 );
not ( \1090_b1 , w_3258 );
not ( \1090_b0 , w_3259 );
and ( w_3258 , w_3259 , \1068_b0 );
buf ( \1091_b1 , \1065_b1 );
not ( \1091_b1 , w_3260 );
not ( \1091_b0 , w_3261 );
and ( w_3260 , w_3261 , \1065_b0 );
or ( \1092_b1 , \1090_b1 , w_3262 );
or ( \1092_b0 , \1090_b0 , \1091_b0 );
not ( \1091_b0 , w_3263 );
and ( w_3263 , w_3262 , \1091_b1 );
or ( \1093_b1 , \a[11]_b1 , \d[1]_b1 );
xor ( \1093_b0 , \a[11]_b0 , w_3264 );
not ( w_3264 , w_3265 );
and ( w_3265 , \d[1]_b1 , \d[1]_b0 );
or ( \1094_b1 , \1093_b1 , w_3267 );
not ( w_3267 , w_3268 );
and ( \1094_b0 , \1093_b0 , w_3269 );
and ( w_3268 ,  , w_3269 );
buf ( w_3267 , \d[0]_b1 );
not ( w_3267 , w_3270 );
not (  , w_3271 );
and ( w_3270 , w_3271 , \d[0]_b0 );
or ( \1095_b1 , \1092_b1 , w_3273 );
not ( w_3273 , w_3274 );
and ( \1095_b0 , \1092_b0 , w_3275 );
and ( w_3274 ,  , w_3275 );
buf ( w_3273 , \1094_b1 );
not ( w_3273 , w_3276 );
not (  , w_3277 );
and ( w_3276 , w_3277 , \1094_b0 );
buf ( \1096_b1 , \1095_b1 );
not ( \1096_b1 , w_3278 );
not ( \1096_b0 , w_3279 );
and ( w_3278 , w_3279 , \1095_b0 );
buf ( \1097_b1 , \1096_b1 );
not ( \1097_b1 , w_3280 );
not ( \1097_b0 , w_3281 );
and ( w_3280 , w_3281 , \1096_b0 );
buf ( \1098_b1 , \1004_b1 );
not ( \1098_b1 , w_3282 );
not ( \1098_b0 , w_3283 );
and ( w_3282 , w_3283 , \1004_b0 );
buf ( \1099_b1 , \1038_b1 );
not ( \1099_b1 , w_3284 );
not ( \1099_b0 , w_3285 );
and ( w_3284 , w_3285 , \1038_b0 );
or ( \1100_b1 , \1098_b1 , w_3286 );
or ( \1100_b0 , \1098_b0 , \1099_b0 );
not ( \1099_b0 , w_3287 );
and ( w_3287 , w_3286 , \1099_b1 );
or ( \1101_b1 , \a[5]_b1 , \d[7]_b1 );
xor ( \1101_b0 , \a[5]_b0 , w_3288 );
not ( w_3288 , w_3289 );
and ( w_3289 , \d[7]_b1 , \d[7]_b0 );
or ( \1102_b1 , \1003_b1 , w_3291 );
not ( w_3291 , w_3292 );
and ( \1102_b0 , \1003_b0 , w_3293 );
and ( w_3292 ,  , w_3293 );
buf ( w_3291 , \1101_b1 );
not ( w_3291 , w_3294 );
not (  , w_3295 );
and ( w_3294 , w_3295 , \1101_b0 );
or ( \1103_b1 , \1100_b1 , w_3297 );
not ( w_3297 , w_3298 );
and ( \1103_b0 , \1100_b0 , w_3299 );
and ( w_3298 ,  , w_3299 );
buf ( w_3297 , \1102_b1 );
not ( w_3297 , w_3300 );
not (  , w_3301 );
and ( w_3300 , w_3301 , \1102_b0 );
buf ( \1104_b1 , \1103_b1 );
not ( \1104_b1 , w_3302 );
not ( \1104_b0 , w_3303 );
and ( w_3302 , w_3303 , \1103_b0 );
or ( \1105_b1 , \1097_b1 , w_3304 );
or ( \1105_b0 , \1097_b0 , \1104_b0 );
not ( \1104_b0 , w_3305 );
and ( w_3305 , w_3304 , \1104_b1 );
buf ( \1106_b1 , \1103_b1 );
not ( \1106_b1 , w_3306 );
not ( \1106_b0 , w_3307 );
and ( w_3306 , w_3307 , \1103_b0 );
or ( \1107_b1 , \1106_b1 , w_3309 );
not ( w_3309 , w_3310 );
and ( \1107_b0 , \1106_b0 , w_3311 );
and ( w_3310 ,  , w_3311 );
buf ( w_3309 , \1095_b1 );
not ( w_3309 , w_3312 );
not (  , w_3313 );
and ( w_3312 , w_3313 , \1095_b0 );
or ( \1108_b1 , \1105_b1 , w_3315 );
not ( w_3315 , w_3316 );
and ( \1108_b0 , \1105_b0 , w_3317 );
and ( w_3316 ,  , w_3317 );
buf ( w_3315 , \1107_b1 );
not ( w_3315 , w_3318 );
not (  , w_3319 );
and ( w_3318 , w_3319 , \1107_b0 );
buf ( \1110_b1 , \1109_b1 );
not ( \1110_b1 , w_3320 );
not ( \1110_b0 , w_3321 );
and ( w_3320 , w_3321 , \1109_b0 );
buf ( \1111_b1 , \1110_b1 );
not ( \1111_b1 , w_3322 );
not ( \1111_b0 , w_3323 );
and ( w_3322 , w_3323 , \1110_b0 );
buf ( \1112_b1 , \1052_b1 );
not ( \1112_b1 , w_3324 );
not ( \1112_b0 , w_3325 );
and ( w_3324 , w_3325 , \1052_b0 );
buf ( \1113_b1 , \1112_b1 );
not ( \1113_b1 , w_3326 );
not ( \1113_b0 , w_3327 );
and ( w_3326 , w_3327 , \1112_b0 );
or ( \1114_b1 , \1111_b1 , \1113_b1 );
not ( \1113_b1 , w_3328 );
and ( \1114_b0 , \1111_b0 , w_3329 );
and ( w_3328 , w_3329 , \1113_b0 );
or ( \1115_b1 , \a[3]_b1 , \d[9]_b1 );
xor ( \1115_b0 , \a[3]_b0 , w_3330 );
not ( w_3330 , w_3331 );
and ( w_3331 , \d[9]_b1 , \d[9]_b0 );
or ( \1116_b1 , \1058_b1 , \1115_b1 );
not ( \1115_b1 , w_3332 );
and ( \1116_b0 , \1058_b0 , w_3333 );
and ( w_3332 , w_3333 , \1115_b0 );
or ( \1117_b1 , \1114_b1 , w_3335 );
not ( w_3335 , w_3336 );
and ( \1117_b0 , \1114_b0 , w_3337 );
and ( w_3336 ,  , w_3337 );
buf ( w_3335 , \1116_b1 );
not ( w_3335 , w_3338 );
not (  , w_3339 );
and ( w_3338 , w_3339 , \1116_b0 );
buf ( \1118_b1 , \1117_b1 );
not ( \1118_b1 , w_3340 );
not ( \1118_b0 , w_3341 );
and ( w_3340 , w_3341 , \1117_b0 );
buf ( \1119_b1 , \1118_b1 );
buf ( \1119_b0 , \1118_b0 );
or ( \1120_b1 , \1108_b1 , \1119_b1 );
not ( \1119_b1 , w_3342 );
and ( \1120_b0 , \1108_b0 , w_3343 );
and ( w_3342 , w_3343 , \1119_b0 );
buf ( \1121_b1 , \1108_b1 );
not ( \1121_b1 , w_3344 );
not ( \1121_b0 , w_3345 );
and ( w_3344 , w_3345 , \1108_b0 );
buf ( \1122_b1 , \1119_b1 );
not ( \1122_b1 , w_3346 );
not ( \1122_b0 , w_3347 );
and ( w_3346 , w_3347 , \1119_b0 );
or ( \1123_b1 , \1121_b1 , \1122_b1 );
not ( \1122_b1 , w_3348 );
and ( \1123_b0 , \1121_b0 , w_3349 );
and ( w_3348 , w_3349 , \1122_b0 );
or ( \1124_b1 , \1120_b1 , w_3351 );
not ( w_3351 , w_3352 );
and ( \1124_b0 , \1120_b0 , w_3353 );
and ( w_3352 ,  , w_3353 );
buf ( w_3351 , \1123_b1 );
not ( w_3351 , w_3354 );
not (  , w_3355 );
and ( w_3354 , w_3355 , \1123_b0 );
or ( \1125_b1 , \1089_b1 , w_3356 );
xor ( \1125_b0 , \1089_b0 , w_3358 );
not ( w_3358 , w_3359 );
and ( w_3359 , w_3356 , w_3357 );
buf ( w_3356 , \1124_b1 );
not ( w_3356 , w_3360 );
not ( w_3357 , w_3361 );
and ( w_3360 , w_3361 , \1124_b0 );
or ( \1126_b1 , \1051_b1 , \1125_b1 );
xor ( \1126_b0 , \1051_b0 , w_3362 );
not ( w_3362 , w_3363 );
and ( w_3363 , \1125_b1 , \1125_b0 );
or ( \1127_b1 , \1062_b1 , \1070_b1 );
xor ( \1127_b0 , \1062_b0 , w_3364 );
not ( w_3364 , w_3365 );
and ( w_3365 , \1070_b1 , \1070_b0 );
or ( \1128_b1 , \1127_b1 , w_3366 );
xor ( \1128_b0 , \1127_b0 , w_3368 );
not ( w_3368 , w_3369 );
and ( w_3369 , w_3366 , w_3367 );
buf ( w_3366 , \1079_b1 );
not ( w_3366 , w_3370 );
not ( w_3367 , w_3371 );
and ( w_3370 , w_3371 , \1079_b0 );
or ( \1129_b1 , \a[4]_b1 , \d[5]_b1 );
xor ( \1129_b0 , \a[4]_b0 , w_3372 );
not ( w_3372 , w_3373 );
and ( w_3373 , \d[5]_b1 , \d[5]_b0 );
or ( \1130_b1 , \933_b1 , \1129_b1 );
not ( \1129_b1 , w_3374 );
and ( \1130_b0 , \933_b0 , w_3375 );
and ( w_3374 , w_3375 , \1129_b0 );
or ( \1131_b1 , \936_b1 , \1074_b1 );
not ( \1074_b1 , w_3376 );
and ( \1131_b0 , \936_b0 , w_3377 );
and ( w_3376 , w_3377 , \1074_b0 );
or ( \1132_b1 , \1130_b1 , w_3379 );
not ( w_3379 , w_3380 );
and ( \1132_b0 , \1130_b0 , w_3381 );
and ( w_3380 ,  , w_3381 );
buf ( w_3379 , \1131_b1 );
not ( w_3379 , w_3382 );
not (  , w_3383 );
and ( w_3382 , w_3383 , \1131_b0 );
buf ( \1133_b1 , \985_b1 );
not ( \1133_b1 , w_3384 );
not ( \1133_b0 , w_3385 );
and ( w_3384 , w_3385 , \985_b0 );
buf ( \1134_b1 , \974_b1 );
not ( \1134_b1 , w_3386 );
not ( \1134_b0 , w_3387 );
and ( w_3386 , w_3387 , \974_b0 );
or ( \1135_b1 , \1133_b1 , \1134_b1 );
not ( \1134_b1 , w_3388 );
and ( \1135_b0 , \1133_b0 , w_3389 );
and ( w_3388 , w_3389 , \1134_b0 );
or ( \1136_b1 , \985_b1 , \974_b1 );
not ( \974_b1 , w_3390 );
and ( \1136_b0 , \985_b0 , w_3391 );
and ( w_3390 , w_3391 , \974_b0 );
or ( \1137_b1 , \1135_b1 , w_3393 );
not ( w_3393 , w_3394 );
and ( \1137_b0 , \1135_b0 , w_3395 );
and ( w_3394 ,  , w_3395 );
buf ( w_3393 , \1136_b1 );
not ( w_3393 , w_3396 );
not (  , w_3397 );
and ( w_3396 , w_3397 , \1136_b0 );
or ( \1138_b1 , \1132_b1 , \1137_b1 );
xor ( \1138_b0 , \1132_b0 , w_3398 );
not ( w_3398 , w_3399 );
and ( w_3399 , \1137_b1 , \1137_b0 );
or ( \1139_b1 , \1029_b1 , w_3401 );
not ( w_3401 , w_3402 );
and ( \1139_b0 , \1029_b0 , w_3403 );
and ( w_3402 ,  , w_3403 );
buf ( w_3401 , \a[0]_b1 );
not ( w_3401 , w_3404 );
not (  , w_3405 );
and ( w_3404 , w_3405 , \a[0]_b0 );
or ( \1140_b1 , \d[1]_b1 , \a[7]_b1 );
xor ( \1140_b0 , \d[1]_b0 , w_3406 );
not ( w_3406 , w_3407 );
and ( w_3407 , \a[7]_b1 , \a[7]_b0 );
or ( \1141_b1 , \1012_b1 , \1140_b1 );
not ( \1140_b1 , w_3408 );
and ( \1141_b0 , \1012_b0 , w_3409 );
and ( w_3408 , w_3409 , \1140_b0 );
or ( \1142_b1 , \1013_b1 , \d[0]_b1 );
not ( \d[0]_b1 , w_3410 );
and ( \1142_b0 , \1013_b0 , w_3411 );
and ( w_3410 , w_3411 , \d[0]_b0 );
or ( \1143_b1 , \1141_b1 , w_3413 );
not ( w_3413 , w_3414 );
and ( \1143_b0 , \1141_b0 , w_3415 );
and ( w_3414 ,  , w_3415 );
buf ( w_3413 , \1142_b1 );
not ( w_3413 , w_3416 );
not (  , w_3417 );
and ( w_3416 , w_3417 , \1142_b0 );
or ( \1144_b1 , \1139_b1 , \1143_b1 );
xor ( \1144_b0 , \1139_b0 , w_3418 );
not ( w_3418 , w_3419 );
and ( w_3419 , \1143_b1 , \1143_b0 );
or ( \1145_b1 , \a[1]_b1 , \d[7]_b1 );
xor ( \1145_b0 , \a[1]_b0 , w_3420 );
not ( w_3420 , w_3421 );
and ( w_3421 , \d[7]_b1 , \d[7]_b0 );
or ( \1146_b1 , \1038_b1 , \1145_b1 );
not ( \1145_b1 , w_3422 );
and ( \1146_b0 , \1038_b0 , w_3423 );
and ( w_3422 , w_3423 , \1145_b0 );
or ( \1147_b1 , \1003_b1 , \1036_b1 );
not ( \1036_b1 , w_3424 );
and ( \1147_b0 , \1003_b0 , w_3425 );
and ( w_3424 , w_3425 , \1036_b0 );
or ( \1148_b1 , \1146_b1 , w_3427 );
not ( w_3427 , w_3428 );
and ( \1148_b0 , \1146_b0 , w_3429 );
and ( w_3428 ,  , w_3429 );
buf ( w_3427 , \1147_b1 );
not ( w_3427 , w_3430 );
not (  , w_3431 );
and ( w_3430 , w_3431 , \1147_b0 );
or ( \1149_b1 , \1144_b1 , \1148_b1 );
not ( \1148_b1 , w_3432 );
and ( \1149_b0 , \1144_b0 , w_3433 );
and ( w_3432 , w_3433 , \1148_b0 );
or ( \1150_b1 , \1139_b1 , \1143_b1 );
not ( \1143_b1 , w_3434 );
and ( \1150_b0 , \1139_b0 , w_3435 );
and ( w_3434 , w_3435 , \1143_b0 );
or ( \1151_b1 , \1149_b1 , w_3436 );
or ( \1151_b0 , \1149_b0 , \1150_b0 );
not ( \1150_b0 , w_3437 );
and ( w_3437 , w_3436 , \1150_b1 );
or ( \1152_b1 , \1138_b1 , \1151_b1 );
not ( \1151_b1 , w_3438 );
and ( \1152_b0 , \1138_b0 , w_3439 );
and ( w_3438 , w_3439 , \1151_b0 );
or ( \1153_b1 , \1132_b1 , \1137_b1 );
not ( \1137_b1 , w_3440 );
and ( \1153_b0 , \1132_b0 , w_3441 );
and ( w_3440 , w_3441 , \1137_b0 );
or ( \1154_b1 , \1152_b1 , w_3442 );
or ( \1154_b0 , \1152_b0 , \1153_b0 );
not ( \1153_b0 , w_3443 );
and ( w_3443 , w_3442 , \1153_b1 );
or ( \1155_b1 , \1128_b1 , \1154_b1 );
xor ( \1155_b0 , \1128_b0 , w_3444 );
not ( w_3444 , w_3445 );
and ( w_3445 , \1154_b1 , \1154_b0 );
or ( \1156_b1 , \986_b1 , \1045_b1 );
xor ( \1156_b0 , \986_b0 , w_3446 );
not ( w_3446 , w_3447 );
and ( w_3447 , \1045_b1 , \1045_b0 );
or ( \1157_b1 , \1156_b1 , \1048_b1 );
xor ( \1157_b0 , \1156_b0 , w_3448 );
not ( w_3448 , w_3449 );
and ( w_3449 , \1048_b1 , \1048_b0 );
or ( \1158_b1 , \1155_b1 , \1157_b1 );
not ( \1157_b1 , w_3450 );
and ( \1158_b0 , \1155_b0 , w_3451 );
and ( w_3450 , w_3451 , \1157_b0 );
or ( \1159_b1 , \1128_b1 , \1154_b1 );
not ( \1154_b1 , w_3452 );
and ( \1159_b0 , \1128_b0 , w_3453 );
and ( w_3452 , w_3453 , \1154_b0 );
or ( \1160_b1 , \1158_b1 , w_3454 );
or ( \1160_b0 , \1158_b0 , \1159_b0 );
not ( \1159_b0 , w_3455 );
and ( w_3455 , w_3454 , \1159_b1 );
or ( \1161_b1 , \1126_b1 , w_3457 );
not ( w_3457 , w_3458 );
and ( \1161_b0 , \1126_b0 , w_3459 );
and ( w_3458 ,  , w_3459 );
buf ( w_3457 , \1160_b1 );
not ( w_3457 , w_3460 );
not (  , w_3461 );
and ( w_3460 , w_3461 , \1160_b0 );
or ( \1162_b1 , \1128_b1 , \1154_b1 );
xor ( \1162_b0 , \1128_b0 , w_3462 );
not ( w_3462 , w_3463 );
and ( w_3463 , \1154_b1 , \1154_b0 );
or ( \1163_b1 , \1162_b1 , \1157_b1 );
xor ( \1163_b0 , \1162_b0 , w_3464 );
not ( w_3464 , w_3465 );
and ( w_3465 , \1157_b1 , \1157_b0 );
buf ( \1164_b1 , \1017_b1 );
not ( \1164_b1 , w_3466 );
not ( \1164_b0 , w_3467 );
and ( w_3466 , w_3467 , \1017_b0 );
buf ( \1165_b1 , \1043_b1 );
not ( \1165_b1 , w_3468 );
not ( \1165_b0 , w_3469 );
and ( w_3468 , w_3469 , \1043_b0 );
or ( \1166_b1 , \1164_b1 , w_3470 );
or ( \1166_b0 , \1164_b0 , \1165_b0 );
not ( \1165_b0 , w_3471 );
and ( w_3471 , w_3470 , \1165_b1 );
buf ( \1167_b1 , \1043_b1 );
not ( \1167_b1 , w_3472 );
not ( \1167_b0 , w_3473 );
and ( w_3472 , w_3473 , \1043_b0 );
or ( \1168_b1 , \1167_b1 , w_3475 );
not ( w_3475 , w_3476 );
and ( \1168_b0 , \1167_b0 , w_3477 );
and ( w_3476 ,  , w_3477 );
buf ( w_3475 , \1018_b1 );
not ( w_3475 , w_3478 );
not (  , w_3479 );
and ( w_3478 , w_3479 , \1018_b0 );
or ( \1169_b1 , \1166_b1 , w_3481 );
not ( w_3481 , w_3482 );
and ( \1169_b0 , \1166_b0 , w_3483 );
and ( w_3482 ,  , w_3483 );
buf ( w_3481 , \1168_b1 );
not ( w_3481 , w_3484 );
not (  , w_3485 );
and ( w_3484 , w_3485 , \1168_b0 );
or ( \1170_b1 , \1169_b1 , \1032_b1 );
xor ( \1170_b0 , \1169_b0 , w_3486 );
not ( w_3486 , w_3487 );
and ( w_3487 , \1032_b1 , \1032_b0 );
buf ( \1171_b1 , \1170_b1 );
not ( \1171_b1 , w_3488 );
not ( \1171_b0 , w_3489 );
and ( w_3488 , w_3489 , \1170_b0 );
buf ( \1172_b1 , \1012_b1 );
not ( \1172_b1 , w_3490 );
not ( \1172_b0 , w_3491 );
and ( w_3490 , w_3491 , \1012_b0 );
or ( \1173_b1 , \d[1]_b1 , \a[6]_b1 );
xor ( \1173_b0 , \d[1]_b0 , w_3492 );
not ( w_3492 , w_3493 );
and ( w_3493 , \a[6]_b1 , \a[6]_b0 );
buf ( \1174_b1 , \1173_b1 );
not ( \1174_b1 , w_3494 );
not ( \1174_b0 , w_3495 );
and ( w_3494 , w_3495 , \1173_b0 );
or ( \1175_b1 , \1172_b1 , w_3496 );
or ( \1175_b0 , \1172_b0 , \1174_b0 );
not ( \1174_b0 , w_3497 );
and ( w_3497 , w_3496 , \1174_b1 );
or ( \1176_b1 , \1140_b1 , w_3499 );
not ( w_3499 , w_3500 );
and ( \1176_b0 , \1140_b0 , w_3501 );
and ( w_3500 ,  , w_3501 );
buf ( w_3499 , \d[0]_b1 );
not ( w_3499 , w_3502 );
not (  , w_3503 );
and ( w_3502 , w_3503 , \d[0]_b0 );
or ( \1177_b1 , \1175_b1 , w_3505 );
not ( w_3505 , w_3506 );
and ( \1177_b0 , \1175_b0 , w_3507 );
and ( w_3506 ,  , w_3507 );
buf ( w_3505 , \1176_b1 );
not ( w_3505 , w_3508 );
not (  , w_3509 );
and ( w_3508 , w_3509 , \1176_b0 );
or ( \1178_b1 , \a[0]_b1 , w_3510 );
or ( \1178_b0 , \a[0]_b0 , \d[6]_b0 );
not ( \d[6]_b0 , w_3511 );
and ( w_3511 , w_3510 , \d[6]_b1 );
or ( \1179_b1 , \1178_b1 , w_3513 );
not ( w_3513 , w_3514 );
and ( \1179_b0 , \1178_b0 , w_3515 );
and ( w_3514 ,  , w_3515 );
buf ( w_3513 , \d[5]_b1 );
not ( w_3513 , w_3516 );
not (  , w_3517 );
and ( w_3516 , w_3517 , \d[5]_b0 );
or ( \1180_b1 , \a[0]_b1 , w_3519 );
not ( w_3519 , w_3520 );
and ( \1180_b0 , \a[0]_b0 , w_3521 );
and ( w_3520 ,  , w_3521 );
buf ( w_3519 , \d[6]_b1 );
not ( w_3519 , w_3522 );
not (  , w_3523 );
and ( w_3522 , w_3523 , \d[6]_b0 );
or ( \1182_b1 , \1177_b1 , w_3525 );
not ( w_3525 , w_3526 );
and ( \1182_b0 , \1177_b0 , w_3527 );
and ( w_3526 ,  , w_3527 );
buf ( w_3525 , \1181_b1 );
not ( w_3525 , w_3528 );
not (  , w_3529 );
and ( w_3528 , w_3529 , \1181_b0 );
or ( \1183_b1 , \a[3]_b1 , \d[5]_b1 );
xor ( \1183_b0 , \a[3]_b0 , w_3530 );
not ( w_3530 , w_3531 );
and ( w_3531 , \d[5]_b1 , \d[5]_b0 );
buf ( \1184_b1 , \1183_b1 );
not ( \1184_b1 , w_3532 );
not ( \1184_b0 , w_3533 );
and ( w_3532 , w_3533 , \1183_b0 );
buf ( \1185_b1 , \930_b1 );
not ( \1185_b1 , w_3534 );
not ( \1185_b0 , w_3535 );
and ( w_3534 , w_3535 , \930_b0 );
or ( \1186_b1 , \1185_b1 , w_3537 );
not ( w_3537 , w_3538 );
and ( \1186_b0 , \1185_b0 , w_3539 );
and ( w_3538 ,  , w_3539 );
buf ( w_3537 , \932_b1 );
not ( w_3537 , w_3540 );
not (  , w_3541 );
and ( w_3540 , w_3541 , \932_b0 );
buf ( \1187_b1 , \1186_b1 );
not ( \1187_b1 , w_3542 );
not ( \1187_b0 , w_3543 );
and ( w_3542 , w_3543 , \1186_b0 );
or ( \1188_b1 , \1184_b1 , w_3544 );
or ( \1188_b0 , \1184_b0 , \1187_b0 );
not ( \1187_b0 , w_3545 );
and ( w_3545 , w_3544 , \1187_b1 );
or ( \1189_b1 , \936_b1 , w_3547 );
not ( w_3547 , w_3548 );
and ( \1189_b0 , \936_b0 , w_3549 );
and ( w_3548 ,  , w_3549 );
buf ( w_3547 , \1129_b1 );
not ( w_3547 , w_3550 );
not (  , w_3551 );
and ( w_3550 , w_3551 , \1129_b0 );
or ( \1190_b1 , \1188_b1 , w_3553 );
not ( w_3553 , w_3554 );
and ( \1190_b0 , \1188_b0 , w_3555 );
and ( w_3554 ,  , w_3555 );
buf ( w_3553 , \1189_b1 );
not ( w_3553 , w_3556 );
not (  , w_3557 );
and ( w_3556 , w_3557 , \1189_b0 );
buf ( \1191_b1 , \1190_b1 );
not ( \1191_b1 , w_3558 );
not ( \1191_b0 , w_3559 );
and ( w_3558 , w_3559 , \1190_b0 );
or ( \1192_b1 , \1182_b1 , w_3561 );
not ( w_3561 , w_3562 );
and ( \1192_b0 , \1182_b0 , w_3563 );
and ( w_3562 ,  , w_3563 );
buf ( w_3561 , \1191_b1 );
not ( w_3561 , w_3564 );
not (  , w_3565 );
and ( w_3564 , w_3565 , \1191_b0 );
or ( \1193_b1 , \a[5]_b1 , \d[3]_b1 );
xor ( \1193_b0 , \a[5]_b0 , w_3566 );
not ( w_3566 , w_3567 );
and ( w_3567 , \d[3]_b1 , \d[3]_b0 );
buf ( \1194_b1 , \1193_b1 );
not ( \1194_b1 , w_3568 );
not ( \1194_b0 , w_3569 );
and ( w_3568 , w_3569 , \1193_b0 );
buf ( \1195_b1 , \962_b1 );
not ( \1195_b1 , w_3570 );
not ( \1195_b0 , w_3571 );
and ( w_3570 , w_3571 , \962_b0 );
or ( \1196_b1 , \1194_b1 , w_3572 );
or ( \1196_b0 , \1194_b0 , \1195_b0 );
not ( \1195_b0 , w_3573 );
and ( w_3573 , w_3572 , \1195_b1 );
or ( \1197_b1 , \965_b1 , w_3575 );
not ( w_3575 , w_3576 );
and ( \1197_b0 , \965_b0 , w_3577 );
and ( w_3576 ,  , w_3577 );
buf ( w_3575 , \976_b1 );
not ( w_3575 , w_3578 );
not (  , w_3579 );
and ( w_3578 , w_3579 , \976_b0 );
or ( \1198_b1 , \1196_b1 , w_3581 );
not ( w_3581 , w_3582 );
and ( \1198_b0 , \1196_b0 , w_3583 );
and ( w_3582 ,  , w_3583 );
buf ( w_3581 , \1197_b1 );
not ( w_3581 , w_3584 );
not (  , w_3585 );
and ( w_3584 , w_3585 , \1197_b0 );
or ( \1199_b1 , \1192_b1 , \1198_b1 );
not ( \1198_b1 , w_3586 );
and ( \1199_b0 , \1192_b0 , w_3587 );
and ( w_3586 , w_3587 , \1198_b0 );
buf ( \1200_b1 , \1182_b1 );
not ( \1200_b1 , w_3588 );
not ( \1200_b0 , w_3589 );
and ( w_3588 , w_3589 , \1182_b0 );
or ( \1201_b1 , \1200_b1 , \1190_b1 );
not ( \1190_b1 , w_3590 );
and ( \1201_b0 , \1200_b0 , w_3591 );
and ( w_3590 , w_3591 , \1190_b0 );
or ( \1202_b1 , \1199_b1 , w_3593 );
not ( w_3593 , w_3594 );
and ( \1202_b0 , \1199_b0 , w_3595 );
and ( w_3594 ,  , w_3595 );
buf ( w_3593 , \1201_b1 );
not ( w_3593 , w_3596 );
not (  , w_3597 );
and ( w_3596 , w_3597 , \1201_b0 );
or ( \1203_b1 , \1171_b1 , w_3599 );
not ( w_3599 , w_3600 );
and ( \1203_b0 , \1171_b0 , w_3601 );
and ( w_3600 ,  , w_3601 );
buf ( w_3599 , \1202_b1 );
not ( w_3599 , w_3602 );
not (  , w_3603 );
and ( w_3602 , w_3603 , \1202_b0 );
buf ( \1204_b1 , \1203_b1 );
not ( \1204_b1 , w_3604 );
not ( \1204_b0 , w_3605 );
and ( w_3604 , w_3605 , \1203_b0 );
or ( \1205_b1 , \1132_b1 , \1137_b1 );
xor ( \1205_b0 , \1132_b0 , w_3606 );
not ( w_3606 , w_3607 );
and ( w_3607 , \1137_b1 , \1137_b0 );
or ( \1206_b1 , \1205_b1 , \1151_b1 );
xor ( \1206_b0 , \1205_b0 , w_3608 );
not ( w_3608 , w_3609 );
and ( w_3609 , \1151_b1 , \1151_b0 );
buf ( \1207_b1 , \1206_b1 );
not ( \1207_b1 , w_3610 );
not ( \1207_b0 , w_3611 );
and ( w_3610 , w_3611 , \1206_b0 );
buf ( \1208_b1 , \1207_b1 );
not ( \1208_b1 , w_3612 );
not ( \1208_b0 , w_3613 );
and ( w_3612 , w_3613 , \1207_b0 );
or ( \1209_b1 , \1204_b1 , w_3614 );
or ( \1209_b0 , \1204_b0 , \1208_b0 );
not ( \1208_b0 , w_3615 );
and ( w_3615 , w_3614 , \1208_b1 );
buf ( \1210_b1 , \1202_b1 );
not ( \1210_b1 , w_3616 );
not ( \1210_b0 , w_3617 );
and ( w_3616 , w_3617 , \1202_b0 );
or ( \1211_b1 , \1210_b1 , w_3619 );
not ( w_3619 , w_3620 );
and ( \1211_b0 , \1210_b0 , w_3621 );
and ( w_3620 ,  , w_3621 );
buf ( w_3619 , \1170_b1 );
not ( w_3619 , w_3622 );
not (  , w_3623 );
and ( w_3622 , w_3623 , \1170_b0 );
or ( \1212_b1 , \1209_b1 , w_3625 );
not ( w_3625 , w_3626 );
and ( \1212_b0 , \1209_b0 , w_3627 );
and ( w_3626 ,  , w_3627 );
buf ( w_3625 , \1211_b1 );
not ( w_3625 , w_3628 );
not (  , w_3629 );
and ( w_3628 , w_3629 , \1211_b0 );
buf ( \1213_b1 , \1212_b1 );
not ( \1213_b1 , w_3630 );
not ( \1213_b0 , w_3631 );
and ( w_3630 , w_3631 , \1212_b0 );
or ( \1214_b1 , \1163_b1 , w_3633 );
not ( w_3633 , w_3634 );
and ( \1214_b0 , \1163_b0 , w_3635 );
and ( w_3634 ,  , w_3635 );
buf ( w_3633 , \1213_b1 );
not ( w_3633 , w_3636 );
not (  , w_3637 );
and ( w_3636 , w_3637 , \1213_b0 );
or ( \1215_b1 , \1139_b1 , \1143_b1 );
xor ( \1215_b0 , \1139_b0 , w_3638 );
not ( w_3638 , w_3639 );
and ( w_3639 , \1143_b1 , \1143_b0 );
or ( \1216_b1 , \1215_b1 , \1148_b1 );
xor ( \1216_b0 , \1215_b0 , w_3640 );
not ( w_3640 , w_3641 );
and ( w_3641 , \1148_b1 , \1148_b0 );
buf ( \1217_b1 , \1216_b1 );
not ( \1217_b1 , w_3642 );
not ( \1217_b0 , w_3643 );
and ( w_3642 , w_3643 , \1216_b0 );
buf ( \1218_b1 , \1217_b1 );
not ( \1218_b1 , w_3644 );
not ( \1218_b0 , w_3645 );
and ( w_3644 , w_3645 , \1217_b0 );
or ( \1219_b1 , \a[4]_b1 , \d[3]_b1 );
xor ( \1219_b0 , \a[4]_b0 , w_3646 );
not ( w_3646 , w_3647 );
and ( w_3647 , \d[3]_b1 , \d[3]_b0 );
buf ( \1220_b1 , \1219_b1 );
not ( \1220_b1 , w_3648 );
not ( \1220_b0 , w_3649 );
and ( w_3648 , w_3649 , \1219_b0 );
buf ( \1221_b1 , \962_b1 );
not ( \1221_b1 , w_3650 );
not ( \1221_b0 , w_3651 );
and ( w_3650 , w_3651 , \962_b0 );
or ( \1222_b1 , \1220_b1 , w_3652 );
or ( \1222_b0 , \1220_b0 , \1221_b0 );
not ( \1221_b0 , w_3653 );
and ( w_3653 , w_3652 , \1221_b1 );
or ( \1223_b1 , \965_b1 , w_3655 );
not ( w_3655 , w_3656 );
and ( \1223_b0 , \965_b0 , w_3657 );
and ( w_3656 ,  , w_3657 );
buf ( w_3655 , \1193_b1 );
not ( w_3655 , w_3658 );
not (  , w_3659 );
and ( w_3658 , w_3659 , \1193_b0 );
or ( \1224_b1 , \1222_b1 , w_3661 );
not ( w_3661 , w_3662 );
and ( \1224_b0 , \1222_b0 , w_3663 );
and ( w_3662 ,  , w_3663 );
buf ( w_3661 , \1223_b1 );
not ( w_3661 , w_3664 );
not (  , w_3665 );
and ( w_3664 , w_3665 , \1223_b0 );
or ( \1225_b1 , \a[2]_b1 , \d[5]_b1 );
xor ( \1225_b0 , \a[2]_b0 , w_3666 );
not ( w_3666 , w_3667 );
and ( w_3667 , \d[5]_b1 , \d[5]_b0 );
buf ( \1226_b1 , \1225_b1 );
not ( \1226_b1 , w_3668 );
not ( \1226_b0 , w_3669 );
and ( w_3668 , w_3669 , \1225_b0 );
buf ( \1227_b1 , \1186_b1 );
not ( \1227_b1 , w_3670 );
not ( \1227_b0 , w_3671 );
and ( w_3670 , w_3671 , \1186_b0 );
or ( \1228_b1 , \1226_b1 , w_3672 );
or ( \1228_b0 , \1226_b0 , \1227_b0 );
not ( \1227_b0 , w_3673 );
and ( w_3673 , w_3672 , \1227_b1 );
or ( \1229_b1 , \936_b1 , w_3675 );
not ( w_3675 , w_3676 );
and ( \1229_b0 , \936_b0 , w_3677 );
and ( w_3676 ,  , w_3677 );
buf ( w_3675 , \1183_b1 );
not ( w_3675 , w_3678 );
not (  , w_3679 );
and ( w_3678 , w_3679 , \1183_b0 );
or ( \1230_b1 , \1228_b1 , w_3681 );
not ( w_3681 , w_3682 );
and ( \1230_b0 , \1228_b0 , w_3683 );
and ( w_3682 ,  , w_3683 );
buf ( w_3681 , \1229_b1 );
not ( w_3681 , w_3684 );
not (  , w_3685 );
and ( w_3684 , w_3685 , \1229_b0 );
or ( \1231_b1 , \1224_b1 , w_3686 );
or ( \1231_b0 , \1224_b0 , \1230_b0 );
not ( \1230_b0 , w_3687 );
and ( w_3687 , w_3686 , \1230_b1 );
or ( \1232_b1 , \a[0]_b1 , \d[7]_b1 );
xor ( \1232_b0 , \a[0]_b0 , w_3688 );
not ( w_3688 , w_3689 );
and ( w_3689 , \d[7]_b1 , \d[7]_b0 );
buf ( \1233_b1 , \1232_b1 );
not ( \1233_b1 , w_3690 );
not ( \1233_b0 , w_3691 );
and ( w_3690 , w_3691 , \1232_b0 );
buf ( \1234_b1 , \999_b1 );
not ( \1234_b1 , w_3692 );
not ( \1234_b0 , w_3693 );
and ( w_3692 , w_3693 , \999_b0 );
or ( \1235_b1 , \1233_b1 , w_3694 );
or ( \1235_b0 , \1233_b0 , \1234_b0 );
not ( \1234_b0 , w_3695 );
and ( w_3695 , w_3694 , \1234_b1 );
or ( \1236_b1 , \1003_b1 , w_3697 );
not ( w_3697 , w_3698 );
and ( \1236_b0 , \1003_b0 , w_3699 );
and ( w_3698 ,  , w_3699 );
buf ( w_3697 , \1145_b1 );
not ( w_3697 , w_3700 );
not (  , w_3701 );
and ( w_3700 , w_3701 , \1145_b0 );
or ( \1237_b1 , \1235_b1 , w_3703 );
not ( w_3703 , w_3704 );
and ( \1237_b0 , \1235_b0 , w_3705 );
and ( w_3704 ,  , w_3705 );
buf ( w_3703 , \1236_b1 );
not ( w_3703 , w_3706 );
not (  , w_3707 );
and ( w_3706 , w_3707 , \1236_b0 );
or ( \1238_b1 , \1231_b1 , w_3709 );
not ( w_3709 , w_3710 );
and ( \1238_b0 , \1231_b0 , w_3711 );
and ( w_3710 ,  , w_3711 );
buf ( w_3709 , \1237_b1 );
not ( w_3709 , w_3712 );
not (  , w_3713 );
and ( w_3712 , w_3713 , \1237_b0 );
or ( \1239_b1 , \1224_b1 , w_3715 );
not ( w_3715 , w_3716 );
and ( \1239_b0 , \1224_b0 , w_3717 );
and ( w_3716 ,  , w_3717 );
buf ( w_3715 , \1230_b1 );
not ( w_3715 , w_3718 );
not (  , w_3719 );
and ( w_3718 , w_3719 , \1230_b0 );
or ( \1240_b1 , \1238_b1 , w_3721 );
not ( w_3721 , w_3722 );
and ( \1240_b0 , \1238_b0 , w_3723 );
and ( w_3722 ,  , w_3723 );
buf ( w_3721 , \1239_b1 );
not ( w_3721 , w_3724 );
not (  , w_3725 );
and ( w_3724 , w_3725 , \1239_b0 );
buf ( \1241_b1 , \1240_b1 );
not ( \1241_b1 , w_3726 );
not ( \1241_b0 , w_3727 );
and ( w_3726 , w_3727 , \1240_b0 );
buf ( \1242_b1 , \1241_b1 );
not ( \1242_b1 , w_3728 );
not ( \1242_b0 , w_3729 );
and ( w_3728 , w_3729 , \1241_b0 );
or ( \1243_b1 , \1218_b1 , w_3730 );
or ( \1243_b0 , \1218_b0 , \1242_b0 );
not ( \1242_b0 , w_3731 );
and ( w_3731 , w_3730 , \1242_b1 );
or ( \1244_b1 , \1240_b1 , w_3733 );
not ( w_3733 , w_3734 );
and ( \1244_b0 , \1240_b0 , w_3735 );
and ( w_3734 ,  , w_3735 );
buf ( w_3733 , \1216_b1 );
not ( w_3733 , w_3736 );
not (  , w_3737 );
and ( w_3736 , w_3737 , \1216_b0 );
or ( \1245_b1 , \1243_b1 , w_3739 );
not ( w_3739 , w_3740 );
and ( \1245_b0 , \1243_b0 , w_3741 );
and ( w_3740 ,  , w_3741 );
buf ( w_3739 , \1244_b1 );
not ( w_3739 , w_3742 );
not (  , w_3743 );
and ( w_3742 , w_3743 , \1244_b0 );
buf ( \1246_b1 , \1191_b1 );
not ( \1246_b1 , w_3744 );
not ( \1246_b0 , w_3745 );
and ( w_3744 , w_3745 , \1191_b0 );
buf ( \1247_b1 , \1200_b1 );
not ( \1247_b1 , w_3746 );
not ( \1247_b0 , w_3747 );
and ( w_3746 , w_3747 , \1200_b0 );
or ( \1248_b1 , \1246_b1 , w_3748 );
or ( \1248_b0 , \1246_b0 , \1247_b0 );
not ( \1247_b0 , w_3749 );
and ( w_3749 , w_3748 , \1247_b1 );
or ( \1249_b1 , \1200_b1 , w_3750 );
or ( \1249_b0 , \1200_b0 , \1191_b0 );
not ( \1191_b0 , w_3751 );
and ( w_3751 , w_3750 , \1191_b1 );
or ( \1250_b1 , \1248_b1 , w_3753 );
not ( w_3753 , w_3754 );
and ( \1250_b0 , \1248_b0 , w_3755 );
and ( w_3754 ,  , w_3755 );
buf ( w_3753 , \1249_b1 );
not ( w_3753 , w_3756 );
not (  , w_3757 );
and ( w_3756 , w_3757 , \1249_b0 );
buf ( \1251_b1 , \1198_b1 );
not ( \1251_b1 , w_3758 );
not ( \1251_b0 , w_3759 );
and ( w_3758 , w_3759 , \1198_b0 );
or ( \1252_b1 , \1250_b1 , \1251_b1 );
not ( \1251_b1 , w_3760 );
and ( \1252_b0 , \1250_b0 , w_3761 );
and ( w_3760 , w_3761 , \1251_b0 );
buf ( \1253_b1 , \1250_b1 );
not ( \1253_b1 , w_3762 );
not ( \1253_b0 , w_3763 );
and ( w_3762 , w_3763 , \1250_b0 );
or ( \1254_b1 , \1253_b1 , \1198_b1 );
not ( \1198_b1 , w_3764 );
and ( \1254_b0 , \1253_b0 , w_3765 );
and ( w_3764 , w_3765 , \1198_b0 );
or ( \1255_b1 , \1252_b1 , w_3767 );
not ( w_3767 , w_3768 );
and ( \1255_b0 , \1252_b0 , w_3769 );
and ( w_3768 ,  , w_3769 );
buf ( w_3767 , \1254_b1 );
not ( w_3767 , w_3770 );
not (  , w_3771 );
and ( w_3770 , w_3771 , \1254_b0 );
or ( \1256_b1 , \1245_b1 , \1255_b1 );
not ( \1255_b1 , w_3772 );
and ( \1256_b0 , \1245_b0 , w_3773 );
and ( w_3772 , w_3773 , \1255_b0 );
buf ( \1257_b1 , \1245_b1 );
not ( \1257_b1 , w_3774 );
not ( \1257_b0 , w_3775 );
and ( w_3774 , w_3775 , \1245_b0 );
buf ( \1258_b1 , \1255_b1 );
not ( \1258_b1 , w_3776 );
not ( \1258_b0 , w_3777 );
and ( w_3776 , w_3777 , \1255_b0 );
or ( \1259_b1 , \1257_b1 , \1258_b1 );
not ( \1258_b1 , w_3778 );
and ( \1259_b0 , \1257_b0 , w_3779 );
and ( w_3778 , w_3779 , \1258_b0 );
or ( \1260_b1 , \1256_b1 , w_3781 );
not ( w_3781 , w_3782 );
and ( \1260_b0 , \1256_b0 , w_3783 );
and ( w_3782 ,  , w_3783 );
buf ( w_3781 , \1259_b1 );
not ( w_3781 , w_3784 );
not (  , w_3785 );
and ( w_3784 , w_3785 , \1259_b0 );
or ( \1261_b1 , \1177_b1 , w_3786 );
xor ( \1261_b0 , \1177_b0 , w_3788 );
not ( w_3788 , w_3789 );
and ( w_3789 , w_3786 , w_3787 );
buf ( w_3786 , \1181_b1 );
not ( w_3786 , w_3790 );
not ( w_3787 , w_3791 );
and ( w_3790 , w_3791 , \1181_b0 );
or ( \1262_b1 , \a[3]_b1 , \d[3]_b1 );
xor ( \1262_b0 , \a[3]_b0 , w_3792 );
not ( w_3792 , w_3793 );
and ( w_3793 , \d[3]_b1 , \d[3]_b0 );
buf ( \1263_b1 , \1262_b1 );
not ( \1263_b1 , w_3794 );
not ( \1263_b0 , w_3795 );
and ( w_3794 , w_3795 , \1262_b0 );
buf ( \1264_b1 , \962_b1 );
not ( \1264_b1 , w_3796 );
not ( \1264_b0 , w_3797 );
and ( w_3796 , w_3797 , \962_b0 );
or ( \1265_b1 , \1263_b1 , w_3798 );
or ( \1265_b0 , \1263_b0 , \1264_b0 );
not ( \1264_b0 , w_3799 );
and ( w_3799 , w_3798 , \1264_b1 );
or ( \1266_b1 , \965_b1 , w_3801 );
not ( w_3801 , w_3802 );
and ( \1266_b0 , \965_b0 , w_3803 );
and ( w_3802 ,  , w_3803 );
buf ( w_3801 , \1219_b1 );
not ( w_3801 , w_3804 );
not (  , w_3805 );
and ( w_3804 , w_3805 , \1219_b0 );
or ( \1267_b1 , \1265_b1 , w_3807 );
not ( w_3807 , w_3808 );
and ( \1267_b0 , \1265_b0 , w_3809 );
and ( w_3808 ,  , w_3809 );
buf ( w_3807 , \1266_b1 );
not ( w_3807 , w_3810 );
not (  , w_3811 );
and ( w_3810 , w_3811 , \1266_b0 );
or ( \1268_b1 , \a[5]_b1 , \d[1]_b1 );
xor ( \1268_b0 , \a[5]_b0 , w_3812 );
not ( w_3812 , w_3813 );
and ( w_3813 , \d[1]_b1 , \d[1]_b0 );
buf ( \1269_b1 , \1268_b1 );
not ( \1269_b1 , w_3814 );
not ( \1269_b0 , w_3815 );
and ( w_3814 , w_3815 , \1268_b0 );
buf ( \1270_b1 , \1065_b1 );
not ( \1270_b1 , w_3816 );
not ( \1270_b0 , w_3817 );
and ( w_3816 , w_3817 , \1065_b0 );
or ( \1271_b1 , \1269_b1 , w_3818 );
or ( \1271_b0 , \1269_b0 , \1270_b0 );
not ( \1270_b0 , w_3819 );
and ( w_3819 , w_3818 , \1270_b1 );
or ( \1272_b1 , \1173_b1 , w_3821 );
not ( w_3821 , w_3822 );
and ( \1272_b0 , \1173_b0 , w_3823 );
and ( w_3822 ,  , w_3823 );
buf ( w_3821 , \d[0]_b1 );
not ( w_3821 , w_3824 );
not (  , w_3825 );
and ( w_3824 , w_3825 , \d[0]_b0 );
or ( \1273_b1 , \1271_b1 , w_3827 );
not ( w_3827 , w_3828 );
and ( \1273_b0 , \1271_b0 , w_3829 );
and ( w_3828 ,  , w_3829 );
buf ( w_3827 , \1272_b1 );
not ( w_3827 , w_3830 );
not (  , w_3831 );
and ( w_3830 , w_3831 , \1272_b0 );
buf ( \1274_b1 , \1273_b1 );
not ( \1274_b1 , w_3832 );
not ( \1274_b0 , w_3833 );
and ( w_3832 , w_3833 , \1273_b0 );
or ( \1275_b1 , \998_b1 , w_3835 );
not ( w_3835 , w_3836 );
and ( \1275_b0 , \998_b0 , w_3837 );
and ( w_3836 ,  , w_3837 );
buf ( w_3835 , \a[0]_b1 );
not ( w_3835 , w_3838 );
not (  , w_3839 );
and ( w_3838 , w_3839 , \a[0]_b0 );
or ( \1276_b1 , \1274_b1 , w_3841 );
not ( w_3841 , w_3842 );
and ( \1276_b0 , \1274_b0 , w_3843 );
and ( w_3842 ,  , w_3843 );
buf ( w_3841 , \1275_b1 );
not ( w_3841 , w_3844 );
not (  , w_3845 );
and ( w_3844 , w_3845 , \1275_b0 );
or ( \1277_b1 , \1267_b1 , \1276_b1 );
not ( \1276_b1 , w_3846 );
and ( \1277_b0 , \1267_b0 , w_3847 );
and ( w_3846 , w_3847 , \1276_b0 );
buf ( \1278_b1 , \1273_b1 );
not ( \1278_b1 , w_3848 );
not ( \1278_b0 , w_3849 );
and ( w_3848 , w_3849 , \1273_b0 );
or ( \1279_b1 , \1278_b1 , w_3851 );
not ( w_3851 , w_3852 );
and ( \1279_b0 , \1278_b0 , w_3853 );
and ( w_3852 ,  , w_3853 );
buf ( w_3851 , \1275_b1 );
not ( w_3851 , w_3854 );
not (  , w_3855 );
and ( w_3854 , w_3855 , \1275_b0 );
or ( \1280_b1 , \1277_b1 , w_3857 );
not ( w_3857 , w_3858 );
and ( \1280_b0 , \1277_b0 , w_3859 );
and ( w_3858 ,  , w_3859 );
buf ( w_3857 , \1279_b1 );
not ( w_3857 , w_3860 );
not (  , w_3861 );
and ( w_3860 , w_3861 , \1279_b0 );
or ( \1281_b1 , \1261_b1 , \1280_b1 );
xor ( \1281_b0 , \1261_b0 , w_3862 );
not ( w_3862 , w_3863 );
and ( w_3863 , \1280_b1 , \1280_b0 );
or ( \1282_b1 , \1237_b1 , \1230_b1 );
xor ( \1282_b0 , \1237_b0 , w_3864 );
not ( w_3864 , w_3865 );
and ( w_3865 , \1230_b1 , \1230_b0 );
or ( \1283_b1 , \1282_b1 , w_3866 );
xor ( \1283_b0 , \1282_b0 , w_3868 );
not ( w_3868 , w_3869 );
and ( w_3869 , w_3866 , w_3867 );
buf ( w_3866 , \1224_b1 );
not ( w_3866 , w_3870 );
not ( w_3867 , w_3871 );
and ( w_3870 , w_3871 , \1224_b0 );
or ( \1284_b1 , \1281_b1 , \1283_b1 );
not ( \1283_b1 , w_3872 );
and ( \1284_b0 , \1281_b0 , w_3873 );
and ( w_3872 , w_3873 , \1283_b0 );
or ( \1285_b1 , \1261_b1 , \1280_b1 );
not ( \1280_b1 , w_3874 );
and ( \1285_b0 , \1261_b0 , w_3875 );
and ( w_3874 , w_3875 , \1280_b0 );
or ( \1286_b1 , \1284_b1 , w_3876 );
or ( \1286_b0 , \1284_b0 , \1285_b0 );
not ( \1285_b0 , w_3877 );
and ( w_3877 , w_3876 , \1285_b1 );
or ( \1287_b1 , \1260_b1 , w_3879 );
not ( w_3879 , w_3880 );
and ( \1287_b0 , \1260_b0 , w_3881 );
and ( w_3880 ,  , w_3881 );
buf ( w_3879 , \1286_b1 );
not ( w_3879 , w_3882 );
not (  , w_3883 );
and ( w_3882 , w_3883 , \1286_b0 );
buf ( \1288_b1 , \1287_b1 );
not ( \1288_b1 , w_3884 );
not ( \1288_b0 , w_3885 );
and ( w_3884 , w_3885 , \1287_b0 );
buf ( \1289_b1 , \1217_b1 );
not ( \1289_b1 , w_3886 );
not ( \1289_b0 , w_3887 );
and ( w_3886 , w_3887 , \1217_b0 );
buf ( \1290_b1 , \1258_b1 );
not ( \1290_b1 , w_3888 );
not ( \1290_b0 , w_3889 );
and ( w_3888 , w_3889 , \1258_b0 );
or ( \1291_b1 , \1289_b1 , w_3890 );
or ( \1291_b0 , \1289_b0 , \1290_b0 );
not ( \1290_b0 , w_3891 );
and ( w_3891 , w_3890 , \1290_b1 );
buf ( \1292_b1 , \1255_b1 );
not ( \1292_b1 , w_3892 );
not ( \1292_b0 , w_3893 );
and ( w_3892 , w_3893 , \1255_b0 );
buf ( \1293_b1 , \1216_b1 );
not ( \1293_b1 , w_3894 );
not ( \1293_b0 , w_3895 );
and ( w_3894 , w_3895 , \1216_b0 );
or ( \1294_b1 , \1292_b1 , w_3896 );
or ( \1294_b0 , \1292_b0 , \1293_b0 );
not ( \1293_b0 , w_3897 );
and ( w_3897 , w_3896 , \1293_b1 );
or ( \1295_b1 , \1294_b1 , w_3899 );
not ( w_3899 , w_3900 );
and ( \1295_b0 , \1294_b0 , w_3901 );
and ( w_3900 ,  , w_3901 );
buf ( w_3899 , \1240_b1 );
not ( w_3899 , w_3902 );
not (  , w_3903 );
and ( w_3902 , w_3903 , \1240_b0 );
or ( \1296_b1 , \1291_b1 , w_3905 );
not ( w_3905 , w_3906 );
and ( \1296_b0 , \1291_b0 , w_3907 );
and ( w_3906 ,  , w_3907 );
buf ( w_3905 , \1295_b1 );
not ( w_3905 , w_3908 );
not (  , w_3909 );
and ( w_3908 , w_3909 , \1295_b0 );
buf ( \1297_b1 , \1202_b1 );
not ( \1297_b1 , w_3910 );
not ( \1297_b0 , w_3911 );
and ( w_3910 , w_3911 , \1202_b0 );
buf ( \1298_b1 , \1170_b1 );
not ( \1298_b1 , w_3912 );
not ( \1298_b0 , w_3913 );
and ( w_3912 , w_3913 , \1170_b0 );
or ( \1299_b1 , \1297_b1 , w_3914 );
or ( \1299_b0 , \1297_b0 , \1298_b0 );
not ( \1298_b0 , w_3915 );
and ( w_3915 , w_3914 , \1298_b1 );
or ( \1300_b1 , \1202_b1 , w_3916 );
or ( \1300_b0 , \1202_b0 , \1170_b0 );
not ( \1170_b0 , w_3917 );
and ( w_3917 , w_3916 , \1170_b1 );
or ( \1301_b1 , \1299_b1 , w_3919 );
not ( w_3919 , w_3920 );
and ( \1301_b0 , \1299_b0 , w_3921 );
and ( w_3920 ,  , w_3921 );
buf ( w_3919 , \1300_b1 );
not ( w_3919 , w_3922 );
not (  , w_3923 );
and ( w_3922 , w_3923 , \1300_b0 );
buf ( \1302_b1 , \1301_b1 );
not ( \1302_b1 , w_3924 );
not ( \1302_b0 , w_3925 );
and ( w_3924 , w_3925 , \1301_b0 );
buf ( \1303_b1 , \1302_b1 );
not ( \1303_b1 , w_3926 );
not ( \1303_b0 , w_3927 );
and ( w_3926 , w_3927 , \1302_b0 );
buf ( \1304_b1 , \1207_b1 );
not ( \1304_b1 , w_3928 );
not ( \1304_b0 , w_3929 );
and ( w_3928 , w_3929 , \1207_b0 );
or ( \1305_b1 , \1303_b1 , w_3930 );
or ( \1305_b0 , \1303_b0 , \1304_b0 );
not ( \1304_b0 , w_3931 );
and ( w_3931 , w_3930 , \1304_b1 );
or ( \1306_b1 , \1206_b1 , w_3933 );
not ( w_3933 , w_3934 );
and ( \1306_b0 , \1206_b0 , w_3935 );
and ( w_3934 ,  , w_3935 );
buf ( w_3933 , \1301_b1 );
not ( w_3933 , w_3936 );
not (  , w_3937 );
and ( w_3936 , w_3937 , \1301_b0 );
or ( \1307_b1 , \1305_b1 , w_3939 );
not ( w_3939 , w_3940 );
and ( \1307_b0 , \1305_b0 , w_3941 );
and ( w_3940 ,  , w_3941 );
buf ( w_3939 , \1306_b1 );
not ( w_3939 , w_3942 );
not (  , w_3943 );
and ( w_3942 , w_3943 , \1306_b0 );
or ( \1308_b1 , \1296_b1 , w_3945 );
not ( w_3945 , w_3946 );
and ( \1308_b0 , \1296_b0 , w_3947 );
and ( w_3946 ,  , w_3947 );
buf ( w_3945 , \1307_b1 );
not ( w_3945 , w_3948 );
not (  , w_3949 );
and ( w_3948 , w_3949 , \1307_b0 );
or ( \1309_b1 , \1288_b1 , w_3951 );
not ( w_3951 , w_3952 );
and ( \1309_b0 , \1288_b0 , w_3953 );
and ( w_3952 ,  , w_3953 );
buf ( w_3951 , \1308_b1 );
not ( w_3951 , w_3954 );
not (  , w_3955 );
and ( w_3954 , w_3955 , \1308_b0 );
buf ( \1311_b1 , \937_b1 );
not ( \1311_b1 , w_3956 );
not ( \1311_b0 , w_3957 );
and ( w_3956 , w_3957 , \937_b0 );
buf ( \1312_b1 , \933_b1 );
buf ( \1312_b0 , \933_b0 );
buf ( \1313_b1 , \1312_b1 );
not ( \1313_b1 , w_3958 );
not ( \1313_b0 , w_3959 );
and ( w_3958 , w_3959 , \1312_b0 );
or ( \1314_b1 , \1311_b1 , w_3960 );
or ( \1314_b0 , \1311_b0 , \1313_b0 );
not ( \1313_b0 , w_3961 );
and ( w_3961 , w_3960 , \1313_b1 );
or ( \1315_b1 , \a[8]_b1 , \d[5]_b1 );
xor ( \1315_b0 , \a[8]_b0 , w_3962 );
not ( w_3962 , w_3963 );
and ( w_3963 , \d[5]_b1 , \d[5]_b0 );
or ( \1316_b1 , \936_b1 , w_3965 );
not ( w_3965 , w_3966 );
and ( \1316_b0 , \936_b0 , w_3967 );
and ( w_3966 ,  , w_3967 );
buf ( w_3965 , \1315_b1 );
not ( w_3965 , w_3968 );
not (  , w_3969 );
and ( w_3968 , w_3969 , \1315_b0 );
or ( \1317_b1 , \1314_b1 , w_3971 );
not ( w_3971 , w_3972 );
and ( \1317_b0 , \1314_b0 , w_3973 );
and ( w_3972 ,  , w_3973 );
buf ( w_3971 , \1316_b1 );
not ( w_3971 , w_3974 );
not (  , w_3975 );
and ( w_3974 , w_3975 , \1316_b0 );
or ( \1318_b1 , \956_b1 , \968_b1 );
not ( \968_b1 , w_3976 );
and ( \1318_b0 , \956_b0 , w_3977 );
and ( w_3976 , w_3977 , \968_b0 );
or ( \1319_b1 , \1317_b1 , \1318_b1 );
xor ( \1319_b0 , \1317_b0 , w_3978 );
not ( w_3978 , w_3979 );
and ( w_3979 , \1318_b1 , \1318_b0 );
buf ( \1320_b1 , \1096_b1 );
not ( \1320_b1 , w_3980 );
not ( \1320_b0 , w_3981 );
and ( w_3980 , w_3981 , \1096_b0 );
buf ( \1321_b1 , \1117_b1 );
not ( \1321_b1 , w_3982 );
not ( \1321_b0 , w_3983 );
and ( w_3982 , w_3983 , \1117_b0 );
or ( \1322_b1 , \1320_b1 , w_3984 );
or ( \1322_b0 , \1320_b0 , \1321_b0 );
not ( \1321_b0 , w_3985 );
and ( w_3985 , w_3984 , \1321_b1 );
or ( \1323_b1 , \1322_b1 , w_3987 );
not ( w_3987 , w_3988 );
and ( \1323_b0 , \1322_b0 , w_3989 );
and ( w_3988 ,  , w_3989 );
buf ( w_3987 , \1103_b1 );
not ( w_3987 , w_3990 );
not (  , w_3991 );
and ( w_3990 , w_3991 , \1103_b0 );
or ( \1324_b1 , \1095_b1 , w_3993 );
not ( w_3993 , w_3994 );
and ( \1324_b0 , \1095_b0 , w_3995 );
and ( w_3994 ,  , w_3995 );
buf ( w_3993 , \1118_b1 );
not ( w_3993 , w_3996 );
not (  , w_3997 );
and ( w_3996 , w_3997 , \1118_b0 );
or ( \1325_b1 , \1323_b1 , w_3999 );
not ( w_3999 , w_4000 );
and ( \1325_b0 , \1323_b0 , w_4001 );
and ( w_4000 ,  , w_4001 );
buf ( w_3999 , \1324_b1 );
not ( w_3999 , w_4002 );
not (  , w_4003 );
and ( w_4002 , w_4003 , \1324_b0 );
or ( \1326_b1 , \1319_b1 , \1325_b1 );
xor ( \1326_b0 , \1319_b0 , w_4004 );
not ( w_4004 , w_4005 );
and ( w_4005 , \1325_b1 , \1325_b0 );
buf ( \1327_b1 , \1081_b1 );
buf ( \1327_b0 , \1081_b0 );
buf ( \1328_b1 , \1327_b1 );
not ( \1328_b1 , w_4006 );
not ( \1328_b0 , w_4007 );
and ( w_4006 , w_4007 , \1327_b0 );
buf ( \1329_b1 , \1124_b1 );
not ( \1329_b1 , w_4008 );
not ( \1329_b0 , w_4009 );
and ( w_4008 , w_4009 , \1124_b0 );
or ( \1330_b1 , \1328_b1 , w_4010 );
or ( \1330_b0 , \1328_b0 , \1329_b0 );
not ( \1329_b0 , w_4011 );
and ( w_4011 , w_4010 , \1329_b1 );
or ( \1331_b1 , \1124_b1 , w_4012 );
or ( \1331_b0 , \1124_b0 , \1327_b0 );
not ( \1327_b0 , w_4013 );
and ( w_4013 , w_4012 , \1327_b1 );
or ( \1332_b1 , \1331_b1 , w_4015 );
not ( w_4015 , w_4016 );
and ( \1332_b0 , \1331_b0 , w_4017 );
and ( w_4016 ,  , w_4017 );
buf ( w_4015 , \1088_b1 );
not ( w_4015 , w_4018 );
not (  , w_4019 );
and ( w_4018 , w_4019 , \1088_b0 );
or ( \1333_b1 , \1330_b1 , w_4021 );
not ( w_4021 , w_4022 );
and ( \1333_b0 , \1330_b0 , w_4023 );
and ( w_4022 ,  , w_4023 );
buf ( w_4021 , \1332_b1 );
not ( w_4021 , w_4024 );
not (  , w_4025 );
and ( w_4024 , w_4025 , \1332_b0 );
or ( \1334_b1 , \1326_b1 , \1333_b1 );
xor ( \1334_b0 , \1326_b0 , w_4026 );
not ( w_4026 , w_4027 );
and ( w_4027 , \1333_b1 , \1333_b0 );
or ( \1335_b1 , \d[12]_b1 , \d[11]_b1 );
xor ( \1335_b0 , \d[12]_b0 , w_4028 );
not ( w_4028 , w_4029 );
and ( w_4029 , \d[11]_b1 , \d[11]_b0 );
or ( \1336_b1 , \1335_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_4030 );
and ( \1336_b0 , \1335_b0 , w_4031 );
and ( w_4030 , w_4031 , \a[0]_b0 );
buf ( \1337_b1 , \1101_b1 );
not ( \1337_b1 , w_4032 );
not ( \1337_b0 , w_4033 );
and ( w_4032 , w_4033 , \1101_b0 );
buf ( \1338_b1 , \1038_b1 );
not ( \1338_b1 , w_4034 );
not ( \1338_b0 , w_4035 );
and ( w_4034 , w_4035 , \1038_b0 );
or ( \1339_b1 , \1337_b1 , w_4036 );
or ( \1339_b0 , \1337_b0 , \1338_b0 );
not ( \1338_b0 , w_4037 );
and ( w_4037 , w_4036 , \1338_b1 );
or ( \1340_b1 , \a[6]_b1 , \d[7]_b1 );
xor ( \1340_b0 , \a[6]_b0 , w_4038 );
not ( w_4038 , w_4039 );
and ( w_4039 , \d[7]_b1 , \d[7]_b0 );
or ( \1341_b1 , \998_b1 , w_4041 );
not ( w_4041 , w_4042 );
and ( \1341_b0 , \998_b0 , w_4043 );
and ( w_4042 ,  , w_4043 );
buf ( w_4041 , \1340_b1 );
not ( w_4041 , w_4044 );
not (  , w_4045 );
and ( w_4044 , w_4045 , \1340_b0 );
or ( \1342_b1 , \1339_b1 , w_4047 );
not ( w_4047 , w_4048 );
and ( \1342_b0 , \1339_b0 , w_4049 );
and ( w_4048 ,  , w_4049 );
buf ( w_4047 , \1341_b1 );
not ( w_4047 , w_4050 );
not (  , w_4051 );
and ( w_4050 , w_4051 , \1341_b0 );
or ( \1343_b1 , \1336_b1 , \1342_b1 );
xor ( \1343_b0 , \1336_b0 , w_4052 );
not ( w_4052 , w_4053 );
and ( w_4053 , \1342_b1 , \1342_b0 );
buf ( \1344_b1 , \966_b1 );
not ( \1344_b1 , w_4054 );
not ( \1344_b0 , w_4055 );
and ( w_4054 , w_4055 , \966_b0 );
buf ( \1345_b1 , \980_b1 );
not ( \1345_b1 , w_4056 );
not ( \1345_b0 , w_4057 );
and ( w_4056 , w_4057 , \980_b0 );
or ( \1346_b1 , \1344_b1 , w_4058 );
or ( \1346_b0 , \1344_b0 , \1345_b0 );
not ( \1345_b0 , w_4059 );
and ( w_4059 , w_4058 , \1345_b1 );
or ( \1347_b1 , \a[10]_b1 , \d[3]_b1 );
xor ( \1347_b0 , \a[10]_b0 , w_4060 );
not ( w_4060 , w_4061 );
and ( w_4061 , \d[3]_b1 , \d[3]_b0 );
or ( \1348_b1 , \965_b1 , w_4063 );
not ( w_4063 , w_4064 );
and ( \1348_b0 , \965_b0 , w_4065 );
and ( w_4064 ,  , w_4065 );
buf ( w_4063 , \1347_b1 );
not ( w_4063 , w_4066 );
not (  , w_4067 );
and ( w_4066 , w_4067 , \1347_b0 );
or ( \1349_b1 , \1346_b1 , w_4069 );
not ( w_4069 , w_4070 );
and ( \1349_b0 , \1346_b0 , w_4071 );
and ( w_4070 ,  , w_4071 );
buf ( w_4069 , \1348_b1 );
not ( w_4069 , w_4072 );
not (  , w_4073 );
and ( w_4072 , w_4073 , \1348_b0 );
or ( \1350_b1 , \1343_b1 , \1349_b1 );
xor ( \1350_b0 , \1343_b0 , w_4074 );
not ( w_4074 , w_4075 );
and ( w_4075 , \1349_b1 , \1349_b0 );
buf ( \1351_b1 , \1109_b1 );
not ( \1351_b1 , w_4076 );
not ( \1351_b0 , w_4077 );
and ( w_4076 , w_4077 , \1109_b0 );
buf ( \1352_b1 , \1115_b1 );
not ( \1352_b1 , w_4078 );
not ( \1352_b0 , w_4079 );
and ( w_4078 , w_4079 , \1115_b0 );
or ( \1353_b1 , \1351_b1 , w_4080 );
or ( \1353_b0 , \1351_b0 , \1352_b0 );
not ( \1352_b0 , w_4081 );
and ( w_4081 , w_4080 , \1352_b1 );
or ( \1354_b1 , \a[4]_b1 , w_4082 );
xor ( \1354_b0 , \a[4]_b0 , w_4084 );
not ( w_4084 , w_4085 );
and ( w_4085 , w_4082 , w_4083 );
buf ( w_4082 , \d[9]_b1 );
not ( w_4082 , w_4086 );
not ( w_4083 , w_4087 );
and ( w_4086 , w_4087 , \d[9]_b0 );
buf ( \1355_b1 , \1354_b1 );
not ( \1355_b1 , w_4088 );
not ( \1355_b0 , w_4089 );
and ( w_4088 , w_4089 , \1354_b0 );
or ( \1356_b1 , \1355_b1 , w_4091 );
not ( w_4091 , w_4092 );
and ( \1356_b0 , \1355_b0 , w_4093 );
and ( w_4092 ,  , w_4093 );
buf ( w_4091 , \1029_b1 );
not ( w_4091 , w_4094 );
not (  , w_4095 );
and ( w_4094 , w_4095 , \1029_b0 );
or ( \1357_b1 , \1353_b1 , w_4097 );
not ( w_4097 , w_4098 );
and ( \1357_b0 , \1353_b0 , w_4099 );
and ( w_4098 ,  , w_4099 );
buf ( w_4097 , \1356_b1 );
not ( w_4097 , w_4100 );
not (  , w_4101 );
and ( w_4100 , w_4101 , \1356_b0 );
buf ( \1358_b1 , \1065_b1 );
not ( \1358_b1 , w_4102 );
not ( \1358_b0 , w_4103 );
and ( w_4102 , w_4103 , \1065_b0 );
buf ( \1359_b1 , \1093_b1 );
not ( \1359_b1 , w_4104 );
not ( \1359_b0 , w_4105 );
and ( w_4104 , w_4105 , \1093_b0 );
or ( \1360_b1 , \1358_b1 , w_4106 );
or ( \1360_b0 , \1358_b0 , \1359_b0 );
not ( \1359_b0 , w_4107 );
and ( w_4107 , w_4106 , \1359_b1 );
or ( \1361_b1 , \d[1]_b1 , \a[12]_b1 );
xor ( \1361_b0 , \d[1]_b0 , w_4108 );
not ( w_4108 , w_4109 );
and ( w_4109 , \a[12]_b1 , \a[12]_b0 );
or ( \1362_b1 , \1361_b1 , w_4111 );
not ( w_4111 , w_4112 );
and ( \1362_b0 , \1361_b0 , w_4113 );
and ( w_4112 ,  , w_4113 );
buf ( w_4111 , \d[0]_b1 );
not ( w_4111 , w_4114 );
not (  , w_4115 );
and ( w_4114 , w_4115 , \d[0]_b0 );
or ( \1363_b1 , \1360_b1 , w_4117 );
not ( w_4117 , w_4118 );
and ( \1363_b0 , \1360_b0 , w_4119 );
and ( w_4118 ,  , w_4119 );
buf ( w_4117 , \1362_b1 );
not ( w_4117 , w_4120 );
not (  , w_4121 );
and ( w_4120 , w_4121 , \1362_b0 );
or ( \1364_b1 , \1357_b1 , \1363_b1 );
xor ( \1364_b0 , \1357_b0 , w_4122 );
not ( w_4122 , w_4123 );
and ( w_4123 , \1363_b1 , \1363_b0 );
buf ( \1365_b1 , \948_b1 );
not ( \1365_b1 , w_4124 );
not ( \1365_b0 , w_4125 );
and ( w_4124 , w_4125 , \948_b0 );
or ( \1366_b1 , \947_b1 , w_4127 );
not ( w_4127 , w_4128 );
and ( \1366_b0 , \947_b0 , w_4129 );
and ( w_4128 ,  , w_4129 );
buf ( w_4127 , \942_b1 );
not ( w_4127 , w_4130 );
not (  , w_4131 );
and ( w_4130 , w_4131 , \942_b0 );
buf ( \1367_b1 , \1366_b1 );
not ( \1367_b1 , w_4132 );
not ( \1367_b0 , w_4133 );
and ( w_4132 , w_4133 , \1366_b0 );
or ( \1368_b1 , \1365_b1 , w_4134 );
or ( \1368_b0 , \1365_b0 , \1367_b0 );
not ( \1367_b0 , w_4135 );
and ( w_4135 , w_4134 , \1367_b1 );
or ( \1369_b1 , \a[2]_b1 , \d[11]_b1 );
xor ( \1369_b0 , \a[2]_b0 , w_4136 );
not ( w_4136 , w_4137 );
and ( w_4137 , \d[11]_b1 , \d[11]_b0 );
or ( \1370_b1 , \947_b1 , w_4139 );
not ( w_4139 , w_4140 );
and ( \1370_b0 , \947_b0 , w_4141 );
and ( w_4140 ,  , w_4141 );
buf ( w_4139 , \1369_b1 );
not ( w_4139 , w_4142 );
not (  , w_4143 );
and ( w_4142 , w_4143 , \1369_b0 );
or ( \1371_b1 , \1368_b1 , w_4145 );
not ( w_4145 , w_4146 );
and ( \1371_b0 , \1368_b0 , w_4147 );
and ( w_4146 ,  , w_4147 );
buf ( w_4145 , \1370_b1 );
not ( w_4145 , w_4148 );
not (  , w_4149 );
and ( w_4148 , w_4149 , \1370_b0 );
or ( \1372_b1 , \1364_b1 , \1371_b1 );
xor ( \1372_b0 , \1364_b0 , w_4150 );
not ( w_4150 , w_4151 );
and ( w_4151 , \1371_b1 , \1371_b0 );
or ( \1373_b1 , \1350_b1 , \1372_b1 );
xor ( \1373_b0 , \1350_b0 , w_4152 );
not ( w_4152 , w_4153 );
and ( w_4153 , \1372_b1 , \1372_b0 );
buf ( \1374_b1 , \939_b1 );
not ( \1374_b1 , w_4154 );
not ( \1374_b0 , w_4155 );
and ( w_4154 , w_4155 , \939_b0 );
or ( \1375_b1 , \1374_b1 , w_4157 );
not ( w_4157 , w_4158 );
and ( \1375_b0 , \1374_b0 , w_4159 );
and ( w_4158 ,  , w_4159 );
buf ( w_4157 , \951_b1 );
not ( w_4157 , w_4160 );
not (  , w_4161 );
and ( w_4160 , w_4161 , \951_b0 );
buf ( \1376_b1 , \1375_b1 );
not ( \1376_b1 , w_4162 );
not ( \1376_b0 , w_4163 );
and ( w_4162 , w_4163 , \1375_b0 );
buf ( \1377_b1 , \969_b1 );
not ( \1377_b1 , w_4164 );
not ( \1377_b0 , w_4165 );
and ( w_4164 , w_4165 , \969_b0 );
or ( \1378_b1 , \1376_b1 , w_4166 );
or ( \1378_b0 , \1376_b0 , \1377_b0 );
not ( \1377_b0 , w_4167 );
and ( w_4167 , w_4166 , \1377_b1 );
or ( \1379_b1 , \939_b1 , w_4169 );
not ( w_4169 , w_4170 );
and ( \1379_b0 , \939_b0 , w_4171 );
and ( w_4170 ,  , w_4171 );
buf ( w_4169 , \950_b1 );
not ( w_4169 , w_4172 );
not (  , w_4173 );
and ( w_4172 , w_4173 , \950_b0 );
or ( \1380_b1 , \1378_b1 , w_4175 );
not ( w_4175 , w_4176 );
and ( \1380_b0 , \1378_b0 , w_4177 );
and ( w_4176 ,  , w_4177 );
buf ( w_4175 , \1379_b1 );
not ( w_4175 , w_4178 );
not (  , w_4179 );
and ( w_4178 , w_4179 , \1379_b0 );
or ( \1381_b1 , \1373_b1 , \1380_b1 );
xor ( \1381_b0 , \1373_b0 , w_4180 );
not ( w_4180 , w_4181 );
and ( w_4181 , \1380_b1 , \1380_b0 );
or ( \1382_b1 , \1334_b1 , \1381_b1 );
xor ( \1382_b0 , \1334_b0 , w_4182 );
not ( w_4182 , w_4183 );
and ( w_4183 , \1381_b1 , \1381_b0 );
or ( \1383_b1 , \1050_b1 , w_4185 );
not ( w_4185 , w_4186 );
and ( \1383_b0 , \1050_b0 , w_4187 );
and ( w_4186 ,  , w_4187 );
buf ( w_4185 , \970_b1 );
not ( w_4185 , w_4188 );
not (  , w_4189 );
and ( w_4188 , w_4189 , \970_b0 );
or ( \1384_b1 , \1125_b1 , w_4190 );
or ( \1384_b0 , \1125_b0 , \1383_b0 );
not ( \1383_b0 , w_4191 );
and ( w_4191 , w_4190 , \1383_b1 );
or ( \1385_b1 , \1050_b1 , w_4193 );
not ( w_4193 , w_4194 );
and ( \1385_b0 , \1050_b0 , w_4195 );
and ( w_4194 ,  , w_4195 );
buf ( w_4193 , \970_b1 );
not ( w_4193 , w_4196 );
not (  , w_4197 );
and ( w_4196 , w_4197 , \970_b0 );
or ( \1386_b1 , \1384_b1 , w_4199 );
not ( w_4199 , w_4200 );
and ( \1386_b0 , \1384_b0 , w_4201 );
and ( w_4200 ,  , w_4201 );
buf ( w_4199 , \1385_b1 );
not ( w_4199 , w_4202 );
not (  , w_4203 );
and ( w_4202 , w_4203 , \1385_b0 );
or ( \1387_b1 , \1382_b1 , w_4205 );
not ( w_4205 , w_4206 );
and ( \1387_b0 , \1382_b0 , w_4207 );
and ( w_4206 ,  , w_4207 );
buf ( w_4205 , \1386_b1 );
not ( w_4205 , w_4208 );
not (  , w_4209 );
and ( w_4208 , w_4209 , \1386_b0 );
buf ( \1388_b1 , \1387_b1 );
not ( \1388_b1 , w_4210 );
not ( \1388_b0 , w_4211 );
and ( w_4210 , w_4211 , \1387_b0 );
or ( \1389_b1 , \1261_b1 , \1280_b1 );
xor ( \1389_b0 , \1261_b0 , w_4212 );
not ( w_4212 , w_4213 );
and ( w_4213 , \1280_b1 , \1280_b0 );
or ( \1390_b1 , \1389_b1 , \1283_b1 );
xor ( \1390_b0 , \1389_b0 , w_4214 );
not ( w_4214 , w_4215 );
and ( w_4215 , \1283_b1 , \1283_b0 );
or ( \1391_b1 , \1275_b1 , \1273_b1 );
xor ( \1391_b0 , \1275_b0 , w_4216 );
not ( w_4216 , w_4217 );
and ( w_4217 , \1273_b1 , \1273_b0 );
or ( \1392_b1 , \1391_b1 , w_4218 );
xor ( \1392_b0 , \1391_b0 , w_4220 );
not ( w_4220 , w_4221 );
and ( w_4221 , w_4218 , w_4219 );
buf ( w_4218 , \1267_b1 );
not ( w_4218 , w_4222 );
not ( w_4219 , w_4223 );
and ( w_4222 , w_4223 , \1267_b0 );
or ( \1393_b1 , \a[0]_b1 , w_4224 );
or ( \1393_b0 , \a[0]_b0 , \d[4]_b0 );
not ( \d[4]_b0 , w_4225 );
and ( w_4225 , w_4224 , \d[4]_b1 );
or ( \1394_b1 , \1393_b1 , w_4227 );
not ( w_4227 , w_4228 );
and ( \1394_b0 , \1393_b0 , w_4229 );
and ( w_4228 ,  , w_4229 );
buf ( w_4227 , \d[3]_b1 );
not ( w_4227 , w_4230 );
not (  , w_4231 );
and ( w_4230 , w_4231 , \d[3]_b0 );
or ( \1395_b1 , \a[0]_b1 , w_4233 );
not ( w_4233 , w_4234 );
and ( \1395_b0 , \a[0]_b0 , w_4235 );
and ( w_4234 ,  , w_4235 );
buf ( w_4233 , \d[4]_b1 );
not ( w_4233 , w_4236 );
not (  , w_4237 );
and ( w_4236 , w_4237 , \d[4]_b0 );
buf ( \1397_b1 , \1396_b1 );
not ( \1397_b1 , w_4238 );
not ( \1397_b0 , w_4239 );
and ( w_4238 , w_4239 , \1396_b0 );
or ( \1398_b1 , \a[4]_b1 , \d[1]_b1 );
xor ( \1398_b0 , \a[4]_b0 , w_4240 );
not ( w_4240 , w_4241 );
and ( w_4241 , \d[1]_b1 , \d[1]_b0 );
buf ( \1399_b1 , \1398_b1 );
not ( \1399_b1 , w_4242 );
not ( \1399_b0 , w_4243 );
and ( w_4242 , w_4243 , \1398_b0 );
buf ( \1400_b1 , \1012_b1 );
not ( \1400_b1 , w_4244 );
not ( \1400_b0 , w_4245 );
and ( w_4244 , w_4245 , \1012_b0 );
or ( \1401_b1 , \1399_b1 , w_4246 );
or ( \1401_b0 , \1399_b0 , \1400_b0 );
not ( \1400_b0 , w_4247 );
and ( w_4247 , w_4246 , \1400_b1 );
or ( \1402_b1 , \1268_b1 , w_4249 );
not ( w_4249 , w_4250 );
and ( \1402_b0 , \1268_b0 , w_4251 );
and ( w_4250 ,  , w_4251 );
buf ( w_4249 , \d[0]_b1 );
not ( w_4249 , w_4252 );
not (  , w_4253 );
and ( w_4252 , w_4253 , \d[0]_b0 );
or ( \1403_b1 , \1401_b1 , w_4255 );
not ( w_4255 , w_4256 );
and ( \1403_b0 , \1401_b0 , w_4257 );
and ( w_4256 ,  , w_4257 );
buf ( w_4255 , \1402_b1 );
not ( w_4255 , w_4258 );
not (  , w_4259 );
and ( w_4258 , w_4259 , \1402_b0 );
or ( \1404_b1 , \1397_b1 , w_4261 );
not ( w_4261 , w_4262 );
and ( \1404_b0 , \1397_b0 , w_4263 );
and ( w_4262 ,  , w_4263 );
buf ( w_4261 , \1403_b1 );
not ( w_4261 , w_4264 );
not (  , w_4265 );
and ( w_4264 , w_4265 , \1403_b0 );
or ( \1405_b1 , \a[1]_b1 , \d[5]_b1 );
xor ( \1405_b0 , \a[1]_b0 , w_4266 );
not ( w_4266 , w_4267 );
and ( w_4267 , \d[5]_b1 , \d[5]_b0 );
buf ( \1406_b1 , \1405_b1 );
not ( \1406_b1 , w_4268 );
not ( \1406_b0 , w_4269 );
and ( w_4268 , w_4269 , \1405_b0 );
buf ( \1407_b1 , \1186_b1 );
not ( \1407_b1 , w_4270 );
not ( \1407_b0 , w_4271 );
and ( w_4270 , w_4271 , \1186_b0 );
or ( \1408_b1 , \1406_b1 , w_4272 );
or ( \1408_b0 , \1406_b0 , \1407_b0 );
not ( \1407_b0 , w_4273 );
and ( w_4273 , w_4272 , \1407_b1 );
or ( \1409_b1 , \936_b1 , w_4275 );
not ( w_4275 , w_4276 );
and ( \1409_b0 , \936_b0 , w_4277 );
and ( w_4276 ,  , w_4277 );
buf ( w_4275 , \1225_b1 );
not ( w_4275 , w_4278 );
not (  , w_4279 );
and ( w_4278 , w_4279 , \1225_b0 );
or ( \1410_b1 , \1408_b1 , w_4281 );
not ( w_4281 , w_4282 );
and ( \1410_b0 , \1408_b0 , w_4283 );
and ( w_4282 ,  , w_4283 );
buf ( w_4281 , \1409_b1 );
not ( w_4281 , w_4284 );
not (  , w_4285 );
and ( w_4284 , w_4285 , \1409_b0 );
buf ( \1411_b1 , \1410_b1 );
not ( \1411_b1 , w_4286 );
not ( \1411_b0 , w_4287 );
and ( w_4286 , w_4287 , \1410_b0 );
or ( \1412_b1 , \1404_b1 , w_4289 );
not ( w_4289 , w_4290 );
and ( \1412_b0 , \1404_b0 , w_4291 );
and ( w_4290 ,  , w_4291 );
buf ( w_4289 , \1411_b1 );
not ( w_4289 , w_4292 );
not (  , w_4293 );
and ( w_4292 , w_4293 , \1411_b0 );
or ( \1413_b1 , \1392_b1 , \1412_b1 );
not ( \1412_b1 , w_4294 );
and ( \1413_b0 , \1392_b0 , w_4295 );
and ( w_4294 , w_4295 , \1412_b0 );
buf ( \1414_b1 , \1404_b1 );
not ( \1414_b1 , w_4296 );
not ( \1414_b0 , w_4297 );
and ( w_4296 , w_4297 , \1404_b0 );
or ( \1415_b1 , \1414_b1 , \1410_b1 );
not ( \1410_b1 , w_4298 );
and ( \1415_b0 , \1414_b0 , w_4299 );
and ( w_4298 , w_4299 , \1410_b0 );
or ( \1416_b1 , \1413_b1 , w_4301 );
not ( w_4301 , w_4302 );
and ( \1416_b0 , \1413_b0 , w_4303 );
and ( w_4302 ,  , w_4303 );
buf ( w_4301 , \1415_b1 );
not ( w_4301 , w_4304 );
not (  , w_4305 );
and ( w_4304 , w_4305 , \1415_b0 );
or ( \1417_b1 , \1390_b1 , w_4307 );
not ( w_4307 , w_4308 );
and ( \1417_b0 , \1390_b0 , w_4309 );
and ( w_4308 ,  , w_4309 );
buf ( w_4307 , \1416_b1 );
not ( w_4307 , w_4310 );
not (  , w_4311 );
and ( w_4310 , w_4311 , \1416_b0 );
buf ( \1418_b1 , \1417_b1 );
not ( \1418_b1 , w_4312 );
not ( \1418_b0 , w_4313 );
and ( w_4312 , w_4313 , \1417_b0 );
buf ( \1419_b1 , \1405_b1 );
not ( \1419_b1 , w_4314 );
not ( \1419_b0 , w_4315 );
and ( w_4314 , w_4315 , \1405_b0 );
buf ( \1420_b1 , \932_b1 );
not ( \1420_b1 , w_4316 );
not ( \1420_b0 , w_4317 );
and ( w_4316 , w_4317 , \932_b0 );
or ( \1421_b1 , \1419_b1 , w_4318 );
or ( \1421_b0 , \1419_b0 , \1420_b0 );
not ( \1420_b0 , w_4319 );
and ( w_4319 , w_4318 , \1420_b1 );
or ( \1422_b1 , \a[0]_b1 , \d[5]_b1 );
xor ( \1422_b0 , \a[0]_b0 , w_4320 );
not ( w_4320 , w_4321 );
and ( w_4321 , \d[5]_b1 , \d[5]_b0 );
or ( \1423_b1 , \930_b1 , w_4323 );
not ( w_4323 , w_4324 );
and ( \1423_b0 , \930_b0 , w_4325 );
and ( w_4324 ,  , w_4325 );
buf ( w_4323 , \1422_b1 );
not ( w_4323 , w_4326 );
not (  , w_4327 );
and ( w_4326 , w_4327 , \1422_b0 );
or ( \1424_b1 , \932_b1 , w_4328 );
or ( \1424_b0 , \932_b0 , \1423_b0 );
not ( \1423_b0 , w_4329 );
and ( w_4329 , w_4328 , \1423_b1 );
or ( \1425_b1 , \1421_b1 , w_4331 );
not ( w_4331 , w_4332 );
and ( \1425_b0 , \1421_b0 , w_4333 );
and ( w_4332 ,  , w_4333 );
buf ( w_4331 , \1424_b1 );
not ( w_4331 , w_4334 );
not (  , w_4335 );
and ( w_4334 , w_4335 , \1424_b0 );
or ( \1426_b1 , \a[2]_b1 , \d[3]_b1 );
xor ( \1426_b0 , \a[2]_b0 , w_4336 );
not ( w_4336 , w_4337 );
and ( w_4337 , \d[3]_b1 , \d[3]_b0 );
buf ( \1427_b1 , \1426_b1 );
not ( \1427_b1 , w_4338 );
not ( \1427_b0 , w_4339 );
and ( w_4338 , w_4339 , \1426_b0 );
buf ( \1428_b1 , \980_b1 );
not ( \1428_b1 , w_4340 );
not ( \1428_b0 , w_4341 );
and ( w_4340 , w_4341 , \980_b0 );
or ( \1429_b1 , \1427_b1 , w_4342 );
or ( \1429_b0 , \1427_b0 , \1428_b0 );
not ( \1428_b0 , w_4343 );
and ( w_4343 , w_4342 , \1428_b1 );
or ( \1430_b1 , \965_b1 , w_4345 );
not ( w_4345 , w_4346 );
and ( \1430_b0 , \965_b0 , w_4347 );
and ( w_4346 ,  , w_4347 );
buf ( w_4345 , \1262_b1 );
not ( w_4345 , w_4348 );
not (  , w_4349 );
and ( w_4348 , w_4349 , \1262_b0 );
or ( \1431_b1 , \1429_b1 , w_4351 );
not ( w_4351 , w_4352 );
and ( \1431_b0 , \1429_b0 , w_4353 );
and ( w_4352 ,  , w_4353 );
buf ( w_4351 , \1430_b1 );
not ( w_4351 , w_4354 );
not (  , w_4355 );
and ( w_4354 , w_4355 , \1430_b0 );
or ( \1432_b1 , \1425_b1 , \1431_b1 );
xor ( \1432_b0 , \1425_b0 , w_4356 );
not ( w_4356 , w_4357 );
and ( w_4357 , \1431_b1 , \1431_b0 );
buf ( \1433_b1 , \1396_b1 );
not ( \1433_b1 , w_4358 );
not ( \1433_b0 , w_4359 );
and ( w_4358 , w_4359 , \1396_b0 );
buf ( \1434_b1 , \1403_b1 );
not ( \1434_b1 , w_4360 );
not ( \1434_b0 , w_4361 );
and ( w_4360 , w_4361 , \1403_b0 );
or ( \1435_b1 , \1433_b1 , w_4362 );
or ( \1435_b0 , \1433_b0 , \1434_b0 );
not ( \1434_b0 , w_4363 );
and ( w_4363 , w_4362 , \1434_b1 );
or ( \1436_b1 , \1403_b1 , w_4364 );
or ( \1436_b0 , \1403_b0 , \1396_b0 );
not ( \1396_b0 , w_4365 );
and ( w_4365 , w_4364 , \1396_b1 );
or ( \1437_b1 , \1435_b1 , w_4367 );
not ( w_4367 , w_4368 );
and ( \1437_b0 , \1435_b0 , w_4369 );
and ( w_4368 ,  , w_4369 );
buf ( w_4367 , \1436_b1 );
not ( w_4367 , w_4370 );
not (  , w_4371 );
and ( w_4370 , w_4371 , \1436_b0 );
or ( \1438_b1 , \1432_b1 , \1437_b1 );
not ( \1437_b1 , w_4372 );
and ( \1438_b0 , \1432_b0 , w_4373 );
and ( w_4372 , w_4373 , \1437_b0 );
or ( \1439_b1 , \1425_b1 , \1431_b1 );
not ( \1431_b1 , w_4374 );
and ( \1439_b0 , \1425_b0 , w_4375 );
and ( w_4374 , w_4375 , \1431_b0 );
or ( \1440_b1 , \1438_b1 , w_4376 );
or ( \1440_b0 , \1438_b0 , \1439_b0 );
not ( \1439_b0 , w_4377 );
and ( w_4377 , w_4376 , \1439_b1 );
or ( \1441_b1 , \1414_b1 , \1411_b1 );
xor ( \1441_b0 , \1414_b0 , w_4378 );
not ( w_4378 , w_4379 );
and ( w_4379 , \1411_b1 , \1411_b0 );
or ( \1442_b1 , \1441_b1 , w_4380 );
xor ( \1442_b0 , \1441_b0 , w_4382 );
not ( w_4382 , w_4383 );
and ( w_4383 , w_4380 , w_4381 );
buf ( w_4380 , \1392_b1 );
not ( w_4380 , w_4384 );
not ( w_4381 , w_4385 );
and ( w_4384 , w_4385 , \1392_b0 );
or ( \1443_b1 , \1440_b1 , \1442_b1 );
xor ( \1443_b0 , \1440_b0 , w_4386 );
not ( w_4386 , w_4387 );
and ( w_4387 , \1442_b1 , \1442_b0 );
or ( \1444_b1 , \1425_b1 , \1431_b1 );
xor ( \1444_b0 , \1425_b0 , w_4388 );
not ( w_4388 , w_4389 );
and ( w_4389 , \1431_b1 , \1431_b0 );
or ( \1445_b1 , \1444_b1 , \1437_b1 );
xor ( \1445_b0 , \1444_b0 , w_4390 );
not ( w_4390 , w_4391 );
and ( w_4391 , \1437_b1 , \1437_b0 );
or ( \1446_b1 , \a[1]_b1 , \d[3]_b1 );
xor ( \1446_b0 , \a[1]_b0 , w_4392 );
not ( w_4392 , w_4393 );
and ( w_4393 , \d[3]_b1 , \d[3]_b0 );
or ( \1447_b1 , \961_b1 , w_4395 );
not ( w_4395 , w_4396 );
and ( \1447_b0 , \961_b0 , w_4397 );
and ( w_4396 ,  , w_4397 );
buf ( w_4395 , \1446_b1 );
not ( w_4395 , w_4398 );
not (  , w_4399 );
and ( w_4398 , w_4399 , \1446_b0 );
or ( \1448_b1 , \1447_b1 , w_4400 );
or ( \1448_b0 , \1447_b0 , \965_b0 );
not ( \965_b0 , w_4401 );
and ( w_4401 , w_4400 , \965_b1 );
or ( \1449_b1 , \959_b1 , w_4403 );
not ( w_4403 , w_4404 );
and ( \1449_b0 , \959_b0 , w_4405 );
and ( w_4404 ,  , w_4405 );
buf ( w_4403 , \1426_b1 );
not ( w_4403 , w_4406 );
not (  , w_4407 );
and ( w_4406 , w_4407 , \1426_b0 );
or ( \1450_b1 , \1448_b1 , w_4409 );
not ( w_4409 , w_4410 );
and ( \1450_b0 , \1448_b0 , w_4411 );
and ( w_4410 ,  , w_4411 );
buf ( w_4409 , \1449_b1 );
not ( w_4409 , w_4412 );
not (  , w_4413 );
and ( w_4412 , w_4413 , \1449_b0 );
buf ( \1451_b1 , \1450_b1 );
not ( \1451_b1 , w_4414 );
not ( \1451_b0 , w_4415 );
and ( w_4414 , w_4415 , \1450_b0 );
or ( \1452_b1 , \d[1]_b1 , \a[3]_b1 );
xor ( \1452_b0 , \d[1]_b0 , w_4416 );
not ( w_4416 , w_4417 );
and ( w_4417 , \a[3]_b1 , \a[3]_b0 );
buf ( \1453_b1 , \1452_b1 );
not ( \1453_b1 , w_4418 );
not ( \1453_b0 , w_4419 );
and ( w_4418 , w_4419 , \1452_b0 );
buf ( \1454_b1 , \1012_b1 );
not ( \1454_b1 , w_4420 );
not ( \1454_b0 , w_4421 );
and ( w_4420 , w_4421 , \1012_b0 );
or ( \1455_b1 , \1453_b1 , w_4422 );
or ( \1455_b0 , \1453_b0 , \1454_b0 );
not ( \1454_b0 , w_4423 );
and ( w_4423 , w_4422 , \1454_b1 );
or ( \1456_b1 , \1398_b1 , w_4425 );
not ( w_4425 , w_4426 );
and ( \1456_b0 , \1398_b0 , w_4427 );
and ( w_4426 ,  , w_4427 );
buf ( w_4425 , \d[0]_b1 );
not ( w_4425 , w_4428 );
not (  , w_4429 );
and ( w_4428 , w_4429 , \d[0]_b0 );
or ( \1457_b1 , \1455_b1 , w_4431 );
not ( w_4431 , w_4432 );
and ( \1457_b0 , \1455_b0 , w_4433 );
and ( w_4432 ,  , w_4433 );
buf ( w_4431 , \1456_b1 );
not ( w_4431 , w_4434 );
not (  , w_4435 );
and ( w_4434 , w_4435 , \1456_b0 );
buf ( \1458_b1 , \1457_b1 );
not ( \1458_b1 , w_4436 );
not ( \1458_b0 , w_4437 );
and ( w_4436 , w_4437 , \1457_b0 );
or ( \1459_b1 , \932_b1 , w_4439 );
not ( w_4439 , w_4440 );
and ( \1459_b0 , \932_b0 , w_4441 );
and ( w_4440 ,  , w_4441 );
buf ( w_4439 , \a[0]_b1 );
not ( w_4439 , w_4442 );
not (  , w_4443 );
and ( w_4442 , w_4443 , \a[0]_b0 );
or ( \1460_b1 , \1458_b1 , w_4445 );
not ( w_4445 , w_4446 );
and ( \1460_b0 , \1458_b0 , w_4447 );
and ( w_4446 ,  , w_4447 );
buf ( w_4445 , \1459_b1 );
not ( w_4445 , w_4448 );
not (  , w_4449 );
and ( w_4448 , w_4449 , \1459_b0 );
buf ( \1461_b1 , \1460_b1 );
not ( \1461_b1 , w_4450 );
not ( \1461_b0 , w_4451 );
and ( w_4450 , w_4451 , \1460_b0 );
or ( \1462_b1 , \1451_b1 , w_4452 );
or ( \1462_b0 , \1451_b0 , \1461_b0 );
not ( \1461_b0 , w_4453 );
and ( w_4453 , w_4452 , \1461_b1 );
buf ( \1463_b1 , \1459_b1 );
not ( \1463_b1 , w_4454 );
not ( \1463_b0 , w_4455 );
and ( w_4454 , w_4455 , \1459_b0 );
or ( \1464_b1 , \1463_b1 , w_4457 );
not ( w_4457 , w_4458 );
and ( \1464_b0 , \1463_b0 , w_4459 );
and ( w_4458 ,  , w_4459 );
buf ( w_4457 , \1457_b1 );
not ( w_4457 , w_4460 );
not (  , w_4461 );
and ( w_4460 , w_4461 , \1457_b0 );
or ( \1465_b1 , \1462_b1 , w_4463 );
not ( w_4463 , w_4464 );
and ( \1465_b0 , \1462_b0 , w_4465 );
and ( w_4464 ,  , w_4465 );
buf ( w_4463 , \1464_b1 );
not ( w_4463 , w_4466 );
not (  , w_4467 );
and ( w_4466 , w_4467 , \1464_b0 );
or ( \1466_b1 , \1445_b1 , w_4469 );
not ( w_4469 , w_4470 );
and ( \1466_b0 , \1445_b0 , w_4471 );
and ( w_4470 ,  , w_4471 );
buf ( w_4469 , \1465_b1 );
not ( w_4469 , w_4472 );
not (  , w_4473 );
and ( w_4472 , w_4473 , \1465_b0 );
or ( \1467_b1 , \d[1]_b1 , \a[2]_b1 );
xor ( \1467_b0 , \d[1]_b0 , w_4474 );
not ( w_4474 , w_4475 );
and ( w_4475 , \a[2]_b1 , \a[2]_b0 );
or ( \1468_b1 , \1065_b1 , \1467_b1 );
not ( \1467_b1 , w_4476 );
and ( \1468_b0 , \1065_b0 , w_4477 );
and ( w_4476 , w_4477 , \1467_b0 );
or ( \1469_b1 , \1452_b1 , \d[0]_b1 );
not ( \d[0]_b1 , w_4478 );
and ( \1469_b0 , \1452_b0 , w_4479 );
and ( w_4478 , w_4479 , \d[0]_b0 );
or ( \1470_b1 , \1468_b1 , w_4481 );
not ( w_4481 , w_4482 );
and ( \1470_b0 , \1468_b0 , w_4483 );
and ( w_4482 ,  , w_4483 );
buf ( w_4481 , \1469_b1 );
not ( w_4481 , w_4484 );
not (  , w_4485 );
and ( w_4484 , w_4485 , \1469_b0 );
or ( \1471_b1 , \a[0]_b1 , w_4486 );
or ( \1471_b0 , \a[0]_b0 , \d[2]_b0 );
not ( \d[2]_b0 , w_4487 );
and ( w_4487 , w_4486 , \d[2]_b1 );
or ( \1472_b1 , \1471_b1 , w_4489 );
not ( w_4489 , w_4490 );
and ( \1472_b0 , \1471_b0 , w_4491 );
and ( w_4490 ,  , w_4491 );
buf ( w_4489 , \d[1]_b1 );
not ( w_4489 , w_4492 );
not (  , w_4493 );
and ( w_4492 , w_4493 , \d[1]_b0 );
or ( \1473_b1 , \a[0]_b1 , w_4495 );
not ( w_4495 , w_4496 );
and ( \1473_b0 , \a[0]_b0 , w_4497 );
and ( w_4496 ,  , w_4497 );
buf ( w_4495 , \d[2]_b1 );
not ( w_4495 , w_4498 );
not (  , w_4499 );
and ( w_4498 , w_4499 , \d[2]_b0 );
buf ( \1475_b1 , \1474_b1 );
not ( \1475_b1 , w_4500 );
not ( \1475_b0 , w_4501 );
and ( w_4500 , w_4501 , \1474_b0 );
or ( \1476_b1 , \1470_b1 , \1475_b1 );
not ( \1475_b1 , w_4502 );
and ( \1476_b0 , \1470_b0 , w_4503 );
and ( w_4502 , w_4503 , \1475_b0 );
buf ( \1477_b1 , \1470_b1 );
not ( \1477_b1 , w_4504 );
not ( \1477_b0 , w_4505 );
and ( w_4504 , w_4505 , \1470_b0 );
or ( \1478_b1 , \1477_b1 , \1474_b1 );
not ( \1474_b1 , w_4506 );
and ( \1478_b0 , \1477_b0 , w_4507 );
and ( w_4506 , w_4507 , \1474_b0 );
or ( \1479_b1 , \1476_b1 , w_4509 );
not ( w_4509 , w_4510 );
and ( \1479_b0 , \1476_b0 , w_4511 );
and ( w_4510 ,  , w_4511 );
buf ( w_4509 , \1478_b1 );
not ( w_4509 , w_4512 );
not (  , w_4513 );
and ( w_4512 , w_4513 , \1478_b0 );
buf ( \1480_b1 , \965_b1 );
not ( \1480_b1 , w_4514 );
not ( \1480_b0 , w_4515 );
and ( w_4514 , w_4515 , \965_b0 );
or ( \1481_b1 , \a[0]_b1 , \d[3]_b1 );
xor ( \1481_b0 , \a[0]_b0 , w_4516 );
not ( w_4516 , w_4517 );
and ( w_4517 , \d[3]_b1 , \d[3]_b0 );
or ( \1482_b1 , \961_b1 , w_4519 );
not ( w_4519 , w_4520 );
and ( \1482_b0 , \961_b0 , w_4521 );
and ( w_4520 ,  , w_4521 );
buf ( w_4519 , \1481_b1 );
not ( w_4519 , w_4522 );
not (  , w_4523 );
and ( w_4522 , w_4523 , \1481_b0 );
buf ( \1483_b1 , \1482_b1 );
not ( \1483_b1 , w_4524 );
not ( \1483_b0 , w_4525 );
and ( w_4524 , w_4525 , \1482_b0 );
or ( \1484_b1 , \1480_b1 , \1483_b1 );
not ( \1483_b1 , w_4526 );
and ( \1484_b0 , \1480_b0 , w_4527 );
and ( w_4526 , w_4527 , \1483_b0 );
or ( \1485_b1 , \965_b1 , \1446_b1 );
not ( \1446_b1 , w_4528 );
and ( \1485_b0 , \965_b0 , w_4529 );
and ( w_4528 , w_4529 , \1446_b0 );
or ( \1486_b1 , \1484_b1 , w_4531 );
not ( w_4531 , w_4532 );
and ( \1486_b0 , \1484_b0 , w_4533 );
and ( w_4532 ,  , w_4533 );
buf ( w_4531 , \1485_b1 );
not ( w_4531 , w_4534 );
not (  , w_4535 );
and ( w_4534 , w_4535 , \1485_b0 );
or ( \1487_b1 , \1479_b1 , w_4536 );
or ( \1487_b0 , \1479_b0 , \1486_b0 );
not ( \1486_b0 , w_4537 );
and ( w_4537 , w_4536 , \1486_b1 );
or ( \1488_b1 , \1479_b1 , w_4539 );
not ( w_4539 , w_4540 );
and ( \1488_b0 , \1479_b0 , w_4541 );
and ( w_4540 ,  , w_4541 );
buf ( w_4539 , \1486_b1 );
not ( w_4539 , w_4542 );
not (  , w_4543 );
and ( w_4542 , w_4543 , \1486_b0 );
or ( \1489_b1 , \d[1]_b1 , \a[1]_b1 );
xor ( \1489_b0 , \d[1]_b0 , w_4544 );
not ( w_4544 , w_4545 );
and ( w_4545 , \a[1]_b1 , \a[1]_b0 );
buf ( \1490_b1 , \1489_b1 );
not ( \1490_b1 , w_4546 );
not ( \1490_b0 , w_4547 );
and ( w_4546 , w_4547 , \1489_b0 );
buf ( \1491_b1 , \1012_b1 );
not ( \1491_b1 , w_4548 );
not ( \1491_b0 , w_4549 );
and ( w_4548 , w_4549 , \1012_b0 );
or ( \1492_b1 , \1490_b1 , w_4550 );
or ( \1492_b0 , \1490_b0 , \1491_b0 );
not ( \1491_b0 , w_4551 );
and ( w_4551 , w_4550 , \1491_b1 );
or ( \1493_b1 , \1467_b1 , w_4553 );
not ( w_4553 , w_4554 );
and ( \1493_b0 , \1467_b0 , w_4555 );
and ( w_4554 ,  , w_4555 );
buf ( w_4553 , \d[0]_b1 );
not ( w_4553 , w_4556 );
not (  , w_4557 );
and ( w_4556 , w_4557 , \d[0]_b0 );
or ( \1494_b1 , \1492_b1 , w_4559 );
not ( w_4559 , w_4560 );
and ( \1494_b0 , \1492_b0 , w_4561 );
and ( w_4560 ,  , w_4561 );
buf ( w_4559 , \1493_b1 );
not ( w_4559 , w_4562 );
not (  , w_4563 );
and ( w_4562 , w_4563 , \1493_b0 );
or ( \1495_b1 , \959_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_4564 );
and ( \1495_b0 , \959_b0 , w_4565 );
and ( w_4564 , w_4565 , \a[0]_b0 );
or ( \1496_b1 , \1494_b1 , w_4567 );
not ( w_4567 , w_4568 );
and ( \1496_b0 , \1494_b0 , w_4569 );
and ( w_4568 ,  , w_4569 );
buf ( w_4567 , \1495_b1 );
not ( w_4567 , w_4570 );
not (  , w_4571 );
and ( w_4570 , w_4571 , \1495_b0 );
or ( \1497_b1 , \a[0]_b1 , \d[1]_b1 );
xor ( \1497_b0 , \a[0]_b0 , w_4572 );
not ( w_4572 , w_4573 );
and ( w_4573 , \d[1]_b1 , \d[1]_b0 );
buf ( \1498_b1 , \1497_b1 );
not ( \1498_b1 , w_4574 );
not ( \1498_b0 , w_4575 );
and ( w_4574 , w_4575 , \1497_b0 );
buf ( \1499_b1 , \1012_b1 );
not ( \1499_b1 , w_4576 );
not ( \1499_b0 , w_4577 );
and ( w_4576 , w_4577 , \1012_b0 );
or ( \1500_b1 , \1498_b1 , w_4578 );
or ( \1500_b0 , \1498_b0 , \1499_b0 );
not ( \1499_b0 , w_4579 );
and ( w_4579 , w_4578 , \1499_b1 );
or ( \1501_b1 , \1489_b1 , w_4581 );
not ( w_4581 , w_4582 );
and ( \1501_b0 , \1489_b0 , w_4583 );
and ( w_4582 ,  , w_4583 );
buf ( w_4581 , \d[0]_b1 );
not ( w_4581 , w_4584 );
not (  , w_4585 );
and ( w_4584 , w_4585 , \d[0]_b0 );
or ( \1502_b1 , \1500_b1 , w_4587 );
not ( w_4587 , w_4588 );
and ( \1502_b0 , \1500_b0 , w_4589 );
and ( w_4588 ,  , w_4589 );
buf ( w_4587 , \1501_b1 );
not ( w_4587 , w_4590 );
not (  , w_4591 );
and ( w_4590 , w_4591 , \1501_b0 );
or ( \1503_b1 , \684_b1 , \d[1]_b1 );
not ( \d[1]_b1 , w_4592 );
and ( \1503_b0 , \684_b0 , w_4593 );
and ( w_4592 , w_4593 , \d[1]_b0 );
or ( \1504_b1 , \1502_b1 , w_4595 );
not ( w_4595 , w_4596 );
and ( \1504_b0 , \1502_b0 , w_4597 );
and ( w_4596 ,  , w_4597 );
buf ( w_4595 , \1503_b1 );
not ( w_4595 , w_4598 );
not (  , w_4599 );
and ( w_4598 , w_4599 , \1503_b0 );
or ( \1505_b1 , \1496_b1 , w_4600 );
or ( \1505_b0 , \1496_b0 , \1504_b0 );
not ( \1504_b0 , w_4601 );
and ( w_4601 , w_4600 , \1504_b1 );
or ( \1506_b1 , \1494_b1 , w_4603 );
not ( w_4603 , w_4604 );
and ( \1506_b0 , \1494_b0 , w_4605 );
and ( w_4604 ,  , w_4605 );
buf ( w_4603 , \1495_b1 );
not ( w_4603 , w_4606 );
not (  , w_4607 );
and ( w_4606 , w_4607 , \1495_b0 );
or ( \1507_b1 , \1505_b1 , w_4609 );
not ( w_4609 , w_4610 );
and ( \1507_b0 , \1505_b0 , w_4611 );
and ( w_4610 ,  , w_4611 );
buf ( w_4609 , \1506_b1 );
not ( w_4609 , w_4612 );
not (  , w_4613 );
and ( w_4612 , w_4613 , \1506_b0 );
or ( \1508_b1 , \1488_b1 , w_4615 );
not ( w_4615 , w_4616 );
and ( \1508_b0 , \1488_b0 , w_4617 );
and ( w_4616 ,  , w_4617 );
buf ( w_4615 , \1507_b1 );
not ( w_4615 , w_4618 );
not (  , w_4619 );
and ( w_4618 , w_4619 , \1507_b0 );
or ( \1509_b1 , \1487_b1 , w_4621 );
not ( w_4621 , w_4622 );
and ( \1509_b0 , \1487_b0 , w_4623 );
and ( w_4622 ,  , w_4623 );
buf ( w_4621 , \1508_b1 );
not ( w_4621 , w_4624 );
not (  , w_4625 );
and ( w_4624 , w_4625 , \1508_b0 );
or ( \1510_b1 , \1459_b1 , \1450_b1 );
xor ( \1510_b0 , \1459_b0 , w_4626 );
not ( w_4626 , w_4627 );
and ( w_4627 , \1450_b1 , \1450_b0 );
or ( \1511_b1 , \1510_b1 , \1457_b1 );
xor ( \1511_b0 , \1510_b0 , w_4628 );
not ( w_4628 , w_4629 );
and ( w_4629 , \1457_b1 , \1457_b0 );
buf ( \1512_b1 , \1470_b1 );
not ( \1512_b1 , w_4630 );
not ( \1512_b0 , w_4631 );
and ( w_4630 , w_4631 , \1470_b0 );
or ( \1513_b1 , \1512_b1 , w_4633 );
not ( w_4633 , w_4634 );
and ( \1513_b0 , \1512_b0 , w_4635 );
and ( w_4634 ,  , w_4635 );
buf ( w_4633 , \1475_b1 );
not ( w_4633 , w_4636 );
not (  , w_4637 );
and ( w_4636 , w_4637 , \1475_b0 );
or ( \1514_b1 , \1511_b1 , w_4639 );
not ( w_4639 , w_4640 );
and ( \1514_b0 , \1511_b0 , w_4641 );
and ( w_4640 ,  , w_4641 );
buf ( w_4639 , \1513_b1 );
not ( w_4639 , w_4642 );
not (  , w_4643 );
and ( w_4642 , w_4643 , \1513_b0 );
or ( \1515_b1 , \1509_b1 , \1514_b1 );
not ( \1514_b1 , w_4644 );
and ( \1515_b0 , \1509_b0 , w_4645 );
and ( w_4644 , w_4645 , \1514_b0 );
or ( \1516_b1 , \1511_b1 , w_4647 );
not ( w_4647 , w_4648 );
and ( \1516_b0 , \1511_b0 , w_4649 );
and ( w_4648 ,  , w_4649 );
buf ( w_4647 , \1513_b1 );
not ( w_4647 , w_4650 );
not (  , w_4651 );
and ( w_4650 , w_4651 , \1513_b0 );
or ( \1517_b1 , \1515_b1 , w_4653 );
not ( w_4653 , w_4654 );
and ( \1517_b0 , \1515_b0 , w_4655 );
and ( w_4654 ,  , w_4655 );
buf ( w_4653 , \1516_b1 );
not ( w_4653 , w_4656 );
not (  , w_4657 );
and ( w_4656 , w_4657 , \1516_b0 );
or ( \1518_b1 , \1466_b1 , w_4658 );
or ( \1518_b0 , \1466_b0 , \1517_b0 );
not ( \1517_b0 , w_4659 );
and ( w_4659 , w_4658 , \1517_b1 );
or ( \1519_b1 , \1445_b1 , w_4661 );
not ( w_4661 , w_4662 );
and ( \1519_b0 , \1445_b0 , w_4663 );
and ( w_4662 ,  , w_4663 );
buf ( w_4661 , \1465_b1 );
not ( w_4661 , w_4664 );
not (  , w_4665 );
and ( w_4664 , w_4665 , \1465_b0 );
or ( \1520_b1 , \1518_b1 , w_4667 );
not ( w_4667 , w_4668 );
and ( \1520_b0 , \1518_b0 , w_4669 );
and ( w_4668 ,  , w_4669 );
buf ( w_4667 , \1519_b1 );
not ( w_4667 , w_4670 );
not (  , w_4671 );
and ( w_4670 , w_4671 , \1519_b0 );
or ( \1521_b1 , \1443_b1 , \1520_b1 );
not ( \1520_b1 , w_4672 );
and ( \1521_b0 , \1443_b0 , w_4673 );
and ( w_4672 , w_4673 , \1520_b0 );
or ( \1522_b1 , \1440_b1 , \1442_b1 );
not ( \1442_b1 , w_4674 );
and ( \1522_b0 , \1440_b0 , w_4675 );
and ( w_4674 , w_4675 , \1442_b0 );
or ( \1523_b1 , \1521_b1 , w_4676 );
or ( \1523_b0 , \1521_b0 , \1522_b0 );
not ( \1522_b0 , w_4677 );
and ( w_4677 , w_4676 , \1522_b1 );
buf ( \1524_b1 , \1523_b1 );
not ( \1524_b1 , w_4678 );
not ( \1524_b0 , w_4679 );
and ( w_4678 , w_4679 , \1523_b0 );
or ( \1525_b1 , \1418_b1 , w_4680 );
or ( \1525_b0 , \1418_b0 , \1524_b0 );
not ( \1524_b0 , w_4681 );
and ( w_4681 , w_4680 , \1524_b1 );
or ( \1526_b1 , \1390_b1 , w_4682 );
or ( \1526_b0 , \1390_b0 , \1416_b0 );
not ( \1416_b0 , w_4683 );
and ( w_4683 , w_4682 , \1416_b1 );
or ( \1527_b1 , \1525_b1 , w_4685 );
not ( w_4685 , w_4686 );
and ( \1527_b0 , \1525_b0 , w_4687 );
and ( w_4686 ,  , w_4687 );
buf ( w_4685 , \1526_b1 );
not ( w_4685 , w_4688 );
not (  , w_4689 );
and ( w_4688 , w_4689 , \1526_b0 );
buf ( \1528_b1 , \1527_b1 );
buf ( \1528_b0 , \1527_b0 );
or ( \1530_b1 , \1160_b1 , w_4691 );
not ( w_4691 , w_4692 );
and ( \1530_b0 , \1160_b0 , w_4693 );
and ( w_4692 ,  , w_4693 );
buf ( w_4691 , \1126_b1 );
not ( w_4691 , w_4694 );
not (  , w_4695 );
and ( w_4694 , w_4695 , \1126_b0 );
or ( \1531_b1 , \1388_b1 , w_4697 );
not ( w_4697 , w_4698 );
and ( \1531_b0 , \1388_b0 , w_4699 );
and ( w_4698 ,  , w_4699 );
buf ( w_4697 , \1530_b1 );
not ( w_4697 , w_4700 );
not (  , w_4701 );
and ( w_4700 , w_4701 , \1530_b0 );
buf ( \1532_b1 , \1260_b1 );
not ( \1532_b1 , w_4702 );
not ( \1532_b0 , w_4703 );
and ( w_4702 , w_4703 , \1260_b0 );
buf ( \1533_b1 , \1286_b1 );
not ( \1533_b1 , w_4704 );
not ( \1533_b0 , w_4705 );
and ( w_4704 , w_4705 , \1286_b0 );
or ( \1534_b1 , \1532_b1 , w_4707 );
not ( w_4707 , w_4708 );
and ( \1534_b0 , \1532_b0 , w_4709 );
and ( w_4708 ,  , w_4709 );
buf ( w_4707 , \1533_b1 );
not ( w_4707 , w_4710 );
not (  , w_4711 );
and ( w_4710 , w_4711 , \1533_b0 );
or ( \1535_b1 , \1308_b1 , w_4712 );
or ( \1535_b0 , \1308_b0 , \1534_b0 );
not ( \1534_b0 , w_4713 );
and ( w_4713 , w_4712 , \1534_b1 );
or ( \1536_b1 , \1307_b1 , w_4715 );
not ( w_4715 , w_4716 );
and ( \1536_b0 , \1307_b0 , w_4717 );
and ( w_4716 ,  , w_4717 );
buf ( w_4715 , \1296_b1 );
not ( w_4715 , w_4718 );
not (  , w_4719 );
and ( w_4718 , w_4719 , \1296_b0 );
or ( \1537_b1 , \1535_b1 , w_4721 );
not ( w_4721 , w_4722 );
and ( \1537_b0 , \1535_b0 , w_4723 );
and ( w_4722 ,  , w_4723 );
buf ( w_4721 , \1536_b1 );
not ( w_4721 , w_4724 );
not (  , w_4725 );
and ( w_4724 , w_4725 , \1536_b0 );
or ( \1538_b1 , \1163_b1 , w_4727 );
not ( w_4727 , w_4728 );
and ( \1538_b0 , \1163_b0 , w_4729 );
and ( w_4728 ,  , w_4729 );
buf ( w_4727 , \1213_b1 );
not ( w_4727 , w_4730 );
not (  , w_4731 );
and ( w_4730 , w_4731 , \1213_b0 );
or ( \1539_b1 , \1537_b1 , w_4733 );
not ( w_4733 , w_4734 );
and ( \1539_b0 , \1537_b0 , w_4735 );
and ( w_4734 ,  , w_4735 );
buf ( w_4733 , \1538_b1 );
not ( w_4733 , w_4736 );
not (  , w_4737 );
and ( w_4736 , w_4737 , \1538_b0 );
buf ( \1540_b1 , \1539_b1 );
not ( \1540_b1 , w_4738 );
not ( \1540_b0 , w_4739 );
and ( w_4738 , w_4739 , \1539_b0 );
buf ( \1541_b1 , \1161_b1 );
buf ( \1541_b0 , \1161_b0 );
or ( \1543_b1 , \1382_b1 , w_4741 );
not ( w_4741 , w_4742 );
and ( \1543_b0 , \1382_b0 , w_4743 );
and ( w_4742 ,  , w_4743 );
buf ( w_4741 , \1386_b1 );
not ( w_4741 , w_4744 );
not (  , w_4745 );
and ( w_4744 , w_4745 , \1386_b0 );
buf ( \1545_b1 , \1361_b1 );
not ( \1545_b1 , w_4746 );
not ( \1545_b0 , w_4747 );
and ( w_4746 , w_4747 , \1361_b0 );
buf ( \1546_b1 , \1065_b1 );
not ( \1546_b1 , w_4748 );
not ( \1546_b0 , w_4749 );
and ( w_4748 , w_4749 , \1065_b0 );
or ( \1547_b1 , \1545_b1 , w_4750 );
or ( \1547_b0 , \1545_b0 , \1546_b0 );
not ( \1546_b0 , w_4751 );
and ( w_4751 , w_4750 , \1546_b1 );
or ( \1548_b1 , \a[13]_b1 , \d[1]_b1 );
xor ( \1548_b0 , \a[13]_b0 , w_4752 );
not ( w_4752 , w_4753 );
and ( w_4753 , \d[1]_b1 , \d[1]_b0 );
or ( \1549_b1 , \1548_b1 , w_4755 );
not ( w_4755 , w_4756 );
and ( \1549_b0 , \1548_b0 , w_4757 );
and ( w_4756 ,  , w_4757 );
buf ( w_4755 , \d[0]_b1 );
not ( w_4755 , w_4758 );
not (  , w_4759 );
and ( w_4758 , w_4759 , \d[0]_b0 );
or ( \1550_b1 , \1547_b1 , w_4761 );
not ( w_4761 , w_4762 );
and ( \1550_b0 , \1547_b0 , w_4763 );
and ( w_4762 ,  , w_4763 );
buf ( w_4761 , \1549_b1 );
not ( w_4761 , w_4764 );
not (  , w_4765 );
and ( w_4764 , w_4765 , \1549_b0 );
buf ( \1551_b1 , \1550_b1 );
not ( \1551_b1 , w_4766 );
not ( \1551_b0 , w_4767 );
and ( w_4766 , w_4767 , \1550_b0 );
or ( \1552_b1 , \a[0]_b1 , w_4768 );
or ( \1552_b0 , \a[0]_b0 , \d[12]_b0 );
not ( \d[12]_b0 , w_4769 );
and ( w_4769 , w_4768 , \d[12]_b1 );
or ( \1553_b1 , \1552_b1 , w_4771 );
not ( w_4771 , w_4772 );
and ( \1553_b0 , \1552_b0 , w_4773 );
and ( w_4772 ,  , w_4773 );
buf ( w_4771 , \d[11]_b1 );
not ( w_4771 , w_4774 );
not (  , w_4775 );
and ( w_4774 , w_4775 , \d[11]_b0 );
or ( \1554_b1 , \a[0]_b1 , w_4777 );
not ( w_4777 , w_4778 );
and ( \1554_b0 , \a[0]_b0 , w_4779 );
and ( w_4778 ,  , w_4779 );
buf ( w_4777 , \d[12]_b1 );
not ( w_4777 , w_4780 );
not (  , w_4781 );
and ( w_4780 , w_4781 , \d[12]_b0 );
buf ( \1556_b1 , \1555_b1 );
not ( \1556_b1 , w_4782 );
not ( \1556_b0 , w_4783 );
and ( w_4782 , w_4783 , \1555_b0 );
or ( \1557_b1 , \1551_b1 , \1556_b1 );
not ( \1556_b1 , w_4784 );
and ( \1557_b0 , \1551_b0 , w_4785 );
and ( w_4784 , w_4785 , \1556_b0 );
or ( \1558_b1 , \1550_b1 , \1555_b1 );
not ( \1555_b1 , w_4786 );
and ( \1558_b0 , \1550_b0 , w_4787 );
and ( w_4786 , w_4787 , \1555_b0 );
or ( \1559_b1 , \1557_b1 , w_4789 );
not ( w_4789 , w_4790 );
and ( \1559_b0 , \1557_b0 , w_4791 );
and ( w_4790 ,  , w_4791 );
buf ( w_4789 , \1558_b1 );
not ( w_4789 , w_4792 );
not (  , w_4793 );
and ( w_4792 , w_4793 , \1558_b0 );
or ( \1560_b1 , \1336_b1 , \1342_b1 );
xor ( \1560_b0 , \1336_b0 , w_4794 );
not ( w_4794 , w_4795 );
and ( w_4795 , \1342_b1 , \1342_b0 );
or ( \1561_b1 , \1560_b1 , \1349_b1 );
not ( \1349_b1 , w_4796 );
and ( \1561_b0 , \1560_b0 , w_4797 );
and ( w_4796 , w_4797 , \1349_b0 );
or ( \1562_b1 , \1336_b1 , \1342_b1 );
not ( \1342_b1 , w_4798 );
and ( \1562_b0 , \1336_b0 , w_4799 );
and ( w_4798 , w_4799 , \1342_b0 );
or ( \1563_b1 , \1561_b1 , w_4800 );
or ( \1563_b0 , \1561_b0 , \1562_b0 );
not ( \1562_b0 , w_4801 );
and ( w_4801 , w_4800 , \1562_b1 );
or ( \1564_b1 , \1559_b1 , \1563_b1 );
xor ( \1564_b0 , \1559_b0 , w_4802 );
not ( w_4802 , w_4803 );
and ( w_4803 , \1563_b1 , \1563_b0 );
or ( \1565_b1 , \1357_b1 , w_4804 );
or ( \1565_b0 , \1357_b0 , \1363_b0 );
not ( \1363_b0 , w_4805 );
and ( w_4805 , w_4804 , \1363_b1 );
or ( \1566_b1 , \1565_b1 , \1371_b1 );
not ( \1371_b1 , w_4806 );
and ( \1566_b0 , \1565_b0 , w_4807 );
and ( w_4806 , w_4807 , \1371_b0 );
or ( \1567_b1 , \1357_b1 , \1363_b1 );
not ( \1363_b1 , w_4808 );
and ( \1567_b0 , \1357_b0 , w_4809 );
and ( w_4808 , w_4809 , \1363_b0 );
or ( \1568_b1 , \1566_b1 , w_4811 );
not ( w_4811 , w_4812 );
and ( \1568_b0 , \1566_b0 , w_4813 );
and ( w_4812 ,  , w_4813 );
buf ( w_4811 , \1567_b1 );
not ( w_4811 , w_4814 );
not (  , w_4815 );
and ( w_4814 , w_4815 , \1567_b0 );
buf ( \1569_b1 , \1568_b1 );
not ( \1569_b1 , w_4816 );
not ( \1569_b0 , w_4817 );
and ( w_4816 , w_4817 , \1568_b0 );
or ( \1570_b1 , \1564_b1 , \1569_b1 );
xor ( \1570_b0 , \1564_b0 , w_4818 );
not ( w_4818 , w_4819 );
and ( w_4819 , \1569_b1 , \1569_b0 );
buf ( \1571_b1 , \1570_b1 );
not ( \1571_b1 , w_4820 );
not ( \1571_b0 , w_4821 );
and ( w_4820 , w_4821 , \1570_b0 );
or ( \1572_b1 , \1350_b1 , \1372_b1 );
xor ( \1572_b0 , \1350_b0 , w_4822 );
not ( w_4822 , w_4823 );
and ( w_4823 , \1372_b1 , \1372_b0 );
or ( \1573_b1 , \1572_b1 , \1380_b1 );
not ( \1380_b1 , w_4824 );
and ( \1573_b0 , \1572_b0 , w_4825 );
and ( w_4824 , w_4825 , \1380_b0 );
or ( \1574_b1 , \1350_b1 , \1372_b1 );
not ( \1372_b1 , w_4826 );
and ( \1574_b0 , \1350_b0 , w_4827 );
and ( w_4826 , w_4827 , \1372_b0 );
or ( \1575_b1 , \1573_b1 , w_4828 );
or ( \1575_b0 , \1573_b0 , \1574_b0 );
not ( \1574_b0 , w_4829 );
and ( w_4829 , w_4828 , \1574_b1 );
buf ( \1576_b1 , \1575_b1 );
not ( \1576_b1 , w_4830 );
not ( \1576_b0 , w_4831 );
and ( w_4830 , w_4831 , \1575_b0 );
or ( \1577_b1 , \1571_b1 , w_4832 );
or ( \1577_b0 , \1571_b0 , \1576_b0 );
not ( \1576_b0 , w_4833 );
and ( w_4833 , w_4832 , \1576_b1 );
or ( \1578_b1 , \1575_b1 , w_4834 );
or ( \1578_b0 , \1575_b0 , \1570_b0 );
not ( \1570_b0 , w_4835 );
and ( w_4835 , w_4834 , \1570_b1 );
or ( \1579_b1 , \1577_b1 , w_4837 );
not ( w_4837 , w_4838 );
and ( \1579_b0 , \1577_b0 , w_4839 );
and ( w_4838 ,  , w_4839 );
buf ( w_4837 , \1578_b1 );
not ( w_4837 , w_4840 );
not (  , w_4841 );
and ( w_4840 , w_4841 , \1578_b0 );
or ( \1580_b1 , \a[0]_b1 , \d[13]_b1 );
xor ( \1580_b0 , \a[0]_b0 , w_4842 );
not ( w_4842 , w_4843 );
and ( w_4843 , \d[13]_b1 , \d[13]_b0 );
buf ( \1581_b1 , \1580_b1 );
not ( \1581_b1 , w_4844 );
not ( \1581_b0 , w_4845 );
and ( w_4844 , w_4845 , \1580_b0 );
or ( \1582_b1 , \d[13]_b1 , w_4846 );
xor ( \1582_b0 , \d[13]_b0 , w_4848 );
not ( w_4848 , w_4849 );
and ( w_4849 , w_4846 , w_4847 );
buf ( w_4846 , \d[12]_b1 );
not ( w_4846 , w_4850 );
not ( w_4847 , w_4851 );
and ( w_4850 , w_4851 , \d[12]_b0 );
or ( \1583_b1 , \1582_b1 , w_4853 );
not ( w_4853 , w_4854 );
and ( \1583_b0 , \1582_b0 , w_4855 );
and ( w_4854 ,  , w_4855 );
buf ( w_4853 , \1335_b1 );
not ( w_4853 , w_4856 );
not (  , w_4857 );
and ( w_4856 , w_4857 , \1335_b0 );
buf ( \1584_b1 , \1583_b1 );
not ( \1584_b1 , w_4858 );
not ( \1584_b0 , w_4859 );
and ( w_4858 , w_4859 , \1583_b0 );
or ( \1585_b1 , \1581_b1 , w_4860 );
or ( \1585_b0 , \1581_b0 , \1584_b0 );
not ( \1584_b0 , w_4861 );
and ( w_4861 , w_4860 , \1584_b1 );
or ( \1586_b1 , \a[1]_b1 , \d[13]_b1 );
xor ( \1586_b0 , \a[1]_b0 , w_4862 );
not ( w_4862 , w_4863 );
and ( w_4863 , \d[13]_b1 , \d[13]_b0 );
or ( \1587_b1 , \1335_b1 , w_4865 );
not ( w_4865 , w_4866 );
and ( \1587_b0 , \1335_b0 , w_4867 );
and ( w_4866 ,  , w_4867 );
buf ( w_4865 , \1586_b1 );
not ( w_4865 , w_4868 );
not (  , w_4869 );
and ( w_4868 , w_4869 , \1586_b0 );
or ( \1588_b1 , \1585_b1 , w_4871 );
not ( w_4871 , w_4872 );
and ( \1588_b0 , \1585_b0 , w_4873 );
and ( w_4872 ,  , w_4873 );
buf ( w_4871 , \1587_b1 );
not ( w_4871 , w_4874 );
not (  , w_4875 );
and ( w_4874 , w_4875 , \1587_b0 );
buf ( \1589_b1 , \1369_b1 );
not ( \1589_b1 , w_4876 );
not ( \1589_b0 , w_4877 );
and ( w_4876 , w_4877 , \1369_b0 );
buf ( \1590_b1 , \944_b1 );
not ( \1590_b1 , w_4878 );
not ( \1590_b0 , w_4879 );
and ( w_4878 , w_4879 , \944_b0 );
or ( \1591_b1 , \1589_b1 , w_4880 );
or ( \1591_b0 , \1589_b0 , \1590_b0 );
not ( \1590_b0 , w_4881 );
and ( w_4881 , w_4880 , \1590_b1 );
or ( \1592_b1 , \a[3]_b1 , \d[11]_b1 );
xor ( \1592_b0 , \a[3]_b0 , w_4882 );
not ( w_4882 , w_4883 );
and ( w_4883 , \d[11]_b1 , \d[11]_b0 );
or ( \1593_b1 , \947_b1 , w_4885 );
not ( w_4885 , w_4886 );
and ( \1593_b0 , \947_b0 , w_4887 );
and ( w_4886 ,  , w_4887 );
buf ( w_4885 , \1592_b1 );
not ( w_4885 , w_4888 );
not (  , w_4889 );
and ( w_4888 , w_4889 , \1592_b0 );
or ( \1594_b1 , \1591_b1 , w_4891 );
not ( w_4891 , w_4892 );
and ( \1594_b0 , \1591_b0 , w_4893 );
and ( w_4892 ,  , w_4893 );
buf ( w_4891 , \1593_b1 );
not ( w_4891 , w_4894 );
not (  , w_4895 );
and ( w_4894 , w_4895 , \1593_b0 );
or ( \1595_b1 , \1588_b1 , \1594_b1 );
xor ( \1595_b0 , \1588_b0 , w_4896 );
not ( w_4896 , w_4897 );
and ( w_4897 , \1594_b1 , \1594_b0 );
buf ( \1596_b1 , \1315_b1 );
not ( \1596_b1 , w_4898 );
not ( \1596_b0 , w_4899 );
and ( w_4898 , w_4899 , \1315_b0 );
buf ( \1597_b1 , \933_b1 );
not ( \1597_b1 , w_4900 );
not ( \1597_b0 , w_4901 );
and ( w_4900 , w_4901 , \933_b0 );
or ( \1598_b1 , \1596_b1 , w_4902 );
or ( \1598_b0 , \1596_b0 , \1597_b0 );
not ( \1597_b0 , w_4903 );
and ( w_4903 , w_4902 , \1597_b1 );
or ( \1599_b1 , \a[9]_b1 , \d[5]_b1 );
xor ( \1599_b0 , \a[9]_b0 , w_4904 );
not ( w_4904 , w_4905 );
and ( w_4905 , \d[5]_b1 , \d[5]_b0 );
or ( \1600_b1 , \936_b1 , w_4907 );
not ( w_4907 , w_4908 );
and ( \1600_b0 , \936_b0 , w_4909 );
and ( w_4908 ,  , w_4909 );
buf ( w_4907 , \1599_b1 );
not ( w_4907 , w_4910 );
not (  , w_4911 );
and ( w_4910 , w_4911 , \1599_b0 );
or ( \1601_b1 , \1598_b1 , w_4913 );
not ( w_4913 , w_4914 );
and ( \1601_b0 , \1598_b0 , w_4915 );
and ( w_4914 ,  , w_4915 );
buf ( w_4913 , \1600_b1 );
not ( w_4913 , w_4916 );
not (  , w_4917 );
and ( w_4916 , w_4917 , \1600_b0 );
or ( \1602_b1 , \1595_b1 , \1601_b1 );
xor ( \1602_b0 , \1595_b0 , w_4918 );
not ( w_4918 , w_4919 );
and ( w_4919 , \1601_b1 , \1601_b0 );
buf ( \1603_b1 , \1602_b1 );
not ( \1603_b1 , w_4920 );
not ( \1603_b0 , w_4921 );
and ( w_4920 , w_4921 , \1602_b0 );
buf ( \1604_b1 , \1603_b1 );
not ( \1604_b1 , w_4922 );
not ( \1604_b0 , w_4923 );
and ( w_4922 , w_4923 , \1603_b0 );
buf ( \1605_b1 , \1110_b1 );
not ( \1605_b1 , w_4924 );
not ( \1605_b0 , w_4925 );
and ( w_4924 , w_4925 , \1110_b0 );
buf ( \1606_b1 , \1354_b1 );
not ( \1606_b1 , w_4926 );
not ( \1606_b0 , w_4927 );
and ( w_4926 , w_4927 , \1354_b0 );
or ( \1607_b1 , \1605_b1 , \1606_b1 );
not ( \1606_b1 , w_4928 );
and ( \1607_b0 , \1605_b0 , w_4929 );
and ( w_4928 , w_4929 , \1606_b0 );
or ( \1608_b1 , \a[5]_b1 , \d[9]_b1 );
xor ( \1608_b0 , \a[5]_b0 , w_4930 );
not ( w_4930 , w_4931 );
and ( w_4931 , \d[9]_b1 , \d[9]_b0 );
or ( \1609_b1 , \1058_b1 , \1608_b1 );
not ( \1608_b1 , w_4932 );
and ( \1609_b0 , \1058_b0 , w_4933 );
and ( w_4932 , w_4933 , \1608_b0 );
or ( \1610_b1 , \1607_b1 , w_4935 );
not ( w_4935 , w_4936 );
and ( \1610_b0 , \1607_b0 , w_4937 );
and ( w_4936 ,  , w_4937 );
buf ( w_4935 , \1609_b1 );
not ( w_4935 , w_4938 );
not (  , w_4939 );
and ( w_4938 , w_4939 , \1609_b0 );
buf ( \1611_b1 , \1610_b1 );
not ( \1611_b1 , w_4940 );
not ( \1611_b0 , w_4941 );
and ( w_4940 , w_4941 , \1610_b0 );
buf ( \1612_b1 , \1611_b1 );
not ( \1612_b1 , w_4942 );
not ( \1612_b0 , w_4943 );
and ( w_4942 , w_4943 , \1611_b0 );
buf ( \1613_b1 , \1340_b1 );
not ( \1613_b1 , w_4944 );
not ( \1613_b0 , w_4945 );
and ( w_4944 , w_4945 , \1340_b0 );
buf ( \1614_b1 , \999_b1 );
not ( \1614_b1 , w_4946 );
not ( \1614_b0 , w_4947 );
and ( w_4946 , w_4947 , \999_b0 );
or ( \1615_b1 , \1613_b1 , w_4948 );
or ( \1615_b0 , \1613_b0 , \1614_b0 );
not ( \1614_b0 , w_4949 );
and ( w_4949 , w_4948 , \1614_b1 );
or ( \1616_b1 , \a[7]_b1 , \d[7]_b1 );
xor ( \1616_b0 , \a[7]_b0 , w_4950 );
not ( w_4950 , w_4951 );
and ( w_4951 , \d[7]_b1 , \d[7]_b0 );
or ( \1617_b1 , \1003_b1 , w_4953 );
not ( w_4953 , w_4954 );
and ( \1617_b0 , \1003_b0 , w_4955 );
and ( w_4954 ,  , w_4955 );
buf ( w_4953 , \1616_b1 );
not ( w_4953 , w_4956 );
not (  , w_4957 );
and ( w_4956 , w_4957 , \1616_b0 );
or ( \1618_b1 , \1615_b1 , w_4959 );
not ( w_4959 , w_4960 );
and ( \1618_b0 , \1615_b0 , w_4961 );
and ( w_4960 ,  , w_4961 );
buf ( w_4959 , \1617_b1 );
not ( w_4959 , w_4962 );
not (  , w_4963 );
and ( w_4962 , w_4963 , \1617_b0 );
buf ( \1619_b1 , \1618_b1 );
not ( \1619_b1 , w_4964 );
not ( \1619_b0 , w_4965 );
and ( w_4964 , w_4965 , \1618_b0 );
buf ( \1620_b1 , \1619_b1 );
not ( \1620_b1 , w_4966 );
not ( \1620_b0 , w_4967 );
and ( w_4966 , w_4967 , \1619_b0 );
or ( \1621_b1 , \1612_b1 , w_4968 );
or ( \1621_b0 , \1612_b0 , \1620_b0 );
not ( \1620_b0 , w_4969 );
and ( w_4969 , w_4968 , \1620_b1 );
or ( \1622_b1 , \1610_b1 , w_4971 );
not ( w_4971 , w_4972 );
and ( \1622_b0 , \1610_b0 , w_4973 );
and ( w_4972 ,  , w_4973 );
buf ( w_4971 , \1618_b1 );
not ( w_4971 , w_4974 );
not (  , w_4975 );
and ( w_4974 , w_4975 , \1618_b0 );
or ( \1623_b1 , \1621_b1 , w_4977 );
not ( w_4977 , w_4978 );
and ( \1623_b0 , \1621_b0 , w_4979 );
and ( w_4978 ,  , w_4979 );
buf ( w_4977 , \1622_b1 );
not ( w_4977 , w_4980 );
not (  , w_4981 );
and ( w_4980 , w_4981 , \1622_b0 );
buf ( \1624_b1 , \1347_b1 );
not ( \1624_b1 , w_4982 );
not ( \1624_b0 , w_4983 );
and ( w_4982 , w_4983 , \1347_b0 );
buf ( \1625_b1 , \962_b1 );
not ( \1625_b1 , w_4984 );
not ( \1625_b0 , w_4985 );
and ( w_4984 , w_4985 , \962_b0 );
or ( \1626_b1 , \1624_b1 , w_4986 );
or ( \1626_b0 , \1624_b0 , \1625_b0 );
not ( \1625_b0 , w_4987 );
and ( w_4987 , w_4986 , \1625_b1 );
or ( \1627_b1 , \a[11]_b1 , \d[3]_b1 );
xor ( \1627_b0 , \a[11]_b0 , w_4988 );
not ( w_4988 , w_4989 );
and ( w_4989 , \d[3]_b1 , \d[3]_b0 );
or ( \1628_b1 , \965_b1 , w_4991 );
not ( w_4991 , w_4992 );
and ( \1628_b0 , \965_b0 , w_4993 );
and ( w_4992 ,  , w_4993 );
buf ( w_4991 , \1627_b1 );
not ( w_4991 , w_4994 );
not (  , w_4995 );
and ( w_4994 , w_4995 , \1627_b0 );
or ( \1629_b1 , \1626_b1 , w_4997 );
not ( w_4997 , w_4998 );
and ( \1629_b0 , \1626_b0 , w_4999 );
and ( w_4998 ,  , w_4999 );
buf ( w_4997 , \1628_b1 );
not ( w_4997 , w_5000 );
not (  , w_5001 );
and ( w_5000 , w_5001 , \1628_b0 );
or ( \1630_b1 , \1623_b1 , w_5002 );
xor ( \1630_b0 , \1623_b0 , w_5004 );
not ( w_5004 , w_5005 );
and ( w_5005 , w_5002 , w_5003 );
buf ( w_5002 , \1629_b1 );
not ( w_5002 , w_5006 );
not ( w_5003 , w_5007 );
and ( w_5006 , w_5007 , \1629_b0 );
buf ( \1631_b1 , \1630_b1 );
not ( \1631_b1 , w_5008 );
not ( \1631_b0 , w_5009 );
and ( w_5008 , w_5009 , \1630_b0 );
buf ( \1632_b1 , \1631_b1 );
not ( \1632_b1 , w_5010 );
not ( \1632_b0 , w_5011 );
and ( w_5010 , w_5011 , \1631_b0 );
or ( \1633_b1 , \1604_b1 , w_5012 );
or ( \1633_b0 , \1604_b0 , \1632_b0 );
not ( \1632_b0 , w_5013 );
and ( w_5013 , w_5012 , \1632_b1 );
or ( \1634_b1 , \1630_b1 , w_5015 );
not ( w_5015 , w_5016 );
and ( \1634_b0 , \1630_b0 , w_5017 );
and ( w_5016 ,  , w_5017 );
buf ( w_5015 , \1602_b1 );
not ( w_5015 , w_5018 );
not (  , w_5019 );
and ( w_5018 , w_5019 , \1602_b0 );
or ( \1635_b1 , \1633_b1 , w_5021 );
not ( w_5021 , w_5022 );
and ( \1635_b0 , \1633_b0 , w_5023 );
and ( w_5022 ,  , w_5023 );
buf ( w_5021 , \1634_b1 );
not ( w_5021 , w_5024 );
not (  , w_5025 );
and ( w_5024 , w_5025 , \1634_b0 );
or ( \1636_b1 , \1317_b1 , \1318_b1 );
xor ( \1636_b0 , \1317_b0 , w_5026 );
not ( w_5026 , w_5027 );
and ( w_5027 , \1318_b1 , \1318_b0 );
or ( \1637_b1 , \1636_b1 , \1325_b1 );
not ( \1325_b1 , w_5028 );
and ( \1637_b0 , \1636_b0 , w_5029 );
and ( w_5028 , w_5029 , \1325_b0 );
or ( \1638_b1 , \1317_b1 , \1318_b1 );
not ( \1318_b1 , w_5030 );
and ( \1638_b0 , \1317_b0 , w_5031 );
and ( w_5030 , w_5031 , \1318_b0 );
or ( \1639_b1 , \1637_b1 , w_5032 );
or ( \1639_b0 , \1637_b0 , \1638_b0 );
not ( \1638_b0 , w_5033 );
and ( w_5033 , w_5032 , \1638_b1 );
buf ( \1640_b1 , \1639_b1 );
not ( \1640_b1 , w_5034 );
not ( \1640_b0 , w_5035 );
and ( w_5034 , w_5035 , \1639_b0 );
or ( \1641_b1 , \1635_b1 , \1640_b1 );
not ( \1640_b1 , w_5036 );
and ( \1641_b0 , \1635_b0 , w_5037 );
and ( w_5036 , w_5037 , \1640_b0 );
buf ( \1642_b1 , \1635_b1 );
not ( \1642_b1 , w_5038 );
not ( \1642_b0 , w_5039 );
and ( w_5038 , w_5039 , \1635_b0 );
or ( \1643_b1 , \1642_b1 , \1639_b1 );
not ( \1639_b1 , w_5040 );
and ( \1643_b0 , \1642_b0 , w_5041 );
and ( w_5040 , w_5041 , \1639_b0 );
or ( \1644_b1 , \1641_b1 , w_5043 );
not ( w_5043 , w_5044 );
and ( \1644_b0 , \1641_b0 , w_5045 );
and ( w_5044 ,  , w_5045 );
buf ( w_5043 , \1643_b1 );
not ( w_5043 , w_5046 );
not (  , w_5047 );
and ( w_5046 , w_5047 , \1643_b0 );
or ( \1645_b1 , \1579_b1 , \1644_b1 );
not ( \1644_b1 , w_5048 );
and ( \1645_b0 , \1579_b0 , w_5049 );
and ( w_5048 , w_5049 , \1644_b0 );
buf ( \1646_b1 , \1579_b1 );
not ( \1646_b1 , w_5050 );
not ( \1646_b0 , w_5051 );
and ( w_5050 , w_5051 , \1579_b0 );
buf ( \1647_b1 , \1644_b1 );
not ( \1647_b1 , w_5052 );
not ( \1647_b0 , w_5053 );
and ( w_5052 , w_5053 , \1644_b0 );
or ( \1648_b1 , \1646_b1 , \1647_b1 );
not ( \1647_b1 , w_5054 );
and ( \1648_b0 , \1646_b0 , w_5055 );
and ( w_5054 , w_5055 , \1647_b0 );
or ( \1649_b1 , \1645_b1 , w_5057 );
not ( w_5057 , w_5058 );
and ( \1649_b0 , \1645_b0 , w_5059 );
and ( w_5058 ,  , w_5059 );
buf ( w_5057 , \1648_b1 );
not ( w_5057 , w_5060 );
not (  , w_5061 );
and ( w_5060 , w_5061 , \1648_b0 );
buf ( \1650_b1 , \1649_b1 );
not ( \1650_b1 , w_5062 );
not ( \1650_b0 , w_5063 );
and ( w_5062 , w_5063 , \1649_b0 );
or ( \1651_b1 , \1326_b1 , \1333_b1 );
xor ( \1651_b0 , \1326_b0 , w_5064 );
not ( w_5064 , w_5065 );
and ( w_5065 , \1333_b1 , \1333_b0 );
or ( \1652_b1 , \1651_b1 , \1381_b1 );
not ( \1381_b1 , w_5066 );
and ( \1652_b0 , \1651_b0 , w_5067 );
and ( w_5066 , w_5067 , \1381_b0 );
or ( \1653_b1 , \1326_b1 , \1333_b1 );
not ( \1333_b1 , w_5068 );
and ( \1653_b0 , \1326_b0 , w_5069 );
and ( w_5068 , w_5069 , \1333_b0 );
or ( \1654_b1 , \1652_b1 , w_5070 );
or ( \1654_b0 , \1652_b0 , \1653_b0 );
not ( \1653_b0 , w_5071 );
and ( w_5071 , w_5070 , \1653_b1 );
or ( \1655_b1 , \1650_b1 , w_5073 );
not ( w_5073 , w_5074 );
and ( \1655_b0 , \1650_b0 , w_5075 );
and ( w_5074 ,  , w_5075 );
buf ( w_5073 , \1654_b1 );
not ( w_5073 , w_5076 );
not (  , w_5077 );
and ( w_5076 , w_5077 , \1654_b0 );
buf ( \1656_b1 , \1654_b1 );
not ( \1656_b1 , w_5078 );
not ( \1656_b0 , w_5079 );
and ( w_5078 , w_5079 , \1654_b0 );
or ( \1657_b1 , \1656_b1 , w_5081 );
not ( w_5081 , w_5082 );
and ( \1657_b0 , \1656_b0 , w_5083 );
and ( w_5082 ,  , w_5083 );
buf ( w_5081 , \1649_b1 );
not ( w_5081 , w_5084 );
not (  , w_5085 );
and ( w_5084 , w_5085 , \1649_b0 );
or ( \1658_b1 , \1655_b1 , w_5087 );
not ( w_5087 , w_5088 );
and ( \1658_b0 , \1655_b0 , w_5089 );
and ( w_5088 ,  , w_5089 );
buf ( w_5087 , \1657_b1 );
not ( w_5087 , w_5090 );
not (  , w_5091 );
and ( w_5090 , w_5091 , \1657_b0 );
buf ( \1659_b1 , \1658_b1 );
not ( \1659_b1 , w_5092 );
not ( \1659_b0 , w_5093 );
and ( w_5092 , w_5093 , \1658_b0 );
or ( \1660_b1 , \1544_b1 , \1659_b1 );
not ( \1659_b1 , w_5094 );
and ( \1660_b0 , \1544_b0 , w_5095 );
and ( w_5094 , w_5095 , \1659_b0 );
buf ( \1661_b1 , \1544_b1 );
not ( \1661_b1 , w_5096 );
not ( \1661_b0 , w_5097 );
and ( w_5096 , w_5097 , \1544_b0 );
or ( \1662_b1 , \1661_b1 , \1658_b1 );
not ( \1658_b1 , w_5098 );
and ( \1662_b0 , \1661_b0 , w_5099 );
and ( w_5098 , w_5099 , \1658_b0 );
or ( \1663_b1 , \1660_b1 , w_5101 );
not ( w_5101 , w_5102 );
and ( \1663_b0 , \1660_b0 , w_5103 );
and ( w_5102 ,  , w_5103 );
buf ( w_5101 , \1662_b1 );
not ( w_5101 , w_5104 );
not (  , w_5105 );
and ( w_5104 , w_5105 , \1662_b0 );
or ( \1664_b1 , \239_b1 , w_5107 );
not ( w_5107 , w_5108 );
and ( \1664_b0 , \239_b0 , w_5109 );
and ( w_5108 ,  , w_5109 );
buf ( w_5107 , \343_b1 );
not ( w_5107 , w_5110 );
not (  , w_5111 );
and ( w_5110 , w_5111 , \343_b0 );
buf ( \1665_b1 , \339_b1 );
buf ( \1665_b0 , \339_b0 );
or ( \1666_b1 , \1664_b1 , w_5112 );
xor ( \1666_b0 , \1664_b0 , w_5114 );
not ( w_5114 , w_5115 );
and ( w_5115 , w_5112 , w_5113 );
buf ( w_5112 , \1665_b1 );
not ( w_5112 , w_5116 );
not ( w_5113 , w_5117 );
and ( w_5116 , w_5117 , \1665_b0 );
buf ( \1667_b1 , \1666_b1 );
not ( \1667_b1 , w_5118 );
not ( \1667_b0 , w_5119 );
and ( w_5118 , w_5119 , \1666_b0 );
buf ( \1668_b1 , \1667_b1 );
not ( \1668_b1 , w_5120 );
not ( \1668_b0 , w_5121 );
and ( w_5120 , w_5121 , \1667_b0 );
or ( \1669_b1 , \1663_b1 , w_5123 );
not ( w_5123 , w_5124 );
and ( \1669_b0 , \1663_b0 , w_5125 );
and ( w_5124 ,  , w_5125 );
buf ( w_5123 , \1668_b1 );
not ( w_5123 , w_5126 );
not (  , w_5127 );
and ( w_5126 , w_5127 , \1668_b0 );
or ( \1670_b1 , \c[5]_b1 , \b[6]_b1 );
xor ( \1670_b0 , \c[5]_b0 , w_5128 );
not ( w_5128 , w_5129 );
and ( w_5129 , \b[6]_b1 , \b[6]_b0 );
buf ( \1671_b1 , \1670_b1 );
not ( \1671_b1 , w_5130 );
not ( \1671_b0 , w_5131 );
and ( w_5130 , w_5131 , \1670_b0 );
or ( \1672_b1 , \c[5]_b1 , \c[4]_b1 );
xor ( \1672_b0 , \c[5]_b0 , w_5132 );
not ( w_5132 , w_5133 );
and ( w_5133 , \c[4]_b1 , \c[4]_b0 );
buf ( \1673_b1 , \1672_b1 );
not ( \1673_b1 , w_5134 );
not ( \1673_b0 , w_5135 );
and ( w_5134 , w_5135 , \1672_b0 );
or ( \1674_b1 , \c[4]_b1 , \c[3]_b1 );
xor ( \1674_b0 , \c[4]_b0 , w_5136 );
not ( w_5136 , w_5137 );
and ( w_5137 , \c[3]_b1 , \c[3]_b0 );
or ( \1675_b1 , \1673_b1 , w_5139 );
not ( w_5139 , w_5140 );
and ( \1675_b0 , \1673_b0 , w_5141 );
and ( w_5140 ,  , w_5141 );
buf ( w_5139 , \1674_b1 );
not ( w_5139 , w_5142 );
not (  , w_5143 );
and ( w_5142 , w_5143 , \1674_b0 );
buf ( \1676_b1 , \1675_b1 );
not ( \1676_b1 , w_5144 );
not ( \1676_b0 , w_5145 );
and ( w_5144 , w_5145 , \1675_b0 );
or ( \1677_b1 , \1671_b1 , w_5146 );
or ( \1677_b0 , \1671_b0 , \1676_b0 );
not ( \1676_b0 , w_5147 );
and ( w_5147 , w_5146 , \1676_b1 );
buf ( \1678_b1 , \1674_b1 );
buf ( \1678_b0 , \1674_b0 );
or ( \1679_b1 , \c[5]_b1 , \b[7]_b1 );
xor ( \1679_b0 , \c[5]_b0 , w_5148 );
not ( w_5148 , w_5149 );
and ( w_5149 , \b[7]_b1 , \b[7]_b0 );
or ( \1680_b1 , \1678_b1 , w_5151 );
not ( w_5151 , w_5152 );
and ( \1680_b0 , \1678_b0 , w_5153 );
and ( w_5152 ,  , w_5153 );
buf ( w_5151 , \1679_b1 );
not ( w_5151 , w_5154 );
not (  , w_5155 );
and ( w_5154 , w_5155 , \1679_b0 );
or ( \1681_b1 , \1677_b1 , w_5157 );
not ( w_5157 , w_5158 );
and ( \1681_b0 , \1677_b0 , w_5159 );
and ( w_5158 ,  , w_5159 );
buf ( w_5157 , \1680_b1 );
not ( w_5157 , w_5160 );
not (  , w_5161 );
and ( w_5160 , w_5161 , \1680_b0 );
or ( \1682_b1 , \b[0]_b1 , \c[11]_b1 );
xor ( \1682_b0 , \b[0]_b0 , w_5162 );
not ( w_5162 , w_5163 );
and ( w_5163 , \c[11]_b1 , \c[11]_b0 );
buf ( \1683_b1 , \1682_b1 );
not ( \1683_b1 , w_5164 );
not ( \1683_b0 , w_5165 );
and ( w_5164 , w_5165 , \1682_b0 );
or ( \1684_b1 , \c[11]_b1 , w_5166 );
xor ( \1684_b0 , \c[11]_b0 , w_5168 );
not ( w_5168 , w_5169 );
and ( w_5169 , w_5166 , w_5167 );
buf ( w_5166 , \c[10]_b1 );
not ( w_5166 , w_5170 );
not ( w_5167 , w_5171 );
and ( w_5170 , w_5171 , \c[10]_b0 );
or ( \1685_b1 , \c[10]_b1 , \c[9]_b1 );
xor ( \1685_b0 , \c[10]_b0 , w_5172 );
not ( w_5172 , w_5173 );
and ( w_5173 , \c[9]_b1 , \c[9]_b0 );
or ( \1686_b1 , \1684_b1 , w_5175 );
not ( w_5175 , w_5176 );
and ( \1686_b0 , \1684_b0 , w_5177 );
and ( w_5176 ,  , w_5177 );
buf ( w_5175 , \1685_b1 );
not ( w_5175 , w_5178 );
not (  , w_5179 );
and ( w_5178 , w_5179 , \1685_b0 );
buf ( \1687_b1 , \1686_b1 );
not ( \1687_b1 , w_5180 );
not ( \1687_b0 , w_5181 );
and ( w_5180 , w_5181 , \1686_b0 );
or ( \1688_b1 , \1683_b1 , w_5182 );
or ( \1688_b0 , \1683_b0 , \1687_b0 );
not ( \1687_b0 , w_5183 );
and ( w_5183 , w_5182 , \1687_b1 );
or ( \1689_b1 , \c[10]_b1 , \c[9]_b1 );
xor ( \1689_b0 , \c[10]_b0 , w_5184 );
not ( w_5184 , w_5185 );
and ( w_5185 , \c[9]_b1 , \c[9]_b0 );
or ( \1690_b1 , \b[1]_b1 , \c[11]_b1 );
xor ( \1690_b0 , \b[1]_b0 , w_5186 );
not ( w_5186 , w_5187 );
and ( w_5187 , \c[11]_b1 , \c[11]_b0 );
or ( \1691_b1 , \1689_b1 , w_5189 );
not ( w_5189 , w_5190 );
and ( \1691_b0 , \1689_b0 , w_5191 );
and ( w_5190 ,  , w_5191 );
buf ( w_5189 , \1690_b1 );
not ( w_5189 , w_5192 );
not (  , w_5193 );
and ( w_5192 , w_5193 , \1690_b0 );
or ( \1692_b1 , \1688_b1 , w_5195 );
not ( w_5195 , w_5196 );
and ( \1692_b0 , \1688_b0 , w_5197 );
and ( w_5196 ,  , w_5197 );
buf ( w_5195 , \1691_b1 );
not ( w_5195 , w_5198 );
not (  , w_5199 );
and ( w_5198 , w_5199 , \1691_b0 );
buf ( \1693_b1 , \1692_b1 );
not ( \1693_b1 , w_5200 );
not ( \1693_b0 , w_5201 );
and ( w_5200 , w_5201 , \1692_b0 );
or ( \1694_b1 , \1681_b1 , \1693_b1 );
xor ( \1694_b0 , \1681_b0 , w_5202 );
not ( w_5202 , w_5203 );
and ( w_5203 , \1693_b1 , \1693_b0 );
or ( \1695_b1 , \b[0]_b1 , w_5204 );
or ( \1695_b0 , \b[0]_b0 , \c[10]_b0 );
not ( \c[10]_b0 , w_5205 );
and ( w_5205 , w_5204 , \c[10]_b1 );
or ( \1696_b1 , \1695_b1 , w_5207 );
not ( w_5207 , w_5208 );
and ( \1696_b0 , \1695_b0 , w_5209 );
and ( w_5208 ,  , w_5209 );
buf ( w_5207 , \c[9]_b1 );
not ( w_5207 , w_5210 );
not (  , w_5211 );
and ( w_5210 , w_5211 , \c[9]_b0 );
or ( \1697_b1 , \b[0]_b1 , w_5213 );
not ( w_5213 , w_5214 );
and ( \1697_b0 , \b[0]_b0 , w_5215 );
and ( w_5214 ,  , w_5215 );
buf ( w_5213 , \c[10]_b1 );
not ( w_5213 , w_5216 );
not (  , w_5217 );
and ( w_5216 , w_5217 , \c[10]_b0 );
or ( \1699_b1 , \b[8]_b1 , \c[3]_b1 );
xor ( \1699_b0 , \b[8]_b0 , w_5218 );
not ( w_5218 , w_5219 );
and ( w_5219 , \c[3]_b1 , \c[3]_b0 );
buf ( \1700_b1 , \1699_b1 );
not ( \1700_b1 , w_5220 );
not ( \1700_b0 , w_5221 );
and ( w_5220 , w_5221 , \1699_b0 );
or ( \1701_b1 , \c[3]_b1 , \c[2]_b1 );
xor ( \1701_b0 , \c[3]_b0 , w_5222 );
not ( w_5222 , w_5223 );
and ( w_5223 , \c[2]_b1 , \c[2]_b0 );
buf ( \1702_b1 , \1701_b1 );
buf ( \1702_b0 , \1701_b0 );
or ( \1703_b1 , \c[2]_b1 , \c[1]_b1 );
xor ( \1703_b0 , \c[2]_b0 , w_5224 );
not ( w_5224 , w_5225 );
and ( w_5225 , \c[1]_b1 , \c[1]_b0 );
buf ( \1704_b1 , \1703_b1 );
not ( \1704_b1 , w_5226 );
not ( \1704_b0 , w_5227 );
and ( w_5226 , w_5227 , \1703_b0 );
or ( \1705_b1 , \1702_b1 , \1704_b1 );
not ( \1704_b1 , w_5228 );
and ( \1705_b0 , \1702_b0 , w_5229 );
and ( w_5228 , w_5229 , \1704_b0 );
buf ( \1706_b1 , \1705_b1 );
not ( \1706_b1 , w_5230 );
not ( \1706_b0 , w_5231 );
and ( w_5230 , w_5231 , \1705_b0 );
or ( \1707_b1 , \1700_b1 , w_5232 );
or ( \1707_b0 , \1700_b0 , \1706_b0 );
not ( \1706_b0 , w_5233 );
and ( w_5233 , w_5232 , \1706_b1 );
buf ( \1708_b1 , \1703_b1 );
buf ( \1708_b0 , \1703_b0 );
or ( \1709_b1 , \b[9]_b1 , \c[3]_b1 );
xor ( \1709_b0 , \b[9]_b0 , w_5234 );
not ( w_5234 , w_5235 );
and ( w_5235 , \c[3]_b1 , \c[3]_b0 );
or ( \1710_b1 , \1708_b1 , w_5237 );
not ( w_5237 , w_5238 );
and ( \1710_b0 , \1708_b0 , w_5239 );
and ( w_5238 ,  , w_5239 );
buf ( w_5237 , \1709_b1 );
not ( w_5237 , w_5240 );
not (  , w_5241 );
and ( w_5240 , w_5241 , \1709_b0 );
or ( \1711_b1 , \1707_b1 , w_5243 );
not ( w_5243 , w_5244 );
and ( \1711_b0 , \1707_b0 , w_5245 );
and ( w_5244 ,  , w_5245 );
buf ( w_5243 , \1710_b1 );
not ( w_5243 , w_5246 );
not (  , w_5247 );
and ( w_5246 , w_5247 , \1710_b0 );
or ( \1712_b1 , \1698_b1 , \1711_b1 );
xor ( \1712_b0 , \1698_b0 , w_5248 );
not ( w_5248 , w_5249 );
and ( w_5249 , \1711_b1 , \1711_b0 );
or ( \1713_b1 , \1694_b1 , w_5250 );
xor ( \1713_b0 , \1694_b0 , w_5252 );
not ( w_5252 , w_5253 );
and ( w_5253 , w_5250 , w_5251 );
buf ( w_5250 , \1712_b1 );
not ( w_5250 , w_5254 );
not ( w_5251 , w_5255 );
and ( w_5254 , w_5255 , \1712_b0 );
or ( \1714_b1 , \b[0]_b1 , w_5256 );
or ( \1714_b0 , \b[0]_b0 , \c[8]_b0 );
not ( \c[8]_b0 , w_5257 );
and ( w_5257 , w_5256 , \c[8]_b1 );
or ( \1715_b1 , \1714_b1 , w_5259 );
not ( w_5259 , w_5260 );
and ( \1715_b0 , \1714_b0 , w_5261 );
and ( w_5260 ,  , w_5261 );
buf ( w_5259 , \c[7]_b1 );
not ( w_5259 , w_5262 );
not (  , w_5263 );
and ( w_5262 , w_5263 , \c[7]_b0 );
or ( \1716_b1 , \b[0]_b1 , w_5265 );
not ( w_5265 , w_5266 );
and ( \1716_b0 , \b[0]_b0 , w_5267 );
and ( w_5266 ,  , w_5267 );
buf ( w_5265 , \c[8]_b1 );
not ( w_5265 , w_5268 );
not (  , w_5269 );
and ( w_5268 , w_5269 , \c[8]_b0 );
buf ( \1718_b1 , \1717_b1 );
not ( \1718_b1 , w_5270 );
not ( \1718_b0 , w_5271 );
and ( w_5270 , w_5271 , \1717_b0 );
or ( \1719_b1 , \b[6]_b1 , \c[3]_b1 );
xor ( \1719_b0 , \b[6]_b0 , w_5272 );
not ( w_5272 , w_5273 );
and ( w_5273 , \c[3]_b1 , \c[3]_b0 );
buf ( \1720_b1 , \1719_b1 );
not ( \1720_b1 , w_5274 );
not ( \1720_b0 , w_5275 );
and ( w_5274 , w_5275 , \1719_b0 );
buf ( \1721_b1 , \1701_b1 );
not ( \1721_b1 , w_5276 );
not ( \1721_b0 , w_5277 );
and ( w_5276 , w_5277 , \1701_b0 );
or ( \1722_b1 , \1721_b1 , w_5279 );
not ( w_5279 , w_5280 );
and ( \1722_b0 , \1721_b0 , w_5281 );
and ( w_5280 ,  , w_5281 );
buf ( w_5279 , \1703_b1 );
not ( w_5279 , w_5282 );
not (  , w_5283 );
and ( w_5282 , w_5283 , \1703_b0 );
buf ( \1723_b1 , \1722_b1 );
not ( \1723_b1 , w_5284 );
not ( \1723_b0 , w_5285 );
and ( w_5284 , w_5285 , \1722_b0 );
or ( \1724_b1 , \1720_b1 , w_5286 );
or ( \1724_b0 , \1720_b0 , \1723_b0 );
not ( \1723_b0 , w_5287 );
and ( w_5287 , w_5286 , \1723_b1 );
buf ( \1725_b1 , \1704_b1 );
not ( \1725_b1 , w_5288 );
not ( \1725_b0 , w_5289 );
and ( w_5288 , w_5289 , \1704_b0 );
or ( \1726_b1 , \b[7]_b1 , \c[3]_b1 );
xor ( \1726_b0 , \b[7]_b0 , w_5290 );
not ( w_5290 , w_5291 );
and ( w_5291 , \c[3]_b1 , \c[3]_b0 );
or ( \1727_b1 , \1725_b1 , w_5293 );
not ( w_5293 , w_5294 );
and ( \1727_b0 , \1725_b0 , w_5295 );
and ( w_5294 ,  , w_5295 );
buf ( w_5293 , \1726_b1 );
not ( w_5293 , w_5296 );
not (  , w_5297 );
and ( w_5296 , w_5297 , \1726_b0 );
or ( \1728_b1 , \1724_b1 , w_5299 );
not ( w_5299 , w_5300 );
and ( \1728_b0 , \1724_b0 , w_5301 );
and ( w_5300 ,  , w_5301 );
buf ( w_5299 , \1727_b1 );
not ( w_5299 , w_5302 );
not (  , w_5303 );
and ( w_5302 , w_5303 , \1727_b0 );
or ( \1729_b1 , \1718_b1 , w_5305 );
not ( w_5305 , w_5306 );
and ( \1729_b0 , \1718_b0 , w_5307 );
and ( w_5306 ,  , w_5307 );
buf ( w_5305 , \1728_b1 );
not ( w_5305 , w_5308 );
not (  , w_5309 );
and ( w_5308 , w_5309 , \1728_b0 );
buf ( \1730_b1 , \1729_b1 );
not ( \1730_b1 , w_5310 );
not ( \1730_b0 , w_5311 );
and ( w_5310 , w_5311 , \1729_b0 );
or ( \1731_b1 , \1685_b1 , w_5313 );
not ( w_5313 , w_5314 );
and ( \1731_b0 , \1685_b0 , w_5315 );
and ( w_5314 ,  , w_5315 );
buf ( w_5313 , \b[0]_b1 );
not ( w_5313 , w_5316 );
not (  , w_5317 );
and ( w_5316 , w_5317 , \b[0]_b0 );
buf ( \1732_b1 , \1731_b1 );
not ( \1732_b1 , w_5318 );
not ( \1732_b0 , w_5319 );
and ( w_5318 , w_5319 , \1731_b0 );
or ( \1733_b1 , \1703_b1 , \1699_b1 );
not ( \1699_b1 , w_5320 );
and ( \1733_b0 , \1703_b0 , w_5321 );
and ( w_5320 , w_5321 , \1699_b0 );
buf ( \1734_b1 , \1703_b1 );
not ( \1734_b1 , w_5322 );
not ( \1734_b0 , w_5323 );
and ( w_5322 , w_5323 , \1703_b0 );
or ( \1735_b1 , \1701_b1 , \1726_b1 );
not ( \1726_b1 , w_5324 );
and ( \1735_b0 , \1701_b0 , w_5325 );
and ( w_5324 , w_5325 , \1726_b0 );
or ( \1736_b1 , \1734_b1 , \1735_b1 );
not ( \1735_b1 , w_5326 );
and ( \1736_b0 , \1734_b0 , w_5327 );
and ( w_5326 , w_5327 , \1735_b0 );
or ( \1737_b1 , \1733_b1 , w_5328 );
or ( \1737_b0 , \1733_b0 , \1736_b0 );
not ( \1736_b0 , w_5329 );
and ( w_5329 , w_5328 , \1736_b1 );
or ( \1738_b1 , \1732_b1 , \1737_b1 );
xor ( \1738_b0 , \1732_b0 , w_5330 );
not ( w_5330 , w_5331 );
and ( w_5331 , \1737_b1 , \1737_b0 );
or ( \1739_b1 , \c[7]_b1 , \b[3]_b1 );
xor ( \1739_b0 , \c[7]_b0 , w_5332 );
not ( w_5332 , w_5333 );
and ( w_5333 , \b[3]_b1 , \b[3]_b0 );
buf ( \1740_b1 , \1739_b1 );
not ( \1740_b1 , w_5334 );
not ( \1740_b0 , w_5335 );
and ( w_5334 , w_5335 , \1739_b0 );
or ( \1741_b1 , \c[7]_b1 , w_5336 );
xor ( \1741_b0 , \c[7]_b0 , w_5338 );
not ( w_5338 , w_5339 );
and ( w_5339 , w_5336 , w_5337 );
buf ( w_5336 , \c[6]_b1 );
not ( w_5336 , w_5340 );
not ( w_5337 , w_5341 );
and ( w_5340 , w_5341 , \c[6]_b0 );
or ( \1742_b1 , \c[6]_b1 , \c[5]_b1 );
xor ( \1742_b0 , \c[6]_b0 , w_5342 );
not ( w_5342 , w_5343 );
and ( w_5343 , \c[5]_b1 , \c[5]_b0 );
or ( \1743_b1 , \1741_b1 , w_5345 );
not ( w_5345 , w_5346 );
and ( \1743_b0 , \1741_b0 , w_5347 );
and ( w_5346 ,  , w_5347 );
buf ( w_5345 , \1742_b1 );
not ( w_5345 , w_5348 );
not (  , w_5349 );
and ( w_5348 , w_5349 , \1742_b0 );
buf ( \1744_b1 , \1743_b1 );
not ( \1744_b1 , w_5350 );
not ( \1744_b0 , w_5351 );
and ( w_5350 , w_5351 , \1743_b0 );
or ( \1745_b1 , \1740_b1 , w_5352 );
or ( \1745_b0 , \1740_b0 , \1744_b0 );
not ( \1744_b0 , w_5353 );
and ( w_5353 , w_5352 , \1744_b1 );
buf ( \1746_b1 , \1742_b1 );
not ( \1746_b1 , w_5354 );
not ( \1746_b0 , w_5355 );
and ( w_5354 , w_5355 , \1742_b0 );
buf ( \1747_b1 , \1746_b1 );
not ( \1747_b1 , w_5356 );
not ( \1747_b0 , w_5357 );
and ( w_5356 , w_5357 , \1746_b0 );
or ( \1748_b1 , \c[7]_b1 , \b[4]_b1 );
xor ( \1748_b0 , \c[7]_b0 , w_5358 );
not ( w_5358 , w_5359 );
and ( w_5359 , \b[4]_b1 , \b[4]_b0 );
or ( \1749_b1 , \1747_b1 , w_5361 );
not ( w_5361 , w_5362 );
and ( \1749_b0 , \1747_b0 , w_5363 );
and ( w_5362 ,  , w_5363 );
buf ( w_5361 , \1748_b1 );
not ( w_5361 , w_5364 );
not (  , w_5365 );
and ( w_5364 , w_5365 , \1748_b0 );
or ( \1750_b1 , \1745_b1 , w_5367 );
not ( w_5367 , w_5368 );
and ( \1750_b0 , \1745_b0 , w_5369 );
and ( w_5368 ,  , w_5369 );
buf ( w_5367 , \1749_b1 );
not ( w_5367 , w_5370 );
not (  , w_5371 );
and ( w_5370 , w_5371 , \1749_b0 );
or ( \1751_b1 , \1738_b1 , w_5372 );
xor ( \1751_b0 , \1738_b0 , w_5374 );
not ( w_5374 , w_5375 );
and ( w_5375 , w_5372 , w_5373 );
buf ( w_5372 , \1750_b1 );
not ( w_5372 , w_5376 );
not ( w_5373 , w_5377 );
and ( w_5376 , w_5377 , \1750_b0 );
buf ( \1752_b1 , \1751_b1 );
not ( \1752_b1 , w_5378 );
not ( \1752_b0 , w_5379 );
and ( w_5378 , w_5379 , \1751_b0 );
or ( \1753_b1 , \1730_b1 , w_5380 );
or ( \1753_b0 , \1730_b0 , \1752_b0 );
not ( \1752_b0 , w_5381 );
and ( w_5381 , w_5380 , \1752_b1 );
buf ( \1754_b1 , \c[0]_b1 );
not ( \1754_b1 , w_5382 );
not ( \1754_b0 , w_5383 );
and ( w_5382 , w_5383 , \c[0]_b0 );
or ( \1755_b1 , \1754_b1 , w_5385 );
not ( w_5385 , w_5386 );
and ( \1755_b0 , \1754_b0 , w_5387 );
and ( w_5386 ,  , w_5387 );
buf ( w_5385 , \c[1]_b1 );
not ( w_5385 , w_5388 );
not (  , w_5389 );
and ( w_5388 , w_5389 , \c[1]_b0 );
buf ( \1756_b1 , \1755_b1 );
not ( \1756_b1 , w_5390 );
not ( \1756_b0 , w_5391 );
and ( w_5390 , w_5391 , \1755_b0 );
or ( \1757_b1 , \c[1]_b1 , \b[8]_b1 );
xor ( \1757_b0 , \c[1]_b0 , w_5392 );
not ( w_5392 , w_5393 );
and ( w_5393 , \b[8]_b1 , \b[8]_b0 );
or ( \1758_b1 , \1756_b1 , \1757_b1 );
not ( \1757_b1 , w_5394 );
and ( \1758_b0 , \1756_b0 , w_5395 );
and ( w_5394 , w_5395 , \1757_b0 );
or ( \1759_b1 , \c[1]_b1 , \b[9]_b1 );
xor ( \1759_b0 , \c[1]_b0 , w_5396 );
not ( w_5396 , w_5397 );
and ( w_5397 , \b[9]_b1 , \b[9]_b0 );
or ( \1760_b1 , \1759_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_5398 );
and ( \1760_b0 , \1759_b0 , w_5399 );
and ( w_5398 , w_5399 , \c[0]_b0 );
or ( \1761_b1 , \1758_b1 , w_5401 );
not ( w_5401 , w_5402 );
and ( \1761_b0 , \1758_b0 , w_5403 );
and ( w_5402 ,  , w_5403 );
buf ( w_5401 , \1760_b1 );
not ( w_5401 , w_5404 );
not (  , w_5405 );
and ( w_5404 , w_5405 , \1760_b0 );
buf ( \1762_b1 , \1761_b1 );
not ( \1762_b1 , w_5406 );
not ( \1762_b0 , w_5407 );
and ( w_5406 , w_5407 , \1761_b0 );
buf ( \1763_b1 , \1762_b1 );
not ( \1763_b1 , w_5408 );
not ( \1763_b0 , w_5409 );
and ( w_5408 , w_5409 , \1762_b0 );
or ( \1764_b1 , \c[9]_b1 , \b[0]_b1 );
xor ( \1764_b0 , \c[9]_b0 , w_5410 );
not ( w_5410 , w_5411 );
and ( w_5411 , \b[0]_b1 , \b[0]_b0 );
buf ( \1765_b1 , \1764_b1 );
not ( \1765_b1 , w_5412 );
not ( \1765_b0 , w_5413 );
and ( w_5412 , w_5413 , \1764_b0 );
buf ( \1766_b1 , \c[7]_b1 );
not ( \1766_b1 , w_5414 );
not ( \1766_b0 , w_5415 );
and ( w_5414 , w_5415 , \c[7]_b0 );
or ( \1767_b1 , \1766_b1 , w_5417 );
not ( w_5417 , w_5418 );
and ( \1767_b0 , \1766_b0 , w_5419 );
and ( w_5418 ,  , w_5419 );
buf ( w_5417 , \c[8]_b1 );
not ( w_5417 , w_5420 );
not (  , w_5421 );
and ( w_5420 , w_5421 , \c[8]_b0 );
or ( \1768_b1 , \c[9]_b1 , w_5422 );
or ( \1768_b0 , \c[9]_b0 , \c[8]_b0 );
not ( \c[8]_b0 , w_5423 );
and ( w_5423 , w_5422 , \c[8]_b1 );
or ( \1769_b1 , \c[9]_b1 , w_5425 );
not ( w_5425 , w_5426 );
and ( \1769_b0 , \c[9]_b0 , w_5427 );
and ( w_5426 ,  , w_5427 );
buf ( w_5425 , \c[7]_b1 );
not ( w_5425 , w_5428 );
not (  , w_5429 );
and ( w_5428 , w_5429 , \c[7]_b0 );
buf ( \1771_b1 , \1770_b1 );
not ( \1771_b1 , w_5430 );
not ( \1771_b0 , w_5431 );
and ( w_5430 , w_5431 , \1770_b0 );
or ( \1772_b1 , \1765_b1 , w_5432 );
or ( \1772_b0 , \1765_b0 , \1771_b0 );
not ( \1771_b0 , w_5433 );
and ( w_5433 , w_5432 , \1771_b1 );
or ( \1773_b1 , \c[8]_b1 , \c[7]_b1 );
xor ( \1773_b0 , \c[8]_b0 , w_5434 );
not ( w_5434 , w_5435 );
and ( w_5435 , \c[7]_b1 , \c[7]_b0 );
or ( \1774_b1 , \c[9]_b1 , \b[1]_b1 );
xor ( \1774_b0 , \c[9]_b0 , w_5436 );
not ( w_5436 , w_5437 );
and ( w_5437 , \b[1]_b1 , \b[1]_b0 );
or ( \1775_b1 , \1773_b1 , w_5439 );
not ( w_5439 , w_5440 );
and ( \1775_b0 , \1773_b0 , w_5441 );
and ( w_5440 ,  , w_5441 );
buf ( w_5439 , \1774_b1 );
not ( w_5439 , w_5442 );
not (  , w_5443 );
and ( w_5442 , w_5443 , \1774_b0 );
or ( \1776_b1 , \1772_b1 , w_5445 );
not ( w_5445 , w_5446 );
and ( \1776_b0 , \1772_b0 , w_5447 );
and ( w_5446 ,  , w_5447 );
buf ( w_5445 , \1775_b1 );
not ( w_5445 , w_5448 );
not (  , w_5449 );
and ( w_5448 , w_5449 , \1775_b0 );
buf ( \1777_b1 , \1776_b1 );
not ( \1777_b1 , w_5450 );
not ( \1777_b0 , w_5451 );
and ( w_5450 , w_5451 , \1776_b0 );
or ( \1778_b1 , \1763_b1 , w_5452 );
or ( \1778_b0 , \1763_b0 , \1777_b0 );
not ( \1777_b0 , w_5453 );
and ( w_5453 , w_5452 , \1777_b1 );
or ( \1779_b1 , \1776_b1 , w_5454 );
or ( \1779_b0 , \1776_b0 , \1762_b0 );
not ( \1762_b0 , w_5455 );
and ( w_5455 , w_5454 , \1762_b1 );
or ( \1780_b1 , \c[7]_b1 , \b[2]_b1 );
xor ( \1780_b0 , \c[7]_b0 , w_5456 );
not ( w_5456 , w_5457 );
and ( w_5457 , \b[2]_b1 , \b[2]_b0 );
buf ( \1781_b1 , \1780_b1 );
not ( \1781_b1 , w_5458 );
not ( \1781_b0 , w_5459 );
and ( w_5458 , w_5459 , \1780_b0 );
or ( \1782_b1 , \1741_b1 , w_5461 );
not ( w_5461 , w_5462 );
and ( \1782_b0 , \1741_b0 , w_5463 );
and ( w_5462 ,  , w_5463 );
buf ( w_5461 , \1742_b1 );
not ( w_5461 , w_5464 );
not (  , w_5465 );
and ( w_5464 , w_5465 , \1742_b0 );
buf ( \1783_b1 , \1782_b1 );
not ( \1783_b1 , w_5466 );
not ( \1783_b0 , w_5467 );
and ( w_5466 , w_5467 , \1782_b0 );
or ( \1784_b1 , \1781_b1 , w_5468 );
or ( \1784_b0 , \1781_b0 , \1783_b0 );
not ( \1783_b0 , w_5469 );
and ( w_5469 , w_5468 , \1783_b1 );
buf ( \1785_b1 , \1746_b1 );
not ( \1785_b1 , w_5470 );
not ( \1785_b0 , w_5471 );
and ( w_5470 , w_5471 , \1746_b0 );
or ( \1786_b1 , \1785_b1 , w_5473 );
not ( w_5473 , w_5474 );
and ( \1786_b0 , \1785_b0 , w_5475 );
and ( w_5474 ,  , w_5475 );
buf ( w_5473 , \1739_b1 );
not ( w_5473 , w_5476 );
not (  , w_5477 );
and ( w_5476 , w_5477 , \1739_b0 );
or ( \1787_b1 , \1784_b1 , w_5479 );
not ( w_5479 , w_5480 );
and ( \1787_b0 , \1784_b0 , w_5481 );
and ( w_5480 ,  , w_5481 );
buf ( w_5479 , \1786_b1 );
not ( w_5479 , w_5482 );
not (  , w_5483 );
and ( w_5482 , w_5483 , \1786_b0 );
or ( \1788_b1 , \1779_b1 , w_5485 );
not ( w_5485 , w_5486 );
and ( \1788_b0 , \1779_b0 , w_5487 );
and ( w_5486 ,  , w_5487 );
buf ( w_5485 , \1787_b1 );
not ( w_5485 , w_5488 );
not (  , w_5489 );
and ( w_5488 , w_5489 , \1787_b0 );
or ( \1789_b1 , \1778_b1 , w_5491 );
not ( w_5491 , w_5492 );
and ( \1789_b0 , \1778_b0 , w_5493 );
and ( w_5492 ,  , w_5493 );
buf ( w_5491 , \1788_b1 );
not ( w_5491 , w_5494 );
not (  , w_5495 );
and ( w_5494 , w_5495 , \1788_b0 );
or ( \1790_b1 , \1753_b1 , w_5497 );
not ( w_5497 , w_5498 );
and ( \1790_b0 , \1753_b0 , w_5499 );
and ( w_5498 ,  , w_5499 );
buf ( w_5497 , \1789_b1 );
not ( w_5497 , w_5500 );
not (  , w_5501 );
and ( w_5500 , w_5501 , \1789_b0 );
buf ( \1791_b1 , \1729_b1 );
not ( \1791_b1 , w_5502 );
not ( \1791_b0 , w_5503 );
and ( w_5502 , w_5503 , \1729_b0 );
buf ( \1792_b1 , \1751_b1 );
not ( \1792_b1 , w_5504 );
not ( \1792_b0 , w_5505 );
and ( w_5504 , w_5505 , \1751_b0 );
or ( \1793_b1 , \1791_b1 , w_5507 );
not ( w_5507 , w_5508 );
and ( \1793_b0 , \1791_b0 , w_5509 );
and ( w_5508 ,  , w_5509 );
buf ( w_5507 , \1792_b1 );
not ( w_5507 , w_5510 );
not (  , w_5511 );
and ( w_5510 , w_5511 , \1792_b0 );
or ( \1794_b1 , \1790_b1 , w_5513 );
not ( w_5513 , w_5514 );
and ( \1794_b0 , \1790_b0 , w_5515 );
and ( w_5514 ,  , w_5515 );
buf ( w_5513 , \1793_b1 );
not ( w_5513 , w_5516 );
not (  , w_5517 );
and ( w_5516 , w_5517 , \1793_b0 );
or ( \1795_b1 , \1713_b1 , \1794_b1 );
xor ( \1795_b0 , \1713_b0 , w_5518 );
not ( w_5518 , w_5519 );
and ( w_5519 , \1794_b1 , \1794_b0 );
or ( \1796_b1 , \b[2]_b1 , \c[9]_b1 );
xor ( \1796_b0 , \b[2]_b0 , w_5520 );
not ( w_5520 , w_5521 );
and ( w_5521 , \c[9]_b1 , \c[9]_b0 );
buf ( \1797_b1 , \1796_b1 );
not ( \1797_b1 , w_5522 );
not ( \1797_b0 , w_5523 );
and ( w_5522 , w_5523 , \1796_b0 );
buf ( \1798_b1 , \c[7]_b1 );
not ( \1798_b1 , w_5524 );
not ( \1798_b0 , w_5525 );
and ( w_5524 , w_5525 , \c[7]_b0 );
buf ( \1799_b1 , \c[8]_b1 );
not ( \1799_b1 , w_5526 );
not ( \1799_b0 , w_5527 );
and ( w_5526 , w_5527 , \c[8]_b0 );
buf ( \1800_b1 , \1799_b1 );
not ( \1800_b1 , w_5528 );
not ( \1800_b0 , w_5529 );
and ( w_5528 , w_5529 , \1799_b0 );
or ( \1801_b1 , \1798_b1 , w_5530 );
or ( \1801_b0 , \1798_b0 , \1800_b0 );
not ( \1800_b0 , w_5531 );
and ( w_5531 , w_5530 , \1800_b1 );
or ( \1802_b1 , \1801_b1 , w_5533 );
not ( w_5533 , w_5534 );
and ( \1802_b0 , \1801_b0 , w_5535 );
and ( w_5534 ,  , w_5535 );
buf ( w_5533 , \1767_b1 );
not ( w_5533 , w_5536 );
not (  , w_5537 );
and ( w_5536 , w_5537 , \1767_b0 );
buf ( \1803_b1 , \1802_b1 );
not ( \1803_b1 , w_5538 );
not ( \1803_b0 , w_5539 );
and ( w_5538 , w_5539 , \1802_b0 );
or ( \1804_b1 , \1797_b1 , w_5540 );
or ( \1804_b0 , \1797_b0 , \1803_b0 );
not ( \1803_b0 , w_5541 );
and ( w_5541 , w_5540 , \1803_b1 );
or ( \1805_b1 , \1770_b1 , w_5543 );
not ( w_5543 , w_5544 );
and ( \1805_b0 , \1770_b0 , w_5545 );
and ( w_5544 ,  , w_5545 );
buf ( w_5543 , \1774_b1 );
not ( w_5543 , w_5546 );
not (  , w_5547 );
and ( w_5546 , w_5547 , \1774_b0 );
or ( \1806_b1 , \1804_b1 , w_5549 );
not ( w_5549 , w_5550 );
and ( \1806_b0 , \1804_b0 , w_5551 );
and ( w_5550 ,  , w_5551 );
buf ( w_5549 , \1805_b1 );
not ( w_5549 , w_5552 );
not (  , w_5553 );
and ( w_5552 , w_5553 , \1805_b0 );
buf ( \1807_b1 , \1759_b1 );
not ( \1807_b1 , w_5554 );
not ( \1807_b0 , w_5555 );
and ( w_5554 , w_5555 , \1759_b0 );
buf ( \1808_b1 , \1756_b1 );
not ( \1808_b1 , w_5556 );
not ( \1808_b0 , w_5557 );
and ( w_5556 , w_5557 , \1756_b0 );
or ( \1809_b1 , \1807_b1 , w_5558 );
or ( \1809_b0 , \1807_b0 , \1808_b0 );
not ( \1808_b0 , w_5559 );
and ( w_5559 , w_5558 , \1808_b1 );
or ( \1810_b1 , \b[10]_b1 , \c[1]_b1 );
xor ( \1810_b0 , \b[10]_b0 , w_5560 );
not ( w_5560 , w_5561 );
and ( w_5561 , \c[1]_b1 , \c[1]_b0 );
or ( \1811_b1 , \1810_b1 , w_5563 );
not ( w_5563 , w_5564 );
and ( \1811_b0 , \1810_b0 , w_5565 );
and ( w_5564 ,  , w_5565 );
buf ( w_5563 , \c[0]_b1 );
not ( w_5563 , w_5566 );
not (  , w_5567 );
and ( w_5566 , w_5567 , \c[0]_b0 );
or ( \1812_b1 , \1809_b1 , w_5569 );
not ( w_5569 , w_5570 );
and ( \1812_b0 , \1809_b0 , w_5571 );
and ( w_5570 ,  , w_5571 );
buf ( w_5569 , \1811_b1 );
not ( w_5569 , w_5572 );
not (  , w_5573 );
and ( w_5572 , w_5573 , \1811_b0 );
or ( \1813_b1 , \1806_b1 , w_5574 );
or ( \1813_b0 , \1806_b0 , \1812_b0 );
not ( \1812_b0 , w_5575 );
and ( w_5575 , w_5574 , \1812_b1 );
or ( \1814_b1 , \b[5]_b1 , \c[5]_b1 );
xor ( \1814_b0 , \b[5]_b0 , w_5576 );
not ( w_5576 , w_5577 );
and ( w_5577 , \c[5]_b1 , \c[5]_b0 );
buf ( \1815_b1 , \1814_b1 );
not ( \1815_b1 , w_5578 );
not ( \1815_b0 , w_5579 );
and ( w_5578 , w_5579 , \1814_b0 );
buf ( \1816_b1 , \1675_b1 );
not ( \1816_b1 , w_5580 );
not ( \1816_b0 , w_5581 );
and ( w_5580 , w_5581 , \1675_b0 );
or ( \1817_b1 , \1815_b1 , w_5582 );
or ( \1817_b0 , \1815_b0 , \1816_b0 );
not ( \1816_b0 , w_5583 );
and ( w_5583 , w_5582 , \1816_b1 );
or ( \1818_b1 , \1678_b1 , w_5585 );
not ( w_5585 , w_5586 );
and ( \1818_b0 , \1678_b0 , w_5587 );
and ( w_5586 ,  , w_5587 );
buf ( w_5585 , \1670_b1 );
not ( w_5585 , w_5588 );
not (  , w_5589 );
and ( w_5588 , w_5589 , \1670_b0 );
or ( \1819_b1 , \1817_b1 , w_5591 );
not ( w_5591 , w_5592 );
and ( \1819_b0 , \1817_b0 , w_5593 );
and ( w_5592 ,  , w_5593 );
buf ( w_5591 , \1818_b1 );
not ( w_5591 , w_5594 );
not (  , w_5595 );
and ( w_5594 , w_5595 , \1818_b0 );
or ( \1820_b1 , \1813_b1 , w_5597 );
not ( w_5597 , w_5598 );
and ( \1820_b0 , \1813_b0 , w_5599 );
and ( w_5598 ,  , w_5599 );
buf ( w_5597 , \1819_b1 );
not ( w_5597 , w_5600 );
not (  , w_5601 );
and ( w_5600 , w_5601 , \1819_b0 );
or ( \1821_b1 , \1806_b1 , w_5603 );
not ( w_5603 , w_5604 );
and ( \1821_b0 , \1806_b0 , w_5605 );
and ( w_5604 ,  , w_5605 );
buf ( w_5603 , \1812_b1 );
not ( w_5603 , w_5606 );
not (  , w_5607 );
and ( w_5606 , w_5607 , \1812_b0 );
or ( \1822_b1 , \1820_b1 , w_5609 );
not ( w_5609 , w_5610 );
and ( \1822_b0 , \1820_b0 , w_5611 );
and ( w_5610 ,  , w_5611 );
buf ( w_5609 , \1821_b1 );
not ( w_5609 , w_5612 );
not (  , w_5613 );
and ( w_5612 , w_5613 , \1821_b0 );
buf ( \1823_b1 , \1737_b1 );
not ( \1823_b1 , w_5614 );
not ( \1823_b0 , w_5615 );
and ( w_5614 , w_5615 , \1737_b0 );
or ( \1824_b1 , \1823_b1 , w_5617 );
not ( w_5617 , w_5618 );
and ( \1824_b0 , \1823_b0 , w_5619 );
and ( w_5618 ,  , w_5619 );
buf ( w_5617 , \1731_b1 );
not ( w_5617 , w_5620 );
not (  , w_5621 );
and ( w_5620 , w_5621 , \1731_b0 );
buf ( \1825_b1 , \1824_b1 );
not ( \1825_b1 , w_5622 );
not ( \1825_b0 , w_5623 );
and ( w_5622 , w_5623 , \1824_b0 );
buf ( \1826_b1 , \1750_b1 );
not ( \1826_b1 , w_5624 );
not ( \1826_b0 , w_5625 );
and ( w_5624 , w_5625 , \1750_b0 );
or ( \1827_b1 , \1825_b1 , w_5626 );
or ( \1827_b0 , \1825_b0 , \1826_b0 );
not ( \1826_b0 , w_5627 );
and ( w_5627 , w_5626 , \1826_b1 );
or ( \1828_b1 , \1737_b1 , w_5629 );
not ( w_5629 , w_5630 );
and ( \1828_b0 , \1737_b0 , w_5631 );
and ( w_5630 ,  , w_5631 );
buf ( w_5629 , \1732_b1 );
not ( w_5629 , w_5632 );
not (  , w_5633 );
and ( w_5632 , w_5633 , \1732_b0 );
or ( \1829_b1 , \1827_b1 , w_5635 );
not ( w_5635 , w_5636 );
and ( \1829_b0 , \1827_b0 , w_5637 );
and ( w_5636 ,  , w_5637 );
buf ( w_5635 , \1828_b1 );
not ( w_5635 , w_5638 );
not (  , w_5639 );
and ( w_5638 , w_5639 , \1828_b0 );
or ( \1830_b1 , \1822_b1 , \1829_b1 );
xor ( \1830_b0 , \1822_b0 , w_5640 );
not ( w_5640 , w_5641 );
and ( w_5641 , \1829_b1 , \1829_b0 );
buf ( \1831_b1 , \1748_b1 );
not ( \1831_b1 , w_5642 );
not ( \1831_b0 , w_5643 );
and ( w_5642 , w_5643 , \1748_b0 );
buf ( \1832_b1 , \1782_b1 );
not ( \1832_b1 , w_5644 );
not ( \1832_b0 , w_5645 );
and ( w_5644 , w_5645 , \1782_b0 );
or ( \1833_b1 , \1831_b1 , w_5646 );
or ( \1833_b0 , \1831_b0 , \1832_b0 );
not ( \1832_b0 , w_5647 );
and ( w_5647 , w_5646 , \1832_b1 );
or ( \1834_b1 , \b[5]_b1 , \c[7]_b1 );
xor ( \1834_b0 , \b[5]_b0 , w_5648 );
not ( w_5648 , w_5649 );
and ( w_5649 , \c[7]_b1 , \c[7]_b0 );
or ( \1835_b1 , \1747_b1 , w_5651 );
not ( w_5651 , w_5652 );
and ( \1835_b0 , \1747_b0 , w_5653 );
and ( w_5652 ,  , w_5653 );
buf ( w_5651 , \1834_b1 );
not ( w_5651 , w_5654 );
not (  , w_5655 );
and ( w_5654 , w_5655 , \1834_b0 );
or ( \1836_b1 , \1833_b1 , w_5657 );
not ( w_5657 , w_5658 );
and ( \1836_b0 , \1833_b0 , w_5659 );
and ( w_5658 ,  , w_5659 );
buf ( w_5657 , \1835_b1 );
not ( w_5657 , w_5660 );
not (  , w_5661 );
and ( w_5660 , w_5661 , \1835_b0 );
buf ( \1837_b1 , \1810_b1 );
not ( \1837_b1 , w_5662 );
not ( \1837_b0 , w_5663 );
and ( w_5662 , w_5663 , \1810_b0 );
buf ( \1838_b1 , \1756_b1 );
not ( \1838_b1 , w_5664 );
not ( \1838_b0 , w_5665 );
and ( w_5664 , w_5665 , \1756_b0 );
or ( \1839_b1 , \1837_b1 , w_5666 );
or ( \1839_b0 , \1837_b0 , \1838_b0 );
not ( \1838_b0 , w_5667 );
and ( w_5667 , w_5666 , \1838_b1 );
or ( \1840_b1 , \b[11]_b1 , \c[1]_b1 );
xor ( \1840_b0 , \b[11]_b0 , w_5668 );
not ( w_5668 , w_5669 );
and ( w_5669 , \c[1]_b1 , \c[1]_b0 );
or ( \1841_b1 , \1840_b1 , w_5671 );
not ( w_5671 , w_5672 );
and ( \1841_b0 , \1840_b0 , w_5673 );
and ( w_5672 ,  , w_5673 );
buf ( w_5671 , \c[0]_b1 );
not ( w_5671 , w_5674 );
not (  , w_5675 );
and ( w_5674 , w_5675 , \c[0]_b0 );
or ( \1842_b1 , \1839_b1 , w_5677 );
not ( w_5677 , w_5678 );
and ( \1842_b0 , \1839_b0 , w_5679 );
and ( w_5678 ,  , w_5679 );
buf ( w_5677 , \1841_b1 );
not ( w_5677 , w_5680 );
not (  , w_5681 );
and ( w_5680 , w_5681 , \1841_b0 );
buf ( \1843_b1 , \1842_b1 );
not ( \1843_b1 , w_5682 );
not ( \1843_b0 , w_5683 );
and ( w_5682 , w_5683 , \1842_b0 );
or ( \1844_b1 , \1836_b1 , \1843_b1 );
not ( \1843_b1 , w_5684 );
and ( \1844_b0 , \1836_b0 , w_5685 );
and ( w_5684 , w_5685 , \1843_b0 );
buf ( \1845_b1 , \1836_b1 );
not ( \1845_b1 , w_5686 );
not ( \1845_b0 , w_5687 );
and ( w_5686 , w_5687 , \1836_b0 );
or ( \1846_b1 , \1845_b1 , \1842_b1 );
not ( \1842_b1 , w_5688 );
and ( \1846_b0 , \1845_b0 , w_5689 );
and ( w_5688 , w_5689 , \1842_b0 );
or ( \1847_b1 , \1844_b1 , w_5690 );
or ( \1847_b0 , \1844_b0 , \1846_b0 );
not ( \1846_b0 , w_5691 );
and ( w_5691 , w_5690 , \1846_b1 );
buf ( \1848_b1 , \1767_b1 );
not ( \1848_b1 , w_5692 );
not ( \1848_b0 , w_5693 );
and ( w_5692 , w_5693 , \1767_b0 );
or ( \1849_b1 , \c[9]_b1 , w_5694 );
or ( \1849_b0 , \c[9]_b0 , \c[8]_b0 );
not ( \c[8]_b0 , w_5695 );
and ( w_5695 , w_5694 , \c[8]_b1 );
or ( \1850_b1 , \1849_b1 , w_5697 );
not ( w_5697 , w_5698 );
and ( \1850_b0 , \1849_b0 , w_5699 );
and ( w_5698 ,  , w_5699 );
buf ( w_5697 , \1769_b1 );
not ( w_5697 , w_5700 );
not (  , w_5701 );
and ( w_5700 , w_5701 , \1769_b0 );
or ( \1851_b1 , \1848_b1 , w_5703 );
not ( w_5703 , w_5704 );
and ( \1851_b0 , \1848_b0 , w_5705 );
and ( w_5704 ,  , w_5705 );
buf ( w_5703 , \1850_b1 );
not ( w_5703 , w_5706 );
not (  , w_5707 );
and ( w_5706 , w_5707 , \1850_b0 );
buf ( \1852_b1 , \1851_b1 );
not ( \1852_b1 , w_5708 );
not ( \1852_b0 , w_5709 );
and ( w_5708 , w_5709 , \1851_b0 );
buf ( \1853_b1 , \1852_b1 );
not ( \1853_b1 , w_5710 );
not ( \1853_b0 , w_5711 );
and ( w_5710 , w_5711 , \1852_b0 );
buf ( \1854_b1 , \1796_b1 );
not ( \1854_b1 , w_5712 );
not ( \1854_b0 , w_5713 );
and ( w_5712 , w_5713 , \1796_b0 );
buf ( \1855_b1 , \1854_b1 );
not ( \1855_b1 , w_5714 );
not ( \1855_b0 , w_5715 );
and ( w_5714 , w_5715 , \1854_b0 );
or ( \1856_b1 , \1853_b1 , \1855_b1 );
not ( \1855_b1 , w_5716 );
and ( \1856_b0 , \1853_b0 , w_5717 );
and ( w_5716 , w_5717 , \1855_b0 );
or ( \1857_b1 , \b[3]_b1 , \c[9]_b1 );
xor ( \1857_b0 , \b[3]_b0 , w_5718 );
not ( w_5718 , w_5719 );
and ( w_5719 , \c[9]_b1 , \c[9]_b0 );
or ( \1858_b1 , \1802_b1 , \1857_b1 );
not ( \1857_b1 , w_5720 );
and ( \1858_b0 , \1802_b0 , w_5721 );
and ( w_5720 , w_5721 , \1857_b0 );
or ( \1859_b1 , \1856_b1 , w_5723 );
not ( w_5723 , w_5724 );
and ( \1859_b0 , \1856_b0 , w_5725 );
and ( w_5724 ,  , w_5725 );
buf ( w_5723 , \1858_b1 );
not ( w_5723 , w_5726 );
not (  , w_5727 );
and ( w_5726 , w_5727 , \1858_b0 );
buf ( \1860_b1 , \1859_b1 );
not ( \1860_b1 , w_5728 );
not ( \1860_b0 , w_5729 );
and ( w_5728 , w_5729 , \1859_b0 );
or ( \1861_b1 , \1847_b1 , \1860_b1 );
not ( \1860_b1 , w_5730 );
and ( \1861_b0 , \1847_b0 , w_5731 );
and ( w_5730 , w_5731 , \1860_b0 );
buf ( \1862_b1 , \1847_b1 );
not ( \1862_b1 , w_5732 );
not ( \1862_b0 , w_5733 );
and ( w_5732 , w_5733 , \1847_b0 );
or ( \1863_b1 , \1862_b1 , \1859_b1 );
not ( \1859_b1 , w_5734 );
and ( \1863_b0 , \1862_b0 , w_5735 );
and ( w_5734 , w_5735 , \1859_b0 );
or ( \1864_b1 , \1861_b1 , w_5737 );
not ( w_5737 , w_5738 );
and ( \1864_b0 , \1861_b0 , w_5739 );
and ( w_5738 ,  , w_5739 );
buf ( w_5737 , \1863_b1 );
not ( w_5737 , w_5740 );
not (  , w_5741 );
and ( w_5740 , w_5741 , \1863_b0 );
or ( \1865_b1 , \1830_b1 , w_5742 );
xor ( \1865_b0 , \1830_b0 , w_5744 );
not ( w_5744 , w_5745 );
and ( w_5745 , w_5742 , w_5743 );
buf ( w_5742 , \1864_b1 );
not ( w_5742 , w_5746 );
not ( w_5743 , w_5747 );
and ( w_5746 , w_5747 , \1864_b0 );
or ( \1866_b1 , \1795_b1 , \1865_b1 );
xor ( \1866_b0 , \1795_b0 , w_5748 );
not ( w_5748 , w_5749 );
and ( w_5749 , \1865_b1 , \1865_b0 );
or ( \1867_b1 , \1806_b1 , \1812_b1 );
xor ( \1867_b0 , \1806_b0 , w_5750 );
not ( w_5750 , w_5751 );
and ( w_5751 , \1812_b1 , \1812_b0 );
or ( \1868_b1 , \1867_b1 , w_5752 );
xor ( \1868_b0 , \1867_b0 , w_5754 );
not ( w_5754 , w_5755 );
and ( w_5755 , w_5752 , w_5753 );
buf ( w_5752 , \1819_b1 );
not ( w_5752 , w_5756 );
not ( w_5753 , w_5757 );
and ( w_5756 , w_5757 , \1819_b0 );
or ( \1869_b1 , \b[4]_b1 , \c[5]_b1 );
xor ( \1869_b0 , \b[4]_b0 , w_5758 );
not ( w_5758 , w_5759 );
and ( w_5759 , \c[5]_b1 , \c[5]_b0 );
or ( \1870_b1 , \1675_b1 , \1869_b1 );
not ( \1869_b1 , w_5760 );
and ( \1870_b0 , \1675_b0 , w_5761 );
and ( w_5760 , w_5761 , \1869_b0 );
or ( \1871_b1 , \1678_b1 , \1814_b1 );
not ( \1814_b1 , w_5762 );
and ( \1871_b0 , \1678_b0 , w_5763 );
and ( w_5762 , w_5763 , \1814_b0 );
or ( \1872_b1 , \1870_b1 , w_5765 );
not ( w_5765 , w_5766 );
and ( \1872_b0 , \1870_b0 , w_5767 );
and ( w_5766 ,  , w_5767 );
buf ( w_5765 , \1871_b1 );
not ( w_5765 , w_5768 );
not (  , w_5769 );
and ( w_5768 , w_5769 , \1871_b0 );
buf ( \1873_b1 , \1728_b1 );
not ( \1873_b1 , w_5770 );
not ( \1873_b0 , w_5771 );
and ( w_5770 , w_5771 , \1728_b0 );
buf ( \1874_b1 , \1717_b1 );
not ( \1874_b1 , w_5772 );
not ( \1874_b0 , w_5773 );
and ( w_5772 , w_5773 , \1717_b0 );
or ( \1875_b1 , \1873_b1 , \1874_b1 );
not ( \1874_b1 , w_5774 );
and ( \1875_b0 , \1873_b0 , w_5775 );
and ( w_5774 , w_5775 , \1874_b0 );
or ( \1876_b1 , \1728_b1 , \1717_b1 );
not ( \1717_b1 , w_5776 );
and ( \1876_b0 , \1728_b0 , w_5777 );
and ( w_5776 , w_5777 , \1717_b0 );
or ( \1877_b1 , \1875_b1 , w_5779 );
not ( w_5779 , w_5780 );
and ( \1877_b0 , \1875_b0 , w_5781 );
and ( w_5780 ,  , w_5781 );
buf ( w_5779 , \1876_b1 );
not ( w_5779 , w_5782 );
not (  , w_5783 );
and ( w_5782 , w_5783 , \1876_b0 );
or ( \1878_b1 , \1872_b1 , \1877_b1 );
xor ( \1878_b0 , \1872_b0 , w_5784 );
not ( w_5784 , w_5785 );
and ( w_5785 , \1877_b1 , \1877_b0 );
or ( \1879_b1 , \1773_b1 , w_5787 );
not ( w_5787 , w_5788 );
and ( \1879_b0 , \1773_b0 , w_5789 );
and ( w_5788 ,  , w_5789 );
buf ( w_5787 , \b[0]_b1 );
not ( w_5787 , w_5790 );
not (  , w_5791 );
and ( w_5790 , w_5791 , \b[0]_b0 );
or ( \1880_b1 , \c[1]_b1 , \b[7]_b1 );
xor ( \1880_b0 , \c[1]_b0 , w_5792 );
not ( w_5792 , w_5793 );
and ( w_5793 , \b[7]_b1 , \b[7]_b0 );
or ( \1881_b1 , \1756_b1 , \1880_b1 );
not ( \1880_b1 , w_5794 );
and ( \1881_b0 , \1756_b0 , w_5795 );
and ( w_5794 , w_5795 , \1880_b0 );
or ( \1882_b1 , \1757_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_5796 );
and ( \1882_b0 , \1757_b0 , w_5797 );
and ( w_5796 , w_5797 , \c[0]_b0 );
or ( \1883_b1 , \1881_b1 , w_5799 );
not ( w_5799 , w_5800 );
and ( \1883_b0 , \1881_b0 , w_5801 );
and ( w_5800 ,  , w_5801 );
buf ( w_5799 , \1882_b1 );
not ( w_5799 , w_5802 );
not (  , w_5803 );
and ( w_5802 , w_5803 , \1882_b0 );
or ( \1884_b1 , \1879_b1 , \1883_b1 );
xor ( \1884_b0 , \1879_b0 , w_5804 );
not ( w_5804 , w_5805 );
and ( w_5805 , \1883_b1 , \1883_b0 );
or ( \1885_b1 , \b[1]_b1 , \c[7]_b1 );
xor ( \1885_b0 , \b[1]_b0 , w_5806 );
not ( w_5806 , w_5807 );
and ( w_5807 , \c[7]_b1 , \c[7]_b0 );
or ( \1886_b1 , \1782_b1 , \1885_b1 );
not ( \1885_b1 , w_5808 );
and ( \1886_b0 , \1782_b0 , w_5809 );
and ( w_5808 , w_5809 , \1885_b0 );
or ( \1887_b1 , \1747_b1 , \1780_b1 );
not ( \1780_b1 , w_5810 );
and ( \1887_b0 , \1747_b0 , w_5811 );
and ( w_5810 , w_5811 , \1780_b0 );
or ( \1888_b1 , \1886_b1 , w_5813 );
not ( w_5813 , w_5814 );
and ( \1888_b0 , \1886_b0 , w_5815 );
and ( w_5814 ,  , w_5815 );
buf ( w_5813 , \1887_b1 );
not ( w_5813 , w_5816 );
not (  , w_5817 );
and ( w_5816 , w_5817 , \1887_b0 );
or ( \1889_b1 , \1884_b1 , \1888_b1 );
not ( \1888_b1 , w_5818 );
and ( \1889_b0 , \1884_b0 , w_5819 );
and ( w_5818 , w_5819 , \1888_b0 );
or ( \1890_b1 , \1879_b1 , \1883_b1 );
not ( \1883_b1 , w_5820 );
and ( \1890_b0 , \1879_b0 , w_5821 );
and ( w_5820 , w_5821 , \1883_b0 );
or ( \1891_b1 , \1889_b1 , w_5822 );
or ( \1891_b0 , \1889_b0 , \1890_b0 );
not ( \1890_b0 , w_5823 );
and ( w_5823 , w_5822 , \1890_b1 );
or ( \1892_b1 , \1878_b1 , \1891_b1 );
not ( \1891_b1 , w_5824 );
and ( \1892_b0 , \1878_b0 , w_5825 );
and ( w_5824 , w_5825 , \1891_b0 );
or ( \1893_b1 , \1872_b1 , \1877_b1 );
not ( \1877_b1 , w_5826 );
and ( \1893_b0 , \1872_b0 , w_5827 );
and ( w_5826 , w_5827 , \1877_b0 );
or ( \1894_b1 , \1892_b1 , w_5828 );
or ( \1894_b0 , \1892_b0 , \1893_b0 );
not ( \1893_b0 , w_5829 );
and ( w_5829 , w_5828 , \1893_b1 );
or ( \1895_b1 , \1868_b1 , \1894_b1 );
xor ( \1895_b0 , \1868_b0 , w_5830 );
not ( w_5830 , w_5831 );
and ( w_5831 , \1894_b1 , \1894_b0 );
or ( \1896_b1 , \1729_b1 , \1789_b1 );
xor ( \1896_b0 , \1729_b0 , w_5832 );
not ( w_5832 , w_5833 );
and ( w_5833 , \1789_b1 , \1789_b0 );
or ( \1897_b1 , \1896_b1 , \1792_b1 );
xor ( \1897_b0 , \1896_b0 , w_5834 );
not ( w_5834 , w_5835 );
and ( w_5835 , \1792_b1 , \1792_b0 );
or ( \1898_b1 , \1895_b1 , \1897_b1 );
not ( \1897_b1 , w_5836 );
and ( \1898_b0 , \1895_b0 , w_5837 );
and ( w_5836 , w_5837 , \1897_b0 );
or ( \1899_b1 , \1868_b1 , \1894_b1 );
not ( \1894_b1 , w_5838 );
and ( \1899_b0 , \1868_b0 , w_5839 );
and ( w_5838 , w_5839 , \1894_b0 );
or ( \1900_b1 , \1898_b1 , w_5840 );
or ( \1900_b0 , \1898_b0 , \1899_b0 );
not ( \1899_b0 , w_5841 );
and ( w_5841 , w_5840 , \1899_b1 );
or ( \1901_b1 , \1866_b1 , w_5843 );
not ( w_5843 , w_5844 );
and ( \1901_b0 , \1866_b0 , w_5845 );
and ( w_5844 ,  , w_5845 );
buf ( w_5843 , \1900_b1 );
not ( w_5843 , w_5846 );
not (  , w_5847 );
and ( w_5846 , w_5847 , \1900_b0 );
or ( \1902_b1 , \1868_b1 , \1894_b1 );
xor ( \1902_b0 , \1868_b0 , w_5848 );
not ( w_5848 , w_5849 );
and ( w_5849 , \1894_b1 , \1894_b0 );
or ( \1903_b1 , \1902_b1 , \1897_b1 );
xor ( \1903_b0 , \1902_b0 , w_5850 );
not ( w_5850 , w_5851 );
and ( w_5851 , \1897_b1 , \1897_b0 );
buf ( \1904_b1 , \1761_b1 );
not ( \1904_b1 , w_5852 );
not ( \1904_b0 , w_5853 );
and ( w_5852 , w_5853 , \1761_b0 );
buf ( \1905_b1 , \1787_b1 );
not ( \1905_b1 , w_5854 );
not ( \1905_b0 , w_5855 );
and ( w_5854 , w_5855 , \1787_b0 );
or ( \1906_b1 , \1904_b1 , w_5856 );
or ( \1906_b0 , \1904_b0 , \1905_b0 );
not ( \1905_b0 , w_5857 );
and ( w_5857 , w_5856 , \1905_b1 );
buf ( \1907_b1 , \1787_b1 );
not ( \1907_b1 , w_5858 );
not ( \1907_b0 , w_5859 );
and ( w_5858 , w_5859 , \1787_b0 );
or ( \1908_b1 , \1907_b1 , w_5861 );
not ( w_5861 , w_5862 );
and ( \1908_b0 , \1907_b0 , w_5863 );
and ( w_5862 ,  , w_5863 );
buf ( w_5861 , \1762_b1 );
not ( w_5861 , w_5864 );
not (  , w_5865 );
and ( w_5864 , w_5865 , \1762_b0 );
or ( \1909_b1 , \1906_b1 , w_5867 );
not ( w_5867 , w_5868 );
and ( \1909_b0 , \1906_b0 , w_5869 );
and ( w_5868 ,  , w_5869 );
buf ( w_5867 , \1908_b1 );
not ( w_5867 , w_5870 );
not (  , w_5871 );
and ( w_5870 , w_5871 , \1908_b0 );
or ( \1910_b1 , \1909_b1 , \1776_b1 );
xor ( \1910_b0 , \1909_b0 , w_5872 );
not ( w_5872 , w_5873 );
and ( w_5873 , \1776_b1 , \1776_b0 );
buf ( \1911_b1 , \1910_b1 );
not ( \1911_b1 , w_5874 );
not ( \1911_b0 , w_5875 );
and ( w_5874 , w_5875 , \1910_b0 );
or ( \1912_b1 , \c[1]_b1 , \b[6]_b1 );
xor ( \1912_b0 , \c[1]_b0 , w_5876 );
not ( w_5876 , w_5877 );
and ( w_5877 , \b[6]_b1 , \b[6]_b0 );
buf ( \1913_b1 , \1912_b1 );
not ( \1913_b1 , w_5878 );
not ( \1913_b0 , w_5879 );
and ( w_5878 , w_5879 , \1912_b0 );
buf ( \1914_b1 , \1756_b1 );
not ( \1914_b1 , w_5880 );
not ( \1914_b0 , w_5881 );
and ( w_5880 , w_5881 , \1756_b0 );
or ( \1915_b1 , \1913_b1 , w_5882 );
or ( \1915_b0 , \1913_b0 , \1914_b0 );
not ( \1914_b0 , w_5883 );
and ( w_5883 , w_5882 , \1914_b1 );
or ( \1916_b1 , \1880_b1 , w_5885 );
not ( w_5885 , w_5886 );
and ( \1916_b0 , \1880_b0 , w_5887 );
and ( w_5886 ,  , w_5887 );
buf ( w_5885 , \c[0]_b1 );
not ( w_5885 , w_5888 );
not (  , w_5889 );
and ( w_5888 , w_5889 , \c[0]_b0 );
or ( \1917_b1 , \1915_b1 , w_5891 );
not ( w_5891 , w_5892 );
and ( \1917_b0 , \1915_b0 , w_5893 );
and ( w_5892 ,  , w_5893 );
buf ( w_5891 , \1916_b1 );
not ( w_5891 , w_5894 );
not (  , w_5895 );
and ( w_5894 , w_5895 , \1916_b0 );
or ( \1918_b1 , \b[0]_b1 , w_5896 );
or ( \1918_b0 , \b[0]_b0 , \c[6]_b0 );
not ( \c[6]_b0 , w_5897 );
and ( w_5897 , w_5896 , \c[6]_b1 );
or ( \1919_b1 , \1918_b1 , w_5899 );
not ( w_5899 , w_5900 );
and ( \1919_b0 , \1918_b0 , w_5901 );
and ( w_5900 ,  , w_5901 );
buf ( w_5899 , \c[5]_b1 );
not ( w_5899 , w_5902 );
not (  , w_5903 );
and ( w_5902 , w_5903 , \c[5]_b0 );
or ( \1920_b1 , \b[0]_b1 , w_5905 );
not ( w_5905 , w_5906 );
and ( \1920_b0 , \b[0]_b0 , w_5907 );
and ( w_5906 ,  , w_5907 );
buf ( w_5905 , \c[6]_b1 );
not ( w_5905 , w_5908 );
not (  , w_5909 );
and ( w_5908 , w_5909 , \c[6]_b0 );
or ( \1922_b1 , \1917_b1 , w_5911 );
not ( w_5911 , w_5912 );
and ( \1922_b0 , \1917_b0 , w_5913 );
and ( w_5912 ,  , w_5913 );
buf ( w_5911 , \1921_b1 );
not ( w_5911 , w_5914 );
not (  , w_5915 );
and ( w_5914 , w_5915 , \1921_b0 );
or ( \1923_b1 , \b[3]_b1 , \c[5]_b1 );
xor ( \1923_b0 , \b[3]_b0 , w_5916 );
not ( w_5916 , w_5917 );
and ( w_5917 , \c[5]_b1 , \c[5]_b0 );
buf ( \1924_b1 , \1923_b1 );
not ( \1924_b1 , w_5918 );
not ( \1924_b0 , w_5919 );
and ( w_5918 , w_5919 , \1923_b0 );
buf ( \1925_b1 , \1672_b1 );
not ( \1925_b1 , w_5920 );
not ( \1925_b0 , w_5921 );
and ( w_5920 , w_5921 , \1672_b0 );
or ( \1926_b1 , \1925_b1 , w_5923 );
not ( w_5923 , w_5924 );
and ( \1926_b0 , \1925_b0 , w_5925 );
and ( w_5924 ,  , w_5925 );
buf ( w_5923 , \1674_b1 );
not ( w_5923 , w_5926 );
not (  , w_5927 );
and ( w_5926 , w_5927 , \1674_b0 );
buf ( \1927_b1 , \1926_b1 );
not ( \1927_b1 , w_5928 );
not ( \1927_b0 , w_5929 );
and ( w_5928 , w_5929 , \1926_b0 );
or ( \1928_b1 , \1924_b1 , w_5930 );
or ( \1928_b0 , \1924_b0 , \1927_b0 );
not ( \1927_b0 , w_5931 );
and ( w_5931 , w_5930 , \1927_b1 );
or ( \1929_b1 , \1678_b1 , w_5933 );
not ( w_5933 , w_5934 );
and ( \1929_b0 , \1678_b0 , w_5935 );
and ( w_5934 ,  , w_5935 );
buf ( w_5933 , \1869_b1 );
not ( w_5933 , w_5936 );
not (  , w_5937 );
and ( w_5936 , w_5937 , \1869_b0 );
or ( \1930_b1 , \1928_b1 , w_5939 );
not ( w_5939 , w_5940 );
and ( \1930_b0 , \1928_b0 , w_5941 );
and ( w_5940 ,  , w_5941 );
buf ( w_5939 , \1929_b1 );
not ( w_5939 , w_5942 );
not (  , w_5943 );
and ( w_5942 , w_5943 , \1929_b0 );
buf ( \1931_b1 , \1930_b1 );
not ( \1931_b1 , w_5944 );
not ( \1931_b0 , w_5945 );
and ( w_5944 , w_5945 , \1930_b0 );
or ( \1932_b1 , \1922_b1 , w_5947 );
not ( w_5947 , w_5948 );
and ( \1932_b0 , \1922_b0 , w_5949 );
and ( w_5948 ,  , w_5949 );
buf ( w_5947 , \1931_b1 );
not ( w_5947 , w_5950 );
not (  , w_5951 );
and ( w_5950 , w_5951 , \1931_b0 );
or ( \1933_b1 , \b[5]_b1 , \c[3]_b1 );
xor ( \1933_b0 , \b[5]_b0 , w_5952 );
not ( w_5952 , w_5953 );
and ( w_5953 , \c[3]_b1 , \c[3]_b0 );
buf ( \1934_b1 , \1933_b1 );
not ( \1934_b1 , w_5954 );
not ( \1934_b0 , w_5955 );
and ( w_5954 , w_5955 , \1933_b0 );
buf ( \1935_b1 , \1705_b1 );
not ( \1935_b1 , w_5956 );
not ( \1935_b0 , w_5957 );
and ( w_5956 , w_5957 , \1705_b0 );
or ( \1936_b1 , \1934_b1 , w_5958 );
or ( \1936_b0 , \1934_b0 , \1935_b0 );
not ( \1935_b0 , w_5959 );
and ( w_5959 , w_5958 , \1935_b1 );
or ( \1937_b1 , \1708_b1 , w_5961 );
not ( w_5961 , w_5962 );
and ( \1937_b0 , \1708_b0 , w_5963 );
and ( w_5962 ,  , w_5963 );
buf ( w_5961 , \1719_b1 );
not ( w_5961 , w_5964 );
not (  , w_5965 );
and ( w_5964 , w_5965 , \1719_b0 );
or ( \1938_b1 , \1936_b1 , w_5967 );
not ( w_5967 , w_5968 );
and ( \1938_b0 , \1936_b0 , w_5969 );
and ( w_5968 ,  , w_5969 );
buf ( w_5967 , \1937_b1 );
not ( w_5967 , w_5970 );
not (  , w_5971 );
and ( w_5970 , w_5971 , \1937_b0 );
or ( \1939_b1 , \1932_b1 , \1938_b1 );
not ( \1938_b1 , w_5972 );
and ( \1939_b0 , \1932_b0 , w_5973 );
and ( w_5972 , w_5973 , \1938_b0 );
buf ( \1940_b1 , \1922_b1 );
not ( \1940_b1 , w_5974 );
not ( \1940_b0 , w_5975 );
and ( w_5974 , w_5975 , \1922_b0 );
or ( \1941_b1 , \1940_b1 , \1930_b1 );
not ( \1930_b1 , w_5976 );
and ( \1941_b0 , \1940_b0 , w_5977 );
and ( w_5976 , w_5977 , \1930_b0 );
or ( \1942_b1 , \1939_b1 , w_5979 );
not ( w_5979 , w_5980 );
and ( \1942_b0 , \1939_b0 , w_5981 );
and ( w_5980 ,  , w_5981 );
buf ( w_5979 , \1941_b1 );
not ( w_5979 , w_5982 );
not (  , w_5983 );
and ( w_5982 , w_5983 , \1941_b0 );
or ( \1943_b1 , \1911_b1 , w_5985 );
not ( w_5985 , w_5986 );
and ( \1943_b0 , \1911_b0 , w_5987 );
and ( w_5986 ,  , w_5987 );
buf ( w_5985 , \1942_b1 );
not ( w_5985 , w_5988 );
not (  , w_5989 );
and ( w_5988 , w_5989 , \1942_b0 );
buf ( \1944_b1 , \1943_b1 );
not ( \1944_b1 , w_5990 );
not ( \1944_b0 , w_5991 );
and ( w_5990 , w_5991 , \1943_b0 );
or ( \1945_b1 , \1872_b1 , \1877_b1 );
xor ( \1945_b0 , \1872_b0 , w_5992 );
not ( w_5992 , w_5993 );
and ( w_5993 , \1877_b1 , \1877_b0 );
or ( \1946_b1 , \1945_b1 , \1891_b1 );
xor ( \1946_b0 , \1945_b0 , w_5994 );
not ( w_5994 , w_5995 );
and ( w_5995 , \1891_b1 , \1891_b0 );
buf ( \1947_b1 , \1946_b1 );
not ( \1947_b1 , w_5996 );
not ( \1947_b0 , w_5997 );
and ( w_5996 , w_5997 , \1946_b0 );
buf ( \1948_b1 , \1947_b1 );
not ( \1948_b1 , w_5998 );
not ( \1948_b0 , w_5999 );
and ( w_5998 , w_5999 , \1947_b0 );
or ( \1949_b1 , \1944_b1 , w_6000 );
or ( \1949_b0 , \1944_b0 , \1948_b0 );
not ( \1948_b0 , w_6001 );
and ( w_6001 , w_6000 , \1948_b1 );
buf ( \1950_b1 , \1942_b1 );
not ( \1950_b1 , w_6002 );
not ( \1950_b0 , w_6003 );
and ( w_6002 , w_6003 , \1942_b0 );
or ( \1951_b1 , \1950_b1 , w_6005 );
not ( w_6005 , w_6006 );
and ( \1951_b0 , \1950_b0 , w_6007 );
and ( w_6006 ,  , w_6007 );
buf ( w_6005 , \1910_b1 );
not ( w_6005 , w_6008 );
not (  , w_6009 );
and ( w_6008 , w_6009 , \1910_b0 );
or ( \1952_b1 , \1949_b1 , w_6011 );
not ( w_6011 , w_6012 );
and ( \1952_b0 , \1949_b0 , w_6013 );
and ( w_6012 ,  , w_6013 );
buf ( w_6011 , \1951_b1 );
not ( w_6011 , w_6014 );
not (  , w_6015 );
and ( w_6014 , w_6015 , \1951_b0 );
buf ( \1953_b1 , \1952_b1 );
not ( \1953_b1 , w_6016 );
not ( \1953_b0 , w_6017 );
and ( w_6016 , w_6017 , \1952_b0 );
or ( \1954_b1 , \1903_b1 , w_6019 );
not ( w_6019 , w_6020 );
and ( \1954_b0 , \1903_b0 , w_6021 );
and ( w_6020 ,  , w_6021 );
buf ( w_6019 , \1953_b1 );
not ( w_6019 , w_6022 );
not (  , w_6023 );
and ( w_6022 , w_6023 , \1953_b0 );
or ( \1955_b1 , \1879_b1 , \1883_b1 );
xor ( \1955_b0 , \1879_b0 , w_6024 );
not ( w_6024 , w_6025 );
and ( w_6025 , \1883_b1 , \1883_b0 );
or ( \1956_b1 , \1955_b1 , \1888_b1 );
xor ( \1956_b0 , \1955_b0 , w_6026 );
not ( w_6026 , w_6027 );
and ( w_6027 , \1888_b1 , \1888_b0 );
buf ( \1957_b1 , \1956_b1 );
not ( \1957_b1 , w_6028 );
not ( \1957_b0 , w_6029 );
and ( w_6028 , w_6029 , \1956_b0 );
buf ( \1958_b1 , \1957_b1 );
not ( \1958_b1 , w_6030 );
not ( \1958_b0 , w_6031 );
and ( w_6030 , w_6031 , \1957_b0 );
or ( \1959_b1 , \b[4]_b1 , \c[3]_b1 );
xor ( \1959_b0 , \b[4]_b0 , w_6032 );
not ( w_6032 , w_6033 );
and ( w_6033 , \c[3]_b1 , \c[3]_b0 );
buf ( \1960_b1 , \1959_b1 );
not ( \1960_b1 , w_6034 );
not ( \1960_b0 , w_6035 );
and ( w_6034 , w_6035 , \1959_b0 );
buf ( \1961_b1 , \1705_b1 );
not ( \1961_b1 , w_6036 );
not ( \1961_b0 , w_6037 );
and ( w_6036 , w_6037 , \1705_b0 );
or ( \1962_b1 , \1960_b1 , w_6038 );
or ( \1962_b0 , \1960_b0 , \1961_b0 );
not ( \1961_b0 , w_6039 );
and ( w_6039 , w_6038 , \1961_b1 );
or ( \1963_b1 , \1708_b1 , w_6041 );
not ( w_6041 , w_6042 );
and ( \1963_b0 , \1708_b0 , w_6043 );
and ( w_6042 ,  , w_6043 );
buf ( w_6041 , \1933_b1 );
not ( w_6041 , w_6044 );
not (  , w_6045 );
and ( w_6044 , w_6045 , \1933_b0 );
or ( \1964_b1 , \1962_b1 , w_6047 );
not ( w_6047 , w_6048 );
and ( \1964_b0 , \1962_b0 , w_6049 );
and ( w_6048 ,  , w_6049 );
buf ( w_6047 , \1963_b1 );
not ( w_6047 , w_6050 );
not (  , w_6051 );
and ( w_6050 , w_6051 , \1963_b0 );
or ( \1965_b1 , \b[2]_b1 , \c[5]_b1 );
xor ( \1965_b0 , \b[2]_b0 , w_6052 );
not ( w_6052 , w_6053 );
and ( w_6053 , \c[5]_b1 , \c[5]_b0 );
buf ( \1966_b1 , \1965_b1 );
not ( \1966_b1 , w_6054 );
not ( \1966_b0 , w_6055 );
and ( w_6054 , w_6055 , \1965_b0 );
buf ( \1967_b1 , \1926_b1 );
not ( \1967_b1 , w_6056 );
not ( \1967_b0 , w_6057 );
and ( w_6056 , w_6057 , \1926_b0 );
or ( \1968_b1 , \1966_b1 , w_6058 );
or ( \1968_b0 , \1966_b0 , \1967_b0 );
not ( \1967_b0 , w_6059 );
and ( w_6059 , w_6058 , \1967_b1 );
or ( \1969_b1 , \1678_b1 , w_6061 );
not ( w_6061 , w_6062 );
and ( \1969_b0 , \1678_b0 , w_6063 );
and ( w_6062 ,  , w_6063 );
buf ( w_6061 , \1923_b1 );
not ( w_6061 , w_6064 );
not (  , w_6065 );
and ( w_6064 , w_6065 , \1923_b0 );
or ( \1970_b1 , \1968_b1 , w_6067 );
not ( w_6067 , w_6068 );
and ( \1970_b0 , \1968_b0 , w_6069 );
and ( w_6068 ,  , w_6069 );
buf ( w_6067 , \1969_b1 );
not ( w_6067 , w_6070 );
not (  , w_6071 );
and ( w_6070 , w_6071 , \1969_b0 );
or ( \1971_b1 , \1964_b1 , w_6072 );
or ( \1971_b0 , \1964_b0 , \1970_b0 );
not ( \1970_b0 , w_6073 );
and ( w_6073 , w_6072 , \1970_b1 );
or ( \1972_b1 , \b[0]_b1 , \c[7]_b1 );
xor ( \1972_b0 , \b[0]_b0 , w_6074 );
not ( w_6074 , w_6075 );
and ( w_6075 , \c[7]_b1 , \c[7]_b0 );
buf ( \1973_b1 , \1972_b1 );
not ( \1973_b1 , w_6076 );
not ( \1973_b0 , w_6077 );
and ( w_6076 , w_6077 , \1972_b0 );
buf ( \1974_b1 , \1743_b1 );
not ( \1974_b1 , w_6078 );
not ( \1974_b0 , w_6079 );
and ( w_6078 , w_6079 , \1743_b0 );
or ( \1975_b1 , \1973_b1 , w_6080 );
or ( \1975_b0 , \1973_b0 , \1974_b0 );
not ( \1974_b0 , w_6081 );
and ( w_6081 , w_6080 , \1974_b1 );
or ( \1976_b1 , \1747_b1 , w_6083 );
not ( w_6083 , w_6084 );
and ( \1976_b0 , \1747_b0 , w_6085 );
and ( w_6084 ,  , w_6085 );
buf ( w_6083 , \1885_b1 );
not ( w_6083 , w_6086 );
not (  , w_6087 );
and ( w_6086 , w_6087 , \1885_b0 );
or ( \1977_b1 , \1975_b1 , w_6089 );
not ( w_6089 , w_6090 );
and ( \1977_b0 , \1975_b0 , w_6091 );
and ( w_6090 ,  , w_6091 );
buf ( w_6089 , \1976_b1 );
not ( w_6089 , w_6092 );
not (  , w_6093 );
and ( w_6092 , w_6093 , \1976_b0 );
or ( \1978_b1 , \1971_b1 , w_6095 );
not ( w_6095 , w_6096 );
and ( \1978_b0 , \1971_b0 , w_6097 );
and ( w_6096 ,  , w_6097 );
buf ( w_6095 , \1977_b1 );
not ( w_6095 , w_6098 );
not (  , w_6099 );
and ( w_6098 , w_6099 , \1977_b0 );
or ( \1979_b1 , \1964_b1 , w_6101 );
not ( w_6101 , w_6102 );
and ( \1979_b0 , \1964_b0 , w_6103 );
and ( w_6102 ,  , w_6103 );
buf ( w_6101 , \1970_b1 );
not ( w_6101 , w_6104 );
not (  , w_6105 );
and ( w_6104 , w_6105 , \1970_b0 );
or ( \1980_b1 , \1978_b1 , w_6107 );
not ( w_6107 , w_6108 );
and ( \1980_b0 , \1978_b0 , w_6109 );
and ( w_6108 ,  , w_6109 );
buf ( w_6107 , \1979_b1 );
not ( w_6107 , w_6110 );
not (  , w_6111 );
and ( w_6110 , w_6111 , \1979_b0 );
buf ( \1981_b1 , \1980_b1 );
not ( \1981_b1 , w_6112 );
not ( \1981_b0 , w_6113 );
and ( w_6112 , w_6113 , \1980_b0 );
buf ( \1982_b1 , \1981_b1 );
not ( \1982_b1 , w_6114 );
not ( \1982_b0 , w_6115 );
and ( w_6114 , w_6115 , \1981_b0 );
or ( \1983_b1 , \1958_b1 , w_6116 );
or ( \1983_b0 , \1958_b0 , \1982_b0 );
not ( \1982_b0 , w_6117 );
and ( w_6117 , w_6116 , \1982_b1 );
or ( \1984_b1 , \1980_b1 , w_6119 );
not ( w_6119 , w_6120 );
and ( \1984_b0 , \1980_b0 , w_6121 );
and ( w_6120 ,  , w_6121 );
buf ( w_6119 , \1956_b1 );
not ( w_6119 , w_6122 );
not (  , w_6123 );
and ( w_6122 , w_6123 , \1956_b0 );
or ( \1985_b1 , \1983_b1 , w_6125 );
not ( w_6125 , w_6126 );
and ( \1985_b0 , \1983_b0 , w_6127 );
and ( w_6126 ,  , w_6127 );
buf ( w_6125 , \1984_b1 );
not ( w_6125 , w_6128 );
not (  , w_6129 );
and ( w_6128 , w_6129 , \1984_b0 );
buf ( \1986_b1 , \1931_b1 );
not ( \1986_b1 , w_6130 );
not ( \1986_b0 , w_6131 );
and ( w_6130 , w_6131 , \1931_b0 );
buf ( \1987_b1 , \1940_b1 );
not ( \1987_b1 , w_6132 );
not ( \1987_b0 , w_6133 );
and ( w_6132 , w_6133 , \1940_b0 );
or ( \1988_b1 , \1986_b1 , w_6134 );
or ( \1988_b0 , \1986_b0 , \1987_b0 );
not ( \1987_b0 , w_6135 );
and ( w_6135 , w_6134 , \1987_b1 );
or ( \1989_b1 , \1940_b1 , w_6136 );
or ( \1989_b0 , \1940_b0 , \1931_b0 );
not ( \1931_b0 , w_6137 );
and ( w_6137 , w_6136 , \1931_b1 );
or ( \1990_b1 , \1988_b1 , w_6139 );
not ( w_6139 , w_6140 );
and ( \1990_b0 , \1988_b0 , w_6141 );
and ( w_6140 ,  , w_6141 );
buf ( w_6139 , \1989_b1 );
not ( w_6139 , w_6142 );
not (  , w_6143 );
and ( w_6142 , w_6143 , \1989_b0 );
buf ( \1991_b1 , \1938_b1 );
not ( \1991_b1 , w_6144 );
not ( \1991_b0 , w_6145 );
and ( w_6144 , w_6145 , \1938_b0 );
or ( \1992_b1 , \1990_b1 , \1991_b1 );
not ( \1991_b1 , w_6146 );
and ( \1992_b0 , \1990_b0 , w_6147 );
and ( w_6146 , w_6147 , \1991_b0 );
buf ( \1993_b1 , \1990_b1 );
not ( \1993_b1 , w_6148 );
not ( \1993_b0 , w_6149 );
and ( w_6148 , w_6149 , \1990_b0 );
or ( \1994_b1 , \1993_b1 , \1938_b1 );
not ( \1938_b1 , w_6150 );
and ( \1994_b0 , \1993_b0 , w_6151 );
and ( w_6150 , w_6151 , \1938_b0 );
or ( \1995_b1 , \1992_b1 , w_6153 );
not ( w_6153 , w_6154 );
and ( \1995_b0 , \1992_b0 , w_6155 );
and ( w_6154 ,  , w_6155 );
buf ( w_6153 , \1994_b1 );
not ( w_6153 , w_6156 );
not (  , w_6157 );
and ( w_6156 , w_6157 , \1994_b0 );
or ( \1996_b1 , \1985_b1 , \1995_b1 );
not ( \1995_b1 , w_6158 );
and ( \1996_b0 , \1985_b0 , w_6159 );
and ( w_6158 , w_6159 , \1995_b0 );
buf ( \1997_b1 , \1985_b1 );
not ( \1997_b1 , w_6160 );
not ( \1997_b0 , w_6161 );
and ( w_6160 , w_6161 , \1985_b0 );
buf ( \1998_b1 , \1995_b1 );
not ( \1998_b1 , w_6162 );
not ( \1998_b0 , w_6163 );
and ( w_6162 , w_6163 , \1995_b0 );
or ( \1999_b1 , \1997_b1 , \1998_b1 );
not ( \1998_b1 , w_6164 );
and ( \1999_b0 , \1997_b0 , w_6165 );
and ( w_6164 , w_6165 , \1998_b0 );
or ( \2000_b1 , \1996_b1 , w_6167 );
not ( w_6167 , w_6168 );
and ( \2000_b0 , \1996_b0 , w_6169 );
and ( w_6168 ,  , w_6169 );
buf ( w_6167 , \1999_b1 );
not ( w_6167 , w_6170 );
not (  , w_6171 );
and ( w_6170 , w_6171 , \1999_b0 );
or ( \2001_b1 , \1917_b1 , w_6172 );
xor ( \2001_b0 , \1917_b0 , w_6174 );
not ( w_6174 , w_6175 );
and ( w_6175 , w_6172 , w_6173 );
buf ( w_6172 , \1921_b1 );
not ( w_6172 , w_6176 );
not ( w_6173 , w_6177 );
and ( w_6176 , w_6177 , \1921_b0 );
or ( \2002_b1 , \b[3]_b1 , \c[3]_b1 );
xor ( \2002_b0 , \b[3]_b0 , w_6178 );
not ( w_6178 , w_6179 );
and ( w_6179 , \c[3]_b1 , \c[3]_b0 );
buf ( \2003_b1 , \2002_b1 );
not ( \2003_b1 , w_6180 );
not ( \2003_b0 , w_6181 );
and ( w_6180 , w_6181 , \2002_b0 );
buf ( \2004_b1 , \1705_b1 );
not ( \2004_b1 , w_6182 );
not ( \2004_b0 , w_6183 );
and ( w_6182 , w_6183 , \1705_b0 );
or ( \2005_b1 , \2003_b1 , w_6184 );
or ( \2005_b0 , \2003_b0 , \2004_b0 );
not ( \2004_b0 , w_6185 );
and ( w_6185 , w_6184 , \2004_b1 );
or ( \2006_b1 , \1725_b1 , w_6187 );
not ( w_6187 , w_6188 );
and ( \2006_b0 , \1725_b0 , w_6189 );
and ( w_6188 ,  , w_6189 );
buf ( w_6187 , \1959_b1 );
not ( w_6187 , w_6190 );
not (  , w_6191 );
and ( w_6190 , w_6191 , \1959_b0 );
or ( \2007_b1 , \2005_b1 , w_6193 );
not ( w_6193 , w_6194 );
and ( \2007_b0 , \2005_b0 , w_6195 );
and ( w_6194 ,  , w_6195 );
buf ( w_6193 , \2006_b1 );
not ( w_6193 , w_6196 );
not (  , w_6197 );
and ( w_6196 , w_6197 , \2006_b0 );
or ( \2008_b1 , \b[5]_b1 , \c[1]_b1 );
xor ( \2008_b0 , \b[5]_b0 , w_6198 );
not ( w_6198 , w_6199 );
and ( w_6199 , \c[1]_b1 , \c[1]_b0 );
buf ( \2009_b1 , \2008_b1 );
not ( \2009_b1 , w_6200 );
not ( \2009_b0 , w_6201 );
and ( w_6200 , w_6201 , \2008_b0 );
buf ( \2010_b1 , \1756_b1 );
not ( \2010_b1 , w_6202 );
not ( \2010_b0 , w_6203 );
and ( w_6202 , w_6203 , \1756_b0 );
or ( \2011_b1 , \2009_b1 , w_6204 );
or ( \2011_b0 , \2009_b0 , \2010_b0 );
not ( \2010_b0 , w_6205 );
and ( w_6205 , w_6204 , \2010_b1 );
or ( \2012_b1 , \1912_b1 , w_6207 );
not ( w_6207 , w_6208 );
and ( \2012_b0 , \1912_b0 , w_6209 );
and ( w_6208 ,  , w_6209 );
buf ( w_6207 , \c[0]_b1 );
not ( w_6207 , w_6210 );
not (  , w_6211 );
and ( w_6210 , w_6211 , \c[0]_b0 );
or ( \2013_b1 , \2011_b1 , w_6213 );
not ( w_6213 , w_6214 );
and ( \2013_b0 , \2011_b0 , w_6215 );
and ( w_6214 ,  , w_6215 );
buf ( w_6213 , \2012_b1 );
not ( w_6213 , w_6216 );
not (  , w_6217 );
and ( w_6216 , w_6217 , \2012_b0 );
buf ( \2014_b1 , \2013_b1 );
not ( \2014_b1 , w_6218 );
not ( \2014_b0 , w_6219 );
and ( w_6218 , w_6219 , \2013_b0 );
or ( \2015_b1 , \1742_b1 , w_6221 );
not ( w_6221 , w_6222 );
and ( \2015_b0 , \1742_b0 , w_6223 );
and ( w_6222 ,  , w_6223 );
buf ( w_6221 , \b[0]_b1 );
not ( w_6221 , w_6224 );
not (  , w_6225 );
and ( w_6224 , w_6225 , \b[0]_b0 );
or ( \2016_b1 , \2014_b1 , w_6227 );
not ( w_6227 , w_6228 );
and ( \2016_b0 , \2014_b0 , w_6229 );
and ( w_6228 ,  , w_6229 );
buf ( w_6227 , \2015_b1 );
not ( w_6227 , w_6230 );
not (  , w_6231 );
and ( w_6230 , w_6231 , \2015_b0 );
or ( \2017_b1 , \2007_b1 , \2016_b1 );
not ( \2016_b1 , w_6232 );
and ( \2017_b0 , \2007_b0 , w_6233 );
and ( w_6232 , w_6233 , \2016_b0 );
buf ( \2018_b1 , \2013_b1 );
not ( \2018_b1 , w_6234 );
not ( \2018_b0 , w_6235 );
and ( w_6234 , w_6235 , \2013_b0 );
or ( \2019_b1 , \2018_b1 , w_6237 );
not ( w_6237 , w_6238 );
and ( \2019_b0 , \2018_b0 , w_6239 );
and ( w_6238 ,  , w_6239 );
buf ( w_6237 , \2015_b1 );
not ( w_6237 , w_6240 );
not (  , w_6241 );
and ( w_6240 , w_6241 , \2015_b0 );
or ( \2020_b1 , \2017_b1 , w_6243 );
not ( w_6243 , w_6244 );
and ( \2020_b0 , \2017_b0 , w_6245 );
and ( w_6244 ,  , w_6245 );
buf ( w_6243 , \2019_b1 );
not ( w_6243 , w_6246 );
not (  , w_6247 );
and ( w_6246 , w_6247 , \2019_b0 );
or ( \2021_b1 , \2001_b1 , \2020_b1 );
xor ( \2021_b0 , \2001_b0 , w_6248 );
not ( w_6248 , w_6249 );
and ( w_6249 , \2020_b1 , \2020_b0 );
or ( \2022_b1 , \1977_b1 , \1970_b1 );
xor ( \2022_b0 , \1977_b0 , w_6250 );
not ( w_6250 , w_6251 );
and ( w_6251 , \1970_b1 , \1970_b0 );
or ( \2023_b1 , \2022_b1 , w_6252 );
xor ( \2023_b0 , \2022_b0 , w_6254 );
not ( w_6254 , w_6255 );
and ( w_6255 , w_6252 , w_6253 );
buf ( w_6252 , \1964_b1 );
not ( w_6252 , w_6256 );
not ( w_6253 , w_6257 );
and ( w_6256 , w_6257 , \1964_b0 );
or ( \2024_b1 , \2021_b1 , \2023_b1 );
not ( \2023_b1 , w_6258 );
and ( \2024_b0 , \2021_b0 , w_6259 );
and ( w_6258 , w_6259 , \2023_b0 );
or ( \2025_b1 , \2001_b1 , \2020_b1 );
not ( \2020_b1 , w_6260 );
and ( \2025_b0 , \2001_b0 , w_6261 );
and ( w_6260 , w_6261 , \2020_b0 );
or ( \2026_b1 , \2024_b1 , w_6262 );
or ( \2026_b0 , \2024_b0 , \2025_b0 );
not ( \2025_b0 , w_6263 );
and ( w_6263 , w_6262 , \2025_b1 );
or ( \2027_b1 , \2000_b1 , w_6265 );
not ( w_6265 , w_6266 );
and ( \2027_b0 , \2000_b0 , w_6267 );
and ( w_6266 ,  , w_6267 );
buf ( w_6265 , \2026_b1 );
not ( w_6265 , w_6268 );
not (  , w_6269 );
and ( w_6268 , w_6269 , \2026_b0 );
buf ( \2028_b1 , \2027_b1 );
not ( \2028_b1 , w_6270 );
not ( \2028_b0 , w_6271 );
and ( w_6270 , w_6271 , \2027_b0 );
buf ( \2029_b1 , \1942_b1 );
not ( \2029_b1 , w_6272 );
not ( \2029_b0 , w_6273 );
and ( w_6272 , w_6273 , \1942_b0 );
buf ( \2030_b1 , \1910_b1 );
not ( \2030_b1 , w_6274 );
not ( \2030_b0 , w_6275 );
and ( w_6274 , w_6275 , \1910_b0 );
or ( \2031_b1 , \2029_b1 , w_6276 );
or ( \2031_b0 , \2029_b0 , \2030_b0 );
not ( \2030_b0 , w_6277 );
and ( w_6277 , w_6276 , \2030_b1 );
or ( \2032_b1 , \1942_b1 , w_6278 );
or ( \2032_b0 , \1942_b0 , \1910_b0 );
not ( \1910_b0 , w_6279 );
and ( w_6279 , w_6278 , \1910_b1 );
or ( \2033_b1 , \2031_b1 , w_6281 );
not ( w_6281 , w_6282 );
and ( \2033_b0 , \2031_b0 , w_6283 );
and ( w_6282 ,  , w_6283 );
buf ( w_6281 , \2032_b1 );
not ( w_6281 , w_6284 );
not (  , w_6285 );
and ( w_6284 , w_6285 , \2032_b0 );
buf ( \2034_b1 , \2033_b1 );
not ( \2034_b1 , w_6286 );
not ( \2034_b0 , w_6287 );
and ( w_6286 , w_6287 , \2033_b0 );
buf ( \2035_b1 , \2034_b1 );
not ( \2035_b1 , w_6288 );
not ( \2035_b0 , w_6289 );
and ( w_6288 , w_6289 , \2034_b0 );
buf ( \2036_b1 , \1947_b1 );
not ( \2036_b1 , w_6290 );
not ( \2036_b0 , w_6291 );
and ( w_6290 , w_6291 , \1947_b0 );
or ( \2037_b1 , \2035_b1 , w_6292 );
or ( \2037_b0 , \2035_b0 , \2036_b0 );
not ( \2036_b0 , w_6293 );
and ( w_6293 , w_6292 , \2036_b1 );
or ( \2038_b1 , \1946_b1 , w_6295 );
not ( w_6295 , w_6296 );
and ( \2038_b0 , \1946_b0 , w_6297 );
and ( w_6296 ,  , w_6297 );
buf ( w_6295 , \2033_b1 );
not ( w_6295 , w_6298 );
not (  , w_6299 );
and ( w_6298 , w_6299 , \2033_b0 );
or ( \2039_b1 , \2037_b1 , w_6301 );
not ( w_6301 , w_6302 );
and ( \2039_b0 , \2037_b0 , w_6303 );
and ( w_6302 ,  , w_6303 );
buf ( w_6301 , \2038_b1 );
not ( w_6301 , w_6304 );
not (  , w_6305 );
and ( w_6304 , w_6305 , \2038_b0 );
buf ( \2040_b1 , \1957_b1 );
not ( \2040_b1 , w_6306 );
not ( \2040_b0 , w_6307 );
and ( w_6306 , w_6307 , \1957_b0 );
buf ( \2041_b1 , \1998_b1 );
not ( \2041_b1 , w_6308 );
not ( \2041_b0 , w_6309 );
and ( w_6308 , w_6309 , \1998_b0 );
or ( \2042_b1 , \2040_b1 , w_6310 );
or ( \2042_b0 , \2040_b0 , \2041_b0 );
not ( \2041_b0 , w_6311 );
and ( w_6311 , w_6310 , \2041_b1 );
buf ( \2043_b1 , \1995_b1 );
not ( \2043_b1 , w_6312 );
not ( \2043_b0 , w_6313 );
and ( w_6312 , w_6313 , \1995_b0 );
buf ( \2044_b1 , \1956_b1 );
not ( \2044_b1 , w_6314 );
not ( \2044_b0 , w_6315 );
and ( w_6314 , w_6315 , \1956_b0 );
or ( \2045_b1 , \2043_b1 , w_6316 );
or ( \2045_b0 , \2043_b0 , \2044_b0 );
not ( \2044_b0 , w_6317 );
and ( w_6317 , w_6316 , \2044_b1 );
or ( \2046_b1 , \2045_b1 , w_6319 );
not ( w_6319 , w_6320 );
and ( \2046_b0 , \2045_b0 , w_6321 );
and ( w_6320 ,  , w_6321 );
buf ( w_6319 , \1980_b1 );
not ( w_6319 , w_6322 );
not (  , w_6323 );
and ( w_6322 , w_6323 , \1980_b0 );
or ( \2047_b1 , \2042_b1 , w_6325 );
not ( w_6325 , w_6326 );
and ( \2047_b0 , \2042_b0 , w_6327 );
and ( w_6326 ,  , w_6327 );
buf ( w_6325 , \2046_b1 );
not ( w_6325 , w_6328 );
not (  , w_6329 );
and ( w_6328 , w_6329 , \2046_b0 );
or ( \2048_b1 , \2039_b1 , w_6331 );
not ( w_6331 , w_6332 );
and ( \2048_b0 , \2039_b0 , w_6333 );
and ( w_6332 ,  , w_6333 );
buf ( w_6331 , \2047_b1 );
not ( w_6331 , w_6334 );
not (  , w_6335 );
and ( w_6334 , w_6335 , \2047_b0 );
or ( \2049_b1 , \2028_b1 , w_6337 );
not ( w_6337 , w_6338 );
and ( \2049_b0 , \2028_b0 , w_6339 );
and ( w_6338 ,  , w_6339 );
buf ( w_6337 , \2048_b1 );
not ( w_6337 , w_6340 );
not (  , w_6341 );
and ( w_6340 , w_6341 , \2048_b0 );
buf ( \2051_b1 , \1679_b1 );
not ( \2051_b1 , w_6342 );
not ( \2051_b0 , w_6343 );
and ( w_6342 , w_6343 , \1679_b0 );
buf ( \2052_b1 , \1675_b1 );
buf ( \2052_b0 , \1675_b0 );
buf ( \2053_b1 , \2052_b1 );
not ( \2053_b1 , w_6344 );
not ( \2053_b0 , w_6345 );
and ( w_6344 , w_6345 , \2052_b0 );
or ( \2054_b1 , \2051_b1 , w_6346 );
or ( \2054_b0 , \2051_b0 , \2053_b0 );
not ( \2053_b0 , w_6347 );
and ( w_6347 , w_6346 , \2053_b1 );
or ( \2055_b1 , \b[8]_b1 , \c[5]_b1 );
xor ( \2055_b0 , \b[8]_b0 , w_6348 );
not ( w_6348 , w_6349 );
and ( w_6349 , \c[5]_b1 , \c[5]_b0 );
or ( \2056_b1 , \1678_b1 , w_6351 );
not ( w_6351 , w_6352 );
and ( \2056_b0 , \1678_b0 , w_6353 );
and ( w_6352 ,  , w_6353 );
buf ( w_6351 , \2055_b1 );
not ( w_6351 , w_6354 );
not (  , w_6355 );
and ( w_6354 , w_6355 , \2055_b0 );
or ( \2057_b1 , \2054_b1 , w_6357 );
not ( w_6357 , w_6358 );
and ( \2057_b0 , \2054_b0 , w_6359 );
and ( w_6358 ,  , w_6359 );
buf ( w_6357 , \2056_b1 );
not ( w_6357 , w_6360 );
not (  , w_6361 );
and ( w_6360 , w_6361 , \2056_b0 );
or ( \2058_b1 , \1698_b1 , \1711_b1 );
not ( \1711_b1 , w_6362 );
and ( \2058_b0 , \1698_b0 , w_6363 );
and ( w_6362 , w_6363 , \1711_b0 );
or ( \2059_b1 , \2057_b1 , \2058_b1 );
xor ( \2059_b0 , \2057_b0 , w_6364 );
not ( w_6364 , w_6365 );
and ( w_6365 , \2058_b1 , \2058_b0 );
buf ( \2060_b1 , \1843_b1 );
not ( \2060_b1 , w_6366 );
not ( \2060_b0 , w_6367 );
and ( w_6366 , w_6367 , \1843_b0 );
buf ( \2061_b1 , \1859_b1 );
not ( \2061_b1 , w_6368 );
not ( \2061_b0 , w_6369 );
and ( w_6368 , w_6369 , \1859_b0 );
or ( \2062_b1 , \2060_b1 , w_6370 );
or ( \2062_b0 , \2060_b0 , \2061_b0 );
not ( \2061_b0 , w_6371 );
and ( w_6371 , w_6370 , \2061_b1 );
or ( \2063_b1 , \2062_b1 , w_6373 );
not ( w_6373 , w_6374 );
and ( \2063_b0 , \2062_b0 , w_6375 );
and ( w_6374 ,  , w_6375 );
buf ( w_6373 , \1836_b1 );
not ( w_6373 , w_6376 );
not (  , w_6377 );
and ( w_6376 , w_6377 , \1836_b0 );
buf ( \2064_b1 , \1859_b1 );
not ( \2064_b1 , w_6378 );
not ( \2064_b0 , w_6379 );
and ( w_6378 , w_6379 , \1859_b0 );
or ( \2065_b1 , \2064_b1 , w_6381 );
not ( w_6381 , w_6382 );
and ( \2065_b0 , \2064_b0 , w_6383 );
and ( w_6382 ,  , w_6383 );
buf ( w_6381 , \1842_b1 );
not ( w_6381 , w_6384 );
not (  , w_6385 );
and ( w_6384 , w_6385 , \1842_b0 );
or ( \2066_b1 , \2063_b1 , w_6387 );
not ( w_6387 , w_6388 );
and ( \2066_b0 , \2063_b0 , w_6389 );
and ( w_6388 ,  , w_6389 );
buf ( w_6387 , \2065_b1 );
not ( w_6387 , w_6390 );
not (  , w_6391 );
and ( w_6390 , w_6391 , \2065_b0 );
or ( \2067_b1 , \2059_b1 , \2066_b1 );
xor ( \2067_b0 , \2059_b0 , w_6392 );
not ( w_6392 , w_6393 );
and ( w_6393 , \2066_b1 , \2066_b0 );
buf ( \2068_b1 , \1822_b1 );
not ( \2068_b1 , w_6394 );
not ( \2068_b0 , w_6395 );
and ( w_6394 , w_6395 , \1822_b0 );
buf ( \2069_b1 , \1864_b1 );
not ( \2069_b1 , w_6396 );
not ( \2069_b0 , w_6397 );
and ( w_6396 , w_6397 , \1864_b0 );
or ( \2070_b1 , \2068_b1 , w_6398 );
or ( \2070_b0 , \2068_b0 , \2069_b0 );
not ( \2069_b0 , w_6399 );
and ( w_6399 , w_6398 , \2069_b1 );
or ( \2071_b1 , \1864_b1 , w_6400 );
or ( \2071_b0 , \1864_b0 , \1822_b0 );
not ( \1822_b0 , w_6401 );
and ( w_6401 , w_6400 , \1822_b1 );
or ( \2072_b1 , \2071_b1 , w_6403 );
not ( w_6403 , w_6404 );
and ( \2072_b0 , \2071_b0 , w_6405 );
and ( w_6404 ,  , w_6405 );
buf ( w_6403 , \1829_b1 );
not ( w_6403 , w_6406 );
not (  , w_6407 );
and ( w_6406 , w_6407 , \1829_b0 );
or ( \2073_b1 , \2070_b1 , w_6409 );
not ( w_6409 , w_6410 );
and ( \2073_b0 , \2070_b0 , w_6411 );
and ( w_6410 ,  , w_6411 );
buf ( w_6409 , \2072_b1 );
not ( w_6409 , w_6412 );
not (  , w_6413 );
and ( w_6412 , w_6413 , \2072_b0 );
or ( \2074_b1 , \2067_b1 , \2073_b1 );
xor ( \2074_b0 , \2067_b0 , w_6414 );
not ( w_6414 , w_6415 );
and ( w_6415 , \2073_b1 , \2073_b0 );
or ( \2075_b1 , \c[12]_b1 , \c[11]_b1 );
xor ( \2075_b0 , \c[12]_b0 , w_6416 );
not ( w_6416 , w_6417 );
and ( w_6417 , \c[11]_b1 , \c[11]_b0 );
or ( \2076_b1 , \2075_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_6418 );
and ( \2076_b0 , \2075_b0 , w_6419 );
and ( w_6418 , w_6419 , \b[0]_b0 );
buf ( \2077_b1 , \1834_b1 );
not ( \2077_b1 , w_6420 );
not ( \2077_b0 , w_6421 );
and ( w_6420 , w_6421 , \1834_b0 );
buf ( \2078_b1 , \1782_b1 );
not ( \2078_b1 , w_6422 );
not ( \2078_b0 , w_6423 );
and ( w_6422 , w_6423 , \1782_b0 );
or ( \2079_b1 , \2077_b1 , w_6424 );
or ( \2079_b0 , \2077_b0 , \2078_b0 );
not ( \2078_b0 , w_6425 );
and ( w_6425 , w_6424 , \2078_b1 );
or ( \2080_b1 , \b[6]_b1 , \c[7]_b1 );
xor ( \2080_b0 , \b[6]_b0 , w_6426 );
not ( w_6426 , w_6427 );
and ( w_6427 , \c[7]_b1 , \c[7]_b0 );
or ( \2081_b1 , \1742_b1 , w_6429 );
not ( w_6429 , w_6430 );
and ( \2081_b0 , \1742_b0 , w_6431 );
and ( w_6430 ,  , w_6431 );
buf ( w_6429 , \2080_b1 );
not ( w_6429 , w_6432 );
not (  , w_6433 );
and ( w_6432 , w_6433 , \2080_b0 );
or ( \2082_b1 , \2079_b1 , w_6435 );
not ( w_6435 , w_6436 );
and ( \2082_b0 , \2079_b0 , w_6437 );
and ( w_6436 ,  , w_6437 );
buf ( w_6435 , \2081_b1 );
not ( w_6435 , w_6438 );
not (  , w_6439 );
and ( w_6438 , w_6439 , \2081_b0 );
or ( \2083_b1 , \2076_b1 , \2082_b1 );
xor ( \2083_b0 , \2076_b0 , w_6440 );
not ( w_6440 , w_6441 );
and ( w_6441 , \2082_b1 , \2082_b0 );
buf ( \2084_b1 , \1709_b1 );
not ( \2084_b1 , w_6442 );
not ( \2084_b0 , w_6443 );
and ( w_6442 , w_6443 , \1709_b0 );
buf ( \2085_b1 , \1722_b1 );
not ( \2085_b1 , w_6444 );
not ( \2085_b0 , w_6445 );
and ( w_6444 , w_6445 , \1722_b0 );
or ( \2086_b1 , \2084_b1 , w_6446 );
or ( \2086_b0 , \2084_b0 , \2085_b0 );
not ( \2085_b0 , w_6447 );
and ( w_6447 , w_6446 , \2085_b1 );
or ( \2087_b1 , \b[10]_b1 , \c[3]_b1 );
xor ( \2087_b0 , \b[10]_b0 , w_6448 );
not ( w_6448 , w_6449 );
and ( w_6449 , \c[3]_b1 , \c[3]_b0 );
or ( \2088_b1 , \1725_b1 , w_6451 );
not ( w_6451 , w_6452 );
and ( \2088_b0 , \1725_b0 , w_6453 );
and ( w_6452 ,  , w_6453 );
buf ( w_6451 , \2087_b1 );
not ( w_6451 , w_6454 );
not (  , w_6455 );
and ( w_6454 , w_6455 , \2087_b0 );
or ( \2089_b1 , \2086_b1 , w_6457 );
not ( w_6457 , w_6458 );
and ( \2089_b0 , \2086_b0 , w_6459 );
and ( w_6458 ,  , w_6459 );
buf ( w_6457 , \2088_b1 );
not ( w_6457 , w_6460 );
not (  , w_6461 );
and ( w_6460 , w_6461 , \2088_b0 );
or ( \2090_b1 , \2083_b1 , \2089_b1 );
xor ( \2090_b0 , \2083_b0 , w_6462 );
not ( w_6462 , w_6463 );
and ( w_6463 , \2089_b1 , \2089_b0 );
buf ( \2091_b1 , \1851_b1 );
not ( \2091_b1 , w_6464 );
not ( \2091_b0 , w_6465 );
and ( w_6464 , w_6465 , \1851_b0 );
buf ( \2092_b1 , \1857_b1 );
not ( \2092_b1 , w_6466 );
not ( \2092_b0 , w_6467 );
and ( w_6466 , w_6467 , \1857_b0 );
or ( \2093_b1 , \2091_b1 , w_6468 );
or ( \2093_b0 , \2091_b0 , \2092_b0 );
not ( \2092_b0 , w_6469 );
and ( w_6469 , w_6468 , \2092_b1 );
buf ( \2094_b1 , \c[9]_b1 );
not ( \2094_b1 , w_6470 );
not ( \2094_b0 , w_6471 );
and ( w_6470 , w_6471 , \c[9]_b0 );
or ( \2095_b1 , \b[4]_b1 , \2094_b1 );
xor ( \2095_b0 , \b[4]_b0 , w_6472 );
not ( w_6472 , w_6473 );
and ( w_6473 , \2094_b1 , \2094_b0 );
buf ( \2096_b1 , \2095_b1 );
not ( \2096_b1 , w_6474 );
not ( \2096_b0 , w_6475 );
and ( w_6474 , w_6475 , \2095_b0 );
or ( \2097_b1 , \2096_b1 , w_6477 );
not ( w_6477 , w_6478 );
and ( \2097_b0 , \2096_b0 , w_6479 );
and ( w_6478 ,  , w_6479 );
buf ( w_6477 , \1773_b1 );
not ( w_6477 , w_6480 );
not (  , w_6481 );
and ( w_6480 , w_6481 , \1773_b0 );
or ( \2098_b1 , \2093_b1 , w_6483 );
not ( w_6483 , w_6484 );
and ( \2098_b0 , \2093_b0 , w_6485 );
and ( w_6484 ,  , w_6485 );
buf ( w_6483 , \2097_b1 );
not ( w_6483 , w_6486 );
not (  , w_6487 );
and ( w_6486 , w_6487 , \2097_b0 );
buf ( \2099_b1 , \1840_b1 );
not ( \2099_b1 , w_6488 );
not ( \2099_b0 , w_6489 );
and ( w_6488 , w_6489 , \1840_b0 );
buf ( \2100_b1 , \1756_b1 );
not ( \2100_b1 , w_6490 );
not ( \2100_b0 , w_6491 );
and ( w_6490 , w_6491 , \1756_b0 );
or ( \2101_b1 , \2099_b1 , w_6492 );
or ( \2101_b0 , \2099_b0 , \2100_b0 );
not ( \2100_b0 , w_6493 );
and ( w_6493 , w_6492 , \2100_b1 );
or ( \2102_b1 , \c[1]_b1 , \b[12]_b1 );
xor ( \2102_b0 , \c[1]_b0 , w_6494 );
not ( w_6494 , w_6495 );
and ( w_6495 , \b[12]_b1 , \b[12]_b0 );
or ( \2103_b1 , \2102_b1 , w_6497 );
not ( w_6497 , w_6498 );
and ( \2103_b0 , \2102_b0 , w_6499 );
and ( w_6498 ,  , w_6499 );
buf ( w_6497 , \c[0]_b1 );
not ( w_6497 , w_6500 );
not (  , w_6501 );
and ( w_6500 , w_6501 , \c[0]_b0 );
or ( \2104_b1 , \2101_b1 , w_6503 );
not ( w_6503 , w_6504 );
and ( \2104_b0 , \2101_b0 , w_6505 );
and ( w_6504 ,  , w_6505 );
buf ( w_6503 , \2103_b1 );
not ( w_6503 , w_6506 );
not (  , w_6507 );
and ( w_6506 , w_6507 , \2103_b0 );
or ( \2105_b1 , \2098_b1 , \2104_b1 );
xor ( \2105_b0 , \2098_b0 , w_6508 );
not ( w_6508 , w_6509 );
and ( w_6509 , \2104_b1 , \2104_b0 );
buf ( \2106_b1 , \1690_b1 );
not ( \2106_b1 , w_6510 );
not ( \2106_b0 , w_6511 );
and ( w_6510 , w_6511 , \1690_b0 );
or ( \2107_b1 , \1689_b1 , w_6513 );
not ( w_6513 , w_6514 );
and ( \2107_b0 , \1689_b0 , w_6515 );
and ( w_6514 ,  , w_6515 );
buf ( w_6513 , \1684_b1 );
not ( w_6513 , w_6516 );
not (  , w_6517 );
and ( w_6516 , w_6517 , \1684_b0 );
buf ( \2108_b1 , \2107_b1 );
not ( \2108_b1 , w_6518 );
not ( \2108_b0 , w_6519 );
and ( w_6518 , w_6519 , \2107_b0 );
or ( \2109_b1 , \2106_b1 , w_6520 );
or ( \2109_b0 , \2106_b0 , \2108_b0 );
not ( \2108_b0 , w_6521 );
and ( w_6521 , w_6520 , \2108_b1 );
or ( \2110_b1 , \b[2]_b1 , \c[11]_b1 );
xor ( \2110_b0 , \b[2]_b0 , w_6522 );
not ( w_6522 , w_6523 );
and ( w_6523 , \c[11]_b1 , \c[11]_b0 );
or ( \2111_b1 , \1689_b1 , w_6525 );
not ( w_6525 , w_6526 );
and ( \2111_b0 , \1689_b0 , w_6527 );
and ( w_6526 ,  , w_6527 );
buf ( w_6525 , \2110_b1 );
not ( w_6525 , w_6528 );
not (  , w_6529 );
and ( w_6528 , w_6529 , \2110_b0 );
or ( \2112_b1 , \2109_b1 , w_6531 );
not ( w_6531 , w_6532 );
and ( \2112_b0 , \2109_b0 , w_6533 );
and ( w_6532 ,  , w_6533 );
buf ( w_6531 , \2111_b1 );
not ( w_6531 , w_6534 );
not (  , w_6535 );
and ( w_6534 , w_6535 , \2111_b0 );
or ( \2113_b1 , \2105_b1 , \2112_b1 );
xor ( \2113_b0 , \2105_b0 , w_6536 );
not ( w_6536 , w_6537 );
and ( w_6537 , \2112_b1 , \2112_b0 );
or ( \2114_b1 , \2090_b1 , \2113_b1 );
xor ( \2114_b0 , \2090_b0 , w_6538 );
not ( w_6538 , w_6539 );
and ( w_6539 , \2113_b1 , \2113_b0 );
buf ( \2115_b1 , \1681_b1 );
not ( \2115_b1 , w_6540 );
not ( \2115_b0 , w_6541 );
and ( w_6540 , w_6541 , \1681_b0 );
or ( \2116_b1 , \2115_b1 , w_6543 );
not ( w_6543 , w_6544 );
and ( \2116_b0 , \2115_b0 , w_6545 );
and ( w_6544 ,  , w_6545 );
buf ( w_6543 , \1693_b1 );
not ( w_6543 , w_6546 );
not (  , w_6547 );
and ( w_6546 , w_6547 , \1693_b0 );
buf ( \2117_b1 , \2116_b1 );
not ( \2117_b1 , w_6548 );
not ( \2117_b0 , w_6549 );
and ( w_6548 , w_6549 , \2116_b0 );
buf ( \2118_b1 , \1712_b1 );
not ( \2118_b1 , w_6550 );
not ( \2118_b0 , w_6551 );
and ( w_6550 , w_6551 , \1712_b0 );
or ( \2119_b1 , \2117_b1 , w_6552 );
or ( \2119_b0 , \2117_b0 , \2118_b0 );
not ( \2118_b0 , w_6553 );
and ( w_6553 , w_6552 , \2118_b1 );
or ( \2120_b1 , \1681_b1 , w_6555 );
not ( w_6555 , w_6556 );
and ( \2120_b0 , \1681_b0 , w_6557 );
and ( w_6556 ,  , w_6557 );
buf ( w_6555 , \1692_b1 );
not ( w_6555 , w_6558 );
not (  , w_6559 );
and ( w_6558 , w_6559 , \1692_b0 );
or ( \2121_b1 , \2119_b1 , w_6561 );
not ( w_6561 , w_6562 );
and ( \2121_b0 , \2119_b0 , w_6563 );
and ( w_6562 ,  , w_6563 );
buf ( w_6561 , \2120_b1 );
not ( w_6561 , w_6564 );
not (  , w_6565 );
and ( w_6564 , w_6565 , \2120_b0 );
or ( \2122_b1 , \2114_b1 , \2121_b1 );
xor ( \2122_b0 , \2114_b0 , w_6566 );
not ( w_6566 , w_6567 );
and ( w_6567 , \2121_b1 , \2121_b0 );
or ( \2123_b1 , \2074_b1 , \2122_b1 );
xor ( \2123_b0 , \2074_b0 , w_6568 );
not ( w_6568 , w_6569 );
and ( w_6569 , \2122_b1 , \2122_b0 );
or ( \2124_b1 , \1794_b1 , w_6571 );
not ( w_6571 , w_6572 );
and ( \2124_b0 , \1794_b0 , w_6573 );
and ( w_6572 ,  , w_6573 );
buf ( w_6571 , \1713_b1 );
not ( w_6571 , w_6574 );
not (  , w_6575 );
and ( w_6574 , w_6575 , \1713_b0 );
or ( \2125_b1 , \2124_b1 , w_6576 );
or ( \2125_b0 , \2124_b0 , \1865_b0 );
not ( \1865_b0 , w_6577 );
and ( w_6577 , w_6576 , \1865_b1 );
or ( \2126_b1 , \1794_b1 , w_6579 );
not ( w_6579 , w_6580 );
and ( \2126_b0 , \1794_b0 , w_6581 );
and ( w_6580 ,  , w_6581 );
buf ( w_6579 , \1713_b1 );
not ( w_6579 , w_6582 );
not (  , w_6583 );
and ( w_6582 , w_6583 , \1713_b0 );
or ( \2127_b1 , \2125_b1 , w_6585 );
not ( w_6585 , w_6586 );
and ( \2127_b0 , \2125_b0 , w_6587 );
and ( w_6586 ,  , w_6587 );
buf ( w_6585 , \2126_b1 );
not ( w_6585 , w_6588 );
not (  , w_6589 );
and ( w_6588 , w_6589 , \2126_b0 );
or ( \2128_b1 , \2123_b1 , w_6591 );
not ( w_6591 , w_6592 );
and ( \2128_b0 , \2123_b0 , w_6593 );
and ( w_6592 ,  , w_6593 );
buf ( w_6591 , \2127_b1 );
not ( w_6591 , w_6594 );
not (  , w_6595 );
and ( w_6594 , w_6595 , \2127_b0 );
buf ( \2129_b1 , \2128_b1 );
not ( \2129_b1 , w_6596 );
not ( \2129_b0 , w_6597 );
and ( w_6596 , w_6597 , \2128_b0 );
or ( \2130_b1 , \2001_b1 , \2020_b1 );
xor ( \2130_b0 , \2001_b0 , w_6598 );
not ( w_6598 , w_6599 );
and ( w_6599 , \2020_b1 , \2020_b0 );
or ( \2131_b1 , \2130_b1 , \2023_b1 );
xor ( \2131_b0 , \2130_b0 , w_6600 );
not ( w_6600 , w_6601 );
and ( w_6601 , \2023_b1 , \2023_b0 );
or ( \2132_b1 , \2015_b1 , \2013_b1 );
xor ( \2132_b0 , \2015_b0 , w_6602 );
not ( w_6602 , w_6603 );
and ( w_6603 , \2013_b1 , \2013_b0 );
or ( \2133_b1 , \2132_b1 , w_6604 );
xor ( \2133_b0 , \2132_b0 , w_6606 );
not ( w_6606 , w_6607 );
and ( w_6607 , w_6604 , w_6605 );
buf ( w_6604 , \2007_b1 );
not ( w_6604 , w_6608 );
not ( w_6605 , w_6609 );
and ( w_6608 , w_6609 , \2007_b0 );
or ( \2134_b1 , \b[0]_b1 , w_6611 );
not ( w_6611 , w_6612 );
and ( \2134_b0 , \b[0]_b0 , w_6613 );
and ( w_6612 ,  , w_6613 );
buf ( w_6611 , \c[4]_b1 );
not ( w_6611 , w_6614 );
not (  , w_6615 );
and ( w_6614 , w_6615 , \c[4]_b0 );
or ( \2135_b1 , \b[0]_b1 , w_6616 );
or ( \2135_b0 , \b[0]_b0 , \c[4]_b0 );
not ( \c[4]_b0 , w_6617 );
and ( w_6617 , w_6616 , \c[4]_b1 );
or ( \2136_b1 , \2135_b1 , w_6619 );
not ( w_6619 , w_6620 );
and ( \2136_b0 , \2135_b0 , w_6621 );
and ( w_6620 ,  , w_6621 );
buf ( w_6619 , \c[3]_b1 );
not ( w_6619 , w_6622 );
not (  , w_6623 );
and ( w_6622 , w_6623 , \c[3]_b0 );
buf ( \2138_b1 , \2137_b1 );
not ( \2138_b1 , w_6624 );
not ( \2138_b0 , w_6625 );
and ( w_6624 , w_6625 , \2137_b0 );
or ( \2139_b1 , \b[4]_b1 , \c[1]_b1 );
xor ( \2139_b0 , \b[4]_b0 , w_6626 );
not ( w_6626 , w_6627 );
and ( w_6627 , \c[1]_b1 , \c[1]_b0 );
buf ( \2140_b1 , \2139_b1 );
not ( \2140_b1 , w_6628 );
not ( \2140_b0 , w_6629 );
and ( w_6628 , w_6629 , \2139_b0 );
buf ( \2141_b1 , \1756_b1 );
not ( \2141_b1 , w_6630 );
not ( \2141_b0 , w_6631 );
and ( w_6630 , w_6631 , \1756_b0 );
or ( \2142_b1 , \2140_b1 , w_6632 );
or ( \2142_b0 , \2140_b0 , \2141_b0 );
not ( \2141_b0 , w_6633 );
and ( w_6633 , w_6632 , \2141_b1 );
or ( \2143_b1 , \2008_b1 , w_6635 );
not ( w_6635 , w_6636 );
and ( \2143_b0 , \2008_b0 , w_6637 );
and ( w_6636 ,  , w_6637 );
buf ( w_6635 , \c[0]_b1 );
not ( w_6635 , w_6638 );
not (  , w_6639 );
and ( w_6638 , w_6639 , \c[0]_b0 );
or ( \2144_b1 , \2142_b1 , w_6641 );
not ( w_6641 , w_6642 );
and ( \2144_b0 , \2142_b0 , w_6643 );
and ( w_6642 ,  , w_6643 );
buf ( w_6641 , \2143_b1 );
not ( w_6641 , w_6644 );
not (  , w_6645 );
and ( w_6644 , w_6645 , \2143_b0 );
or ( \2145_b1 , \2138_b1 , w_6647 );
not ( w_6647 , w_6648 );
and ( \2145_b0 , \2138_b0 , w_6649 );
and ( w_6648 ,  , w_6649 );
buf ( w_6647 , \2144_b1 );
not ( w_6647 , w_6650 );
not (  , w_6651 );
and ( w_6650 , w_6651 , \2144_b0 );
or ( \2146_b1 , \b[1]_b1 , \c[5]_b1 );
xor ( \2146_b0 , \b[1]_b0 , w_6652 );
not ( w_6652 , w_6653 );
and ( w_6653 , \c[5]_b1 , \c[5]_b0 );
buf ( \2147_b1 , \2146_b1 );
not ( \2147_b1 , w_6654 );
not ( \2147_b0 , w_6655 );
and ( w_6654 , w_6655 , \2146_b0 );
buf ( \2148_b1 , \1926_b1 );
not ( \2148_b1 , w_6656 );
not ( \2148_b0 , w_6657 );
and ( w_6656 , w_6657 , \1926_b0 );
or ( \2149_b1 , \2147_b1 , w_6658 );
or ( \2149_b0 , \2147_b0 , \2148_b0 );
not ( \2148_b0 , w_6659 );
and ( w_6659 , w_6658 , \2148_b1 );
or ( \2150_b1 , \1678_b1 , w_6661 );
not ( w_6661 , w_6662 );
and ( \2150_b0 , \1678_b0 , w_6663 );
and ( w_6662 ,  , w_6663 );
buf ( w_6661 , \1965_b1 );
not ( w_6661 , w_6664 );
not (  , w_6665 );
and ( w_6664 , w_6665 , \1965_b0 );
or ( \2151_b1 , \2149_b1 , w_6667 );
not ( w_6667 , w_6668 );
and ( \2151_b0 , \2149_b0 , w_6669 );
and ( w_6668 ,  , w_6669 );
buf ( w_6667 , \2150_b1 );
not ( w_6667 , w_6670 );
not (  , w_6671 );
and ( w_6670 , w_6671 , \2150_b0 );
buf ( \2152_b1 , \2151_b1 );
not ( \2152_b1 , w_6672 );
not ( \2152_b0 , w_6673 );
and ( w_6672 , w_6673 , \2151_b0 );
or ( \2153_b1 , \2145_b1 , w_6675 );
not ( w_6675 , w_6676 );
and ( \2153_b0 , \2145_b0 , w_6677 );
and ( w_6676 ,  , w_6677 );
buf ( w_6675 , \2152_b1 );
not ( w_6675 , w_6678 );
not (  , w_6679 );
and ( w_6678 , w_6679 , \2152_b0 );
or ( \2154_b1 , \2133_b1 , \2153_b1 );
not ( \2153_b1 , w_6680 );
and ( \2154_b0 , \2133_b0 , w_6681 );
and ( w_6680 , w_6681 , \2153_b0 );
buf ( \2155_b1 , \2145_b1 );
not ( \2155_b1 , w_6682 );
not ( \2155_b0 , w_6683 );
and ( w_6682 , w_6683 , \2145_b0 );
or ( \2156_b1 , \2155_b1 , \2151_b1 );
not ( \2151_b1 , w_6684 );
and ( \2156_b0 , \2155_b0 , w_6685 );
and ( w_6684 , w_6685 , \2151_b0 );
or ( \2157_b1 , \2154_b1 , w_6687 );
not ( w_6687 , w_6688 );
and ( \2157_b0 , \2154_b0 , w_6689 );
and ( w_6688 ,  , w_6689 );
buf ( w_6687 , \2156_b1 );
not ( w_6687 , w_6690 );
not (  , w_6691 );
and ( w_6690 , w_6691 , \2156_b0 );
or ( \2158_b1 , \2131_b1 , w_6693 );
not ( w_6693 , w_6694 );
and ( \2158_b0 , \2131_b0 , w_6695 );
and ( w_6694 ,  , w_6695 );
buf ( w_6693 , \2157_b1 );
not ( w_6693 , w_6696 );
not (  , w_6697 );
and ( w_6696 , w_6697 , \2157_b0 );
buf ( \2159_b1 , \2158_b1 );
not ( \2159_b1 , w_6698 );
not ( \2159_b0 , w_6699 );
and ( w_6698 , w_6699 , \2158_b0 );
buf ( \2160_b1 , \2146_b1 );
not ( \2160_b1 , w_6700 );
not ( \2160_b0 , w_6701 );
and ( w_6700 , w_6701 , \2146_b0 );
buf ( \2161_b1 , \1674_b1 );
not ( \2161_b1 , w_6702 );
not ( \2161_b0 , w_6703 );
and ( w_6702 , w_6703 , \1674_b0 );
or ( \2162_b1 , \2160_b1 , w_6704 );
or ( \2162_b0 , \2160_b0 , \2161_b0 );
not ( \2161_b0 , w_6705 );
and ( w_6705 , w_6704 , \2161_b1 );
or ( \2163_b1 , \b[0]_b1 , \c[5]_b1 );
xor ( \2163_b0 , \b[0]_b0 , w_6706 );
not ( w_6706 , w_6707 );
and ( w_6707 , \c[5]_b1 , \c[5]_b0 );
or ( \2164_b1 , \1672_b1 , w_6709 );
not ( w_6709 , w_6710 );
and ( \2164_b0 , \1672_b0 , w_6711 );
and ( w_6710 ,  , w_6711 );
buf ( w_6709 , \2163_b1 );
not ( w_6709 , w_6712 );
not (  , w_6713 );
and ( w_6712 , w_6713 , \2163_b0 );
or ( \2165_b1 , \2164_b1 , w_6714 );
or ( \2165_b0 , \2164_b0 , \1674_b0 );
not ( \1674_b0 , w_6715 );
and ( w_6715 , w_6714 , \1674_b1 );
or ( \2166_b1 , \2162_b1 , w_6717 );
not ( w_6717 , w_6718 );
and ( \2166_b0 , \2162_b0 , w_6719 );
and ( w_6718 ,  , w_6719 );
buf ( w_6717 , \2165_b1 );
not ( w_6717 , w_6720 );
not (  , w_6721 );
and ( w_6720 , w_6721 , \2165_b0 );
or ( \2167_b1 , \b[2]_b1 , \c[3]_b1 );
xor ( \2167_b0 , \b[2]_b0 , w_6722 );
not ( w_6722 , w_6723 );
and ( w_6723 , \c[3]_b1 , \c[3]_b0 );
buf ( \2168_b1 , \2167_b1 );
not ( \2168_b1 , w_6724 );
not ( \2168_b0 , w_6725 );
and ( w_6724 , w_6725 , \2167_b0 );
buf ( \2169_b1 , \1722_b1 );
not ( \2169_b1 , w_6726 );
not ( \2169_b0 , w_6727 );
and ( w_6726 , w_6727 , \1722_b0 );
or ( \2170_b1 , \2168_b1 , w_6728 );
or ( \2170_b0 , \2168_b0 , \2169_b0 );
not ( \2169_b0 , w_6729 );
and ( w_6729 , w_6728 , \2169_b1 );
or ( \2171_b1 , \1725_b1 , w_6731 );
not ( w_6731 , w_6732 );
and ( \2171_b0 , \1725_b0 , w_6733 );
and ( w_6732 ,  , w_6733 );
buf ( w_6731 , \2002_b1 );
not ( w_6731 , w_6734 );
not (  , w_6735 );
and ( w_6734 , w_6735 , \2002_b0 );
or ( \2172_b1 , \2170_b1 , w_6737 );
not ( w_6737 , w_6738 );
and ( \2172_b0 , \2170_b0 , w_6739 );
and ( w_6738 ,  , w_6739 );
buf ( w_6737 , \2171_b1 );
not ( w_6737 , w_6740 );
not (  , w_6741 );
and ( w_6740 , w_6741 , \2171_b0 );
or ( \2173_b1 , \2166_b1 , \2172_b1 );
xor ( \2173_b0 , \2166_b0 , w_6742 );
not ( w_6742 , w_6743 );
and ( w_6743 , \2172_b1 , \2172_b0 );
buf ( \2174_b1 , \2144_b1 );
not ( \2174_b1 , w_6744 );
not ( \2174_b0 , w_6745 );
and ( w_6744 , w_6745 , \2144_b0 );
or ( \2175_b1 , \2137_b1 , \2174_b1 );
xor ( \2175_b0 , \2137_b0 , w_6746 );
not ( w_6746 , w_6747 );
and ( w_6747 , \2174_b1 , \2174_b0 );
or ( \2176_b1 , \2173_b1 , \2175_b1 );
not ( \2175_b1 , w_6748 );
and ( \2176_b0 , \2173_b0 , w_6749 );
and ( w_6748 , w_6749 , \2175_b0 );
or ( \2177_b1 , \2166_b1 , \2172_b1 );
not ( \2172_b1 , w_6750 );
and ( \2177_b0 , \2166_b0 , w_6751 );
and ( w_6750 , w_6751 , \2172_b0 );
or ( \2178_b1 , \2176_b1 , w_6752 );
or ( \2178_b0 , \2176_b0 , \2177_b0 );
not ( \2177_b0 , w_6753 );
and ( w_6753 , w_6752 , \2177_b1 );
or ( \2179_b1 , \2155_b1 , \2152_b1 );
xor ( \2179_b0 , \2155_b0 , w_6754 );
not ( w_6754 , w_6755 );
and ( w_6755 , \2152_b1 , \2152_b0 );
or ( \2180_b1 , \2179_b1 , w_6756 );
xor ( \2180_b0 , \2179_b0 , w_6758 );
not ( w_6758 , w_6759 );
and ( w_6759 , w_6756 , w_6757 );
buf ( w_6756 , \2133_b1 );
not ( w_6756 , w_6760 );
not ( w_6757 , w_6761 );
and ( w_6760 , w_6761 , \2133_b0 );
or ( \2181_b1 , \2178_b1 , \2180_b1 );
xor ( \2181_b0 , \2178_b0 , w_6762 );
not ( w_6762 , w_6763 );
and ( w_6763 , \2180_b1 , \2180_b0 );
or ( \2182_b1 , \c[1]_b1 , \b[2]_b1 );
xor ( \2182_b0 , \c[1]_b0 , w_6764 );
not ( w_6764 , w_6765 );
and ( w_6765 , \b[2]_b1 , \b[2]_b0 );
or ( \2183_b1 , \1756_b1 , \2182_b1 );
not ( \2182_b1 , w_6766 );
and ( \2183_b0 , \1756_b0 , w_6767 );
and ( w_6766 , w_6767 , \2182_b0 );
or ( \2184_b1 , \c[1]_b1 , \b[3]_b1 );
xor ( \2184_b0 , \c[1]_b0 , w_6768 );
not ( w_6768 , w_6769 );
and ( w_6769 , \b[3]_b1 , \b[3]_b0 );
or ( \2185_b1 , \2184_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_6770 );
and ( \2185_b0 , \2184_b0 , w_6771 );
and ( w_6770 , w_6771 , \c[0]_b0 );
or ( \2186_b1 , \2183_b1 , w_6773 );
not ( w_6773 , w_6774 );
and ( \2186_b0 , \2183_b0 , w_6775 );
and ( w_6774 ,  , w_6775 );
buf ( w_6773 , \2185_b1 );
not ( w_6773 , w_6776 );
not (  , w_6777 );
and ( w_6776 , w_6777 , \2185_b0 );
or ( \2187_b1 , \b[0]_b1 , w_6778 );
or ( \2187_b0 , \b[0]_b0 , \c[2]_b0 );
not ( \c[2]_b0 , w_6779 );
and ( w_6779 , w_6778 , \c[2]_b1 );
or ( \2188_b1 , \2187_b1 , w_6781 );
not ( w_6781 , w_6782 );
and ( \2188_b0 , \2187_b0 , w_6783 );
and ( w_6782 ,  , w_6783 );
buf ( w_6781 , \c[1]_b1 );
not ( w_6781 , w_6784 );
not (  , w_6785 );
and ( w_6784 , w_6785 , \c[1]_b0 );
or ( \2189_b1 , \b[0]_b1 , w_6787 );
not ( w_6787 , w_6788 );
and ( \2189_b0 , \b[0]_b0 , w_6789 );
and ( w_6788 ,  , w_6789 );
buf ( w_6787 , \c[2]_b1 );
not ( w_6787 , w_6790 );
not (  , w_6791 );
and ( w_6790 , w_6791 , \c[2]_b0 );
buf ( \2191_b1 , \2190_b1 );
not ( \2191_b1 , w_6792 );
not ( \2191_b0 , w_6793 );
and ( w_6792 , w_6793 , \2190_b0 );
or ( \2192_b1 , \2186_b1 , \2191_b1 );
not ( \2191_b1 , w_6794 );
and ( \2192_b0 , \2186_b0 , w_6795 );
and ( w_6794 , w_6795 , \2191_b0 );
buf ( \2193_b1 , \2186_b1 );
not ( \2193_b1 , w_6796 );
not ( \2193_b0 , w_6797 );
and ( w_6796 , w_6797 , \2186_b0 );
or ( \2194_b1 , \2193_b1 , \2190_b1 );
not ( \2190_b1 , w_6798 );
and ( \2194_b0 , \2193_b0 , w_6799 );
and ( w_6798 , w_6799 , \2190_b0 );
or ( \2195_b1 , \2192_b1 , w_6801 );
not ( w_6801 , w_6802 );
and ( \2195_b0 , \2192_b0 , w_6803 );
and ( w_6802 ,  , w_6803 );
buf ( w_6801 , \2194_b1 );
not ( w_6801 , w_6804 );
not (  , w_6805 );
and ( w_6804 , w_6805 , \2194_b0 );
buf ( \2196_b1 , \1708_b1 );
not ( \2196_b1 , w_6806 );
not ( \2196_b0 , w_6807 );
and ( w_6806 , w_6807 , \1708_b0 );
or ( \2197_b1 , \b[0]_b1 , \c[3]_b1 );
xor ( \2197_b0 , \b[0]_b0 , w_6808 );
not ( w_6808 , w_6809 );
and ( w_6809 , \c[3]_b1 , \c[3]_b0 );
or ( \2198_b1 , \1702_b1 , w_6811 );
not ( w_6811 , w_6812 );
and ( \2198_b0 , \1702_b0 , w_6813 );
and ( w_6812 ,  , w_6813 );
buf ( w_6811 , \2197_b1 );
not ( w_6811 , w_6814 );
not (  , w_6815 );
and ( w_6814 , w_6815 , \2197_b0 );
buf ( \2199_b1 , \2198_b1 );
not ( \2199_b1 , w_6816 );
not ( \2199_b0 , w_6817 );
and ( w_6816 , w_6817 , \2198_b0 );
or ( \2200_b1 , \2196_b1 , \2199_b1 );
not ( \2199_b1 , w_6818 );
and ( \2200_b0 , \2196_b0 , w_6819 );
and ( w_6818 , w_6819 , \2199_b0 );
or ( \2201_b1 , \b[1]_b1 , \c[3]_b1 );
xor ( \2201_b0 , \b[1]_b0 , w_6820 );
not ( w_6820 , w_6821 );
and ( w_6821 , \c[3]_b1 , \c[3]_b0 );
or ( \2202_b1 , \1708_b1 , \2201_b1 );
not ( \2201_b1 , w_6822 );
and ( \2202_b0 , \1708_b0 , w_6823 );
and ( w_6822 , w_6823 , \2201_b0 );
or ( \2203_b1 , \2200_b1 , w_6825 );
not ( w_6825 , w_6826 );
and ( \2203_b0 , \2200_b0 , w_6827 );
and ( w_6826 ,  , w_6827 );
buf ( w_6825 , \2202_b1 );
not ( w_6825 , w_6828 );
not (  , w_6829 );
and ( w_6828 , w_6829 , \2202_b0 );
or ( \2204_b1 , \2195_b1 , w_6831 );
not ( w_6831 , w_6832 );
and ( \2204_b0 , \2195_b0 , w_6833 );
and ( w_6832 ,  , w_6833 );
buf ( w_6831 , \2203_b1 );
not ( w_6831 , w_6834 );
not (  , w_6835 );
and ( w_6834 , w_6835 , \2203_b0 );
buf ( \2205_b1 , \2204_b1 );
not ( \2205_b1 , w_6836 );
not ( \2205_b0 , w_6837 );
and ( w_6836 , w_6837 , \2204_b0 );
or ( \2206_b1 , \1725_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_6838 );
and ( \2206_b0 , \1725_b0 , w_6839 );
and ( w_6838 , w_6839 , \b[0]_b0 );
or ( \2207_b1 , \c[1]_b1 , \b[1]_b1 );
xor ( \2207_b0 , \c[1]_b0 , w_6840 );
not ( w_6840 , w_6841 );
and ( w_6841 , \b[1]_b1 , \b[1]_b0 );
buf ( \2208_b1 , \2207_b1 );
not ( \2208_b1 , w_6842 );
not ( \2208_b0 , w_6843 );
and ( w_6842 , w_6843 , \2207_b0 );
buf ( \2209_b1 , \1756_b1 );
not ( \2209_b1 , w_6844 );
not ( \2209_b0 , w_6845 );
and ( w_6844 , w_6845 , \1756_b0 );
or ( \2210_b1 , \2208_b1 , w_6846 );
or ( \2210_b0 , \2208_b0 , \2209_b0 );
not ( \2209_b0 , w_6847 );
and ( w_6847 , w_6846 , \2209_b1 );
or ( \2211_b1 , \2182_b1 , w_6849 );
not ( w_6849 , w_6850 );
and ( \2211_b0 , \2182_b0 , w_6851 );
and ( w_6850 ,  , w_6851 );
buf ( w_6849 , \c[0]_b1 );
not ( w_6849 , w_6852 );
not (  , w_6853 );
and ( w_6852 , w_6853 , \c[0]_b0 );
or ( \2212_b1 , \2210_b1 , w_6855 );
not ( w_6855 , w_6856 );
and ( \2212_b0 , \2210_b0 , w_6857 );
and ( w_6856 ,  , w_6857 );
buf ( w_6855 , \2211_b1 );
not ( w_6855 , w_6858 );
not (  , w_6859 );
and ( w_6858 , w_6859 , \2211_b0 );
or ( \2213_b1 , \2206_b1 , w_6861 );
not ( w_6861 , w_6862 );
and ( \2213_b0 , \2206_b0 , w_6863 );
and ( w_6862 ,  , w_6863 );
buf ( w_6861 , \2212_b1 );
not ( w_6861 , w_6864 );
not (  , w_6865 );
and ( w_6864 , w_6865 , \2212_b0 );
or ( \2214_b1 , \b[0]_b1 , \c[1]_b1 );
xor ( \2214_b0 , \b[0]_b0 , w_6866 );
not ( w_6866 , w_6867 );
and ( w_6867 , \c[1]_b1 , \c[1]_b0 );
buf ( \2215_b1 , \2214_b1 );
not ( \2215_b1 , w_6868 );
not ( \2215_b0 , w_6869 );
and ( w_6868 , w_6869 , \2214_b0 );
buf ( \2216_b1 , \1756_b1 );
not ( \2216_b1 , w_6870 );
not ( \2216_b0 , w_6871 );
and ( w_6870 , w_6871 , \1756_b0 );
or ( \2217_b1 , \2215_b1 , w_6872 );
or ( \2217_b0 , \2215_b0 , \2216_b0 );
not ( \2216_b0 , w_6873 );
and ( w_6873 , w_6872 , \2216_b1 );
or ( \2218_b1 , \2207_b1 , w_6875 );
not ( w_6875 , w_6876 );
and ( \2218_b0 , \2207_b0 , w_6877 );
and ( w_6876 ,  , w_6877 );
buf ( w_6875 , \c[0]_b1 );
not ( w_6875 , w_6878 );
not (  , w_6879 );
and ( w_6878 , w_6879 , \c[0]_b0 );
or ( \2219_b1 , \2217_b1 , w_6881 );
not ( w_6881 , w_6882 );
and ( \2219_b0 , \2217_b0 , w_6883 );
and ( w_6882 ,  , w_6883 );
buf ( w_6881 , \2218_b1 );
not ( w_6881 , w_6884 );
not (  , w_6885 );
and ( w_6884 , w_6885 , \2218_b0 );
or ( \2220_b1 , \b[0]_b1 , w_6887 );
not ( w_6887 , w_6888 );
and ( \2220_b0 , \b[0]_b0 , w_6889 );
and ( w_6888 ,  , w_6889 );
buf ( w_6887 , \c[0]_b1 );
not ( w_6887 , w_6890 );
not (  , w_6891 );
and ( w_6890 , w_6891 , \c[0]_b0 );
or ( \2221_b1 , \2220_b1 , \c[1]_b1 );
not ( \c[1]_b1 , w_6892 );
and ( \2221_b0 , \2220_b0 , w_6893 );
and ( w_6892 , w_6893 , \c[1]_b0 );
or ( \2222_b1 , \2219_b1 , w_6895 );
not ( w_6895 , w_6896 );
and ( \2222_b0 , \2219_b0 , w_6897 );
and ( w_6896 ,  , w_6897 );
buf ( w_6895 , \2221_b1 );
not ( w_6895 , w_6898 );
not (  , w_6899 );
and ( w_6898 , w_6899 , \2221_b0 );
or ( \2223_b1 , \2213_b1 , w_6900 );
or ( \2223_b0 , \2213_b0 , \2222_b0 );
not ( \2222_b0 , w_6901 );
and ( w_6901 , w_6900 , \2222_b1 );
or ( \2224_b1 , \2212_b1 , w_6903 );
not ( w_6903 , w_6904 );
and ( \2224_b0 , \2212_b0 , w_6905 );
and ( w_6904 ,  , w_6905 );
buf ( w_6903 , \2206_b1 );
not ( w_6903 , w_6906 );
not (  , w_6907 );
and ( w_6906 , w_6907 , \2206_b0 );
or ( \2225_b1 , \2223_b1 , w_6909 );
not ( w_6909 , w_6910 );
and ( \2225_b0 , \2223_b0 , w_6911 );
and ( w_6910 ,  , w_6911 );
buf ( w_6909 , \2224_b1 );
not ( w_6909 , w_6912 );
not (  , w_6913 );
and ( w_6912 , w_6913 , \2224_b0 );
buf ( \2226_b1 , \2225_b1 );
not ( \2226_b1 , w_6914 );
not ( \2226_b0 , w_6915 );
and ( w_6914 , w_6915 , \2225_b0 );
or ( \2227_b1 , \2205_b1 , w_6916 );
or ( \2227_b0 , \2205_b0 , \2226_b0 );
not ( \2226_b0 , w_6917 );
and ( w_6917 , w_6916 , \2226_b1 );
or ( \2228_b1 , \2195_b1 , w_6918 );
or ( \2228_b0 , \2195_b0 , \2203_b0 );
not ( \2203_b0 , w_6919 );
and ( w_6919 , w_6918 , \2203_b1 );
or ( \2229_b1 , \2227_b1 , w_6921 );
not ( w_6921 , w_6922 );
and ( \2229_b0 , \2227_b0 , w_6923 );
and ( w_6922 ,  , w_6923 );
buf ( w_6921 , \2228_b1 );
not ( w_6921 , w_6924 );
not (  , w_6925 );
and ( w_6924 , w_6925 , \2228_b0 );
or ( \2230_b1 , \1674_b1 , w_6927 );
not ( w_6927 , w_6928 );
and ( \2230_b0 , \1674_b0 , w_6929 );
and ( w_6928 ,  , w_6929 );
buf ( w_6927 , \b[0]_b1 );
not ( w_6927 , w_6930 );
not (  , w_6931 );
and ( w_6930 , w_6931 , \b[0]_b0 );
or ( \2231_b1 , \1702_b1 , w_6933 );
not ( w_6933 , w_6934 );
and ( \2231_b0 , \1702_b0 , w_6935 );
and ( w_6934 ,  , w_6935 );
buf ( w_6933 , \2201_b1 );
not ( w_6933 , w_6936 );
not (  , w_6937 );
and ( w_6936 , w_6937 , \2201_b0 );
or ( \2232_b1 , \2231_b1 , w_6938 );
or ( \2232_b0 , \2231_b0 , \1725_b0 );
not ( \1725_b0 , w_6939 );
and ( w_6939 , w_6938 , \1725_b1 );
or ( \2233_b1 , \2167_b1 , w_6941 );
not ( w_6941 , w_6942 );
and ( \2233_b0 , \2167_b0 , w_6943 );
and ( w_6942 ,  , w_6943 );
buf ( w_6941 , \1703_b1 );
not ( w_6941 , w_6944 );
not (  , w_6945 );
and ( w_6944 , w_6945 , \1703_b0 );
or ( \2234_b1 , \2232_b1 , w_6947 );
not ( w_6947 , w_6948 );
and ( \2234_b0 , \2232_b0 , w_6949 );
and ( w_6948 ,  , w_6949 );
buf ( w_6947 , \2233_b1 );
not ( w_6947 , w_6950 );
not (  , w_6951 );
and ( w_6950 , w_6951 , \2233_b0 );
buf ( \2235_b1 , \2234_b1 );
not ( \2235_b1 , w_6952 );
not ( \2235_b0 , w_6953 );
and ( w_6952 , w_6953 , \2234_b0 );
or ( \2236_b1 , \2230_b1 , \2235_b1 );
xor ( \2236_b0 , \2230_b0 , w_6954 );
not ( w_6954 , w_6955 );
and ( w_6955 , \2235_b1 , \2235_b0 );
buf ( \2237_b1 , \2184_b1 );
not ( \2237_b1 , w_6956 );
not ( \2237_b0 , w_6957 );
and ( w_6956 , w_6957 , \2184_b0 );
buf ( \2238_b1 , \1756_b1 );
not ( \2238_b1 , w_6958 );
not ( \2238_b0 , w_6959 );
and ( w_6958 , w_6959 , \1756_b0 );
or ( \2239_b1 , \2237_b1 , w_6960 );
or ( \2239_b0 , \2237_b0 , \2238_b0 );
not ( \2238_b0 , w_6961 );
and ( w_6961 , w_6960 , \2238_b1 );
or ( \2240_b1 , \2139_b1 , w_6963 );
not ( w_6963 , w_6964 );
and ( \2240_b0 , \2139_b0 , w_6965 );
and ( w_6964 ,  , w_6965 );
buf ( w_6963 , \c[0]_b1 );
not ( w_6963 , w_6966 );
not (  , w_6967 );
and ( w_6966 , w_6967 , \c[0]_b0 );
or ( \2241_b1 , \2239_b1 , w_6969 );
not ( w_6969 , w_6970 );
and ( \2241_b0 , \2239_b0 , w_6971 );
and ( w_6970 ,  , w_6971 );
buf ( w_6969 , \2240_b1 );
not ( w_6969 , w_6972 );
not (  , w_6973 );
and ( w_6972 , w_6973 , \2240_b0 );
or ( \2242_b1 , \2236_b1 , w_6974 );
xor ( \2242_b0 , \2236_b0 , w_6976 );
not ( w_6976 , w_6977 );
and ( w_6977 , w_6974 , w_6975 );
buf ( w_6974 , \2241_b1 );
not ( w_6974 , w_6978 );
not ( w_6975 , w_6979 );
and ( w_6978 , w_6979 , \2241_b0 );
buf ( \2243_b1 , \2186_b1 );
not ( \2243_b1 , w_6980 );
not ( \2243_b0 , w_6981 );
and ( w_6980 , w_6981 , \2186_b0 );
or ( \2244_b1 , \2243_b1 , w_6983 );
not ( w_6983 , w_6984 );
and ( \2244_b0 , \2243_b0 , w_6985 );
and ( w_6984 ,  , w_6985 );
buf ( w_6983 , \2191_b1 );
not ( w_6983 , w_6986 );
not (  , w_6987 );
and ( w_6986 , w_6987 , \2191_b0 );
or ( \2245_b1 , \2242_b1 , w_6989 );
not ( w_6989 , w_6990 );
and ( \2245_b0 , \2242_b0 , w_6991 );
and ( w_6990 ,  , w_6991 );
buf ( w_6989 , \2244_b1 );
not ( w_6989 , w_6992 );
not (  , w_6993 );
and ( w_6992 , w_6993 , \2244_b0 );
or ( \2246_b1 , \2229_b1 , \2245_b1 );
not ( \2245_b1 , w_6994 );
and ( \2246_b0 , \2229_b0 , w_6995 );
and ( w_6994 , w_6995 , \2245_b0 );
or ( \2247_b1 , \2242_b1 , w_6997 );
not ( w_6997 , w_6998 );
and ( \2247_b0 , \2242_b0 , w_6999 );
and ( w_6998 ,  , w_6999 );
buf ( w_6997 , \2244_b1 );
not ( w_6997 , w_7000 );
not (  , w_7001 );
and ( w_7000 , w_7001 , \2244_b0 );
or ( \2248_b1 , \2246_b1 , w_7003 );
not ( w_7003 , w_7004 );
and ( \2248_b0 , \2246_b0 , w_7005 );
and ( w_7004 ,  , w_7005 );
buf ( w_7003 , \2247_b1 );
not ( w_7003 , w_7006 );
not (  , w_7007 );
and ( w_7006 , w_7007 , \2247_b0 );
or ( \2249_b1 , \2166_b1 , \2172_b1 );
xor ( \2249_b0 , \2166_b0 , w_7008 );
not ( w_7008 , w_7009 );
and ( w_7009 , \2172_b1 , \2172_b0 );
or ( \2250_b1 , \2249_b1 , \2175_b1 );
xor ( \2250_b0 , \2249_b0 , w_7010 );
not ( w_7010 , w_7011 );
and ( w_7011 , \2175_b1 , \2175_b0 );
buf ( \2251_b1 , \2235_b1 );
not ( \2251_b1 , w_7012 );
not ( \2251_b0 , w_7013 );
and ( w_7012 , w_7013 , \2235_b0 );
buf ( \2252_b1 , \2241_b1 );
not ( \2252_b1 , w_7014 );
not ( \2252_b0 , w_7015 );
and ( w_7014 , w_7015 , \2241_b0 );
or ( \2253_b1 , \2252_b1 , w_7017 );
not ( w_7017 , w_7018 );
and ( \2253_b0 , \2252_b0 , w_7019 );
and ( w_7018 ,  , w_7019 );
buf ( w_7017 , \2230_b1 );
not ( w_7017 , w_7020 );
not (  , w_7021 );
and ( w_7020 , w_7021 , \2230_b0 );
or ( \2254_b1 , \2251_b1 , w_7023 );
not ( w_7023 , w_7024 );
and ( \2254_b0 , \2251_b0 , w_7025 );
and ( w_7024 ,  , w_7025 );
buf ( w_7023 , \2253_b1 );
not ( w_7023 , w_7026 );
not (  , w_7027 );
and ( w_7026 , w_7027 , \2253_b0 );
buf ( \2255_b1 , \2230_b1 );
not ( \2255_b1 , w_7028 );
not ( \2255_b0 , w_7029 );
and ( w_7028 , w_7029 , \2230_b0 );
or ( \2256_b1 , \2255_b1 , w_7031 );
not ( w_7031 , w_7032 );
and ( \2256_b0 , \2255_b0 , w_7033 );
and ( w_7032 ,  , w_7033 );
buf ( w_7031 , \2241_b1 );
not ( w_7031 , w_7034 );
not (  , w_7035 );
and ( w_7034 , w_7035 , \2241_b0 );
or ( \2257_b1 , \2254_b1 , w_7037 );
not ( w_7037 , w_7038 );
and ( \2257_b0 , \2254_b0 , w_7039 );
and ( w_7038 ,  , w_7039 );
buf ( w_7037 , \2256_b1 );
not ( w_7037 , w_7040 );
not (  , w_7041 );
and ( w_7040 , w_7041 , \2256_b0 );
or ( \2258_b1 , \2250_b1 , w_7043 );
not ( w_7043 , w_7044 );
and ( \2258_b0 , \2250_b0 , w_7045 );
and ( w_7044 ,  , w_7045 );
buf ( w_7043 , \2257_b1 );
not ( w_7043 , w_7046 );
not (  , w_7047 );
and ( w_7046 , w_7047 , \2257_b0 );
or ( \2259_b1 , \2248_b1 , w_7048 );
or ( \2259_b0 , \2248_b0 , \2258_b0 );
not ( \2258_b0 , w_7049 );
and ( w_7049 , w_7048 , \2258_b1 );
or ( \2260_b1 , \2250_b1 , w_7051 );
not ( w_7051 , w_7052 );
and ( \2260_b0 , \2250_b0 , w_7053 );
and ( w_7052 ,  , w_7053 );
buf ( w_7051 , \2257_b1 );
not ( w_7051 , w_7054 );
not (  , w_7055 );
and ( w_7054 , w_7055 , \2257_b0 );
or ( \2261_b1 , \2259_b1 , w_7057 );
not ( w_7057 , w_7058 );
and ( \2261_b0 , \2259_b0 , w_7059 );
and ( w_7058 ,  , w_7059 );
buf ( w_7057 , \2260_b1 );
not ( w_7057 , w_7060 );
not (  , w_7061 );
and ( w_7060 , w_7061 , \2260_b0 );
or ( \2262_b1 , \2181_b1 , \2261_b1 );
not ( \2261_b1 , w_7062 );
and ( \2262_b0 , \2181_b0 , w_7063 );
and ( w_7062 , w_7063 , \2261_b0 );
or ( \2263_b1 , \2178_b1 , \2180_b1 );
not ( \2180_b1 , w_7064 );
and ( \2263_b0 , \2178_b0 , w_7065 );
and ( w_7064 , w_7065 , \2180_b0 );
or ( \2264_b1 , \2262_b1 , w_7066 );
or ( \2264_b0 , \2262_b0 , \2263_b0 );
not ( \2263_b0 , w_7067 );
and ( w_7067 , w_7066 , \2263_b1 );
buf ( \2265_b1 , \2264_b1 );
not ( \2265_b1 , w_7068 );
not ( \2265_b0 , w_7069 );
and ( w_7068 , w_7069 , \2264_b0 );
or ( \2266_b1 , \2159_b1 , w_7070 );
or ( \2266_b0 , \2159_b0 , \2265_b0 );
not ( \2265_b0 , w_7071 );
and ( w_7071 , w_7070 , \2265_b1 );
buf ( \2267_b1 , \2131_b1 );
not ( \2267_b1 , w_7072 );
not ( \2267_b0 , w_7073 );
and ( w_7072 , w_7073 , \2131_b0 );
buf ( \2268_b1 , \2157_b1 );
not ( \2268_b1 , w_7074 );
not ( \2268_b0 , w_7075 );
and ( w_7074 , w_7075 , \2157_b0 );
or ( \2269_b1 , \2267_b1 , w_7077 );
not ( w_7077 , w_7078 );
and ( \2269_b0 , \2267_b0 , w_7079 );
and ( w_7078 ,  , w_7079 );
buf ( w_7077 , \2268_b1 );
not ( w_7077 , w_7080 );
not (  , w_7081 );
and ( w_7080 , w_7081 , \2268_b0 );
or ( \2270_b1 , \2266_b1 , w_7083 );
not ( w_7083 , w_7084 );
and ( \2270_b0 , \2266_b0 , w_7085 );
and ( w_7084 ,  , w_7085 );
buf ( w_7083 , \2269_b1 );
not ( w_7083 , w_7086 );
not (  , w_7087 );
and ( w_7086 , w_7087 , \2269_b0 );
buf ( \2271_b1 , \2270_b1 );
buf ( \2271_b0 , \2270_b0 );
or ( \2273_b1 , \1866_b1 , w_7089 );
not ( w_7089 , w_7090 );
and ( \2273_b0 , \1866_b0 , w_7091 );
and ( w_7090 ,  , w_7091 );
buf ( w_7089 , \1900_b1 );
not ( w_7089 , w_7092 );
not (  , w_7093 );
and ( w_7092 , w_7093 , \1900_b0 );
or ( \2274_b1 , \2129_b1 , w_7095 );
not ( w_7095 , w_7096 );
and ( \2274_b0 , \2129_b0 , w_7097 );
and ( w_7096 ,  , w_7097 );
buf ( w_7095 , \2273_b1 );
not ( w_7095 , w_7098 );
not (  , w_7099 );
and ( w_7098 , w_7099 , \2273_b0 );
buf ( \2275_b1 , \2000_b1 );
not ( \2275_b1 , w_7100 );
not ( \2275_b0 , w_7101 );
and ( w_7100 , w_7101 , \2000_b0 );
buf ( \2276_b1 , \2026_b1 );
not ( \2276_b1 , w_7102 );
not ( \2276_b0 , w_7103 );
and ( w_7102 , w_7103 , \2026_b0 );
or ( \2277_b1 , \2275_b1 , w_7105 );
not ( w_7105 , w_7106 );
and ( \2277_b0 , \2275_b0 , w_7107 );
and ( w_7106 ,  , w_7107 );
buf ( w_7105 , \2276_b1 );
not ( w_7105 , w_7108 );
not (  , w_7109 );
and ( w_7108 , w_7109 , \2276_b0 );
or ( \2278_b1 , \2048_b1 , w_7110 );
or ( \2278_b0 , \2048_b0 , \2277_b0 );
not ( \2277_b0 , w_7111 );
and ( w_7111 , w_7110 , \2277_b1 );
or ( \2279_b1 , \2039_b1 , w_7113 );
not ( w_7113 , w_7114 );
and ( \2279_b0 , \2039_b0 , w_7115 );
and ( w_7114 ,  , w_7115 );
buf ( w_7113 , \2047_b1 );
not ( w_7113 , w_7116 );
not (  , w_7117 );
and ( w_7116 , w_7117 , \2047_b0 );
or ( \2280_b1 , \2278_b1 , w_7119 );
not ( w_7119 , w_7120 );
and ( \2280_b0 , \2278_b0 , w_7121 );
and ( w_7120 ,  , w_7121 );
buf ( w_7119 , \2279_b1 );
not ( w_7119 , w_7122 );
not (  , w_7123 );
and ( w_7122 , w_7123 , \2279_b0 );
or ( \2281_b1 , \1903_b1 , w_7125 );
not ( w_7125 , w_7126 );
and ( \2281_b0 , \1903_b0 , w_7127 );
and ( w_7126 ,  , w_7127 );
buf ( w_7125 , \1953_b1 );
not ( w_7125 , w_7128 );
not (  , w_7129 );
and ( w_7128 , w_7129 , \1953_b0 );
or ( \2282_b1 , \2280_b1 , w_7131 );
not ( w_7131 , w_7132 );
and ( \2282_b0 , \2280_b0 , w_7133 );
and ( w_7132 ,  , w_7133 );
buf ( w_7131 , \2281_b1 );
not ( w_7131 , w_7134 );
not (  , w_7135 );
and ( w_7134 , w_7135 , \2281_b0 );
buf ( \2283_b1 , \2282_b1 );
not ( \2283_b1 , w_7136 );
not ( \2283_b0 , w_7137 );
and ( w_7136 , w_7137 , \2282_b0 );
or ( \2284_b1 , \1866_b1 , w_7139 );
not ( w_7139 , w_7140 );
and ( \2284_b0 , \1866_b0 , w_7141 );
and ( w_7140 ,  , w_7141 );
buf ( w_7139 , \1900_b1 );
not ( w_7139 , w_7142 );
not (  , w_7143 );
and ( w_7142 , w_7143 , \1900_b0 );
buf ( \2285_b1 , \1954_b1 );
buf ( \2285_b0 , \1954_b0 );
or ( \2287_b1 , \2123_b1 , \2127_b1 );
not ( \2127_b1 , w_7144 );
and ( \2287_b0 , \2123_b0 , w_7145 );
and ( w_7144 , w_7145 , \2127_b0 );
buf ( \2288_b1 , \2287_b1 );
not ( \2288_b1 , w_7146 );
not ( \2288_b0 , w_7147 );
and ( w_7146 , w_7147 , \2287_b0 );
buf ( \2290_b1 , \2102_b1 );
not ( \2290_b1 , w_7148 );
not ( \2290_b0 , w_7149 );
and ( w_7148 , w_7149 , \2102_b0 );
buf ( \2291_b1 , \1756_b1 );
not ( \2291_b1 , w_7150 );
not ( \2291_b0 , w_7151 );
and ( w_7150 , w_7151 , \1756_b0 );
or ( \2292_b1 , \2290_b1 , w_7152 );
or ( \2292_b0 , \2290_b0 , \2291_b0 );
not ( \2291_b0 , w_7153 );
and ( w_7153 , w_7152 , \2291_b1 );
or ( \2293_b1 , \b[13]_b1 , \c[1]_b1 );
xor ( \2293_b0 , \b[13]_b0 , w_7154 );
not ( w_7154 , w_7155 );
and ( w_7155 , \c[1]_b1 , \c[1]_b0 );
or ( \2294_b1 , \2293_b1 , w_7157 );
not ( w_7157 , w_7158 );
and ( \2294_b0 , \2293_b0 , w_7159 );
and ( w_7158 ,  , w_7159 );
buf ( w_7157 , \c[0]_b1 );
not ( w_7157 , w_7160 );
not (  , w_7161 );
and ( w_7160 , w_7161 , \c[0]_b0 );
or ( \2295_b1 , \2292_b1 , w_7163 );
not ( w_7163 , w_7164 );
and ( \2295_b0 , \2292_b0 , w_7165 );
and ( w_7164 ,  , w_7165 );
buf ( w_7163 , \2294_b1 );
not ( w_7163 , w_7166 );
not (  , w_7167 );
and ( w_7166 , w_7167 , \2294_b0 );
buf ( \2296_b1 , \2295_b1 );
not ( \2296_b1 , w_7168 );
not ( \2296_b0 , w_7169 );
and ( w_7168 , w_7169 , \2295_b0 );
or ( \2297_b1 , \b[0]_b1 , w_7170 );
or ( \2297_b0 , \b[0]_b0 , \c[12]_b0 );
not ( \c[12]_b0 , w_7171 );
and ( w_7171 , w_7170 , \c[12]_b1 );
or ( \2298_b1 , \2297_b1 , w_7173 );
not ( w_7173 , w_7174 );
and ( \2298_b0 , \2297_b0 , w_7175 );
and ( w_7174 ,  , w_7175 );
buf ( w_7173 , \c[11]_b1 );
not ( w_7173 , w_7176 );
not (  , w_7177 );
and ( w_7176 , w_7177 , \c[11]_b0 );
or ( \2299_b1 , \b[0]_b1 , w_7179 );
not ( w_7179 , w_7180 );
and ( \2299_b0 , \b[0]_b0 , w_7181 );
and ( w_7180 ,  , w_7181 );
buf ( w_7179 , \c[12]_b1 );
not ( w_7179 , w_7182 );
not (  , w_7183 );
and ( w_7182 , w_7183 , \c[12]_b0 );
buf ( \2301_b1 , \2300_b1 );
not ( \2301_b1 , w_7184 );
not ( \2301_b0 , w_7185 );
and ( w_7184 , w_7185 , \2300_b0 );
or ( \2302_b1 , \2296_b1 , \2301_b1 );
not ( \2301_b1 , w_7186 );
and ( \2302_b0 , \2296_b0 , w_7187 );
and ( w_7186 , w_7187 , \2301_b0 );
or ( \2303_b1 , \2295_b1 , \2300_b1 );
not ( \2300_b1 , w_7188 );
and ( \2303_b0 , \2295_b0 , w_7189 );
and ( w_7188 , w_7189 , \2300_b0 );
or ( \2304_b1 , \2302_b1 , w_7191 );
not ( w_7191 , w_7192 );
and ( \2304_b0 , \2302_b0 , w_7193 );
and ( w_7192 ,  , w_7193 );
buf ( w_7191 , \2303_b1 );
not ( w_7191 , w_7194 );
not (  , w_7195 );
and ( w_7194 , w_7195 , \2303_b0 );
or ( \2305_b1 , \2076_b1 , \2082_b1 );
xor ( \2305_b0 , \2076_b0 , w_7196 );
not ( w_7196 , w_7197 );
and ( w_7197 , \2082_b1 , \2082_b0 );
or ( \2306_b1 , \2305_b1 , \2089_b1 );
not ( \2089_b1 , w_7198 );
and ( \2306_b0 , \2305_b0 , w_7199 );
and ( w_7198 , w_7199 , \2089_b0 );
or ( \2307_b1 , \2076_b1 , \2082_b1 );
not ( \2082_b1 , w_7200 );
and ( \2307_b0 , \2076_b0 , w_7201 );
and ( w_7200 , w_7201 , \2082_b0 );
or ( \2308_b1 , \2306_b1 , w_7202 );
or ( \2308_b0 , \2306_b0 , \2307_b0 );
not ( \2307_b0 , w_7203 );
and ( w_7203 , w_7202 , \2307_b1 );
or ( \2309_b1 , \2304_b1 , \2308_b1 );
xor ( \2309_b0 , \2304_b0 , w_7204 );
not ( w_7204 , w_7205 );
and ( w_7205 , \2308_b1 , \2308_b0 );
or ( \2310_b1 , \2098_b1 , w_7206 );
or ( \2310_b0 , \2098_b0 , \2104_b0 );
not ( \2104_b0 , w_7207 );
and ( w_7207 , w_7206 , \2104_b1 );
or ( \2311_b1 , \2310_b1 , \2112_b1 );
not ( \2112_b1 , w_7208 );
and ( \2311_b0 , \2310_b0 , w_7209 );
and ( w_7208 , w_7209 , \2112_b0 );
or ( \2312_b1 , \2098_b1 , \2104_b1 );
not ( \2104_b1 , w_7210 );
and ( \2312_b0 , \2098_b0 , w_7211 );
and ( w_7210 , w_7211 , \2104_b0 );
or ( \2313_b1 , \2311_b1 , w_7213 );
not ( w_7213 , w_7214 );
and ( \2313_b0 , \2311_b0 , w_7215 );
and ( w_7214 ,  , w_7215 );
buf ( w_7213 , \2312_b1 );
not ( w_7213 , w_7216 );
not (  , w_7217 );
and ( w_7216 , w_7217 , \2312_b0 );
buf ( \2314_b1 , \2313_b1 );
not ( \2314_b1 , w_7218 );
not ( \2314_b0 , w_7219 );
and ( w_7218 , w_7219 , \2313_b0 );
or ( \2315_b1 , \2309_b1 , \2314_b1 );
xor ( \2315_b0 , \2309_b0 , w_7220 );
not ( w_7220 , w_7221 );
and ( w_7221 , \2314_b1 , \2314_b0 );
buf ( \2316_b1 , \2315_b1 );
not ( \2316_b1 , w_7222 );
not ( \2316_b0 , w_7223 );
and ( w_7222 , w_7223 , \2315_b0 );
or ( \2317_b1 , \2090_b1 , \2113_b1 );
xor ( \2317_b0 , \2090_b0 , w_7224 );
not ( w_7224 , w_7225 );
and ( w_7225 , \2113_b1 , \2113_b0 );
or ( \2318_b1 , \2317_b1 , \2121_b1 );
not ( \2121_b1 , w_7226 );
and ( \2318_b0 , \2317_b0 , w_7227 );
and ( w_7226 , w_7227 , \2121_b0 );
or ( \2319_b1 , \2090_b1 , \2113_b1 );
not ( \2113_b1 , w_7228 );
and ( \2319_b0 , \2090_b0 , w_7229 );
and ( w_7228 , w_7229 , \2113_b0 );
or ( \2320_b1 , \2318_b1 , w_7230 );
or ( \2320_b0 , \2318_b0 , \2319_b0 );
not ( \2319_b0 , w_7231 );
and ( w_7231 , w_7230 , \2319_b1 );
buf ( \2321_b1 , \2320_b1 );
not ( \2321_b1 , w_7232 );
not ( \2321_b0 , w_7233 );
and ( w_7232 , w_7233 , \2320_b0 );
or ( \2322_b1 , \2316_b1 , w_7234 );
or ( \2322_b0 , \2316_b0 , \2321_b0 );
not ( \2321_b0 , w_7235 );
and ( w_7235 , w_7234 , \2321_b1 );
or ( \2323_b1 , \2320_b1 , w_7236 );
or ( \2323_b0 , \2320_b0 , \2315_b0 );
not ( \2315_b0 , w_7237 );
and ( w_7237 , w_7236 , \2315_b1 );
or ( \2324_b1 , \2322_b1 , w_7239 );
not ( w_7239 , w_7240 );
and ( \2324_b0 , \2322_b0 , w_7241 );
and ( w_7240 ,  , w_7241 );
buf ( w_7239 , \2323_b1 );
not ( w_7239 , w_7242 );
not (  , w_7243 );
and ( w_7242 , w_7243 , \2323_b0 );
buf ( \2325_b1 , \2055_b1 );
not ( \2325_b1 , w_7244 );
not ( \2325_b0 , w_7245 );
and ( w_7244 , w_7245 , \2055_b0 );
buf ( \2326_b1 , \1675_b1 );
not ( \2326_b1 , w_7246 );
not ( \2326_b0 , w_7247 );
and ( w_7246 , w_7247 , \1675_b0 );
or ( \2327_b1 , \2325_b1 , w_7248 );
or ( \2327_b0 , \2325_b0 , \2326_b0 );
not ( \2326_b0 , w_7249 );
and ( w_7249 , w_7248 , \2326_b1 );
or ( \2328_b1 , \b[9]_b1 , \c[5]_b1 );
xor ( \2328_b0 , \b[9]_b0 , w_7250 );
not ( w_7250 , w_7251 );
and ( w_7251 , \c[5]_b1 , \c[5]_b0 );
or ( \2329_b1 , \1678_b1 , w_7253 );
not ( w_7253 , w_7254 );
and ( \2329_b0 , \1678_b0 , w_7255 );
and ( w_7254 ,  , w_7255 );
buf ( w_7253 , \2328_b1 );
not ( w_7253 , w_7256 );
not (  , w_7257 );
and ( w_7256 , w_7257 , \2328_b0 );
or ( \2330_b1 , \2327_b1 , w_7259 );
not ( w_7259 , w_7260 );
and ( \2330_b0 , \2327_b0 , w_7261 );
and ( w_7260 ,  , w_7261 );
buf ( w_7259 , \2329_b1 );
not ( w_7259 , w_7262 );
not (  , w_7263 );
and ( w_7262 , w_7263 , \2329_b0 );
buf ( \2331_b1 , \2110_b1 );
not ( \2331_b1 , w_7264 );
not ( \2331_b0 , w_7265 );
and ( w_7264 , w_7265 , \2110_b0 );
buf ( \2332_b1 , \1686_b1 );
not ( \2332_b1 , w_7266 );
not ( \2332_b0 , w_7267 );
and ( w_7266 , w_7267 , \1686_b0 );
or ( \2333_b1 , \2331_b1 , w_7268 );
or ( \2333_b0 , \2331_b0 , \2332_b0 );
not ( \2332_b0 , w_7269 );
and ( w_7269 , w_7268 , \2332_b1 );
or ( \2334_b1 , \b[3]_b1 , \c[11]_b1 );
xor ( \2334_b0 , \b[3]_b0 , w_7270 );
not ( w_7270 , w_7271 );
and ( w_7271 , \c[11]_b1 , \c[11]_b0 );
or ( \2335_b1 , \1689_b1 , w_7273 );
not ( w_7273 , w_7274 );
and ( \2335_b0 , \1689_b0 , w_7275 );
and ( w_7274 ,  , w_7275 );
buf ( w_7273 , \2334_b1 );
not ( w_7273 , w_7276 );
not (  , w_7277 );
and ( w_7276 , w_7277 , \2334_b0 );
or ( \2336_b1 , \2333_b1 , w_7279 );
not ( w_7279 , w_7280 );
and ( \2336_b0 , \2333_b0 , w_7281 );
and ( w_7280 ,  , w_7281 );
buf ( w_7279 , \2335_b1 );
not ( w_7279 , w_7282 );
not (  , w_7283 );
and ( w_7282 , w_7283 , \2335_b0 );
or ( \2337_b1 , \2330_b1 , \2336_b1 );
xor ( \2337_b0 , \2330_b0 , w_7284 );
not ( w_7284 , w_7285 );
and ( w_7285 , \2336_b1 , \2336_b0 );
or ( \2338_b1 , \b[0]_b1 , \c[13]_b1 );
xor ( \2338_b0 , \b[0]_b0 , w_7286 );
not ( w_7286 , w_7287 );
and ( w_7287 , \c[13]_b1 , \c[13]_b0 );
buf ( \2339_b1 , \2338_b1 );
not ( \2339_b1 , w_7288 );
not ( \2339_b0 , w_7289 );
and ( w_7288 , w_7289 , \2338_b0 );
or ( \2340_b1 , \c[13]_b1 , w_7290 );
xor ( \2340_b0 , \c[13]_b0 , w_7292 );
not ( w_7292 , w_7293 );
and ( w_7293 , w_7290 , w_7291 );
buf ( w_7290 , \c[12]_b1 );
not ( w_7290 , w_7294 );
not ( w_7291 , w_7295 );
and ( w_7294 , w_7295 , \c[12]_b0 );
or ( \2341_b1 , \2340_b1 , w_7297 );
not ( w_7297 , w_7298 );
and ( \2341_b0 , \2340_b0 , w_7299 );
and ( w_7298 ,  , w_7299 );
buf ( w_7297 , \2075_b1 );
not ( w_7297 , w_7300 );
not (  , w_7301 );
and ( w_7300 , w_7301 , \2075_b0 );
buf ( \2342_b1 , \2341_b1 );
not ( \2342_b1 , w_7302 );
not ( \2342_b0 , w_7303 );
and ( w_7302 , w_7303 , \2341_b0 );
or ( \2343_b1 , \2339_b1 , w_7304 );
or ( \2343_b0 , \2339_b0 , \2342_b0 );
not ( \2342_b0 , w_7305 );
and ( w_7305 , w_7304 , \2342_b1 );
or ( \2344_b1 , \b[1]_b1 , \c[13]_b1 );
xor ( \2344_b0 , \b[1]_b0 , w_7306 );
not ( w_7306 , w_7307 );
and ( w_7307 , \c[13]_b1 , \c[13]_b0 );
or ( \2345_b1 , \2075_b1 , w_7309 );
not ( w_7309 , w_7310 );
and ( \2345_b0 , \2075_b0 , w_7311 );
and ( w_7310 ,  , w_7311 );
buf ( w_7309 , \2344_b1 );
not ( w_7309 , w_7312 );
not (  , w_7313 );
and ( w_7312 , w_7313 , \2344_b0 );
or ( \2346_b1 , \2343_b1 , w_7315 );
not ( w_7315 , w_7316 );
and ( \2346_b0 , \2343_b0 , w_7317 );
and ( w_7316 ,  , w_7317 );
buf ( w_7315 , \2345_b1 );
not ( w_7315 , w_7318 );
not (  , w_7319 );
and ( w_7318 , w_7319 , \2345_b0 );
or ( \2347_b1 , \2337_b1 , \2346_b1 );
xor ( \2347_b0 , \2337_b0 , w_7320 );
not ( w_7320 , w_7321 );
and ( w_7321 , \2346_b1 , \2346_b0 );
buf ( \2348_b1 , \2347_b1 );
not ( \2348_b1 , w_7322 );
not ( \2348_b0 , w_7323 );
and ( w_7322 , w_7323 , \2347_b0 );
buf ( \2349_b1 , \2348_b1 );
not ( \2349_b1 , w_7324 );
not ( \2349_b0 , w_7325 );
and ( w_7324 , w_7325 , \2348_b0 );
buf ( \2350_b1 , \1852_b1 );
not ( \2350_b1 , w_7326 );
not ( \2350_b0 , w_7327 );
and ( w_7326 , w_7327 , \1852_b0 );
buf ( \2351_b1 , \2095_b1 );
not ( \2351_b1 , w_7328 );
not ( \2351_b0 , w_7329 );
and ( w_7328 , w_7329 , \2095_b0 );
or ( \2352_b1 , \2350_b1 , \2351_b1 );
not ( \2351_b1 , w_7330 );
and ( \2352_b0 , \2350_b0 , w_7331 );
and ( w_7330 , w_7331 , \2351_b0 );
or ( \2353_b1 , \b[5]_b1 , \c[9]_b1 );
xor ( \2353_b0 , \b[5]_b0 , w_7332 );
not ( w_7332 , w_7333 );
and ( w_7333 , \c[9]_b1 , \c[9]_b0 );
or ( \2354_b1 , \1802_b1 , \2353_b1 );
not ( \2353_b1 , w_7334 );
and ( \2354_b0 , \1802_b0 , w_7335 );
and ( w_7334 , w_7335 , \2353_b0 );
or ( \2355_b1 , \2352_b1 , w_7337 );
not ( w_7337 , w_7338 );
and ( \2355_b0 , \2352_b0 , w_7339 );
and ( w_7338 ,  , w_7339 );
buf ( w_7337 , \2354_b1 );
not ( w_7337 , w_7340 );
not (  , w_7341 );
and ( w_7340 , w_7341 , \2354_b0 );
buf ( \2356_b1 , \2355_b1 );
not ( \2356_b1 , w_7342 );
not ( \2356_b0 , w_7343 );
and ( w_7342 , w_7343 , \2355_b0 );
buf ( \2357_b1 , \2356_b1 );
not ( \2357_b1 , w_7344 );
not ( \2357_b0 , w_7345 );
and ( w_7344 , w_7345 , \2356_b0 );
buf ( \2358_b1 , \2080_b1 );
not ( \2358_b1 , w_7346 );
not ( \2358_b0 , w_7347 );
and ( w_7346 , w_7347 , \2080_b0 );
buf ( \2359_b1 , \1743_b1 );
not ( \2359_b1 , w_7348 );
not ( \2359_b0 , w_7349 );
and ( w_7348 , w_7349 , \1743_b0 );
or ( \2360_b1 , \2358_b1 , w_7350 );
or ( \2360_b0 , \2358_b0 , \2359_b0 );
not ( \2359_b0 , w_7351 );
and ( w_7351 , w_7350 , \2359_b1 );
or ( \2361_b1 , \b[7]_b1 , \c[7]_b1 );
xor ( \2361_b0 , \b[7]_b0 , w_7352 );
not ( w_7352 , w_7353 );
and ( w_7353 , \c[7]_b1 , \c[7]_b0 );
or ( \2362_b1 , \1747_b1 , w_7355 );
not ( w_7355 , w_7356 );
and ( \2362_b0 , \1747_b0 , w_7357 );
and ( w_7356 ,  , w_7357 );
buf ( w_7355 , \2361_b1 );
not ( w_7355 , w_7358 );
not (  , w_7359 );
and ( w_7358 , w_7359 , \2361_b0 );
or ( \2363_b1 , \2360_b1 , w_7361 );
not ( w_7361 , w_7362 );
and ( \2363_b0 , \2360_b0 , w_7363 );
and ( w_7362 ,  , w_7363 );
buf ( w_7361 , \2362_b1 );
not ( w_7361 , w_7364 );
not (  , w_7365 );
and ( w_7364 , w_7365 , \2362_b0 );
buf ( \2364_b1 , \2363_b1 );
not ( \2364_b1 , w_7366 );
not ( \2364_b0 , w_7367 );
and ( w_7366 , w_7367 , \2363_b0 );
buf ( \2365_b1 , \2364_b1 );
not ( \2365_b1 , w_7368 );
not ( \2365_b0 , w_7369 );
and ( w_7368 , w_7369 , \2364_b0 );
or ( \2366_b1 , \2357_b1 , w_7370 );
or ( \2366_b0 , \2357_b0 , \2365_b0 );
not ( \2365_b0 , w_7371 );
and ( w_7371 , w_7370 , \2365_b1 );
or ( \2367_b1 , \2355_b1 , w_7373 );
not ( w_7373 , w_7374 );
and ( \2367_b0 , \2355_b0 , w_7375 );
and ( w_7374 ,  , w_7375 );
buf ( w_7373 , \2363_b1 );
not ( w_7373 , w_7376 );
not (  , w_7377 );
and ( w_7376 , w_7377 , \2363_b0 );
or ( \2368_b1 , \2366_b1 , w_7379 );
not ( w_7379 , w_7380 );
and ( \2368_b0 , \2366_b0 , w_7381 );
and ( w_7380 ,  , w_7381 );
buf ( w_7379 , \2367_b1 );
not ( w_7379 , w_7382 );
not (  , w_7383 );
and ( w_7382 , w_7383 , \2367_b0 );
buf ( \2369_b1 , \2087_b1 );
not ( \2369_b1 , w_7384 );
not ( \2369_b0 , w_7385 );
and ( w_7384 , w_7385 , \2087_b0 );
buf ( \2370_b1 , \1705_b1 );
buf ( \2370_b0 , \1705_b0 );
buf ( \2371_b1 , \2370_b1 );
not ( \2371_b1 , w_7386 );
not ( \2371_b0 , w_7387 );
and ( w_7386 , w_7387 , \2370_b0 );
or ( \2372_b1 , \2369_b1 , w_7388 );
or ( \2372_b0 , \2369_b0 , \2371_b0 );
not ( \2371_b0 , w_7389 );
and ( w_7389 , w_7388 , \2371_b1 );
or ( \2373_b1 , \b[11]_b1 , \c[3]_b1 );
xor ( \2373_b0 , \b[11]_b0 , w_7390 );
not ( w_7390 , w_7391 );
and ( w_7391 , \c[3]_b1 , \c[3]_b0 );
or ( \2374_b1 , \1708_b1 , w_7393 );
not ( w_7393 , w_7394 );
and ( \2374_b0 , \1708_b0 , w_7395 );
and ( w_7394 ,  , w_7395 );
buf ( w_7393 , \2373_b1 );
not ( w_7393 , w_7396 );
not (  , w_7397 );
and ( w_7396 , w_7397 , \2373_b0 );
or ( \2375_b1 , \2372_b1 , w_7399 );
not ( w_7399 , w_7400 );
and ( \2375_b0 , \2372_b0 , w_7401 );
and ( w_7400 ,  , w_7401 );
buf ( w_7399 , \2374_b1 );
not ( w_7399 , w_7402 );
not (  , w_7403 );
and ( w_7402 , w_7403 , \2374_b0 );
or ( \2376_b1 , \2368_b1 , w_7404 );
xor ( \2376_b0 , \2368_b0 , w_7406 );
not ( w_7406 , w_7407 );
and ( w_7407 , w_7404 , w_7405 );
buf ( w_7404 , \2375_b1 );
not ( w_7404 , w_7408 );
not ( w_7405 , w_7409 );
and ( w_7408 , w_7409 , \2375_b0 );
buf ( \2377_b1 , \2376_b1 );
not ( \2377_b1 , w_7410 );
not ( \2377_b0 , w_7411 );
and ( w_7410 , w_7411 , \2376_b0 );
buf ( \2378_b1 , \2377_b1 );
not ( \2378_b1 , w_7412 );
not ( \2378_b0 , w_7413 );
and ( w_7412 , w_7413 , \2377_b0 );
or ( \2379_b1 , \2349_b1 , w_7414 );
or ( \2379_b0 , \2349_b0 , \2378_b0 );
not ( \2378_b0 , w_7415 );
and ( w_7415 , w_7414 , \2378_b1 );
or ( \2380_b1 , \2376_b1 , w_7417 );
not ( w_7417 , w_7418 );
and ( \2380_b0 , \2376_b0 , w_7419 );
and ( w_7418 ,  , w_7419 );
buf ( w_7417 , \2347_b1 );
not ( w_7417 , w_7420 );
not (  , w_7421 );
and ( w_7420 , w_7421 , \2347_b0 );
or ( \2381_b1 , \2379_b1 , w_7423 );
not ( w_7423 , w_7424 );
and ( \2381_b0 , \2379_b0 , w_7425 );
and ( w_7424 ,  , w_7425 );
buf ( w_7423 , \2380_b1 );
not ( w_7423 , w_7426 );
not (  , w_7427 );
and ( w_7426 , w_7427 , \2380_b0 );
or ( \2382_b1 , \2057_b1 , \2058_b1 );
xor ( \2382_b0 , \2057_b0 , w_7428 );
not ( w_7428 , w_7429 );
and ( w_7429 , \2058_b1 , \2058_b0 );
or ( \2383_b1 , \2382_b1 , \2066_b1 );
not ( \2066_b1 , w_7430 );
and ( \2383_b0 , \2382_b0 , w_7431 );
and ( w_7430 , w_7431 , \2066_b0 );
or ( \2384_b1 , \2057_b1 , \2058_b1 );
not ( \2058_b1 , w_7432 );
and ( \2384_b0 , \2057_b0 , w_7433 );
and ( w_7432 , w_7433 , \2058_b0 );
or ( \2385_b1 , \2383_b1 , w_7434 );
or ( \2385_b0 , \2383_b0 , \2384_b0 );
not ( \2384_b0 , w_7435 );
and ( w_7435 , w_7434 , \2384_b1 );
buf ( \2386_b1 , \2385_b1 );
not ( \2386_b1 , w_7436 );
not ( \2386_b0 , w_7437 );
and ( w_7436 , w_7437 , \2385_b0 );
or ( \2387_b1 , \2381_b1 , \2386_b1 );
not ( \2386_b1 , w_7438 );
and ( \2387_b0 , \2381_b0 , w_7439 );
and ( w_7438 , w_7439 , \2386_b0 );
buf ( \2388_b1 , \2381_b1 );
not ( \2388_b1 , w_7440 );
not ( \2388_b0 , w_7441 );
and ( w_7440 , w_7441 , \2381_b0 );
or ( \2389_b1 , \2388_b1 , \2385_b1 );
not ( \2385_b1 , w_7442 );
and ( \2389_b0 , \2388_b0 , w_7443 );
and ( w_7442 , w_7443 , \2385_b0 );
or ( \2390_b1 , \2387_b1 , w_7445 );
not ( w_7445 , w_7446 );
and ( \2390_b0 , \2387_b0 , w_7447 );
and ( w_7446 ,  , w_7447 );
buf ( w_7445 , \2389_b1 );
not ( w_7445 , w_7448 );
not (  , w_7449 );
and ( w_7448 , w_7449 , \2389_b0 );
or ( \2391_b1 , \2324_b1 , \2390_b1 );
not ( \2390_b1 , w_7450 );
and ( \2391_b0 , \2324_b0 , w_7451 );
and ( w_7450 , w_7451 , \2390_b0 );
buf ( \2392_b1 , \2324_b1 );
not ( \2392_b1 , w_7452 );
not ( \2392_b0 , w_7453 );
and ( w_7452 , w_7453 , \2324_b0 );
buf ( \2393_b1 , \2390_b1 );
not ( \2393_b1 , w_7454 );
not ( \2393_b0 , w_7455 );
and ( w_7454 , w_7455 , \2390_b0 );
or ( \2394_b1 , \2392_b1 , \2393_b1 );
not ( \2393_b1 , w_7456 );
and ( \2394_b0 , \2392_b0 , w_7457 );
and ( w_7456 , w_7457 , \2393_b0 );
or ( \2395_b1 , \2391_b1 , w_7459 );
not ( w_7459 , w_7460 );
and ( \2395_b0 , \2391_b0 , w_7461 );
and ( w_7460 ,  , w_7461 );
buf ( w_7459 , \2394_b1 );
not ( w_7459 , w_7462 );
not (  , w_7463 );
and ( w_7462 , w_7463 , \2394_b0 );
buf ( \2396_b1 , \2395_b1 );
not ( \2396_b1 , w_7464 );
not ( \2396_b0 , w_7465 );
and ( w_7464 , w_7465 , \2395_b0 );
or ( \2397_b1 , \2067_b1 , \2073_b1 );
xor ( \2397_b0 , \2067_b0 , w_7466 );
not ( w_7466 , w_7467 );
and ( w_7467 , \2073_b1 , \2073_b0 );
or ( \2398_b1 , \2397_b1 , \2122_b1 );
not ( \2122_b1 , w_7468 );
and ( \2398_b0 , \2397_b0 , w_7469 );
and ( w_7468 , w_7469 , \2122_b0 );
or ( \2399_b1 , \2067_b1 , \2073_b1 );
not ( \2073_b1 , w_7470 );
and ( \2399_b0 , \2067_b0 , w_7471 );
and ( w_7470 , w_7471 , \2073_b0 );
or ( \2400_b1 , \2398_b1 , w_7472 );
or ( \2400_b0 , \2398_b0 , \2399_b0 );
not ( \2399_b0 , w_7473 );
and ( w_7473 , w_7472 , \2399_b1 );
or ( \2401_b1 , \2396_b1 , w_7475 );
not ( w_7475 , w_7476 );
and ( \2401_b0 , \2396_b0 , w_7477 );
and ( w_7476 ,  , w_7477 );
buf ( w_7475 , \2400_b1 );
not ( w_7475 , w_7478 );
not (  , w_7479 );
and ( w_7478 , w_7479 , \2400_b0 );
buf ( \2402_b1 , \2400_b1 );
not ( \2402_b1 , w_7480 );
not ( \2402_b0 , w_7481 );
and ( w_7480 , w_7481 , \2400_b0 );
or ( \2403_b1 , \2402_b1 , w_7483 );
not ( w_7483 , w_7484 );
and ( \2403_b0 , \2402_b0 , w_7485 );
and ( w_7484 ,  , w_7485 );
buf ( w_7483 , \2395_b1 );
not ( w_7483 , w_7486 );
not (  , w_7487 );
and ( w_7486 , w_7487 , \2395_b0 );
or ( \2404_b1 , \2401_b1 , w_7489 );
not ( w_7489 , w_7490 );
and ( \2404_b0 , \2401_b0 , w_7491 );
and ( w_7490 ,  , w_7491 );
buf ( w_7489 , \2403_b1 );
not ( w_7489 , w_7492 );
not (  , w_7493 );
and ( w_7492 , w_7493 , \2403_b0 );
buf ( \2405_b1 , \2404_b1 );
not ( \2405_b1 , w_7494 );
not ( \2405_b0 , w_7495 );
and ( w_7494 , w_7495 , \2404_b0 );
or ( \2406_b1 , \2289_b1 , \2405_b1 );
not ( \2405_b1 , w_7496 );
and ( \2406_b0 , \2289_b0 , w_7497 );
and ( w_7496 , w_7497 , \2405_b0 );
buf ( \2407_b1 , \2289_b1 );
not ( \2407_b1 , w_7498 );
not ( \2407_b0 , w_7499 );
and ( w_7498 , w_7499 , \2289_b0 );
or ( \2408_b1 , \2407_b1 , \2404_b1 );
not ( \2404_b1 , w_7500 );
and ( \2408_b0 , \2407_b0 , w_7501 );
and ( w_7500 , w_7501 , \2404_b0 );
or ( \2409_b1 , \2406_b1 , w_7503 );
not ( w_7503 , w_7504 );
and ( \2409_b0 , \2406_b0 , w_7505 );
and ( w_7504 ,  , w_7505 );
buf ( w_7503 , \2408_b1 );
not ( w_7503 , w_7506 );
not (  , w_7507 );
and ( w_7506 , w_7507 , \2408_b0 );
or ( \2410_b1 , \155_b1 , \202_b1 );
xor ( \2410_b0 , \155_b0 , w_7508 );
not ( w_7508 , w_7509 );
and ( w_7509 , \202_b1 , \202_b0 );
or ( \2411_b1 , \2410_b1 , \344_b1 );
xor ( \2411_b0 , \2410_b0 , w_7510 );
not ( w_7510 , w_7511 );
and ( w_7511 , \344_b1 , \344_b0 );
buf ( \2412_b1 , \2411_b1 );
not ( \2412_b1 , w_7512 );
not ( \2412_b0 , w_7513 );
and ( w_7512 , w_7513 , \2411_b0 );
buf ( \2413_b1 , \2412_b1 );
not ( \2413_b1 , w_7514 );
not ( \2413_b0 , w_7515 );
and ( w_7514 , w_7515 , \2412_b0 );
or ( \2414_b1 , \2409_b1 , w_7517 );
not ( w_7517 , w_7518 );
and ( \2414_b0 , \2409_b0 , w_7519 );
and ( w_7518 ,  , w_7519 );
buf ( w_7517 , \2413_b1 );
not ( w_7517 , w_7520 );
not (  , w_7521 );
and ( w_7520 , w_7521 , \2413_b0 );
or ( \2415_b1 , \a[13]_b1 , w_7522 );
or ( \2415_b0 , \a[13]_b0 , \d[13]_b0 );
not ( \d[13]_b0 , w_7523 );
and ( w_7523 , w_7522 , \d[13]_b1 );
buf ( \2416_b1 , \2415_b1 );
not ( \2416_b1 , w_7524 );
not ( \2416_b0 , w_7525 );
and ( w_7524 , w_7525 , \2415_b0 );
buf ( \2417_b1 , \648_b1 );
not ( \2417_b1 , w_7526 );
not ( \2417_b0 , w_7527 );
and ( w_7526 , w_7527 , \648_b0 );
or ( \2418_b1 , \2416_b1 , w_7528 );
or ( \2418_b0 , \2416_b0 , \2417_b0 );
not ( \2417_b0 , w_7529 );
and ( w_7529 , w_7528 , \2417_b1 );
or ( \2419_b1 , \a[13]_b1 , w_7530 );
or ( \2419_b0 , \a[13]_b0 , \b[13]_b0 );
not ( \b[13]_b0 , w_7531 );
and ( w_7531 , w_7530 , \b[13]_b1 );
or ( \2420_b1 , \667_b1 , w_7533 );
not ( w_7533 , w_7534 );
and ( \2420_b0 , \667_b0 , w_7535 );
and ( w_7534 ,  , w_7535 );
buf ( w_7533 , \2419_b1 );
not ( w_7533 , w_7536 );
not (  , w_7537 );
and ( w_7536 , w_7537 , \2419_b0 );
or ( \2421_b1 , \2418_b1 , w_7539 );
not ( w_7539 , w_7540 );
and ( \2421_b0 , \2418_b0 , w_7541 );
and ( w_7540 ,  , w_7541 );
buf ( w_7539 , \2420_b1 );
not ( w_7539 , w_7542 );
not (  , w_7543 );
and ( w_7542 , w_7543 , \2420_b0 );
or ( \2422_b1 , \b[13]_b1 , \c[13]_b1 );
not ( \c[13]_b1 , w_7544 );
and ( \2422_b0 , \b[13]_b0 , w_7545 );
and ( w_7544 , w_7545 , \c[13]_b0 );
buf ( \2423_b1 , \2422_b1 );
not ( \2423_b1 , w_7546 );
not ( \2423_b0 , w_7547 );
and ( w_7546 , w_7547 , \2422_b0 );
buf ( \2424_b1 , \922_b1 );
not ( \2424_b1 , w_7548 );
not ( \2424_b0 , w_7549 );
and ( w_7548 , w_7549 , \922_b0 );
or ( \2425_b1 , \2423_b1 , w_7550 );
or ( \2425_b0 , \2423_b0 , \2424_b0 );
not ( \2424_b0 , w_7551 );
and ( w_7551 , w_7550 , \2424_b1 );
or ( \2426_b1 , \c[13]_b1 , \d[13]_b1 );
xor ( \2426_b0 , \c[13]_b0 , w_7552 );
not ( w_7552 , w_7553 );
and ( w_7553 , \d[13]_b1 , \d[13]_b0 );
or ( \2427_b1 , \697_b1 , \2426_b1 );
not ( \2426_b1 , w_7554 );
and ( \2427_b0 , \697_b0 , w_7555 );
and ( w_7554 , w_7555 , \2426_b0 );
buf ( \2428_b1 , \757_b1 );
not ( \2428_b1 , w_7556 );
not ( \2428_b0 , w_7557 );
and ( w_7556 , w_7557 , \757_b0 );
or ( \2429_b1 , \2428_b1 , w_7559 );
not ( w_7559 , w_7560 );
and ( \2429_b0 , \2428_b0 , w_7561 );
and ( w_7560 ,  , w_7561 );
buf ( w_7559 , \781_b1 );
not ( w_7559 , w_7562 );
not (  , w_7563 );
and ( w_7562 , w_7563 , \781_b0 );
buf ( \2430_b1 , \2429_b1 );
not ( \2430_b1 , w_7564 );
not ( \2430_b0 , w_7565 );
and ( w_7564 , w_7565 , \2429_b0 );
or ( \2431_b1 , \777_b1 , w_7566 );
or ( \2431_b0 , \777_b0 , \758_b0 );
not ( \758_b0 , w_7567 );
and ( w_7567 , w_7566 , \758_b1 );
buf ( \2432_b1 , \758_b1 );
not ( \2432_b1 , w_7568 );
not ( \2432_b0 , w_7569 );
and ( w_7568 , w_7569 , \758_b0 );
buf ( \2435_b1 , \2434_b1 );
not ( \2435_b1 , w_7570 );
not ( \2435_b0 , w_7571 );
and ( w_7570 , w_7571 , \2434_b0 );
or ( \2436_b1 , \2430_b1 , w_7572 );
or ( \2436_b0 , \2430_b0 , \2435_b0 );
not ( \2435_b0 , w_7573 );
and ( w_7573 , w_7572 , \2435_b1 );
or ( \2437_b1 , \2434_b1 , w_7574 );
or ( \2437_b0 , \2434_b0 , \2429_b0 );
not ( \2429_b0 , w_7575 );
and ( w_7575 , w_7574 , \2429_b1 );
or ( \2438_b1 , \2436_b1 , w_7577 );
not ( w_7577 , w_7578 );
and ( \2438_b0 , \2436_b0 , w_7579 );
and ( w_7578 ,  , w_7579 );
buf ( w_7577 , \2437_b1 );
not ( w_7577 , w_7580 );
not (  , w_7581 );
and ( w_7580 , w_7581 , \2437_b0 );
buf ( \2439_b1 , \2438_b1 );
not ( \2439_b1 , w_7582 );
not ( \2439_b0 , w_7583 );
and ( w_7582 , w_7583 , \2438_b0 );
buf ( \2440_b1 , \707_b1 );
not ( \2440_b1 , w_7584 );
not ( \2440_b0 , w_7585 );
and ( w_7584 , w_7585 , \707_b0 );
or ( \2441_b1 , \2439_b1 , w_7586 );
or ( \2441_b0 , \2439_b0 , \2440_b0 );
not ( \2440_b0 , w_7587 );
and ( w_7587 , w_7586 , \2440_b1 );
buf ( \2442_b1 , \842_b1 );
not ( \2442_b1 , w_7588 );
not ( \2442_b0 , w_7589 );
and ( w_7588 , w_7589 , \842_b0 );
or ( \2443_b1 , \2442_b1 , w_7591 );
not ( w_7591 , w_7592 );
and ( \2443_b0 , \2442_b0 , w_7593 );
and ( w_7592 ,  , w_7593 );
buf ( w_7591 , \866_b1 );
not ( w_7591 , w_7594 );
not (  , w_7595 );
and ( w_7594 , w_7595 , \866_b0 );
buf ( \2444_b1 , \2443_b1 );
not ( \2444_b1 , w_7596 );
not ( \2444_b0 , w_7597 );
and ( w_7596 , w_7597 , \2443_b0 );
or ( \2445_b1 , \862_b1 , w_7598 );
or ( \2445_b0 , \862_b0 , \843_b0 );
not ( \843_b0 , w_7599 );
and ( w_7599 , w_7598 , \843_b1 );
buf ( \2446_b1 , \843_b1 );
not ( \2446_b1 , w_7600 );
not ( \2446_b0 , w_7601 );
and ( w_7600 , w_7601 , \843_b0 );
buf ( \2449_b1 , \2448_b1 );
not ( \2449_b1 , w_7602 );
not ( \2449_b0 , w_7603 );
and ( w_7602 , w_7603 , \2448_b0 );
or ( \2450_b1 , \2444_b1 , w_7604 );
or ( \2450_b0 , \2444_b0 , \2449_b0 );
not ( \2449_b0 , w_7605 );
and ( w_7605 , w_7604 , \2449_b1 );
or ( \2451_b1 , \2448_b1 , w_7606 );
or ( \2451_b0 , \2448_b0 , \2443_b0 );
not ( \2443_b0 , w_7607 );
and ( w_7607 , w_7606 , \2443_b1 );
or ( \2452_b1 , \2450_b1 , w_7609 );
not ( w_7609 , w_7610 );
and ( \2452_b0 , \2450_b0 , w_7611 );
and ( w_7610 ,  , w_7611 );
buf ( w_7609 , \2451_b1 );
not ( w_7609 , w_7612 );
not (  , w_7613 );
and ( w_7612 , w_7613 , \2451_b0 );
or ( \2453_b1 , \880_b1 , \2452_b1 );
not ( \2452_b1 , w_7614 );
and ( \2453_b0 , \880_b0 , w_7615 );
and ( w_7614 , w_7615 , \2452_b0 );
buf ( \2454_b1 , \d[13]_b1 );
not ( \2454_b1 , w_7616 );
not ( \2454_b0 , w_7617 );
and ( w_7616 , w_7617 , \d[13]_b0 );
buf ( \2455_b1 , \894_b1 );
not ( \2455_b1 , w_7618 );
not ( \2455_b0 , w_7619 );
and ( w_7618 , w_7619 , \894_b0 );
or ( \2456_b1 , \2454_b1 , w_7620 );
or ( \2456_b0 , \2454_b0 , \2455_b0 );
not ( \2455_b0 , w_7621 );
and ( w_7621 , w_7620 , \2455_b1 );
or ( \2457_b1 , \885_b1 , \b[13]_b1 );
not ( \b[13]_b1 , w_7622 );
and ( \2457_b0 , \885_b0 , w_7623 );
and ( w_7622 , w_7623 , \b[13]_b0 );
or ( \2458_b1 , \907_b1 , \c[13]_b1 );
not ( \c[13]_b1 , w_7624 );
and ( \2458_b0 , \907_b0 , w_7625 );
and ( w_7624 , w_7625 , \c[13]_b0 );
or ( \2459_b1 , \2457_b1 , w_7627 );
not ( w_7627 , w_7628 );
and ( \2459_b0 , \2457_b0 , w_7629 );
and ( w_7628 ,  , w_7629 );
buf ( w_7627 , \2458_b1 );
not ( w_7627 , w_7630 );
not (  , w_7631 );
and ( w_7630 , w_7631 , \2458_b0 );
or ( \2460_b1 , \2456_b1 , w_7633 );
not ( w_7633 , w_7634 );
and ( \2460_b0 , \2456_b0 , w_7635 );
and ( w_7634 ,  , w_7635 );
buf ( w_7633 , \2459_b1 );
not ( w_7633 , w_7636 );
not (  , w_7637 );
and ( w_7636 , w_7637 , \2459_b0 );
or ( \2461_b1 , \2453_b1 , w_7639 );
not ( w_7639 , w_7640 );
and ( \2461_b0 , \2453_b0 , w_7641 );
and ( w_7640 ,  , w_7641 );
buf ( w_7639 , \2460_b1 );
not ( w_7639 , w_7642 );
not (  , w_7643 );
and ( w_7642 , w_7643 , \2460_b0 );
or ( \2462_b1 , \2441_b1 , w_7645 );
not ( w_7645 , w_7646 );
and ( \2462_b0 , \2441_b0 , w_7647 );
and ( w_7646 ,  , w_7647 );
buf ( w_7645 , \2461_b1 );
not ( w_7645 , w_7648 );
not (  , w_7649 );
and ( w_7648 , w_7649 , \2461_b0 );
or ( \2463_b1 , \2427_b1 , w_7651 );
not ( w_7651 , w_7652 );
and ( \2463_b0 , \2427_b0 , w_7653 );
and ( w_7652 ,  , w_7653 );
buf ( w_7651 , \2462_b1 );
not ( w_7651 , w_7654 );
not (  , w_7655 );
and ( w_7654 , w_7655 , \2462_b0 );
or ( \2464_b1 , \2425_b1 , w_7657 );
not ( w_7657 , w_7658 );
and ( \2464_b0 , \2425_b0 , w_7659 );
and ( w_7658 ,  , w_7659 );
buf ( w_7657 , \2463_b1 );
not ( w_7657 , w_7660 );
not (  , w_7661 );
and ( w_7660 , w_7661 , \2463_b0 );
or ( \2465_b1 , \2421_b1 , w_7663 );
not ( w_7663 , w_7664 );
and ( \2465_b0 , \2421_b0 , w_7665 );
and ( w_7664 ,  , w_7665 );
buf ( w_7663 , \2464_b1 );
not ( w_7663 , w_7666 );
not (  , w_7667 );
and ( w_7666 , w_7667 , \2464_b0 );
or ( \2466_b1 , \915_b1 , \916_b1 );
xor ( \2466_b0 , \915_b0 , w_7668 );
not ( w_7668 , w_7669 );
and ( w_7669 , \916_b1 , \916_b0 );
buf ( \2467_b1 , \705_b1 );
not ( \2467_b1 , w_7670 );
not ( \2467_b0 , w_7671 );
and ( w_7670 , w_7671 , \705_b0 );
or ( \2468_b1 , \907_b1 , w_7673 );
not ( w_7673 , w_7674 );
and ( \2468_b0 , \907_b0 , w_7675 );
and ( w_7674 ,  , w_7675 );
buf ( w_7673 , \885_b1 );
not ( w_7673 , w_7676 );
not (  , w_7677 );
and ( w_7676 , w_7677 , \885_b0 );
or ( \2469_b1 , \893_b1 , w_7679 );
not ( w_7679 , w_7680 );
and ( \2469_b0 , \893_b0 , w_7681 );
and ( w_7680 ,  , w_7681 );
buf ( w_7679 , \2468_b1 );
not ( w_7679 , w_7682 );
not (  , w_7683 );
and ( w_7682 , w_7683 , \2468_b0 );
or ( \2470_b1 , \879_b1 , w_7685 );
not ( w_7685 , w_7686 );
and ( \2470_b0 , \879_b0 , w_7687 );
and ( w_7686 ,  , w_7687 );
buf ( w_7685 , \2469_b1 );
not ( w_7685 , w_7688 );
not (  , w_7689 );
and ( w_7688 , w_7689 , \2469_b0 );
or ( \2471_b1 , \2467_b1 , w_7691 );
not ( w_7691 , w_7692 );
and ( \2471_b0 , \2467_b0 , w_7693 );
and ( w_7692 ,  , w_7693 );
buf ( w_7691 , \2470_b1 );
not ( w_7691 , w_7694 );
not (  , w_7695 );
and ( w_7694 , w_7695 , \2470_b0 );
or ( \2472_b1 , \1666_b1 , w_7697 );
not ( w_7697 , w_7698 );
and ( \2472_b0 , \1666_b0 , w_7699 );
and ( w_7698 ,  , w_7699 );
buf ( w_7697 , \2471_b1 );
not ( w_7697 , w_7700 );
not (  , w_7701 );
and ( w_7700 , w_7701 , \2471_b0 );
or ( \2473_b1 , \2412_b1 , w_7703 );
not ( w_7703 , w_7704 );
and ( \2473_b0 , \2412_b0 , w_7705 );
and ( w_7704 ,  , w_7705 );
buf ( w_7703 , \2472_b1 );
not ( w_7703 , w_7706 );
not (  , w_7707 );
and ( w_7706 , w_7707 , \2472_b0 );
or ( \2474_b1 , \2473_b1 , w_7709 );
not ( w_7709 , w_7710 );
and ( \2474_b0 , \2473_b0 , w_7711 );
and ( w_7710 ,  , w_7711 );
buf ( w_7709 , \695_b1 );
not ( w_7709 , w_7712 );
not (  , w_7713 );
and ( w_7712 , w_7713 , \695_b0 );
or ( \2475_b1 , \2466_b1 , \2474_b1 );
not ( \2474_b1 , w_7714 );
and ( \2475_b0 , \2466_b0 , w_7715 );
and ( w_7714 , w_7715 , \2474_b0 );
or ( \2476_b1 , \2475_b1 , w_7717 );
not ( w_7717 , w_7718 );
and ( \2476_b0 , \2475_b0 , w_7719 );
and ( w_7718 ,  , w_7719 );
buf ( w_7717 , \a[13]_b1 );
not ( w_7717 , w_7720 );
not (  , w_7721 );
and ( w_7720 , w_7721 , \a[13]_b0 );
buf ( \2478_b1 , \2344_b1 );
not ( \2478_b1 , w_7722 );
not ( \2478_b0 , w_7723 );
and ( w_7722 , w_7723 , \2344_b0 );
buf ( \2479_b1 , \2341_b1 );
not ( \2479_b1 , w_7724 );
not ( \2479_b0 , w_7725 );
and ( w_7724 , w_7725 , \2341_b0 );
or ( \2480_b1 , \2478_b1 , w_7726 );
or ( \2480_b0 , \2478_b0 , \2479_b0 );
not ( \2479_b0 , w_7727 );
and ( w_7727 , w_7726 , \2479_b1 );
or ( \2481_b1 , \b[2]_b1 , \c[13]_b1 );
xor ( \2481_b0 , \b[2]_b0 , w_7728 );
not ( w_7728 , w_7729 );
and ( w_7729 , \c[13]_b1 , \c[13]_b0 );
or ( \2482_b1 , \2075_b1 , w_7731 );
not ( w_7731 , w_7732 );
and ( \2482_b0 , \2075_b0 , w_7733 );
and ( w_7732 ,  , w_7733 );
buf ( w_7731 , \2481_b1 );
not ( w_7731 , w_7734 );
not (  , w_7735 );
and ( w_7734 , w_7735 , \2481_b0 );
or ( \2483_b1 , \2480_b1 , w_7737 );
not ( w_7737 , w_7738 );
and ( \2483_b0 , \2480_b0 , w_7739 );
and ( w_7738 ,  , w_7739 );
buf ( w_7737 , \2482_b1 );
not ( w_7737 , w_7740 );
not (  , w_7741 );
and ( w_7740 , w_7741 , \2482_b0 );
buf ( \2484_b1 , \2300_b1 );
not ( \2484_b1 , w_7742 );
not ( \2484_b0 , w_7743 );
and ( w_7742 , w_7743 , \2300_b0 );
or ( \2485_b1 , \2484_b1 , w_7745 );
not ( w_7745 , w_7746 );
and ( \2485_b0 , \2484_b0 , w_7747 );
and ( w_7746 ,  , w_7747 );
buf ( w_7745 , \2295_b1 );
not ( w_7745 , w_7748 );
not (  , w_7749 );
and ( w_7748 , w_7749 , \2295_b0 );
or ( \2486_b1 , \2483_b1 , \2485_b1 );
xor ( \2486_b0 , \2483_b0 , w_7750 );
not ( w_7750 , w_7751 );
and ( w_7751 , \2485_b1 , \2485_b0 );
buf ( \2487_b1 , \2334_b1 );
not ( \2487_b1 , w_7752 );
not ( \2487_b0 , w_7753 );
and ( w_7752 , w_7753 , \2334_b0 );
buf ( \2488_b1 , \2107_b1 );
not ( \2488_b1 , w_7754 );
not ( \2488_b0 , w_7755 );
and ( w_7754 , w_7755 , \2107_b0 );
or ( \2489_b1 , \2487_b1 , w_7756 );
or ( \2489_b0 , \2487_b0 , \2488_b0 );
not ( \2488_b0 , w_7757 );
and ( w_7757 , w_7756 , \2488_b1 );
or ( \2490_b1 , \b[4]_b1 , \c[11]_b1 );
xor ( \2490_b0 , \b[4]_b0 , w_7758 );
not ( w_7758 , w_7759 );
and ( w_7759 , \c[11]_b1 , \c[11]_b0 );
or ( \2491_b1 , \1689_b1 , w_7761 );
not ( w_7761 , w_7762 );
and ( \2491_b0 , \1689_b0 , w_7763 );
and ( w_7762 ,  , w_7763 );
buf ( w_7761 , \2490_b1 );
not ( w_7761 , w_7764 );
not (  , w_7765 );
and ( w_7764 , w_7765 , \2490_b0 );
or ( \2492_b1 , \2489_b1 , w_7767 );
not ( w_7767 , w_7768 );
and ( \2492_b0 , \2489_b0 , w_7769 );
and ( w_7768 ,  , w_7769 );
buf ( w_7767 , \2491_b1 );
not ( w_7767 , w_7770 );
not (  , w_7771 );
and ( w_7770 , w_7771 , \2491_b0 );
or ( \2493_b1 , \2486_b1 , \2492_b1 );
xor ( \2493_b0 , \2486_b0 , w_7772 );
not ( w_7772 , w_7773 );
and ( w_7773 , \2492_b1 , \2492_b0 );
buf ( \2494_b1 , \2493_b1 );
not ( \2494_b1 , w_7774 );
not ( \2494_b0 , w_7775 );
and ( w_7774 , w_7775 , \2493_b0 );
buf ( \2495_b1 , \2494_b1 );
not ( \2495_b1 , w_7776 );
not ( \2495_b0 , w_7777 );
and ( w_7776 , w_7777 , \2494_b0 );
buf ( \2496_b1 , \1773_b1 );
not ( \2496_b1 , w_7778 );
not ( \2496_b0 , w_7779 );
and ( w_7778 , w_7779 , \1773_b0 );
or ( \2497_b1 , \b[6]_b1 , \c[9]_b1 );
xor ( \2497_b0 , \b[6]_b0 , w_7780 );
not ( w_7780 , w_7781 );
and ( w_7781 , \c[9]_b1 , \c[9]_b0 );
buf ( \2498_b1 , \2497_b1 );
not ( \2498_b1 , w_7782 );
not ( \2498_b0 , w_7783 );
and ( w_7782 , w_7783 , \2497_b0 );
or ( \2499_b1 , \2496_b1 , w_7784 );
or ( \2499_b0 , \2496_b0 , \2498_b0 );
not ( \2498_b0 , w_7785 );
and ( w_7785 , w_7784 , \2498_b1 );
or ( \2500_b1 , \1770_b1 , w_7787 );
not ( w_7787 , w_7788 );
and ( \2500_b0 , \1770_b0 , w_7789 );
and ( w_7788 ,  , w_7789 );
buf ( w_7787 , \2353_b1 );
not ( w_7787 , w_7790 );
not (  , w_7791 );
and ( w_7790 , w_7791 , \2353_b0 );
or ( \2501_b1 , \2499_b1 , w_7793 );
not ( w_7793 , w_7794 );
and ( \2501_b0 , \2499_b0 , w_7795 );
and ( w_7794 ,  , w_7795 );
buf ( w_7793 , \2500_b1 );
not ( w_7793 , w_7796 );
not (  , w_7797 );
and ( w_7796 , w_7797 , \2500_b0 );
buf ( \2502_b1 , \2361_b1 );
not ( \2502_b1 , w_7798 );
not ( \2502_b0 , w_7799 );
and ( w_7798 , w_7799 , \2361_b0 );
buf ( \2503_b1 , \1743_b1 );
not ( \2503_b1 , w_7800 );
not ( \2503_b0 , w_7801 );
and ( w_7800 , w_7801 , \1743_b0 );
or ( \2504_b1 , \2502_b1 , w_7802 );
or ( \2504_b0 , \2502_b0 , \2503_b0 );
not ( \2503_b0 , w_7803 );
and ( w_7803 , w_7802 , \2503_b1 );
or ( \2505_b1 , \b[8]_b1 , \c[7]_b1 );
xor ( \2505_b0 , \b[8]_b0 , w_7804 );
not ( w_7804 , w_7805 );
and ( w_7805 , \c[7]_b1 , \c[7]_b0 );
or ( \2506_b1 , \1747_b1 , w_7807 );
not ( w_7807 , w_7808 );
and ( \2506_b0 , \1747_b0 , w_7809 );
and ( w_7808 ,  , w_7809 );
buf ( w_7807 , \2505_b1 );
not ( w_7807 , w_7810 );
not (  , w_7811 );
and ( w_7810 , w_7811 , \2505_b0 );
or ( \2507_b1 , \2504_b1 , w_7813 );
not ( w_7813 , w_7814 );
and ( \2507_b0 , \2504_b0 , w_7815 );
and ( w_7814 ,  , w_7815 );
buf ( w_7813 , \2506_b1 );
not ( w_7813 , w_7816 );
not (  , w_7817 );
and ( w_7816 , w_7817 , \2506_b0 );
or ( \2508_b1 , \2501_b1 , \2507_b1 );
xor ( \2508_b0 , \2501_b0 , w_7818 );
not ( w_7818 , w_7819 );
and ( w_7819 , \2507_b1 , \2507_b0 );
buf ( \2509_b1 , \2328_b1 );
not ( \2509_b1 , w_7820 );
not ( \2509_b0 , w_7821 );
and ( w_7820 , w_7821 , \2328_b0 );
buf ( \2510_b1 , \2052_b1 );
not ( \2510_b1 , w_7822 );
not ( \2510_b0 , w_7823 );
and ( w_7822 , w_7823 , \2052_b0 );
or ( \2511_b1 , \2509_b1 , w_7824 );
or ( \2511_b0 , \2509_b0 , \2510_b0 );
not ( \2510_b0 , w_7825 );
and ( w_7825 , w_7824 , \2510_b1 );
or ( \2512_b1 , \b[10]_b1 , \c[5]_b1 );
xor ( \2512_b0 , \b[10]_b0 , w_7826 );
not ( w_7826 , w_7827 );
and ( w_7827 , \c[5]_b1 , \c[5]_b0 );
or ( \2513_b1 , \1678_b1 , w_7829 );
not ( w_7829 , w_7830 );
and ( \2513_b0 , \1678_b0 , w_7831 );
and ( w_7830 ,  , w_7831 );
buf ( w_7829 , \2512_b1 );
not ( w_7829 , w_7832 );
not (  , w_7833 );
and ( w_7832 , w_7833 , \2512_b0 );
or ( \2514_b1 , \2511_b1 , w_7835 );
not ( w_7835 , w_7836 );
and ( \2514_b0 , \2511_b0 , w_7837 );
and ( w_7836 ,  , w_7837 );
buf ( w_7835 , \2513_b1 );
not ( w_7835 , w_7838 );
not (  , w_7839 );
and ( w_7838 , w_7839 , \2513_b0 );
or ( \2515_b1 , \2508_b1 , \2514_b1 );
xor ( \2515_b0 , \2508_b0 , w_7840 );
not ( w_7840 , w_7841 );
and ( w_7841 , \2514_b1 , \2514_b0 );
buf ( \2516_b1 , \2515_b1 );
not ( \2516_b1 , w_7842 );
not ( \2516_b0 , w_7843 );
and ( w_7842 , w_7843 , \2515_b0 );
buf ( \2517_b1 , \2516_b1 );
not ( \2517_b1 , w_7844 );
not ( \2517_b0 , w_7845 );
and ( w_7844 , w_7845 , \2516_b0 );
or ( \2518_b1 , \2495_b1 , w_7846 );
or ( \2518_b0 , \2495_b0 , \2517_b0 );
not ( \2517_b0 , w_7847 );
and ( w_7847 , w_7846 , \2517_b1 );
or ( \2519_b1 , \2493_b1 , w_7849 );
not ( w_7849 , w_7850 );
and ( \2519_b0 , \2493_b0 , w_7851 );
and ( w_7850 ,  , w_7851 );
buf ( w_7849 , \2515_b1 );
not ( w_7849 , w_7852 );
not (  , w_7853 );
and ( w_7852 , w_7853 , \2515_b0 );
or ( \2520_b1 , \2518_b1 , w_7855 );
not ( w_7855 , w_7856 );
and ( \2520_b0 , \2518_b0 , w_7857 );
and ( w_7856 ,  , w_7857 );
buf ( w_7855 , \2519_b1 );
not ( w_7855 , w_7858 );
not (  , w_7859 );
and ( w_7858 , w_7859 , \2519_b0 );
buf ( \2521_b1 , \2304_b1 );
not ( \2521_b1 , w_7860 );
not ( \2521_b0 , w_7861 );
and ( w_7860 , w_7861 , \2304_b0 );
buf ( \2522_b1 , \2313_b1 );
not ( \2522_b1 , w_7862 );
not ( \2522_b0 , w_7863 );
and ( w_7862 , w_7863 , \2313_b0 );
or ( \2523_b1 , \2521_b1 , w_7864 );
or ( \2523_b0 , \2521_b0 , \2522_b0 );
not ( \2522_b0 , w_7865 );
and ( w_7865 , w_7864 , \2522_b1 );
or ( \2524_b1 , \2523_b1 , w_7867 );
not ( w_7867 , w_7868 );
and ( \2524_b0 , \2523_b0 , w_7869 );
and ( w_7868 ,  , w_7869 );
buf ( w_7867 , \2308_b1 );
not ( w_7867 , w_7870 );
not (  , w_7871 );
and ( w_7870 , w_7871 , \2308_b0 );
buf ( \2525_b1 , \2304_b1 );
not ( \2525_b1 , w_7872 );
not ( \2525_b0 , w_7873 );
and ( w_7872 , w_7873 , \2304_b0 );
or ( \2526_b1 , \2525_b1 , w_7875 );
not ( w_7875 , w_7876 );
and ( \2526_b0 , \2525_b0 , w_7877 );
and ( w_7876 ,  , w_7877 );
buf ( w_7875 , \2314_b1 );
not ( w_7875 , w_7878 );
not (  , w_7879 );
and ( w_7878 , w_7879 , \2314_b0 );
or ( \2527_b1 , \2524_b1 , w_7881 );
not ( w_7881 , w_7882 );
and ( \2527_b0 , \2524_b0 , w_7883 );
and ( w_7882 ,  , w_7883 );
buf ( w_7881 , \2526_b1 );
not ( w_7881 , w_7884 );
not (  , w_7885 );
and ( w_7884 , w_7885 , \2526_b0 );
or ( \2528_b1 , \2520_b1 , w_7886 );
xor ( \2528_b0 , \2520_b0 , w_7888 );
not ( w_7888 , w_7889 );
and ( w_7889 , w_7886 , w_7887 );
buf ( w_7886 , \2527_b1 );
not ( w_7886 , w_7890 );
not ( w_7887 , w_7891 );
and ( w_7890 , w_7891 , \2527_b0 );
buf ( \2529_b1 , \2528_b1 );
not ( \2529_b1 , w_7892 );
not ( \2529_b0 , w_7893 );
and ( w_7892 , w_7893 , \2528_b0 );
or ( \2530_b1 , \2330_b1 , \2336_b1 );
xor ( \2530_b0 , \2330_b0 , w_7894 );
not ( w_7894 , w_7895 );
and ( w_7895 , \2336_b1 , \2336_b0 );
or ( \2531_b1 , \2530_b1 , \2346_b1 );
not ( \2346_b1 , w_7896 );
and ( \2531_b0 , \2530_b0 , w_7897 );
and ( w_7896 , w_7897 , \2346_b0 );
or ( \2532_b1 , \2330_b1 , \2336_b1 );
not ( \2336_b1 , w_7898 );
and ( \2532_b0 , \2330_b0 , w_7899 );
and ( w_7898 , w_7899 , \2336_b0 );
or ( \2533_b1 , \2531_b1 , w_7900 );
or ( \2533_b0 , \2531_b0 , \2532_b0 );
not ( \2532_b0 , w_7901 );
and ( w_7901 , w_7900 , \2532_b1 );
or ( \2534_b1 , \c[14]_b1 , \c[13]_b1 );
xor ( \2534_b0 , \c[14]_b0 , w_7902 );
not ( w_7902 , w_7903 );
and ( w_7903 , \c[13]_b1 , \c[13]_b0 );
or ( \2535_b1 , \2534_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_7904 );
and ( \2535_b0 , \2534_b0 , w_7905 );
and ( w_7904 , w_7905 , \b[0]_b0 );
buf ( \2536_b1 , \1756_b1 );
not ( \2536_b1 , w_7906 );
not ( \2536_b0 , w_7907 );
and ( w_7906 , w_7907 , \1756_b0 );
buf ( \2537_b1 , \2293_b1 );
not ( \2537_b1 , w_7908 );
not ( \2537_b0 , w_7909 );
and ( w_7908 , w_7909 , \2293_b0 );
or ( \2538_b1 , \2536_b1 , w_7910 );
or ( \2538_b0 , \2536_b0 , \2537_b0 );
not ( \2537_b0 , w_7911 );
and ( w_7911 , w_7910 , \2537_b1 );
or ( \2539_b1 , \c[1]_b1 , \b[14]_b1 );
xor ( \2539_b0 , \c[1]_b0 , w_7912 );
not ( w_7912 , w_7913 );
and ( w_7913 , \b[14]_b1 , \b[14]_b0 );
or ( \2540_b1 , \2539_b1 , w_7915 );
not ( w_7915 , w_7916 );
and ( \2540_b0 , \2539_b0 , w_7917 );
and ( w_7916 ,  , w_7917 );
buf ( w_7915 , \c[0]_b1 );
not ( w_7915 , w_7918 );
not (  , w_7919 );
and ( w_7918 , w_7919 , \c[0]_b0 );
or ( \2541_b1 , \2538_b1 , w_7921 );
not ( w_7921 , w_7922 );
and ( \2541_b0 , \2538_b0 , w_7923 );
and ( w_7922 ,  , w_7923 );
buf ( w_7921 , \2540_b1 );
not ( w_7921 , w_7924 );
not (  , w_7925 );
and ( w_7924 , w_7925 , \2540_b0 );
or ( \2542_b1 , \2535_b1 , \2541_b1 );
xor ( \2542_b0 , \2535_b0 , w_7926 );
not ( w_7926 , w_7927 );
and ( w_7927 , \2541_b1 , \2541_b0 );
buf ( \2543_b1 , \2373_b1 );
not ( \2543_b1 , w_7928 );
not ( \2543_b0 , w_7929 );
and ( w_7928 , w_7929 , \2373_b0 );
buf ( \2544_b1 , \1705_b1 );
not ( \2544_b1 , w_7930 );
not ( \2544_b0 , w_7931 );
and ( w_7930 , w_7931 , \1705_b0 );
or ( \2545_b1 , \2543_b1 , w_7932 );
or ( \2545_b0 , \2543_b0 , \2544_b0 );
not ( \2544_b0 , w_7933 );
and ( w_7933 , w_7932 , \2544_b1 );
or ( \2546_b1 , \b[12]_b1 , \c[3]_b1 );
xor ( \2546_b0 , \b[12]_b0 , w_7934 );
not ( w_7934 , w_7935 );
and ( w_7935 , \c[3]_b1 , \c[3]_b0 );
or ( \2547_b1 , \1708_b1 , w_7937 );
not ( w_7937 , w_7938 );
and ( \2547_b0 , \1708_b0 , w_7939 );
and ( w_7938 ,  , w_7939 );
buf ( w_7937 , \2546_b1 );
not ( w_7937 , w_7940 );
not (  , w_7941 );
and ( w_7940 , w_7941 , \2546_b0 );
or ( \2548_b1 , \2545_b1 , w_7943 );
not ( w_7943 , w_7944 );
and ( \2548_b0 , \2545_b0 , w_7945 );
and ( w_7944 ,  , w_7945 );
buf ( w_7943 , \2547_b1 );
not ( w_7943 , w_7946 );
not (  , w_7947 );
and ( w_7946 , w_7947 , \2547_b0 );
or ( \2549_b1 , \2542_b1 , \2548_b1 );
xor ( \2549_b0 , \2542_b0 , w_7948 );
not ( w_7948 , w_7949 );
and ( w_7949 , \2548_b1 , \2548_b0 );
or ( \2550_b1 , \2533_b1 , \2549_b1 );
xor ( \2550_b0 , \2533_b0 , w_7950 );
not ( w_7950 , w_7951 );
and ( w_7951 , \2549_b1 , \2549_b0 );
or ( \2551_b1 , \2375_b1 , w_7952 );
or ( \2551_b0 , \2375_b0 , \2356_b0 );
not ( \2356_b0 , w_7953 );
and ( w_7953 , w_7952 , \2356_b1 );
or ( \2552_b1 , \2551_b1 , w_7955 );
not ( w_7955 , w_7956 );
and ( \2552_b0 , \2551_b0 , w_7957 );
and ( w_7956 ,  , w_7957 );
buf ( w_7955 , \2363_b1 );
not ( w_7955 , w_7958 );
not (  , w_7959 );
and ( w_7958 , w_7959 , \2363_b0 );
or ( \2553_b1 , \2375_b1 , w_7961 );
not ( w_7961 , w_7962 );
and ( \2553_b0 , \2375_b0 , w_7963 );
and ( w_7962 ,  , w_7963 );
buf ( w_7961 , \2356_b1 );
not ( w_7961 , w_7964 );
not (  , w_7965 );
and ( w_7964 , w_7965 , \2356_b0 );
or ( \2554_b1 , \2552_b1 , w_7967 );
not ( w_7967 , w_7968 );
and ( \2554_b0 , \2552_b0 , w_7969 );
and ( w_7968 ,  , w_7969 );
buf ( w_7967 , \2553_b1 );
not ( w_7967 , w_7970 );
not (  , w_7971 );
and ( w_7970 , w_7971 , \2553_b0 );
or ( \2555_b1 , \2550_b1 , \2554_b1 );
xor ( \2555_b0 , \2550_b0 , w_7972 );
not ( w_7972 , w_7973 );
and ( w_7973 , \2554_b1 , \2554_b0 );
buf ( \2556_b1 , \2555_b1 );
not ( \2556_b1 , w_7974 );
not ( \2556_b0 , w_7975 );
and ( w_7974 , w_7975 , \2555_b0 );
or ( \2557_b1 , \2529_b1 , \2556_b1 );
not ( \2556_b1 , w_7976 );
and ( \2557_b0 , \2529_b0 , w_7977 );
and ( w_7976 , w_7977 , \2556_b0 );
or ( \2558_b1 , \2528_b1 , \2555_b1 );
not ( \2555_b1 , w_7978 );
and ( \2558_b0 , \2528_b0 , w_7979 );
and ( w_7978 , w_7979 , \2555_b0 );
or ( \2559_b1 , \2557_b1 , w_7981 );
not ( w_7981 , w_7982 );
and ( \2559_b0 , \2557_b0 , w_7983 );
and ( w_7982 ,  , w_7983 );
buf ( w_7981 , \2558_b1 );
not ( w_7981 , w_7984 );
not (  , w_7985 );
and ( w_7984 , w_7985 , \2558_b0 );
buf ( \2560_b1 , \2559_b1 );
not ( \2560_b1 , w_7986 );
not ( \2560_b0 , w_7987 );
and ( w_7986 , w_7987 , \2559_b0 );
buf ( \2561_b1 , \2347_b1 );
not ( \2561_b1 , w_7988 );
not ( \2561_b0 , w_7989 );
and ( w_7988 , w_7989 , \2347_b0 );
buf ( \2562_b1 , \2385_b1 );
not ( \2562_b1 , w_7990 );
not ( \2562_b0 , w_7991 );
and ( w_7990 , w_7991 , \2385_b0 );
or ( \2563_b1 , \2561_b1 , w_7992 );
or ( \2563_b0 , \2561_b0 , \2562_b0 );
not ( \2562_b0 , w_7993 );
and ( w_7993 , w_7992 , \2562_b1 );
or ( \2564_b1 , \2385_b1 , w_7994 );
or ( \2564_b0 , \2385_b0 , \2347_b0 );
not ( \2347_b0 , w_7995 );
and ( w_7995 , w_7994 , \2347_b1 );
or ( \2565_b1 , \2564_b1 , w_7997 );
not ( w_7997 , w_7998 );
and ( \2565_b0 , \2564_b0 , w_7999 );
and ( w_7998 ,  , w_7999 );
buf ( w_7997 , \2377_b1 );
not ( w_7997 , w_8000 );
not (  , w_8001 );
and ( w_8000 , w_8001 , \2377_b0 );
or ( \2566_b1 , \2563_b1 , w_8003 );
not ( w_8003 , w_8004 );
and ( \2566_b0 , \2563_b0 , w_8005 );
and ( w_8004 ,  , w_8005 );
buf ( w_8003 , \2565_b1 );
not ( w_8003 , w_8006 );
not (  , w_8007 );
and ( w_8006 , w_8007 , \2565_b0 );
buf ( \2567_b1 , \2566_b1 );
not ( \2567_b1 , w_8008 );
not ( \2567_b0 , w_8009 );
and ( w_8008 , w_8009 , \2566_b0 );
or ( \2568_b1 , \2560_b1 , \2567_b1 );
not ( \2567_b1 , w_8010 );
and ( \2568_b0 , \2560_b0 , w_8011 );
and ( w_8010 , w_8011 , \2567_b0 );
or ( \2569_b1 , \2559_b1 , \2566_b1 );
not ( \2566_b1 , w_8012 );
and ( \2569_b0 , \2559_b0 , w_8013 );
and ( w_8012 , w_8013 , \2566_b0 );
or ( \2570_b1 , \2568_b1 , w_8015 );
not ( w_8015 , w_8016 );
and ( \2570_b0 , \2568_b0 , w_8017 );
and ( w_8016 ,  , w_8017 );
buf ( w_8015 , \2569_b1 );
not ( w_8015 , w_8018 );
not (  , w_8019 );
and ( w_8018 , w_8019 , \2569_b0 );
buf ( \2571_b1 , \2570_b1 );
not ( \2571_b1 , w_8020 );
not ( \2571_b0 , w_8021 );
and ( w_8020 , w_8021 , \2570_b0 );
buf ( \2572_b1 , \2315_b1 );
not ( \2572_b1 , w_8022 );
not ( \2572_b0 , w_8023 );
and ( w_8022 , w_8023 , \2315_b0 );
buf ( \2573_b1 , \2390_b1 );
not ( \2573_b1 , w_8024 );
not ( \2573_b0 , w_8025 );
and ( w_8024 , w_8025 , \2390_b0 );
or ( \2574_b1 , \2572_b1 , w_8026 );
or ( \2574_b0 , \2572_b0 , \2573_b0 );
not ( \2573_b0 , w_8027 );
and ( w_8027 , w_8026 , \2573_b1 );
or ( \2575_b1 , \2574_b1 , w_8029 );
not ( w_8029 , w_8030 );
and ( \2575_b0 , \2574_b0 , w_8031 );
and ( w_8030 ,  , w_8031 );
buf ( w_8029 , \2320_b1 );
not ( w_8029 , w_8032 );
not (  , w_8033 );
and ( w_8032 , w_8033 , \2320_b0 );
buf ( \2576_b1 , \2315_b1 );
not ( \2576_b1 , w_8034 );
not ( \2576_b0 , w_8035 );
and ( w_8034 , w_8035 , \2315_b0 );
or ( \2577_b1 , \2576_b1 , w_8037 );
not ( w_8037 , w_8038 );
and ( \2577_b0 , \2576_b0 , w_8039 );
and ( w_8038 ,  , w_8039 );
buf ( w_8037 , \2393_b1 );
not ( w_8037 , w_8040 );
not (  , w_8041 );
and ( w_8040 , w_8041 , \2393_b0 );
or ( \2578_b1 , \2575_b1 , w_8043 );
not ( w_8043 , w_8044 );
and ( \2578_b0 , \2575_b0 , w_8045 );
and ( w_8044 ,  , w_8045 );
buf ( w_8043 , \2577_b1 );
not ( w_8043 , w_8046 );
not (  , w_8047 );
and ( w_8046 , w_8047 , \2577_b0 );
or ( \2579_b1 , \2571_b1 , w_8049 );
not ( w_8049 , w_8050 );
and ( \2579_b0 , \2571_b0 , w_8051 );
and ( w_8050 ,  , w_8051 );
buf ( w_8049 , \2578_b1 );
not ( w_8049 , w_8052 );
not (  , w_8053 );
and ( w_8052 , w_8053 , \2578_b0 );
buf ( \2580_b1 , \2578_b1 );
not ( \2580_b1 , w_8054 );
not ( \2580_b0 , w_8055 );
and ( w_8054 , w_8055 , \2578_b0 );
or ( \2581_b1 , \2580_b1 , w_8057 );
not ( w_8057 , w_8058 );
and ( \2581_b0 , \2580_b0 , w_8059 );
and ( w_8058 ,  , w_8059 );
buf ( w_8057 , \2570_b1 );
not ( w_8057 , w_8060 );
not (  , w_8061 );
and ( w_8060 , w_8061 , \2570_b0 );
or ( \2582_b1 , \2579_b1 , w_8063 );
not ( w_8063 , w_8064 );
and ( \2582_b0 , \2579_b0 , w_8065 );
and ( w_8064 ,  , w_8065 );
buf ( w_8063 , \2581_b1 );
not ( w_8063 , w_8066 );
not (  , w_8067 );
and ( w_8066 , w_8067 , \2581_b0 );
buf ( \2583_b1 , \2582_b1 );
not ( \2583_b1 , w_8068 );
not ( \2583_b0 , w_8069 );
and ( w_8068 , w_8069 , \2582_b0 );
buf ( \2585_b1 , \2584_b1 );
not ( \2585_b1 , w_8070 );
not ( \2585_b0 , w_8071 );
and ( w_8070 , w_8071 , \2584_b0 );
buf ( \2586_b1 , \2273_b1 );
not ( \2586_b1 , w_8072 );
not ( \2586_b0 , w_8073 );
and ( w_8072 , w_8073 , \2273_b0 );
or ( \2587_b1 , \2270_b1 , w_8075 );
not ( w_8075 , w_8076 );
and ( \2587_b0 , \2270_b0 , w_8077 );
and ( w_8076 ,  , w_8077 );
buf ( w_8075 , \2049_b1 );
not ( w_8075 , w_8078 );
not (  , w_8079 );
and ( w_8078 , w_8079 , \2049_b0 );
buf ( \2588_b1 , \2587_b1 );
not ( \2588_b1 , w_8080 );
not ( \2588_b0 , w_8081 );
and ( w_8080 , w_8081 , \2587_b0 );
buf ( \2589_b1 , \2282_b1 );
not ( \2589_b1 , w_8082 );
not ( \2589_b0 , w_8083 );
and ( w_8082 , w_8083 , \2282_b0 );
or ( \2590_b1 , \2588_b1 , w_8084 );
or ( \2590_b0 , \2588_b0 , \2589_b0 );
not ( \2589_b0 , w_8085 );
and ( w_8085 , w_8084 , \2589_b1 );
or ( \2591_b1 , \2590_b1 , w_8087 );
not ( w_8087 , w_8088 );
and ( \2591_b0 , \2590_b0 , w_8089 );
and ( w_8088 ,  , w_8089 );
buf ( w_8087 , \2285_b1 );
not ( w_8087 , w_8090 );
not (  , w_8091 );
and ( w_8090 , w_8091 , \2285_b0 );
or ( \2592_b1 , \2586_b1 , w_8093 );
not ( w_8093 , w_8094 );
and ( \2592_b0 , \2586_b0 , w_8095 );
and ( w_8094 ,  , w_8095 );
buf ( w_8093 , \2591_b1 );
not ( w_8093 , w_8096 );
not (  , w_8097 );
and ( w_8096 , w_8097 , \2591_b0 );
buf ( \2593_b1 , \2592_b1 );
not ( \2593_b1 , w_8098 );
not ( \2593_b0 , w_8099 );
and ( w_8098 , w_8099 , \2592_b0 );
or ( \2594_b1 , \2585_b1 , w_8100 );
or ( \2594_b0 , \2585_b0 , \2593_b0 );
not ( \2593_b0 , w_8101 );
and ( w_8101 , w_8100 , \2593_b1 );
or ( \2595_b1 , \2287_b1 , w_8103 );
not ( w_8103 , w_8104 );
and ( \2595_b0 , \2287_b0 , w_8105 );
and ( w_8104 ,  , w_8105 );
buf ( w_8103 , \2403_b1 );
not ( w_8103 , w_8106 );
not (  , w_8107 );
and ( w_8106 , w_8107 , \2403_b0 );
or ( \2596_b1 , \2595_b1 , w_8109 );
not ( w_8109 , w_8110 );
and ( \2596_b0 , \2595_b0 , w_8111 );
and ( w_8110 ,  , w_8111 );
buf ( w_8109 , \2401_b1 );
not ( w_8109 , w_8112 );
not (  , w_8113 );
and ( w_8112 , w_8113 , \2401_b0 );
buf ( \2597_b1 , \2596_b1 );
not ( \2597_b1 , w_8114 );
not ( \2597_b0 , w_8115 );
and ( w_8114 , w_8115 , \2596_b0 );
or ( \2598_b1 , \2594_b1 , w_8117 );
not ( w_8117 , w_8118 );
and ( \2598_b0 , \2594_b0 , w_8119 );
and ( w_8118 ,  , w_8119 );
buf ( w_8117 , \2597_b1 );
not ( w_8117 , w_8120 );
not (  , w_8121 );
and ( w_8120 , w_8121 , \2597_b0 );
buf ( \2599_b1 , \2598_b1 );
not ( \2599_b1 , w_8122 );
not ( \2599_b0 , w_8123 );
and ( w_8122 , w_8123 , \2598_b0 );
or ( \2600_b1 , \2583_b1 , w_8124 );
or ( \2600_b0 , \2583_b0 , \2599_b0 );
not ( \2599_b0 , w_8125 );
and ( w_8125 , w_8124 , \2599_b1 );
or ( \2601_b1 , \2582_b1 , w_8126 );
or ( \2601_b0 , \2582_b0 , \2598_b0 );
not ( \2598_b0 , w_8127 );
and ( w_8127 , w_8126 , \2598_b1 );
or ( \2602_b1 , \2600_b1 , w_8129 );
not ( w_8129 , w_8130 );
and ( \2602_b0 , \2600_b0 , w_8131 );
and ( w_8130 ,  , w_8131 );
buf ( w_8129 , \2601_b1 );
not ( w_8129 , w_8132 );
not (  , w_8133 );
and ( w_8132 , w_8133 , \2601_b0 );
or ( \2603_b1 , \2602_b1 , w_8135 );
not ( w_8135 , w_8136 );
and ( \2603_b0 , \2602_b0 , w_8137 );
and ( w_8136 ,  , w_8137 );
buf ( w_8135 , \2413_b1 );
not ( w_8135 , w_8138 );
not (  , w_8139 );
and ( w_8138 , w_8139 , \2413_b0 );
buf ( \2604_b1 , \686_b1 );
not ( \2604_b1 , w_8140 );
not ( \2604_b0 , w_8141 );
and ( w_8140 , w_8141 , \686_b0 );
buf ( \2605_b1 , \648_b1 );
not ( \2605_b1 , w_8142 );
not ( \2605_b0 , w_8143 );
and ( w_8142 , w_8143 , \648_b0 );
or ( \2606_b1 , \2604_b1 , w_8144 );
or ( \2606_b0 , \2604_b0 , \2605_b0 );
not ( \2605_b0 , w_8145 );
and ( w_8145 , w_8144 , \2605_b1 );
or ( \2607_b1 , \a[14]_b1 , w_8146 );
or ( \2607_b0 , \a[14]_b0 , \b[14]_b0 );
not ( \b[14]_b0 , w_8147 );
and ( w_8147 , w_8146 , \b[14]_b1 );
or ( \2608_b1 , \2607_b1 , w_8149 );
not ( w_8149 , w_8150 );
and ( \2608_b0 , \2607_b0 , w_8151 );
and ( w_8150 ,  , w_8151 );
buf ( w_8149 , \667_b1 );
not ( w_8149 , w_8152 );
not (  , w_8153 );
and ( w_8152 , w_8153 , \667_b0 );
or ( \2609_b1 , \2606_b1 , w_8155 );
not ( w_8155 , w_8156 );
and ( \2609_b0 , \2606_b0 , w_8157 );
and ( w_8156 ,  , w_8157 );
buf ( w_8155 , \2608_b1 );
not ( w_8155 , w_8158 );
not (  , w_8159 );
and ( w_8158 , w_8159 , \2608_b0 );
or ( \2610_b1 , \b[14]_b1 , \c[14]_b1 );
not ( \c[14]_b1 , w_8160 );
and ( \2610_b0 , \b[14]_b0 , w_8161 );
and ( w_8160 , w_8161 , \c[14]_b0 );
buf ( \2611_b1 , \2610_b1 );
not ( \2611_b1 , w_8162 );
not ( \2611_b0 , w_8163 );
and ( w_8162 , w_8163 , \2610_b0 );
buf ( \2612_b1 , \922_b1 );
not ( \2612_b1 , w_8164 );
not ( \2612_b0 , w_8165 );
and ( w_8164 , w_8165 , \922_b0 );
or ( \2613_b1 , \2611_b1 , w_8166 );
or ( \2613_b0 , \2611_b0 , \2612_b0 );
not ( \2612_b0 , w_8167 );
and ( w_8167 , w_8166 , \2612_b1 );
buf ( \2614_b1 , \696_b1 );
not ( \2614_b1 , w_8168 );
not ( \2614_b0 , w_8169 );
and ( w_8168 , w_8169 , \696_b0 );
buf ( \2615_b1 , \2614_b1 );
buf ( \2615_b0 , \2614_b0 );
or ( \2616_b1 , \c[14]_b1 , \d[14]_b1 );
xor ( \2616_b0 , \c[14]_b0 , w_8170 );
not ( w_8170 , w_8171 );
and ( w_8171 , \d[14]_b1 , \d[14]_b0 );
or ( \2617_b1 , \2615_b1 , \2616_b1 );
not ( \2616_b1 , w_8172 );
and ( \2617_b0 , \2615_b0 , w_8173 );
and ( w_8172 , w_8173 , \2616_b0 );
buf ( \2618_b1 , \785_b1 );
not ( \2618_b1 , w_8174 );
not ( \2618_b0 , w_8175 );
and ( w_8174 , w_8175 , \785_b0 );
or ( \2619_b1 , \2618_b1 , w_8177 );
not ( w_8177 , w_8178 );
and ( \2619_b0 , \2618_b0 , w_8179 );
and ( w_8178 ,  , w_8179 );
buf ( w_8177 , \755_b1 );
not ( w_8177 , w_8180 );
not (  , w_8181 );
and ( w_8180 , w_8181 , \755_b0 );
buf ( \2620_b1 , \2619_b1 );
not ( \2620_b1 , w_8182 );
not ( \2620_b0 , w_8183 );
and ( w_8182 , w_8183 , \2619_b0 );
buf ( \2622_b1 , \782_b1 );
not ( \2622_b1 , w_8184 );
not ( \2622_b0 , w_8185 );
and ( w_8184 , w_8185 , \782_b0 );
or ( \2623_b1 , \776_b1 , w_8187 );
not ( w_8187 , w_8188 );
and ( \2623_b0 , \776_b0 , w_8189 );
and ( w_8188 ,  , w_8189 );
buf ( w_8187 , \759_b1 );
not ( w_8187 , w_8190 );
not (  , w_8191 );
and ( w_8190 , w_8191 , \759_b0 );
or ( \2624_b1 , \2622_b1 , w_8193 );
not ( w_8193 , w_8194 );
and ( \2624_b0 , \2622_b0 , w_8195 );
and ( w_8194 ,  , w_8195 );
buf ( w_8193 , \2623_b1 );
not ( w_8193 , w_8196 );
not (  , w_8197 );
and ( w_8196 , w_8197 , \2623_b0 );
or ( \2625_b1 , \2621_b1 , w_8199 );
not ( w_8199 , w_8200 );
and ( \2625_b0 , \2621_b0 , w_8201 );
and ( w_8200 ,  , w_8201 );
buf ( w_8199 , \2624_b1 );
not ( w_8199 , w_8202 );
not (  , w_8203 );
and ( w_8202 , w_8203 , \2624_b0 );
buf ( \2626_b1 , \2625_b1 );
not ( \2626_b1 , w_8204 );
not ( \2626_b0 , w_8205 );
and ( w_8204 , w_8205 , \2625_b0 );
or ( \2627_b1 , \2620_b1 , w_8206 );
or ( \2627_b0 , \2620_b0 , \2626_b0 );
not ( \2626_b0 , w_8207 );
and ( w_8207 , w_8206 , \2626_b1 );
or ( \2628_b1 , \2625_b1 , w_8208 );
or ( \2628_b0 , \2625_b0 , \2619_b0 );
not ( \2619_b0 , w_8209 );
and ( w_8209 , w_8208 , \2619_b1 );
or ( \2629_b1 , \2627_b1 , w_8211 );
not ( w_8211 , w_8212 );
and ( \2629_b0 , \2627_b0 , w_8213 );
and ( w_8212 ,  , w_8213 );
buf ( w_8211 , \2628_b1 );
not ( w_8211 , w_8214 );
not (  , w_8215 );
and ( w_8214 , w_8215 , \2628_b0 );
buf ( \2630_b1 , \2629_b1 );
not ( \2630_b1 , w_8216 );
not ( \2630_b0 , w_8217 );
and ( w_8216 , w_8217 , \2629_b0 );
buf ( \2631_b1 , \707_b1 );
not ( \2631_b1 , w_8218 );
not ( \2631_b0 , w_8219 );
and ( w_8218 , w_8219 , \707_b0 );
or ( \2632_b1 , \2630_b1 , w_8220 );
or ( \2632_b0 , \2630_b0 , \2631_b0 );
not ( \2631_b0 , w_8221 );
and ( w_8221 , w_8220 , \2631_b1 );
buf ( \2633_b1 , \870_b1 );
not ( \2633_b1 , w_8222 );
not ( \2633_b0 , w_8223 );
and ( w_8222 , w_8223 , \870_b0 );
or ( \2634_b1 , \2633_b1 , w_8225 );
not ( w_8225 , w_8226 );
and ( \2634_b0 , \2633_b0 , w_8227 );
and ( w_8226 ,  , w_8227 );
buf ( w_8225 , \840_b1 );
not ( w_8225 , w_8228 );
not (  , w_8229 );
and ( w_8228 , w_8229 , \840_b0 );
buf ( \2635_b1 , \2634_b1 );
not ( \2635_b1 , w_8230 );
not ( \2635_b0 , w_8231 );
and ( w_8230 , w_8231 , \2634_b0 );
buf ( \2637_b1 , \867_b1 );
not ( \2637_b1 , w_8232 );
not ( \2637_b0 , w_8233 );
and ( w_8232 , w_8233 , \867_b0 );
or ( \2638_b1 , \861_b1 , w_8235 );
not ( w_8235 , w_8236 );
and ( \2638_b0 , \861_b0 , w_8237 );
and ( w_8236 ,  , w_8237 );
buf ( w_8235 , \844_b1 );
not ( w_8235 , w_8238 );
not (  , w_8239 );
and ( w_8238 , w_8239 , \844_b0 );
or ( \2639_b1 , \2637_b1 , w_8241 );
not ( w_8241 , w_8242 );
and ( \2639_b0 , \2637_b0 , w_8243 );
and ( w_8242 ,  , w_8243 );
buf ( w_8241 , \2638_b1 );
not ( w_8241 , w_8244 );
not (  , w_8245 );
and ( w_8244 , w_8245 , \2638_b0 );
or ( \2640_b1 , \2636_b1 , w_8247 );
not ( w_8247 , w_8248 );
and ( \2640_b0 , \2636_b0 , w_8249 );
and ( w_8248 ,  , w_8249 );
buf ( w_8247 , \2639_b1 );
not ( w_8247 , w_8250 );
not (  , w_8251 );
and ( w_8250 , w_8251 , \2639_b0 );
buf ( \2641_b1 , \2640_b1 );
not ( \2641_b1 , w_8252 );
not ( \2641_b0 , w_8253 );
and ( w_8252 , w_8253 , \2640_b0 );
or ( \2642_b1 , \2635_b1 , w_8254 );
or ( \2642_b0 , \2635_b0 , \2641_b0 );
not ( \2641_b0 , w_8255 );
and ( w_8255 , w_8254 , \2641_b1 );
or ( \2643_b1 , \2640_b1 , w_8256 );
or ( \2643_b0 , \2640_b0 , \2634_b0 );
not ( \2634_b0 , w_8257 );
and ( w_8257 , w_8256 , \2634_b1 );
or ( \2644_b1 , \2642_b1 , w_8259 );
not ( w_8259 , w_8260 );
and ( \2644_b0 , \2642_b0 , w_8261 );
and ( w_8260 ,  , w_8261 );
buf ( w_8259 , \2643_b1 );
not ( w_8259 , w_8262 );
not (  , w_8263 );
and ( w_8262 , w_8263 , \2643_b0 );
or ( \2645_b1 , \880_b1 , \2644_b1 );
not ( \2644_b1 , w_8264 );
and ( \2645_b0 , \880_b0 , w_8265 );
and ( w_8264 , w_8265 , \2644_b0 );
buf ( \2646_b1 , \d[14]_b1 );
not ( \2646_b1 , w_8266 );
not ( \2646_b0 , w_8267 );
and ( w_8266 , w_8267 , \d[14]_b0 );
buf ( \2647_b1 , \894_b1 );
not ( \2647_b1 , w_8268 );
not ( \2647_b0 , w_8269 );
and ( w_8268 , w_8269 , \894_b0 );
or ( \2648_b1 , \2646_b1 , w_8270 );
or ( \2648_b0 , \2646_b0 , \2647_b0 );
not ( \2647_b0 , w_8271 );
and ( w_8271 , w_8270 , \2647_b1 );
or ( \2649_b1 , \885_b1 , \b[14]_b1 );
not ( \b[14]_b1 , w_8272 );
and ( \2649_b0 , \885_b0 , w_8273 );
and ( w_8272 , w_8273 , \b[14]_b0 );
or ( \2650_b1 , \907_b1 , \c[14]_b1 );
not ( \c[14]_b1 , w_8274 );
and ( \2650_b0 , \907_b0 , w_8275 );
and ( w_8274 , w_8275 , \c[14]_b0 );
or ( \2651_b1 , \2649_b1 , w_8277 );
not ( w_8277 , w_8278 );
and ( \2651_b0 , \2649_b0 , w_8279 );
and ( w_8278 ,  , w_8279 );
buf ( w_8277 , \2650_b1 );
not ( w_8277 , w_8280 );
not (  , w_8281 );
and ( w_8280 , w_8281 , \2650_b0 );
or ( \2652_b1 , \2648_b1 , w_8283 );
not ( w_8283 , w_8284 );
and ( \2652_b0 , \2648_b0 , w_8285 );
and ( w_8284 ,  , w_8285 );
buf ( w_8283 , \2651_b1 );
not ( w_8283 , w_8286 );
not (  , w_8287 );
and ( w_8286 , w_8287 , \2651_b0 );
or ( \2653_b1 , \2645_b1 , w_8289 );
not ( w_8289 , w_8290 );
and ( \2653_b0 , \2645_b0 , w_8291 );
and ( w_8290 ,  , w_8291 );
buf ( w_8289 , \2652_b1 );
not ( w_8289 , w_8292 );
not (  , w_8293 );
and ( w_8292 , w_8293 , \2652_b0 );
or ( \2654_b1 , \2632_b1 , w_8295 );
not ( w_8295 , w_8296 );
and ( \2654_b0 , \2632_b0 , w_8297 );
and ( w_8296 ,  , w_8297 );
buf ( w_8295 , \2653_b1 );
not ( w_8295 , w_8298 );
not (  , w_8299 );
and ( w_8298 , w_8299 , \2653_b0 );
or ( \2655_b1 , \2617_b1 , w_8301 );
not ( w_8301 , w_8302 );
and ( \2655_b0 , \2617_b0 , w_8303 );
and ( w_8302 ,  , w_8303 );
buf ( w_8301 , \2654_b1 );
not ( w_8301 , w_8304 );
not (  , w_8305 );
and ( w_8304 , w_8305 , \2654_b0 );
or ( \2656_b1 , \2613_b1 , w_8307 );
not ( w_8307 , w_8308 );
and ( \2656_b0 , \2613_b0 , w_8309 );
and ( w_8308 ,  , w_8309 );
buf ( w_8307 , \2655_b1 );
not ( w_8307 , w_8310 );
not (  , w_8311 );
and ( w_8310 , w_8311 , \2655_b0 );
or ( \2657_b1 , \2609_b1 , w_8313 );
not ( w_8313 , w_8314 );
and ( \2657_b0 , \2609_b0 , w_8315 );
and ( w_8314 ,  , w_8315 );
buf ( w_8313 , \2656_b1 );
not ( w_8313 , w_8316 );
not (  , w_8317 );
and ( w_8316 , w_8317 , \2656_b0 );
buf ( \2658_b1 , \1586_b1 );
not ( \2658_b1 , w_8318 );
not ( \2658_b0 , w_8319 );
and ( w_8318 , w_8319 , \1586_b0 );
or ( \2659_b1 , \1582_b1 , w_8321 );
not ( w_8321 , w_8322 );
and ( \2659_b0 , \1582_b0 , w_8323 );
and ( w_8322 ,  , w_8323 );
buf ( w_8321 , \1335_b1 );
not ( w_8321 , w_8324 );
not (  , w_8325 );
and ( w_8324 , w_8325 , \1335_b0 );
buf ( \2660_b1 , \2659_b1 );
not ( \2660_b1 , w_8326 );
not ( \2660_b0 , w_8327 );
and ( w_8326 , w_8327 , \2659_b0 );
or ( \2661_b1 , \2658_b1 , w_8328 );
or ( \2661_b0 , \2658_b0 , \2660_b0 );
not ( \2660_b0 , w_8329 );
and ( w_8329 , w_8328 , \2660_b1 );
or ( \2662_b1 , \a[2]_b1 , \d[13]_b1 );
xor ( \2662_b0 , \a[2]_b0 , w_8330 );
not ( w_8330 , w_8331 );
and ( w_8331 , \d[13]_b1 , \d[13]_b0 );
or ( \2663_b1 , \1335_b1 , w_8333 );
not ( w_8333 , w_8334 );
and ( \2663_b0 , \1335_b0 , w_8335 );
and ( w_8334 ,  , w_8335 );
buf ( w_8333 , \2662_b1 );
not ( w_8333 , w_8336 );
not (  , w_8337 );
and ( w_8336 , w_8337 , \2662_b0 );
or ( \2664_b1 , \2661_b1 , w_8339 );
not ( w_8339 , w_8340 );
and ( \2664_b0 , \2661_b0 , w_8341 );
and ( w_8340 ,  , w_8341 );
buf ( w_8339 , \2663_b1 );
not ( w_8339 , w_8342 );
not (  , w_8343 );
and ( w_8342 , w_8343 , \2663_b0 );
buf ( \2665_b1 , \1555_b1 );
not ( \2665_b1 , w_8344 );
not ( \2665_b0 , w_8345 );
and ( w_8344 , w_8345 , \1555_b0 );
or ( \2666_b1 , \2665_b1 , w_8347 );
not ( w_8347 , w_8348 );
and ( \2666_b0 , \2665_b0 , w_8349 );
and ( w_8348 ,  , w_8349 );
buf ( w_8347 , \1550_b1 );
not ( w_8347 , w_8350 );
not (  , w_8351 );
and ( w_8350 , w_8351 , \1550_b0 );
or ( \2667_b1 , \2664_b1 , \2666_b1 );
xor ( \2667_b0 , \2664_b0 , w_8352 );
not ( w_8352 , w_8353 );
and ( w_8353 , \2666_b1 , \2666_b0 );
buf ( \2668_b1 , \1592_b1 );
not ( \2668_b1 , w_8354 );
not ( \2668_b0 , w_8355 );
and ( w_8354 , w_8355 , \1592_b0 );
buf ( \2669_b1 , \1366_b1 );
not ( \2669_b1 , w_8356 );
not ( \2669_b0 , w_8357 );
and ( w_8356 , w_8357 , \1366_b0 );
or ( \2670_b1 , \2668_b1 , w_8358 );
or ( \2670_b0 , \2668_b0 , \2669_b0 );
not ( \2669_b0 , w_8359 );
and ( w_8359 , w_8358 , \2669_b1 );
or ( \2671_b1 , \a[4]_b1 , \d[11]_b1 );
xor ( \2671_b0 , \a[4]_b0 , w_8360 );
not ( w_8360 , w_8361 );
and ( w_8361 , \d[11]_b1 , \d[11]_b0 );
or ( \2672_b1 , \947_b1 , w_8363 );
not ( w_8363 , w_8364 );
and ( \2672_b0 , \947_b0 , w_8365 );
and ( w_8364 ,  , w_8365 );
buf ( w_8363 , \2671_b1 );
not ( w_8363 , w_8366 );
not (  , w_8367 );
and ( w_8366 , w_8367 , \2671_b0 );
or ( \2673_b1 , \2670_b1 , w_8369 );
not ( w_8369 , w_8370 );
and ( \2673_b0 , \2670_b0 , w_8371 );
and ( w_8370 ,  , w_8371 );
buf ( w_8369 , \2672_b1 );
not ( w_8369 , w_8372 );
not (  , w_8373 );
and ( w_8372 , w_8373 , \2672_b0 );
or ( \2674_b1 , \2667_b1 , \2673_b1 );
xor ( \2674_b0 , \2667_b0 , w_8374 );
not ( w_8374 , w_8375 );
and ( w_8375 , \2673_b1 , \2673_b0 );
buf ( \2675_b1 , \2674_b1 );
not ( \2675_b1 , w_8376 );
not ( \2675_b0 , w_8377 );
and ( w_8376 , w_8377 , \2674_b0 );
buf ( \2676_b1 , \2675_b1 );
not ( \2676_b1 , w_8378 );
not ( \2676_b0 , w_8379 );
and ( w_8378 , w_8379 , \2675_b0 );
buf ( \2677_b1 , \1026_b1 );
not ( \2677_b1 , w_8380 );
not ( \2677_b0 , w_8381 );
and ( w_8380 , w_8381 , \1026_b0 );
buf ( \2678_b1 , \1608_b1 );
not ( \2678_b1 , w_8382 );
not ( \2678_b0 , w_8383 );
and ( w_8382 , w_8383 , \1608_b0 );
or ( \2679_b1 , \2677_b1 , w_8384 );
or ( \2679_b0 , \2677_b0 , \2678_b0 );
not ( \2678_b0 , w_8385 );
and ( w_8385 , w_8384 , \2678_b1 );
or ( \2680_b1 , \a[6]_b1 , \d[9]_b1 );
xor ( \2680_b0 , \a[6]_b0 , w_8386 );
not ( w_8386 , w_8387 );
and ( w_8387 , \d[9]_b1 , \d[9]_b0 );
or ( \2681_b1 , \1029_b1 , w_8389 );
not ( w_8389 , w_8390 );
and ( \2681_b0 , \1029_b0 , w_8391 );
and ( w_8390 ,  , w_8391 );
buf ( w_8389 , \2680_b1 );
not ( w_8389 , w_8392 );
not (  , w_8393 );
and ( w_8392 , w_8393 , \2680_b0 );
or ( \2682_b1 , \2679_b1 , w_8395 );
not ( w_8395 , w_8396 );
and ( \2682_b0 , \2679_b0 , w_8397 );
and ( w_8396 ,  , w_8397 );
buf ( w_8395 , \2681_b1 );
not ( w_8395 , w_8398 );
not (  , w_8399 );
and ( w_8398 , w_8399 , \2681_b0 );
buf ( \2683_b1 , \1616_b1 );
not ( \2683_b1 , w_8400 );
not ( \2683_b0 , w_8401 );
and ( w_8400 , w_8401 , \1616_b0 );
buf ( \2684_b1 , \999_b1 );
not ( \2684_b1 , w_8402 );
not ( \2684_b0 , w_8403 );
and ( w_8402 , w_8403 , \999_b0 );
or ( \2685_b1 , \2683_b1 , w_8404 );
or ( \2685_b0 , \2683_b0 , \2684_b0 );
not ( \2684_b0 , w_8405 );
and ( w_8405 , w_8404 , \2684_b1 );
or ( \2686_b1 , \a[8]_b1 , \d[7]_b1 );
xor ( \2686_b0 , \a[8]_b0 , w_8406 );
not ( w_8406 , w_8407 );
and ( w_8407 , \d[7]_b1 , \d[7]_b0 );
or ( \2687_b1 , \1003_b1 , w_8409 );
not ( w_8409 , w_8410 );
and ( \2687_b0 , \1003_b0 , w_8411 );
and ( w_8410 ,  , w_8411 );
buf ( w_8409 , \2686_b1 );
not ( w_8409 , w_8412 );
not (  , w_8413 );
and ( w_8412 , w_8413 , \2686_b0 );
or ( \2688_b1 , \2685_b1 , w_8415 );
not ( w_8415 , w_8416 );
and ( \2688_b0 , \2685_b0 , w_8417 );
and ( w_8416 ,  , w_8417 );
buf ( w_8415 , \2687_b1 );
not ( w_8415 , w_8418 );
not (  , w_8419 );
and ( w_8418 , w_8419 , \2687_b0 );
or ( \2689_b1 , \2682_b1 , \2688_b1 );
xor ( \2689_b0 , \2682_b0 , w_8420 );
not ( w_8420 , w_8421 );
and ( w_8421 , \2688_b1 , \2688_b0 );
buf ( \2690_b1 , \1599_b1 );
not ( \2690_b1 , w_8422 );
not ( \2690_b0 , w_8423 );
and ( w_8422 , w_8423 , \1599_b0 );
buf ( \2691_b1 , \1312_b1 );
not ( \2691_b1 , w_8424 );
not ( \2691_b0 , w_8425 );
and ( w_8424 , w_8425 , \1312_b0 );
or ( \2692_b1 , \2690_b1 , w_8426 );
or ( \2692_b0 , \2690_b0 , \2691_b0 );
not ( \2691_b0 , w_8427 );
and ( w_8427 , w_8426 , \2691_b1 );
or ( \2693_b1 , \a[10]_b1 , \d[5]_b1 );
xor ( \2693_b0 , \a[10]_b0 , w_8428 );
not ( w_8428 , w_8429 );
and ( w_8429 , \d[5]_b1 , \d[5]_b0 );
or ( \2694_b1 , \936_b1 , w_8431 );
not ( w_8431 , w_8432 );
and ( \2694_b0 , \936_b0 , w_8433 );
and ( w_8432 ,  , w_8433 );
buf ( w_8431 , \2693_b1 );
not ( w_8431 , w_8434 );
not (  , w_8435 );
and ( w_8434 , w_8435 , \2693_b0 );
or ( \2695_b1 , \2692_b1 , w_8437 );
not ( w_8437 , w_8438 );
and ( \2695_b0 , \2692_b0 , w_8439 );
and ( w_8438 ,  , w_8439 );
buf ( w_8437 , \2694_b1 );
not ( w_8437 , w_8440 );
not (  , w_8441 );
and ( w_8440 , w_8441 , \2694_b0 );
or ( \2696_b1 , \2689_b1 , \2695_b1 );
xor ( \2696_b0 , \2689_b0 , w_8442 );
not ( w_8442 , w_8443 );
and ( w_8443 , \2695_b1 , \2695_b0 );
buf ( \2697_b1 , \2696_b1 );
not ( \2697_b1 , w_8444 );
not ( \2697_b0 , w_8445 );
and ( w_8444 , w_8445 , \2696_b0 );
buf ( \2698_b1 , \2697_b1 );
not ( \2698_b1 , w_8446 );
not ( \2698_b0 , w_8447 );
and ( w_8446 , w_8447 , \2697_b0 );
or ( \2699_b1 , \2676_b1 , w_8448 );
or ( \2699_b0 , \2676_b0 , \2698_b0 );
not ( \2698_b0 , w_8449 );
and ( w_8449 , w_8448 , \2698_b1 );
or ( \2700_b1 , \2674_b1 , w_8451 );
not ( w_8451 , w_8452 );
and ( \2700_b0 , \2674_b0 , w_8453 );
and ( w_8452 ,  , w_8453 );
buf ( w_8451 , \2696_b1 );
not ( w_8451 , w_8454 );
not (  , w_8455 );
and ( w_8454 , w_8455 , \2696_b0 );
or ( \2701_b1 , \2699_b1 , w_8457 );
not ( w_8457 , w_8458 );
and ( \2701_b0 , \2699_b0 , w_8459 );
and ( w_8458 ,  , w_8459 );
buf ( w_8457 , \2700_b1 );
not ( w_8457 , w_8460 );
not (  , w_8461 );
and ( w_8460 , w_8461 , \2700_b0 );
buf ( \2702_b1 , \1559_b1 );
not ( \2702_b1 , w_8462 );
not ( \2702_b0 , w_8463 );
and ( w_8462 , w_8463 , \1559_b0 );
buf ( \2703_b1 , \1568_b1 );
not ( \2703_b1 , w_8464 );
not ( \2703_b0 , w_8465 );
and ( w_8464 , w_8465 , \1568_b0 );
or ( \2704_b1 , \2702_b1 , w_8466 );
or ( \2704_b0 , \2702_b0 , \2703_b0 );
not ( \2703_b0 , w_8467 );
and ( w_8467 , w_8466 , \2703_b1 );
or ( \2705_b1 , \2704_b1 , w_8469 );
not ( w_8469 , w_8470 );
and ( \2705_b0 , \2704_b0 , w_8471 );
and ( w_8470 ,  , w_8471 );
buf ( w_8469 , \1563_b1 );
not ( w_8469 , w_8472 );
not (  , w_8473 );
and ( w_8472 , w_8473 , \1563_b0 );
buf ( \2706_b1 , \1559_b1 );
not ( \2706_b1 , w_8474 );
not ( \2706_b0 , w_8475 );
and ( w_8474 , w_8475 , \1559_b0 );
or ( \2707_b1 , \2706_b1 , w_8477 );
not ( w_8477 , w_8478 );
and ( \2707_b0 , \2706_b0 , w_8479 );
and ( w_8478 ,  , w_8479 );
buf ( w_8477 , \1569_b1 );
not ( w_8477 , w_8480 );
not (  , w_8481 );
and ( w_8480 , w_8481 , \1569_b0 );
or ( \2708_b1 , \2705_b1 , w_8483 );
not ( w_8483 , w_8484 );
and ( \2708_b0 , \2705_b0 , w_8485 );
and ( w_8484 ,  , w_8485 );
buf ( w_8483 , \2707_b1 );
not ( w_8483 , w_8486 );
not (  , w_8487 );
and ( w_8486 , w_8487 , \2707_b0 );
or ( \2709_b1 , \2701_b1 , w_8488 );
xor ( \2709_b0 , \2701_b0 , w_8490 );
not ( w_8490 , w_8491 );
and ( w_8491 , w_8488 , w_8489 );
buf ( w_8488 , \2708_b1 );
not ( w_8488 , w_8492 );
not ( w_8489 , w_8493 );
and ( w_8492 , w_8493 , \2708_b0 );
buf ( \2710_b1 , \2709_b1 );
not ( \2710_b1 , w_8494 );
not ( \2710_b0 , w_8495 );
and ( w_8494 , w_8495 , \2709_b0 );
or ( \2711_b1 , \1588_b1 , \1594_b1 );
xor ( \2711_b0 , \1588_b0 , w_8496 );
not ( w_8496 , w_8497 );
and ( w_8497 , \1594_b1 , \1594_b0 );
or ( \2712_b1 , \2711_b1 , \1601_b1 );
not ( \1601_b1 , w_8498 );
and ( \2712_b0 , \2711_b0 , w_8499 );
and ( w_8498 , w_8499 , \1601_b0 );
or ( \2713_b1 , \1588_b1 , \1594_b1 );
not ( \1594_b1 , w_8500 );
and ( \2713_b0 , \1588_b0 , w_8501 );
and ( w_8500 , w_8501 , \1594_b0 );
or ( \2714_b1 , \2712_b1 , w_8502 );
or ( \2714_b0 , \2712_b0 , \2713_b0 );
not ( \2713_b0 , w_8503 );
and ( w_8503 , w_8502 , \2713_b1 );
or ( \2715_b1 , \d[14]_b1 , \d[13]_b1 );
xor ( \2715_b0 , \d[14]_b0 , w_8504 );
not ( w_8504 , w_8505 );
and ( w_8505 , \d[13]_b1 , \d[13]_b0 );
or ( \2716_b1 , \2715_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_8506 );
and ( \2716_b0 , \2715_b0 , w_8507 );
and ( w_8506 , w_8507 , \a[0]_b0 );
buf ( \2717_b1 , \1012_b1 );
not ( \2717_b1 , w_8508 );
not ( \2717_b0 , w_8509 );
and ( w_8508 , w_8509 , \1012_b0 );
buf ( \2718_b1 , \1548_b1 );
not ( \2718_b1 , w_8510 );
not ( \2718_b0 , w_8511 );
and ( w_8510 , w_8511 , \1548_b0 );
or ( \2719_b1 , \2717_b1 , w_8512 );
or ( \2719_b0 , \2717_b0 , \2718_b0 );
not ( \2718_b0 , w_8513 );
and ( w_8513 , w_8512 , \2718_b1 );
or ( \2720_b1 , \d[1]_b1 , \a[14]_b1 );
xor ( \2720_b0 , \d[1]_b0 , w_8514 );
not ( w_8514 , w_8515 );
and ( w_8515 , \a[14]_b1 , \a[14]_b0 );
or ( \2721_b1 , \2720_b1 , w_8517 );
not ( w_8517 , w_8518 );
and ( \2721_b0 , \2720_b0 , w_8519 );
and ( w_8518 ,  , w_8519 );
buf ( w_8517 , \d[0]_b1 );
not ( w_8517 , w_8520 );
not (  , w_8521 );
and ( w_8520 , w_8521 , \d[0]_b0 );
or ( \2722_b1 , \2719_b1 , w_8523 );
not ( w_8523 , w_8524 );
and ( \2722_b0 , \2719_b0 , w_8525 );
and ( w_8524 ,  , w_8525 );
buf ( w_8523 , \2721_b1 );
not ( w_8523 , w_8526 );
not (  , w_8527 );
and ( w_8526 , w_8527 , \2721_b0 );
or ( \2723_b1 , \2716_b1 , \2722_b1 );
xor ( \2723_b0 , \2716_b0 , w_8528 );
not ( w_8528 , w_8529 );
and ( w_8529 , \2722_b1 , \2722_b0 );
buf ( \2724_b1 , \1627_b1 );
not ( \2724_b1 , w_8530 );
not ( \2724_b0 , w_8531 );
and ( w_8530 , w_8531 , \1627_b0 );
buf ( \2725_b1 , \962_b1 );
not ( \2725_b1 , w_8532 );
not ( \2725_b0 , w_8533 );
and ( w_8532 , w_8533 , \962_b0 );
or ( \2726_b1 , \2724_b1 , w_8534 );
or ( \2726_b0 , \2724_b0 , \2725_b0 );
not ( \2725_b0 , w_8535 );
and ( w_8535 , w_8534 , \2725_b1 );
or ( \2727_b1 , \a[12]_b1 , \d[3]_b1 );
xor ( \2727_b0 , \a[12]_b0 , w_8536 );
not ( w_8536 , w_8537 );
and ( w_8537 , \d[3]_b1 , \d[3]_b0 );
or ( \2728_b1 , \965_b1 , w_8539 );
not ( w_8539 , w_8540 );
and ( \2728_b0 , \965_b0 , w_8541 );
and ( w_8540 ,  , w_8541 );
buf ( w_8539 , \2727_b1 );
not ( w_8539 , w_8542 );
not (  , w_8543 );
and ( w_8542 , w_8543 , \2727_b0 );
or ( \2729_b1 , \2726_b1 , w_8545 );
not ( w_8545 , w_8546 );
and ( \2729_b0 , \2726_b0 , w_8547 );
and ( w_8546 ,  , w_8547 );
buf ( w_8545 , \2728_b1 );
not ( w_8545 , w_8548 );
not (  , w_8549 );
and ( w_8548 , w_8549 , \2728_b0 );
or ( \2730_b1 , \2723_b1 , \2729_b1 );
xor ( \2730_b0 , \2723_b0 , w_8550 );
not ( w_8550 , w_8551 );
and ( w_8551 , \2729_b1 , \2729_b0 );
or ( \2731_b1 , \2714_b1 , \2730_b1 );
xor ( \2731_b0 , \2714_b0 , w_8552 );
not ( w_8552 , w_8553 );
and ( w_8553 , \2730_b1 , \2730_b0 );
buf ( \2732_b1 , \1610_b1 );
not ( \2732_b1 , w_8554 );
not ( \2732_b0 , w_8555 );
and ( w_8554 , w_8555 , \1610_b0 );
or ( \2733_b1 , \1629_b1 , w_8557 );
not ( w_8557 , w_8558 );
and ( \2733_b0 , \1629_b0 , w_8559 );
and ( w_8558 ,  , w_8559 );
buf ( w_8557 , \2732_b1 );
not ( w_8557 , w_8560 );
not (  , w_8561 );
and ( w_8560 , w_8561 , \2732_b0 );
or ( \2734_b1 , \1629_b1 , w_8562 );
or ( \2734_b0 , \1629_b0 , \2732_b0 );
not ( \2732_b0 , w_8563 );
and ( w_8563 , w_8562 , \2732_b1 );
or ( \2735_b1 , \2734_b1 , w_8565 );
not ( w_8565 , w_8566 );
and ( \2735_b0 , \2734_b0 , w_8567 );
and ( w_8566 ,  , w_8567 );
buf ( w_8565 , \1618_b1 );
not ( w_8565 , w_8568 );
not (  , w_8569 );
and ( w_8568 , w_8569 , \1618_b0 );
or ( \2736_b1 , \2733_b1 , w_8571 );
not ( w_8571 , w_8572 );
and ( \2736_b0 , \2733_b0 , w_8573 );
and ( w_8572 ,  , w_8573 );
buf ( w_8571 , \2735_b1 );
not ( w_8571 , w_8574 );
not (  , w_8575 );
and ( w_8574 , w_8575 , \2735_b0 );
or ( \2737_b1 , \2731_b1 , \2736_b1 );
xor ( \2737_b0 , \2731_b0 , w_8576 );
not ( w_8576 , w_8577 );
and ( w_8577 , \2736_b1 , \2736_b0 );
buf ( \2738_b1 , \2737_b1 );
not ( \2738_b1 , w_8578 );
not ( \2738_b0 , w_8579 );
and ( w_8578 , w_8579 , \2737_b0 );
or ( \2739_b1 , \2710_b1 , \2738_b1 );
not ( \2738_b1 , w_8580 );
and ( \2739_b0 , \2710_b0 , w_8581 );
and ( w_8580 , w_8581 , \2738_b0 );
or ( \2740_b1 , \2709_b1 , \2737_b1 );
not ( \2737_b1 , w_8582 );
and ( \2740_b0 , \2709_b0 , w_8583 );
and ( w_8582 , w_8583 , \2737_b0 );
or ( \2741_b1 , \2739_b1 , w_8585 );
not ( w_8585 , w_8586 );
and ( \2741_b0 , \2739_b0 , w_8587 );
and ( w_8586 ,  , w_8587 );
buf ( w_8585 , \2740_b1 );
not ( w_8585 , w_8588 );
not (  , w_8589 );
and ( w_8588 , w_8589 , \2740_b0 );
buf ( \2742_b1 , \2741_b1 );
not ( \2742_b1 , w_8590 );
not ( \2742_b0 , w_8591 );
and ( w_8590 , w_8591 , \2741_b0 );
buf ( \2743_b1 , \1602_b1 );
not ( \2743_b1 , w_8592 );
not ( \2743_b0 , w_8593 );
and ( w_8592 , w_8593 , \1602_b0 );
buf ( \2744_b1 , \1639_b1 );
not ( \2744_b1 , w_8594 );
not ( \2744_b0 , w_8595 );
and ( w_8594 , w_8595 , \1639_b0 );
or ( \2745_b1 , \2743_b1 , w_8596 );
or ( \2745_b0 , \2743_b0 , \2744_b0 );
not ( \2744_b0 , w_8597 );
and ( w_8597 , w_8596 , \2744_b1 );
or ( \2746_b1 , \1639_b1 , w_8598 );
or ( \2746_b0 , \1639_b0 , \1602_b0 );
not ( \1602_b0 , w_8599 );
and ( w_8599 , w_8598 , \1602_b1 );
or ( \2747_b1 , \2746_b1 , w_8601 );
not ( w_8601 , w_8602 );
and ( \2747_b0 , \2746_b0 , w_8603 );
and ( w_8602 ,  , w_8603 );
buf ( w_8601 , \1631_b1 );
not ( w_8601 , w_8604 );
not (  , w_8605 );
and ( w_8604 , w_8605 , \1631_b0 );
or ( \2748_b1 , \2745_b1 , w_8607 );
not ( w_8607 , w_8608 );
and ( \2748_b0 , \2745_b0 , w_8609 );
and ( w_8608 ,  , w_8609 );
buf ( w_8607 , \2747_b1 );
not ( w_8607 , w_8610 );
not (  , w_8611 );
and ( w_8610 , w_8611 , \2747_b0 );
buf ( \2749_b1 , \2748_b1 );
not ( \2749_b1 , w_8612 );
not ( \2749_b0 , w_8613 );
and ( w_8612 , w_8613 , \2748_b0 );
or ( \2750_b1 , \2742_b1 , \2749_b1 );
not ( \2749_b1 , w_8614 );
and ( \2750_b0 , \2742_b0 , w_8615 );
and ( w_8614 , w_8615 , \2749_b0 );
or ( \2751_b1 , \2741_b1 , \2748_b1 );
not ( \2748_b1 , w_8616 );
and ( \2751_b0 , \2741_b0 , w_8617 );
and ( w_8616 , w_8617 , \2748_b0 );
or ( \2752_b1 , \2750_b1 , w_8619 );
not ( w_8619 , w_8620 );
and ( \2752_b0 , \2750_b0 , w_8621 );
and ( w_8620 ,  , w_8621 );
buf ( w_8619 , \2751_b1 );
not ( w_8619 , w_8622 );
not (  , w_8623 );
and ( w_8622 , w_8623 , \2751_b0 );
buf ( \2753_b1 , \2752_b1 );
not ( \2753_b1 , w_8624 );
not ( \2753_b0 , w_8625 );
and ( w_8624 , w_8625 , \2752_b0 );
buf ( \2754_b1 , \1570_b1 );
not ( \2754_b1 , w_8626 );
not ( \2754_b0 , w_8627 );
and ( w_8626 , w_8627 , \1570_b0 );
buf ( \2755_b1 , \1644_b1 );
not ( \2755_b1 , w_8628 );
not ( \2755_b0 , w_8629 );
and ( w_8628 , w_8629 , \1644_b0 );
or ( \2756_b1 , \2754_b1 , w_8630 );
or ( \2756_b0 , \2754_b0 , \2755_b0 );
not ( \2755_b0 , w_8631 );
and ( w_8631 , w_8630 , \2755_b1 );
or ( \2757_b1 , \2756_b1 , w_8633 );
not ( w_8633 , w_8634 );
and ( \2757_b0 , \2756_b0 , w_8635 );
and ( w_8634 ,  , w_8635 );
buf ( w_8633 , \1575_b1 );
not ( w_8633 , w_8636 );
not (  , w_8637 );
and ( w_8636 , w_8637 , \1575_b0 );
buf ( \2758_b1 , \1570_b1 );
not ( \2758_b1 , w_8638 );
not ( \2758_b0 , w_8639 );
and ( w_8638 , w_8639 , \1570_b0 );
or ( \2759_b1 , \2758_b1 , w_8641 );
not ( w_8641 , w_8642 );
and ( \2759_b0 , \2758_b0 , w_8643 );
and ( w_8642 ,  , w_8643 );
buf ( w_8641 , \1647_b1 );
not ( w_8641 , w_8644 );
not (  , w_8645 );
and ( w_8644 , w_8645 , \1647_b0 );
or ( \2760_b1 , \2757_b1 , w_8647 );
not ( w_8647 , w_8648 );
and ( \2760_b0 , \2757_b0 , w_8649 );
and ( w_8648 ,  , w_8649 );
buf ( w_8647 , \2759_b1 );
not ( w_8647 , w_8650 );
not (  , w_8651 );
and ( w_8650 , w_8651 , \2759_b0 );
or ( \2761_b1 , \2753_b1 , w_8653 );
not ( w_8653 , w_8654 );
and ( \2761_b0 , \2753_b0 , w_8655 );
and ( w_8654 ,  , w_8655 );
buf ( w_8653 , \2760_b1 );
not ( w_8653 , w_8656 );
not (  , w_8657 );
and ( w_8656 , w_8657 , \2760_b0 );
buf ( \2762_b1 , \2760_b1 );
not ( \2762_b1 , w_8658 );
not ( \2762_b0 , w_8659 );
and ( w_8658 , w_8659 , \2760_b0 );
or ( \2763_b1 , \2762_b1 , w_8661 );
not ( w_8661 , w_8662 );
and ( \2763_b0 , \2762_b0 , w_8663 );
and ( w_8662 ,  , w_8663 );
buf ( w_8661 , \2752_b1 );
not ( w_8661 , w_8664 );
not (  , w_8665 );
and ( w_8664 , w_8665 , \2752_b0 );
or ( \2764_b1 , \2761_b1 , w_8667 );
not ( w_8667 , w_8668 );
and ( \2764_b0 , \2761_b0 , w_8669 );
and ( w_8668 ,  , w_8669 );
buf ( w_8667 , \2763_b1 );
not ( w_8667 , w_8670 );
not (  , w_8671 );
and ( w_8670 , w_8671 , \2763_b0 );
buf ( \2765_b1 , \2764_b1 );
not ( \2765_b1 , w_8672 );
not ( \2765_b0 , w_8673 );
and ( w_8672 , w_8673 , \2764_b0 );
buf ( \2767_b1 , \2766_b1 );
not ( \2767_b1 , w_8674 );
not ( \2767_b0 , w_8675 );
and ( w_8674 , w_8675 , \2766_b0 );
buf ( \2768_b1 , \1530_b1 );
not ( \2768_b1 , w_8676 );
not ( \2768_b0 , w_8677 );
and ( w_8676 , w_8677 , \1530_b0 );
buf ( \2769_b1 , \1539_b1 );
not ( \2769_b1 , w_8678 );
not ( \2769_b0 , w_8679 );
and ( w_8678 , w_8679 , \1539_b0 );
or ( \2770_b1 , \1309_b1 , w_8681 );
not ( w_8681 , w_8682 );
and ( \2770_b0 , \1309_b0 , w_8683 );
and ( w_8682 ,  , w_8683 );
buf ( w_8681 , \1527_b1 );
not ( w_8681 , w_8684 );
not (  , w_8685 );
and ( w_8684 , w_8685 , \1527_b0 );
buf ( \2771_b1 , \2770_b1 );
not ( \2771_b1 , w_8686 );
not ( \2771_b0 , w_8687 );
and ( w_8686 , w_8687 , \2770_b0 );
or ( \2772_b1 , \2769_b1 , w_8688 );
or ( \2772_b0 , \2769_b0 , \2771_b0 );
not ( \2771_b0 , w_8689 );
and ( w_8689 , w_8688 , \2771_b1 );
or ( \2773_b1 , \2772_b1 , w_8691 );
not ( w_8691 , w_8692 );
and ( \2773_b0 , \2772_b0 , w_8693 );
and ( w_8692 ,  , w_8693 );
buf ( w_8691 , \1214_b1 );
not ( w_8691 , w_8694 );
not (  , w_8695 );
and ( w_8694 , w_8695 , \1214_b0 );
or ( \2774_b1 , \2768_b1 , w_8697 );
not ( w_8697 , w_8698 );
and ( \2774_b0 , \2768_b0 , w_8699 );
and ( w_8698 ,  , w_8699 );
buf ( w_8697 , \2773_b1 );
not ( w_8697 , w_8700 );
not (  , w_8701 );
and ( w_8700 , w_8701 , \2773_b0 );
buf ( \2775_b1 , \2774_b1 );
not ( \2775_b1 , w_8702 );
not ( \2775_b0 , w_8703 );
and ( w_8702 , w_8703 , \2774_b0 );
or ( \2776_b1 , \2767_b1 , w_8704 );
or ( \2776_b0 , \2767_b0 , \2775_b0 );
not ( \2775_b0 , w_8705 );
and ( w_8705 , w_8704 , \2775_b1 );
buf ( \2777_b1 , \1543_b1 );
not ( \2777_b1 , w_8706 );
not ( \2777_b0 , w_8707 );
and ( w_8706 , w_8707 , \1543_b0 );
buf ( \2778_b1 , \2777_b1 );
not ( \2778_b1 , w_8708 );
not ( \2778_b0 , w_8709 );
and ( w_8708 , w_8709 , \2777_b0 );
buf ( \2779_b1 , \1657_b1 );
not ( \2779_b1 , w_8710 );
not ( \2779_b0 , w_8711 );
and ( w_8710 , w_8711 , \1657_b0 );
or ( \2780_b1 , \2778_b1 , w_8712 );
or ( \2780_b0 , \2778_b0 , \2779_b0 );
not ( \2779_b0 , w_8713 );
and ( w_8713 , w_8712 , \2779_b1 );
or ( \2781_b1 , \2780_b1 , w_8715 );
not ( w_8715 , w_8716 );
and ( \2781_b0 , \2780_b0 , w_8717 );
and ( w_8716 ,  , w_8717 );
buf ( w_8715 , \1655_b1 );
not ( w_8715 , w_8718 );
not (  , w_8719 );
and ( w_8718 , w_8719 , \1655_b0 );
buf ( \2782_b1 , \2781_b1 );
not ( \2782_b1 , w_8720 );
not ( \2782_b0 , w_8721 );
and ( w_8720 , w_8721 , \2781_b0 );
or ( \2783_b1 , \2776_b1 , w_8723 );
not ( w_8723 , w_8724 );
and ( \2783_b0 , \2776_b0 , w_8725 );
and ( w_8724 ,  , w_8725 );
buf ( w_8723 , \2782_b1 );
not ( w_8723 , w_8726 );
not (  , w_8727 );
and ( w_8726 , w_8727 , \2782_b0 );
buf ( \2784_b1 , \2783_b1 );
not ( \2784_b1 , w_8728 );
not ( \2784_b0 , w_8729 );
and ( w_8728 , w_8729 , \2783_b0 );
or ( \2785_b1 , \2765_b1 , w_8730 );
or ( \2785_b0 , \2765_b0 , \2784_b0 );
not ( \2784_b0 , w_8731 );
and ( w_8731 , w_8730 , \2784_b1 );
or ( \2786_b1 , \2764_b1 , w_8732 );
or ( \2786_b0 , \2764_b0 , \2783_b0 );
not ( \2783_b0 , w_8733 );
and ( w_8733 , w_8732 , \2783_b1 );
or ( \2787_b1 , \2785_b1 , w_8735 );
not ( w_8735 , w_8736 );
and ( \2787_b0 , \2785_b0 , w_8737 );
and ( w_8736 ,  , w_8737 );
buf ( w_8735 , \2786_b1 );
not ( w_8735 , w_8738 );
not (  , w_8739 );
and ( w_8738 , w_8739 , \2786_b0 );
or ( \2788_b1 , \2787_b1 , w_8741 );
not ( w_8741 , w_8742 );
and ( \2788_b0 , \2787_b0 , w_8743 );
and ( w_8742 ,  , w_8743 );
buf ( w_8741 , \1668_b1 );
not ( w_8741 , w_8744 );
not (  , w_8745 );
and ( w_8744 , w_8745 , \1668_b0 );
or ( \2789_b1 , \2475_b1 , w_8747 );
not ( w_8747 , w_8748 );
and ( \2789_b0 , \2475_b0 , w_8749 );
and ( w_8748 ,  , w_8749 );
buf ( w_8747 , \a[14]_b1 );
not ( w_8747 , w_8750 );
not (  , w_8751 );
and ( w_8750 , w_8751 , \a[14]_b0 );
buf ( \2791_b1 , \667_b1 );
buf ( \2791_b0 , \667_b0 );
or ( \2792_b1 , \a[11]_b1 , w_8752 );
or ( \2792_b0 , \a[11]_b0 , \b[11]_b0 );
not ( \b[11]_b0 , w_8753 );
and ( w_8753 , w_8752 , \b[11]_b1 );
or ( \2793_b1 , \2791_b1 , \2792_b1 );
not ( \2792_b1 , w_8754 );
and ( \2793_b0 , \2791_b0 , w_8755 );
and ( w_8754 , w_8755 , \2792_b0 );
or ( \2794_b1 , \b[11]_b1 , \c[11]_b1 );
not ( \c[11]_b1 , w_8756 );
and ( \2794_b0 , \b[11]_b0 , w_8757 );
and ( w_8756 , w_8757 , \c[11]_b0 );
buf ( \2795_b1 , \2794_b1 );
not ( \2795_b1 , w_8758 );
not ( \2795_b0 , w_8759 );
and ( w_8758 , w_8759 , \2794_b0 );
buf ( \2796_b1 , \922_b1 );
not ( \2796_b1 , w_8760 );
not ( \2796_b0 , w_8761 );
and ( w_8760 , w_8761 , \922_b0 );
or ( \2797_b1 , \2795_b1 , w_8762 );
or ( \2797_b0 , \2795_b0 , \2796_b0 );
not ( \2796_b0 , w_8763 );
and ( w_8763 , w_8762 , \2796_b1 );
or ( \2798_b1 , \c[11]_b1 , \d[11]_b1 );
xor ( \2798_b0 , \c[11]_b0 , w_8764 );
not ( w_8764 , w_8765 );
and ( w_8765 , \d[11]_b1 , \d[11]_b0 );
or ( \2799_b1 , \2615_b1 , \2798_b1 );
not ( \2798_b1 , w_8766 );
and ( \2799_b0 , \2615_b0 , w_8767 );
and ( w_8766 , w_8767 , \2798_b0 );
or ( \2800_b1 , \748_b1 , w_8769 );
not ( w_8769 , w_8770 );
and ( \2800_b0 , \748_b0 , w_8771 );
and ( w_8770 ,  , w_8771 );
buf ( w_8769 , \774_b1 );
not ( w_8769 , w_8772 );
not (  , w_8773 );
and ( w_8772 , w_8773 , \774_b0 );
buf ( \2801_b1 , \2800_b1 );
not ( \2801_b1 , w_8774 );
not ( \2801_b0 , w_8775 );
and ( w_8774 , w_8775 , \2800_b0 );
buf ( \2802_b1 , \749_b1 );
not ( \2802_b1 , w_8776 );
not ( \2802_b0 , w_8777 );
and ( w_8776 , w_8777 , \749_b0 );
buf ( \2804_b1 , \2802_b1 );
not ( \2804_b1 , w_8778 );
not ( \2804_b0 , w_8779 );
and ( w_8778 , w_8779 , \2802_b0 );
buf ( \2805_b1 , \766_b1 );
not ( \2805_b1 , w_8780 );
not ( \2805_b0 , w_8781 );
and ( w_8780 , w_8781 , \766_b0 );
or ( \2806_b1 , \2804_b1 , w_8782 );
or ( \2806_b0 , \2804_b0 , \2805_b0 );
not ( \2805_b0 , w_8783 );
and ( w_8783 , w_8782 , \2805_b1 );
or ( \2807_b1 , \2806_b1 , w_8785 );
not ( w_8785 , w_8786 );
and ( \2807_b0 , \2806_b0 , w_8787 );
and ( w_8786 ,  , w_8787 );
buf ( w_8785 , \771_b1 );
not ( w_8785 , w_8788 );
not (  , w_8789 );
and ( w_8788 , w_8789 , \771_b0 );
or ( \2808_b1 , \2803_b1 , w_8791 );
not ( w_8791 , w_8792 );
and ( \2808_b0 , \2803_b0 , w_8793 );
and ( w_8792 ,  , w_8793 );
buf ( w_8791 , \2807_b1 );
not ( w_8791 , w_8794 );
not (  , w_8795 );
and ( w_8794 , w_8795 , \2807_b0 );
buf ( \2809_b1 , \2808_b1 );
not ( \2809_b1 , w_8796 );
not ( \2809_b0 , w_8797 );
and ( w_8796 , w_8797 , \2808_b0 );
or ( \2810_b1 , \2801_b1 , w_8798 );
or ( \2810_b0 , \2801_b0 , \2809_b0 );
not ( \2809_b0 , w_8799 );
and ( w_8799 , w_8798 , \2809_b1 );
or ( \2811_b1 , \2808_b1 , w_8800 );
or ( \2811_b0 , \2808_b0 , \2800_b0 );
not ( \2800_b0 , w_8801 );
and ( w_8801 , w_8800 , \2800_b1 );
or ( \2812_b1 , \2810_b1 , w_8803 );
not ( w_8803 , w_8804 );
and ( \2812_b0 , \2810_b0 , w_8805 );
and ( w_8804 ,  , w_8805 );
buf ( w_8803 , \2811_b1 );
not ( w_8803 , w_8806 );
not (  , w_8807 );
and ( w_8806 , w_8807 , \2811_b0 );
buf ( \2813_b1 , \2812_b1 );
not ( \2813_b1 , w_8808 );
not ( \2813_b0 , w_8809 );
and ( w_8808 , w_8809 , \2812_b0 );
buf ( \2814_b1 , \707_b1 );
not ( \2814_b1 , w_8810 );
not ( \2814_b0 , w_8811 );
and ( w_8810 , w_8811 , \707_b0 );
or ( \2815_b1 , \2813_b1 , w_8812 );
or ( \2815_b0 , \2813_b0 , \2814_b0 );
not ( \2814_b0 , w_8813 );
and ( w_8813 , w_8812 , \2814_b1 );
or ( \2816_b1 , \833_b1 , w_8815 );
not ( w_8815 , w_8816 );
and ( \2816_b0 , \833_b0 , w_8817 );
and ( w_8816 ,  , w_8817 );
buf ( w_8815 , \859_b1 );
not ( w_8815 , w_8818 );
not (  , w_8819 );
and ( w_8818 , w_8819 , \859_b0 );
buf ( \2817_b1 , \2816_b1 );
not ( \2817_b1 , w_8820 );
not ( \2817_b0 , w_8821 );
and ( w_8820 , w_8821 , \2816_b0 );
buf ( \2818_b1 , \834_b1 );
not ( \2818_b1 , w_8822 );
not ( \2818_b0 , w_8823 );
and ( w_8822 , w_8823 , \834_b0 );
buf ( \2820_b1 , \2818_b1 );
not ( \2820_b1 , w_8824 );
not ( \2820_b0 , w_8825 );
and ( w_8824 , w_8825 , \2818_b0 );
buf ( \2821_b1 , \851_b1 );
not ( \2821_b1 , w_8826 );
not ( \2821_b0 , w_8827 );
and ( w_8826 , w_8827 , \851_b0 );
or ( \2822_b1 , \2820_b1 , w_8828 );
or ( \2822_b0 , \2820_b0 , \2821_b0 );
not ( \2821_b0 , w_8829 );
and ( w_8829 , w_8828 , \2821_b1 );
or ( \2823_b1 , \2822_b1 , w_8831 );
not ( w_8831 , w_8832 );
and ( \2823_b0 , \2822_b0 , w_8833 );
and ( w_8832 ,  , w_8833 );
buf ( w_8831 , \856_b1 );
not ( w_8831 , w_8834 );
not (  , w_8835 );
and ( w_8834 , w_8835 , \856_b0 );
or ( \2824_b1 , \2819_b1 , w_8837 );
not ( w_8837 , w_8838 );
and ( \2824_b0 , \2819_b0 , w_8839 );
and ( w_8838 ,  , w_8839 );
buf ( w_8837 , \2823_b1 );
not ( w_8837 , w_8840 );
not (  , w_8841 );
and ( w_8840 , w_8841 , \2823_b0 );
buf ( \2825_b1 , \2824_b1 );
not ( \2825_b1 , w_8842 );
not ( \2825_b0 , w_8843 );
and ( w_8842 , w_8843 , \2824_b0 );
or ( \2826_b1 , \2817_b1 , w_8844 );
or ( \2826_b0 , \2817_b0 , \2825_b0 );
not ( \2825_b0 , w_8845 );
and ( w_8845 , w_8844 , \2825_b1 );
or ( \2827_b1 , \2824_b1 , w_8846 );
or ( \2827_b0 , \2824_b0 , \2816_b0 );
not ( \2816_b0 , w_8847 );
and ( w_8847 , w_8846 , \2816_b1 );
or ( \2828_b1 , \2826_b1 , w_8849 );
not ( w_8849 , w_8850 );
and ( \2828_b0 , \2826_b0 , w_8851 );
and ( w_8850 ,  , w_8851 );
buf ( w_8849 , \2827_b1 );
not ( w_8849 , w_8852 );
not (  , w_8853 );
and ( w_8852 , w_8853 , \2827_b0 );
or ( \2829_b1 , \880_b1 , \2828_b1 );
not ( \2828_b1 , w_8854 );
and ( \2829_b0 , \880_b0 , w_8855 );
and ( w_8854 , w_8855 , \2828_b0 );
buf ( \2830_b1 , \d[11]_b1 );
not ( \2830_b1 , w_8856 );
not ( \2830_b0 , w_8857 );
and ( w_8856 , w_8857 , \d[11]_b0 );
buf ( \2831_b1 , \894_b1 );
not ( \2831_b1 , w_8858 );
not ( \2831_b0 , w_8859 );
and ( w_8858 , w_8859 , \894_b0 );
or ( \2832_b1 , \2830_b1 , w_8860 );
or ( \2832_b0 , \2830_b0 , \2831_b0 );
not ( \2831_b0 , w_8861 );
and ( w_8861 , w_8860 , \2831_b1 );
or ( \2833_b1 , \885_b1 , \b[11]_b1 );
not ( \b[11]_b1 , w_8862 );
and ( \2833_b0 , \885_b0 , w_8863 );
and ( w_8862 , w_8863 , \b[11]_b0 );
or ( \2834_b1 , \909_b1 , \c[11]_b1 );
not ( \c[11]_b1 , w_8864 );
and ( \2834_b0 , \909_b0 , w_8865 );
and ( w_8864 , w_8865 , \c[11]_b0 );
or ( \2835_b1 , \2833_b1 , w_8867 );
not ( w_8867 , w_8868 );
and ( \2835_b0 , \2833_b0 , w_8869 );
and ( w_8868 ,  , w_8869 );
buf ( w_8867 , \2834_b1 );
not ( w_8867 , w_8870 );
not (  , w_8871 );
and ( w_8870 , w_8871 , \2834_b0 );
or ( \2836_b1 , \2832_b1 , w_8873 );
not ( w_8873 , w_8874 );
and ( \2836_b0 , \2832_b0 , w_8875 );
and ( w_8874 ,  , w_8875 );
buf ( w_8873 , \2835_b1 );
not ( w_8873 , w_8876 );
not (  , w_8877 );
and ( w_8876 , w_8877 , \2835_b0 );
or ( \2837_b1 , \2829_b1 , w_8879 );
not ( w_8879 , w_8880 );
and ( \2837_b0 , \2829_b0 , w_8881 );
and ( w_8880 ,  , w_8881 );
buf ( w_8879 , \2836_b1 );
not ( w_8879 , w_8882 );
not (  , w_8883 );
and ( w_8882 , w_8883 , \2836_b0 );
or ( \2838_b1 , \2815_b1 , w_8885 );
not ( w_8885 , w_8886 );
and ( \2838_b0 , \2815_b0 , w_8887 );
and ( w_8886 ,  , w_8887 );
buf ( w_8885 , \2837_b1 );
not ( w_8885 , w_8888 );
not (  , w_8889 );
and ( w_8888 , w_8889 , \2837_b0 );
or ( \2839_b1 , \2799_b1 , w_8891 );
not ( w_8891 , w_8892 );
and ( \2839_b0 , \2799_b0 , w_8893 );
and ( w_8892 ,  , w_8893 );
buf ( w_8891 , \2838_b1 );
not ( w_8891 , w_8894 );
not (  , w_8895 );
and ( w_8894 , w_8895 , \2838_b0 );
or ( \2840_b1 , \2797_b1 , w_8897 );
not ( w_8897 , w_8898 );
and ( \2840_b0 , \2797_b0 , w_8899 );
and ( w_8898 ,  , w_8899 );
buf ( w_8897 , \2839_b1 );
not ( w_8897 , w_8900 );
not (  , w_8901 );
and ( w_8900 , w_8901 , \2839_b0 );
or ( \2841_b1 , \2793_b1 , w_8903 );
not ( w_8903 , w_8904 );
and ( \2841_b0 , \2793_b0 , w_8905 );
and ( w_8904 ,  , w_8905 );
buf ( w_8903 , \2840_b1 );
not ( w_8903 , w_8906 );
not (  , w_8907 );
and ( w_8906 , w_8907 , \2840_b0 );
or ( \2842_b1 , \a[11]_b1 , w_8908 );
or ( \2842_b0 , \a[11]_b0 , \d[11]_b0 );
not ( \d[11]_b0 , w_8909 );
and ( w_8909 , w_8908 , \d[11]_b1 );
buf ( \2843_b1 , \648_b1 );
buf ( \2843_b0 , \648_b0 );
or ( \2844_b1 , \2842_b1 , \2843_b1 );
not ( \2843_b1 , w_8910 );
and ( \2844_b0 , \2842_b0 , w_8911 );
and ( w_8910 , w_8911 , \2843_b0 );
buf ( \2845_b1 , \1537_b1 );
not ( \2845_b1 , w_8912 );
not ( \2845_b0 , w_8913 );
and ( w_8912 , w_8913 , \1537_b0 );
or ( \2846_b1 , \2845_b1 , w_8915 );
not ( w_8915 , w_8916 );
and ( \2846_b0 , \2845_b0 , w_8917 );
and ( w_8916 ,  , w_8917 );
buf ( w_8915 , \2770_b1 );
not ( w_8915 , w_8918 );
not (  , w_8919 );
and ( w_8918 , w_8919 , \2770_b0 );
buf ( \2847_b1 , \2846_b1 );
not ( \2847_b1 , w_8920 );
not ( \2847_b0 , w_8921 );
and ( w_8920 , w_8921 , \2846_b0 );
buf ( \2848_b1 , \1214_b1 );
not ( \2848_b1 , w_8922 );
not ( \2848_b0 , w_8923 );
and ( w_8922 , w_8923 , \1214_b0 );
or ( \2849_b1 , \2847_b1 , w_8924 );
or ( \2849_b0 , \2847_b0 , \2848_b0 );
not ( \2848_b0 , w_8925 );
and ( w_8925 , w_8924 , \2848_b1 );
buf ( \2850_b1 , \1538_b1 );
not ( \2850_b1 , w_8926 );
not ( \2850_b0 , w_8927 );
and ( w_8926 , w_8927 , \1538_b0 );
or ( \2851_b1 , \2849_b1 , w_8929 );
not ( w_8929 , w_8930 );
and ( \2851_b0 , \2849_b0 , w_8931 );
and ( w_8930 ,  , w_8931 );
buf ( w_8929 , \2850_b1 );
not ( w_8929 , w_8932 );
not (  , w_8933 );
and ( w_8932 , w_8933 , \2850_b0 );
buf ( \2852_b1 , \1530_b1 );
not ( \2852_b1 , w_8934 );
not ( \2852_b0 , w_8935 );
and ( w_8934 , w_8935 , \1530_b0 );
or ( \2853_b1 , \2852_b1 , w_8937 );
not ( w_8937 , w_8938 );
and ( \2853_b0 , \2852_b0 , w_8939 );
and ( w_8938 ,  , w_8939 );
buf ( w_8937 , \1541_b1 );
not ( w_8937 , w_8940 );
not (  , w_8941 );
and ( w_8940 , w_8941 , \1541_b0 );
or ( \2854_b1 , \2851_b1 , \2853_b1 );
xor ( \2854_b0 , \2851_b0 , w_8942 );
not ( w_8942 , w_8943 );
and ( w_8943 , \2853_b1 , \2853_b0 );
or ( \2855_b1 , \2854_b1 , w_8945 );
not ( w_8945 , w_8946 );
and ( \2855_b0 , \2854_b0 , w_8947 );
and ( w_8946 ,  , w_8947 );
buf ( w_8945 , \1667_b1 );
not ( w_8945 , w_8948 );
not (  , w_8949 );
and ( w_8948 , w_8949 , \1667_b0 );
or ( \2856_b1 , \2844_b1 , w_8951 );
not ( w_8951 , w_8952 );
and ( \2856_b0 , \2844_b0 , w_8953 );
and ( w_8952 ,  , w_8953 );
buf ( w_8951 , \2855_b1 );
not ( w_8951 , w_8954 );
not (  , w_8955 );
and ( w_8954 , w_8955 , \2855_b0 );
or ( \2857_b1 , \2466_b1 , w_8957 );
not ( w_8957 , w_8958 );
and ( \2857_b0 , \2466_b0 , w_8959 );
and ( w_8958 ,  , w_8959 );
buf ( w_8957 , \2474_b1 );
not ( w_8957 , w_8960 );
not (  , w_8961 );
and ( w_8960 , w_8961 , \2474_b0 );
buf ( \2858_b1 , \2857_b1 );
not ( \2858_b1 , w_8962 );
not ( \2858_b0 , w_8963 );
and ( w_8962 , w_8963 , \2857_b0 );
buf ( \2859_b1 , \2858_b1 );
buf ( \2859_b0 , \2858_b0 );
or ( \2860_b1 , \2859_b1 , w_8965 );
not ( w_8965 , w_8966 );
and ( \2860_b0 , \2859_b0 , w_8967 );
and ( w_8966 ,  , w_8967 );
buf ( w_8965 , \a[11]_b1 );
not ( w_8965 , w_8968 );
not (  , w_8969 );
and ( w_8968 , w_8969 , \a[11]_b0 );
buf ( \2861_b1 , \2285_b1 );
not ( \2861_b1 , w_8970 );
not ( \2861_b0 , w_8971 );
and ( w_8970 , w_8971 , \2285_b0 );
buf ( \2862_b1 , \2280_b1 );
not ( \2862_b1 , w_8972 );
not ( \2862_b0 , w_8973 );
and ( w_8972 , w_8973 , \2280_b0 );
or ( \2863_b1 , \2862_b1 , w_8975 );
not ( w_8975 , w_8976 );
and ( \2863_b0 , \2862_b0 , w_8977 );
and ( w_8976 ,  , w_8977 );
buf ( w_8975 , \2587_b1 );
not ( w_8975 , w_8978 );
not (  , w_8979 );
and ( w_8978 , w_8979 , \2587_b0 );
buf ( \2864_b1 , \2863_b1 );
not ( \2864_b1 , w_8980 );
not ( \2864_b0 , w_8981 );
and ( w_8980 , w_8981 , \2863_b0 );
or ( \2865_b1 , \2861_b1 , w_8982 );
or ( \2865_b0 , \2861_b0 , \2864_b0 );
not ( \2864_b0 , w_8983 );
and ( w_8983 , w_8982 , \2864_b1 );
buf ( \2866_b1 , \2281_b1 );
not ( \2866_b1 , w_8984 );
not ( \2866_b0 , w_8985 );
and ( w_8984 , w_8985 , \2281_b0 );
or ( \2867_b1 , \2865_b1 , w_8987 );
not ( w_8987 , w_8988 );
and ( \2867_b0 , \2865_b0 , w_8989 );
and ( w_8988 ,  , w_8989 );
buf ( w_8987 , \2866_b1 );
not ( w_8987 , w_8990 );
not (  , w_8991 );
and ( w_8990 , w_8991 , \2866_b0 );
buf ( \2868_b1 , \2273_b1 );
not ( \2868_b1 , w_8992 );
not ( \2868_b0 , w_8993 );
and ( w_8992 , w_8993 , \2273_b0 );
or ( \2869_b1 , \2868_b1 , w_8995 );
not ( w_8995 , w_8996 );
and ( \2869_b0 , \2868_b0 , w_8997 );
and ( w_8996 ,  , w_8997 );
buf ( w_8995 , \2284_b1 );
not ( w_8995 , w_8998 );
not (  , w_8999 );
and ( w_8998 , w_8999 , \2284_b0 );
buf ( \2870_b1 , \2869_b1 );
not ( \2870_b1 , w_9000 );
not ( \2870_b0 , w_9001 );
and ( w_9000 , w_9001 , \2869_b0 );
or ( \2871_b1 , \2867_b1 , \2870_b1 );
not ( \2870_b1 , w_9002 );
and ( \2871_b0 , \2867_b0 , w_9003 );
and ( w_9002 , w_9003 , \2870_b0 );
buf ( \2872_b1 , \2867_b1 );
not ( \2872_b1 , w_9004 );
not ( \2872_b0 , w_9005 );
and ( w_9004 , w_9005 , \2867_b0 );
or ( \2873_b1 , \2872_b1 , \2869_b1 );
not ( \2869_b1 , w_9006 );
and ( \2873_b0 , \2872_b0 , w_9007 );
and ( w_9006 , w_9007 , \2869_b0 );
or ( \2874_b1 , \2871_b1 , w_9009 );
not ( w_9009 , w_9010 );
and ( \2874_b0 , \2871_b0 , w_9011 );
and ( w_9010 ,  , w_9011 );
buf ( w_9009 , \2873_b1 );
not ( w_9009 , w_9012 );
not (  , w_9013 );
and ( w_9012 , w_9013 , \2873_b0 );
or ( \2875_b1 , \2874_b1 , w_9015 );
not ( w_9015 , w_9016 );
and ( \2875_b0 , \2874_b0 , w_9017 );
and ( w_9016 ,  , w_9017 );
buf ( w_9015 , \2413_b1 );
not ( w_9015 , w_9018 );
not (  , w_9019 );
and ( w_9018 , w_9019 , \2413_b0 );
buf ( \2877_b1 , \666_b1 );
not ( \2877_b1 , w_9020 );
not ( \2877_b0 , w_9021 );
and ( w_9020 , w_9021 , \666_b0 );
buf ( \2878_b1 , \2877_b1 );
not ( \2878_b1 , w_9022 );
not ( \2878_b0 , w_9023 );
and ( w_9022 , w_9023 , \2877_b0 );
or ( \2879_b1 , \a[3]_b1 , w_9025 );
not ( w_9025 , w_9026 );
and ( \2879_b0 , \a[3]_b0 , w_9027 );
and ( w_9026 ,  , w_9027 );
buf ( w_9025 , \b[3]_b1 );
not ( w_9025 , w_9028 );
not (  , w_9029 );
and ( w_9028 , w_9029 , \b[3]_b0 );
buf ( \2880_b1 , \2879_b1 );
not ( \2880_b1 , w_9030 );
not ( \2880_b0 , w_9031 );
and ( w_9030 , w_9031 , \2879_b0 );
or ( \2881_b1 , \2878_b1 , \2880_b1 );
not ( \2880_b1 , w_9032 );
and ( \2881_b0 , \2878_b0 , w_9033 );
and ( w_9032 , w_9033 , \2880_b0 );
buf ( \2882_b1 , \674_b1 );
not ( \2882_b1 , w_9034 );
not ( \2882_b0 , w_9035 );
and ( w_9034 , w_9035 , \674_b0 );
or ( \2883_b1 , \648_b1 , \2882_b1 );
not ( \2882_b1 , w_9036 );
and ( \2883_b0 , \648_b0 , w_9037 );
and ( w_9036 , w_9037 , \2882_b0 );
or ( \2884_b1 , \2881_b1 , w_9039 );
not ( w_9039 , w_9040 );
and ( \2884_b0 , \2881_b0 , w_9041 );
and ( w_9040 ,  , w_9041 );
buf ( w_9039 , \2883_b1 );
not ( w_9039 , w_9042 );
not (  , w_9043 );
and ( w_9042 , w_9043 , \2883_b0 );
or ( \2885_b1 , \2858_b1 , w_9045 );
not ( w_9045 , w_9046 );
and ( \2885_b0 , \2858_b0 , w_9047 );
and ( w_9046 ,  , w_9047 );
buf ( w_9045 , \a[3]_b1 );
not ( w_9045 , w_9048 );
not (  , w_9049 );
and ( w_9048 , w_9049 , \a[3]_b0 );
buf ( \2886_b1 , \921_b1 );
not ( \2886_b1 , w_9050 );
not ( \2886_b0 , w_9051 );
and ( w_9050 , w_9051 , \921_b0 );
buf ( \2887_b1 , \2886_b1 );
not ( \2887_b1 , w_9052 );
not ( \2887_b0 , w_9053 );
and ( w_9052 , w_9053 , \2886_b0 );
or ( \2888_b1 , \b[3]_b1 , \c[3]_b1 );
not ( \c[3]_b1 , w_9054 );
and ( \2888_b0 , \b[3]_b0 , w_9055 );
and ( w_9054 , w_9055 , \c[3]_b0 );
or ( \2889_b1 , \2887_b1 , \2888_b1 );
not ( \2888_b1 , w_9056 );
and ( \2889_b0 , \2887_b0 , w_9057 );
and ( w_9056 , w_9057 , \2888_b0 );
or ( \2890_b1 , \c[3]_b1 , \d[3]_b1 );
xor ( \2890_b0 , \c[3]_b0 , w_9058 );
not ( w_9058 , w_9059 );
and ( w_9059 , \d[3]_b1 , \d[3]_b0 );
buf ( \2891_b1 , \2890_b1 );
not ( \2891_b1 , w_9060 );
not ( \2891_b0 , w_9061 );
and ( w_9060 , w_9061 , \2890_b0 );
buf ( \2892_b1 , \697_b1 );
not ( \2892_b1 , w_9062 );
not ( \2892_b0 , w_9063 );
and ( w_9062 , w_9063 , \697_b0 );
or ( \2893_b1 , \2891_b1 , w_9064 );
or ( \2893_b0 , \2891_b0 , \2892_b0 );
not ( \2892_b0 , w_9065 );
and ( w_9065 , w_9064 , \2892_b1 );
buf ( \2894_b1 , \2225_b1 );
not ( \2894_b1 , w_9066 );
not ( \2894_b0 , w_9067 );
and ( w_9066 , w_9067 , \2225_b0 );
or ( \2895_b1 , \2228_b1 , w_9069 );
not ( w_9069 , w_9070 );
and ( \2895_b0 , \2228_b0 , w_9071 );
and ( w_9070 ,  , w_9071 );
buf ( w_9069 , \2204_b1 );
not ( w_9069 , w_9072 );
not (  , w_9073 );
and ( w_9072 , w_9073 , \2204_b0 );
buf ( \2896_b1 , \2895_b1 );
not ( \2896_b1 , w_9074 );
not ( \2896_b0 , w_9075 );
and ( w_9074 , w_9075 , \2895_b0 );
or ( \2897_b1 , \2894_b1 , w_9076 );
or ( \2897_b0 , \2894_b0 , \2896_b0 );
not ( \2896_b0 , w_9077 );
and ( w_9077 , w_9076 , \2896_b1 );
or ( \2898_b1 , \2895_b1 , w_9078 );
or ( \2898_b0 , \2895_b0 , \2225_b0 );
not ( \2225_b0 , w_9079 );
and ( w_9079 , w_9078 , \2225_b1 );
or ( \2899_b1 , \2897_b1 , w_9081 );
not ( w_9081 , w_9082 );
and ( \2899_b0 , \2897_b0 , w_9083 );
and ( w_9082 ,  , w_9083 );
buf ( w_9081 , \2898_b1 );
not ( w_9081 , w_9084 );
not (  , w_9085 );
and ( w_9084 , w_9085 , \2898_b0 );
or ( \2900_b1 , \2413_b1 , \2899_b1 );
not ( \2899_b1 , w_9086 );
and ( \2900_b0 , \2413_b0 , w_9087 );
and ( w_9086 , w_9087 , \2899_b0 );
buf ( \2901_b1 , \1507_b1 );
not ( \2901_b1 , w_9088 );
not ( \2901_b0 , w_9089 );
and ( w_9088 , w_9089 , \1507_b0 );
or ( \2902_b1 , \1487_b1 , w_9091 );
not ( w_9091 , w_9092 );
and ( \2902_b0 , \1487_b0 , w_9093 );
and ( w_9092 ,  , w_9093 );
buf ( w_9091 , \1488_b1 );
not ( w_9091 , w_9094 );
not (  , w_9095 );
and ( w_9094 , w_9095 , \1488_b0 );
buf ( \2903_b1 , \2902_b1 );
not ( \2903_b1 , w_9096 );
not ( \2903_b0 , w_9097 );
and ( w_9096 , w_9097 , \2902_b0 );
or ( \2904_b1 , \2901_b1 , w_9098 );
or ( \2904_b0 , \2901_b0 , \2903_b0 );
not ( \2903_b0 , w_9099 );
and ( w_9099 , w_9098 , \2903_b1 );
or ( \2905_b1 , \2902_b1 , w_9100 );
or ( \2905_b0 , \2902_b0 , \1507_b0 );
not ( \1507_b0 , w_9101 );
and ( w_9101 , w_9100 , \1507_b1 );
or ( \2906_b1 , \2904_b1 , w_9103 );
not ( w_9103 , w_9104 );
and ( \2906_b0 , \2904_b0 , w_9105 );
and ( w_9104 ,  , w_9105 );
buf ( w_9103 , \2905_b1 );
not ( w_9103 , w_9106 );
not (  , w_9107 );
and ( w_9106 , w_9107 , \2905_b0 );
buf ( \2907_b1 , \2906_b1 );
not ( \2907_b1 , w_9108 );
not ( \2907_b0 , w_9109 );
and ( w_9108 , w_9109 , \2906_b0 );
buf ( \2908_b1 , \1667_b1 );
not ( \2908_b1 , w_9110 );
not ( \2908_b0 , w_9111 );
and ( w_9110 , w_9111 , \1667_b0 );
buf ( \2909_b1 , \2908_b1 );
not ( \2909_b1 , w_9112 );
not ( \2909_b0 , w_9113 );
and ( w_9112 , w_9113 , \2908_b0 );
or ( \2910_b1 , \2907_b1 , w_9114 );
or ( \2910_b0 , \2907_b0 , \2909_b0 );
not ( \2909_b0 , w_9115 );
and ( w_9115 , w_9114 , \2909_b1 );
buf ( \2911_b1 , \732_b1 );
not ( \2911_b1 , w_9116 );
not ( \2911_b0 , w_9117 );
and ( w_9116 , w_9117 , \732_b0 );
or ( \2912_b1 , \2911_b1 , w_9119 );
not ( w_9119 , w_9120 );
and ( \2912_b0 , \2911_b0 , w_9121 );
and ( w_9120 ,  , w_9121 );
buf ( w_9119 , \721_b1 );
not ( w_9119 , w_9122 );
not (  , w_9123 );
and ( w_9122 , w_9123 , \721_b0 );
buf ( \2913_b1 , \2912_b1 );
not ( \2913_b1 , w_9124 );
not ( \2913_b0 , w_9125 );
and ( w_9124 , w_9125 , \2912_b0 );
or ( \2914_b1 , \720_b1 , w_9127 );
not ( w_9127 , w_9128 );
and ( \2914_b0 , \720_b0 , w_9129 );
and ( w_9128 ,  , w_9129 );
buf ( w_9127 , \722_b1 );
not ( w_9127 , w_9130 );
not (  , w_9131 );
and ( w_9130 , w_9131 , \722_b0 );
buf ( \2915_b1 , \2914_b1 );
not ( \2915_b1 , w_9132 );
not ( \2915_b0 , w_9133 );
and ( w_9132 , w_9133 , \2914_b0 );
or ( \2916_b1 , \2913_b1 , w_9134 );
or ( \2916_b0 , \2913_b0 , \2915_b0 );
not ( \2915_b0 , w_9135 );
and ( w_9135 , w_9134 , \2915_b1 );
or ( \2917_b1 , \2914_b1 , w_9136 );
or ( \2917_b0 , \2914_b0 , \2912_b0 );
not ( \2912_b0 , w_9137 );
and ( w_9137 , w_9136 , \2912_b1 );
or ( \2918_b1 , \2916_b1 , w_9139 );
not ( w_9139 , w_9140 );
and ( \2918_b0 , \2916_b0 , w_9141 );
and ( w_9140 ,  , w_9141 );
buf ( w_9139 , \2917_b1 );
not ( w_9139 , w_9142 );
not (  , w_9143 );
and ( w_9142 , w_9143 , \2917_b0 );
or ( \2919_b1 , \707_b1 , \2918_b1 );
not ( \2918_b1 , w_9144 );
and ( \2919_b0 , \707_b0 , w_9145 );
and ( w_9144 , w_9145 , \2918_b0 );
buf ( \2920_b1 , \817_b1 );
not ( \2920_b1 , w_9146 );
not ( \2920_b0 , w_9147 );
and ( w_9146 , w_9147 , \817_b0 );
or ( \2921_b1 , \2920_b1 , w_9149 );
not ( w_9149 , w_9150 );
and ( \2921_b0 , \2920_b0 , w_9151 );
and ( w_9150 ,  , w_9151 );
buf ( w_9149 , \806_b1 );
not ( w_9149 , w_9152 );
not (  , w_9153 );
and ( w_9152 , w_9153 , \806_b0 );
buf ( \2922_b1 , \2921_b1 );
not ( \2922_b1 , w_9154 );
not ( \2922_b0 , w_9155 );
and ( w_9154 , w_9155 , \2921_b0 );
or ( \2923_b1 , \805_b1 , w_9157 );
not ( w_9157 , w_9158 );
and ( \2923_b0 , \805_b0 , w_9159 );
and ( w_9158 ,  , w_9159 );
buf ( w_9157 , \807_b1 );
not ( w_9157 , w_9160 );
not (  , w_9161 );
and ( w_9160 , w_9161 , \807_b0 );
buf ( \2924_b1 , \2923_b1 );
not ( \2924_b1 , w_9162 );
not ( \2924_b0 , w_9163 );
and ( w_9162 , w_9163 , \2923_b0 );
or ( \2925_b1 , \2922_b1 , w_9164 );
or ( \2925_b0 , \2922_b0 , \2924_b0 );
not ( \2924_b0 , w_9165 );
and ( w_9165 , w_9164 , \2924_b1 );
or ( \2926_b1 , \2923_b1 , w_9166 );
or ( \2926_b0 , \2923_b0 , \2921_b0 );
not ( \2921_b0 , w_9167 );
and ( w_9167 , w_9166 , \2921_b1 );
or ( \2927_b1 , \2925_b1 , w_9169 );
not ( w_9169 , w_9170 );
and ( \2927_b0 , \2925_b0 , w_9171 );
and ( w_9170 ,  , w_9171 );
buf ( w_9169 , \2926_b1 );
not ( w_9169 , w_9172 );
not (  , w_9173 );
and ( w_9172 , w_9173 , \2926_b0 );
buf ( \2928_b1 , \2927_b1 );
not ( \2928_b1 , w_9174 );
not ( \2928_b0 , w_9175 );
and ( w_9174 , w_9175 , \2927_b0 );
buf ( \2929_b1 , \879_b1 );
not ( \2929_b1 , w_9176 );
not ( \2929_b0 , w_9177 );
and ( w_9176 , w_9177 , \879_b0 );
or ( \2930_b1 , \2928_b1 , w_9178 );
or ( \2930_b0 , \2928_b0 , \2929_b0 );
not ( \2929_b0 , w_9179 );
and ( w_9179 , w_9178 , \2929_b1 );
or ( \2931_b1 , \894_b1 , \d[3]_b1 );
not ( \d[3]_b1 , w_9180 );
and ( \2931_b0 , \894_b0 , w_9181 );
and ( w_9180 , w_9181 , \d[3]_b0 );
buf ( \2932_b1 , \c[3]_b1 );
not ( \2932_b1 , w_9182 );
not ( \2932_b0 , w_9183 );
and ( w_9182 , w_9183 , \c[3]_b0 );
buf ( \2933_b1 , \907_b1 );
not ( \2933_b1 , w_9184 );
not ( \2933_b0 , w_9185 );
and ( w_9184 , w_9185 , \907_b0 );
or ( \2934_b1 , \2932_b1 , w_9186 );
or ( \2934_b0 , \2932_b0 , \2933_b0 );
not ( \2933_b0 , w_9187 );
and ( w_9187 , w_9186 , \2933_b1 );
or ( \2935_b1 , \885_b1 , w_9189 );
not ( w_9189 , w_9190 );
and ( \2935_b0 , \885_b0 , w_9191 );
and ( w_9190 ,  , w_9191 );
buf ( w_9189 , \b[3]_b1 );
not ( w_9189 , w_9192 );
not (  , w_9193 );
and ( w_9192 , w_9193 , \b[3]_b0 );
or ( \2936_b1 , \2934_b1 , w_9195 );
not ( w_9195 , w_9196 );
and ( \2936_b0 , \2934_b0 , w_9197 );
and ( w_9196 ,  , w_9197 );
buf ( w_9195 , \2935_b1 );
not ( w_9195 , w_9198 );
not (  , w_9199 );
and ( w_9198 , w_9199 , \2935_b0 );
or ( \2937_b1 , \2931_b1 , w_9201 );
not ( w_9201 , w_9202 );
and ( \2937_b0 , \2931_b0 , w_9203 );
and ( w_9202 ,  , w_9203 );
buf ( w_9201 , \2936_b1 );
not ( w_9201 , w_9204 );
not (  , w_9205 );
and ( w_9204 , w_9205 , \2936_b0 );
or ( \2938_b1 , \2930_b1 , w_9207 );
not ( w_9207 , w_9208 );
and ( \2938_b0 , \2930_b0 , w_9209 );
and ( w_9208 ,  , w_9209 );
buf ( w_9207 , \2937_b1 );
not ( w_9207 , w_9210 );
not (  , w_9211 );
and ( w_9210 , w_9211 , \2937_b0 );
or ( \2939_b1 , \2919_b1 , w_9213 );
not ( w_9213 , w_9214 );
and ( \2939_b0 , \2919_b0 , w_9215 );
and ( w_9214 ,  , w_9215 );
buf ( w_9213 , \2938_b1 );
not ( w_9213 , w_9216 );
not (  , w_9217 );
and ( w_9216 , w_9217 , \2938_b0 );
or ( \2940_b1 , \2910_b1 , w_9219 );
not ( w_9219 , w_9220 );
and ( \2940_b0 , \2910_b0 , w_9221 );
and ( w_9220 ,  , w_9221 );
buf ( w_9219 , \2939_b1 );
not ( w_9219 , w_9222 );
not (  , w_9223 );
and ( w_9222 , w_9223 , \2939_b0 );
or ( \2941_b1 , \2900_b1 , w_9225 );
not ( w_9225 , w_9226 );
and ( \2941_b0 , \2900_b0 , w_9227 );
and ( w_9226 ,  , w_9227 );
buf ( w_9225 , \2940_b1 );
not ( w_9225 , w_9228 );
not (  , w_9229 );
and ( w_9228 , w_9229 , \2940_b0 );
or ( \2942_b1 , \2893_b1 , w_9231 );
not ( w_9231 , w_9232 );
and ( \2942_b0 , \2893_b0 , w_9233 );
and ( w_9232 ,  , w_9233 );
buf ( w_9231 , \2941_b1 );
not ( w_9231 , w_9234 );
not (  , w_9235 );
and ( w_9234 , w_9235 , \2941_b0 );
or ( \2943_b1 , \2889_b1 , w_9237 );
not ( w_9237 , w_9238 );
and ( \2943_b0 , \2889_b0 , w_9239 );
and ( w_9238 ,  , w_9239 );
buf ( w_9237 , \2942_b1 );
not ( w_9237 , w_9240 );
not (  , w_9241 );
and ( w_9240 , w_9241 , \2942_b0 );
buf ( \2945_b1 , \2944_b1 );
buf ( \2945_b0 , \2944_b0 );
buf ( \2946_b1 , \922_b1 );
not ( \2946_b1 , w_9242 );
not ( \2946_b0 , w_9243 );
and ( w_9242 , w_9243 , \922_b0 );
or ( \2947_b1 , \2474_b1 , \a[2]_b1 );
not ( \a[2]_b1 , w_9244 );
and ( \2947_b0 , \2474_b0 , w_9245 );
and ( w_9244 , w_9245 , \a[2]_b0 );
or ( \2948_b1 , \2946_b1 , w_9247 );
not ( w_9247 , w_9248 );
and ( \2948_b0 , \2946_b0 , w_9249 );
and ( w_9248 ,  , w_9249 );
buf ( w_9247 , \2947_b1 );
not ( w_9247 , w_9250 );
not (  , w_9251 );
and ( w_9250 , w_9251 , \2947_b0 );
or ( \2949_b1 , \b[2]_b1 , \c[2]_b1 );
not ( \c[2]_b1 , w_9252 );
and ( \2949_b0 , \b[2]_b0 , w_9253 );
and ( w_9252 , w_9253 , \c[2]_b0 );
or ( \2950_b1 , \2887_b1 , \2949_b1 );
not ( \2949_b1 , w_9254 );
and ( \2950_b0 , \2887_b0 , w_9255 );
and ( w_9254 , w_9255 , \2949_b0 );
or ( \2951_b1 , \c[2]_b1 , \d[2]_b1 );
xor ( \2951_b0 , \c[2]_b0 , w_9256 );
not ( w_9256 , w_9257 );
and ( w_9257 , \d[2]_b1 , \d[2]_b0 );
buf ( \2952_b1 , \2951_b1 );
not ( \2952_b1 , w_9258 );
not ( \2952_b0 , w_9259 );
and ( w_9258 , w_9259 , \2951_b0 );
buf ( \2953_b1 , \2614_b1 );
not ( \2953_b1 , w_9260 );
not ( \2953_b0 , w_9261 );
and ( w_9260 , w_9261 , \2614_b0 );
or ( \2954_b1 , \2952_b1 , w_9262 );
or ( \2954_b0 , \2952_b0 , \2953_b0 );
not ( \2953_b0 , w_9263 );
and ( w_9263 , w_9262 , \2953_b1 );
buf ( \2955_b1 , \2222_b1 );
not ( \2955_b1 , w_9264 );
not ( \2955_b0 , w_9265 );
and ( w_9264 , w_9265 , \2222_b0 );
buf ( \2956_b1 , \2224_b1 );
not ( \2956_b1 , w_9266 );
not ( \2956_b0 , w_9267 );
and ( w_9266 , w_9267 , \2224_b0 );
or ( \2957_b1 , \2956_b1 , w_9269 );
not ( w_9269 , w_9270 );
and ( \2957_b0 , \2956_b0 , w_9271 );
and ( w_9270 ,  , w_9271 );
buf ( w_9269 , \2213_b1 );
not ( w_9269 , w_9272 );
not (  , w_9273 );
and ( w_9272 , w_9273 , \2213_b0 );
buf ( \2958_b1 , \2957_b1 );
not ( \2958_b1 , w_9274 );
not ( \2958_b0 , w_9275 );
and ( w_9274 , w_9275 , \2957_b0 );
or ( \2959_b1 , \2955_b1 , w_9276 );
or ( \2959_b0 , \2955_b0 , \2958_b0 );
not ( \2958_b0 , w_9277 );
and ( w_9277 , w_9276 , \2958_b1 );
or ( \2960_b1 , \2957_b1 , w_9278 );
or ( \2960_b0 , \2957_b0 , \2222_b0 );
not ( \2222_b0 , w_9279 );
and ( w_9279 , w_9278 , \2222_b1 );
or ( \2961_b1 , \2959_b1 , w_9281 );
not ( w_9281 , w_9282 );
and ( \2961_b0 , \2959_b0 , w_9283 );
and ( w_9282 ,  , w_9283 );
buf ( w_9281 , \2960_b1 );
not ( w_9281 , w_9284 );
not (  , w_9285 );
and ( w_9284 , w_9285 , \2960_b0 );
or ( \2962_b1 , \2413_b1 , \2961_b1 );
not ( \2961_b1 , w_9286 );
and ( \2962_b0 , \2413_b0 , w_9287 );
and ( w_9286 , w_9287 , \2961_b0 );
buf ( \2963_b1 , \1504_b1 );
not ( \2963_b1 , w_9288 );
not ( \2963_b0 , w_9289 );
and ( w_9288 , w_9289 , \1504_b0 );
buf ( \2964_b1 , \1506_b1 );
not ( \2964_b1 , w_9290 );
not ( \2964_b0 , w_9291 );
and ( w_9290 , w_9291 , \1506_b0 );
or ( \2965_b1 , \2964_b1 , w_9293 );
not ( w_9293 , w_9294 );
and ( \2965_b0 , \2964_b0 , w_9295 );
and ( w_9294 ,  , w_9295 );
buf ( w_9293 , \1496_b1 );
not ( w_9293 , w_9296 );
not (  , w_9297 );
and ( w_9296 , w_9297 , \1496_b0 );
buf ( \2966_b1 , \2965_b1 );
not ( \2966_b1 , w_9298 );
not ( \2966_b0 , w_9299 );
and ( w_9298 , w_9299 , \2965_b0 );
or ( \2967_b1 , \2963_b1 , w_9300 );
or ( \2967_b0 , \2963_b0 , \2966_b0 );
not ( \2966_b0 , w_9301 );
and ( w_9301 , w_9300 , \2966_b1 );
or ( \2968_b1 , \2965_b1 , w_9302 );
or ( \2968_b0 , \2965_b0 , \1504_b0 );
not ( \1504_b0 , w_9303 );
and ( w_9303 , w_9302 , \1504_b1 );
or ( \2969_b1 , \2967_b1 , w_9305 );
not ( w_9305 , w_9306 );
and ( \2969_b0 , \2967_b0 , w_9307 );
and ( w_9306 ,  , w_9307 );
buf ( w_9305 , \2968_b1 );
not ( w_9305 , w_9308 );
not (  , w_9309 );
and ( w_9308 , w_9309 , \2968_b0 );
buf ( \2970_b1 , \2969_b1 );
not ( \2970_b1 , w_9310 );
not ( \2970_b0 , w_9311 );
and ( w_9310 , w_9311 , \2969_b0 );
buf ( \2971_b1 , \2908_b1 );
not ( \2971_b1 , w_9312 );
not ( \2971_b0 , w_9313 );
and ( w_9312 , w_9313 , \2908_b0 );
or ( \2972_b1 , \2970_b1 , w_9314 );
or ( \2972_b0 , \2970_b0 , \2971_b0 );
not ( \2971_b0 , w_9315 );
and ( w_9315 , w_9314 , \2971_b1 );
or ( \2973_b1 , \719_b1 , w_9317 );
not ( w_9317 , w_9318 );
and ( \2973_b0 , \719_b0 , w_9319 );
and ( w_9318 ,  , w_9319 );
buf ( w_9317 , \722_b1 );
not ( w_9317 , w_9320 );
not (  , w_9321 );
and ( w_9320 , w_9321 , \722_b0 );
buf ( \2974_b1 , \2973_b1 );
not ( \2974_b1 , w_9322 );
not ( \2974_b0 , w_9323 );
and ( w_9322 , w_9323 , \2973_b0 );
buf ( \2975_b1 , \714_b1 );
not ( \2975_b1 , w_9324 );
not ( \2975_b0 , w_9325 );
and ( w_9324 , w_9325 , \714_b0 );
buf ( \2976_b1 , \2975_b1 );
not ( \2976_b1 , w_9326 );
not ( \2976_b0 , w_9327 );
and ( w_9326 , w_9327 , \2975_b0 );
buf ( \2977_b1 , \717_b1 );
not ( \2977_b1 , w_9328 );
not ( \2977_b0 , w_9329 );
and ( w_9328 , w_9329 , \717_b0 );
or ( \2978_b1 , \2976_b1 , w_9330 );
or ( \2978_b0 , \2976_b0 , \2977_b0 );
not ( \2977_b0 , w_9331 );
and ( w_9331 , w_9330 , \2977_b1 );
or ( \2979_b1 , \2978_b1 , w_9333 );
not ( w_9333 , w_9334 );
and ( \2979_b0 , \2978_b0 , w_9335 );
and ( w_9334 ,  , w_9335 );
buf ( w_9333 , \715_b1 );
not ( w_9333 , w_9336 );
not (  , w_9337 );
and ( w_9336 , w_9337 , \715_b0 );
buf ( \2980_b1 , \2979_b1 );
not ( \2980_b1 , w_9338 );
not ( \2980_b0 , w_9339 );
and ( w_9338 , w_9339 , \2979_b0 );
or ( \2981_b1 , \2974_b1 , w_9340 );
or ( \2981_b0 , \2974_b0 , \2980_b0 );
not ( \2980_b0 , w_9341 );
and ( w_9341 , w_9340 , \2980_b1 );
or ( \2982_b1 , \2979_b1 , w_9342 );
or ( \2982_b0 , \2979_b0 , \2973_b0 );
not ( \2973_b0 , w_9343 );
and ( w_9343 , w_9342 , \2973_b1 );
or ( \2983_b1 , \2981_b1 , w_9345 );
not ( w_9345 , w_9346 );
and ( \2983_b0 , \2981_b0 , w_9347 );
and ( w_9346 ,  , w_9347 );
buf ( w_9345 , \2982_b1 );
not ( w_9345 , w_9348 );
not (  , w_9349 );
and ( w_9348 , w_9349 , \2982_b0 );
or ( \2984_b1 , \707_b1 , \2983_b1 );
not ( \2983_b1 , w_9350 );
and ( \2984_b0 , \707_b0 , w_9351 );
and ( w_9350 , w_9351 , \2983_b0 );
or ( \2985_b1 , \804_b1 , w_9353 );
not ( w_9353 , w_9354 );
and ( \2985_b0 , \804_b0 , w_9355 );
and ( w_9354 ,  , w_9355 );
buf ( w_9353 , \807_b1 );
not ( w_9353 , w_9356 );
not (  , w_9357 );
and ( w_9356 , w_9357 , \807_b0 );
buf ( \2986_b1 , \2985_b1 );
not ( \2986_b1 , w_9358 );
not ( \2986_b0 , w_9359 );
and ( w_9358 , w_9359 , \2985_b0 );
buf ( \2987_b1 , \799_b1 );
not ( \2987_b1 , w_9360 );
not ( \2987_b0 , w_9361 );
and ( w_9360 , w_9361 , \799_b0 );
buf ( \2988_b1 , \2987_b1 );
not ( \2988_b1 , w_9362 );
not ( \2988_b0 , w_9363 );
and ( w_9362 , w_9363 , \2987_b0 );
buf ( \2989_b1 , \802_b1 );
not ( \2989_b1 , w_9364 );
not ( \2989_b0 , w_9365 );
and ( w_9364 , w_9365 , \802_b0 );
or ( \2990_b1 , \2988_b1 , w_9366 );
or ( \2990_b0 , \2988_b0 , \2989_b0 );
not ( \2989_b0 , w_9367 );
and ( w_9367 , w_9366 , \2989_b1 );
or ( \2991_b1 , \2990_b1 , w_9369 );
not ( w_9369 , w_9370 );
and ( \2991_b0 , \2990_b0 , w_9371 );
and ( w_9370 ,  , w_9371 );
buf ( w_9369 , \800_b1 );
not ( w_9369 , w_9372 );
not (  , w_9373 );
and ( w_9372 , w_9373 , \800_b0 );
buf ( \2992_b1 , \2991_b1 );
not ( \2992_b1 , w_9374 );
not ( \2992_b0 , w_9375 );
and ( w_9374 , w_9375 , \2991_b0 );
or ( \2993_b1 , \2986_b1 , w_9376 );
or ( \2993_b0 , \2986_b0 , \2992_b0 );
not ( \2992_b0 , w_9377 );
and ( w_9377 , w_9376 , \2992_b1 );
or ( \2994_b1 , \2991_b1 , w_9378 );
or ( \2994_b0 , \2991_b0 , \2985_b0 );
not ( \2985_b0 , w_9379 );
and ( w_9379 , w_9378 , \2985_b1 );
or ( \2995_b1 , \2993_b1 , w_9381 );
not ( w_9381 , w_9382 );
and ( \2995_b0 , \2993_b0 , w_9383 );
and ( w_9382 ,  , w_9383 );
buf ( w_9381 , \2994_b1 );
not ( w_9381 , w_9384 );
not (  , w_9385 );
and ( w_9384 , w_9385 , \2994_b0 );
buf ( \2996_b1 , \2995_b1 );
not ( \2996_b1 , w_9386 );
not ( \2996_b0 , w_9387 );
and ( w_9386 , w_9387 , \2995_b0 );
buf ( \2997_b1 , \879_b1 );
not ( \2997_b1 , w_9388 );
not ( \2997_b0 , w_9389 );
and ( w_9388 , w_9389 , \879_b0 );
or ( \2998_b1 , \2996_b1 , w_9390 );
or ( \2998_b0 , \2996_b0 , \2997_b0 );
not ( \2997_b0 , w_9391 );
and ( w_9391 , w_9390 , \2997_b1 );
or ( \2999_b1 , \894_b1 , \d[2]_b1 );
not ( \d[2]_b1 , w_9392 );
and ( \2999_b0 , \894_b0 , w_9393 );
and ( w_9392 , w_9393 , \d[2]_b0 );
buf ( \3000_b1 , \c[2]_b1 );
not ( \3000_b1 , w_9394 );
not ( \3000_b0 , w_9395 );
and ( w_9394 , w_9395 , \c[2]_b0 );
buf ( \3001_b1 , \907_b1 );
not ( \3001_b1 , w_9396 );
not ( \3001_b0 , w_9397 );
and ( w_9396 , w_9397 , \907_b0 );
or ( \3002_b1 , \3000_b1 , w_9398 );
or ( \3002_b0 , \3000_b0 , \3001_b0 );
not ( \3001_b0 , w_9399 );
and ( w_9399 , w_9398 , \3001_b1 );
or ( \3003_b1 , \885_b1 , w_9401 );
not ( w_9401 , w_9402 );
and ( \3003_b0 , \885_b0 , w_9403 );
and ( w_9402 ,  , w_9403 );
buf ( w_9401 , \b[2]_b1 );
not ( w_9401 , w_9404 );
not (  , w_9405 );
and ( w_9404 , w_9405 , \b[2]_b0 );
or ( \3004_b1 , \3002_b1 , w_9407 );
not ( w_9407 , w_9408 );
and ( \3004_b0 , \3002_b0 , w_9409 );
and ( w_9408 ,  , w_9409 );
buf ( w_9407 , \3003_b1 );
not ( w_9407 , w_9410 );
not (  , w_9411 );
and ( w_9410 , w_9411 , \3003_b0 );
or ( \3005_b1 , \2999_b1 , w_9413 );
not ( w_9413 , w_9414 );
and ( \3005_b0 , \2999_b0 , w_9415 );
and ( w_9414 ,  , w_9415 );
buf ( w_9413 , \3004_b1 );
not ( w_9413 , w_9416 );
not (  , w_9417 );
and ( w_9416 , w_9417 , \3004_b0 );
or ( \3006_b1 , \2998_b1 , w_9419 );
not ( w_9419 , w_9420 );
and ( \3006_b0 , \2998_b0 , w_9421 );
and ( w_9420 ,  , w_9421 );
buf ( w_9419 , \3005_b1 );
not ( w_9419 , w_9422 );
not (  , w_9423 );
and ( w_9422 , w_9423 , \3005_b0 );
or ( \3007_b1 , \2984_b1 , w_9425 );
not ( w_9425 , w_9426 );
and ( \3007_b0 , \2984_b0 , w_9427 );
and ( w_9426 ,  , w_9427 );
buf ( w_9425 , \3006_b1 );
not ( w_9425 , w_9428 );
not (  , w_9429 );
and ( w_9428 , w_9429 , \3006_b0 );
or ( \3008_b1 , \2972_b1 , w_9431 );
not ( w_9431 , w_9432 );
and ( \3008_b0 , \2972_b0 , w_9433 );
and ( w_9432 ,  , w_9433 );
buf ( w_9431 , \3007_b1 );
not ( w_9431 , w_9434 );
not (  , w_9435 );
and ( w_9434 , w_9435 , \3007_b0 );
or ( \3009_b1 , \2962_b1 , w_9437 );
not ( w_9437 , w_9438 );
and ( \3009_b0 , \2962_b0 , w_9439 );
and ( w_9438 ,  , w_9439 );
buf ( w_9437 , \3008_b1 );
not ( w_9437 , w_9440 );
not (  , w_9441 );
and ( w_9440 , w_9441 , \3008_b0 );
or ( \3010_b1 , \2954_b1 , w_9443 );
not ( w_9443 , w_9444 );
and ( \3010_b0 , \2954_b0 , w_9445 );
and ( w_9444 ,  , w_9445 );
buf ( w_9443 , \3009_b1 );
not ( w_9443 , w_9446 );
not (  , w_9447 );
and ( w_9446 , w_9447 , \3009_b0 );
or ( \3011_b1 , \2950_b1 , w_9449 );
not ( w_9449 , w_9450 );
and ( \3011_b0 , \2950_b0 , w_9451 );
and ( w_9450 ,  , w_9451 );
buf ( w_9449 , \3010_b1 );
not ( w_9449 , w_9452 );
not (  , w_9453 );
and ( w_9452 , w_9453 , \3010_b0 );
buf ( \3012_b1 , \683_b1 );
not ( \3012_b1 , w_9454 );
not ( \3012_b0 , w_9455 );
and ( w_9454 , w_9455 , \683_b0 );
or ( \3013_b1 , \3012_b1 , w_9457 );
not ( w_9457 , w_9458 );
and ( \3013_b0 , \3012_b0 , w_9459 );
and ( w_9458 ,  , w_9459 );
buf ( w_9457 , \648_b1 );
not ( w_9457 , w_9460 );
not (  , w_9461 );
and ( w_9460 , w_9461 , \648_b0 );
or ( \3014_b1 , \b[2]_b1 , w_9462 );
or ( \3014_b0 , \b[2]_b0 , \a[2]_b0 );
not ( \a[2]_b0 , w_9463 );
and ( w_9463 , w_9462 , \a[2]_b1 );
or ( \3015_b1 , \3014_b1 , w_9465 );
not ( w_9465 , w_9466 );
and ( \3015_b0 , \3014_b0 , w_9467 );
and ( w_9466 ,  , w_9467 );
buf ( w_9465 , \667_b1 );
not ( w_9465 , w_9468 );
not (  , w_9469 );
and ( w_9468 , w_9469 , \667_b0 );
or ( \3017_b1 , \b[1]_b1 , \c[1]_b1 );
not ( \c[1]_b1 , w_9470 );
and ( \3017_b0 , \b[1]_b0 , w_9471 );
and ( w_9470 , w_9471 , \c[1]_b0 );
or ( \3018_b1 , \922_b1 , \3017_b1 );
not ( \3017_b1 , w_9472 );
and ( \3018_b0 , \922_b0 , w_9473 );
and ( w_9472 , w_9473 , \3017_b0 );
or ( \3019_b1 , \c[1]_b1 , \d[1]_b1 );
xor ( \3019_b0 , \c[1]_b0 , w_9474 );
not ( w_9474 , w_9475 );
and ( w_9475 , \d[1]_b1 , \d[1]_b0 );
buf ( \3020_b1 , \3019_b1 );
not ( \3020_b1 , w_9476 );
not ( \3020_b0 , w_9477 );
and ( w_9476 , w_9477 , \3019_b0 );
buf ( \3021_b1 , \2614_b1 );
not ( \3021_b1 , w_9478 );
not ( \3021_b0 , w_9479 );
and ( w_9478 , w_9479 , \2614_b0 );
or ( \3022_b1 , \3020_b1 , w_9480 );
or ( \3022_b0 , \3020_b0 , \3021_b0 );
not ( \3021_b0 , w_9481 );
and ( w_9481 , w_9480 , \3021_b1 );
or ( \3023_b1 , \2219_b1 , w_9482 );
or ( \3023_b0 , \2219_b0 , \2221_b0 );
not ( \2221_b0 , w_9483 );
and ( w_9483 , w_9482 , \2221_b1 );
or ( \3024_b1 , \2222_b1 , \3023_b1 );
not ( \3023_b1 , w_9484 );
and ( \3024_b0 , \2222_b0 , w_9485 );
and ( w_9484 , w_9485 , \3023_b0 );
or ( \3025_b1 , \2413_b1 , \3024_b1 );
not ( \3024_b1 , w_9486 );
and ( \3025_b0 , \2413_b0 , w_9487 );
and ( w_9486 , w_9487 , \3024_b0 );
or ( \3026_b1 , \1502_b1 , w_9488 );
or ( \3026_b0 , \1502_b0 , \1503_b0 );
not ( \1503_b0 , w_9489 );
and ( w_9489 , w_9488 , \1503_b1 );
or ( \3027_b1 , \1504_b1 , \3026_b1 );
not ( \3026_b1 , w_9490 );
and ( \3027_b0 , \1504_b0 , w_9491 );
and ( w_9490 , w_9491 , \3026_b0 );
buf ( \3028_b1 , \3027_b1 );
not ( \3028_b1 , w_9492 );
not ( \3028_b0 , w_9493 );
and ( w_9492 , w_9493 , \3027_b0 );
buf ( \3029_b1 , \2908_b1 );
not ( \3029_b1 , w_9494 );
not ( \3029_b0 , w_9495 );
and ( w_9494 , w_9495 , \2908_b0 );
or ( \3030_b1 , \3028_b1 , w_9496 );
or ( \3030_b0 , \3028_b0 , \3029_b0 );
not ( \3029_b0 , w_9497 );
and ( w_9497 , w_9496 , \3029_b1 );
buf ( \3031_b1 , \2975_b1 );
not ( \3031_b1 , w_9498 );
not ( \3031_b0 , w_9499 );
and ( w_9498 , w_9499 , \2975_b0 );
or ( \3032_b1 , \717_b1 , w_9501 );
not ( w_9501 , w_9502 );
and ( \3032_b0 , \717_b0 , w_9503 );
and ( w_9502 ,  , w_9503 );
buf ( w_9501 , \715_b1 );
not ( w_9501 , w_9504 );
not (  , w_9505 );
and ( w_9504 , w_9505 , \715_b0 );
buf ( \3033_b1 , \3032_b1 );
not ( \3033_b1 , w_9506 );
not ( \3033_b0 , w_9507 );
and ( w_9506 , w_9507 , \3032_b0 );
or ( \3034_b1 , \3031_b1 , w_9508 );
or ( \3034_b0 , \3031_b0 , \3033_b0 );
not ( \3033_b0 , w_9509 );
and ( w_9509 , w_9508 , \3033_b1 );
or ( \3035_b1 , \3032_b1 , w_9510 );
or ( \3035_b0 , \3032_b0 , \2975_b0 );
not ( \2975_b0 , w_9511 );
and ( w_9511 , w_9510 , \2975_b1 );
or ( \3036_b1 , \3034_b1 , w_9513 );
not ( w_9513 , w_9514 );
and ( \3036_b0 , \3034_b0 , w_9515 );
and ( w_9514 ,  , w_9515 );
buf ( w_9513 , \3035_b1 );
not ( w_9513 , w_9516 );
not (  , w_9517 );
and ( w_9516 , w_9517 , \3035_b0 );
or ( \3037_b1 , \707_b1 , \3036_b1 );
not ( \3036_b1 , w_9518 );
and ( \3037_b0 , \707_b0 , w_9519 );
and ( w_9518 , w_9519 , \3036_b0 );
buf ( \3038_b1 , \2987_b1 );
not ( \3038_b1 , w_9520 );
not ( \3038_b0 , w_9521 );
and ( w_9520 , w_9521 , \2987_b0 );
or ( \3039_b1 , \802_b1 , w_9523 );
not ( w_9523 , w_9524 );
and ( \3039_b0 , \802_b0 , w_9525 );
and ( w_9524 ,  , w_9525 );
buf ( w_9523 , \800_b1 );
not ( w_9523 , w_9526 );
not (  , w_9527 );
and ( w_9526 , w_9527 , \800_b0 );
buf ( \3040_b1 , \3039_b1 );
not ( \3040_b1 , w_9528 );
not ( \3040_b0 , w_9529 );
and ( w_9528 , w_9529 , \3039_b0 );
or ( \3041_b1 , \3038_b1 , w_9530 );
or ( \3041_b0 , \3038_b0 , \3040_b0 );
not ( \3040_b0 , w_9531 );
and ( w_9531 , w_9530 , \3040_b1 );
or ( \3042_b1 , \3039_b1 , w_9532 );
or ( \3042_b0 , \3039_b0 , \2987_b0 );
not ( \2987_b0 , w_9533 );
and ( w_9533 , w_9532 , \2987_b1 );
or ( \3043_b1 , \3041_b1 , w_9535 );
not ( w_9535 , w_9536 );
and ( \3043_b0 , \3041_b0 , w_9537 );
and ( w_9536 ,  , w_9537 );
buf ( w_9535 , \3042_b1 );
not ( w_9535 , w_9538 );
not (  , w_9539 );
and ( w_9538 , w_9539 , \3042_b0 );
buf ( \3044_b1 , \3043_b1 );
not ( \3044_b1 , w_9540 );
not ( \3044_b0 , w_9541 );
and ( w_9540 , w_9541 , \3043_b0 );
buf ( \3045_b1 , \879_b1 );
not ( \3045_b1 , w_9542 );
not ( \3045_b0 , w_9543 );
and ( w_9542 , w_9543 , \879_b0 );
or ( \3046_b1 , \3044_b1 , w_9544 );
or ( \3046_b0 , \3044_b0 , \3045_b0 );
not ( \3045_b0 , w_9545 );
and ( w_9545 , w_9544 , \3045_b1 );
or ( \3047_b1 , \894_b1 , \d[1]_b1 );
not ( \d[1]_b1 , w_9546 );
and ( \3047_b0 , \894_b0 , w_9547 );
and ( w_9546 , w_9547 , \d[1]_b0 );
buf ( \3048_b1 , \c[1]_b1 );
not ( \3048_b1 , w_9548 );
not ( \3048_b0 , w_9549 );
and ( w_9548 , w_9549 , \c[1]_b0 );
buf ( \3049_b1 , \907_b1 );
not ( \3049_b1 , w_9550 );
not ( \3049_b0 , w_9551 );
and ( w_9550 , w_9551 , \907_b0 );
or ( \3050_b1 , \3048_b1 , w_9552 );
or ( \3050_b0 , \3048_b0 , \3049_b0 );
not ( \3049_b0 , w_9553 );
and ( w_9553 , w_9552 , \3049_b1 );
or ( \3051_b1 , \885_b1 , w_9555 );
not ( w_9555 , w_9556 );
and ( \3051_b0 , \885_b0 , w_9557 );
and ( w_9556 ,  , w_9557 );
buf ( w_9555 , \b[1]_b1 );
not ( w_9555 , w_9558 );
not (  , w_9559 );
and ( w_9558 , w_9559 , \b[1]_b0 );
or ( \3052_b1 , \3050_b1 , w_9561 );
not ( w_9561 , w_9562 );
and ( \3052_b0 , \3050_b0 , w_9563 );
and ( w_9562 ,  , w_9563 );
buf ( w_9561 , \3051_b1 );
not ( w_9561 , w_9564 );
not (  , w_9565 );
and ( w_9564 , w_9565 , \3051_b0 );
or ( \3053_b1 , \3047_b1 , w_9567 );
not ( w_9567 , w_9568 );
and ( \3053_b0 , \3047_b0 , w_9569 );
and ( w_9568 ,  , w_9569 );
buf ( w_9567 , \3052_b1 );
not ( w_9567 , w_9570 );
not (  , w_9571 );
and ( w_9570 , w_9571 , \3052_b0 );
or ( \3054_b1 , \3046_b1 , w_9573 );
not ( w_9573 , w_9574 );
and ( \3054_b0 , \3046_b0 , w_9575 );
and ( w_9574 ,  , w_9575 );
buf ( w_9573 , \3053_b1 );
not ( w_9573 , w_9576 );
not (  , w_9577 );
and ( w_9576 , w_9577 , \3053_b0 );
or ( \3055_b1 , \3037_b1 , w_9579 );
not ( w_9579 , w_9580 );
and ( \3055_b0 , \3037_b0 , w_9581 );
and ( w_9580 ,  , w_9581 );
buf ( w_9579 , \3054_b1 );
not ( w_9579 , w_9582 );
not (  , w_9583 );
and ( w_9582 , w_9583 , \3054_b0 );
or ( \3056_b1 , \3030_b1 , w_9585 );
not ( w_9585 , w_9586 );
and ( \3056_b0 , \3030_b0 , w_9587 );
and ( w_9586 ,  , w_9587 );
buf ( w_9585 , \3055_b1 );
not ( w_9585 , w_9588 );
not (  , w_9589 );
and ( w_9588 , w_9589 , \3055_b0 );
or ( \3057_b1 , \3025_b1 , w_9591 );
not ( w_9591 , w_9592 );
and ( \3057_b0 , \3025_b0 , w_9593 );
and ( w_9592 ,  , w_9593 );
buf ( w_9591 , \3056_b1 );
not ( w_9591 , w_9594 );
not (  , w_9595 );
and ( w_9594 , w_9595 , \3056_b0 );
or ( \3058_b1 , \3022_b1 , w_9597 );
not ( w_9597 , w_9598 );
and ( \3058_b0 , \3022_b0 , w_9599 );
and ( w_9598 ,  , w_9599 );
buf ( w_9597 , \3057_b1 );
not ( w_9597 , w_9600 );
not (  , w_9601 );
and ( w_9600 , w_9601 , \3057_b0 );
or ( \3059_b1 , \3018_b1 , w_9603 );
not ( w_9603 , w_9604 );
and ( \3059_b0 , \3018_b0 , w_9605 );
and ( w_9604 ,  , w_9605 );
buf ( w_9603 , \3058_b1 );
not ( w_9603 , w_9606 );
not (  , w_9607 );
and ( w_9606 , w_9607 , \3058_b0 );
or ( \3060_b1 , \2474_b1 , \a[1]_b1 );
not ( \a[1]_b1 , w_9608 );
and ( \3060_b0 , \2474_b0 , w_9609 );
and ( w_9608 , w_9609 , \a[1]_b0 );
or ( \3061_b1 , \3060_b1 , w_9611 );
not ( w_9611 , w_9612 );
and ( \3061_b0 , \3060_b0 , w_9613 );
and ( w_9612 ,  , w_9613 );
buf ( w_9611 , \2886_b1 );
not ( w_9611 , w_9614 );
not (  , w_9615 );
and ( w_9614 , w_9615 , \2886_b0 );
buf ( \3062_b1 , \b[1]_b1 );
not ( \3062_b1 , w_9616 );
not ( \3062_b0 , w_9617 );
and ( w_9616 , w_9617 , \b[1]_b0 );
buf ( \3063_b1 , \3062_b1 );
not ( \3063_b1 , w_9618 );
not ( \3063_b0 , w_9619 );
and ( w_9618 , w_9619 , \3062_b0 );
buf ( \3064_b1 , \a[1]_b1 );
not ( \3064_b1 , w_9620 );
not ( \3064_b0 , w_9621 );
and ( w_9620 , w_9621 , \a[1]_b0 );
buf ( \3065_b1 , \3064_b1 );
not ( \3065_b1 , w_9622 );
not ( \3065_b0 , w_9623 );
and ( w_9622 , w_9623 , \3064_b0 );
or ( \3066_b1 , \3063_b1 , w_9624 );
or ( \3066_b0 , \3063_b0 , \3065_b0 );
not ( \3065_b0 , w_9625 );
and ( w_9625 , w_9624 , \3065_b1 );
or ( \3067_b1 , \3066_b1 , w_9627 );
not ( w_9627 , w_9628 );
and ( \3067_b0 , \3066_b0 , w_9629 );
and ( w_9628 ,  , w_9629 );
buf ( w_9627 , \667_b1 );
not ( w_9627 , w_9630 );
not (  , w_9631 );
and ( w_9630 , w_9631 , \667_b0 );
buf ( \3068_b1 , \680_b1 );
not ( \3068_b1 , w_9632 );
not ( \3068_b0 , w_9633 );
and ( w_9632 , w_9633 , \680_b0 );
or ( \3069_b1 , \3068_b1 , w_9635 );
not ( w_9635 , w_9636 );
and ( \3069_b0 , \3068_b0 , w_9637 );
and ( w_9636 ,  , w_9637 );
buf ( w_9635 , \648_b1 );
not ( w_9635 , w_9638 );
not (  , w_9639 );
and ( w_9638 , w_9639 , \648_b0 );
buf ( \3071_b1 , \a[8]_b1 );
not ( \3071_b1 , w_9640 );
not ( \3071_b0 , w_9641 );
and ( w_9640 , w_9641 , \a[8]_b0 );
buf ( \3072_b1 , \2857_b1 );
not ( \3072_b1 , w_9642 );
not ( \3072_b0 , w_9643 );
and ( w_9642 , w_9643 , \2857_b0 );
buf ( \3073_b1 , \3072_b1 );
not ( \3073_b1 , w_9644 );
not ( \3073_b0 , w_9645 );
and ( w_9644 , w_9645 , \3072_b0 );
or ( \3074_b1 , \648_b1 , w_9647 );
not ( w_9647 , w_9648 );
and ( \3074_b0 , \648_b0 , w_9649 );
and ( w_9648 ,  , w_9649 );
buf ( w_9647 , \666_b1 );
not ( w_9647 , w_9650 );
not (  , w_9651 );
and ( w_9650 , w_9651 , \666_b0 );
or ( \3075_b1 , \3073_b1 , w_9653 );
not ( w_9653 , w_9654 );
and ( \3075_b0 , \3073_b0 , w_9655 );
and ( w_9654 ,  , w_9655 );
buf ( w_9653 , \3074_b1 );
not ( w_9653 , w_9656 );
not (  , w_9657 );
and ( w_9656 , w_9657 , \3074_b0 );
buf ( \3076_b1 , \3075_b1 );
not ( \3076_b1 , w_9658 );
not ( \3076_b0 , w_9659 );
and ( w_9658 , w_9659 , \3075_b0 );
or ( \3077_b1 , \3071_b1 , w_9660 );
or ( \3077_b0 , \3071_b0 , \3076_b0 );
not ( \3076_b0 , w_9661 );
and ( w_9661 , w_9660 , \3076_b1 );
buf ( \3078_b1 , \c[8]_b1 );
not ( \3078_b1 , w_9662 );
not ( \3078_b0 , w_9663 );
and ( w_9662 , w_9663 , \c[8]_b0 );
buf ( \3079_b1 , \922_b1 );
not ( \3079_b1 , w_9664 );
not ( \3079_b0 , w_9665 );
and ( w_9664 , w_9665 , \922_b0 );
or ( \3080_b1 , \3078_b1 , w_9666 );
or ( \3080_b0 , \3078_b0 , \3079_b0 );
not ( \3079_b0 , w_9667 );
and ( w_9667 , w_9666 , \3079_b1 );
buf ( \3081_b1 , \667_b1 );
not ( \3081_b1 , w_9668 );
not ( \3081_b0 , w_9669 );
and ( w_9668 , w_9669 , \667_b0 );
or ( \3082_b1 , \3080_b1 , w_9671 );
not ( w_9671 , w_9672 );
and ( \3082_b0 , \3080_b0 , w_9673 );
and ( w_9672 ,  , w_9673 );
buf ( w_9671 , \3081_b1 );
not ( w_9671 , w_9674 );
not (  , w_9675 );
and ( w_9674 , w_9675 , \3081_b0 );
or ( \3083_b1 , \3082_b1 , \b[8]_b1 );
not ( \b[8]_b1 , w_9676 );
and ( \3083_b0 , \3082_b0 , w_9677 );
and ( w_9676 , w_9677 , \b[8]_b0 );
buf ( \3084_b1 , \d[8]_b1 );
not ( \3084_b1 , w_9678 );
not ( \3084_b0 , w_9679 );
and ( w_9678 , w_9679 , \d[8]_b0 );
buf ( \3085_b1 , \648_b1 );
not ( \3085_b1 , w_9680 );
not ( \3085_b0 , w_9681 );
and ( w_9680 , w_9681 , \648_b0 );
or ( \3086_b1 , \3084_b1 , w_9682 );
or ( \3086_b0 , \3084_b0 , \3085_b0 );
not ( \3085_b0 , w_9683 );
and ( w_9683 , w_9682 , \3085_b1 );
buf ( \3087_b1 , \1527_b1 );
not ( \3087_b1 , w_9684 );
not ( \3087_b0 , w_9685 );
and ( w_9684 , w_9685 , \1527_b0 );
buf ( \3088_b1 , \1287_b1 );
buf ( \3088_b0 , \1287_b0 );
buf ( \3089_b1 , \1534_b1 );
buf ( \3089_b0 , \1534_b0 );
or ( \3090_b1 , \3088_b1 , w_9687 );
not ( w_9687 , w_9688 );
and ( \3090_b0 , \3088_b0 , w_9689 );
and ( w_9688 ,  , w_9689 );
buf ( w_9687 , \3089_b1 );
not ( w_9687 , w_9690 );
not (  , w_9691 );
and ( w_9690 , w_9691 , \3089_b0 );
buf ( \3091_b1 , \3090_b1 );
not ( \3091_b1 , w_9692 );
not ( \3091_b0 , w_9693 );
and ( w_9692 , w_9693 , \3090_b0 );
or ( \3092_b1 , \3087_b1 , w_9694 );
or ( \3092_b0 , \3087_b0 , \3091_b0 );
not ( \3091_b0 , w_9695 );
and ( w_9695 , w_9694 , \3091_b1 );
or ( \3093_b1 , \1528_b1 , w_9696 );
or ( \3093_b0 , \1528_b0 , \3090_b0 );
not ( \3090_b0 , w_9697 );
and ( w_9697 , w_9696 , \3090_b1 );
or ( \3094_b1 , \3092_b1 , w_9699 );
not ( w_9699 , w_9700 );
and ( \3094_b0 , \3092_b0 , w_9701 );
and ( w_9700 ,  , w_9701 );
buf ( w_9699 , \3093_b1 );
not ( w_9699 , w_9702 );
not (  , w_9703 );
and ( w_9702 , w_9703 , \3093_b0 );
or ( \3095_b1 , \3094_b1 , \2908_b1 );
not ( \2908_b1 , w_9704 );
and ( \3095_b0 , \3094_b0 , w_9705 );
and ( w_9704 , w_9705 , \2908_b0 );
buf ( \3096_b1 , \837_b1 );
not ( \3096_b1 , w_9706 );
not ( \3096_b0 , w_9707 );
and ( w_9706 , w_9707 , \837_b0 );
or ( \3097_b1 , \3096_b1 , w_9709 );
not ( w_9709 , w_9710 );
and ( \3097_b0 , \3096_b0 , w_9711 );
and ( w_9710 ,  , w_9711 );
buf ( w_9709 , \848_b1 );
not ( w_9709 , w_9712 );
not (  , w_9713 );
and ( w_9712 , w_9713 , \848_b0 );
buf ( \3098_b1 , \3097_b1 );
not ( \3098_b1 , w_9714 );
not ( \3098_b0 , w_9715 );
and ( w_9714 , w_9715 , \3097_b0 );
buf ( \3099_b1 , \832_b1 );
not ( \3099_b1 , w_9716 );
not ( \3099_b0 , w_9717 );
and ( w_9716 , w_9717 , \832_b0 );
or ( \3100_b1 , \3098_b1 , w_9718 );
or ( \3100_b0 , \3098_b0 , \3099_b0 );
not ( \3099_b0 , w_9719 );
and ( w_9719 , w_9718 , \3099_b1 );
or ( \3101_b1 , \832_b1 , w_9720 );
or ( \3101_b0 , \832_b0 , \3097_b0 );
not ( \3097_b0 , w_9721 );
and ( w_9721 , w_9720 , \3097_b1 );
or ( \3102_b1 , \3100_b1 , w_9723 );
not ( w_9723 , w_9724 );
and ( \3102_b0 , \3100_b0 , w_9725 );
and ( w_9724 ,  , w_9725 );
buf ( w_9723 , \3101_b1 );
not ( w_9723 , w_9726 );
not (  , w_9727 );
and ( w_9726 , w_9727 , \3101_b0 );
buf ( \3103_b1 , \3102_b1 );
not ( \3103_b1 , w_9728 );
not ( \3103_b0 , w_9729 );
and ( w_9728 , w_9729 , \3102_b0 );
buf ( \3104_b1 , \880_b1 );
not ( \3104_b1 , w_9730 );
not ( \3104_b0 , w_9731 );
and ( w_9730 , w_9731 , \880_b0 );
or ( \3105_b1 , \3103_b1 , w_9732 );
or ( \3105_b0 , \3103_b0 , \3104_b0 );
not ( \3104_b0 , w_9733 );
and ( w_9733 , w_9732 , \3104_b1 );
or ( \3106_b1 , \894_b1 , \d[8]_b1 );
not ( \d[8]_b1 , w_9734 );
and ( \3106_b0 , \894_b0 , w_9735 );
and ( w_9734 , w_9735 , \d[8]_b0 );
or ( \3107_b1 , \c[8]_b1 , \909_b1 );
not ( \909_b1 , w_9736 );
and ( \3107_b0 , \c[8]_b0 , w_9737 );
and ( w_9736 , w_9737 , \909_b0 );
or ( \3108_b1 , \885_b1 , \b[8]_b1 );
not ( \b[8]_b1 , w_9738 );
and ( \3108_b0 , \885_b0 , w_9739 );
and ( w_9738 , w_9739 , \b[8]_b0 );
or ( \3110_b1 , \3105_b1 , w_9741 );
not ( w_9741 , w_9742 );
and ( \3110_b0 , \3105_b0 , w_9743 );
and ( w_9742 ,  , w_9743 );
buf ( w_9741 , \3109_b1 );
not ( w_9741 , w_9744 );
not (  , w_9745 );
and ( w_9744 , w_9745 , \3109_b0 );
buf ( \3111_b1 , \3110_b1 );
not ( \3111_b1 , w_9746 );
not ( \3111_b0 , w_9747 );
and ( w_9746 , w_9747 , \3110_b0 );
buf ( \3112_b1 , \752_b1 );
not ( \3112_b1 , w_9748 );
not ( \3112_b0 , w_9749 );
and ( w_9748 , w_9749 , \752_b0 );
or ( \3113_b1 , \3112_b1 , w_9751 );
not ( w_9751 , w_9752 );
and ( \3113_b0 , \3112_b0 , w_9753 );
and ( w_9752 ,  , w_9753 );
buf ( w_9751 , \763_b1 );
not ( w_9751 , w_9754 );
not (  , w_9755 );
and ( w_9754 , w_9755 , \763_b0 );
buf ( \3114_b1 , \3113_b1 );
not ( \3114_b1 , w_9756 );
not ( \3114_b0 , w_9757 );
and ( w_9756 , w_9757 , \3113_b0 );
buf ( \3115_b1 , \747_b1 );
not ( \3115_b1 , w_9758 );
not ( \3115_b0 , w_9759 );
and ( w_9758 , w_9759 , \747_b0 );
or ( \3116_b1 , \3114_b1 , w_9760 );
or ( \3116_b0 , \3114_b0 , \3115_b0 );
not ( \3115_b0 , w_9761 );
and ( w_9761 , w_9760 , \3115_b1 );
or ( \3117_b1 , \747_b1 , w_9762 );
or ( \3117_b0 , \747_b0 , \3113_b0 );
not ( \3113_b0 , w_9763 );
and ( w_9763 , w_9762 , \3113_b1 );
or ( \3118_b1 , \3116_b1 , w_9765 );
not ( w_9765 , w_9766 );
and ( \3118_b0 , \3116_b0 , w_9767 );
and ( w_9766 ,  , w_9767 );
buf ( w_9765 , \3117_b1 );
not ( w_9765 , w_9768 );
not (  , w_9769 );
and ( w_9768 , w_9769 , \3117_b0 );
or ( \3119_b1 , \3118_b1 , w_9771 );
not ( w_9771 , w_9772 );
and ( \3119_b0 , \3118_b0 , w_9773 );
and ( w_9772 ,  , w_9773 );
buf ( w_9771 , \707_b1 );
not ( w_9771 , w_9774 );
not (  , w_9775 );
and ( w_9774 , w_9775 , \707_b0 );
or ( \3120_b1 , \3111_b1 , w_9777 );
not ( w_9777 , w_9778 );
and ( \3120_b0 , \3111_b0 , w_9779 );
and ( w_9778 ,  , w_9779 );
buf ( w_9777 , \3119_b1 );
not ( w_9777 , w_9780 );
not (  , w_9781 );
and ( w_9780 , w_9781 , \3119_b0 );
or ( \3121_b1 , \3095_b1 , w_9783 );
not ( w_9783 , w_9784 );
and ( \3121_b0 , \3095_b0 , w_9785 );
and ( w_9784 ,  , w_9785 );
buf ( w_9783 , \3120_b1 );
not ( w_9783 , w_9786 );
not (  , w_9787 );
and ( w_9786 , w_9787 , \3120_b0 );
or ( \3122_b1 , \c[8]_b1 , \d[8]_b1 );
xor ( \3122_b0 , \c[8]_b0 , w_9788 );
not ( w_9788 , w_9789 );
and ( w_9789 , \d[8]_b1 , \d[8]_b0 );
or ( \3123_b1 , \2614_b1 , w_9791 );
not ( w_9791 , w_9792 );
and ( \3123_b0 , \2614_b0 , w_9793 );
and ( w_9792 ,  , w_9793 );
buf ( w_9791 , \3122_b1 );
not ( w_9791 , w_9794 );
not (  , w_9795 );
and ( w_9794 , w_9795 , \3122_b0 );
buf ( \3124_b1 , \2027_b1 );
buf ( \3124_b0 , \2027_b0 );
buf ( \3125_b1 , \2277_b1 );
buf ( \3125_b0 , \2277_b0 );
or ( \3126_b1 , \3124_b1 , w_9797 );
not ( w_9797 , w_9798 );
and ( \3126_b0 , \3124_b0 , w_9799 );
and ( w_9798 ,  , w_9799 );
buf ( w_9797 , \3125_b1 );
not ( w_9797 , w_9800 );
not (  , w_9801 );
and ( w_9800 , w_9801 , \3125_b0 );
buf ( \3127_b1 , \3126_b1 );
not ( \3127_b1 , w_9802 );
not ( \3127_b0 , w_9803 );
and ( w_9802 , w_9803 , \3126_b0 );
buf ( \3128_b1 , \2270_b1 );
not ( \3128_b1 , w_9804 );
not ( \3128_b0 , w_9805 );
and ( w_9804 , w_9805 , \2270_b0 );
or ( \3129_b1 , \3127_b1 , w_9806 );
or ( \3129_b0 , \3127_b0 , \3128_b0 );
not ( \3128_b0 , w_9807 );
and ( w_9807 , w_9806 , \3128_b1 );
or ( \3130_b1 , \2271_b1 , w_9808 );
or ( \3130_b0 , \2271_b0 , \3126_b0 );
not ( \3126_b0 , w_9809 );
and ( w_9809 , w_9808 , \3126_b1 );
or ( \3131_b1 , \3129_b1 , w_9811 );
not ( w_9811 , w_9812 );
and ( \3131_b0 , \3129_b0 , w_9813 );
and ( w_9812 ,  , w_9813 );
buf ( w_9811 , \3130_b1 );
not ( w_9811 , w_9814 );
not (  , w_9815 );
and ( w_9814 , w_9815 , \3130_b0 );
or ( \3132_b1 , \3131_b1 , w_9817 );
not ( w_9817 , w_9818 );
and ( \3132_b0 , \3131_b0 , w_9819 );
and ( w_9818 ,  , w_9819 );
buf ( w_9817 , \2413_b1 );
not ( w_9817 , w_9820 );
not (  , w_9821 );
and ( w_9820 , w_9821 , \2413_b0 );
or ( \3134_b1 , \3086_b1 , w_9823 );
not ( w_9823 , w_9824 );
and ( \3134_b0 , \3086_b0 , w_9825 );
and ( w_9824 ,  , w_9825 );
buf ( w_9823 , \3133_b1 );
not ( w_9823 , w_9826 );
not (  , w_9827 );
and ( w_9826 , w_9827 , \3133_b0 );
or ( \3135_b1 , \3083_b1 , w_9829 );
not ( w_9829 , w_9830 );
and ( \3135_b0 , \3083_b0 , w_9831 );
and ( w_9830 ,  , w_9831 );
buf ( w_9829 , \3134_b1 );
not ( w_9829 , w_9832 );
not (  , w_9833 );
and ( w_9832 , w_9833 , \3134_b0 );
or ( \3136_b1 , \3077_b1 , w_9835 );
not ( w_9835 , w_9836 );
and ( \3136_b0 , \3077_b0 , w_9837 );
and ( w_9836 ,  , w_9837 );
buf ( w_9835 , \3135_b1 );
not ( w_9835 , w_9838 );
not (  , w_9839 );
and ( w_9838 , w_9839 , \3135_b0 );
buf ( \3137_b1 , \689_b1 );
not ( \3137_b1 , w_9840 );
not ( \3137_b0 , w_9841 );
and ( w_9840 , w_9841 , \689_b0 );
buf ( \3138_b1 , \649_b1 );
not ( \3138_b1 , w_9842 );
not ( \3138_b0 , w_9843 );
and ( w_9842 , w_9843 , \649_b0 );
or ( \3139_b1 , \3137_b1 , w_9844 );
or ( \3139_b0 , \3137_b0 , \3138_b0 );
not ( \3138_b0 , w_9845 );
and ( w_9845 , w_9844 , \3138_b1 );
buf ( \3140_b1 , \b[12]_b1 );
not ( \3140_b1 , w_9846 );
not ( \3140_b0 , w_9847 );
and ( w_9846 , w_9847 , \b[12]_b0 );
buf ( \3141_b1 , \922_b1 );
not ( \3141_b1 , w_9848 );
not ( \3141_b0 , w_9849 );
and ( w_9848 , w_9849 , \922_b0 );
or ( \3142_b1 , \3140_b1 , w_9850 );
or ( \3142_b0 , \3140_b0 , \3141_b0 );
not ( \3141_b0 , w_9851 );
and ( w_9851 , w_9850 , \3141_b1 );
or ( \3143_b1 , \697_b1 , \687_b1 );
not ( \687_b1 , w_9852 );
and ( \3143_b0 , \697_b0 , w_9853 );
and ( w_9852 , w_9853 , \687_b0 );
or ( \3144_b1 , \3143_b1 , w_9855 );
not ( w_9855 , w_9856 );
and ( \3144_b0 , \3143_b0 , w_9857 );
and ( w_9856 ,  , w_9857 );
buf ( w_9855 , \909_b1 );
not ( w_9855 , w_9858 );
not (  , w_9859 );
and ( w_9858 , w_9859 , \909_b0 );
or ( \3145_b1 , \3142_b1 , w_9861 );
not ( w_9861 , w_9862 );
and ( \3145_b0 , \3142_b0 , w_9863 );
and ( w_9862 ,  , w_9863 );
buf ( w_9861 , \3144_b1 );
not ( w_9861 , w_9864 );
not (  , w_9865 );
and ( w_9864 , w_9865 , \3144_b0 );
or ( \3146_b1 , \3145_b1 , w_9867 );
not ( w_9867 , w_9868 );
and ( \3146_b0 , \3145_b0 , w_9869 );
and ( w_9868 ,  , w_9869 );
buf ( w_9867 , \c[12]_b1 );
not ( w_9867 , w_9870 );
not (  , w_9871 );
and ( w_9870 , w_9871 , \c[12]_b0 );
or ( \3147_b1 , \3139_b1 , w_9873 );
not ( w_9873 , w_9874 );
and ( \3147_b0 , \3139_b0 , w_9875 );
and ( w_9874 ,  , w_9875 );
buf ( w_9873 , \3146_b1 );
not ( w_9873 , w_9876 );
not (  , w_9877 );
and ( w_9876 , w_9877 , \3146_b0 );
or ( \3148_b1 , \2475_b1 , w_9879 );
not ( w_9879 , w_9880 );
and ( \3148_b0 , \2475_b0 , w_9881 );
and ( w_9880 ,  , w_9881 );
buf ( w_9879 , \a[12]_b1 );
not ( w_9879 , w_9882 );
not (  , w_9883 );
and ( w_9882 , w_9883 , \a[12]_b0 );
buf ( \3149_b1 , \b[12]_b1 );
not ( \3149_b1 , w_9884 );
not ( \3149_b0 , w_9885 );
and ( w_9884 , w_9885 , \b[12]_b0 );
buf ( \3150_b1 , \3149_b1 );
not ( \3150_b1 , w_9886 );
not ( \3150_b0 , w_9887 );
and ( w_9886 , w_9887 , \3149_b0 );
buf ( \3151_b1 , \688_b1 );
not ( \3151_b1 , w_9888 );
not ( \3151_b0 , w_9889 );
and ( w_9888 , w_9889 , \688_b0 );
or ( \3152_b1 , \3150_b1 , w_9890 );
or ( \3152_b0 , \3150_b0 , \3151_b0 );
not ( \3151_b0 , w_9891 );
and ( w_9891 , w_9890 , \3151_b1 );
or ( \3153_b1 , \3152_b1 , w_9893 );
not ( w_9893 , w_9894 );
and ( \3153_b0 , \3152_b0 , w_9895 );
and ( w_9894 ,  , w_9895 );
buf ( w_9893 , \667_b1 );
not ( w_9893 , w_9896 );
not (  , w_9897 );
and ( w_9896 , w_9897 , \667_b0 );
buf ( \3154_b1 , \c[12]_b1 );
not ( \3154_b1 , w_9898 );
not ( \3154_b0 , w_9899 );
and ( w_9898 , w_9899 , \c[12]_b0 );
buf ( \3155_b1 , \3154_b1 );
not ( \3155_b1 , w_9900 );
not ( \3155_b0 , w_9901 );
and ( w_9900 , w_9901 , \3154_b0 );
buf ( \3156_b1 , \697_b1 );
not ( \3156_b1 , w_9902 );
not ( \3156_b0 , w_9903 );
and ( w_9902 , w_9903 , \697_b0 );
or ( \3157_b1 , \3155_b1 , w_9904 );
or ( \3157_b0 , \3155_b0 , \3156_b0 );
not ( \3156_b0 , w_9905 );
and ( w_9905 , w_9904 , \3156_b1 );
or ( \3158_b1 , \3157_b1 , w_9907 );
not ( w_9907 , w_9908 );
and ( \3158_b0 , \3157_b0 , w_9909 );
and ( w_9908 ,  , w_9909 );
buf ( w_9907 , \893_b1 );
not ( w_9907 , w_9910 );
not (  , w_9911 );
and ( w_9910 , w_9911 , \893_b0 );
or ( \3159_b1 , \3158_b1 , \d[12]_b1 );
not ( \d[12]_b1 , w_9912 );
and ( \3159_b0 , \3158_b0 , w_9913 );
and ( w_9912 , w_9913 , \d[12]_b0 );
buf ( \3160_b1 , \758_b1 );
not ( \3160_b1 , w_9914 );
not ( \3160_b0 , w_9915 );
and ( w_9914 , w_9915 , \758_b0 );
or ( \3161_b1 , \3160_b1 , w_9917 );
not ( w_9917 , w_9918 );
and ( \3161_b0 , \3160_b0 , w_9919 );
and ( w_9918 ,  , w_9919 );
buf ( w_9917 , \779_b1 );
not ( w_9917 , w_9920 );
not (  , w_9921 );
and ( w_9920 , w_9921 , \779_b0 );
buf ( \3162_b1 , \3161_b1 );
not ( \3162_b1 , w_9922 );
not ( \3162_b0 , w_9923 );
and ( w_9922 , w_9923 , \3161_b0 );
buf ( \3163_b1 , \754_b1 );
not ( \3163_b1 , w_9924 );
not ( \3163_b0 , w_9925 );
and ( w_9924 , w_9925 , \754_b0 );
buf ( \3164_b1 , \747_b1 );
not ( \3164_b1 , w_9926 );
not ( \3164_b0 , w_9927 );
and ( w_9926 , w_9927 , \747_b0 );
or ( \3165_b1 , \3163_b1 , w_9928 );
or ( \3165_b0 , \3163_b0 , \3164_b0 );
not ( \3164_b0 , w_9929 );
and ( w_9929 , w_9928 , \3164_b1 );
or ( \3166_b1 , \3165_b1 , w_9931 );
not ( w_9931 , w_9932 );
and ( \3166_b0 , \3165_b0 , w_9933 );
and ( w_9932 ,  , w_9933 );
buf ( w_9931 , \777_b1 );
not ( w_9931 , w_9934 );
not (  , w_9935 );
and ( w_9934 , w_9935 , \777_b0 );
buf ( \3167_b1 , \3166_b1 );
not ( \3167_b1 , w_9936 );
not ( \3167_b0 , w_9937 );
and ( w_9936 , w_9937 , \3166_b0 );
or ( \3168_b1 , \3162_b1 , w_9938 );
or ( \3168_b0 , \3162_b0 , \3167_b0 );
not ( \3167_b0 , w_9939 );
and ( w_9939 , w_9938 , \3167_b1 );
or ( \3169_b1 , \3166_b1 , w_9940 );
or ( \3169_b0 , \3166_b0 , \3161_b0 );
not ( \3161_b0 , w_9941 );
and ( w_9941 , w_9940 , \3161_b1 );
or ( \3170_b1 , \3168_b1 , w_9943 );
not ( w_9943 , w_9944 );
and ( \3170_b0 , \3168_b0 , w_9945 );
and ( w_9944 ,  , w_9945 );
buf ( w_9943 , \3169_b1 );
not ( w_9943 , w_9946 );
not (  , w_9947 );
and ( w_9946 , w_9947 , \3169_b0 );
buf ( \3171_b1 , \3170_b1 );
not ( \3171_b1 , w_9948 );
not ( \3171_b0 , w_9949 );
and ( w_9948 , w_9949 , \3170_b0 );
buf ( \3172_b1 , \707_b1 );
not ( \3172_b1 , w_9950 );
not ( \3172_b0 , w_9951 );
and ( w_9950 , w_9951 , \707_b0 );
or ( \3173_b1 , \3171_b1 , w_9952 );
or ( \3173_b0 , \3171_b0 , \3172_b0 );
not ( \3172_b0 , w_9953 );
and ( w_9953 , w_9952 , \3172_b1 );
buf ( \3174_b1 , \886_b1 );
not ( \3174_b1 , w_9954 );
not ( \3174_b0 , w_9955 );
and ( w_9954 , w_9955 , \886_b0 );
buf ( \3175_b1 , \3149_b1 );
not ( \3175_b1 , w_9956 );
not ( \3175_b0 , w_9957 );
and ( w_9956 , w_9957 , \3149_b0 );
or ( \3176_b1 , \3174_b1 , \3175_b1 );
not ( \3175_b1 , w_9958 );
and ( \3176_b0 , \3174_b0 , w_9959 );
and ( w_9958 , w_9959 , \3175_b0 );
buf ( \3177_b1 , \843_b1 );
not ( \3177_b1 , w_9960 );
not ( \3177_b0 , w_9961 );
and ( w_9960 , w_9961 , \843_b0 );
or ( \3178_b1 , \3177_b1 , w_9963 );
not ( w_9963 , w_9964 );
and ( \3178_b0 , \3177_b0 , w_9965 );
and ( w_9964 ,  , w_9965 );
buf ( w_9963 , \864_b1 );
not ( w_9963 , w_9966 );
not (  , w_9967 );
and ( w_9966 , w_9967 , \864_b0 );
buf ( \3179_b1 , \3178_b1 );
not ( \3179_b1 , w_9968 );
not ( \3179_b0 , w_9969 );
and ( w_9968 , w_9969 , \3178_b0 );
buf ( \3180_b1 , \839_b1 );
not ( \3180_b1 , w_9970 );
not ( \3180_b0 , w_9971 );
and ( w_9970 , w_9971 , \839_b0 );
buf ( \3181_b1 , \832_b1 );
not ( \3181_b1 , w_9972 );
not ( \3181_b0 , w_9973 );
and ( w_9972 , w_9973 , \832_b0 );
or ( \3182_b1 , \3180_b1 , w_9974 );
or ( \3182_b0 , \3180_b0 , \3181_b0 );
not ( \3181_b0 , w_9975 );
and ( w_9975 , w_9974 , \3181_b1 );
or ( \3183_b1 , \3182_b1 , w_9977 );
not ( w_9977 , w_9978 );
and ( \3183_b0 , \3182_b0 , w_9979 );
and ( w_9978 ,  , w_9979 );
buf ( w_9977 , \862_b1 );
not ( w_9977 , w_9980 );
not (  , w_9981 );
and ( w_9980 , w_9981 , \862_b0 );
buf ( \3184_b1 , \3183_b1 );
not ( \3184_b1 , w_9982 );
not ( \3184_b0 , w_9983 );
and ( w_9982 , w_9983 , \3183_b0 );
or ( \3185_b1 , \3179_b1 , w_9984 );
or ( \3185_b0 , \3179_b0 , \3184_b0 );
not ( \3184_b0 , w_9985 );
and ( w_9985 , w_9984 , \3184_b1 );
or ( \3186_b1 , \3183_b1 , w_9986 );
or ( \3186_b0 , \3183_b0 , \3178_b0 );
not ( \3178_b0 , w_9987 );
and ( w_9987 , w_9986 , \3178_b1 );
or ( \3187_b1 , \3185_b1 , w_9989 );
not ( w_9989 , w_9990 );
and ( \3187_b0 , \3185_b0 , w_9991 );
and ( w_9990 ,  , w_9991 );
buf ( w_9989 , \3186_b1 );
not ( w_9989 , w_9992 );
not (  , w_9993 );
and ( w_9992 , w_9993 , \3186_b0 );
or ( \3188_b1 , \880_b1 , \3187_b1 );
not ( \3187_b1 , w_9994 );
and ( \3188_b0 , \880_b0 , w_9995 );
and ( w_9994 , w_9995 , \3187_b0 );
or ( \3189_b1 , \3176_b1 , w_9997 );
not ( w_9997 , w_9998 );
and ( \3189_b0 , \3176_b0 , w_9999 );
and ( w_9998 ,  , w_9999 );
buf ( w_9997 , \3188_b1 );
not ( w_9997 , w_10000 );
not (  , w_10001 );
and ( w_10000 , w_10001 , \3188_b0 );
or ( \3190_b1 , \3173_b1 , w_10003 );
not ( w_10003 , w_10004 );
and ( \3190_b0 , \3173_b0 , w_10005 );
and ( w_10004 ,  , w_10005 );
buf ( w_10003 , \3189_b1 );
not ( w_10003 , w_10006 );
not (  , w_10007 );
and ( w_10006 , w_10007 , \3189_b0 );
or ( \3191_b1 , \3159_b1 , w_10009 );
not ( w_10009 , w_10010 );
and ( \3191_b0 , \3159_b0 , w_10011 );
and ( w_10010 ,  , w_10011 );
buf ( w_10009 , \3190_b1 );
not ( w_10009 , w_10012 );
not (  , w_10013 );
and ( w_10012 , w_10013 , \3190_b0 );
or ( \3193_b1 , \3147_b1 , w_10015 );
not ( w_10015 , w_10016 );
and ( \3193_b0 , \3147_b0 , w_10017 );
and ( w_10016 ,  , w_10017 );
buf ( w_10015 , \3192_b1 );
not ( w_10015 , w_10018 );
not (  , w_10019 );
and ( w_10018 , w_10019 , \3192_b0 );
buf ( \3194_b1 , \a[0]_b1 );
not ( \3194_b1 , w_10020 );
not ( \3194_b0 , w_10021 );
and ( w_10020 , w_10021 , \a[0]_b0 );
buf ( \3195_b1 , \3072_b1 );
not ( \3195_b1 , w_10022 );
not ( \3195_b0 , w_10023 );
and ( w_10022 , w_10023 , \3072_b0 );
or ( \3196_b1 , \3195_b1 , w_10025 );
not ( w_10025 , w_10026 );
and ( \3196_b0 , \3195_b0 , w_10027 );
and ( w_10026 ,  , w_10027 );
buf ( w_10025 , \3074_b1 );
not ( w_10025 , w_10028 );
not (  , w_10029 );
and ( w_10028 , w_10029 , \3074_b0 );
buf ( \3197_b1 , \3196_b1 );
not ( \3197_b1 , w_10030 );
not ( \3197_b0 , w_10031 );
and ( w_10030 , w_10031 , \3196_b0 );
or ( \3198_b1 , \3194_b1 , w_10032 );
or ( \3198_b0 , \3194_b0 , \3197_b0 );
not ( \3197_b0 , w_10033 );
and ( w_10033 , w_10032 , \3197_b1 );
buf ( \3199_b1 , \c[0]_b1 );
not ( \3199_b1 , w_10034 );
not ( \3199_b0 , w_10035 );
and ( w_10034 , w_10035 , \c[0]_b0 );
buf ( \3200_b1 , \b[0]_b1 );
not ( \3200_b1 , w_10036 );
not ( \3200_b0 , w_10037 );
and ( w_10036 , w_10037 , \b[0]_b0 );
buf ( \3201_b1 , \2887_b1 );
not ( \3201_b1 , w_10038 );
not ( \3201_b0 , w_10039 );
and ( w_10038 , w_10039 , \2887_b0 );
or ( \3202_b1 , \3200_b1 , w_10040 );
or ( \3202_b0 , \3200_b0 , \3201_b0 );
not ( \3201_b0 , w_10041 );
and ( w_10041 , w_10040 , \3201_b1 );
buf ( \3203_b1 , \d[0]_b1 );
not ( \3203_b1 , w_10042 );
not ( \3203_b0 , w_10043 );
and ( w_10042 , w_10043 , \d[0]_b0 );
or ( \3204_b1 , \903_b1 , \3203_b1 );
not ( \3203_b1 , w_10044 );
and ( \3204_b0 , \903_b0 , w_10045 );
and ( w_10044 , w_10045 , \3203_b0 );
or ( \3205_b1 , \3204_b1 , w_10047 );
not ( w_10047 , w_10048 );
and ( \3205_b0 , \3204_b0 , w_10049 );
and ( w_10048 ,  , w_10049 );
buf ( w_10047 , \909_b1 );
not ( w_10047 , w_10050 );
not (  , w_10051 );
and ( w_10050 , w_10051 , \909_b0 );
or ( \3206_b1 , \3202_b1 , w_10053 );
not ( w_10053 , w_10054 );
and ( \3206_b0 , \3202_b0 , w_10055 );
and ( w_10054 ,  , w_10055 );
buf ( w_10053 , \3205_b1 );
not ( w_10053 , w_10056 );
not (  , w_10057 );
and ( w_10056 , w_10057 , \3205_b0 );
buf ( \3207_b1 , \3206_b1 );
not ( \3207_b1 , w_10058 );
not ( \3207_b0 , w_10059 );
and ( w_10058 , w_10059 , \3206_b0 );
or ( \3208_b1 , \3199_b1 , w_10060 );
or ( \3208_b0 , \3199_b0 , \3207_b0 );
not ( \3207_b0 , w_10061 );
and ( w_10061 , w_10060 , \3207_b1 );
buf ( \3209_b1 , \c[0]_b1 );
not ( \3209_b1 , w_10062 );
not ( \3209_b0 , w_10063 );
and ( w_10062 , w_10063 , \c[0]_b0 );
buf ( \3210_b1 , \3209_b1 );
not ( \3210_b1 , w_10064 );
not ( \3210_b0 , w_10065 );
and ( w_10064 , w_10065 , \3209_b0 );
buf ( \3211_b1 , \903_b1 );
not ( \3211_b1 , w_10066 );
not ( \3211_b0 , w_10067 );
and ( w_10066 , w_10067 , \903_b0 );
or ( \3212_b1 , \3210_b1 , w_10068 );
or ( \3212_b0 , \3210_b0 , \3211_b0 );
not ( \3211_b0 , w_10069 );
and ( w_10069 , w_10068 , \3211_b1 );
or ( \3213_b1 , \3212_b1 , w_10071 );
not ( w_10071 , w_10072 );
and ( \3213_b0 , \3212_b0 , w_10073 );
and ( w_10072 ,  , w_10073 );
buf ( w_10071 , \893_b1 );
not ( w_10071 , w_10074 );
not (  , w_10075 );
and ( w_10074 , w_10075 , \893_b0 );
or ( \3214_b1 , \3213_b1 , \d[0]_b1 );
not ( \d[0]_b1 , w_10076 );
and ( \3214_b0 , \3213_b0 , w_10077 );
and ( w_10076 , w_10077 , \d[0]_b0 );
buf ( \3215_b1 , \2220_b1 );
not ( \3215_b1 , w_10078 );
not ( \3215_b0 , w_10079 );
and ( w_10078 , w_10079 , \2220_b0 );
buf ( \3216_b1 , \3215_b1 );
not ( \3216_b1 , w_10080 );
not ( \3216_b0 , w_10081 );
and ( w_10080 , w_10081 , \3215_b0 );
buf ( \3217_b1 , \2413_b1 );
not ( \3217_b1 , w_10082 );
not ( \3217_b0 , w_10083 );
and ( w_10082 , w_10083 , \2413_b0 );
or ( \3218_b1 , \3216_b1 , w_10084 );
or ( \3218_b0 , \3216_b0 , \3217_b0 );
not ( \3217_b0 , w_10085 );
and ( w_10085 , w_10084 , \3217_b1 );
buf ( \3219_b1 , \684_b1 );
not ( \3219_b1 , w_10086 );
not ( \3219_b0 , w_10087 );
and ( w_10086 , w_10087 , \684_b0 );
or ( \3220_b1 , \1668_b1 , \3219_b1 );
not ( \3219_b1 , w_10088 );
and ( \3220_b0 , \1668_b0 , w_10089 );
and ( w_10088 , w_10089 , \3219_b0 );
or ( \3221_b1 , \b[0]_b1 , \d[0]_b1 );
xor ( \3221_b0 , \b[0]_b0 , w_10090 );
not ( w_10090 , w_10091 );
and ( w_10091 , \d[0]_b1 , \d[0]_b0 );
buf ( \3222_b1 , \3221_b1 );
not ( \3222_b1 , w_10092 );
not ( \3222_b0 , w_10093 );
and ( w_10092 , w_10093 , \3221_b0 );
buf ( \3223_b1 , \707_b1 );
not ( \3223_b1 , w_10094 );
not ( \3223_b0 , w_10095 );
and ( w_10094 , w_10095 , \707_b0 );
or ( \3224_b1 , \3222_b1 , w_10096 );
or ( \3224_b0 , \3222_b0 , \3223_b0 );
not ( \3223_b0 , w_10097 );
and ( w_10097 , w_10096 , \3223_b1 );
or ( \3225_b1 , \a[0]_b1 , \c[0]_b1 );
xor ( \3225_b0 , \a[0]_b0 , w_10098 );
not ( w_10098 , w_10099 );
and ( w_10099 , \c[0]_b1 , \c[0]_b0 );
or ( \3226_b1 , \880_b1 , \3225_b1 );
not ( \3225_b1 , w_10100 );
and ( \3226_b0 , \880_b0 , w_10101 );
and ( w_10100 , w_10101 , \3225_b0 );
or ( \3227_b1 , \885_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_10102 );
and ( \3227_b0 , \885_b0 , w_10103 );
and ( w_10102 , w_10103 , \b[0]_b0 );
or ( \3228_b1 , \3226_b1 , w_10105 );
not ( w_10105 , w_10106 );
and ( \3228_b0 , \3226_b0 , w_10107 );
and ( w_10106 ,  , w_10107 );
buf ( w_10105 , \3227_b1 );
not ( w_10105 , w_10108 );
not (  , w_10109 );
and ( w_10108 , w_10109 , \3227_b0 );
or ( \3229_b1 , \3224_b1 , w_10111 );
not ( w_10111 , w_10112 );
and ( \3229_b0 , \3224_b0 , w_10113 );
and ( w_10112 ,  , w_10113 );
buf ( w_10111 , \3228_b1 );
not ( w_10111 , w_10114 );
not (  , w_10115 );
and ( w_10114 , w_10115 , \3228_b0 );
or ( \3230_b1 , \3220_b1 , w_10117 );
not ( w_10117 , w_10118 );
and ( \3230_b0 , \3220_b0 , w_10119 );
and ( w_10118 ,  , w_10119 );
buf ( w_10117 , \3229_b1 );
not ( w_10117 , w_10120 );
not (  , w_10121 );
and ( w_10120 , w_10121 , \3229_b0 );
or ( \3231_b1 , \3218_b1 , w_10123 );
not ( w_10123 , w_10124 );
and ( \3231_b0 , \3218_b0 , w_10125 );
and ( w_10124 ,  , w_10125 );
buf ( w_10123 , \3230_b1 );
not ( w_10123 , w_10126 );
not (  , w_10127 );
and ( w_10126 , w_10127 , \3230_b0 );
or ( \3232_b1 , \3214_b1 , w_10129 );
not ( w_10129 , w_10130 );
and ( \3232_b0 , \3214_b0 , w_10131 );
and ( w_10130 ,  , w_10131 );
buf ( w_10129 , \3231_b1 );
not ( w_10129 , w_10132 );
not (  , w_10133 );
and ( w_10132 , w_10133 , \3231_b0 );
or ( \3233_b1 , \3208_b1 , w_10135 );
not ( w_10135 , w_10136 );
and ( \3233_b0 , \3208_b0 , w_10137 );
and ( w_10136 ,  , w_10137 );
buf ( w_10135 , \3232_b1 );
not ( w_10135 , w_10138 );
not (  , w_10139 );
and ( w_10138 , w_10139 , \3232_b0 );
buf ( \3234_b1 , \d[0]_b1 );
not ( \3234_b1 , w_10140 );
not ( \3234_b0 , w_10141 );
and ( w_10140 , w_10141 , \d[0]_b0 );
buf ( \3235_b1 , \648_b1 );
buf ( \3235_b0 , \648_b0 );
buf ( \3236_b1 , \3235_b1 );
not ( \3236_b1 , w_10142 );
not ( \3236_b0 , w_10143 );
and ( w_10142 , w_10143 , \3235_b0 );
or ( \3237_b1 , \3234_b1 , w_10144 );
or ( \3237_b0 , \3234_b0 , \3236_b0 );
not ( \3236_b0 , w_10145 );
and ( w_10145 , w_10144 , \3236_b1 );
or ( \3238_b1 , \2791_b1 , w_10147 );
not ( w_10147 , w_10148 );
and ( \3238_b0 , \2791_b0 , w_10149 );
and ( w_10148 ,  , w_10149 );
buf ( w_10147 , \b[0]_b1 );
not ( w_10147 , w_10150 );
not (  , w_10151 );
and ( w_10150 , w_10151 , \b[0]_b0 );
or ( \3239_b1 , \3237_b1 , w_10153 );
not ( w_10153 , w_10154 );
and ( \3239_b0 , \3237_b0 , w_10155 );
and ( w_10154 ,  , w_10155 );
buf ( w_10153 , \3238_b1 );
not ( w_10153 , w_10156 );
not (  , w_10157 );
and ( w_10156 , w_10157 , \3238_b0 );
or ( \3240_b1 , \3233_b1 , w_10159 );
not ( w_10159 , w_10160 );
and ( \3240_b0 , \3233_b0 , w_10161 );
and ( w_10160 ,  , w_10161 );
buf ( w_10159 , \3239_b1 );
not ( w_10159 , w_10162 );
not (  , w_10163 );
and ( w_10162 , w_10163 , \3239_b0 );
or ( \3241_b1 , \3198_b1 , w_10165 );
not ( w_10165 , w_10166 );
and ( \3241_b0 , \3198_b0 , w_10167 );
and ( w_10166 ,  , w_10167 );
buf ( w_10165 , \3240_b1 );
not ( w_10165 , w_10168 );
not (  , w_10169 );
and ( w_10168 , w_10169 , \3240_b0 );
buf ( \3242_b1 , \a[7]_b1 );
not ( \3242_b1 , w_10170 );
not ( \3242_b0 , w_10171 );
and ( w_10170 , w_10171 , \a[7]_b0 );
buf ( \3243_b1 , \3075_b1 );
not ( \3243_b1 , w_10172 );
not ( \3243_b0 , w_10173 );
and ( w_10172 , w_10173 , \3075_b0 );
or ( \3244_b1 , \3242_b1 , w_10174 );
or ( \3244_b0 , \3242_b0 , \3243_b0 );
not ( \3243_b0 , w_10175 );
and ( w_10175 , w_10174 , \3243_b1 );
buf ( \3245_b1 , \d[7]_b1 );
not ( \3245_b1 , w_10176 );
not ( \3245_b0 , w_10177 );
and ( w_10176 , w_10177 , \d[7]_b0 );
buf ( \3246_b1 , \648_b1 );
not ( \3246_b1 , w_10178 );
not ( \3246_b0 , w_10179 );
and ( w_10178 , w_10179 , \648_b0 );
or ( \3247_b1 , \3245_b1 , w_10180 );
or ( \3247_b0 , \3245_b0 , \3246_b0 );
not ( \3246_b0 , w_10181 );
and ( w_10181 , w_10180 , \3246_b1 );
or ( \3248_b1 , \667_b1 , w_10183 );
not ( w_10183 , w_10184 );
and ( \3248_b0 , \667_b0 , w_10185 );
and ( w_10184 ,  , w_10185 );
buf ( w_10183 , \b[7]_b1 );
not ( w_10183 , w_10186 );
not (  , w_10187 );
and ( w_10186 , w_10187 , \b[7]_b0 );
or ( \3249_b1 , \3247_b1 , w_10189 );
not ( w_10189 , w_10190 );
and ( \3249_b0 , \3247_b0 , w_10191 );
and ( w_10190 ,  , w_10191 );
buf ( w_10189 , \3248_b1 );
not ( w_10189 , w_10192 );
not (  , w_10193 );
and ( w_10192 , w_10193 , \3248_b0 );
or ( \3250_b1 , \b[7]_b1 , \c[7]_b1 );
not ( \c[7]_b1 , w_10194 );
and ( \3250_b0 , \b[7]_b0 , w_10195 );
and ( w_10194 , w_10195 , \c[7]_b0 );
buf ( \3251_b1 , \3250_b1 );
not ( \3251_b1 , w_10196 );
not ( \3251_b0 , w_10197 );
and ( w_10196 , w_10197 , \3250_b0 );
buf ( \3252_b1 , \922_b1 );
not ( \3252_b1 , w_10198 );
not ( \3252_b0 , w_10199 );
and ( w_10198 , w_10199 , \922_b0 );
or ( \3253_b1 , \3251_b1 , w_10200 );
or ( \3253_b0 , \3251_b0 , \3252_b0 );
not ( \3252_b0 , w_10201 );
and ( w_10201 , w_10200 , \3252_b1 );
or ( \3254_b1 , \c[7]_b1 , \d[7]_b1 );
xor ( \3254_b0 , \c[7]_b0 , w_10202 );
not ( w_10202 , w_10203 );
and ( w_10203 , \d[7]_b1 , \d[7]_b0 );
or ( \3255_b1 , \2615_b1 , \3254_b1 );
not ( \3254_b1 , w_10204 );
and ( \3255_b0 , \2615_b0 , w_10205 );
and ( w_10204 , w_10205 , \3254_b0 );
or ( \3256_b1 , \2269_b1 , w_10207 );
not ( w_10207 , w_10208 );
and ( \3256_b0 , \2269_b0 , w_10209 );
and ( w_10208 ,  , w_10209 );
buf ( w_10207 , \2158_b1 );
not ( w_10207 , w_10210 );
not (  , w_10211 );
and ( w_10210 , w_10211 , \2158_b0 );
or ( \3257_b1 , \2264_b1 , w_10212 );
xor ( \3257_b0 , \2264_b0 , w_10214 );
not ( w_10214 , w_10215 );
and ( w_10215 , w_10212 , w_10213 );
buf ( w_10212 , \3256_b1 );
not ( w_10212 , w_10216 );
not ( w_10213 , w_10217 );
and ( w_10216 , w_10217 , \3256_b0 );
buf ( \3258_b1 , \3257_b1 );
not ( \3258_b1 , w_10218 );
not ( \3258_b0 , w_10219 );
and ( w_10218 , w_10219 , \3257_b0 );
buf ( \3259_b1 , \2413_b1 );
not ( \3259_b1 , w_10220 );
not ( \3259_b0 , w_10221 );
and ( w_10220 , w_10221 , \2413_b0 );
or ( \3260_b1 , \3258_b1 , w_10222 );
or ( \3260_b0 , \3258_b0 , \3259_b0 );
not ( \3259_b0 , w_10223 );
and ( w_10223 , w_10222 , \3259_b1 );
buf ( \3261_b1 , \1523_b1 );
buf ( \3261_b0 , \1523_b0 );
buf ( \3262_b1 , \3261_b1 );
not ( \3262_b1 , w_10224 );
not ( \3262_b0 , w_10225 );
and ( w_10224 , w_10225 , \3261_b0 );
or ( \3263_b1 , \1526_b1 , w_10227 );
not ( w_10227 , w_10228 );
and ( \3263_b0 , \1526_b0 , w_10229 );
and ( w_10228 ,  , w_10229 );
buf ( w_10227 , \1417_b1 );
not ( w_10227 , w_10230 );
not (  , w_10231 );
and ( w_10230 , w_10231 , \1417_b0 );
buf ( \3264_b1 , \3263_b1 );
not ( \3264_b1 , w_10232 );
not ( \3264_b0 , w_10233 );
and ( w_10232 , w_10233 , \3263_b0 );
or ( \3265_b1 , \3262_b1 , w_10234 );
or ( \3265_b0 , \3262_b0 , \3264_b0 );
not ( \3264_b0 , w_10235 );
and ( w_10235 , w_10234 , \3264_b1 );
or ( \3266_b1 , \3263_b1 , w_10236 );
or ( \3266_b0 , \3263_b0 , \3261_b0 );
not ( \3261_b0 , w_10237 );
and ( w_10237 , w_10236 , \3261_b1 );
or ( \3267_b1 , \3265_b1 , w_10239 );
not ( w_10239 , w_10240 );
and ( \3267_b0 , \3265_b0 , w_10241 );
and ( w_10240 ,  , w_10241 );
buf ( w_10239 , \3266_b1 );
not ( w_10239 , w_10242 );
not (  , w_10243 );
and ( w_10242 , w_10243 , \3266_b0 );
or ( \3268_b1 , \2908_b1 , \3267_b1 );
not ( \3267_b1 , w_10244 );
and ( \3268_b0 , \2908_b0 , w_10245 );
and ( w_10244 , w_10245 , \3267_b0 );
buf ( \3269_b1 , \729_b1 );
not ( \3269_b1 , w_10246 );
not ( \3269_b0 , w_10247 );
and ( w_10246 , w_10247 , \729_b0 );
or ( \3270_b1 , \3269_b1 , w_10249 );
not ( w_10249 , w_10250 );
and ( \3270_b0 , \3269_b0 , w_10251 );
and ( w_10250 ,  , w_10251 );
buf ( w_10249 , \736_b1 );
not ( w_10249 , w_10252 );
not (  , w_10253 );
and ( w_10252 , w_10253 , \736_b0 );
buf ( \3271_b1 , \3270_b1 );
not ( \3271_b1 , w_10254 );
not ( \3271_b0 , w_10255 );
and ( w_10254 , w_10255 , \3270_b0 );
or ( \3272_b1 , \732_b1 , w_10257 );
not ( w_10257 , w_10258 );
and ( \3272_b0 , \732_b0 , w_10259 );
and ( w_10258 ,  , w_10259 );
buf ( w_10257 , \718_b1 );
not ( w_10257 , w_10260 );
not (  , w_10261 );
and ( w_10260 , w_10261 , \718_b0 );
or ( \3273_b1 , \2979_b1 , \3272_b1 );
not ( \3272_b1 , w_10262 );
and ( \3273_b0 , \2979_b0 , w_10263 );
and ( w_10262 , w_10263 , \3272_b0 );
or ( \3274_b1 , \732_b1 , w_10264 );
or ( \3274_b0 , \732_b0 , \722_b0 );
not ( \722_b0 , w_10265 );
and ( w_10265 , w_10264 , \722_b1 );
or ( \3275_b1 , \3274_b1 , w_10267 );
not ( w_10267 , w_10268 );
and ( \3275_b0 , \3274_b0 , w_10269 );
and ( w_10268 ,  , w_10269 );
buf ( w_10267 , \721_b1 );
not ( w_10267 , w_10270 );
not (  , w_10271 );
and ( w_10270 , w_10271 , \721_b0 );
or ( \3276_b1 , \3273_b1 , w_10273 );
not ( w_10273 , w_10274 );
and ( \3276_b0 , \3273_b0 , w_10275 );
and ( w_10274 ,  , w_10275 );
buf ( w_10273 , \3275_b1 );
not ( w_10273 , w_10276 );
not (  , w_10277 );
and ( w_10276 , w_10277 , \3275_b0 );
buf ( \3277_b1 , \728_b1 );
not ( \3277_b1 , w_10278 );
not ( \3277_b0 , w_10279 );
and ( w_10278 , w_10279 , \728_b0 );
or ( \3278_b1 , \3277_b1 , w_10281 );
not ( w_10281 , w_10282 );
and ( \3278_b0 , \3277_b0 , w_10283 );
and ( w_10282 ,  , w_10283 );
buf ( w_10281 , \727_b1 );
not ( w_10281 , w_10284 );
not (  , w_10285 );
and ( w_10284 , w_10285 , \727_b0 );
or ( \3279_b1 , \3276_b1 , w_10286 );
or ( \3279_b0 , \3276_b0 , \3278_b0 );
not ( \3278_b0 , w_10287 );
and ( w_10287 , w_10286 , \3278_b1 );
or ( \3280_b1 , \744_b1 , \742_b1 );
not ( \742_b1 , w_10288 );
and ( \3280_b0 , \744_b0 , w_10289 );
and ( w_10288 , w_10289 , \742_b0 );
or ( \3281_b1 , \728_b1 , w_10290 );
or ( \3281_b0 , \728_b0 , \3280_b0 );
not ( \3280_b0 , w_10291 );
and ( w_10291 , w_10290 , \3280_b1 );
buf ( \3283_b1 , \3282_b1 );
not ( \3283_b1 , w_10292 );
not ( \3283_b0 , w_10293 );
and ( w_10292 , w_10293 , \3282_b0 );
or ( \3284_b1 , \3271_b1 , w_10294 );
or ( \3284_b0 , \3271_b0 , \3283_b0 );
not ( \3283_b0 , w_10295 );
and ( w_10295 , w_10294 , \3283_b1 );
or ( \3285_b1 , \3282_b1 , w_10296 );
or ( \3285_b0 , \3282_b0 , \3270_b0 );
not ( \3270_b0 , w_10297 );
and ( w_10297 , w_10296 , \3270_b1 );
or ( \3286_b1 , \3284_b1 , w_10299 );
not ( w_10299 , w_10300 );
and ( \3286_b0 , \3284_b0 , w_10301 );
and ( w_10300 ,  , w_10301 );
buf ( w_10299 , \3285_b1 );
not ( w_10299 , w_10302 );
not (  , w_10303 );
and ( w_10302 , w_10303 , \3285_b0 );
buf ( \3287_b1 , \3286_b1 );
not ( \3287_b1 , w_10304 );
not ( \3287_b0 , w_10305 );
and ( w_10304 , w_10305 , \3286_b0 );
buf ( \3288_b1 , \707_b1 );
not ( \3288_b1 , w_10306 );
not ( \3288_b0 , w_10307 );
and ( w_10306 , w_10307 , \707_b0 );
or ( \3289_b1 , \3287_b1 , w_10308 );
or ( \3289_b0 , \3287_b0 , \3288_b0 );
not ( \3288_b0 , w_10309 );
and ( w_10309 , w_10308 , \3288_b1 );
buf ( \3290_b1 , \814_b1 );
not ( \3290_b1 , w_10310 );
not ( \3290_b0 , w_10311 );
and ( w_10310 , w_10311 , \814_b0 );
or ( \3291_b1 , \3290_b1 , w_10313 );
not ( w_10313 , w_10314 );
and ( \3291_b0 , \3290_b0 , w_10315 );
and ( w_10314 ,  , w_10315 );
buf ( w_10313 , \821_b1 );
not ( w_10313 , w_10316 );
not (  , w_10317 );
and ( w_10316 , w_10317 , \821_b0 );
buf ( \3292_b1 , \3291_b1 );
not ( \3292_b1 , w_10318 );
not ( \3292_b0 , w_10319 );
and ( w_10318 , w_10319 , \3291_b0 );
or ( \3293_b1 , \817_b1 , w_10321 );
not ( w_10321 , w_10322 );
and ( \3293_b0 , \817_b0 , w_10323 );
and ( w_10322 ,  , w_10323 );
buf ( w_10321 , \803_b1 );
not ( w_10321 , w_10324 );
not (  , w_10325 );
and ( w_10324 , w_10325 , \803_b0 );
or ( \3294_b1 , \2991_b1 , \3293_b1 );
not ( \3293_b1 , w_10326 );
and ( \3294_b0 , \2991_b0 , w_10327 );
and ( w_10326 , w_10327 , \3293_b0 );
or ( \3295_b1 , \817_b1 , w_10328 );
or ( \3295_b0 , \817_b0 , \807_b0 );
not ( \807_b0 , w_10329 );
and ( w_10329 , w_10328 , \807_b1 );
or ( \3296_b1 , \3295_b1 , w_10331 );
not ( w_10331 , w_10332 );
and ( \3296_b0 , \3295_b0 , w_10333 );
and ( w_10332 ,  , w_10333 );
buf ( w_10331 , \806_b1 );
not ( w_10331 , w_10334 );
not (  , w_10335 );
and ( w_10334 , w_10335 , \806_b0 );
or ( \3297_b1 , \3294_b1 , w_10337 );
not ( w_10337 , w_10338 );
and ( \3297_b0 , \3294_b0 , w_10339 );
and ( w_10338 ,  , w_10339 );
buf ( w_10337 , \3296_b1 );
not ( w_10337 , w_10340 );
not (  , w_10341 );
and ( w_10340 , w_10341 , \3296_b0 );
buf ( \3298_b1 , \813_b1 );
not ( \3298_b1 , w_10342 );
not ( \3298_b0 , w_10343 );
and ( w_10342 , w_10343 , \813_b0 );
or ( \3299_b1 , \3298_b1 , w_10345 );
not ( w_10345 , w_10346 );
and ( \3299_b0 , \3298_b0 , w_10347 );
and ( w_10346 ,  , w_10347 );
buf ( w_10345 , \812_b1 );
not ( w_10345 , w_10348 );
not (  , w_10349 );
and ( w_10348 , w_10349 , \812_b0 );
or ( \3300_b1 , \3297_b1 , w_10350 );
or ( \3300_b0 , \3297_b0 , \3299_b0 );
not ( \3299_b0 , w_10351 );
and ( w_10351 , w_10350 , \3299_b1 );
or ( \3301_b1 , \829_b1 , \827_b1 );
not ( \827_b1 , w_10352 );
and ( \3301_b0 , \829_b0 , w_10353 );
and ( w_10352 , w_10353 , \827_b0 );
or ( \3302_b1 , \813_b1 , w_10354 );
or ( \3302_b0 , \813_b0 , \3301_b0 );
not ( \3301_b0 , w_10355 );
and ( w_10355 , w_10354 , \3301_b1 );
buf ( \3304_b1 , \3303_b1 );
not ( \3304_b1 , w_10356 );
not ( \3304_b0 , w_10357 );
and ( w_10356 , w_10357 , \3303_b0 );
or ( \3305_b1 , \3292_b1 , w_10358 );
or ( \3305_b0 , \3292_b0 , \3304_b0 );
not ( \3304_b0 , w_10359 );
and ( w_10359 , w_10358 , \3304_b1 );
or ( \3306_b1 , \3303_b1 , w_10360 );
or ( \3306_b0 , \3303_b0 , \3291_b0 );
not ( \3291_b0 , w_10361 );
and ( w_10361 , w_10360 , \3291_b1 );
or ( \3307_b1 , \3305_b1 , w_10363 );
not ( w_10363 , w_10364 );
and ( \3307_b0 , \3305_b0 , w_10365 );
and ( w_10364 ,  , w_10365 );
buf ( w_10363 , \3306_b1 );
not ( w_10363 , w_10366 );
not (  , w_10367 );
and ( w_10366 , w_10367 , \3306_b0 );
or ( \3308_b1 , \880_b1 , \3307_b1 );
not ( \3307_b1 , w_10368 );
and ( \3308_b0 , \880_b0 , w_10369 );
and ( w_10368 , w_10369 , \3307_b0 );
buf ( \3309_b1 , \d[7]_b1 );
not ( \3309_b1 , w_10370 );
not ( \3309_b0 , w_10371 );
and ( w_10370 , w_10371 , \d[7]_b0 );
buf ( \3310_b1 , \894_b1 );
not ( \3310_b1 , w_10372 );
not ( \3310_b0 , w_10373 );
and ( w_10372 , w_10373 , \894_b0 );
or ( \3311_b1 , \3309_b1 , w_10374 );
or ( \3311_b0 , \3309_b0 , \3310_b0 );
not ( \3310_b0 , w_10375 );
and ( w_10375 , w_10374 , \3310_b1 );
buf ( \3312_b1 , \886_b1 );
not ( \3312_b1 , w_10376 );
not ( \3312_b0 , w_10377 );
and ( w_10376 , w_10377 , \886_b0 );
buf ( \3313_b1 , \b[7]_b1 );
not ( \3313_b1 , w_10378 );
not ( \3313_b0 , w_10379 );
and ( w_10378 , w_10379 , \b[7]_b0 );
buf ( \3314_b1 , \3313_b1 );
not ( \3314_b1 , w_10380 );
not ( \3314_b0 , w_10381 );
and ( w_10380 , w_10381 , \3313_b0 );
or ( \3315_b1 , \3312_b1 , \3314_b1 );
not ( \3314_b1 , w_10382 );
and ( \3315_b0 , \3312_b0 , w_10383 );
and ( w_10382 , w_10383 , \3314_b0 );
or ( \3316_b1 , \907_b1 , \c[7]_b1 );
not ( \c[7]_b1 , w_10384 );
and ( \3316_b0 , \907_b0 , w_10385 );
and ( w_10384 , w_10385 , \c[7]_b0 );
or ( \3317_b1 , \3315_b1 , w_10387 );
not ( w_10387 , w_10388 );
and ( \3317_b0 , \3315_b0 , w_10389 );
and ( w_10388 ,  , w_10389 );
buf ( w_10387 , \3316_b1 );
not ( w_10387 , w_10390 );
not (  , w_10391 );
and ( w_10390 , w_10391 , \3316_b0 );
or ( \3318_b1 , \3311_b1 , w_10393 );
not ( w_10393 , w_10394 );
and ( \3318_b0 , \3311_b0 , w_10395 );
and ( w_10394 ,  , w_10395 );
buf ( w_10393 , \3317_b1 );
not ( w_10393 , w_10396 );
not (  , w_10397 );
and ( w_10396 , w_10397 , \3317_b0 );
or ( \3319_b1 , \3308_b1 , w_10399 );
not ( w_10399 , w_10400 );
and ( \3319_b0 , \3308_b0 , w_10401 );
and ( w_10400 ,  , w_10401 );
buf ( w_10399 , \3318_b1 );
not ( w_10399 , w_10402 );
not (  , w_10403 );
and ( w_10402 , w_10403 , \3318_b0 );
or ( \3320_b1 , \3289_b1 , w_10405 );
not ( w_10405 , w_10406 );
and ( \3320_b0 , \3289_b0 , w_10407 );
and ( w_10406 ,  , w_10407 );
buf ( w_10405 , \3319_b1 );
not ( w_10405 , w_10408 );
not (  , w_10409 );
and ( w_10408 , w_10409 , \3319_b0 );
or ( \3321_b1 , \3268_b1 , w_10411 );
not ( w_10411 , w_10412 );
and ( \3321_b0 , \3268_b0 , w_10413 );
and ( w_10412 ,  , w_10413 );
buf ( w_10411 , \3320_b1 );
not ( w_10411 , w_10414 );
not (  , w_10415 );
and ( w_10414 , w_10415 , \3320_b0 );
or ( \3322_b1 , \3260_b1 , w_10417 );
not ( w_10417 , w_10418 );
and ( \3322_b0 , \3260_b0 , w_10419 );
and ( w_10418 ,  , w_10419 );
buf ( w_10417 , \3321_b1 );
not ( w_10417 , w_10420 );
not (  , w_10421 );
and ( w_10420 , w_10421 , \3321_b0 );
or ( \3323_b1 , \3255_b1 , w_10423 );
not ( w_10423 , w_10424 );
and ( \3323_b0 , \3255_b0 , w_10425 );
and ( w_10424 ,  , w_10425 );
buf ( w_10423 , \3322_b1 );
not ( w_10423 , w_10426 );
not (  , w_10427 );
and ( w_10426 , w_10427 , \3322_b0 );
or ( \3324_b1 , \3253_b1 , w_10429 );
not ( w_10429 , w_10430 );
and ( \3324_b0 , \3253_b0 , w_10431 );
and ( w_10430 ,  , w_10431 );
buf ( w_10429 , \3323_b1 );
not ( w_10429 , w_10432 );
not (  , w_10433 );
and ( w_10432 , w_10433 , \3323_b0 );
or ( \3325_b1 , \3249_b1 , w_10435 );
not ( w_10435 , w_10436 );
and ( \3325_b0 , \3249_b0 , w_10437 );
and ( w_10436 ,  , w_10437 );
buf ( w_10435 , \3324_b1 );
not ( w_10435 , w_10438 );
not (  , w_10439 );
and ( w_10438 , w_10439 , \3324_b0 );
or ( \3326_b1 , \3244_b1 , w_10441 );
not ( w_10441 , w_10442 );
and ( \3326_b0 , \3244_b0 , w_10443 );
and ( w_10442 ,  , w_10443 );
buf ( w_10441 , \3325_b1 );
not ( w_10441 , w_10444 );
not (  , w_10445 );
and ( w_10444 , w_10445 , \3325_b0 );
buf ( \3327_b1 , \a[6]_b1 );
not ( \3327_b1 , w_10446 );
not ( \3327_b0 , w_10447 );
and ( w_10446 , w_10447 , \a[6]_b0 );
buf ( \3328_b1 , \3196_b1 );
not ( \3328_b1 , w_10448 );
not ( \3328_b0 , w_10449 );
and ( w_10448 , w_10449 , \3196_b0 );
or ( \3329_b1 , \3327_b1 , w_10450 );
or ( \3329_b0 , \3327_b0 , \3328_b0 );
not ( \3328_b0 , w_10451 );
and ( w_10451 , w_10450 , \3328_b1 );
buf ( \3330_b1 , \d[6]_b1 );
not ( \3330_b1 , w_10452 );
not ( \3330_b0 , w_10453 );
and ( w_10452 , w_10453 , \d[6]_b0 );
buf ( \3331_b1 , \649_b1 );
not ( \3331_b1 , w_10454 );
not ( \3331_b0 , w_10455 );
and ( w_10454 , w_10455 , \649_b0 );
or ( \3332_b1 , \3330_b1 , w_10456 );
or ( \3332_b0 , \3330_b0 , \3331_b0 );
not ( \3331_b0 , w_10457 );
and ( w_10457 , w_10456 , \3331_b1 );
or ( \3333_b1 , \667_b1 , w_10459 );
not ( w_10459 , w_10460 );
and ( \3333_b0 , \667_b0 , w_10461 );
and ( w_10460 ,  , w_10461 );
buf ( w_10459 , \b[6]_b1 );
not ( w_10459 , w_10462 );
not (  , w_10463 );
and ( w_10462 , w_10463 , \b[6]_b0 );
or ( \3334_b1 , \3332_b1 , w_10465 );
not ( w_10465 , w_10466 );
and ( \3334_b0 , \3332_b0 , w_10467 );
and ( w_10466 ,  , w_10467 );
buf ( w_10465 , \3333_b1 );
not ( w_10465 , w_10468 );
not (  , w_10469 );
and ( w_10468 , w_10469 , \3333_b0 );
or ( \3335_b1 , \b[6]_b1 , \c[6]_b1 );
not ( \c[6]_b1 , w_10470 );
and ( \3335_b0 , \b[6]_b0 , w_10471 );
and ( w_10470 , w_10471 , \c[6]_b0 );
buf ( \3336_b1 , \3335_b1 );
not ( \3336_b1 , w_10472 );
not ( \3336_b0 , w_10473 );
and ( w_10472 , w_10473 , \3335_b0 );
buf ( \3337_b1 , \922_b1 );
not ( \3337_b1 , w_10474 );
not ( \3337_b0 , w_10475 );
and ( w_10474 , w_10475 , \922_b0 );
or ( \3338_b1 , \3336_b1 , w_10476 );
or ( \3338_b0 , \3336_b0 , \3337_b0 );
not ( \3337_b0 , w_10477 );
and ( w_10477 , w_10476 , \3337_b1 );
or ( \3339_b1 , \c[6]_b1 , \d[6]_b1 );
xor ( \3339_b0 , \c[6]_b0 , w_10478 );
not ( w_10478 , w_10479 );
and ( w_10479 , \d[6]_b1 , \d[6]_b0 );
or ( \3340_b1 , \903_b1 , \3339_b1 );
not ( \3339_b1 , w_10480 );
and ( \3340_b0 , \903_b0 , w_10481 );
and ( w_10480 , w_10481 , \3339_b0 );
or ( \3341_b1 , \2178_b1 , \2180_b1 );
xor ( \3341_b0 , \2178_b0 , w_10482 );
not ( w_10482 , w_10483 );
and ( w_10483 , \2180_b1 , \2180_b0 );
or ( \3342_b1 , \3341_b1 , \2261_b1 );
xor ( \3342_b0 , \3341_b0 , w_10484 );
not ( w_10484 , w_10485 );
and ( w_10485 , \2261_b1 , \2261_b0 );
buf ( \3343_b1 , \3342_b1 );
not ( \3343_b1 , w_10486 );
not ( \3343_b0 , w_10487 );
and ( w_10486 , w_10487 , \3342_b0 );
buf ( \3344_b1 , \2413_b1 );
not ( \3344_b1 , w_10488 );
not ( \3344_b0 , w_10489 );
and ( w_10488 , w_10489 , \2413_b0 );
or ( \3345_b1 , \3343_b1 , w_10490 );
or ( \3345_b0 , \3343_b0 , \3344_b0 );
not ( \3344_b0 , w_10491 );
and ( w_10491 , w_10490 , \3344_b1 );
or ( \3346_b1 , \1440_b1 , \1442_b1 );
xor ( \3346_b0 , \1440_b0 , w_10492 );
not ( w_10492 , w_10493 );
and ( w_10493 , \1442_b1 , \1442_b0 );
or ( \3347_b1 , \3346_b1 , \1520_b1 );
xor ( \3347_b0 , \3346_b0 , w_10494 );
not ( w_10494 , w_10495 );
and ( w_10495 , \1520_b1 , \1520_b0 );
or ( \3348_b1 , \2908_b1 , \3347_b1 );
not ( \3347_b1 , w_10496 );
and ( \3348_b0 , \2908_b0 , w_10497 );
and ( w_10496 , w_10497 , \3347_b0 );
buf ( \3349_b1 , \728_b1 );
not ( \3349_b1 , w_10498 );
not ( \3349_b0 , w_10499 );
and ( w_10498 , w_10499 , \728_b0 );
or ( \3350_b1 , \3349_b1 , w_10501 );
not ( w_10501 , w_10502 );
and ( \3350_b0 , \3349_b0 , w_10503 );
and ( w_10502 ,  , w_10503 );
buf ( w_10501 , \741_b1 );
not ( w_10501 , w_10504 );
not (  , w_10505 );
and ( w_10504 , w_10505 , \741_b0 );
buf ( \3351_b1 , \3350_b1 );
not ( \3351_b1 , w_10506 );
not ( \3351_b0 , w_10507 );
and ( w_10506 , w_10507 , \3350_b0 );
buf ( \3352_b1 , \727_b1 );
not ( \3352_b1 , w_10508 );
not ( \3352_b0 , w_10509 );
and ( w_10508 , w_10509 , \727_b0 );
or ( \3353_b1 , \3276_b1 , w_10510 );
or ( \3353_b0 , \3276_b0 , \3352_b0 );
not ( \3352_b0 , w_10511 );
and ( w_10511 , w_10510 , \3352_b1 );
or ( \3354_b1 , \3353_b1 , w_10513 );
not ( w_10513 , w_10514 );
and ( \3354_b0 , \3353_b0 , w_10515 );
and ( w_10514 ,  , w_10515 );
buf ( w_10513 , \3280_b1 );
not ( w_10513 , w_10516 );
not (  , w_10517 );
and ( w_10516 , w_10517 , \3280_b0 );
buf ( \3355_b1 , \3354_b1 );
not ( \3355_b1 , w_10518 );
not ( \3355_b0 , w_10519 );
and ( w_10518 , w_10519 , \3354_b0 );
or ( \3356_b1 , \3351_b1 , w_10520 );
or ( \3356_b0 , \3351_b0 , \3355_b0 );
not ( \3355_b0 , w_10521 );
and ( w_10521 , w_10520 , \3355_b1 );
or ( \3357_b1 , \3354_b1 , w_10522 );
or ( \3357_b0 , \3354_b0 , \3350_b0 );
not ( \3350_b0 , w_10523 );
and ( w_10523 , w_10522 , \3350_b1 );
or ( \3358_b1 , \3356_b1 , w_10525 );
not ( w_10525 , w_10526 );
and ( \3358_b0 , \3356_b0 , w_10527 );
and ( w_10526 ,  , w_10527 );
buf ( w_10525 , \3357_b1 );
not ( w_10525 , w_10528 );
not (  , w_10529 );
and ( w_10528 , w_10529 , \3357_b0 );
buf ( \3359_b1 , \3358_b1 );
not ( \3359_b1 , w_10530 );
not ( \3359_b0 , w_10531 );
and ( w_10530 , w_10531 , \3358_b0 );
buf ( \3360_b1 , \707_b1 );
not ( \3360_b1 , w_10532 );
not ( \3360_b0 , w_10533 );
and ( w_10532 , w_10533 , \707_b0 );
or ( \3361_b1 , \3359_b1 , w_10534 );
or ( \3361_b0 , \3359_b0 , \3360_b0 );
not ( \3360_b0 , w_10535 );
and ( w_10535 , w_10534 , \3360_b1 );
buf ( \3362_b1 , \813_b1 );
not ( \3362_b1 , w_10536 );
not ( \3362_b0 , w_10537 );
and ( w_10536 , w_10537 , \813_b0 );
or ( \3363_b1 , \3362_b1 , w_10539 );
not ( w_10539 , w_10540 );
and ( \3363_b0 , \3362_b0 , w_10541 );
and ( w_10540 ,  , w_10541 );
buf ( w_10539 , \826_b1 );
not ( w_10539 , w_10542 );
not (  , w_10543 );
and ( w_10542 , w_10543 , \826_b0 );
buf ( \3364_b1 , \3363_b1 );
not ( \3364_b1 , w_10544 );
not ( \3364_b0 , w_10545 );
and ( w_10544 , w_10545 , \3363_b0 );
buf ( \3365_b1 , \812_b1 );
not ( \3365_b1 , w_10546 );
not ( \3365_b0 , w_10547 );
and ( w_10546 , w_10547 , \812_b0 );
or ( \3366_b1 , \3297_b1 , w_10548 );
or ( \3366_b0 , \3297_b0 , \3365_b0 );
not ( \3365_b0 , w_10549 );
and ( w_10549 , w_10548 , \3365_b1 );
or ( \3367_b1 , \3366_b1 , w_10551 );
not ( w_10551 , w_10552 );
and ( \3367_b0 , \3366_b0 , w_10553 );
and ( w_10552 ,  , w_10553 );
buf ( w_10551 , \3301_b1 );
not ( w_10551 , w_10554 );
not (  , w_10555 );
and ( w_10554 , w_10555 , \3301_b0 );
buf ( \3368_b1 , \3367_b1 );
not ( \3368_b1 , w_10556 );
not ( \3368_b0 , w_10557 );
and ( w_10556 , w_10557 , \3367_b0 );
or ( \3369_b1 , \3364_b1 , w_10558 );
or ( \3369_b0 , \3364_b0 , \3368_b0 );
not ( \3368_b0 , w_10559 );
and ( w_10559 , w_10558 , \3368_b1 );
or ( \3370_b1 , \3367_b1 , w_10560 );
or ( \3370_b0 , \3367_b0 , \3363_b0 );
not ( \3363_b0 , w_10561 );
and ( w_10561 , w_10560 , \3363_b1 );
or ( \3371_b1 , \3369_b1 , w_10563 );
not ( w_10563 , w_10564 );
and ( \3371_b0 , \3369_b0 , w_10565 );
and ( w_10564 ,  , w_10565 );
buf ( w_10563 , \3370_b1 );
not ( w_10563 , w_10566 );
not (  , w_10567 );
and ( w_10566 , w_10567 , \3370_b0 );
or ( \3372_b1 , \880_b1 , \3371_b1 );
not ( \3371_b1 , w_10568 );
and ( \3372_b0 , \880_b0 , w_10569 );
and ( w_10568 , w_10569 , \3371_b0 );
buf ( \3373_b1 , \d[6]_b1 );
not ( \3373_b1 , w_10570 );
not ( \3373_b0 , w_10571 );
and ( w_10570 , w_10571 , \d[6]_b0 );
buf ( \3374_b1 , \894_b1 );
not ( \3374_b1 , w_10572 );
not ( \3374_b0 , w_10573 );
and ( w_10572 , w_10573 , \894_b0 );
or ( \3375_b1 , \3373_b1 , w_10574 );
or ( \3375_b0 , \3373_b0 , \3374_b0 );
not ( \3374_b0 , w_10575 );
and ( w_10575 , w_10574 , \3374_b1 );
or ( \3376_b1 , \885_b1 , \b[6]_b1 );
not ( \b[6]_b1 , w_10576 );
and ( \3376_b0 , \885_b0 , w_10577 );
and ( w_10576 , w_10577 , \b[6]_b0 );
or ( \3377_b1 , \909_b1 , \c[6]_b1 );
not ( \c[6]_b1 , w_10578 );
and ( \3377_b0 , \909_b0 , w_10579 );
and ( w_10578 , w_10579 , \c[6]_b0 );
or ( \3378_b1 , \3376_b1 , w_10581 );
not ( w_10581 , w_10582 );
and ( \3378_b0 , \3376_b0 , w_10583 );
and ( w_10582 ,  , w_10583 );
buf ( w_10581 , \3377_b1 );
not ( w_10581 , w_10584 );
not (  , w_10585 );
and ( w_10584 , w_10585 , \3377_b0 );
or ( \3379_b1 , \3375_b1 , w_10587 );
not ( w_10587 , w_10588 );
and ( \3379_b0 , \3375_b0 , w_10589 );
and ( w_10588 ,  , w_10589 );
buf ( w_10587 , \3378_b1 );
not ( w_10587 , w_10590 );
not (  , w_10591 );
and ( w_10590 , w_10591 , \3378_b0 );
or ( \3380_b1 , \3372_b1 , w_10593 );
not ( w_10593 , w_10594 );
and ( \3380_b0 , \3372_b0 , w_10595 );
and ( w_10594 ,  , w_10595 );
buf ( w_10593 , \3379_b1 );
not ( w_10593 , w_10596 );
not (  , w_10597 );
and ( w_10596 , w_10597 , \3379_b0 );
or ( \3381_b1 , \3361_b1 , w_10599 );
not ( w_10599 , w_10600 );
and ( \3381_b0 , \3361_b0 , w_10601 );
and ( w_10600 ,  , w_10601 );
buf ( w_10599 , \3380_b1 );
not ( w_10599 , w_10602 );
not (  , w_10603 );
and ( w_10602 , w_10603 , \3380_b0 );
or ( \3382_b1 , \3348_b1 , w_10605 );
not ( w_10605 , w_10606 );
and ( \3382_b0 , \3348_b0 , w_10607 );
and ( w_10606 ,  , w_10607 );
buf ( w_10605 , \3381_b1 );
not ( w_10605 , w_10608 );
not (  , w_10609 );
and ( w_10608 , w_10609 , \3381_b0 );
or ( \3383_b1 , \3345_b1 , w_10611 );
not ( w_10611 , w_10612 );
and ( \3383_b0 , \3345_b0 , w_10613 );
and ( w_10612 ,  , w_10613 );
buf ( w_10611 , \3382_b1 );
not ( w_10611 , w_10614 );
not (  , w_10615 );
and ( w_10614 , w_10615 , \3382_b0 );
or ( \3384_b1 , \3340_b1 , w_10617 );
not ( w_10617 , w_10618 );
and ( \3384_b0 , \3340_b0 , w_10619 );
and ( w_10618 ,  , w_10619 );
buf ( w_10617 , \3383_b1 );
not ( w_10617 , w_10620 );
not (  , w_10621 );
and ( w_10620 , w_10621 , \3383_b0 );
or ( \3385_b1 , \3338_b1 , w_10623 );
not ( w_10623 , w_10624 );
and ( \3385_b0 , \3338_b0 , w_10625 );
and ( w_10624 ,  , w_10625 );
buf ( w_10623 , \3384_b1 );
not ( w_10623 , w_10626 );
not (  , w_10627 );
and ( w_10626 , w_10627 , \3384_b0 );
or ( \3386_b1 , \3334_b1 , w_10629 );
not ( w_10629 , w_10630 );
and ( \3386_b0 , \3334_b0 , w_10631 );
and ( w_10630 ,  , w_10631 );
buf ( w_10629 , \3385_b1 );
not ( w_10629 , w_10632 );
not (  , w_10633 );
and ( w_10632 , w_10633 , \3385_b0 );
or ( \3387_b1 , \3329_b1 , w_10635 );
not ( w_10635 , w_10636 );
and ( \3387_b0 , \3329_b0 , w_10637 );
and ( w_10636 ,  , w_10637 );
buf ( w_10635 , \3386_b1 );
not ( w_10635 , w_10638 );
not (  , w_10639 );
and ( w_10638 , w_10639 , \3386_b0 );
buf ( \3388_b1 , \a[5]_b1 );
not ( \3388_b1 , w_10640 );
not ( \3388_b0 , w_10641 );
and ( w_10640 , w_10641 , \a[5]_b0 );
buf ( \3389_b1 , \3075_b1 );
not ( \3389_b1 , w_10642 );
not ( \3389_b0 , w_10643 );
and ( w_10642 , w_10643 , \3075_b0 );
or ( \3390_b1 , \3388_b1 , w_10644 );
or ( \3390_b0 , \3388_b0 , \3389_b0 );
not ( \3389_b0 , w_10645 );
and ( w_10645 , w_10644 , \3389_b1 );
buf ( \3391_b1 , \d[5]_b1 );
not ( \3391_b1 , w_10646 );
not ( \3391_b0 , w_10647 );
and ( w_10646 , w_10647 , \d[5]_b0 );
buf ( \3392_b1 , \649_b1 );
not ( \3392_b1 , w_10648 );
not ( \3392_b0 , w_10649 );
and ( w_10648 , w_10649 , \649_b0 );
or ( \3393_b1 , \3391_b1 , w_10650 );
or ( \3393_b0 , \3391_b0 , \3392_b0 );
not ( \3392_b0 , w_10651 );
and ( w_10651 , w_10650 , \3392_b1 );
or ( \3394_b1 , \667_b1 , w_10653 );
not ( w_10653 , w_10654 );
and ( \3394_b0 , \667_b0 , w_10655 );
and ( w_10654 ,  , w_10655 );
buf ( w_10653 , \b[5]_b1 );
not ( w_10653 , w_10656 );
not (  , w_10657 );
and ( w_10656 , w_10657 , \b[5]_b0 );
or ( \3395_b1 , \3393_b1 , w_10659 );
not ( w_10659 , w_10660 );
and ( \3395_b0 , \3393_b0 , w_10661 );
and ( w_10660 ,  , w_10661 );
buf ( w_10659 , \3394_b1 );
not ( w_10659 , w_10662 );
not (  , w_10663 );
and ( w_10662 , w_10663 , \3394_b0 );
or ( \3396_b1 , \b[5]_b1 , \c[5]_b1 );
not ( \c[5]_b1 , w_10664 );
and ( \3396_b0 , \b[5]_b0 , w_10665 );
and ( w_10664 , w_10665 , \c[5]_b0 );
buf ( \3397_b1 , \3396_b1 );
not ( \3397_b1 , w_10666 );
not ( \3397_b0 , w_10667 );
and ( w_10666 , w_10667 , \3396_b0 );
buf ( \3398_b1 , \922_b1 );
not ( \3398_b1 , w_10668 );
not ( \3398_b0 , w_10669 );
and ( w_10668 , w_10669 , \922_b0 );
or ( \3399_b1 , \3397_b1 , w_10670 );
or ( \3399_b0 , \3397_b0 , \3398_b0 );
not ( \3398_b0 , w_10671 );
and ( w_10671 , w_10670 , \3398_b1 );
or ( \3400_b1 , \c[5]_b1 , \d[5]_b1 );
xor ( \3400_b0 , \c[5]_b0 , w_10672 );
not ( w_10672 , w_10673 );
and ( w_10673 , \d[5]_b1 , \d[5]_b0 );
or ( \3401_b1 , \3400_b1 , \903_b1 );
not ( \903_b1 , w_10674 );
and ( \3401_b0 , \3400_b0 , w_10675 );
and ( w_10674 , w_10675 , \903_b0 );
buf ( \3402_b1 , \2258_b1 );
not ( \3402_b1 , w_10676 );
not ( \3402_b0 , w_10677 );
and ( w_10676 , w_10677 , \2258_b0 );
or ( \3403_b1 , \3402_b1 , w_10679 );
not ( w_10679 , w_10680 );
and ( \3403_b0 , \3402_b0 , w_10681 );
and ( w_10680 ,  , w_10681 );
buf ( w_10679 , \2260_b1 );
not ( w_10679 , w_10682 );
not (  , w_10683 );
and ( w_10682 , w_10683 , \2260_b0 );
or ( \3404_b1 , \3403_b1 , \2248_b1 );
xor ( \3404_b0 , \3403_b0 , w_10684 );
not ( w_10684 , w_10685 );
and ( w_10685 , \2248_b1 , \2248_b0 );
buf ( \3405_b1 , \3404_b1 );
not ( \3405_b1 , w_10686 );
not ( \3405_b0 , w_10687 );
and ( w_10686 , w_10687 , \3404_b0 );
buf ( \3406_b1 , \2413_b1 );
not ( \3406_b1 , w_10688 );
not ( \3406_b0 , w_10689 );
and ( w_10688 , w_10689 , \2413_b0 );
or ( \3407_b1 , \3405_b1 , w_10690 );
or ( \3407_b0 , \3405_b0 , \3406_b0 );
not ( \3406_b0 , w_10691 );
and ( w_10691 , w_10690 , \3406_b1 );
buf ( \3408_b1 , \1466_b1 );
not ( \3408_b1 , w_10692 );
not ( \3408_b0 , w_10693 );
and ( w_10692 , w_10693 , \1466_b0 );
or ( \3409_b1 , \3408_b1 , w_10695 );
not ( w_10695 , w_10696 );
and ( \3409_b0 , \3408_b0 , w_10697 );
and ( w_10696 ,  , w_10697 );
buf ( w_10695 , \1519_b1 );
not ( w_10695 , w_10698 );
not (  , w_10699 );
and ( w_10698 , w_10699 , \1519_b0 );
or ( \3410_b1 , \1517_b1 , \3409_b1 );
xor ( \3410_b0 , \1517_b0 , w_10700 );
not ( w_10700 , w_10701 );
and ( w_10701 , \3409_b1 , \3409_b0 );
or ( \3411_b1 , \2908_b1 , \3410_b1 );
not ( \3410_b1 , w_10702 );
and ( \3411_b0 , \2908_b0 , w_10703 );
and ( w_10702 , w_10703 , \3410_b0 );
buf ( \3412_b1 , \725_b1 );
not ( \3412_b1 , w_10704 );
not ( \3412_b0 , w_10705 );
and ( w_10704 , w_10705 , \725_b0 );
or ( \3413_b1 , \3412_b1 , w_10707 );
not ( w_10707 , w_10708 );
and ( \3413_b0 , \3412_b0 , w_10709 );
and ( w_10708 ,  , w_10709 );
buf ( w_10707 , \742_b1 );
not ( w_10707 , w_10710 );
not (  , w_10711 );
and ( w_10710 , w_10711 , \742_b0 );
buf ( \3414_b1 , \3413_b1 );
not ( \3414_b1 , w_10712 );
not ( \3414_b0 , w_10713 );
and ( w_10712 , w_10713 , \3413_b0 );
or ( \3415_b1 , \3276_b1 , w_10714 );
or ( \3415_b0 , \3276_b0 , \726_b0 );
not ( \726_b0 , w_10715 );
and ( w_10715 , w_10714 , \726_b1 );
or ( \3416_b1 , \3415_b1 , w_10717 );
not ( w_10717 , w_10718 );
and ( \3416_b0 , \3415_b0 , w_10719 );
and ( w_10718 ,  , w_10719 );
buf ( w_10717 , \743_b1 );
not ( w_10717 , w_10720 );
not (  , w_10721 );
and ( w_10720 , w_10721 , \743_b0 );
buf ( \3417_b1 , \3416_b1 );
not ( \3417_b1 , w_10722 );
not ( \3417_b0 , w_10723 );
and ( w_10722 , w_10723 , \3416_b0 );
or ( \3418_b1 , \3414_b1 , w_10724 );
or ( \3418_b0 , \3414_b0 , \3417_b0 );
not ( \3417_b0 , w_10725 );
and ( w_10725 , w_10724 , \3417_b1 );
or ( \3419_b1 , \3416_b1 , w_10726 );
or ( \3419_b0 , \3416_b0 , \3413_b0 );
not ( \3413_b0 , w_10727 );
and ( w_10727 , w_10726 , \3413_b1 );
or ( \3420_b1 , \3418_b1 , w_10729 );
not ( w_10729 , w_10730 );
and ( \3420_b0 , \3418_b0 , w_10731 );
and ( w_10730 ,  , w_10731 );
buf ( w_10729 , \3419_b1 );
not ( w_10729 , w_10732 );
not (  , w_10733 );
and ( w_10732 , w_10733 , \3419_b0 );
buf ( \3421_b1 , \3420_b1 );
not ( \3421_b1 , w_10734 );
not ( \3421_b0 , w_10735 );
and ( w_10734 , w_10735 , \3420_b0 );
buf ( \3422_b1 , \707_b1 );
not ( \3422_b1 , w_10736 );
not ( \3422_b0 , w_10737 );
and ( w_10736 , w_10737 , \707_b0 );
or ( \3423_b1 , \3421_b1 , w_10738 );
or ( \3423_b0 , \3421_b0 , \3422_b0 );
not ( \3422_b0 , w_10739 );
and ( w_10739 , w_10738 , \3422_b1 );
buf ( \3424_b1 , \810_b1 );
not ( \3424_b1 , w_10740 );
not ( \3424_b0 , w_10741 );
and ( w_10740 , w_10741 , \810_b0 );
or ( \3425_b1 , \3424_b1 , w_10743 );
not ( w_10743 , w_10744 );
and ( \3425_b0 , \3424_b0 , w_10745 );
and ( w_10744 ,  , w_10745 );
buf ( w_10743 , \827_b1 );
not ( w_10743 , w_10746 );
not (  , w_10747 );
and ( w_10746 , w_10747 , \827_b0 );
buf ( \3426_b1 , \3425_b1 );
not ( \3426_b1 , w_10748 );
not ( \3426_b0 , w_10749 );
and ( w_10748 , w_10749 , \3425_b0 );
or ( \3427_b1 , \811_b1 , w_10750 );
or ( \3427_b0 , \811_b0 , \3297_b0 );
not ( \3297_b0 , w_10751 );
and ( w_10751 , w_10750 , \3297_b1 );
or ( \3428_b1 , \3427_b1 , w_10753 );
not ( w_10753 , w_10754 );
and ( \3428_b0 , \3427_b0 , w_10755 );
and ( w_10754 ,  , w_10755 );
buf ( w_10753 , \828_b1 );
not ( w_10753 , w_10756 );
not (  , w_10757 );
and ( w_10756 , w_10757 , \828_b0 );
buf ( \3429_b1 , \3428_b1 );
not ( \3429_b1 , w_10758 );
not ( \3429_b0 , w_10759 );
and ( w_10758 , w_10759 , \3428_b0 );
or ( \3430_b1 , \3426_b1 , w_10760 );
or ( \3430_b0 , \3426_b0 , \3429_b0 );
not ( \3429_b0 , w_10761 );
and ( w_10761 , w_10760 , \3429_b1 );
or ( \3431_b1 , \3428_b1 , w_10762 );
or ( \3431_b0 , \3428_b0 , \3425_b0 );
not ( \3425_b0 , w_10763 );
and ( w_10763 , w_10762 , \3425_b1 );
or ( \3432_b1 , \3430_b1 , w_10765 );
not ( w_10765 , w_10766 );
and ( \3432_b0 , \3430_b0 , w_10767 );
and ( w_10766 ,  , w_10767 );
buf ( w_10765 , \3431_b1 );
not ( w_10765 , w_10768 );
not (  , w_10769 );
and ( w_10768 , w_10769 , \3431_b0 );
or ( \3433_b1 , \880_b1 , \3432_b1 );
not ( \3432_b1 , w_10770 );
and ( \3433_b0 , \880_b0 , w_10771 );
and ( w_10770 , w_10771 , \3432_b0 );
buf ( \3434_b1 , \d[5]_b1 );
not ( \3434_b1 , w_10772 );
not ( \3434_b0 , w_10773 );
and ( w_10772 , w_10773 , \d[5]_b0 );
buf ( \3435_b1 , \894_b1 );
not ( \3435_b1 , w_10774 );
not ( \3435_b0 , w_10775 );
and ( w_10774 , w_10775 , \894_b0 );
or ( \3436_b1 , \3434_b1 , w_10776 );
or ( \3436_b0 , \3434_b0 , \3435_b0 );
not ( \3435_b0 , w_10777 );
and ( w_10777 , w_10776 , \3435_b1 );
or ( \3437_b1 , \885_b1 , \b[5]_b1 );
not ( \b[5]_b1 , w_10778 );
and ( \3437_b0 , \885_b0 , w_10779 );
and ( w_10778 , w_10779 , \b[5]_b0 );
or ( \3438_b1 , \909_b1 , \c[5]_b1 );
not ( \c[5]_b1 , w_10780 );
and ( \3438_b0 , \909_b0 , w_10781 );
and ( w_10780 , w_10781 , \c[5]_b0 );
or ( \3439_b1 , \3437_b1 , w_10783 );
not ( w_10783 , w_10784 );
and ( \3439_b0 , \3437_b0 , w_10785 );
and ( w_10784 ,  , w_10785 );
buf ( w_10783 , \3438_b1 );
not ( w_10783 , w_10786 );
not (  , w_10787 );
and ( w_10786 , w_10787 , \3438_b0 );
or ( \3440_b1 , \3436_b1 , w_10789 );
not ( w_10789 , w_10790 );
and ( \3440_b0 , \3436_b0 , w_10791 );
and ( w_10790 ,  , w_10791 );
buf ( w_10789 , \3439_b1 );
not ( w_10789 , w_10792 );
not (  , w_10793 );
and ( w_10792 , w_10793 , \3439_b0 );
or ( \3441_b1 , \3433_b1 , w_10795 );
not ( w_10795 , w_10796 );
and ( \3441_b0 , \3433_b0 , w_10797 );
and ( w_10796 ,  , w_10797 );
buf ( w_10795 , \3440_b1 );
not ( w_10795 , w_10798 );
not (  , w_10799 );
and ( w_10798 , w_10799 , \3440_b0 );
or ( \3442_b1 , \3423_b1 , w_10801 );
not ( w_10801 , w_10802 );
and ( \3442_b0 , \3423_b0 , w_10803 );
and ( w_10802 ,  , w_10803 );
buf ( w_10801 , \3441_b1 );
not ( w_10801 , w_10804 );
not (  , w_10805 );
and ( w_10804 , w_10805 , \3441_b0 );
or ( \3443_b1 , \3411_b1 , w_10807 );
not ( w_10807 , w_10808 );
and ( \3443_b0 , \3411_b0 , w_10809 );
and ( w_10808 ,  , w_10809 );
buf ( w_10807 , \3442_b1 );
not ( w_10807 , w_10810 );
not (  , w_10811 );
and ( w_10810 , w_10811 , \3442_b0 );
or ( \3444_b1 , \3407_b1 , w_10813 );
not ( w_10813 , w_10814 );
and ( \3444_b0 , \3407_b0 , w_10815 );
and ( w_10814 ,  , w_10815 );
buf ( w_10813 , \3443_b1 );
not ( w_10813 , w_10816 );
not (  , w_10817 );
and ( w_10816 , w_10817 , \3443_b0 );
or ( \3445_b1 , \3401_b1 , w_10819 );
not ( w_10819 , w_10820 );
and ( \3445_b0 , \3401_b0 , w_10821 );
and ( w_10820 ,  , w_10821 );
buf ( w_10819 , \3444_b1 );
not ( w_10819 , w_10822 );
not (  , w_10823 );
and ( w_10822 , w_10823 , \3444_b0 );
or ( \3446_b1 , \3399_b1 , w_10825 );
not ( w_10825 , w_10826 );
and ( \3446_b0 , \3399_b0 , w_10827 );
and ( w_10826 ,  , w_10827 );
buf ( w_10825 , \3445_b1 );
not ( w_10825 , w_10828 );
not (  , w_10829 );
and ( w_10828 , w_10829 , \3445_b0 );
or ( \3447_b1 , \3395_b1 , w_10831 );
not ( w_10831 , w_10832 );
and ( \3447_b0 , \3395_b0 , w_10833 );
and ( w_10832 ,  , w_10833 );
buf ( w_10831 , \3446_b1 );
not ( w_10831 , w_10834 );
not (  , w_10835 );
and ( w_10834 , w_10835 , \3446_b0 );
or ( \3448_b1 , \3390_b1 , w_10837 );
not ( w_10837 , w_10838 );
and ( \3448_b0 , \3390_b0 , w_10839 );
and ( w_10838 ,  , w_10839 );
buf ( w_10837 , \3447_b1 );
not ( w_10837 , w_10840 );
not (  , w_10841 );
and ( w_10840 , w_10841 , \3447_b0 );
buf ( \3449_b1 , \a[4]_b1 );
not ( \3449_b1 , w_10842 );
not ( \3449_b0 , w_10843 );
and ( w_10842 , w_10843 , \a[4]_b0 );
buf ( \3450_b1 , \3075_b1 );
not ( \3450_b1 , w_10844 );
not ( \3450_b0 , w_10845 );
and ( w_10844 , w_10845 , \3075_b0 );
or ( \3451_b1 , \3449_b1 , w_10846 );
or ( \3451_b0 , \3449_b0 , \3450_b0 );
not ( \3450_b0 , w_10847 );
and ( w_10847 , w_10846 , \3450_b1 );
buf ( \3452_b1 , \d[4]_b1 );
not ( \3452_b1 , w_10848 );
not ( \3452_b0 , w_10849 );
and ( w_10848 , w_10849 , \d[4]_b0 );
buf ( \3453_b1 , \648_b1 );
not ( \3453_b1 , w_10850 );
not ( \3453_b0 , w_10851 );
and ( w_10850 , w_10851 , \648_b0 );
or ( \3454_b1 , \3452_b1 , w_10852 );
or ( \3454_b0 , \3452_b0 , \3453_b0 );
not ( \3453_b0 , w_10853 );
and ( w_10853 , w_10852 , \3453_b1 );
or ( \3455_b1 , \667_b1 , w_10855 );
not ( w_10855 , w_10856 );
and ( \3455_b0 , \667_b0 , w_10857 );
and ( w_10856 ,  , w_10857 );
buf ( w_10855 , \b[4]_b1 );
not ( w_10855 , w_10858 );
not (  , w_10859 );
and ( w_10858 , w_10859 , \b[4]_b0 );
or ( \3456_b1 , \3454_b1 , w_10861 );
not ( w_10861 , w_10862 );
and ( \3456_b0 , \3454_b0 , w_10863 );
and ( w_10862 ,  , w_10863 );
buf ( w_10861 , \3455_b1 );
not ( w_10861 , w_10864 );
not (  , w_10865 );
and ( w_10864 , w_10865 , \3455_b0 );
or ( \3457_b1 , \b[4]_b1 , \c[4]_b1 );
not ( \c[4]_b1 , w_10866 );
and ( \3457_b0 , \b[4]_b0 , w_10867 );
and ( w_10866 , w_10867 , \c[4]_b0 );
buf ( \3458_b1 , \3457_b1 );
not ( \3458_b1 , w_10868 );
not ( \3458_b0 , w_10869 );
and ( w_10868 , w_10869 , \3457_b0 );
buf ( \3459_b1 , \2887_b1 );
not ( \3459_b1 , w_10870 );
not ( \3459_b0 , w_10871 );
and ( w_10870 , w_10871 , \2887_b0 );
or ( \3460_b1 , \3458_b1 , w_10872 );
or ( \3460_b0 , \3458_b0 , \3459_b0 );
not ( \3459_b0 , w_10873 );
and ( w_10873 , w_10872 , \3459_b1 );
or ( \3461_b1 , \c[4]_b1 , \d[4]_b1 );
xor ( \3461_b0 , \c[4]_b0 , w_10874 );
not ( w_10874 , w_10875 );
and ( w_10875 , \d[4]_b1 , \d[4]_b0 );
or ( \3462_b1 , \903_b1 , \3461_b1 );
not ( \3461_b1 , w_10876 );
and ( \3462_b0 , \903_b0 , w_10877 );
and ( w_10876 , w_10877 , \3461_b0 );
buf ( \3463_b1 , \2229_b1 );
not ( \3463_b1 , w_10878 );
not ( \3463_b0 , w_10879 );
and ( w_10878 , w_10879 , \2229_b0 );
buf ( \3464_b1 , \2247_b1 );
not ( \3464_b1 , w_10880 );
not ( \3464_b0 , w_10881 );
and ( w_10880 , w_10881 , \2247_b0 );
or ( \3465_b1 , \3464_b1 , w_10883 );
not ( w_10883 , w_10884 );
and ( \3465_b0 , \3464_b0 , w_10885 );
and ( w_10884 ,  , w_10885 );
buf ( w_10883 , \2245_b1 );
not ( w_10883 , w_10886 );
not (  , w_10887 );
and ( w_10886 , w_10887 , \2245_b0 );
buf ( \3466_b1 , \3465_b1 );
not ( \3466_b1 , w_10888 );
not ( \3466_b0 , w_10889 );
and ( w_10888 , w_10889 , \3465_b0 );
or ( \3467_b1 , \3463_b1 , w_10890 );
or ( \3467_b0 , \3463_b0 , \3466_b0 );
not ( \3466_b0 , w_10891 );
and ( w_10891 , w_10890 , \3466_b1 );
or ( \3468_b1 , \3465_b1 , w_10892 );
or ( \3468_b0 , \3465_b0 , \2229_b0 );
not ( \2229_b0 , w_10893 );
and ( w_10893 , w_10892 , \2229_b1 );
or ( \3469_b1 , \3467_b1 , w_10895 );
not ( w_10895 , w_10896 );
and ( \3469_b0 , \3467_b0 , w_10897 );
and ( w_10896 ,  , w_10897 );
buf ( w_10895 , \3468_b1 );
not ( w_10895 , w_10898 );
not (  , w_10899 );
and ( w_10898 , w_10899 , \3468_b0 );
buf ( \3470_b1 , \3469_b1 );
not ( \3470_b1 , w_10900 );
not ( \3470_b0 , w_10901 );
and ( w_10900 , w_10901 , \3469_b0 );
buf ( \3471_b1 , \2413_b1 );
not ( \3471_b1 , w_10902 );
not ( \3471_b0 , w_10903 );
and ( w_10902 , w_10903 , \2413_b0 );
or ( \3472_b1 , \3470_b1 , w_10904 );
or ( \3472_b0 , \3470_b0 , \3471_b0 );
not ( \3471_b0 , w_10905 );
and ( w_10905 , w_10904 , \3471_b1 );
buf ( \3473_b1 , \1509_b1 );
not ( \3473_b1 , w_10906 );
not ( \3473_b0 , w_10907 );
and ( w_10906 , w_10907 , \1509_b0 );
buf ( \3474_b1 , \1516_b1 );
not ( \3474_b1 , w_10908 );
not ( \3474_b0 , w_10909 );
and ( w_10908 , w_10909 , \1516_b0 );
or ( \3475_b1 , \3474_b1 , w_10911 );
not ( w_10911 , w_10912 );
and ( \3475_b0 , \3474_b0 , w_10913 );
and ( w_10912 ,  , w_10913 );
buf ( w_10911 , \1514_b1 );
not ( w_10911 , w_10914 );
not (  , w_10915 );
and ( w_10914 , w_10915 , \1514_b0 );
buf ( \3476_b1 , \3475_b1 );
not ( \3476_b1 , w_10916 );
not ( \3476_b0 , w_10917 );
and ( w_10916 , w_10917 , \3475_b0 );
or ( \3477_b1 , \3473_b1 , w_10918 );
or ( \3477_b0 , \3473_b0 , \3476_b0 );
not ( \3476_b0 , w_10919 );
and ( w_10919 , w_10918 , \3476_b1 );
or ( \3478_b1 , \3475_b1 , w_10920 );
or ( \3478_b0 , \3475_b0 , \1509_b0 );
not ( \1509_b0 , w_10921 );
and ( w_10921 , w_10920 , \1509_b1 );
or ( \3479_b1 , \3477_b1 , w_10923 );
not ( w_10923 , w_10924 );
and ( \3479_b0 , \3477_b0 , w_10925 );
and ( w_10924 ,  , w_10925 );
buf ( w_10923 , \3478_b1 );
not ( w_10923 , w_10926 );
not (  , w_10927 );
and ( w_10926 , w_10927 , \3478_b0 );
or ( \3480_b1 , \2908_b1 , \3479_b1 );
not ( \3479_b1 , w_10928 );
and ( \3480_b0 , \2908_b0 , w_10929 );
and ( w_10928 , w_10929 , \3479_b0 );
buf ( \3481_b1 , \743_b1 );
not ( \3481_b1 , w_10930 );
not ( \3481_b0 , w_10931 );
and ( w_10930 , w_10931 , \743_b0 );
or ( \3482_b1 , \3481_b1 , w_10933 );
not ( w_10933 , w_10934 );
and ( \3482_b0 , \3481_b0 , w_10935 );
and ( w_10934 ,  , w_10935 );
buf ( w_10933 , \726_b1 );
not ( w_10933 , w_10936 );
not (  , w_10937 );
and ( w_10936 , w_10937 , \726_b0 );
buf ( \3483_b1 , \3482_b1 );
not ( \3483_b1 , w_10938 );
not ( \3483_b0 , w_10939 );
and ( w_10938 , w_10939 , \3482_b0 );
buf ( \3484_b1 , \3276_b1 );
not ( \3484_b1 , w_10940 );
not ( \3484_b0 , w_10941 );
and ( w_10940 , w_10941 , \3276_b0 );
or ( \3485_b1 , \3483_b1 , w_10942 );
or ( \3485_b0 , \3483_b0 , \3484_b0 );
not ( \3484_b0 , w_10943 );
and ( w_10943 , w_10942 , \3484_b1 );
or ( \3486_b1 , \3276_b1 , w_10944 );
or ( \3486_b0 , \3276_b0 , \3482_b0 );
not ( \3482_b0 , w_10945 );
and ( w_10945 , w_10944 , \3482_b1 );
or ( \3487_b1 , \3485_b1 , w_10947 );
not ( w_10947 , w_10948 );
and ( \3487_b0 , \3485_b0 , w_10949 );
and ( w_10948 ,  , w_10949 );
buf ( w_10947 , \3486_b1 );
not ( w_10947 , w_10950 );
not (  , w_10951 );
and ( w_10950 , w_10951 , \3486_b0 );
buf ( \3488_b1 , \3487_b1 );
not ( \3488_b1 , w_10952 );
not ( \3488_b0 , w_10953 );
and ( w_10952 , w_10953 , \3487_b0 );
buf ( \3489_b1 , \707_b1 );
not ( \3489_b1 , w_10954 );
not ( \3489_b0 , w_10955 );
and ( w_10954 , w_10955 , \707_b0 );
or ( \3490_b1 , \3488_b1 , w_10956 );
or ( \3490_b0 , \3488_b0 , \3489_b0 );
not ( \3489_b0 , w_10957 );
and ( w_10957 , w_10956 , \3489_b1 );
buf ( \3491_b1 , \828_b1 );
not ( \3491_b1 , w_10958 );
not ( \3491_b0 , w_10959 );
and ( w_10958 , w_10959 , \828_b0 );
or ( \3492_b1 , \3491_b1 , w_10961 );
not ( w_10961 , w_10962 );
and ( \3492_b0 , \3491_b0 , w_10963 );
and ( w_10962 ,  , w_10963 );
buf ( w_10961 , \811_b1 );
not ( w_10961 , w_10964 );
not (  , w_10965 );
and ( w_10964 , w_10965 , \811_b0 );
buf ( \3493_b1 , \3492_b1 );
not ( \3493_b1 , w_10966 );
not ( \3493_b0 , w_10967 );
and ( w_10966 , w_10967 , \3492_b0 );
buf ( \3494_b1 , \3297_b1 );
not ( \3494_b1 , w_10968 );
not ( \3494_b0 , w_10969 );
and ( w_10968 , w_10969 , \3297_b0 );
or ( \3495_b1 , \3493_b1 , w_10970 );
or ( \3495_b0 , \3493_b0 , \3494_b0 );
not ( \3494_b0 , w_10971 );
and ( w_10971 , w_10970 , \3494_b1 );
or ( \3496_b1 , \3297_b1 , w_10972 );
or ( \3496_b0 , \3297_b0 , \3492_b0 );
not ( \3492_b0 , w_10973 );
and ( w_10973 , w_10972 , \3492_b1 );
or ( \3497_b1 , \3495_b1 , w_10975 );
not ( w_10975 , w_10976 );
and ( \3497_b0 , \3495_b0 , w_10977 );
and ( w_10976 ,  , w_10977 );
buf ( w_10975 , \3496_b1 );
not ( w_10975 , w_10978 );
not (  , w_10979 );
and ( w_10978 , w_10979 , \3496_b0 );
or ( \3498_b1 , \880_b1 , \3497_b1 );
not ( \3497_b1 , w_10980 );
and ( \3498_b0 , \880_b0 , w_10981 );
and ( w_10980 , w_10981 , \3497_b0 );
buf ( \3499_b1 , \d[4]_b1 );
not ( \3499_b1 , w_10982 );
not ( \3499_b0 , w_10983 );
and ( w_10982 , w_10983 , \d[4]_b0 );
buf ( \3500_b1 , \894_b1 );
not ( \3500_b1 , w_10984 );
not ( \3500_b0 , w_10985 );
and ( w_10984 , w_10985 , \894_b0 );
or ( \3501_b1 , \3499_b1 , w_10986 );
or ( \3501_b0 , \3499_b0 , \3500_b0 );
not ( \3500_b0 , w_10987 );
and ( w_10987 , w_10986 , \3500_b1 );
buf ( \3502_b1 , \886_b1 );
not ( \3502_b1 , w_10988 );
not ( \3502_b0 , w_10989 );
and ( w_10988 , w_10989 , \886_b0 );
buf ( \3503_b1 , \b[4]_b1 );
not ( \3503_b1 , w_10990 );
not ( \3503_b0 , w_10991 );
and ( w_10990 , w_10991 , \b[4]_b0 );
buf ( \3504_b1 , \3503_b1 );
not ( \3504_b1 , w_10992 );
not ( \3504_b0 , w_10993 );
and ( w_10992 , w_10993 , \3503_b0 );
or ( \3505_b1 , \3502_b1 , \3504_b1 );
not ( \3504_b1 , w_10994 );
and ( \3505_b0 , \3502_b0 , w_10995 );
and ( w_10994 , w_10995 , \3504_b0 );
or ( \3506_b1 , \907_b1 , \c[4]_b1 );
not ( \c[4]_b1 , w_10996 );
and ( \3506_b0 , \907_b0 , w_10997 );
and ( w_10996 , w_10997 , \c[4]_b0 );
or ( \3507_b1 , \3505_b1 , w_10999 );
not ( w_10999 , w_11000 );
and ( \3507_b0 , \3505_b0 , w_11001 );
and ( w_11000 ,  , w_11001 );
buf ( w_10999 , \3506_b1 );
not ( w_10999 , w_11002 );
not (  , w_11003 );
and ( w_11002 , w_11003 , \3506_b0 );
or ( \3508_b1 , \3501_b1 , w_11005 );
not ( w_11005 , w_11006 );
and ( \3508_b0 , \3501_b0 , w_11007 );
and ( w_11006 ,  , w_11007 );
buf ( w_11005 , \3507_b1 );
not ( w_11005 , w_11008 );
not (  , w_11009 );
and ( w_11008 , w_11009 , \3507_b0 );
or ( \3509_b1 , \3498_b1 , w_11011 );
not ( w_11011 , w_11012 );
and ( \3509_b0 , \3498_b0 , w_11013 );
and ( w_11012 ,  , w_11013 );
buf ( w_11011 , \3508_b1 );
not ( w_11011 , w_11014 );
not (  , w_11015 );
and ( w_11014 , w_11015 , \3508_b0 );
or ( \3510_b1 , \3490_b1 , w_11017 );
not ( w_11017 , w_11018 );
and ( \3510_b0 , \3490_b0 , w_11019 );
and ( w_11018 ,  , w_11019 );
buf ( w_11017 , \3509_b1 );
not ( w_11017 , w_11020 );
not (  , w_11021 );
and ( w_11020 , w_11021 , \3509_b0 );
or ( \3511_b1 , \3480_b1 , w_11023 );
not ( w_11023 , w_11024 );
and ( \3511_b0 , \3480_b0 , w_11025 );
and ( w_11024 ,  , w_11025 );
buf ( w_11023 , \3510_b1 );
not ( w_11023 , w_11026 );
not (  , w_11027 );
and ( w_11026 , w_11027 , \3510_b0 );
or ( \3512_b1 , \3472_b1 , w_11029 );
not ( w_11029 , w_11030 );
and ( \3512_b0 , \3472_b0 , w_11031 );
and ( w_11030 ,  , w_11031 );
buf ( w_11029 , \3511_b1 );
not ( w_11029 , w_11032 );
not (  , w_11033 );
and ( w_11032 , w_11033 , \3511_b0 );
or ( \3513_b1 , \3462_b1 , w_11035 );
not ( w_11035 , w_11036 );
and ( \3513_b0 , \3462_b0 , w_11037 );
and ( w_11036 ,  , w_11037 );
buf ( w_11035 , \3512_b1 );
not ( w_11035 , w_11038 );
not (  , w_11039 );
and ( w_11038 , w_11039 , \3512_b0 );
or ( \3514_b1 , \3460_b1 , w_11041 );
not ( w_11041 , w_11042 );
and ( \3514_b0 , \3460_b0 , w_11043 );
and ( w_11042 ,  , w_11043 );
buf ( w_11041 , \3513_b1 );
not ( w_11041 , w_11044 );
not (  , w_11045 );
and ( w_11044 , w_11045 , \3513_b0 );
or ( \3515_b1 , \3456_b1 , w_11047 );
not ( w_11047 , w_11048 );
and ( \3515_b0 , \3456_b0 , w_11049 );
and ( w_11048 ,  , w_11049 );
buf ( w_11047 , \3514_b1 );
not ( w_11047 , w_11050 );
not (  , w_11051 );
and ( w_11050 , w_11051 , \3514_b0 );
or ( \3516_b1 , \3451_b1 , w_11053 );
not ( w_11053 , w_11054 );
and ( \3516_b0 , \3451_b0 , w_11055 );
and ( w_11054 ,  , w_11055 );
buf ( w_11053 , \3515_b1 );
not ( w_11053 , w_11056 );
not (  , w_11057 );
and ( w_11056 , w_11057 , \3515_b0 );
or ( \3517_b1 , \3196_b1 , w_11059 );
not ( w_11059 , w_11060 );
and ( \3517_b0 , \3196_b0 , w_11061 );
and ( w_11060 ,  , w_11061 );
buf ( w_11059 , \a[15]_b1 );
not ( w_11059 , w_11062 );
not (  , w_11063 );
and ( w_11062 , w_11063 , \a[15]_b0 );
buf ( \3518_b1 , \2281_b1 );
not ( \3518_b1 , w_11064 );
not ( \3518_b0 , w_11065 );
and ( w_11064 , w_11065 , \2281_b0 );
or ( \3519_b1 , \3518_b1 , w_11067 );
not ( w_11067 , w_11068 );
and ( \3519_b0 , \3518_b0 , w_11069 );
and ( w_11068 ,  , w_11069 );
buf ( w_11067 , \1954_b1 );
not ( w_11067 , w_11070 );
not (  , w_11071 );
and ( w_11070 , w_11071 , \1954_b0 );
or ( \3520_b1 , \2863_b1 , w_11072 );
xor ( \3520_b0 , \2863_b0 , w_11074 );
not ( w_11074 , w_11075 );
and ( w_11075 , w_11072 , w_11073 );
buf ( w_11072 , \3519_b1 );
not ( w_11072 , w_11076 );
not ( w_11073 , w_11077 );
and ( w_11076 , w_11077 , \3519_b0 );
or ( \3521_b1 , \3520_b1 , \2413_b1 );
not ( \2413_b1 , w_11078 );
and ( \3521_b0 , \3520_b0 , w_11079 );
and ( w_11078 , w_11079 , \2413_b0 );
buf ( \3522_b1 , \1538_b1 );
not ( \3522_b1 , w_11080 );
not ( \3522_b0 , w_11081 );
and ( w_11080 , w_11081 , \1538_b0 );
or ( \3523_b1 , \3522_b1 , w_11083 );
not ( w_11083 , w_11084 );
and ( \3523_b0 , \3522_b0 , w_11085 );
and ( w_11084 ,  , w_11085 );
buf ( w_11083 , \1214_b1 );
not ( w_11083 , w_11086 );
not (  , w_11087 );
and ( w_11086 , w_11087 , \1214_b0 );
buf ( \3524_b1 , \3523_b1 );
not ( \3524_b1 , w_11088 );
not ( \3524_b0 , w_11089 );
and ( w_11088 , w_11089 , \3523_b0 );
buf ( \3525_b1 , \2846_b1 );
not ( \3525_b1 , w_11090 );
not ( \3525_b0 , w_11091 );
and ( w_11090 , w_11091 , \2846_b0 );
or ( \3526_b1 , \3524_b1 , w_11092 );
or ( \3526_b0 , \3524_b0 , \3525_b0 );
not ( \3525_b0 , w_11093 );
and ( w_11093 , w_11092 , \3525_b1 );
or ( \3527_b1 , \2846_b1 , w_11094 );
or ( \3527_b0 , \2846_b0 , \3523_b0 );
not ( \3523_b0 , w_11095 );
and ( w_11095 , w_11094 , \3523_b1 );
or ( \3528_b1 , \3526_b1 , w_11097 );
not ( w_11097 , w_11098 );
and ( \3528_b0 , \3526_b0 , w_11099 );
and ( w_11098 ,  , w_11099 );
buf ( w_11097 , \3527_b1 );
not ( w_11097 , w_11100 );
not (  , w_11101 );
and ( w_11100 , w_11101 , \3527_b0 );
or ( \3529_b1 , \3528_b1 , \1668_b1 );
not ( \1668_b1 , w_11102 );
and ( \3529_b0 , \3528_b0 , w_11103 );
and ( w_11102 , w_11103 , \1668_b0 );
or ( \3530_b1 , \3521_b1 , w_11105 );
not ( w_11105 , w_11106 );
and ( \3530_b0 , \3521_b0 , w_11107 );
and ( w_11106 ,  , w_11107 );
buf ( w_11105 , \3529_b1 );
not ( w_11105 , w_11108 );
not (  , w_11109 );
and ( w_11108 , w_11109 , \3529_b0 );
or ( \3531_b1 , \b[10]_b1 , \c[10]_b1 );
not ( \c[10]_b1 , w_11110 );
and ( \3531_b0 , \b[10]_b0 , w_11111 );
and ( w_11110 , w_11111 , \c[10]_b0 );
or ( \3532_b1 , \922_b1 , w_11113 );
not ( w_11113 , w_11114 );
and ( \3532_b0 , \922_b0 , w_11115 );
and ( w_11114 ,  , w_11115 );
buf ( w_11113 , \3531_b1 );
not ( w_11113 , w_11116 );
not (  , w_11117 );
and ( w_11116 , w_11117 , \3531_b0 );
or ( \3533_b1 , \c[10]_b1 , \d[10]_b1 );
xor ( \3533_b0 , \c[10]_b0 , w_11118 );
not ( w_11118 , w_11119 );
and ( w_11119 , \d[10]_b1 , \d[10]_b0 );
or ( \3534_b1 , \2615_b1 , \3533_b1 );
not ( \3533_b1 , w_11120 );
and ( \3534_b0 , \2615_b0 , w_11121 );
and ( w_11120 , w_11121 , \3533_b0 );
buf ( \3535_b1 , \771_b1 );
not ( \3535_b1 , w_11122 );
not ( \3535_b0 , w_11123 );
and ( w_11122 , w_11123 , \771_b0 );
or ( \3536_b1 , \3535_b1 , w_11125 );
not ( w_11125 , w_11126 );
and ( \3536_b0 , \3535_b0 , w_11127 );
and ( w_11126 ,  , w_11127 );
buf ( w_11125 , \749_b1 );
not ( w_11125 , w_11128 );
not (  , w_11129 );
and ( w_11128 , w_11129 , \749_b0 );
buf ( \3537_b1 , \3536_b1 );
not ( \3537_b1 , w_11130 );
not ( \3537_b0 , w_11131 );
and ( w_11130 , w_11131 , \3536_b0 );
or ( \3538_b1 , \747_b1 , \753_b1 );
not ( \753_b1 , w_11132 );
and ( \3538_b0 , \747_b0 , w_11133 );
and ( w_11132 , w_11133 , \753_b0 );
or ( \3539_b1 , \3538_b1 , w_11135 );
not ( w_11135 , w_11136 );
and ( \3539_b0 , \3538_b0 , w_11137 );
and ( w_11136 ,  , w_11137 );
buf ( w_11135 , \766_b1 );
not ( w_11135 , w_11138 );
not (  , w_11139 );
and ( w_11138 , w_11139 , \766_b0 );
buf ( \3540_b1 , \3539_b1 );
not ( \3540_b1 , w_11140 );
not ( \3540_b0 , w_11141 );
and ( w_11140 , w_11141 , \3539_b0 );
or ( \3541_b1 , \3537_b1 , w_11142 );
or ( \3541_b0 , \3537_b0 , \3540_b0 );
not ( \3540_b0 , w_11143 );
and ( w_11143 , w_11142 , \3540_b1 );
or ( \3542_b1 , \3539_b1 , w_11144 );
or ( \3542_b0 , \3539_b0 , \3536_b0 );
not ( \3536_b0 , w_11145 );
and ( w_11145 , w_11144 , \3536_b1 );
or ( \3543_b1 , \3541_b1 , w_11147 );
not ( w_11147 , w_11148 );
and ( \3543_b0 , \3541_b0 , w_11149 );
and ( w_11148 ,  , w_11149 );
buf ( w_11147 , \3542_b1 );
not ( w_11147 , w_11150 );
not (  , w_11151 );
and ( w_11150 , w_11151 , \3542_b0 );
buf ( \3544_b1 , \3543_b1 );
not ( \3544_b1 , w_11152 );
not ( \3544_b0 , w_11153 );
and ( w_11152 , w_11153 , \3543_b0 );
buf ( \3545_b1 , \707_b1 );
not ( \3545_b1 , w_11154 );
not ( \3545_b0 , w_11155 );
and ( w_11154 , w_11155 , \707_b0 );
or ( \3546_b1 , \3544_b1 , w_11156 );
or ( \3546_b0 , \3544_b0 , \3545_b0 );
not ( \3545_b0 , w_11157 );
and ( w_11157 , w_11156 , \3545_b1 );
buf ( \3547_b1 , \856_b1 );
not ( \3547_b1 , w_11158 );
not ( \3547_b0 , w_11159 );
and ( w_11158 , w_11159 , \856_b0 );
or ( \3548_b1 , \3547_b1 , w_11161 );
not ( w_11161 , w_11162 );
and ( \3548_b0 , \3547_b0 , w_11163 );
and ( w_11162 ,  , w_11163 );
buf ( w_11161 , \834_b1 );
not ( w_11161 , w_11164 );
not (  , w_11165 );
and ( w_11164 , w_11165 , \834_b0 );
buf ( \3549_b1 , \3548_b1 );
not ( \3549_b1 , w_11166 );
not ( \3549_b0 , w_11167 );
and ( w_11166 , w_11167 , \3548_b0 );
or ( \3550_b1 , \832_b1 , \838_b1 );
not ( \838_b1 , w_11168 );
and ( \3550_b0 , \832_b0 , w_11169 );
and ( w_11168 , w_11169 , \838_b0 );
or ( \3551_b1 , \3550_b1 , w_11171 );
not ( w_11171 , w_11172 );
and ( \3551_b0 , \3550_b0 , w_11173 );
and ( w_11172 ,  , w_11173 );
buf ( w_11171 , \851_b1 );
not ( w_11171 , w_11174 );
not (  , w_11175 );
and ( w_11174 , w_11175 , \851_b0 );
buf ( \3552_b1 , \3551_b1 );
not ( \3552_b1 , w_11176 );
not ( \3552_b0 , w_11177 );
and ( w_11176 , w_11177 , \3551_b0 );
or ( \3553_b1 , \3549_b1 , w_11178 );
or ( \3553_b0 , \3549_b0 , \3552_b0 );
not ( \3552_b0 , w_11179 );
and ( w_11179 , w_11178 , \3552_b1 );
or ( \3554_b1 , \3551_b1 , w_11180 );
or ( \3554_b0 , \3551_b0 , \3548_b0 );
not ( \3548_b0 , w_11181 );
and ( w_11181 , w_11180 , \3548_b1 );
or ( \3555_b1 , \3553_b1 , w_11183 );
not ( w_11183 , w_11184 );
and ( \3555_b0 , \3553_b0 , w_11185 );
and ( w_11184 ,  , w_11185 );
buf ( w_11183 , \3554_b1 );
not ( w_11183 , w_11186 );
not (  , w_11187 );
and ( w_11186 , w_11187 , \3554_b0 );
or ( \3556_b1 , \880_b1 , \3555_b1 );
not ( \3555_b1 , w_11188 );
and ( \3556_b0 , \880_b0 , w_11189 );
and ( w_11188 , w_11189 , \3555_b0 );
buf ( \3557_b1 , \d[10]_b1 );
not ( \3557_b1 , w_11190 );
not ( \3557_b0 , w_11191 );
and ( w_11190 , w_11191 , \d[10]_b0 );
buf ( \3558_b1 , \894_b1 );
not ( \3558_b1 , w_11192 );
not ( \3558_b0 , w_11193 );
and ( w_11192 , w_11193 , \894_b0 );
or ( \3559_b1 , \3557_b1 , w_11194 );
or ( \3559_b0 , \3557_b0 , \3558_b0 );
not ( \3558_b0 , w_11195 );
and ( w_11195 , w_11194 , \3558_b1 );
or ( \3560_b1 , \885_b1 , \b[10]_b1 );
not ( \b[10]_b1 , w_11196 );
and ( \3560_b0 , \885_b0 , w_11197 );
and ( w_11196 , w_11197 , \b[10]_b0 );
or ( \3561_b1 , \907_b1 , \c[10]_b1 );
not ( \c[10]_b1 , w_11198 );
and ( \3561_b0 , \907_b0 , w_11199 );
and ( w_11198 , w_11199 , \c[10]_b0 );
or ( \3562_b1 , \3560_b1 , w_11201 );
not ( w_11201 , w_11202 );
and ( \3562_b0 , \3560_b0 , w_11203 );
and ( w_11202 ,  , w_11203 );
buf ( w_11201 , \3561_b1 );
not ( w_11201 , w_11204 );
not (  , w_11205 );
and ( w_11204 , w_11205 , \3561_b0 );
or ( \3563_b1 , \3559_b1 , w_11207 );
not ( w_11207 , w_11208 );
and ( \3563_b0 , \3559_b0 , w_11209 );
and ( w_11208 ,  , w_11209 );
buf ( w_11207 , \3562_b1 );
not ( w_11207 , w_11210 );
not (  , w_11211 );
and ( w_11210 , w_11211 , \3562_b0 );
or ( \3564_b1 , \3556_b1 , w_11213 );
not ( w_11213 , w_11214 );
and ( \3564_b0 , \3556_b0 , w_11215 );
and ( w_11214 ,  , w_11215 );
buf ( w_11213 , \3563_b1 );
not ( w_11213 , w_11216 );
not (  , w_11217 );
and ( w_11216 , w_11217 , \3563_b0 );
or ( \3565_b1 , \3546_b1 , w_11219 );
not ( w_11219 , w_11220 );
and ( \3565_b0 , \3546_b0 , w_11221 );
and ( w_11220 ,  , w_11221 );
buf ( w_11219 , \3564_b1 );
not ( w_11219 , w_11222 );
not (  , w_11223 );
and ( w_11222 , w_11223 , \3564_b0 );
or ( \3566_b1 , \3534_b1 , w_11225 );
not ( w_11225 , w_11226 );
and ( \3566_b0 , \3534_b0 , w_11227 );
and ( w_11226 ,  , w_11227 );
buf ( w_11225 , \3565_b1 );
not ( w_11225 , w_11228 );
not (  , w_11229 );
and ( w_11228 , w_11229 , \3565_b0 );
buf ( \3568_b1 , \672_b1 );
not ( \3568_b1 , w_11230 );
not ( \3568_b0 , w_11231 );
and ( w_11230 , w_11231 , \672_b0 );
or ( \3569_b1 , \3568_b1 , w_11233 );
not ( w_11233 , w_11234 );
and ( \3569_b0 , \3568_b0 , w_11235 );
and ( w_11234 ,  , w_11235 );
buf ( w_11233 , \3235_b1 );
not ( w_11233 , w_11236 );
not (  , w_11237 );
and ( w_11236 , w_11237 , \3235_b0 );
or ( \3570_b1 , \2859_b1 , w_11239 );
not ( w_11239 , w_11240 );
and ( \3570_b0 , \2859_b0 , w_11241 );
and ( w_11240 ,  , w_11241 );
buf ( w_11239 , \a[10]_b1 );
not ( w_11239 , w_11242 );
not (  , w_11243 );
and ( w_11242 , w_11243 , \a[10]_b0 );
or ( \3571_b1 , \a[10]_b1 , w_11244 );
or ( \3571_b0 , \a[10]_b0 , \b[10]_b0 );
not ( \b[10]_b0 , w_11245 );
and ( w_11245 , w_11244 , \b[10]_b1 );
or ( \3572_b1 , \2791_b1 , w_11247 );
not ( w_11247 , w_11248 );
and ( \3572_b0 , \2791_b0 , w_11249 );
and ( w_11248 ,  , w_11249 );
buf ( w_11247 , \3571_b1 );
not ( w_11247 , w_11250 );
not (  , w_11251 );
and ( w_11250 , w_11251 , \3571_b0 );
or ( \3574_b1 , \b[9]_b1 , \c[9]_b1 );
not ( \c[9]_b1 , w_11252 );
and ( \3574_b0 , \b[9]_b0 , w_11253 );
and ( w_11252 , w_11253 , \c[9]_b0 );
or ( \3575_b1 , \2887_b1 , \3574_b1 );
not ( \3574_b1 , w_11254 );
and ( \3575_b0 , \2887_b0 , w_11255 );
and ( w_11254 , w_11255 , \3574_b0 );
buf ( \3576_b1 , \3124_b1 );
not ( \3576_b1 , w_11256 );
not ( \3576_b0 , w_11257 );
and ( w_11256 , w_11257 , \3124_b0 );
buf ( \3577_b1 , \2270_b1 );
not ( \3577_b1 , w_11258 );
not ( \3577_b0 , w_11259 );
and ( w_11258 , w_11259 , \2270_b0 );
or ( \3578_b1 , \3576_b1 , w_11260 );
or ( \3578_b0 , \3576_b0 , \3577_b0 );
not ( \3577_b0 , w_11261 );
and ( w_11261 , w_11260 , \3577_b1 );
or ( \3579_b1 , \3578_b1 , w_11263 );
not ( w_11263 , w_11264 );
and ( \3579_b0 , \3578_b0 , w_11265 );
and ( w_11264 ,  , w_11265 );
buf ( w_11263 , \3125_b1 );
not ( w_11263 , w_11266 );
not (  , w_11267 );
and ( w_11266 , w_11267 , \3125_b0 );
buf ( \3580_b1 , \2048_b1 );
not ( \3580_b1 , w_11268 );
not ( \3580_b0 , w_11269 );
and ( w_11268 , w_11269 , \2048_b0 );
or ( \3581_b1 , \3580_b1 , w_11271 );
not ( w_11271 , w_11272 );
and ( \3581_b0 , \3580_b0 , w_11273 );
and ( w_11272 ,  , w_11273 );
buf ( w_11271 , \2279_b1 );
not ( w_11271 , w_11274 );
not (  , w_11275 );
and ( w_11274 , w_11275 , \2279_b0 );
or ( \3582_b1 , \3579_b1 , w_11276 );
xor ( \3582_b0 , \3579_b0 , w_11278 );
not ( w_11278 , w_11279 );
and ( w_11279 , w_11276 , w_11277 );
buf ( w_11276 , \3581_b1 );
not ( w_11276 , w_11280 );
not ( w_11277 , w_11281 );
and ( w_11280 , w_11281 , \3581_b0 );
buf ( \3583_b1 , \3582_b1 );
not ( \3583_b1 , w_11282 );
not ( \3583_b0 , w_11283 );
and ( w_11282 , w_11283 , \3582_b0 );
or ( \3584_b1 , \3583_b1 , w_11285 );
not ( w_11285 , w_11286 );
and ( \3584_b0 , \3583_b0 , w_11287 );
and ( w_11286 ,  , w_11287 );
buf ( w_11285 , \2412_b1 );
not ( w_11285 , w_11288 );
not (  , w_11289 );
and ( w_11288 , w_11289 , \2412_b0 );
or ( \3585_b1 , \3575_b1 , w_11291 );
not ( w_11291 , w_11292 );
and ( \3585_b0 , \3575_b0 , w_11293 );
and ( w_11292 ,  , w_11293 );
buf ( w_11291 , \3584_b1 );
not ( w_11291 , w_11294 );
not (  , w_11295 );
and ( w_11294 , w_11295 , \3584_b0 );
or ( \3586_b1 , \a[9]_b1 , w_11296 );
or ( \3586_b0 , \a[9]_b0 , \b[9]_b0 );
not ( \b[9]_b0 , w_11297 );
and ( w_11297 , w_11296 , \b[9]_b1 );
or ( \3587_b1 , \667_b1 , \3586_b1 );
not ( \3586_b1 , w_11298 );
and ( \3587_b0 , \667_b0 , w_11299 );
and ( w_11298 , w_11299 , \3586_b0 );
buf ( \3588_b1 , \1308_b1 );
not ( \3588_b1 , w_11300 );
not ( \3588_b0 , w_11301 );
and ( w_11300 , w_11301 , \1308_b0 );
or ( \3589_b1 , \3588_b1 , w_11303 );
not ( w_11303 , w_11304 );
and ( \3589_b0 , \3588_b0 , w_11305 );
and ( w_11304 ,  , w_11305 );
buf ( w_11303 , \1536_b1 );
not ( w_11303 , w_11306 );
not (  , w_11307 );
and ( w_11306 , w_11307 , \1536_b0 );
buf ( \3590_b1 , \3589_b1 );
not ( \3590_b1 , w_11308 );
not ( \3590_b0 , w_11309 );
and ( w_11308 , w_11309 , \3589_b0 );
buf ( \3591_b1 , \3088_b1 );
not ( \3591_b1 , w_11310 );
not ( \3591_b0 , w_11311 );
and ( w_11310 , w_11311 , \3088_b0 );
buf ( \3592_b1 , \1527_b1 );
not ( \3592_b1 , w_11312 );
not ( \3592_b0 , w_11313 );
and ( w_11312 , w_11313 , \1527_b0 );
or ( \3593_b1 , \3591_b1 , w_11314 );
or ( \3593_b0 , \3591_b0 , \3592_b0 );
not ( \3592_b0 , w_11315 );
and ( w_11315 , w_11314 , \3592_b1 );
or ( \3594_b1 , \3593_b1 , w_11317 );
not ( w_11317 , w_11318 );
and ( \3594_b0 , \3593_b0 , w_11319 );
and ( w_11318 ,  , w_11319 );
buf ( w_11317 , \3089_b1 );
not ( w_11317 , w_11320 );
not (  , w_11321 );
and ( w_11320 , w_11321 , \3089_b0 );
buf ( \3595_b1 , \3594_b1 );
not ( \3595_b1 , w_11322 );
not ( \3595_b0 , w_11323 );
and ( w_11322 , w_11323 , \3594_b0 );
or ( \3596_b1 , \3590_b1 , w_11324 );
or ( \3596_b0 , \3590_b0 , \3595_b0 );
not ( \3595_b0 , w_11325 );
and ( w_11325 , w_11324 , \3595_b1 );
or ( \3597_b1 , \3594_b1 , w_11326 );
or ( \3597_b0 , \3594_b0 , \3589_b0 );
not ( \3589_b0 , w_11327 );
and ( w_11327 , w_11326 , \3589_b1 );
or ( \3598_b1 , \3596_b1 , w_11329 );
not ( w_11329 , w_11330 );
and ( \3598_b0 , \3596_b0 , w_11331 );
and ( w_11330 ,  , w_11331 );
buf ( w_11329 , \3597_b1 );
not ( w_11329 , w_11332 );
not (  , w_11333 );
and ( w_11332 , w_11333 , \3597_b0 );
or ( \3599_b1 , \3598_b1 , w_11335 );
not ( w_11335 , w_11336 );
and ( \3599_b0 , \3598_b0 , w_11337 );
and ( w_11336 ,  , w_11337 );
buf ( w_11335 , \1668_b1 );
not ( w_11335 , w_11338 );
not (  , w_11339 );
and ( w_11338 , w_11339 , \1668_b0 );
or ( \3600_b1 , \c[9]_b1 , \d[9]_b1 );
xor ( \3600_b0 , \c[9]_b0 , w_11340 );
not ( w_11340 , w_11341 );
and ( w_11341 , \d[9]_b1 , \d[9]_b0 );
or ( \3601_b1 , \2614_b1 , w_11343 );
not ( w_11343 , w_11344 );
and ( \3601_b0 , \2614_b0 , w_11345 );
and ( w_11344 ,  , w_11345 );
buf ( w_11343 , \3600_b1 );
not ( w_11343 , w_11346 );
not (  , w_11347 );
and ( w_11346 , w_11347 , \3600_b0 );
buf ( \3602_b1 , \751_b1 );
not ( \3602_b1 , w_11348 );
not ( \3602_b0 , w_11349 );
and ( w_11348 , w_11349 , \751_b0 );
or ( \3603_b1 , \3602_b1 , w_11351 );
not ( w_11351 , w_11352 );
and ( \3603_b0 , \3602_b0 , w_11353 );
and ( w_11352 ,  , w_11353 );
buf ( w_11351 , \765_b1 );
not ( w_11351 , w_11354 );
not (  , w_11355 );
and ( w_11354 , w_11355 , \765_b0 );
buf ( \3604_b1 , \3603_b1 );
not ( \3604_b1 , w_11356 );
not ( \3604_b0 , w_11357 );
and ( w_11356 , w_11357 , \3603_b0 );
buf ( \3605_b1 , \747_b1 );
not ( \3605_b1 , w_11358 );
not ( \3605_b0 , w_11359 );
and ( w_11358 , w_11359 , \747_b0 );
or ( \3606_b1 , \3605_b1 , w_11360 );
or ( \3606_b0 , \3605_b0 , \752_b0 );
not ( \752_b0 , w_11361 );
and ( w_11361 , w_11360 , \752_b1 );
or ( \3607_b1 , \3606_b1 , w_11363 );
not ( w_11363 , w_11364 );
and ( \3607_b0 , \3606_b0 , w_11365 );
and ( w_11364 ,  , w_11365 );
buf ( w_11363 , \763_b1 );
not ( w_11363 , w_11366 );
not (  , w_11367 );
and ( w_11366 , w_11367 , \763_b0 );
buf ( \3608_b1 , \3607_b1 );
not ( \3608_b1 , w_11368 );
not ( \3608_b0 , w_11369 );
and ( w_11368 , w_11369 , \3607_b0 );
or ( \3609_b1 , \3604_b1 , w_11370 );
or ( \3609_b0 , \3604_b0 , \3608_b0 );
not ( \3608_b0 , w_11371 );
and ( w_11371 , w_11370 , \3608_b1 );
or ( \3610_b1 , \3607_b1 , w_11372 );
or ( \3610_b0 , \3607_b0 , \3603_b0 );
not ( \3603_b0 , w_11373 );
and ( w_11373 , w_11372 , \3603_b1 );
or ( \3611_b1 , \3609_b1 , w_11375 );
not ( w_11375 , w_11376 );
and ( \3611_b0 , \3609_b0 , w_11377 );
and ( w_11376 ,  , w_11377 );
buf ( w_11375 , \3610_b1 );
not ( w_11375 , w_11378 );
not (  , w_11379 );
and ( w_11378 , w_11379 , \3610_b0 );
or ( \3612_b1 , \707_b1 , \3611_b1 );
not ( \3611_b1 , w_11380 );
and ( \3612_b0 , \707_b0 , w_11381 );
and ( w_11380 , w_11381 , \3611_b0 );
buf ( \3613_b1 , \836_b1 );
not ( \3613_b1 , w_11382 );
not ( \3613_b0 , w_11383 );
and ( w_11382 , w_11383 , \836_b0 );
or ( \3614_b1 , \3613_b1 , w_11385 );
not ( w_11385 , w_11386 );
and ( \3614_b0 , \3613_b0 , w_11387 );
and ( w_11386 ,  , w_11387 );
buf ( w_11385 , \850_b1 );
not ( w_11385 , w_11388 );
not (  , w_11389 );
and ( w_11388 , w_11389 , \850_b0 );
buf ( \3615_b1 , \3614_b1 );
not ( \3615_b1 , w_11390 );
not ( \3615_b0 , w_11391 );
and ( w_11390 , w_11391 , \3614_b0 );
buf ( \3616_b1 , \832_b1 );
not ( \3616_b1 , w_11392 );
not ( \3616_b0 , w_11393 );
and ( w_11392 , w_11393 , \832_b0 );
or ( \3617_b1 , \3616_b1 , w_11394 );
or ( \3617_b0 , \3616_b0 , \837_b0 );
not ( \837_b0 , w_11395 );
and ( w_11395 , w_11394 , \837_b1 );
or ( \3618_b1 , \3617_b1 , w_11397 );
not ( w_11397 , w_11398 );
and ( \3618_b0 , \3617_b0 , w_11399 );
and ( w_11398 ,  , w_11399 );
buf ( w_11397 , \848_b1 );
not ( w_11397 , w_11400 );
not (  , w_11401 );
and ( w_11400 , w_11401 , \848_b0 );
buf ( \3619_b1 , \3618_b1 );
not ( \3619_b1 , w_11402 );
not ( \3619_b0 , w_11403 );
and ( w_11402 , w_11403 , \3618_b0 );
or ( \3620_b1 , \3615_b1 , w_11404 );
or ( \3620_b0 , \3615_b0 , \3619_b0 );
not ( \3619_b0 , w_11405 );
and ( w_11405 , w_11404 , \3619_b1 );
or ( \3621_b1 , \3618_b1 , w_11406 );
or ( \3621_b0 , \3618_b0 , \3614_b0 );
not ( \3614_b0 , w_11407 );
and ( w_11407 , w_11406 , \3614_b1 );
or ( \3622_b1 , \3620_b1 , w_11409 );
not ( w_11409 , w_11410 );
and ( \3622_b0 , \3620_b0 , w_11411 );
and ( w_11410 ,  , w_11411 );
buf ( w_11409 , \3621_b1 );
not ( w_11409 , w_11412 );
not (  , w_11413 );
and ( w_11412 , w_11413 , \3621_b0 );
buf ( \3623_b1 , \3622_b1 );
not ( \3623_b1 , w_11414 );
not ( \3623_b0 , w_11415 );
and ( w_11414 , w_11415 , \3622_b0 );
buf ( \3624_b1 , \880_b1 );
not ( \3624_b1 , w_11416 );
not ( \3624_b0 , w_11417 );
and ( w_11416 , w_11417 , \880_b0 );
or ( \3625_b1 , \3623_b1 , w_11418 );
or ( \3625_b0 , \3623_b0 , \3624_b0 );
not ( \3624_b0 , w_11419 );
and ( w_11419 , w_11418 , \3624_b1 );
or ( \3626_b1 , \894_b1 , \d[9]_b1 );
not ( \d[9]_b1 , w_11420 );
and ( \3626_b0 , \894_b0 , w_11421 );
and ( w_11420 , w_11421 , \d[9]_b0 );
or ( \3627_b1 , \b[9]_b1 , \885_b1 );
not ( \885_b1 , w_11422 );
and ( \3627_b0 , \b[9]_b0 , w_11423 );
and ( w_11422 , w_11423 , \885_b0 );
or ( \3628_b1 , \907_b1 , \c[9]_b1 );
not ( \c[9]_b1 , w_11424 );
and ( \3628_b0 , \907_b0 , w_11425 );
and ( w_11424 , w_11425 , \c[9]_b0 );
or ( \3630_b1 , \3625_b1 , w_11427 );
not ( w_11427 , w_11428 );
and ( \3630_b0 , \3625_b0 , w_11429 );
and ( w_11428 ,  , w_11429 );
buf ( w_11427 , \3629_b1 );
not ( w_11427 , w_11430 );
not (  , w_11431 );
and ( w_11430 , w_11431 , \3629_b0 );
or ( \3631_b1 , \3612_b1 , w_11433 );
not ( w_11433 , w_11434 );
and ( \3631_b0 , \3612_b0 , w_11435 );
and ( w_11434 ,  , w_11435 );
buf ( w_11433 , \3630_b1 );
not ( w_11433 , w_11436 );
not (  , w_11437 );
and ( w_11436 , w_11437 , \3630_b0 );
or ( \3633_b1 , \3587_b1 , w_11439 );
not ( w_11439 , w_11440 );
and ( \3633_b0 , \3587_b0 , w_11441 );
and ( w_11440 ,  , w_11441 );
buf ( w_11439 , \3632_b1 );
not ( w_11439 , w_11442 );
not (  , w_11443 );
and ( w_11442 , w_11443 , \3632_b0 );
or ( \3634_b1 , \2858_b1 , w_11445 );
not ( w_11445 , w_11446 );
and ( \3634_b0 , \2858_b0 , w_11447 );
and ( w_11446 ,  , w_11447 );
buf ( w_11445 , \a[9]_b1 );
not ( w_11445 , w_11448 );
not (  , w_11449 );
and ( w_11448 , w_11449 , \a[9]_b0 );
buf ( \3635_b1 , \673_b1 );
not ( \3635_b1 , w_11450 );
not ( \3635_b0 , w_11451 );
and ( w_11450 , w_11451 , \673_b0 );
or ( \3636_b1 , \2843_b1 , w_11453 );
not ( w_11453 , w_11454 );
and ( \3636_b0 , \2843_b0 , w_11455 );
and ( w_11454 ,  , w_11455 );
buf ( w_11453 , \3635_b1 );
not ( w_11453 , w_11456 );
not (  , w_11457 );
and ( w_11456 , w_11457 , \3635_b0 );
buf ( \3638_b1 , \2129_b1 );
not ( \3638_b1 , w_11458 );
not ( \3638_b0 , w_11459 );
and ( w_11458 , w_11459 , \2129_b0 );
or ( \3639_b1 , \3638_b1 , w_11461 );
not ( w_11461 , w_11462 );
and ( \3639_b0 , \3638_b0 , w_11463 );
and ( w_11462 ,  , w_11463 );
buf ( w_11461 , \2287_b1 );
not ( w_11461 , w_11464 );
not (  , w_11465 );
and ( w_11464 , w_11465 , \2287_b0 );
buf ( \3640_b1 , \3639_b1 );
not ( \3640_b1 , w_11466 );
not ( \3640_b0 , w_11467 );
and ( w_11466 , w_11467 , \3639_b0 );
or ( \3641_b1 , \2592_b1 , w_11469 );
not ( w_11469 , w_11470 );
and ( \3641_b0 , \2592_b0 , w_11471 );
and ( w_11470 ,  , w_11471 );
buf ( w_11469 , \2284_b1 );
not ( w_11469 , w_11472 );
not (  , w_11473 );
and ( w_11472 , w_11473 , \2284_b0 );
buf ( \3642_b1 , \3641_b1 );
not ( \3642_b1 , w_11474 );
not ( \3642_b0 , w_11475 );
and ( w_11474 , w_11475 , \3641_b0 );
or ( \3643_b1 , \3640_b1 , w_11476 );
or ( \3643_b0 , \3640_b0 , \3642_b0 );
not ( \3642_b0 , w_11477 );
and ( w_11477 , w_11476 , \3642_b1 );
or ( \3644_b1 , \3641_b1 , w_11478 );
or ( \3644_b0 , \3641_b0 , \3639_b0 );
not ( \3639_b0 , w_11479 );
and ( w_11479 , w_11478 , \3639_b1 );
or ( \3645_b1 , \3643_b1 , w_11481 );
not ( w_11481 , w_11482 );
and ( \3645_b0 , \3643_b0 , w_11483 );
and ( w_11482 ,  , w_11483 );
buf ( w_11481 , \3644_b1 );
not ( w_11481 , w_11484 );
not (  , w_11485 );
and ( w_11484 , w_11485 , \3644_b0 );
or ( \3646_b1 , \3645_b1 , \2413_b1 );
not ( \2413_b1 , w_11486 );
and ( \3646_b0 , \3645_b0 , w_11487 );
and ( w_11486 , w_11487 , \2413_b0 );
buf ( \3647_b1 , \1388_b1 );
not ( \3647_b1 , w_11488 );
not ( \3647_b0 , w_11489 );
and ( w_11488 , w_11489 , \1388_b0 );
or ( \3648_b1 , \3647_b1 , w_11491 );
not ( w_11491 , w_11492 );
and ( \3648_b0 , \3647_b0 , w_11493 );
and ( w_11492 ,  , w_11493 );
buf ( w_11491 , \2777_b1 );
not ( w_11491 , w_11494 );
not (  , w_11495 );
and ( w_11494 , w_11495 , \2777_b0 );
buf ( \3649_b1 , \3648_b1 );
not ( \3649_b1 , w_11496 );
not ( \3649_b0 , w_11497 );
and ( w_11496 , w_11497 , \3648_b0 );
or ( \3650_b1 , \2774_b1 , w_11499 );
not ( w_11499 , w_11500 );
and ( \3650_b0 , \2774_b0 , w_11501 );
and ( w_11500 ,  , w_11501 );
buf ( w_11499 , \1541_b1 );
not ( w_11499 , w_11502 );
not (  , w_11503 );
and ( w_11502 , w_11503 , \1541_b0 );
buf ( \3651_b1 , \3650_b1 );
not ( \3651_b1 , w_11504 );
not ( \3651_b0 , w_11505 );
and ( w_11504 , w_11505 , \3650_b0 );
or ( \3652_b1 , \3649_b1 , w_11506 );
or ( \3652_b0 , \3649_b0 , \3651_b0 );
not ( \3651_b0 , w_11507 );
and ( w_11507 , w_11506 , \3651_b1 );
or ( \3653_b1 , \3650_b1 , w_11508 );
or ( \3653_b0 , \3650_b0 , \3648_b0 );
not ( \3648_b0 , w_11509 );
and ( w_11509 , w_11508 , \3648_b1 );
or ( \3654_b1 , \3652_b1 , w_11511 );
not ( w_11511 , w_11512 );
and ( \3654_b0 , \3652_b0 , w_11513 );
and ( w_11512 ,  , w_11513 );
buf ( w_11511 , \3653_b1 );
not ( w_11511 , w_11514 );
not (  , w_11515 );
and ( w_11514 , w_11515 , \3653_b0 );
or ( \3655_b1 , \3654_b1 , \1668_b1 );
not ( \1668_b1 , w_11516 );
and ( \3655_b0 , \3654_b0 , w_11517 );
and ( w_11516 , w_11517 , \1668_b0 );
or ( \3656_b1 , \3646_b1 , w_11519 );
not ( w_11519 , w_11520 );
and ( \3656_b0 , \3646_b0 , w_11521 );
and ( w_11520 ,  , w_11521 );
buf ( w_11519 , \3655_b1 );
not ( w_11519 , w_11522 );
not (  , w_11523 );
and ( w_11522 , w_11523 , \3655_b0 );
or ( \3658_b1 , \1539_b1 , \2770_b1 );
not ( \2770_b1 , w_11524 );
and ( \3658_b0 , \1539_b0 , w_11525 );
and ( w_11524 , w_11525 , \2770_b0 );
or ( \3659_b1 , \1388_b1 , w_11527 );
not ( w_11527 , w_11528 );
and ( \3659_b0 , \1388_b0 , w_11529 );
and ( w_11528 ,  , w_11529 );
buf ( w_11527 , \1214_b1 );
not ( w_11527 , w_11530 );
not (  , w_11531 );
and ( w_11530 , w_11531 , \1214_b0 );
or ( \3660_b1 , \3658_b1 , w_11532 );
or ( \3660_b0 , \3658_b0 , \3659_b0 );
not ( \3659_b0 , w_11533 );
and ( w_11533 , w_11532 , \3659_b1 );
or ( \3661_b1 , \1388_b1 , w_11535 );
not ( w_11535 , w_11536 );
and ( \3661_b0 , \1388_b0 , w_11537 );
and ( w_11536 ,  , w_11537 );
buf ( w_11535 , \1530_b1 );
not ( w_11535 , w_11538 );
not (  , w_11539 );
and ( w_11538 , w_11539 , \1530_b0 );
or ( \3662_b1 , \3660_b1 , w_11541 );
not ( w_11541 , w_11542 );
and ( \3662_b0 , \3660_b0 , w_11543 );
and ( w_11542 ,  , w_11543 );
buf ( w_11541 , \3661_b1 );
not ( w_11541 , w_11544 );
not (  , w_11545 );
and ( w_11544 , w_11545 , \3661_b0 );
or ( \3663_b1 , \3657_b1 , \3662_b1 );
not ( \3662_b1 , w_11546 );
and ( \3663_b0 , \3657_b0 , w_11547 );
and ( w_11546 , w_11547 , \3662_b0 );
buf ( \3664_b1 , \2781_b1 );
not ( \3664_b1 , w_11548 );
not ( \3664_b0 , w_11549 );
and ( w_11548 , w_11549 , \2781_b0 );
buf ( \3665_b1 , \2763_b1 );
not ( \3665_b1 , w_11550 );
not ( \3665_b0 , w_11551 );
and ( w_11550 , w_11551 , \2763_b0 );
or ( \3666_b1 , \3664_b1 , w_11552 );
or ( \3666_b0 , \3664_b0 , \3665_b0 );
not ( \3665_b0 , w_11553 );
and ( w_11553 , w_11552 , \3665_b1 );
or ( \3667_b1 , \3666_b1 , w_11555 );
not ( w_11555 , w_11556 );
and ( \3667_b0 , \3666_b0 , w_11557 );
and ( w_11556 ,  , w_11557 );
buf ( w_11555 , \2761_b1 );
not ( w_11555 , w_11558 );
not (  , w_11559 );
and ( w_11558 , w_11559 , \2761_b0 );
or ( \3668_b1 , \3663_b1 , w_11561 );
not ( w_11561 , w_11562 );
and ( \3668_b0 , \3663_b0 , w_11563 );
and ( w_11562 ,  , w_11563 );
buf ( w_11561 , \3667_b1 );
not ( w_11561 , w_11564 );
not (  , w_11565 );
and ( w_11564 , w_11565 , \3667_b0 );
buf ( \3669_b1 , \2737_b1 );
not ( \3669_b1 , w_11566 );
not ( \3669_b0 , w_11567 );
and ( w_11566 , w_11567 , \2737_b0 );
buf ( \3670_b1 , \3669_b1 );
not ( \3670_b1 , w_11568 );
not ( \3670_b0 , w_11569 );
and ( w_11568 , w_11569 , \3669_b0 );
buf ( \3671_b1 , \2709_b1 );
not ( \3671_b1 , w_11570 );
not ( \3671_b0 , w_11571 );
and ( w_11570 , w_11571 , \2709_b0 );
or ( \3672_b1 , \3670_b1 , w_11572 );
or ( \3672_b0 , \3670_b0 , \3671_b0 );
not ( \3671_b0 , w_11573 );
and ( w_11573 , w_11572 , \3671_b1 );
or ( \3673_b1 , \3672_b1 , w_11575 );
not ( w_11575 , w_11576 );
and ( \3673_b0 , \3672_b0 , w_11577 );
and ( w_11576 ,  , w_11577 );
buf ( w_11575 , \2748_b1 );
not ( w_11575 , w_11578 );
not (  , w_11579 );
and ( w_11578 , w_11579 , \2748_b0 );
buf ( \3674_b1 , \2709_b1 );
not ( \3674_b1 , w_11580 );
not ( \3674_b0 , w_11581 );
and ( w_11580 , w_11581 , \2709_b0 );
or ( \3675_b1 , \3674_b1 , w_11583 );
not ( w_11583 , w_11584 );
and ( \3675_b0 , \3674_b0 , w_11585 );
and ( w_11584 ,  , w_11585 );
buf ( w_11583 , \2737_b1 );
not ( w_11583 , w_11586 );
not (  , w_11587 );
and ( w_11586 , w_11587 , \2737_b0 );
or ( \3676_b1 , \3673_b1 , w_11589 );
not ( w_11589 , w_11590 );
and ( \3676_b0 , \3673_b0 , w_11591 );
and ( w_11590 ,  , w_11591 );
buf ( w_11589 , \3675_b1 );
not ( w_11589 , w_11592 );
not (  , w_11593 );
and ( w_11592 , w_11593 , \3675_b0 );
buf ( \3677_b1 , \2708_b1 );
not ( \3677_b1 , w_11594 );
not ( \3677_b0 , w_11595 );
and ( w_11594 , w_11595 , \2708_b0 );
or ( \3678_b1 , \2674_b1 , w_11597 );
not ( w_11597 , w_11598 );
and ( \3678_b0 , \2674_b0 , w_11599 );
and ( w_11598 ,  , w_11599 );
buf ( w_11597 , \2697_b1 );
not ( w_11597 , w_11600 );
not (  , w_11601 );
and ( w_11600 , w_11601 , \2697_b0 );
buf ( \3679_b1 , \3678_b1 );
not ( \3679_b1 , w_11602 );
not ( \3679_b0 , w_11603 );
and ( w_11602 , w_11603 , \3678_b0 );
or ( \3680_b1 , \3677_b1 , w_11604 );
or ( \3680_b0 , \3677_b0 , \3679_b0 );
not ( \3679_b0 , w_11605 );
and ( w_11605 , w_11604 , \3679_b1 );
buf ( \3681_b1 , \2674_b1 );
not ( \3681_b1 , w_11606 );
not ( \3681_b0 , w_11607 );
and ( w_11606 , w_11607 , \2674_b0 );
or ( \3682_b1 , \3681_b1 , w_11609 );
not ( w_11609 , w_11610 );
and ( \3682_b0 , \3681_b0 , w_11611 );
and ( w_11610 ,  , w_11611 );
buf ( w_11609 , \2696_b1 );
not ( w_11609 , w_11612 );
not (  , w_11613 );
and ( w_11612 , w_11613 , \2696_b0 );
or ( \3683_b1 , \3680_b1 , w_11615 );
not ( w_11615 , w_11616 );
and ( \3683_b0 , \3680_b0 , w_11617 );
and ( w_11616 ,  , w_11617 );
buf ( w_11615 , \3682_b1 );
not ( w_11615 , w_11618 );
not (  , w_11619 );
and ( w_11618 , w_11619 , \3682_b0 );
buf ( \3684_b1 , \2693_b1 );
not ( \3684_b1 , w_11620 );
not ( \3684_b0 , w_11621 );
and ( w_11620 , w_11621 , \2693_b0 );
buf ( \3685_b1 , \1312_b1 );
not ( \3685_b1 , w_11622 );
not ( \3685_b0 , w_11623 );
and ( w_11622 , w_11623 , \1312_b0 );
or ( \3686_b1 , \3684_b1 , w_11624 );
or ( \3686_b0 , \3684_b0 , \3685_b0 );
not ( \3685_b0 , w_11625 );
and ( w_11625 , w_11624 , \3685_b1 );
or ( \3687_b1 , \d[5]_b1 , \a[11]_b1 );
xor ( \3687_b0 , \d[5]_b0 , w_11626 );
not ( w_11626 , w_11627 );
and ( w_11627 , \a[11]_b1 , \a[11]_b0 );
or ( \3688_b1 , \936_b1 , w_11629 );
not ( w_11629 , w_11630 );
and ( \3688_b0 , \936_b0 , w_11631 );
and ( w_11630 ,  , w_11631 );
buf ( w_11629 , \3687_b1 );
not ( w_11629 , w_11632 );
not (  , w_11633 );
and ( w_11632 , w_11633 , \3687_b0 );
or ( \3689_b1 , \3686_b1 , w_11635 );
not ( w_11635 , w_11636 );
and ( \3689_b0 , \3686_b0 , w_11637 );
and ( w_11636 ,  , w_11637 );
buf ( w_11635 , \3688_b1 );
not ( w_11635 , w_11638 );
not (  , w_11639 );
and ( w_11638 , w_11639 , \3688_b0 );
or ( \3690_b1 , \1366_b1 , \2671_b1 );
not ( \2671_b1 , w_11640 );
and ( \3690_b0 , \1366_b0 , w_11641 );
and ( w_11640 , w_11641 , \2671_b0 );
or ( \3691_b1 , \d[11]_b1 , \a[5]_b1 );
xor ( \3691_b0 , \d[11]_b0 , w_11642 );
not ( w_11642 , w_11643 );
and ( w_11643 , \a[5]_b1 , \a[5]_b0 );
or ( \3692_b1 , \947_b1 , \3691_b1 );
not ( \3691_b1 , w_11644 );
and ( \3692_b0 , \947_b0 , w_11645 );
and ( w_11644 , w_11645 , \3691_b0 );
or ( \3693_b1 , \3690_b1 , w_11647 );
not ( w_11647 , w_11648 );
and ( \3693_b0 , \3690_b0 , w_11649 );
and ( w_11648 ,  , w_11649 );
buf ( w_11647 , \3692_b1 );
not ( w_11647 , w_11650 );
not (  , w_11651 );
and ( w_11650 , w_11651 , \3692_b0 );
or ( \3694_b1 , \3689_b1 , \3693_b1 );
xor ( \3694_b0 , \3689_b0 , w_11652 );
not ( w_11652 , w_11653 );
and ( w_11653 , \3693_b1 , \3693_b0 );
buf ( \3695_b1 , \2664_b1 );
not ( \3695_b1 , w_11654 );
not ( \3695_b0 , w_11655 );
and ( w_11654 , w_11655 , \2664_b0 );
buf ( \3696_b1 , \2666_b1 );
not ( \3696_b1 , w_11656 );
not ( \3696_b0 , w_11657 );
and ( w_11656 , w_11657 , \2666_b0 );
buf ( \3697_b1 , \3696_b1 );
not ( \3697_b1 , w_11658 );
not ( \3697_b0 , w_11659 );
and ( w_11658 , w_11659 , \3696_b0 );
or ( \3698_b1 , \3695_b1 , w_11660 );
or ( \3698_b0 , \3695_b0 , \3697_b0 );
not ( \3697_b0 , w_11661 );
and ( w_11661 , w_11660 , \3697_b1 );
buf ( \3699_b1 , \2664_b1 );
not ( \3699_b1 , w_11662 );
not ( \3699_b0 , w_11663 );
and ( w_11662 , w_11663 , \2664_b0 );
buf ( \3700_b1 , \3699_b1 );
not ( \3700_b1 , w_11664 );
not ( \3700_b0 , w_11665 );
and ( w_11664 , w_11665 , \3699_b0 );
buf ( \3701_b1 , \2666_b1 );
not ( \3701_b1 , w_11666 );
not ( \3701_b0 , w_11667 );
and ( w_11666 , w_11667 , \2666_b0 );
or ( \3702_b1 , \3700_b1 , w_11668 );
or ( \3702_b0 , \3700_b0 , \3701_b0 );
not ( \3701_b0 , w_11669 );
and ( w_11669 , w_11668 , \3701_b1 );
or ( \3703_b1 , \3702_b1 , w_11671 );
not ( w_11671 , w_11672 );
and ( \3703_b0 , \3702_b0 , w_11673 );
and ( w_11672 ,  , w_11673 );
buf ( w_11671 , \2673_b1 );
not ( w_11671 , w_11674 );
not (  , w_11675 );
and ( w_11674 , w_11675 , \2673_b0 );
or ( \3704_b1 , \3698_b1 , w_11677 );
not ( w_11677 , w_11678 );
and ( \3704_b0 , \3698_b0 , w_11679 );
and ( w_11678 ,  , w_11679 );
buf ( w_11677 , \3703_b1 );
not ( w_11677 , w_11680 );
not (  , w_11681 );
and ( w_11680 , w_11681 , \3703_b0 );
or ( \3705_b1 , \3694_b1 , w_11682 );
xor ( \3705_b0 , \3694_b0 , w_11684 );
not ( w_11684 , w_11685 );
and ( w_11685 , w_11682 , w_11683 );
buf ( w_11682 , \3704_b1 );
not ( w_11682 , w_11686 );
not ( w_11683 , w_11687 );
and ( w_11686 , w_11687 , \3704_b0 );
or ( \3706_b1 , \2716_b1 , \2722_b1 );
xor ( \3706_b0 , \2716_b0 , w_11688 );
not ( w_11688 , w_11689 );
and ( w_11689 , \2722_b1 , \2722_b0 );
or ( \3707_b1 , \3706_b1 , \2729_b1 );
not ( \2729_b1 , w_11690 );
and ( \3707_b0 , \3706_b0 , w_11691 );
and ( w_11690 , w_11691 , \2729_b0 );
or ( \3708_b1 , \2716_b1 , \2722_b1 );
not ( \2722_b1 , w_11692 );
and ( \3708_b0 , \2716_b0 , w_11693 );
and ( w_11692 , w_11693 , \2722_b0 );
or ( \3709_b1 , \3707_b1 , w_11694 );
or ( \3709_b0 , \3707_b0 , \3708_b0 );
not ( \3708_b0 , w_11695 );
and ( w_11695 , w_11694 , \3708_b1 );
or ( \3710_b1 , \1583_b1 , \2662_b1 );
not ( \2662_b1 , w_11696 );
and ( \3710_b0 , \1583_b0 , w_11697 );
and ( w_11696 , w_11697 , \2662_b0 );
or ( \3711_b1 , \d[13]_b1 , \a[3]_b1 );
xor ( \3711_b0 , \d[13]_b0 , w_11698 );
not ( w_11698 , w_11699 );
and ( w_11699 , \a[3]_b1 , \a[3]_b0 );
or ( \3712_b1 , \1335_b1 , \3711_b1 );
not ( \3711_b1 , w_11700 );
and ( \3712_b0 , \1335_b0 , w_11701 );
and ( w_11700 , w_11701 , \3711_b0 );
or ( \3713_b1 , \3710_b1 , w_11703 );
not ( w_11703 , w_11704 );
and ( \3713_b0 , \3710_b0 , w_11705 );
and ( w_11704 ,  , w_11705 );
buf ( w_11703 , \3712_b1 );
not ( w_11703 , w_11706 );
not (  , w_11707 );
and ( w_11706 , w_11707 , \3712_b0 );
or ( \3714_b1 , \d[15]_b1 , \d[14]_b1 );
xor ( \3714_b0 , \d[15]_b0 , w_11708 );
not ( w_11708 , w_11709 );
and ( w_11709 , \d[14]_b1 , \d[14]_b0 );
or ( \3715_b1 , \a[0]_b1 , \d[15]_b1 );
xor ( \3715_b0 , \a[0]_b0 , w_11710 );
not ( w_11710 , w_11711 );
and ( w_11711 , \d[15]_b1 , \d[15]_b0 );
or ( \3716_b1 , \3714_b1 , w_11713 );
not ( w_11713 , w_11714 );
and ( \3716_b0 , \3714_b0 , w_11715 );
and ( w_11714 ,  , w_11715 );
buf ( w_11713 , \3715_b1 );
not ( w_11713 , w_11716 );
not (  , w_11717 );
and ( w_11716 , w_11717 , \3715_b0 );
or ( \3717_b1 , \3716_b1 , w_11718 );
or ( \3717_b0 , \3716_b0 , \2715_b0 );
not ( \2715_b0 , w_11719 );
and ( w_11719 , w_11718 , \2715_b1 );
or ( \3718_b1 , \a[1]_b1 , \d[15]_b1 );
xor ( \3718_b0 , \a[1]_b0 , w_11720 );
not ( w_11720 , w_11721 );
and ( w_11721 , \d[15]_b1 , \d[15]_b0 );
or ( \3719_b1 , \2715_b1 , w_11723 );
not ( w_11723 , w_11724 );
and ( \3719_b0 , \2715_b0 , w_11725 );
and ( w_11724 ,  , w_11725 );
buf ( w_11723 , \3718_b1 );
not ( w_11723 , w_11726 );
not (  , w_11727 );
and ( w_11726 , w_11727 , \3718_b0 );
or ( \3720_b1 , \3717_b1 , w_11729 );
not ( w_11729 , w_11730 );
and ( \3720_b0 , \3717_b0 , w_11731 );
and ( w_11730 ,  , w_11731 );
buf ( w_11729 , \3719_b1 );
not ( w_11729 , w_11732 );
not (  , w_11733 );
and ( w_11732 , w_11733 , \3719_b0 );
or ( \3721_b1 , \3713_b1 , \3720_b1 );
xor ( \3721_b0 , \3713_b0 , w_11734 );
not ( w_11734 , w_11735 );
and ( w_11735 , \3720_b1 , \3720_b0 );
buf ( \3722_b1 , \2686_b1 );
not ( \3722_b1 , w_11736 );
not ( \3722_b0 , w_11737 );
and ( w_11736 , w_11737 , \2686_b0 );
buf ( \3723_b1 , \999_b1 );
not ( \3723_b1 , w_11738 );
not ( \3723_b0 , w_11739 );
and ( w_11738 , w_11739 , \999_b0 );
or ( \3724_b1 , \3722_b1 , w_11740 );
or ( \3724_b0 , \3722_b0 , \3723_b0 );
not ( \3723_b0 , w_11741 );
and ( w_11741 , w_11740 , \3723_b1 );
buf ( \3725_b1 , \d[7]_b1 );
not ( \3725_b1 , w_11742 );
not ( \3725_b0 , w_11743 );
and ( w_11742 , w_11743 , \d[7]_b0 );
or ( \3726_b1 , \3725_b1 , w_11745 );
not ( w_11745 , w_11746 );
and ( \3726_b0 , \3725_b0 , w_11747 );
and ( w_11746 ,  , w_11747 );
buf ( w_11745 , \a[9]_b1 );
not ( w_11745 , w_11748 );
not (  , w_11749 );
and ( w_11748 , w_11749 , \a[9]_b0 );
buf ( \3727_b1 , \3726_b1 );
not ( \3727_b1 , w_11750 );
not ( \3727_b0 , w_11751 );
and ( w_11750 , w_11751 , \3726_b0 );
buf ( \3728_b1 , \a[9]_b1 );
not ( \3728_b1 , w_11752 );
not ( \3728_b0 , w_11753 );
and ( w_11752 , w_11753 , \a[9]_b0 );
or ( \3729_b1 , \3728_b1 , w_11755 );
not ( w_11755 , w_11756 );
and ( \3729_b0 , \3728_b0 , w_11757 );
and ( w_11756 ,  , w_11757 );
buf ( w_11755 , \d[7]_b1 );
not ( w_11755 , w_11758 );
not (  , w_11759 );
and ( w_11758 , w_11759 , \d[7]_b0 );
buf ( \3730_b1 , \3729_b1 );
not ( \3730_b1 , w_11760 );
not ( \3730_b0 , w_11761 );
and ( w_11760 , w_11761 , \3729_b0 );
or ( \3731_b1 , \3727_b1 , w_11762 );
or ( \3731_b0 , \3727_b0 , \3730_b0 );
not ( \3730_b0 , w_11763 );
and ( w_11763 , w_11762 , \3730_b1 );
or ( \3732_b1 , \3731_b1 , w_11765 );
not ( w_11765 , w_11766 );
and ( \3732_b0 , \3731_b0 , w_11767 );
and ( w_11766 ,  , w_11767 );
buf ( w_11765 , \1003_b1 );
not ( w_11765 , w_11768 );
not (  , w_11769 );
and ( w_11768 , w_11769 , \1003_b0 );
or ( \3733_b1 , \3724_b1 , w_11771 );
not ( w_11771 , w_11772 );
and ( \3733_b0 , \3724_b0 , w_11773 );
and ( w_11772 ,  , w_11773 );
buf ( w_11771 , \3732_b1 );
not ( w_11771 , w_11774 );
not (  , w_11775 );
and ( w_11774 , w_11775 , \3732_b0 );
or ( \3734_b1 , \3721_b1 , w_11776 );
xor ( \3734_b0 , \3721_b0 , w_11778 );
not ( w_11778 , w_11779 );
and ( w_11779 , w_11776 , w_11777 );
buf ( w_11776 , \3733_b1 );
not ( w_11776 , w_11780 );
not ( w_11777 , w_11781 );
and ( w_11780 , w_11781 , \3733_b0 );
buf ( \3735_b1 , \3734_b1 );
not ( \3735_b1 , w_11782 );
not ( \3735_b0 , w_11783 );
and ( w_11782 , w_11783 , \3734_b0 );
or ( \3736_b1 , \3709_b1 , \3735_b1 );
xor ( \3736_b0 , \3709_b0 , w_11784 );
not ( w_11784 , w_11785 );
and ( w_11785 , \3735_b1 , \3735_b0 );
or ( \3737_b1 , \3705_b1 , \3736_b1 );
xor ( \3737_b0 , \3705_b0 , w_11786 );
not ( w_11786 , w_11787 );
and ( w_11787 , \3736_b1 , \3736_b0 );
or ( \3738_b1 , \3683_b1 , \3737_b1 );
xor ( \3738_b0 , \3683_b0 , w_11788 );
not ( w_11788 , w_11789 );
and ( w_11789 , \3737_b1 , \3737_b0 );
buf ( \3739_b1 , \2680_b1 );
not ( \3739_b1 , w_11790 );
not ( \3739_b0 , w_11791 );
and ( w_11790 , w_11791 , \2680_b0 );
buf ( \3740_b1 , \1026_b1 );
not ( \3740_b1 , w_11792 );
not ( \3740_b0 , w_11793 );
and ( w_11792 , w_11793 , \1026_b0 );
or ( \3741_b1 , \3739_b1 , w_11794 );
or ( \3741_b0 , \3739_b0 , \3740_b0 );
not ( \3740_b0 , w_11795 );
and ( w_11795 , w_11794 , \3740_b1 );
or ( \3742_b1 , \d[9]_b1 , \a[7]_b1 );
xor ( \3742_b0 , \d[9]_b0 , w_11796 );
not ( w_11796 , w_11797 );
and ( w_11797 , \a[7]_b1 , \a[7]_b0 );
or ( \3743_b1 , \1058_b1 , w_11799 );
not ( w_11799 , w_11800 );
and ( \3743_b0 , \1058_b0 , w_11801 );
and ( w_11800 ,  , w_11801 );
buf ( w_11799 , \3742_b1 );
not ( w_11799 , w_11802 );
not (  , w_11803 );
and ( w_11802 , w_11803 , \3742_b0 );
or ( \3744_b1 , \3741_b1 , w_11805 );
not ( w_11805 , w_11806 );
and ( \3744_b0 , \3741_b0 , w_11807 );
and ( w_11806 ,  , w_11807 );
buf ( w_11805 , \3743_b1 );
not ( w_11805 , w_11808 );
not (  , w_11809 );
and ( w_11808 , w_11809 , \3743_b0 );
buf ( \3745_b1 , \2727_b1 );
not ( \3745_b1 , w_11810 );
not ( \3745_b0 , w_11811 );
and ( w_11810 , w_11811 , \2727_b0 );
buf ( \3746_b1 , \962_b1 );
not ( \3746_b1 , w_11812 );
not ( \3746_b0 , w_11813 );
and ( w_11812 , w_11813 , \962_b0 );
or ( \3747_b1 , \3745_b1 , w_11814 );
or ( \3747_b0 , \3745_b0 , \3746_b0 );
not ( \3746_b0 , w_11815 );
and ( w_11815 , w_11814 , \3746_b1 );
or ( \3748_b1 , \d[3]_b1 , \a[13]_b1 );
xor ( \3748_b0 , \d[3]_b0 , w_11816 );
not ( w_11816 , w_11817 );
and ( w_11817 , \a[13]_b1 , \a[13]_b0 );
or ( \3749_b1 , \965_b1 , w_11819 );
not ( w_11819 , w_11820 );
and ( \3749_b0 , \965_b0 , w_11821 );
and ( w_11820 ,  , w_11821 );
buf ( w_11819 , \3748_b1 );
not ( w_11819 , w_11822 );
not (  , w_11823 );
and ( w_11822 , w_11823 , \3748_b0 );
or ( \3750_b1 , \3747_b1 , w_11825 );
not ( w_11825 , w_11826 );
and ( \3750_b0 , \3747_b0 , w_11827 );
and ( w_11826 ,  , w_11827 );
buf ( w_11825 , \3749_b1 );
not ( w_11825 , w_11828 );
not (  , w_11829 );
and ( w_11828 , w_11829 , \3749_b0 );
or ( \3751_b1 , \3744_b1 , \3750_b1 );
xor ( \3751_b0 , \3744_b0 , w_11830 );
not ( w_11830 , w_11831 );
and ( w_11831 , \3750_b1 , \3750_b0 );
or ( \3752_b1 , \1065_b1 , \2720_b1 );
not ( \2720_b1 , w_11832 );
and ( \3752_b0 , \1065_b0 , w_11833 );
and ( w_11832 , w_11833 , \2720_b0 );
buf ( \3753_b1 , \d[0]_b1 );
not ( \3753_b1 , w_11834 );
not ( \3753_b0 , w_11835 );
and ( w_11834 , w_11835 , \d[0]_b0 );
or ( \3754_b1 , \d[1]_b1 , w_11836 );
xor ( \3754_b0 , \d[1]_b0 , w_11838 );
not ( w_11838 , w_11839 );
and ( w_11839 , w_11836 , w_11837 );
buf ( w_11836 , \a[15]_b1 );
not ( w_11836 , w_11840 );
not ( w_11837 , w_11841 );
and ( w_11840 , w_11841 , \a[15]_b0 );
or ( \3755_b1 , \3753_b1 , w_11843 );
not ( w_11843 , w_11844 );
and ( \3755_b0 , \3753_b0 , w_11845 );
and ( w_11844 ,  , w_11845 );
buf ( w_11843 , \3754_b1 );
not ( w_11843 , w_11846 );
not (  , w_11847 );
and ( w_11846 , w_11847 , \3754_b0 );
or ( \3756_b1 , \3752_b1 , w_11849 );
not ( w_11849 , w_11850 );
and ( \3756_b0 , \3752_b0 , w_11851 );
and ( w_11850 ,  , w_11851 );
buf ( w_11849 , \3755_b1 );
not ( w_11849 , w_11852 );
not (  , w_11853 );
and ( w_11852 , w_11853 , \3755_b0 );
buf ( \3757_b1 , \3756_b1 );
not ( \3757_b1 , w_11854 );
not ( \3757_b0 , w_11855 );
and ( w_11854 , w_11855 , \3756_b0 );
or ( \3758_b1 , \a[0]_b1 , w_11856 );
or ( \3758_b0 , \a[0]_b0 , \d[14]_b0 );
not ( \d[14]_b0 , w_11857 );
and ( w_11857 , w_11856 , \d[14]_b1 );
or ( \3759_b1 , \3758_b1 , w_11859 );
not ( w_11859 , w_11860 );
and ( \3759_b0 , \3758_b0 , w_11861 );
and ( w_11860 ,  , w_11861 );
buf ( w_11859 , \d[13]_b1 );
not ( w_11859 , w_11862 );
not (  , w_11863 );
and ( w_11862 , w_11863 , \d[13]_b0 );
or ( \3760_b1 , \a[0]_b1 , w_11865 );
not ( w_11865 , w_11866 );
and ( \3760_b0 , \a[0]_b0 , w_11867 );
and ( w_11866 ,  , w_11867 );
buf ( w_11865 , \d[14]_b1 );
not ( w_11865 , w_11868 );
not (  , w_11869 );
and ( w_11868 , w_11869 , \d[14]_b0 );
buf ( \3762_b1 , \3761_b1 );
not ( \3762_b1 , w_11870 );
not ( \3762_b0 , w_11871 );
and ( w_11870 , w_11871 , \3761_b0 );
or ( \3763_b1 , \3757_b1 , \3762_b1 );
not ( \3762_b1 , w_11872 );
and ( \3763_b0 , \3757_b0 , w_11873 );
and ( w_11872 , w_11873 , \3762_b0 );
or ( \3764_b1 , \3756_b1 , \3761_b1 );
not ( \3761_b1 , w_11874 );
and ( \3764_b0 , \3756_b0 , w_11875 );
and ( w_11874 , w_11875 , \3761_b0 );
or ( \3765_b1 , \3763_b1 , w_11877 );
not ( w_11877 , w_11878 );
and ( \3765_b0 , \3763_b0 , w_11879 );
and ( w_11878 ,  , w_11879 );
buf ( w_11877 , \3764_b1 );
not ( w_11877 , w_11880 );
not (  , w_11881 );
and ( w_11880 , w_11881 , \3764_b0 );
or ( \3766_b1 , \3751_b1 , w_11882 );
xor ( \3766_b0 , \3751_b0 , w_11884 );
not ( w_11884 , w_11885 );
and ( w_11885 , w_11882 , w_11883 );
buf ( w_11882 , \3765_b1 );
not ( w_11882 , w_11886 );
not ( w_11883 , w_11887 );
and ( w_11886 , w_11887 , \3765_b0 );
or ( \3767_b1 , \2682_b1 , \2688_b1 );
xor ( \3767_b0 , \2682_b0 , w_11888 );
not ( w_11888 , w_11889 );
and ( w_11889 , \2688_b1 , \2688_b0 );
or ( \3768_b1 , \3767_b1 , \2695_b1 );
not ( \2695_b1 , w_11890 );
and ( \3768_b0 , \3767_b0 , w_11891 );
and ( w_11890 , w_11891 , \2695_b0 );
or ( \3769_b1 , \2682_b1 , \2688_b1 );
not ( \2688_b1 , w_11892 );
and ( \3769_b0 , \2682_b0 , w_11893 );
and ( w_11892 , w_11893 , \2688_b0 );
or ( \3770_b1 , \3768_b1 , w_11894 );
or ( \3770_b0 , \3768_b0 , \3769_b0 );
not ( \3769_b0 , w_11895 );
and ( w_11895 , w_11894 , \3769_b1 );
or ( \3771_b1 , \3766_b1 , w_11896 );
xor ( \3771_b0 , \3766_b0 , w_11898 );
not ( w_11898 , w_11899 );
and ( w_11899 , w_11896 , w_11897 );
buf ( w_11896 , \3770_b1 );
not ( w_11896 , w_11900 );
not ( w_11897 , w_11901 );
and ( w_11900 , w_11901 , \3770_b0 );
buf ( \3772_b1 , \3771_b1 );
not ( \3772_b1 , w_11902 );
not ( \3772_b0 , w_11903 );
and ( w_11902 , w_11903 , \3771_b0 );
or ( \3773_b1 , \2714_b1 , \2730_b1 );
xor ( \3773_b0 , \2714_b0 , w_11904 );
not ( w_11904 , w_11905 );
and ( w_11905 , \2730_b1 , \2730_b0 );
or ( \3774_b1 , \3773_b1 , \2736_b1 );
not ( \2736_b1 , w_11906 );
and ( \3774_b0 , \3773_b0 , w_11907 );
and ( w_11906 , w_11907 , \2736_b0 );
or ( \3775_b1 , \2714_b1 , \2730_b1 );
not ( \2730_b1 , w_11908 );
and ( \3775_b0 , \2714_b0 , w_11909 );
and ( w_11908 , w_11909 , \2730_b0 );
or ( \3776_b1 , \3774_b1 , w_11910 );
or ( \3776_b0 , \3774_b0 , \3775_b0 );
not ( \3775_b0 , w_11911 );
and ( w_11911 , w_11910 , \3775_b1 );
buf ( \3777_b1 , \3776_b1 );
not ( \3777_b1 , w_11912 );
not ( \3777_b0 , w_11913 );
and ( w_11912 , w_11913 , \3776_b0 );
or ( \3778_b1 , \3772_b1 , \3777_b1 );
not ( \3777_b1 , w_11914 );
and ( \3778_b0 , \3772_b0 , w_11915 );
and ( w_11914 , w_11915 , \3777_b0 );
or ( \3779_b1 , \3776_b1 , \3771_b1 );
not ( \3771_b1 , w_11916 );
and ( \3779_b0 , \3776_b0 , w_11917 );
and ( w_11916 , w_11917 , \3771_b0 );
or ( \3780_b1 , \3778_b1 , w_11919 );
not ( w_11919 , w_11920 );
and ( \3780_b0 , \3778_b0 , w_11921 );
and ( w_11920 ,  , w_11921 );
buf ( w_11919 , \3779_b1 );
not ( w_11919 , w_11922 );
not (  , w_11923 );
and ( w_11922 , w_11923 , \3779_b0 );
or ( \3781_b1 , \3738_b1 , w_11924 );
xor ( \3781_b0 , \3738_b0 , w_11926 );
not ( w_11926 , w_11927 );
and ( w_11927 , w_11924 , w_11925 );
buf ( w_11924 , \3780_b1 );
not ( w_11924 , w_11928 );
not ( w_11925 , w_11929 );
and ( w_11928 , w_11929 , \3780_b0 );
or ( \3782_b1 , \3676_b1 , w_11930 );
xor ( \3782_b0 , \3676_b0 , w_11932 );
not ( w_11932 , w_11933 );
and ( w_11933 , w_11930 , w_11931 );
buf ( w_11930 , \3781_b1 );
not ( w_11930 , w_11934 );
not ( w_11931 , w_11935 );
and ( w_11934 , w_11935 , \3781_b0 );
buf ( \3783_b1 , \3782_b1 );
not ( \3783_b1 , w_11936 );
not ( \3783_b0 , w_11937 );
and ( w_11936 , w_11937 , \3782_b0 );
or ( \3784_b1 , \3668_b1 , \3783_b1 );
not ( \3783_b1 , w_11938 );
and ( \3784_b0 , \3668_b0 , w_11939 );
and ( w_11938 , w_11939 , \3783_b0 );
buf ( \3785_b1 , \3668_b1 );
not ( \3785_b1 , w_11940 );
not ( \3785_b0 , w_11941 );
and ( w_11940 , w_11941 , \3668_b0 );
or ( \3786_b1 , \3785_b1 , \3782_b1 );
not ( \3782_b1 , w_11942 );
and ( \3786_b0 , \3785_b0 , w_11943 );
and ( w_11942 , w_11943 , \3782_b0 );
or ( \3787_b1 , \3784_b1 , w_11945 );
not ( w_11945 , w_11946 );
and ( \3787_b0 , \3784_b0 , w_11947 );
and ( w_11946 ,  , w_11947 );
buf ( w_11945 , \3786_b1 );
not ( w_11945 , w_11948 );
not (  , w_11949 );
and ( w_11948 , w_11949 , \3786_b0 );
or ( \3788_b1 , \3787_b1 , w_11951 );
not ( w_11951 , w_11952 );
and ( \3788_b0 , \3787_b0 , w_11953 );
and ( w_11952 ,  , w_11953 );
buf ( w_11951 , \1668_b1 );
not ( w_11951 , w_11954 );
not (  , w_11955 );
and ( w_11954 , w_11955 , \1668_b0 );
buf ( \3789_b1 , \2581_b1 );
not ( \3789_b1 , w_11956 );
not ( \3789_b0 , w_11957 );
and ( w_11956 , w_11957 , \2581_b0 );
or ( \3790_b1 , \2403_b1 , w_11959 );
not ( w_11959 , w_11960 );
and ( \3790_b0 , \2403_b0 , w_11961 );
and ( w_11960 ,  , w_11961 );
buf ( w_11959 , \2284_b1 );
not ( w_11959 , w_11962 );
not (  , w_11963 );
and ( w_11962 , w_11963 , \2284_b0 );
or ( \3791_b1 , \3789_b1 , w_11965 );
not ( w_11965 , w_11966 );
and ( \3791_b0 , \3789_b0 , w_11967 );
and ( w_11966 ,  , w_11967 );
buf ( w_11965 , \3790_b1 );
not ( w_11965 , w_11968 );
not (  , w_11969 );
and ( w_11968 , w_11969 , \3790_b0 );
or ( \3792_b1 , \2282_b1 , \2587_b1 );
not ( \2587_b1 , w_11970 );
and ( \3792_b0 , \2282_b0 , w_11971 );
and ( w_11970 , w_11971 , \2587_b0 );
or ( \3793_b1 , \2129_b1 , w_11973 );
not ( w_11973 , w_11974 );
and ( \3793_b0 , \2129_b0 , w_11975 );
and ( w_11974 ,  , w_11975 );
buf ( w_11973 , \2285_b1 );
not ( w_11973 , w_11976 );
not (  , w_11977 );
and ( w_11976 , w_11977 , \2285_b0 );
or ( \3794_b1 , \3792_b1 , w_11978 );
or ( \3794_b0 , \3792_b0 , \3793_b0 );
not ( \3793_b0 , w_11979 );
and ( w_11979 , w_11978 , \3793_b1 );
or ( \3795_b1 , \2129_b1 , w_11981 );
not ( w_11981 , w_11982 );
and ( \3795_b0 , \2129_b0 , w_11983 );
and ( w_11982 ,  , w_11983 );
buf ( w_11981 , \2273_b1 );
not ( w_11981 , w_11984 );
not (  , w_11985 );
and ( w_11984 , w_11985 , \2273_b0 );
or ( \3796_b1 , \3794_b1 , w_11987 );
not ( w_11987 , w_11988 );
and ( \3796_b0 , \3794_b0 , w_11989 );
and ( w_11988 ,  , w_11989 );
buf ( w_11987 , \3795_b1 );
not ( w_11987 , w_11990 );
not (  , w_11991 );
and ( w_11990 , w_11991 , \3795_b0 );
or ( \3797_b1 , \3791_b1 , \3796_b1 );
not ( \3796_b1 , w_11992 );
and ( \3797_b0 , \3791_b0 , w_11993 );
and ( w_11992 , w_11993 , \3796_b0 );
buf ( \3798_b1 , \2596_b1 );
not ( \3798_b1 , w_11994 );
not ( \3798_b0 , w_11995 );
and ( w_11994 , w_11995 , \2596_b0 );
buf ( \3799_b1 , \2581_b1 );
not ( \3799_b1 , w_11996 );
not ( \3799_b0 , w_11997 );
and ( w_11996 , w_11997 , \2581_b0 );
or ( \3800_b1 , \3798_b1 , w_11998 );
or ( \3800_b0 , \3798_b0 , \3799_b0 );
not ( \3799_b0 , w_11999 );
and ( w_11999 , w_11998 , \3799_b1 );
or ( \3801_b1 , \3800_b1 , w_12001 );
not ( w_12001 , w_12002 );
and ( \3801_b0 , \3800_b0 , w_12003 );
and ( w_12002 ,  , w_12003 );
buf ( w_12001 , \2579_b1 );
not ( w_12001 , w_12004 );
not (  , w_12005 );
and ( w_12004 , w_12005 , \2579_b0 );
or ( \3802_b1 , \3797_b1 , w_12007 );
not ( w_12007 , w_12008 );
and ( \3802_b0 , \3797_b0 , w_12009 );
and ( w_12008 ,  , w_12009 );
buf ( w_12007 , \3801_b1 );
not ( w_12007 , w_12010 );
not (  , w_12011 );
and ( w_12010 , w_12011 , \3801_b0 );
buf ( \3803_b1 , \2555_b1 );
not ( \3803_b1 , w_12012 );
not ( \3803_b0 , w_12013 );
and ( w_12012 , w_12013 , \2555_b0 );
buf ( \3804_b1 , \3803_b1 );
not ( \3804_b1 , w_12014 );
not ( \3804_b0 , w_12015 );
and ( w_12014 , w_12015 , \3803_b0 );
buf ( \3805_b1 , \2528_b1 );
not ( \3805_b1 , w_12016 );
not ( \3805_b0 , w_12017 );
and ( w_12016 , w_12017 , \2528_b0 );
or ( \3806_b1 , \3804_b1 , w_12018 );
or ( \3806_b0 , \3804_b0 , \3805_b0 );
not ( \3805_b0 , w_12019 );
and ( w_12019 , w_12018 , \3805_b1 );
or ( \3807_b1 , \3806_b1 , w_12021 );
not ( w_12021 , w_12022 );
and ( \3807_b0 , \3806_b0 , w_12023 );
and ( w_12022 ,  , w_12023 );
buf ( w_12021 , \2566_b1 );
not ( w_12021 , w_12024 );
not (  , w_12025 );
and ( w_12024 , w_12025 , \2566_b0 );
buf ( \3808_b1 , \2528_b1 );
not ( \3808_b1 , w_12026 );
not ( \3808_b0 , w_12027 );
and ( w_12026 , w_12027 , \2528_b0 );
or ( \3809_b1 , \3808_b1 , w_12029 );
not ( w_12029 , w_12030 );
and ( \3809_b0 , \3808_b0 , w_12031 );
and ( w_12030 ,  , w_12031 );
buf ( w_12029 , \2555_b1 );
not ( w_12029 , w_12032 );
not (  , w_12033 );
and ( w_12032 , w_12033 , \2555_b0 );
or ( \3810_b1 , \3807_b1 , w_12035 );
not ( w_12035 , w_12036 );
and ( \3810_b0 , \3807_b0 , w_12037 );
and ( w_12036 ,  , w_12037 );
buf ( w_12035 , \3809_b1 );
not ( w_12035 , w_12038 );
not (  , w_12039 );
and ( w_12038 , w_12039 , \3809_b0 );
buf ( \3811_b1 , \2497_b1 );
not ( \3811_b1 , w_12040 );
not ( \3811_b0 , w_12041 );
and ( w_12040 , w_12041 , \2497_b0 );
buf ( \3812_b1 , \1770_b1 );
not ( \3812_b1 , w_12042 );
not ( \3812_b0 , w_12043 );
and ( w_12042 , w_12043 , \1770_b0 );
or ( \3813_b1 , \3811_b1 , w_12044 );
or ( \3813_b0 , \3811_b0 , \3812_b0 );
not ( \3812_b0 , w_12045 );
and ( w_12045 , w_12044 , \3812_b1 );
or ( \3814_b1 , \c[9]_b1 , \b[7]_b1 );
xor ( \3814_b0 , \c[9]_b0 , w_12046 );
not ( w_12046 , w_12047 );
and ( w_12047 , \b[7]_b1 , \b[7]_b0 );
or ( \3815_b1 , \1802_b1 , w_12049 );
not ( w_12049 , w_12050 );
and ( \3815_b0 , \1802_b0 , w_12051 );
and ( w_12050 ,  , w_12051 );
buf ( w_12049 , \3814_b1 );
not ( w_12049 , w_12052 );
not (  , w_12053 );
and ( w_12052 , w_12053 , \3814_b0 );
or ( \3816_b1 , \3813_b1 , w_12055 );
not ( w_12055 , w_12056 );
and ( \3816_b0 , \3813_b0 , w_12057 );
and ( w_12056 ,  , w_12057 );
buf ( w_12055 , \3815_b1 );
not ( w_12055 , w_12058 );
not (  , w_12059 );
and ( w_12058 , w_12059 , \3815_b0 );
buf ( \3817_b1 , \2546_b1 );
not ( \3817_b1 , w_12060 );
not ( \3817_b0 , w_12061 );
and ( w_12060 , w_12061 , \2546_b0 );
buf ( \3818_b1 , \2370_b1 );
not ( \3818_b1 , w_12062 );
not ( \3818_b0 , w_12063 );
and ( w_12062 , w_12063 , \2370_b0 );
or ( \3819_b1 , \3817_b1 , w_12064 );
or ( \3819_b0 , \3817_b0 , \3818_b0 );
not ( \3818_b0 , w_12065 );
and ( w_12065 , w_12064 , \3818_b1 );
or ( \3820_b1 , \c[3]_b1 , \b[13]_b1 );
xor ( \3820_b0 , \c[3]_b0 , w_12066 );
not ( w_12066 , w_12067 );
and ( w_12067 , \b[13]_b1 , \b[13]_b0 );
or ( \3821_b1 , \1708_b1 , w_12069 );
not ( w_12069 , w_12070 );
and ( \3821_b0 , \1708_b0 , w_12071 );
and ( w_12070 ,  , w_12071 );
buf ( w_12069 , \3820_b1 );
not ( w_12069 , w_12072 );
not (  , w_12073 );
and ( w_12072 , w_12073 , \3820_b0 );
or ( \3822_b1 , \3819_b1 , w_12075 );
not ( w_12075 , w_12076 );
and ( \3822_b0 , \3819_b0 , w_12077 );
and ( w_12076 ,  , w_12077 );
buf ( w_12075 , \3821_b1 );
not ( w_12075 , w_12078 );
not (  , w_12079 );
and ( w_12078 , w_12079 , \3821_b0 );
or ( \3823_b1 , \3816_b1 , \3822_b1 );
xor ( \3823_b0 , \3816_b0 , w_12080 );
not ( w_12080 , w_12081 );
and ( w_12081 , \3822_b1 , \3822_b0 );
or ( \3824_b1 , \1756_b1 , \2539_b1 );
not ( \2539_b1 , w_12082 );
and ( \3824_b0 , \1756_b0 , w_12083 );
and ( w_12082 , w_12083 , \2539_b0 );
buf ( \3825_b1 , \c[0]_b1 );
not ( \3825_b1 , w_12084 );
not ( \3825_b0 , w_12085 );
and ( w_12084 , w_12085 , \c[0]_b0 );
or ( \3826_b1 , \c[1]_b1 , w_12086 );
xor ( \3826_b0 , \c[1]_b0 , w_12088 );
not ( w_12088 , w_12089 );
and ( w_12089 , w_12086 , w_12087 );
buf ( w_12086 , \b[15]_b1 );
not ( w_12086 , w_12090 );
not ( w_12087 , w_12091 );
and ( w_12090 , w_12091 , \b[15]_b0 );
or ( \3827_b1 , \3825_b1 , w_12093 );
not ( w_12093 , w_12094 );
and ( \3827_b0 , \3825_b0 , w_12095 );
and ( w_12094 ,  , w_12095 );
buf ( w_12093 , \3826_b1 );
not ( w_12093 , w_12096 );
not (  , w_12097 );
and ( w_12096 , w_12097 , \3826_b0 );
or ( \3828_b1 , \3824_b1 , w_12099 );
not ( w_12099 , w_12100 );
and ( \3828_b0 , \3824_b0 , w_12101 );
and ( w_12100 ,  , w_12101 );
buf ( w_12099 , \3827_b1 );
not ( w_12099 , w_12102 );
not (  , w_12103 );
and ( w_12102 , w_12103 , \3827_b0 );
buf ( \3829_b1 , \3828_b1 );
not ( \3829_b1 , w_12104 );
not ( \3829_b0 , w_12105 );
and ( w_12104 , w_12105 , \3828_b0 );
or ( \3830_b1 , \b[0]_b1 , w_12106 );
or ( \3830_b0 , \b[0]_b0 , \c[14]_b0 );
not ( \c[14]_b0 , w_12107 );
and ( w_12107 , w_12106 , \c[14]_b1 );
or ( \3831_b1 , \3830_b1 , w_12109 );
not ( w_12109 , w_12110 );
and ( \3831_b0 , \3830_b0 , w_12111 );
and ( w_12110 ,  , w_12111 );
buf ( w_12109 , \c[13]_b1 );
not ( w_12109 , w_12112 );
not (  , w_12113 );
and ( w_12112 , w_12113 , \c[13]_b0 );
or ( \3832_b1 , \b[0]_b1 , w_12115 );
not ( w_12115 , w_12116 );
and ( \3832_b0 , \b[0]_b0 , w_12117 );
and ( w_12116 ,  , w_12117 );
buf ( w_12115 , \c[14]_b1 );
not ( w_12115 , w_12118 );
not (  , w_12119 );
and ( w_12118 , w_12119 , \c[14]_b0 );
buf ( \3834_b1 , \3833_b1 );
not ( \3834_b1 , w_12120 );
not ( \3834_b0 , w_12121 );
and ( w_12120 , w_12121 , \3833_b0 );
or ( \3835_b1 , \3829_b1 , \3834_b1 );
not ( \3834_b1 , w_12122 );
and ( \3835_b0 , \3829_b0 , w_12123 );
and ( w_12122 , w_12123 , \3834_b0 );
or ( \3836_b1 , \3828_b1 , \3833_b1 );
not ( \3833_b1 , w_12124 );
and ( \3836_b0 , \3828_b0 , w_12125 );
and ( w_12124 , w_12125 , \3833_b0 );
or ( \3837_b1 , \3835_b1 , w_12127 );
not ( w_12127 , w_12128 );
and ( \3837_b0 , \3835_b0 , w_12129 );
and ( w_12128 ,  , w_12129 );
buf ( w_12127 , \3836_b1 );
not ( w_12127 , w_12130 );
not (  , w_12131 );
and ( w_12130 , w_12131 , \3836_b0 );
or ( \3838_b1 , \3823_b1 , w_12132 );
xor ( \3838_b0 , \3823_b0 , w_12134 );
not ( w_12134 , w_12135 );
and ( w_12135 , w_12132 , w_12133 );
buf ( w_12132 , \3837_b1 );
not ( w_12132 , w_12136 );
not ( w_12133 , w_12137 );
and ( w_12136 , w_12137 , \3837_b0 );
or ( \3839_b1 , \2501_b1 , \2507_b1 );
xor ( \3839_b0 , \2501_b0 , w_12138 );
not ( w_12138 , w_12139 );
and ( w_12139 , \2507_b1 , \2507_b0 );
or ( \3840_b1 , \3839_b1 , \2514_b1 );
not ( \2514_b1 , w_12140 );
and ( \3840_b0 , \3839_b0 , w_12141 );
and ( w_12140 , w_12141 , \2514_b0 );
or ( \3841_b1 , \2501_b1 , \2507_b1 );
not ( \2507_b1 , w_12142 );
and ( \3841_b0 , \2501_b0 , w_12143 );
and ( w_12142 , w_12143 , \2507_b0 );
or ( \3842_b1 , \3840_b1 , w_12144 );
or ( \3842_b0 , \3840_b0 , \3841_b0 );
not ( \3841_b0 , w_12145 );
and ( w_12145 , w_12144 , \3841_b1 );
or ( \3843_b1 , \3838_b1 , w_12146 );
xor ( \3843_b0 , \3838_b0 , w_12148 );
not ( w_12148 , w_12149 );
and ( w_12149 , w_12146 , w_12147 );
buf ( w_12146 , \3842_b1 );
not ( w_12146 , w_12150 );
not ( w_12147 , w_12151 );
and ( w_12150 , w_12151 , \3842_b0 );
buf ( \3844_b1 , \3843_b1 );
not ( \3844_b1 , w_12152 );
not ( \3844_b0 , w_12153 );
and ( w_12152 , w_12153 , \3843_b0 );
or ( \3845_b1 , \2533_b1 , \2549_b1 );
xor ( \3845_b0 , \2533_b0 , w_12154 );
not ( w_12154 , w_12155 );
and ( w_12155 , \2549_b1 , \2549_b0 );
or ( \3846_b1 , \3845_b1 , \2554_b1 );
not ( \2554_b1 , w_12156 );
and ( \3846_b0 , \3845_b0 , w_12157 );
and ( w_12156 , w_12157 , \2554_b0 );
or ( \3847_b1 , \2533_b1 , \2549_b1 );
not ( \2549_b1 , w_12158 );
and ( \3847_b0 , \2533_b0 , w_12159 );
and ( w_12158 , w_12159 , \2549_b0 );
or ( \3848_b1 , \3846_b1 , w_12160 );
or ( \3848_b0 , \3846_b0 , \3847_b0 );
not ( \3847_b0 , w_12161 );
and ( w_12161 , w_12160 , \3847_b1 );
buf ( \3849_b1 , \3848_b1 );
not ( \3849_b1 , w_12162 );
not ( \3849_b0 , w_12163 );
and ( w_12162 , w_12163 , \3848_b0 );
or ( \3850_b1 , \3844_b1 , \3849_b1 );
not ( \3849_b1 , w_12164 );
and ( \3850_b0 , \3844_b0 , w_12165 );
and ( w_12164 , w_12165 , \3849_b0 );
or ( \3851_b1 , \3848_b1 , \3843_b1 );
not ( \3843_b1 , w_12166 );
and ( \3851_b0 , \3848_b0 , w_12167 );
and ( w_12166 , w_12167 , \3843_b0 );
or ( \3852_b1 , \3850_b1 , w_12169 );
not ( w_12169 , w_12170 );
and ( \3852_b0 , \3850_b0 , w_12171 );
and ( w_12170 ,  , w_12171 );
buf ( w_12169 , \3851_b1 );
not ( w_12169 , w_12172 );
not (  , w_12173 );
and ( w_12172 , w_12173 , \3851_b0 );
or ( \3853_b1 , \2493_b1 , w_12175 );
not ( w_12175 , w_12176 );
and ( \3853_b0 , \2493_b0 , w_12177 );
and ( w_12176 ,  , w_12177 );
buf ( w_12175 , \2516_b1 );
not ( w_12175 , w_12178 );
not (  , w_12179 );
and ( w_12178 , w_12179 , \2516_b0 );
buf ( \3854_b1 , \3853_b1 );
not ( \3854_b1 , w_12180 );
not ( \3854_b0 , w_12181 );
and ( w_12180 , w_12181 , \3853_b0 );
buf ( \3855_b1 , \2527_b1 );
not ( \3855_b1 , w_12182 );
not ( \3855_b0 , w_12183 );
and ( w_12182 , w_12183 , \2527_b0 );
or ( \3856_b1 , \3854_b1 , w_12184 );
or ( \3856_b0 , \3854_b0 , \3855_b0 );
not ( \3855_b0 , w_12185 );
and ( w_12185 , w_12184 , \3855_b1 );
buf ( \3857_b1 , \2493_b1 );
not ( \3857_b1 , w_12186 );
not ( \3857_b0 , w_12187 );
and ( w_12186 , w_12187 , \2493_b0 );
or ( \3858_b1 , \3857_b1 , w_12189 );
not ( w_12189 , w_12190 );
and ( \3858_b0 , \3857_b0 , w_12191 );
and ( w_12190 ,  , w_12191 );
buf ( w_12189 , \2515_b1 );
not ( w_12189 , w_12192 );
not (  , w_12193 );
and ( w_12192 , w_12193 , \2515_b0 );
or ( \3859_b1 , \3856_b1 , w_12195 );
not ( w_12195 , w_12196 );
and ( \3859_b0 , \3856_b0 , w_12197 );
and ( w_12196 ,  , w_12197 );
buf ( w_12195 , \3858_b1 );
not ( w_12195 , w_12198 );
not (  , w_12199 );
and ( w_12198 , w_12199 , \3858_b0 );
buf ( \3860_b1 , \2512_b1 );
not ( \3860_b1 , w_12200 );
not ( \3860_b0 , w_12201 );
and ( w_12200 , w_12201 , \2512_b0 );
buf ( \3861_b1 , \2052_b1 );
not ( \3861_b1 , w_12202 );
not ( \3861_b0 , w_12203 );
and ( w_12202 , w_12203 , \2052_b0 );
or ( \3862_b1 , \3860_b1 , w_12204 );
or ( \3862_b0 , \3860_b0 , \3861_b0 );
not ( \3861_b0 , w_12205 );
and ( w_12205 , w_12204 , \3861_b1 );
or ( \3863_b1 , \c[5]_b1 , \b[11]_b1 );
xor ( \3863_b0 , \c[5]_b0 , w_12206 );
not ( w_12206 , w_12207 );
and ( w_12207 , \b[11]_b1 , \b[11]_b0 );
or ( \3864_b1 , \1678_b1 , w_12209 );
not ( w_12209 , w_12210 );
and ( \3864_b0 , \1678_b0 , w_12211 );
and ( w_12210 ,  , w_12211 );
buf ( w_12209 , \3863_b1 );
not ( w_12209 , w_12212 );
not (  , w_12213 );
and ( w_12212 , w_12213 , \3863_b0 );
or ( \3865_b1 , \3862_b1 , w_12215 );
not ( w_12215 , w_12216 );
and ( \3865_b0 , \3862_b0 , w_12217 );
and ( w_12216 ,  , w_12217 );
buf ( w_12215 , \3864_b1 );
not ( w_12215 , w_12218 );
not (  , w_12219 );
and ( w_12218 , w_12219 , \3864_b0 );
buf ( \3866_b1 , \3865_b1 );
not ( \3866_b1 , w_12220 );
not ( \3866_b0 , w_12221 );
and ( w_12220 , w_12221 , \3865_b0 );
or ( \3867_b1 , \2107_b1 , \2490_b1 );
not ( \2490_b1 , w_12222 );
and ( \3867_b0 , \2107_b0 , w_12223 );
and ( w_12222 , w_12223 , \2490_b0 );
or ( \3868_b1 , \c[11]_b1 , \b[5]_b1 );
xor ( \3868_b0 , \c[11]_b0 , w_12224 );
not ( w_12224 , w_12225 );
and ( w_12225 , \b[5]_b1 , \b[5]_b0 );
or ( \3869_b1 , \1689_b1 , \3868_b1 );
not ( \3868_b1 , w_12226 );
and ( \3869_b0 , \1689_b0 , w_12227 );
and ( w_12226 , w_12227 , \3868_b0 );
or ( \3870_b1 , \3867_b1 , w_12229 );
not ( w_12229 , w_12230 );
and ( \3870_b0 , \3867_b0 , w_12231 );
and ( w_12230 ,  , w_12231 );
buf ( w_12229 , \3869_b1 );
not ( w_12229 , w_12232 );
not (  , w_12233 );
and ( w_12232 , w_12233 , \3869_b0 );
buf ( \3871_b1 , \3870_b1 );
not ( \3871_b1 , w_12234 );
not ( \3871_b0 , w_12235 );
and ( w_12234 , w_12235 , \3870_b0 );
or ( \3872_b1 , \3866_b1 , \3871_b1 );
not ( \3871_b1 , w_12236 );
and ( \3872_b0 , \3866_b0 , w_12237 );
and ( w_12236 , w_12237 , \3871_b0 );
or ( \3873_b1 , \3865_b1 , \3870_b1 );
not ( \3870_b1 , w_12238 );
and ( \3873_b0 , \3865_b0 , w_12239 );
and ( w_12238 , w_12239 , \3870_b0 );
or ( \3874_b1 , \3872_b1 , w_12241 );
not ( w_12241 , w_12242 );
and ( \3874_b0 , \3872_b0 , w_12243 );
and ( w_12242 ,  , w_12243 );
buf ( w_12241 , \3873_b1 );
not ( w_12241 , w_12244 );
not (  , w_12245 );
and ( w_12244 , w_12245 , \3873_b0 );
buf ( \3875_b1 , \2483_b1 );
not ( \3875_b1 , w_12246 );
not ( \3875_b0 , w_12247 );
and ( w_12246 , w_12247 , \2483_b0 );
buf ( \3876_b1 , \2485_b1 );
not ( \3876_b1 , w_12248 );
not ( \3876_b0 , w_12249 );
and ( w_12248 , w_12249 , \2485_b0 );
buf ( \3877_b1 , \3876_b1 );
not ( \3877_b1 , w_12250 );
not ( \3877_b0 , w_12251 );
and ( w_12250 , w_12251 , \3876_b0 );
or ( \3878_b1 , \3875_b1 , w_12252 );
or ( \3878_b0 , \3875_b0 , \3877_b0 );
not ( \3877_b0 , w_12253 );
and ( w_12253 , w_12252 , \3877_b1 );
buf ( \3879_b1 , \2483_b1 );
not ( \3879_b1 , w_12254 );
not ( \3879_b0 , w_12255 );
and ( w_12254 , w_12255 , \2483_b0 );
buf ( \3880_b1 , \3879_b1 );
not ( \3880_b1 , w_12256 );
not ( \3880_b0 , w_12257 );
and ( w_12256 , w_12257 , \3879_b0 );
buf ( \3881_b1 , \2485_b1 );
not ( \3881_b1 , w_12258 );
not ( \3881_b0 , w_12259 );
and ( w_12258 , w_12259 , \2485_b0 );
or ( \3882_b1 , \3880_b1 , w_12260 );
or ( \3882_b0 , \3880_b0 , \3881_b0 );
not ( \3881_b0 , w_12261 );
and ( w_12261 , w_12260 , \3881_b1 );
or ( \3883_b1 , \3882_b1 , w_12263 );
not ( w_12263 , w_12264 );
and ( \3883_b0 , \3882_b0 , w_12265 );
and ( w_12264 ,  , w_12265 );
buf ( w_12263 , \2492_b1 );
not ( w_12263 , w_12266 );
not (  , w_12267 );
and ( w_12266 , w_12267 , \2492_b0 );
or ( \3884_b1 , \3878_b1 , w_12269 );
not ( w_12269 , w_12270 );
and ( \3884_b0 , \3878_b0 , w_12271 );
and ( w_12270 ,  , w_12271 );
buf ( w_12269 , \3883_b1 );
not ( w_12269 , w_12272 );
not (  , w_12273 );
and ( w_12272 , w_12273 , \3883_b0 );
or ( \3885_b1 , \3874_b1 , \3884_b1 );
xor ( \3885_b0 , \3874_b0 , w_12274 );
not ( w_12274 , w_12275 );
and ( w_12275 , \3884_b1 , \3884_b0 );
or ( \3886_b1 , \2535_b1 , \2541_b1 );
xor ( \3886_b0 , \2535_b0 , w_12276 );
not ( w_12276 , w_12277 );
and ( w_12277 , \2541_b1 , \2541_b0 );
or ( \3887_b1 , \3886_b1 , \2548_b1 );
not ( \2548_b1 , w_12278 );
and ( \3887_b0 , \3886_b0 , w_12279 );
and ( w_12278 , w_12279 , \2548_b0 );
or ( \3888_b1 , \2535_b1 , \2541_b1 );
not ( \2541_b1 , w_12280 );
and ( \3888_b0 , \2535_b0 , w_12281 );
and ( w_12280 , w_12281 , \2541_b0 );
or ( \3889_b1 , \3887_b1 , w_12282 );
or ( \3889_b0 , \3887_b0 , \3888_b0 );
not ( \3888_b0 , w_12283 );
and ( w_12283 , w_12282 , \3888_b1 );
or ( \3890_b1 , \2341_b1 , \2481_b1 );
not ( \2481_b1 , w_12284 );
and ( \3890_b0 , \2341_b0 , w_12285 );
and ( w_12284 , w_12285 , \2481_b0 );
or ( \3891_b1 , \c[13]_b1 , \b[3]_b1 );
xor ( \3891_b0 , \c[13]_b0 , w_12286 );
not ( w_12286 , w_12287 );
and ( w_12287 , \b[3]_b1 , \b[3]_b0 );
or ( \3892_b1 , \2075_b1 , \3891_b1 );
not ( \3891_b1 , w_12288 );
and ( \3892_b0 , \2075_b0 , w_12289 );
and ( w_12288 , w_12289 , \3891_b0 );
or ( \3893_b1 , \3890_b1 , w_12291 );
not ( w_12291 , w_12292 );
and ( \3893_b0 , \3890_b0 , w_12293 );
and ( w_12292 ,  , w_12293 );
buf ( w_12291 , \3892_b1 );
not ( w_12291 , w_12294 );
not (  , w_12295 );
and ( w_12294 , w_12295 , \3892_b0 );
or ( \3894_b1 , \c[15]_b1 , \c[14]_b1 );
xor ( \3894_b0 , \c[15]_b0 , w_12296 );
not ( w_12296 , w_12297 );
and ( w_12297 , \c[14]_b1 , \c[14]_b0 );
or ( \3895_b1 , \b[0]_b1 , \c[15]_b1 );
xor ( \3895_b0 , \b[0]_b0 , w_12298 );
not ( w_12298 , w_12299 );
and ( w_12299 , \c[15]_b1 , \c[15]_b0 );
or ( \3896_b1 , \3894_b1 , w_12301 );
not ( w_12301 , w_12302 );
and ( \3896_b0 , \3894_b0 , w_12303 );
and ( w_12302 ,  , w_12303 );
buf ( w_12301 , \3895_b1 );
not ( w_12301 , w_12304 );
not (  , w_12305 );
and ( w_12304 , w_12305 , \3895_b0 );
or ( \3897_b1 , \3896_b1 , w_12306 );
or ( \3897_b0 , \3896_b0 , \2534_b0 );
not ( \2534_b0 , w_12307 );
and ( w_12307 , w_12306 , \2534_b1 );
or ( \3898_b1 , \b[1]_b1 , \c[15]_b1 );
xor ( \3898_b0 , \b[1]_b0 , w_12308 );
not ( w_12308 , w_12309 );
and ( w_12309 , \c[15]_b1 , \c[15]_b0 );
or ( \3899_b1 , \2534_b1 , w_12311 );
not ( w_12311 , w_12312 );
and ( \3899_b0 , \2534_b0 , w_12313 );
and ( w_12312 ,  , w_12313 );
buf ( w_12311 , \3898_b1 );
not ( w_12311 , w_12314 );
not (  , w_12315 );
and ( w_12314 , w_12315 , \3898_b0 );
or ( \3900_b1 , \3897_b1 , w_12317 );
not ( w_12317 , w_12318 );
and ( \3900_b0 , \3897_b0 , w_12319 );
and ( w_12318 ,  , w_12319 );
buf ( w_12317 , \3899_b1 );
not ( w_12317 , w_12320 );
not (  , w_12321 );
and ( w_12320 , w_12321 , \3899_b0 );
or ( \3901_b1 , \3893_b1 , \3900_b1 );
xor ( \3901_b0 , \3893_b0 , w_12322 );
not ( w_12322 , w_12323 );
and ( w_12323 , \3900_b1 , \3900_b0 );
buf ( \3902_b1 , \2505_b1 );
not ( \3902_b1 , w_12324 );
not ( \3902_b0 , w_12325 );
and ( w_12324 , w_12325 , \2505_b0 );
buf ( \3903_b1 , \1743_b1 );
not ( \3903_b1 , w_12326 );
not ( \3903_b0 , w_12327 );
and ( w_12326 , w_12327 , \1743_b0 );
or ( \3904_b1 , \3902_b1 , w_12328 );
or ( \3904_b0 , \3902_b0 , \3903_b0 );
not ( \3903_b0 , w_12329 );
and ( w_12329 , w_12328 , \3903_b1 );
buf ( \3905_b1 , \c[7]_b1 );
not ( \3905_b1 , w_12330 );
not ( \3905_b0 , w_12331 );
and ( w_12330 , w_12331 , \c[7]_b0 );
or ( \3906_b1 , \3905_b1 , w_12333 );
not ( w_12333 , w_12334 );
and ( \3906_b0 , \3905_b0 , w_12335 );
and ( w_12334 ,  , w_12335 );
buf ( w_12333 , \b[9]_b1 );
not ( w_12333 , w_12336 );
not (  , w_12337 );
and ( w_12336 , w_12337 , \b[9]_b0 );
buf ( \3907_b1 , \3906_b1 );
not ( \3907_b1 , w_12338 );
not ( \3907_b0 , w_12339 );
and ( w_12338 , w_12339 , \3906_b0 );
buf ( \3908_b1 , \b[9]_b1 );
not ( \3908_b1 , w_12340 );
not ( \3908_b0 , w_12341 );
and ( w_12340 , w_12341 , \b[9]_b0 );
or ( \3909_b1 , \3908_b1 , w_12343 );
not ( w_12343 , w_12344 );
and ( \3909_b0 , \3908_b0 , w_12345 );
and ( w_12344 ,  , w_12345 );
buf ( w_12343 , \c[7]_b1 );
not ( w_12343 , w_12346 );
not (  , w_12347 );
and ( w_12346 , w_12347 , \c[7]_b0 );
buf ( \3910_b1 , \3909_b1 );
not ( \3910_b1 , w_12348 );
not ( \3910_b0 , w_12349 );
and ( w_12348 , w_12349 , \3909_b0 );
or ( \3911_b1 , \3907_b1 , w_12350 );
or ( \3911_b0 , \3907_b0 , \3910_b0 );
not ( \3910_b0 , w_12351 );
and ( w_12351 , w_12350 , \3910_b1 );
or ( \3912_b1 , \3911_b1 , w_12353 );
not ( w_12353 , w_12354 );
and ( \3912_b0 , \3911_b0 , w_12355 );
and ( w_12354 ,  , w_12355 );
buf ( w_12353 , \1747_b1 );
not ( w_12353 , w_12356 );
not (  , w_12357 );
and ( w_12356 , w_12357 , \1747_b0 );
or ( \3913_b1 , \3904_b1 , w_12359 );
not ( w_12359 , w_12360 );
and ( \3913_b0 , \3904_b0 , w_12361 );
and ( w_12360 ,  , w_12361 );
buf ( w_12359 , \3912_b1 );
not ( w_12359 , w_12362 );
not (  , w_12363 );
and ( w_12362 , w_12363 , \3912_b0 );
or ( \3914_b1 , \3901_b1 , w_12364 );
xor ( \3914_b0 , \3901_b0 , w_12366 );
not ( w_12366 , w_12367 );
and ( w_12367 , w_12364 , w_12365 );
buf ( w_12364 , \3913_b1 );
not ( w_12364 , w_12368 );
not ( w_12365 , w_12369 );
and ( w_12368 , w_12369 , \3913_b0 );
buf ( \3915_b1 , \3914_b1 );
not ( \3915_b1 , w_12370 );
not ( \3915_b0 , w_12371 );
and ( w_12370 , w_12371 , \3914_b0 );
or ( \3916_b1 , \3889_b1 , \3915_b1 );
xor ( \3916_b0 , \3889_b0 , w_12372 );
not ( w_12372 , w_12373 );
and ( w_12373 , \3915_b1 , \3915_b0 );
or ( \3917_b1 , \3885_b1 , w_12374 );
xor ( \3917_b0 , \3885_b0 , w_12376 );
not ( w_12376 , w_12377 );
and ( w_12377 , w_12374 , w_12375 );
buf ( w_12374 , \3916_b1 );
not ( w_12374 , w_12378 );
not ( w_12375 , w_12379 );
and ( w_12378 , w_12379 , \3916_b0 );
or ( \3918_b1 , \3859_b1 , w_12380 );
xor ( \3918_b0 , \3859_b0 , w_12382 );
not ( w_12382 , w_12383 );
and ( w_12383 , w_12380 , w_12381 );
buf ( w_12380 , \3917_b1 );
not ( w_12380 , w_12384 );
not ( w_12381 , w_12385 );
and ( w_12384 , w_12385 , \3917_b0 );
or ( \3919_b1 , \3852_b1 , \3918_b1 );
xor ( \3919_b0 , \3852_b0 , w_12386 );
not ( w_12386 , w_12387 );
and ( w_12387 , \3918_b1 , \3918_b0 );
or ( \3920_b1 , \3810_b1 , w_12388 );
xor ( \3920_b0 , \3810_b0 , w_12390 );
not ( w_12390 , w_12391 );
and ( w_12391 , w_12388 , w_12389 );
buf ( w_12388 , \3919_b1 );
not ( w_12388 , w_12392 );
not ( w_12389 , w_12393 );
and ( w_12392 , w_12393 , \3919_b0 );
buf ( \3921_b1 , \3920_b1 );
not ( \3921_b1 , w_12394 );
not ( \3921_b0 , w_12395 );
and ( w_12394 , w_12395 , \3920_b0 );
or ( \3922_b1 , \3802_b1 , \3921_b1 );
not ( \3921_b1 , w_12396 );
and ( \3922_b0 , \3802_b0 , w_12397 );
and ( w_12396 , w_12397 , \3921_b0 );
buf ( \3923_b1 , \3802_b1 );
not ( \3923_b1 , w_12398 );
not ( \3923_b0 , w_12399 );
and ( w_12398 , w_12399 , \3802_b0 );
or ( \3924_b1 , \3923_b1 , \3920_b1 );
not ( \3920_b1 , w_12400 );
and ( \3924_b0 , \3923_b0 , w_12401 );
and ( w_12400 , w_12401 , \3920_b0 );
or ( \3925_b1 , \3922_b1 , w_12403 );
not ( w_12403 , w_12404 );
and ( \3925_b0 , \3922_b0 , w_12405 );
and ( w_12404 ,  , w_12405 );
buf ( w_12403 , \3924_b1 );
not ( w_12403 , w_12406 );
not (  , w_12407 );
and ( w_12406 , w_12407 , \3924_b0 );
or ( \3926_b1 , \3925_b1 , w_12409 );
not ( w_12409 , w_12410 );
and ( \3926_b0 , \3925_b0 , w_12411 );
and ( w_12410 ,  , w_12411 );
buf ( w_12409 , \2413_b1 );
not ( w_12409 , w_12412 );
not (  , w_12413 );
and ( w_12412 , w_12413 , \2413_b0 );
or ( \3927_b1 , \c[15]_b1 , w_12415 );
not ( w_12415 , w_12416 );
and ( \3927_b0 , \c[15]_b0 , w_12417 );
and ( w_12416 ,  , w_12417 );
buf ( w_12415 , \d[15]_b1 );
not ( w_12415 , w_12418 );
not (  , w_12419 );
and ( w_12418 , w_12419 , \d[15]_b0 );
buf ( \3928_b1 , \3927_b1 );
not ( \3928_b1 , w_12420 );
not ( \3928_b0 , w_12421 );
and ( w_12420 , w_12421 , \3927_b0 );
or ( \3929_b1 , \c[15]_b1 , w_12423 );
not ( w_12423 , w_12424 );
and ( \3929_b0 , \c[15]_b0 , w_12425 );
and ( w_12424 ,  , w_12425 );
buf ( w_12423 , \d[15]_b1 );
not ( w_12423 , w_12426 );
not (  , w_12427 );
and ( w_12426 , w_12427 , \d[15]_b0 );
or ( \3930_b1 , \3928_b1 , w_12429 );
not ( w_12429 , w_12430 );
and ( \3930_b0 , \3928_b0 , w_12431 );
and ( w_12430 ,  , w_12431 );
buf ( w_12429 , \3929_b1 );
not ( w_12429 , w_12432 );
not (  , w_12433 );
and ( w_12432 , w_12433 , \3929_b0 );
or ( \3931_b1 , \c[1]_b1 , w_12435 );
not ( w_12435 , w_12436 );
and ( \3931_b0 , \c[1]_b0 , w_12437 );
and ( w_12436 ,  , w_12437 );
buf ( w_12435 , \d[1]_b1 );
not ( w_12435 , w_12438 );
not (  , w_12439 );
and ( w_12438 , w_12439 , \d[1]_b0 );
or ( \3932_b1 , \c[0]_b1 , w_12441 );
not ( w_12441 , w_12442 );
and ( \3932_b0 , \c[0]_b0 , w_12443 );
and ( w_12442 ,  , w_12443 );
buf ( w_12441 , \d[0]_b1 );
not ( w_12441 , w_12444 );
not (  , w_12445 );
and ( w_12444 , w_12445 , \d[0]_b0 );
or ( \3933_b1 , \3931_b1 , \3932_b1 );
not ( \3932_b1 , w_12446 );
and ( \3933_b0 , \3931_b0 , w_12447 );
and ( w_12446 , w_12447 , \3932_b0 );
or ( \3934_b1 , \c[1]_b1 , w_12449 );
not ( w_12449 , w_12450 );
and ( \3934_b0 , \c[1]_b0 , w_12451 );
and ( w_12450 ,  , w_12451 );
buf ( w_12449 , \d[1]_b1 );
not ( w_12449 , w_12452 );
not (  , w_12453 );
and ( w_12452 , w_12453 , \d[1]_b0 );
or ( \3935_b1 , \c[2]_b1 , w_12455 );
not ( w_12455 , w_12456 );
and ( \3935_b0 , \c[2]_b0 , w_12457 );
and ( w_12456 ,  , w_12457 );
buf ( w_12455 , \d[2]_b1 );
not ( w_12455 , w_12458 );
not (  , w_12459 );
and ( w_12458 , w_12459 , \d[2]_b0 );
buf ( \3937_b1 , \3936_b1 );
not ( \3937_b1 , w_12460 );
not ( \3937_b0 , w_12461 );
and ( w_12460 , w_12461 , \3936_b0 );
or ( \3938_b1 , \c[3]_b1 , w_12463 );
not ( w_12463 , w_12464 );
and ( \3938_b0 , \c[3]_b0 , w_12465 );
and ( w_12464 ,  , w_12465 );
buf ( w_12463 , \d[3]_b1 );
not ( w_12463 , w_12466 );
not (  , w_12467 );
and ( w_12466 , w_12467 , \d[3]_b0 );
or ( \3939_b1 , \c[2]_b1 , w_12469 );
not ( w_12469 , w_12470 );
and ( \3939_b0 , \c[2]_b0 , w_12471 );
and ( w_12470 ,  , w_12471 );
buf ( w_12469 , \d[2]_b1 );
not ( w_12469 , w_12472 );
not (  , w_12473 );
and ( w_12472 , w_12473 , \d[2]_b0 );
or ( \3941_b1 , \c[5]_b1 , w_12475 );
not ( w_12475 , w_12476 );
and ( \3941_b0 , \c[5]_b0 , w_12477 );
and ( w_12476 ,  , w_12477 );
buf ( w_12475 , \d[5]_b1 );
not ( w_12475 , w_12478 );
not (  , w_12479 );
and ( w_12478 , w_12479 , \d[5]_b0 );
or ( \3942_b1 , \c[4]_b1 , w_12481 );
not ( w_12481 , w_12482 );
and ( \3942_b0 , \c[4]_b0 , w_12483 );
and ( w_12482 ,  , w_12483 );
buf ( w_12481 , \d[4]_b1 );
not ( w_12481 , w_12484 );
not (  , w_12485 );
and ( w_12484 , w_12485 , \d[4]_b0 );
or ( \3943_b1 , \3941_b1 , w_12487 );
not ( w_12487 , w_12488 );
and ( \3943_b0 , \3941_b0 , w_12489 );
and ( w_12488 ,  , w_12489 );
buf ( w_12487 , \3942_b1 );
not ( w_12487 , w_12490 );
not (  , w_12491 );
and ( w_12490 , w_12491 , \3942_b0 );
or ( \3944_b1 , \c[7]_b1 , w_12493 );
not ( w_12493 , w_12494 );
and ( \3944_b0 , \c[7]_b0 , w_12495 );
and ( w_12494 ,  , w_12495 );
buf ( w_12493 , \d[7]_b1 );
not ( w_12493 , w_12496 );
not (  , w_12497 );
and ( w_12496 , w_12497 , \d[7]_b0 );
or ( \3945_b1 , \c[6]_b1 , w_12499 );
not ( w_12499 , w_12500 );
and ( \3945_b0 , \c[6]_b0 , w_12501 );
and ( w_12500 ,  , w_12501 );
buf ( w_12499 , \d[6]_b1 );
not ( w_12499 , w_12502 );
not (  , w_12503 );
and ( w_12502 , w_12503 , \d[6]_b0 );
or ( \3946_b1 , \3944_b1 , w_12505 );
not ( w_12505 , w_12506 );
and ( \3946_b0 , \3944_b0 , w_12507 );
and ( w_12506 ,  , w_12507 );
buf ( w_12505 , \3945_b1 );
not ( w_12505 , w_12508 );
not (  , w_12509 );
and ( w_12508 , w_12509 , \3945_b0 );
or ( \3947_b1 , \c[3]_b1 , w_12511 );
not ( w_12511 , w_12512 );
and ( \3947_b0 , \c[3]_b0 , w_12513 );
and ( w_12512 ,  , w_12513 );
buf ( w_12511 , \d[3]_b1 );
not ( w_12511 , w_12514 );
not (  , w_12515 );
and ( w_12514 , w_12515 , \d[3]_b0 );
buf ( \3948_b1 , \3947_b1 );
not ( \3948_b1 , w_12516 );
not ( \3948_b0 , w_12517 );
and ( w_12516 , w_12517 , \3947_b0 );
or ( \3950_b1 , \c[4]_b1 , w_12519 );
not ( w_12519 , w_12520 );
and ( \3950_b0 , \c[4]_b0 , w_12521 );
and ( w_12520 ,  , w_12521 );
buf ( w_12519 , \d[4]_b1 );
not ( w_12519 , w_12522 );
not (  , w_12523 );
and ( w_12522 , w_12523 , \d[4]_b0 );
or ( \3951_b1 , \3941_b1 , w_12525 );
not ( w_12525 , w_12526 );
and ( \3951_b0 , \3941_b0 , w_12527 );
and ( w_12526 ,  , w_12527 );
buf ( w_12525 , \3950_b1 );
not ( w_12525 , w_12528 );
not (  , w_12529 );
and ( w_12528 , w_12529 , \3950_b0 );
or ( \3952_b1 , \c[6]_b1 , w_12531 );
not ( w_12531 , w_12532 );
and ( \3952_b0 , \c[6]_b0 , w_12533 );
and ( w_12532 ,  , w_12533 );
buf ( w_12531 , \d[6]_b1 );
not ( w_12531 , w_12534 );
not (  , w_12535 );
and ( w_12534 , w_12535 , \d[6]_b0 );
or ( \3953_b1 , \c[7]_b1 , w_12537 );
not ( w_12537 , w_12538 );
and ( \3953_b0 , \c[7]_b0 , w_12539 );
and ( w_12538 ,  , w_12539 );
buf ( w_12537 , \d[7]_b1 );
not ( w_12537 , w_12540 );
not (  , w_12541 );
and ( w_12540 , w_12541 , \d[7]_b0 );
or ( \3954_b1 , \c[5]_b1 , w_12543 );
not ( w_12543 , w_12544 );
and ( \3954_b0 , \c[5]_b0 , w_12545 );
and ( w_12544 ,  , w_12545 );
buf ( w_12543 , \d[5]_b1 );
not ( w_12543 , w_12546 );
not (  , w_12547 );
and ( w_12546 , w_12547 , \d[5]_b0 );
or ( \3956_b1 , \3951_b1 , w_12548 );
or ( \3956_b0 , \3951_b0 , \3955_b0 );
not ( \3955_b0 , w_12549 );
and ( w_12549 , w_12548 , \3955_b1 );
buf ( \3957_b1 , \3953_b1 );
not ( \3957_b1 , w_12550 );
not ( \3957_b0 , w_12551 );
and ( w_12550 , w_12551 , \3953_b0 );
or ( \3958_b1 , \3946_b1 , w_12552 );
or ( \3958_b0 , \3946_b0 , \3957_b0 );
not ( \3957_b0 , w_12553 );
and ( w_12553 , w_12552 , \3957_b1 );
or ( \3959_b1 , \3956_b1 , w_12555 );
not ( w_12555 , w_12556 );
and ( \3959_b0 , \3956_b0 , w_12557 );
and ( w_12556 ,  , w_12557 );
buf ( w_12555 , \3958_b1 );
not ( w_12555 , w_12558 );
not (  , w_12559 );
and ( w_12558 , w_12559 , \3958_b0 );
or ( \3960_b1 , \3949_b1 , w_12561 );
not ( w_12561 , w_12562 );
and ( \3960_b0 , \3949_b0 , w_12563 );
and ( w_12562 ,  , w_12563 );
buf ( w_12561 , \3959_b1 );
not ( w_12561 , w_12564 );
not (  , w_12565 );
and ( w_12564 , w_12565 , \3959_b0 );
or ( \3961_b1 , \c[11]_b1 , w_12567 );
not ( w_12567 , w_12568 );
and ( \3961_b0 , \c[11]_b0 , w_12569 );
and ( w_12568 ,  , w_12569 );
buf ( w_12567 , \d[11]_b1 );
not ( w_12567 , w_12570 );
not (  , w_12571 );
and ( w_12570 , w_12571 , \d[11]_b0 );
or ( \3962_b1 , \c[10]_b1 , w_12573 );
not ( w_12573 , w_12574 );
and ( \3962_b0 , \c[10]_b0 , w_12575 );
and ( w_12574 ,  , w_12575 );
buf ( w_12573 , \d[10]_b1 );
not ( w_12573 , w_12576 );
not (  , w_12577 );
and ( w_12576 , w_12577 , \d[10]_b0 );
or ( \3963_b1 , \3961_b1 , w_12579 );
not ( w_12579 , w_12580 );
and ( \3963_b0 , \3961_b0 , w_12581 );
and ( w_12580 ,  , w_12581 );
buf ( w_12579 , \3962_b1 );
not ( w_12579 , w_12582 );
not (  , w_12583 );
and ( w_12582 , w_12583 , \3962_b0 );
or ( \3964_b1 , \c[9]_b1 , w_12585 );
not ( w_12585 , w_12586 );
and ( \3964_b0 , \c[9]_b0 , w_12587 );
and ( w_12586 ,  , w_12587 );
buf ( w_12585 , \d[9]_b1 );
not ( w_12585 , w_12588 );
not (  , w_12589 );
and ( w_12588 , w_12589 , \d[9]_b0 );
or ( \3965_b1 , \c[8]_b1 , w_12591 );
not ( w_12591 , w_12592 );
and ( \3965_b0 , \c[8]_b0 , w_12593 );
and ( w_12592 ,  , w_12593 );
buf ( w_12591 , \d[8]_b1 );
not ( w_12591 , w_12594 );
not (  , w_12595 );
and ( w_12594 , w_12595 , \d[8]_b0 );
or ( \3966_b1 , \3964_b1 , w_12597 );
not ( w_12597 , w_12598 );
and ( \3966_b0 , \3964_b0 , w_12599 );
and ( w_12598 ,  , w_12599 );
buf ( w_12597 , \3965_b1 );
not ( w_12597 , w_12600 );
not (  , w_12601 );
and ( w_12600 , w_12601 , \3965_b0 );
or ( \3967_b1 , \3963_b1 , w_12603 );
not ( w_12603 , w_12604 );
and ( \3967_b0 , \3963_b0 , w_12605 );
and ( w_12604 ,  , w_12605 );
buf ( w_12603 , \3966_b1 );
not ( w_12603 , w_12606 );
not (  , w_12607 );
and ( w_12606 , w_12607 , \3966_b0 );
buf ( \3968_b1 , \3967_b1 );
not ( \3968_b1 , w_12608 );
not ( \3968_b0 , w_12609 );
and ( w_12608 , w_12609 , \3967_b0 );
or ( \3969_b1 , \c[14]_b1 , w_12611 );
not ( w_12611 , w_12612 );
and ( \3969_b0 , \c[14]_b0 , w_12613 );
and ( w_12612 ,  , w_12613 );
buf ( w_12611 , \d[14]_b1 );
not ( w_12611 , w_12614 );
not (  , w_12615 );
and ( w_12614 , w_12615 , \d[14]_b0 );
buf ( \3970_b1 , \3969_b1 );
not ( \3970_b1 , w_12616 );
not ( \3970_b0 , w_12617 );
and ( w_12616 , w_12617 , \3969_b0 );
or ( \3971_b1 , \c[13]_b1 , w_12619 );
not ( w_12619 , w_12620 );
and ( \3971_b0 , \c[13]_b0 , w_12621 );
and ( w_12620 ,  , w_12621 );
buf ( w_12619 , \d[13]_b1 );
not ( w_12619 , w_12622 );
not (  , w_12623 );
and ( w_12622 , w_12623 , \d[13]_b0 );
or ( \3972_b1 , \c[12]_b1 , w_12625 );
not ( w_12625 , w_12626 );
and ( \3972_b0 , \c[12]_b0 , w_12627 );
and ( w_12626 ,  , w_12627 );
buf ( w_12625 , \d[12]_b1 );
not ( w_12625 , w_12628 );
not (  , w_12629 );
and ( w_12628 , w_12629 , \d[12]_b0 );
or ( \3973_b1 , \3971_b1 , w_12631 );
not ( w_12631 , w_12632 );
and ( \3973_b0 , \3971_b0 , w_12633 );
and ( w_12632 ,  , w_12633 );
buf ( w_12631 , \3972_b1 );
not ( w_12631 , w_12634 );
not (  , w_12635 );
and ( w_12634 , w_12635 , \3972_b0 );
or ( \3974_b1 , \3970_b1 , w_12637 );
not ( w_12637 , w_12638 );
and ( \3974_b0 , \3970_b0 , w_12639 );
and ( w_12638 ,  , w_12639 );
buf ( w_12637 , \3973_b1 );
not ( w_12637 , w_12640 );
not (  , w_12641 );
and ( w_12640 , w_12641 , \3973_b0 );
buf ( \3975_b1 , \3974_b1 );
not ( \3975_b1 , w_12642 );
not ( \3975_b0 , w_12643 );
and ( w_12642 , w_12643 , \3974_b0 );
or ( \3977_b1 , \c[8]_b1 , w_12645 );
not ( w_12645 , w_12646 );
and ( \3977_b0 , \c[8]_b0 , w_12647 );
and ( w_12646 ,  , w_12647 );
buf ( w_12645 , \d[8]_b1 );
not ( w_12645 , w_12648 );
not (  , w_12649 );
and ( w_12648 , w_12649 , \d[8]_b0 );
or ( \3978_b1 , \3964_b1 , w_12650 );
or ( \3978_b0 , \3964_b0 , \3977_b0 );
not ( \3977_b0 , w_12651 );
and ( w_12651 , w_12650 , \3977_b1 );
or ( \3979_b1 , \c[9]_b1 , w_12653 );
not ( w_12653 , w_12654 );
and ( \3979_b0 , \c[9]_b0 , w_12655 );
and ( w_12654 ,  , w_12655 );
buf ( w_12653 , \d[9]_b1 );
not ( w_12653 , w_12656 );
not (  , w_12657 );
and ( w_12656 , w_12657 , \d[9]_b0 );
or ( \3980_b1 , \3978_b1 , w_12659 );
not ( w_12659 , w_12660 );
and ( \3980_b0 , \3978_b0 , w_12661 );
and ( w_12660 ,  , w_12661 );
buf ( w_12659 , \3979_b1 );
not ( w_12659 , w_12662 );
not (  , w_12663 );
and ( w_12662 , w_12663 , \3979_b0 );
or ( \3981_b1 , \3963_b1 , \3980_b1 );
not ( \3980_b1 , w_12664 );
and ( \3981_b0 , \3963_b0 , w_12665 );
and ( w_12664 , w_12665 , \3980_b0 );
or ( \3982_b1 , \c[10]_b1 , w_12667 );
not ( w_12667 , w_12668 );
and ( \3982_b0 , \c[10]_b0 , w_12669 );
and ( w_12668 ,  , w_12669 );
buf ( w_12667 , \d[10]_b1 );
not ( w_12667 , w_12670 );
not (  , w_12671 );
and ( w_12670 , w_12671 , \d[10]_b0 );
or ( \3983_b1 , \3961_b1 , w_12672 );
or ( \3983_b0 , \3961_b0 , \3982_b0 );
not ( \3982_b0 , w_12673 );
and ( w_12673 , w_12672 , \3982_b1 );
or ( \3984_b1 , \c[11]_b1 , w_12675 );
not ( w_12675 , w_12676 );
and ( \3984_b0 , \c[11]_b0 , w_12677 );
and ( w_12676 ,  , w_12677 );
buf ( w_12675 , \d[11]_b1 );
not ( w_12675 , w_12678 );
not (  , w_12679 );
and ( w_12678 , w_12679 , \d[11]_b0 );
or ( \3985_b1 , \3983_b1 , w_12681 );
not ( w_12681 , w_12682 );
and ( \3985_b0 , \3983_b0 , w_12683 );
and ( w_12682 ,  , w_12683 );
buf ( w_12681 , \3984_b1 );
not ( w_12681 , w_12684 );
not (  , w_12685 );
and ( w_12684 , w_12685 , \3984_b0 );
or ( \3986_b1 , \3981_b1 , w_12687 );
not ( w_12687 , w_12688 );
and ( \3986_b0 , \3981_b0 , w_12689 );
and ( w_12688 ,  , w_12689 );
buf ( w_12687 , \3985_b1 );
not ( w_12687 , w_12690 );
not (  , w_12691 );
and ( w_12690 , w_12691 , \3985_b0 );
or ( \3987_b1 , \3986_b1 , w_12692 );
or ( \3987_b0 , \3986_b0 , \3974_b0 );
not ( \3974_b0 , w_12693 );
and ( w_12693 , w_12692 , \3974_b1 );
or ( \3988_b1 , \c[12]_b1 , w_12695 );
not ( w_12695 , w_12696 );
and ( \3988_b0 , \c[12]_b0 , w_12697 );
and ( w_12696 ,  , w_12697 );
buf ( w_12695 , \d[12]_b1 );
not ( w_12695 , w_12698 );
not (  , w_12699 );
and ( w_12698 , w_12699 , \d[12]_b0 );
or ( \3989_b1 , \3971_b1 , w_12700 );
or ( \3989_b0 , \3971_b0 , \3988_b0 );
not ( \3988_b0 , w_12701 );
and ( w_12701 , w_12700 , \3988_b1 );
or ( \3990_b1 , \c[13]_b1 , w_12703 );
not ( w_12703 , w_12704 );
and ( \3990_b0 , \c[13]_b0 , w_12705 );
and ( w_12704 ,  , w_12705 );
buf ( w_12703 , \d[13]_b1 );
not ( w_12703 , w_12706 );
not (  , w_12707 );
and ( w_12706 , w_12707 , \d[13]_b0 );
or ( \3991_b1 , \3989_b1 , w_12709 );
not ( w_12709 , w_12710 );
and ( \3991_b0 , \3989_b0 , w_12711 );
and ( w_12710 ,  , w_12711 );
buf ( w_12709 , \3990_b1 );
not ( w_12709 , w_12712 );
not (  , w_12713 );
and ( w_12712 , w_12713 , \3990_b0 );
buf ( \3992_b1 , \3991_b1 );
not ( \3992_b1 , w_12714 );
not ( \3992_b0 , w_12715 );
and ( w_12714 , w_12715 , \3991_b0 );
or ( \3993_b1 , \3969_b1 , w_12716 );
or ( \3993_b0 , \3969_b0 , \3992_b0 );
not ( \3992_b0 , w_12717 );
and ( w_12717 , w_12716 , \3992_b1 );
or ( \3994_b1 , \c[14]_b1 , w_12719 );
not ( w_12719 , w_12720 );
and ( \3994_b0 , \c[14]_b0 , w_12721 );
and ( w_12720 ,  , w_12721 );
buf ( w_12719 , \d[14]_b1 );
not ( w_12719 , w_12722 );
not (  , w_12723 );
and ( w_12722 , w_12723 , \d[14]_b0 );
or ( \3996_b1 , \3976_b1 , w_12725 );
not ( w_12725 , w_12726 );
and ( \3996_b0 , \3976_b0 , w_12727 );
and ( w_12726 ,  , w_12727 );
buf ( w_12725 , \3995_b1 );
not ( w_12725 , w_12728 );
not (  , w_12729 );
and ( w_12728 , w_12729 , \3995_b0 );
or ( \3997_b1 , \3930_b1 , \3996_b1 );
xor ( \3997_b0 , \3930_b0 , w_12730 );
not ( w_12730 , w_12731 );
and ( w_12731 , \3996_b1 , \3996_b0 );
buf ( \3998_b1 , \3944_b1 );
not ( \3998_b1 , w_12732 );
not ( \3998_b0 , w_12733 );
and ( w_12732 , w_12733 , \3944_b0 );
or ( \3999_b1 , \3998_b1 , w_12735 );
not ( w_12735 , w_12736 );
and ( \3999_b0 , \3998_b0 , w_12737 );
and ( w_12736 ,  , w_12737 );
buf ( w_12735 , \3953_b1 );
not ( w_12735 , w_12738 );
not (  , w_12739 );
and ( w_12738 , w_12739 , \3953_b0 );
or ( \4000_b1 , \3934_b1 , w_12740 );
or ( \4000_b0 , \3934_b0 , \3932_b0 );
not ( \3932_b0 , w_12741 );
and ( w_12741 , w_12740 , \3932_b1 );
or ( \4001_b1 , \4000_b1 , w_12743 );
not ( w_12743 , w_12744 );
and ( \4001_b0 , \4000_b0 , w_12745 );
and ( w_12744 ,  , w_12745 );
buf ( w_12743 , \3931_b1 );
not ( w_12743 , w_12746 );
not (  , w_12747 );
and ( w_12746 , w_12747 , \3931_b0 );
or ( \4002_b1 , \3947_b1 , w_12749 );
not ( w_12749 , w_12750 );
and ( \4002_b0 , \3947_b0 , w_12751 );
and ( w_12750 ,  , w_12751 );
buf ( w_12749 , \3935_b1 );
not ( w_12749 , w_12752 );
not (  , w_12753 );
and ( w_12752 , w_12753 , \3935_b0 );
or ( \4003_b1 , \4001_b1 , \4002_b1 );
not ( \4002_b1 , w_12754 );
and ( \4003_b0 , \4001_b0 , w_12755 );
and ( w_12754 , w_12755 , \4002_b0 );
or ( \4004_b1 , \3947_b1 , w_12756 );
or ( \4004_b0 , \3947_b0 , \3939_b0 );
not ( \3939_b0 , w_12757 );
and ( w_12757 , w_12756 , \3939_b1 );
or ( \4005_b1 , \4004_b1 , w_12759 );
not ( w_12759 , w_12760 );
and ( \4005_b0 , \4004_b0 , w_12761 );
and ( w_12760 ,  , w_12761 );
buf ( w_12759 , \3938_b1 );
not ( w_12759 , w_12762 );
not (  , w_12763 );
and ( w_12762 , w_12763 , \3938_b0 );
or ( \4006_b1 , \4003_b1 , w_12765 );
not ( w_12765 , w_12766 );
and ( \4006_b0 , \4003_b0 , w_12767 );
and ( w_12766 ,  , w_12767 );
buf ( w_12765 , \4005_b1 );
not ( w_12765 , w_12768 );
not (  , w_12769 );
and ( w_12768 , w_12769 , \4005_b0 );
buf ( \4007_b1 , \4006_b1 );
not ( \4007_b1 , w_12770 );
not ( \4007_b0 , w_12771 );
and ( w_12770 , w_12771 , \4006_b0 );
buf ( \4008_b1 , \3945_b1 );
not ( \4008_b1 , w_12772 );
not ( \4008_b0 , w_12773 );
and ( w_12772 , w_12773 , \3945_b0 );
buf ( \4010_b1 , \4008_b1 );
not ( \4010_b1 , w_12774 );
not ( \4010_b0 , w_12775 );
and ( w_12774 , w_12775 , \4008_b0 );
buf ( \4011_b1 , \3951_b1 );
not ( \4011_b1 , w_12776 );
not ( \4011_b0 , w_12777 );
and ( w_12776 , w_12777 , \3951_b0 );
or ( \4012_b1 , \4011_b1 , w_12779 );
not ( w_12779 , w_12780 );
and ( \4012_b0 , \4011_b0 , w_12781 );
and ( w_12780 ,  , w_12781 );
buf ( w_12779 , \3954_b1 );
not ( w_12779 , w_12782 );
not (  , w_12783 );
and ( w_12782 , w_12783 , \3954_b0 );
buf ( \4013_b1 , \4012_b1 );
not ( \4013_b1 , w_12784 );
not ( \4013_b0 , w_12785 );
and ( w_12784 , w_12785 , \4012_b0 );
or ( \4014_b1 , \4010_b1 , w_12786 );
or ( \4014_b0 , \4010_b0 , \4013_b0 );
not ( \4013_b0 , w_12787 );
and ( w_12787 , w_12786 , \4013_b1 );
or ( \4015_b1 , \4014_b1 , w_12789 );
not ( w_12789 , w_12790 );
and ( \4015_b0 , \4014_b0 , w_12791 );
and ( w_12790 ,  , w_12791 );
buf ( w_12789 , \3952_b1 );
not ( w_12789 , w_12792 );
not (  , w_12793 );
and ( w_12792 , w_12793 , \3952_b0 );
or ( \4016_b1 , \4009_b1 , w_12795 );
not ( w_12795 , w_12796 );
and ( \4016_b0 , \4009_b0 , w_12797 );
and ( w_12796 ,  , w_12797 );
buf ( w_12795 , \4015_b1 );
not ( w_12795 , w_12798 );
not (  , w_12799 );
and ( w_12798 , w_12799 , \4015_b0 );
or ( \4017_b1 , \3999_b1 , \4016_b1 );
xor ( \4017_b0 , \3999_b0 , w_12800 );
not ( w_12800 , w_12801 );
and ( w_12801 , \4016_b1 , \4016_b0 );
or ( \4018_b1 , \4008_b1 , w_12803 );
not ( w_12803 , w_12804 );
and ( \4018_b0 , \4008_b0 , w_12805 );
and ( w_12804 ,  , w_12805 );
buf ( w_12803 , \3952_b1 );
not ( w_12803 , w_12806 );
not (  , w_12807 );
and ( w_12806 , w_12807 , \3952_b0 );
or ( \4019_b1 , \4007_b1 , \3943_b1 );
not ( \3943_b1 , w_12808 );
and ( \4019_b0 , \4007_b0 , w_12809 );
and ( w_12808 , w_12809 , \3943_b0 );
or ( \4020_b1 , \4019_b1 , w_12811 );
not ( w_12811 , w_12812 );
and ( \4020_b0 , \4019_b0 , w_12813 );
and ( w_12812 ,  , w_12813 );
buf ( w_12811 , \4012_b1 );
not ( w_12811 , w_12814 );
not (  , w_12815 );
and ( w_12814 , w_12815 , \4012_b0 );
or ( \4021_b1 , \4018_b1 , \4020_b1 );
xor ( \4021_b0 , \4018_b0 , w_12816 );
not ( w_12816 , w_12817 );
and ( w_12817 , \4020_b1 , \4020_b0 );
buf ( \4022_b1 , \3954_b1 );
not ( \4022_b1 , w_12818 );
not ( \4022_b0 , w_12819 );
and ( w_12818 , w_12819 , \3954_b0 );
or ( \4023_b1 , \4022_b1 , w_12821 );
not ( w_12821 , w_12822 );
and ( \4023_b0 , \4022_b0 , w_12823 );
and ( w_12822 ,  , w_12823 );
buf ( w_12821 , \3941_b1 );
not ( w_12821 , w_12824 );
not (  , w_12825 );
and ( w_12824 , w_12825 , \3941_b0 );
or ( \4024_b1 , \4006_b1 , w_12826 );
or ( \4024_b0 , \4006_b0 , \3942_b0 );
not ( \3942_b0 , w_12827 );
and ( w_12827 , w_12826 , \3942_b1 );
or ( \4025_b1 , \4024_b1 , w_12829 );
not ( w_12829 , w_12830 );
and ( \4025_b0 , \4024_b0 , w_12831 );
and ( w_12830 ,  , w_12831 );
buf ( w_12829 , \3950_b1 );
not ( w_12829 , w_12832 );
not (  , w_12833 );
and ( w_12832 , w_12833 , \3950_b0 );
or ( \4026_b1 , \4023_b1 , \4025_b1 );
xor ( \4026_b0 , \4023_b0 , w_12834 );
not ( w_12834 , w_12835 );
and ( w_12835 , \4025_b1 , \4025_b0 );
or ( \4027_b1 , \3960_b1 , \3966_b1 );
not ( \3966_b1 , w_12836 );
and ( \4027_b0 , \3960_b0 , w_12837 );
and ( w_12836 , w_12837 , \3966_b0 );
or ( \4028_b1 , \4027_b1 , w_12839 );
not ( w_12839 , w_12840 );
and ( \4028_b0 , \4027_b0 , w_12841 );
and ( w_12840 ,  , w_12841 );
buf ( w_12839 , \3980_b1 );
not ( w_12839 , w_12842 );
not (  , w_12843 );
and ( w_12842 , w_12843 , \3980_b0 );
buf ( \4029_b1 , \3972_b1 );
not ( \4029_b1 , w_12844 );
not ( \4029_b0 , w_12845 );
and ( w_12844 , w_12845 , \3972_b0 );
or ( \4031_b1 , \3986_b1 , w_12846 );
or ( \4031_b0 , \3986_b0 , \3972_b0 );
not ( \3972_b0 , w_12847 );
and ( w_12847 , w_12846 , \3972_b1 );
or ( \4032_b1 , \4031_b1 , w_12849 );
not ( w_12849 , w_12850 );
and ( \4032_b0 , \4031_b0 , w_12851 );
and ( w_12850 ,  , w_12851 );
buf ( w_12849 , \3988_b1 );
not ( w_12849 , w_12852 );
not (  , w_12853 );
and ( w_12852 , w_12853 , \3988_b0 );
or ( \4033_b1 , \4030_b1 , w_12855 );
not ( w_12855 , w_12856 );
and ( \4033_b0 , \4030_b0 , w_12857 );
and ( w_12856 ,  , w_12857 );
buf ( w_12855 , \4032_b1 );
not ( w_12855 , w_12858 );
not (  , w_12859 );
and ( w_12858 , w_12859 , \4032_b0 );
buf ( \4035_b1 , \3991_b1 );
not ( \4035_b1 , w_12860 );
not ( \4035_b0 , w_12861 );
and ( w_12860 , w_12861 , \3991_b0 );
buf ( \4036_b1 , \3986_b1 );
not ( \4036_b1 , w_12862 );
not ( \4036_b0 , w_12863 );
and ( w_12862 , w_12863 , \3986_b0 );
or ( \4037_b1 , \4036_b1 , w_12865 );
not ( w_12865 , w_12866 );
and ( \4037_b0 , \4036_b0 , w_12867 );
and ( w_12866 ,  , w_12867 );
buf ( w_12865 , \3973_b1 );
not ( w_12865 , w_12868 );
not (  , w_12869 );
and ( w_12868 , w_12869 , \3973_b0 );
or ( \4038_b1 , \4035_b1 , w_12871 );
not ( w_12871 , w_12872 );
and ( \4038_b0 , \4035_b0 , w_12873 );
and ( w_12872 ,  , w_12873 );
buf ( w_12871 , \4037_b1 );
not ( w_12871 , w_12874 );
not (  , w_12875 );
and ( w_12874 , w_12875 , \4037_b0 );
or ( \4039_b1 , \4034_b1 , w_12877 );
not ( w_12877 , w_12878 );
and ( \4039_b0 , \4034_b0 , w_12879 );
and ( w_12878 ,  , w_12879 );
buf ( w_12877 , \4038_b1 );
not ( w_12877 , w_12880 );
not (  , w_12881 );
and ( w_12880 , w_12881 , \4038_b0 );
buf ( \4040_b1 , \3960_b1 );
not ( \4040_b1 , w_12882 );
not ( \4040_b0 , w_12883 );
and ( w_12882 , w_12883 , \3960_b0 );
or ( \4041_b1 , \4040_b1 , w_12884 );
or ( \4041_b0 , \4040_b0 , \3965_b0 );
not ( \3965_b0 , w_12885 );
and ( w_12885 , w_12884 , \3965_b1 );
or ( \4042_b1 , \4041_b1 , w_12887 );
not ( w_12887 , w_12888 );
and ( \4042_b0 , \4041_b0 , w_12889 );
and ( w_12888 ,  , w_12889 );
buf ( w_12887 , \3977_b1 );
not ( w_12887 , w_12890 );
not (  , w_12891 );
and ( w_12890 , w_12891 , \3977_b0 );
or ( \4043_b1 , \3969_b1 , w_12893 );
not ( w_12893 , w_12894 );
and ( \4043_b0 , \3969_b0 , w_12895 );
and ( w_12894 ,  , w_12895 );
buf ( w_12893 , \3927_b1 );
not ( w_12893 , w_12896 );
not (  , w_12897 );
and ( w_12896 , w_12897 , \3927_b0 );
or ( \4044_b1 , \4043_b1 , w_12899 );
not ( w_12899 , w_12900 );
and ( \4044_b0 , \4043_b0 , w_12901 );
and ( w_12900 ,  , w_12901 );
buf ( w_12899 , \3973_b1 );
not ( w_12899 , w_12902 );
not (  , w_12903 );
and ( w_12902 , w_12903 , \3973_b0 );
or ( \4046_b1 , \3991_b1 , \4043_b1 );
not ( \4043_b1 , w_12904 );
and ( \4046_b0 , \3991_b0 , w_12905 );
and ( w_12904 , w_12905 , \4043_b0 );
or ( \4047_b1 , \3986_b1 , w_12907 );
not ( w_12907 , w_12908 );
and ( \4047_b0 , \3986_b0 , w_12909 );
and ( w_12908 ,  , w_12909 );
buf ( w_12907 , \4044_b1 );
not ( w_12907 , w_12910 );
not (  , w_12911 );
and ( w_12910 , w_12911 , \4044_b0 );
or ( \4048_b1 , \3927_b1 , w_12912 );
or ( \4048_b0 , \3927_b0 , \3994_b0 );
not ( \3994_b0 , w_12913 );
and ( w_12913 , w_12912 , \3994_b1 );
or ( \4049_b1 , \4048_b1 , w_12915 );
not ( w_12915 , w_12916 );
and ( \4049_b0 , \4048_b0 , w_12917 );
and ( w_12916 ,  , w_12917 );
buf ( w_12915 , \3929_b1 );
not ( w_12915 , w_12918 );
not (  , w_12919 );
and ( w_12918 , w_12919 , \3929_b0 );
or ( \4051_b1 , \4045_b1 , w_12921 );
not ( w_12921 , w_12922 );
and ( \4051_b0 , \4045_b0 , w_12923 );
and ( w_12922 ,  , w_12923 );
buf ( w_12921 , \4050_b1 );
not ( w_12921 , w_12924 );
not (  , w_12925 );
and ( w_12924 , w_12925 , \4050_b0 );
buf ( \4052_b1 , \3962_b1 );
not ( \4052_b1 , w_12926 );
not ( \4052_b0 , w_12927 );
and ( w_12926 , w_12927 , \3962_b0 );
buf ( \4054_b1 , \4052_b1 );
not ( \4054_b1 , w_12928 );
not ( \4054_b0 , w_12929 );
and ( w_12928 , w_12929 , \4052_b0 );
buf ( \4055_b1 , \3980_b1 );
not ( \4055_b1 , w_12930 );
not ( \4055_b0 , w_12931 );
and ( w_12930 , w_12931 , \3980_b0 );
or ( \4056_b1 , \4054_b1 , w_12932 );
or ( \4056_b0 , \4054_b0 , \4055_b0 );
not ( \4055_b0 , w_12933 );
and ( w_12933 , w_12932 , \4055_b1 );
or ( \4057_b1 , \4056_b1 , w_12935 );
not ( w_12935 , w_12936 );
and ( \4057_b0 , \4056_b0 , w_12937 );
and ( w_12936 ,  , w_12937 );
buf ( w_12935 , \3982_b1 );
not ( w_12935 , w_12938 );
not (  , w_12939 );
and ( w_12938 , w_12939 , \3982_b0 );
or ( \4058_b1 , \4053_b1 , w_12941 );
not ( w_12941 , w_12942 );
and ( \4058_b0 , \4053_b0 , w_12943 );
and ( w_12942 ,  , w_12943 );
buf ( w_12941 , \4057_b1 );
not ( w_12941 , w_12944 );
not (  , w_12945 );
and ( w_12944 , w_12945 , \4057_b0 );
or ( \4059_b1 , \4040_b1 , w_12946 );
or ( \4059_b0 , \4040_b0 , \3967_b0 );
not ( \3967_b0 , w_12947 );
and ( w_12947 , w_12946 , \3967_b1 );
or ( \4060_b1 , \4059_b1 , w_12949 );
not ( w_12949 , w_12950 );
and ( \4060_b0 , \4059_b0 , w_12951 );
and ( w_12950 ,  , w_12951 );
buf ( w_12949 , \3986_b1 );
not ( w_12949 , w_12952 );
not (  , w_12953 );
and ( w_12952 , w_12953 , \3986_b0 );
buf ( \4061_b1 , \3965_b1 );
not ( \4061_b1 , w_12954 );
not ( \4061_b0 , w_12955 );
and ( w_12954 , w_12955 , \3965_b0 );
or ( \4062_b1 , \4061_b1 , w_12957 );
not ( w_12957 , w_12958 );
and ( \4062_b0 , \4061_b0 , w_12959 );
and ( w_12958 ,  , w_12959 );
buf ( w_12957 , \3977_b1 );
not ( w_12957 , w_12960 );
not (  , w_12961 );
and ( w_12960 , w_12961 , \3977_b0 );
or ( \4063_b1 , \4062_b1 , \3960_b1 );
not ( \3960_b1 , w_12962 );
and ( \4063_b0 , \4062_b0 , w_12963 );
and ( w_12962 , w_12963 , \3960_b0 );
buf ( \4064_b1 , \4062_b1 );
not ( \4064_b1 , w_12964 );
not ( \4064_b0 , w_12965 );
and ( w_12964 , w_12965 , \4062_b0 );
or ( \4065_b1 , \4064_b1 , \4040_b1 );
not ( \4040_b1 , w_12966 );
and ( \4065_b0 , \4064_b0 , w_12967 );
and ( w_12966 , w_12967 , \4040_b0 );
or ( \4066_b1 , \4063_b1 , w_12968 );
or ( \4066_b0 , \4063_b0 , \4065_b0 );
not ( \4065_b0 , w_12969 );
and ( w_12969 , w_12968 , \4065_b1 );
buf ( \4067_b1 , \3942_b1 );
not ( \4067_b1 , w_12970 );
not ( \4067_b0 , w_12971 );
and ( w_12970 , w_12971 , \3942_b0 );
or ( \4068_b1 , \4067_b1 , w_12973 );
not ( w_12973 , w_12974 );
and ( \4068_b0 , \4067_b0 , w_12975 );
and ( w_12974 ,  , w_12975 );
buf ( w_12973 , \3950_b1 );
not ( w_12973 , w_12976 );
not (  , w_12977 );
and ( w_12976 , w_12977 , \3950_b0 );
or ( \4069_b1 , \4068_b1 , \4007_b1 );
not ( \4007_b1 , w_12978 );
and ( \4069_b0 , \4068_b0 , w_12979 );
and ( w_12978 , w_12979 , \4007_b0 );
buf ( \4070_b1 , \4068_b1 );
not ( \4070_b1 , w_12980 );
not ( \4070_b0 , w_12981 );
and ( w_12980 , w_12981 , \4068_b0 );
or ( \4071_b1 , \4070_b1 , \4006_b1 );
not ( \4006_b1 , w_12982 );
and ( \4071_b0 , \4070_b0 , w_12983 );
and ( w_12982 , w_12983 , \4006_b0 );
or ( \4072_b1 , \4069_b1 , w_12984 );
or ( \4072_b0 , \4069_b0 , \4071_b0 );
not ( \4071_b0 , w_12985 );
and ( w_12985 , w_12984 , \4071_b1 );
or ( \4073_b1 , \3948_b1 , w_12987 );
not ( w_12987 , w_12988 );
and ( \4073_b0 , \3948_b0 , w_12989 );
and ( w_12988 ,  , w_12989 );
buf ( w_12987 , \3938_b1 );
not ( w_12987 , w_12990 );
not (  , w_12991 );
and ( w_12990 , w_12991 , \3938_b0 );
buf ( \4074_b1 , \3939_b1 );
not ( \4074_b1 , w_12992 );
not ( \4074_b0 , w_12993 );
and ( w_12992 , w_12993 , \3939_b0 );
or ( \4075_b1 , \4074_b1 , w_12995 );
not ( w_12995 , w_12996 );
and ( \4075_b0 , \4074_b0 , w_12997 );
and ( w_12996 ,  , w_12997 );
buf ( w_12995 , \3936_b1 );
not ( w_12995 , w_12998 );
not (  , w_12999 );
and ( w_12998 , w_12999 , \3936_b0 );
or ( \4076_b1 , \4073_b1 , \4075_b1 );
xor ( \4076_b0 , \4073_b0 , w_13000 );
not ( w_13000 , w_13001 );
and ( w_13001 , \4075_b1 , \4075_b0 );
buf ( \4077_b1 , \3939_b1 );
not ( \4077_b1 , w_13002 );
not ( \4077_b0 , w_13003 );
and ( w_13002 , w_13003 , \3939_b0 );
or ( \4078_b1 , \4077_b1 , w_13005 );
not ( w_13005 , w_13006 );
and ( \4078_b0 , \4077_b0 , w_13007 );
and ( w_13006 ,  , w_13007 );
buf ( w_13005 , \3935_b1 );
not ( w_13005 , w_13008 );
not (  , w_13009 );
and ( w_13008 , w_13009 , \3935_b0 );
or ( \4079_b1 , \4078_b1 , \4001_b1 );
xor ( \4079_b0 , \4078_b0 , w_13010 );
not ( w_13010 , w_13011 );
and ( w_13011 , \4001_b1 , \4001_b0 );
buf ( \4080_b1 , \3934_b1 );
not ( \4080_b1 , w_13012 );
not ( \4080_b0 , w_13013 );
and ( w_13012 , w_13013 , \3934_b0 );
or ( \4081_b1 , \4080_b1 , w_13015 );
not ( w_13015 , w_13016 );
and ( \4081_b0 , \4080_b0 , w_13017 );
and ( w_13016 ,  , w_13017 );
buf ( w_13015 , \3931_b1 );
not ( w_13015 , w_13018 );
not (  , w_13019 );
and ( w_13018 , w_13019 , \3931_b0 );
or ( \4082_b1 , \3932_b1 , \4081_b1 );
xor ( \4082_b0 , \3932_b0 , w_13020 );
not ( w_13020 , w_13021 );
and ( w_13021 , \4081_b1 , \4081_b0 );
or ( \4083_b1 , \4029_b1 , w_13023 );
not ( w_13023 , w_13024 );
and ( \4083_b0 , \4029_b0 , w_13025 );
and ( w_13024 ,  , w_13025 );
buf ( w_13023 , \3988_b1 );
not ( w_13023 , w_13026 );
not (  , w_13027 );
and ( w_13026 , w_13027 , \3988_b0 );
buf ( \4084_b1 , \3961_b1 );
not ( \4084_b1 , w_13028 );
not ( \4084_b0 , w_13029 );
and ( w_13028 , w_13029 , \3961_b0 );
or ( \4085_b1 , \4084_b1 , w_13031 );
not ( w_13031 , w_13032 );
and ( \4085_b0 , \4084_b0 , w_13033 );
and ( w_13032 ,  , w_13033 );
buf ( w_13031 , \3984_b1 );
not ( w_13031 , w_13034 );
not (  , w_13035 );
and ( w_13034 , w_13035 , \3984_b0 );
or ( \4086_b1 , \4052_b1 , w_13037 );
not ( w_13037 , w_13038 );
and ( \4086_b0 , \4052_b0 , w_13039 );
and ( w_13038 ,  , w_13039 );
buf ( w_13037 , \3982_b1 );
not ( w_13037 , w_13040 );
not (  , w_13041 );
and ( w_13040 , w_13041 , \3982_b0 );
buf ( \4087_b1 , \3979_b1 );
not ( \4087_b1 , w_13042 );
not ( \4087_b0 , w_13043 );
and ( w_13042 , w_13043 , \3979_b0 );
or ( \4088_b1 , \4087_b1 , w_13045 );
not ( w_13045 , w_13046 );
and ( \4088_b0 , \4087_b0 , w_13047 );
and ( w_13046 ,  , w_13047 );
buf ( w_13045 , \3964_b1 );
not ( w_13045 , w_13048 );
not (  , w_13049 );
and ( w_13048 , w_13049 , \3964_b0 );
buf ( \4089_b1 , \3969_b1 );
not ( \4089_b1 , w_13050 );
not ( \4089_b0 , w_13051 );
and ( w_13050 , w_13051 , \3969_b0 );
or ( \4090_b1 , \4089_b1 , w_13053 );
not ( w_13053 , w_13054 );
and ( \4090_b0 , \4089_b0 , w_13055 );
and ( w_13054 ,  , w_13055 );
buf ( w_13053 , \3994_b1 );
not ( w_13053 , w_13056 );
not (  , w_13057 );
and ( w_13056 , w_13057 , \3994_b0 );
buf ( \4091_b1 , \3971_b1 );
not ( \4091_b1 , w_13058 );
not ( \4091_b0 , w_13059 );
and ( w_13058 , w_13059 , \3971_b0 );
or ( \4092_b1 , \4091_b1 , w_13061 );
not ( w_13061 , w_13062 );
and ( \4092_b0 , \4091_b0 , w_13063 );
and ( w_13062 ,  , w_13063 );
buf ( w_13061 , \3990_b1 );
not ( w_13061 , w_13064 );
not (  , w_13065 );
and ( w_13064 , w_13065 , \3990_b0 );
or ( \4093_b1 , \4086_b1 , \4028_b1 );
xor ( \4093_b0 , \4086_b0 , w_13066 );
not ( w_13066 , w_13067 );
and ( w_13067 , \4028_b1 , \4028_b0 );
or ( \4094_b1 , \4092_b1 , \4033_b1 );
xor ( \4094_b0 , \4092_b0 , w_13068 );
not ( w_13068 , w_13069 );
and ( w_13069 , \4033_b1 , \4033_b0 );
or ( \4095_b1 , \4088_b1 , \4042_b1 );
xor ( \4095_b0 , \4088_b0 , w_13070 );
not ( w_13070 , w_13071 );
and ( w_13071 , \4042_b1 , \4042_b0 );
or ( \4096_b1 , \4060_b1 , w_13072 );
xor ( \4096_b0 , \4060_b0 , w_13074 );
not ( w_13074 , w_13075 );
and ( w_13075 , w_13072 , w_13073 );
buf ( w_13072 , \4083_b1 );
not ( w_13072 , w_13076 );
not ( w_13073 , w_13077 );
and ( w_13076 , w_13077 , \4083_b0 );
or ( \4097_b1 , \4058_b1 , \4085_b1 );
xor ( \4097_b0 , \4058_b0 , w_13078 );
not ( w_13078 , w_13079 );
and ( w_13079 , \4085_b1 , \4085_b0 );
or ( \4098_b1 , \d[0]_b1 , \c[0]_b1 );
xor ( \4098_b0 , \d[0]_b0 , w_13080 );
not ( w_13080 , w_13081 );
and ( w_13081 , \c[0]_b1 , \c[0]_b0 );
buf ( \4100_b1 , \4099_b1 );
buf ( \4100_b0 , \4099_b0 );
buf ( \4101_b1 , \4100_b1 );
not ( \4101_b1 , w_13082 );
not ( \4101_b0 , w_13083 );
and ( w_13082 , w_13083 , \4100_b0 );
buf ( \4102_b1 , \4101_b1 );
not ( \4102_b1 , w_13084 );
not ( \4102_b0 , w_13085 );
and ( w_13084 , w_13085 , \4101_b0 );
or ( \4103_b1 , \4102_b1 , \4096_b1 );
not ( \4096_b1 , w_13086 );
and ( \4103_b0 , \4102_b0 , w_13087 );
and ( w_13086 , w_13087 , \4096_b0 );
buf ( \4104_b1 , \3997_b1 );
not ( \4104_b1 , w_13088 );
not ( \4104_b0 , w_13089 );
and ( w_13088 , w_13089 , \3997_b0 );
buf ( \4105_b1 , \2477_b1 );
buf ( \4105_b0 , \2477_b0 );
buf ( \4106_b1 , \4105_b1 );
buf ( \4106_b0 , \4105_b0 );
buf ( \4107_b1 , \4106_b1 );
not ( \4107_b1 , w_13090 );
not ( \4107_b0 , w_13091 );
and ( w_13090 , w_13091 , \4106_b0 );
buf ( \4108_b1 , \4107_b1 );
not ( \4108_b1 , w_13092 );
not ( \4108_b0 , w_13093 );
and ( w_13092 , w_13093 , \4107_b0 );
or ( \4109_b1 , \4104_b1 , w_13094 );
or ( \4109_b0 , \4104_b0 , \4108_b0 );
not ( \4108_b0 , w_13095 );
and ( w_13095 , w_13094 , \4108_b1 );
buf ( \4110_b1 , \4105_b1 );
buf ( \4110_b0 , \4105_b0 );
buf ( \4111_b1 , \3997_b1 );
not ( \4111_b1 , w_13096 );
not ( \4111_b0 , w_13097 );
and ( w_13096 , w_13097 , \3997_b0 );
or ( \4112_b1 , \4110_b1 , w_13099 );
not ( w_13099 , w_13100 );
and ( \4112_b0 , \4110_b0 , w_13101 );
and ( w_13100 ,  , w_13101 );
buf ( w_13099 , \4111_b1 );
not ( w_13099 , w_13102 );
not (  , w_13103 );
and ( w_13102 , w_13103 , \4111_b0 );
or ( \4113_b1 , \4109_b1 , w_13105 );
not ( w_13105 , w_13106 );
and ( \4113_b0 , \4109_b0 , w_13107 );
and ( w_13106 ,  , w_13107 );
buf ( w_13105 , \4112_b1 );
not ( w_13105 , w_13108 );
not (  , w_13109 );
and ( w_13108 , w_13109 , \4112_b0 );
buf ( \4114_b1 , \4113_b1 );
not ( \4114_b1 , w_13110 );
not ( \4114_b0 , w_13111 );
and ( w_13110 , w_13111 , \4113_b0 );
or ( \4115_b1 , \3193_b1 , w_13113 );
not ( w_13113 , w_13114 );
and ( \4115_b0 , \3193_b0 , w_13115 );
and ( w_13114 ,  , w_13115 );
buf ( w_13113 , \3656_b1 );
not ( w_13113 , w_13116 );
not (  , w_13117 );
and ( w_13116 , w_13117 , \3656_b0 );
buf ( \4116_b1 , \4115_b1 );
not ( \4116_b1 , w_13118 );
not ( \4116_b0 , w_13119 );
and ( w_13118 , w_13119 , \4115_b0 );
buf ( \4117_b1 , \4116_b1 );
not ( \4117_b1 , w_13120 );
not ( \4117_b0 , w_13121 );
and ( w_13120 , w_13121 , \4116_b0 );
buf ( \4118_b1 , \4105_b1 );
not ( \4118_b1 , w_13122 );
not ( \4118_b0 , w_13123 );
and ( w_13122 , w_13123 , \4105_b0 );
or ( \4119_b1 , \4117_b1 , w_13124 );
or ( \4119_b0 , \4117_b0 , \4118_b0 );
not ( \4118_b0 , w_13125 );
and ( w_13125 , w_13124 , \4118_b1 );
buf ( \4120_b1 , \3656_b1 );
not ( \4120_b1 , w_13126 );
not ( \4120_b0 , w_13127 );
and ( w_13126 , w_13127 , \3656_b0 );
buf ( \4121_b1 , \3193_b1 );
not ( \4121_b1 , w_13128 );
not ( \4121_b0 , w_13129 );
and ( w_13128 , w_13129 , \3193_b0 );
or ( \4122_b1 , \4120_b1 , w_13130 );
or ( \4122_b0 , \4120_b0 , \4121_b0 );
not ( \4121_b0 , w_13131 );
and ( w_13131 , w_13130 , \4121_b1 );
buf ( \4123_b1 , \4105_b1 );
not ( \4123_b1 , w_13132 );
not ( \4123_b0 , w_13133 );
and ( w_13132 , w_13133 , \4105_b0 );
or ( \4124_b1 , \4122_b1 , w_13135 );
not ( w_13135 , w_13136 );
and ( \4124_b0 , \4122_b0 , w_13137 );
and ( w_13136 ,  , w_13137 );
buf ( w_13135 , \4123_b1 );
not ( w_13135 , w_13138 );
not (  , w_13139 );
and ( w_13138 , w_13139 , \4123_b0 );
or ( \4125_b1 , \4119_b1 , w_13141 );
not ( w_13141 , w_13142 );
and ( \4125_b0 , \4119_b0 , w_13143 );
and ( w_13142 ,  , w_13143 );
buf ( w_13141 , \4124_b1 );
not ( w_13141 , w_13144 );
not (  , w_13145 );
and ( w_13144 , w_13145 , \4124_b0 );
or ( \4126_b1 , \2876_b1 , w_13146 );
xor ( \4126_b0 , \2876_b0 , w_13148 );
not ( w_13148 , w_13149 );
and ( w_13149 , w_13146 , w_13147 );
buf ( w_13146 , \4115_b1 );
not ( w_13146 , w_13150 );
not ( w_13147 , w_13151 );
and ( w_13150 , w_13151 , \4115_b0 );
or ( \4127_b1 , \4125_b1 , w_13153 );
not ( w_13153 , w_13154 );
and ( \4127_b0 , \4125_b0 , w_13155 );
and ( w_13154 ,  , w_13155 );
buf ( w_13153 , \4126_b1 );
not ( w_13153 , w_13156 );
not (  , w_13157 );
and ( w_13156 , w_13157 , \4126_b0 );
buf ( \4128_b1 , \4127_b1 );
not ( \4128_b1 , w_13158 );
not ( \4128_b0 , w_13159 );
and ( w_13158 , w_13159 , \4127_b0 );
buf ( \4129_b1 , \4128_b1 );
buf ( \4129_b0 , \4128_b0 );
buf ( \4130_b1 , \4129_b1 );
not ( \4130_b1 , w_13160 );
not ( \4130_b0 , w_13161 );
and ( w_13160 , w_13161 , \4129_b0 );
or ( \4131_b1 , \4114_b1 , w_13162 );
or ( \4131_b0 , \4114_b0 , \4130_b0 );
not ( \4130_b0 , w_13163 );
and ( w_13163 , w_13162 , \4130_b1 );
buf ( \4132_b1 , \4126_b1 );
not ( \4132_b1 , w_13164 );
not ( \4132_b0 , w_13165 );
and ( w_13164 , w_13165 , \4126_b0 );
buf ( \4133_b1 , \4132_b1 );
buf ( \4133_b0 , \4132_b0 );
buf ( \4134_b1 , \4110_b1 );
not ( \4134_b1 , w_13166 );
not ( \4134_b0 , w_13167 );
and ( w_13166 , w_13167 , \4110_b0 );
buf ( \4135_b1 , \4051_b1 );
not ( \4135_b1 , w_13168 );
not ( \4135_b0 , w_13169 );
and ( w_13168 , w_13169 , \4051_b0 );
or ( \4136_b1 , \4134_b1 , \4135_b1 );
not ( \4135_b1 , w_13170 );
and ( \4136_b0 , \4134_b0 , w_13171 );
and ( w_13170 , w_13171 , \4135_b0 );
buf ( \4137_b1 , \4134_b1 );
not ( \4137_b1 , w_13172 );
not ( \4137_b0 , w_13173 );
and ( w_13172 , w_13173 , \4134_b0 );
or ( \4138_b1 , \4137_b1 , \4051_b1 );
not ( \4051_b1 , w_13174 );
and ( \4138_b0 , \4137_b0 , w_13175 );
and ( w_13174 , w_13175 , \4051_b0 );
or ( \4139_b1 , \4136_b1 , w_13177 );
not ( w_13177 , w_13178 );
and ( \4139_b0 , \4136_b0 , w_13179 );
and ( w_13178 ,  , w_13179 );
buf ( w_13177 , \4138_b1 );
not ( w_13177 , w_13180 );
not (  , w_13181 );
and ( w_13180 , w_13181 , \4138_b0 );
or ( \4140_b1 , \4133_b1 , w_13183 );
not ( w_13183 , w_13184 );
and ( \4140_b0 , \4133_b0 , w_13185 );
and ( w_13184 ,  , w_13185 );
buf ( w_13183 , \4139_b1 );
not ( w_13183 , w_13186 );
not (  , w_13187 );
and ( w_13186 , w_13187 , \4139_b0 );
or ( \4141_b1 , \4131_b1 , w_13189 );
not ( w_13189 , w_13190 );
and ( \4141_b0 , \4131_b0 , w_13191 );
and ( w_13190 ,  , w_13191 );
buf ( w_13189 , \4140_b1 );
not ( w_13189 , w_13192 );
not (  , w_13193 );
and ( w_13192 , w_13193 , \4140_b0 );
or ( \4142_b1 , \4103_b1 , \4141_b1 );
xor ( \4142_b0 , \4103_b0 , w_13194 );
not ( w_13194 , w_13195 );
and ( w_13195 , \4141_b1 , \4141_b0 );
buf ( \4143_b1 , \3637_b1 );
not ( \4143_b1 , w_13196 );
not ( \4143_b0 , w_13197 );
and ( w_13196 , w_13197 , \3637_b0 );
buf ( \4144_b1 , \4143_b1 );
not ( \4144_b1 , w_13198 );
not ( \4144_b0 , w_13199 );
and ( w_13198 , w_13199 , \4143_b0 );
buf ( \4145_b1 , \3573_b1 );
not ( \4145_b1 , w_13200 );
not ( \4145_b0 , w_13201 );
and ( w_13200 , w_13201 , \3573_b0 );
or ( \4146_b1 , \4144_b1 , w_13202 );
or ( \4146_b0 , \4144_b0 , \4145_b0 );
not ( \4145_b0 , w_13203 );
and ( w_13203 , w_13202 , \4145_b1 );
buf ( \4147_b1 , \3573_b1 );
not ( \4147_b1 , w_13204 );
not ( \4147_b0 , w_13205 );
and ( w_13204 , w_13205 , \3573_b0 );
or ( \4148_b1 , \4147_b1 , w_13207 );
not ( w_13207 , w_13208 );
and ( \4148_b0 , \4147_b0 , w_13209 );
and ( w_13208 ,  , w_13209 );
buf ( w_13207 , \3637_b1 );
not ( w_13207 , w_13210 );
not (  , w_13211 );
and ( w_13210 , w_13211 , \3637_b0 );
or ( \4149_b1 , \4146_b1 , w_13213 );
not ( w_13213 , w_13214 );
and ( \4149_b0 , \4146_b0 , w_13215 );
and ( w_13214 ,  , w_13215 );
buf ( w_13213 , \4148_b1 );
not ( w_13213 , w_13216 );
not (  , w_13217 );
and ( w_13216 , w_13217 , \4148_b0 );
buf ( \4150_b1 , \4149_b1 );
buf ( \4150_b0 , \4149_b0 );
buf ( \4151_b1 , \4150_b1 );
not ( \4151_b1 , w_13218 );
not ( \4151_b0 , w_13219 );
and ( w_13218 , w_13219 , \4150_b0 );
buf ( \4152_b1 , \4151_b1 );
not ( \4152_b1 , w_13220 );
not ( \4152_b0 , w_13221 );
and ( w_13220 , w_13221 , \4151_b0 );
buf ( \4153_b1 , \2876_b1 );
not ( \4153_b1 , w_13222 );
not ( \4153_b0 , w_13223 );
and ( w_13222 , w_13223 , \2876_b0 );
buf ( \4154_b1 , \4153_b1 );
not ( \4154_b1 , w_13224 );
not ( \4154_b0 , w_13225 );
and ( w_13224 , w_13225 , \4153_b0 );
or ( \4155_b1 , \4154_b1 , \4147_b1 );
not ( \4147_b1 , w_13226 );
and ( \4155_b0 , \4154_b0 , w_13227 );
and ( w_13226 , w_13227 , \4147_b0 );
or ( \4156_b1 , \4153_b1 , \3573_b1 );
not ( \3573_b1 , w_13228 );
and ( \4156_b0 , \4153_b0 , w_13229 );
and ( w_13228 , w_13229 , \3573_b0 );
or ( \4157_b1 , \4155_b1 , w_13231 );
not ( w_13231 , w_13232 );
and ( \4157_b0 , \4155_b0 , w_13233 );
and ( w_13232 ,  , w_13233 );
buf ( w_13231 , \4156_b1 );
not ( w_13231 , w_13234 );
not (  , w_13235 );
and ( w_13234 , w_13235 , \4156_b0 );
or ( \4158_b1 , \4157_b1 , w_13237 );
not ( w_13237 , w_13238 );
and ( \4158_b0 , \4157_b0 , w_13239 );
and ( w_13238 ,  , w_13239 );
buf ( w_13237 , \4149_b1 );
not ( w_13237 , w_13240 );
not (  , w_13241 );
and ( w_13240 , w_13241 , \4149_b0 );
buf ( \4159_b1 , \4158_b1 );
buf ( \4159_b0 , \4158_b0 );
buf ( \4160_b1 , \4159_b1 );
not ( \4160_b1 , w_13242 );
not ( \4160_b0 , w_13243 );
and ( w_13242 , w_13243 , \4159_b0 );
buf ( \4161_b1 , \4160_b1 );
not ( \4161_b1 , w_13244 );
not ( \4161_b0 , w_13245 );
and ( w_13244 , w_13245 , \4160_b0 );
or ( \4162_b1 , \4152_b1 , w_13246 );
or ( \4162_b0 , \4152_b0 , \4161_b0 );
not ( \4161_b0 , w_13247 );
and ( w_13247 , w_13246 , \4161_b1 );
buf ( \4163_b1 , \4153_b1 );
buf ( \4163_b0 , \4153_b0 );
buf ( \4164_b1 , \4163_b1 );
not ( \4164_b1 , w_13248 );
not ( \4164_b0 , w_13249 );
and ( w_13248 , w_13249 , \4163_b0 );
or ( \4165_b1 , \4162_b1 , w_13251 );
not ( w_13251 , w_13252 );
and ( \4165_b0 , \4162_b0 , w_13253 );
and ( w_13252 ,  , w_13253 );
buf ( w_13251 , \4164_b1 );
not ( w_13251 , w_13254 );
not (  , w_13255 );
and ( w_13254 , w_13255 , \4164_b0 );
or ( \4166_b1 , \4142_b1 , \4165_b1 );
xor ( \4166_b0 , \4142_b0 , w_13256 );
not ( w_13256 , w_13257 );
and ( w_13257 , \4165_b1 , \4165_b0 );
buf ( \4167_b1 , \4051_b1 );
not ( \4167_b1 , w_13258 );
not ( \4167_b0 , w_13259 );
and ( w_13258 , w_13259 , \4051_b0 );
buf ( \4168_b1 , \4163_b1 );
not ( \4168_b1 , w_13260 );
not ( \4168_b0 , w_13261 );
and ( w_13260 , w_13261 , \4163_b0 );
or ( \4169_b1 , \4167_b1 , w_13262 );
or ( \4169_b0 , \4167_b0 , \4168_b0 );
not ( \4168_b0 , w_13263 );
and ( w_13263 , w_13262 , \4168_b1 );
buf ( \4170_b1 , \4163_b1 );
not ( \4170_b1 , w_13264 );
not ( \4170_b0 , w_13265 );
and ( w_13264 , w_13265 , \4163_b0 );
or ( \4171_b1 , \4135_b1 , w_13267 );
not ( w_13267 , w_13268 );
and ( \4171_b0 , \4135_b0 , w_13269 );
and ( w_13268 ,  , w_13269 );
buf ( w_13267 , \4170_b1 );
not ( w_13267 , w_13270 );
not (  , w_13271 );
and ( w_13270 , w_13271 , \4170_b0 );
or ( \4172_b1 , \4169_b1 , w_13273 );
not ( w_13273 , w_13274 );
and ( \4172_b0 , \4169_b0 , w_13275 );
and ( w_13274 ,  , w_13275 );
buf ( w_13273 , \4171_b1 );
not ( w_13273 , w_13276 );
not (  , w_13277 );
and ( w_13276 , w_13277 , \4171_b0 );
buf ( \4173_b1 , \4172_b1 );
not ( \4173_b1 , w_13278 );
not ( \4173_b0 , w_13279 );
and ( w_13278 , w_13279 , \4172_b0 );
buf ( \4174_b1 , \4159_b1 );
not ( \4174_b1 , w_13280 );
not ( \4174_b0 , w_13281 );
and ( w_13280 , w_13281 , \4159_b0 );
or ( \4175_b1 , \4173_b1 , w_13282 );
or ( \4175_b0 , \4173_b0 , \4174_b0 );
not ( \4174_b0 , w_13283 );
and ( w_13283 , w_13282 , \4174_b1 );
or ( \4176_b1 , \4150_b1 , w_13285 );
not ( w_13285 , w_13286 );
and ( \4176_b0 , \4150_b0 , w_13287 );
and ( w_13286 ,  , w_13287 );
buf ( w_13285 , \4164_b1 );
not ( w_13285 , w_13288 );
not (  , w_13289 );
and ( w_13288 , w_13289 , \4164_b0 );
or ( \4177_b1 , \4175_b1 , w_13291 );
not ( w_13291 , w_13292 );
and ( \4177_b0 , \4175_b0 , w_13293 );
and ( w_13292 ,  , w_13293 );
buf ( w_13291 , \4176_b1 );
not ( w_13291 , w_13294 );
not (  , w_13295 );
and ( w_13294 , w_13295 , \4176_b0 );
or ( \4178_b1 , \4094_b1 , \4100_b1 );
xor ( \4178_b0 , \4094_b0 , w_13296 );
not ( w_13296 , w_13297 );
and ( w_13297 , \4100_b1 , \4100_b0 );
buf ( \4179_b1 , \4178_b1 );
not ( \4179_b1 , w_13298 );
not ( \4179_b0 , w_13299 );
and ( w_13298 , w_13299 , \4178_b0 );
buf ( \4180_b1 , \2790_b1 );
not ( \4180_b1 , w_13300 );
not ( \4180_b0 , w_13301 );
and ( w_13300 , w_13301 , \2790_b0 );
buf ( \4181_b1 , \4180_b1 );
not ( \4181_b1 , w_13302 );
not ( \4181_b0 , w_13303 );
and ( w_13302 , w_13303 , \4180_b0 );
buf ( \4182_b1 , \4181_b1 );
not ( \4182_b1 , w_13304 );
not ( \4182_b0 , w_13305 );
and ( w_13304 , w_13305 , \4181_b0 );
or ( \4183_b1 , \4099_b1 , w_13307 );
not ( w_13307 , w_13308 );
and ( \4183_b0 , \4099_b0 , w_13309 );
and ( w_13308 ,  , w_13309 );
buf ( w_13307 , \4182_b1 );
not ( w_13307 , w_13310 );
not (  , w_13311 );
and ( w_13310 , w_13311 , \4182_b0 );
buf ( \4184_b1 , \4183_b1 );
not ( \4184_b1 , w_13312 );
not ( \4184_b0 , w_13313 );
and ( w_13312 , w_13313 , \4183_b0 );
or ( \4186_b1 , \4181_b1 , w_13315 );
not ( w_13315 , w_13316 );
and ( \4186_b0 , \4181_b0 , w_13317 );
and ( w_13316 ,  , w_13317 );
buf ( w_13315 , \4185_b1 );
not ( w_13315 , w_13318 );
not (  , w_13319 );
and ( w_13318 , w_13319 , \4185_b0 );
buf ( \4187_b1 , \4186_b1 );
not ( \4187_b1 , w_13320 );
not ( \4187_b0 , w_13321 );
and ( w_13320 , w_13321 , \4186_b0 );
or ( \4188_b1 , \4184_b1 , w_13322 );
or ( \4188_b0 , \4184_b0 , \4187_b0 );
not ( \4187_b0 , w_13323 );
and ( w_13323 , w_13322 , \4187_b1 );
or ( \4189_b1 , \2477_b1 , \2790_b1 );
not ( \2790_b1 , w_13324 );
and ( \4189_b0 , \2477_b0 , w_13325 );
and ( w_13324 , w_13325 , \2790_b0 );
buf ( \4190_b1 , \2477_b1 );
not ( \4190_b1 , w_13326 );
not ( \4190_b0 , w_13327 );
and ( w_13326 , w_13327 , \2477_b0 );
or ( \4191_b1 , \4190_b1 , \4180_b1 );
not ( \4180_b1 , w_13328 );
and ( \4191_b0 , \4190_b0 , w_13329 );
and ( w_13328 , w_13329 , \4180_b0 );
or ( \4192_b1 , \4189_b1 , w_13330 );
or ( \4192_b0 , \4189_b0 , \4191_b0 );
not ( \4191_b0 , w_13331 );
and ( w_13331 , w_13330 , \4191_b1 );
or ( \4193_b1 , \4188_b1 , w_13333 );
not ( w_13333 , w_13334 );
and ( \4193_b0 , \4188_b0 , w_13335 );
and ( w_13334 ,  , w_13335 );
buf ( w_13333 , \4192_b1 );
not ( w_13333 , w_13336 );
not (  , w_13337 );
and ( w_13336 , w_13337 , \4192_b0 );
buf ( \4194_b1 , \4193_b1 );
not ( \4194_b1 , w_13338 );
not ( \4194_b0 , w_13339 );
and ( w_13338 , w_13339 , \4193_b0 );
buf ( \4195_b1 , \4194_b1 );
buf ( \4195_b0 , \4194_b0 );
buf ( \4196_b1 , \4195_b1 );
not ( \4196_b1 , w_13340 );
not ( \4196_b0 , w_13341 );
and ( w_13340 , w_13341 , \4195_b0 );
or ( \4197_b1 , \4179_b1 , w_13342 );
or ( \4197_b0 , \4179_b0 , \4196_b0 );
not ( \4196_b0 , w_13343 );
and ( w_13343 , w_13342 , \4196_b1 );
or ( \4198_b1 , \4039_b1 , \4090_b1 );
xor ( \4198_b0 , \4039_b0 , w_13344 );
not ( w_13344 , w_13345 );
and ( w_13345 , \4090_b1 , \4090_b0 );
or ( \4199_b1 , \4198_b1 , \4102_b1 );
xor ( \4199_b0 , \4198_b0 , w_13346 );
not ( w_13346 , w_13347 );
and ( w_13347 , \4102_b1 , \4102_b0 );
buf ( \4200_b1 , \4192_b1 );
not ( \4200_b1 , w_13348 );
not ( \4200_b0 , w_13349 );
and ( w_13348 , w_13349 , \4192_b0 );
or ( \4201_b1 , \4199_b1 , w_13351 );
not ( w_13351 , w_13352 );
and ( \4201_b0 , \4199_b0 , w_13353 );
and ( w_13352 ,  , w_13353 );
buf ( w_13351 , \4200_b1 );
not ( w_13351 , w_13354 );
not (  , w_13355 );
and ( w_13354 , w_13355 , \4200_b0 );
or ( \4202_b1 , \4197_b1 , w_13357 );
not ( w_13357 , w_13358 );
and ( \4202_b0 , \4197_b0 , w_13359 );
and ( w_13358 ,  , w_13359 );
buf ( w_13357 , \4201_b1 );
not ( w_13357 , w_13360 );
not (  , w_13361 );
and ( w_13360 , w_13361 , \4201_b0 );
or ( \4203_b1 , \4177_b1 , \4202_b1 );
xor ( \4203_b0 , \4177_b0 , w_13362 );
not ( w_13362 , w_13363 );
and ( w_13363 , \4202_b1 , \4202_b0 );
or ( \4204_b1 , \4102_b1 , \4097_b1 );
not ( \4097_b1 , w_13364 );
and ( \4204_b0 , \4102_b0 , w_13365 );
and ( w_13364 , w_13365 , \4097_b0 );
buf ( \4205_b1 , \4198_b1 );
not ( \4205_b1 , w_13366 );
not ( \4205_b0 , w_13367 );
and ( w_13366 , w_13367 , \4198_b0 );
buf ( \4206_b1 , \4106_b1 );
not ( \4206_b1 , w_13368 );
not ( \4206_b0 , w_13369 );
and ( w_13368 , w_13369 , \4106_b0 );
buf ( \4207_b1 , \4206_b1 );
not ( \4207_b1 , w_13370 );
not ( \4207_b0 , w_13371 );
and ( w_13370 , w_13371 , \4206_b0 );
or ( \4208_b1 , \4205_b1 , w_13372 );
or ( \4208_b0 , \4205_b0 , \4207_b0 );
not ( \4207_b0 , w_13373 );
and ( w_13373 , w_13372 , \4207_b1 );
buf ( \4209_b1 , \4198_b1 );
not ( \4209_b1 , w_13374 );
not ( \4209_b0 , w_13375 );
and ( w_13374 , w_13375 , \4198_b0 );
or ( \4210_b1 , \4110_b1 , w_13377 );
not ( w_13377 , w_13378 );
and ( \4210_b0 , \4110_b0 , w_13379 );
and ( w_13378 ,  , w_13379 );
buf ( w_13377 , \4209_b1 );
not ( w_13377 , w_13380 );
not (  , w_13381 );
and ( w_13380 , w_13381 , \4209_b0 );
or ( \4211_b1 , \4208_b1 , w_13383 );
not ( w_13383 , w_13384 );
and ( \4211_b0 , \4208_b0 , w_13385 );
and ( w_13384 ,  , w_13385 );
buf ( w_13383 , \4210_b1 );
not ( w_13383 , w_13386 );
not (  , w_13387 );
and ( w_13386 , w_13387 , \4210_b0 );
buf ( \4212_b1 , \4211_b1 );
not ( \4212_b1 , w_13388 );
not ( \4212_b0 , w_13389 );
and ( w_13388 , w_13389 , \4211_b0 );
buf ( \4213_b1 , \4129_b1 );
not ( \4213_b1 , w_13390 );
not ( \4213_b0 , w_13391 );
and ( w_13390 , w_13391 , \4129_b0 );
or ( \4214_b1 , \4212_b1 , w_13392 );
or ( \4214_b0 , \4212_b0 , \4213_b0 );
not ( \4213_b0 , w_13393 );
and ( w_13393 , w_13392 , \4213_b1 );
or ( \4215_b1 , \4133_b1 , w_13395 );
not ( w_13395 , w_13396 );
and ( \4215_b0 , \4133_b0 , w_13397 );
and ( w_13396 ,  , w_13397 );
buf ( w_13395 , \4113_b1 );
not ( w_13395 , w_13398 );
not (  , w_13399 );
and ( w_13398 , w_13399 , \4113_b0 );
or ( \4216_b1 , \4214_b1 , w_13401 );
not ( w_13401 , w_13402 );
and ( \4216_b0 , \4214_b0 , w_13403 );
and ( w_13402 ,  , w_13403 );
buf ( w_13401 , \4215_b1 );
not ( w_13401 , w_13404 );
not (  , w_13405 );
and ( w_13404 , w_13405 , \4215_b0 );
or ( \4217_b1 , \4204_b1 , \4216_b1 );
xor ( \4217_b0 , \4204_b0 , w_13406 );
not ( w_13406 , w_13407 );
and ( w_13407 , \4216_b1 , \4216_b0 );
or ( \4218_b1 , \4096_b1 , \4100_b1 );
not ( \4100_b1 , w_13408 );
and ( \4218_b0 , \4096_b0 , w_13409 );
and ( w_13408 , w_13409 , \4100_b0 );
buf ( \4219_b1 , \4096_b1 );
not ( \4219_b1 , w_13410 );
not ( \4219_b0 , w_13411 );
and ( w_13410 , w_13411 , \4096_b0 );
or ( \4220_b1 , \4219_b1 , \4101_b1 );
not ( \4101_b1 , w_13412 );
and ( \4220_b0 , \4219_b0 , w_13413 );
and ( w_13412 , w_13413 , \4101_b0 );
or ( \4221_b1 , \4218_b1 , w_13415 );
not ( w_13415 , w_13416 );
and ( \4221_b0 , \4218_b0 , w_13417 );
and ( w_13416 ,  , w_13417 );
buf ( w_13415 , \4220_b1 );
not ( w_13415 , w_13418 );
not (  , w_13419 );
and ( w_13418 , w_13419 , \4220_b0 );
buf ( \4222_b1 , \4221_b1 );
not ( \4222_b1 , w_13420 );
not ( \4222_b0 , w_13421 );
and ( w_13420 , w_13421 , \4221_b0 );
buf ( \4223_b1 , \4195_b1 );
not ( \4223_b1 , w_13422 );
not ( \4223_b0 , w_13423 );
and ( w_13422 , w_13423 , \4195_b0 );
or ( \4224_b1 , \4222_b1 , w_13424 );
or ( \4224_b0 , \4222_b0 , \4223_b0 );
not ( \4223_b0 , w_13425 );
and ( w_13425 , w_13424 , \4223_b1 );
or ( \4225_b1 , \4178_b1 , w_13427 );
not ( w_13427 , w_13428 );
and ( \4225_b0 , \4178_b0 , w_13429 );
and ( w_13428 ,  , w_13429 );
buf ( w_13427 , \4200_b1 );
not ( w_13427 , w_13430 );
not (  , w_13431 );
and ( w_13430 , w_13431 , \4200_b0 );
or ( \4226_b1 , \4224_b1 , w_13433 );
not ( w_13433 , w_13434 );
and ( \4226_b0 , \4224_b0 , w_13435 );
and ( w_13434 ,  , w_13435 );
buf ( w_13433 , \4225_b1 );
not ( w_13433 , w_13436 );
not (  , w_13437 );
and ( w_13436 , w_13437 , \4225_b0 );
or ( \4227_b1 , \4217_b1 , \4226_b1 );
not ( \4226_b1 , w_13438 );
and ( \4227_b0 , \4217_b0 , w_13439 );
and ( w_13438 , w_13439 , \4226_b0 );
or ( \4228_b1 , \4204_b1 , \4216_b1 );
not ( \4216_b1 , w_13440 );
and ( \4228_b0 , \4204_b0 , w_13441 );
and ( w_13440 , w_13441 , \4216_b0 );
or ( \4229_b1 , \4227_b1 , w_13442 );
or ( \4229_b0 , \4227_b0 , \4228_b0 );
not ( \4228_b0 , w_13443 );
and ( w_13443 , w_13442 , \4228_b1 );
or ( \4230_b1 , \4203_b1 , \4229_b1 );
xor ( \4230_b0 , \4203_b0 , w_13444 );
not ( w_13444 , w_13445 );
and ( w_13445 , \4229_b1 , \4229_b0 );
or ( \4231_b1 , \4166_b1 , \4230_b1 );
xor ( \4231_b0 , \4166_b0 , w_13446 );
not ( w_13446 , w_13447 );
and ( w_13447 , \4230_b1 , \4230_b0 );
buf ( \4232_b1 , \4177_b1 );
not ( \4232_b1 , w_13448 );
not ( \4232_b0 , w_13449 );
and ( w_13448 , w_13449 , \4177_b0 );
or ( \4233_b1 , \4204_b1 , \4216_b1 );
xor ( \4233_b0 , \4204_b0 , w_13450 );
not ( w_13450 , w_13451 );
and ( w_13451 , \4216_b1 , \4216_b0 );
or ( \4234_b1 , \4233_b1 , \4226_b1 );
xor ( \4234_b0 , \4233_b0 , w_13452 );
not ( w_13452 , w_13453 );
and ( w_13453 , \4226_b1 , \4226_b0 );
buf ( \4235_b1 , \4234_b1 );
not ( \4235_b1 , w_13454 );
not ( \4235_b0 , w_13455 );
and ( w_13454 , w_13455 , \4234_b0 );
buf ( \4236_b1 , \4235_b1 );
not ( \4236_b1 , w_13456 );
not ( \4236_b0 , w_13457 );
and ( w_13456 , w_13457 , \4235_b0 );
or ( \4237_b1 , \4232_b1 , w_13458 );
or ( \4237_b0 , \4232_b0 , \4236_b0 );
not ( \4236_b0 , w_13459 );
and ( w_13459 , w_13458 , \4236_b1 );
buf ( \4238_b1 , \3997_b1 );
not ( \4238_b1 , w_13460 );
not ( \4238_b0 , w_13461 );
and ( w_13460 , w_13461 , \3997_b0 );
buf ( \4239_b1 , \4163_b1 );
not ( \4239_b1 , w_13462 );
not ( \4239_b0 , w_13463 );
and ( w_13462 , w_13463 , \4163_b0 );
or ( \4240_b1 , \4238_b1 , w_13464 );
or ( \4240_b0 , \4238_b0 , \4239_b0 );
not ( \4239_b0 , w_13465 );
and ( w_13465 , w_13464 , \4239_b1 );
or ( \4241_b1 , \4170_b1 , w_13467 );
not ( w_13467 , w_13468 );
and ( \4241_b0 , \4170_b0 , w_13469 );
and ( w_13468 ,  , w_13469 );
buf ( w_13467 , \4111_b1 );
not ( w_13467 , w_13470 );
not (  , w_13471 );
and ( w_13470 , w_13471 , \4111_b0 );
or ( \4242_b1 , \4240_b1 , w_13473 );
not ( w_13473 , w_13474 );
and ( \4242_b0 , \4240_b0 , w_13475 );
and ( w_13474 ,  , w_13475 );
buf ( w_13473 , \4241_b1 );
not ( w_13473 , w_13476 );
not (  , w_13477 );
and ( w_13476 , w_13477 , \4241_b0 );
buf ( \4243_b1 , \4242_b1 );
not ( \4243_b1 , w_13478 );
not ( \4243_b0 , w_13479 );
and ( w_13478 , w_13479 , \4242_b0 );
buf ( \4244_b1 , \4159_b1 );
not ( \4244_b1 , w_13480 );
not ( \4244_b0 , w_13481 );
and ( w_13480 , w_13481 , \4159_b0 );
or ( \4245_b1 , \4243_b1 , w_13482 );
or ( \4245_b0 , \4243_b0 , \4244_b0 );
not ( \4244_b0 , w_13483 );
and ( w_13483 , w_13482 , \4244_b1 );
or ( \4246_b1 , \4150_b1 , w_13485 );
not ( w_13485 , w_13486 );
and ( \4246_b0 , \4150_b0 , w_13487 );
and ( w_13486 ,  , w_13487 );
buf ( w_13485 , \4172_b1 );
not ( w_13485 , w_13488 );
not (  , w_13489 );
and ( w_13488 , w_13489 , \4172_b0 );
or ( \4247_b1 , \4245_b1 , w_13491 );
not ( w_13491 , w_13492 );
and ( \4247_b0 , \4245_b0 , w_13493 );
and ( w_13492 ,  , w_13493 );
buf ( w_13491 , \4246_b1 );
not ( w_13491 , w_13494 );
not (  , w_13495 );
and ( w_13494 , w_13495 , \4246_b0 );
buf ( \4248_b1 , \4247_b1 );
not ( \4248_b1 , w_13496 );
not ( \4248_b0 , w_13497 );
and ( w_13496 , w_13497 , \4247_b0 );
buf ( \4249_b1 , \4097_b1 );
not ( \4249_b1 , w_13498 );
not ( \4249_b0 , w_13499 );
and ( w_13498 , w_13499 , \4097_b0 );
buf ( \4250_b1 , \4100_b1 );
not ( \4250_b1 , w_13500 );
not ( \4250_b0 , w_13501 );
and ( w_13500 , w_13501 , \4100_b0 );
buf ( \4251_b1 , \4250_b1 );
not ( \4251_b1 , w_13502 );
not ( \4251_b0 , w_13503 );
and ( w_13502 , w_13503 , \4250_b0 );
or ( \4252_b1 , \4249_b1 , w_13504 );
or ( \4252_b0 , \4249_b0 , \4251_b0 );
not ( \4251_b0 , w_13505 );
and ( w_13505 , w_13504 , \4251_b1 );
buf ( \4253_b1 , \4101_b1 );
not ( \4253_b1 , w_13506 );
not ( \4253_b0 , w_13507 );
and ( w_13506 , w_13507 , \4101_b0 );
buf ( \4254_b1 , \4097_b1 );
not ( \4254_b1 , w_13508 );
not ( \4254_b0 , w_13509 );
and ( w_13508 , w_13509 , \4097_b0 );
or ( \4255_b1 , \4253_b1 , w_13511 );
not ( w_13511 , w_13512 );
and ( \4255_b0 , \4253_b0 , w_13513 );
and ( w_13512 ,  , w_13513 );
buf ( w_13511 , \4254_b1 );
not ( w_13511 , w_13514 );
not (  , w_13515 );
and ( w_13514 , w_13515 , \4254_b0 );
or ( \4256_b1 , \4252_b1 , w_13517 );
not ( w_13517 , w_13518 );
and ( \4256_b0 , \4252_b0 , w_13519 );
and ( w_13518 ,  , w_13519 );
buf ( w_13517 , \4255_b1 );
not ( w_13517 , w_13520 );
not (  , w_13521 );
and ( w_13520 , w_13521 , \4255_b0 );
buf ( \4257_b1 , \4256_b1 );
not ( \4257_b1 , w_13522 );
not ( \4257_b0 , w_13523 );
and ( w_13522 , w_13523 , \4256_b0 );
buf ( \4258_b1 , \4195_b1 );
not ( \4258_b1 , w_13524 );
not ( \4258_b0 , w_13525 );
and ( w_13524 , w_13525 , \4195_b0 );
or ( \4259_b1 , \4257_b1 , w_13526 );
or ( \4259_b0 , \4257_b0 , \4258_b0 );
not ( \4258_b0 , w_13527 );
and ( w_13527 , w_13526 , \4258_b1 );
or ( \4260_b1 , \4221_b1 , w_13529 );
not ( w_13529 , w_13530 );
and ( \4260_b0 , \4221_b0 , w_13531 );
and ( w_13530 ,  , w_13531 );
buf ( w_13529 , \4200_b1 );
not ( w_13529 , w_13532 );
not (  , w_13533 );
and ( w_13532 , w_13533 , \4200_b0 );
or ( \4261_b1 , \4259_b1 , w_13535 );
not ( w_13535 , w_13536 );
and ( \4261_b0 , \4259_b0 , w_13537 );
and ( w_13536 ,  , w_13537 );
buf ( w_13535 , \4260_b1 );
not ( w_13535 , w_13538 );
not (  , w_13539 );
and ( w_13538 , w_13539 , \4260_b0 );
buf ( \4262_b1 , \4261_b1 );
not ( \4262_b1 , w_13540 );
not ( \4262_b0 , w_13541 );
and ( w_13540 , w_13541 , \4261_b0 );
or ( \4263_b1 , \4248_b1 , w_13542 );
or ( \4263_b0 , \4248_b0 , \4262_b0 );
not ( \4262_b0 , w_13543 );
and ( w_13543 , w_13542 , \4262_b1 );
or ( \4264_b1 , \4261_b1 , w_13544 );
or ( \4264_b0 , \4261_b0 , \4247_b0 );
not ( \4247_b0 , w_13545 );
and ( w_13545 , w_13544 , \4247_b1 );
or ( \4265_b1 , \3136_b1 , w_13546 );
xor ( \4265_b0 , \3136_b0 , w_13548 );
not ( w_13548 , w_13549 );
and ( w_13549 , w_13546 , w_13547 );
buf ( w_13546 , \3326_b1 );
not ( w_13546 , w_13550 );
not ( w_13547 , w_13551 );
and ( w_13550 , w_13551 , \3326_b0 );
buf ( \4266_b1 , \4265_b1 );
not ( \4266_b1 , w_13552 );
not ( \4266_b0 , w_13553 );
and ( w_13552 , w_13553 , \4265_b0 );
buf ( \4267_b1 , \4266_b1 );
not ( \4267_b1 , w_13554 );
not ( \4267_b0 , w_13555 );
and ( w_13554 , w_13555 , \4266_b0 );
buf ( \4268_b1 , \4267_b1 );
buf ( \4268_b0 , \4267_b0 );
buf ( \4269_b1 , \4268_b1 );
not ( \4269_b1 , w_13556 );
not ( \4269_b0 , w_13557 );
and ( w_13556 , w_13557 , \4268_b0 );
buf ( \4270_b1 , \3136_b1 );
not ( \4270_b1 , w_13558 );
not ( \4270_b0 , w_13559 );
and ( w_13558 , w_13559 , \3136_b0 );
or ( \4271_b1 , \4270_b1 , w_13561 );
not ( w_13561 , w_13562 );
and ( \4271_b0 , \4270_b0 , w_13563 );
and ( w_13562 ,  , w_13563 );
buf ( w_13561 , \3637_b1 );
not ( w_13561 , w_13564 );
not (  , w_13565 );
and ( w_13564 , w_13565 , \3637_b0 );
buf ( \4272_b1 , \4271_b1 );
not ( \4272_b1 , w_13566 );
not ( \4272_b0 , w_13567 );
and ( w_13566 , w_13567 , \4271_b0 );
buf ( \4273_b1 , \3637_b1 );
not ( \4273_b1 , w_13568 );
not ( \4273_b0 , w_13569 );
and ( w_13568 , w_13569 , \3637_b0 );
buf ( \4274_b1 , \4270_b1 );
not ( \4274_b1 , w_13570 );
not ( \4274_b0 , w_13571 );
and ( w_13570 , w_13571 , \4270_b0 );
or ( \4275_b1 , \4273_b1 , w_13573 );
not ( w_13573 , w_13574 );
and ( \4275_b0 , \4273_b0 , w_13575 );
and ( w_13574 ,  , w_13575 );
buf ( w_13573 , \4274_b1 );
not ( w_13573 , w_13576 );
not (  , w_13577 );
and ( w_13576 , w_13577 , \4274_b0 );
buf ( \4276_b1 , \4275_b1 );
not ( \4276_b1 , w_13578 );
not ( \4276_b0 , w_13579 );
and ( w_13578 , w_13579 , \4275_b0 );
or ( \4277_b1 , \4272_b1 , w_13580 );
or ( \4277_b0 , \4272_b0 , \4276_b0 );
not ( \4276_b0 , w_13581 );
and ( w_13581 , w_13580 , \4276_b1 );
or ( \4278_b1 , \4277_b1 , w_13583 );
not ( w_13583 , w_13584 );
and ( \4278_b0 , \4277_b0 , w_13585 );
and ( w_13584 ,  , w_13585 );
buf ( w_13583 , \4265_b1 );
not ( w_13583 , w_13586 );
not (  , w_13587 );
and ( w_13586 , w_13587 , \4265_b0 );
buf ( \4279_b1 , \4278_b1 );
not ( \4279_b1 , w_13588 );
not ( \4279_b0 , w_13589 );
and ( w_13588 , w_13589 , \4278_b0 );
buf ( \4280_b1 , \4279_b1 );
not ( \4280_b1 , w_13590 );
not ( \4280_b0 , w_13591 );
and ( w_13590 , w_13591 , \4279_b0 );
buf ( \4281_b1 , \4280_b1 );
not ( \4281_b1 , w_13592 );
not ( \4281_b0 , w_13593 );
and ( w_13592 , w_13593 , \4280_b0 );
or ( \4282_b1 , \4269_b1 , w_13594 );
or ( \4282_b0 , \4269_b0 , \4281_b0 );
not ( \4281_b0 , w_13595 );
and ( w_13595 , w_13594 , \4281_b1 );
buf ( \4283_b1 , \3637_b1 );
buf ( \4283_b0 , \3637_b0 );
buf ( \4284_b1 , \4283_b1 );
not ( \4284_b1 , w_13596 );
not ( \4284_b0 , w_13597 );
and ( w_13596 , w_13597 , \4283_b0 );
buf ( \4285_b1 , \4284_b1 );
not ( \4285_b1 , w_13598 );
not ( \4285_b0 , w_13599 );
and ( w_13598 , w_13599 , \4284_b0 );
or ( \4286_b1 , \4282_b1 , w_13601 );
not ( w_13601 , w_13602 );
and ( \4286_b0 , \4282_b0 , w_13603 );
and ( w_13602 ,  , w_13603 );
buf ( w_13601 , \4285_b1 );
not ( w_13601 , w_13604 );
not (  , w_13605 );
and ( w_13604 , w_13605 , \4285_b0 );
or ( \4287_b1 , \4264_b1 , w_13607 );
not ( w_13607 , w_13608 );
and ( \4287_b0 , \4264_b0 , w_13609 );
and ( w_13608 ,  , w_13609 );
buf ( w_13607 , \4286_b1 );
not ( w_13607 , w_13610 );
not (  , w_13611 );
and ( w_13610 , w_13611 , \4286_b0 );
or ( \4288_b1 , \4263_b1 , w_13613 );
not ( w_13613 , w_13614 );
and ( \4288_b0 , \4263_b0 , w_13615 );
and ( w_13614 ,  , w_13615 );
buf ( w_13613 , \4287_b1 );
not ( w_13613 , w_13616 );
not (  , w_13617 );
and ( w_13616 , w_13617 , \4287_b0 );
or ( \4289_b1 , \4237_b1 , w_13619 );
not ( w_13619 , w_13620 );
and ( \4289_b0 , \4237_b0 , w_13621 );
and ( w_13620 ,  , w_13621 );
buf ( w_13619 , \4288_b1 );
not ( w_13619 , w_13622 );
not (  , w_13623 );
and ( w_13622 , w_13623 , \4288_b0 );
buf ( \4290_b1 , \4177_b1 );
not ( \4290_b1 , w_13624 );
not ( \4290_b0 , w_13625 );
and ( w_13624 , w_13625 , \4177_b0 );
or ( \4291_b1 , \4290_b1 , w_13627 );
not ( w_13627 , w_13628 );
and ( \4291_b0 , \4290_b0 , w_13629 );
and ( w_13628 ,  , w_13629 );
buf ( w_13627 , \4234_b1 );
not ( w_13627 , w_13630 );
not (  , w_13631 );
and ( w_13630 , w_13631 , \4234_b0 );
or ( \4292_b1 , \4289_b1 , w_13633 );
not ( w_13633 , w_13634 );
and ( \4292_b0 , \4289_b0 , w_13635 );
and ( w_13634 ,  , w_13635 );
buf ( w_13633 , \4291_b1 );
not ( w_13633 , w_13636 );
not (  , w_13637 );
and ( w_13636 , w_13637 , \4291_b0 );
or ( \4293_b1 , \4231_b1 , w_13638 );
xor ( \4293_b0 , \4231_b0 , w_13640 );
not ( w_13640 , w_13641 );
and ( w_13641 , w_13638 , w_13639 );
buf ( w_13638 , \4292_b1 );
not ( w_13638 , w_13642 );
not ( w_13639 , w_13643 );
and ( w_13642 , w_13643 , \4292_b0 );
or ( \4294_b1 , \4102_b1 , \4093_b1 );
not ( \4093_b1 , w_13644 );
and ( \4294_b0 , \4102_b0 , w_13645 );
and ( w_13644 , w_13645 , \4093_b0 );
buf ( \4295_b1 , \4094_b1 );
not ( \4295_b1 , w_13646 );
not ( \4295_b0 , w_13647 );
and ( w_13646 , w_13647 , \4094_b0 );
buf ( \4296_b1 , \4206_b1 );
not ( \4296_b1 , w_13648 );
not ( \4296_b0 , w_13649 );
and ( w_13648 , w_13649 , \4206_b0 );
or ( \4297_b1 , \4295_b1 , w_13650 );
or ( \4297_b0 , \4295_b0 , \4296_b0 );
not ( \4296_b0 , w_13651 );
and ( w_13651 , w_13650 , \4296_b1 );
buf ( \4298_b1 , \4094_b1 );
not ( \4298_b1 , w_13652 );
not ( \4298_b0 , w_13653 );
and ( w_13652 , w_13653 , \4094_b0 );
or ( \4299_b1 , \4106_b1 , w_13655 );
not ( w_13655 , w_13656 );
and ( \4299_b0 , \4106_b0 , w_13657 );
and ( w_13656 ,  , w_13657 );
buf ( w_13655 , \4298_b1 );
not ( w_13655 , w_13658 );
not (  , w_13659 );
and ( w_13658 , w_13659 , \4298_b0 );
or ( \4300_b1 , \4297_b1 , w_13661 );
not ( w_13661 , w_13662 );
and ( \4300_b0 , \4297_b0 , w_13663 );
and ( w_13662 ,  , w_13663 );
buf ( w_13661 , \4299_b1 );
not ( w_13661 , w_13664 );
not (  , w_13665 );
and ( w_13664 , w_13665 , \4299_b0 );
buf ( \4301_b1 , \4300_b1 );
not ( \4301_b1 , w_13666 );
not ( \4301_b0 , w_13667 );
and ( w_13666 , w_13667 , \4300_b0 );
buf ( \4302_b1 , \4128_b1 );
buf ( \4302_b0 , \4128_b0 );
buf ( \4303_b1 , \4302_b1 );
not ( \4303_b1 , w_13668 );
not ( \4303_b0 , w_13669 );
and ( w_13668 , w_13669 , \4302_b0 );
or ( \4304_b1 , \4301_b1 , w_13670 );
or ( \4304_b0 , \4301_b0 , \4303_b0 );
not ( \4303_b0 , w_13671 );
and ( w_13671 , w_13670 , \4303_b1 );
or ( \4305_b1 , \4133_b1 , w_13673 );
not ( w_13673 , w_13674 );
and ( \4305_b0 , \4133_b0 , w_13675 );
and ( w_13674 ,  , w_13675 );
buf ( w_13673 , \4211_b1 );
not ( w_13673 , w_13676 );
not (  , w_13677 );
and ( w_13676 , w_13677 , \4211_b0 );
or ( \4306_b1 , \4304_b1 , w_13679 );
not ( w_13679 , w_13680 );
and ( \4306_b0 , \4304_b0 , w_13681 );
and ( w_13680 ,  , w_13681 );
buf ( w_13679 , \4305_b1 );
not ( w_13679 , w_13682 );
not (  , w_13683 );
and ( w_13682 , w_13683 , \4305_b0 );
or ( \4307_b1 , \4294_b1 , \4306_b1 );
xor ( \4307_b0 , \4294_b0 , w_13684 );
not ( w_13684 , w_13685 );
and ( w_13685 , \4306_b1 , \4306_b0 );
buf ( \4308_b1 , \4198_b1 );
not ( \4308_b1 , w_13686 );
not ( \4308_b0 , w_13687 );
and ( w_13686 , w_13687 , \4198_b0 );
buf ( \4309_b1 , \4163_b1 );
not ( \4309_b1 , w_13688 );
not ( \4309_b0 , w_13689 );
and ( w_13688 , w_13689 , \4163_b0 );
or ( \4310_b1 , \4308_b1 , w_13690 );
or ( \4310_b0 , \4308_b0 , \4309_b0 );
not ( \4309_b0 , w_13691 );
and ( w_13691 , w_13690 , \4309_b1 );
buf ( \4311_b1 , \4163_b1 );
not ( \4311_b1 , w_13692 );
not ( \4311_b0 , w_13693 );
and ( w_13692 , w_13693 , \4163_b0 );
or ( \4312_b1 , \4311_b1 , w_13695 );
not ( w_13695 , w_13696 );
and ( \4312_b0 , \4311_b0 , w_13697 );
and ( w_13696 ,  , w_13697 );
buf ( w_13695 , \4209_b1 );
not ( w_13695 , w_13698 );
not (  , w_13699 );
and ( w_13698 , w_13699 , \4209_b0 );
or ( \4313_b1 , \4310_b1 , w_13701 );
not ( w_13701 , w_13702 );
and ( \4313_b0 , \4310_b0 , w_13703 );
and ( w_13702 ,  , w_13703 );
buf ( w_13701 , \4312_b1 );
not ( w_13701 , w_13704 );
not (  , w_13705 );
and ( w_13704 , w_13705 , \4312_b0 );
buf ( \4314_b1 , \4313_b1 );
not ( \4314_b1 , w_13706 );
not ( \4314_b0 , w_13707 );
and ( w_13706 , w_13707 , \4313_b0 );
buf ( \4315_b1 , \4159_b1 );
not ( \4315_b1 , w_13708 );
not ( \4315_b0 , w_13709 );
and ( w_13708 , w_13709 , \4159_b0 );
or ( \4316_b1 , \4314_b1 , w_13710 );
or ( \4316_b0 , \4314_b0 , \4315_b0 );
not ( \4315_b0 , w_13711 );
and ( w_13711 , w_13710 , \4315_b1 );
buf ( \4317_b1 , \4150_b1 );
buf ( \4317_b0 , \4150_b0 );
or ( \4318_b1 , \4317_b1 , w_13713 );
not ( w_13713 , w_13714 );
and ( \4318_b0 , \4317_b0 , w_13715 );
and ( w_13714 ,  , w_13715 );
buf ( w_13713 , \4242_b1 );
not ( w_13713 , w_13716 );
not (  , w_13717 );
and ( w_13716 , w_13717 , \4242_b0 );
or ( \4319_b1 , \4316_b1 , w_13719 );
not ( w_13719 , w_13720 );
and ( \4319_b0 , \4316_b0 , w_13721 );
and ( w_13720 ,  , w_13721 );
buf ( w_13719 , \4318_b1 );
not ( w_13719 , w_13722 );
not (  , w_13723 );
and ( w_13722 , w_13723 , \4318_b0 );
or ( \4320_b1 , \4307_b1 , \4319_b1 );
not ( \4319_b1 , w_13724 );
and ( \4320_b0 , \4307_b0 , w_13725 );
and ( w_13724 , w_13725 , \4319_b0 );
or ( \4321_b1 , \4294_b1 , \4306_b1 );
not ( \4306_b1 , w_13726 );
and ( \4321_b0 , \4294_b0 , w_13727 );
and ( w_13726 , w_13727 , \4306_b0 );
or ( \4322_b1 , \4320_b1 , w_13728 );
or ( \4322_b0 , \4320_b0 , \4321_b0 );
not ( \4321_b0 , w_13729 );
and ( w_13729 , w_13728 , \4321_b1 );
buf ( \4323_b1 , \4322_b1 );
not ( \4323_b1 , w_13730 );
not ( \4323_b0 , w_13731 );
and ( w_13730 , w_13731 , \4322_b0 );
or ( \4324_b1 , \4177_b1 , \4288_b1 );
xor ( \4324_b0 , \4177_b0 , w_13732 );
not ( w_13732 , w_13733 );
and ( w_13733 , \4288_b1 , \4288_b0 );
or ( \4325_b1 , \4324_b1 , w_13734 );
xor ( \4325_b0 , \4324_b0 , w_13736 );
not ( w_13736 , w_13737 );
and ( w_13737 , w_13734 , w_13735 );
buf ( w_13734 , \4234_b1 );
not ( w_13734 , w_13738 );
not ( w_13735 , w_13739 );
and ( w_13738 , w_13739 , \4234_b0 );
buf ( \4326_b1 , \4325_b1 );
not ( \4326_b1 , w_13740 );
not ( \4326_b0 , w_13741 );
and ( w_13740 , w_13741 , \4325_b0 );
or ( \4327_b1 , \4323_b1 , w_13743 );
not ( w_13743 , w_13744 );
and ( \4327_b0 , \4323_b0 , w_13745 );
and ( w_13744 ,  , w_13745 );
buf ( w_13743 , \4326_b1 );
not ( w_13743 , w_13746 );
not (  , w_13747 );
and ( w_13746 , w_13747 , \4326_b0 );
or ( \4328_b1 , \4294_b1 , \4306_b1 );
xor ( \4328_b0 , \4294_b0 , w_13748 );
not ( w_13748 , w_13749 );
and ( w_13749 , \4306_b1 , \4306_b0 );
or ( \4329_b1 , \4328_b1 , \4319_b1 );
xor ( \4329_b0 , \4328_b0 , w_13750 );
not ( w_13750 , w_13751 );
and ( w_13751 , \4319_b1 , \4319_b0 );
or ( \4330_b1 , \4102_b1 , \4095_b1 );
not ( \4095_b1 , w_13752 );
and ( \4330_b0 , \4102_b0 , w_13753 );
and ( w_13752 , w_13753 , \4095_b0 );
buf ( \4331_b1 , \4051_b1 );
not ( \4331_b1 , w_13754 );
not ( \4331_b0 , w_13755 );
and ( w_13754 , w_13755 , \4051_b0 );
buf ( \4332_b1 , \3637_b1 );
not ( \4332_b1 , w_13756 );
not ( \4332_b0 , w_13757 );
and ( w_13756 , w_13757 , \3637_b0 );
buf ( \4333_b1 , \4332_b1 );
not ( \4333_b1 , w_13758 );
not ( \4333_b0 , w_13759 );
and ( w_13758 , w_13759 , \4332_b0 );
or ( \4334_b1 , \4331_b1 , w_13760 );
or ( \4334_b0 , \4331_b0 , \4333_b0 );
not ( \4333_b0 , w_13761 );
and ( w_13761 , w_13760 , \4333_b1 );
or ( \4335_b1 , \4283_b1 , w_13763 );
not ( w_13763 , w_13764 );
and ( \4335_b0 , \4283_b0 , w_13765 );
and ( w_13764 ,  , w_13765 );
buf ( w_13763 , \4135_b1 );
not ( w_13763 , w_13766 );
not (  , w_13767 );
and ( w_13766 , w_13767 , \4135_b0 );
or ( \4336_b1 , \4334_b1 , w_13769 );
not ( w_13769 , w_13770 );
and ( \4336_b0 , \4334_b0 , w_13771 );
and ( w_13770 ,  , w_13771 );
buf ( w_13769 , \4335_b1 );
not ( w_13769 , w_13772 );
not (  , w_13773 );
and ( w_13772 , w_13773 , \4335_b0 );
buf ( \4337_b1 , \4336_b1 );
not ( \4337_b1 , w_13774 );
not ( \4337_b0 , w_13775 );
and ( w_13774 , w_13775 , \4336_b0 );
buf ( \4338_b1 , \4280_b1 );
not ( \4338_b1 , w_13776 );
not ( \4338_b0 , w_13777 );
and ( w_13776 , w_13777 , \4280_b0 );
buf ( \4339_b1 , \4338_b1 );
not ( \4339_b1 , w_13778 );
not ( \4339_b0 , w_13779 );
and ( w_13778 , w_13779 , \4338_b0 );
or ( \4340_b1 , \4337_b1 , w_13780 );
or ( \4340_b0 , \4337_b0 , \4339_b0 );
not ( \4339_b0 , w_13781 );
and ( w_13781 , w_13780 , \4339_b1 );
buf ( \4341_b1 , \4268_b1 );
not ( \4341_b1 , w_13782 );
not ( \4341_b0 , w_13783 );
and ( w_13782 , w_13783 , \4268_b0 );
or ( \4342_b1 , \4341_b1 , w_13785 );
not ( w_13785 , w_13786 );
and ( \4342_b0 , \4341_b0 , w_13787 );
and ( w_13786 ,  , w_13787 );
buf ( w_13785 , \4285_b1 );
not ( w_13785 , w_13788 );
not (  , w_13789 );
and ( w_13788 , w_13789 , \4285_b0 );
or ( \4343_b1 , \4340_b1 , w_13791 );
not ( w_13791 , w_13792 );
and ( \4343_b0 , \4340_b0 , w_13793 );
and ( w_13792 ,  , w_13793 );
buf ( w_13791 , \4342_b1 );
not ( w_13791 , w_13794 );
not (  , w_13795 );
and ( w_13794 , w_13795 , \4342_b0 );
or ( \4344_b1 , \4330_b1 , \4343_b1 );
xor ( \4344_b0 , \4330_b0 , w_13796 );
not ( w_13796 , w_13797 );
and ( w_13797 , \4343_b1 , \4343_b0 );
buf ( \4345_b1 , \4093_b1 );
not ( \4345_b1 , w_13798 );
not ( \4345_b0 , w_13799 );
and ( w_13798 , w_13799 , \4093_b0 );
buf ( \4346_b1 , \4100_b1 );
not ( \4346_b1 , w_13800 );
not ( \4346_b0 , w_13801 );
and ( w_13800 , w_13801 , \4100_b0 );
buf ( \4347_b1 , \4346_b1 );
not ( \4347_b1 , w_13802 );
not ( \4347_b0 , w_13803 );
and ( w_13802 , w_13803 , \4346_b0 );
or ( \4348_b1 , \4345_b1 , w_13804 );
or ( \4348_b0 , \4345_b0 , \4347_b0 );
not ( \4347_b0 , w_13805 );
and ( w_13805 , w_13804 , \4347_b1 );
buf ( \4349_b1 , \4093_b1 );
not ( \4349_b1 , w_13806 );
not ( \4349_b0 , w_13807 );
and ( w_13806 , w_13807 , \4093_b0 );
or ( \4350_b1 , \4100_b1 , w_13809 );
not ( w_13809 , w_13810 );
and ( \4350_b0 , \4100_b0 , w_13811 );
and ( w_13810 ,  , w_13811 );
buf ( w_13809 , \4349_b1 );
not ( w_13809 , w_13812 );
not (  , w_13813 );
and ( w_13812 , w_13813 , \4349_b0 );
or ( \4351_b1 , \4348_b1 , w_13815 );
not ( w_13815 , w_13816 );
and ( \4351_b0 , \4348_b0 , w_13817 );
and ( w_13816 ,  , w_13817 );
buf ( w_13815 , \4350_b1 );
not ( w_13815 , w_13818 );
not (  , w_13819 );
and ( w_13818 , w_13819 , \4350_b0 );
buf ( \4352_b1 , \4351_b1 );
not ( \4352_b1 , w_13820 );
not ( \4352_b0 , w_13821 );
and ( w_13820 , w_13821 , \4351_b0 );
buf ( \4353_b1 , \4195_b1 );
not ( \4353_b1 , w_13822 );
not ( \4353_b0 , w_13823 );
and ( w_13822 , w_13823 , \4195_b0 );
or ( \4354_b1 , \4352_b1 , w_13824 );
or ( \4354_b0 , \4352_b0 , \4353_b0 );
not ( \4353_b0 , w_13825 );
and ( w_13825 , w_13824 , \4353_b1 );
or ( \4355_b1 , \4256_b1 , w_13827 );
not ( w_13827 , w_13828 );
and ( \4355_b0 , \4256_b0 , w_13829 );
and ( w_13828 ,  , w_13829 );
buf ( w_13827 , \4200_b1 );
not ( w_13827 , w_13830 );
not (  , w_13831 );
and ( w_13830 , w_13831 , \4200_b0 );
or ( \4356_b1 , \4354_b1 , w_13833 );
not ( w_13833 , w_13834 );
and ( \4356_b0 , \4354_b0 , w_13835 );
and ( w_13834 ,  , w_13835 );
buf ( w_13833 , \4355_b1 );
not ( w_13833 , w_13836 );
not (  , w_13837 );
and ( w_13836 , w_13837 , \4355_b0 );
or ( \4357_b1 , \4344_b1 , \4356_b1 );
not ( \4356_b1 , w_13838 );
and ( \4357_b0 , \4344_b0 , w_13839 );
and ( w_13838 , w_13839 , \4356_b0 );
or ( \4358_b1 , \4330_b1 , \4343_b1 );
not ( \4343_b1 , w_13840 );
and ( \4358_b0 , \4330_b0 , w_13841 );
and ( w_13840 , w_13841 , \4343_b0 );
or ( \4359_b1 , \4357_b1 , w_13842 );
or ( \4359_b0 , \4357_b0 , \4358_b0 );
not ( \4358_b0 , w_13843 );
and ( w_13843 , w_13842 , \4358_b1 );
or ( \4360_b1 , \4329_b1 , \4359_b1 );
xor ( \4360_b0 , \4329_b0 , w_13844 );
not ( w_13844 , w_13845 );
and ( w_13845 , \4359_b1 , \4359_b0 );
or ( \4361_b1 , \4286_b1 , \4247_b1 );
xor ( \4361_b0 , \4286_b0 , w_13846 );
not ( w_13846 , w_13847 );
and ( w_13847 , \4247_b1 , \4247_b0 );
or ( \4362_b1 , \4361_b1 , \4261_b1 );
xor ( \4362_b0 , \4361_b0 , w_13848 );
not ( w_13848 , w_13849 );
and ( w_13849 , \4261_b1 , \4261_b0 );
or ( \4363_b1 , \4360_b1 , \4362_b1 );
not ( \4362_b1 , w_13850 );
and ( \4363_b0 , \4360_b0 , w_13851 );
and ( w_13850 , w_13851 , \4362_b0 );
or ( \4364_b1 , \4329_b1 , \4359_b1 );
not ( \4359_b1 , w_13852 );
and ( \4364_b0 , \4329_b0 , w_13853 );
and ( w_13852 , w_13853 , \4359_b0 );
or ( \4365_b1 , \4363_b1 , w_13854 );
or ( \4365_b0 , \4363_b0 , \4364_b0 );
not ( \4364_b0 , w_13855 );
and ( w_13855 , w_13854 , \4364_b1 );
or ( \4366_b1 , \4327_b1 , \4365_b1 );
not ( \4365_b1 , w_13856 );
and ( \4366_b0 , \4327_b0 , w_13857 );
and ( w_13856 , w_13857 , \4365_b0 );
buf ( \4367_b1 , \4322_b1 );
not ( \4367_b1 , w_13858 );
not ( \4367_b0 , w_13859 );
and ( w_13858 , w_13859 , \4322_b0 );
or ( \4368_b1 , \4367_b1 , w_13861 );
not ( w_13861 , w_13862 );
and ( \4368_b0 , \4367_b0 , w_13863 );
and ( w_13862 ,  , w_13863 );
buf ( w_13861 , \4326_b1 );
not ( w_13861 , w_13864 );
not (  , w_13865 );
and ( w_13864 , w_13865 , \4326_b0 );
or ( \4369_b1 , \4366_b1 , w_13867 );
not ( w_13867 , w_13868 );
and ( \4369_b0 , \4366_b0 , w_13869 );
and ( w_13868 ,  , w_13869 );
buf ( w_13867 , \4368_b1 );
not ( w_13867 , w_13870 );
not (  , w_13871 );
and ( w_13870 , w_13871 , \4368_b0 );
or ( \4370_b1 , \4293_b1 , w_13873 );
not ( w_13873 , w_13874 );
and ( \4370_b0 , \4293_b0 , w_13875 );
and ( w_13874 ,  , w_13875 );
buf ( w_13873 , \4369_b1 );
not ( w_13873 , w_13876 );
not (  , w_13877 );
and ( w_13876 , w_13877 , \4369_b0 );
buf ( \4371_b1 , \4370_b1 );
not ( \4371_b1 , w_13878 );
not ( \4371_b0 , w_13879 );
and ( w_13878 , w_13879 , \4370_b0 );
buf ( \4372_b1 , \4096_b1 );
not ( \4372_b1 , w_13880 );
not ( \4372_b0 , w_13881 );
and ( w_13880 , w_13881 , \4096_b0 );
buf ( \4373_b1 , \4372_b1 );
not ( \4373_b1 , w_13882 );
not ( \4373_b0 , w_13883 );
and ( w_13882 , w_13883 , \4372_b0 );
buf ( \4374_b1 , \4106_b1 );
not ( \4374_b1 , w_13884 );
not ( \4374_b0 , w_13885 );
and ( w_13884 , w_13885 , \4106_b0 );
or ( \4375_b1 , \4373_b1 , w_13886 );
or ( \4375_b0 , \4373_b0 , \4374_b0 );
not ( \4374_b0 , w_13887 );
and ( w_13887 , w_13886 , \4374_b1 );
or ( \4376_b1 , \4206_b1 , w_13889 );
not ( w_13889 , w_13890 );
and ( \4376_b0 , \4206_b0 , w_13891 );
and ( w_13890 ,  , w_13891 );
buf ( w_13889 , \4096_b1 );
not ( w_13889 , w_13892 );
not (  , w_13893 );
and ( w_13892 , w_13893 , \4096_b0 );
or ( \4377_b1 , \4375_b1 , w_13895 );
not ( w_13895 , w_13896 );
and ( \4377_b0 , \4375_b0 , w_13897 );
and ( w_13896 ,  , w_13897 );
buf ( w_13895 , \4376_b1 );
not ( w_13895 , w_13898 );
not (  , w_13899 );
and ( w_13898 , w_13899 , \4376_b0 );
buf ( \4378_b1 , \4377_b1 );
not ( \4378_b1 , w_13900 );
not ( \4378_b0 , w_13901 );
and ( w_13900 , w_13901 , \4377_b0 );
buf ( \4379_b1 , \4302_b1 );
not ( \4379_b1 , w_13902 );
not ( \4379_b0 , w_13903 );
and ( w_13902 , w_13903 , \4302_b0 );
or ( \4380_b1 , \4378_b1 , w_13904 );
or ( \4380_b0 , \4378_b0 , \4379_b0 );
not ( \4379_b0 , w_13905 );
and ( w_13905 , w_13904 , \4379_b1 );
or ( \4381_b1 , \4133_b1 , w_13907 );
not ( w_13907 , w_13908 );
and ( \4381_b0 , \4133_b0 , w_13909 );
and ( w_13908 ,  , w_13909 );
buf ( w_13907 , \4300_b1 );
not ( w_13907 , w_13910 );
not (  , w_13911 );
and ( w_13910 , w_13911 , \4300_b0 );
or ( \4382_b1 , \4380_b1 , w_13913 );
not ( w_13913 , w_13914 );
and ( \4382_b0 , \4380_b0 , w_13915 );
and ( w_13914 ,  , w_13915 );
buf ( w_13913 , \4381_b1 );
not ( w_13913 , w_13916 );
not (  , w_13917 );
and ( w_13916 , w_13917 , \4381_b0 );
buf ( \4383_b1 , \4382_b1 );
not ( \4383_b1 , w_13918 );
not ( \4383_b0 , w_13919 );
and ( w_13918 , w_13919 , \4382_b0 );
or ( \4384_b1 , \4383_b1 , w_13921 );
not ( w_13921 , w_13922 );
and ( \4384_b0 , \4383_b0 , w_13923 );
and ( w_13922 ,  , w_13923 );
buf ( w_13921 , \4319_b1 );
not ( w_13921 , w_13924 );
not (  , w_13925 );
and ( w_13924 , w_13925 , \4319_b0 );
buf ( \4385_b1 , \4384_b1 );
not ( \4385_b1 , w_13926 );
not ( \4385_b0 , w_13927 );
and ( w_13926 , w_13927 , \4384_b0 );
or ( \4386_b1 , \4100_b1 , \4066_b1 );
not ( \4066_b1 , w_13928 );
and ( \4386_b0 , \4100_b0 , w_13929 );
and ( w_13928 , w_13929 , \4066_b0 );
buf ( \4387_b1 , \4095_b1 );
not ( \4387_b1 , w_13930 );
not ( \4387_b0 , w_13931 );
and ( w_13930 , w_13931 , \4095_b0 );
buf ( \4388_b1 , \4100_b1 );
not ( \4388_b1 , w_13932 );
not ( \4388_b0 , w_13933 );
and ( w_13932 , w_13933 , \4100_b0 );
buf ( \4389_b1 , \4388_b1 );
not ( \4389_b1 , w_13934 );
not ( \4389_b0 , w_13935 );
and ( w_13934 , w_13935 , \4388_b0 );
or ( \4390_b1 , \4387_b1 , w_13936 );
or ( \4390_b0 , \4387_b0 , \4389_b0 );
not ( \4389_b0 , w_13937 );
and ( w_13937 , w_13936 , \4389_b1 );
buf ( \4391_b1 , \4095_b1 );
not ( \4391_b1 , w_13938 );
not ( \4391_b0 , w_13939 );
and ( w_13938 , w_13939 , \4095_b0 );
or ( \4392_b1 , \4100_b1 , w_13941 );
not ( w_13941 , w_13942 );
and ( \4392_b0 , \4100_b0 , w_13943 );
and ( w_13942 ,  , w_13943 );
buf ( w_13941 , \4391_b1 );
not ( w_13941 , w_13944 );
not (  , w_13945 );
and ( w_13944 , w_13945 , \4391_b0 );
or ( \4393_b1 , \4390_b1 , w_13947 );
not ( w_13947 , w_13948 );
and ( \4393_b0 , \4390_b0 , w_13949 );
and ( w_13948 ,  , w_13949 );
buf ( w_13947 , \4392_b1 );
not ( w_13947 , w_13950 );
not (  , w_13951 );
and ( w_13950 , w_13951 , \4392_b0 );
buf ( \4394_b1 , \4393_b1 );
not ( \4394_b1 , w_13952 );
not ( \4394_b0 , w_13953 );
and ( w_13952 , w_13953 , \4393_b0 );
buf ( \4395_b1 , \4193_b1 );
not ( \4395_b1 , w_13954 );
not ( \4395_b0 , w_13955 );
and ( w_13954 , w_13955 , \4193_b0 );
buf ( \4396_b1 , \4395_b1 );
not ( \4396_b1 , w_13956 );
not ( \4396_b0 , w_13957 );
and ( w_13956 , w_13957 , \4395_b0 );
or ( \4397_b1 , \4394_b1 , w_13958 );
or ( \4397_b0 , \4394_b0 , \4396_b0 );
not ( \4396_b0 , w_13959 );
and ( w_13959 , w_13958 , \4396_b1 );
or ( \4398_b1 , \4200_b1 , w_13961 );
not ( w_13961 , w_13962 );
and ( \4398_b0 , \4200_b0 , w_13963 );
and ( w_13962 ,  , w_13963 );
buf ( w_13961 , \4351_b1 );
not ( w_13961 , w_13964 );
not (  , w_13965 );
and ( w_13964 , w_13965 , \4351_b0 );
or ( \4399_b1 , \4397_b1 , w_13967 );
not ( w_13967 , w_13968 );
and ( \4399_b0 , \4397_b0 , w_13969 );
and ( w_13968 ,  , w_13969 );
buf ( w_13967 , \4398_b1 );
not ( w_13967 , w_13970 );
not (  , w_13971 );
and ( w_13970 , w_13971 , \4398_b0 );
or ( \4400_b1 , \4386_b1 , \4399_b1 );
xor ( \4400_b0 , \4386_b0 , w_13972 );
not ( w_13972 , w_13973 );
and ( w_13973 , \4399_b1 , \4399_b0 );
buf ( \4401_b1 , \4159_b1 );
not ( \4401_b1 , w_13974 );
not ( \4401_b0 , w_13975 );
and ( w_13974 , w_13975 , \4159_b0 );
buf ( \4402_b1 , \4094_b1 );
not ( \4402_b1 , w_13976 );
not ( \4402_b0 , w_13977 );
and ( w_13976 , w_13977 , \4094_b0 );
buf ( \4403_b1 , \4163_b1 );
not ( \4403_b1 , w_13978 );
not ( \4403_b0 , w_13979 );
and ( w_13978 , w_13979 , \4163_b0 );
or ( \4404_b1 , \4402_b1 , w_13980 );
or ( \4404_b0 , \4402_b0 , \4403_b0 );
not ( \4403_b0 , w_13981 );
and ( w_13981 , w_13980 , \4403_b1 );
or ( \4405_b1 , \4170_b1 , w_13983 );
not ( w_13983 , w_13984 );
and ( \4405_b0 , \4170_b0 , w_13985 );
and ( w_13984 ,  , w_13985 );
buf ( w_13983 , \4298_b1 );
not ( w_13983 , w_13986 );
not (  , w_13987 );
and ( w_13986 , w_13987 , \4298_b0 );
or ( \4406_b1 , \4404_b1 , w_13989 );
not ( w_13989 , w_13990 );
and ( \4406_b0 , \4404_b0 , w_13991 );
and ( w_13990 ,  , w_13991 );
buf ( w_13989 , \4405_b1 );
not ( w_13989 , w_13992 );
not (  , w_13993 );
and ( w_13992 , w_13993 , \4405_b0 );
buf ( \4407_b1 , \4406_b1 );
not ( \4407_b1 , w_13994 );
not ( \4407_b0 , w_13995 );
and ( w_13994 , w_13995 , \4406_b0 );
or ( \4408_b1 , \4401_b1 , w_13996 );
or ( \4408_b0 , \4401_b0 , \4407_b0 );
not ( \4407_b0 , w_13997 );
and ( w_13997 , w_13996 , \4407_b1 );
or ( \4409_b1 , \4150_b1 , w_13999 );
not ( w_13999 , w_14000 );
and ( \4409_b0 , \4150_b0 , w_14001 );
and ( w_14000 ,  , w_14001 );
buf ( w_13999 , \4313_b1 );
not ( w_13999 , w_14002 );
not (  , w_14003 );
and ( w_14002 , w_14003 , \4313_b0 );
or ( \4410_b1 , \4408_b1 , w_14005 );
not ( w_14005 , w_14006 );
and ( \4410_b0 , \4408_b0 , w_14007 );
and ( w_14006 ,  , w_14007 );
buf ( w_14005 , \4409_b1 );
not ( w_14005 , w_14008 );
not (  , w_14009 );
and ( w_14008 , w_14009 , \4409_b0 );
or ( \4411_b1 , \4400_b1 , \4410_b1 );
not ( \4410_b1 , w_14010 );
and ( \4411_b0 , \4400_b0 , w_14011 );
and ( w_14010 , w_14011 , \4410_b0 );
or ( \4412_b1 , \4386_b1 , \4399_b1 );
not ( \4399_b1 , w_14012 );
and ( \4412_b0 , \4386_b0 , w_14013 );
and ( w_14012 , w_14013 , \4399_b0 );
or ( \4413_b1 , \4411_b1 , w_14014 );
or ( \4413_b0 , \4411_b0 , \4412_b0 );
not ( \4412_b0 , w_14015 );
and ( w_14015 , w_14014 , \4412_b1 );
buf ( \4414_b1 , \4413_b1 );
not ( \4414_b1 , w_14016 );
not ( \4414_b0 , w_14017 );
and ( w_14016 , w_14017 , \4413_b0 );
or ( \4415_b1 , \4385_b1 , w_14018 );
or ( \4415_b0 , \4385_b0 , \4414_b0 );
not ( \4414_b0 , w_14019 );
and ( w_14019 , w_14018 , \4414_b1 );
buf ( \4416_b1 , \4319_b1 );
not ( \4416_b1 , w_14020 );
not ( \4416_b0 , w_14021 );
and ( w_14020 , w_14021 , \4319_b0 );
or ( \4417_b1 , \4416_b1 , w_14023 );
not ( w_14023 , w_14024 );
and ( \4417_b0 , \4416_b0 , w_14025 );
and ( w_14024 ,  , w_14025 );
buf ( w_14023 , \4382_b1 );
not ( w_14023 , w_14026 );
not (  , w_14027 );
and ( w_14026 , w_14027 , \4382_b0 );
or ( \4418_b1 , \4415_b1 , w_14029 );
not ( w_14029 , w_14030 );
and ( \4418_b0 , \4415_b0 , w_14031 );
and ( w_14030 ,  , w_14031 );
buf ( w_14029 , \4417_b1 );
not ( w_14029 , w_14032 );
not (  , w_14033 );
and ( w_14032 , w_14033 , \4417_b0 );
or ( \4419_b1 , \4329_b1 , \4359_b1 );
xor ( \4419_b0 , \4329_b0 , w_14034 );
not ( w_14034 , w_14035 );
and ( w_14035 , \4359_b1 , \4359_b0 );
or ( \4420_b1 , \4419_b1 , \4362_b1 );
xor ( \4420_b0 , \4419_b0 , w_14036 );
not ( w_14036 , w_14037 );
and ( w_14037 , \4362_b1 , \4362_b0 );
or ( \4421_b1 , \4418_b1 , \4420_b1 );
xor ( \4421_b0 , \4418_b0 , w_14038 );
not ( w_14038 , w_14039 );
and ( w_14039 , \4420_b1 , \4420_b0 );
or ( \4422_b1 , \4330_b1 , \4343_b1 );
xor ( \4422_b0 , \4330_b0 , w_14040 );
not ( w_14040 , w_14041 );
and ( w_14041 , \4343_b1 , \4343_b0 );
or ( \4423_b1 , \4422_b1 , \4356_b1 );
xor ( \4423_b0 , \4422_b0 , w_14042 );
not ( w_14042 , w_14043 );
and ( w_14043 , \4356_b1 , \4356_b0 );
buf ( \4424_b1 , \3997_b1 );
not ( \4424_b1 , w_14044 );
not ( \4424_b0 , w_14045 );
and ( w_14044 , w_14045 , \3997_b0 );
buf ( \4425_b1 , \4332_b1 );
not ( \4425_b1 , w_14046 );
not ( \4425_b0 , w_14047 );
and ( w_14046 , w_14047 , \4332_b0 );
or ( \4426_b1 , \4424_b1 , w_14048 );
or ( \4426_b0 , \4424_b0 , \4425_b0 );
not ( \4425_b0 , w_14049 );
and ( w_14049 , w_14048 , \4425_b1 );
or ( \4427_b1 , \4283_b1 , w_14051 );
not ( w_14051 , w_14052 );
and ( \4427_b0 , \4283_b0 , w_14053 );
and ( w_14052 ,  , w_14053 );
buf ( w_14051 , \4111_b1 );
not ( w_14051 , w_14054 );
not (  , w_14055 );
and ( w_14054 , w_14055 , \4111_b0 );
or ( \4428_b1 , \4426_b1 , w_14057 );
not ( w_14057 , w_14058 );
and ( \4428_b0 , \4426_b0 , w_14059 );
and ( w_14058 ,  , w_14059 );
buf ( w_14057 , \4427_b1 );
not ( w_14057 , w_14060 );
not (  , w_14061 );
and ( w_14060 , w_14061 , \4427_b0 );
buf ( \4429_b1 , \4428_b1 );
not ( \4429_b1 , w_14062 );
not ( \4429_b0 , w_14063 );
and ( w_14062 , w_14063 , \4428_b0 );
buf ( \4430_b1 , \4279_b1 );
buf ( \4430_b0 , \4279_b0 );
buf ( \4431_b1 , \4430_b1 );
not ( \4431_b1 , w_14064 );
not ( \4431_b0 , w_14065 );
and ( w_14064 , w_14065 , \4430_b0 );
or ( \4432_b1 , \4429_b1 , w_14066 );
or ( \4432_b0 , \4429_b0 , \4431_b0 );
not ( \4431_b0 , w_14067 );
and ( w_14067 , w_14066 , \4431_b1 );
or ( \4433_b1 , \4341_b1 , w_14069 );
not ( w_14069 , w_14070 );
and ( \4433_b0 , \4341_b0 , w_14071 );
and ( w_14070 ,  , w_14071 );
buf ( w_14069 , \4336_b1 );
not ( w_14069 , w_14072 );
not (  , w_14073 );
and ( w_14072 , w_14073 , \4336_b0 );
or ( \4434_b1 , \4432_b1 , w_14075 );
not ( w_14075 , w_14076 );
and ( \4434_b0 , \4432_b0 , w_14077 );
and ( w_14076 ,  , w_14077 );
buf ( w_14075 , \4433_b1 );
not ( w_14075 , w_14078 );
not (  , w_14079 );
and ( w_14078 , w_14079 , \4433_b0 );
buf ( \4435_b1 , \3326_b1 );
not ( \4435_b1 , w_14080 );
not ( \4435_b0 , w_14081 );
and ( w_14080 , w_14081 , \3326_b0 );
buf ( \4436_b1 , \4435_b1 );
not ( \4436_b1 , w_14082 );
not ( \4436_b0 , w_14083 );
and ( w_14082 , w_14083 , \4435_b0 );
buf ( \4437_b1 , \3387_b1 );
not ( \4437_b1 , w_14084 );
not ( \4437_b0 , w_14085 );
and ( w_14084 , w_14085 , \3387_b0 );
or ( \4438_b1 , \4436_b1 , \4437_b1 );
not ( \4437_b1 , w_14086 );
and ( \4438_b0 , \4436_b0 , w_14087 );
and ( w_14086 , w_14087 , \4437_b0 );
or ( \4439_b1 , \3387_b1 , \4435_b1 );
not ( \4435_b1 , w_14088 );
and ( \4439_b0 , \3387_b0 , w_14089 );
and ( w_14088 , w_14089 , \4435_b0 );
or ( \4440_b1 , \4438_b1 , w_14091 );
not ( w_14091 , w_14092 );
and ( \4440_b0 , \4438_b0 , w_14093 );
and ( w_14092 ,  , w_14093 );
buf ( w_14091 , \4439_b1 );
not ( w_14091 , w_14094 );
not (  , w_14095 );
and ( w_14094 , w_14095 , \4439_b0 );
buf ( \4441_b1 , \3387_b1 );
not ( \4441_b1 , w_14096 );
not ( \4441_b0 , w_14097 );
and ( w_14096 , w_14097 , \3387_b0 );
buf ( \4442_b1 , \3448_b1 );
not ( \4442_b1 , w_14098 );
not ( \4442_b0 , w_14099 );
and ( w_14098 , w_14099 , \3448_b0 );
buf ( \4443_b1 , \4442_b1 );
not ( \4443_b1 , w_14100 );
not ( \4443_b0 , w_14101 );
and ( w_14100 , w_14101 , \4442_b0 );
or ( \4444_b1 , \4441_b1 , w_14102 );
or ( \4444_b0 , \4441_b0 , \4443_b0 );
not ( \4443_b0 , w_14103 );
and ( w_14103 , w_14102 , \4443_b1 );
buf ( \4445_b1 , \3387_b1 );
not ( \4445_b1 , w_14104 );
not ( \4445_b0 , w_14105 );
and ( w_14104 , w_14105 , \3387_b0 );
or ( \4446_b1 , \4445_b1 , w_14107 );
not ( w_14107 , w_14108 );
and ( \4446_b0 , \4445_b0 , w_14109 );
and ( w_14108 ,  , w_14109 );
buf ( w_14107 , \3448_b1 );
not ( w_14107 , w_14110 );
not (  , w_14111 );
and ( w_14110 , w_14111 , \3448_b0 );
or ( \4447_b1 , \4444_b1 , w_14113 );
not ( w_14113 , w_14114 );
and ( \4447_b0 , \4444_b0 , w_14115 );
and ( w_14114 ,  , w_14115 );
buf ( w_14113 , \4446_b1 );
not ( w_14113 , w_14116 );
not (  , w_14117 );
and ( w_14116 , w_14117 , \4446_b0 );
or ( \4448_b1 , \4440_b1 , w_14119 );
not ( w_14119 , w_14120 );
and ( \4448_b0 , \4440_b0 , w_14121 );
and ( w_14120 ,  , w_14121 );
buf ( w_14119 , \4447_b1 );
not ( w_14119 , w_14122 );
not (  , w_14123 );
and ( w_14122 , w_14123 , \4447_b0 );
buf ( \4449_b1 , \4448_b1 );
buf ( \4449_b0 , \4448_b0 );
buf ( \4450_b1 , \4449_b1 );
not ( \4450_b1 , w_14124 );
not ( \4450_b0 , w_14125 );
and ( w_14124 , w_14125 , \4449_b0 );
buf ( \4451_b1 , \4450_b1 );
not ( \4451_b1 , w_14126 );
not ( \4451_b0 , w_14127 );
and ( w_14126 , w_14127 , \4450_b0 );
buf ( \4452_b1 , \4447_b1 );
buf ( \4452_b0 , \4447_b0 );
buf ( \4453_b1 , \4452_b1 );
buf ( \4453_b0 , \4452_b0 );
buf ( \4454_b1 , \4453_b1 );
not ( \4454_b1 , w_14128 );
not ( \4454_b0 , w_14129 );
and ( w_14128 , w_14129 , \4453_b0 );
buf ( \4455_b1 , \4454_b1 );
not ( \4455_b1 , w_14130 );
not ( \4455_b0 , w_14131 );
and ( w_14130 , w_14131 , \4454_b0 );
or ( \4456_b1 , \4451_b1 , w_14132 );
or ( \4456_b0 , \4451_b0 , \4455_b0 );
not ( \4455_b0 , w_14133 );
and ( w_14133 , w_14132 , \4455_b1 );
buf ( \4457_b1 , \4435_b1 );
buf ( \4457_b0 , \4435_b0 );
buf ( \4458_b1 , \4457_b1 );
not ( \4458_b1 , w_14134 );
not ( \4458_b0 , w_14135 );
and ( w_14134 , w_14135 , \4457_b0 );
or ( \4459_b1 , \4456_b1 , w_14137 );
not ( w_14137 , w_14138 );
and ( \4459_b0 , \4456_b0 , w_14139 );
and ( w_14138 ,  , w_14139 );
buf ( w_14137 , \4458_b1 );
not ( w_14137 , w_14140 );
not (  , w_14141 );
and ( w_14140 , w_14141 , \4458_b0 );
or ( \4460_b1 , \4434_b1 , \4459_b1 );
xor ( \4460_b0 , \4434_b0 , w_14142 );
not ( w_14142 , w_14143 );
and ( w_14143 , \4459_b1 , \4459_b0 );
or ( \4461_b1 , \4097_b1 , \4107_b1 );
not ( \4107_b1 , w_14144 );
and ( \4461_b0 , \4097_b0 , w_14145 );
and ( w_14144 , w_14145 , \4107_b0 );
buf ( \4462_b1 , \4097_b1 );
not ( \4462_b1 , w_14146 );
not ( \4462_b0 , w_14147 );
and ( w_14146 , w_14147 , \4097_b0 );
or ( \4463_b1 , \4462_b1 , \4106_b1 );
not ( \4106_b1 , w_14148 );
and ( \4463_b0 , \4462_b0 , w_14149 );
and ( w_14148 , w_14149 , \4106_b0 );
or ( \4464_b1 , \4461_b1 , w_14151 );
not ( w_14151 , w_14152 );
and ( \4464_b0 , \4461_b0 , w_14153 );
and ( w_14152 ,  , w_14153 );
buf ( w_14151 , \4463_b1 );
not ( w_14151 , w_14154 );
not (  , w_14155 );
and ( w_14154 , w_14155 , \4463_b0 );
buf ( \4465_b1 , \4464_b1 );
not ( \4465_b1 , w_14156 );
not ( \4465_b0 , w_14157 );
and ( w_14156 , w_14157 , \4464_b0 );
buf ( \4466_b1 , \4465_b1 );
not ( \4466_b1 , w_14158 );
not ( \4466_b0 , w_14159 );
and ( w_14158 , w_14159 , \4465_b0 );
buf ( \4467_b1 , \4129_b1 );
not ( \4467_b1 , w_14160 );
not ( \4467_b0 , w_14161 );
and ( w_14160 , w_14161 , \4129_b0 );
or ( \4468_b1 , \4466_b1 , w_14162 );
or ( \4468_b0 , \4466_b0 , \4467_b0 );
not ( \4467_b0 , w_14163 );
and ( w_14163 , w_14162 , \4467_b1 );
or ( \4469_b1 , \4133_b1 , w_14165 );
not ( w_14165 , w_14166 );
and ( \4469_b0 , \4133_b0 , w_14167 );
and ( w_14166 ,  , w_14167 );
buf ( w_14165 , \4377_b1 );
not ( w_14165 , w_14168 );
not (  , w_14169 );
and ( w_14168 , w_14169 , \4377_b0 );
or ( \4470_b1 , \4468_b1 , w_14171 );
not ( w_14171 , w_14172 );
and ( \4470_b0 , \4468_b0 , w_14173 );
and ( w_14172 ,  , w_14173 );
buf ( w_14171 , \4469_b1 );
not ( w_14171 , w_14174 );
not (  , w_14175 );
and ( w_14174 , w_14175 , \4469_b0 );
or ( \4471_b1 , \4460_b1 , \4470_b1 );
not ( \4470_b1 , w_14176 );
and ( \4471_b0 , \4460_b0 , w_14177 );
and ( w_14176 , w_14177 , \4470_b0 );
or ( \4472_b1 , \4434_b1 , \4459_b1 );
not ( \4459_b1 , w_14178 );
and ( \4472_b0 , \4434_b0 , w_14179 );
and ( w_14178 , w_14179 , \4459_b0 );
or ( \4473_b1 , \4471_b1 , w_14180 );
or ( \4473_b0 , \4471_b0 , \4472_b0 );
not ( \4472_b0 , w_14181 );
and ( w_14181 , w_14180 , \4472_b1 );
or ( \4474_b1 , \4423_b1 , \4473_b1 );
xor ( \4474_b0 , \4423_b0 , w_14182 );
not ( w_14182 , w_14183 );
and ( w_14183 , \4473_b1 , \4473_b0 );
buf ( \4475_b1 , \4382_b1 );
not ( \4475_b1 , w_14184 );
not ( \4475_b0 , w_14185 );
and ( w_14184 , w_14185 , \4382_b0 );
buf ( \4476_b1 , \4319_b1 );
not ( \4476_b1 , w_14186 );
not ( \4476_b0 , w_14187 );
and ( w_14186 , w_14187 , \4319_b0 );
or ( \4477_b1 , \4475_b1 , \4476_b1 );
not ( \4476_b1 , w_14188 );
and ( \4477_b0 , \4475_b0 , w_14189 );
and ( w_14188 , w_14189 , \4476_b0 );
or ( \4478_b1 , \4382_b1 , \4319_b1 );
not ( \4319_b1 , w_14190 );
and ( \4478_b0 , \4382_b0 , w_14191 );
and ( w_14190 , w_14191 , \4319_b0 );
or ( \4479_b1 , \4477_b1 , w_14193 );
not ( w_14193 , w_14194 );
and ( \4479_b0 , \4477_b0 , w_14195 );
and ( w_14194 ,  , w_14195 );
buf ( w_14193 , \4478_b1 );
not ( w_14193 , w_14196 );
not (  , w_14197 );
and ( w_14196 , w_14197 , \4478_b0 );
buf ( \4480_b1 , \4479_b1 );
not ( \4480_b1 , w_14198 );
not ( \4480_b0 , w_14199 );
and ( w_14198 , w_14199 , \4479_b0 );
buf ( \4481_b1 , \4413_b1 );
not ( \4481_b1 , w_14200 );
not ( \4481_b0 , w_14201 );
and ( w_14200 , w_14201 , \4413_b0 );
or ( \4482_b1 , \4480_b1 , w_14202 );
or ( \4482_b0 , \4480_b0 , \4481_b0 );
not ( \4481_b0 , w_14203 );
and ( w_14203 , w_14202 , \4481_b1 );
or ( \4483_b1 , \4413_b1 , w_14204 );
or ( \4483_b0 , \4413_b0 , \4479_b0 );
not ( \4479_b0 , w_14205 );
and ( w_14205 , w_14204 , \4479_b1 );
or ( \4484_b1 , \4482_b1 , w_14207 );
not ( w_14207 , w_14208 );
and ( \4484_b0 , \4482_b0 , w_14209 );
and ( w_14208 ,  , w_14209 );
buf ( w_14207 , \4483_b1 );
not ( w_14207 , w_14210 );
not (  , w_14211 );
and ( w_14210 , w_14211 , \4483_b0 );
or ( \4485_b1 , \4474_b1 , \4484_b1 );
not ( \4484_b1 , w_14212 );
and ( \4485_b0 , \4474_b0 , w_14213 );
and ( w_14212 , w_14213 , \4484_b0 );
or ( \4486_b1 , \4423_b1 , \4473_b1 );
not ( \4473_b1 , w_14214 );
and ( \4486_b0 , \4423_b0 , w_14215 );
and ( w_14214 , w_14215 , \4473_b0 );
or ( \4487_b1 , \4485_b1 , w_14216 );
or ( \4487_b0 , \4485_b0 , \4486_b0 );
not ( \4486_b0 , w_14217 );
and ( w_14217 , w_14216 , \4486_b1 );
or ( \4488_b1 , \4421_b1 , \4487_b1 );
xor ( \4488_b0 , \4421_b0 , w_14218 );
not ( w_14218 , w_14219 );
and ( w_14219 , \4487_b1 , \4487_b0 );
buf ( \4489_b1 , \4488_b1 );
not ( \4489_b1 , w_14220 );
not ( \4489_b0 , w_14221 );
and ( w_14220 , w_14221 , \4488_b0 );
or ( \4490_b1 , \4386_b1 , \4399_b1 );
xor ( \4490_b0 , \4386_b0 , w_14222 );
not ( w_14222 , w_14223 );
and ( w_14223 , \4399_b1 , \4399_b0 );
or ( \4491_b1 , \4490_b1 , \4410_b1 );
xor ( \4491_b0 , \4490_b0 , w_14224 );
not ( w_14224 , w_14225 );
and ( w_14225 , \4410_b1 , \4410_b0 );
buf ( \4492_b1 , \4198_b1 );
not ( \4492_b1 , w_14226 );
not ( \4492_b0 , w_14227 );
and ( w_14226 , w_14227 , \4198_b0 );
buf ( \4493_b1 , \4283_b1 );
not ( \4493_b1 , w_14228 );
not ( \4493_b0 , w_14229 );
and ( w_14228 , w_14229 , \4283_b0 );
buf ( \4494_b1 , \4493_b1 );
not ( \4494_b1 , w_14230 );
not ( \4494_b0 , w_14231 );
and ( w_14230 , w_14231 , \4493_b0 );
or ( \4495_b1 , \4492_b1 , w_14232 );
or ( \4495_b0 , \4492_b0 , \4494_b0 );
not ( \4494_b0 , w_14233 );
and ( w_14233 , w_14232 , \4494_b1 );
or ( \4496_b1 , \4285_b1 , w_14235 );
not ( w_14235 , w_14236 );
and ( \4496_b0 , \4285_b0 , w_14237 );
and ( w_14236 ,  , w_14237 );
buf ( w_14235 , \4209_b1 );
not ( w_14235 , w_14238 );
not (  , w_14239 );
and ( w_14238 , w_14239 , \4209_b0 );
or ( \4497_b1 , \4495_b1 , w_14241 );
not ( w_14241 , w_14242 );
and ( \4497_b0 , \4495_b0 , w_14243 );
and ( w_14242 ,  , w_14243 );
buf ( w_14241 , \4496_b1 );
not ( w_14241 , w_14244 );
not (  , w_14245 );
and ( w_14244 , w_14245 , \4496_b0 );
buf ( \4498_b1 , \4497_b1 );
not ( \4498_b1 , w_14246 );
not ( \4498_b0 , w_14247 );
and ( w_14246 , w_14247 , \4497_b0 );
buf ( \4499_b1 , \4338_b1 );
not ( \4499_b1 , w_14248 );
not ( \4499_b0 , w_14249 );
and ( w_14248 , w_14249 , \4338_b0 );
or ( \4500_b1 , \4498_b1 , w_14250 );
or ( \4500_b0 , \4498_b0 , \4499_b0 );
not ( \4499_b0 , w_14251 );
and ( w_14251 , w_14250 , \4499_b1 );
or ( \4501_b1 , \4341_b1 , w_14253 );
not ( w_14253 , w_14254 );
and ( \4501_b0 , \4341_b0 , w_14255 );
and ( w_14254 ,  , w_14255 );
buf ( w_14253 , \4428_b1 );
not ( w_14253 , w_14256 );
not (  , w_14257 );
and ( w_14256 , w_14257 , \4428_b0 );
or ( \4502_b1 , \4500_b1 , w_14259 );
not ( w_14259 , w_14260 );
and ( \4502_b0 , \4500_b0 , w_14261 );
and ( w_14260 ,  , w_14261 );
buf ( w_14259 , \4501_b1 );
not ( w_14259 , w_14262 );
not (  , w_14263 );
and ( w_14262 , w_14263 , \4501_b0 );
or ( \4503_b1 , \4491_b1 , w_14264 );
or ( \4503_b0 , \4491_b0 , \4502_b0 );
not ( \4502_b0 , w_14265 );
and ( w_14265 , w_14264 , \4502_b1 );
or ( \4504_b1 , \4093_b1 , \4134_b1 );
not ( \4134_b1 , w_14266 );
and ( \4504_b0 , \4093_b0 , w_14267 );
and ( w_14266 , w_14267 , \4134_b0 );
buf ( \4505_b1 , \4093_b1 );
not ( \4505_b1 , w_14268 );
not ( \4505_b0 , w_14269 );
and ( w_14268 , w_14269 , \4093_b0 );
or ( \4506_b1 , \4505_b1 , \4106_b1 );
not ( \4106_b1 , w_14270 );
and ( \4506_b0 , \4505_b0 , w_14271 );
and ( w_14270 , w_14271 , \4106_b0 );
or ( \4507_b1 , \4504_b1 , w_14273 );
not ( w_14273 , w_14274 );
and ( \4507_b0 , \4504_b0 , w_14275 );
and ( w_14274 ,  , w_14275 );
buf ( w_14273 , \4506_b1 );
not ( w_14273 , w_14276 );
not (  , w_14277 );
and ( w_14276 , w_14277 , \4506_b0 );
buf ( \4508_b1 , \4507_b1 );
not ( \4508_b1 , w_14278 );
not ( \4508_b0 , w_14279 );
and ( w_14278 , w_14279 , \4507_b0 );
buf ( \4509_b1 , \4127_b1 );
not ( \4509_b1 , w_14280 );
not ( \4509_b0 , w_14281 );
and ( w_14280 , w_14281 , \4127_b0 );
or ( \4510_b1 , \4508_b1 , \4509_b1 );
not ( \4509_b1 , w_14282 );
and ( \4510_b0 , \4508_b0 , w_14283 );
and ( w_14282 , w_14283 , \4509_b0 );
buf ( \4511_b1 , \4132_b1 );
not ( \4511_b1 , w_14284 );
not ( \4511_b0 , w_14285 );
and ( w_14284 , w_14285 , \4132_b0 );
or ( \4512_b1 , \4511_b1 , w_14287 );
not ( w_14287 , w_14288 );
and ( \4512_b0 , \4511_b0 , w_14289 );
and ( w_14288 ,  , w_14289 );
buf ( w_14287 , \4464_b1 );
not ( w_14287 , w_14290 );
not (  , w_14291 );
and ( w_14290 , w_14291 , \4464_b0 );
or ( \4513_b1 , \4510_b1 , w_14293 );
not ( w_14293 , w_14294 );
and ( \4513_b0 , \4510_b0 , w_14295 );
and ( w_14294 ,  , w_14295 );
buf ( w_14293 , \4512_b1 );
not ( w_14293 , w_14296 );
not (  , w_14297 );
and ( w_14296 , w_14297 , \4512_b0 );
buf ( \4514_b1 , \4513_b1 );
not ( \4514_b1 , w_14298 );
not ( \4514_b0 , w_14299 );
and ( w_14298 , w_14299 , \4513_b0 );
buf ( \4515_b1 , \4514_b1 );
not ( \4515_b1 , w_14300 );
not ( \4515_b0 , w_14301 );
and ( w_14300 , w_14301 , \4514_b0 );
buf ( \4516_b1 , \4066_b1 );
not ( \4516_b1 , w_14302 );
not ( \4516_b0 , w_14303 );
and ( w_14302 , w_14303 , \4066_b0 );
buf ( \4517_b1 , \4388_b1 );
not ( \4517_b1 , w_14304 );
not ( \4517_b0 , w_14305 );
and ( w_14304 , w_14305 , \4388_b0 );
or ( \4518_b1 , \4516_b1 , w_14306 );
or ( \4518_b0 , \4516_b0 , \4517_b0 );
not ( \4517_b0 , w_14307 );
and ( w_14307 , w_14306 , \4517_b1 );
buf ( \4519_b1 , \4066_b1 );
not ( \4519_b1 , w_14308 );
not ( \4519_b0 , w_14309 );
and ( w_14308 , w_14309 , \4066_b0 );
or ( \4520_b1 , \4100_b1 , w_14311 );
not ( w_14311 , w_14312 );
and ( \4520_b0 , \4100_b0 , w_14313 );
and ( w_14312 ,  , w_14313 );
buf ( w_14311 , \4519_b1 );
not ( w_14311 , w_14314 );
not (  , w_14315 );
and ( w_14314 , w_14315 , \4519_b0 );
or ( \4521_b1 , \4518_b1 , w_14317 );
not ( w_14317 , w_14318 );
and ( \4521_b0 , \4518_b0 , w_14319 );
and ( w_14318 ,  , w_14319 );
buf ( w_14317 , \4520_b1 );
not ( w_14317 , w_14320 );
not (  , w_14321 );
and ( w_14320 , w_14321 , \4520_b0 );
buf ( \4522_b1 , \4521_b1 );
not ( \4522_b1 , w_14322 );
not ( \4522_b0 , w_14323 );
and ( w_14322 , w_14323 , \4521_b0 );
buf ( \4523_b1 , \4193_b1 );
not ( \4523_b1 , w_14324 );
not ( \4523_b0 , w_14325 );
and ( w_14324 , w_14325 , \4193_b0 );
buf ( \4524_b1 , \4523_b1 );
not ( \4524_b1 , w_14326 );
not ( \4524_b0 , w_14327 );
and ( w_14326 , w_14327 , \4523_b0 );
or ( \4525_b1 , \4522_b1 , w_14328 );
or ( \4525_b0 , \4522_b0 , \4524_b0 );
not ( \4524_b0 , w_14329 );
and ( w_14329 , w_14328 , \4524_b1 );
or ( \4526_b1 , \4393_b1 , w_14331 );
not ( w_14331 , w_14332 );
and ( \4526_b0 , \4393_b0 , w_14333 );
and ( w_14332 ,  , w_14333 );
buf ( w_14331 , \4200_b1 );
not ( w_14331 , w_14334 );
not (  , w_14335 );
and ( w_14334 , w_14335 , \4200_b0 );
or ( \4527_b1 , \4525_b1 , w_14337 );
not ( w_14337 , w_14338 );
and ( \4527_b0 , \4525_b0 , w_14339 );
and ( w_14338 ,  , w_14339 );
buf ( w_14337 , \4526_b1 );
not ( w_14337 , w_14340 );
not (  , w_14341 );
and ( w_14340 , w_14341 , \4526_b0 );
buf ( \4528_b1 , \4527_b1 );
not ( \4528_b1 , w_14342 );
not ( \4528_b0 , w_14343 );
and ( w_14342 , w_14343 , \4527_b0 );
or ( \4529_b1 , \4515_b1 , w_14344 );
or ( \4529_b0 , \4515_b0 , \4528_b0 );
not ( \4528_b0 , w_14345 );
and ( w_14345 , w_14344 , \4528_b1 );
or ( \4530_b1 , \4514_b1 , w_14346 );
or ( \4530_b0 , \4514_b0 , \4527_b0 );
not ( \4527_b0 , w_14347 );
and ( w_14347 , w_14346 , \4527_b1 );
buf ( \4531_b1 , \4051_b1 );
not ( \4531_b1 , w_14348 );
not ( \4531_b0 , w_14349 );
and ( w_14348 , w_14349 , \4051_b0 );
buf ( \4532_b1 , \4458_b1 );
not ( \4532_b1 , w_14350 );
not ( \4532_b0 , w_14351 );
and ( w_14350 , w_14351 , \4458_b0 );
buf ( \4533_b1 , \4532_b1 );
not ( \4533_b1 , w_14352 );
not ( \4533_b0 , w_14353 );
and ( w_14352 , w_14353 , \4532_b0 );
or ( \4534_b1 , \4531_b1 , w_14354 );
or ( \4534_b0 , \4531_b0 , \4533_b0 );
not ( \4533_b0 , w_14355 );
and ( w_14355 , w_14354 , \4533_b1 );
buf ( \4535_b1 , \4436_b1 );
not ( \4535_b1 , w_14356 );
not ( \4535_b0 , w_14357 );
and ( w_14356 , w_14357 , \4436_b0 );
buf ( \4536_b1 , \4535_b1 );
not ( \4536_b1 , w_14358 );
not ( \4536_b0 , w_14359 );
and ( w_14358 , w_14359 , \4535_b0 );
or ( \4537_b1 , \4536_b1 , w_14361 );
not ( w_14361 , w_14362 );
and ( \4537_b0 , \4536_b0 , w_14363 );
and ( w_14362 ,  , w_14363 );
buf ( w_14361 , \4135_b1 );
not ( w_14361 , w_14364 );
not (  , w_14365 );
and ( w_14364 , w_14365 , \4135_b0 );
or ( \4538_b1 , \4534_b1 , w_14367 );
not ( w_14367 , w_14368 );
and ( \4538_b0 , \4534_b0 , w_14369 );
and ( w_14368 ,  , w_14369 );
buf ( w_14367 , \4537_b1 );
not ( w_14367 , w_14370 );
not (  , w_14371 );
and ( w_14370 , w_14371 , \4537_b0 );
buf ( \4539_b1 , \4538_b1 );
not ( \4539_b1 , w_14372 );
not ( \4539_b0 , w_14373 );
and ( w_14372 , w_14373 , \4538_b0 );
buf ( \4540_b1 , \4450_b1 );
not ( \4540_b1 , w_14374 );
not ( \4540_b0 , w_14375 );
and ( w_14374 , w_14375 , \4450_b0 );
buf ( \4541_b1 , \4540_b1 );
not ( \4541_b1 , w_14376 );
not ( \4541_b0 , w_14377 );
and ( w_14376 , w_14377 , \4540_b0 );
or ( \4542_b1 , \4539_b1 , w_14378 );
or ( \4542_b0 , \4539_b0 , \4541_b0 );
not ( \4541_b0 , w_14379 );
and ( w_14379 , w_14378 , \4541_b1 );
buf ( \4543_b1 , \4532_b1 );
not ( \4543_b1 , w_14380 );
not ( \4543_b0 , w_14381 );
and ( w_14380 , w_14381 , \4532_b0 );
or ( \4544_b1 , \4543_b1 , w_14383 );
not ( w_14383 , w_14384 );
and ( \4544_b0 , \4543_b0 , w_14385 );
and ( w_14384 ,  , w_14385 );
buf ( w_14383 , \4453_b1 );
not ( w_14383 , w_14386 );
not (  , w_14387 );
and ( w_14386 , w_14387 , \4453_b0 );
or ( \4545_b1 , \4542_b1 , w_14389 );
not ( w_14389 , w_14390 );
and ( \4545_b0 , \4542_b0 , w_14391 );
and ( w_14390 ,  , w_14391 );
buf ( w_14389 , \4544_b1 );
not ( w_14389 , w_14392 );
not (  , w_14393 );
and ( w_14392 , w_14393 , \4544_b0 );
or ( \4546_b1 , \4530_b1 , w_14395 );
not ( w_14395 , w_14396 );
and ( \4546_b0 , \4530_b0 , w_14397 );
and ( w_14396 ,  , w_14397 );
buf ( w_14395 , \4545_b1 );
not ( w_14395 , w_14398 );
not (  , w_14399 );
and ( w_14398 , w_14399 , \4545_b0 );
or ( \4547_b1 , \4529_b1 , w_14401 );
not ( w_14401 , w_14402 );
and ( \4547_b0 , \4529_b0 , w_14403 );
and ( w_14402 ,  , w_14403 );
buf ( w_14401 , \4546_b1 );
not ( w_14401 , w_14404 );
not (  , w_14405 );
and ( w_14404 , w_14405 , \4546_b0 );
or ( \4548_b1 , \4503_b1 , w_14407 );
not ( w_14407 , w_14408 );
and ( \4548_b0 , \4503_b0 , w_14409 );
and ( w_14408 ,  , w_14409 );
buf ( w_14407 , \4547_b1 );
not ( w_14407 , w_14410 );
not (  , w_14411 );
and ( w_14410 , w_14411 , \4547_b0 );
or ( \4549_b1 , \4491_b1 , w_14413 );
not ( w_14413 , w_14414 );
and ( \4549_b0 , \4491_b0 , w_14415 );
and ( w_14414 ,  , w_14415 );
buf ( w_14413 , \4502_b1 );
not ( w_14413 , w_14416 );
not (  , w_14417 );
and ( w_14416 , w_14417 , \4502_b0 );
or ( \4550_b1 , \4548_b1 , w_14419 );
not ( w_14419 , w_14420 );
and ( \4550_b0 , \4548_b0 , w_14421 );
and ( w_14420 ,  , w_14421 );
buf ( w_14419 , \4549_b1 );
not ( w_14419 , w_14422 );
not (  , w_14423 );
and ( w_14422 , w_14423 , \4549_b0 );
or ( \4551_b1 , \4423_b1 , \4473_b1 );
xor ( \4551_b0 , \4423_b0 , w_14424 );
not ( w_14424 , w_14425 );
and ( w_14425 , \4473_b1 , \4473_b0 );
or ( \4552_b1 , \4551_b1 , \4484_b1 );
xor ( \4552_b0 , \4551_b0 , w_14426 );
not ( w_14426 , w_14427 );
and ( w_14427 , \4484_b1 , \4484_b0 );
or ( \4553_b1 , \4550_b1 , \4552_b1 );
xor ( \4553_b0 , \4550_b0 , w_14428 );
not ( w_14428 , w_14429 );
and ( w_14429 , \4552_b1 , \4552_b0 );
or ( \4554_b1 , \4434_b1 , \4459_b1 );
xor ( \4554_b0 , \4434_b0 , w_14430 );
not ( w_14430 , w_14431 );
and ( w_14431 , \4459_b1 , \4459_b0 );
or ( \4555_b1 , \4554_b1 , \4470_b1 );
xor ( \4555_b0 , \4554_b0 , w_14432 );
not ( w_14432 , w_14433 );
and ( w_14433 , \4470_b1 , \4470_b0 );
buf ( \4556_b1 , \4555_b1 );
not ( \4556_b1 , w_14434 );
not ( \4556_b0 , w_14435 );
and ( w_14434 , w_14435 , \4555_b0 );
buf ( \4557_b1 , \4096_b1 );
not ( \4557_b1 , w_14436 );
not ( \4557_b0 , w_14437 );
and ( w_14436 , w_14437 , \4096_b0 );
buf ( \4558_b1 , \4163_b1 );
not ( \4558_b1 , w_14438 );
not ( \4558_b0 , w_14439 );
and ( w_14438 , w_14439 , \4163_b0 );
or ( \4559_b1 , \4557_b1 , w_14440 );
or ( \4559_b0 , \4557_b0 , \4558_b0 );
not ( \4558_b0 , w_14441 );
and ( w_14441 , w_14440 , \4558_b1 );
or ( \4560_b1 , \4170_b1 , w_14443 );
not ( w_14443 , w_14444 );
and ( \4560_b0 , \4170_b0 , w_14445 );
and ( w_14444 ,  , w_14445 );
buf ( w_14443 , \4372_b1 );
not ( w_14443 , w_14446 );
not (  , w_14447 );
and ( w_14446 , w_14447 , \4372_b0 );
or ( \4561_b1 , \4559_b1 , w_14449 );
not ( w_14449 , w_14450 );
and ( \4561_b0 , \4559_b0 , w_14451 );
and ( w_14450 ,  , w_14451 );
buf ( w_14449 , \4560_b1 );
not ( w_14449 , w_14452 );
not (  , w_14453 );
and ( w_14452 , w_14453 , \4560_b0 );
buf ( \4562_b1 , \4561_b1 );
not ( \4562_b1 , w_14454 );
not ( \4562_b0 , w_14455 );
and ( w_14454 , w_14455 , \4561_b0 );
buf ( \4563_b1 , \4159_b1 );
not ( \4563_b1 , w_14456 );
not ( \4563_b0 , w_14457 );
and ( w_14456 , w_14457 , \4159_b0 );
or ( \4564_b1 , \4562_b1 , w_14458 );
or ( \4564_b0 , \4562_b0 , \4563_b0 );
not ( \4563_b0 , w_14459 );
and ( w_14459 , w_14458 , \4563_b1 );
or ( \4565_b1 , \4150_b1 , w_14461 );
not ( w_14461 , w_14462 );
and ( \4565_b0 , \4150_b0 , w_14463 );
and ( w_14462 ,  , w_14463 );
buf ( w_14461 , \4406_b1 );
not ( w_14461 , w_14464 );
not (  , w_14465 );
and ( w_14464 , w_14465 , \4406_b0 );
or ( \4566_b1 , \4564_b1 , w_14467 );
not ( w_14467 , w_14468 );
and ( \4566_b0 , \4564_b0 , w_14469 );
and ( w_14468 ,  , w_14469 );
buf ( w_14467 , \4565_b1 );
not ( w_14467 , w_14470 );
not (  , w_14471 );
and ( w_14470 , w_14471 , \4565_b0 );
buf ( \4567_b1 , \4566_b1 );
not ( \4567_b1 , w_14472 );
not ( \4567_b0 , w_14473 );
and ( w_14472 , w_14473 , \4566_b0 );
or ( \4568_b1 , \4102_b1 , w_14475 );
not ( w_14475 , w_14476 );
and ( \4568_b0 , \4102_b0 , w_14477 );
and ( w_14476 ,  , w_14477 );
buf ( w_14475 , \4017_b1 );
not ( w_14475 , w_14478 );
not (  , w_14479 );
and ( w_14478 , w_14479 , \4017_b0 );
or ( \4569_b1 , \4567_b1 , w_14481 );
not ( w_14481 , w_14482 );
and ( \4569_b0 , \4567_b0 , w_14483 );
and ( w_14482 ,  , w_14483 );
buf ( w_14481 , \4568_b1 );
not ( w_14481 , w_14484 );
not (  , w_14485 );
and ( w_14484 , w_14485 , \4568_b0 );
buf ( \4570_b1 , \4502_b1 );
not ( \4570_b1 , w_14486 );
not ( \4570_b0 , w_14487 );
and ( w_14486 , w_14487 , \4502_b0 );
or ( \4571_b1 , \4569_b1 , \4570_b1 );
not ( \4570_b1 , w_14488 );
and ( \4571_b0 , \4569_b0 , w_14489 );
and ( w_14488 , w_14489 , \4570_b0 );
or ( \4572_b1 , \4567_b1 , w_14491 );
not ( w_14491 , w_14492 );
and ( \4572_b0 , \4567_b0 , w_14493 );
and ( w_14492 ,  , w_14493 );
buf ( w_14491 , \4568_b1 );
not ( w_14491 , w_14494 );
not (  , w_14495 );
and ( w_14494 , w_14495 , \4568_b0 );
or ( \4573_b1 , \4571_b1 , w_14497 );
not ( w_14497 , w_14498 );
and ( \4573_b0 , \4571_b0 , w_14499 );
and ( w_14498 ,  , w_14499 );
buf ( w_14497 , \4572_b1 );
not ( w_14497 , w_14500 );
not (  , w_14501 );
and ( w_14500 , w_14501 , \4572_b0 );
or ( \4574_b1 , \4556_b1 , w_14503 );
not ( w_14503 , w_14504 );
and ( \4574_b0 , \4556_b0 , w_14505 );
and ( w_14504 ,  , w_14505 );
buf ( w_14503 , \4573_b1 );
not ( w_14503 , w_14506 );
not (  , w_14507 );
and ( w_14506 , w_14507 , \4573_b0 );
buf ( \4575_b1 , \4574_b1 );
not ( \4575_b1 , w_14508 );
not ( \4575_b0 , w_14509 );
and ( w_14508 , w_14509 , \4574_b0 );
or ( \4576_b1 , \4502_b1 , \4547_b1 );
xor ( \4576_b0 , \4502_b0 , w_14510 );
not ( w_14510 , w_14511 );
and ( w_14511 , \4547_b1 , \4547_b0 );
or ( \4577_b1 , \4576_b1 , w_14512 );
xor ( \4577_b0 , \4576_b0 , w_14514 );
not ( w_14514 , w_14515 );
and ( w_14515 , w_14512 , w_14513 );
buf ( w_14512 , \4491_b1 );
not ( w_14512 , w_14516 );
not ( w_14513 , w_14517 );
and ( w_14516 , w_14517 , \4491_b0 );
buf ( \4578_b1 , \4577_b1 );
not ( \4578_b1 , w_14518 );
not ( \4578_b0 , w_14519 );
and ( w_14518 , w_14519 , \4577_b0 );
buf ( \4579_b1 , \4578_b1 );
not ( \4579_b1 , w_14520 );
not ( \4579_b0 , w_14521 );
and ( w_14520 , w_14521 , \4578_b0 );
or ( \4580_b1 , \4575_b1 , w_14522 );
or ( \4580_b0 , \4575_b0 , \4579_b0 );
not ( \4579_b0 , w_14523 );
and ( w_14523 , w_14522 , \4579_b1 );
buf ( \4581_b1 , \4573_b1 );
not ( \4581_b1 , w_14524 );
not ( \4581_b0 , w_14525 );
and ( w_14524 , w_14525 , \4573_b0 );
or ( \4582_b1 , \4581_b1 , w_14527 );
not ( w_14527 , w_14528 );
and ( \4582_b0 , \4581_b0 , w_14529 );
and ( w_14528 ,  , w_14529 );
buf ( w_14527 , \4555_b1 );
not ( w_14527 , w_14530 );
not (  , w_14531 );
and ( w_14530 , w_14531 , \4555_b0 );
or ( \4583_b1 , \4580_b1 , w_14533 );
not ( w_14533 , w_14534 );
and ( \4583_b0 , \4580_b0 , w_14535 );
and ( w_14534 ,  , w_14535 );
buf ( w_14533 , \4582_b1 );
not ( w_14533 , w_14536 );
not (  , w_14537 );
and ( w_14536 , w_14537 , \4582_b0 );
or ( \4584_b1 , \4553_b1 , \4583_b1 );
not ( \4583_b1 , w_14538 );
and ( \4584_b0 , \4553_b0 , w_14539 );
and ( w_14538 , w_14539 , \4583_b0 );
or ( \4585_b1 , \4550_b1 , \4552_b1 );
not ( \4552_b1 , w_14540 );
and ( \4585_b0 , \4550_b0 , w_14541 );
and ( w_14540 , w_14541 , \4552_b0 );
or ( \4586_b1 , \4584_b1 , w_14542 );
or ( \4586_b0 , \4584_b0 , \4585_b0 );
not ( \4585_b0 , w_14543 );
and ( w_14543 , w_14542 , \4585_b1 );
buf ( \4587_b1 , \4586_b1 );
not ( \4587_b1 , w_14544 );
not ( \4587_b0 , w_14545 );
and ( w_14544 , w_14545 , \4586_b0 );
or ( \4588_b1 , \4489_b1 , w_14547 );
not ( w_14547 , w_14548 );
and ( \4588_b0 , \4489_b0 , w_14549 );
and ( w_14548 ,  , w_14549 );
buf ( w_14547 , \4587_b1 );
not ( w_14547 , w_14550 );
not (  , w_14551 );
and ( w_14550 , w_14551 , \4587_b0 );
buf ( \4589_b1 , \4588_b1 );
buf ( \4589_b0 , \4588_b0 );
buf ( \4590_b1 , \4589_b1 );
not ( \4590_b1 , w_14552 );
not ( \4590_b0 , w_14553 );
and ( w_14552 , w_14553 , \4589_b0 );
buf ( \4591_b1 , \4513_b1 );
not ( \4591_b1 , w_14554 );
not ( \4591_b0 , w_14555 );
and ( w_14554 , w_14555 , \4513_b0 );
buf ( \4592_b1 , \4527_b1 );
not ( \4592_b1 , w_14556 );
not ( \4592_b0 , w_14557 );
and ( w_14556 , w_14557 , \4527_b0 );
or ( \4593_b1 , \4591_b1 , w_14558 );
or ( \4593_b0 , \4591_b0 , \4592_b0 );
not ( \4592_b0 , w_14559 );
and ( w_14559 , w_14558 , \4592_b1 );
or ( \4594_b1 , \4527_b1 , w_14560 );
or ( \4594_b0 , \4527_b0 , \4513_b0 );
not ( \4513_b0 , w_14561 );
and ( w_14561 , w_14560 , \4513_b1 );
or ( \4595_b1 , \4593_b1 , w_14563 );
not ( w_14563 , w_14564 );
and ( \4595_b0 , \4593_b0 , w_14565 );
and ( w_14564 ,  , w_14565 );
buf ( w_14563 , \4594_b1 );
not ( w_14563 , w_14566 );
not (  , w_14567 );
and ( w_14566 , w_14567 , \4594_b0 );
or ( \4596_b1 , \4595_b1 , \4545_b1 );
xor ( \4596_b0 , \4595_b0 , w_14568 );
not ( w_14568 , w_14569 );
and ( w_14569 , \4545_b1 , \4545_b0 );
buf ( \4597_b1 , \3516_b1 );
not ( \4597_b1 , w_14570 );
not ( \4597_b0 , w_14571 );
and ( w_14570 , w_14571 , \3516_b0 );
or ( \4598_b1 , \2945_b1 , \4597_b1 );
not ( \4597_b1 , w_14572 );
and ( \4598_b0 , \2945_b0 , w_14573 );
and ( w_14572 , w_14573 , \4597_b0 );
buf ( \4599_b1 , \2945_b1 );
not ( \4599_b1 , w_14574 );
not ( \4599_b0 , w_14575 );
and ( w_14574 , w_14575 , \2945_b0 );
or ( \4600_b1 , \4599_b1 , \3516_b1 );
not ( \3516_b1 , w_14576 );
and ( \4600_b0 , \4599_b0 , w_14577 );
and ( w_14576 , w_14577 , \3516_b0 );
or ( \4601_b1 , \4598_b1 , w_14579 );
not ( w_14579 , w_14580 );
and ( \4601_b0 , \4598_b0 , w_14581 );
and ( w_14580 ,  , w_14581 );
buf ( w_14579 , \4600_b1 );
not ( w_14579 , w_14582 );
not (  , w_14583 );
and ( w_14582 , w_14583 , \4600_b0 );
buf ( \4602_b1 , \4601_b1 );
buf ( \4602_b0 , \4601_b0 );
buf ( \4603_b1 , \4602_b1 );
not ( \4603_b1 , w_14584 );
not ( \4603_b0 , w_14585 );
and ( w_14584 , w_14585 , \4602_b0 );
buf ( \4604_b1 , \4442_b1 );
not ( \4604_b1 , w_14586 );
not ( \4604_b0 , w_14587 );
and ( w_14586 , w_14587 , \4442_b0 );
buf ( \4605_b1 , \3516_b1 );
not ( \4605_b1 , w_14588 );
not ( \4605_b0 , w_14589 );
and ( w_14588 , w_14589 , \3516_b0 );
or ( \4606_b1 , \4604_b1 , w_14590 );
or ( \4606_b0 , \4604_b0 , \4605_b0 );
not ( \4605_b0 , w_14591 );
and ( w_14591 , w_14590 , \4605_b1 );
or ( \4607_b1 , \4597_b1 , w_14593 );
not ( w_14593 , w_14594 );
and ( \4607_b0 , \4597_b0 , w_14595 );
and ( w_14594 ,  , w_14595 );
buf ( w_14593 , \3448_b1 );
not ( w_14593 , w_14596 );
not (  , w_14597 );
and ( w_14596 , w_14597 , \3448_b0 );
or ( \4608_b1 , \4606_b1 , w_14599 );
not ( w_14599 , w_14600 );
and ( \4608_b0 , \4606_b0 , w_14601 );
and ( w_14600 ,  , w_14601 );
buf ( w_14599 , \4607_b1 );
not ( w_14599 , w_14602 );
not (  , w_14603 );
and ( w_14602 , w_14603 , \4607_b0 );
or ( \4609_b1 , \4608_b1 , w_14605 );
not ( w_14605 , w_14606 );
and ( \4609_b0 , \4608_b0 , w_14607 );
and ( w_14606 ,  , w_14607 );
buf ( w_14605 , \4601_b1 );
not ( w_14605 , w_14608 );
not (  , w_14609 );
and ( w_14608 , w_14609 , \4601_b0 );
buf ( \4610_b1 , \4609_b1 );
not ( \4610_b1 , w_14610 );
not ( \4610_b0 , w_14611 );
and ( w_14610 , w_14611 , \4609_b0 );
buf ( \4611_b1 , \4610_b1 );
buf ( \4611_b0 , \4610_b0 );
buf ( \4612_b1 , \4611_b1 );
not ( \4612_b1 , w_14612 );
not ( \4612_b0 , w_14613 );
and ( w_14612 , w_14613 , \4611_b0 );
buf ( \4613_b1 , \4612_b1 );
not ( \4613_b1 , w_14614 );
not ( \4613_b0 , w_14615 );
and ( w_14614 , w_14615 , \4612_b0 );
or ( \4614_b1 , \4603_b1 , w_14616 );
or ( \4614_b0 , \4603_b0 , \4613_b0 );
not ( \4613_b0 , w_14617 );
and ( w_14617 , w_14616 , \4613_b1 );
buf ( \4615_b1 , \3448_b1 );
buf ( \4615_b0 , \3448_b0 );
buf ( \4616_b1 , \4615_b1 );
buf ( \4616_b0 , \4615_b0 );
or ( \4617_b1 , \4614_b1 , w_14619 );
not ( w_14619 , w_14620 );
and ( \4617_b0 , \4614_b0 , w_14621 );
and ( w_14620 ,  , w_14621 );
buf ( w_14619 , \4616_b1 );
not ( w_14619 , w_14622 );
not (  , w_14623 );
and ( w_14622 , w_14623 , \4616_b0 );
buf ( \4618_b1 , \4617_b1 );
not ( \4618_b1 , w_14624 );
not ( \4618_b0 , w_14625 );
and ( w_14624 , w_14625 , \4617_b0 );
buf ( \4619_b1 , \4159_b1 );
not ( \4619_b1 , w_14626 );
not ( \4619_b0 , w_14627 );
and ( w_14626 , w_14627 , \4159_b0 );
buf ( \4620_b1 , \4097_b1 );
not ( \4620_b1 , w_14628 );
not ( \4620_b0 , w_14629 );
and ( w_14628 , w_14629 , \4097_b0 );
buf ( \4621_b1 , \4163_b1 );
not ( \4621_b1 , w_14630 );
not ( \4621_b0 , w_14631 );
and ( w_14630 , w_14631 , \4163_b0 );
or ( \4622_b1 , \4620_b1 , w_14632 );
or ( \4622_b0 , \4620_b0 , \4621_b0 );
not ( \4621_b0 , w_14633 );
and ( w_14633 , w_14632 , \4621_b1 );
or ( \4623_b1 , \4170_b1 , w_14635 );
not ( w_14635 , w_14636 );
and ( \4623_b0 , \4170_b0 , w_14637 );
and ( w_14636 ,  , w_14637 );
buf ( w_14635 , \4254_b1 );
not ( w_14635 , w_14638 );
not (  , w_14639 );
and ( w_14638 , w_14639 , \4254_b0 );
or ( \4624_b1 , \4622_b1 , w_14641 );
not ( w_14641 , w_14642 );
and ( \4624_b0 , \4622_b0 , w_14643 );
and ( w_14642 ,  , w_14643 );
buf ( w_14641 , \4623_b1 );
not ( w_14641 , w_14644 );
not (  , w_14645 );
and ( w_14644 , w_14645 , \4623_b0 );
buf ( \4625_b1 , \4624_b1 );
not ( \4625_b1 , w_14646 );
not ( \4625_b0 , w_14647 );
and ( w_14646 , w_14647 , \4624_b0 );
or ( \4626_b1 , \4619_b1 , w_14648 );
or ( \4626_b0 , \4619_b0 , \4625_b0 );
not ( \4625_b0 , w_14649 );
and ( w_14649 , w_14648 , \4625_b1 );
or ( \4627_b1 , \4561_b1 , w_14651 );
not ( w_14651 , w_14652 );
and ( \4627_b0 , \4561_b0 , w_14653 );
and ( w_14652 ,  , w_14653 );
buf ( w_14651 , \4150_b1 );
not ( w_14651 , w_14654 );
not (  , w_14655 );
and ( w_14654 , w_14655 , \4150_b0 );
or ( \4628_b1 , \4626_b1 , w_14657 );
not ( w_14657 , w_14658 );
and ( \4628_b0 , \4626_b0 , w_14659 );
and ( w_14658 ,  , w_14659 );
buf ( w_14657 , \4627_b1 );
not ( w_14657 , w_14660 );
not (  , w_14661 );
and ( w_14660 , w_14661 , \4627_b0 );
buf ( \4629_b1 , \4628_b1 );
not ( \4629_b1 , w_14662 );
not ( \4629_b0 , w_14663 );
and ( w_14662 , w_14663 , \4628_b0 );
or ( \4630_b1 , \4618_b1 , w_14664 );
or ( \4630_b0 , \4618_b0 , \4629_b0 );
not ( \4629_b0 , w_14665 );
and ( w_14665 , w_14664 , \4629_b1 );
or ( \4631_b1 , \4628_b1 , w_14666 );
or ( \4631_b0 , \4628_b0 , \4617_b0 );
not ( \4617_b0 , w_14667 );
and ( w_14667 , w_14666 , \4617_b1 );
buf ( \4632_b1 , \4449_b1 );
buf ( \4632_b0 , \4449_b0 );
buf ( \4633_b1 , \3997_b1 );
not ( \4633_b1 , w_14668 );
not ( \4633_b0 , w_14669 );
and ( w_14668 , w_14669 , \3997_b0 );
buf ( \4634_b1 , \4535_b1 );
not ( \4634_b1 , w_14670 );
not ( \4634_b0 , w_14671 );
and ( w_14670 , w_14671 , \4535_b0 );
or ( \4635_b1 , \4633_b1 , w_14672 );
or ( \4635_b0 , \4633_b0 , \4634_b0 );
not ( \4634_b0 , w_14673 );
and ( w_14673 , w_14672 , \4634_b1 );
or ( \4636_b1 , \4536_b1 , w_14675 );
not ( w_14675 , w_14676 );
and ( \4636_b0 , \4536_b0 , w_14677 );
and ( w_14676 ,  , w_14677 );
buf ( w_14675 , \4111_b1 );
not ( w_14675 , w_14678 );
not (  , w_14679 );
and ( w_14678 , w_14679 , \4111_b0 );
or ( \4637_b1 , \4635_b1 , w_14681 );
not ( w_14681 , w_14682 );
and ( \4637_b0 , \4635_b0 , w_14683 );
and ( w_14682 ,  , w_14683 );
buf ( w_14681 , \4636_b1 );
not ( w_14681 , w_14684 );
not (  , w_14685 );
and ( w_14684 , w_14685 , \4636_b0 );
or ( \4638_b1 , \4632_b1 , \4637_b1 );
not ( \4637_b1 , w_14686 );
and ( \4638_b0 , \4632_b0 , w_14687 );
and ( w_14686 , w_14687 , \4637_b0 );
or ( \4639_b1 , \4538_b1 , \4453_b1 );
not ( \4453_b1 , w_14688 );
and ( \4639_b0 , \4538_b0 , w_14689 );
and ( w_14688 , w_14689 , \4453_b0 );
or ( \4640_b1 , \4638_b1 , w_14691 );
not ( w_14691 , w_14692 );
and ( \4640_b0 , \4638_b0 , w_14693 );
and ( w_14692 ,  , w_14693 );
buf ( w_14691 , \4639_b1 );
not ( w_14691 , w_14694 );
not (  , w_14695 );
and ( w_14694 , w_14695 , \4639_b0 );
buf ( \4641_b1 , \4640_b1 );
not ( \4641_b1 , w_14696 );
not ( \4641_b0 , w_14697 );
and ( w_14696 , w_14697 , \4640_b0 );
or ( \4642_b1 , \4631_b1 , w_14699 );
not ( w_14699 , w_14700 );
and ( \4642_b0 , \4631_b0 , w_14701 );
and ( w_14700 ,  , w_14701 );
buf ( w_14699 , \4641_b1 );
not ( w_14699 , w_14702 );
not (  , w_14703 );
and ( w_14702 , w_14703 , \4641_b0 );
or ( \4643_b1 , \4630_b1 , w_14705 );
not ( w_14705 , w_14706 );
and ( \4643_b0 , \4630_b0 , w_14707 );
and ( w_14706 ,  , w_14707 );
buf ( w_14705 , \4642_b1 );
not ( w_14705 , w_14708 );
not (  , w_14709 );
and ( w_14708 , w_14709 , \4642_b0 );
or ( \4644_b1 , \4596_b1 , \4643_b1 );
xor ( \4644_b0 , \4596_b0 , w_14710 );
not ( w_14710 , w_14711 );
and ( w_14711 , \4643_b1 , \4643_b0 );
buf ( \4645_b1 , \4095_b1 );
not ( \4645_b1 , w_14712 );
not ( \4645_b0 , w_14713 );
and ( w_14712 , w_14713 , \4095_b0 );
buf ( \4646_b1 , \4134_b1 );
not ( \4646_b1 , w_14714 );
not ( \4646_b0 , w_14715 );
and ( w_14714 , w_14715 , \4134_b0 );
or ( \4647_b1 , \4645_b1 , w_14716 );
or ( \4647_b0 , \4645_b0 , \4646_b0 );
not ( \4646_b0 , w_14717 );
and ( w_14717 , w_14716 , \4646_b1 );
or ( \4648_b1 , \4106_b1 , w_14719 );
not ( w_14719 , w_14720 );
and ( \4648_b0 , \4106_b0 , w_14721 );
and ( w_14720 ,  , w_14721 );
buf ( w_14719 , \4391_b1 );
not ( w_14719 , w_14722 );
not (  , w_14723 );
and ( w_14722 , w_14723 , \4391_b0 );
or ( \4649_b1 , \4647_b1 , w_14725 );
not ( w_14725 , w_14726 );
and ( \4649_b0 , \4647_b0 , w_14727 );
and ( w_14726 ,  , w_14727 );
buf ( w_14725 , \4648_b1 );
not ( w_14725 , w_14728 );
not (  , w_14729 );
and ( w_14728 , w_14729 , \4648_b0 );
buf ( \4650_b1 , \4649_b1 );
not ( \4650_b1 , w_14730 );
not ( \4650_b0 , w_14731 );
and ( w_14730 , w_14731 , \4649_b0 );
buf ( \4651_b1 , \4302_b1 );
not ( \4651_b1 , w_14732 );
not ( \4651_b0 , w_14733 );
and ( w_14732 , w_14733 , \4302_b0 );
or ( \4652_b1 , \4650_b1 , w_14734 );
or ( \4652_b0 , \4650_b0 , \4651_b0 );
not ( \4651_b0 , w_14735 );
and ( w_14735 , w_14734 , \4651_b1 );
buf ( \4653_b1 , \4507_b1 );
not ( \4653_b1 , w_14736 );
not ( \4653_b0 , w_14737 );
and ( w_14736 , w_14737 , \4507_b0 );
buf ( \4654_b1 , \4511_b1 );
not ( \4654_b1 , w_14738 );
not ( \4654_b0 , w_14739 );
and ( w_14738 , w_14739 , \4511_b0 );
or ( \4655_b1 , \4653_b1 , w_14741 );
not ( w_14741 , w_14742 );
and ( \4655_b0 , \4653_b0 , w_14743 );
and ( w_14742 ,  , w_14743 );
buf ( w_14741 , \4654_b1 );
not ( w_14741 , w_14744 );
not (  , w_14745 );
and ( w_14744 , w_14745 , \4654_b0 );
or ( \4656_b1 , \4652_b1 , w_14747 );
not ( w_14747 , w_14748 );
and ( \4656_b0 , \4652_b0 , w_14749 );
and ( w_14748 ,  , w_14749 );
buf ( w_14747 , \4655_b1 );
not ( w_14747 , w_14750 );
not (  , w_14751 );
and ( w_14750 , w_14751 , \4655_b0 );
buf ( \4657_b1 , \4395_b1 );
not ( \4657_b1 , w_14752 );
not ( \4657_b0 , w_14753 );
and ( w_14752 , w_14753 , \4395_b0 );
buf ( \4658_b1 , \4017_b1 );
not ( \4658_b1 , w_14754 );
not ( \4658_b0 , w_14755 );
and ( w_14754 , w_14755 , \4017_b0 );
buf ( \4659_b1 , \4101_b1 );
not ( \4659_b1 , w_14756 );
not ( \4659_b0 , w_14757 );
and ( w_14756 , w_14757 , \4101_b0 );
or ( \4660_b1 , \4658_b1 , w_14758 );
or ( \4660_b0 , \4658_b0 , \4659_b0 );
not ( \4659_b0 , w_14759 );
and ( w_14759 , w_14758 , \4659_b1 );
buf ( \4661_b1 , \4346_b1 );
not ( \4661_b1 , w_14760 );
not ( \4661_b0 , w_14761 );
and ( w_14760 , w_14761 , \4346_b0 );
buf ( \4662_b1 , \4017_b1 );
not ( \4662_b1 , w_14762 );
not ( \4662_b0 , w_14763 );
and ( w_14762 , w_14763 , \4017_b0 );
or ( \4663_b1 , \4661_b1 , w_14765 );
not ( w_14765 , w_14766 );
and ( \4663_b0 , \4661_b0 , w_14767 );
and ( w_14766 ,  , w_14767 );
buf ( w_14765 , \4662_b1 );
not ( w_14765 , w_14768 );
not (  , w_14769 );
and ( w_14768 , w_14769 , \4662_b0 );
or ( \4664_b1 , \4660_b1 , w_14771 );
not ( w_14771 , w_14772 );
and ( \4664_b0 , \4660_b0 , w_14773 );
and ( w_14772 ,  , w_14773 );
buf ( w_14771 , \4663_b1 );
not ( w_14771 , w_14774 );
not (  , w_14775 );
and ( w_14774 , w_14775 , \4663_b0 );
buf ( \4665_b1 , \4664_b1 );
not ( \4665_b1 , w_14776 );
not ( \4665_b0 , w_14777 );
and ( w_14776 , w_14777 , \4664_b0 );
or ( \4666_b1 , \4657_b1 , w_14778 );
or ( \4666_b0 , \4657_b0 , \4665_b0 );
not ( \4665_b0 , w_14779 );
and ( w_14779 , w_14778 , \4665_b1 );
or ( \4667_b1 , \4521_b1 , w_14781 );
not ( w_14781 , w_14782 );
and ( \4667_b0 , \4521_b0 , w_14783 );
and ( w_14782 ,  , w_14783 );
buf ( w_14781 , \4200_b1 );
not ( w_14781 , w_14784 );
not (  , w_14785 );
and ( w_14784 , w_14785 , \4200_b0 );
or ( \4668_b1 , \4666_b1 , w_14787 );
not ( w_14787 , w_14788 );
and ( \4668_b0 , \4666_b0 , w_14789 );
and ( w_14788 ,  , w_14789 );
buf ( w_14787 , \4667_b1 );
not ( w_14787 , w_14790 );
not (  , w_14791 );
and ( w_14790 , w_14791 , \4667_b0 );
or ( \4669_b1 , \4656_b1 , w_14792 );
or ( \4669_b0 , \4656_b0 , \4668_b0 );
not ( \4668_b0 , w_14793 );
and ( w_14793 , w_14792 , \4668_b1 );
buf ( \4670_b1 , \4094_b1 );
not ( \4670_b1 , w_14794 );
not ( \4670_b0 , w_14795 );
and ( w_14794 , w_14795 , \4094_b0 );
buf ( \4671_b1 , \4284_b1 );
not ( \4671_b1 , w_14796 );
not ( \4671_b0 , w_14797 );
and ( w_14796 , w_14797 , \4284_b0 );
or ( \4672_b1 , \4670_b1 , w_14798 );
or ( \4672_b0 , \4670_b0 , \4671_b0 );
not ( \4671_b0 , w_14799 );
and ( w_14799 , w_14798 , \4671_b1 );
buf ( \4673_b1 , \4332_b1 );
not ( \4673_b1 , w_14800 );
not ( \4673_b0 , w_14801 );
and ( w_14800 , w_14801 , \4332_b0 );
or ( \4674_b1 , \4673_b1 , w_14803 );
not ( w_14803 , w_14804 );
and ( \4674_b0 , \4673_b0 , w_14805 );
and ( w_14804 ,  , w_14805 );
buf ( w_14803 , \4298_b1 );
not ( w_14803 , w_14806 );
not (  , w_14807 );
and ( w_14806 , w_14807 , \4298_b0 );
or ( \4675_b1 , \4672_b1 , w_14809 );
not ( w_14809 , w_14810 );
and ( \4675_b0 , \4672_b0 , w_14811 );
and ( w_14810 ,  , w_14811 );
buf ( w_14809 , \4674_b1 );
not ( w_14809 , w_14812 );
not (  , w_14813 );
and ( w_14812 , w_14813 , \4674_b0 );
buf ( \4676_b1 , \4675_b1 );
not ( \4676_b1 , w_14814 );
not ( \4676_b0 , w_14815 );
and ( w_14814 , w_14815 , \4675_b0 );
buf ( \4677_b1 , \4430_b1 );
not ( \4677_b1 , w_14816 );
not ( \4677_b0 , w_14817 );
and ( w_14816 , w_14817 , \4430_b0 );
or ( \4678_b1 , \4676_b1 , w_14818 );
or ( \4678_b0 , \4676_b0 , \4677_b0 );
not ( \4677_b0 , w_14819 );
and ( w_14819 , w_14818 , \4677_b1 );
or ( \4679_b1 , \4497_b1 , w_14821 );
not ( w_14821 , w_14822 );
and ( \4679_b0 , \4497_b0 , w_14823 );
and ( w_14822 ,  , w_14823 );
buf ( w_14821 , \4341_b1 );
not ( w_14821 , w_14824 );
not (  , w_14825 );
and ( w_14824 , w_14825 , \4341_b0 );
or ( \4680_b1 , \4678_b1 , w_14827 );
not ( w_14827 , w_14828 );
and ( \4680_b0 , \4678_b0 , w_14829 );
and ( w_14828 ,  , w_14829 );
buf ( w_14827 , \4679_b1 );
not ( w_14827 , w_14830 );
not (  , w_14831 );
and ( w_14830 , w_14831 , \4679_b0 );
or ( \4681_b1 , \4669_b1 , w_14833 );
not ( w_14833 , w_14834 );
and ( \4681_b0 , \4669_b0 , w_14835 );
and ( w_14834 ,  , w_14835 );
buf ( w_14833 , \4680_b1 );
not ( w_14833 , w_14836 );
not (  , w_14837 );
and ( w_14836 , w_14837 , \4680_b0 );
buf ( \4682_b1 , \4656_b1 );
not ( \4682_b1 , w_14838 );
not ( \4682_b0 , w_14839 );
and ( w_14838 , w_14839 , \4656_b0 );
buf ( \4683_b1 , \4682_b1 );
not ( \4683_b1 , w_14840 );
not ( \4683_b0 , w_14841 );
and ( w_14840 , w_14841 , \4682_b0 );
or ( \4684_b1 , \4683_b1 , w_14843 );
not ( w_14843 , w_14844 );
and ( \4684_b0 , \4683_b0 , w_14845 );
and ( w_14844 ,  , w_14845 );
buf ( w_14843 , \4668_b1 );
not ( w_14843 , w_14846 );
not (  , w_14847 );
and ( w_14846 , w_14847 , \4668_b0 );
or ( \4685_b1 , \4681_b1 , w_14849 );
not ( w_14849 , w_14850 );
and ( \4685_b0 , \4681_b0 , w_14851 );
and ( w_14850 ,  , w_14851 );
buf ( w_14849 , \4684_b1 );
not ( w_14849 , w_14852 );
not (  , w_14853 );
and ( w_14852 , w_14853 , \4684_b0 );
or ( \4686_b1 , \4644_b1 , \4685_b1 );
not ( \4685_b1 , w_14854 );
and ( \4686_b0 , \4644_b0 , w_14855 );
and ( w_14854 , w_14855 , \4685_b0 );
or ( \4687_b1 , \4596_b1 , \4643_b1 );
not ( \4643_b1 , w_14856 );
and ( \4687_b0 , \4596_b0 , w_14857 );
and ( w_14856 , w_14857 , \4643_b0 );
or ( \4688_b1 , \4686_b1 , w_14858 );
or ( \4688_b0 , \4686_b0 , \4687_b0 );
not ( \4687_b0 , w_14859 );
and ( w_14859 , w_14858 , \4687_b1 );
buf ( \4689_b1 , \4573_b1 );
not ( \4689_b1 , w_14860 );
not ( \4689_b0 , w_14861 );
and ( w_14860 , w_14861 , \4573_b0 );
buf ( \4690_b1 , \4555_b1 );
not ( \4690_b1 , w_14862 );
not ( \4690_b0 , w_14863 );
and ( w_14862 , w_14863 , \4555_b0 );
or ( \4691_b1 , \4689_b1 , w_14864 );
or ( \4691_b0 , \4689_b0 , \4690_b0 );
not ( \4690_b0 , w_14865 );
and ( w_14865 , w_14864 , \4690_b1 );
or ( \4692_b1 , \4573_b1 , w_14866 );
or ( \4692_b0 , \4573_b0 , \4555_b0 );
not ( \4555_b0 , w_14867 );
and ( w_14867 , w_14866 , \4555_b1 );
or ( \4693_b1 , \4691_b1 , w_14869 );
not ( w_14869 , w_14870 );
and ( \4693_b0 , \4691_b0 , w_14871 );
and ( w_14870 ,  , w_14871 );
buf ( w_14869 , \4692_b1 );
not ( w_14869 , w_14872 );
not (  , w_14873 );
and ( w_14872 , w_14873 , \4692_b0 );
buf ( \4694_b1 , \4693_b1 );
not ( \4694_b1 , w_14874 );
not ( \4694_b0 , w_14875 );
and ( w_14874 , w_14875 , \4693_b0 );
buf ( \4695_b1 , \4694_b1 );
not ( \4695_b1 , w_14876 );
not ( \4695_b0 , w_14877 );
and ( w_14876 , w_14877 , \4694_b0 );
buf ( \4696_b1 , \4578_b1 );
not ( \4696_b1 , w_14878 );
not ( \4696_b0 , w_14879 );
and ( w_14878 , w_14879 , \4578_b0 );
or ( \4697_b1 , \4695_b1 , w_14880 );
or ( \4697_b0 , \4695_b0 , \4696_b0 );
not ( \4696_b0 , w_14881 );
and ( w_14881 , w_14880 , \4696_b1 );
or ( \4698_b1 , \4577_b1 , w_14883 );
not ( w_14883 , w_14884 );
and ( \4698_b0 , \4577_b0 , w_14885 );
and ( w_14884 ,  , w_14885 );
buf ( w_14883 , \4693_b1 );
not ( w_14883 , w_14886 );
not (  , w_14887 );
and ( w_14886 , w_14887 , \4693_b0 );
or ( \4699_b1 , \4697_b1 , w_14889 );
not ( w_14889 , w_14890 );
and ( \4699_b0 , \4697_b0 , w_14891 );
and ( w_14890 ,  , w_14891 );
buf ( w_14889 , \4698_b1 );
not ( w_14889 , w_14892 );
not (  , w_14893 );
and ( w_14892 , w_14893 , \4698_b0 );
or ( \4700_b1 , \4688_b1 , \4699_b1 );
xor ( \4700_b0 , \4688_b0 , w_14894 );
not ( w_14894 , w_14895 );
and ( w_14895 , \4699_b1 , \4699_b0 );
or ( \4701_b1 , \4568_b1 , \4566_b1 );
xor ( \4701_b0 , \4568_b0 , w_14896 );
not ( w_14896 , w_14897 );
and ( w_14897 , \4566_b1 , \4566_b0 );
or ( \4702_b1 , \4701_b1 , w_14898 );
xor ( \4702_b0 , \4701_b0 , w_14900 );
not ( w_14900 , w_14901 );
and ( w_14901 , w_14898 , w_14899 );
buf ( w_14898 , \4570_b1 );
not ( w_14898 , w_14902 );
not ( w_14899 , w_14903 );
and ( w_14902 , w_14903 , \4570_b0 );
buf ( \4703_b1 , \4702_b1 );
not ( \4703_b1 , w_14904 );
not ( \4703_b0 , w_14905 );
and ( w_14904 , w_14905 , \4702_b0 );
buf ( \4704_b1 , \4066_b1 );
not ( \4704_b1 , w_14906 );
not ( \4704_b0 , w_14907 );
and ( w_14906 , w_14907 , \4066_b0 );
buf ( \4705_b1 , \4134_b1 );
not ( \4705_b1 , w_14908 );
not ( \4705_b0 , w_14909 );
and ( w_14908 , w_14909 , \4134_b0 );
or ( \4706_b1 , \4704_b1 , w_14910 );
or ( \4706_b0 , \4704_b0 , \4705_b0 );
not ( \4705_b0 , w_14911 );
and ( w_14911 , w_14910 , \4705_b1 );
or ( \4707_b1 , \4106_b1 , w_14913 );
not ( w_14913 , w_14914 );
and ( \4707_b0 , \4106_b0 , w_14915 );
and ( w_14914 ,  , w_14915 );
buf ( w_14913 , \4519_b1 );
not ( w_14913 , w_14916 );
not (  , w_14917 );
and ( w_14916 , w_14917 , \4519_b0 );
or ( \4708_b1 , \4706_b1 , w_14919 );
not ( w_14919 , w_14920 );
and ( \4708_b0 , \4706_b0 , w_14921 );
and ( w_14920 ,  , w_14921 );
buf ( w_14919 , \4707_b1 );
not ( w_14919 , w_14922 );
not (  , w_14923 );
and ( w_14922 , w_14923 , \4707_b0 );
buf ( \4709_b1 , \4708_b1 );
not ( \4709_b1 , w_14924 );
not ( \4709_b0 , w_14925 );
and ( w_14924 , w_14925 , \4708_b0 );
buf ( \4710_b1 , \4127_b1 );
not ( \4710_b1 , w_14926 );
not ( \4710_b0 , w_14927 );
and ( w_14926 , w_14927 , \4127_b0 );
buf ( \4711_b1 , \4710_b1 );
not ( \4711_b1 , w_14928 );
not ( \4711_b0 , w_14929 );
and ( w_14928 , w_14929 , \4710_b0 );
or ( \4712_b1 , \4709_b1 , w_14930 );
or ( \4712_b0 , \4709_b0 , \4711_b0 );
not ( \4711_b0 , w_14931 );
and ( w_14931 , w_14930 , \4711_b1 );
or ( \4713_b1 , \4654_b1 , w_14933 );
not ( w_14933 , w_14934 );
and ( \4713_b0 , \4654_b0 , w_14935 );
and ( w_14934 ,  , w_14935 );
buf ( w_14933 , \4649_b1 );
not ( w_14933 , w_14936 );
not (  , w_14937 );
and ( w_14936 , w_14937 , \4649_b0 );
or ( \4714_b1 , \4712_b1 , w_14939 );
not ( w_14939 , w_14940 );
and ( \4714_b0 , \4712_b0 , w_14941 );
and ( w_14940 ,  , w_14941 );
buf ( w_14939 , \4713_b1 );
not ( w_14939 , w_14942 );
not (  , w_14943 );
and ( w_14942 , w_14943 , \4713_b0 );
buf ( \4715_b1 , \4714_b1 );
not ( \4715_b1 , w_14944 );
not ( \4715_b0 , w_14945 );
and ( w_14944 , w_14945 , \4714_b0 );
buf ( \4716_b1 , \4093_b1 );
not ( \4716_b1 , w_14946 );
not ( \4716_b0 , w_14947 );
and ( w_14946 , w_14947 , \4093_b0 );
buf ( \4717_b1 , \4163_b1 );
not ( \4717_b1 , w_14948 );
not ( \4717_b0 , w_14949 );
and ( w_14948 , w_14949 , \4163_b0 );
or ( \4718_b1 , \4716_b1 , w_14950 );
or ( \4718_b0 , \4716_b0 , \4717_b0 );
not ( \4717_b0 , w_14951 );
and ( w_14951 , w_14950 , \4717_b1 );
or ( \4719_b1 , \4170_b1 , w_14953 );
not ( w_14953 , w_14954 );
and ( \4719_b0 , \4170_b0 , w_14955 );
and ( w_14954 ,  , w_14955 );
buf ( w_14953 , \4349_b1 );
not ( w_14953 , w_14956 );
not (  , w_14957 );
and ( w_14956 , w_14957 , \4349_b0 );
or ( \4720_b1 , \4718_b1 , w_14959 );
not ( w_14959 , w_14960 );
and ( \4720_b0 , \4718_b0 , w_14961 );
and ( w_14960 ,  , w_14961 );
buf ( w_14959 , \4719_b1 );
not ( w_14959 , w_14962 );
not (  , w_14963 );
and ( w_14962 , w_14963 , \4719_b0 );
buf ( \4721_b1 , \4720_b1 );
not ( \4721_b1 , w_14964 );
not ( \4721_b0 , w_14965 );
and ( w_14964 , w_14965 , \4720_b0 );
buf ( \4722_b1 , \4159_b1 );
not ( \4722_b1 , w_14966 );
not ( \4722_b0 , w_14967 );
and ( w_14966 , w_14967 , \4159_b0 );
or ( \4723_b1 , \4721_b1 , w_14968 );
or ( \4723_b0 , \4721_b0 , \4722_b0 );
not ( \4722_b0 , w_14969 );
and ( w_14969 , w_14968 , \4722_b1 );
or ( \4724_b1 , \4624_b1 , w_14971 );
not ( w_14971 , w_14972 );
and ( \4724_b0 , \4624_b0 , w_14973 );
and ( w_14972 ,  , w_14973 );
buf ( w_14971 , \4317_b1 );
not ( w_14971 , w_14974 );
not (  , w_14975 );
and ( w_14974 , w_14975 , \4317_b0 );
or ( \4725_b1 , \4723_b1 , w_14977 );
not ( w_14977 , w_14978 );
and ( \4725_b0 , \4723_b0 , w_14979 );
and ( w_14978 ,  , w_14979 );
buf ( w_14977 , \4724_b1 );
not ( w_14977 , w_14980 );
not (  , w_14981 );
and ( w_14980 , w_14981 , \4724_b0 );
buf ( \4726_b1 , \4725_b1 );
not ( \4726_b1 , w_14982 );
not ( \4726_b0 , w_14983 );
and ( w_14982 , w_14983 , \4725_b0 );
or ( \4727_b1 , \4715_b1 , w_14984 );
or ( \4727_b0 , \4715_b0 , \4726_b0 );
not ( \4726_b0 , w_14985 );
and ( w_14985 , w_14984 , \4726_b1 );
or ( \4728_b1 , \4714_b1 , w_14986 );
or ( \4728_b0 , \4714_b0 , \4725_b0 );
not ( \4725_b0 , w_14987 );
and ( w_14987 , w_14986 , \4725_b1 );
buf ( \4729_b1 , \4436_b1 );
buf ( \4729_b0 , \4436_b0 );
or ( \4730_b1 , \4198_b1 , \4729_b1 );
not ( \4729_b1 , w_14988 );
and ( \4730_b0 , \4198_b0 , w_14989 );
and ( w_14988 , w_14989 , \4729_b0 );
buf ( \4731_b1 , \4198_b1 );
not ( \4731_b1 , w_14990 );
not ( \4731_b0 , w_14991 );
and ( w_14990 , w_14991 , \4198_b0 );
buf ( \4732_b1 , \4457_b1 );
buf ( \4732_b0 , \4457_b0 );
or ( \4733_b1 , \4731_b1 , \4732_b1 );
not ( \4732_b1 , w_14992 );
and ( \4733_b0 , \4731_b0 , w_14993 );
and ( w_14992 , w_14993 , \4732_b0 );
or ( \4734_b1 , \4730_b1 , w_14995 );
not ( w_14995 , w_14996 );
and ( \4734_b0 , \4730_b0 , w_14997 );
and ( w_14996 ,  , w_14997 );
buf ( w_14995 , \4733_b1 );
not ( w_14995 , w_14998 );
not (  , w_14999 );
and ( w_14998 , w_14999 , \4733_b0 );
buf ( \4735_b1 , \4734_b1 );
not ( \4735_b1 , w_15000 );
not ( \4735_b0 , w_15001 );
and ( w_15000 , w_15001 , \4734_b0 );
buf ( \4736_b1 , \4540_b1 );
not ( \4736_b1 , w_15002 );
not ( \4736_b0 , w_15003 );
and ( w_15002 , w_15003 , \4540_b0 );
or ( \4737_b1 , \4735_b1 , w_15004 );
or ( \4737_b0 , \4735_b0 , \4736_b0 );
not ( \4736_b0 , w_15005 );
and ( w_15005 , w_15004 , \4736_b1 );
or ( \4738_b1 , \4637_b1 , w_15007 );
not ( w_15007 , w_15008 );
and ( \4738_b0 , \4637_b0 , w_15009 );
and ( w_15008 ,  , w_15009 );
buf ( w_15007 , \4453_b1 );
not ( w_15007 , w_15010 );
not (  , w_15011 );
and ( w_15010 , w_15011 , \4453_b0 );
or ( \4739_b1 , \4737_b1 , w_15013 );
not ( w_15013 , w_15014 );
and ( \4739_b0 , \4737_b0 , w_15015 );
and ( w_15014 ,  , w_15015 );
buf ( w_15013 , \4738_b1 );
not ( w_15013 , w_15016 );
not (  , w_15017 );
and ( w_15016 , w_15017 , \4738_b0 );
or ( \4740_b1 , \4728_b1 , w_15019 );
not ( w_15019 , w_15020 );
and ( \4740_b0 , \4728_b0 , w_15021 );
and ( w_15020 ,  , w_15021 );
buf ( w_15019 , \4739_b1 );
not ( w_15019 , w_15022 );
not (  , w_15023 );
and ( w_15022 , w_15023 , \4739_b0 );
or ( \4741_b1 , \4727_b1 , w_15025 );
not ( w_15025 , w_15026 );
and ( \4741_b0 , \4727_b0 , w_15027 );
and ( w_15026 ,  , w_15027 );
buf ( w_15025 , \4740_b1 );
not ( w_15025 , w_15028 );
not (  , w_15029 );
and ( w_15028 , w_15029 , \4740_b0 );
or ( \4742_b1 , \4102_b1 , \4021_b1 );
not ( \4021_b1 , w_15030 );
and ( \4742_b0 , \4102_b0 , w_15031 );
and ( w_15030 , w_15031 , \4021_b0 );
buf ( \4743_b1 , \4742_b1 );
not ( \4743_b1 , w_15032 );
not ( \4743_b0 , w_15033 );
and ( w_15032 , w_15033 , \4742_b0 );
buf ( \4744_b1 , \4051_b1 );
not ( \4744_b1 , w_15034 );
not ( \4744_b0 , w_15035 );
and ( w_15034 , w_15035 , \4051_b0 );
buf ( \4745_b1 , \3448_b1 );
buf ( \4745_b0 , \3448_b0 );
buf ( \4746_b1 , \4745_b1 );
not ( \4746_b1 , w_15036 );
not ( \4746_b0 , w_15037 );
and ( w_15036 , w_15037 , \4745_b0 );
buf ( \4747_b1 , \4746_b1 );
not ( \4747_b1 , w_15038 );
not ( \4747_b0 , w_15039 );
and ( w_15038 , w_15039 , \4746_b0 );
or ( \4748_b1 , \4744_b1 , w_15040 );
or ( \4748_b0 , \4744_b0 , \4747_b0 );
not ( \4747_b0 , w_15041 );
and ( w_15041 , w_15040 , \4747_b1 );
or ( \4749_b1 , \4745_b1 , w_15043 );
not ( w_15043 , w_15044 );
and ( \4749_b0 , \4745_b0 , w_15045 );
and ( w_15044 ,  , w_15045 );
buf ( w_15043 , \4135_b1 );
not ( w_15043 , w_15046 );
not (  , w_15047 );
and ( w_15046 , w_15047 , \4135_b0 );
or ( \4750_b1 , \4748_b1 , w_15049 );
not ( w_15049 , w_15050 );
and ( \4750_b0 , \4748_b0 , w_15051 );
and ( w_15050 ,  , w_15051 );
buf ( w_15049 , \4749_b1 );
not ( w_15049 , w_15052 );
not (  , w_15053 );
and ( w_15052 , w_15053 , \4749_b0 );
buf ( \4751_b1 , \4750_b1 );
not ( \4751_b1 , w_15054 );
not ( \4751_b0 , w_15055 );
and ( w_15054 , w_15055 , \4750_b0 );
buf ( \4752_b1 , \4611_b1 );
not ( \4752_b1 , w_15056 );
not ( \4752_b0 , w_15057 );
and ( w_15056 , w_15057 , \4611_b0 );
or ( \4753_b1 , \4751_b1 , w_15058 );
or ( \4753_b0 , \4751_b0 , \4752_b0 );
not ( \4752_b0 , w_15059 );
and ( w_15059 , w_15058 , \4752_b1 );
buf ( \4754_b1 , \4602_b1 );
not ( \4754_b1 , w_15060 );
not ( \4754_b0 , w_15061 );
and ( w_15060 , w_15061 , \4602_b0 );
or ( \4755_b1 , \4754_b1 , w_15063 );
not ( w_15063 , w_15064 );
and ( \4755_b0 , \4754_b0 , w_15065 );
and ( w_15064 ,  , w_15065 );
buf ( w_15063 , \4616_b1 );
not ( w_15063 , w_15066 );
not (  , w_15067 );
and ( w_15066 , w_15067 , \4616_b0 );
or ( \4756_b1 , \4753_b1 , w_15069 );
not ( w_15069 , w_15070 );
and ( \4756_b0 , \4753_b0 , w_15071 );
and ( w_15070 ,  , w_15071 );
buf ( w_15069 , \4755_b1 );
not ( w_15069 , w_15072 );
not (  , w_15073 );
and ( w_15072 , w_15073 , \4755_b0 );
buf ( \4757_b1 , \4756_b1 );
not ( \4757_b1 , w_15074 );
not ( \4757_b0 , w_15075 );
and ( w_15074 , w_15075 , \4756_b0 );
or ( \4758_b1 , \4743_b1 , w_15077 );
not ( w_15077 , w_15078 );
and ( \4758_b0 , \4743_b0 , w_15079 );
and ( w_15078 ,  , w_15079 );
buf ( w_15077 , \4757_b1 );
not ( w_15077 , w_15080 );
not (  , w_15081 );
and ( w_15080 , w_15081 , \4757_b0 );
or ( \4759_b1 , \4741_b1 , \4758_b1 );
not ( \4758_b1 , w_15082 );
and ( \4759_b0 , \4741_b0 , w_15083 );
and ( w_15082 , w_15083 , \4758_b0 );
or ( \4760_b1 , \4742_b1 , \4756_b1 );
not ( \4756_b1 , w_15084 );
and ( \4760_b0 , \4742_b0 , w_15085 );
and ( w_15084 , w_15085 , \4756_b0 );
or ( \4761_b1 , \4759_b1 , w_15087 );
not ( w_15087 , w_15088 );
and ( \4761_b0 , \4759_b0 , w_15089 );
and ( w_15088 ,  , w_15089 );
buf ( w_15087 , \4760_b1 );
not ( w_15087 , w_15090 );
not (  , w_15091 );
and ( w_15090 , w_15091 , \4760_b0 );
or ( \4762_b1 , \4703_b1 , w_15093 );
not ( w_15093 , w_15094 );
and ( \4762_b0 , \4703_b0 , w_15095 );
and ( w_15094 ,  , w_15095 );
buf ( w_15093 , \4761_b1 );
not ( w_15093 , w_15096 );
not (  , w_15097 );
and ( w_15096 , w_15097 , \4761_b0 );
buf ( \4763_b1 , \4762_b1 );
not ( \4763_b1 , w_15098 );
not ( \4763_b0 , w_15099 );
and ( w_15098 , w_15099 , \4762_b0 );
or ( \4764_b1 , \4680_b1 , \4656_b1 );
not ( \4656_b1 , w_15100 );
and ( \4764_b0 , \4680_b0 , w_15101 );
and ( w_15100 , w_15101 , \4656_b0 );
buf ( \4765_b1 , \4680_b1 );
not ( \4765_b1 , w_15102 );
not ( \4765_b0 , w_15103 );
and ( w_15102 , w_15103 , \4680_b0 );
or ( \4766_b1 , \4765_b1 , \4682_b1 );
not ( \4682_b1 , w_15104 );
and ( \4766_b0 , \4765_b0 , w_15105 );
and ( w_15104 , w_15105 , \4682_b0 );
or ( \4767_b1 , \4764_b1 , w_15107 );
not ( w_15107 , w_15108 );
and ( \4767_b0 , \4764_b0 , w_15109 );
and ( w_15108 ,  , w_15109 );
buf ( w_15107 , \4766_b1 );
not ( w_15107 , w_15110 );
not (  , w_15111 );
and ( w_15110 , w_15111 , \4766_b0 );
buf ( \4768_b1 , \4668_b1 );
not ( \4768_b1 , w_15112 );
not ( \4768_b0 , w_15113 );
and ( w_15112 , w_15113 , \4668_b0 );
or ( \4769_b1 , \4767_b1 , \4768_b1 );
not ( \4768_b1 , w_15114 );
and ( \4769_b0 , \4767_b0 , w_15115 );
and ( w_15114 , w_15115 , \4768_b0 );
buf ( \4770_b1 , \4767_b1 );
not ( \4770_b1 , w_15116 );
not ( \4770_b0 , w_15117 );
and ( w_15116 , w_15117 , \4767_b0 );
or ( \4771_b1 , \4770_b1 , \4668_b1 );
not ( \4668_b1 , w_15118 );
and ( \4771_b0 , \4770_b0 , w_15119 );
and ( w_15118 , w_15119 , \4668_b0 );
or ( \4772_b1 , \4769_b1 , w_15121 );
not ( w_15121 , w_15122 );
and ( \4772_b0 , \4769_b0 , w_15123 );
and ( w_15122 ,  , w_15123 );
buf ( w_15121 , \4771_b1 );
not ( w_15121 , w_15124 );
not (  , w_15125 );
and ( w_15124 , w_15125 , \4771_b0 );
buf ( \4773_b1 , \4772_b1 );
not ( \4773_b1 , w_15126 );
not ( \4773_b0 , w_15127 );
and ( w_15126 , w_15127 , \4772_b0 );
buf ( \4774_b1 , \4773_b1 );
not ( \4774_b1 , w_15128 );
not ( \4774_b0 , w_15129 );
and ( w_15128 , w_15129 , \4773_b0 );
or ( \4775_b1 , \4100_b1 , \4026_b1 );
not ( \4026_b1 , w_15130 );
and ( \4775_b0 , \4100_b0 , w_15131 );
and ( w_15130 , w_15131 , \4026_b0 );
buf ( \4776_b1 , \4775_b1 );
not ( \4776_b1 , w_15132 );
not ( \4776_b0 , w_15133 );
and ( w_15132 , w_15133 , \4775_b0 );
buf ( \4777_b1 , \4021_b1 );
not ( \4777_b1 , w_15134 );
not ( \4777_b0 , w_15135 );
and ( w_15134 , w_15135 , \4021_b0 );
buf ( \4778_b1 , \4101_b1 );
not ( \4778_b1 , w_15136 );
not ( \4778_b0 , w_15137 );
and ( w_15136 , w_15137 , \4101_b0 );
or ( \4779_b1 , \4777_b1 , w_15138 );
or ( \4779_b0 , \4777_b0 , \4778_b0 );
not ( \4778_b0 , w_15139 );
and ( w_15139 , w_15138 , \4778_b1 );
buf ( \4780_b1 , \4021_b1 );
not ( \4780_b1 , w_15140 );
not ( \4780_b0 , w_15141 );
and ( w_15140 , w_15141 , \4021_b0 );
or ( \4781_b1 , \4100_b1 , w_15143 );
not ( w_15143 , w_15144 );
and ( \4781_b0 , \4100_b0 , w_15145 );
and ( w_15144 ,  , w_15145 );
buf ( w_15143 , \4780_b1 );
not ( w_15143 , w_15146 );
not (  , w_15147 );
and ( w_15146 , w_15147 , \4780_b0 );
or ( \4782_b1 , \4779_b1 , w_15149 );
not ( w_15149 , w_15150 );
and ( \4782_b0 , \4779_b0 , w_15151 );
and ( w_15150 ,  , w_15151 );
buf ( w_15149 , \4781_b1 );
not ( w_15149 , w_15152 );
not (  , w_15153 );
and ( w_15152 , w_15153 , \4781_b0 );
buf ( \4783_b1 , \4782_b1 );
not ( \4783_b1 , w_15154 );
not ( \4783_b0 , w_15155 );
and ( w_15154 , w_15155 , \4782_b0 );
buf ( \4784_b1 , \4395_b1 );
not ( \4784_b1 , w_15156 );
not ( \4784_b0 , w_15157 );
and ( w_15156 , w_15157 , \4395_b0 );
or ( \4785_b1 , \4783_b1 , w_15158 );
or ( \4785_b0 , \4783_b0 , \4784_b0 );
not ( \4784_b0 , w_15159 );
and ( w_15159 , w_15158 , \4784_b1 );
or ( \4786_b1 , \4664_b1 , w_15161 );
not ( w_15161 , w_15162 );
and ( \4786_b0 , \4664_b0 , w_15163 );
and ( w_15162 ,  , w_15163 );
buf ( w_15161 , \4200_b1 );
not ( w_15161 , w_15164 );
not (  , w_15165 );
and ( w_15164 , w_15165 , \4200_b0 );
or ( \4787_b1 , \4785_b1 , w_15167 );
not ( w_15167 , w_15168 );
and ( \4787_b0 , \4785_b0 , w_15169 );
and ( w_15168 ,  , w_15169 );
buf ( w_15167 , \4786_b1 );
not ( w_15167 , w_15170 );
not (  , w_15171 );
and ( w_15170 , w_15171 , \4786_b0 );
buf ( \4788_b1 , \4787_b1 );
not ( \4788_b1 , w_15172 );
not ( \4788_b0 , w_15173 );
and ( w_15172 , w_15173 , \4787_b0 );
or ( \4789_b1 , \4776_b1 , w_15174 );
or ( \4789_b0 , \4776_b0 , \4788_b0 );
not ( \4788_b0 , w_15175 );
and ( w_15175 , w_15174 , \4788_b1 );
or ( \4790_b1 , \4787_b1 , w_15176 );
or ( \4790_b0 , \4787_b0 , \4775_b0 );
not ( \4775_b0 , w_15177 );
and ( w_15177 , w_15176 , \4775_b1 );
buf ( \4791_b1 , \4096_b1 );
not ( \4791_b1 , w_15178 );
not ( \4791_b0 , w_15179 );
and ( w_15178 , w_15179 , \4096_b0 );
buf ( \4792_b1 , \4284_b1 );
not ( \4792_b1 , w_15180 );
not ( \4792_b0 , w_15181 );
and ( w_15180 , w_15181 , \4284_b0 );
or ( \4793_b1 , \4791_b1 , w_15182 );
or ( \4793_b0 , \4791_b0 , \4792_b0 );
not ( \4792_b0 , w_15183 );
and ( w_15183 , w_15182 , \4792_b1 );
or ( \4794_b1 , \4283_b1 , w_15185 );
not ( w_15185 , w_15186 );
and ( \4794_b0 , \4283_b0 , w_15187 );
and ( w_15186 ,  , w_15187 );
buf ( w_15185 , \4372_b1 );
not ( w_15185 , w_15188 );
not (  , w_15189 );
and ( w_15188 , w_15189 , \4372_b0 );
or ( \4795_b1 , \4793_b1 , w_15191 );
not ( w_15191 , w_15192 );
and ( \4795_b0 , \4793_b0 , w_15193 );
and ( w_15192 ,  , w_15193 );
buf ( w_15191 , \4794_b1 );
not ( w_15191 , w_15194 );
not (  , w_15195 );
and ( w_15194 , w_15195 , \4794_b0 );
buf ( \4796_b1 , \4795_b1 );
not ( \4796_b1 , w_15196 );
not ( \4796_b0 , w_15197 );
and ( w_15196 , w_15197 , \4795_b0 );
buf ( \4797_b1 , \4278_b1 );
not ( \4797_b1 , w_15198 );
not ( \4797_b0 , w_15199 );
and ( w_15198 , w_15199 , \4278_b0 );
buf ( \4798_b1 , \4797_b1 );
not ( \4798_b1 , w_15200 );
not ( \4798_b0 , w_15201 );
and ( w_15200 , w_15201 , \4797_b0 );
or ( \4799_b1 , \4796_b1 , w_15202 );
or ( \4799_b0 , \4796_b0 , \4798_b0 );
not ( \4798_b0 , w_15203 );
and ( w_15203 , w_15202 , \4798_b1 );
buf ( \4800_b1 , \4265_b1 );
not ( \4800_b1 , w_15204 );
not ( \4800_b0 , w_15205 );
and ( w_15204 , w_15205 , \4265_b0 );
or ( \4801_b1 , \4675_b1 , w_15207 );
not ( w_15207 , w_15208 );
and ( \4801_b0 , \4675_b0 , w_15209 );
and ( w_15208 ,  , w_15209 );
buf ( w_15207 , \4800_b1 );
not ( w_15207 , w_15210 );
not (  , w_15211 );
and ( w_15210 , w_15211 , \4800_b0 );
or ( \4802_b1 , \4799_b1 , w_15213 );
not ( w_15213 , w_15214 );
and ( \4802_b0 , \4799_b0 , w_15215 );
and ( w_15214 ,  , w_15215 );
buf ( w_15213 , \4801_b1 );
not ( w_15213 , w_15216 );
not (  , w_15217 );
and ( w_15216 , w_15217 , \4801_b0 );
or ( \4803_b1 , \4790_b1 , w_15219 );
not ( w_15219 , w_15220 );
and ( \4803_b0 , \4790_b0 , w_15221 );
and ( w_15220 ,  , w_15221 );
buf ( w_15219 , \4802_b1 );
not ( w_15219 , w_15222 );
not (  , w_15223 );
and ( w_15222 , w_15223 , \4802_b0 );
or ( \4804_b1 , \4789_b1 , w_15225 );
not ( w_15225 , w_15226 );
and ( \4804_b0 , \4789_b0 , w_15227 );
and ( w_15226 ,  , w_15227 );
buf ( w_15225 , \4803_b1 );
not ( w_15225 , w_15228 );
not (  , w_15229 );
and ( w_15228 , w_15229 , \4803_b0 );
buf ( \4805_b1 , \4804_b1 );
not ( \4805_b1 , w_15230 );
not ( \4805_b0 , w_15231 );
and ( w_15230 , w_15231 , \4804_b0 );
or ( \4806_b1 , \4774_b1 , w_15232 );
or ( \4806_b0 , \4774_b0 , \4805_b0 );
not ( \4805_b0 , w_15233 );
and ( w_15233 , w_15232 , \4805_b1 );
buf ( \4807_b1 , \4804_b1 );
not ( \4807_b1 , w_15234 );
not ( \4807_b0 , w_15235 );
and ( w_15234 , w_15235 , \4804_b0 );
buf ( \4808_b1 , \4807_b1 );
not ( \4808_b1 , w_15236 );
not ( \4808_b0 , w_15237 );
and ( w_15236 , w_15237 , \4807_b0 );
buf ( \4809_b1 , \4772_b1 );
not ( \4809_b1 , w_15238 );
not ( \4809_b0 , w_15239 );
and ( w_15238 , w_15239 , \4772_b0 );
or ( \4810_b1 , \4808_b1 , w_15240 );
or ( \4810_b0 , \4808_b0 , \4809_b0 );
not ( \4809_b0 , w_15241 );
and ( w_15241 , w_15240 , \4809_b1 );
or ( \4811_b1 , \4617_b1 , \4640_b1 );
xor ( \4811_b0 , \4617_b0 , w_15242 );
not ( w_15242 , w_15243 );
and ( w_15243 , \4640_b1 , \4640_b0 );
or ( \4812_b1 , \4811_b1 , w_15244 );
xor ( \4812_b0 , \4811_b0 , w_15246 );
not ( w_15246 , w_15247 );
and ( w_15247 , w_15244 , w_15245 );
buf ( w_15244 , \4628_b1 );
not ( w_15244 , w_15248 );
not ( w_15245 , w_15249 );
and ( w_15248 , w_15249 , \4628_b0 );
or ( \4813_b1 , \4810_b1 , w_15251 );
not ( w_15251 , w_15252 );
and ( \4813_b0 , \4810_b0 , w_15253 );
and ( w_15252 ,  , w_15253 );
buf ( w_15251 , \4812_b1 );
not ( w_15251 , w_15254 );
not (  , w_15255 );
and ( w_15254 , w_15255 , \4812_b0 );
or ( \4814_b1 , \4806_b1 , w_15257 );
not ( w_15257 , w_15258 );
and ( \4814_b0 , \4806_b0 , w_15259 );
and ( w_15258 ,  , w_15259 );
buf ( w_15257 , \4813_b1 );
not ( w_15257 , w_15260 );
not (  , w_15261 );
and ( w_15260 , w_15261 , \4813_b0 );
buf ( \4815_b1 , \4814_b1 );
not ( \4815_b1 , w_15262 );
not ( \4815_b0 , w_15263 );
and ( w_15262 , w_15263 , \4814_b0 );
or ( \4816_b1 , \4763_b1 , w_15264 );
or ( \4816_b0 , \4763_b0 , \4815_b0 );
not ( \4815_b0 , w_15265 );
and ( w_15265 , w_15264 , \4815_b1 );
buf ( \4817_b1 , \4761_b1 );
not ( \4817_b1 , w_15266 );
not ( \4817_b0 , w_15267 );
and ( w_15266 , w_15267 , \4761_b0 );
or ( \4818_b1 , \4817_b1 , w_15269 );
not ( w_15269 , w_15270 );
and ( \4818_b0 , \4817_b0 , w_15271 );
and ( w_15270 ,  , w_15271 );
buf ( w_15269 , \4702_b1 );
not ( w_15269 , w_15272 );
not (  , w_15273 );
and ( w_15272 , w_15273 , \4702_b0 );
or ( \4819_b1 , \4816_b1 , w_15275 );
not ( w_15275 , w_15276 );
and ( \4819_b0 , \4816_b0 , w_15277 );
and ( w_15276 ,  , w_15277 );
buf ( w_15275 , \4818_b1 );
not ( w_15275 , w_15278 );
not (  , w_15279 );
and ( w_15278 , w_15279 , \4818_b0 );
or ( \4820_b1 , \4700_b1 , \4819_b1 );
not ( \4819_b1 , w_15280 );
and ( \4820_b0 , \4700_b0 , w_15281 );
and ( w_15280 , w_15281 , \4819_b0 );
or ( \4821_b1 , \4688_b1 , \4699_b1 );
not ( \4699_b1 , w_15282 );
and ( \4821_b0 , \4688_b0 , w_15283 );
and ( w_15282 , w_15283 , \4699_b0 );
or ( \4822_b1 , \4820_b1 , w_15284 );
or ( \4822_b0 , \4820_b0 , \4821_b0 );
not ( \4821_b0 , w_15285 );
and ( w_15285 , w_15284 , \4821_b1 );
or ( \4823_b1 , \4550_b1 , \4552_b1 );
xor ( \4823_b0 , \4550_b0 , w_15286 );
not ( w_15286 , w_15287 );
and ( w_15287 , \4552_b1 , \4552_b0 );
or ( \4824_b1 , \4823_b1 , \4583_b1 );
xor ( \4824_b0 , \4823_b0 , w_15288 );
not ( w_15288 , w_15289 );
and ( w_15289 , \4583_b1 , \4583_b0 );
or ( \4825_b1 , \4822_b1 , w_15291 );
not ( w_15291 , w_15292 );
and ( \4825_b0 , \4822_b0 , w_15293 );
and ( w_15292 ,  , w_15293 );
buf ( w_15291 , \4824_b1 );
not ( w_15291 , w_15294 );
not (  , w_15295 );
and ( w_15294 , w_15295 , \4824_b0 );
buf ( \4826_b1 , \4825_b1 );
not ( \4826_b1 , w_15296 );
not ( \4826_b0 , w_15297 );
and ( w_15296 , w_15297 , \4825_b0 );
or ( \4827_b1 , \4688_b1 , \4699_b1 );
xor ( \4827_b0 , \4688_b0 , w_15298 );
not ( w_15298 , w_15299 );
and ( w_15299 , \4699_b1 , \4699_b0 );
or ( \4828_b1 , \4827_b1 , \4819_b1 );
xor ( \4828_b0 , \4827_b0 , w_15300 );
not ( w_15300 , w_15301 );
and ( w_15301 , \4819_b1 , \4819_b0 );
buf ( \4829_b1 , \4761_b1 );
not ( \4829_b1 , w_15302 );
not ( \4829_b0 , w_15303 );
and ( w_15302 , w_15303 , \4761_b0 );
buf ( \4830_b1 , \4702_b1 );
not ( \4830_b1 , w_15304 );
not ( \4830_b0 , w_15305 );
and ( w_15304 , w_15305 , \4702_b0 );
or ( \4831_b1 , \4829_b1 , w_15306 );
or ( \4831_b0 , \4829_b0 , \4830_b0 );
not ( \4830_b0 , w_15307 );
and ( w_15307 , w_15306 , \4830_b1 );
or ( \4832_b1 , \4761_b1 , w_15308 );
or ( \4832_b0 , \4761_b0 , \4702_b0 );
not ( \4702_b0 , w_15309 );
and ( w_15309 , w_15308 , \4702_b1 );
or ( \4833_b1 , \4831_b1 , w_15311 );
not ( w_15311 , w_15312 );
and ( \4833_b0 , \4831_b0 , w_15313 );
and ( w_15312 ,  , w_15313 );
buf ( w_15311 , \4832_b1 );
not ( w_15311 , w_15314 );
not (  , w_15315 );
and ( w_15314 , w_15315 , \4832_b0 );
or ( \4834_b1 , \4814_b1 , \4833_b1 );
xor ( \4834_b0 , \4814_b0 , w_15316 );
not ( w_15316 , w_15317 );
and ( w_15317 , \4833_b1 , \4833_b0 );
buf ( \4835_b1 , \4834_b1 );
not ( \4835_b1 , w_15318 );
not ( \4835_b0 , w_15319 );
and ( w_15318 , w_15319 , \4834_b0 );
or ( \4836_b1 , \4596_b1 , \4643_b1 );
xor ( \4836_b0 , \4596_b0 , w_15320 );
not ( w_15320 , w_15321 );
and ( w_15321 , \4643_b1 , \4643_b0 );
or ( \4837_b1 , \4836_b1 , \4685_b1 );
xor ( \4837_b0 , \4836_b0 , w_15322 );
not ( w_15322 , w_15323 );
and ( w_15323 , \4685_b1 , \4685_b0 );
buf ( \4838_b1 , \4837_b1 );
buf ( \4838_b0 , \4837_b0 );
buf ( \4839_b1 , \4838_b1 );
not ( \4839_b1 , w_15324 );
not ( \4839_b0 , w_15325 );
and ( w_15324 , w_15325 , \4838_b0 );
or ( \4840_b1 , \4835_b1 , w_15326 );
or ( \4840_b0 , \4835_b0 , \4839_b0 );
not ( \4839_b0 , w_15327 );
and ( w_15327 , w_15326 , \4839_b1 );
or ( \4841_b1 , \4838_b1 , w_15328 );
or ( \4841_b0 , \4838_b0 , \4834_b0 );
not ( \4834_b0 , w_15329 );
and ( w_15329 , w_15328 , \4834_b1 );
or ( \4842_b1 , \4742_b1 , \4756_b1 );
xor ( \4842_b0 , \4742_b0 , w_15330 );
not ( w_15330 , w_15331 );
and ( w_15331 , \4756_b1 , \4756_b0 );
or ( \4843_b1 , \4741_b1 , \4842_b1 );
not ( \4842_b1 , w_15332 );
and ( \4843_b0 , \4741_b0 , w_15333 );
and ( w_15332 , w_15333 , \4842_b0 );
buf ( \4844_b1 , \4741_b1 );
not ( \4844_b1 , w_15334 );
not ( \4844_b0 , w_15335 );
and ( w_15334 , w_15335 , \4741_b0 );
buf ( \4845_b1 , \4842_b1 );
not ( \4845_b1 , w_15336 );
not ( \4845_b0 , w_15337 );
and ( w_15336 , w_15337 , \4842_b0 );
or ( \4846_b1 , \4844_b1 , \4845_b1 );
not ( \4845_b1 , w_15338 );
and ( \4846_b0 , \4844_b0 , w_15339 );
and ( w_15338 , w_15339 , \4845_b0 );
or ( \4847_b1 , \4843_b1 , w_15341 );
not ( w_15341 , w_15342 );
and ( \4847_b0 , \4843_b0 , w_15343 );
and ( w_15342 ,  , w_15343 );
buf ( w_15341 , \4846_b1 );
not ( w_15341 , w_15344 );
not (  , w_15345 );
and ( w_15344 , w_15345 , \4846_b0 );
buf ( \4848_b1 , \4847_b1 );
buf ( \4848_b0 , \4847_b0 );
buf ( \4849_b1 , \4848_b1 );
not ( \4849_b1 , w_15346 );
not ( \4849_b0 , w_15347 );
and ( w_15346 , w_15347 , \4848_b0 );
buf ( \4850_b1 , \4757_b1 );
not ( \4850_b1 , w_15348 );
not ( \4850_b0 , w_15349 );
and ( w_15348 , w_15349 , \4757_b0 );
buf ( \4851_b1 , \3016_b1 );
buf ( \4851_b0 , \3016_b0 );
buf ( \4852_b1 , \4851_b1 );
not ( \4852_b1 , w_15350 );
not ( \4852_b0 , w_15351 );
and ( w_15350 , w_15351 , \4851_b0 );
buf ( \4853_b1 , \2945_b1 );
not ( \4853_b1 , w_15352 );
not ( \4853_b0 , w_15353 );
and ( w_15352 , w_15353 , \2945_b0 );
buf ( \4854_b1 , \4853_b1 );
not ( \4854_b1 , w_15354 );
not ( \4854_b0 , w_15355 );
and ( w_15354 , w_15355 , \4853_b0 );
or ( \4855_b1 , \4852_b1 , w_15356 );
or ( \4855_b0 , \4852_b0 , \4854_b0 );
not ( \4854_b0 , w_15357 );
and ( w_15357 , w_15356 , \4854_b1 );
buf ( \4856_b1 , \4851_b1 );
not ( \4856_b1 , w_15358 );
not ( \4856_b0 , w_15359 );
and ( w_15358 , w_15359 , \4851_b0 );
or ( \4857_b1 , \4856_b1 , w_15361 );
not ( w_15361 , w_15362 );
and ( \4857_b0 , \4856_b0 , w_15363 );
and ( w_15362 ,  , w_15363 );
buf ( w_15361 , \2945_b1 );
not ( w_15361 , w_15364 );
not (  , w_15365 );
and ( w_15364 , w_15365 , \2945_b0 );
or ( \4858_b1 , \4855_b1 , w_15367 );
not ( w_15367 , w_15368 );
and ( \4858_b0 , \4855_b0 , w_15369 );
and ( w_15368 ,  , w_15369 );
buf ( w_15367 , \4857_b1 );
not ( w_15367 , w_15370 );
not (  , w_15371 );
and ( w_15370 , w_15371 , \4857_b0 );
buf ( \4859_b1 , \4858_b1 );
buf ( \4859_b0 , \4858_b0 );
buf ( \4860_b1 , \4859_b1 );
not ( \4860_b1 , w_15372 );
not ( \4860_b0 , w_15373 );
and ( w_15372 , w_15373 , \4859_b0 );
or ( \4861_b1 , \3016_b1 , w_15374 );
xor ( \4861_b0 , \3016_b0 , w_15376 );
not ( w_15376 , w_15377 );
and ( w_15377 , w_15374 , w_15375 );
buf ( w_15374 , \3070_b1 );
not ( w_15374 , w_15378 );
not ( w_15375 , w_15379 );
and ( w_15378 , w_15379 , \3070_b0 );
buf ( \4862_b1 , \4861_b1 );
buf ( \4862_b0 , \4861_b0 );
buf ( \4863_b1 , \4862_b1 );
not ( \4863_b1 , w_15380 );
not ( \4863_b0 , w_15381 );
and ( w_15380 , w_15381 , \4862_b0 );
buf ( \4864_b1 , \4863_b1 );
not ( \4864_b1 , w_15382 );
not ( \4864_b0 , w_15383 );
and ( w_15382 , w_15383 , \4863_b0 );
or ( \4865_b1 , \4860_b1 , \4864_b1 );
not ( \4864_b1 , w_15384 );
and ( \4865_b0 , \4860_b0 , w_15385 );
and ( w_15384 , w_15385 , \4864_b0 );
buf ( \4866_b1 , \4853_b1 );
buf ( \4866_b0 , \4853_b0 );
buf ( \4867_b1 , \4866_b1 );
not ( \4867_b1 , w_15386 );
not ( \4867_b0 , w_15387 );
and ( w_15386 , w_15387 , \4866_b0 );
buf ( \4868_b1 , \4867_b1 );
buf ( \4868_b0 , \4867_b0 );
buf ( \4869_b1 , \4868_b1 );
not ( \4869_b1 , w_15388 );
not ( \4869_b0 , w_15389 );
and ( w_15388 , w_15389 , \4868_b0 );
or ( \4870_b1 , \4865_b1 , w_15391 );
not ( w_15391 , w_15392 );
and ( \4870_b0 , \4865_b0 , w_15393 );
and ( w_15392 ,  , w_15393 );
buf ( w_15391 , \4869_b1 );
not ( w_15391 , w_15394 );
not (  , w_15395 );
and ( w_15394 , w_15395 , \4869_b0 );
buf ( \4871_b1 , \4870_b1 );
not ( \4871_b1 , w_15396 );
not ( \4871_b0 , w_15397 );
and ( w_15396 , w_15397 , \4870_b0 );
buf ( \4872_b1 , \4871_b1 );
not ( \4872_b1 , w_15398 );
not ( \4872_b0 , w_15399 );
and ( w_15398 , w_15399 , \4871_b0 );
buf ( \4873_b1 , \4610_b1 );
not ( \4873_b1 , w_15400 );
not ( \4873_b0 , w_15401 );
and ( w_15400 , w_15401 , \4610_b0 );
buf ( \4874_b1 , \3997_b1 );
not ( \4874_b1 , w_15402 );
not ( \4874_b0 , w_15403 );
and ( w_15402 , w_15403 , \3997_b0 );
buf ( \4875_b1 , \4746_b1 );
not ( \4875_b1 , w_15404 );
not ( \4875_b0 , w_15405 );
and ( w_15404 , w_15405 , \4746_b0 );
or ( \4876_b1 , \4874_b1 , w_15406 );
or ( \4876_b0 , \4874_b0 , \4875_b0 );
not ( \4875_b0 , w_15407 );
and ( w_15407 , w_15406 , \4875_b1 );
or ( \4877_b1 , \4745_b1 , w_15409 );
not ( w_15409 , w_15410 );
and ( \4877_b0 , \4745_b0 , w_15411 );
and ( w_15410 ,  , w_15411 );
buf ( w_15409 , \4111_b1 );
not ( w_15409 , w_15412 );
not (  , w_15413 );
and ( w_15412 , w_15413 , \4111_b0 );
or ( \4878_b1 , \4876_b1 , w_15415 );
not ( w_15415 , w_15416 );
and ( \4878_b0 , \4876_b0 , w_15417 );
and ( w_15416 ,  , w_15417 );
buf ( w_15415 , \4877_b1 );
not ( w_15415 , w_15418 );
not (  , w_15419 );
and ( w_15418 , w_15419 , \4877_b0 );
buf ( \4879_b1 , \4878_b1 );
not ( \4879_b1 , w_15420 );
not ( \4879_b0 , w_15421 );
and ( w_15420 , w_15421 , \4878_b0 );
or ( \4880_b1 , \4873_b1 , w_15422 );
or ( \4880_b0 , \4873_b0 , \4879_b0 );
not ( \4879_b0 , w_15423 );
and ( w_15423 , w_15422 , \4879_b1 );
buf ( \4881_b1 , \4602_b1 );
not ( \4881_b1 , w_15424 );
not ( \4881_b0 , w_15425 );
and ( w_15424 , w_15425 , \4602_b0 );
or ( \4882_b1 , \4881_b1 , w_15427 );
not ( w_15427 , w_15428 );
and ( \4882_b0 , \4881_b0 , w_15429 );
and ( w_15428 ,  , w_15429 );
buf ( w_15427 , \4750_b1 );
not ( w_15427 , w_15430 );
not (  , w_15431 );
and ( w_15430 , w_15431 , \4750_b0 );
or ( \4883_b1 , \4880_b1 , w_15433 );
not ( w_15433 , w_15434 );
and ( \4883_b0 , \4880_b0 , w_15435 );
and ( w_15434 ,  , w_15435 );
buf ( w_15433 , \4882_b1 );
not ( w_15433 , w_15436 );
not (  , w_15437 );
and ( w_15436 , w_15437 , \4882_b0 );
buf ( \4884_b1 , \4883_b1 );
not ( \4884_b1 , w_15438 );
not ( \4884_b0 , w_15439 );
and ( w_15438 , w_15439 , \4883_b0 );
or ( \4885_b1 , \4872_b1 , w_15440 );
or ( \4885_b0 , \4872_b0 , \4884_b0 );
not ( \4884_b0 , w_15441 );
and ( w_15441 , w_15440 , \4884_b1 );
or ( \4886_b1 , \4871_b1 , w_15442 );
or ( \4886_b0 , \4871_b0 , \4883_b0 );
not ( \4883_b0 , w_15443 );
and ( w_15443 , w_15442 , \4883_b1 );
buf ( \4887_b1 , \4097_b1 );
not ( \4887_b1 , w_15444 );
not ( \4887_b0 , w_15445 );
and ( w_15444 , w_15445 , \4097_b0 );
buf ( \4888_b1 , \4493_b1 );
not ( \4888_b1 , w_15446 );
not ( \4888_b0 , w_15447 );
and ( w_15446 , w_15447 , \4493_b0 );
or ( \4889_b1 , \4887_b1 , w_15448 );
or ( \4889_b0 , \4887_b0 , \4888_b0 );
not ( \4888_b0 , w_15449 );
and ( w_15449 , w_15448 , \4888_b1 );
or ( \4890_b1 , \4285_b1 , w_15451 );
not ( w_15451 , w_15452 );
and ( \4890_b0 , \4285_b0 , w_15453 );
and ( w_15452 ,  , w_15453 );
buf ( w_15451 , \4254_b1 );
not ( w_15451 , w_15454 );
not (  , w_15455 );
and ( w_15454 , w_15455 , \4254_b0 );
or ( \4891_b1 , \4889_b1 , w_15457 );
not ( w_15457 , w_15458 );
and ( \4891_b0 , \4889_b0 , w_15459 );
and ( w_15458 ,  , w_15459 );
buf ( w_15457 , \4890_b1 );
not ( w_15457 , w_15460 );
not (  , w_15461 );
and ( w_15460 , w_15461 , \4890_b0 );
buf ( \4892_b1 , \4891_b1 );
not ( \4892_b1 , w_15462 );
not ( \4892_b0 , w_15463 );
and ( w_15462 , w_15463 , \4891_b0 );
buf ( \4893_b1 , \4430_b1 );
not ( \4893_b1 , w_15464 );
not ( \4893_b0 , w_15465 );
and ( w_15464 , w_15465 , \4430_b0 );
or ( \4894_b1 , \4892_b1 , w_15466 );
or ( \4894_b0 , \4892_b0 , \4893_b0 );
not ( \4893_b0 , w_15467 );
and ( w_15467 , w_15466 , \4893_b1 );
or ( \4895_b1 , \4341_b1 , w_15469 );
not ( w_15469 , w_15470 );
and ( \4895_b0 , \4341_b0 , w_15471 );
and ( w_15470 ,  , w_15471 );
buf ( w_15469 , \4795_b1 );
not ( w_15469 , w_15472 );
not (  , w_15473 );
and ( w_15472 , w_15473 , \4795_b0 );
or ( \4896_b1 , \4894_b1 , w_15475 );
not ( w_15475 , w_15476 );
and ( \4896_b0 , \4894_b0 , w_15477 );
and ( w_15476 ,  , w_15477 );
buf ( w_15475 , \4895_b1 );
not ( w_15475 , w_15478 );
not (  , w_15479 );
and ( w_15478 , w_15479 , \4895_b0 );
or ( \4897_b1 , \4886_b1 , w_15481 );
not ( w_15481 , w_15482 );
and ( \4897_b0 , \4886_b0 , w_15483 );
and ( w_15482 ,  , w_15483 );
buf ( w_15481 , \4896_b1 );
not ( w_15481 , w_15484 );
not (  , w_15485 );
and ( w_15484 , w_15485 , \4896_b0 );
or ( \4898_b1 , \4885_b1 , w_15487 );
not ( w_15487 , w_15488 );
and ( \4898_b0 , \4885_b0 , w_15489 );
and ( w_15488 ,  , w_15489 );
buf ( w_15487 , \4897_b1 );
not ( w_15487 , w_15490 );
not (  , w_15491 );
and ( w_15490 , w_15491 , \4897_b0 );
buf ( \4899_b1 , \4898_b1 );
not ( \4899_b1 , w_15492 );
not ( \4899_b0 , w_15493 );
and ( w_15492 , w_15493 , \4898_b0 );
or ( \4900_b1 , \4850_b1 , w_15494 );
or ( \4900_b0 , \4850_b0 , \4899_b0 );
not ( \4899_b0 , w_15495 );
and ( w_15495 , w_15494 , \4899_b1 );
or ( \4901_b1 , \4757_b1 , w_15496 );
or ( \4901_b0 , \4757_b0 , \4898_b0 );
not ( \4898_b0 , w_15497 );
and ( w_15497 , w_15496 , \4898_b1 );
or ( \4902_b1 , \4102_b1 , \4072_b1 );
not ( \4072_b1 , w_15498 );
and ( \4902_b0 , \4102_b0 , w_15499 );
and ( w_15498 , w_15499 , \4072_b0 );
buf ( \4903_b1 , \4902_b1 );
not ( \4903_b1 , w_15500 );
not ( \4903_b0 , w_15501 );
and ( w_15500 , w_15501 , \4902_b0 );
buf ( \4904_b1 , \4095_b1 );
not ( \4904_b1 , w_15502 );
not ( \4904_b0 , w_15503 );
and ( w_15502 , w_15503 , \4095_b0 );
buf ( \4905_b1 , \4163_b1 );
not ( \4905_b1 , w_15504 );
not ( \4905_b0 , w_15505 );
and ( w_15504 , w_15505 , \4163_b0 );
or ( \4906_b1 , \4904_b1 , w_15506 );
or ( \4906_b0 , \4904_b0 , \4905_b0 );
not ( \4905_b0 , w_15507 );
and ( w_15507 , w_15506 , \4905_b1 );
or ( \4907_b1 , \4164_b1 , w_15509 );
not ( w_15509 , w_15510 );
and ( \4907_b0 , \4164_b0 , w_15511 );
and ( w_15510 ,  , w_15511 );
buf ( w_15509 , \4391_b1 );
not ( w_15509 , w_15512 );
not (  , w_15513 );
and ( w_15512 , w_15513 , \4391_b0 );
or ( \4908_b1 , \4906_b1 , w_15515 );
not ( w_15515 , w_15516 );
and ( \4908_b0 , \4906_b0 , w_15517 );
and ( w_15516 ,  , w_15517 );
buf ( w_15515 , \4907_b1 );
not ( w_15515 , w_15518 );
not (  , w_15519 );
and ( w_15518 , w_15519 , \4907_b0 );
buf ( \4909_b1 , \4908_b1 );
not ( \4909_b1 , w_15520 );
not ( \4909_b0 , w_15521 );
and ( w_15520 , w_15521 , \4908_b0 );
buf ( \4910_b1 , \4159_b1 );
not ( \4910_b1 , w_15522 );
not ( \4910_b0 , w_15523 );
and ( w_15522 , w_15523 , \4159_b0 );
or ( \4911_b1 , \4909_b1 , w_15524 );
or ( \4911_b0 , \4909_b0 , \4910_b0 );
not ( \4910_b0 , w_15525 );
and ( w_15525 , w_15524 , \4910_b1 );
or ( \4912_b1 , \4150_b1 , w_15527 );
not ( w_15527 , w_15528 );
and ( \4912_b0 , \4150_b0 , w_15529 );
and ( w_15528 ,  , w_15529 );
buf ( w_15527 , \4720_b1 );
not ( w_15527 , w_15530 );
not (  , w_15531 );
and ( w_15530 , w_15531 , \4720_b0 );
or ( \4913_b1 , \4911_b1 , w_15533 );
not ( w_15533 , w_15534 );
and ( \4913_b0 , \4911_b0 , w_15535 );
and ( w_15534 ,  , w_15535 );
buf ( w_15533 , \4912_b1 );
not ( w_15533 , w_15536 );
not (  , w_15537 );
and ( w_15536 , w_15537 , \4912_b0 );
buf ( \4914_b1 , \4913_b1 );
not ( \4914_b1 , w_15538 );
not ( \4914_b0 , w_15539 );
and ( w_15538 , w_15539 , \4913_b0 );
or ( \4915_b1 , \4903_b1 , w_15540 );
or ( \4915_b0 , \4903_b0 , \4914_b0 );
not ( \4914_b0 , w_15541 );
and ( w_15541 , w_15540 , \4914_b1 );
or ( \4916_b1 , \4913_b1 , w_15542 );
or ( \4916_b0 , \4913_b0 , \4902_b0 );
not ( \4902_b0 , w_15543 );
and ( w_15543 , w_15542 , \4902_b1 );
buf ( \4917_b1 , \4732_b1 );
not ( \4917_b1 , w_15544 );
not ( \4917_b0 , w_15545 );
and ( w_15544 , w_15545 , \4732_b0 );
or ( \4918_b1 , \4094_b1 , \4917_b1 );
not ( \4917_b1 , w_15546 );
and ( \4918_b0 , \4094_b0 , w_15547 );
and ( w_15546 , w_15547 , \4917_b0 );
buf ( \4919_b1 , \4094_b1 );
not ( \4919_b1 , w_15548 );
not ( \4919_b0 , w_15549 );
and ( w_15548 , w_15549 , \4094_b0 );
or ( \4920_b1 , \4919_b1 , \4535_b1 );
not ( \4535_b1 , w_15550 );
and ( \4920_b0 , \4919_b0 , w_15551 );
and ( w_15550 , w_15551 , \4535_b0 );
or ( \4921_b1 , \4918_b1 , w_15553 );
not ( w_15553 , w_15554 );
and ( \4921_b0 , \4918_b0 , w_15555 );
and ( w_15554 ,  , w_15555 );
buf ( w_15553 , \4920_b1 );
not ( w_15553 , w_15556 );
not (  , w_15557 );
and ( w_15556 , w_15557 , \4920_b0 );
buf ( \4922_b1 , \4921_b1 );
not ( \4922_b1 , w_15558 );
not ( \4922_b0 , w_15559 );
and ( w_15558 , w_15559 , \4921_b0 );
buf ( \4923_b1 , \4632_b1 );
not ( \4923_b1 , w_15560 );
not ( \4923_b0 , w_15561 );
and ( w_15560 , w_15561 , \4632_b0 );
or ( \4924_b1 , \4922_b1 , w_15562 );
or ( \4924_b0 , \4922_b0 , \4923_b0 );
not ( \4923_b0 , w_15563 );
and ( w_15563 , w_15562 , \4923_b1 );
or ( \4925_b1 , \4453_b1 , w_15565 );
not ( w_15565 , w_15566 );
and ( \4925_b0 , \4453_b0 , w_15567 );
and ( w_15566 ,  , w_15567 );
buf ( w_15565 , \4734_b1 );
not ( w_15565 , w_15568 );
not (  , w_15569 );
and ( w_15568 , w_15569 , \4734_b0 );
or ( \4926_b1 , \4924_b1 , w_15571 );
not ( w_15571 , w_15572 );
and ( \4926_b0 , \4924_b0 , w_15573 );
and ( w_15572 ,  , w_15573 );
buf ( w_15571 , \4925_b1 );
not ( w_15571 , w_15574 );
not (  , w_15575 );
and ( w_15574 , w_15575 , \4925_b0 );
or ( \4927_b1 , \4916_b1 , w_15577 );
not ( w_15577 , w_15578 );
and ( \4927_b0 , \4916_b0 , w_15579 );
and ( w_15578 ,  , w_15579 );
buf ( w_15577 , \4926_b1 );
not ( w_15577 , w_15580 );
not (  , w_15581 );
and ( w_15580 , w_15581 , \4926_b0 );
or ( \4928_b1 , \4915_b1 , w_15583 );
not ( w_15583 , w_15584 );
and ( \4928_b0 , \4915_b0 , w_15585 );
and ( w_15584 ,  , w_15585 );
buf ( w_15583 , \4927_b1 );
not ( w_15583 , w_15586 );
not (  , w_15587 );
and ( w_15586 , w_15587 , \4927_b0 );
or ( \4929_b1 , \4901_b1 , w_15589 );
not ( w_15589 , w_15590 );
and ( \4929_b0 , \4901_b0 , w_15591 );
and ( w_15590 ,  , w_15591 );
buf ( w_15589 , \4928_b1 );
not ( w_15589 , w_15592 );
not (  , w_15593 );
and ( w_15592 , w_15593 , \4928_b0 );
or ( \4930_b1 , \4900_b1 , w_15595 );
not ( w_15595 , w_15596 );
and ( \4930_b0 , \4900_b0 , w_15597 );
and ( w_15596 ,  , w_15597 );
buf ( w_15595 , \4929_b1 );
not ( w_15595 , w_15598 );
not (  , w_15599 );
and ( w_15598 , w_15599 , \4929_b0 );
buf ( \4931_b1 , \4930_b1 );
not ( \4931_b1 , w_15600 );
not ( \4931_b0 , w_15601 );
and ( w_15600 , w_15601 , \4930_b0 );
or ( \4932_b1 , \4849_b1 , w_15602 );
or ( \4932_b0 , \4849_b0 , \4931_b0 );
not ( \4931_b0 , w_15603 );
and ( w_15603 , w_15602 , \4931_b1 );
or ( \4933_b1 , \4848_b1 , w_15604 );
or ( \4933_b0 , \4848_b0 , \4930_b0 );
not ( \4930_b0 , w_15605 );
and ( w_15605 , w_15604 , \4930_b1 );
buf ( \4934_b1 , \2945_b1 );
buf ( \4934_b0 , \2945_b0 );
buf ( \4935_b1 , \4934_b1 );
not ( \4935_b1 , w_15606 );
not ( \4935_b0 , w_15607 );
and ( w_15606 , w_15607 , \4934_b0 );
buf ( \4936_b1 , \4935_b1 );
not ( \4936_b1 , w_15608 );
not ( \4936_b0 , w_15609 );
and ( w_15608 , w_15609 , \4935_b0 );
or ( \4937_b1 , \4051_b1 , \4936_b1 );
not ( \4936_b1 , w_15610 );
and ( \4937_b0 , \4051_b0 , w_15611 );
and ( w_15610 , w_15611 , \4936_b0 );
buf ( \4938_b1 , \4051_b1 );
not ( \4938_b1 , w_15612 );
not ( \4938_b0 , w_15613 );
and ( w_15612 , w_15613 , \4051_b0 );
buf ( \4939_b1 , \4934_b1 );
not ( \4939_b1 , w_15614 );
not ( \4939_b0 , w_15615 );
and ( w_15614 , w_15615 , \4934_b0 );
or ( \4940_b1 , \4938_b1 , \4939_b1 );
not ( \4939_b1 , w_15616 );
and ( \4940_b0 , \4938_b0 , w_15617 );
and ( w_15616 , w_15617 , \4939_b0 );
or ( \4941_b1 , \4937_b1 , w_15619 );
not ( w_15619 , w_15620 );
and ( \4941_b0 , \4937_b0 , w_15621 );
and ( w_15620 ,  , w_15621 );
buf ( w_15619 , \4940_b1 );
not ( w_15619 , w_15622 );
not (  , w_15623 );
and ( w_15622 , w_15623 , \4940_b0 );
buf ( \4942_b1 , \4941_b1 );
not ( \4942_b1 , w_15624 );
not ( \4942_b0 , w_15625 );
and ( w_15624 , w_15625 , \4941_b0 );
or ( \4943_b1 , \4858_b1 , w_15627 );
not ( w_15627 , w_15628 );
and ( \4943_b0 , \4858_b0 , w_15629 );
and ( w_15628 ,  , w_15629 );
buf ( w_15627 , \4862_b1 );
not ( w_15627 , w_15630 );
not (  , w_15631 );
and ( w_15630 , w_15631 , \4862_b0 );
buf ( \4944_b1 , \4943_b1 );
not ( \4944_b1 , w_15632 );
not ( \4944_b0 , w_15633 );
and ( w_15632 , w_15633 , \4943_b0 );
buf ( \4945_b1 , \4944_b1 );
buf ( \4945_b0 , \4944_b0 );
buf ( \4946_b1 , \4945_b1 );
not ( \4946_b1 , w_15634 );
not ( \4946_b0 , w_15635 );
and ( w_15634 , w_15635 , \4945_b0 );
or ( \4947_b1 , \4942_b1 , w_15636 );
or ( \4947_b0 , \4942_b0 , \4946_b0 );
not ( \4946_b0 , w_15637 );
and ( w_15637 , w_15636 , \4946_b1 );
buf ( \4948_b1 , \4862_b1 );
not ( \4948_b1 , w_15638 );
not ( \4948_b0 , w_15639 );
and ( w_15638 , w_15639 , \4862_b0 );
buf ( \4949_b1 , \4939_b1 );
not ( \4949_b1 , w_15640 );
not ( \4949_b0 , w_15641 );
and ( w_15640 , w_15641 , \4939_b0 );
or ( \4950_b1 , \4948_b1 , w_15643 );
not ( w_15643 , w_15644 );
and ( \4950_b0 , \4948_b0 , w_15645 );
and ( w_15644 ,  , w_15645 );
buf ( w_15643 , \4949_b1 );
not ( w_15643 , w_15646 );
not (  , w_15647 );
and ( w_15646 , w_15647 , \4949_b0 );
or ( \4951_b1 , \4947_b1 , w_15649 );
not ( w_15649 , w_15650 );
and ( \4951_b0 , \4947_b0 , w_15651 );
and ( w_15650 ,  , w_15651 );
buf ( w_15649 , \4950_b1 );
not ( w_15649 , w_15652 );
not (  , w_15653 );
and ( w_15652 , w_15653 , \4950_b0 );
buf ( \4952_b1 , \4951_b1 );
not ( \4952_b1 , w_15654 );
not ( \4952_b0 , w_15655 );
and ( w_15654 , w_15655 , \4951_b0 );
buf ( \4953_b1 , \4017_b1 );
not ( \4953_b1 , w_15656 );
not ( \4953_b0 , w_15657 );
and ( w_15656 , w_15657 , \4017_b0 );
buf ( \4954_b1 , \4134_b1 );
not ( \4954_b1 , w_15658 );
not ( \4954_b0 , w_15659 );
and ( w_15658 , w_15659 , \4134_b0 );
or ( \4955_b1 , \4953_b1 , w_15660 );
or ( \4955_b0 , \4953_b0 , \4954_b0 );
not ( \4954_b0 , w_15661 );
and ( w_15661 , w_15660 , \4954_b1 );
or ( \4956_b1 , \4106_b1 , w_15663 );
not ( w_15663 , w_15664 );
and ( \4956_b0 , \4106_b0 , w_15665 );
and ( w_15664 ,  , w_15665 );
buf ( w_15663 , \4662_b1 );
not ( w_15663 , w_15666 );
not (  , w_15667 );
and ( w_15666 , w_15667 , \4662_b0 );
or ( \4957_b1 , \4955_b1 , w_15669 );
not ( w_15669 , w_15670 );
and ( \4957_b0 , \4955_b0 , w_15671 );
and ( w_15670 ,  , w_15671 );
buf ( w_15669 , \4956_b1 );
not ( w_15669 , w_15672 );
not (  , w_15673 );
and ( w_15672 , w_15673 , \4956_b0 );
buf ( \4958_b1 , \4957_b1 );
not ( \4958_b1 , w_15674 );
not ( \4958_b0 , w_15675 );
and ( w_15674 , w_15675 , \4957_b0 );
buf ( \4959_b1 , \4302_b1 );
not ( \4959_b1 , w_15676 );
not ( \4959_b0 , w_15677 );
and ( w_15676 , w_15677 , \4302_b0 );
or ( \4960_b1 , \4958_b1 , w_15678 );
or ( \4960_b0 , \4958_b0 , \4959_b0 );
not ( \4959_b0 , w_15679 );
and ( w_15679 , w_15678 , \4959_b1 );
or ( \4961_b1 , \4654_b1 , w_15681 );
not ( w_15681 , w_15682 );
and ( \4961_b0 , \4654_b0 , w_15683 );
and ( w_15682 ,  , w_15683 );
buf ( w_15681 , \4708_b1 );
not ( w_15681 , w_15684 );
not (  , w_15685 );
and ( w_15684 , w_15685 , \4708_b0 );
or ( \4962_b1 , \4960_b1 , w_15687 );
not ( w_15687 , w_15688 );
and ( \4962_b0 , \4960_b0 , w_15689 );
and ( w_15688 ,  , w_15689 );
buf ( w_15687 , \4961_b1 );
not ( w_15687 , w_15690 );
not (  , w_15691 );
and ( w_15690 , w_15691 , \4961_b0 );
buf ( \4963_b1 , \4962_b1 );
not ( \4963_b1 , w_15692 );
not ( \4963_b0 , w_15693 );
and ( w_15692 , w_15693 , \4962_b0 );
or ( \4964_b1 , \4952_b1 , w_15694 );
or ( \4964_b0 , \4952_b0 , \4963_b0 );
not ( \4963_b0 , w_15695 );
and ( w_15695 , w_15694 , \4963_b1 );
or ( \4965_b1 , \4951_b1 , w_15696 );
or ( \4965_b0 , \4951_b0 , \4962_b0 );
not ( \4962_b0 , w_15697 );
and ( w_15697 , w_15696 , \4962_b1 );
buf ( \4966_b1 , \4026_b1 );
not ( \4966_b1 , w_15698 );
not ( \4966_b0 , w_15699 );
and ( w_15698 , w_15699 , \4026_b0 );
buf ( \4967_b1 , \4250_b1 );
not ( \4967_b1 , w_15700 );
not ( \4967_b0 , w_15701 );
and ( w_15700 , w_15701 , \4250_b0 );
or ( \4968_b1 , \4966_b1 , w_15702 );
or ( \4968_b0 , \4966_b0 , \4967_b0 );
not ( \4967_b0 , w_15703 );
and ( w_15703 , w_15702 , \4967_b1 );
buf ( \4969_b1 , \4026_b1 );
not ( \4969_b1 , w_15704 );
not ( \4969_b0 , w_15705 );
and ( w_15704 , w_15705 , \4026_b0 );
or ( \4970_b1 , \4661_b1 , w_15707 );
not ( w_15707 , w_15708 );
and ( \4970_b0 , \4661_b0 , w_15709 );
and ( w_15708 ,  , w_15709 );
buf ( w_15707 , \4969_b1 );
not ( w_15707 , w_15710 );
not (  , w_15711 );
and ( w_15710 , w_15711 , \4969_b0 );
or ( \4971_b1 , \4968_b1 , w_15713 );
not ( w_15713 , w_15714 );
and ( \4971_b0 , \4968_b0 , w_15715 );
and ( w_15714 ,  , w_15715 );
buf ( w_15713 , \4970_b1 );
not ( w_15713 , w_15716 );
not (  , w_15717 );
and ( w_15716 , w_15717 , \4970_b0 );
buf ( \4972_b1 , \4971_b1 );
not ( \4972_b1 , w_15718 );
not ( \4972_b0 , w_15719 );
and ( w_15718 , w_15719 , \4971_b0 );
buf ( \4973_b1 , \4395_b1 );
not ( \4973_b1 , w_15720 );
not ( \4973_b0 , w_15721 );
and ( w_15720 , w_15721 , \4395_b0 );
or ( \4974_b1 , \4972_b1 , w_15722 );
or ( \4974_b0 , \4972_b0 , \4973_b0 );
not ( \4973_b0 , w_15723 );
and ( w_15723 , w_15722 , \4973_b1 );
or ( \4975_b1 , \4782_b1 , w_15725 );
not ( w_15725 , w_15726 );
and ( \4975_b0 , \4782_b0 , w_15727 );
and ( w_15726 ,  , w_15727 );
buf ( w_15725 , \4200_b1 );
not ( w_15725 , w_15728 );
not (  , w_15729 );
and ( w_15728 , w_15729 , \4200_b0 );
or ( \4976_b1 , \4974_b1 , w_15731 );
not ( w_15731 , w_15732 );
and ( \4976_b0 , \4974_b0 , w_15733 );
and ( w_15732 ,  , w_15733 );
buf ( w_15731 , \4975_b1 );
not ( w_15731 , w_15734 );
not (  , w_15735 );
and ( w_15734 , w_15735 , \4975_b0 );
or ( \4977_b1 , \4965_b1 , w_15737 );
not ( w_15737 , w_15738 );
and ( \4977_b0 , \4965_b0 , w_15739 );
and ( w_15738 ,  , w_15739 );
buf ( w_15737 , \4976_b1 );
not ( w_15737 , w_15740 );
not (  , w_15741 );
and ( w_15740 , w_15741 , \4976_b0 );
or ( \4978_b1 , \4964_b1 , w_15743 );
not ( w_15743 , w_15744 );
and ( \4978_b0 , \4964_b0 , w_15745 );
and ( w_15744 ,  , w_15745 );
buf ( w_15743 , \4977_b1 );
not ( w_15743 , w_15746 );
not (  , w_15747 );
and ( w_15746 , w_15747 , \4977_b0 );
buf ( \4979_b1 , \4978_b1 );
not ( \4979_b1 , w_15748 );
not ( \4979_b0 , w_15749 );
and ( w_15748 , w_15749 , \4978_b0 );
buf ( \4980_b1 , \4979_b1 );
not ( \4980_b1 , w_15750 );
not ( \4980_b0 , w_15751 );
and ( w_15750 , w_15751 , \4979_b0 );
or ( \4981_b1 , \4775_b1 , \4802_b1 );
xor ( \4981_b0 , \4775_b0 , w_15752 );
not ( w_15752 , w_15753 );
and ( w_15753 , \4802_b1 , \4802_b0 );
or ( \4982_b1 , \4981_b1 , w_15754 );
xor ( \4982_b0 , \4981_b0 , w_15756 );
not ( w_15756 , w_15757 );
and ( w_15757 , w_15754 , w_15755 );
buf ( w_15754 , \4787_b1 );
not ( w_15754 , w_15758 );
not ( w_15755 , w_15759 );
and ( w_15758 , w_15759 , \4787_b0 );
buf ( \4983_b1 , \4982_b1 );
not ( \4983_b1 , w_15760 );
not ( \4983_b0 , w_15761 );
and ( w_15760 , w_15761 , \4982_b0 );
or ( \4984_b1 , \4980_b1 , w_15762 );
or ( \4984_b0 , \4980_b0 , \4983_b0 );
not ( \4983_b0 , w_15763 );
and ( w_15763 , w_15762 , \4983_b1 );
buf ( \4985_b1 , \4725_b1 );
not ( \4985_b1 , w_15764 );
not ( \4985_b0 , w_15765 );
and ( w_15764 , w_15765 , \4725_b0 );
buf ( \4986_b1 , \4714_b1 );
not ( \4986_b1 , w_15766 );
not ( \4986_b0 , w_15767 );
and ( w_15766 , w_15767 , \4714_b0 );
buf ( \4987_b1 , \4986_b1 );
not ( \4987_b1 , w_15768 );
not ( \4987_b0 , w_15769 );
and ( w_15768 , w_15769 , \4986_b0 );
or ( \4988_b1 , \4985_b1 , w_15770 );
or ( \4988_b0 , \4985_b0 , \4987_b0 );
not ( \4987_b0 , w_15771 );
and ( w_15771 , w_15770 , \4987_b1 );
buf ( \4989_b1 , \4725_b1 );
not ( \4989_b1 , w_15772 );
not ( \4989_b0 , w_15773 );
and ( w_15772 , w_15773 , \4725_b0 );
or ( \4990_b1 , \4989_b1 , w_15775 );
not ( w_15775 , w_15776 );
and ( \4990_b0 , \4989_b0 , w_15777 );
and ( w_15776 ,  , w_15777 );
buf ( w_15775 , \4714_b1 );
not ( w_15775 , w_15778 );
not (  , w_15779 );
and ( w_15778 , w_15779 , \4714_b0 );
or ( \4991_b1 , \4988_b1 , w_15781 );
not ( w_15781 , w_15782 );
and ( \4991_b0 , \4988_b0 , w_15783 );
and ( w_15782 ,  , w_15783 );
buf ( w_15781 , \4990_b1 );
not ( w_15781 , w_15784 );
not (  , w_15785 );
and ( w_15784 , w_15785 , \4990_b0 );
or ( \4992_b1 , \4991_b1 , \4739_b1 );
not ( \4739_b1 , w_15786 );
and ( \4992_b0 , \4991_b0 , w_15787 );
and ( w_15786 , w_15787 , \4739_b0 );
buf ( \4993_b1 , \4991_b1 );
not ( \4993_b1 , w_15788 );
not ( \4993_b0 , w_15789 );
and ( w_15788 , w_15789 , \4991_b0 );
buf ( \4994_b1 , \4739_b1 );
not ( \4994_b1 , w_15790 );
not ( \4994_b0 , w_15791 );
and ( w_15790 , w_15791 , \4739_b0 );
or ( \4995_b1 , \4993_b1 , \4994_b1 );
not ( \4994_b1 , w_15792 );
and ( \4995_b0 , \4993_b0 , w_15793 );
and ( w_15792 , w_15793 , \4994_b0 );
or ( \4996_b1 , \4992_b1 , w_15795 );
not ( w_15795 , w_15796 );
and ( \4996_b0 , \4992_b0 , w_15797 );
and ( w_15796 ,  , w_15797 );
buf ( w_15795 , \4995_b1 );
not ( w_15795 , w_15798 );
not (  , w_15799 );
and ( w_15798 , w_15799 , \4995_b0 );
or ( \4997_b1 , \4984_b1 , w_15801 );
not ( w_15801 , w_15802 );
and ( \4997_b0 , \4984_b0 , w_15803 );
and ( w_15802 ,  , w_15803 );
buf ( w_15801 , \4996_b1 );
not ( w_15801 , w_15804 );
not (  , w_15805 );
and ( w_15804 , w_15805 , \4996_b0 );
or ( \4998_b1 , \4982_b1 , w_15806 );
or ( \4998_b0 , \4982_b0 , \4979_b0 );
not ( \4979_b0 , w_15807 );
and ( w_15807 , w_15806 , \4979_b1 );
or ( \4999_b1 , \4997_b1 , w_15809 );
not ( w_15809 , w_15810 );
and ( \4999_b0 , \4997_b0 , w_15811 );
and ( w_15810 ,  , w_15811 );
buf ( w_15809 , \4998_b1 );
not ( w_15809 , w_15812 );
not (  , w_15813 );
and ( w_15812 , w_15813 , \4998_b0 );
or ( \5000_b1 , \4933_b1 , w_15815 );
not ( w_15815 , w_15816 );
and ( \5000_b0 , \4933_b0 , w_15817 );
and ( w_15816 ,  , w_15817 );
buf ( w_15815 , \4999_b1 );
not ( w_15815 , w_15818 );
not (  , w_15819 );
and ( w_15818 , w_15819 , \4999_b0 );
or ( \5001_b1 , \4932_b1 , w_15821 );
not ( w_15821 , w_15822 );
and ( \5001_b0 , \4932_b0 , w_15823 );
and ( w_15822 ,  , w_15823 );
buf ( w_15821 , \5000_b1 );
not ( w_15821 , w_15824 );
not (  , w_15825 );
and ( w_15824 , w_15825 , \5000_b0 );
or ( \5002_b1 , \4841_b1 , w_15827 );
not ( w_15827 , w_15828 );
and ( \5002_b0 , \4841_b0 , w_15829 );
and ( w_15828 ,  , w_15829 );
buf ( w_15827 , \5001_b1 );
not ( w_15827 , w_15830 );
not (  , w_15831 );
and ( w_15830 , w_15831 , \5001_b0 );
or ( \5003_b1 , \4840_b1 , w_15833 );
not ( w_15833 , w_15834 );
and ( \5003_b0 , \4840_b0 , w_15835 );
and ( w_15834 ,  , w_15835 );
buf ( w_15833 , \5002_b1 );
not ( w_15833 , w_15836 );
not (  , w_15837 );
and ( w_15836 , w_15837 , \5002_b0 );
or ( \5004_b1 , \4828_b1 , w_15838 );
or ( \5004_b0 , \4828_b0 , \5003_b0 );
not ( \5003_b0 , w_15839 );
and ( w_15839 , w_15838 , \5003_b1 );
or ( \5005_b1 , \4826_b1 , w_15841 );
not ( w_15841 , w_15842 );
and ( \5005_b0 , \4826_b0 , w_15843 );
and ( w_15842 ,  , w_15843 );
buf ( w_15841 , \5004_b1 );
not ( w_15841 , w_15844 );
not (  , w_15845 );
and ( w_15844 , w_15845 , \5004_b0 );
or ( \5006_b1 , \4590_b1 , w_15847 );
not ( w_15847 , w_15848 );
and ( \5006_b0 , \4590_b0 , w_15849 );
and ( w_15848 ,  , w_15849 );
buf ( w_15847 , \5005_b1 );
not ( w_15847 , w_15850 );
not (  , w_15851 );
and ( w_15850 , w_15851 , \5005_b0 );
or ( \5007_b1 , \4418_b1 , \4420_b1 );
xor ( \5007_b0 , \4418_b0 , w_15852 );
not ( w_15852 , w_15853 );
and ( w_15853 , \4420_b1 , \4420_b0 );
or ( \5008_b1 , \5007_b1 , \4487_b1 );
not ( \4487_b1 , w_15854 );
and ( \5008_b0 , \5007_b0 , w_15855 );
and ( w_15854 , w_15855 , \4487_b0 );
or ( \5009_b1 , \4418_b1 , \4420_b1 );
not ( \4420_b1 , w_15856 );
and ( \5009_b0 , \4418_b0 , w_15857 );
and ( w_15856 , w_15857 , \4420_b0 );
or ( \5010_b1 , \5008_b1 , w_15858 );
or ( \5010_b0 , \5008_b0 , \5009_b0 );
not ( \5009_b0 , w_15859 );
and ( w_15859 , w_15858 , \5009_b1 );
or ( \5011_b1 , \4322_b1 , \4325_b1 );
xor ( \5011_b0 , \4322_b0 , w_15860 );
not ( w_15860 , w_15861 );
and ( w_15861 , \4325_b1 , \4325_b0 );
or ( \5012_b1 , \5011_b1 , \4365_b1 );
xor ( \5012_b0 , \5011_b0 , w_15862 );
not ( w_15862 , w_15863 );
and ( w_15863 , \4365_b1 , \4365_b0 );
or ( \5013_b1 , \5010_b1 , w_15864 );
or ( \5013_b0 , \5010_b0 , \5012_b0 );
not ( \5012_b0 , w_15865 );
and ( w_15865 , w_15864 , \5012_b1 );
or ( \5014_b1 , \5006_b1 , w_15867 );
not ( w_15867 , w_15868 );
and ( \5014_b0 , \5006_b0 , w_15869 );
and ( w_15868 ,  , w_15869 );
buf ( w_15867 , \5013_b1 );
not ( w_15867 , w_15870 );
not (  , w_15871 );
and ( w_15870 , w_15871 , \5013_b0 );
or ( \5015_b1 , \4371_b1 , w_15873 );
not ( w_15873 , w_15874 );
and ( \5015_b0 , \4371_b0 , w_15875 );
and ( w_15874 ,  , w_15875 );
buf ( w_15873 , \5014_b1 );
not ( w_15873 , w_15876 );
not (  , w_15877 );
and ( w_15876 , w_15877 , \5014_b0 );
or ( \5016_b1 , \4230_b1 , w_15878 );
or ( \5016_b0 , \4230_b0 , \4166_b0 );
not ( \4166_b0 , w_15879 );
and ( w_15879 , w_15878 , \4166_b1 );
or ( \5017_b1 , \5016_b1 , w_15881 );
not ( w_15881 , w_15882 );
and ( \5017_b0 , \5016_b0 , w_15883 );
and ( w_15882 ,  , w_15883 );
buf ( w_15881 , \4292_b1 );
not ( w_15881 , w_15884 );
not (  , w_15885 );
and ( w_15884 , w_15885 , \4292_b0 );
or ( \5018_b1 , \4166_b1 , w_15887 );
not ( w_15887 , w_15888 );
and ( \5018_b0 , \4166_b0 , w_15889 );
and ( w_15888 ,  , w_15889 );
buf ( w_15887 , \4230_b1 );
not ( w_15887 , w_15890 );
not (  , w_15891 );
and ( w_15890 , w_15891 , \4230_b0 );
or ( \5019_b1 , \5017_b1 , w_15893 );
not ( w_15893 , w_15894 );
and ( \5019_b0 , \5017_b0 , w_15895 );
and ( w_15894 ,  , w_15895 );
buf ( w_15893 , \5018_b1 );
not ( w_15893 , w_15896 );
not (  , w_15897 );
and ( w_15896 , w_15897 , \5018_b0 );
or ( \5020_b1 , \4103_b1 , \4141_b1 );
xor ( \5020_b0 , \4103_b0 , w_15898 );
not ( w_15898 , w_15899 );
and ( w_15899 , \4141_b1 , \4141_b0 );
or ( \5021_b1 , \5020_b1 , \4165_b1 );
not ( \4165_b1 , w_15900 );
and ( \5021_b0 , \5020_b0 , w_15901 );
and ( w_15900 , w_15901 , \4165_b0 );
or ( \5022_b1 , \4103_b1 , \4141_b1 );
not ( \4141_b1 , w_15902 );
and ( \5022_b0 , \4103_b0 , w_15903 );
and ( w_15902 , w_15903 , \4141_b0 );
or ( \5023_b1 , \5021_b1 , w_15904 );
or ( \5023_b0 , \5021_b0 , \5022_b0 );
not ( \5022_b0 , w_15905 );
and ( w_15905 , w_15904 , \5022_b1 );
or ( \5024_b1 , \4094_b1 , \4100_b1 );
not ( \4100_b1 , w_15906 );
and ( \5024_b0 , \4094_b0 , w_15907 );
and ( w_15906 , w_15907 , \4100_b0 );
or ( \5025_b1 , \4129_b1 , w_15909 );
not ( w_15909 , w_15910 );
and ( \5025_b0 , \4129_b0 , w_15911 );
and ( w_15910 ,  , w_15911 );
buf ( w_15909 , \4139_b1 );
not ( w_15909 , w_15912 );
not (  , w_15913 );
and ( w_15912 , w_15913 , \4139_b0 );
or ( \5026_b1 , \4133_b1 , w_15915 );
not ( w_15915 , w_15916 );
and ( \5026_b0 , \4133_b0 , w_15917 );
and ( w_15916 ,  , w_15917 );
buf ( w_15915 , \4106_b1 );
not ( w_15915 , w_15918 );
not (  , w_15919 );
and ( w_15918 , w_15919 , \4106_b0 );
or ( \5027_b1 , \5025_b1 , \5026_b1 );
not ( \5026_b1 , w_15920 );
and ( \5027_b0 , \5025_b0 , w_15921 );
and ( w_15920 , w_15921 , \5026_b0 );
or ( \5028_b1 , \5024_b1 , \5027_b1 );
xor ( \5028_b0 , \5024_b0 , w_15922 );
not ( w_15922 , w_15923 );
and ( w_15923 , \5027_b1 , \5027_b0 );
buf ( \5029_b1 , \4195_b1 );
not ( \5029_b1 , w_15924 );
not ( \5029_b0 , w_15925 );
and ( w_15924 , w_15925 , \4195_b0 );
buf ( \5030_b1 , \4199_b1 );
not ( \5030_b1 , w_15926 );
not ( \5030_b0 , w_15927 );
and ( w_15926 , w_15927 , \4199_b0 );
or ( \5031_b1 , \5029_b1 , w_15928 );
or ( \5031_b0 , \5029_b0 , \5030_b0 );
not ( \5030_b0 , w_15929 );
and ( w_15929 , w_15928 , \5030_b1 );
or ( \5032_b1 , \4102_b1 , \4111_b1 );
not ( \4111_b1 , w_15930 );
and ( \5032_b0 , \4102_b0 , w_15931 );
and ( w_15930 , w_15931 , \4111_b0 );
buf ( \5033_b1 , \4102_b1 );
not ( \5033_b1 , w_15932 );
not ( \5033_b0 , w_15933 );
and ( w_15932 , w_15933 , \4102_b0 );
or ( \5034_b1 , \5033_b1 , \3997_b1 );
not ( \3997_b1 , w_15934 );
and ( \5034_b0 , \5033_b0 , w_15935 );
and ( w_15934 , w_15935 , \3997_b0 );
or ( \5035_b1 , \5032_b1 , w_15937 );
not ( w_15937 , w_15938 );
and ( \5035_b0 , \5032_b0 , w_15939 );
and ( w_15938 ,  , w_15939 );
buf ( w_15937 , \5034_b1 );
not ( w_15937 , w_15940 );
not (  , w_15941 );
and ( w_15940 , w_15941 , \5034_b0 );
or ( \5036_b1 , \5035_b1 , w_15942 );
or ( \5036_b0 , \5035_b0 , \4192_b0 );
not ( \4192_b0 , w_15943 );
and ( w_15943 , w_15942 , \4192_b1 );
or ( \5037_b1 , \5031_b1 , w_15945 );
not ( w_15945 , w_15946 );
and ( \5037_b0 , \5031_b0 , w_15947 );
and ( w_15946 ,  , w_15947 );
buf ( w_15945 , \5036_b1 );
not ( w_15945 , w_15948 );
not (  , w_15949 );
and ( w_15948 , w_15949 , \5036_b0 );
or ( \5038_b1 , \5028_b1 , \5037_b1 );
xor ( \5038_b0 , \5028_b0 , w_15950 );
not ( w_15950 , w_15951 );
and ( w_15951 , \5037_b1 , \5037_b0 );
or ( \5039_b1 , \5023_b1 , \5038_b1 );
xor ( \5039_b0 , \5023_b0 , w_15952 );
not ( w_15952 , w_15953 );
and ( w_15953 , \5038_b1 , \5038_b0 );
or ( \5040_b1 , \4177_b1 , \4202_b1 );
xor ( \5040_b0 , \4177_b0 , w_15954 );
not ( w_15954 , w_15955 );
and ( w_15955 , \4202_b1 , \4202_b0 );
or ( \5041_b1 , \5040_b1 , \4229_b1 );
not ( \4229_b1 , w_15956 );
and ( \5041_b0 , \5040_b0 , w_15957 );
and ( w_15956 , w_15957 , \4229_b0 );
or ( \5042_b1 , \4177_b1 , \4202_b1 );
not ( \4202_b1 , w_15958 );
and ( \5042_b0 , \4177_b0 , w_15959 );
and ( w_15958 , w_15959 , \4202_b0 );
or ( \5043_b1 , \5041_b1 , w_15960 );
or ( \5043_b0 , \5041_b0 , \5042_b0 );
not ( \5042_b0 , w_15961 );
and ( w_15961 , w_15960 , \5042_b1 );
or ( \5044_b1 , \5039_b1 , \5043_b1 );
xor ( \5044_b0 , \5039_b0 , w_15962 );
not ( w_15962 , w_15963 );
and ( w_15963 , \5043_b1 , \5043_b0 );
or ( \5045_b1 , \5019_b1 , w_15964 );
or ( \5045_b0 , \5019_b0 , \5044_b0 );
not ( \5044_b0 , w_15965 );
and ( w_15965 , w_15964 , \5044_b1 );
or ( \5046_b1 , \5015_b1 , w_15967 );
not ( w_15967 , w_15968 );
and ( \5046_b0 , \5015_b0 , w_15969 );
and ( w_15968 ,  , w_15969 );
buf ( w_15967 , \5045_b1 );
not ( w_15967 , w_15970 );
not (  , w_15971 );
and ( w_15970 , w_15971 , \5045_b0 );
or ( \5047_b1 , \5023_b1 , \5038_b1 );
xor ( \5047_b0 , \5023_b0 , w_15972 );
not ( w_15972 , w_15973 );
and ( w_15973 , \5038_b1 , \5038_b0 );
or ( \5048_b1 , \5047_b1 , \5043_b1 );
not ( \5043_b1 , w_15974 );
and ( \5048_b0 , \5047_b0 , w_15975 );
and ( w_15974 , w_15975 , \5043_b0 );
or ( \5049_b1 , \5023_b1 , \5038_b1 );
not ( \5038_b1 , w_15976 );
and ( \5049_b0 , \5023_b0 , w_15977 );
and ( w_15976 , w_15977 , \5038_b0 );
or ( \5050_b1 , \5048_b1 , w_15978 );
or ( \5050_b0 , \5048_b0 , \5049_b0 );
not ( \5049_b0 , w_15979 );
and ( w_15979 , w_15978 , \5049_b1 );
buf ( \5051_b1 , \5027_b1 );
not ( \5051_b1 , w_15980 );
not ( \5051_b0 , w_15981 );
and ( w_15980 , w_15981 , \5027_b0 );
or ( \5052_b1 , \5024_b1 , \5027_b1 );
xor ( \5052_b0 , \5024_b0 , w_15982 );
not ( w_15982 , w_15983 );
and ( w_15983 , \5027_b1 , \5027_b0 );
or ( \5053_b1 , \5052_b1 , \5037_b1 );
not ( \5037_b1 , w_15984 );
and ( \5053_b0 , \5052_b0 , w_15985 );
and ( w_15984 , w_15985 , \5037_b0 );
or ( \5054_b1 , \5024_b1 , \5027_b1 );
not ( \5027_b1 , w_15986 );
and ( \5054_b0 , \5024_b0 , w_15987 );
and ( w_15986 , w_15987 , \5027_b0 );
or ( \5055_b1 , \5053_b1 , w_15988 );
or ( \5055_b0 , \5053_b0 , \5054_b0 );
not ( \5054_b0 , w_15989 );
and ( w_15989 , w_15988 , \5054_b1 );
or ( \5056_b1 , \5051_b1 , \5055_b1 );
xor ( \5056_b0 , \5051_b0 , w_15990 );
not ( w_15990 , w_15991 );
and ( w_15991 , \5055_b1 , \5055_b0 );
or ( \5057_b1 , \4198_b1 , \4102_b1 );
not ( \4102_b1 , w_15992 );
and ( \5057_b0 , \4198_b0 , w_15993 );
and ( w_15992 , w_15993 , \4102_b0 );
or ( \5058_b1 , \4133_b1 , w_15994 );
or ( \5058_b0 , \4133_b0 , \4302_b0 );
not ( \4302_b0 , w_15995 );
and ( w_15995 , w_15994 , \4302_b1 );
or ( \5059_b1 , \5058_b1 , w_15997 );
not ( w_15997 , w_15998 );
and ( \5059_b0 , \5058_b0 , w_15999 );
and ( w_15998 ,  , w_15999 );
buf ( w_15997 , \4106_b1 );
not ( w_15997 , w_16000 );
not (  , w_16001 );
and ( w_16000 , w_16001 , \4106_b0 );
or ( \5060_b1 , \5057_b1 , \5059_b1 );
xor ( \5060_b0 , \5057_b0 , w_16002 );
not ( w_16002 , w_16003 );
and ( w_16003 , \5059_b1 , \5059_b0 );
or ( \5061_b1 , \5029_b1 , w_16004 );
or ( \5061_b0 , \5029_b0 , \5035_b0 );
not ( \5035_b0 , w_16005 );
and ( w_16005 , w_16004 , \5035_b1 );
or ( \5062_b1 , \4101_b1 , \4051_b1 );
not ( \4051_b1 , w_16006 );
and ( \5062_b0 , \4101_b0 , w_16007 );
and ( w_16006 , w_16007 , \4051_b0 );
or ( \5063_b1 , \4102_b1 , \4135_b1 );
not ( \4135_b1 , w_16008 );
and ( \5063_b0 , \4102_b0 , w_16009 );
and ( w_16008 , w_16009 , \4135_b0 );
or ( \5064_b1 , \5062_b1 , w_16011 );
not ( w_16011 , w_16012 );
and ( \5064_b0 , \5062_b0 , w_16013 );
and ( w_16012 ,  , w_16013 );
buf ( w_16011 , \5063_b1 );
not ( w_16011 , w_16014 );
not (  , w_16015 );
and ( w_16014 , w_16015 , \5063_b0 );
or ( \5065_b1 , \5064_b1 , w_16016 );
or ( \5065_b0 , \5064_b0 , \4192_b0 );
not ( \4192_b0 , w_16017 );
and ( w_16017 , w_16016 , \4192_b1 );
or ( \5066_b1 , \5061_b1 , w_16019 );
not ( w_16019 , w_16020 );
and ( \5066_b0 , \5061_b0 , w_16021 );
and ( w_16020 ,  , w_16021 );
buf ( w_16019 , \5065_b1 );
not ( w_16019 , w_16022 );
not (  , w_16023 );
and ( w_16022 , w_16023 , \5065_b0 );
or ( \5067_b1 , \5060_b1 , \5066_b1 );
xor ( \5067_b0 , \5060_b0 , w_16024 );
not ( w_16024 , w_16025 );
and ( w_16025 , \5066_b1 , \5066_b0 );
or ( \5068_b1 , \5056_b1 , \5067_b1 );
xor ( \5068_b0 , \5056_b0 , w_16026 );
not ( w_16026 , w_16027 );
and ( w_16027 , \5067_b1 , \5067_b0 );
or ( \5069_b1 , \5050_b1 , w_16029 );
not ( w_16029 , w_16030 );
and ( \5069_b0 , \5050_b0 , w_16031 );
and ( w_16030 ,  , w_16031 );
buf ( w_16029 , \5068_b1 );
not ( w_16029 , w_16032 );
not (  , w_16033 );
and ( w_16032 , w_16033 , \5068_b0 );
or ( \5070_b1 , \5046_b1 , w_16035 );
not ( w_16035 , w_16036 );
and ( \5070_b0 , \5046_b0 , w_16037 );
and ( w_16036 ,  , w_16037 );
buf ( w_16035 , \5069_b1 );
not ( w_16035 , w_16038 );
not (  , w_16039 );
and ( w_16038 , w_16039 , \5069_b0 );
buf ( \5071_b1 , \5070_b1 );
not ( \5071_b1 , w_16040 );
not ( \5071_b0 , w_16041 );
and ( w_16040 , w_16041 , \5070_b0 );
or ( \5072_b1 , \4962_b1 , \4976_b1 );
xor ( \5072_b0 , \4962_b0 , w_16042 );
not ( w_16042 , w_16043 );
and ( w_16043 , \4976_b1 , \4976_b0 );
buf ( \5073_b1 , \4951_b1 );
buf ( \5073_b0 , \4951_b0 );
buf ( \5074_b1 , \5073_b1 );
not ( \5074_b1 , w_16044 );
not ( \5074_b0 , w_16045 );
and ( w_16044 , w_16045 , \5073_b0 );
or ( \5075_b1 , \5072_b1 , \5074_b1 );
not ( \5074_b1 , w_16046 );
and ( \5075_b0 , \5072_b0 , w_16047 );
and ( w_16046 , w_16047 , \5074_b0 );
buf ( \5076_b1 , \5072_b1 );
not ( \5076_b1 , w_16048 );
not ( \5076_b0 , w_16049 );
and ( w_16048 , w_16049 , \5072_b0 );
or ( \5077_b1 , \5076_b1 , \5073_b1 );
not ( \5073_b1 , w_16050 );
and ( \5077_b0 , \5076_b0 , w_16051 );
and ( w_16050 , w_16051 , \5073_b0 );
or ( \5078_b1 , \5075_b1 , w_16053 );
not ( w_16053 , w_16054 );
and ( \5078_b0 , \5075_b0 , w_16055 );
and ( w_16054 ,  , w_16055 );
buf ( w_16053 , \5077_b1 );
not ( w_16053 , w_16056 );
not (  , w_16057 );
and ( w_16056 , w_16057 , \5077_b0 );
buf ( \5079_b1 , \5078_b1 );
not ( \5079_b1 , w_16058 );
not ( \5079_b0 , w_16059 );
and ( w_16058 , w_16059 , \5078_b0 );
buf ( \5080_b1 , \5079_b1 );
not ( \5080_b1 , w_16060 );
not ( \5080_b0 , w_16061 );
and ( w_16060 , w_16061 , \5079_b0 );
or ( \5081_b1 , \4913_b1 , \4902_b1 );
xor ( \5081_b0 , \4913_b0 , w_16062 );
not ( w_16062 , w_16063 );
and ( w_16063 , \4902_b1 , \4902_b0 );
buf ( \5082_b1 , \4926_b1 );
buf ( \5082_b0 , \4926_b0 );
or ( \5083_b1 , \5081_b1 , w_16064 );
xor ( \5083_b0 , \5081_b0 , w_16066 );
not ( w_16066 , w_16067 );
and ( w_16067 , w_16064 , w_16065 );
buf ( w_16064 , \5082_b1 );
not ( w_16064 , w_16068 );
not ( w_16065 , w_16069 );
and ( w_16068 , w_16069 , \5082_b0 );
or ( \5084_b1 , \5080_b1 , w_16071 );
not ( w_16071 , w_16072 );
and ( \5084_b0 , \5080_b0 , w_16073 );
and ( w_16072 ,  , w_16073 );
buf ( w_16071 , \5083_b1 );
not ( w_16071 , w_16074 );
not (  , w_16075 );
and ( w_16074 , w_16075 , \5083_b0 );
buf ( \5085_b1 , \5074_b1 );
not ( \5085_b1 , w_16076 );
not ( \5085_b0 , w_16077 );
and ( w_16076 , w_16077 , \5074_b0 );
buf ( \5086_b1 , \4072_b1 );
not ( \5086_b1 , w_16078 );
not ( \5086_b0 , w_16079 );
and ( w_16078 , w_16079 , \4072_b0 );
buf ( \5087_b1 , \4250_b1 );
not ( \5087_b1 , w_16080 );
not ( \5087_b0 , w_16081 );
and ( w_16080 , w_16081 , \4250_b0 );
or ( \5088_b1 , \5086_b1 , w_16082 );
or ( \5088_b0 , \5086_b0 , \5087_b0 );
not ( \5087_b0 , w_16083 );
and ( w_16083 , w_16082 , \5087_b1 );
buf ( \5089_b1 , \4072_b1 );
not ( \5089_b1 , w_16084 );
not ( \5089_b0 , w_16085 );
and ( w_16084 , w_16085 , \4072_b0 );
or ( \5090_b1 , \4661_b1 , w_16087 );
not ( w_16087 , w_16088 );
and ( \5090_b0 , \4661_b0 , w_16089 );
and ( w_16088 ,  , w_16089 );
buf ( w_16087 , \5089_b1 );
not ( w_16087 , w_16090 );
not (  , w_16091 );
and ( w_16090 , w_16091 , \5089_b0 );
or ( \5091_b1 , \5088_b1 , w_16093 );
not ( w_16093 , w_16094 );
and ( \5091_b0 , \5088_b0 , w_16095 );
and ( w_16094 ,  , w_16095 );
buf ( w_16093 , \5090_b1 );
not ( w_16093 , w_16096 );
not (  , w_16097 );
and ( w_16096 , w_16097 , \5090_b0 );
buf ( \5092_b1 , \5091_b1 );
not ( \5092_b1 , w_16098 );
not ( \5092_b0 , w_16099 );
and ( w_16098 , w_16099 , \5091_b0 );
buf ( \5093_b1 , \4395_b1 );
not ( \5093_b1 , w_16100 );
not ( \5093_b0 , w_16101 );
and ( w_16100 , w_16101 , \4395_b0 );
or ( \5094_b1 , \5092_b1 , w_16102 );
or ( \5094_b0 , \5092_b0 , \5093_b0 );
not ( \5093_b0 , w_16103 );
and ( w_16103 , w_16102 , \5093_b1 );
or ( \5095_b1 , \4971_b1 , w_16105 );
not ( w_16105 , w_16106 );
and ( \5095_b0 , \4971_b0 , w_16107 );
and ( w_16106 ,  , w_16107 );
buf ( w_16105 , \4200_b1 );
not ( w_16105 , w_16108 );
not (  , w_16109 );
and ( w_16108 , w_16109 , \4200_b0 );
or ( \5096_b1 , \5094_b1 , w_16111 );
not ( w_16111 , w_16112 );
and ( \5096_b0 , \5094_b0 , w_16113 );
and ( w_16112 ,  , w_16113 );
buf ( w_16111 , \5095_b1 );
not ( w_16111 , w_16114 );
not (  , w_16115 );
and ( w_16114 , w_16115 , \5095_b0 );
buf ( \5097_b1 , \5096_b1 );
not ( \5097_b1 , w_16116 );
not ( \5097_b0 , w_16117 );
and ( w_16116 , w_16117 , \5096_b0 );
or ( \5098_b1 , \5085_b1 , w_16118 );
or ( \5098_b0 , \5085_b0 , \5097_b0 );
not ( \5097_b0 , w_16119 );
and ( w_16119 , w_16118 , \5097_b1 );
buf ( \5099_b1 , \4951_b1 );
not ( \5099_b1 , w_16120 );
not ( \5099_b0 , w_16121 );
and ( w_16120 , w_16121 , \4951_b0 );
buf ( \5100_b1 , \5096_b1 );
not ( \5100_b1 , w_16122 );
not ( \5100_b0 , w_16123 );
and ( w_16122 , w_16123 , \5096_b0 );
buf ( \5101_b1 , \5100_b1 );
not ( \5101_b1 , w_16124 );
not ( \5101_b0 , w_16125 );
and ( w_16124 , w_16125 , \5100_b0 );
or ( \5102_b1 , \5099_b1 , w_16126 );
or ( \5102_b0 , \5099_b0 , \5101_b0 );
not ( \5101_b0 , w_16127 );
and ( w_16127 , w_16126 , \5101_b1 );
buf ( \5103_b1 , \3997_b1 );
not ( \5103_b1 , w_16128 );
not ( \5103_b0 , w_16129 );
and ( w_16128 , w_16129 , \3997_b0 );
buf ( \5104_b1 , \4939_b1 );
not ( \5104_b1 , w_16130 );
not ( \5104_b0 , w_16131 );
and ( w_16130 , w_16131 , \4939_b0 );
or ( \5105_b1 , \5103_b1 , w_16132 );
or ( \5105_b0 , \5103_b0 , \5104_b0 );
not ( \5104_b0 , w_16133 );
and ( w_16133 , w_16132 , \5104_b1 );
or ( \5106_b1 , \4867_b1 , w_16135 );
not ( w_16135 , w_16136 );
and ( \5106_b0 , \4867_b0 , w_16137 );
and ( w_16136 ,  , w_16137 );
buf ( w_16135 , \4111_b1 );
not ( w_16135 , w_16138 );
not (  , w_16139 );
and ( w_16138 , w_16139 , \4111_b0 );
or ( \5107_b1 , \5105_b1 , w_16141 );
not ( w_16141 , w_16142 );
and ( \5107_b0 , \5105_b0 , w_16143 );
and ( w_16142 ,  , w_16143 );
buf ( w_16141 , \5106_b1 );
not ( w_16141 , w_16144 );
not (  , w_16145 );
and ( w_16144 , w_16145 , \5106_b0 );
or ( \5108_b1 , \4945_b1 , \5107_b1 );
not ( \5107_b1 , w_16146 );
and ( \5108_b0 , \4945_b0 , w_16147 );
and ( w_16146 , w_16147 , \5107_b0 );
or ( \5109_b1 , \4863_b1 , \4941_b1 );
not ( \4941_b1 , w_16148 );
and ( \5109_b0 , \4863_b0 , w_16149 );
and ( w_16148 , w_16149 , \4941_b0 );
or ( \5110_b1 , \5108_b1 , w_16151 );
not ( w_16151 , w_16152 );
and ( \5110_b0 , \5108_b0 , w_16153 );
and ( w_16152 ,  , w_16153 );
buf ( w_16151 , \5109_b1 );
not ( w_16151 , w_16154 );
not (  , w_16155 );
and ( w_16154 , w_16155 , \5109_b0 );
buf ( \5111_b1 , \4097_b1 );
not ( \5111_b1 , w_16156 );
not ( \5111_b0 , w_16157 );
and ( w_16156 , w_16157 , \4097_b0 );
buf ( \5112_b1 , \4729_b1 );
not ( \5112_b1 , w_16158 );
not ( \5112_b0 , w_16159 );
and ( w_16158 , w_16159 , \4729_b0 );
buf ( \5113_b1 , \5112_b1 );
not ( \5113_b1 , w_16160 );
not ( \5113_b0 , w_16161 );
and ( w_16160 , w_16161 , \5112_b0 );
or ( \5114_b1 , \5111_b1 , w_16162 );
or ( \5114_b0 , \5111_b0 , \5113_b0 );
not ( \5113_b0 , w_16163 );
and ( w_16163 , w_16162 , \5113_b1 );
or ( \5115_b1 , \4458_b1 , w_16165 );
not ( w_16165 , w_16166 );
and ( \5115_b0 , \4458_b0 , w_16167 );
and ( w_16166 ,  , w_16167 );
buf ( w_16165 , \4254_b1 );
not ( w_16165 , w_16168 );
not (  , w_16169 );
and ( w_16168 , w_16169 , \4254_b0 );
or ( \5116_b1 , \5114_b1 , w_16171 );
not ( w_16171 , w_16172 );
and ( \5116_b0 , \5114_b0 , w_16173 );
and ( w_16172 ,  , w_16173 );
buf ( w_16171 , \5115_b1 );
not ( w_16171 , w_16174 );
not (  , w_16175 );
and ( w_16174 , w_16175 , \5115_b0 );
or ( \5117_b1 , \5116_b1 , \4632_b1 );
not ( \4632_b1 , w_16176 );
and ( \5117_b0 , \5116_b0 , w_16177 );
and ( w_16176 , w_16177 , \4632_b0 );
buf ( \5118_b1 , \4096_b1 );
not ( \5118_b1 , w_16178 );
not ( \5118_b0 , w_16179 );
and ( w_16178 , w_16179 , \4096_b0 );
buf ( \5119_b1 , \4535_b1 );
not ( \5119_b1 , w_16180 );
not ( \5119_b0 , w_16181 );
and ( w_16180 , w_16181 , \4535_b0 );
or ( \5120_b1 , \5118_b1 , w_16182 );
or ( \5120_b0 , \5118_b0 , \5119_b0 );
not ( \5119_b0 , w_16183 );
and ( w_16183 , w_16182 , \5119_b1 );
or ( \5121_b1 , \4536_b1 , w_16185 );
not ( w_16185 , w_16186 );
and ( \5121_b0 , \4536_b0 , w_16187 );
and ( w_16186 ,  , w_16187 );
buf ( w_16185 , \4372_b1 );
not ( w_16185 , w_16188 );
not (  , w_16189 );
and ( w_16188 , w_16189 , \4372_b0 );
or ( \5122_b1 , \5120_b1 , w_16191 );
not ( w_16191 , w_16192 );
and ( \5122_b0 , \5120_b0 , w_16193 );
and ( w_16192 ,  , w_16193 );
buf ( w_16191 , \5121_b1 );
not ( w_16191 , w_16194 );
not (  , w_16195 );
and ( w_16194 , w_16195 , \5121_b0 );
or ( \5123_b1 , \5122_b1 , \4453_b1 );
not ( \4453_b1 , w_16196 );
and ( \5123_b0 , \5122_b0 , w_16197 );
and ( w_16196 , w_16197 , \4453_b0 );
or ( \5124_b1 , \5117_b1 , w_16199 );
not ( w_16199 , w_16200 );
and ( \5124_b0 , \5117_b0 , w_16201 );
and ( w_16200 ,  , w_16201 );
buf ( w_16199 , \5123_b1 );
not ( w_16199 , w_16202 );
not (  , w_16203 );
and ( w_16202 , w_16203 , \5123_b0 );
or ( \5125_b1 , \5110_b1 , w_16205 );
not ( w_16205 , w_16206 );
and ( \5125_b0 , \5110_b0 , w_16207 );
and ( w_16206 ,  , w_16207 );
buf ( w_16205 , \5124_b1 );
not ( w_16205 , w_16208 );
not (  , w_16209 );
and ( w_16208 , w_16209 , \5124_b0 );
or ( \5126_b1 , \5102_b1 , w_16211 );
not ( w_16211 , w_16212 );
and ( \5126_b0 , \5102_b0 , w_16213 );
and ( w_16212 ,  , w_16213 );
buf ( w_16211 , \5125_b1 );
not ( w_16211 , w_16214 );
not (  , w_16215 );
and ( w_16214 , w_16215 , \5125_b0 );
or ( \5127_b1 , \5098_b1 , w_16217 );
not ( w_16217 , w_16218 );
and ( \5127_b0 , \5098_b0 , w_16219 );
and ( w_16218 ,  , w_16219 );
buf ( w_16217 , \5126_b1 );
not ( w_16217 , w_16220 );
not (  , w_16221 );
and ( w_16220 , w_16221 , \5126_b0 );
or ( \5128_b1 , \5084_b1 , \5127_b1 );
not ( \5127_b1 , w_16222 );
and ( \5128_b0 , \5084_b0 , w_16223 );
and ( w_16222 , w_16223 , \5127_b0 );
or ( \5129_b1 , \5080_b1 , w_16225 );
not ( w_16225 , w_16226 );
and ( \5129_b0 , \5080_b0 , w_16227 );
and ( w_16226 ,  , w_16227 );
buf ( w_16225 , \5083_b1 );
not ( w_16225 , w_16228 );
not (  , w_16229 );
and ( w_16228 , w_16229 , \5083_b0 );
or ( \5130_b1 , \5128_b1 , w_16231 );
not ( w_16231 , w_16232 );
and ( \5130_b0 , \5128_b0 , w_16233 );
and ( w_16232 ,  , w_16233 );
buf ( w_16231 , \5129_b1 );
not ( w_16231 , w_16234 );
not (  , w_16235 );
and ( w_16234 , w_16235 , \5129_b0 );
or ( \5131_b1 , \4757_b1 , \4898_b1 );
xor ( \5131_b0 , \4757_b0 , w_16236 );
not ( w_16236 , w_16237 );
and ( w_16237 , \4898_b1 , \4898_b0 );
or ( \5132_b1 , \5131_b1 , w_16238 );
xor ( \5132_b0 , \5131_b0 , w_16240 );
not ( w_16240 , w_16241 );
and ( w_16241 , w_16238 , w_16239 );
buf ( w_16238 , \4928_b1 );
not ( w_16238 , w_16242 );
not ( w_16239 , w_16243 );
and ( w_16242 , w_16243 , \4928_b0 );
buf ( \5133_b1 , \4250_b1 );
not ( \5133_b1 , w_16244 );
not ( \5133_b0 , w_16245 );
and ( w_16244 , w_16245 , \4250_b0 );
or ( \5134_b1 , \5133_b1 , w_16247 );
not ( w_16247 , w_16248 );
and ( \5134_b0 , \5133_b0 , w_16249 );
and ( w_16248 ,  , w_16249 );
buf ( w_16247 , \4076_b1 );
not ( w_16247 , w_16250 );
not (  , w_16251 );
and ( w_16250 , w_16251 , \4076_b0 );
buf ( \5135_b1 , \5134_b1 );
not ( \5135_b1 , w_16252 );
not ( \5135_b0 , w_16253 );
and ( w_16252 , w_16253 , \5134_b0 );
buf ( \5136_b1 , \5135_b1 );
not ( \5136_b1 , w_16254 );
not ( \5136_b0 , w_16255 );
and ( w_16254 , w_16255 , \5135_b0 );
buf ( \5137_b1 , \4198_b1 );
not ( \5137_b1 , w_16256 );
not ( \5137_b0 , w_16257 );
and ( w_16256 , w_16257 , \4198_b0 );
buf ( \5138_b1 , \4615_b1 );
not ( \5138_b1 , w_16258 );
not ( \5138_b0 , w_16259 );
and ( w_16258 , w_16259 , \4615_b0 );
buf ( \5139_b1 , \5138_b1 );
not ( \5139_b1 , w_16260 );
not ( \5139_b0 , w_16261 );
and ( w_16260 , w_16261 , \5138_b0 );
or ( \5140_b1 , \5137_b1 , w_16262 );
or ( \5140_b0 , \5137_b0 , \5139_b0 );
not ( \5139_b0 , w_16263 );
and ( w_16263 , w_16262 , \5139_b1 );
or ( \5141_b1 , \4616_b1 , w_16265 );
not ( w_16265 , w_16266 );
and ( \5141_b0 , \4616_b0 , w_16267 );
and ( w_16266 ,  , w_16267 );
buf ( w_16265 , \4209_b1 );
not ( w_16265 , w_16268 );
not (  , w_16269 );
and ( w_16268 , w_16269 , \4209_b0 );
or ( \5142_b1 , \5140_b1 , w_16271 );
not ( w_16271 , w_16272 );
and ( \5142_b0 , \5140_b0 , w_16273 );
and ( w_16272 ,  , w_16273 );
buf ( w_16271 , \5141_b1 );
not ( w_16271 , w_16274 );
not (  , w_16275 );
and ( w_16274 , w_16275 , \5141_b0 );
buf ( \5143_b1 , \5142_b1 );
not ( \5143_b1 , w_16276 );
not ( \5143_b0 , w_16277 );
and ( w_16276 , w_16277 , \5142_b0 );
buf ( \5144_b1 , \4611_b1 );
not ( \5144_b1 , w_16278 );
not ( \5144_b0 , w_16279 );
and ( w_16278 , w_16279 , \4611_b0 );
or ( \5145_b1 , \5143_b1 , w_16280 );
or ( \5145_b0 , \5143_b0 , \5144_b0 );
not ( \5144_b0 , w_16281 );
and ( w_16281 , w_16280 , \5144_b1 );
buf ( \5146_b1 , \4602_b1 );
not ( \5146_b1 , w_16282 );
not ( \5146_b0 , w_16283 );
and ( w_16282 , w_16283 , \4602_b0 );
or ( \5147_b1 , \4878_b1 , w_16285 );
not ( w_16285 , w_16286 );
and ( \5147_b0 , \4878_b0 , w_16287 );
and ( w_16286 ,  , w_16287 );
buf ( w_16285 , \5146_b1 );
not ( w_16285 , w_16288 );
not (  , w_16289 );
and ( w_16288 , w_16289 , \5146_b0 );
or ( \5148_b1 , \5145_b1 , w_16291 );
not ( w_16291 , w_16292 );
and ( \5148_b0 , \5145_b0 , w_16293 );
and ( w_16292 ,  , w_16293 );
buf ( w_16291 , \5147_b1 );
not ( w_16291 , w_16294 );
not (  , w_16295 );
and ( w_16294 , w_16295 , \5147_b0 );
buf ( \5149_b1 , \5148_b1 );
not ( \5149_b1 , w_16296 );
not ( \5149_b0 , w_16297 );
and ( w_16296 , w_16297 , \5148_b0 );
or ( \5150_b1 , \5136_b1 , w_16298 );
or ( \5150_b0 , \5136_b0 , \5149_b0 );
not ( \5149_b0 , w_16299 );
and ( w_16299 , w_16298 , \5149_b1 );
or ( \5151_b1 , \5148_b1 , w_16300 );
or ( \5151_b0 , \5148_b0 , \5135_b0 );
not ( \5135_b0 , w_16301 );
and ( w_16301 , w_16300 , \5135_b1 );
buf ( \5152_b1 , \4093_b1 );
not ( \5152_b1 , w_16302 );
not ( \5152_b0 , w_16303 );
and ( w_16302 , w_16303 , \4093_b0 );
buf ( \5153_b1 , \4493_b1 );
not ( \5153_b1 , w_16304 );
not ( \5153_b0 , w_16305 );
and ( w_16304 , w_16305 , \4493_b0 );
or ( \5154_b1 , \5152_b1 , w_16306 );
or ( \5154_b0 , \5152_b0 , \5153_b0 );
not ( \5153_b0 , w_16307 );
and ( w_16307 , w_16306 , \5153_b1 );
or ( \5155_b1 , \4285_b1 , w_16309 );
not ( w_16309 , w_16310 );
and ( \5155_b0 , \4285_b0 , w_16311 );
and ( w_16310 ,  , w_16311 );
buf ( w_16309 , \4349_b1 );
not ( w_16309 , w_16312 );
not (  , w_16313 );
and ( w_16312 , w_16313 , \4349_b0 );
or ( \5156_b1 , \5154_b1 , w_16315 );
not ( w_16315 , w_16316 );
and ( \5156_b0 , \5154_b0 , w_16317 );
and ( w_16316 ,  , w_16317 );
buf ( w_16315 , \5155_b1 );
not ( w_16315 , w_16318 );
not (  , w_16319 );
and ( w_16318 , w_16319 , \5155_b0 );
buf ( \5157_b1 , \5156_b1 );
not ( \5157_b1 , w_16320 );
not ( \5157_b0 , w_16321 );
and ( w_16320 , w_16321 , \5156_b0 );
buf ( \5158_b1 , \4430_b1 );
not ( \5158_b1 , w_16322 );
not ( \5158_b0 , w_16323 );
and ( w_16322 , w_16323 , \4430_b0 );
or ( \5159_b1 , \5157_b1 , w_16324 );
or ( \5159_b0 , \5157_b0 , \5158_b0 );
not ( \5158_b0 , w_16325 );
and ( w_16325 , w_16324 , \5158_b1 );
buf ( \5160_b1 , \4800_b1 );
buf ( \5160_b0 , \4800_b0 );
or ( \5161_b1 , \4891_b1 , w_16327 );
not ( w_16327 , w_16328 );
and ( \5161_b0 , \4891_b0 , w_16329 );
and ( w_16328 ,  , w_16329 );
buf ( w_16327 , \5160_b1 );
not ( w_16327 , w_16330 );
not (  , w_16331 );
and ( w_16330 , w_16331 , \5160_b0 );
or ( \5162_b1 , \5159_b1 , w_16333 );
not ( w_16333 , w_16334 );
and ( \5162_b0 , \5159_b0 , w_16335 );
and ( w_16334 ,  , w_16335 );
buf ( w_16333 , \5161_b1 );
not ( w_16333 , w_16336 );
not (  , w_16337 );
and ( w_16336 , w_16337 , \5161_b0 );
or ( \5163_b1 , \5151_b1 , w_16339 );
not ( w_16339 , w_16340 );
and ( \5163_b0 , \5151_b0 , w_16341 );
and ( w_16340 ,  , w_16341 );
buf ( w_16339 , \5162_b1 );
not ( w_16339 , w_16342 );
not (  , w_16343 );
and ( w_16342 , w_16343 , \5162_b0 );
or ( \5164_b1 , \5150_b1 , w_16345 );
not ( w_16345 , w_16346 );
and ( \5164_b0 , \5150_b0 , w_16347 );
and ( w_16346 ,  , w_16347 );
buf ( w_16345 , \5163_b1 );
not ( w_16345 , w_16348 );
not (  , w_16349 );
and ( w_16348 , w_16349 , \5163_b0 );
buf ( \5165_b1 , \5164_b1 );
not ( \5165_b1 , w_16350 );
not ( \5165_b0 , w_16351 );
and ( w_16350 , w_16351 , \5164_b0 );
buf ( \5166_b1 , \5165_b1 );
not ( \5166_b1 , w_16352 );
not ( \5166_b0 , w_16353 );
and ( w_16352 , w_16353 , \5165_b0 );
or ( \5167_b1 , \4870_b1 , \4883_b1 );
xor ( \5167_b0 , \4870_b0 , w_16354 );
not ( w_16354 , w_16355 );
and ( w_16355 , \4883_b1 , \4883_b0 );
or ( \5168_b1 , \5167_b1 , \4896_b1 );
xor ( \5168_b0 , \5167_b0 , w_16356 );
not ( w_16356 , w_16357 );
and ( w_16357 , \4896_b1 , \4896_b0 );
buf ( \5169_b1 , \5168_b1 );
not ( \5169_b1 , w_16358 );
not ( \5169_b0 , w_16359 );
and ( w_16358 , w_16359 , \5168_b0 );
or ( \5170_b1 , \5166_b1 , w_16360 );
or ( \5170_b0 , \5166_b0 , \5169_b0 );
not ( \5169_b0 , w_16361 );
and ( w_16361 , w_16360 , \5169_b1 );
buf ( \5171_b1 , \4066_b1 );
not ( \5171_b1 , w_16362 );
not ( \5171_b0 , w_16363 );
and ( w_16362 , w_16363 , \4066_b0 );
buf ( \5172_b1 , \4163_b1 );
not ( \5172_b1 , w_16364 );
not ( \5172_b0 , w_16365 );
and ( w_16364 , w_16365 , \4163_b0 );
or ( \5173_b1 , \5171_b1 , w_16366 );
or ( \5173_b0 , \5171_b0 , \5172_b0 );
not ( \5172_b0 , w_16367 );
and ( w_16367 , w_16366 , \5172_b1 );
or ( \5174_b1 , \4311_b1 , w_16369 );
not ( w_16369 , w_16370 );
and ( \5174_b0 , \4311_b0 , w_16371 );
and ( w_16370 ,  , w_16371 );
buf ( w_16369 , \4519_b1 );
not ( w_16369 , w_16372 );
not (  , w_16373 );
and ( w_16372 , w_16373 , \4519_b0 );
or ( \5175_b1 , \5173_b1 , w_16375 );
not ( w_16375 , w_16376 );
and ( \5175_b0 , \5173_b0 , w_16377 );
and ( w_16376 ,  , w_16377 );
buf ( w_16375 , \5174_b1 );
not ( w_16375 , w_16378 );
not (  , w_16379 );
and ( w_16378 , w_16379 , \5174_b0 );
buf ( \5176_b1 , \5175_b1 );
not ( \5176_b1 , w_16380 );
not ( \5176_b0 , w_16381 );
and ( w_16380 , w_16381 , \5175_b0 );
buf ( \5177_b1 , \4159_b1 );
not ( \5177_b1 , w_16382 );
not ( \5177_b0 , w_16383 );
and ( w_16382 , w_16383 , \4159_b0 );
or ( \5178_b1 , \5176_b1 , w_16384 );
or ( \5178_b0 , \5176_b0 , \5177_b0 );
not ( \5177_b0 , w_16385 );
and ( w_16385 , w_16384 , \5177_b1 );
or ( \5179_b1 , \4150_b1 , w_16387 );
not ( w_16387 , w_16388 );
and ( \5179_b0 , \4150_b0 , w_16389 );
and ( w_16388 ,  , w_16389 );
buf ( w_16387 , \4908_b1 );
not ( w_16387 , w_16390 );
not (  , w_16391 );
and ( w_16390 , w_16391 , \4908_b0 );
or ( \5180_b1 , \5178_b1 , w_16393 );
not ( w_16393 , w_16394 );
and ( \5180_b0 , \5178_b0 , w_16395 );
and ( w_16394 ,  , w_16395 );
buf ( w_16393 , \5179_b1 );
not ( w_16393 , w_16396 );
not (  , w_16397 );
and ( w_16396 , w_16397 , \5179_b0 );
buf ( \5181_b1 , \5180_b1 );
not ( \5181_b1 , w_16398 );
not ( \5181_b0 , w_16399 );
and ( w_16398 , w_16399 , \5180_b0 );
buf ( \5182_b1 , \4021_b1 );
not ( \5182_b1 , w_16400 );
not ( \5182_b0 , w_16401 );
and ( w_16400 , w_16401 , \4021_b0 );
buf ( \5183_b1 , \4110_b1 );
not ( \5183_b1 , w_16402 );
not ( \5183_b0 , w_16403 );
and ( w_16402 , w_16403 , \4110_b0 );
buf ( \5184_b1 , \5183_b1 );
not ( \5184_b1 , w_16404 );
not ( \5184_b0 , w_16405 );
and ( w_16404 , w_16405 , \5183_b0 );
or ( \5185_b1 , \5182_b1 , w_16406 );
or ( \5185_b0 , \5182_b0 , \5184_b0 );
not ( \5184_b0 , w_16407 );
and ( w_16407 , w_16406 , \5184_b1 );
or ( \5186_b1 , \4106_b1 , w_16409 );
not ( w_16409 , w_16410 );
and ( \5186_b0 , \4106_b0 , w_16411 );
and ( w_16410 ,  , w_16411 );
buf ( w_16409 , \4780_b1 );
not ( w_16409 , w_16412 );
not (  , w_16413 );
and ( w_16412 , w_16413 , \4780_b0 );
or ( \5187_b1 , \5185_b1 , w_16415 );
not ( w_16415 , w_16416 );
and ( \5187_b0 , \5185_b0 , w_16417 );
and ( w_16416 ,  , w_16417 );
buf ( w_16415 , \5186_b1 );
not ( w_16415 , w_16418 );
not (  , w_16419 );
and ( w_16418 , w_16419 , \5186_b0 );
buf ( \5188_b1 , \5187_b1 );
not ( \5188_b1 , w_16420 );
not ( \5188_b0 , w_16421 );
and ( w_16420 , w_16421 , \5187_b0 );
buf ( \5189_b1 , \4710_b1 );
not ( \5189_b1 , w_16422 );
not ( \5189_b0 , w_16423 );
and ( w_16422 , w_16423 , \4710_b0 );
or ( \5190_b1 , \5188_b1 , w_16424 );
or ( \5190_b0 , \5188_b0 , \5189_b0 );
not ( \5189_b0 , w_16425 );
and ( w_16425 , w_16424 , \5189_b1 );
or ( \5191_b1 , \4957_b1 , w_16427 );
not ( w_16427 , w_16428 );
and ( \5191_b0 , \4957_b0 , w_16429 );
and ( w_16428 ,  , w_16429 );
buf ( w_16427 , \4132_b1 );
not ( w_16427 , w_16430 );
not (  , w_16431 );
and ( w_16430 , w_16431 , \4132_b0 );
or ( \5192_b1 , \5190_b1 , w_16433 );
not ( w_16433 , w_16434 );
and ( \5192_b0 , \5190_b0 , w_16435 );
and ( w_16434 ,  , w_16435 );
buf ( w_16433 , \5191_b1 );
not ( w_16433 , w_16436 );
not (  , w_16437 );
and ( w_16436 , w_16437 , \5191_b0 );
buf ( \5193_b1 , \5192_b1 );
not ( \5193_b1 , w_16438 );
not ( \5193_b0 , w_16439 );
and ( w_16438 , w_16439 , \5192_b0 );
or ( \5194_b1 , \5181_b1 , w_16440 );
or ( \5194_b0 , \5181_b0 , \5193_b0 );
not ( \5193_b0 , w_16441 );
and ( w_16441 , w_16440 , \5193_b1 );
or ( \5195_b1 , \5192_b1 , w_16442 );
or ( \5195_b0 , \5192_b0 , \5180_b0 );
not ( \5180_b0 , w_16443 );
and ( w_16443 , w_16442 , \5180_b1 );
buf ( \5196_b1 , \5122_b1 );
not ( \5196_b1 , w_16444 );
not ( \5196_b0 , w_16445 );
and ( w_16444 , w_16445 , \5122_b0 );
buf ( \5197_b1 , \4632_b1 );
not ( \5197_b1 , w_16446 );
not ( \5197_b0 , w_16447 );
and ( w_16446 , w_16447 , \4632_b0 );
or ( \5198_b1 , \5196_b1 , w_16448 );
or ( \5198_b0 , \5196_b0 , \5197_b0 );
not ( \5197_b0 , w_16449 );
and ( w_16449 , w_16448 , \5197_b1 );
or ( \5199_b1 , \4453_b1 , w_16451 );
not ( w_16451 , w_16452 );
and ( \5199_b0 , \4453_b0 , w_16453 );
and ( w_16452 ,  , w_16453 );
buf ( w_16451 , \4921_b1 );
not ( w_16451 , w_16454 );
not (  , w_16455 );
and ( w_16454 , w_16455 , \4921_b0 );
or ( \5200_b1 , \5198_b1 , w_16457 );
not ( w_16457 , w_16458 );
and ( \5200_b0 , \5198_b0 , w_16459 );
and ( w_16458 ,  , w_16459 );
buf ( w_16457 , \5199_b1 );
not ( w_16457 , w_16460 );
not (  , w_16461 );
and ( w_16460 , w_16461 , \5199_b0 );
or ( \5201_b1 , \5195_b1 , w_16463 );
not ( w_16463 , w_16464 );
and ( \5201_b0 , \5195_b0 , w_16465 );
and ( w_16464 ,  , w_16465 );
buf ( w_16463 , \5200_b1 );
not ( w_16463 , w_16466 );
not (  , w_16467 );
and ( w_16466 , w_16467 , \5200_b0 );
or ( \5202_b1 , \5194_b1 , w_16469 );
not ( w_16469 , w_16470 );
and ( \5202_b0 , \5194_b0 , w_16471 );
and ( w_16470 ,  , w_16471 );
buf ( w_16469 , \5201_b1 );
not ( w_16469 , w_16472 );
not (  , w_16473 );
and ( w_16472 , w_16473 , \5201_b0 );
or ( \5203_b1 , \5170_b1 , w_16475 );
not ( w_16475 , w_16476 );
and ( \5203_b0 , \5170_b0 , w_16477 );
and ( w_16476 ,  , w_16477 );
buf ( w_16475 , \5202_b1 );
not ( w_16475 , w_16478 );
not (  , w_16479 );
and ( w_16478 , w_16479 , \5202_b0 );
buf ( \5204_b1 , \5165_b1 );
not ( \5204_b1 , w_16480 );
not ( \5204_b0 , w_16481 );
and ( w_16480 , w_16481 , \5165_b0 );
buf ( \5205_b1 , \5168_b1 );
not ( \5205_b1 , w_16482 );
not ( \5205_b0 , w_16483 );
and ( w_16482 , w_16483 , \5168_b0 );
or ( \5206_b1 , \5204_b1 , w_16485 );
not ( w_16485 , w_16486 );
and ( \5206_b0 , \5204_b0 , w_16487 );
and ( w_16486 ,  , w_16487 );
buf ( w_16485 , \5205_b1 );
not ( w_16485 , w_16488 );
not (  , w_16489 );
and ( w_16488 , w_16489 , \5205_b0 );
or ( \5207_b1 , \5203_b1 , \5206_b1 );
not ( \5206_b1 , w_16490 );
and ( \5207_b0 , \5203_b0 , w_16491 );
and ( w_16490 , w_16491 , \5206_b0 );
or ( \5208_b1 , \5132_b1 , \5207_b1 );
xor ( \5208_b0 , \5132_b0 , w_16492 );
not ( w_16492 , w_16493 );
and ( w_16493 , \5207_b1 , \5207_b0 );
buf ( \5209_b1 , \4982_b1 );
not ( \5209_b1 , w_16494 );
not ( \5209_b0 , w_16495 );
and ( w_16494 , w_16495 , \4982_b0 );
buf ( \5210_b1 , \4978_b1 );
not ( \5210_b1 , w_16496 );
not ( \5210_b0 , w_16497 );
and ( w_16496 , w_16497 , \4978_b0 );
or ( \5211_b1 , \5209_b1 , w_16498 );
or ( \5211_b0 , \5209_b0 , \5210_b0 );
not ( \5210_b0 , w_16499 );
and ( w_16499 , w_16498 , \5210_b1 );
or ( \5212_b1 , \4978_b1 , w_16500 );
or ( \5212_b0 , \4978_b0 , \4982_b0 );
not ( \4982_b0 , w_16501 );
and ( w_16501 , w_16500 , \4982_b1 );
or ( \5213_b1 , \5211_b1 , w_16503 );
not ( w_16503 , w_16504 );
and ( \5213_b0 , \5211_b0 , w_16505 );
and ( w_16504 ,  , w_16505 );
buf ( w_16503 , \5212_b1 );
not ( w_16503 , w_16506 );
not (  , w_16507 );
and ( w_16506 , w_16507 , \5212_b0 );
buf ( \5214_b1 , \4996_b1 );
not ( \5214_b1 , w_16508 );
not ( \5214_b0 , w_16509 );
and ( w_16508 , w_16509 , \4996_b0 );
or ( \5215_b1 , \5213_b1 , \5214_b1 );
not ( \5214_b1 , w_16510 );
and ( \5215_b0 , \5213_b0 , w_16511 );
and ( w_16510 , w_16511 , \5214_b0 );
buf ( \5216_b1 , \5213_b1 );
not ( \5216_b1 , w_16512 );
not ( \5216_b0 , w_16513 );
and ( w_16512 , w_16513 , \5213_b0 );
or ( \5217_b1 , \5216_b1 , \4996_b1 );
not ( \4996_b1 , w_16514 );
and ( \5217_b0 , \5216_b0 , w_16515 );
and ( w_16514 , w_16515 , \4996_b0 );
or ( \5218_b1 , \5215_b1 , w_16517 );
not ( w_16517 , w_16518 );
and ( \5218_b0 , \5215_b0 , w_16519 );
and ( w_16518 ,  , w_16519 );
buf ( w_16517 , \5217_b1 );
not ( w_16517 , w_16520 );
not (  , w_16521 );
and ( w_16520 , w_16521 , \5217_b0 );
or ( \5219_b1 , \5208_b1 , \5218_b1 );
xor ( \5219_b0 , \5208_b0 , w_16522 );
not ( w_16522 , w_16523 );
and ( w_16523 , \5218_b1 , \5218_b0 );
or ( \5220_b1 , \5130_b1 , \5219_b1 );
xor ( \5220_b0 , \5130_b0 , w_16524 );
not ( w_16524 , w_16525 );
and ( w_16525 , \5219_b1 , \5219_b0 );
buf ( \5221_b1 , \4951_b1 );
not ( \5221_b1 , w_16526 );
not ( \5221_b0 , w_16527 );
and ( w_16526 , w_16527 , \4951_b0 );
buf ( \5222_b1 , \5221_b1 );
not ( \5222_b1 , w_16528 );
not ( \5222_b0 , w_16529 );
and ( w_16528 , w_16529 , \5221_b0 );
buf ( \5223_b1 , \5100_b1 );
not ( \5223_b1 , w_16530 );
not ( \5223_b0 , w_16531 );
and ( w_16530 , w_16531 , \5100_b0 );
or ( \5224_b1 , \5222_b1 , w_16532 );
or ( \5224_b0 , \5222_b0 , \5223_b0 );
not ( \5223_b0 , w_16533 );
and ( w_16533 , w_16532 , \5223_b1 );
or ( \5225_b1 , \5100_b1 , w_16534 );
or ( \5225_b0 , \5100_b0 , \5221_b0 );
not ( \5221_b0 , w_16535 );
and ( w_16535 , w_16534 , \5221_b1 );
or ( \5226_b1 , \5224_b1 , w_16537 );
not ( w_16537 , w_16538 );
and ( \5226_b0 , \5224_b0 , w_16539 );
and ( w_16538 ,  , w_16539 );
buf ( w_16537 , \5225_b1 );
not ( w_16537 , w_16540 );
not (  , w_16541 );
and ( w_16540 , w_16541 , \5225_b0 );
buf ( \5227_b1 , \5125_b1 );
not ( \5227_b1 , w_16542 );
not ( \5227_b0 , w_16543 );
and ( w_16542 , w_16543 , \5125_b0 );
or ( \5228_b1 , \5226_b1 , \5227_b1 );
not ( \5227_b1 , w_16544 );
and ( \5228_b0 , \5226_b0 , w_16545 );
and ( w_16544 , w_16545 , \5227_b0 );
buf ( \5229_b1 , \5226_b1 );
not ( \5229_b1 , w_16546 );
not ( \5229_b0 , w_16547 );
and ( w_16546 , w_16547 , \5226_b0 );
or ( \5230_b1 , \5229_b1 , \5125_b1 );
not ( \5125_b1 , w_16548 );
and ( \5230_b0 , \5229_b0 , w_16549 );
and ( w_16548 , w_16549 , \5125_b0 );
or ( \5231_b1 , \5228_b1 , w_16551 );
not ( w_16551 , w_16552 );
and ( \5231_b0 , \5228_b0 , w_16553 );
and ( w_16552 ,  , w_16553 );
buf ( w_16551 , \5230_b1 );
not ( w_16551 , w_16554 );
not (  , w_16555 );
and ( w_16554 , w_16555 , \5230_b0 );
buf ( \5232_b1 , \5231_b1 );
not ( \5232_b1 , w_16556 );
not ( \5232_b0 , w_16557 );
and ( w_16556 , w_16557 , \5231_b0 );
buf ( \5233_b1 , \5232_b1 );
not ( \5233_b1 , w_16558 );
not ( \5233_b0 , w_16559 );
and ( w_16558 , w_16559 , \5232_b0 );
buf ( \5234_b1 , \5162_b1 );
buf ( \5234_b0 , \5162_b0 );
or ( \5235_b1 , \5148_b1 , \5135_b1 );
not ( \5135_b1 , w_16560 );
and ( \5235_b0 , \5148_b0 , w_16561 );
and ( w_16560 , w_16561 , \5135_b0 );
buf ( \5236_b1 , \5148_b1 );
not ( \5236_b1 , w_16562 );
not ( \5236_b0 , w_16563 );
and ( w_16562 , w_16563 , \5148_b0 );
or ( \5237_b1 , \5236_b1 , \5134_b1 );
not ( \5134_b1 , w_16564 );
and ( \5237_b0 , \5236_b0 , w_16565 );
and ( w_16564 , w_16565 , \5134_b0 );
or ( \5238_b1 , \5235_b1 , w_16567 );
not ( w_16567 , w_16568 );
and ( \5238_b0 , \5235_b0 , w_16569 );
and ( w_16568 ,  , w_16569 );
buf ( w_16567 , \5237_b1 );
not ( w_16567 , w_16570 );
not (  , w_16571 );
and ( w_16570 , w_16571 , \5237_b0 );
or ( \5239_b1 , \5234_b1 , \5238_b1 );
xor ( \5239_b0 , \5234_b0 , w_16572 );
not ( w_16572 , w_16573 );
and ( w_16573 , \5238_b1 , \5238_b0 );
buf ( \5240_b1 , \5239_b1 );
not ( \5240_b1 , w_16574 );
not ( \5240_b0 , w_16575 );
and ( w_16574 , w_16575 , \5239_b0 );
or ( \5241_b1 , \5233_b1 , w_16576 );
or ( \5241_b0 , \5233_b0 , \5240_b0 );
not ( \5240_b0 , w_16577 );
and ( w_16577 , w_16576 , \5240_b1 );
buf ( \5242_b1 , \5231_b1 );
not ( \5242_b1 , w_16578 );
not ( \5242_b0 , w_16579 );
and ( w_16578 , w_16579 , \5231_b0 );
buf ( \5243_b1 , \5239_b1 );
not ( \5243_b1 , w_16580 );
not ( \5243_b0 , w_16581 );
and ( w_16580 , w_16581 , \5239_b0 );
buf ( \5244_b1 , \5243_b1 );
not ( \5244_b1 , w_16582 );
not ( \5244_b0 , w_16583 );
and ( w_16582 , w_16583 , \5243_b0 );
or ( \5245_b1 , \5242_b1 , w_16584 );
or ( \5245_b0 , \5242_b0 , \5244_b0 );
not ( \5244_b0 , w_16585 );
and ( w_16585 , w_16584 , \5244_b1 );
or ( \5246_b1 , \5124_b1 , w_16587 );
not ( w_16587 , w_16588 );
and ( \5246_b0 , \5124_b0 , w_16589 );
and ( w_16588 ,  , w_16589 );
buf ( w_16587 , \5110_b1 );
not ( w_16587 , w_16590 );
not (  , w_16591 );
and ( w_16590 , w_16591 , \5110_b0 );
buf ( \5247_b1 , \5246_b1 );
not ( \5247_b1 , w_16592 );
not ( \5247_b0 , w_16593 );
and ( w_16592 , w_16593 , \5246_b0 );
or ( \5248_b1 , \5247_b1 , w_16595 );
not ( w_16595 , w_16596 );
and ( \5248_b0 , \5247_b0 , w_16597 );
and ( w_16596 ,  , w_16597 );
buf ( w_16595 , \5125_b1 );
not ( w_16595 , w_16598 );
not (  , w_16599 );
and ( w_16598 , w_16599 , \5125_b0 );
buf ( \5249_b1 , \4026_b1 );
not ( \5249_b1 , w_16600 );
not ( \5249_b0 , w_16601 );
and ( w_16600 , w_16601 , \4026_b0 );
buf ( \5250_b1 , \5183_b1 );
not ( \5250_b1 , w_16602 );
not ( \5250_b0 , w_16603 );
and ( w_16602 , w_16603 , \5183_b0 );
or ( \5251_b1 , \5249_b1 , w_16604 );
or ( \5251_b0 , \5249_b0 , \5250_b0 );
not ( \5250_b0 , w_16605 );
and ( w_16605 , w_16604 , \5250_b1 );
or ( \5252_b1 , \4106_b1 , w_16607 );
not ( w_16607 , w_16608 );
and ( \5252_b0 , \4106_b0 , w_16609 );
and ( w_16608 ,  , w_16609 );
buf ( w_16607 , \4969_b1 );
not ( w_16607 , w_16610 );
not (  , w_16611 );
and ( w_16610 , w_16611 , \4969_b0 );
or ( \5253_b1 , \5251_b1 , w_16613 );
not ( w_16613 , w_16614 );
and ( \5253_b0 , \5251_b0 , w_16615 );
and ( w_16614 ,  , w_16615 );
buf ( w_16613 , \5252_b1 );
not ( w_16613 , w_16616 );
not (  , w_16617 );
and ( w_16616 , w_16617 , \5252_b0 );
buf ( \5254_b1 , \5253_b1 );
not ( \5254_b1 , w_16618 );
not ( \5254_b0 , w_16619 );
and ( w_16618 , w_16619 , \5253_b0 );
buf ( \5255_b1 , \4129_b1 );
not ( \5255_b1 , w_16620 );
not ( \5255_b0 , w_16621 );
and ( w_16620 , w_16621 , \4129_b0 );
or ( \5256_b1 , \5254_b1 , w_16622 );
or ( \5256_b0 , \5254_b0 , \5255_b0 );
not ( \5255_b0 , w_16623 );
and ( w_16623 , w_16622 , \5255_b1 );
or ( \5257_b1 , \4133_b1 , w_16625 );
not ( w_16625 , w_16626 );
and ( \5257_b0 , \4133_b0 , w_16627 );
and ( w_16626 ,  , w_16627 );
buf ( w_16625 , \5187_b1 );
not ( w_16625 , w_16628 );
not (  , w_16629 );
and ( w_16628 , w_16629 , \5187_b0 );
or ( \5258_b1 , \5256_b1 , w_16631 );
not ( w_16631 , w_16632 );
and ( \5258_b0 , \5256_b0 , w_16633 );
and ( w_16632 ,  , w_16633 );
buf ( w_16631 , \5257_b1 );
not ( w_16631 , w_16634 );
not (  , w_16635 );
and ( w_16634 , w_16635 , \5257_b0 );
or ( \5259_b1 , \5248_b1 , \5258_b1 );
not ( \5258_b1 , w_16636 );
and ( \5259_b0 , \5248_b0 , w_16637 );
and ( w_16636 , w_16637 , \5258_b0 );
or ( \5260_b1 , \5245_b1 , w_16639 );
not ( w_16639 , w_16640 );
and ( \5260_b0 , \5245_b0 , w_16641 );
and ( w_16640 ,  , w_16641 );
buf ( w_16639 , \5259_b1 );
not ( w_16639 , w_16642 );
not (  , w_16643 );
and ( w_16642 , w_16643 , \5259_b0 );
or ( \5261_b1 , \5241_b1 , w_16645 );
not ( w_16645 , w_16646 );
and ( \5261_b0 , \5241_b0 , w_16647 );
and ( w_16646 ,  , w_16647 );
buf ( w_16645 , \5260_b1 );
not ( w_16645 , w_16648 );
not (  , w_16649 );
and ( w_16648 , w_16649 , \5260_b0 );
buf ( \5262_b1 , \5261_b1 );
not ( \5262_b1 , w_16650 );
not ( \5262_b0 , w_16651 );
and ( w_16650 , w_16651 , \5261_b0 );
or ( \5263_b1 , \5164_b1 , \5202_b1 );
xor ( \5263_b0 , \5164_b0 , w_16652 );
not ( w_16652 , w_16653 );
and ( w_16653 , \5202_b1 , \5202_b0 );
or ( \5264_b1 , \5263_b1 , w_16654 );
xor ( \5264_b0 , \5263_b0 , w_16656 );
not ( w_16656 , w_16657 );
and ( w_16657 , w_16654 , w_16655 );
buf ( w_16654 , \5205_b1 );
not ( w_16654 , w_16658 );
not ( w_16655 , w_16659 );
and ( w_16658 , w_16659 , \5205_b0 );
or ( \5265_b1 , \5262_b1 , w_16661 );
not ( w_16661 , w_16662 );
and ( \5265_b0 , \5262_b0 , w_16663 );
and ( w_16662 ,  , w_16663 );
buf ( w_16661 , \5264_b1 );
not ( w_16661 , w_16664 );
not (  , w_16665 );
and ( w_16664 , w_16665 , \5264_b0 );
buf ( \5266_b1 , \3241_b1 );
buf ( \5266_b0 , \3241_b0 );
buf ( \5267_b1 , \5266_b1 );
not ( \5267_b1 , w_16666 );
not ( \5267_b0 , w_16667 );
and ( w_16666 , w_16667 , \5266_b0 );
buf ( \5268_b1 , \3070_b1 );
buf ( \5268_b0 , \3070_b0 );
buf ( \5269_b1 , \5268_b1 );
not ( \5269_b1 , w_16668 );
not ( \5269_b0 , w_16669 );
and ( w_16668 , w_16669 , \5268_b0 );
or ( \5270_b1 , \5269_b1 , w_16671 );
not ( w_16671 , w_16672 );
and ( \5270_b0 , \5269_b0 , w_16673 );
and ( w_16672 ,  , w_16673 );
buf ( w_16671 , \3241_b1 );
not ( w_16671 , w_16674 );
not (  , w_16675 );
and ( w_16674 , w_16675 , \3241_b0 );
buf ( \5271_b1 , \5270_b1 );
buf ( \5271_b0 , \5270_b0 );
buf ( \5272_b1 , \5271_b1 );
not ( \5272_b1 , w_16676 );
not ( \5272_b0 , w_16677 );
and ( w_16676 , w_16677 , \5271_b0 );
or ( \5273_b1 , \5267_b1 , w_16679 );
not ( w_16679 , w_16680 );
and ( \5273_b0 , \5267_b0 , w_16681 );
and ( w_16680 ,  , w_16681 );
buf ( w_16679 , \5272_b1 );
not ( w_16679 , w_16682 );
not (  , w_16683 );
and ( w_16682 , w_16683 , \5272_b0 );
buf ( \5274_b1 , \5268_b1 );
not ( \5274_b1 , w_16684 );
not ( \5274_b0 , w_16685 );
and ( w_16684 , w_16685 , \5268_b0 );
buf ( \5275_b1 , \5274_b1 );
not ( \5275_b1 , w_16686 );
not ( \5275_b0 , w_16687 );
and ( w_16686 , w_16687 , \5274_b0 );
or ( \5276_b1 , \5273_b1 , w_16689 );
not ( w_16689 , w_16690 );
and ( \5276_b0 , \5273_b0 , w_16691 );
and ( w_16690 ,  , w_16691 );
buf ( w_16689 , \5275_b1 );
not ( w_16689 , w_16692 );
not (  , w_16693 );
and ( w_16692 , w_16693 , \5275_b0 );
buf ( \5277_b1 , \5276_b1 );
not ( \5277_b1 , w_16694 );
not ( \5277_b0 , w_16695 );
and ( w_16694 , w_16695 , \5276_b0 );
or ( \5278_b1 , \4253_b1 , w_16697 );
not ( w_16697 , w_16698 );
and ( \5278_b0 , \4253_b0 , w_16699 );
and ( w_16698 ,  , w_16699 );
buf ( w_16697 , \4079_b1 );
not ( w_16697 , w_16700 );
not (  , w_16701 );
and ( w_16700 , w_16701 , \4079_b0 );
or ( \5279_b1 , \5277_b1 , w_16703 );
not ( w_16703 , w_16704 );
and ( \5279_b0 , \5277_b0 , w_16705 );
and ( w_16704 ,  , w_16705 );
buf ( w_16703 , \5278_b1 );
not ( w_16703 , w_16706 );
not (  , w_16707 );
and ( w_16706 , w_16707 , \5278_b0 );
buf ( \5280_b1 , \5279_b1 );
not ( \5280_b1 , w_16708 );
not ( \5280_b0 , w_16709 );
and ( w_16708 , w_16709 , \5279_b0 );
buf ( \5281_b1 , \4076_b1 );
not ( \5281_b1 , w_16710 );
not ( \5281_b0 , w_16711 );
and ( w_16710 , w_16711 , \4076_b0 );
buf ( \5282_b1 , \4250_b1 );
not ( \5282_b1 , w_16712 );
not ( \5282_b0 , w_16713 );
and ( w_16712 , w_16713 , \4250_b0 );
or ( \5283_b1 , \5281_b1 , w_16714 );
or ( \5283_b0 , \5281_b0 , \5282_b0 );
not ( \5282_b0 , w_16715 );
and ( w_16715 , w_16714 , \5282_b1 );
buf ( \5284_b1 , \4076_b1 );
not ( \5284_b1 , w_16716 );
not ( \5284_b0 , w_16717 );
and ( w_16716 , w_16717 , \4076_b0 );
or ( \5285_b1 , \5133_b1 , w_16719 );
not ( w_16719 , w_16720 );
and ( \5285_b0 , \5133_b0 , w_16721 );
and ( w_16720 ,  , w_16721 );
buf ( w_16719 , \5284_b1 );
not ( w_16719 , w_16722 );
not (  , w_16723 );
and ( w_16722 , w_16723 , \5284_b0 );
or ( \5286_b1 , \5283_b1 , w_16725 );
not ( w_16725 , w_16726 );
and ( \5286_b0 , \5283_b0 , w_16727 );
and ( w_16726 ,  , w_16727 );
buf ( w_16725 , \5285_b1 );
not ( w_16725 , w_16728 );
not (  , w_16729 );
and ( w_16728 , w_16729 , \5285_b0 );
buf ( \5287_b1 , \5286_b1 );
not ( \5287_b1 , w_16730 );
not ( \5287_b0 , w_16731 );
and ( w_16730 , w_16731 , \5286_b0 );
buf ( \5288_b1 , \4395_b1 );
not ( \5288_b1 , w_16732 );
not ( \5288_b0 , w_16733 );
and ( w_16732 , w_16733 , \4395_b0 );
or ( \5289_b1 , \5287_b1 , w_16734 );
or ( \5289_b0 , \5287_b0 , \5288_b0 );
not ( \5288_b0 , w_16735 );
and ( w_16735 , w_16734 , \5288_b1 );
or ( \5290_b1 , \5091_b1 , w_16737 );
not ( w_16737 , w_16738 );
and ( \5290_b0 , \5091_b0 , w_16739 );
and ( w_16738 ,  , w_16739 );
buf ( w_16737 , \4200_b1 );
not ( w_16737 , w_16740 );
not (  , w_16741 );
and ( w_16740 , w_16741 , \4200_b0 );
or ( \5291_b1 , \5289_b1 , w_16743 );
not ( w_16743 , w_16744 );
and ( \5291_b0 , \5289_b0 , w_16745 );
and ( w_16744 ,  , w_16745 );
buf ( w_16743 , \5290_b1 );
not ( w_16743 , w_16746 );
not (  , w_16747 );
and ( w_16746 , w_16747 , \5290_b0 );
buf ( \5292_b1 , \5291_b1 );
not ( \5292_b1 , w_16748 );
not ( \5292_b0 , w_16749 );
and ( w_16748 , w_16749 , \5291_b0 );
or ( \5293_b1 , \5280_b1 , w_16750 );
or ( \5293_b0 , \5280_b0 , \5292_b0 );
not ( \5292_b0 , w_16751 );
and ( w_16751 , w_16750 , \5292_b1 );
buf ( \5294_b1 , \5278_b1 );
not ( \5294_b1 , w_16752 );
not ( \5294_b0 , w_16753 );
and ( w_16752 , w_16753 , \5278_b0 );
or ( \5295_b1 , \5294_b1 , w_16755 );
not ( w_16755 , w_16756 );
and ( \5295_b0 , \5294_b0 , w_16757 );
and ( w_16756 ,  , w_16757 );
buf ( w_16755 , \5276_b1 );
not ( w_16755 , w_16758 );
not (  , w_16759 );
and ( w_16758 , w_16759 , \5276_b0 );
or ( \5296_b1 , \5293_b1 , w_16761 );
not ( w_16761 , w_16762 );
and ( \5296_b0 , \5293_b0 , w_16763 );
and ( w_16762 ,  , w_16763 );
buf ( w_16761 , \5295_b1 );
not ( w_16761 , w_16764 );
not (  , w_16765 );
and ( w_16764 , w_16765 , \5295_b0 );
buf ( \5297_b1 , \5296_b1 );
not ( \5297_b1 , w_16766 );
not ( \5297_b0 , w_16767 );
and ( w_16766 , w_16767 , \5296_b0 );
buf ( \5298_b1 , \5297_b1 );
not ( \5298_b1 , w_16768 );
not ( \5298_b0 , w_16769 );
and ( w_16768 , w_16769 , \5297_b0 );
buf ( \5299_b1 , \4611_b1 );
not ( \5299_b1 , w_16770 );
not ( \5299_b0 , w_16771 );
and ( w_16770 , w_16771 , \4611_b0 );
buf ( \5300_b1 , \4094_b1 );
not ( \5300_b1 , w_16772 );
not ( \5300_b0 , w_16773 );
and ( w_16772 , w_16773 , \4094_b0 );
buf ( \5301_b1 , \4616_b1 );
not ( \5301_b1 , w_16774 );
not ( \5301_b0 , w_16775 );
and ( w_16774 , w_16775 , \4616_b0 );
buf ( \5302_b1 , \5301_b1 );
not ( \5302_b1 , w_16776 );
not ( \5302_b0 , w_16777 );
and ( w_16776 , w_16777 , \5301_b0 );
or ( \5303_b1 , \5300_b1 , w_16778 );
or ( \5303_b0 , \5300_b0 , \5302_b0 );
not ( \5302_b0 , w_16779 );
and ( w_16779 , w_16778 , \5302_b1 );
or ( \5304_b1 , \4616_b1 , w_16781 );
not ( w_16781 , w_16782 );
and ( \5304_b0 , \4616_b0 , w_16783 );
and ( w_16782 ,  , w_16783 );
buf ( w_16781 , \4298_b1 );
not ( w_16781 , w_16784 );
not (  , w_16785 );
and ( w_16784 , w_16785 , \4298_b0 );
or ( \5305_b1 , \5303_b1 , w_16787 );
not ( w_16787 , w_16788 );
and ( \5305_b0 , \5303_b0 , w_16789 );
and ( w_16788 ,  , w_16789 );
buf ( w_16787 , \5304_b1 );
not ( w_16787 , w_16790 );
not (  , w_16791 );
and ( w_16790 , w_16791 , \5304_b0 );
buf ( \5306_b1 , \5305_b1 );
not ( \5306_b1 , w_16792 );
not ( \5306_b0 , w_16793 );
and ( w_16792 , w_16793 , \5305_b0 );
or ( \5307_b1 , \5299_b1 , w_16794 );
or ( \5307_b0 , \5299_b0 , \5306_b0 );
not ( \5306_b0 , w_16795 );
and ( w_16795 , w_16794 , \5306_b1 );
or ( \5308_b1 , \5142_b1 , w_16797 );
not ( w_16797 , w_16798 );
and ( \5308_b0 , \5142_b0 , w_16799 );
and ( w_16798 ,  , w_16799 );
buf ( w_16797 , \4881_b1 );
not ( w_16797 , w_16800 );
not (  , w_16801 );
and ( w_16800 , w_16801 , \4881_b0 );
or ( \5309_b1 , \5307_b1 , w_16803 );
not ( w_16803 , w_16804 );
and ( \5309_b0 , \5307_b0 , w_16805 );
and ( w_16804 ,  , w_16805 );
buf ( w_16803 , \5308_b1 );
not ( w_16803 , w_16806 );
not (  , w_16807 );
and ( w_16806 , w_16807 , \5308_b0 );
buf ( \5310_b1 , \5309_b1 );
not ( \5310_b1 , w_16808 );
not ( \5310_b0 , w_16809 );
and ( w_16808 , w_16809 , \5309_b0 );
buf ( \5311_b1 , \4017_b1 );
not ( \5311_b1 , w_16810 );
not ( \5311_b0 , w_16811 );
and ( w_16810 , w_16811 , \4017_b0 );
buf ( \5312_b1 , \4163_b1 );
not ( \5312_b1 , w_16812 );
not ( \5312_b0 , w_16813 );
and ( w_16812 , w_16813 , \4163_b0 );
or ( \5313_b1 , \5311_b1 , w_16814 );
or ( \5313_b0 , \5311_b0 , \5312_b0 );
not ( \5312_b0 , w_16815 );
and ( w_16815 , w_16814 , \5312_b1 );
or ( \5314_b1 , \4164_b1 , w_16817 );
not ( w_16817 , w_16818 );
and ( \5314_b0 , \4164_b0 , w_16819 );
and ( w_16818 ,  , w_16819 );
buf ( w_16817 , \4662_b1 );
not ( w_16817 , w_16820 );
not (  , w_16821 );
and ( w_16820 , w_16821 , \4662_b0 );
or ( \5315_b1 , \5313_b1 , w_16823 );
not ( w_16823 , w_16824 );
and ( \5315_b0 , \5313_b0 , w_16825 );
and ( w_16824 ,  , w_16825 );
buf ( w_16823 , \5314_b1 );
not ( w_16823 , w_16826 );
not (  , w_16827 );
and ( w_16826 , w_16827 , \5314_b0 );
buf ( \5316_b1 , \5315_b1 );
not ( \5316_b1 , w_16828 );
not ( \5316_b0 , w_16829 );
and ( w_16828 , w_16829 , \5315_b0 );
buf ( \5317_b1 , \4159_b1 );
not ( \5317_b1 , w_16830 );
not ( \5317_b0 , w_16831 );
and ( w_16830 , w_16831 , \4159_b0 );
or ( \5318_b1 , \5316_b1 , w_16832 );
or ( \5318_b0 , \5316_b0 , \5317_b0 );
not ( \5317_b0 , w_16833 );
and ( w_16833 , w_16832 , \5317_b1 );
or ( \5319_b1 , \4317_b1 , w_16835 );
not ( w_16835 , w_16836 );
and ( \5319_b0 , \4317_b0 , w_16837 );
and ( w_16836 ,  , w_16837 );
buf ( w_16835 , \5175_b1 );
not ( w_16835 , w_16838 );
not (  , w_16839 );
and ( w_16838 , w_16839 , \5175_b0 );
or ( \5320_b1 , \5318_b1 , w_16841 );
not ( w_16841 , w_16842 );
and ( \5320_b0 , \5318_b0 , w_16843 );
and ( w_16842 ,  , w_16843 );
buf ( w_16841 , \5319_b1 );
not ( w_16841 , w_16844 );
not (  , w_16845 );
and ( w_16844 , w_16845 , \5319_b0 );
buf ( \5321_b1 , \5320_b1 );
not ( \5321_b1 , w_16846 );
not ( \5321_b0 , w_16847 );
and ( w_16846 , w_16847 , \5320_b0 );
or ( \5322_b1 , \5310_b1 , w_16848 );
or ( \5322_b0 , \5310_b0 , \5321_b0 );
not ( \5321_b0 , w_16849 );
and ( w_16849 , w_16848 , \5321_b1 );
or ( \5323_b1 , \5309_b1 , w_16850 );
or ( \5323_b0 , \5309_b0 , \5320_b0 );
not ( \5320_b0 , w_16851 );
and ( w_16851 , w_16850 , \5320_b1 );
buf ( \5324_b1 , \4095_b1 );
not ( \5324_b1 , w_16852 );
not ( \5324_b0 , w_16853 );
and ( w_16852 , w_16853 , \4095_b0 );
buf ( \5325_b1 , \4332_b1 );
not ( \5325_b1 , w_16854 );
not ( \5325_b0 , w_16855 );
and ( w_16854 , w_16855 , \4332_b0 );
or ( \5326_b1 , \5324_b1 , w_16856 );
or ( \5326_b0 , \5324_b0 , \5325_b0 );
not ( \5325_b0 , w_16857 );
and ( w_16857 , w_16856 , \5325_b1 );
or ( \5327_b1 , \4283_b1 , w_16859 );
not ( w_16859 , w_16860 );
and ( \5327_b0 , \4283_b0 , w_16861 );
and ( w_16860 ,  , w_16861 );
buf ( w_16859 , \4391_b1 );
not ( w_16859 , w_16862 );
not (  , w_16863 );
and ( w_16862 , w_16863 , \4391_b0 );
or ( \5328_b1 , \5326_b1 , w_16865 );
not ( w_16865 , w_16866 );
and ( \5328_b0 , \5326_b0 , w_16867 );
and ( w_16866 ,  , w_16867 );
buf ( w_16865 , \5327_b1 );
not ( w_16865 , w_16868 );
not (  , w_16869 );
and ( w_16868 , w_16869 , \5327_b0 );
buf ( \5329_b1 , \5328_b1 );
not ( \5329_b1 , w_16870 );
not ( \5329_b0 , w_16871 );
and ( w_16870 , w_16871 , \5328_b0 );
buf ( \5330_b1 , \4430_b1 );
not ( \5330_b1 , w_16872 );
not ( \5330_b0 , w_16873 );
and ( w_16872 , w_16873 , \4430_b0 );
or ( \5331_b1 , \5329_b1 , w_16874 );
or ( \5331_b0 , \5329_b0 , \5330_b0 );
not ( \5330_b0 , w_16875 );
and ( w_16875 , w_16874 , \5330_b1 );
or ( \5332_b1 , \5156_b1 , w_16877 );
not ( w_16877 , w_16878 );
and ( \5332_b0 , \5156_b0 , w_16879 );
and ( w_16878 ,  , w_16879 );
buf ( w_16877 , \4341_b1 );
not ( w_16877 , w_16880 );
not (  , w_16881 );
and ( w_16880 , w_16881 , \4341_b0 );
or ( \5333_b1 , \5331_b1 , w_16883 );
not ( w_16883 , w_16884 );
and ( \5333_b0 , \5331_b0 , w_16885 );
and ( w_16884 ,  , w_16885 );
buf ( w_16883 , \5332_b1 );
not ( w_16883 , w_16886 );
not (  , w_16887 );
and ( w_16886 , w_16887 , \5332_b0 );
or ( \5334_b1 , \5323_b1 , w_16889 );
not ( w_16889 , w_16890 );
and ( \5334_b0 , \5323_b0 , w_16891 );
and ( w_16890 ,  , w_16891 );
buf ( w_16889 , \5333_b1 );
not ( w_16889 , w_16892 );
not (  , w_16893 );
and ( w_16892 , w_16893 , \5333_b0 );
or ( \5335_b1 , \5322_b1 , w_16895 );
not ( w_16895 , w_16896 );
and ( \5335_b0 , \5322_b0 , w_16897 );
and ( w_16896 ,  , w_16897 );
buf ( w_16895 , \5334_b1 );
not ( w_16895 , w_16898 );
not (  , w_16899 );
and ( w_16898 , w_16899 , \5334_b0 );
buf ( \5336_b1 , \5335_b1 );
not ( \5336_b1 , w_16900 );
not ( \5336_b0 , w_16901 );
and ( w_16900 , w_16901 , \5335_b0 );
buf ( \5337_b1 , \5336_b1 );
not ( \5337_b1 , w_16902 );
not ( \5337_b0 , w_16903 );
and ( w_16902 , w_16903 , \5336_b0 );
or ( \5338_b1 , \5298_b1 , w_16904 );
or ( \5338_b0 , \5298_b0 , \5337_b0 );
not ( \5337_b0 , w_16905 );
and ( w_16905 , w_16904 , \5337_b1 );
or ( \5339_b1 , \5192_b1 , \5180_b1 );
xor ( \5339_b0 , \5192_b0 , w_16906 );
not ( w_16906 , w_16907 );
and ( w_16907 , \5180_b1 , \5180_b0 );
or ( \5340_b1 , \5339_b1 , \5200_b1 );
not ( \5200_b1 , w_16908 );
and ( \5340_b0 , \5339_b0 , w_16909 );
and ( w_16908 , w_16909 , \5200_b0 );
buf ( \5341_b1 , \5339_b1 );
not ( \5341_b1 , w_16910 );
not ( \5341_b0 , w_16911 );
and ( w_16910 , w_16911 , \5339_b0 );
buf ( \5342_b1 , \5200_b1 );
not ( \5342_b1 , w_16912 );
not ( \5342_b0 , w_16913 );
and ( w_16912 , w_16913 , \5200_b0 );
or ( \5343_b1 , \5341_b1 , \5342_b1 );
not ( \5342_b1 , w_16914 );
and ( \5343_b0 , \5341_b0 , w_16915 );
and ( w_16914 , w_16915 , \5342_b0 );
or ( \5344_b1 , \5340_b1 , w_16917 );
not ( w_16917 , w_16918 );
and ( \5344_b0 , \5340_b0 , w_16919 );
and ( w_16918 ,  , w_16919 );
buf ( w_16917 , \5343_b1 );
not ( w_16917 , w_16920 );
not (  , w_16921 );
and ( w_16920 , w_16921 , \5343_b0 );
or ( \5345_b1 , \5338_b1 , w_16923 );
not ( w_16923 , w_16924 );
and ( \5345_b0 , \5338_b0 , w_16925 );
and ( w_16924 ,  , w_16925 );
buf ( w_16923 , \5344_b1 );
not ( w_16923 , w_16926 );
not (  , w_16927 );
and ( w_16926 , w_16927 , \5344_b0 );
buf ( \5346_b1 , \5336_b1 );
not ( \5346_b1 , w_16928 );
not ( \5346_b0 , w_16929 );
and ( w_16928 , w_16929 , \5336_b0 );
buf ( \5347_b1 , \5296_b1 );
buf ( \5347_b0 , \5296_b0 );
or ( \5348_b1 , \5346_b1 , w_16931 );
not ( w_16931 , w_16932 );
and ( \5348_b0 , \5346_b0 , w_16933 );
and ( w_16932 ,  , w_16933 );
buf ( w_16931 , \5347_b1 );
not ( w_16931 , w_16934 );
not (  , w_16935 );
and ( w_16934 , w_16935 , \5347_b0 );
or ( \5349_b1 , \5345_b1 , w_16937 );
not ( w_16937 , w_16938 );
and ( \5349_b0 , \5345_b0 , w_16939 );
and ( w_16938 ,  , w_16939 );
buf ( w_16937 , \5348_b1 );
not ( w_16937 , w_16940 );
not (  , w_16941 );
and ( w_16940 , w_16941 , \5348_b0 );
buf ( \5350_b1 , \5349_b1 );
buf ( \5350_b0 , \5349_b0 );
or ( \5351_b1 , \5265_b1 , \5350_b1 );
not ( \5350_b1 , w_16942 );
and ( \5351_b0 , \5265_b0 , w_16943 );
and ( w_16942 , w_16943 , \5350_b0 );
or ( \5352_b1 , \5262_b1 , w_16945 );
not ( w_16945 , w_16946 );
and ( \5352_b0 , \5262_b0 , w_16947 );
and ( w_16946 ,  , w_16947 );
buf ( w_16945 , \5264_b1 );
not ( w_16945 , w_16948 );
not (  , w_16949 );
and ( w_16948 , w_16949 , \5264_b0 );
or ( \5353_b1 , \5351_b1 , w_16951 );
not ( w_16951 , w_16952 );
and ( \5353_b0 , \5351_b0 , w_16953 );
and ( w_16952 ,  , w_16953 );
buf ( w_16951 , \5352_b1 );
not ( w_16951 , w_16954 );
not (  , w_16955 );
and ( w_16954 , w_16955 , \5352_b0 );
or ( \5354_b1 , \5220_b1 , \5353_b1 );
xor ( \5354_b0 , \5220_b0 , w_16956 );
not ( w_16956 , w_16957 );
and ( w_16957 , \5353_b1 , \5353_b0 );
or ( \5355_b1 , \5349_b1 , \5264_b1 );
xor ( \5355_b0 , \5349_b0 , w_16958 );
not ( w_16958 , w_16959 );
and ( w_16959 , \5264_b1 , \5264_b0 );
or ( \5356_b1 , \5355_b1 , w_16960 );
xor ( \5356_b0 , \5355_b0 , w_16962 );
not ( w_16962 , w_16963 );
and ( w_16963 , w_16960 , w_16961 );
buf ( w_16960 , \5261_b1 );
not ( w_16960 , w_16964 );
not ( w_16961 , w_16965 );
and ( w_16964 , w_16965 , \5261_b0 );
buf ( \5357_b1 , \5356_b1 );
not ( \5357_b1 , w_16966 );
not ( \5357_b0 , w_16967 );
and ( w_16966 , w_16967 , \5356_b0 );
buf ( \5358_b1 , \5079_b1 );
not ( \5358_b1 , w_16968 );
not ( \5358_b0 , w_16969 );
and ( w_16968 , w_16969 , \5079_b0 );
buf ( \5359_b1 , \5127_b1 );
not ( \5359_b1 , w_16970 );
not ( \5359_b0 , w_16971 );
and ( w_16970 , w_16971 , \5127_b0 );
buf ( \5360_b1 , \5359_b1 );
not ( \5360_b1 , w_16972 );
not ( \5360_b0 , w_16973 );
and ( w_16972 , w_16973 , \5359_b0 );
or ( \5361_b1 , \5358_b1 , w_16974 );
or ( \5361_b0 , \5358_b0 , \5360_b0 );
not ( \5360_b0 , w_16975 );
and ( w_16975 , w_16974 , \5360_b1 );
or ( \5362_b1 , \5078_b1 , w_16977 );
not ( w_16977 , w_16978 );
and ( \5362_b0 , \5078_b0 , w_16979 );
and ( w_16978 ,  , w_16979 );
buf ( w_16977 , \5127_b1 );
not ( w_16977 , w_16980 );
not (  , w_16981 );
and ( w_16980 , w_16981 , \5127_b0 );
or ( \5363_b1 , \5361_b1 , w_16983 );
not ( w_16983 , w_16984 );
and ( \5363_b0 , \5361_b0 , w_16985 );
and ( w_16984 ,  , w_16985 );
buf ( w_16983 , \5362_b1 );
not ( w_16983 , w_16986 );
not (  , w_16987 );
and ( w_16986 , w_16987 , \5362_b0 );
buf ( \5364_b1 , \5083_b1 );
not ( \5364_b1 , w_16988 );
not ( \5364_b0 , w_16989 );
and ( w_16988 , w_16989 , \5083_b0 );
or ( \5365_b1 , \5363_b1 , \5364_b1 );
not ( \5364_b1 , w_16990 );
and ( \5365_b0 , \5363_b0 , w_16991 );
and ( w_16990 , w_16991 , \5364_b0 );
buf ( \5366_b1 , \5363_b1 );
not ( \5366_b1 , w_16992 );
not ( \5366_b0 , w_16993 );
and ( w_16992 , w_16993 , \5363_b0 );
or ( \5367_b1 , \5366_b1 , \5083_b1 );
not ( \5083_b1 , w_16994 );
and ( \5367_b0 , \5366_b0 , w_16995 );
and ( w_16994 , w_16995 , \5083_b0 );
or ( \5368_b1 , \5365_b1 , w_16997 );
not ( w_16997 , w_16998 );
and ( \5368_b0 , \5365_b0 , w_16999 );
and ( w_16998 ,  , w_16999 );
buf ( w_16997 , \5367_b1 );
not ( w_16997 , w_17000 );
not (  , w_17001 );
and ( w_17000 , w_17001 , \5367_b0 );
buf ( \5369_b1 , \5368_b1 );
buf ( \5369_b0 , \5368_b0 );
buf ( \5370_b1 , \5369_b1 );
not ( \5370_b1 , w_17002 );
not ( \5370_b0 , w_17003 );
and ( w_17002 , w_17003 , \5369_b0 );
or ( \5371_b1 , \5357_b1 , w_17005 );
not ( w_17005 , w_17006 );
and ( \5371_b0 , \5357_b0 , w_17007 );
and ( w_17006 ,  , w_17007 );
buf ( w_17005 , \5370_b1 );
not ( w_17005 , w_17008 );
not (  , w_17009 );
and ( w_17008 , w_17009 , \5370_b0 );
buf ( \5372_b1 , \4198_b1 );
not ( \5372_b1 , w_17010 );
not ( \5372_b0 , w_17011 );
and ( w_17010 , w_17011 , \4198_b0 );
buf ( \5373_b1 , \4935_b1 );
not ( \5373_b1 , w_17012 );
not ( \5373_b0 , w_17013 );
and ( w_17012 , w_17013 , \4935_b0 );
or ( \5374_b1 , \5372_b1 , w_17014 );
or ( \5374_b0 , \5372_b0 , \5373_b0 );
not ( \5373_b0 , w_17015 );
and ( w_17015 , w_17014 , \5373_b1 );
or ( \5375_b1 , \4934_b1 , w_17017 );
not ( w_17017 , w_17018 );
and ( \5375_b0 , \4934_b0 , w_17019 );
and ( w_17018 ,  , w_17019 );
buf ( w_17017 , \4209_b1 );
not ( w_17017 , w_17020 );
not (  , w_17021 );
and ( w_17020 , w_17021 , \4209_b0 );
or ( \5376_b1 , \5374_b1 , w_17023 );
not ( w_17023 , w_17024 );
and ( \5376_b0 , \5374_b0 , w_17025 );
and ( w_17024 ,  , w_17025 );
buf ( w_17023 , \5375_b1 );
not ( w_17023 , w_17026 );
not (  , w_17027 );
and ( w_17026 , w_17027 , \5375_b0 );
buf ( \5377_b1 , \5376_b1 );
not ( \5377_b1 , w_17028 );
not ( \5377_b0 , w_17029 );
and ( w_17028 , w_17029 , \5376_b0 );
buf ( \5378_b1 , \4944_b1 );
not ( \5378_b1 , w_17030 );
not ( \5378_b0 , w_17031 );
and ( w_17030 , w_17031 , \4944_b0 );
or ( \5379_b1 , \5377_b1 , w_17032 );
or ( \5379_b0 , \5377_b0 , \5378_b0 );
not ( \5378_b0 , w_17033 );
and ( w_17033 , w_17032 , \5378_b1 );
or ( \5380_b1 , \4863_b1 , w_17035 );
not ( w_17035 , w_17036 );
and ( \5380_b0 , \4863_b0 , w_17037 );
and ( w_17036 ,  , w_17037 );
buf ( w_17035 , \5107_b1 );
not ( w_17035 , w_17038 );
not (  , w_17039 );
and ( w_17038 , w_17039 , \5107_b0 );
or ( \5381_b1 , \5379_b1 , w_17041 );
not ( w_17041 , w_17042 );
and ( \5381_b0 , \5379_b0 , w_17043 );
and ( w_17042 ,  , w_17043 );
buf ( w_17041 , \5380_b1 );
not ( w_17041 , w_17044 );
not (  , w_17045 );
and ( w_17044 , w_17045 , \5380_b0 );
buf ( \5382_b1 , \5381_b1 );
not ( \5382_b1 , w_17046 );
not ( \5382_b0 , w_17047 );
and ( w_17046 , w_17047 , \5381_b0 );
buf ( \5383_b1 , \4072_b1 );
not ( \5383_b1 , w_17048 );
not ( \5383_b0 , w_17049 );
and ( w_17048 , w_17049 , \4072_b0 );
buf ( \5384_b1 , \5183_b1 );
not ( \5384_b1 , w_17050 );
not ( \5384_b0 , w_17051 );
and ( w_17050 , w_17051 , \5183_b0 );
or ( \5385_b1 , \5383_b1 , w_17052 );
or ( \5385_b0 , \5383_b0 , \5384_b0 );
not ( \5384_b0 , w_17053 );
and ( w_17053 , w_17052 , \5384_b1 );
or ( \5386_b1 , \4110_b1 , w_17055 );
not ( w_17055 , w_17056 );
and ( \5386_b0 , \4110_b0 , w_17057 );
and ( w_17056 ,  , w_17057 );
buf ( w_17055 , \5089_b1 );
not ( w_17055 , w_17058 );
not (  , w_17059 );
and ( w_17058 , w_17059 , \5089_b0 );
or ( \5387_b1 , \5385_b1 , w_17061 );
not ( w_17061 , w_17062 );
and ( \5387_b0 , \5385_b0 , w_17063 );
and ( w_17062 ,  , w_17063 );
buf ( w_17061 , \5386_b1 );
not ( w_17061 , w_17064 );
not (  , w_17065 );
and ( w_17064 , w_17065 , \5386_b0 );
buf ( \5388_b1 , \5387_b1 );
not ( \5388_b1 , w_17066 );
not ( \5388_b0 , w_17067 );
and ( w_17066 , w_17067 , \5387_b0 );
buf ( \5389_b1 , \4128_b1 );
not ( \5389_b1 , w_17068 );
not ( \5389_b0 , w_17069 );
and ( w_17068 , w_17069 , \4128_b0 );
or ( \5390_b1 , \5388_b1 , w_17070 );
or ( \5390_b0 , \5388_b0 , \5389_b0 );
not ( \5389_b0 , w_17071 );
and ( w_17071 , w_17070 , \5389_b1 );
or ( \5391_b1 , \4132_b1 , w_17073 );
not ( w_17073 , w_17074 );
and ( \5391_b0 , \4132_b0 , w_17075 );
and ( w_17074 ,  , w_17075 );
buf ( w_17073 , \5253_b1 );
not ( w_17073 , w_17076 );
not (  , w_17077 );
and ( w_17076 , w_17077 , \5253_b0 );
or ( \5392_b1 , \5390_b1 , w_17079 );
not ( w_17079 , w_17080 );
and ( \5392_b0 , \5390_b0 , w_17081 );
and ( w_17080 ,  , w_17081 );
buf ( w_17079 , \5391_b1 );
not ( w_17079 , w_17082 );
not (  , w_17083 );
and ( w_17082 , w_17083 , \5391_b0 );
buf ( \5393_b1 , \5392_b1 );
not ( \5393_b1 , w_17084 );
not ( \5393_b0 , w_17085 );
and ( w_17084 , w_17085 , \5392_b0 );
buf ( \5394_b1 , \5393_b1 );
not ( \5394_b1 , w_17086 );
not ( \5394_b0 , w_17087 );
and ( w_17086 , w_17087 , \5393_b0 );
buf ( \5395_b1 , \5394_b1 );
not ( \5395_b1 , w_17088 );
not ( \5395_b0 , w_17089 );
and ( w_17088 , w_17089 , \5394_b0 );
or ( \5396_b1 , \5382_b1 , w_17090 );
or ( \5396_b0 , \5382_b0 , \5395_b0 );
not ( \5395_b0 , w_17091 );
and ( w_17091 , w_17090 , \5395_b1 );
buf ( \5397_b1 , \5381_b1 );
not ( \5397_b1 , w_17092 );
not ( \5397_b0 , w_17093 );
and ( w_17092 , w_17093 , \5381_b0 );
buf ( \5398_b1 , \5397_b1 );
not ( \5398_b1 , w_17094 );
not ( \5398_b0 , w_17095 );
and ( w_17094 , w_17095 , \5397_b0 );
buf ( \5399_b1 , \5393_b1 );
not ( \5399_b1 , w_17096 );
not ( \5399_b0 , w_17097 );
and ( w_17096 , w_17097 , \5393_b0 );
or ( \5400_b1 , \5398_b1 , w_17098 );
or ( \5400_b0 , \5398_b0 , \5399_b0 );
not ( \5399_b0 , w_17099 );
and ( w_17099 , w_17098 , \5399_b1 );
buf ( \5401_b1 , \4780_b1 );
not ( \5401_b1 , w_17100 );
not ( \5401_b0 , w_17101 );
and ( w_17100 , w_17101 , \4780_b0 );
buf ( \5402_b1 , \4311_b1 );
not ( \5402_b1 , w_17102 );
not ( \5402_b0 , w_17103 );
and ( w_17102 , w_17103 , \4311_b0 );
or ( \5403_b1 , \5401_b1 , w_17104 );
or ( \5403_b0 , \5401_b0 , \5402_b0 );
not ( \5402_b0 , w_17105 );
and ( w_17105 , w_17104 , \5402_b1 );
or ( \5404_b1 , \4163_b1 , w_17107 );
not ( w_17107 , w_17108 );
and ( \5404_b0 , \4163_b0 , w_17109 );
and ( w_17108 ,  , w_17109 );
buf ( w_17107 , \4021_b1 );
not ( w_17107 , w_17110 );
not (  , w_17111 );
and ( w_17110 , w_17111 , \4021_b0 );
or ( \5405_b1 , \5403_b1 , w_17113 );
not ( w_17113 , w_17114 );
and ( \5405_b0 , \5403_b0 , w_17115 );
and ( w_17114 ,  , w_17115 );
buf ( w_17113 , \5404_b1 );
not ( w_17113 , w_17116 );
not (  , w_17117 );
and ( w_17116 , w_17117 , \5404_b0 );
buf ( \5406_b1 , \5405_b1 );
not ( \5406_b1 , w_17118 );
not ( \5406_b0 , w_17119 );
and ( w_17118 , w_17119 , \5405_b0 );
buf ( \5407_b1 , \4159_b1 );
not ( \5407_b1 , w_17120 );
not ( \5407_b0 , w_17121 );
and ( w_17120 , w_17121 , \4159_b0 );
or ( \5408_b1 , \5406_b1 , w_17122 );
or ( \5408_b0 , \5406_b0 , \5407_b0 );
not ( \5407_b0 , w_17123 );
and ( w_17123 , w_17122 , \5407_b1 );
or ( \5409_b1 , \4317_b1 , w_17125 );
not ( w_17125 , w_17126 );
and ( \5409_b0 , \4317_b0 , w_17127 );
and ( w_17126 ,  , w_17127 );
buf ( w_17125 , \5315_b1 );
not ( w_17125 , w_17128 );
not (  , w_17129 );
and ( w_17128 , w_17129 , \5315_b0 );
or ( \5410_b1 , \5408_b1 , w_17131 );
not ( w_17131 , w_17132 );
and ( \5410_b0 , \5408_b0 , w_17133 );
and ( w_17132 ,  , w_17133 );
buf ( w_17131 , \5409_b1 );
not ( w_17131 , w_17134 );
not (  , w_17135 );
and ( w_17134 , w_17135 , \5409_b0 );
or ( \5411_b1 , \5400_b1 , w_17137 );
not ( w_17137 , w_17138 );
and ( \5411_b0 , \5400_b0 , w_17139 );
and ( w_17138 ,  , w_17139 );
buf ( w_17137 , \5410_b1 );
not ( w_17137 , w_17140 );
not (  , w_17141 );
and ( w_17140 , w_17141 , \5410_b0 );
or ( \5412_b1 , \5396_b1 , w_17143 );
not ( w_17143 , w_17144 );
and ( \5412_b0 , \5396_b0 , w_17145 );
and ( w_17144 ,  , w_17145 );
buf ( w_17143 , \5411_b1 );
not ( w_17143 , w_17146 );
not (  , w_17147 );
and ( w_17146 , w_17147 , \5411_b0 );
buf ( \5413_b1 , \5412_b1 );
not ( \5413_b1 , w_17148 );
not ( \5413_b0 , w_17149 );
and ( w_17148 , w_17149 , \5412_b0 );
or ( \5414_b1 , \5276_b1 , \5294_b1 );
xor ( \5414_b0 , \5276_b0 , w_17150 );
not ( w_17150 , w_17151 );
and ( w_17151 , \5294_b1 , \5294_b0 );
or ( \5415_b1 , \5414_b1 , w_17152 );
xor ( \5415_b0 , \5414_b0 , w_17154 );
not ( w_17154 , w_17155 );
and ( w_17155 , w_17152 , w_17153 );
buf ( w_17152 , \5291_b1 );
not ( w_17152 , w_17156 );
not ( w_17153 , w_17157 );
and ( w_17156 , w_17157 , \5291_b0 );
or ( \5416_b1 , \5413_b1 , w_17159 );
not ( w_17159 , w_17160 );
and ( \5416_b0 , \5413_b0 , w_17161 );
and ( w_17160 ,  , w_17161 );
buf ( w_17159 , \5415_b1 );
not ( w_17159 , w_17162 );
not (  , w_17163 );
and ( w_17162 , w_17163 , \5415_b0 );
buf ( \5417_b1 , \5416_b1 );
not ( \5417_b1 , w_17164 );
not ( \5417_b0 , w_17165 );
and ( w_17164 , w_17165 , \5416_b0 );
buf ( \5418_b1 , \4098_b1 );
not ( \5418_b1 , w_17166 );
not ( \5418_b0 , w_17167 );
and ( w_17166 , w_17167 , \4098_b0 );
or ( \5419_b1 , \4388_b1 , w_17169 );
not ( w_17169 , w_17170 );
and ( \5419_b0 , \4388_b0 , w_17171 );
and ( w_17170 ,  , w_17171 );
buf ( w_17169 , \5418_b1 );
not ( w_17169 , w_17172 );
not (  , w_17173 );
and ( w_17172 , w_17173 , \5418_b0 );
buf ( \5420_b1 , \5271_b1 );
not ( \5420_b1 , w_17174 );
not ( \5420_b0 , w_17175 );
and ( w_17174 , w_17175 , \5271_b0 );
buf ( \5421_b1 , \3997_b1 );
not ( \5421_b1 , w_17176 );
not ( \5421_b0 , w_17177 );
and ( w_17176 , w_17177 , \3997_b0 );
buf ( \5422_b1 , \5268_b1 );
not ( \5422_b1 , w_17178 );
not ( \5422_b0 , w_17179 );
and ( w_17178 , w_17179 , \5268_b0 );
buf ( \5423_b1 , \5422_b1 );
not ( \5423_b1 , w_17180 );
not ( \5423_b0 , w_17181 );
and ( w_17180 , w_17181 , \5422_b0 );
or ( \5424_b1 , \5421_b1 , w_17182 );
or ( \5424_b0 , \5421_b0 , \5423_b0 );
not ( \5423_b0 , w_17183 );
and ( w_17183 , w_17182 , \5423_b1 );
buf ( \5425_b1 , \5422_b1 );
not ( \5425_b1 , w_17184 );
not ( \5425_b0 , w_17185 );
and ( w_17184 , w_17185 , \5422_b0 );
or ( \5426_b1 , \5425_b1 , w_17187 );
not ( w_17187 , w_17188 );
and ( \5426_b0 , \5425_b0 , w_17189 );
and ( w_17188 ,  , w_17189 );
buf ( w_17187 , \4111_b1 );
not ( w_17187 , w_17190 );
not (  , w_17191 );
and ( w_17190 , w_17191 , \4111_b0 );
or ( \5427_b1 , \5424_b1 , w_17193 );
not ( w_17193 , w_17194 );
and ( \5427_b0 , \5424_b0 , w_17195 );
and ( w_17194 ,  , w_17195 );
buf ( w_17193 , \5426_b1 );
not ( w_17193 , w_17196 );
not (  , w_17197 );
and ( w_17196 , w_17197 , \5426_b0 );
buf ( \5428_b1 , \5427_b1 );
not ( \5428_b1 , w_17198 );
not ( \5428_b0 , w_17199 );
and ( w_17198 , w_17199 , \5427_b0 );
or ( \5429_b1 , \5420_b1 , w_17200 );
or ( \5429_b0 , \5420_b0 , \5428_b0 );
not ( \5428_b0 , w_17201 );
and ( w_17201 , w_17200 , \5428_b1 );
buf ( \5430_b1 , \4051_b1 );
not ( \5430_b1 , w_17202 );
not ( \5430_b0 , w_17203 );
and ( w_17202 , w_17203 , \4051_b0 );
buf ( \5431_b1 , \5422_b1 );
not ( \5431_b1 , w_17204 );
not ( \5431_b0 , w_17205 );
and ( w_17204 , w_17205 , \5422_b0 );
or ( \5432_b1 , \5430_b1 , w_17206 );
or ( \5432_b0 , \5430_b0 , \5431_b0 );
not ( \5431_b0 , w_17207 );
and ( w_17207 , w_17206 , \5431_b1 );
buf ( \5433_b1 , \5268_b1 );
buf ( \5433_b0 , \5268_b0 );
or ( \5434_b1 , \5433_b1 , w_17209 );
not ( w_17209 , w_17210 );
and ( \5434_b0 , \5433_b0 , w_17211 );
and ( w_17210 ,  , w_17211 );
buf ( w_17209 , \4135_b1 );
not ( w_17209 , w_17212 );
not (  , w_17213 );
and ( w_17212 , w_17213 , \4135_b0 );
or ( \5435_b1 , \5432_b1 , w_17215 );
not ( w_17215 , w_17216 );
and ( \5435_b0 , \5432_b0 , w_17217 );
and ( w_17216 ,  , w_17217 );
buf ( w_17215 , \5434_b1 );
not ( w_17215 , w_17218 );
not (  , w_17219 );
and ( w_17218 , w_17219 , \5434_b0 );
or ( \5436_b1 , \5435_b1 , w_17221 );
not ( w_17221 , w_17222 );
and ( \5436_b0 , \5435_b0 , w_17223 );
and ( w_17222 ,  , w_17223 );
buf ( w_17221 , \5266_b1 );
not ( w_17221 , w_17224 );
not (  , w_17225 );
and ( w_17224 , w_17225 , \5266_b0 );
or ( \5437_b1 , \5429_b1 , w_17227 );
not ( w_17227 , w_17228 );
and ( \5437_b0 , \5429_b0 , w_17229 );
and ( w_17228 ,  , w_17229 );
buf ( w_17227 , \5436_b1 );
not ( w_17227 , w_17230 );
not (  , w_17231 );
and ( w_17230 , w_17231 , \5436_b0 );
or ( \5438_b1 , \5419_b1 , \5437_b1 );
xor ( \5438_b0 , \5419_b0 , w_17232 );
not ( w_17232 , w_17233 );
and ( w_17233 , \5437_b1 , \5437_b0 );
or ( \5439_b1 , \4935_b1 , \4094_b1 );
not ( \4094_b1 , w_17234 );
and ( \5439_b0 , \4935_b0 , w_17235 );
and ( w_17234 , w_17235 , \4094_b0 );
or ( \5440_b1 , \4934_b1 , \4298_b1 );
not ( \4298_b1 , w_17236 );
and ( \5440_b0 , \4934_b0 , w_17237 );
and ( w_17236 , w_17237 , \4298_b0 );
or ( \5441_b1 , \5439_b1 , w_17239 );
not ( w_17239 , w_17240 );
and ( \5441_b0 , \5439_b0 , w_17241 );
and ( w_17240 ,  , w_17241 );
buf ( w_17239 , \5440_b1 );
not ( w_17239 , w_17242 );
not (  , w_17243 );
and ( w_17242 , w_17243 , \5440_b0 );
or ( \5442_b1 , \4943_b1 , w_17244 );
or ( \5442_b0 , \4943_b0 , \5441_b0 );
not ( \5441_b0 , w_17245 );
and ( w_17245 , w_17244 , \5441_b1 );
buf ( \5443_b1 , \5376_b1 );
not ( \5443_b1 , w_17246 );
not ( \5443_b0 , w_17247 );
and ( w_17246 , w_17247 , \5376_b0 );
or ( \5444_b1 , \5443_b1 , w_17248 );
or ( \5444_b0 , \5443_b0 , \4862_b0 );
not ( \4862_b0 , w_17249 );
and ( w_17249 , w_17248 , \4862_b1 );
or ( \5445_b1 , \5442_b1 , w_17251 );
not ( w_17251 , w_17252 );
and ( \5445_b0 , \5442_b0 , w_17253 );
and ( w_17252 ,  , w_17253 );
buf ( w_17251 , \5444_b1 );
not ( w_17251 , w_17254 );
not (  , w_17255 );
and ( w_17254 , w_17255 , \5444_b0 );
or ( \5446_b1 , \5438_b1 , \5445_b1 );
not ( \5445_b1 , w_17256 );
and ( \5446_b0 , \5438_b0 , w_17257 );
and ( w_17256 , w_17257 , \5445_b0 );
or ( \5447_b1 , \5419_b1 , \5437_b1 );
not ( \5437_b1 , w_17258 );
and ( \5447_b0 , \5419_b0 , w_17259 );
and ( w_17258 , w_17259 , \5437_b0 );
or ( \5448_b1 , \5446_b1 , w_17260 );
or ( \5448_b0 , \5446_b0 , \5447_b0 );
not ( \5447_b0 , w_17261 );
and ( w_17261 , w_17260 , \5447_b1 );
buf ( \5449_b1 , \4969_b1 );
not ( \5449_b1 , w_17262 );
not ( \5449_b0 , w_17263 );
and ( w_17262 , w_17263 , \4969_b0 );
buf ( \5450_b1 , \4311_b1 );
not ( \5450_b1 , w_17264 );
not ( \5450_b0 , w_17265 );
and ( w_17264 , w_17265 , \4311_b0 );
or ( \5451_b1 , \5449_b1 , w_17266 );
or ( \5451_b0 , \5449_b0 , \5450_b0 );
not ( \5450_b0 , w_17267 );
and ( w_17267 , w_17266 , \5450_b1 );
or ( \5452_b1 , \4163_b1 , w_17269 );
not ( w_17269 , w_17270 );
and ( \5452_b0 , \4163_b0 , w_17271 );
and ( w_17270 ,  , w_17271 );
buf ( w_17269 , \4026_b1 );
not ( w_17269 , w_17272 );
not (  , w_17273 );
and ( w_17272 , w_17273 , \4026_b0 );
or ( \5453_b1 , \5451_b1 , w_17275 );
not ( w_17275 , w_17276 );
and ( \5453_b0 , \5451_b0 , w_17277 );
and ( w_17276 ,  , w_17277 );
buf ( w_17275 , \5452_b1 );
not ( w_17275 , w_17278 );
not (  , w_17279 );
and ( w_17278 , w_17279 , \5452_b0 );
buf ( \5454_b1 , \5453_b1 );
not ( \5454_b1 , w_17280 );
not ( \5454_b0 , w_17281 );
and ( w_17280 , w_17281 , \5453_b0 );
buf ( \5455_b1 , \4158_b1 );
not ( \5455_b1 , w_17282 );
not ( \5455_b0 , w_17283 );
and ( w_17282 , w_17283 , \4158_b0 );
or ( \5456_b1 , \5454_b1 , w_17284 );
or ( \5456_b0 , \5454_b0 , \5455_b0 );
not ( \5455_b0 , w_17285 );
and ( w_17285 , w_17284 , \5455_b1 );
or ( \5457_b1 , \5405_b1 , w_17287 );
not ( w_17287 , w_17288 );
and ( \5457_b0 , \5405_b0 , w_17289 );
and ( w_17288 ,  , w_17289 );
buf ( w_17287 , \4150_b1 );
not ( w_17287 , w_17290 );
not (  , w_17291 );
and ( w_17290 , w_17291 , \4150_b0 );
or ( \5458_b1 , \5456_b1 , w_17293 );
not ( w_17293 , w_17294 );
and ( \5458_b0 , \5456_b0 , w_17295 );
and ( w_17294 ,  , w_17295 );
buf ( w_17293 , \5457_b1 );
not ( w_17293 , w_17296 );
not (  , w_17297 );
and ( w_17296 , w_17297 , \5457_b0 );
buf ( \5459_b1 , \5458_b1 );
not ( \5459_b1 , w_17298 );
not ( \5459_b0 , w_17299 );
and ( w_17298 , w_17299 , \5458_b0 );
buf ( \5460_b1 , \4610_b1 );
not ( \5460_b1 , w_17300 );
not ( \5460_b0 , w_17301 );
and ( w_17300 , w_17301 , \4610_b0 );
buf ( \5461_b1 , \4097_b1 );
not ( \5461_b1 , w_17302 );
not ( \5461_b0 , w_17303 );
and ( w_17302 , w_17303 , \4097_b0 );
buf ( \5462_b1 , \4746_b1 );
not ( \5462_b1 , w_17304 );
not ( \5462_b0 , w_17305 );
and ( w_17304 , w_17305 , \4746_b0 );
or ( \5463_b1 , \5461_b1 , w_17306 );
or ( \5463_b0 , \5461_b0 , \5462_b0 );
not ( \5462_b0 , w_17307 );
and ( w_17307 , w_17306 , \5462_b1 );
or ( \5464_b1 , \4745_b1 , w_17309 );
not ( w_17309 , w_17310 );
and ( \5464_b0 , \4745_b0 , w_17311 );
and ( w_17310 ,  , w_17311 );
buf ( w_17309 , \4254_b1 );
not ( w_17309 , w_17312 );
not (  , w_17313 );
and ( w_17312 , w_17313 , \4254_b0 );
or ( \5465_b1 , \5463_b1 , w_17315 );
not ( w_17315 , w_17316 );
and ( \5465_b0 , \5463_b0 , w_17317 );
and ( w_17316 ,  , w_17317 );
buf ( w_17315 , \5464_b1 );
not ( w_17315 , w_17318 );
not (  , w_17319 );
and ( w_17318 , w_17319 , \5464_b0 );
buf ( \5466_b1 , \5465_b1 );
not ( \5466_b1 , w_17320 );
not ( \5466_b0 , w_17321 );
and ( w_17320 , w_17321 , \5465_b0 );
or ( \5467_b1 , \5460_b1 , w_17322 );
or ( \5467_b0 , \5460_b0 , \5466_b0 );
not ( \5466_b0 , w_17323 );
and ( w_17323 , w_17322 , \5466_b1 );
buf ( \5468_b1 , \4096_b1 );
not ( \5468_b1 , w_17324 );
not ( \5468_b0 , w_17325 );
and ( w_17324 , w_17325 , \4096_b0 );
buf ( \5469_b1 , \5138_b1 );
not ( \5469_b1 , w_17326 );
not ( \5469_b0 , w_17327 );
and ( w_17326 , w_17327 , \5138_b0 );
or ( \5470_b1 , \5468_b1 , w_17328 );
or ( \5470_b0 , \5468_b0 , \5469_b0 );
not ( \5469_b0 , w_17329 );
and ( w_17329 , w_17328 , \5469_b1 );
or ( \5471_b1 , \4615_b1 , w_17331 );
not ( w_17331 , w_17332 );
and ( \5471_b0 , \4615_b0 , w_17333 );
and ( w_17332 ,  , w_17333 );
buf ( w_17331 , \4372_b1 );
not ( w_17331 , w_17334 );
not (  , w_17335 );
and ( w_17334 , w_17335 , \4372_b0 );
or ( \5472_b1 , \5470_b1 , w_17337 );
not ( w_17337 , w_17338 );
and ( \5472_b0 , \5470_b0 , w_17339 );
and ( w_17338 ,  , w_17339 );
buf ( w_17337 , \5471_b1 );
not ( w_17337 , w_17340 );
not (  , w_17341 );
and ( w_17340 , w_17341 , \5471_b0 );
or ( \5473_b1 , \4754_b1 , w_17343 );
not ( w_17343 , w_17344 );
and ( \5473_b0 , \4754_b0 , w_17345 );
and ( w_17344 ,  , w_17345 );
buf ( w_17343 , \5472_b1 );
not ( w_17343 , w_17346 );
not (  , w_17347 );
and ( w_17346 , w_17347 , \5472_b0 );
or ( \5474_b1 , \5467_b1 , w_17349 );
not ( w_17349 , w_17350 );
and ( \5474_b0 , \5467_b0 , w_17351 );
and ( w_17350 ,  , w_17351 );
buf ( w_17349 , \5473_b1 );
not ( w_17349 , w_17352 );
not (  , w_17353 );
and ( w_17352 , w_17353 , \5473_b0 );
buf ( \5475_b1 , \5474_b1 );
not ( \5475_b1 , w_17354 );
not ( \5475_b0 , w_17355 );
and ( w_17354 , w_17355 , \5474_b0 );
or ( \5476_b1 , \5459_b1 , w_17356 );
or ( \5476_b0 , \5459_b0 , \5475_b0 );
not ( \5475_b0 , w_17357 );
and ( w_17357 , w_17356 , \5475_b1 );
or ( \5477_b1 , \5474_b1 , w_17358 );
or ( \5477_b0 , \5474_b0 , \5458_b0 );
not ( \5458_b0 , w_17359 );
and ( w_17359 , w_17358 , \5458_b1 );
buf ( \5478_b1 , \4076_b1 );
not ( \5478_b1 , w_17360 );
not ( \5478_b0 , w_17361 );
and ( w_17360 , w_17361 , \4076_b0 );
buf ( \5479_b1 , \4134_b1 );
not ( \5479_b1 , w_17362 );
not ( \5479_b0 , w_17363 );
and ( w_17362 , w_17363 , \4134_b0 );
or ( \5480_b1 , \5478_b1 , w_17364 );
or ( \5480_b0 , \5478_b0 , \5479_b0 );
not ( \5479_b0 , w_17365 );
and ( w_17365 , w_17364 , \5479_b1 );
or ( \5481_b1 , \4106_b1 , w_17367 );
not ( w_17367 , w_17368 );
and ( \5481_b0 , \4106_b0 , w_17369 );
and ( w_17368 ,  , w_17369 );
buf ( w_17367 , \5284_b1 );
not ( w_17367 , w_17370 );
not (  , w_17371 );
and ( w_17370 , w_17371 , \5284_b0 );
or ( \5482_b1 , \5480_b1 , w_17373 );
not ( w_17373 , w_17374 );
and ( \5482_b0 , \5480_b0 , w_17375 );
and ( w_17374 ,  , w_17375 );
buf ( w_17373 , \5481_b1 );
not ( w_17373 , w_17376 );
not (  , w_17377 );
and ( w_17376 , w_17377 , \5481_b0 );
buf ( \5483_b1 , \5482_b1 );
not ( \5483_b1 , w_17378 );
not ( \5483_b0 , w_17379 );
and ( w_17378 , w_17379 , \5482_b0 );
buf ( \5484_b1 , \4710_b1 );
not ( \5484_b1 , w_17380 );
not ( \5484_b0 , w_17381 );
and ( w_17380 , w_17381 , \4710_b0 );
or ( \5485_b1 , \5483_b1 , w_17382 );
or ( \5485_b0 , \5483_b0 , \5484_b0 );
not ( \5484_b0 , w_17383 );
and ( w_17383 , w_17382 , \5484_b1 );
or ( \5486_b1 , \5387_b1 , w_17385 );
not ( w_17385 , w_17386 );
and ( \5486_b0 , \5387_b0 , w_17387 );
and ( w_17386 ,  , w_17387 );
buf ( w_17385 , \4132_b1 );
not ( w_17385 , w_17388 );
not (  , w_17389 );
and ( w_17388 , w_17389 , \4132_b0 );
or ( \5487_b1 , \5485_b1 , w_17391 );
not ( w_17391 , w_17392 );
and ( \5487_b0 , \5485_b0 , w_17393 );
and ( w_17392 ,  , w_17393 );
buf ( w_17391 , \5486_b1 );
not ( w_17391 , w_17394 );
not (  , w_17395 );
and ( w_17394 , w_17395 , \5486_b0 );
or ( \5488_b1 , \5477_b1 , w_17397 );
not ( w_17397 , w_17398 );
and ( \5488_b0 , \5477_b0 , w_17399 );
and ( w_17398 ,  , w_17399 );
buf ( w_17397 , \5487_b1 );
not ( w_17397 , w_17400 );
not (  , w_17401 );
and ( w_17400 , w_17401 , \5487_b0 );
or ( \5489_b1 , \5476_b1 , w_17403 );
not ( w_17403 , w_17404 );
and ( \5489_b0 , \5476_b0 , w_17405 );
and ( w_17404 ,  , w_17405 );
buf ( w_17403 , \5488_b1 );
not ( w_17403 , w_17406 );
not (  , w_17407 );
and ( w_17406 , w_17407 , \5488_b0 );
or ( \5490_b1 , \5448_b1 , \5489_b1 );
xor ( \5490_b0 , \5448_b0 , w_17408 );
not ( w_17408 , w_17409 );
and ( w_17409 , \5489_b1 , \5489_b0 );
buf ( \5491_b1 , \4017_b1 );
not ( \5491_b1 , w_17410 );
not ( \5491_b0 , w_17411 );
and ( w_17410 , w_17411 , \4017_b0 );
buf ( \5492_b1 , \4332_b1 );
not ( \5492_b1 , w_17412 );
not ( \5492_b0 , w_17413 );
and ( w_17412 , w_17413 , \4332_b0 );
or ( \5493_b1 , \5491_b1 , w_17414 );
or ( \5493_b0 , \5491_b0 , \5492_b0 );
not ( \5492_b0 , w_17415 );
and ( w_17415 , w_17414 , \5492_b1 );
or ( \5494_b1 , \4283_b1 , w_17417 );
not ( w_17417 , w_17418 );
and ( \5494_b0 , \4283_b0 , w_17419 );
and ( w_17418 ,  , w_17419 );
buf ( w_17417 , \4662_b1 );
not ( w_17417 , w_17420 );
not (  , w_17421 );
and ( w_17420 , w_17421 , \4662_b0 );
or ( \5495_b1 , \5493_b1 , w_17423 );
not ( w_17423 , w_17424 );
and ( \5495_b0 , \5493_b0 , w_17425 );
and ( w_17424 ,  , w_17425 );
buf ( w_17423 , \5494_b1 );
not ( w_17423 , w_17426 );
not (  , w_17427 );
and ( w_17426 , w_17427 , \5494_b0 );
buf ( \5496_b1 , \5495_b1 );
not ( \5496_b1 , w_17428 );
not ( \5496_b0 , w_17429 );
and ( w_17428 , w_17429 , \5495_b0 );
buf ( \5497_b1 , \4278_b1 );
not ( \5497_b1 , w_17430 );
not ( \5497_b0 , w_17431 );
and ( w_17430 , w_17431 , \4278_b0 );
buf ( \5498_b1 , \5497_b1 );
not ( \5498_b1 , w_17432 );
not ( \5498_b0 , w_17433 );
and ( w_17432 , w_17433 , \5497_b0 );
or ( \5499_b1 , \5496_b1 , w_17434 );
or ( \5499_b0 , \5496_b0 , \5498_b0 );
not ( \5498_b0 , w_17435 );
and ( w_17435 , w_17434 , \5498_b1 );
buf ( \5500_b1 , \4066_b1 );
not ( \5500_b1 , w_17436 );
not ( \5500_b0 , w_17437 );
and ( w_17436 , w_17437 , \4066_b0 );
buf ( \5501_b1 , \4493_b1 );
not ( \5501_b1 , w_17438 );
not ( \5501_b0 , w_17439 );
and ( w_17438 , w_17439 , \4493_b0 );
or ( \5502_b1 , \5500_b1 , w_17440 );
or ( \5502_b0 , \5500_b0 , \5501_b0 );
not ( \5501_b0 , w_17441 );
and ( w_17441 , w_17440 , \5501_b1 );
or ( \5503_b1 , \4283_b1 , w_17443 );
not ( w_17443 , w_17444 );
and ( \5503_b0 , \4283_b0 , w_17445 );
and ( w_17444 ,  , w_17445 );
buf ( w_17443 , \4519_b1 );
not ( w_17443 , w_17446 );
not (  , w_17447 );
and ( w_17446 , w_17447 , \4519_b0 );
or ( \5504_b1 , \5502_b1 , w_17449 );
not ( w_17449 , w_17450 );
and ( \5504_b0 , \5502_b0 , w_17451 );
and ( w_17450 ,  , w_17451 );
buf ( w_17449 , \5503_b1 );
not ( w_17449 , w_17452 );
not (  , w_17453 );
and ( w_17452 , w_17453 , \5503_b0 );
or ( \5505_b1 , \5504_b1 , w_17455 );
not ( w_17455 , w_17456 );
and ( \5505_b0 , \5504_b0 , w_17457 );
and ( w_17456 ,  , w_17457 );
buf ( w_17455 , \4800_b1 );
not ( w_17455 , w_17458 );
not (  , w_17459 );
and ( w_17458 , w_17459 , \4800_b0 );
or ( \5506_b1 , \5499_b1 , w_17461 );
not ( w_17461 , w_17462 );
and ( \5506_b0 , \5499_b0 , w_17463 );
and ( w_17462 ,  , w_17463 );
buf ( w_17461 , \5505_b1 );
not ( w_17461 , w_17464 );
not (  , w_17465 );
and ( w_17464 , w_17465 , \5505_b0 );
buf ( \5507_b1 , \4449_b1 );
not ( \5507_b1 , w_17466 );
not ( \5507_b0 , w_17467 );
and ( w_17466 , w_17467 , \4449_b0 );
buf ( \5508_b1 , \4095_b1 );
not ( \5508_b1 , w_17468 );
not ( \5508_b0 , w_17469 );
and ( w_17468 , w_17469 , \4095_b0 );
buf ( \5509_b1 , \5112_b1 );
not ( \5509_b1 , w_17470 );
not ( \5509_b0 , w_17471 );
and ( w_17470 , w_17471 , \5112_b0 );
or ( \5510_b1 , \5508_b1 , w_17472 );
or ( \5510_b0 , \5508_b0 , \5509_b0 );
not ( \5509_b0 , w_17473 );
and ( w_17473 , w_17472 , \5509_b1 );
or ( \5511_b1 , \4536_b1 , w_17475 );
not ( w_17475 , w_17476 );
and ( \5511_b0 , \4536_b0 , w_17477 );
and ( w_17476 ,  , w_17477 );
buf ( w_17475 , \4391_b1 );
not ( w_17475 , w_17478 );
not (  , w_17479 );
and ( w_17478 , w_17479 , \4391_b0 );
or ( \5512_b1 , \5510_b1 , w_17481 );
not ( w_17481 , w_17482 );
and ( \5512_b0 , \5510_b0 , w_17483 );
and ( w_17482 ,  , w_17483 );
buf ( w_17481 , \5511_b1 );
not ( w_17481 , w_17484 );
not (  , w_17485 );
and ( w_17484 , w_17485 , \5511_b0 );
buf ( \5513_b1 , \5512_b1 );
not ( \5513_b1 , w_17486 );
not ( \5513_b0 , w_17487 );
and ( w_17486 , w_17487 , \5512_b0 );
or ( \5514_b1 , \5507_b1 , w_17488 );
or ( \5514_b0 , \5507_b0 , \5513_b0 );
not ( \5513_b0 , w_17489 );
and ( w_17489 , w_17488 , \5513_b1 );
buf ( \5515_b1 , \4093_b1 );
not ( \5515_b1 , w_17490 );
not ( \5515_b0 , w_17491 );
and ( w_17490 , w_17491 , \4093_b0 );
buf ( \5516_b1 , \5112_b1 );
not ( \5516_b1 , w_17492 );
not ( \5516_b0 , w_17493 );
and ( w_17492 , w_17493 , \5112_b0 );
or ( \5517_b1 , \5515_b1 , w_17494 );
or ( \5517_b0 , \5515_b0 , \5516_b0 );
not ( \5516_b0 , w_17495 );
and ( w_17495 , w_17494 , \5516_b1 );
or ( \5518_b1 , \4729_b1 , w_17497 );
not ( w_17497 , w_17498 );
and ( \5518_b0 , \4729_b0 , w_17499 );
and ( w_17498 ,  , w_17499 );
buf ( w_17497 , \4349_b1 );
not ( w_17497 , w_17500 );
not (  , w_17501 );
and ( w_17500 , w_17501 , \4349_b0 );
or ( \5519_b1 , \5517_b1 , w_17503 );
not ( w_17503 , w_17504 );
and ( \5519_b0 , \5517_b0 , w_17505 );
and ( w_17504 ,  , w_17505 );
buf ( w_17503 , \5518_b1 );
not ( w_17503 , w_17506 );
not (  , w_17507 );
and ( w_17506 , w_17507 , \5518_b0 );
or ( \5520_b1 , \5519_b1 , w_17509 );
not ( w_17509 , w_17510 );
and ( \5520_b0 , \5519_b0 , w_17511 );
and ( w_17510 ,  , w_17511 );
buf ( w_17509 , \4452_b1 );
not ( w_17509 , w_17512 );
not (  , w_17513 );
and ( w_17512 , w_17513 , \4452_b0 );
or ( \5521_b1 , \5514_b1 , w_17515 );
not ( w_17515 , w_17516 );
and ( \5521_b0 , \5514_b0 , w_17517 );
and ( w_17516 ,  , w_17517 );
buf ( w_17515 , \5520_b1 );
not ( w_17515 , w_17518 );
not (  , w_17519 );
and ( w_17518 , w_17519 , \5520_b0 );
or ( \5522_b1 , \5506_b1 , \5521_b1 );
xor ( \5522_b0 , \5506_b0 , w_17520 );
not ( w_17520 , w_17521 );
and ( w_17521 , \5521_b1 , \5521_b0 );
buf ( \5523_b1 , \4082_b1 );
not ( \5523_b1 , w_17522 );
not ( \5523_b0 , w_17523 );
and ( w_17522 , w_17523 , \4082_b0 );
buf ( \5524_b1 , \4388_b1 );
not ( \5524_b1 , w_17524 );
not ( \5524_b0 , w_17525 );
and ( w_17524 , w_17525 , \4388_b0 );
or ( \5525_b1 , \5523_b1 , w_17526 );
or ( \5525_b0 , \5523_b0 , \5524_b0 );
not ( \5524_b0 , w_17527 );
and ( w_17527 , w_17526 , \5524_b1 );
buf ( \5526_b1 , \4082_b1 );
not ( \5526_b1 , w_17528 );
not ( \5526_b0 , w_17529 );
and ( w_17528 , w_17529 , \4082_b0 );
or ( \5527_b1 , \4100_b1 , w_17531 );
not ( w_17531 , w_17532 );
and ( \5527_b0 , \4100_b0 , w_17533 );
and ( w_17532 ,  , w_17533 );
buf ( w_17531 , \5526_b1 );
not ( w_17531 , w_17534 );
not (  , w_17535 );
and ( w_17534 , w_17535 , \5526_b0 );
or ( \5528_b1 , \5525_b1 , w_17537 );
not ( w_17537 , w_17538 );
and ( \5528_b0 , \5525_b0 , w_17539 );
and ( w_17538 ,  , w_17539 );
buf ( w_17537 , \5527_b1 );
not ( w_17537 , w_17540 );
not (  , w_17541 );
and ( w_17540 , w_17541 , \5527_b0 );
buf ( \5529_b1 , \5528_b1 );
not ( \5529_b1 , w_17542 );
not ( \5529_b0 , w_17543 );
and ( w_17542 , w_17543 , \5528_b0 );
buf ( \5530_b1 , \4395_b1 );
not ( \5530_b1 , w_17544 );
not ( \5530_b0 , w_17545 );
and ( w_17544 , w_17545 , \4395_b0 );
or ( \5531_b1 , \5529_b1 , w_17546 );
or ( \5531_b0 , \5529_b0 , \5530_b0 );
not ( \5530_b0 , w_17547 );
and ( w_17547 , w_17546 , \5530_b1 );
buf ( \5532_b1 , \4079_b1 );
not ( \5532_b1 , w_17548 );
not ( \5532_b0 , w_17549 );
and ( w_17548 , w_17549 , \4079_b0 );
buf ( \5533_b1 , \4101_b1 );
not ( \5533_b1 , w_17550 );
not ( \5533_b0 , w_17551 );
and ( w_17550 , w_17551 , \4101_b0 );
or ( \5534_b1 , \5532_b1 , w_17552 );
or ( \5534_b0 , \5532_b0 , \5533_b0 );
not ( \5533_b0 , w_17553 );
and ( w_17553 , w_17552 , \5533_b1 );
buf ( \5535_b1 , \4079_b1 );
not ( \5535_b1 , w_17554 );
not ( \5535_b0 , w_17555 );
and ( w_17554 , w_17555 , \4079_b0 );
or ( \5536_b1 , \4100_b1 , w_17557 );
not ( w_17557 , w_17558 );
and ( \5536_b0 , \4100_b0 , w_17559 );
and ( w_17558 ,  , w_17559 );
buf ( w_17557 , \5535_b1 );
not ( w_17557 , w_17560 );
not (  , w_17561 );
and ( w_17560 , w_17561 , \5535_b0 );
or ( \5537_b1 , \5534_b1 , w_17563 );
not ( w_17563 , w_17564 );
and ( \5537_b0 , \5534_b0 , w_17565 );
and ( w_17564 ,  , w_17565 );
buf ( w_17563 , \5536_b1 );
not ( w_17563 , w_17566 );
not (  , w_17567 );
and ( w_17566 , w_17567 , \5536_b0 );
or ( \5538_b1 , \5537_b1 , w_17569 );
not ( w_17569 , w_17570 );
and ( \5538_b0 , \5537_b0 , w_17571 );
and ( w_17570 ,  , w_17571 );
buf ( w_17569 , \4200_b1 );
not ( w_17569 , w_17572 );
not (  , w_17573 );
and ( w_17572 , w_17573 , \4200_b0 );
or ( \5539_b1 , \5531_b1 , w_17575 );
not ( w_17575 , w_17576 );
and ( \5539_b0 , \5531_b0 , w_17577 );
and ( w_17576 ,  , w_17577 );
buf ( w_17575 , \5538_b1 );
not ( w_17575 , w_17578 );
not (  , w_17579 );
and ( w_17578 , w_17579 , \5538_b0 );
or ( \5540_b1 , \5522_b1 , \5539_b1 );
not ( \5539_b1 , w_17580 );
and ( \5540_b0 , \5522_b0 , w_17581 );
and ( w_17580 , w_17581 , \5539_b0 );
or ( \5541_b1 , \5506_b1 , \5521_b1 );
not ( \5521_b1 , w_17582 );
and ( \5541_b0 , \5506_b0 , w_17583 );
and ( w_17582 , w_17583 , \5521_b0 );
or ( \5542_b1 , \5540_b1 , w_17584 );
or ( \5542_b0 , \5540_b0 , \5541_b0 );
not ( \5541_b0 , w_17585 );
and ( w_17585 , w_17584 , \5541_b1 );
or ( \5543_b1 , \5490_b1 , \5542_b1 );
not ( \5542_b1 , w_17586 );
and ( \5543_b0 , \5490_b0 , w_17587 );
and ( w_17586 , w_17587 , \5542_b0 );
or ( \5544_b1 , \5448_b1 , \5489_b1 );
not ( \5489_b1 , w_17588 );
and ( \5544_b0 , \5448_b0 , w_17589 );
and ( w_17588 , w_17589 , \5489_b0 );
or ( \5545_b1 , \5543_b1 , w_17590 );
or ( \5545_b0 , \5543_b0 , \5544_b0 );
not ( \5544_b0 , w_17591 );
and ( w_17591 , w_17590 , \5544_b1 );
buf ( \5546_b1 , \5545_b1 );
not ( \5546_b1 , w_17592 );
not ( \5546_b0 , w_17593 );
and ( w_17592 , w_17593 , \5545_b0 );
or ( \5547_b1 , \5417_b1 , w_17594 );
or ( \5547_b0 , \5417_b0 , \5546_b0 );
not ( \5546_b0 , w_17595 );
and ( w_17595 , w_17594 , \5546_b1 );
buf ( \5548_b1 , \5415_b1 );
not ( \5548_b1 , w_17596 );
not ( \5548_b0 , w_17597 );
and ( w_17596 , w_17597 , \5415_b0 );
or ( \5549_b1 , \5548_b1 , w_17599 );
not ( w_17599 , w_17600 );
and ( \5549_b0 , \5548_b0 , w_17601 );
and ( w_17600 ,  , w_17601 );
buf ( w_17599 , \5412_b1 );
not ( w_17599 , w_17602 );
not (  , w_17603 );
and ( w_17602 , w_17603 , \5412_b0 );
or ( \5550_b1 , \5547_b1 , w_17605 );
not ( w_17605 , w_17606 );
and ( \5550_b0 , \5547_b0 , w_17607 );
and ( w_17606 ,  , w_17607 );
buf ( w_17605 , \5549_b1 );
not ( w_17605 , w_17608 );
not (  , w_17609 );
and ( w_17608 , w_17609 , \5549_b0 );
buf ( \5551_b1 , \5550_b1 );
not ( \5551_b1 , w_17610 );
not ( \5551_b0 , w_17611 );
and ( w_17610 , w_17611 , \5550_b0 );
or ( \5552_b1 , \5296_b1 , \5336_b1 );
not ( \5336_b1 , w_17612 );
and ( \5552_b0 , \5296_b0 , w_17613 );
and ( w_17612 , w_17613 , \5336_b0 );
buf ( \5553_b1 , \5296_b1 );
not ( \5553_b1 , w_17614 );
not ( \5553_b0 , w_17615 );
and ( w_17614 , w_17615 , \5296_b0 );
or ( \5554_b1 , \5553_b1 , \5335_b1 );
not ( \5335_b1 , w_17616 );
and ( \5554_b0 , \5553_b0 , w_17617 );
and ( w_17616 , w_17617 , \5335_b0 );
or ( \5555_b1 , \5552_b1 , w_17618 );
or ( \5555_b0 , \5552_b0 , \5554_b0 );
not ( \5554_b0 , w_17619 );
and ( w_17619 , w_17618 , \5554_b1 );
or ( \5556_b1 , \5555_b1 , \5344_b1 );
not ( \5344_b1 , w_17620 );
and ( \5556_b0 , \5555_b0 , w_17621 );
and ( w_17620 , w_17621 , \5344_b0 );
buf ( \5557_b1 , \5555_b1 );
not ( \5557_b1 , w_17622 );
not ( \5557_b0 , w_17623 );
and ( w_17622 , w_17623 , \5555_b0 );
buf ( \5558_b1 , \5344_b1 );
not ( \5558_b1 , w_17624 );
not ( \5558_b0 , w_17625 );
and ( w_17624 , w_17625 , \5344_b0 );
or ( \5559_b1 , \5557_b1 , \5558_b1 );
not ( \5558_b1 , w_17626 );
and ( \5559_b0 , \5557_b0 , w_17627 );
and ( w_17626 , w_17627 , \5558_b0 );
or ( \5560_b1 , \5556_b1 , w_17629 );
not ( w_17629 , w_17630 );
and ( \5560_b0 , \5556_b0 , w_17631 );
and ( w_17630 ,  , w_17631 );
buf ( w_17629 , \5559_b1 );
not ( w_17629 , w_17632 );
not (  , w_17633 );
and ( w_17632 , w_17633 , \5559_b0 );
buf ( \5561_b1 , \5560_b1 );
not ( \5561_b1 , w_17634 );
not ( \5561_b0 , w_17635 );
and ( w_17634 , w_17635 , \5560_b0 );
buf ( \5562_b1 , \5435_b1 );
not ( \5562_b1 , w_17636 );
not ( \5562_b0 , w_17637 );
and ( w_17636 , w_17637 , \5435_b0 );
buf ( \5563_b1 , \5271_b1 );
not ( \5563_b1 , w_17638 );
not ( \5563_b0 , w_17639 );
and ( w_17638 , w_17639 , \5271_b0 );
or ( \5564_b1 , \5562_b1 , w_17640 );
or ( \5564_b0 , \5562_b0 , \5563_b0 );
not ( \5563_b0 , w_17641 );
and ( w_17641 , w_17640 , \5563_b1 );
or ( \5565_b1 , \5275_b1 , w_17643 );
not ( w_17643 , w_17644 );
and ( \5565_b0 , \5275_b0 , w_17645 );
and ( w_17644 ,  , w_17645 );
buf ( w_17643 , \5266_b1 );
not ( w_17643 , w_17646 );
not (  , w_17647 );
and ( w_17646 , w_17647 , \5266_b0 );
or ( \5566_b1 , \5564_b1 , w_17649 );
not ( w_17649 , w_17650 );
and ( \5566_b0 , \5564_b0 , w_17651 );
and ( w_17650 ,  , w_17651 );
buf ( w_17649 , \5565_b1 );
not ( w_17649 , w_17652 );
not (  , w_17653 );
and ( w_17652 , w_17653 , \5565_b0 );
buf ( \5567_b1 , \5504_b1 );
not ( \5567_b1 , w_17654 );
not ( \5567_b0 , w_17655 );
and ( w_17654 , w_17655 , \5504_b0 );
buf ( \5568_b1 , \4797_b1 );
not ( \5568_b1 , w_17656 );
not ( \5568_b0 , w_17657 );
and ( w_17656 , w_17657 , \4797_b0 );
or ( \5569_b1 , \5567_b1 , w_17658 );
or ( \5569_b0 , \5567_b0 , \5568_b0 );
not ( \5568_b0 , w_17659 );
and ( w_17659 , w_17658 , \5568_b1 );
or ( \5570_b1 , \5328_b1 , w_17661 );
not ( w_17661 , w_17662 );
and ( \5570_b0 , \5328_b0 , w_17663 );
and ( w_17662 ,  , w_17663 );
buf ( w_17661 , \4800_b1 );
not ( w_17661 , w_17664 );
not (  , w_17665 );
and ( w_17664 , w_17665 , \4800_b0 );
or ( \5571_b1 , \5569_b1 , w_17667 );
not ( w_17667 , w_17668 );
and ( \5571_b0 , \5569_b0 , w_17669 );
and ( w_17668 ,  , w_17669 );
buf ( w_17667 , \5570_b1 );
not ( w_17667 , w_17670 );
not (  , w_17671 );
and ( w_17670 , w_17671 , \5570_b0 );
or ( \5572_b1 , \5566_b1 , \5571_b1 );
xor ( \5572_b0 , \5566_b0 , w_17672 );
not ( w_17672 , w_17673 );
and ( w_17673 , \5571_b1 , \5571_b0 );
buf ( \5573_b1 , \5472_b1 );
not ( \5573_b1 , w_17674 );
not ( \5573_b0 , w_17675 );
and ( w_17674 , w_17675 , \5472_b0 );
buf ( \5574_b1 , \4611_b1 );
not ( \5574_b1 , w_17676 );
not ( \5574_b0 , w_17677 );
and ( w_17676 , w_17677 , \4611_b0 );
or ( \5575_b1 , \5573_b1 , w_17678 );
or ( \5575_b0 , \5573_b0 , \5574_b0 );
not ( \5574_b0 , w_17679 );
and ( w_17679 , w_17678 , \5574_b1 );
or ( \5576_b1 , \5305_b1 , w_17681 );
not ( w_17681 , w_17682 );
and ( \5576_b0 , \5305_b0 , w_17683 );
and ( w_17682 ,  , w_17683 );
buf ( w_17681 , \4881_b1 );
not ( w_17681 , w_17684 );
not (  , w_17685 );
and ( w_17684 , w_17685 , \4881_b0 );
or ( \5577_b1 , \5575_b1 , w_17687 );
not ( w_17687 , w_17688 );
and ( \5577_b0 , \5575_b0 , w_17689 );
and ( w_17688 ,  , w_17689 );
buf ( w_17687 , \5576_b1 );
not ( w_17687 , w_17690 );
not (  , w_17691 );
and ( w_17690 , w_17691 , \5576_b0 );
or ( \5578_b1 , \5572_b1 , \5577_b1 );
not ( \5577_b1 , w_17692 );
and ( \5578_b0 , \5572_b0 , w_17693 );
and ( w_17692 , w_17693 , \5577_b0 );
or ( \5579_b1 , \5566_b1 , \5571_b1 );
not ( \5571_b1 , w_17694 );
and ( \5579_b0 , \5566_b0 , w_17695 );
and ( w_17694 , w_17695 , \5571_b0 );
or ( \5580_b1 , \5578_b1 , w_17696 );
or ( \5580_b0 , \5578_b0 , \5579_b0 );
not ( \5579_b0 , w_17697 );
and ( w_17697 , w_17696 , \5579_b1 );
buf ( \5581_b1 , \5580_b1 );
not ( \5581_b1 , w_17698 );
not ( \5581_b0 , w_17699 );
and ( w_17698 , w_17699 , \5580_b0 );
or ( \5582_b1 , \5309_b1 , \5320_b1 );
xor ( \5582_b0 , \5309_b0 , w_17700 );
not ( w_17700 , w_17701 );
and ( w_17701 , \5320_b1 , \5320_b0 );
or ( \5583_b1 , \5582_b1 , \5333_b1 );
xor ( \5583_b0 , \5582_b0 , w_17702 );
not ( w_17702 , w_17703 );
and ( w_17703 , \5333_b1 , \5333_b0 );
buf ( \5584_b1 , \5583_b1 );
not ( \5584_b1 , w_17704 );
not ( \5584_b0 , w_17705 );
and ( w_17704 , w_17705 , \5583_b0 );
or ( \5585_b1 , \5581_b1 , w_17706 );
or ( \5585_b0 , \5581_b0 , \5584_b0 );
not ( \5584_b0 , w_17707 );
and ( w_17707 , w_17706 , \5584_b1 );
or ( \5586_b1 , \5583_b1 , w_17708 );
or ( \5586_b0 , \5583_b0 , \5580_b0 );
not ( \5580_b0 , w_17709 );
and ( w_17709 , w_17708 , \5580_b1 );
or ( \5587_b1 , \4100_b1 , \4082_b1 );
not ( \4082_b1 , w_17710 );
and ( \5587_b0 , \4100_b0 , w_17711 );
and ( w_17710 , w_17711 , \4082_b0 );
buf ( \5588_b1 , \5587_b1 );
not ( \5588_b1 , w_17712 );
not ( \5588_b0 , w_17713 );
and ( w_17712 , w_17713 , \5587_b0 );
buf ( \5589_b1 , \5537_b1 );
not ( \5589_b1 , w_17714 );
not ( \5589_b0 , w_17715 );
and ( w_17714 , w_17715 , \5537_b0 );
buf ( \5590_b1 , \4395_b1 );
not ( \5590_b1 , w_17716 );
not ( \5590_b0 , w_17717 );
and ( w_17716 , w_17717 , \4395_b0 );
or ( \5591_b1 , \5589_b1 , w_17718 );
or ( \5591_b0 , \5589_b0 , \5590_b0 );
not ( \5590_b0 , w_17719 );
and ( w_17719 , w_17718 , \5590_b1 );
or ( \5592_b1 , \5286_b1 , w_17721 );
not ( w_17721 , w_17722 );
and ( \5592_b0 , \5286_b0 , w_17723 );
and ( w_17722 ,  , w_17723 );
buf ( w_17721 , \4200_b1 );
not ( w_17721 , w_17724 );
not (  , w_17725 );
and ( w_17724 , w_17725 , \4200_b0 );
or ( \5593_b1 , \5591_b1 , w_17727 );
not ( w_17727 , w_17728 );
and ( \5593_b0 , \5591_b0 , w_17729 );
and ( w_17728 ,  , w_17729 );
buf ( w_17727 , \5592_b1 );
not ( w_17727 , w_17730 );
not (  , w_17731 );
and ( w_17730 , w_17731 , \5592_b0 );
buf ( \5594_b1 , \5593_b1 );
not ( \5594_b1 , w_17732 );
not ( \5594_b0 , w_17733 );
and ( w_17732 , w_17733 , \5593_b0 );
or ( \5595_b1 , \5588_b1 , w_17734 );
or ( \5595_b0 , \5588_b0 , \5594_b0 );
not ( \5594_b0 , w_17735 );
and ( w_17735 , w_17734 , \5594_b1 );
or ( \5596_b1 , \5593_b1 , w_17736 );
or ( \5596_b0 , \5593_b0 , \5587_b0 );
not ( \5587_b0 , w_17737 );
and ( w_17737 , w_17736 , \5587_b1 );
buf ( \5597_b1 , \4449_b1 );
not ( \5597_b1 , w_17738 );
not ( \5597_b0 , w_17739 );
and ( w_17738 , w_17739 , \4449_b0 );
buf ( \5598_b1 , \5519_b1 );
not ( \5598_b1 , w_17740 );
not ( \5598_b0 , w_17741 );
and ( w_17740 , w_17741 , \5519_b0 );
or ( \5599_b1 , \5597_b1 , w_17742 );
or ( \5599_b0 , \5597_b0 , \5598_b0 );
not ( \5598_b0 , w_17743 );
and ( w_17743 , w_17742 , \5598_b1 );
or ( \5600_b1 , \4452_b1 , w_17745 );
not ( w_17745 , w_17746 );
and ( \5600_b0 , \4452_b0 , w_17747 );
and ( w_17746 ,  , w_17747 );
buf ( w_17745 , \5116_b1 );
not ( w_17745 , w_17748 );
not (  , w_17749 );
and ( w_17748 , w_17749 , \5116_b0 );
or ( \5601_b1 , \5599_b1 , w_17751 );
not ( w_17751 , w_17752 );
and ( \5601_b0 , \5599_b0 , w_17753 );
and ( w_17752 ,  , w_17753 );
buf ( w_17751 , \5600_b1 );
not ( w_17751 , w_17754 );
not (  , w_17755 );
and ( w_17754 , w_17755 , \5600_b0 );
or ( \5602_b1 , \5596_b1 , w_17757 );
not ( w_17757 , w_17758 );
and ( \5602_b0 , \5596_b0 , w_17759 );
and ( w_17758 ,  , w_17759 );
buf ( w_17757 , \5601_b1 );
not ( w_17757 , w_17760 );
not (  , w_17761 );
and ( w_17760 , w_17761 , \5601_b0 );
or ( \5603_b1 , \5595_b1 , w_17763 );
not ( w_17763 , w_17764 );
and ( \5603_b0 , \5595_b0 , w_17765 );
and ( w_17764 ,  , w_17765 );
buf ( w_17763 , \5602_b1 );
not ( w_17763 , w_17766 );
not (  , w_17767 );
and ( w_17766 , w_17767 , \5602_b0 );
or ( \5604_b1 , \5586_b1 , w_17769 );
not ( w_17769 , w_17770 );
and ( \5604_b0 , \5586_b0 , w_17771 );
and ( w_17770 ,  , w_17771 );
buf ( w_17769 , \5603_b1 );
not ( w_17769 , w_17772 );
not (  , w_17773 );
and ( w_17772 , w_17773 , \5603_b0 );
or ( \5605_b1 , \5585_b1 , w_17775 );
not ( w_17775 , w_17776 );
and ( \5605_b0 , \5585_b0 , w_17777 );
and ( w_17776 ,  , w_17777 );
buf ( w_17775 , \5604_b1 );
not ( w_17775 , w_17778 );
not (  , w_17779 );
and ( w_17778 , w_17779 , \5604_b0 );
buf ( \5606_b1 , \5605_b1 );
not ( \5606_b1 , w_17780 );
not ( \5606_b0 , w_17781 );
and ( w_17780 , w_17781 , \5605_b0 );
or ( \5607_b1 , \5561_b1 , w_17783 );
not ( w_17783 , w_17784 );
and ( \5607_b0 , \5561_b0 , w_17785 );
and ( w_17784 ,  , w_17785 );
buf ( w_17783 , \5606_b1 );
not ( w_17783 , w_17786 );
not (  , w_17787 );
and ( w_17786 , w_17787 , \5606_b0 );
buf ( \5608_b1 , \5607_b1 );
not ( \5608_b1 , w_17788 );
not ( \5608_b0 , w_17789 );
and ( w_17788 , w_17789 , \5607_b0 );
or ( \5609_b1 , \5551_b1 , w_17790 );
or ( \5609_b0 , \5551_b0 , \5608_b0 );
not ( \5608_b0 , w_17791 );
and ( w_17791 , w_17790 , \5608_b1 );
buf ( \5610_b1 , \5561_b1 );
not ( \5610_b1 , w_17792 );
not ( \5610_b0 , w_17793 );
and ( w_17792 , w_17793 , \5561_b0 );
or ( \5611_b1 , \5610_b1 , w_17795 );
not ( w_17795 , w_17796 );
and ( \5611_b0 , \5610_b0 , w_17797 );
and ( w_17796 ,  , w_17797 );
buf ( w_17795 , \5605_b1 );
not ( w_17795 , w_17798 );
not (  , w_17799 );
and ( w_17798 , w_17799 , \5605_b0 );
or ( \5612_b1 , \5609_b1 , w_17801 );
not ( w_17801 , w_17802 );
and ( \5612_b0 , \5609_b0 , w_17803 );
and ( w_17802 ,  , w_17803 );
buf ( w_17801 , \5611_b1 );
not ( w_17801 , w_17804 );
not (  , w_17805 );
and ( w_17804 , w_17805 , \5611_b0 );
buf ( \5613_b1 , \5612_b1 );
buf ( \5613_b0 , \5612_b0 );
or ( \5614_b1 , \5371_b1 , \5613_b1 );
not ( \5613_b1 , w_17806 );
and ( \5614_b0 , \5371_b0 , w_17807 );
and ( w_17806 , w_17807 , \5613_b0 );
buf ( \5615_b1 , \5369_b1 );
not ( \5615_b1 , w_17808 );
not ( \5615_b0 , w_17809 );
and ( w_17808 , w_17809 , \5369_b0 );
or ( \5616_b1 , \5357_b1 , w_17811 );
not ( w_17811 , w_17812 );
and ( \5616_b0 , \5357_b0 , w_17813 );
and ( w_17812 ,  , w_17813 );
buf ( w_17811 , \5615_b1 );
not ( w_17811 , w_17814 );
not (  , w_17815 );
and ( w_17814 , w_17815 , \5615_b0 );
or ( \5617_b1 , \5614_b1 , w_17817 );
not ( w_17817 , w_17818 );
and ( \5617_b0 , \5614_b0 , w_17819 );
and ( w_17818 ,  , w_17819 );
buf ( w_17817 , \5616_b1 );
not ( w_17817 , w_17820 );
not (  , w_17821 );
and ( w_17820 , w_17821 , \5616_b0 );
or ( \5618_b1 , \5354_b1 , w_17823 );
not ( w_17823 , w_17824 );
and ( \5618_b0 , \5354_b0 , w_17825 );
and ( w_17824 ,  , w_17825 );
buf ( w_17823 , \5617_b1 );
not ( w_17823 , w_17826 );
not (  , w_17827 );
and ( w_17826 , w_17827 , \5617_b0 );
or ( \5619_b1 , \5130_b1 , \5219_b1 );
xor ( \5619_b0 , \5130_b0 , w_17828 );
not ( w_17828 , w_17829 );
and ( w_17829 , \5219_b1 , \5219_b0 );
or ( \5620_b1 , \5619_b1 , \5353_b1 );
not ( \5353_b1 , w_17830 );
and ( \5620_b0 , \5619_b0 , w_17831 );
and ( w_17830 , w_17831 , \5353_b0 );
or ( \5621_b1 , \5130_b1 , \5219_b1 );
not ( \5219_b1 , w_17832 );
and ( \5621_b0 , \5130_b0 , w_17833 );
and ( w_17832 , w_17833 , \5219_b0 );
or ( \5622_b1 , \5620_b1 , w_17834 );
or ( \5622_b0 , \5620_b0 , \5621_b0 );
not ( \5621_b0 , w_17835 );
and ( w_17835 , w_17834 , \5621_b1 );
buf ( \5623_b1 , \4807_b1 );
not ( \5623_b1 , w_17836 );
not ( \5623_b0 , w_17837 );
and ( w_17836 , w_17837 , \4807_b0 );
buf ( \5624_b1 , \4773_b1 );
not ( \5624_b1 , w_17838 );
not ( \5624_b0 , w_17839 );
and ( w_17838 , w_17839 , \4773_b0 );
or ( \5625_b1 , \5623_b1 , w_17840 );
or ( \5625_b0 , \5623_b0 , \5624_b0 );
not ( \5624_b0 , w_17841 );
and ( w_17841 , w_17840 , \5624_b1 );
or ( \5626_b1 , \4804_b1 , w_17843 );
not ( w_17843 , w_17844 );
and ( \5626_b0 , \4804_b0 , w_17845 );
and ( w_17844 ,  , w_17845 );
buf ( w_17843 , \4772_b1 );
not ( w_17843 , w_17846 );
not (  , w_17847 );
and ( w_17846 , w_17847 , \4772_b0 );
or ( \5627_b1 , \5625_b1 , w_17849 );
not ( w_17849 , w_17850 );
and ( \5627_b0 , \5625_b0 , w_17851 );
and ( w_17850 ,  , w_17851 );
buf ( w_17849 , \5626_b1 );
not ( w_17849 , w_17852 );
not (  , w_17853 );
and ( w_17852 , w_17853 , \5626_b0 );
buf ( \5628_b1 , \4812_b1 );
not ( \5628_b1 , w_17854 );
not ( \5628_b0 , w_17855 );
and ( w_17854 , w_17855 , \4812_b0 );
or ( \5629_b1 , \5627_b1 , \5628_b1 );
not ( \5628_b1 , w_17856 );
and ( \5629_b0 , \5627_b0 , w_17857 );
and ( w_17856 , w_17857 , \5628_b0 );
buf ( \5630_b1 , \5627_b1 );
not ( \5630_b1 , w_17858 );
not ( \5630_b0 , w_17859 );
and ( w_17858 , w_17859 , \5627_b0 );
or ( \5631_b1 , \5630_b1 , \4812_b1 );
not ( \4812_b1 , w_17860 );
and ( \5631_b0 , \5630_b0 , w_17861 );
and ( w_17860 , w_17861 , \4812_b0 );
or ( \5632_b1 , \5629_b1 , w_17863 );
not ( w_17863 , w_17864 );
and ( \5632_b0 , \5629_b0 , w_17865 );
and ( w_17864 ,  , w_17865 );
buf ( w_17863 , \5631_b1 );
not ( w_17863 , w_17866 );
not (  , w_17867 );
and ( w_17866 , w_17867 , \5631_b0 );
or ( \5633_b1 , \4847_b1 , \4930_b1 );
xor ( \5633_b0 , \4847_b0 , w_17868 );
not ( w_17868 , w_17869 );
and ( w_17869 , \4930_b1 , \4930_b0 );
or ( \5634_b1 , \5633_b1 , w_17870 );
xor ( \5634_b0 , \5633_b0 , w_17872 );
not ( w_17872 , w_17873 );
and ( w_17873 , w_17870 , w_17871 );
buf ( w_17870 , \4999_b1 );
not ( w_17870 , w_17874 );
not ( w_17871 , w_17875 );
and ( w_17874 , w_17875 , \4999_b0 );
or ( \5635_b1 , \5632_b1 , \5634_b1 );
xor ( \5635_b0 , \5632_b0 , w_17876 );
not ( w_17876 , w_17877 );
and ( w_17877 , \5634_b1 , \5634_b0 );
or ( \5636_b1 , \5132_b1 , \5207_b1 );
xor ( \5636_b0 , \5132_b0 , w_17878 );
not ( w_17878 , w_17879 );
and ( w_17879 , \5207_b1 , \5207_b0 );
or ( \5637_b1 , \5636_b1 , \5218_b1 );
not ( \5218_b1 , w_17880 );
and ( \5637_b0 , \5636_b0 , w_17881 );
and ( w_17880 , w_17881 , \5218_b0 );
or ( \5638_b1 , \5132_b1 , \5207_b1 );
not ( \5207_b1 , w_17882 );
and ( \5638_b0 , \5132_b0 , w_17883 );
and ( w_17882 , w_17883 , \5207_b0 );
or ( \5639_b1 , \5637_b1 , w_17884 );
or ( \5639_b0 , \5637_b0 , \5638_b0 );
not ( \5638_b0 , w_17885 );
and ( w_17885 , w_17884 , \5638_b1 );
or ( \5640_b1 , \5635_b1 , \5639_b1 );
xor ( \5640_b0 , \5635_b0 , w_17886 );
not ( w_17886 , w_17887 );
and ( w_17887 , \5639_b1 , \5639_b0 );
or ( \5641_b1 , \5622_b1 , w_17889 );
not ( w_17889 , w_17890 );
and ( \5641_b0 , \5622_b0 , w_17891 );
and ( w_17890 ,  , w_17891 );
buf ( w_17889 , \5640_b1 );
not ( w_17889 , w_17892 );
not (  , w_17893 );
and ( w_17892 , w_17893 , \5640_b0 );
or ( \5642_b1 , \5632_b1 , \5634_b1 );
xor ( \5642_b0 , \5632_b0 , w_17894 );
not ( w_17894 , w_17895 );
and ( w_17895 , \5634_b1 , \5634_b0 );
or ( \5643_b1 , \5642_b1 , \5639_b1 );
not ( \5639_b1 , w_17896 );
and ( \5643_b0 , \5642_b0 , w_17897 );
and ( w_17896 , w_17897 , \5639_b0 );
or ( \5644_b1 , \5632_b1 , \5634_b1 );
not ( \5634_b1 , w_17898 );
and ( \5644_b0 , \5632_b0 , w_17899 );
and ( w_17898 , w_17899 , \5634_b0 );
or ( \5645_b1 , \5643_b1 , w_17900 );
or ( \5645_b0 , \5643_b0 , \5644_b0 );
not ( \5644_b0 , w_17901 );
and ( w_17901 , w_17900 , \5644_b1 );
or ( \5646_b1 , \4837_b1 , \5001_b1 );
xor ( \5646_b0 , \4837_b0 , w_17902 );
not ( w_17902 , w_17903 );
and ( w_17903 , \5001_b1 , \5001_b0 );
or ( \5647_b1 , \5646_b1 , w_17904 );
xor ( \5647_b0 , \5646_b0 , w_17906 );
not ( w_17906 , w_17907 );
and ( w_17907 , w_17904 , w_17905 );
buf ( w_17904 , \4834_b1 );
not ( w_17904 , w_17908 );
not ( w_17905 , w_17909 );
and ( w_17908 , w_17909 , \4834_b0 );
or ( \5648_b1 , \5645_b1 , w_17911 );
not ( w_17911 , w_17912 );
and ( \5648_b0 , \5645_b0 , w_17913 );
and ( w_17912 ,  , w_17913 );
buf ( w_17911 , \5647_b1 );
not ( w_17911 , w_17914 );
not (  , w_17915 );
and ( w_17914 , w_17915 , \5647_b0 );
or ( \5650_b1 , \5368_b1 , \5612_b1 );
xor ( \5650_b0 , \5368_b0 , w_17916 );
not ( w_17916 , w_17917 );
and ( w_17917 , \5612_b1 , \5612_b0 );
or ( \5651_b1 , \5650_b1 , w_17918 );
xor ( \5651_b0 , \5650_b0 , w_17920 );
not ( w_17920 , w_17921 );
and ( w_17921 , w_17918 , w_17919 );
buf ( w_17918 , \5356_b1 );
not ( w_17918 , w_17922 );
not ( w_17919 , w_17923 );
and ( w_17922 , w_17923 , \5356_b0 );
or ( \5652_b1 , \5239_b1 , \5232_b1 );
xor ( \5652_b0 , \5239_b0 , w_17924 );
not ( w_17924 , w_17925 );
and ( w_17925 , \5232_b1 , \5232_b0 );
or ( \5653_b1 , \5652_b1 , w_17926 );
xor ( \5653_b0 , \5652_b0 , w_17928 );
not ( w_17928 , w_17929 );
and ( w_17929 , w_17926 , w_17927 );
buf ( w_17926 , \5259_b1 );
not ( w_17926 , w_17930 );
not ( w_17927 , w_17931 );
and ( w_17930 , w_17931 , \5259_b0 );
or ( \5654_b1 , \5580_b1 , \5603_b1 );
xor ( \5654_b0 , \5580_b0 , w_17932 );
not ( w_17932 , w_17933 );
and ( w_17933 , \5603_b1 , \5603_b0 );
or ( \5655_b1 , \5654_b1 , w_17934 );
xor ( \5655_b0 , \5654_b0 , w_17936 );
not ( w_17936 , w_17937 );
and ( w_17937 , w_17934 , w_17935 );
buf ( w_17934 , \5583_b1 );
not ( w_17934 , w_17938 );
not ( w_17935 , w_17939 );
and ( w_17938 , w_17939 , \5583_b0 );
buf ( \5656_b1 , \5248_b1 );
not ( \5656_b1 , w_17940 );
not ( \5656_b0 , w_17941 );
and ( w_17940 , w_17941 , \5248_b0 );
buf ( \5657_b1 , \5258_b1 );
not ( \5657_b1 , w_17942 );
not ( \5657_b0 , w_17943 );
and ( w_17942 , w_17943 , \5258_b0 );
buf ( \5658_b1 , \5657_b1 );
not ( \5658_b1 , w_17944 );
not ( \5658_b0 , w_17945 );
and ( w_17944 , w_17945 , \5657_b0 );
or ( \5659_b1 , \5656_b1 , \5658_b1 );
not ( \5658_b1 , w_17946 );
and ( \5659_b0 , \5656_b0 , w_17947 );
and ( w_17946 , w_17947 , \5658_b0 );
or ( \5660_b1 , \5248_b1 , \5657_b1 );
not ( \5657_b1 , w_17948 );
and ( \5660_b0 , \5248_b0 , w_17949 );
and ( w_17948 , w_17949 , \5657_b0 );
or ( \5661_b1 , \5659_b1 , w_17951 );
not ( w_17951 , w_17952 );
and ( \5661_b0 , \5659_b0 , w_17953 );
and ( w_17952 ,  , w_17953 );
buf ( w_17951 , \5660_b1 );
not ( w_17951 , w_17954 );
not (  , w_17955 );
and ( w_17954 , w_17955 , \5660_b0 );
buf ( \5662_b1 , \5661_b1 );
buf ( \5662_b0 , \5661_b0 );
or ( \5663_b1 , \5655_b1 , w_17957 );
not ( w_17957 , w_17958 );
and ( \5663_b0 , \5655_b0 , w_17959 );
and ( w_17958 ,  , w_17959 );
buf ( w_17957 , \5662_b1 );
not ( w_17957 , w_17960 );
not (  , w_17961 );
and ( w_17960 , w_17961 , \5662_b0 );
or ( \5664_b1 , \5566_b1 , \5571_b1 );
xor ( \5664_b0 , \5566_b0 , w_17962 );
not ( w_17962 , w_17963 );
and ( w_17963 , \5571_b1 , \5571_b0 );
or ( \5665_b1 , \5664_b1 , \5577_b1 );
xor ( \5665_b0 , \5664_b0 , w_17964 );
not ( w_17964 , w_17965 );
and ( w_17965 , \5577_b1 , \5577_b0 );
buf ( \5666_b1 , \5665_b1 );
not ( \5666_b1 , w_17966 );
not ( \5666_b0 , w_17967 );
and ( w_17966 , w_17967 , \5665_b0 );
or ( \5667_b1 , \5587_b1 , \5601_b1 );
xor ( \5667_b0 , \5587_b0 , w_17968 );
not ( w_17968 , w_17969 );
and ( w_17969 , \5601_b1 , \5601_b0 );
or ( \5668_b1 , \5667_b1 , w_17970 );
xor ( \5668_b0 , \5667_b0 , w_17972 );
not ( w_17972 , w_17973 );
and ( w_17973 , w_17970 , w_17971 );
buf ( w_17970 , \5593_b1 );
not ( w_17970 , w_17974 );
not ( w_17971 , w_17975 );
and ( w_17974 , w_17975 , \5593_b0 );
buf ( \5669_b1 , \5668_b1 );
not ( \5669_b1 , w_17976 );
not ( \5669_b0 , w_17977 );
and ( w_17976 , w_17977 , \5668_b0 );
buf ( \5670_b1 , \5669_b1 );
not ( \5670_b1 , w_17978 );
not ( \5670_b0 , w_17979 );
and ( w_17978 , w_17979 , \5669_b0 );
or ( \5671_b1 , \5666_b1 , w_17980 );
or ( \5671_b0 , \5666_b0 , \5670_b0 );
not ( \5670_b0 , w_17981 );
and ( w_17981 , w_17980 , \5670_b1 );
buf ( \5672_b1 , \5668_b1 );
not ( \5672_b1 , w_17982 );
not ( \5672_b0 , w_17983 );
and ( w_17982 , w_17983 , \5668_b0 );
buf ( \5673_b1 , \5665_b1 );
not ( \5673_b1 , w_17984 );
not ( \5673_b0 , w_17985 );
and ( w_17984 , w_17985 , \5665_b0 );
buf ( \5674_b1 , \5673_b1 );
not ( \5674_b1 , w_17986 );
not ( \5674_b0 , w_17987 );
and ( w_17986 , w_17987 , \5673_b0 );
or ( \5675_b1 , \5672_b1 , w_17988 );
or ( \5675_b0 , \5672_b0 , \5674_b0 );
not ( \5674_b0 , w_17989 );
and ( w_17989 , w_17988 , \5674_b1 );
buf ( \5676_b1 , \5397_b1 );
not ( \5676_b1 , w_17990 );
not ( \5676_b0 , w_17991 );
and ( w_17990 , w_17991 , \5397_b0 );
buf ( \5677_b1 , \5392_b1 );
not ( \5677_b1 , w_17992 );
not ( \5677_b0 , w_17993 );
and ( w_17992 , w_17993 , \5392_b0 );
or ( \5678_b1 , \5676_b1 , w_17994 );
or ( \5678_b0 , \5676_b0 , \5677_b0 );
not ( \5677_b0 , w_17995 );
and ( w_17995 , w_17994 , \5677_b1 );
or ( \5679_b1 , \5397_b1 , w_17996 );
or ( \5679_b0 , \5397_b0 , \5392_b0 );
not ( \5392_b0 , w_17997 );
and ( w_17997 , w_17996 , \5392_b1 );
or ( \5680_b1 , \5678_b1 , w_17999 );
not ( w_17999 , w_18000 );
and ( \5680_b0 , \5678_b0 , w_18001 );
and ( w_18000 ,  , w_18001 );
buf ( w_17999 , \5679_b1 );
not ( w_17999 , w_18002 );
not (  , w_18003 );
and ( w_18002 , w_18003 , \5679_b0 );
buf ( \5681_b1 , \5410_b1 );
not ( \5681_b1 , w_18004 );
not ( \5681_b0 , w_18005 );
and ( w_18004 , w_18005 , \5410_b0 );
or ( \5682_b1 , \5680_b1 , \5681_b1 );
not ( \5681_b1 , w_18006 );
and ( \5682_b0 , \5680_b0 , w_18007 );
and ( w_18006 , w_18007 , \5681_b0 );
buf ( \5683_b1 , \5680_b1 );
not ( \5683_b1 , w_18008 );
not ( \5683_b0 , w_18009 );
and ( w_18008 , w_18009 , \5680_b0 );
or ( \5684_b1 , \5683_b1 , \5410_b1 );
not ( \5410_b1 , w_18010 );
and ( \5684_b0 , \5683_b0 , w_18011 );
and ( w_18010 , w_18011 , \5410_b0 );
or ( \5685_b1 , \5682_b1 , w_18013 );
not ( w_18013 , w_18014 );
and ( \5685_b0 , \5682_b0 , w_18015 );
and ( w_18014 ,  , w_18015 );
buf ( w_18013 , \5684_b1 );
not ( w_18013 , w_18016 );
not (  , w_18017 );
and ( w_18016 , w_18017 , \5684_b0 );
buf ( \5686_b1 , \5685_b1 );
not ( \5686_b1 , w_18018 );
not ( \5686_b0 , w_18019 );
and ( w_18018 , w_18019 , \5685_b0 );
or ( \5687_b1 , \5675_b1 , w_18021 );
not ( w_18021 , w_18022 );
and ( \5687_b0 , \5675_b0 , w_18023 );
and ( w_18022 ,  , w_18023 );
buf ( w_18021 , \5686_b1 );
not ( w_18021 , w_18024 );
not (  , w_18025 );
and ( w_18024 , w_18025 , \5686_b0 );
or ( \5688_b1 , \5671_b1 , w_18027 );
not ( w_18027 , w_18028 );
and ( \5688_b0 , \5671_b0 , w_18029 );
and ( w_18028 ,  , w_18029 );
buf ( w_18027 , \5687_b1 );
not ( w_18027 , w_18030 );
not (  , w_18031 );
and ( w_18030 , w_18031 , \5687_b0 );
or ( \5689_b1 , \5663_b1 , \5688_b1 );
not ( \5688_b1 , w_18032 );
and ( \5689_b0 , \5663_b0 , w_18033 );
and ( w_18032 , w_18033 , \5688_b0 );
or ( \5690_b1 , \5655_b1 , w_18035 );
not ( w_18035 , w_18036 );
and ( \5690_b0 , \5655_b0 , w_18037 );
and ( w_18036 ,  , w_18037 );
buf ( w_18035 , \5662_b1 );
not ( w_18035 , w_18038 );
not (  , w_18039 );
and ( w_18038 , w_18039 , \5662_b0 );
or ( \5691_b1 , \5689_b1 , w_18041 );
not ( w_18041 , w_18042 );
and ( \5691_b0 , \5689_b0 , w_18043 );
and ( w_18042 ,  , w_18043 );
buf ( w_18041 , \5690_b1 );
not ( w_18041 , w_18044 );
not (  , w_18045 );
and ( w_18044 , w_18045 , \5690_b0 );
or ( \5692_b1 , \5653_b1 , \5691_b1 );
xor ( \5692_b0 , \5653_b0 , w_18046 );
not ( w_18046 , w_18047 );
and ( w_18047 , \5691_b1 , \5691_b0 );
buf ( \5693_b1 , \5605_b1 );
not ( \5693_b1 , w_18048 );
not ( \5693_b0 , w_18049 );
and ( w_18048 , w_18049 , \5605_b0 );
buf ( \5694_b1 , \5561_b1 );
not ( \5694_b1 , w_18050 );
not ( \5694_b0 , w_18051 );
and ( w_18050 , w_18051 , \5561_b0 );
or ( \5695_b1 , \5693_b1 , w_18052 );
or ( \5695_b0 , \5693_b0 , \5694_b0 );
not ( \5694_b0 , w_18053 );
and ( w_18053 , w_18052 , \5694_b1 );
or ( \5696_b1 , \5606_b1 , w_18055 );
not ( w_18055 , w_18056 );
and ( \5696_b0 , \5606_b0 , w_18057 );
and ( w_18056 ,  , w_18057 );
buf ( w_18055 , \5560_b1 );
not ( w_18055 , w_18058 );
not (  , w_18059 );
and ( w_18058 , w_18059 , \5560_b0 );
or ( \5697_b1 , \5695_b1 , w_18061 );
not ( w_18061 , w_18062 );
and ( \5697_b0 , \5695_b0 , w_18063 );
and ( w_18062 ,  , w_18063 );
buf ( w_18061 , \5696_b1 );
not ( w_18061 , w_18064 );
not (  , w_18065 );
and ( w_18064 , w_18065 , \5696_b0 );
buf ( \5698_b1 , \5550_b1 );
not ( \5698_b1 , w_18066 );
not ( \5698_b0 , w_18067 );
and ( w_18066 , w_18067 , \5550_b0 );
or ( \5699_b1 , \5697_b1 , \5698_b1 );
not ( \5698_b1 , w_18068 );
and ( \5699_b0 , \5697_b0 , w_18069 );
and ( w_18068 , w_18069 , \5698_b0 );
buf ( \5700_b1 , \5697_b1 );
not ( \5700_b1 , w_18070 );
not ( \5700_b0 , w_18071 );
and ( w_18070 , w_18071 , \5697_b0 );
or ( \5701_b1 , \5700_b1 , \5550_b1 );
not ( \5550_b1 , w_18072 );
and ( \5701_b0 , \5700_b0 , w_18073 );
and ( w_18072 , w_18073 , \5550_b0 );
or ( \5702_b1 , \5699_b1 , w_18075 );
not ( w_18075 , w_18076 );
and ( \5702_b0 , \5699_b0 , w_18077 );
and ( w_18076 ,  , w_18077 );
buf ( w_18075 , \5701_b1 );
not ( w_18075 , w_18078 );
not (  , w_18079 );
and ( w_18078 , w_18079 , \5701_b0 );
or ( \5703_b1 , \5692_b1 , \5702_b1 );
not ( \5702_b1 , w_18080 );
and ( \5703_b0 , \5692_b0 , w_18081 );
and ( w_18080 , w_18081 , \5702_b0 );
or ( \5704_b1 , \5653_b1 , \5691_b1 );
not ( \5691_b1 , w_18082 );
and ( \5704_b0 , \5653_b0 , w_18083 );
and ( w_18082 , w_18083 , \5691_b0 );
or ( \5705_b1 , \5703_b1 , w_18084 );
or ( \5705_b0 , \5703_b0 , \5704_b0 );
not ( \5704_b0 , w_18085 );
and ( w_18085 , w_18084 , \5704_b1 );
or ( \5706_b1 , \5651_b1 , w_18087 );
not ( w_18087 , w_18088 );
and ( \5706_b0 , \5651_b0 , w_18089 );
and ( w_18088 ,  , w_18089 );
buf ( w_18087 , \5705_b1 );
not ( w_18087 , w_18090 );
not (  , w_18091 );
and ( w_18090 , w_18091 , \5705_b0 );
or ( \5707_b1 , \5649_b1 , \5706_b1 );
not ( \5706_b1 , w_18092 );
and ( \5707_b0 , \5649_b0 , w_18093 );
and ( w_18092 , w_18093 , \5706_b0 );
buf ( \5708_b1 , \5655_b1 );
not ( \5708_b1 , w_18094 );
not ( \5708_b0 , w_18095 );
and ( w_18094 , w_18095 , \5655_b0 );
buf ( \5709_b1 , \5661_b1 );
not ( \5709_b1 , w_18096 );
not ( \5709_b0 , w_18097 );
and ( w_18096 , w_18097 , \5661_b0 );
buf ( \5710_b1 , \5688_b1 );
not ( \5710_b1 , w_18098 );
not ( \5710_b0 , w_18099 );
and ( w_18098 , w_18099 , \5688_b0 );
or ( \5711_b1 , \5709_b1 , w_18100 );
or ( \5711_b0 , \5709_b0 , \5710_b0 );
not ( \5710_b0 , w_18101 );
and ( w_18101 , w_18100 , \5710_b1 );
or ( \5712_b1 , \5661_b1 , w_18102 );
or ( \5712_b0 , \5661_b0 , \5688_b0 );
not ( \5688_b0 , w_18103 );
and ( w_18103 , w_18102 , \5688_b1 );
or ( \5713_b1 , \5711_b1 , w_18105 );
not ( w_18105 , w_18106 );
and ( \5713_b0 , \5711_b0 , w_18107 );
and ( w_18106 ,  , w_18107 );
buf ( w_18105 , \5712_b1 );
not ( w_18105 , w_18108 );
not (  , w_18109 );
and ( w_18108 , w_18109 , \5712_b0 );
buf ( \5714_b1 , \5713_b1 );
not ( \5714_b1 , w_18110 );
not ( \5714_b0 , w_18111 );
and ( w_18110 , w_18111 , \5713_b0 );
or ( \5715_b1 , \5708_b1 , w_18112 );
or ( \5715_b0 , \5708_b0 , \5714_b0 );
not ( \5714_b0 , w_18113 );
and ( w_18113 , w_18112 , \5714_b1 );
or ( \5716_b1 , \5655_b1 , w_18114 );
or ( \5716_b0 , \5655_b0 , \5713_b0 );
not ( \5713_b0 , w_18115 );
and ( w_18115 , w_18114 , \5713_b1 );
or ( \5717_b1 , \5715_b1 , w_18117 );
not ( w_18117 , w_18118 );
and ( \5717_b0 , \5715_b0 , w_18119 );
and ( w_18118 ,  , w_18119 );
buf ( w_18117 , \5716_b1 );
not ( w_18117 , w_18120 );
not (  , w_18121 );
and ( w_18120 , w_18121 , \5716_b0 );
buf ( \5718_b1 , \5717_b1 );
not ( \5718_b1 , w_18122 );
not ( \5718_b0 , w_18123 );
and ( w_18122 , w_18123 , \5717_b0 );
buf ( \5719_b1 , \5718_b1 );
not ( \5719_b1 , w_18124 );
not ( \5719_b0 , w_18125 );
and ( w_18124 , w_18125 , \5718_b0 );
or ( \5720_b1 , \5412_b1 , \5415_b1 );
xor ( \5720_b0 , \5412_b0 , w_18126 );
not ( w_18126 , w_18127 );
and ( w_18127 , \5415_b1 , \5415_b0 );
or ( \5721_b1 , \5720_b1 , w_18128 );
xor ( \5721_b0 , \5720_b0 , w_18130 );
not ( w_18130 , w_18131 );
and ( w_18131 , w_18128 , w_18129 );
buf ( w_18128 , \5545_b1 );
not ( w_18128 , w_18132 );
not ( w_18129 , w_18133 );
and ( w_18132 , w_18133 , \5545_b0 );
buf ( \5722_b1 , \5721_b1 );
not ( \5722_b1 , w_18134 );
not ( \5722_b0 , w_18135 );
and ( w_18134 , w_18135 , \5721_b0 );
or ( \5723_b1 , \5448_b1 , \5489_b1 );
xor ( \5723_b0 , \5448_b0 , w_18136 );
not ( w_18136 , w_18137 );
and ( w_18137 , \5489_b1 , \5489_b0 );
or ( \5724_b1 , \5723_b1 , \5542_b1 );
xor ( \5724_b0 , \5723_b0 , w_18138 );
not ( w_18138 , w_18139 );
and ( w_18139 , \5542_b1 , \5542_b0 );
buf ( \5725_b1 , \5724_b1 );
not ( \5725_b1 , w_18140 );
not ( \5725_b0 , w_18141 );
and ( w_18140 , w_18141 , \5724_b0 );
buf ( \5726_b1 , \5418_b1 );
not ( \5726_b1 , w_18142 );
not ( \5726_b0 , w_18143 );
and ( w_18142 , w_18143 , \5418_b0 );
buf ( \5727_b1 , \4182_b1 );
not ( \5727_b1 , w_18144 );
not ( \5727_b0 , w_18145 );
and ( w_18144 , w_18145 , \4182_b0 );
or ( \5728_b1 , \5726_b1 , w_18146 );
or ( \5728_b0 , \5726_b0 , \5727_b0 );
not ( \5727_b0 , w_18147 );
and ( w_18147 , w_18146 , \5727_b1 );
or ( \5729_b1 , \5728_b1 , w_18149 );
not ( w_18149 , w_18150 );
and ( \5729_b0 , \5728_b0 , w_18151 );
and ( w_18150 ,  , w_18151 );
buf ( w_18149 , \4110_b1 );
not ( w_18149 , w_18152 );
not (  , w_18153 );
and ( w_18152 , w_18153 , \4110_b0 );
buf ( \5730_b1 , \4182_b1 );
not ( \5730_b1 , w_18154 );
not ( \5730_b0 , w_18155 );
and ( w_18154 , w_18155 , \4182_b0 );
or ( \5731_b1 , \5730_b1 , w_18157 );
not ( w_18157 , w_18158 );
and ( \5731_b0 , \5730_b0 , w_18159 );
and ( w_18158 ,  , w_18159 );
buf ( w_18157 , \4098_b1 );
not ( w_18157 , w_18160 );
not (  , w_18161 );
and ( w_18160 , w_18161 , \4098_b0 );
buf ( \5733_b1 , \4096_b1 );
not ( \5733_b1 , w_18162 );
not ( \5733_b0 , w_18163 );
and ( w_18162 , w_18163 , \4096_b0 );
buf ( \5734_b1 , \4935_b1 );
not ( \5734_b1 , w_18164 );
not ( \5734_b0 , w_18165 );
and ( w_18164 , w_18165 , \4935_b0 );
or ( \5735_b1 , \5733_b1 , w_18166 );
or ( \5735_b0 , \5733_b0 , \5734_b0 );
not ( \5734_b0 , w_18167 );
and ( w_18167 , w_18166 , \5734_b1 );
or ( \5736_b1 , \2945_b1 , w_18169 );
not ( w_18169 , w_18170 );
and ( \5736_b0 , \2945_b0 , w_18171 );
and ( w_18170 ,  , w_18171 );
buf ( w_18169 , \4372_b1 );
not ( w_18169 , w_18172 );
not (  , w_18173 );
and ( w_18172 , w_18173 , \4372_b0 );
or ( \5737_b1 , \5735_b1 , w_18175 );
not ( w_18175 , w_18176 );
and ( \5737_b0 , \5735_b0 , w_18177 );
and ( w_18176 ,  , w_18177 );
buf ( w_18175 , \5736_b1 );
not ( w_18175 , w_18178 );
not (  , w_18179 );
and ( w_18178 , w_18179 , \5736_b0 );
buf ( \5738_b1 , \5737_b1 );
not ( \5738_b1 , w_18180 );
not ( \5738_b0 , w_18181 );
and ( w_18180 , w_18181 , \5737_b0 );
buf ( \5739_b1 , \4944_b1 );
not ( \5739_b1 , w_18182 );
not ( \5739_b0 , w_18183 );
and ( w_18182 , w_18183 , \4944_b0 );
or ( \5740_b1 , \5738_b1 , w_18184 );
or ( \5740_b0 , \5738_b0 , \5739_b0 );
not ( \5739_b0 , w_18185 );
and ( w_18185 , w_18184 , \5739_b1 );
buf ( \5741_b1 , \5441_b1 );
not ( \5741_b1 , w_18186 );
not ( \5741_b0 , w_18187 );
and ( w_18186 , w_18187 , \5441_b0 );
or ( \5742_b1 , \5741_b1 , w_18189 );
not ( w_18189 , w_18190 );
and ( \5742_b0 , \5741_b0 , w_18191 );
and ( w_18190 ,  , w_18191 );
buf ( w_18189 , \4863_b1 );
not ( w_18189 , w_18192 );
not (  , w_18193 );
and ( w_18192 , w_18193 , \4863_b0 );
or ( \5743_b1 , \5740_b1 , w_18195 );
not ( w_18195 , w_18196 );
and ( \5743_b0 , \5740_b0 , w_18197 );
and ( w_18196 ,  , w_18197 );
buf ( w_18195 , \5742_b1 );
not ( w_18195 , w_18198 );
not (  , w_18199 );
and ( w_18198 , w_18199 , \5742_b0 );
buf ( \5744_b1 , \5743_b1 );
not ( \5744_b1 , w_18200 );
not ( \5744_b0 , w_18201 );
and ( w_18200 , w_18201 , \5743_b0 );
or ( \5745_b1 , \5732_b1 , w_18203 );
not ( w_18203 , w_18204 );
and ( \5745_b0 , \5732_b0 , w_18205 );
and ( w_18204 ,  , w_18205 );
buf ( w_18203 , \5744_b1 );
not ( w_18203 , w_18206 );
not (  , w_18207 );
and ( w_18206 , w_18207 , \5744_b0 );
or ( \5746_b1 , \5419_b1 , \5437_b1 );
xor ( \5746_b0 , \5419_b0 , w_18208 );
not ( w_18208 , w_18209 );
and ( w_18209 , \5437_b1 , \5437_b0 );
or ( \5747_b1 , \5746_b1 , \5445_b1 );
xor ( \5747_b0 , \5746_b0 , w_18210 );
not ( w_18210 , w_18211 );
and ( w_18211 , \5445_b1 , \5445_b0 );
or ( \5748_b1 , \5745_b1 , \5747_b1 );
xor ( \5748_b0 , \5745_b0 , w_18212 );
not ( w_18212 , w_18213 );
and ( w_18213 , \5747_b1 , \5747_b0 );
buf ( \5749_b1 , \4198_b1 );
not ( \5749_b1 , w_18214 );
not ( \5749_b0 , w_18215 );
and ( w_18214 , w_18215 , \4198_b0 );
buf ( \5750_b1 , \5422_b1 );
not ( \5750_b1 , w_18216 );
not ( \5750_b0 , w_18217 );
and ( w_18216 , w_18217 , \5422_b0 );
or ( \5751_b1 , \5749_b1 , w_18218 );
or ( \5751_b0 , \5749_b0 , \5750_b0 );
not ( \5750_b0 , w_18219 );
and ( w_18219 , w_18218 , \5750_b1 );
or ( \5752_b1 , \5433_b1 , w_18221 );
not ( w_18221 , w_18222 );
and ( \5752_b0 , \5433_b0 , w_18223 );
and ( w_18222 ,  , w_18223 );
buf ( w_18221 , \4209_b1 );
not ( w_18221 , w_18224 );
not (  , w_18225 );
and ( w_18224 , w_18225 , \4209_b0 );
or ( \5753_b1 , \5751_b1 , w_18227 );
not ( w_18227 , w_18228 );
and ( \5753_b0 , \5751_b0 , w_18229 );
and ( w_18228 ,  , w_18229 );
buf ( w_18227 , \5752_b1 );
not ( w_18227 , w_18230 );
not (  , w_18231 );
and ( w_18230 , w_18231 , \5752_b0 );
buf ( \5754_b1 , \5753_b1 );
not ( \5754_b1 , w_18232 );
not ( \5754_b0 , w_18233 );
and ( w_18232 , w_18233 , \5753_b0 );
buf ( \5755_b1 , \5271_b1 );
not ( \5755_b1 , w_18234 );
not ( \5755_b0 , w_18235 );
and ( w_18234 , w_18235 , \5271_b0 );
or ( \5756_b1 , \5754_b1 , w_18236 );
or ( \5756_b0 , \5754_b0 , \5755_b0 );
not ( \5755_b0 , w_18237 );
and ( w_18237 , w_18236 , \5755_b1 );
or ( \5757_b1 , \5427_b1 , w_18239 );
not ( w_18239 , w_18240 );
and ( \5757_b0 , \5427_b0 , w_18241 );
and ( w_18240 ,  , w_18241 );
buf ( w_18239 , \5266_b1 );
not ( w_18239 , w_18242 );
not (  , w_18243 );
and ( w_18242 , w_18243 , \5266_b0 );
or ( \5758_b1 , \5756_b1 , w_18245 );
not ( w_18245 , w_18246 );
and ( \5758_b0 , \5756_b0 , w_18247 );
and ( w_18246 ,  , w_18247 );
buf ( w_18245 , \5757_b1 );
not ( w_18245 , w_18248 );
not (  , w_18249 );
and ( w_18248 , w_18249 , \5757_b0 );
buf ( \5759_b1 , \4098_b1 );
not ( \5759_b1 , w_18250 );
not ( \5759_b0 , w_18251 );
and ( w_18250 , w_18251 , \4098_b0 );
buf ( \5760_b1 , \4346_b1 );
not ( \5760_b1 , w_18252 );
not ( \5760_b0 , w_18253 );
and ( w_18252 , w_18253 , \4346_b0 );
or ( \5761_b1 , \5759_b1 , w_18254 );
or ( \5761_b0 , \5759_b0 , \5760_b0 );
not ( \5760_b0 , w_18255 );
and ( w_18255 , w_18254 , \5760_b1 );
or ( \5762_b1 , \4100_b1 , w_18257 );
not ( w_18257 , w_18258 );
and ( \5762_b0 , \4100_b0 , w_18259 );
and ( w_18258 ,  , w_18259 );
buf ( w_18257 , \5418_b1 );
not ( w_18257 , w_18260 );
not (  , w_18261 );
and ( w_18260 , w_18261 , \5418_b0 );
or ( \5763_b1 , \5761_b1 , w_18263 );
not ( w_18263 , w_18264 );
and ( \5763_b0 , \5761_b0 , w_18265 );
and ( w_18264 ,  , w_18265 );
buf ( w_18263 , \5762_b1 );
not ( w_18263 , w_18266 );
not (  , w_18267 );
and ( w_18266 , w_18267 , \5762_b0 );
buf ( \5764_b1 , \5763_b1 );
not ( \5764_b1 , w_18268 );
not ( \5764_b0 , w_18269 );
and ( w_18268 , w_18269 , \5763_b0 );
buf ( \5765_b1 , \4194_b1 );
not ( \5765_b1 , w_18270 );
not ( \5765_b0 , w_18271 );
and ( w_18270 , w_18271 , \4194_b0 );
or ( \5766_b1 , \5764_b1 , w_18272 );
or ( \5766_b0 , \5764_b0 , \5765_b0 );
not ( \5765_b0 , w_18273 );
and ( w_18273 , w_18272 , \5765_b1 );
or ( \5767_b1 , \5528_b1 , w_18275 );
not ( w_18275 , w_18276 );
and ( \5767_b0 , \5528_b0 , w_18277 );
and ( w_18276 ,  , w_18277 );
buf ( w_18275 , \4200_b1 );
not ( w_18275 , w_18278 );
not (  , w_18279 );
and ( w_18278 , w_18279 , \4200_b0 );
or ( \5768_b1 , \5766_b1 , w_18281 );
not ( w_18281 , w_18282 );
and ( \5768_b0 , \5766_b0 , w_18283 );
and ( w_18282 ,  , w_18283 );
buf ( w_18281 , \5767_b1 );
not ( w_18281 , w_18284 );
not (  , w_18285 );
and ( w_18284 , w_18285 , \5767_b0 );
or ( \5769_b1 , \5758_b1 , \5768_b1 );
xor ( \5769_b0 , \5758_b0 , w_18286 );
not ( w_18286 , w_18287 );
and ( w_18287 , \5768_b1 , \5768_b0 );
or ( \5770_b1 , \4519_b1 , \4458_b1 );
not ( \4458_b1 , w_18288 );
and ( \5770_b0 , \4519_b0 , w_18289 );
and ( w_18288 , w_18289 , \4458_b0 );
buf ( \5771_b1 , \4519_b1 );
not ( \5771_b1 , w_18290 );
not ( \5771_b0 , w_18291 );
and ( w_18290 , w_18291 , \4519_b0 );
or ( \5772_b1 , \5771_b1 , \4535_b1 );
not ( \4535_b1 , w_18292 );
and ( \5772_b0 , \5771_b0 , w_18293 );
and ( w_18292 , w_18293 , \4535_b0 );
or ( \5773_b1 , \5770_b1 , w_18295 );
not ( w_18295 , w_18296 );
and ( \5773_b0 , \5770_b0 , w_18297 );
and ( w_18296 ,  , w_18297 );
buf ( w_18295 , \5772_b1 );
not ( w_18295 , w_18298 );
not (  , w_18299 );
and ( w_18298 , w_18299 , \5772_b0 );
buf ( \5774_b1 , \5773_b1 );
not ( \5774_b1 , w_18300 );
not ( \5774_b0 , w_18301 );
and ( w_18300 , w_18301 , \5773_b0 );
buf ( \5775_b1 , \5774_b1 );
not ( \5775_b1 , w_18302 );
not ( \5775_b0 , w_18303 );
and ( w_18302 , w_18303 , \5774_b0 );
buf ( \5776_b1 , \4632_b1 );
not ( \5776_b1 , w_18304 );
not ( \5776_b0 , w_18305 );
and ( w_18304 , w_18305 , \4632_b0 );
or ( \5777_b1 , \5775_b1 , w_18306 );
or ( \5777_b0 , \5775_b0 , \5776_b0 );
not ( \5776_b0 , w_18307 );
and ( w_18307 , w_18306 , \5776_b1 );
or ( \5778_b1 , \4453_b1 , w_18309 );
not ( w_18309 , w_18310 );
and ( \5778_b0 , \4453_b0 , w_18311 );
and ( w_18310 ,  , w_18311 );
buf ( w_18309 , \5512_b1 );
not ( w_18309 , w_18312 );
not (  , w_18313 );
and ( w_18312 , w_18313 , \5512_b0 );
or ( \5779_b1 , \5777_b1 , w_18315 );
not ( w_18315 , w_18316 );
and ( \5779_b0 , \5777_b0 , w_18317 );
and ( w_18316 ,  , w_18317 );
buf ( w_18315 , \5778_b1 );
not ( w_18315 , w_18318 );
not (  , w_18319 );
and ( w_18318 , w_18319 , \5778_b0 );
or ( \5780_b1 , \5769_b1 , \5779_b1 );
not ( \5779_b1 , w_18320 );
and ( \5780_b0 , \5769_b0 , w_18321 );
and ( w_18320 , w_18321 , \5779_b0 );
or ( \5781_b1 , \5758_b1 , \5768_b1 );
not ( \5768_b1 , w_18322 );
and ( \5781_b0 , \5758_b0 , w_18323 );
and ( w_18322 , w_18323 , \5768_b0 );
or ( \5782_b1 , \5780_b1 , w_18324 );
or ( \5782_b0 , \5780_b0 , \5781_b0 );
not ( \5781_b0 , w_18325 );
and ( w_18325 , w_18324 , \5781_b1 );
or ( \5783_b1 , \5748_b1 , \5782_b1 );
not ( \5782_b1 , w_18326 );
and ( \5783_b0 , \5748_b0 , w_18327 );
and ( w_18326 , w_18327 , \5782_b0 );
or ( \5784_b1 , \5745_b1 , \5747_b1 );
not ( \5747_b1 , w_18328 );
and ( \5784_b0 , \5745_b0 , w_18329 );
and ( w_18328 , w_18329 , \5747_b0 );
or ( \5785_b1 , \5783_b1 , w_18330 );
or ( \5785_b0 , \5783_b0 , \5784_b0 );
not ( \5784_b0 , w_18331 );
and ( w_18331 , w_18330 , \5784_b1 );
buf ( \5786_b1 , \5785_b1 );
not ( \5786_b1 , w_18332 );
not ( \5786_b0 , w_18333 );
and ( w_18332 , w_18333 , \5785_b0 );
or ( \5787_b1 , \5725_b1 , w_18335 );
not ( w_18335 , w_18336 );
and ( \5787_b0 , \5725_b0 , w_18337 );
and ( w_18336 ,  , w_18337 );
buf ( w_18335 , \5786_b1 );
not ( w_18335 , w_18338 );
not (  , w_18339 );
and ( w_18338 , w_18339 , \5786_b0 );
or ( \5788_b1 , \5506_b1 , \5521_b1 );
xor ( \5788_b0 , \5506_b0 , w_18340 );
not ( w_18340 , w_18341 );
and ( w_18341 , \5521_b1 , \5521_b0 );
or ( \5789_b1 , \5788_b1 , \5539_b1 );
xor ( \5789_b0 , \5788_b0 , w_18342 );
not ( w_18342 , w_18343 );
and ( w_18343 , \5539_b1 , \5539_b0 );
buf ( \5790_b1 , \5789_b1 );
not ( \5790_b1 , w_18344 );
not ( \5790_b0 , w_18345 );
and ( w_18344 , w_18345 , \5789_b0 );
buf ( \5791_b1 , \4093_b1 );
not ( \5791_b1 , w_18346 );
not ( \5791_b0 , w_18347 );
and ( w_18346 , w_18347 , \4093_b0 );
buf ( \5792_b1 , \4746_b1 );
not ( \5792_b1 , w_18348 );
not ( \5792_b0 , w_18349 );
and ( w_18348 , w_18349 , \4746_b0 );
or ( \5793_b1 , \5791_b1 , w_18350 );
or ( \5793_b0 , \5791_b0 , \5792_b0 );
not ( \5792_b0 , w_18351 );
and ( w_18351 , w_18350 , \5792_b1 );
or ( \5794_b1 , \4615_b1 , w_18353 );
not ( w_18353 , w_18354 );
and ( \5794_b0 , \4615_b0 , w_18355 );
and ( w_18354 ,  , w_18355 );
buf ( w_18353 , \4349_b1 );
not ( w_18353 , w_18356 );
not (  , w_18357 );
and ( w_18356 , w_18357 , \4349_b0 );
or ( \5795_b1 , \5793_b1 , w_18359 );
not ( w_18359 , w_18360 );
and ( \5795_b0 , \5793_b0 , w_18361 );
and ( w_18360 ,  , w_18361 );
buf ( w_18359 , \5794_b1 );
not ( w_18359 , w_18362 );
not (  , w_18363 );
and ( w_18362 , w_18363 , \5794_b0 );
buf ( \5796_b1 , \5795_b1 );
not ( \5796_b1 , w_18364 );
not ( \5796_b0 , w_18365 );
and ( w_18364 , w_18365 , \5795_b0 );
buf ( \5797_b1 , \4610_b1 );
not ( \5797_b1 , w_18366 );
not ( \5797_b0 , w_18367 );
and ( w_18366 , w_18367 , \4610_b0 );
or ( \5798_b1 , \5796_b1 , w_18368 );
or ( \5798_b0 , \5796_b0 , \5797_b0 );
not ( \5797_b0 , w_18369 );
and ( w_18369 , w_18368 , \5797_b1 );
or ( \5799_b1 , \5465_b1 , w_18371 );
not ( w_18371 , w_18372 );
and ( \5799_b0 , \5465_b0 , w_18373 );
and ( w_18372 ,  , w_18373 );
buf ( w_18371 , \5146_b1 );
not ( w_18371 , w_18374 );
not (  , w_18375 );
and ( w_18374 , w_18375 , \5146_b0 );
or ( \5800_b1 , \5798_b1 , w_18377 );
not ( w_18377 , w_18378 );
and ( \5800_b0 , \5798_b0 , w_18379 );
and ( w_18378 ,  , w_18379 );
buf ( w_18377 , \5799_b1 );
not ( w_18377 , w_18380 );
not (  , w_18381 );
and ( w_18380 , w_18381 , \5799_b0 );
buf ( \5801_b1 , \5800_b1 );
buf ( \5801_b0 , \5800_b0 );
buf ( \5802_b1 , \5801_b1 );
not ( \5802_b1 , w_18382 );
not ( \5802_b0 , w_18383 );
and ( w_18382 , w_18383 , \5801_b0 );
buf ( \5803_b1 , \4158_b1 );
not ( \5803_b1 , w_18384 );
not ( \5803_b0 , w_18385 );
and ( w_18384 , w_18385 , \4158_b0 );
buf ( \5804_b1 , \5803_b1 );
not ( \5804_b1 , w_18386 );
not ( \5804_b0 , w_18387 );
and ( w_18386 , w_18387 , \5803_b0 );
or ( \5805_b1 , \5089_b1 , \4170_b1 );
not ( \4170_b1 , w_18388 );
and ( \5805_b0 , \5089_b0 , w_18389 );
and ( w_18388 , w_18389 , \4170_b0 );
buf ( \5806_b1 , \5089_b1 );
not ( \5806_b1 , w_18390 );
not ( \5806_b0 , w_18391 );
and ( w_18390 , w_18391 , \5089_b0 );
or ( \5807_b1 , \5806_b1 , \4163_b1 );
not ( \4163_b1 , w_18392 );
and ( \5807_b0 , \5806_b0 , w_18393 );
and ( w_18392 , w_18393 , \4163_b0 );
or ( \5808_b1 , \5805_b1 , w_18395 );
not ( w_18395 , w_18396 );
and ( \5808_b0 , \5805_b0 , w_18397 );
and ( w_18396 ,  , w_18397 );
buf ( w_18395 , \5807_b1 );
not ( w_18395 , w_18398 );
not (  , w_18399 );
and ( w_18398 , w_18399 , \5807_b0 );
buf ( \5809_b1 , \5808_b1 );
not ( \5809_b1 , w_18400 );
not ( \5809_b0 , w_18401 );
and ( w_18400 , w_18401 , \5808_b0 );
or ( \5810_b1 , \5804_b1 , \5809_b1 );
not ( \5809_b1 , w_18402 );
and ( \5810_b0 , \5804_b0 , w_18403 );
and ( w_18402 , w_18403 , \5809_b0 );
buf ( \5811_b1 , \5453_b1 );
not ( \5811_b1 , w_18404 );
not ( \5811_b0 , w_18405 );
and ( w_18404 , w_18405 , \5453_b0 );
or ( \5812_b1 , \5811_b1 , w_18407 );
not ( w_18407 , w_18408 );
and ( \5812_b0 , \5811_b0 , w_18409 );
and ( w_18408 ,  , w_18409 );
buf ( w_18407 , \4151_b1 );
not ( w_18407 , w_18410 );
not (  , w_18411 );
and ( w_18410 , w_18411 , \4151_b0 );
or ( \5813_b1 , \5810_b1 , w_18413 );
not ( w_18413 , w_18414 );
and ( \5813_b0 , \5810_b0 , w_18415 );
and ( w_18414 ,  , w_18415 );
buf ( w_18413 , \5812_b1 );
not ( w_18413 , w_18416 );
not (  , w_18417 );
and ( w_18416 , w_18417 , \5812_b0 );
buf ( \5814_b1 , \5813_b1 );
not ( \5814_b1 , w_18418 );
not ( \5814_b0 , w_18419 );
and ( w_18418 , w_18419 , \5813_b0 );
buf ( \5815_b1 , \5814_b1 );
not ( \5815_b1 , w_18420 );
not ( \5815_b0 , w_18421 );
and ( w_18420 , w_18421 , \5814_b0 );
or ( \5816_b1 , \5802_b1 , w_18422 );
or ( \5816_b0 , \5802_b0 , \5815_b0 );
not ( \5815_b0 , w_18423 );
and ( w_18423 , w_18422 , \5815_b1 );
or ( \5817_b1 , \5814_b1 , w_18424 );
or ( \5817_b0 , \5814_b0 , \5801_b0 );
not ( \5801_b0 , w_18425 );
and ( w_18425 , w_18424 , \5801_b1 );
buf ( \5818_b1 , \4278_b1 );
not ( \5818_b1 , w_18426 );
not ( \5818_b0 , w_18427 );
and ( w_18426 , w_18427 , \4278_b0 );
or ( \5819_b1 , \4021_b1 , \4332_b1 );
not ( \4332_b1 , w_18428 );
and ( \5819_b0 , \4021_b0 , w_18429 );
and ( w_18428 , w_18429 , \4332_b0 );
buf ( \5820_b1 , \4021_b1 );
not ( \5820_b1 , w_18430 );
not ( \5820_b0 , w_18431 );
and ( w_18430 , w_18431 , \4021_b0 );
or ( \5821_b1 , \5820_b1 , \4283_b1 );
not ( \4283_b1 , w_18432 );
and ( \5821_b0 , \5820_b0 , w_18433 );
and ( w_18432 , w_18433 , \4283_b0 );
or ( \5822_b1 , \5819_b1 , w_18435 );
not ( w_18435 , w_18436 );
and ( \5822_b0 , \5819_b0 , w_18437 );
and ( w_18436 ,  , w_18437 );
buf ( w_18435 , \5821_b1 );
not ( w_18435 , w_18438 );
not (  , w_18439 );
and ( w_18438 , w_18439 , \5821_b0 );
buf ( \5823_b1 , \5822_b1 );
not ( \5823_b1 , w_18440 );
not ( \5823_b0 , w_18441 );
and ( w_18440 , w_18441 , \5822_b0 );
or ( \5824_b1 , \5818_b1 , \5823_b1 );
not ( \5823_b1 , w_18442 );
and ( \5824_b0 , \5818_b0 , w_18443 );
and ( w_18442 , w_18443 , \5823_b0 );
or ( \5825_b1 , \5495_b1 , \4266_b1 );
not ( \4266_b1 , w_18444 );
and ( \5825_b0 , \5495_b0 , w_18445 );
and ( w_18444 , w_18445 , \4266_b0 );
or ( \5826_b1 , \5824_b1 , w_18447 );
not ( w_18447 , w_18448 );
and ( \5826_b0 , \5824_b0 , w_18449 );
and ( w_18448 ,  , w_18449 );
buf ( w_18447 , \5825_b1 );
not ( w_18447 , w_18450 );
not (  , w_18451 );
and ( w_18450 , w_18451 , \5825_b0 );
buf ( \5827_b1 , \5826_b1 );
not ( \5827_b1 , w_18452 );
not ( \5827_b0 , w_18453 );
and ( w_18452 , w_18453 , \5826_b0 );
or ( \5828_b1 , \5817_b1 , w_18455 );
not ( w_18455 , w_18456 );
and ( \5828_b0 , \5817_b0 , w_18457 );
and ( w_18456 ,  , w_18457 );
buf ( w_18455 , \5827_b1 );
not ( w_18455 , w_18458 );
not (  , w_18459 );
and ( w_18458 , w_18459 , \5827_b0 );
or ( \5829_b1 , \5816_b1 , w_18461 );
not ( w_18461 , w_18462 );
and ( \5829_b0 , \5816_b0 , w_18463 );
and ( w_18462 ,  , w_18463 );
buf ( w_18461 , \5828_b1 );
not ( w_18461 , w_18464 );
not (  , w_18465 );
and ( w_18464 , w_18465 , \5828_b0 );
buf ( \5830_b1 , \5829_b1 );
not ( \5830_b1 , w_18466 );
not ( \5830_b0 , w_18467 );
and ( w_18466 , w_18467 , \5829_b0 );
or ( \5831_b1 , \5790_b1 , w_18468 );
or ( \5831_b0 , \5790_b0 , \5830_b0 );
not ( \5830_b0 , w_18469 );
and ( w_18469 , w_18468 , \5830_b1 );
or ( \5832_b1 , \5789_b1 , w_18470 );
or ( \5832_b0 , \5789_b0 , \5829_b0 );
not ( \5829_b0 , w_18471 );
and ( w_18471 , w_18470 , \5829_b1 );
or ( \5833_b1 , \5474_b1 , \5458_b1 );
xor ( \5833_b0 , \5474_b0 , w_18472 );
not ( w_18472 , w_18473 );
and ( w_18473 , \5458_b1 , \5458_b0 );
or ( \5834_b1 , \5833_b1 , w_18474 );
xor ( \5834_b0 , \5833_b0 , w_18476 );
not ( w_18476 , w_18477 );
and ( w_18477 , w_18474 , w_18475 );
buf ( w_18474 , \5487_b1 );
not ( w_18474 , w_18478 );
not ( w_18475 , w_18479 );
and ( w_18478 , w_18479 , \5487_b0 );
buf ( \5835_b1 , \5834_b1 );
not ( \5835_b1 , w_18480 );
not ( \5835_b0 , w_18481 );
and ( w_18480 , w_18481 , \5834_b0 );
or ( \5836_b1 , \5832_b1 , w_18483 );
not ( w_18483 , w_18484 );
and ( \5836_b0 , \5832_b0 , w_18485 );
and ( w_18484 ,  , w_18485 );
buf ( w_18483 , \5835_b1 );
not ( w_18483 , w_18486 );
not (  , w_18487 );
and ( w_18486 , w_18487 , \5835_b0 );
or ( \5837_b1 , \5831_b1 , w_18489 );
not ( w_18489 , w_18490 );
and ( \5837_b0 , \5831_b0 , w_18491 );
and ( w_18490 ,  , w_18491 );
buf ( w_18489 , \5836_b1 );
not ( w_18489 , w_18492 );
not (  , w_18493 );
and ( w_18492 , w_18493 , \5836_b0 );
or ( \5838_b1 , \5787_b1 , \5837_b1 );
not ( \5837_b1 , w_18494 );
and ( \5838_b0 , \5787_b0 , w_18495 );
and ( w_18494 , w_18495 , \5837_b0 );
or ( \5839_b1 , \5785_b1 , \5724_b1 );
not ( \5724_b1 , w_18496 );
and ( \5839_b0 , \5785_b0 , w_18497 );
and ( w_18496 , w_18497 , \5724_b0 );
or ( \5840_b1 , \5838_b1 , w_18499 );
not ( w_18499 , w_18500 );
and ( \5840_b0 , \5838_b0 , w_18501 );
and ( w_18500 ,  , w_18501 );
buf ( w_18499 , \5839_b1 );
not ( w_18499 , w_18502 );
not (  , w_18503 );
and ( w_18502 , w_18503 , \5839_b0 );
buf ( \5841_b1 , \5840_b1 );
not ( \5841_b1 , w_18504 );
not ( \5841_b0 , w_18505 );
and ( w_18504 , w_18505 , \5840_b0 );
or ( \5842_b1 , \5722_b1 , w_18506 );
or ( \5842_b0 , \5722_b0 , \5841_b0 );
not ( \5841_b0 , w_18507 );
and ( w_18507 , w_18506 , \5841_b1 );
or ( \5843_b1 , \5721_b1 , w_18508 );
or ( \5843_b0 , \5721_b0 , \5840_b0 );
not ( \5840_b0 , w_18509 );
and ( w_18509 , w_18508 , \5840_b1 );
or ( \5844_b1 , \5842_b1 , w_18511 );
not ( w_18511 , w_18512 );
and ( \5844_b0 , \5842_b0 , w_18513 );
and ( w_18512 ,  , w_18513 );
buf ( w_18511 , \5843_b1 );
not ( w_18511 , w_18514 );
not (  , w_18515 );
and ( w_18514 , w_18515 , \5843_b0 );
buf ( \5845_b1 , \5844_b1 );
not ( \5845_b1 , w_18516 );
not ( \5845_b0 , w_18517 );
and ( w_18516 , w_18517 , \5844_b0 );
or ( \5846_b1 , \5719_b1 , w_18518 );
or ( \5846_b0 , \5719_b0 , \5845_b0 );
not ( \5845_b0 , w_18519 );
and ( w_18519 , w_18518 , \5845_b1 );
buf ( \5847_b1 , \5717_b1 );
not ( \5847_b1 , w_18520 );
not ( \5847_b0 , w_18521 );
and ( w_18520 , w_18521 , \5717_b0 );
or ( \5848_b1 , \5847_b1 , w_18522 );
or ( \5848_b0 , \5847_b0 , \5844_b0 );
not ( \5844_b0 , w_18523 );
and ( w_18523 , w_18522 , \5844_b1 );
or ( \5849_b1 , \5846_b1 , w_18525 );
not ( w_18525 , w_18526 );
and ( \5849_b0 , \5846_b0 , w_18527 );
and ( w_18526 ,  , w_18527 );
buf ( w_18525 , \5848_b1 );
not ( w_18525 , w_18528 );
not (  , w_18529 );
and ( w_18528 , w_18529 , \5848_b0 );
buf ( \5850_b1 , \5665_b1 );
not ( \5850_b1 , w_18530 );
not ( \5850_b0 , w_18531 );
and ( w_18530 , w_18531 , \5665_b0 );
buf ( \5851_b1 , \5685_b1 );
not ( \5851_b1 , w_18532 );
not ( \5851_b0 , w_18533 );
and ( w_18532 , w_18533 , \5685_b0 );
or ( \5852_b1 , \5850_b1 , w_18534 );
or ( \5852_b0 , \5850_b0 , \5851_b0 );
not ( \5851_b0 , w_18535 );
and ( w_18535 , w_18534 , \5851_b1 );
or ( \5853_b1 , \5665_b1 , w_18536 );
or ( \5853_b0 , \5665_b0 , \5685_b0 );
not ( \5685_b0 , w_18537 );
and ( w_18537 , w_18536 , \5685_b1 );
or ( \5854_b1 , \5852_b1 , w_18539 );
not ( w_18539 , w_18540 );
and ( \5854_b0 , \5852_b0 , w_18541 );
and ( w_18540 ,  , w_18541 );
buf ( w_18539 , \5853_b1 );
not ( w_18539 , w_18542 );
not (  , w_18543 );
and ( w_18542 , w_18543 , \5853_b0 );
or ( \5855_b1 , \5854_b1 , \5669_b1 );
not ( \5669_b1 , w_18544 );
and ( \5855_b0 , \5854_b0 , w_18545 );
and ( w_18544 , w_18545 , \5669_b0 );
buf ( \5856_b1 , \5854_b1 );
not ( \5856_b1 , w_18546 );
not ( \5856_b0 , w_18547 );
and ( w_18546 , w_18547 , \5854_b0 );
buf ( \5857_b1 , \5668_b1 );
buf ( \5857_b0 , \5668_b0 );
or ( \5858_b1 , \5856_b1 , \5857_b1 );
not ( \5857_b1 , w_18548 );
and ( \5858_b0 , \5856_b0 , w_18549 );
and ( w_18548 , w_18549 , \5857_b0 );
or ( \5859_b1 , \5855_b1 , w_18551 );
not ( w_18551 , w_18552 );
and ( \5859_b0 , \5855_b0 , w_18553 );
and ( w_18552 ,  , w_18553 );
buf ( w_18551 , \5858_b1 );
not ( w_18551 , w_18554 );
not (  , w_18555 );
and ( w_18554 , w_18555 , \5858_b0 );
buf ( \5860_b1 , \5859_b1 );
not ( \5860_b1 , w_18556 );
not ( \5860_b0 , w_18557 );
and ( w_18556 , w_18557 , \5859_b0 );
buf ( \5861_b1 , \5860_b1 );
not ( \5861_b1 , w_18558 );
not ( \5861_b0 , w_18559 );
and ( w_18558 , w_18559 , \5860_b0 );
buf ( \5862_b1 , \5861_b1 );
not ( \5862_b1 , w_18560 );
not ( \5862_b0 , w_18561 );
and ( w_18560 , w_18561 , \5861_b0 );
or ( \5863_b1 , \5785_b1 , \5724_b1 );
xor ( \5863_b0 , \5785_b0 , w_18562 );
not ( w_18562 , w_18563 );
and ( w_18563 , \5724_b1 , \5724_b0 );
buf ( \5864_b1 , \5837_b1 );
not ( \5864_b1 , w_18564 );
not ( \5864_b0 , w_18565 );
and ( w_18564 , w_18565 , \5837_b0 );
or ( \5865_b1 , \5863_b1 , \5864_b1 );
not ( \5864_b1 , w_18566 );
and ( \5865_b0 , \5863_b0 , w_18567 );
and ( w_18566 , w_18567 , \5864_b0 );
buf ( \5866_b1 , \5863_b1 );
not ( \5866_b1 , w_18568 );
not ( \5866_b0 , w_18569 );
and ( w_18568 , w_18569 , \5863_b0 );
or ( \5867_b1 , \5866_b1 , \5837_b1 );
not ( \5837_b1 , w_18570 );
and ( \5867_b0 , \5866_b0 , w_18571 );
and ( w_18570 , w_18571 , \5837_b0 );
or ( \5868_b1 , \5865_b1 , w_18573 );
not ( w_18573 , w_18574 );
and ( \5868_b0 , \5865_b0 , w_18575 );
and ( w_18574 ,  , w_18575 );
buf ( w_18573 , \5867_b1 );
not ( w_18573 , w_18576 );
not (  , w_18577 );
and ( w_18576 , w_18577 , \5867_b0 );
buf ( \5869_b1 , \5868_b1 );
not ( \5869_b1 , w_18578 );
not ( \5869_b0 , w_18579 );
and ( w_18578 , w_18579 , \5868_b0 );
buf ( \5870_b1 , \5869_b1 );
not ( \5870_b1 , w_18580 );
not ( \5870_b0 , w_18581 );
and ( w_18580 , w_18581 , \5869_b0 );
or ( \5871_b1 , \5862_b1 , w_18582 );
or ( \5871_b0 , \5862_b0 , \5870_b0 );
not ( \5870_b0 , w_18583 );
and ( w_18583 , w_18582 , \5870_b1 );
buf ( \5872_b1 , \5860_b1 );
not ( \5872_b1 , w_18584 );
not ( \5872_b0 , w_18585 );
and ( w_18584 , w_18585 , \5860_b0 );
buf ( \5873_b1 , \5868_b1 );
not ( \5873_b1 , w_18586 );
not ( \5873_b0 , w_18587 );
and ( w_18586 , w_18587 , \5868_b0 );
or ( \5874_b1 , \5872_b1 , w_18588 );
or ( \5874_b0 , \5872_b0 , \5873_b0 );
not ( \5873_b0 , w_18589 );
and ( w_18589 , w_18588 , \5873_b1 );
or ( \5875_b1 , \5744_b1 , w_18590 );
xor ( \5875_b0 , \5744_b0 , w_18592 );
not ( w_18592 , w_18593 );
and ( w_18593 , w_18590 , w_18591 );
buf ( w_18590 , \5732_b1 );
not ( w_18590 , w_18594 );
not ( w_18591 , w_18595 );
and ( w_18594 , w_18595 , \5732_b0 );
buf ( \5876_b1 , \4079_b1 );
not ( \5876_b1 , w_18596 );
not ( \5876_b0 , w_18597 );
and ( w_18596 , w_18597 , \4079_b0 );
buf ( \5877_b1 , \4107_b1 );
not ( \5877_b1 , w_18598 );
not ( \5877_b0 , w_18599 );
and ( w_18598 , w_18599 , \4107_b0 );
or ( \5878_b1 , \5876_b1 , w_18600 );
or ( \5878_b0 , \5876_b0 , \5877_b0 );
not ( \5877_b0 , w_18601 );
and ( w_18601 , w_18600 , \5877_b1 );
or ( \5879_b1 , \4110_b1 , w_18603 );
not ( w_18603 , w_18604 );
and ( \5879_b0 , \4110_b0 , w_18605 );
and ( w_18604 ,  , w_18605 );
buf ( w_18603 , \5535_b1 );
not ( w_18603 , w_18606 );
not (  , w_18607 );
and ( w_18606 , w_18607 , \5535_b0 );
or ( \5880_b1 , \5878_b1 , w_18609 );
not ( w_18609 , w_18610 );
and ( \5880_b0 , \5878_b0 , w_18611 );
and ( w_18610 ,  , w_18611 );
buf ( w_18609 , \5879_b1 );
not ( w_18609 , w_18612 );
not (  , w_18613 );
and ( w_18612 , w_18613 , \5879_b0 );
buf ( \5881_b1 , \5880_b1 );
not ( \5881_b1 , w_18614 );
not ( \5881_b0 , w_18615 );
and ( w_18614 , w_18615 , \5880_b0 );
buf ( \5882_b1 , \4302_b1 );
not ( \5882_b1 , w_18616 );
not ( \5882_b0 , w_18617 );
and ( w_18616 , w_18617 , \4302_b0 );
or ( \5883_b1 , \5881_b1 , w_18618 );
or ( \5883_b0 , \5881_b0 , \5882_b0 );
not ( \5882_b0 , w_18619 );
and ( w_18619 , w_18618 , \5882_b1 );
or ( \5884_b1 , \4133_b1 , w_18621 );
not ( w_18621 , w_18622 );
and ( \5884_b0 , \4133_b0 , w_18623 );
and ( w_18622 ,  , w_18623 );
buf ( w_18621 , \5482_b1 );
not ( w_18621 , w_18624 );
not (  , w_18625 );
and ( w_18624 , w_18625 , \5482_b0 );
or ( \5885_b1 , \5883_b1 , w_18627 );
not ( w_18627 , w_18628 );
and ( \5885_b0 , \5883_b0 , w_18629 );
and ( w_18628 ,  , w_18629 );
buf ( w_18627 , \5884_b1 );
not ( w_18627 , w_18630 );
not (  , w_18631 );
and ( w_18630 , w_18631 , \5884_b0 );
buf ( \5886_b1 , \5885_b1 );
not ( \5886_b1 , w_18632 );
not ( \5886_b0 , w_18633 );
and ( w_18632 , w_18633 , \5885_b0 );
or ( \5887_b1 , \5875_b1 , w_18635 );
not ( w_18635 , w_18636 );
and ( \5887_b0 , \5875_b0 , w_18637 );
and ( w_18636 ,  , w_18637 );
buf ( w_18635 , \5886_b1 );
not ( w_18635 , w_18638 );
not (  , w_18639 );
and ( w_18638 , w_18639 , \5886_b0 );
or ( \5888_b1 , \4192_b1 , w_18641 );
not ( w_18641 , w_18642 );
and ( \5888_b0 , \4192_b0 , w_18643 );
and ( w_18642 ,  , w_18643 );
buf ( w_18641 , \5418_b1 );
not ( w_18641 , w_18644 );
not (  , w_18645 );
and ( w_18644 , w_18645 , \5418_b0 );
buf ( \5889_b1 , \5266_b1 );
not ( \5889_b1 , w_18646 );
not ( \5889_b0 , w_18647 );
and ( w_18646 , w_18647 , \5266_b0 );
buf ( \5890_b1 , \5753_b1 );
not ( \5890_b1 , w_18648 );
not ( \5890_b0 , w_18649 );
and ( w_18648 , w_18649 , \5753_b0 );
or ( \5891_b1 , \5889_b1 , w_18650 );
or ( \5891_b0 , \5889_b0 , \5890_b0 );
not ( \5890_b0 , w_18651 );
and ( w_18651 , w_18650 , \5890_b1 );
buf ( \5892_b1 , \4094_b1 );
not ( \5892_b1 , w_18652 );
not ( \5892_b0 , w_18653 );
and ( w_18652 , w_18653 , \4094_b0 );
buf ( \5893_b1 , \5274_b1 );
not ( \5893_b1 , w_18654 );
not ( \5893_b0 , w_18655 );
and ( w_18654 , w_18655 , \5274_b0 );
or ( \5894_b1 , \5892_b1 , w_18656 );
or ( \5894_b0 , \5892_b0 , \5893_b0 );
not ( \5893_b0 , w_18657 );
and ( w_18657 , w_18656 , \5893_b1 );
or ( \5895_b1 , \5268_b1 , w_18659 );
not ( w_18659 , w_18660 );
and ( \5895_b0 , \5268_b0 , w_18661 );
and ( w_18660 ,  , w_18661 );
buf ( w_18659 , \4298_b1 );
not ( w_18659 , w_18662 );
not (  , w_18663 );
and ( w_18662 , w_18663 , \4298_b0 );
or ( \5896_b1 , \5894_b1 , w_18665 );
not ( w_18665 , w_18666 );
and ( \5896_b0 , \5894_b0 , w_18667 );
and ( w_18666 ,  , w_18667 );
buf ( w_18665 , \5895_b1 );
not ( w_18665 , w_18668 );
not (  , w_18669 );
and ( w_18668 , w_18669 , \5895_b0 );
or ( \5897_b1 , \5271_b1 , w_18671 );
not ( w_18671 , w_18672 );
and ( \5897_b0 , \5271_b0 , w_18673 );
and ( w_18672 ,  , w_18673 );
buf ( w_18671 , \5896_b1 );
not ( w_18671 , w_18674 );
not (  , w_18675 );
and ( w_18674 , w_18675 , \5896_b0 );
or ( \5898_b1 , \5891_b1 , w_18677 );
not ( w_18677 , w_18678 );
and ( \5898_b0 , \5891_b0 , w_18679 );
and ( w_18678 ,  , w_18679 );
buf ( w_18677 , \5897_b1 );
not ( w_18677 , w_18680 );
not (  , w_18681 );
and ( w_18680 , w_18681 , \5897_b0 );
or ( \5899_b1 , \5888_b1 , \5898_b1 );
xor ( \5899_b0 , \5888_b0 , w_18682 );
not ( w_18682 , w_18683 );
and ( w_18683 , \5898_b1 , \5898_b0 );
buf ( \5900_b1 , \4948_b1 );
not ( \5900_b1 , w_18684 );
not ( \5900_b0 , w_18685 );
and ( w_18684 , w_18685 , \4948_b0 );
buf ( \5901_b1 , \5737_b1 );
not ( \5901_b1 , w_18686 );
not ( \5901_b0 , w_18687 );
and ( w_18686 , w_18687 , \5737_b0 );
or ( \5902_b1 , \5900_b1 , w_18688 );
or ( \5902_b0 , \5900_b0 , \5901_b0 );
not ( \5901_b0 , w_18689 );
and ( w_18689 , w_18688 , \5901_b1 );
buf ( \5903_b1 , \2945_b1 );
not ( \5903_b1 , w_18690 );
not ( \5903_b0 , w_18691 );
and ( w_18690 , w_18691 , \2945_b0 );
or ( \5904_b1 , \5903_b1 , \4097_b1 );
not ( \4097_b1 , w_18692 );
and ( \5904_b0 , \5903_b0 , w_18693 );
and ( w_18692 , w_18693 , \4097_b0 );
buf ( \5905_b1 , \4853_b1 );
not ( \5905_b1 , w_18694 );
not ( \5905_b0 , w_18695 );
and ( w_18694 , w_18695 , \4853_b0 );
or ( \5906_b1 , \5905_b1 , \4254_b1 );
not ( \4254_b1 , w_18696 );
and ( \5906_b0 , \5905_b0 , w_18697 );
and ( w_18696 , w_18697 , \4254_b0 );
or ( \5907_b1 , \5904_b1 , w_18699 );
not ( w_18699 , w_18700 );
and ( \5907_b0 , \5904_b0 , w_18701 );
and ( w_18700 ,  , w_18701 );
buf ( w_18699 , \5906_b1 );
not ( w_18699 , w_18702 );
not (  , w_18703 );
and ( w_18702 , w_18703 , \5906_b0 );
buf ( \5908_b1 , \5907_b1 );
not ( \5908_b1 , w_18704 );
not ( \5908_b0 , w_18705 );
and ( w_18704 , w_18705 , \5907_b0 );
or ( \5909_b1 , \5908_b1 , w_18707 );
not ( w_18707 , w_18708 );
and ( \5909_b0 , \5908_b0 , w_18709 );
and ( w_18708 ,  , w_18709 );
buf ( w_18707 , \4944_b1 );
not ( w_18707 , w_18710 );
not (  , w_18711 );
and ( w_18710 , w_18711 , \4944_b0 );
or ( \5910_b1 , \5902_b1 , w_18713 );
not ( w_18713 , w_18714 );
and ( \5910_b0 , \5902_b0 , w_18715 );
and ( w_18714 ,  , w_18715 );
buf ( w_18713 , \5909_b1 );
not ( w_18713 , w_18716 );
not (  , w_18717 );
and ( w_18716 , w_18717 , \5909_b0 );
or ( \5911_b1 , \5899_b1 , \5910_b1 );
not ( \5910_b1 , w_18718 );
and ( \5911_b0 , \5899_b0 , w_18719 );
and ( w_18718 , w_18719 , \5910_b0 );
or ( \5912_b1 , \5888_b1 , \5898_b1 );
not ( \5898_b1 , w_18720 );
and ( \5912_b0 , \5888_b0 , w_18721 );
and ( w_18720 , w_18721 , \5898_b0 );
or ( \5913_b1 , \5911_b1 , w_18722 );
or ( \5913_b0 , \5911_b0 , \5912_b0 );
not ( \5912_b0 , w_18723 );
and ( w_18723 , w_18722 , \5912_b1 );
or ( \5914_b1 , \5887_b1 , \5913_b1 );
not ( \5913_b1 , w_18724 );
and ( \5914_b0 , \5887_b0 , w_18725 );
and ( w_18724 , w_18725 , \5913_b0 );
or ( \5915_b1 , \5875_b1 , w_18727 );
not ( w_18727 , w_18728 );
and ( \5915_b0 , \5875_b0 , w_18729 );
and ( w_18728 ,  , w_18729 );
buf ( w_18727 , \5886_b1 );
not ( w_18727 , w_18730 );
not (  , w_18731 );
and ( w_18730 , w_18731 , \5886_b0 );
or ( \5916_b1 , \5914_b1 , w_18733 );
not ( w_18733 , w_18734 );
and ( \5916_b0 , \5914_b0 , w_18735 );
and ( w_18734 ,  , w_18735 );
buf ( w_18733 , \5915_b1 );
not ( w_18733 , w_18736 );
not (  , w_18737 );
and ( w_18736 , w_18737 , \5915_b0 );
buf ( \5917_b1 , \5916_b1 );
not ( \5917_b1 , w_18738 );
not ( \5917_b0 , w_18739 );
and ( w_18738 , w_18739 , \5916_b0 );
buf ( \5918_b1 , \5917_b1 );
not ( \5918_b1 , w_18740 );
not ( \5918_b0 , w_18741 );
and ( w_18740 , w_18741 , \5917_b0 );
buf ( \5919_b1 , \4610_b1 );
not ( \5919_b1 , w_18742 );
not ( \5919_b0 , w_18743 );
and ( w_18742 , w_18743 , \4610_b0 );
buf ( \5920_b1 , \4095_b1 );
not ( \5920_b1 , w_18744 );
not ( \5920_b0 , w_18745 );
and ( w_18744 , w_18745 , \4095_b0 );
buf ( \5921_b1 , \5138_b1 );
not ( \5921_b1 , w_18746 );
not ( \5921_b0 , w_18747 );
and ( w_18746 , w_18747 , \5138_b0 );
or ( \5922_b1 , \5920_b1 , w_18748 );
or ( \5922_b0 , \5920_b0 , \5921_b0 );
not ( \5921_b0 , w_18749 );
and ( w_18749 , w_18748 , \5921_b1 );
or ( \5923_b1 , \4745_b1 , w_18751 );
not ( w_18751 , w_18752 );
and ( \5923_b0 , \4745_b0 , w_18753 );
and ( w_18752 ,  , w_18753 );
buf ( w_18751 , \4391_b1 );
not ( w_18751 , w_18754 );
not (  , w_18755 );
and ( w_18754 , w_18755 , \4391_b0 );
or ( \5924_b1 , \5922_b1 , w_18757 );
not ( w_18757 , w_18758 );
and ( \5924_b0 , \5922_b0 , w_18759 );
and ( w_18758 ,  , w_18759 );
buf ( w_18757 , \5923_b1 );
not ( w_18757 , w_18760 );
not (  , w_18761 );
and ( w_18760 , w_18761 , \5923_b0 );
buf ( \5925_b1 , \5924_b1 );
not ( \5925_b1 , w_18762 );
not ( \5925_b0 , w_18763 );
and ( w_18762 , w_18763 , \5924_b0 );
or ( \5926_b1 , \5919_b1 , w_18764 );
or ( \5926_b0 , \5919_b0 , \5925_b0 );
not ( \5925_b0 , w_18765 );
and ( w_18765 , w_18764 , \5925_b1 );
or ( \5927_b1 , \5795_b1 , w_18767 );
not ( w_18767 , w_18768 );
and ( \5927_b0 , \5795_b0 , w_18769 );
and ( w_18768 ,  , w_18769 );
buf ( w_18767 , \5146_b1 );
not ( w_18767 , w_18770 );
not (  , w_18771 );
and ( w_18770 , w_18771 , \5146_b0 );
or ( \5928_b1 , \5926_b1 , w_18773 );
not ( w_18773 , w_18774 );
and ( \5928_b0 , \5926_b0 , w_18775 );
and ( w_18774 ,  , w_18775 );
buf ( w_18773 , \5927_b1 );
not ( w_18773 , w_18776 );
not (  , w_18777 );
and ( w_18776 , w_18777 , \5927_b0 );
buf ( \5929_b1 , \5928_b1 );
not ( \5929_b1 , w_18778 );
not ( \5929_b0 , w_18779 );
and ( w_18778 , w_18779 , \5928_b0 );
buf ( \5930_b1 , \4450_b1 );
not ( \5930_b1 , w_18780 );
not ( \5930_b0 , w_18781 );
and ( w_18780 , w_18781 , \4450_b0 );
or ( \5931_b1 , \4662_b1 , \4458_b1 );
not ( \4458_b1 , w_18782 );
and ( \5931_b0 , \4662_b0 , w_18783 );
and ( w_18782 , w_18783 , \4458_b0 );
buf ( \5932_b1 , \4662_b1 );
not ( \5932_b1 , w_18784 );
not ( \5932_b0 , w_18785 );
and ( w_18784 , w_18785 , \4662_b0 );
or ( \5933_b1 , \5932_b1 , \4535_b1 );
not ( \4535_b1 , w_18786 );
and ( \5933_b0 , \5932_b0 , w_18787 );
and ( w_18786 , w_18787 , \4535_b0 );
or ( \5934_b1 , \5931_b1 , w_18789 );
not ( w_18789 , w_18790 );
and ( \5934_b0 , \5931_b0 , w_18791 );
and ( w_18790 ,  , w_18791 );
buf ( w_18789 , \5933_b1 );
not ( w_18789 , w_18792 );
not (  , w_18793 );
and ( w_18792 , w_18793 , \5933_b0 );
buf ( \5935_b1 , \5934_b1 );
not ( \5935_b1 , w_18794 );
not ( \5935_b0 , w_18795 );
and ( w_18794 , w_18795 , \5934_b0 );
or ( \5936_b1 , \5930_b1 , \5935_b1 );
not ( \5935_b1 , w_18796 );
and ( \5936_b0 , \5930_b0 , w_18797 );
and ( w_18796 , w_18797 , \5935_b0 );
buf ( \5937_b1 , \4452_b1 );
not ( \5937_b1 , w_18798 );
not ( \5937_b0 , w_18799 );
and ( w_18798 , w_18799 , \4452_b0 );
or ( \5938_b1 , \5937_b1 , w_18801 );
not ( w_18801 , w_18802 );
and ( \5938_b0 , \5937_b0 , w_18803 );
and ( w_18802 ,  , w_18803 );
buf ( w_18801 , \5773_b1 );
not ( w_18801 , w_18804 );
not (  , w_18805 );
and ( w_18804 , w_18805 , \5773_b0 );
or ( \5939_b1 , \5936_b1 , w_18807 );
not ( w_18807 , w_18808 );
and ( \5939_b0 , \5936_b0 , w_18809 );
and ( w_18808 ,  , w_18809 );
buf ( w_18807 , \5938_b1 );
not ( w_18807 , w_18810 );
not (  , w_18811 );
and ( w_18810 , w_18811 , \5938_b0 );
buf ( \5940_b1 , \5939_b1 );
not ( \5940_b1 , w_18812 );
not ( \5940_b0 , w_18813 );
and ( w_18812 , w_18813 , \5939_b0 );
buf ( \5941_b1 , \5940_b1 );
not ( \5941_b1 , w_18814 );
not ( \5941_b0 , w_18815 );
and ( w_18814 , w_18815 , \5940_b0 );
or ( \5942_b1 , \5929_b1 , w_18816 );
or ( \5942_b0 , \5929_b0 , \5941_b0 );
not ( \5941_b0 , w_18817 );
and ( w_18817 , w_18816 , \5941_b1 );
buf ( \5943_b1 , \5928_b1 );
not ( \5943_b1 , w_18818 );
not ( \5943_b0 , w_18819 );
and ( w_18818 , w_18819 , \5928_b0 );
buf ( \5944_b1 , \5943_b1 );
not ( \5944_b1 , w_18820 );
not ( \5944_b0 , w_18821 );
and ( w_18820 , w_18821 , \5943_b0 );
buf ( \5945_b1 , \5939_b1 );
not ( \5945_b1 , w_18822 );
not ( \5945_b0 , w_18823 );
and ( w_18822 , w_18823 , \5939_b0 );
or ( \5946_b1 , \5944_b1 , w_18824 );
or ( \5946_b0 , \5944_b0 , \5945_b0 );
not ( \5945_b0 , w_18825 );
and ( w_18825 , w_18824 , \5945_b1 );
buf ( \5947_b1 , \4026_b1 );
not ( \5947_b1 , w_18826 );
not ( \5947_b0 , w_18827 );
and ( w_18826 , w_18827 , \4026_b0 );
buf ( \5948_b1 , \4332_b1 );
not ( \5948_b1 , w_18828 );
not ( \5948_b0 , w_18829 );
and ( w_18828 , w_18829 , \4332_b0 );
or ( \5949_b1 , \5947_b1 , w_18830 );
or ( \5949_b0 , \5947_b0 , \5948_b0 );
not ( \5948_b0 , w_18831 );
and ( w_18831 , w_18830 , \5948_b1 );
or ( \5950_b1 , \4673_b1 , w_18833 );
not ( w_18833 , w_18834 );
and ( \5950_b0 , \4673_b0 , w_18835 );
and ( w_18834 ,  , w_18835 );
buf ( w_18833 , \4969_b1 );
not ( w_18833 , w_18836 );
not (  , w_18837 );
and ( w_18836 , w_18837 , \4969_b0 );
or ( \5951_b1 , \5949_b1 , w_18839 );
not ( w_18839 , w_18840 );
and ( \5951_b0 , \5949_b0 , w_18841 );
and ( w_18840 ,  , w_18841 );
buf ( w_18839 , \5950_b1 );
not ( w_18839 , w_18842 );
not (  , w_18843 );
and ( w_18842 , w_18843 , \5950_b0 );
buf ( \5952_b1 , \5951_b1 );
not ( \5952_b1 , w_18844 );
not ( \5952_b0 , w_18845 );
and ( w_18844 , w_18845 , \5951_b0 );
buf ( \5953_b1 , \5497_b1 );
not ( \5953_b1 , w_18846 );
not ( \5953_b0 , w_18847 );
and ( w_18846 , w_18847 , \5497_b0 );
or ( \5954_b1 , \5952_b1 , w_18848 );
or ( \5954_b0 , \5952_b0 , \5953_b0 );
not ( \5953_b0 , w_18849 );
and ( w_18849 , w_18848 , \5953_b1 );
buf ( \5955_b1 , \5822_b1 );
not ( \5955_b1 , w_18850 );
not ( \5955_b0 , w_18851 );
and ( w_18850 , w_18851 , \5822_b0 );
or ( \5956_b1 , \5955_b1 , w_18853 );
not ( w_18853 , w_18854 );
and ( \5956_b0 , \5955_b0 , w_18855 );
and ( w_18854 ,  , w_18855 );
buf ( w_18853 , \4800_b1 );
not ( w_18853 , w_18856 );
not (  , w_18857 );
and ( w_18856 , w_18857 , \4800_b0 );
or ( \5957_b1 , \5954_b1 , w_18859 );
not ( w_18859 , w_18860 );
and ( \5957_b0 , \5954_b0 , w_18861 );
and ( w_18860 ,  , w_18861 );
buf ( w_18859 , \5956_b1 );
not ( w_18859 , w_18862 );
not (  , w_18863 );
and ( w_18862 , w_18863 , \5956_b0 );
or ( \5958_b1 , \5946_b1 , w_18865 );
not ( w_18865 , w_18866 );
and ( \5958_b0 , \5946_b0 , w_18867 );
and ( w_18866 ,  , w_18867 );
buf ( w_18865 , \5957_b1 );
not ( w_18865 , w_18868 );
not (  , w_18869 );
and ( w_18868 , w_18869 , \5957_b0 );
or ( \5959_b1 , \5942_b1 , w_18871 );
not ( w_18871 , w_18872 );
and ( \5959_b0 , \5942_b0 , w_18873 );
and ( w_18872 ,  , w_18873 );
buf ( w_18871 , \5958_b1 );
not ( w_18871 , w_18874 );
not (  , w_18875 );
and ( w_18874 , w_18875 , \5958_b0 );
buf ( \5960_b1 , \5959_b1 );
not ( \5960_b1 , w_18876 );
not ( \5960_b0 , w_18877 );
and ( w_18876 , w_18877 , \5959_b0 );
buf ( \5961_b1 , \5800_b1 );
not ( \5961_b1 , w_18878 );
not ( \5961_b0 , w_18879 );
and ( w_18878 , w_18879 , \5800_b0 );
buf ( \5962_b1 , \5961_b1 );
not ( \5962_b1 , w_18880 );
not ( \5962_b0 , w_18881 );
and ( w_18880 , w_18881 , \5961_b0 );
buf ( \5963_b1 , \5827_b1 );
not ( \5963_b1 , w_18882 );
not ( \5963_b0 , w_18883 );
and ( w_18882 , w_18883 , \5827_b0 );
or ( \5964_b1 , \5962_b1 , w_18884 );
or ( \5964_b0 , \5962_b0 , \5963_b0 );
not ( \5963_b0 , w_18885 );
and ( w_18885 , w_18884 , \5963_b1 );
or ( \5965_b1 , \5826_b1 , w_18887 );
not ( w_18887 , w_18888 );
and ( \5965_b0 , \5826_b0 , w_18889 );
and ( w_18888 ,  , w_18889 );
buf ( w_18887 , \5800_b1 );
not ( w_18887 , w_18890 );
not (  , w_18891 );
and ( w_18890 , w_18891 , \5800_b0 );
or ( \5966_b1 , \5964_b1 , w_18893 );
not ( w_18893 , w_18894 );
and ( \5966_b0 , \5964_b0 , w_18895 );
and ( w_18894 ,  , w_18895 );
buf ( w_18893 , \5965_b1 );
not ( w_18893 , w_18896 );
not (  , w_18897 );
and ( w_18896 , w_18897 , \5965_b0 );
or ( \5967_b1 , \5966_b1 , \5813_b1 );
not ( \5813_b1 , w_18898 );
and ( \5967_b0 , \5966_b0 , w_18899 );
and ( w_18898 , w_18899 , \5813_b0 );
buf ( \5968_b1 , \5966_b1 );
not ( \5968_b1 , w_18900 );
not ( \5968_b0 , w_18901 );
and ( w_18900 , w_18901 , \5966_b0 );
or ( \5969_b1 , \5968_b1 , \5814_b1 );
not ( \5814_b1 , w_18902 );
and ( \5969_b0 , \5968_b0 , w_18903 );
and ( w_18902 , w_18903 , \5814_b0 );
or ( \5970_b1 , \5967_b1 , w_18905 );
not ( w_18905 , w_18906 );
and ( \5970_b0 , \5967_b0 , w_18907 );
and ( w_18906 ,  , w_18907 );
buf ( w_18905 , \5969_b1 );
not ( w_18905 , w_18908 );
not (  , w_18909 );
and ( w_18908 , w_18909 , \5969_b0 );
or ( \5971_b1 , \5960_b1 , w_18911 );
not ( w_18911 , w_18912 );
and ( \5971_b0 , \5960_b0 , w_18913 );
and ( w_18912 ,  , w_18913 );
buf ( w_18911 , \5970_b1 );
not ( w_18911 , w_18914 );
not (  , w_18915 );
and ( w_18914 , w_18915 , \5970_b0 );
or ( \5972_b1 , \5907_b1 , w_18916 );
or ( \5972_b0 , \5907_b0 , \4862_b0 );
not ( \4862_b0 , w_18917 );
and ( w_18917 , w_18916 , \4862_b1 );
buf ( \5973_b1 , \4093_b1 );
not ( \5973_b1 , w_18918 );
not ( \5973_b0 , w_18919 );
and ( w_18918 , w_18919 , \4093_b0 );
buf ( \5974_b1 , \5905_b1 );
not ( \5974_b1 , w_18920 );
not ( \5974_b0 , w_18921 );
and ( w_18920 , w_18921 , \5905_b0 );
buf ( \5975_b1 , \5974_b1 );
not ( \5975_b1 , w_18922 );
not ( \5975_b0 , w_18923 );
and ( w_18922 , w_18923 , \5974_b0 );
or ( \5976_b1 , \5973_b1 , w_18924 );
or ( \5976_b0 , \5973_b0 , \5975_b0 );
not ( \5975_b0 , w_18925 );
and ( w_18925 , w_18924 , \5975_b1 );
or ( \5977_b1 , \5905_b1 , w_18927 );
not ( w_18927 , w_18928 );
and ( \5977_b0 , \5905_b0 , w_18929 );
and ( w_18928 ,  , w_18929 );
buf ( w_18927 , \4349_b1 );
not ( w_18927 , w_18930 );
not (  , w_18931 );
and ( w_18930 , w_18931 , \4349_b0 );
or ( \5978_b1 , \5976_b1 , w_18933 );
not ( w_18933 , w_18934 );
and ( \5978_b0 , \5976_b0 , w_18935 );
and ( w_18934 ,  , w_18935 );
buf ( w_18933 , \5977_b1 );
not ( w_18933 , w_18936 );
not (  , w_18937 );
and ( w_18936 , w_18937 , \5977_b0 );
or ( \5980_b1 , \5972_b1 , w_18939 );
not ( w_18939 , w_18940 );
and ( \5980_b0 , \5972_b0 , w_18941 );
and ( w_18940 ,  , w_18941 );
buf ( w_18939 , \5979_b1 );
not ( w_18939 , w_18942 );
not (  , w_18943 );
and ( w_18942 , w_18943 , \5979_b0 );
or ( \5981_b1 , \4116_b1 , w_18945 );
not ( w_18945 , w_18946 );
and ( \5981_b0 , \4116_b0 , w_18947 );
and ( w_18946 ,  , w_18947 );
buf ( w_18945 , \5418_b1 );
not ( w_18945 , w_18948 );
not (  , w_18949 );
and ( w_18948 , w_18949 , \5418_b0 );
or ( \5982_b1 , \4170_b1 , \5981_b1 );
not ( \5981_b1 , w_18950 );
and ( \5982_b0 , \4170_b0 , w_18951 );
and ( w_18950 , w_18951 , \5981_b0 );
buf ( \5983_b1 , \4098_b1 );
not ( \5983_b1 , w_18952 );
not ( \5983_b0 , w_18953 );
and ( w_18952 , w_18953 , \4098_b0 );
buf ( \5984_b1 , \4115_b1 );
not ( \5984_b1 , w_18954 );
not ( \5984_b0 , w_18955 );
and ( w_18954 , w_18955 , \4115_b0 );
or ( \5985_b1 , \5983_b1 , w_18956 );
or ( \5985_b0 , \5983_b0 , \5984_b0 );
not ( \5984_b0 , w_18957 );
and ( w_18957 , w_18956 , \5984_b1 );
or ( \5986_b1 , \5985_b1 , w_18959 );
not ( w_18959 , w_18960 );
and ( \5986_b0 , \5985_b0 , w_18961 );
and ( w_18960 ,  , w_18961 );
buf ( w_18959 , \4106_b1 );
not ( w_18959 , w_18962 );
not (  , w_18963 );
and ( w_18962 , w_18963 , \4106_b0 );
or ( \5987_b1 , \5982_b1 , w_18965 );
not ( w_18965 , w_18966 );
and ( \5987_b0 , \5982_b0 , w_18967 );
and ( w_18966 ,  , w_18967 );
buf ( w_18965 , \5986_b1 );
not ( w_18965 , w_18968 );
not (  , w_18969 );
and ( w_18968 , w_18969 , \5986_b0 );
or ( \5988_b1 , \5980_b1 , w_18971 );
not ( w_18971 , w_18972 );
and ( \5988_b0 , \5980_b0 , w_18973 );
and ( w_18972 ,  , w_18973 );
buf ( w_18971 , \5987_b1 );
not ( w_18971 , w_18974 );
not (  , w_18975 );
and ( w_18974 , w_18975 , \5987_b0 );
buf ( \5989_b1 , \5988_b1 );
not ( \5989_b1 , w_18976 );
not ( \5989_b0 , w_18977 );
and ( w_18976 , w_18977 , \5988_b0 );
buf ( \5990_b1 , \4082_b1 );
not ( \5990_b1 , w_18978 );
not ( \5990_b0 , w_18979 );
and ( w_18978 , w_18979 , \4082_b0 );
buf ( \5991_b1 , \4107_b1 );
not ( \5991_b1 , w_18980 );
not ( \5991_b0 , w_18981 );
and ( w_18980 , w_18981 , \4107_b0 );
or ( \5992_b1 , \5990_b1 , w_18982 );
or ( \5992_b0 , \5990_b0 , \5991_b0 );
not ( \5991_b0 , w_18983 );
and ( w_18983 , w_18982 , \5991_b1 );
or ( \5993_b1 , \4110_b1 , w_18985 );
not ( w_18985 , w_18986 );
and ( \5993_b0 , \4110_b0 , w_18987 );
and ( w_18986 ,  , w_18987 );
buf ( w_18985 , \5526_b1 );
not ( w_18985 , w_18988 );
not (  , w_18989 );
and ( w_18988 , w_18989 , \5526_b0 );
or ( \5994_b1 , \5992_b1 , w_18991 );
not ( w_18991 , w_18992 );
and ( \5994_b0 , \5992_b0 , w_18993 );
and ( w_18992 ,  , w_18993 );
buf ( w_18991 , \5993_b1 );
not ( w_18991 , w_18994 );
not (  , w_18995 );
and ( w_18994 , w_18995 , \5993_b0 );
buf ( \5995_b1 , \5994_b1 );
not ( \5995_b1 , w_18996 );
not ( \5995_b0 , w_18997 );
and ( w_18996 , w_18997 , \5994_b0 );
buf ( \5996_b1 , \4128_b1 );
not ( \5996_b1 , w_18998 );
not ( \5996_b0 , w_18999 );
and ( w_18998 , w_18999 , \4128_b0 );
or ( \5997_b1 , \5995_b1 , w_19000 );
or ( \5997_b0 , \5995_b0 , \5996_b0 );
not ( \5996_b0 , w_19001 );
and ( w_19001 , w_19000 , \5996_b1 );
or ( \5998_b1 , \5880_b1 , w_19003 );
not ( w_19003 , w_19004 );
and ( \5998_b0 , \5880_b0 , w_19005 );
and ( w_19004 ,  , w_19005 );
buf ( w_19003 , \4132_b1 );
not ( w_19003 , w_19006 );
not (  , w_19007 );
and ( w_19006 , w_19007 , \4132_b0 );
or ( \5999_b1 , \5997_b1 , w_19009 );
not ( w_19009 , w_19010 );
and ( \5999_b0 , \5997_b0 , w_19011 );
and ( w_19010 ,  , w_19011 );
buf ( w_19009 , \5998_b1 );
not ( w_19009 , w_19012 );
not (  , w_19013 );
and ( w_19012 , w_19013 , \5998_b0 );
buf ( \6000_b1 , \5999_b1 );
not ( \6000_b1 , w_19014 );
not ( \6000_b0 , w_19015 );
and ( w_19014 , w_19015 , \5999_b0 );
buf ( \6001_b1 , \6000_b1 );
not ( \6001_b1 , w_19016 );
not ( \6001_b0 , w_19017 );
and ( w_19016 , w_19017 , \6000_b0 );
or ( \6002_b1 , \5989_b1 , w_19018 );
or ( \6002_b0 , \5989_b0 , \6001_b0 );
not ( \6001_b0 , w_19019 );
and ( w_19019 , w_19018 , \6001_b1 );
buf ( \6003_b1 , \4076_b1 );
not ( \6003_b1 , w_19020 );
not ( \6003_b0 , w_19021 );
and ( w_19020 , w_19021 , \4076_b0 );
buf ( \6004_b1 , \4163_b1 );
not ( \6004_b1 , w_19022 );
not ( \6004_b0 , w_19023 );
and ( w_19022 , w_19023 , \4163_b0 );
or ( \6005_b1 , \6003_b1 , w_19024 );
or ( \6005_b0 , \6003_b0 , \6004_b0 );
not ( \6004_b0 , w_19025 );
and ( w_19025 , w_19024 , \6004_b1 );
or ( \6006_b1 , \4311_b1 , w_19027 );
not ( w_19027 , w_19028 );
and ( \6006_b0 , \4311_b0 , w_19029 );
and ( w_19028 ,  , w_19029 );
buf ( w_19027 , \5284_b1 );
not ( w_19027 , w_19030 );
not (  , w_19031 );
and ( w_19030 , w_19031 , \5284_b0 );
or ( \6007_b1 , \6005_b1 , w_19033 );
not ( w_19033 , w_19034 );
and ( \6007_b0 , \6005_b0 , w_19035 );
and ( w_19034 ,  , w_19035 );
buf ( w_19033 , \6006_b1 );
not ( w_19033 , w_19036 );
not (  , w_19037 );
and ( w_19036 , w_19037 , \6006_b0 );
buf ( \6008_b1 , \6007_b1 );
not ( \6008_b1 , w_19038 );
not ( \6008_b0 , w_19039 );
and ( w_19038 , w_19039 , \6007_b0 );
buf ( \6009_b1 , \4159_b1 );
not ( \6009_b1 , w_19040 );
not ( \6009_b0 , w_19041 );
and ( w_19040 , w_19041 , \4159_b0 );
or ( \6010_b1 , \6008_b1 , w_19042 );
or ( \6010_b0 , \6008_b0 , \6009_b0 );
not ( \6009_b0 , w_19043 );
and ( w_19043 , w_19042 , \6009_b1 );
buf ( \6011_b1 , \5808_b1 );
not ( \6011_b1 , w_19044 );
not ( \6011_b0 , w_19045 );
and ( w_19044 , w_19045 , \5808_b0 );
or ( \6012_b1 , \6011_b1 , w_19047 );
not ( w_19047 , w_19048 );
and ( \6012_b0 , \6011_b0 , w_19049 );
and ( w_19048 ,  , w_19049 );
buf ( w_19047 , \4317_b1 );
not ( w_19047 , w_19050 );
not (  , w_19051 );
and ( w_19050 , w_19051 , \4317_b0 );
or ( \6013_b1 , \6010_b1 , w_19053 );
not ( w_19053 , w_19054 );
and ( \6013_b0 , \6010_b0 , w_19055 );
and ( w_19054 ,  , w_19055 );
buf ( w_19053 , \6012_b1 );
not ( w_19053 , w_19056 );
not (  , w_19057 );
and ( w_19056 , w_19057 , \6012_b0 );
or ( \6014_b1 , \6002_b1 , w_19059 );
not ( w_19059 , w_19060 );
and ( \6014_b0 , \6002_b0 , w_19061 );
and ( w_19060 ,  , w_19061 );
buf ( w_19059 , \6013_b1 );
not ( w_19059 , w_19062 );
not (  , w_19063 );
and ( w_19062 , w_19063 , \6013_b0 );
buf ( \6015_b1 , \5988_b1 );
not ( \6015_b1 , w_19064 );
not ( \6015_b0 , w_19065 );
and ( w_19064 , w_19065 , \5988_b0 );
or ( \6016_b1 , \6015_b1 , w_19067 );
not ( w_19067 , w_19068 );
and ( \6016_b0 , \6015_b0 , w_19069 );
and ( w_19068 ,  , w_19069 );
buf ( w_19067 , \5999_b1 );
not ( w_19067 , w_19070 );
not (  , w_19071 );
and ( w_19070 , w_19071 , \5999_b0 );
or ( \6017_b1 , \6014_b1 , w_19073 );
not ( w_19073 , w_19074 );
and ( \6017_b0 , \6014_b0 , w_19075 );
and ( w_19074 ,  , w_19075 );
buf ( w_19073 , \6016_b1 );
not ( w_19073 , w_19076 );
not (  , w_19077 );
and ( w_19076 , w_19077 , \6016_b0 );
or ( \6018_b1 , \5971_b1 , \6017_b1 );
not ( \6017_b1 , w_19078 );
and ( \6018_b0 , \5971_b0 , w_19079 );
and ( w_19078 , w_19079 , \6017_b0 );
or ( \6019_b1 , \5970_b1 , w_19081 );
not ( w_19081 , w_19082 );
and ( \6019_b0 , \5970_b0 , w_19083 );
and ( w_19082 ,  , w_19083 );
buf ( w_19081 , \5960_b1 );
not ( w_19081 , w_19084 );
not (  , w_19085 );
and ( w_19084 , w_19085 , \5960_b0 );
or ( \6020_b1 , \6018_b1 , w_19087 );
not ( w_19087 , w_19088 );
and ( \6020_b0 , \6018_b0 , w_19089 );
and ( w_19088 ,  , w_19089 );
buf ( w_19087 , \6019_b1 );
not ( w_19087 , w_19090 );
not (  , w_19091 );
and ( w_19090 , w_19091 , \6019_b0 );
buf ( \6021_b1 , \6020_b1 );
not ( \6021_b1 , w_19092 );
not ( \6021_b0 , w_19093 );
and ( w_19092 , w_19093 , \6020_b0 );
buf ( \6022_b1 , \6021_b1 );
not ( \6022_b1 , w_19094 );
not ( \6022_b0 , w_19095 );
and ( w_19094 , w_19095 , \6021_b0 );
or ( \6023_b1 , \5918_b1 , w_19096 );
or ( \6023_b0 , \5918_b0 , \6022_b0 );
not ( \6022_b0 , w_19097 );
and ( w_19097 , w_19096 , \6022_b1 );
buf ( \6024_b1 , \5916_b1 );
not ( \6024_b1 , w_19098 );
not ( \6024_b0 , w_19099 );
and ( w_19098 , w_19099 , \5916_b0 );
buf ( \6025_b1 , \6020_b1 );
not ( \6025_b1 , w_19100 );
not ( \6025_b0 , w_19101 );
and ( w_19100 , w_19101 , \6020_b0 );
or ( \6026_b1 , \6024_b1 , w_19102 );
or ( \6026_b0 , \6024_b0 , \6025_b0 );
not ( \6025_b0 , w_19103 );
and ( w_19103 , w_19102 , \6025_b1 );
or ( \6027_b1 , \5745_b1 , \5747_b1 );
xor ( \6027_b0 , \5745_b0 , w_19104 );
not ( w_19104 , w_19105 );
and ( w_19105 , \5747_b1 , \5747_b0 );
or ( \6028_b1 , \6027_b1 , \5782_b1 );
xor ( \6028_b0 , \6027_b0 , w_19106 );
not ( w_19106 , w_19107 );
and ( w_19107 , \5782_b1 , \5782_b0 );
or ( \6029_b1 , \6026_b1 , w_19109 );
not ( w_19109 , w_19110 );
and ( \6029_b0 , \6026_b0 , w_19111 );
and ( w_19110 ,  , w_19111 );
buf ( w_19109 , \6028_b1 );
not ( w_19109 , w_19112 );
not (  , w_19113 );
and ( w_19112 , w_19113 , \6028_b0 );
or ( \6030_b1 , \6023_b1 , w_19115 );
not ( w_19115 , w_19116 );
and ( \6030_b0 , \6023_b0 , w_19117 );
and ( w_19116 ,  , w_19117 );
buf ( w_19115 , \6029_b1 );
not ( w_19115 , w_19118 );
not (  , w_19119 );
and ( w_19118 , w_19119 , \6029_b0 );
or ( \6031_b1 , \5874_b1 , w_19121 );
not ( w_19121 , w_19122 );
and ( \6031_b0 , \5874_b0 , w_19123 );
and ( w_19122 ,  , w_19123 );
buf ( w_19121 , \6030_b1 );
not ( w_19121 , w_19124 );
not (  , w_19125 );
and ( w_19124 , w_19125 , \6030_b0 );
or ( \6032_b1 , \5871_b1 , w_19127 );
not ( w_19127 , w_19128 );
and ( \6032_b0 , \5871_b0 , w_19129 );
and ( w_19128 ,  , w_19129 );
buf ( w_19127 , \6031_b1 );
not ( w_19127 , w_19130 );
not (  , w_19131 );
and ( w_19130 , w_19131 , \6031_b0 );
or ( \6033_b1 , \5849_b1 , w_19133 );
not ( w_19133 , w_19134 );
and ( \6033_b0 , \5849_b0 , w_19135 );
and ( w_19134 ,  , w_19135 );
buf ( w_19133 , \6032_b1 );
not ( w_19133 , w_19136 );
not (  , w_19137 );
and ( w_19136 , w_19137 , \6032_b0 );
buf ( \6034_b1 , \6033_b1 );
not ( \6034_b1 , w_19138 );
not ( \6034_b0 , w_19139 );
and ( w_19138 , w_19139 , \6033_b0 );
buf ( \6035_b1 , \5868_b1 );
not ( \6035_b1 , w_19140 );
not ( \6035_b0 , w_19141 );
and ( w_19140 , w_19141 , \5868_b0 );
or ( \6036_b1 , \5859_b1 , \6030_b1 );
not ( \6030_b1 , w_19142 );
and ( \6036_b0 , \5859_b0 , w_19143 );
and ( w_19142 , w_19143 , \6030_b0 );
buf ( \6037_b1 , \5859_b1 );
not ( \6037_b1 , w_19144 );
not ( \6037_b0 , w_19145 );
and ( w_19144 , w_19145 , \5859_b0 );
buf ( \6038_b1 , \6030_b1 );
not ( \6038_b1 , w_19146 );
not ( \6038_b0 , w_19147 );
and ( w_19146 , w_19147 , \6030_b0 );
or ( \6039_b1 , \6037_b1 , \6038_b1 );
not ( \6038_b1 , w_19148 );
and ( \6039_b0 , \6037_b0 , w_19149 );
and ( w_19148 , w_19149 , \6038_b0 );
or ( \6040_b1 , \6036_b1 , w_19151 );
not ( w_19151 , w_19152 );
and ( \6040_b0 , \6036_b0 , w_19153 );
and ( w_19152 ,  , w_19153 );
buf ( w_19151 , \6039_b1 );
not ( w_19151 , w_19154 );
not (  , w_19155 );
and ( w_19154 , w_19155 , \6039_b0 );
buf ( \6041_b1 , \6040_b1 );
not ( \6041_b1 , w_19156 );
not ( \6041_b0 , w_19157 );
and ( w_19156 , w_19157 , \6040_b0 );
or ( \6042_b1 , \6035_b1 , w_19158 );
or ( \6042_b0 , \6035_b0 , \6041_b0 );
not ( \6041_b0 , w_19159 );
and ( w_19159 , w_19158 , \6041_b1 );
or ( \6043_b1 , \5868_b1 , w_19160 );
or ( \6043_b0 , \5868_b0 , \6040_b0 );
not ( \6040_b0 , w_19161 );
and ( w_19161 , w_19160 , \6040_b1 );
or ( \6044_b1 , \6042_b1 , w_19163 );
not ( w_19163 , w_19164 );
and ( \6044_b0 , \6042_b0 , w_19165 );
and ( w_19164 ,  , w_19165 );
buf ( w_19163 , \6043_b1 );
not ( w_19163 , w_19166 );
not (  , w_19167 );
and ( w_19166 , w_19167 , \6043_b0 );
buf ( \6045_b1 , \6044_b1 );
not ( \6045_b1 , w_19168 );
not ( \6045_b0 , w_19169 );
and ( w_19168 , w_19169 , \6044_b0 );
or ( \6046_b1 , \5829_b1 , \5834_b1 );
xor ( \6046_b0 , \5829_b0 , w_19170 );
not ( w_19170 , w_19171 );
and ( w_19171 , \5834_b1 , \5834_b0 );
or ( \6047_b1 , \6046_b1 , w_19172 );
xor ( \6047_b0 , \6046_b0 , w_19174 );
not ( w_19174 , w_19175 );
and ( w_19175 , w_19172 , w_19173 );
buf ( w_19172 , \5789_b1 );
not ( w_19172 , w_19176 );
not ( w_19173 , w_19177 );
and ( w_19176 , w_19177 , \5789_b0 );
or ( \6048_b1 , \5758_b1 , \5768_b1 );
xor ( \6048_b0 , \5758_b0 , w_19178 );
not ( w_19178 , w_19179 );
and ( w_19179 , \5768_b1 , \5768_b0 );
or ( \6049_b1 , \6048_b1 , \5779_b1 );
xor ( \6049_b0 , \6048_b0 , w_19180 );
not ( w_19180 , w_19181 );
and ( w_19181 , \5779_b1 , \5779_b0 );
or ( \6050_b1 , \5888_b1 , \5898_b1 );
xor ( \6050_b0 , \5888_b0 , w_19182 );
not ( w_19182 , w_19183 );
and ( w_19183 , \5898_b1 , \5898_b0 );
or ( \6051_b1 , \6050_b1 , \5910_b1 );
xor ( \6051_b0 , \6050_b0 , w_19184 );
not ( w_19184 , w_19185 );
and ( w_19185 , \5910_b1 , \5910_b0 );
buf ( \6052_b1 , \6051_b1 );
not ( \6052_b1 , w_19186 );
not ( \6052_b0 , w_19187 );
and ( w_19186 , w_19187 , \6051_b0 );
buf ( \6053_b1 , \5271_b1 );
not ( \6053_b1 , w_19188 );
not ( \6053_b0 , w_19189 );
and ( w_19188 , w_19189 , \5271_b0 );
buf ( \6054_b1 , \4096_b1 );
not ( \6054_b1 , w_19190 );
not ( \6054_b0 , w_19191 );
and ( w_19190 , w_19191 , \4096_b0 );
buf ( \6055_b1 , \5422_b1 );
not ( \6055_b1 , w_19192 );
not ( \6055_b0 , w_19193 );
and ( w_19192 , w_19193 , \5422_b0 );
or ( \6056_b1 , \6054_b1 , w_19194 );
or ( \6056_b0 , \6054_b0 , \6055_b0 );
not ( \6055_b0 , w_19195 );
and ( w_19195 , w_19194 , \6055_b1 );
or ( \6057_b1 , \4372_b1 , w_19197 );
not ( w_19197 , w_19198 );
and ( \6057_b0 , \4372_b0 , w_19199 );
and ( w_19198 ,  , w_19199 );
buf ( w_19197 , \5268_b1 );
not ( w_19197 , w_19200 );
not (  , w_19201 );
and ( w_19200 , w_19201 , \5268_b0 );
or ( \6058_b1 , \6056_b1 , w_19203 );
not ( w_19203 , w_19204 );
and ( \6058_b0 , \6056_b0 , w_19205 );
and ( w_19204 ,  , w_19205 );
buf ( w_19203 , \6057_b1 );
not ( w_19203 , w_19206 );
not (  , w_19207 );
and ( w_19206 , w_19207 , \6057_b0 );
buf ( \6059_b1 , \6058_b1 );
not ( \6059_b1 , w_19208 );
not ( \6059_b0 , w_19209 );
and ( w_19208 , w_19209 , \6058_b0 );
or ( \6060_b1 , \6053_b1 , w_19210 );
or ( \6060_b0 , \6053_b0 , \6059_b0 );
not ( \6059_b0 , w_19211 );
and ( w_19211 , w_19210 , \6059_b1 );
or ( \6061_b1 , \5896_b1 , w_19213 );
not ( w_19213 , w_19214 );
and ( \6061_b0 , \5896_b0 , w_19215 );
and ( w_19214 ,  , w_19215 );
buf ( w_19213 , \5266_b1 );
not ( w_19213 , w_19216 );
not (  , w_19217 );
and ( w_19216 , w_19217 , \5266_b0 );
or ( \6062_b1 , \6060_b1 , w_19219 );
not ( w_19219 , w_19220 );
and ( \6062_b0 , \6060_b0 , w_19221 );
and ( w_19220 ,  , w_19221 );
buf ( w_19219 , \6061_b1 );
not ( w_19219 , w_19222 );
not (  , w_19223 );
and ( w_19222 , w_19223 , \6061_b0 );
buf ( \6063_b1 , \6062_b1 );
not ( \6063_b1 , w_19224 );
not ( \6063_b0 , w_19225 );
and ( w_19224 , w_19225 , \6062_b0 );
buf ( \6064_b1 , \4449_b1 );
not ( \6064_b1 , w_19226 );
not ( \6064_b0 , w_19227 );
and ( w_19226 , w_19227 , \4449_b0 );
buf ( \6065_b1 , \4021_b1 );
not ( \6065_b1 , w_19228 );
not ( \6065_b0 , w_19229 );
and ( w_19228 , w_19229 , \4021_b0 );
buf ( \6066_b1 , \4532_b1 );
not ( \6066_b1 , w_19230 );
not ( \6066_b0 , w_19231 );
and ( w_19230 , w_19231 , \4532_b0 );
or ( \6067_b1 , \6065_b1 , w_19232 );
or ( \6067_b0 , \6065_b0 , \6066_b0 );
not ( \6066_b0 , w_19233 );
and ( w_19233 , w_19232 , \6066_b1 );
or ( \6068_b1 , \4458_b1 , w_19235 );
not ( w_19235 , w_19236 );
and ( \6068_b0 , \4458_b0 , w_19237 );
and ( w_19236 ,  , w_19237 );
buf ( w_19235 , \4780_b1 );
not ( w_19235 , w_19238 );
not (  , w_19239 );
and ( w_19238 , w_19239 , \4780_b0 );
or ( \6069_b1 , \6067_b1 , w_19241 );
not ( w_19241 , w_19242 );
and ( \6069_b0 , \6067_b0 , w_19243 );
and ( w_19242 ,  , w_19243 );
buf ( w_19241 , \6068_b1 );
not ( w_19241 , w_19244 );
not (  , w_19245 );
and ( w_19244 , w_19245 , \6068_b0 );
buf ( \6070_b1 , \6069_b1 );
not ( \6070_b1 , w_19246 );
not ( \6070_b0 , w_19247 );
and ( w_19246 , w_19247 , \6069_b0 );
or ( \6071_b1 , \6064_b1 , w_19248 );
or ( \6071_b0 , \6064_b0 , \6070_b0 );
not ( \6070_b0 , w_19249 );
and ( w_19249 , w_19248 , \6070_b1 );
buf ( \6072_b1 , \5934_b1 );
not ( \6072_b1 , w_19250 );
not ( \6072_b0 , w_19251 );
and ( w_19250 , w_19251 , \5934_b0 );
or ( \6073_b1 , \6072_b1 , w_19253 );
not ( w_19253 , w_19254 );
and ( \6073_b0 , \6072_b0 , w_19255 );
and ( w_19254 ,  , w_19255 );
buf ( w_19253 , \4452_b1 );
not ( w_19253 , w_19256 );
not (  , w_19257 );
and ( w_19256 , w_19257 , \4452_b0 );
or ( \6074_b1 , \6071_b1 , w_19259 );
not ( w_19259 , w_19260 );
and ( \6074_b0 , \6071_b0 , w_19261 );
and ( w_19260 ,  , w_19261 );
buf ( w_19259 , \6073_b1 );
not ( w_19259 , w_19262 );
not (  , w_19263 );
and ( w_19262 , w_19263 , \6073_b0 );
buf ( \6075_b1 , \6074_b1 );
not ( \6075_b1 , w_19264 );
not ( \6075_b0 , w_19265 );
and ( w_19264 , w_19265 , \6074_b0 );
or ( \6076_b1 , \6063_b1 , w_19266 );
or ( \6076_b0 , \6063_b0 , \6075_b0 );
not ( \6075_b0 , w_19267 );
and ( w_19267 , w_19266 , \6075_b1 );
or ( \6077_b1 , \6074_b1 , w_19268 );
or ( \6077_b0 , \6074_b0 , \6062_b0 );
not ( \6062_b0 , w_19269 );
and ( w_19269 , w_19268 , \6062_b1 );
buf ( \6078_b1 , \4072_b1 );
not ( \6078_b1 , w_19270 );
not ( \6078_b0 , w_19271 );
and ( w_19270 , w_19271 , \4072_b0 );
buf ( \6079_b1 , \4284_b1 );
not ( \6079_b1 , w_19272 );
not ( \6079_b0 , w_19273 );
and ( w_19272 , w_19273 , \4284_b0 );
or ( \6080_b1 , \6078_b1 , w_19274 );
or ( \6080_b0 , \6078_b0 , \6079_b0 );
not ( \6079_b0 , w_19275 );
and ( w_19275 , w_19274 , \6079_b1 );
or ( \6081_b1 , \4283_b1 , w_19277 );
not ( w_19277 , w_19278 );
and ( \6081_b0 , \4283_b0 , w_19279 );
and ( w_19278 ,  , w_19279 );
buf ( w_19277 , \5089_b1 );
not ( w_19277 , w_19280 );
not (  , w_19281 );
and ( w_19280 , w_19281 , \5089_b0 );
or ( \6082_b1 , \6080_b1 , w_19283 );
not ( w_19283 , w_19284 );
and ( \6082_b0 , \6080_b0 , w_19285 );
and ( w_19284 ,  , w_19285 );
buf ( w_19283 , \6081_b1 );
not ( w_19283 , w_19286 );
not (  , w_19287 );
and ( w_19286 , w_19287 , \6081_b0 );
buf ( \6083_b1 , \6082_b1 );
not ( \6083_b1 , w_19288 );
not ( \6083_b0 , w_19289 );
and ( w_19288 , w_19289 , \6082_b0 );
buf ( \6084_b1 , \4797_b1 );
not ( \6084_b1 , w_19290 );
not ( \6084_b0 , w_19291 );
and ( w_19290 , w_19291 , \4797_b0 );
or ( \6085_b1 , \6083_b1 , w_19292 );
or ( \6085_b0 , \6083_b0 , \6084_b0 );
not ( \6084_b0 , w_19293 );
and ( w_19293 , w_19292 , \6084_b1 );
buf ( \6086_b1 , \4267_b1 );
not ( \6086_b1 , w_19294 );
not ( \6086_b0 , w_19295 );
and ( w_19294 , w_19295 , \4267_b0 );
or ( \6087_b1 , \6086_b1 , w_19297 );
not ( w_19297 , w_19298 );
and ( \6087_b0 , \6086_b0 , w_19299 );
and ( w_19298 ,  , w_19299 );
buf ( w_19297 , \5951_b1 );
not ( w_19297 , w_19300 );
not (  , w_19301 );
and ( w_19300 , w_19301 , \5951_b0 );
or ( \6088_b1 , \6085_b1 , w_19303 );
not ( w_19303 , w_19304 );
and ( \6088_b0 , \6085_b0 , w_19305 );
and ( w_19304 ,  , w_19305 );
buf ( w_19303 , \6087_b1 );
not ( w_19303 , w_19306 );
not (  , w_19307 );
and ( w_19306 , w_19307 , \6087_b0 );
or ( \6089_b1 , \6077_b1 , w_19309 );
not ( w_19309 , w_19310 );
and ( \6089_b0 , \6077_b0 , w_19311 );
and ( w_19310 ,  , w_19311 );
buf ( w_19309 , \6088_b1 );
not ( w_19309 , w_19312 );
not (  , w_19313 );
and ( w_19312 , w_19313 , \6088_b0 );
or ( \6090_b1 , \6076_b1 , w_19315 );
not ( w_19315 , w_19316 );
and ( \6090_b0 , \6076_b0 , w_19317 );
and ( w_19316 ,  , w_19317 );
buf ( w_19315 , \6089_b1 );
not ( w_19315 , w_19318 );
not (  , w_19319 );
and ( w_19318 , w_19319 , \6089_b0 );
buf ( \6091_b1 , \6090_b1 );
not ( \6091_b1 , w_19320 );
not ( \6091_b0 , w_19321 );
and ( w_19320 , w_19321 , \6090_b0 );
or ( \6092_b1 , \6052_b1 , w_19322 );
or ( \6092_b0 , \6052_b0 , \6091_b0 );
not ( \6091_b0 , w_19323 );
and ( w_19323 , w_19322 , \6091_b1 );
or ( \6093_b1 , \6051_b1 , w_19324 );
or ( \6093_b0 , \6051_b0 , \6090_b0 );
not ( \6090_b0 , w_19325 );
and ( w_19325 , w_19324 , \6090_b1 );
buf ( \6094_b1 , \4079_b1 );
not ( \6094_b1 , w_19326 );
not ( \6094_b0 , w_19327 );
and ( w_19326 , w_19327 , \4079_b0 );
buf ( \6095_b1 , \4163_b1 );
not ( \6095_b1 , w_19328 );
not ( \6095_b0 , w_19329 );
and ( w_19328 , w_19329 , \4163_b0 );
or ( \6096_b1 , \6094_b1 , w_19330 );
or ( \6096_b0 , \6094_b0 , \6095_b0 );
not ( \6095_b0 , w_19331 );
and ( w_19331 , w_19330 , \6095_b1 );
or ( \6097_b1 , \4170_b1 , w_19333 );
not ( w_19333 , w_19334 );
and ( \6097_b0 , \4170_b0 , w_19335 );
and ( w_19334 ,  , w_19335 );
buf ( w_19333 , \5535_b1 );
not ( w_19333 , w_19336 );
not (  , w_19337 );
and ( w_19336 , w_19337 , \5535_b0 );
or ( \6098_b1 , \6096_b1 , w_19339 );
not ( w_19339 , w_19340 );
and ( \6098_b0 , \6096_b0 , w_19341 );
and ( w_19340 ,  , w_19341 );
buf ( w_19339 , \6097_b1 );
not ( w_19339 , w_19342 );
not (  , w_19343 );
and ( w_19342 , w_19343 , \6097_b0 );
buf ( \6099_b1 , \6098_b1 );
not ( \6099_b1 , w_19344 );
not ( \6099_b0 , w_19345 );
and ( w_19344 , w_19345 , \6098_b0 );
buf ( \6100_b1 , \4159_b1 );
not ( \6100_b1 , w_19346 );
not ( \6100_b0 , w_19347 );
and ( w_19346 , w_19347 , \4159_b0 );
or ( \6101_b1 , \6099_b1 , w_19348 );
or ( \6101_b0 , \6099_b0 , \6100_b0 );
not ( \6100_b0 , w_19349 );
and ( w_19349 , w_19348 , \6100_b1 );
or ( \6102_b1 , \6007_b1 , w_19351 );
not ( w_19351 , w_19352 );
and ( \6102_b0 , \6007_b0 , w_19353 );
and ( w_19352 ,  , w_19353 );
buf ( w_19351 , \4317_b1 );
not ( w_19351 , w_19354 );
not (  , w_19355 );
and ( w_19354 , w_19355 , \4317_b0 );
or ( \6103_b1 , \6101_b1 , w_19357 );
not ( w_19357 , w_19358 );
and ( \6103_b0 , \6101_b0 , w_19359 );
and ( w_19358 ,  , w_19359 );
buf ( w_19357 , \6102_b1 );
not ( w_19357 , w_19360 );
not (  , w_19361 );
and ( w_19360 , w_19361 , \6102_b0 );
buf ( \6104_b1 , \4066_b1 );
not ( \6104_b1 , w_19362 );
not ( \6104_b0 , w_19363 );
and ( w_19362 , w_19363 , \4066_b0 );
buf ( \6105_b1 , \5138_b1 );
not ( \6105_b1 , w_19364 );
not ( \6105_b0 , w_19365 );
and ( w_19364 , w_19365 , \5138_b0 );
or ( \6106_b1 , \6104_b1 , w_19366 );
or ( \6106_b0 , \6104_b0 , \6105_b0 );
not ( \6105_b0 , w_19367 );
and ( w_19367 , w_19366 , \6105_b1 );
or ( \6107_b1 , \4616_b1 , w_19369 );
not ( w_19369 , w_19370 );
and ( \6107_b0 , \4616_b0 , w_19371 );
and ( w_19370 ,  , w_19371 );
buf ( w_19369 , \4519_b1 );
not ( w_19369 , w_19372 );
not (  , w_19373 );
and ( w_19372 , w_19373 , \4519_b0 );
or ( \6108_b1 , \6106_b1 , w_19375 );
not ( w_19375 , w_19376 );
and ( \6108_b0 , \6106_b0 , w_19377 );
and ( w_19376 ,  , w_19377 );
buf ( w_19375 , \6107_b1 );
not ( w_19375 , w_19378 );
not (  , w_19379 );
and ( w_19378 , w_19379 , \6107_b0 );
buf ( \6109_b1 , \6108_b1 );
not ( \6109_b1 , w_19380 );
not ( \6109_b0 , w_19381 );
and ( w_19380 , w_19381 , \6108_b0 );
buf ( \6110_b1 , \4611_b1 );
not ( \6110_b1 , w_19382 );
not ( \6110_b0 , w_19383 );
and ( w_19382 , w_19383 , \4611_b0 );
or ( \6111_b1 , \6109_b1 , w_19384 );
or ( \6111_b0 , \6109_b0 , \6110_b0 );
not ( \6110_b0 , w_19385 );
and ( w_19385 , w_19384 , \6110_b1 );
or ( \6112_b1 , \5924_b1 , w_19387 );
not ( w_19387 , w_19388 );
and ( \6112_b0 , \5924_b0 , w_19389 );
and ( w_19388 ,  , w_19389 );
buf ( w_19387 , \4881_b1 );
not ( w_19387 , w_19390 );
not (  , w_19391 );
and ( w_19390 , w_19391 , \4881_b0 );
or ( \6113_b1 , \6111_b1 , w_19393 );
not ( w_19393 , w_19394 );
and ( \6113_b0 , \6111_b0 , w_19395 );
and ( w_19394 ,  , w_19395 );
buf ( w_19393 , \6112_b1 );
not ( w_19393 , w_19396 );
not (  , w_19397 );
and ( w_19396 , w_19397 , \6112_b0 );
or ( \6114_b1 , \6103_b1 , w_19398 );
or ( \6114_b0 , \6103_b0 , \6113_b0 );
not ( \6113_b0 , w_19399 );
and ( w_19399 , w_19398 , \6113_b1 );
buf ( \6115_b1 , \4098_b1 );
not ( \6115_b1 , w_19400 );
not ( \6115_b0 , w_19401 );
and ( w_19400 , w_19401 , \4098_b0 );
buf ( \6116_b1 , \4206_b1 );
not ( \6116_b1 , w_19402 );
not ( \6116_b0 , w_19403 );
and ( w_19402 , w_19403 , \4206_b0 );
or ( \6117_b1 , \6115_b1 , w_19404 );
or ( \6117_b0 , \6115_b0 , \6116_b0 );
not ( \6116_b0 , w_19405 );
and ( w_19405 , w_19404 , \6116_b1 );
or ( \6118_b1 , \4110_b1 , w_19407 );
not ( w_19407 , w_19408 );
and ( \6118_b0 , \4110_b0 , w_19409 );
and ( w_19408 ,  , w_19409 );
buf ( w_19407 , \5418_b1 );
not ( w_19407 , w_19410 );
not (  , w_19411 );
and ( w_19410 , w_19411 , \5418_b0 );
or ( \6119_b1 , \6117_b1 , w_19413 );
not ( w_19413 , w_19414 );
and ( \6119_b0 , \6117_b0 , w_19415 );
and ( w_19414 ,  , w_19415 );
buf ( w_19413 , \6118_b1 );
not ( w_19413 , w_19416 );
not (  , w_19417 );
and ( w_19416 , w_19417 , \6118_b0 );
buf ( \6120_b1 , \6119_b1 );
not ( \6120_b1 , w_19418 );
not ( \6120_b0 , w_19419 );
and ( w_19418 , w_19419 , \6119_b0 );
buf ( \6121_b1 , \4710_b1 );
not ( \6121_b1 , w_19420 );
not ( \6121_b0 , w_19421 );
and ( w_19420 , w_19421 , \4710_b0 );
or ( \6122_b1 , \6120_b1 , w_19422 );
or ( \6122_b0 , \6120_b0 , \6121_b0 );
not ( \6121_b0 , w_19423 );
and ( w_19423 , w_19422 , \6121_b1 );
or ( \6123_b1 , \5994_b1 , w_19425 );
not ( w_19425 , w_19426 );
and ( \6123_b0 , \5994_b0 , w_19427 );
and ( w_19426 ,  , w_19427 );
buf ( w_19425 , \4654_b1 );
not ( w_19425 , w_19428 );
not (  , w_19429 );
and ( w_19428 , w_19429 , \4654_b0 );
or ( \6124_b1 , \6122_b1 , w_19431 );
not ( w_19431 , w_19432 );
and ( \6124_b0 , \6122_b0 , w_19433 );
and ( w_19432 ,  , w_19433 );
buf ( w_19431 , \6123_b1 );
not ( w_19431 , w_19434 );
not (  , w_19435 );
and ( w_19434 , w_19435 , \6123_b0 );
or ( \6125_b1 , \6114_b1 , w_19437 );
not ( w_19437 , w_19438 );
and ( \6125_b0 , \6114_b0 , w_19439 );
and ( w_19438 ,  , w_19439 );
buf ( w_19437 , \6124_b1 );
not ( w_19437 , w_19440 );
not (  , w_19441 );
and ( w_19440 , w_19441 , \6124_b0 );
or ( \6126_b1 , \6103_b1 , w_19443 );
not ( w_19443 , w_19444 );
and ( \6126_b0 , \6103_b0 , w_19445 );
and ( w_19444 ,  , w_19445 );
buf ( w_19443 , \6113_b1 );
not ( w_19443 , w_19446 );
not (  , w_19447 );
and ( w_19446 , w_19447 , \6113_b0 );
or ( \6127_b1 , \6125_b1 , w_19449 );
not ( w_19449 , w_19450 );
and ( \6127_b0 , \6125_b0 , w_19451 );
and ( w_19450 ,  , w_19451 );
buf ( w_19449 , \6126_b1 );
not ( w_19449 , w_19452 );
not (  , w_19453 );
and ( w_19452 , w_19453 , \6126_b0 );
or ( \6128_b1 , \6093_b1 , w_19455 );
not ( w_19455 , w_19456 );
and ( \6128_b0 , \6093_b0 , w_19457 );
and ( w_19456 ,  , w_19457 );
buf ( w_19455 , \6127_b1 );
not ( w_19455 , w_19458 );
not (  , w_19459 );
and ( w_19458 , w_19459 , \6127_b0 );
or ( \6129_b1 , \6092_b1 , w_19461 );
not ( w_19461 , w_19462 );
and ( \6129_b0 , \6092_b0 , w_19463 );
and ( w_19462 ,  , w_19463 );
buf ( w_19461 , \6128_b1 );
not ( w_19461 , w_19464 );
not (  , w_19465 );
and ( w_19464 , w_19465 , \6128_b0 );
or ( \6130_b1 , \6049_b1 , \6129_b1 );
xor ( \6130_b0 , \6049_b0 , w_19466 );
not ( w_19466 , w_19467 );
and ( w_19467 , \6129_b1 , \6129_b0 );
or ( \6131_b1 , \5885_b1 , \5913_b1 );
xor ( \6131_b0 , \5885_b0 , w_19468 );
not ( w_19468 , w_19469 );
and ( w_19469 , \5913_b1 , \5913_b0 );
or ( \6132_b1 , \6131_b1 , w_19470 );
xor ( \6132_b0 , \6131_b0 , w_19472 );
not ( w_19472 , w_19473 );
and ( w_19473 , w_19470 , w_19471 );
buf ( w_19470 , \5875_b1 );
not ( w_19470 , w_19474 );
not ( w_19471 , w_19475 );
and ( w_19474 , w_19475 , \5875_b0 );
or ( \6133_b1 , \6130_b1 , \6132_b1 );
not ( \6132_b1 , w_19476 );
and ( \6133_b0 , \6130_b0 , w_19477 );
and ( w_19476 , w_19477 , \6132_b0 );
or ( \6134_b1 , \6049_b1 , \6129_b1 );
not ( \6129_b1 , w_19478 );
and ( \6134_b0 , \6049_b0 , w_19479 );
and ( w_19478 , w_19479 , \6129_b0 );
or ( \6135_b1 , \6133_b1 , w_19480 );
or ( \6135_b0 , \6133_b0 , \6134_b0 );
not ( \6134_b0 , w_19481 );
and ( w_19481 , w_19480 , \6134_b1 );
or ( \6136_b1 , \6047_b1 , \6135_b1 );
xor ( \6136_b0 , \6047_b0 , w_19482 );
not ( w_19482 , w_19483 );
and ( w_19483 , \6135_b1 , \6135_b0 );
buf ( \6137_b1 , \5916_b1 );
not ( \6137_b1 , w_19484 );
not ( \6137_b0 , w_19485 );
and ( w_19484 , w_19485 , \5916_b0 );
buf ( \6138_b1 , \6021_b1 );
not ( \6138_b1 , w_19486 );
not ( \6138_b0 , w_19487 );
and ( w_19486 , w_19487 , \6021_b0 );
or ( \6139_b1 , \6137_b1 , w_19488 );
or ( \6139_b0 , \6137_b0 , \6138_b0 );
not ( \6138_b0 , w_19489 );
and ( w_19489 , w_19488 , \6138_b1 );
or ( \6140_b1 , \6020_b1 , w_19491 );
not ( w_19491 , w_19492 );
and ( \6140_b0 , \6020_b0 , w_19493 );
and ( w_19492 ,  , w_19493 );
buf ( w_19491 , \5917_b1 );
not ( w_19491 , w_19494 );
not (  , w_19495 );
and ( w_19494 , w_19495 , \5917_b0 );
or ( \6141_b1 , \6139_b1 , w_19497 );
not ( w_19497 , w_19498 );
and ( \6141_b0 , \6139_b0 , w_19499 );
and ( w_19498 ,  , w_19499 );
buf ( w_19497 , \6140_b1 );
not ( w_19497 , w_19500 );
not (  , w_19501 );
and ( w_19500 , w_19501 , \6140_b0 );
or ( \6142_b1 , \6141_b1 , \6028_b1 );
not ( \6028_b1 , w_19502 );
and ( \6142_b0 , \6141_b0 , w_19503 );
and ( w_19502 , w_19503 , \6028_b0 );
buf ( \6143_b1 , \6141_b1 );
not ( \6143_b1 , w_19504 );
not ( \6143_b0 , w_19505 );
and ( w_19504 , w_19505 , \6141_b0 );
buf ( \6144_b1 , \6028_b1 );
not ( \6144_b1 , w_19506 );
not ( \6144_b0 , w_19507 );
and ( w_19506 , w_19507 , \6028_b0 );
or ( \6145_b1 , \6143_b1 , \6144_b1 );
not ( \6144_b1 , w_19508 );
and ( \6145_b0 , \6143_b0 , w_19509 );
and ( w_19508 , w_19509 , \6144_b0 );
or ( \6146_b1 , \6142_b1 , w_19511 );
not ( w_19511 , w_19512 );
and ( \6146_b0 , \6142_b0 , w_19513 );
and ( w_19512 ,  , w_19513 );
buf ( w_19511 , \6145_b1 );
not ( w_19511 , w_19514 );
not (  , w_19515 );
and ( w_19514 , w_19515 , \6145_b0 );
or ( \6147_b1 , \6136_b1 , \6146_b1 );
not ( \6146_b1 , w_19516 );
and ( \6147_b0 , \6136_b0 , w_19517 );
and ( w_19516 , w_19517 , \6146_b0 );
or ( \6148_b1 , \6047_b1 , \6135_b1 );
not ( \6135_b1 , w_19518 );
and ( \6148_b0 , \6047_b0 , w_19519 );
and ( w_19518 , w_19519 , \6135_b0 );
or ( \6149_b1 , \6147_b1 , w_19520 );
or ( \6149_b0 , \6147_b0 , \6148_b0 );
not ( \6148_b0 , w_19521 );
and ( w_19521 , w_19520 , \6148_b1 );
buf ( \6150_b1 , \6149_b1 );
not ( \6150_b1 , w_19522 );
not ( \6150_b0 , w_19523 );
and ( w_19522 , w_19523 , \6149_b0 );
or ( \6151_b1 , \6045_b1 , w_19525 );
not ( w_19525 , w_19526 );
and ( \6151_b0 , \6045_b0 , w_19527 );
and ( w_19526 ,  , w_19527 );
buf ( w_19525 , \6150_b1 );
not ( w_19525 , w_19528 );
not (  , w_19529 );
and ( w_19528 , w_19529 , \6150_b0 );
or ( \6152_b1 , \6017_b1 , \5959_b1 );
not ( \5959_b1 , w_19530 );
and ( \6152_b0 , \6017_b0 , w_19531 );
and ( w_19530 , w_19531 , \5959_b0 );
buf ( \6153_b1 , \6017_b1 );
not ( \6153_b1 , w_19532 );
not ( \6153_b0 , w_19533 );
and ( w_19532 , w_19533 , \6017_b0 );
or ( \6154_b1 , \6153_b1 , \5960_b1 );
not ( \5960_b1 , w_19534 );
and ( \6154_b0 , \6153_b0 , w_19535 );
and ( w_19534 , w_19535 , \5960_b0 );
or ( \6155_b1 , \6152_b1 , w_19537 );
not ( w_19537 , w_19538 );
and ( \6155_b0 , \6152_b0 , w_19539 );
and ( w_19538 ,  , w_19539 );
buf ( w_19537 , \6154_b1 );
not ( w_19537 , w_19540 );
not (  , w_19541 );
and ( w_19540 , w_19541 , \6154_b0 );
buf ( \6156_b1 , \5970_b1 );
buf ( \6156_b0 , \5970_b0 );
buf ( \6157_b1 , \6156_b1 );
not ( \6157_b1 , w_19542 );
not ( \6157_b0 , w_19543 );
and ( w_19542 , w_19543 , \6156_b0 );
or ( \6158_b1 , \6155_b1 , \6157_b1 );
not ( \6157_b1 , w_19544 );
and ( \6158_b0 , \6155_b0 , w_19545 );
and ( w_19544 , w_19545 , \6157_b0 );
buf ( \6159_b1 , \6155_b1 );
not ( \6159_b1 , w_19546 );
not ( \6159_b0 , w_19547 );
and ( w_19546 , w_19547 , \6155_b0 );
or ( \6160_b1 , \6159_b1 , \6156_b1 );
not ( \6156_b1 , w_19548 );
and ( \6160_b0 , \6159_b0 , w_19549 );
and ( w_19548 , w_19549 , \6156_b0 );
or ( \6161_b1 , \6158_b1 , w_19551 );
not ( w_19551 , w_19552 );
and ( \6161_b0 , \6158_b0 , w_19553 );
and ( w_19552 ,  , w_19553 );
buf ( w_19551 , \6160_b1 );
not ( w_19551 , w_19554 );
not (  , w_19555 );
and ( w_19554 , w_19555 , \6160_b0 );
or ( \6162_b1 , \5987_b1 , \5980_b1 );
xor ( \6162_b0 , \5987_b0 , w_19556 );
not ( w_19556 , w_19557 );
and ( w_19557 , \5980_b1 , \5980_b0 );
buf ( \6163_b1 , \6162_b1 );
not ( \6163_b1 , w_19558 );
not ( \6163_b0 , w_19559 );
and ( w_19558 , w_19559 , \6162_b0 );
buf ( \6164_b1 , \4097_b1 );
not ( \6164_b1 , w_19560 );
not ( \6164_b0 , w_19561 );
and ( w_19560 , w_19561 , \4097_b0 );
buf ( \6165_b1 , \5422_b1 );
not ( \6165_b1 , w_19562 );
not ( \6165_b0 , w_19563 );
and ( w_19562 , w_19563 , \5422_b0 );
or ( \6166_b1 , \6164_b1 , w_19564 );
or ( \6166_b0 , \6164_b0 , \6165_b0 );
not ( \6165_b0 , w_19565 );
and ( w_19565 , w_19564 , \6165_b1 );
or ( \6167_b1 , \5268_b1 , w_19567 );
not ( w_19567 , w_19568 );
and ( \6167_b0 , \5268_b0 , w_19569 );
and ( w_19568 ,  , w_19569 );
buf ( w_19567 , \4254_b1 );
not ( w_19567 , w_19570 );
not (  , w_19571 );
and ( w_19570 , w_19571 , \4254_b0 );
or ( \6168_b1 , \6166_b1 , w_19573 );
not ( w_19573 , w_19574 );
and ( \6168_b0 , \6166_b0 , w_19575 );
and ( w_19574 ,  , w_19575 );
buf ( w_19573 , \6167_b1 );
not ( w_19573 , w_19576 );
not (  , w_19577 );
and ( w_19576 , w_19577 , \6167_b0 );
buf ( \6169_b1 , \6168_b1 );
not ( \6169_b1 , w_19578 );
not ( \6169_b0 , w_19579 );
and ( w_19578 , w_19579 , \6168_b0 );
buf ( \6170_b1 , \5270_b1 );
not ( \6170_b1 , w_19580 );
not ( \6170_b0 , w_19581 );
and ( w_19580 , w_19581 , \5270_b0 );
or ( \6171_b1 , \6169_b1 , w_19582 );
or ( \6171_b0 , \6169_b0 , \6170_b0 );
not ( \6170_b0 , w_19583 );
and ( w_19583 , w_19582 , \6170_b1 );
or ( \6172_b1 , \6058_b1 , w_19585 );
not ( w_19585 , w_19586 );
and ( \6172_b0 , \6058_b0 , w_19587 );
and ( w_19586 ,  , w_19587 );
buf ( w_19585 , \5266_b1 );
not ( w_19585 , w_19588 );
not (  , w_19589 );
and ( w_19588 , w_19589 , \5266_b0 );
or ( \6173_b1 , \6171_b1 , w_19591 );
not ( w_19591 , w_19592 );
and ( \6173_b0 , \6171_b0 , w_19593 );
and ( w_19592 ,  , w_19593 );
buf ( w_19591 , \6172_b1 );
not ( w_19591 , w_19594 );
not (  , w_19595 );
and ( w_19594 , w_19595 , \6172_b0 );
buf ( \6174_b1 , \6173_b1 );
not ( \6174_b1 , w_19596 );
not ( \6174_b0 , w_19597 );
and ( w_19596 , w_19597 , \6173_b0 );
or ( \6175_b1 , \4132_b1 , w_19599 );
not ( w_19599 , w_19600 );
and ( \6175_b0 , \4132_b0 , w_19601 );
and ( w_19600 ,  , w_19601 );
buf ( w_19599 , \4098_b1 );
not ( w_19599 , w_19602 );
not (  , w_19603 );
and ( w_19602 , w_19603 , \4098_b0 );
or ( \6176_b1 , \6174_b1 , w_19605 );
not ( w_19605 , w_19606 );
and ( \6176_b0 , \6174_b0 , w_19607 );
and ( w_19606 ,  , w_19607 );
buf ( w_19605 , \6175_b1 );
not ( w_19605 , w_19608 );
not (  , w_19609 );
and ( w_19608 , w_19609 , \6175_b0 );
buf ( \6177_b1 , \6176_b1 );
not ( \6177_b1 , w_19610 );
not ( \6177_b0 , w_19611 );
and ( w_19610 , w_19611 , \6176_b0 );
or ( \6178_b1 , \4866_b1 , \4095_b1 );
not ( \4095_b1 , w_19612 );
and ( \6178_b0 , \4866_b0 , w_19613 );
and ( w_19612 , w_19613 , \4095_b0 );
or ( \6179_b1 , \4934_b1 , \4391_b1 );
not ( \4391_b1 , w_19614 );
and ( \6179_b0 , \4934_b0 , w_19615 );
and ( w_19614 , w_19615 , \4391_b0 );
or ( \6180_b1 , \6178_b1 , w_19617 );
not ( w_19617 , w_19618 );
and ( \6180_b0 , \6178_b0 , w_19619 );
and ( w_19618 ,  , w_19619 );
buf ( w_19617 , \6179_b1 );
not ( w_19617 , w_19620 );
not (  , w_19621 );
and ( w_19620 , w_19621 , \6179_b0 );
buf ( \6181_b1 , \6180_b1 );
not ( \6181_b1 , w_19622 );
not ( \6181_b0 , w_19623 );
and ( w_19622 , w_19623 , \6180_b0 );
buf ( \6182_b1 , \6181_b1 );
not ( \6182_b1 , w_19624 );
not ( \6182_b0 , w_19625 );
and ( w_19624 , w_19625 , \6181_b0 );
buf ( \6183_b1 , \4944_b1 );
not ( \6183_b1 , w_19626 );
not ( \6183_b0 , w_19627 );
and ( w_19626 , w_19627 , \4944_b0 );
or ( \6184_b1 , \6182_b1 , w_19628 );
or ( \6184_b0 , \6182_b0 , \6183_b0 );
not ( \6183_b0 , w_19629 );
and ( w_19629 , w_19628 , \6183_b1 );
or ( \6185_b1 , \4863_b1 , w_19631 );
not ( w_19631 , w_19632 );
and ( \6185_b0 , \4863_b0 , w_19633 );
and ( w_19632 ,  , w_19633 );
buf ( w_19631 , \5978_b1 );
not ( w_19631 , w_19634 );
not (  , w_19635 );
and ( w_19634 , w_19635 , \5978_b0 );
or ( \6186_b1 , \6184_b1 , w_19637 );
not ( w_19637 , w_19638 );
and ( \6186_b0 , \6184_b0 , w_19639 );
and ( w_19638 ,  , w_19639 );
buf ( w_19637 , \6185_b1 );
not ( w_19637 , w_19640 );
not (  , w_19641 );
and ( w_19640 , w_19641 , \6185_b0 );
buf ( \6187_b1 , \6186_b1 );
not ( \6187_b1 , w_19642 );
not ( \6187_b0 , w_19643 );
and ( w_19642 , w_19643 , \6186_b0 );
or ( \6188_b1 , \6177_b1 , w_19644 );
or ( \6188_b0 , \6177_b0 , \6187_b0 );
not ( \6187_b0 , w_19645 );
and ( w_19645 , w_19644 , \6187_b1 );
buf ( \6189_b1 , \6175_b1 );
not ( \6189_b1 , w_19646 );
not ( \6189_b0 , w_19647 );
and ( w_19646 , w_19647 , \6175_b0 );
or ( \6190_b1 , \6189_b1 , w_19649 );
not ( w_19649 , w_19650 );
and ( \6190_b0 , \6189_b0 , w_19651 );
and ( w_19650 ,  , w_19651 );
buf ( w_19649 , \6173_b1 );
not ( w_19649 , w_19652 );
not (  , w_19653 );
and ( w_19652 , w_19653 , \6173_b0 );
or ( \6191_b1 , \6188_b1 , w_19655 );
not ( w_19655 , w_19656 );
and ( \6191_b0 , \6188_b0 , w_19657 );
and ( w_19656 ,  , w_19657 );
buf ( w_19655 , \6190_b1 );
not ( w_19655 , w_19658 );
not (  , w_19659 );
and ( w_19658 , w_19659 , \6190_b0 );
buf ( \6192_b1 , \6191_b1 );
not ( \6192_b1 , w_19660 );
not ( \6192_b0 , w_19661 );
and ( w_19660 , w_19661 , \6191_b0 );
or ( \6193_b1 , \6163_b1 , w_19663 );
not ( w_19663 , w_19664 );
and ( \6193_b0 , \6163_b0 , w_19665 );
and ( w_19664 ,  , w_19665 );
buf ( w_19663 , \6192_b1 );
not ( w_19663 , w_19666 );
not (  , w_19667 );
and ( w_19666 , w_19667 , \6192_b0 );
buf ( \6194_b1 , \6193_b1 );
not ( \6194_b1 , w_19668 );
not ( \6194_b0 , w_19669 );
and ( w_19668 , w_19669 , \6193_b0 );
buf ( \6195_b1 , \4449_b1 );
not ( \6195_b1 , w_19670 );
not ( \6195_b0 , w_19671 );
and ( w_19670 , w_19671 , \4449_b0 );
buf ( \6196_b1 , \4026_b1 );
not ( \6196_b1 , w_19672 );
not ( \6196_b0 , w_19673 );
and ( w_19672 , w_19673 , \4026_b0 );
buf ( \6197_b1 , \5112_b1 );
not ( \6197_b1 , w_19674 );
not ( \6197_b0 , w_19675 );
and ( w_19674 , w_19675 , \5112_b0 );
or ( \6198_b1 , \6196_b1 , w_19676 );
or ( \6198_b0 , \6196_b0 , \6197_b0 );
not ( \6197_b0 , w_19677 );
and ( w_19677 , w_19676 , \6197_b1 );
or ( \6199_b1 , \4729_b1 , w_19679 );
not ( w_19679 , w_19680 );
and ( \6199_b0 , \4729_b0 , w_19681 );
and ( w_19680 ,  , w_19681 );
buf ( w_19679 , \4969_b1 );
not ( w_19679 , w_19682 );
not (  , w_19683 );
and ( w_19682 , w_19683 , \4969_b0 );
or ( \6200_b1 , \6198_b1 , w_19685 );
not ( w_19685 , w_19686 );
and ( \6200_b0 , \6198_b0 , w_19687 );
and ( w_19686 ,  , w_19687 );
buf ( w_19685 , \6199_b1 );
not ( w_19685 , w_19688 );
not (  , w_19689 );
and ( w_19688 , w_19689 , \6199_b0 );
buf ( \6201_b1 , \6200_b1 );
not ( \6201_b1 , w_19690 );
not ( \6201_b0 , w_19691 );
and ( w_19690 , w_19691 , \6200_b0 );
or ( \6202_b1 , \6195_b1 , w_19692 );
or ( \6202_b0 , \6195_b0 , \6201_b0 );
not ( \6201_b0 , w_19693 );
and ( w_19693 , w_19692 , \6201_b1 );
or ( \6203_b1 , \4452_b1 , w_19695 );
not ( w_19695 , w_19696 );
and ( \6203_b0 , \4452_b0 , w_19697 );
and ( w_19696 ,  , w_19697 );
buf ( w_19695 , \6069_b1 );
not ( w_19695 , w_19698 );
not (  , w_19699 );
and ( w_19698 , w_19699 , \6069_b0 );
or ( \6204_b1 , \6202_b1 , w_19701 );
not ( w_19701 , w_19702 );
and ( \6204_b0 , \6202_b0 , w_19703 );
and ( w_19702 ,  , w_19703 );
buf ( w_19701 , \6203_b1 );
not ( w_19701 , w_19704 );
not (  , w_19705 );
and ( w_19704 , w_19705 , \6203_b0 );
buf ( \6205_b1 , \6204_b1 );
not ( \6205_b1 , w_19706 );
not ( \6205_b0 , w_19707 );
and ( w_19706 , w_19707 , \6204_b0 );
buf ( \6206_b1 , \6205_b1 );
not ( \6206_b1 , w_19708 );
not ( \6206_b0 , w_19709 );
and ( w_19708 , w_19709 , \6205_b0 );
buf ( \6207_b1 , \4082_b1 );
not ( \6207_b1 , w_19710 );
not ( \6207_b0 , w_19711 );
and ( w_19710 , w_19711 , \4082_b0 );
buf ( \6208_b1 , \4163_b1 );
not ( \6208_b1 , w_19712 );
not ( \6208_b0 , w_19713 );
and ( w_19712 , w_19713 , \4163_b0 );
or ( \6209_b1 , \6207_b1 , w_19714 );
or ( \6209_b0 , \6207_b0 , \6208_b0 );
not ( \6208_b0 , w_19715 );
and ( w_19715 , w_19714 , \6208_b1 );
or ( \6210_b1 , \4170_b1 , w_19717 );
not ( w_19717 , w_19718 );
and ( \6210_b0 , \4170_b0 , w_19719 );
and ( w_19718 ,  , w_19719 );
buf ( w_19717 , \5526_b1 );
not ( w_19717 , w_19720 );
not (  , w_19721 );
and ( w_19720 , w_19721 , \5526_b0 );
or ( \6211_b1 , \6209_b1 , w_19723 );
not ( w_19723 , w_19724 );
and ( \6211_b0 , \6209_b0 , w_19725 );
and ( w_19724 ,  , w_19725 );
buf ( w_19723 , \6210_b1 );
not ( w_19723 , w_19726 );
not (  , w_19727 );
and ( w_19726 , w_19727 , \6210_b0 );
buf ( \6212_b1 , \6211_b1 );
not ( \6212_b1 , w_19728 );
not ( \6212_b0 , w_19729 );
and ( w_19728 , w_19729 , \6211_b0 );
buf ( \6213_b1 , \4159_b1 );
not ( \6213_b1 , w_19730 );
not ( \6213_b0 , w_19731 );
and ( w_19730 , w_19731 , \4159_b0 );
or ( \6214_b1 , \6212_b1 , w_19732 );
or ( \6214_b0 , \6212_b0 , \6213_b0 );
not ( \6213_b0 , w_19733 );
and ( w_19733 , w_19732 , \6213_b1 );
or ( \6215_b1 , \4317_b1 , w_19735 );
not ( w_19735 , w_19736 );
and ( \6215_b0 , \4317_b0 , w_19737 );
and ( w_19736 ,  , w_19737 );
buf ( w_19735 , \6098_b1 );
not ( w_19735 , w_19738 );
not (  , w_19739 );
and ( w_19738 , w_19739 , \6098_b0 );
or ( \6216_b1 , \6214_b1 , w_19741 );
not ( w_19741 , w_19742 );
and ( \6216_b0 , \6214_b0 , w_19743 );
and ( w_19742 ,  , w_19743 );
buf ( w_19741 , \6215_b1 );
not ( w_19741 , w_19744 );
not (  , w_19745 );
and ( w_19744 , w_19745 , \6215_b0 );
buf ( \6217_b1 , \6216_b1 );
not ( \6217_b1 , w_19746 );
not ( \6217_b0 , w_19747 );
and ( w_19746 , w_19747 , \6216_b0 );
buf ( \6218_b1 , \6217_b1 );
not ( \6218_b1 , w_19748 );
not ( \6218_b0 , w_19749 );
and ( w_19748 , w_19749 , \6217_b0 );
or ( \6219_b1 , \6206_b1 , w_19750 );
or ( \6219_b0 , \6206_b0 , \6218_b0 );
not ( \6218_b0 , w_19751 );
and ( w_19751 , w_19750 , \6218_b1 );
buf ( \6220_b1 , \4076_b1 );
not ( \6220_b1 , w_19752 );
not ( \6220_b0 , w_19753 );
and ( w_19752 , w_19753 , \4076_b0 );
buf ( \6221_b1 , \4493_b1 );
not ( \6221_b1 , w_19754 );
not ( \6221_b0 , w_19755 );
and ( w_19754 , w_19755 , \4493_b0 );
or ( \6222_b1 , \6220_b1 , w_19756 );
or ( \6222_b0 , \6220_b0 , \6221_b0 );
not ( \6221_b0 , w_19757 );
and ( w_19757 , w_19756 , \6221_b1 );
or ( \6223_b1 , \4283_b1 , w_19759 );
not ( w_19759 , w_19760 );
and ( \6223_b0 , \4283_b0 , w_19761 );
and ( w_19760 ,  , w_19761 );
buf ( w_19759 , \5284_b1 );
not ( w_19759 , w_19762 );
not (  , w_19763 );
and ( w_19762 , w_19763 , \5284_b0 );
or ( \6224_b1 , \6222_b1 , w_19765 );
not ( w_19765 , w_19766 );
and ( \6224_b0 , \6222_b0 , w_19767 );
and ( w_19766 ,  , w_19767 );
buf ( w_19765 , \6223_b1 );
not ( w_19765 , w_19768 );
not (  , w_19769 );
and ( w_19768 , w_19769 , \6223_b0 );
buf ( \6225_b1 , \6224_b1 );
not ( \6225_b1 , w_19770 );
not ( \6225_b0 , w_19771 );
and ( w_19770 , w_19771 , \6224_b0 );
buf ( \6226_b1 , \4797_b1 );
not ( \6226_b1 , w_19772 );
not ( \6226_b0 , w_19773 );
and ( w_19772 , w_19773 , \4797_b0 );
or ( \6227_b1 , \6225_b1 , w_19774 );
or ( \6227_b0 , \6225_b0 , \6226_b0 );
not ( \6226_b0 , w_19775 );
and ( w_19775 , w_19774 , \6226_b1 );
or ( \6228_b1 , \6082_b1 , w_19777 );
not ( w_19777 , w_19778 );
and ( \6228_b0 , \6082_b0 , w_19779 );
and ( w_19778 ,  , w_19779 );
buf ( w_19777 , \4800_b1 );
not ( w_19777 , w_19780 );
not (  , w_19781 );
and ( w_19780 , w_19781 , \4800_b0 );
or ( \6229_b1 , \6227_b1 , w_19783 );
not ( w_19783 , w_19784 );
and ( \6229_b0 , \6227_b0 , w_19785 );
and ( w_19784 ,  , w_19785 );
buf ( w_19783 , \6228_b1 );
not ( w_19783 , w_19786 );
not (  , w_19787 );
and ( w_19786 , w_19787 , \6228_b0 );
or ( \6230_b1 , \6219_b1 , w_19789 );
not ( w_19789 , w_19790 );
and ( \6230_b0 , \6219_b0 , w_19791 );
and ( w_19790 ,  , w_19791 );
buf ( w_19789 , \6229_b1 );
not ( w_19789 , w_19792 );
not (  , w_19793 );
and ( w_19792 , w_19793 , \6229_b0 );
or ( \6231_b1 , \6204_b1 , w_19795 );
not ( w_19795 , w_19796 );
and ( \6231_b0 , \6204_b0 , w_19797 );
and ( w_19796 ,  , w_19797 );
buf ( w_19795 , \6216_b1 );
not ( w_19795 , w_19798 );
not (  , w_19799 );
and ( w_19798 , w_19799 , \6216_b0 );
or ( \6232_b1 , \6230_b1 , w_19801 );
not ( w_19801 , w_19802 );
and ( \6232_b0 , \6230_b0 , w_19803 );
and ( w_19802 ,  , w_19803 );
buf ( w_19801 , \6231_b1 );
not ( w_19801 , w_19804 );
not (  , w_19805 );
and ( w_19804 , w_19805 , \6231_b0 );
buf ( \6233_b1 , \6232_b1 );
not ( \6233_b1 , w_19806 );
not ( \6233_b0 , w_19807 );
and ( w_19806 , w_19807 , \6232_b0 );
or ( \6234_b1 , \6194_b1 , w_19808 );
or ( \6234_b0 , \6194_b0 , \6233_b0 );
not ( \6233_b0 , w_19809 );
and ( w_19809 , w_19808 , \6233_b1 );
or ( \6235_b1 , \6191_b1 , w_19811 );
not ( w_19811 , w_19812 );
and ( \6235_b0 , \6191_b0 , w_19813 );
and ( w_19812 ,  , w_19813 );
buf ( w_19811 , \6162_b1 );
not ( w_19811 , w_19814 );
not (  , w_19815 );
and ( w_19814 , w_19815 , \6162_b0 );
or ( \6236_b1 , \6234_b1 , w_19817 );
not ( w_19817 , w_19818 );
and ( \6236_b0 , \6234_b0 , w_19819 );
and ( w_19818 ,  , w_19819 );
buf ( w_19817 , \6235_b1 );
not ( w_19817 , w_19820 );
not (  , w_19821 );
and ( w_19820 , w_19821 , \6235_b0 );
buf ( \6237_b1 , \6236_b1 );
not ( \6237_b1 , w_19822 );
not ( \6237_b0 , w_19823 );
and ( w_19822 , w_19823 , \6236_b0 );
buf ( \6238_b1 , \5940_b1 );
not ( \6238_b1 , w_19824 );
not ( \6238_b0 , w_19825 );
and ( w_19824 , w_19825 , \5940_b0 );
buf ( \6239_b1 , \6238_b1 );
not ( \6239_b1 , w_19826 );
not ( \6239_b0 , w_19827 );
and ( w_19826 , w_19827 , \6238_b0 );
buf ( \6240_b1 , \5928_b1 );
not ( \6240_b1 , w_19828 );
not ( \6240_b0 , w_19829 );
and ( w_19828 , w_19829 , \5928_b0 );
buf ( \6241_b1 , \5957_b1 );
not ( \6241_b1 , w_19830 );
not ( \6241_b0 , w_19831 );
and ( w_19830 , w_19831 , \5957_b0 );
buf ( \6242_b1 , \6241_b1 );
not ( \6242_b1 , w_19832 );
not ( \6242_b0 , w_19833 );
and ( w_19832 , w_19833 , \6241_b0 );
or ( \6243_b1 , \6240_b1 , w_19834 );
or ( \6243_b0 , \6240_b0 , \6242_b0 );
not ( \6242_b0 , w_19835 );
and ( w_19835 , w_19834 , \6242_b1 );
or ( \6244_b1 , \5928_b1 , w_19836 );
or ( \6244_b0 , \5928_b0 , \6241_b0 );
not ( \6241_b0 , w_19837 );
and ( w_19837 , w_19836 , \6241_b1 );
or ( \6245_b1 , \6243_b1 , w_19839 );
not ( w_19839 , w_19840 );
and ( \6245_b0 , \6243_b0 , w_19841 );
and ( w_19840 ,  , w_19841 );
buf ( w_19839 , \6244_b1 );
not ( w_19839 , w_19842 );
not (  , w_19843 );
and ( w_19842 , w_19843 , \6244_b0 );
buf ( \6246_b1 , \6245_b1 );
not ( \6246_b1 , w_19844 );
not ( \6246_b0 , w_19845 );
and ( w_19844 , w_19845 , \6245_b0 );
or ( \6247_b1 , \6239_b1 , w_19846 );
or ( \6247_b0 , \6239_b0 , \6246_b0 );
not ( \6246_b0 , w_19847 );
and ( w_19847 , w_19846 , \6246_b1 );
buf ( \6248_b1 , \6245_b1 );
not ( \6248_b1 , w_19848 );
not ( \6248_b0 , w_19849 );
and ( w_19848 , w_19849 , \6245_b0 );
buf ( \6249_b1 , \6238_b1 );
not ( \6249_b1 , w_19850 );
not ( \6249_b0 , w_19851 );
and ( w_19850 , w_19851 , \6238_b0 );
or ( \6250_b1 , \6248_b1 , w_19853 );
not ( w_19853 , w_19854 );
and ( \6250_b0 , \6248_b0 , w_19855 );
and ( w_19854 ,  , w_19855 );
buf ( w_19853 , \6249_b1 );
not ( w_19853 , w_19856 );
not (  , w_19857 );
and ( w_19856 , w_19857 , \6249_b0 );
or ( \6251_b1 , \6247_b1 , w_19859 );
not ( w_19859 , w_19860 );
and ( \6251_b0 , \6247_b0 , w_19861 );
and ( w_19860 ,  , w_19861 );
buf ( w_19859 , \6250_b1 );
not ( w_19859 , w_19862 );
not (  , w_19863 );
and ( w_19862 , w_19863 , \6250_b0 );
buf ( \6252_b1 , \6251_b1 );
not ( \6252_b1 , w_19864 );
not ( \6252_b0 , w_19865 );
and ( w_19864 , w_19865 , \6251_b0 );
or ( \6253_b1 , \5988_b1 , \5999_b1 );
not ( \5999_b1 , w_19866 );
and ( \6253_b0 , \5988_b0 , w_19867 );
and ( w_19866 , w_19867 , \5999_b0 );
buf ( \6254_b1 , \5988_b1 );
not ( \6254_b1 , w_19868 );
not ( \6254_b0 , w_19869 );
and ( w_19868 , w_19869 , \5988_b0 );
or ( \6255_b1 , \6254_b1 , \6000_b1 );
not ( \6000_b1 , w_19870 );
and ( \6255_b0 , \6254_b0 , w_19871 );
and ( w_19870 , w_19871 , \6000_b0 );
or ( \6256_b1 , \6253_b1 , w_19872 );
or ( \6256_b0 , \6253_b0 , \6255_b0 );
not ( \6255_b0 , w_19873 );
and ( w_19873 , w_19872 , \6255_b1 );
buf ( \6257_b1 , \6013_b1 );
not ( \6257_b1 , w_19874 );
not ( \6257_b0 , w_19875 );
and ( w_19874 , w_19875 , \6013_b0 );
or ( \6258_b1 , \6256_b1 , \6257_b1 );
not ( \6257_b1 , w_19876 );
and ( \6258_b0 , \6256_b0 , w_19877 );
and ( w_19876 , w_19877 , \6257_b0 );
buf ( \6259_b1 , \6256_b1 );
not ( \6259_b1 , w_19878 );
not ( \6259_b0 , w_19879 );
and ( w_19878 , w_19879 , \6256_b0 );
or ( \6260_b1 , \6259_b1 , \6013_b1 );
not ( \6013_b1 , w_19880 );
and ( \6260_b0 , \6259_b0 , w_19881 );
and ( w_19880 , w_19881 , \6013_b0 );
or ( \6261_b1 , \6258_b1 , w_19883 );
not ( w_19883 , w_19884 );
and ( \6261_b0 , \6258_b0 , w_19885 );
and ( w_19884 ,  , w_19885 );
buf ( w_19883 , \6260_b1 );
not ( w_19883 , w_19886 );
not (  , w_19887 );
and ( w_19886 , w_19887 , \6260_b0 );
or ( \6262_b1 , \6252_b1 , w_19889 );
not ( w_19889 , w_19890 );
and ( \6262_b0 , \6252_b0 , w_19891 );
and ( w_19890 ,  , w_19891 );
buf ( w_19889 , \6261_b1 );
not ( w_19889 , w_19892 );
not (  , w_19893 );
and ( w_19892 , w_19893 , \6261_b0 );
buf ( \6263_b1 , \6262_b1 );
not ( \6263_b1 , w_19894 );
not ( \6263_b0 , w_19895 );
and ( w_19894 , w_19895 , \6262_b0 );
or ( \6264_b1 , \6237_b1 , w_19896 );
or ( \6264_b0 , \6237_b0 , \6263_b0 );
not ( \6263_b0 , w_19897 );
and ( w_19897 , w_19896 , \6263_b1 );
buf ( \6265_b1 , \6261_b1 );
not ( \6265_b1 , w_19898 );
not ( \6265_b0 , w_19899 );
and ( w_19898 , w_19899 , \6261_b0 );
or ( \6266_b1 , \6265_b1 , w_19901 );
not ( w_19901 , w_19902 );
and ( \6266_b0 , \6265_b0 , w_19903 );
and ( w_19902 ,  , w_19903 );
buf ( w_19901 , \6251_b1 );
not ( w_19901 , w_19904 );
not (  , w_19905 );
and ( w_19904 , w_19905 , \6251_b0 );
or ( \6267_b1 , \6264_b1 , w_19907 );
not ( w_19907 , w_19908 );
and ( \6267_b0 , \6264_b0 , w_19909 );
and ( w_19908 ,  , w_19909 );
buf ( w_19907 , \6266_b1 );
not ( w_19907 , w_19910 );
not (  , w_19911 );
and ( w_19910 , w_19911 , \6266_b0 );
or ( \6268_b1 , \6161_b1 , \6267_b1 );
xor ( \6268_b0 , \6161_b0 , w_19912 );
not ( w_19912 , w_19913 );
and ( w_19913 , \6267_b1 , \6267_b0 );
or ( \6269_b1 , \6049_b1 , \6129_b1 );
xor ( \6269_b0 , \6049_b0 , w_19914 );
not ( w_19914 , w_19915 );
and ( w_19915 , \6129_b1 , \6129_b0 );
or ( \6270_b1 , \6269_b1 , \6132_b1 );
xor ( \6270_b0 , \6269_b0 , w_19916 );
not ( w_19916 , w_19917 );
and ( w_19917 , \6132_b1 , \6132_b0 );
or ( \6271_b1 , \6268_b1 , \6270_b1 );
not ( \6270_b1 , w_19918 );
and ( \6271_b0 , \6268_b0 , w_19919 );
and ( w_19918 , w_19919 , \6270_b0 );
or ( \6272_b1 , \6161_b1 , \6267_b1 );
not ( \6267_b1 , w_19920 );
and ( \6272_b0 , \6161_b0 , w_19921 );
and ( w_19920 , w_19921 , \6267_b0 );
or ( \6273_b1 , \6271_b1 , w_19922 );
or ( \6273_b0 , \6271_b0 , \6272_b0 );
not ( \6272_b0 , w_19923 );
and ( w_19923 , w_19922 , \6272_b1 );
buf ( \6274_b1 , \6273_b1 );
not ( \6274_b1 , w_19924 );
not ( \6274_b0 , w_19925 );
and ( w_19924 , w_19925 , \6273_b0 );
or ( \6275_b1 , \6047_b1 , \6135_b1 );
xor ( \6275_b0 , \6047_b0 , w_19926 );
not ( w_19926 , w_19927 );
and ( w_19927 , \6135_b1 , \6135_b0 );
or ( \6276_b1 , \6275_b1 , \6146_b1 );
xor ( \6276_b0 , \6275_b0 , w_19928 );
not ( w_19928 , w_19929 );
and ( w_19929 , \6146_b1 , \6146_b0 );
buf ( \6277_b1 , \6276_b1 );
not ( \6277_b1 , w_19930 );
not ( \6277_b0 , w_19931 );
and ( w_19930 , w_19931 , \6276_b0 );
or ( \6278_b1 , \6274_b1 , w_19933 );
not ( w_19933 , w_19934 );
and ( \6278_b0 , \6274_b0 , w_19935 );
and ( w_19934 ,  , w_19935 );
buf ( w_19933 , \6277_b1 );
not ( w_19933 , w_19936 );
not (  , w_19937 );
and ( w_19936 , w_19937 , \6277_b0 );
or ( \6279_b1 , \6151_b1 , \6278_b1 );
not ( \6278_b1 , w_19938 );
and ( \6279_b0 , \6151_b0 , w_19939 );
and ( w_19938 , w_19939 , \6278_b0 );
or ( \6280_b1 , \5653_b1 , \5691_b1 );
xor ( \6280_b0 , \5653_b0 , w_19940 );
not ( w_19940 , w_19941 );
and ( w_19941 , \5691_b1 , \5691_b0 );
or ( \6281_b1 , \6280_b1 , \5702_b1 );
xor ( \6281_b0 , \6280_b0 , w_19942 );
not ( w_19942 , w_19943 );
and ( w_19943 , \5702_b1 , \5702_b0 );
buf ( \6282_b1 , \5721_b1 );
not ( \6282_b1 , w_19944 );
not ( \6282_b0 , w_19945 );
and ( w_19944 , w_19945 , \5721_b0 );
or ( \6283_b1 , \5847_b1 , w_19947 );
not ( w_19947 , w_19948 );
and ( \6283_b0 , \5847_b0 , w_19949 );
and ( w_19948 ,  , w_19949 );
buf ( w_19947 , \6282_b1 );
not ( w_19947 , w_19950 );
not (  , w_19951 );
and ( w_19950 , w_19951 , \6282_b0 );
buf ( \6284_b1 , \5840_b1 );
not ( \6284_b1 , w_19952 );
not ( \6284_b0 , w_19953 );
and ( w_19952 , w_19953 , \5840_b0 );
or ( \6285_b1 , \6283_b1 , \6284_b1 );
not ( \6284_b1 , w_19954 );
and ( \6285_b0 , \6283_b0 , w_19955 );
and ( w_19954 , w_19955 , \6284_b0 );
or ( \6286_b1 , \5847_b1 , w_19957 );
not ( w_19957 , w_19958 );
and ( \6286_b0 , \5847_b0 , w_19959 );
and ( w_19958 ,  , w_19959 );
buf ( w_19957 , \6282_b1 );
not ( w_19957 , w_19960 );
not (  , w_19961 );
and ( w_19960 , w_19961 , \6282_b0 );
or ( \6287_b1 , \6285_b1 , w_19963 );
not ( w_19963 , w_19964 );
and ( \6287_b0 , \6285_b0 , w_19965 );
and ( w_19964 ,  , w_19965 );
buf ( w_19963 , \6286_b1 );
not ( w_19963 , w_19966 );
not (  , w_19967 );
and ( w_19966 , w_19967 , \6286_b0 );
or ( \6288_b1 , \6281_b1 , w_19969 );
not ( w_19969 , w_19970 );
and ( \6288_b0 , \6281_b0 , w_19971 );
and ( w_19970 ,  , w_19971 );
buf ( w_19969 , \6287_b1 );
not ( w_19969 , w_19972 );
not (  , w_19973 );
and ( w_19972 , w_19973 , \6287_b0 );
buf ( \6290_b1 , \6289_b1 );
not ( \6290_b1 , w_19974 );
not ( \6290_b0 , w_19975 );
and ( w_19974 , w_19975 , \6289_b0 );
buf ( \6291_b1 , \4082_b1 );
not ( \6291_b1 , w_19976 );
not ( \6291_b0 , w_19977 );
and ( w_19976 , w_19977 , \4082_b0 );
buf ( \6292_b1 , \5301_b1 );
not ( \6292_b1 , w_19978 );
not ( \6292_b0 , w_19979 );
and ( w_19978 , w_19979 , \5301_b0 );
or ( \6293_b1 , \6291_b1 , w_19980 );
or ( \6293_b0 , \6291_b0 , \6292_b0 );
not ( \6292_b0 , w_19981 );
and ( w_19981 , w_19980 , \6292_b1 );
or ( \6294_b1 , \4616_b1 , w_19983 );
not ( w_19983 , w_19984 );
and ( \6294_b0 , \4616_b0 , w_19985 );
and ( w_19984 ,  , w_19985 );
buf ( w_19983 , \5526_b1 );
not ( w_19983 , w_19986 );
not (  , w_19987 );
and ( w_19986 , w_19987 , \5526_b0 );
or ( \6295_b1 , \6293_b1 , w_19989 );
not ( w_19989 , w_19990 );
and ( \6295_b0 , \6293_b0 , w_19991 );
and ( w_19990 ,  , w_19991 );
buf ( w_19989 , \6294_b1 );
not ( w_19989 , w_19992 );
not (  , w_19993 );
and ( w_19992 , w_19993 , \6294_b0 );
buf ( \6296_b1 , \6295_b1 );
not ( \6296_b1 , w_19994 );
not ( \6296_b0 , w_19995 );
and ( w_19994 , w_19995 , \6295_b0 );
buf ( \6297_b1 , \4611_b1 );
not ( \6297_b1 , w_19996 );
not ( \6297_b0 , w_19997 );
and ( w_19996 , w_19997 , \4611_b0 );
or ( \6298_b1 , \6296_b1 , w_19998 );
or ( \6298_b0 , \6296_b0 , \6297_b0 );
not ( \6297_b0 , w_19999 );
and ( w_19999 , w_19998 , \6297_b1 );
buf ( \6299_b1 , \4079_b1 );
not ( \6299_b1 , w_20000 );
not ( \6299_b0 , w_20001 );
and ( w_20000 , w_20001 , \4079_b0 );
buf ( \6300_b1 , \5301_b1 );
not ( \6300_b1 , w_20002 );
not ( \6300_b0 , w_20003 );
and ( w_20002 , w_20003 , \5301_b0 );
or ( \6301_b1 , \6299_b1 , w_20004 );
or ( \6301_b0 , \6299_b0 , \6300_b0 );
not ( \6300_b0 , w_20005 );
and ( w_20005 , w_20004 , \6300_b1 );
buf ( \6302_b1 , \5138_b1 );
not ( \6302_b1 , w_20006 );
not ( \6302_b0 , w_20007 );
and ( w_20006 , w_20007 , \5138_b0 );
or ( \6303_b1 , \6302_b1 , w_20009 );
not ( w_20009 , w_20010 );
and ( \6303_b0 , \6302_b0 , w_20011 );
and ( w_20010 ,  , w_20011 );
buf ( w_20009 , \5535_b1 );
not ( w_20009 , w_20012 );
not (  , w_20013 );
and ( w_20012 , w_20013 , \5535_b0 );
or ( \6304_b1 , \6301_b1 , w_20015 );
not ( w_20015 , w_20016 );
and ( \6304_b0 , \6301_b0 , w_20017 );
and ( w_20016 ,  , w_20017 );
buf ( w_20015 , \6303_b1 );
not ( w_20015 , w_20018 );
not (  , w_20019 );
and ( w_20018 , w_20019 , \6303_b0 );
or ( \6305_b1 , \6304_b1 , w_20021 );
not ( w_20021 , w_20022 );
and ( \6305_b0 , \6304_b0 , w_20023 );
and ( w_20022 ,  , w_20023 );
buf ( w_20021 , \5146_b1 );
not ( w_20021 , w_20024 );
not (  , w_20025 );
and ( w_20024 , w_20025 , \5146_b0 );
or ( \6306_b1 , \6298_b1 , w_20027 );
not ( w_20027 , w_20028 );
and ( \6306_b0 , \6298_b0 , w_20029 );
and ( w_20028 ,  , w_20029 );
buf ( w_20027 , \6305_b1 );
not ( w_20027 , w_20030 );
not (  , w_20031 );
and ( w_20030 , w_20031 , \6305_b0 );
buf ( \6307_b1 , \6306_b1 );
not ( \6307_b1 , w_20032 );
not ( \6307_b0 , w_20033 );
and ( w_20032 , w_20033 , \6306_b0 );
buf ( \6308_b1 , \4079_b1 );
not ( \6308_b1 , w_20034 );
not ( \6308_b0 , w_20035 );
and ( w_20034 , w_20035 , \4079_b0 );
buf ( \6309_b1 , \4939_b1 );
not ( \6309_b1 , w_20036 );
not ( \6309_b0 , w_20037 );
and ( w_20036 , w_20037 , \4939_b0 );
or ( \6310_b1 , \6308_b1 , w_20038 );
or ( \6310_b0 , \6308_b0 , \6309_b0 );
not ( \6309_b0 , w_20039 );
and ( w_20039 , w_20038 , \6309_b1 );
or ( \6311_b1 , \4936_b1 , w_20041 );
not ( w_20041 , w_20042 );
and ( \6311_b0 , \4936_b0 , w_20043 );
and ( w_20042 ,  , w_20043 );
buf ( w_20041 , \5535_b1 );
not ( w_20041 , w_20044 );
not (  , w_20045 );
and ( w_20044 , w_20045 , \5535_b0 );
or ( \6312_b1 , \6310_b1 , w_20047 );
not ( w_20047 , w_20048 );
and ( \6312_b0 , \6310_b0 , w_20049 );
and ( w_20048 ,  , w_20049 );
buf ( w_20047 , \6311_b1 );
not ( w_20047 , w_20050 );
not (  , w_20051 );
and ( w_20050 , w_20051 , \6311_b0 );
buf ( \6313_b1 , \6312_b1 );
not ( \6313_b1 , w_20052 );
not ( \6313_b0 , w_20053 );
and ( w_20052 , w_20053 , \6312_b0 );
buf ( \6314_b1 , \4945_b1 );
not ( \6314_b1 , w_20054 );
not ( \6314_b0 , w_20055 );
and ( w_20054 , w_20055 , \4945_b0 );
or ( \6315_b1 , \6313_b1 , w_20056 );
or ( \6315_b0 , \6313_b0 , \6314_b0 );
not ( \6314_b0 , w_20057 );
and ( w_20057 , w_20056 , \6314_b1 );
or ( \6316_b1 , \4076_b1 , \4949_b1 );
not ( \4949_b1 , w_20058 );
and ( \6316_b0 , \4076_b0 , w_20059 );
and ( w_20058 , w_20059 , \4949_b0 );
buf ( \6317_b1 , \4076_b1 );
not ( \6317_b1 , w_20060 );
not ( \6317_b0 , w_20061 );
and ( w_20060 , w_20061 , \4076_b0 );
or ( \6318_b1 , \6317_b1 , \4935_b1 );
not ( \4935_b1 , w_20062 );
and ( \6318_b0 , \6317_b0 , w_20063 );
and ( w_20062 , w_20063 , \4935_b0 );
or ( \6319_b1 , \6316_b1 , w_20065 );
not ( w_20065 , w_20066 );
and ( \6319_b0 , \6316_b0 , w_20067 );
and ( w_20066 ,  , w_20067 );
buf ( w_20065 , \6318_b1 );
not ( w_20065 , w_20068 );
not (  , w_20069 );
and ( w_20068 , w_20069 , \6318_b0 );
or ( \6320_b1 , \4948_b1 , w_20071 );
not ( w_20071 , w_20072 );
and ( \6320_b0 , \4948_b0 , w_20073 );
and ( w_20072 ,  , w_20073 );
buf ( w_20071 , \6319_b1 );
not ( w_20071 , w_20074 );
not (  , w_20075 );
and ( w_20074 , w_20075 , \6319_b0 );
or ( \6321_b1 , \6315_b1 , w_20077 );
not ( w_20077 , w_20078 );
and ( \6321_b0 , \6315_b0 , w_20079 );
and ( w_20078 ,  , w_20079 );
buf ( w_20077 , \6320_b1 );
not ( w_20077 , w_20080 );
not (  , w_20081 );
and ( w_20080 , w_20081 , \6320_b0 );
buf ( \6322_b1 , \5418_b1 );
not ( \6322_b1 , w_20082 );
not ( \6322_b0 , w_20083 );
and ( w_20082 , w_20083 , \5418_b0 );
buf ( \6323_b1 , \4597_b1 );
not ( \6323_b1 , w_20084 );
not ( \6323_b0 , w_20085 );
and ( w_20084 , w_20085 , \4597_b0 );
or ( \6324_b1 , \6322_b1 , w_20086 );
or ( \6324_b0 , \6322_b0 , \6323_b0 );
not ( \6323_b0 , w_20087 );
and ( w_20087 , w_20086 , \6323_b1 );
or ( \6325_b1 , \6324_b1 , w_20089 );
not ( w_20089 , w_20090 );
and ( \6325_b0 , \6324_b0 , w_20091 );
and ( w_20090 ,  , w_20091 );
buf ( w_20089 , \4868_b1 );
not ( w_20089 , w_20092 );
not (  , w_20093 );
and ( w_20092 , w_20093 , \4868_b0 );
or ( \6326_b1 , \3516_b1 , w_20095 );
not ( w_20095 , w_20096 );
and ( \6326_b0 , \3516_b0 , w_20097 );
and ( w_20096 ,  , w_20097 );
buf ( w_20095 , \4098_b1 );
not ( w_20095 , w_20098 );
not (  , w_20099 );
and ( w_20098 , w_20099 , \4098_b0 );
or ( \6328_b1 , \6321_b1 , w_20101 );
not ( w_20101 , w_20102 );
and ( \6328_b0 , \6321_b0 , w_20103 );
and ( w_20102 ,  , w_20103 );
buf ( w_20101 , \6327_b1 );
not ( w_20101 , w_20104 );
not (  , w_20105 );
and ( w_20104 , w_20105 , \6327_b0 );
or ( \6329_b1 , \6307_b1 , w_20107 );
not ( w_20107 , w_20108 );
and ( \6329_b0 , \6307_b0 , w_20109 );
and ( w_20108 ,  , w_20109 );
buf ( w_20107 , \6328_b1 );
not ( w_20107 , w_20110 );
not (  , w_20111 );
and ( w_20110 , w_20111 , \6328_b0 );
buf ( \6330_b1 , \6329_b1 );
not ( \6330_b1 , w_20112 );
not ( \6330_b0 , w_20113 );
and ( w_20112 , w_20113 , \6329_b0 );
buf ( \6331_b1 , \4026_b1 );
not ( \6331_b1 , w_20114 );
not ( \6331_b0 , w_20115 );
and ( w_20114 , w_20115 , \4026_b0 );
buf ( \6332_b1 , \5274_b1 );
not ( \6332_b1 , w_20116 );
not ( \6332_b0 , w_20117 );
and ( w_20116 , w_20117 , \5274_b0 );
or ( \6333_b1 , \6331_b1 , w_20118 );
or ( \6333_b0 , \6331_b0 , \6332_b0 );
not ( \6332_b0 , w_20119 );
and ( w_20119 , w_20118 , \6332_b1 );
or ( \6334_b1 , \5425_b1 , w_20121 );
not ( w_20121 , w_20122 );
and ( \6334_b0 , \5425_b0 , w_20123 );
and ( w_20122 ,  , w_20123 );
buf ( w_20121 , \4969_b1 );
not ( w_20121 , w_20124 );
not (  , w_20125 );
and ( w_20124 , w_20125 , \4969_b0 );
or ( \6335_b1 , \6333_b1 , w_20127 );
not ( w_20127 , w_20128 );
and ( \6335_b0 , \6333_b0 , w_20129 );
and ( w_20128 ,  , w_20129 );
buf ( w_20127 , \6334_b1 );
not ( w_20127 , w_20130 );
not (  , w_20131 );
and ( w_20130 , w_20131 , \6334_b0 );
buf ( \6336_b1 , \6335_b1 );
not ( \6336_b1 , w_20132 );
not ( \6336_b0 , w_20133 );
and ( w_20132 , w_20133 , \6335_b0 );
buf ( \6337_b1 , \5272_b1 );
not ( \6337_b1 , w_20134 );
not ( \6337_b0 , w_20135 );
and ( w_20134 , w_20135 , \5272_b0 );
buf ( \6338_b1 , \6337_b1 );
not ( \6338_b1 , w_20136 );
not ( \6338_b0 , w_20137 );
and ( w_20136 , w_20137 , \6337_b0 );
or ( \6339_b1 , \6336_b1 , w_20138 );
or ( \6339_b0 , \6336_b0 , \6338_b0 );
not ( \6338_b0 , w_20139 );
and ( w_20139 , w_20138 , \6338_b1 );
buf ( \6340_b1 , \4021_b1 );
not ( \6340_b1 , w_20140 );
not ( \6340_b0 , w_20141 );
and ( w_20140 , w_20141 , \4021_b0 );
buf ( \6341_b1 , \5274_b1 );
not ( \6341_b1 , w_20142 );
not ( \6341_b0 , w_20143 );
and ( w_20142 , w_20143 , \5274_b0 );
or ( \6342_b1 , \6340_b1 , w_20144 );
or ( \6342_b0 , \6340_b0 , \6341_b0 );
not ( \6341_b0 , w_20145 );
and ( w_20145 , w_20144 , \6341_b1 );
or ( \6343_b1 , \5425_b1 , w_20147 );
not ( w_20147 , w_20148 );
and ( \6343_b0 , \5425_b0 , w_20149 );
and ( w_20148 ,  , w_20149 );
buf ( w_20147 , \4780_b1 );
not ( w_20147 , w_20150 );
not (  , w_20151 );
and ( w_20150 , w_20151 , \4780_b0 );
or ( \6344_b1 , \6342_b1 , w_20153 );
not ( w_20153 , w_20154 );
and ( \6344_b0 , \6342_b0 , w_20155 );
and ( w_20154 ,  , w_20155 );
buf ( w_20153 , \6343_b1 );
not ( w_20153 , w_20156 );
not (  , w_20157 );
and ( w_20156 , w_20157 , \6343_b0 );
or ( \6345_b1 , \6344_b1 , w_20159 );
not ( w_20159 , w_20160 );
and ( \6345_b0 , \6344_b0 , w_20161 );
and ( w_20160 ,  , w_20161 );
buf ( w_20159 , \5266_b1 );
not ( w_20159 , w_20162 );
not (  , w_20163 );
and ( w_20162 , w_20163 , \5266_b0 );
or ( \6346_b1 , \6339_b1 , w_20165 );
not ( w_20165 , w_20166 );
and ( \6346_b0 , \6339_b0 , w_20167 );
and ( w_20166 ,  , w_20167 );
buf ( w_20165 , \6345_b1 );
not ( w_20165 , w_20168 );
not (  , w_20169 );
and ( w_20168 , w_20169 , \6345_b0 );
or ( \6347_b1 , \4454_b1 , w_20171 );
not ( w_20171 , w_20172 );
and ( \6347_b0 , \4454_b0 , w_20173 );
and ( w_20172 ,  , w_20173 );
buf ( w_20171 , \5418_b1 );
not ( w_20171 , w_20174 );
not (  , w_20175 );
and ( w_20174 , w_20175 , \5418_b0 );
or ( \6348_b1 , \6346_b1 , \6347_b1 );
xor ( \6348_b0 , \6346_b0 , w_20176 );
not ( w_20176 , w_20177 );
and ( w_20177 , \6347_b1 , \6347_b0 );
buf ( \6349_b1 , \4945_b1 );
not ( \6349_b1 , w_20178 );
not ( \6349_b0 , w_20179 );
and ( w_20178 , w_20179 , \4945_b0 );
buf ( \6350_b1 , \6319_b1 );
not ( \6350_b1 , w_20180 );
not ( \6350_b0 , w_20181 );
and ( w_20180 , w_20181 , \6319_b0 );
or ( \6351_b1 , \6349_b1 , w_20182 );
or ( \6351_b0 , \6349_b0 , \6350_b0 );
not ( \6350_b0 , w_20183 );
and ( w_20183 , w_20182 , \6350_b1 );
buf ( \6352_b1 , \4072_b1 );
not ( \6352_b1 , w_20184 );
not ( \6352_b0 , w_20185 );
and ( w_20184 , w_20185 , \4072_b0 );
buf ( \6353_b1 , \4869_b1 );
not ( \6353_b1 , w_20186 );
not ( \6353_b0 , w_20187 );
and ( w_20186 , w_20187 , \4869_b0 );
or ( \6354_b1 , \6352_b1 , w_20188 );
or ( \6354_b0 , \6352_b0 , \6353_b0 );
not ( \6353_b0 , w_20189 );
and ( w_20189 , w_20188 , \6353_b1 );
or ( \6355_b1 , \4868_b1 , w_20191 );
not ( w_20191 , w_20192 );
and ( \6355_b0 , \4868_b0 , w_20193 );
and ( w_20192 ,  , w_20193 );
buf ( w_20191 , \5089_b1 );
not ( w_20191 , w_20194 );
not (  , w_20195 );
and ( w_20194 , w_20195 , \5089_b0 );
or ( \6356_b1 , \6354_b1 , w_20197 );
not ( w_20197 , w_20198 );
and ( \6356_b0 , \6354_b0 , w_20199 );
and ( w_20198 ,  , w_20199 );
buf ( w_20197 , \6355_b1 );
not ( w_20197 , w_20200 );
not (  , w_20201 );
and ( w_20200 , w_20201 , \6355_b0 );
or ( \6357_b1 , \4948_b1 , w_20203 );
not ( w_20203 , w_20204 );
and ( \6357_b0 , \4948_b0 , w_20205 );
and ( w_20204 ,  , w_20205 );
buf ( w_20203 , \6356_b1 );
not ( w_20203 , w_20206 );
not (  , w_20207 );
and ( w_20206 , w_20207 , \6356_b0 );
or ( \6358_b1 , \6351_b1 , w_20209 );
not ( w_20209 , w_20210 );
and ( \6358_b0 , \6351_b0 , w_20211 );
and ( w_20210 ,  , w_20211 );
buf ( w_20209 , \6357_b1 );
not ( w_20209 , w_20212 );
not (  , w_20213 );
and ( w_20212 , w_20213 , \6357_b0 );
or ( \6359_b1 , \6348_b1 , \6358_b1 );
xor ( \6359_b0 , \6348_b0 , w_20214 );
not ( w_20214 , w_20215 );
and ( w_20215 , \6358_b1 , \6358_b0 );
buf ( \6360_b1 , \6359_b1 );
not ( \6360_b1 , w_20216 );
not ( \6360_b0 , w_20217 );
and ( w_20216 , w_20217 , \6359_b0 );
or ( \6361_b1 , \6330_b1 , w_20218 );
or ( \6361_b0 , \6330_b0 , \6360_b0 );
not ( \6360_b0 , w_20219 );
and ( w_20219 , w_20218 , \6360_b1 );
buf ( \6362_b1 , \6328_b1 );
not ( \6362_b1 , w_20220 );
not ( \6362_b0 , w_20221 );
and ( w_20220 , w_20221 , \6328_b0 );
or ( \6363_b1 , \6362_b1 , w_20223 );
not ( w_20223 , w_20224 );
and ( \6363_b0 , \6362_b0 , w_20225 );
and ( w_20224 ,  , w_20225 );
buf ( w_20223 , \6306_b1 );
not ( w_20223 , w_20226 );
not (  , w_20227 );
and ( w_20226 , w_20227 , \6306_b0 );
or ( \6364_b1 , \6361_b1 , w_20229 );
not ( w_20229 , w_20230 );
and ( \6364_b0 , \6361_b0 , w_20231 );
and ( w_20230 ,  , w_20231 );
buf ( w_20229 , \6363_b1 );
not ( w_20229 , w_20232 );
not (  , w_20233 );
and ( w_20232 , w_20233 , \6363_b0 );
or ( \6365_b1 , \4437_b1 , w_20235 );
not ( w_20235 , w_20236 );
and ( \6365_b0 , \4437_b0 , w_20237 );
and ( w_20236 ,  , w_20237 );
buf ( w_20235 , \5418_b1 );
not ( w_20235 , w_20238 );
not (  , w_20239 );
and ( w_20238 , w_20239 , \5418_b0 );
or ( \6366_b1 , \4616_b1 , \6365_b1 );
not ( \6365_b1 , w_20240 );
and ( \6366_b0 , \4616_b0 , w_20241 );
and ( w_20240 , w_20241 , \6365_b0 );
buf ( \6367_b1 , \4098_b1 );
not ( \6367_b1 , w_20242 );
not ( \6367_b0 , w_20243 );
and ( w_20242 , w_20243 , \4098_b0 );
buf ( \6368_b1 , \4437_b1 );
not ( \6368_b1 , w_20244 );
not ( \6368_b0 , w_20245 );
and ( w_20244 , w_20245 , \4437_b0 );
buf ( \6369_b1 , \6368_b1 );
not ( \6369_b1 , w_20246 );
not ( \6369_b0 , w_20247 );
and ( w_20246 , w_20247 , \6368_b0 );
or ( \6370_b1 , \6367_b1 , w_20248 );
or ( \6370_b0 , \6367_b0 , \6369_b0 );
not ( \6369_b0 , w_20249 );
and ( w_20249 , w_20248 , \6369_b1 );
or ( \6371_b1 , \6370_b1 , w_20251 );
not ( w_20251 , w_20252 );
and ( \6371_b0 , \6370_b0 , w_20253 );
and ( w_20252 ,  , w_20253 );
buf ( w_20251 , \4729_b1 );
not ( w_20251 , w_20254 );
not (  , w_20255 );
and ( w_20254 , w_20255 , \4729_b0 );
or ( \6372_b1 , \6366_b1 , w_20257 );
not ( w_20257 , w_20258 );
and ( \6372_b0 , \6366_b0 , w_20259 );
and ( w_20258 ,  , w_20259 );
buf ( w_20257 , \6371_b1 );
not ( w_20257 , w_20260 );
not (  , w_20261 );
and ( w_20260 , w_20261 , \6371_b0 );
buf ( \6373_b1 , \6372_b1 );
not ( \6373_b1 , w_20262 );
not ( \6373_b0 , w_20263 );
and ( w_20262 , w_20263 , \6372_b0 );
buf ( \6374_b1 , \6373_b1 );
not ( \6374_b1 , w_20264 );
not ( \6374_b0 , w_20265 );
and ( w_20264 , w_20265 , \6373_b0 );
buf ( \6375_b1 , \6356_b1 );
not ( \6375_b1 , w_20266 );
not ( \6375_b0 , w_20267 );
and ( w_20266 , w_20267 , \6356_b0 );
buf ( \6376_b1 , \4945_b1 );
not ( \6376_b1 , w_20268 );
not ( \6376_b0 , w_20269 );
and ( w_20268 , w_20269 , \4945_b0 );
or ( \6377_b1 , \6375_b1 , w_20270 );
or ( \6377_b0 , \6375_b0 , \6376_b0 );
not ( \6376_b0 , w_20271 );
and ( w_20271 , w_20270 , \6376_b1 );
buf ( \6378_b1 , \4026_b1 );
not ( \6378_b1 , w_20272 );
not ( \6378_b0 , w_20273 );
and ( w_20272 , w_20273 , \4026_b0 );
buf ( \6379_b1 , \4935_b1 );
not ( \6379_b1 , w_20274 );
not ( \6379_b0 , w_20275 );
and ( w_20274 , w_20275 , \4935_b0 );
or ( \6380_b1 , \6378_b1 , w_20276 );
or ( \6380_b0 , \6378_b0 , \6379_b0 );
not ( \6379_b0 , w_20277 );
and ( w_20277 , w_20276 , \6379_b1 );
or ( \6381_b1 , \2945_b1 , w_20279 );
not ( w_20279 , w_20280 );
and ( \6381_b0 , \2945_b0 , w_20281 );
and ( w_20280 ,  , w_20281 );
buf ( w_20279 , \4969_b1 );
not ( w_20279 , w_20282 );
not (  , w_20283 );
and ( w_20282 , w_20283 , \4969_b0 );
or ( \6382_b1 , \6380_b1 , w_20285 );
not ( w_20285 , w_20286 );
and ( \6382_b0 , \6380_b0 , w_20287 );
and ( w_20286 ,  , w_20287 );
buf ( w_20285 , \6381_b1 );
not ( w_20285 , w_20288 );
not (  , w_20289 );
and ( w_20288 , w_20289 , \6381_b0 );
or ( \6383_b1 , \4863_b1 , w_20291 );
not ( w_20291 , w_20292 );
and ( \6383_b0 , \4863_b0 , w_20293 );
and ( w_20292 ,  , w_20293 );
buf ( w_20291 , \6382_b1 );
not ( w_20291 , w_20294 );
not (  , w_20295 );
and ( w_20294 , w_20295 , \6382_b0 );
or ( \6384_b1 , \6377_b1 , w_20297 );
not ( w_20297 , w_20298 );
and ( \6384_b0 , \6377_b0 , w_20299 );
and ( w_20298 ,  , w_20299 );
buf ( w_20297 , \6383_b1 );
not ( w_20297 , w_20300 );
not (  , w_20301 );
and ( w_20300 , w_20301 , \6383_b0 );
buf ( \6385_b1 , \6384_b1 );
not ( \6385_b1 , w_20302 );
not ( \6385_b0 , w_20303 );
and ( w_20302 , w_20303 , \6384_b0 );
or ( \6386_b1 , \6374_b1 , w_20304 );
or ( \6386_b0 , \6374_b0 , \6385_b0 );
not ( \6385_b0 , w_20305 );
and ( w_20305 , w_20304 , \6385_b1 );
or ( \6387_b1 , \6384_b1 , w_20306 );
or ( \6387_b0 , \6384_b0 , \6373_b0 );
not ( \6373_b0 , w_20307 );
and ( w_20307 , w_20306 , \6373_b1 );
or ( \6388_b1 , \6386_b1 , w_20309 );
not ( w_20309 , w_20310 );
and ( \6388_b0 , \6386_b0 , w_20311 );
and ( w_20310 ,  , w_20311 );
buf ( w_20309 , \6387_b1 );
not ( w_20309 , w_20312 );
not (  , w_20313 );
and ( w_20312 , w_20313 , \6387_b0 );
or ( \6389_b1 , \6346_b1 , \6347_b1 );
xor ( \6389_b0 , \6346_b0 , w_20314 );
not ( w_20314 , w_20315 );
and ( w_20315 , \6347_b1 , \6347_b0 );
or ( \6390_b1 , \6389_b1 , \6358_b1 );
not ( \6358_b1 , w_20316 );
and ( \6390_b0 , \6389_b0 , w_20317 );
and ( w_20316 , w_20317 , \6358_b0 );
or ( \6391_b1 , \6346_b1 , \6347_b1 );
not ( \6347_b1 , w_20318 );
and ( \6391_b0 , \6346_b0 , w_20319 );
and ( w_20318 , w_20319 , \6347_b0 );
or ( \6392_b1 , \6390_b1 , w_20320 );
or ( \6392_b0 , \6390_b0 , \6391_b0 );
not ( \6391_b0 , w_20321 );
and ( w_20321 , w_20320 , \6391_b1 );
or ( \6393_b1 , \6388_b1 , \6392_b1 );
xor ( \6393_b0 , \6388_b0 , w_20322 );
not ( w_20322 , w_20323 );
and ( w_20323 , \6392_b1 , \6392_b0 );
buf ( \6394_b1 , \6344_b1 );
not ( \6394_b1 , w_20324 );
not ( \6394_b0 , w_20325 );
and ( w_20324 , w_20325 , \6344_b0 );
buf ( \6395_b1 , \6337_b1 );
not ( \6395_b1 , w_20326 );
not ( \6395_b0 , w_20327 );
and ( w_20326 , w_20327 , \6337_b0 );
or ( \6396_b1 , \6394_b1 , w_20328 );
or ( \6396_b0 , \6394_b0 , \6395_b0 );
not ( \6395_b0 , w_20329 );
and ( w_20329 , w_20328 , \6395_b1 );
buf ( \6397_b1 , \4017_b1 );
not ( \6397_b1 , w_20330 );
not ( \6397_b0 , w_20331 );
and ( w_20330 , w_20331 , \4017_b0 );
buf ( \6398_b1 , \5422_b1 );
not ( \6398_b1 , w_20332 );
not ( \6398_b0 , w_20333 );
and ( w_20332 , w_20333 , \5422_b0 );
or ( \6399_b1 , \6397_b1 , w_20334 );
or ( \6399_b0 , \6397_b0 , \6398_b0 );
not ( \6398_b0 , w_20335 );
and ( w_20335 , w_20334 , \6398_b1 );
or ( \6400_b1 , \4662_b1 , w_20337 );
not ( w_20337 , w_20338 );
and ( \6400_b0 , \4662_b0 , w_20339 );
and ( w_20338 ,  , w_20339 );
buf ( w_20337 , \5275_b1 );
not ( w_20337 , w_20340 );
not (  , w_20341 );
and ( w_20340 , w_20341 , \5275_b0 );
or ( \6401_b1 , \6399_b1 , w_20343 );
not ( w_20343 , w_20344 );
and ( \6401_b0 , \6399_b0 , w_20345 );
and ( w_20344 ,  , w_20345 );
buf ( w_20343 , \6400_b1 );
not ( w_20343 , w_20346 );
not (  , w_20347 );
and ( w_20346 , w_20347 , \6400_b0 );
or ( \6402_b1 , \6401_b1 , w_20349 );
not ( w_20349 , w_20350 );
and ( \6402_b0 , \6401_b0 , w_20351 );
and ( w_20350 ,  , w_20351 );
buf ( w_20349 , \5266_b1 );
not ( w_20349 , w_20352 );
not (  , w_20353 );
and ( w_20352 , w_20353 , \5266_b0 );
or ( \6403_b1 , \6396_b1 , w_20355 );
not ( w_20355 , w_20356 );
and ( \6403_b0 , \6396_b0 , w_20357 );
and ( w_20356 ,  , w_20357 );
buf ( w_20355 , \6402_b1 );
not ( w_20355 , w_20358 );
not (  , w_20359 );
and ( w_20358 , w_20359 , \6402_b0 );
buf ( \6404_b1 , \6304_b1 );
not ( \6404_b1 , w_20360 );
not ( \6404_b0 , w_20361 );
and ( w_20360 , w_20361 , \6304_b0 );
buf ( \6405_b1 , \4611_b1 );
not ( \6405_b1 , w_20362 );
not ( \6405_b0 , w_20363 );
and ( w_20362 , w_20363 , \4611_b0 );
or ( \6406_b1 , \6404_b1 , w_20364 );
or ( \6406_b0 , \6404_b0 , \6405_b0 );
not ( \6405_b0 , w_20365 );
and ( w_20365 , w_20364 , \6405_b1 );
or ( \6407_b1 , \4076_b1 , \4616_b1 );
not ( \4616_b1 , w_20366 );
and ( \6407_b0 , \4076_b0 , w_20367 );
and ( w_20366 , w_20367 , \4616_b0 );
buf ( \6408_b1 , \4076_b1 );
not ( \6408_b1 , w_20368 );
not ( \6408_b0 , w_20369 );
and ( w_20368 , w_20369 , \4076_b0 );
or ( \6409_b1 , \6408_b1 , \5138_b1 );
not ( \5138_b1 , w_20370 );
and ( \6409_b0 , \6408_b0 , w_20371 );
and ( w_20370 , w_20371 , \5138_b0 );
or ( \6410_b1 , \6407_b1 , w_20373 );
not ( w_20373 , w_20374 );
and ( \6410_b0 , \6407_b0 , w_20375 );
and ( w_20374 ,  , w_20375 );
buf ( w_20373 , \6409_b1 );
not ( w_20373 , w_20376 );
not (  , w_20377 );
and ( w_20376 , w_20377 , \6409_b0 );
or ( \6411_b1 , \6410_b1 , w_20379 );
not ( w_20379 , w_20380 );
and ( \6411_b0 , \6410_b0 , w_20381 );
and ( w_20380 ,  , w_20381 );
buf ( w_20379 , \4754_b1 );
not ( w_20379 , w_20382 );
not (  , w_20383 );
and ( w_20382 , w_20383 , \4754_b0 );
or ( \6412_b1 , \6406_b1 , w_20385 );
not ( w_20385 , w_20386 );
and ( \6412_b0 , \6406_b0 , w_20387 );
and ( w_20386 ,  , w_20387 );
buf ( w_20385 , \6411_b1 );
not ( w_20385 , w_20388 );
not (  , w_20389 );
and ( w_20388 , w_20389 , \6411_b0 );
or ( \6413_b1 , \6403_b1 , \6412_b1 );
xor ( \6413_b0 , \6403_b0 , w_20390 );
not ( w_20390 , w_20391 );
and ( w_20391 , \6412_b1 , \6412_b0 );
or ( \6414_b1 , \4098_b1 , \4532_b1 );
not ( \4532_b1 , w_20392 );
and ( \6414_b0 , \4098_b0 , w_20393 );
and ( w_20392 , w_20393 , \4532_b0 );
buf ( \6415_b1 , \4098_b1 );
not ( \6415_b1 , w_20394 );
not ( \6415_b0 , w_20395 );
and ( w_20394 , w_20395 , \4098_b0 );
or ( \6416_b1 , \6415_b1 , \4458_b1 );
not ( \4458_b1 , w_20396 );
and ( \6416_b0 , \6415_b0 , w_20397 );
and ( w_20396 , w_20397 , \4458_b0 );
or ( \6417_b1 , \6414_b1 , w_20399 );
not ( w_20399 , w_20400 );
and ( \6417_b0 , \6414_b0 , w_20401 );
and ( w_20400 ,  , w_20401 );
buf ( w_20399 , \6416_b1 );
not ( w_20399 , w_20402 );
not (  , w_20403 );
and ( w_20402 , w_20403 , \6416_b0 );
buf ( \6418_b1 , \4632_b1 );
not ( \6418_b1 , w_20404 );
not ( \6418_b0 , w_20405 );
and ( w_20404 , w_20405 , \4632_b0 );
or ( \6419_b1 , \6417_b1 , w_20406 );
or ( \6419_b0 , \6417_b0 , \6418_b0 );
not ( \6418_b0 , w_20407 );
and ( w_20407 , w_20406 , \6418_b1 );
or ( \6420_b1 , \4082_b1 , \4917_b1 );
not ( \4917_b1 , w_20408 );
and ( \6420_b0 , \4082_b0 , w_20409 );
and ( w_20408 , w_20409 , \4917_b0 );
buf ( \6421_b1 , \4082_b1 );
not ( \6421_b1 , w_20410 );
not ( \6421_b0 , w_20411 );
and ( w_20410 , w_20411 , \4082_b0 );
or ( \6422_b1 , \6421_b1 , \4535_b1 );
not ( \4535_b1 , w_20412 );
and ( \6422_b0 , \6421_b0 , w_20413 );
and ( w_20412 , w_20413 , \4535_b0 );
or ( \6423_b1 , \6420_b1 , w_20415 );
not ( w_20415 , w_20416 );
and ( \6423_b0 , \6420_b0 , w_20417 );
and ( w_20416 ,  , w_20417 );
buf ( w_20415 , \6422_b1 );
not ( w_20415 , w_20418 );
not (  , w_20419 );
and ( w_20418 , w_20419 , \6422_b0 );
buf ( \6424_b1 , \6423_b1 );
not ( \6424_b1 , w_20420 );
not ( \6424_b0 , w_20421 );
and ( w_20420 , w_20421 , \6423_b0 );
or ( \6425_b1 , \4454_b1 , w_20422 );
or ( \6425_b0 , \4454_b0 , \6424_b0 );
not ( \6424_b0 , w_20423 );
and ( w_20423 , w_20422 , \6424_b1 );
or ( \6426_b1 , \6419_b1 , w_20425 );
not ( w_20425 , w_20426 );
and ( \6426_b0 , \6419_b0 , w_20427 );
and ( w_20426 ,  , w_20427 );
buf ( w_20425 , \6425_b1 );
not ( w_20425 , w_20428 );
not (  , w_20429 );
and ( w_20428 , w_20429 , \6425_b0 );
or ( \6427_b1 , \6413_b1 , \6426_b1 );
xor ( \6427_b0 , \6413_b0 , w_20430 );
not ( w_20430 , w_20431 );
and ( w_20431 , \6426_b1 , \6426_b0 );
or ( \6428_b1 , \6393_b1 , \6427_b1 );
xor ( \6428_b0 , \6393_b0 , w_20432 );
not ( w_20432 , w_20433 );
and ( w_20433 , \6427_b1 , \6427_b0 );
or ( \6429_b1 , \6364_b1 , \6428_b1 );
xor ( \6429_b0 , \6364_b0 , w_20434 );
not ( w_20434 , w_20435 );
and ( w_20435 , \6428_b1 , \6428_b0 );
buf ( \6430_b1 , \5418_b1 );
not ( \6430_b1 , w_20436 );
not ( \6430_b0 , w_20437 );
and ( w_20436 , w_20437 , \5418_b0 );
buf ( \6431_b1 , \4616_b1 );
not ( \6431_b1 , w_20438 );
not ( \6431_b0 , w_20439 );
and ( w_20438 , w_20439 , \4616_b0 );
or ( \6432_b1 , \6430_b1 , w_20440 );
or ( \6432_b0 , \6430_b0 , \6431_b0 );
not ( \6431_b0 , w_20441 );
and ( w_20441 , w_20440 , \6431_b1 );
or ( \6433_b1 , \5301_b1 , w_20443 );
not ( w_20443 , w_20444 );
and ( \6433_b0 , \5301_b0 , w_20445 );
and ( w_20444 ,  , w_20445 );
buf ( w_20443 , \4098_b1 );
not ( w_20443 , w_20446 );
not (  , w_20447 );
and ( w_20446 , w_20447 , \4098_b0 );
or ( \6434_b1 , \6432_b1 , w_20449 );
not ( w_20449 , w_20450 );
and ( \6434_b0 , \6432_b0 , w_20451 );
and ( w_20450 ,  , w_20451 );
buf ( w_20449 , \6433_b1 );
not ( w_20449 , w_20452 );
not (  , w_20453 );
and ( w_20452 , w_20453 , \6433_b0 );
buf ( \6435_b1 , \6434_b1 );
not ( \6435_b1 , w_20454 );
not ( \6435_b0 , w_20455 );
and ( w_20454 , w_20455 , \6434_b0 );
buf ( \6436_b1 , \4611_b1 );
not ( \6436_b1 , w_20456 );
not ( \6436_b0 , w_20457 );
and ( w_20456 , w_20457 , \4611_b0 );
or ( \6437_b1 , \6435_b1 , w_20458 );
or ( \6437_b0 , \6435_b0 , \6436_b0 );
not ( \6436_b0 , w_20459 );
and ( w_20459 , w_20458 , \6436_b1 );
or ( \6438_b1 , \6295_b1 , w_20461 );
not ( w_20461 , w_20462 );
and ( \6438_b0 , \6295_b0 , w_20463 );
and ( w_20462 ,  , w_20463 );
buf ( w_20461 , \4754_b1 );
not ( w_20461 , w_20464 );
not (  , w_20465 );
and ( w_20464 , w_20465 , \4754_b0 );
or ( \6439_b1 , \6437_b1 , w_20467 );
not ( w_20467 , w_20468 );
and ( \6439_b0 , \6437_b0 , w_20469 );
and ( w_20468 ,  , w_20469 );
buf ( w_20467 , \6438_b1 );
not ( w_20467 , w_20470 );
not (  , w_20471 );
and ( w_20470 , w_20471 , \6438_b0 );
buf ( \6440_b1 , \6439_b1 );
not ( \6440_b1 , w_20472 );
not ( \6440_b0 , w_20473 );
and ( w_20472 , w_20473 , \6439_b0 );
buf ( \6441_b1 , \4072_b1 );
not ( \6441_b1 , w_20474 );
not ( \6441_b0 , w_20475 );
and ( w_20474 , w_20475 , \4072_b0 );
buf ( \6442_b1 , \5422_b1 );
not ( \6442_b1 , w_20476 );
not ( \6442_b0 , w_20477 );
and ( w_20476 , w_20477 , \5422_b0 );
or ( \6443_b1 , \6441_b1 , w_20478 );
or ( \6443_b0 , \6441_b0 , \6442_b0 );
not ( \6442_b0 , w_20479 );
and ( w_20479 , w_20478 , \6442_b1 );
or ( \6444_b1 , \5275_b1 , w_20481 );
not ( w_20481 , w_20482 );
and ( \6444_b0 , \5275_b0 , w_20483 );
and ( w_20482 ,  , w_20483 );
buf ( w_20481 , \5089_b1 );
not ( w_20481 , w_20484 );
not (  , w_20485 );
and ( w_20484 , w_20485 , \5089_b0 );
or ( \6445_b1 , \6443_b1 , w_20487 );
not ( w_20487 , w_20488 );
and ( \6445_b0 , \6443_b0 , w_20489 );
and ( w_20488 ,  , w_20489 );
buf ( w_20487 , \6444_b1 );
not ( w_20487 , w_20490 );
not (  , w_20491 );
and ( w_20490 , w_20491 , \6444_b0 );
buf ( \6446_b1 , \6445_b1 );
not ( \6446_b1 , w_20492 );
not ( \6446_b0 , w_20493 );
and ( w_20492 , w_20493 , \6445_b0 );
buf ( \6447_b1 , \6337_b1 );
not ( \6447_b1 , w_20494 );
not ( \6447_b0 , w_20495 );
and ( w_20494 , w_20495 , \6337_b0 );
or ( \6448_b1 , \6446_b1 , w_20496 );
or ( \6448_b0 , \6446_b0 , \6447_b0 );
not ( \6447_b0 , w_20497 );
and ( w_20497 , w_20496 , \6447_b1 );
or ( \6449_b1 , \6335_b1 , w_20499 );
not ( w_20499 , w_20500 );
and ( \6449_b0 , \6335_b0 , w_20501 );
and ( w_20500 ,  , w_20501 );
buf ( w_20499 , \5266_b1 );
not ( w_20499 , w_20502 );
not (  , w_20503 );
and ( w_20502 , w_20503 , \5266_b0 );
or ( \6450_b1 , \6448_b1 , w_20505 );
not ( w_20505 , w_20506 );
and ( \6450_b0 , \6448_b0 , w_20507 );
and ( w_20506 ,  , w_20507 );
buf ( w_20505 , \6449_b1 );
not ( w_20505 , w_20508 );
not (  , w_20509 );
and ( w_20508 , w_20509 , \6449_b0 );
buf ( \6451_b1 , \6450_b1 );
not ( \6451_b1 , w_20510 );
not ( \6451_b0 , w_20511 );
and ( w_20510 , w_20511 , \6450_b0 );
or ( \6452_b1 , \6440_b1 , w_20513 );
not ( w_20513 , w_20514 );
and ( \6452_b0 , \6440_b0 , w_20515 );
and ( w_20514 ,  , w_20515 );
buf ( w_20513 , \6451_b1 );
not ( w_20513 , w_20516 );
not (  , w_20517 );
and ( w_20516 , w_20517 , \6451_b0 );
buf ( \6453_b1 , \6452_b1 );
not ( \6453_b1 , w_20518 );
not ( \6453_b0 , w_20519 );
and ( w_20518 , w_20519 , \6452_b0 );
buf ( \6454_b1 , \6327_b1 );
not ( \6454_b1 , w_20520 );
not ( \6454_b0 , w_20521 );
and ( w_20520 , w_20521 , \6327_b0 );
buf ( \6455_b1 , \6321_b1 );
not ( \6455_b1 , w_20522 );
not ( \6455_b0 , w_20523 );
and ( w_20522 , w_20523 , \6321_b0 );
buf ( \6456_b1 , \6455_b1 );
not ( \6456_b1 , w_20524 );
not ( \6456_b0 , w_20525 );
and ( w_20524 , w_20525 , \6455_b0 );
or ( \6457_b1 , \6454_b1 , w_20526 );
or ( \6457_b0 , \6454_b0 , \6456_b0 );
not ( \6456_b0 , w_20527 );
and ( w_20527 , w_20526 , \6456_b1 );
or ( \6458_b1 , \6455_b1 , w_20528 );
or ( \6458_b0 , \6455_b0 , \6327_b0 );
not ( \6327_b0 , w_20529 );
and ( w_20529 , w_20528 , \6327_b1 );
or ( \6459_b1 , \6457_b1 , w_20531 );
not ( w_20531 , w_20532 );
and ( \6459_b0 , \6457_b0 , w_20533 );
and ( w_20532 ,  , w_20533 );
buf ( w_20531 , \6458_b1 );
not ( w_20531 , w_20534 );
not (  , w_20535 );
and ( w_20534 , w_20535 , \6458_b0 );
buf ( \6460_b1 , \6459_b1 );
not ( \6460_b1 , w_20536 );
not ( \6460_b0 , w_20537 );
and ( w_20536 , w_20537 , \6459_b0 );
or ( \6461_b1 , \6453_b1 , w_20538 );
or ( \6461_b0 , \6453_b0 , \6460_b0 );
not ( \6460_b0 , w_20539 );
and ( w_20539 , w_20538 , \6460_b1 );
or ( \6462_b1 , \6439_b1 , w_20541 );
not ( w_20541 , w_20542 );
and ( \6462_b0 , \6439_b0 , w_20543 );
and ( w_20542 ,  , w_20543 );
buf ( w_20541 , \6450_b1 );
not ( w_20541 , w_20544 );
not (  , w_20545 );
and ( w_20544 , w_20545 , \6450_b0 );
or ( \6463_b1 , \6461_b1 , w_20547 );
not ( w_20547 , w_20548 );
and ( \6463_b0 , \6461_b0 , w_20549 );
and ( w_20548 ,  , w_20549 );
buf ( w_20547 , \6462_b1 );
not ( w_20547 , w_20550 );
not (  , w_20551 );
and ( w_20550 , w_20551 , \6462_b0 );
buf ( \6464_b1 , \6463_b1 );
not ( \6464_b1 , w_20552 );
not ( \6464_b0 , w_20553 );
and ( w_20552 , w_20553 , \6463_b0 );
buf ( \6465_b1 , \6328_b1 );
not ( \6465_b1 , w_20554 );
not ( \6465_b0 , w_20555 );
and ( w_20554 , w_20555 , \6328_b0 );
buf ( \6466_b1 , \6306_b1 );
not ( \6466_b1 , w_20556 );
not ( \6466_b0 , w_20557 );
and ( w_20556 , w_20557 , \6306_b0 );
or ( \6467_b1 , \6465_b1 , \6466_b1 );
not ( \6466_b1 , w_20558 );
and ( \6467_b0 , \6465_b0 , w_20559 );
and ( w_20558 , w_20559 , \6466_b0 );
or ( \6468_b1 , \6328_b1 , \6306_b1 );
not ( \6306_b1 , w_20560 );
and ( \6468_b0 , \6328_b0 , w_20561 );
and ( w_20560 , w_20561 , \6306_b0 );
or ( \6469_b1 , \6467_b1 , w_20563 );
not ( w_20563 , w_20564 );
and ( \6469_b0 , \6467_b0 , w_20565 );
and ( w_20564 ,  , w_20565 );
buf ( w_20563 , \6468_b1 );
not ( w_20563 , w_20566 );
not (  , w_20567 );
and ( w_20566 , w_20567 , \6468_b0 );
or ( \6470_b1 , \6359_b1 , \6469_b1 );
xor ( \6470_b0 , \6359_b0 , w_20568 );
not ( w_20568 , w_20569 );
and ( w_20569 , \6469_b1 , \6469_b0 );
or ( \6471_b1 , \6464_b1 , w_20571 );
not ( w_20571 , w_20572 );
and ( \6471_b0 , \6464_b0 , w_20573 );
and ( w_20572 ,  , w_20573 );
buf ( w_20571 , \6470_b1 );
not ( w_20571 , w_20574 );
not (  , w_20575 );
and ( w_20574 , w_20575 , \6470_b0 );
buf ( \6472_b1 , \6471_b1 );
not ( \6472_b1 , w_20576 );
not ( \6472_b0 , w_20577 );
and ( w_20576 , w_20577 , \6471_b0 );
buf ( \6473_b1 , \4602_b1 );
not ( \6473_b1 , w_20578 );
not ( \6473_b0 , w_20579 );
and ( w_20578 , w_20579 , \4602_b0 );
or ( \6474_b1 , \6473_b1 , w_20581 );
not ( w_20581 , w_20582 );
and ( \6474_b0 , \6473_b0 , w_20583 );
and ( w_20582 ,  , w_20583 );
buf ( w_20581 , \4098_b1 );
not ( w_20581 , w_20584 );
not (  , w_20585 );
and ( w_20584 , w_20585 , \4098_b0 );
buf ( \6475_b1 , \4082_b1 );
not ( \6475_b1 , w_20586 );
not ( \6475_b0 , w_20587 );
and ( w_20586 , w_20587 , \4082_b0 );
buf ( \6476_b1 , \4939_b1 );
not ( \6476_b1 , w_20588 );
not ( \6476_b0 , w_20589 );
and ( w_20588 , w_20589 , \4939_b0 );
or ( \6477_b1 , \6475_b1 , w_20590 );
or ( \6477_b0 , \6475_b0 , \6476_b0 );
not ( \6476_b0 , w_20591 );
and ( w_20591 , w_20590 , \6476_b1 );
or ( \6478_b1 , \4936_b1 , w_20593 );
not ( w_20593 , w_20594 );
and ( \6478_b0 , \4936_b0 , w_20595 );
and ( w_20594 ,  , w_20595 );
buf ( w_20593 , \5526_b1 );
not ( w_20593 , w_20596 );
not (  , w_20597 );
and ( w_20596 , w_20597 , \5526_b0 );
or ( \6479_b1 , \6477_b1 , w_20599 );
not ( w_20599 , w_20600 );
and ( \6479_b0 , \6477_b0 , w_20601 );
and ( w_20600 ,  , w_20601 );
buf ( w_20599 , \6478_b1 );
not ( w_20599 , w_20602 );
not (  , w_20603 );
and ( w_20602 , w_20603 , \6478_b0 );
buf ( \6480_b1 , \6479_b1 );
not ( \6480_b1 , w_20604 );
not ( \6480_b0 , w_20605 );
and ( w_20604 , w_20605 , \6479_b0 );
buf ( \6481_b1 , \4945_b1 );
not ( \6481_b1 , w_20606 );
not ( \6481_b0 , w_20607 );
and ( w_20606 , w_20607 , \4945_b0 );
or ( \6482_b1 , \6480_b1 , w_20608 );
or ( \6482_b0 , \6480_b0 , \6481_b0 );
not ( \6481_b0 , w_20609 );
and ( w_20609 , w_20608 , \6481_b1 );
or ( \6483_b1 , \6312_b1 , w_20611 );
not ( w_20611 , w_20612 );
and ( \6483_b0 , \6312_b0 , w_20613 );
and ( w_20612 ,  , w_20613 );
buf ( w_20611 , \4863_b1 );
not ( w_20611 , w_20614 );
not (  , w_20615 );
and ( w_20614 , w_20615 , \4863_b0 );
or ( \6484_b1 , \6482_b1 , w_20617 );
not ( w_20617 , w_20618 );
and ( \6484_b0 , \6482_b0 , w_20619 );
and ( w_20618 ,  , w_20619 );
buf ( w_20617 , \6483_b1 );
not ( w_20617 , w_20620 );
not (  , w_20621 );
and ( w_20620 , w_20621 , \6483_b0 );
or ( \6485_b1 , \6474_b1 , \6484_b1 );
xor ( \6485_b0 , \6474_b0 , w_20622 );
not ( w_20622 , w_20623 );
and ( w_20623 , \6484_b1 , \6484_b0 );
buf ( \6486_b1 , \4076_b1 );
not ( \6486_b1 , w_20624 );
not ( \6486_b0 , w_20625 );
and ( w_20624 , w_20625 , \4076_b0 );
buf ( \6487_b1 , \5422_b1 );
not ( \6487_b1 , w_20626 );
not ( \6487_b0 , w_20627 );
and ( w_20626 , w_20627 , \5422_b0 );
or ( \6488_b1 , \6486_b1 , w_20628 );
or ( \6488_b0 , \6486_b0 , \6487_b0 );
not ( \6487_b0 , w_20629 );
and ( w_20629 , w_20628 , \6487_b1 );
or ( \6489_b1 , \5425_b1 , w_20631 );
not ( w_20631 , w_20632 );
and ( \6489_b0 , \5425_b0 , w_20633 );
and ( w_20632 ,  , w_20633 );
buf ( w_20631 , \5284_b1 );
not ( w_20631 , w_20634 );
not (  , w_20635 );
and ( w_20634 , w_20635 , \5284_b0 );
or ( \6490_b1 , \6488_b1 , w_20637 );
not ( w_20637 , w_20638 );
and ( \6490_b0 , \6488_b0 , w_20639 );
and ( w_20638 ,  , w_20639 );
buf ( w_20637 , \6489_b1 );
not ( w_20637 , w_20640 );
not (  , w_20641 );
and ( w_20640 , w_20641 , \6489_b0 );
buf ( \6491_b1 , \5270_b1 );
not ( \6491_b1 , w_20642 );
not ( \6491_b0 , w_20643 );
and ( w_20642 , w_20643 , \5270_b0 );
buf ( \6492_b1 , \6491_b1 );
not ( \6492_b1 , w_20644 );
not ( \6492_b0 , w_20645 );
and ( w_20644 , w_20645 , \6491_b0 );
or ( \6493_b1 , \6490_b1 , w_20647 );
not ( w_20647 , w_20648 );
and ( \6493_b0 , \6490_b0 , w_20649 );
and ( w_20648 ,  , w_20649 );
buf ( w_20647 , \6492_b1 );
not ( w_20647 , w_20650 );
not (  , w_20651 );
and ( w_20650 , w_20651 , \6492_b0 );
or ( \6494_b1 , \5266_b1 , w_20653 );
not ( w_20653 , w_20654 );
and ( \6494_b0 , \5266_b0 , w_20655 );
and ( w_20654 ,  , w_20655 );
buf ( w_20653 , \6445_b1 );
not ( w_20653 , w_20656 );
not (  , w_20657 );
and ( w_20656 , w_20657 , \6445_b0 );
or ( \6495_b1 , \6493_b1 , \6494_b1 );
not ( \6494_b1 , w_20658 );
and ( \6495_b0 , \6493_b0 , w_20659 );
and ( w_20658 , w_20659 , \6494_b0 );
or ( \6496_b1 , \6485_b1 , w_20660 );
xor ( \6496_b0 , \6485_b0 , w_20662 );
not ( w_20662 , w_20663 );
and ( w_20663 , w_20660 , w_20661 );
buf ( w_20660 , \6495_b1 );
not ( w_20660 , w_20664 );
not ( w_20661 , w_20665 );
and ( w_20664 , w_20665 , \6495_b0 );
or ( \6497_b1 , \4851_b1 , w_20667 );
not ( w_20667 , w_20668 );
and ( \6497_b0 , \4851_b0 , w_20669 );
and ( w_20668 ,  , w_20669 );
buf ( w_20667 , \4098_b1 );
not ( w_20667 , w_20670 );
not (  , w_20671 );
and ( w_20670 , w_20671 , \4098_b0 );
or ( \6498_b1 , \4934_b1 , \6497_b1 );
not ( \6497_b1 , w_20672 );
and ( \6498_b0 , \4934_b0 , w_20673 );
and ( w_20672 , w_20673 , \6497_b0 );
buf ( \6499_b1 , \5418_b1 );
not ( \6499_b1 , w_20674 );
not ( \6499_b0 , w_20675 );
and ( w_20674 , w_20675 , \5418_b0 );
buf ( \6500_b1 , \4856_b1 );
not ( \6500_b1 , w_20676 );
not ( \6500_b0 , w_20677 );
and ( w_20676 , w_20677 , \4856_b0 );
or ( \6501_b1 , \6499_b1 , w_20678 );
or ( \6501_b0 , \6499_b0 , \6500_b0 );
not ( \6500_b0 , w_20679 );
and ( w_20679 , w_20678 , \6500_b1 );
or ( \6502_b1 , \6501_b1 , w_20681 );
not ( w_20681 , w_20682 );
and ( \6502_b0 , \6501_b0 , w_20683 );
and ( w_20682 ,  , w_20683 );
buf ( w_20681 , \5275_b1 );
not ( w_20681 , w_20684 );
not (  , w_20685 );
and ( w_20684 , w_20685 , \5275_b0 );
or ( \6503_b1 , \6498_b1 , w_20687 );
not ( w_20687 , w_20688 );
and ( \6503_b0 , \6498_b0 , w_20689 );
and ( w_20688 ,  , w_20689 );
buf ( w_20687 , \6502_b1 );
not ( w_20687 , w_20690 );
not (  , w_20691 );
and ( w_20690 , w_20691 , \6502_b0 );
buf ( \6504_b1 , \6503_b1 );
not ( \6504_b1 , w_20692 );
not ( \6504_b0 , w_20693 );
and ( w_20692 , w_20693 , \6503_b0 );
or ( \6505_b1 , \5418_b1 , \4935_b1 );
not ( \4935_b1 , w_20694 );
and ( \6505_b0 , \5418_b0 , w_20695 );
and ( w_20694 , w_20695 , \4935_b0 );
buf ( \6506_b1 , \5418_b1 );
not ( \6506_b1 , w_20696 );
not ( \6506_b0 , w_20697 );
and ( w_20696 , w_20697 , \5418_b0 );
or ( \6507_b1 , \6506_b1 , \4949_b1 );
not ( \4949_b1 , w_20698 );
and ( \6507_b0 , \6506_b0 , w_20699 );
and ( w_20698 , w_20699 , \4949_b0 );
or ( \6508_b1 , \6505_b1 , w_20701 );
not ( w_20701 , w_20702 );
and ( \6508_b0 , \6505_b0 , w_20703 );
and ( w_20702 ,  , w_20703 );
buf ( w_20701 , \6507_b1 );
not ( w_20701 , w_20704 );
not (  , w_20705 );
and ( w_20704 , w_20705 , \6507_b0 );
buf ( \6509_b1 , \6508_b1 );
not ( \6509_b1 , w_20706 );
not ( \6509_b0 , w_20707 );
and ( w_20706 , w_20707 , \6508_b0 );
buf ( \6510_b1 , \4945_b1 );
not ( \6510_b1 , w_20708 );
not ( \6510_b0 , w_20709 );
and ( w_20708 , w_20709 , \4945_b0 );
or ( \6511_b1 , \6509_b1 , w_20710 );
or ( \6511_b0 , \6509_b0 , \6510_b0 );
not ( \6510_b0 , w_20711 );
and ( w_20711 , w_20710 , \6510_b1 );
or ( \6512_b1 , \4948_b1 , w_20713 );
not ( w_20713 , w_20714 );
and ( \6512_b0 , \4948_b0 , w_20715 );
and ( w_20714 ,  , w_20715 );
buf ( w_20713 , \6479_b1 );
not ( w_20713 , w_20716 );
not (  , w_20717 );
and ( w_20716 , w_20717 , \6479_b0 );
or ( \6513_b1 , \6511_b1 , w_20719 );
not ( w_20719 , w_20720 );
and ( \6513_b0 , \6511_b0 , w_20721 );
and ( w_20720 ,  , w_20721 );
buf ( w_20719 , \6512_b1 );
not ( w_20719 , w_20722 );
not (  , w_20723 );
and ( w_20722 , w_20723 , \6512_b0 );
or ( \6514_b1 , \6504_b1 , w_20725 );
not ( w_20725 , w_20726 );
and ( \6514_b0 , \6504_b0 , w_20727 );
and ( w_20726 ,  , w_20727 );
buf ( w_20725 , \6513_b1 );
not ( w_20725 , w_20728 );
not (  , w_20729 );
and ( w_20728 , w_20729 , \6513_b0 );
or ( \6515_b1 , \6496_b1 , w_20731 );
not ( w_20731 , w_20732 );
and ( \6515_b0 , \6496_b0 , w_20733 );
and ( w_20732 ,  , w_20733 );
buf ( w_20731 , \6514_b1 );
not ( w_20731 , w_20734 );
not (  , w_20735 );
and ( w_20734 , w_20735 , \6514_b0 );
buf ( \6516_b1 , \6515_b1 );
not ( \6516_b1 , w_20736 );
not ( \6516_b0 , w_20737 );
and ( w_20736 , w_20737 , \6515_b0 );
buf ( \6517_b1 , \5535_b1 );
not ( \6517_b1 , w_20738 );
not ( \6517_b0 , w_20739 );
and ( w_20738 , w_20739 , \5535_b0 );
buf ( \6518_b1 , \5275_b1 );
not ( \6518_b1 , w_20740 );
not ( \6518_b0 , w_20741 );
and ( w_20740 , w_20741 , \5275_b0 );
or ( \6519_b1 , \6517_b1 , w_20742 );
or ( \6519_b0 , \6517_b0 , \6518_b0 );
not ( \6518_b0 , w_20743 );
and ( w_20743 , w_20742 , \6518_b1 );
or ( \6520_b1 , \5422_b1 , w_20745 );
not ( w_20745 , w_20746 );
and ( \6520_b0 , \5422_b0 , w_20747 );
and ( w_20746 ,  , w_20747 );
buf ( w_20745 , \4079_b1 );
not ( w_20745 , w_20748 );
not (  , w_20749 );
and ( w_20748 , w_20749 , \4079_b0 );
or ( \6521_b1 , \6519_b1 , w_20751 );
not ( w_20751 , w_20752 );
and ( \6521_b0 , \6519_b0 , w_20753 );
and ( w_20752 ,  , w_20753 );
buf ( w_20751 , \6520_b1 );
not ( w_20751 , w_20754 );
not (  , w_20755 );
and ( w_20754 , w_20755 , \6520_b0 );
buf ( \6522_b1 , \6521_b1 );
not ( \6522_b1 , w_20756 );
not ( \6522_b0 , w_20757 );
and ( w_20756 , w_20757 , \6521_b0 );
buf ( \6523_b1 , \6337_b1 );
not ( \6523_b1 , w_20758 );
not ( \6523_b0 , w_20759 );
and ( w_20758 , w_20759 , \6337_b0 );
or ( \6524_b1 , \6522_b1 , w_20760 );
or ( \6524_b0 , \6522_b0 , \6523_b0 );
not ( \6523_b0 , w_20761 );
and ( w_20761 , w_20760 , \6523_b1 );
or ( \6525_b1 , \6490_b1 , w_20763 );
not ( w_20763 , w_20764 );
and ( \6525_b0 , \6490_b0 , w_20765 );
and ( w_20764 ,  , w_20765 );
buf ( w_20763 , \5266_b1 );
not ( w_20763 , w_20766 );
not (  , w_20767 );
and ( w_20766 , w_20767 , \5266_b0 );
or ( \6526_b1 , \6524_b1 , w_20769 );
not ( w_20769 , w_20770 );
and ( \6526_b0 , \6524_b0 , w_20771 );
and ( w_20770 ,  , w_20771 );
buf ( w_20769 , \6525_b1 );
not ( w_20769 , w_20772 );
not (  , w_20773 );
and ( w_20772 , w_20773 , \6525_b0 );
buf ( \6527_b1 , \4082_b1 );
not ( \6527_b1 , w_20774 );
not ( \6527_b0 , w_20775 );
and ( w_20774 , w_20775 , \4082_b0 );
buf ( \6528_b1 , \5274_b1 );
not ( \6528_b1 , w_20776 );
not ( \6528_b0 , w_20777 );
and ( w_20776 , w_20777 , \5274_b0 );
or ( \6529_b1 , \6527_b1 , w_20778 );
or ( \6529_b0 , \6527_b0 , \6528_b0 );
not ( \6528_b0 , w_20779 );
and ( w_20779 , w_20778 , \6528_b1 );
or ( \6530_b1 , \5433_b1 , w_20781 );
not ( w_20781 , w_20782 );
and ( \6530_b0 , \5433_b0 , w_20783 );
and ( w_20782 ,  , w_20783 );
buf ( w_20781 , \5526_b1 );
not ( w_20781 , w_20784 );
not (  , w_20785 );
and ( w_20784 , w_20785 , \5526_b0 );
or ( \6531_b1 , \6529_b1 , w_20787 );
not ( w_20787 , w_20788 );
and ( \6531_b0 , \6529_b0 , w_20789 );
and ( w_20788 ,  , w_20789 );
buf ( w_20787 , \6530_b1 );
not ( w_20787 , w_20790 );
not (  , w_20791 );
and ( w_20790 , w_20791 , \6530_b0 );
buf ( \6532_b1 , \6531_b1 );
not ( \6532_b1 , w_20792 );
not ( \6532_b0 , w_20793 );
and ( w_20792 , w_20793 , \6531_b0 );
buf ( \6533_b1 , \6532_b1 );
not ( \6533_b1 , w_20794 );
not ( \6533_b0 , w_20795 );
and ( w_20794 , w_20795 , \6532_b0 );
buf ( \6534_b1 , \6491_b1 );
not ( \6534_b1 , w_20796 );
not ( \6534_b0 , w_20797 );
and ( w_20796 , w_20797 , \6491_b0 );
or ( \6535_b1 , \6533_b1 , \6534_b1 );
not ( \6534_b1 , w_20798 );
and ( \6535_b0 , \6533_b0 , w_20799 );
and ( w_20798 , w_20799 , \6534_b0 );
or ( \6536_b1 , \6521_b1 , \5266_b1 );
not ( \5266_b1 , w_20800 );
and ( \6536_b0 , \6521_b0 , w_20801 );
and ( w_20800 , w_20801 , \5266_b0 );
or ( \6537_b1 , \6535_b1 , w_20803 );
not ( w_20803 , w_20804 );
and ( \6537_b0 , \6535_b0 , w_20805 );
and ( w_20804 ,  , w_20805 );
buf ( w_20803 , \6536_b1 );
not ( w_20803 , w_20806 );
not (  , w_20807 );
and ( w_20806 , w_20807 , \6536_b0 );
or ( \6538_b1 , \4863_b1 , w_20809 );
not ( w_20809 , w_20810 );
and ( \6538_b0 , \4863_b0 , w_20811 );
and ( w_20810 ,  , w_20811 );
buf ( w_20809 , \4098_b1 );
not ( w_20809 , w_20812 );
not (  , w_20813 );
and ( w_20812 , w_20813 , \4098_b0 );
or ( \6539_b1 , \6537_b1 , w_20815 );
not ( w_20815 , w_20816 );
and ( \6539_b0 , \6537_b0 , w_20817 );
and ( w_20816 ,  , w_20817 );
buf ( w_20815 , \6538_b1 );
not ( w_20815 , w_20818 );
not (  , w_20819 );
and ( w_20818 , w_20819 , \6538_b0 );
buf ( \6540_b1 , \5271_b1 );
not ( \6540_b1 , w_20820 );
not ( \6540_b0 , w_20821 );
and ( w_20820 , w_20821 , \5271_b0 );
buf ( \6541_b1 , \5433_b1 );
not ( \6541_b1 , w_20822 );
not ( \6541_b0 , w_20823 );
and ( w_20822 , w_20823 , \5433_b0 );
or ( \6542_b1 , \5418_b1 , \6541_b1 );
not ( \6541_b1 , w_20824 );
and ( \6542_b0 , \5418_b0 , w_20825 );
and ( w_20824 , w_20825 , \6541_b0 );
buf ( \6543_b1 , \5418_b1 );
not ( \6543_b1 , w_20826 );
not ( \6543_b0 , w_20827 );
and ( w_20826 , w_20827 , \5418_b0 );
or ( \6544_b1 , \6543_b1 , \5275_b1 );
not ( \5275_b1 , w_20828 );
and ( \6544_b0 , \6543_b0 , w_20829 );
and ( w_20828 , w_20829 , \5275_b0 );
or ( \6545_b1 , \6542_b1 , w_20831 );
not ( w_20831 , w_20832 );
and ( \6545_b0 , \6542_b0 , w_20833 );
and ( w_20832 ,  , w_20833 );
buf ( w_20831 , \6544_b1 );
not ( w_20831 , w_20834 );
not (  , w_20835 );
and ( w_20834 , w_20835 , \6544_b0 );
buf ( \6546_b1 , \6545_b1 );
not ( \6546_b1 , w_20836 );
not ( \6546_b0 , w_20837 );
and ( w_20836 , w_20837 , \6545_b0 );
or ( \6547_b1 , \6540_b1 , w_20838 );
or ( \6547_b0 , \6540_b0 , \6546_b0 );
not ( \6546_b0 , w_20839 );
and ( w_20839 , w_20838 , \6546_b1 );
or ( \6548_b1 , \6531_b1 , w_20841 );
not ( w_20841 , w_20842 );
and ( \6548_b0 , \6531_b0 , w_20843 );
and ( w_20842 ,  , w_20843 );
buf ( w_20841 , \5266_b1 );
not ( w_20841 , w_20844 );
not (  , w_20845 );
and ( w_20844 , w_20845 , \5266_b0 );
or ( \6549_b1 , \6547_b1 , w_20847 );
not ( w_20847 , w_20848 );
and ( \6549_b0 , \6547_b0 , w_20849 );
and ( w_20848 ,  , w_20849 );
buf ( w_20847 , \6548_b1 );
not ( w_20847 , w_20850 );
not (  , w_20851 );
and ( w_20850 , w_20851 , \6548_b0 );
or ( \6550_b1 , \5266_b1 , w_20853 );
not ( w_20853 , w_20854 );
and ( \6550_b0 , \5266_b0 , w_20855 );
and ( w_20854 ,  , w_20855 );
buf ( w_20853 , \4098_b1 );
not ( w_20853 , w_20856 );
not (  , w_20857 );
and ( w_20856 , w_20857 , \4098_b0 );
or ( \6551_b1 , \6550_b1 , \5425_b1 );
not ( \5425_b1 , w_20858 );
and ( \6551_b0 , \6550_b0 , w_20859 );
and ( w_20858 , w_20859 , \5425_b0 );
or ( \6552_b1 , \6549_b1 , w_20861 );
not ( w_20861 , w_20862 );
and ( \6552_b0 , \6549_b0 , w_20863 );
and ( w_20862 ,  , w_20863 );
buf ( w_20861 , \6551_b1 );
not ( w_20861 , w_20864 );
not (  , w_20865 );
and ( w_20864 , w_20865 , \6551_b0 );
buf ( \6553_b1 , \6552_b1 );
not ( \6553_b1 , w_20866 );
not ( \6553_b0 , w_20867 );
and ( w_20866 , w_20867 , \6552_b0 );
or ( \6554_b1 , \6539_b1 , w_20869 );
not ( w_20869 , w_20870 );
and ( \6554_b0 , \6539_b0 , w_20871 );
and ( w_20870 ,  , w_20871 );
buf ( w_20869 , \6553_b1 );
not ( w_20869 , w_20872 );
not (  , w_20873 );
and ( w_20872 , w_20873 , \6553_b0 );
buf ( \6555_b1 , \6537_b1 );
not ( \6555_b1 , w_20874 );
not ( \6555_b0 , w_20875 );
and ( w_20874 , w_20875 , \6537_b0 );
buf ( \6556_b1 , \6538_b1 );
not ( \6556_b1 , w_20876 );
not ( \6556_b0 , w_20877 );
and ( w_20876 , w_20877 , \6538_b0 );
or ( \6557_b1 , \6555_b1 , w_20879 );
not ( w_20879 , w_20880 );
and ( \6557_b0 , \6555_b0 , w_20881 );
and ( w_20880 ,  , w_20881 );
buf ( w_20879 , \6556_b1 );
not ( w_20879 , w_20882 );
not (  , w_20883 );
and ( w_20882 , w_20883 , \6556_b0 );
or ( \6558_b1 , \6554_b1 , w_20885 );
not ( w_20885 , w_20886 );
and ( \6558_b0 , \6554_b0 , w_20887 );
and ( w_20886 ,  , w_20887 );
buf ( w_20885 , \6557_b1 );
not ( w_20885 , w_20888 );
not (  , w_20889 );
and ( w_20888 , w_20889 , \6557_b0 );
or ( \6559_b1 , \6526_b1 , \6558_b1 );
xor ( \6559_b0 , \6526_b0 , w_20890 );
not ( w_20890 , w_20891 );
and ( w_20891 , \6558_b1 , \6558_b0 );
buf ( \6560_b1 , \6503_b1 );
not ( \6560_b1 , w_20892 );
not ( \6560_b0 , w_20893 );
and ( w_20892 , w_20893 , \6503_b0 );
buf ( \6561_b1 , \6513_b1 );
not ( \6561_b1 , w_20894 );
not ( \6561_b0 , w_20895 );
and ( w_20894 , w_20895 , \6513_b0 );
or ( \6562_b1 , \6560_b1 , w_20896 );
or ( \6562_b0 , \6560_b0 , \6561_b0 );
not ( \6561_b0 , w_20897 );
and ( w_20897 , w_20896 , \6561_b1 );
or ( \6563_b1 , \6513_b1 , w_20898 );
or ( \6563_b0 , \6513_b0 , \6503_b0 );
not ( \6503_b0 , w_20899 );
and ( w_20899 , w_20898 , \6503_b1 );
or ( \6564_b1 , \6562_b1 , w_20901 );
not ( w_20901 , w_20902 );
and ( \6564_b0 , \6562_b0 , w_20903 );
and ( w_20902 ,  , w_20903 );
buf ( w_20901 , \6563_b1 );
not ( w_20901 , w_20904 );
not (  , w_20905 );
and ( w_20904 , w_20905 , \6563_b0 );
or ( \6565_b1 , \6559_b1 , \6564_b1 );
not ( \6564_b1 , w_20906 );
and ( \6565_b0 , \6559_b0 , w_20907 );
and ( w_20906 , w_20907 , \6564_b0 );
or ( \6566_b1 , \6526_b1 , \6558_b1 );
not ( \6558_b1 , w_20908 );
and ( \6566_b0 , \6526_b0 , w_20909 );
and ( w_20908 , w_20909 , \6558_b0 );
or ( \6567_b1 , \6565_b1 , w_20910 );
or ( \6567_b0 , \6565_b0 , \6566_b0 );
not ( \6566_b0 , w_20911 );
and ( w_20911 , w_20910 , \6566_b1 );
buf ( \6568_b1 , \6567_b1 );
not ( \6568_b1 , w_20912 );
not ( \6568_b0 , w_20913 );
and ( w_20912 , w_20913 , \6567_b0 );
or ( \6569_b1 , \6516_b1 , w_20914 );
or ( \6569_b0 , \6516_b0 , \6568_b0 );
not ( \6568_b0 , w_20915 );
and ( w_20915 , w_20914 , \6568_b1 );
or ( \6570_b1 , \6496_b1 , w_20916 );
or ( \6570_b0 , \6496_b0 , \6514_b0 );
not ( \6514_b0 , w_20917 );
and ( w_20917 , w_20916 , \6514_b1 );
or ( \6571_b1 , \6569_b1 , w_20919 );
not ( w_20919 , w_20920 );
and ( \6571_b0 , \6569_b0 , w_20921 );
and ( w_20920 ,  , w_20921 );
buf ( w_20919 , \6570_b1 );
not ( w_20919 , w_20922 );
not (  , w_20923 );
and ( w_20922 , w_20923 , \6570_b0 );
buf ( \6572_b1 , \6474_b1 );
not ( \6572_b1 , w_20924 );
not ( \6572_b0 , w_20925 );
and ( w_20924 , w_20925 , \6474_b0 );
buf ( \6573_b1 , \6495_b1 );
not ( \6573_b1 , w_20926 );
not ( \6573_b0 , w_20927 );
and ( w_20926 , w_20927 , \6495_b0 );
or ( \6574_b1 , \6572_b1 , w_20928 );
or ( \6574_b0 , \6572_b0 , \6573_b0 );
not ( \6573_b0 , w_20929 );
and ( w_20929 , w_20928 , \6573_b1 );
or ( \6575_b1 , \6574_b1 , w_20931 );
not ( w_20931 , w_20932 );
and ( \6575_b0 , \6574_b0 , w_20933 );
and ( w_20932 ,  , w_20933 );
buf ( w_20931 , \6484_b1 );
not ( w_20931 , w_20934 );
not (  , w_20935 );
and ( w_20934 , w_20935 , \6484_b0 );
or ( \6576_b1 , \6495_b1 , w_20936 );
or ( \6576_b0 , \6495_b0 , \6474_b0 );
not ( \6474_b0 , w_20937 );
and ( w_20937 , w_20936 , \6474_b1 );
or ( \6577_b1 , \6575_b1 , w_20939 );
not ( w_20939 , w_20940 );
and ( \6577_b0 , \6575_b0 , w_20941 );
and ( w_20940 ,  , w_20941 );
buf ( w_20939 , \6576_b1 );
not ( w_20939 , w_20942 );
not (  , w_20943 );
and ( w_20942 , w_20943 , \6576_b0 );
buf ( \6578_b1 , \6577_b1 );
not ( \6578_b1 , w_20944 );
not ( \6578_b0 , w_20945 );
and ( w_20944 , w_20945 , \6577_b0 );
buf ( \6579_b1 , \6459_b1 );
not ( \6579_b1 , w_20946 );
not ( \6579_b0 , w_20947 );
and ( w_20946 , w_20947 , \6459_b0 );
buf ( \6580_b1 , \6439_b1 );
not ( \6580_b1 , w_20948 );
not ( \6580_b0 , w_20949 );
and ( w_20948 , w_20949 , \6439_b0 );
buf ( \6581_b1 , \6451_b1 );
not ( \6581_b1 , w_20950 );
not ( \6581_b0 , w_20951 );
and ( w_20950 , w_20951 , \6451_b0 );
or ( \6582_b1 , \6580_b1 , \6581_b1 );
not ( \6581_b1 , w_20952 );
and ( \6582_b0 , \6580_b0 , w_20953 );
and ( w_20952 , w_20953 , \6581_b0 );
or ( \6583_b1 , \6439_b1 , \6451_b1 );
not ( \6451_b1 , w_20954 );
and ( \6583_b0 , \6439_b0 , w_20955 );
and ( w_20954 , w_20955 , \6451_b0 );
or ( \6584_b1 , \6582_b1 , w_20957 );
not ( w_20957 , w_20958 );
and ( \6584_b0 , \6582_b0 , w_20959 );
and ( w_20958 ,  , w_20959 );
buf ( w_20957 , \6583_b1 );
not ( w_20957 , w_20960 );
not (  , w_20961 );
and ( w_20960 , w_20961 , \6583_b0 );
buf ( \6585_b1 , \6584_b1 );
not ( \6585_b1 , w_20962 );
not ( \6585_b0 , w_20963 );
and ( w_20962 , w_20963 , \6584_b0 );
or ( \6586_b1 , \6579_b1 , \6585_b1 );
not ( \6585_b1 , w_20964 );
and ( \6586_b0 , \6579_b0 , w_20965 );
and ( w_20964 , w_20965 , \6585_b0 );
or ( \6587_b1 , \6459_b1 , \6584_b1 );
not ( \6584_b1 , w_20966 );
and ( \6587_b0 , \6459_b0 , w_20967 );
and ( w_20966 , w_20967 , \6584_b0 );
or ( \6588_b1 , \6586_b1 , w_20969 );
not ( w_20969 , w_20970 );
and ( \6588_b0 , \6586_b0 , w_20971 );
and ( w_20970 ,  , w_20971 );
buf ( w_20969 , \6587_b1 );
not ( w_20969 , w_20972 );
not (  , w_20973 );
and ( w_20972 , w_20973 , \6587_b0 );
or ( \6589_b1 , \6578_b1 , w_20975 );
not ( w_20975 , w_20976 );
and ( \6589_b0 , \6578_b0 , w_20977 );
and ( w_20976 ,  , w_20977 );
buf ( w_20975 , \6588_b1 );
not ( w_20975 , w_20978 );
not (  , w_20979 );
and ( w_20978 , w_20979 , \6588_b0 );
or ( \6590_b1 , \6571_b1 , w_20981 );
not ( w_20981 , w_20982 );
and ( \6590_b0 , \6571_b0 , w_20983 );
and ( w_20982 ,  , w_20983 );
buf ( w_20981 , \6589_b1 );
not ( w_20981 , w_20984 );
not (  , w_20985 );
and ( w_20984 , w_20985 , \6589_b0 );
buf ( \6591_b1 , \6588_b1 );
not ( \6591_b1 , w_20986 );
not ( \6591_b0 , w_20987 );
and ( w_20986 , w_20987 , \6588_b0 );
or ( \6592_b1 , \6591_b1 , w_20989 );
not ( w_20989 , w_20990 );
and ( \6592_b0 , \6591_b0 , w_20991 );
and ( w_20990 ,  , w_20991 );
buf ( w_20989 , \6577_b1 );
not ( w_20989 , w_20992 );
not (  , w_20993 );
and ( w_20992 , w_20993 , \6577_b0 );
or ( \6593_b1 , \6590_b1 , w_20995 );
not ( w_20995 , w_20996 );
and ( \6593_b0 , \6590_b0 , w_20997 );
and ( w_20996 ,  , w_20997 );
buf ( w_20995 , \6592_b1 );
not ( w_20995 , w_20998 );
not (  , w_20999 );
and ( w_20998 , w_20999 , \6592_b0 );
buf ( \6594_b1 , \6593_b1 );
not ( \6594_b1 , w_21000 );
not ( \6594_b0 , w_21001 );
and ( w_21000 , w_21001 , \6593_b0 );
or ( \6595_b1 , \6472_b1 , w_21002 );
or ( \6595_b0 , \6472_b0 , \6594_b0 );
not ( \6594_b0 , w_21003 );
and ( w_21003 , w_21002 , \6594_b1 );
buf ( \6596_b1 , \6470_b1 );
not ( \6596_b1 , w_21004 );
not ( \6596_b0 , w_21005 );
and ( w_21004 , w_21005 , \6470_b0 );
or ( \6597_b1 , \6596_b1 , w_21007 );
not ( w_21007 , w_21008 );
and ( \6597_b0 , \6596_b0 , w_21009 );
and ( w_21008 ,  , w_21009 );
buf ( w_21007 , \6463_b1 );
not ( w_21007 , w_21010 );
not (  , w_21011 );
and ( w_21010 , w_21011 , \6463_b0 );
or ( \6598_b1 , \6595_b1 , w_21013 );
not ( w_21013 , w_21014 );
and ( \6598_b0 , \6595_b0 , w_21015 );
and ( w_21014 ,  , w_21015 );
buf ( w_21013 , \6597_b1 );
not ( w_21013 , w_21016 );
not (  , w_21017 );
and ( w_21016 , w_21017 , \6597_b0 );
or ( \6599_b1 , \6429_b1 , \6598_b1 );
not ( \6598_b1 , w_21018 );
and ( \6599_b0 , \6429_b0 , w_21019 );
and ( w_21018 , w_21019 , \6598_b0 );
or ( \6600_b1 , \6364_b1 , \6428_b1 );
not ( \6428_b1 , w_21020 );
and ( \6600_b0 , \6364_b0 , w_21021 );
and ( w_21020 , w_21021 , \6428_b0 );
or ( \6601_b1 , \6599_b1 , w_21022 );
or ( \6601_b0 , \6599_b0 , \6600_b0 );
not ( \6600_b0 , w_21023 );
and ( w_21023 , w_21022 , \6600_b1 );
buf ( \6602_b1 , \6601_b1 );
not ( \6602_b1 , w_21024 );
not ( \6602_b0 , w_21025 );
and ( w_21024 , w_21025 , \6601_b0 );
buf ( \6603_b1 , \5089_b1 );
not ( \6603_b1 , w_21026 );
not ( \6603_b0 , w_21027 );
and ( w_21026 , w_21027 , \5089_b0 );
buf ( \6604_b1 , \4729_b1 );
not ( \6604_b1 , w_21028 );
not ( \6604_b0 , w_21029 );
and ( w_21028 , w_21029 , \4729_b0 );
or ( \6605_b1 , \6603_b1 , w_21030 );
or ( \6605_b0 , \6603_b0 , \6604_b0 );
not ( \6604_b0 , w_21031 );
and ( w_21031 , w_21030 , \6604_b1 );
or ( \6606_b1 , \4457_b1 , w_21033 );
not ( w_21033 , w_21034 );
and ( \6606_b0 , \4457_b0 , w_21035 );
and ( w_21034 ,  , w_21035 );
buf ( w_21033 , \4072_b1 );
not ( w_21033 , w_21036 );
not (  , w_21037 );
and ( w_21036 , w_21037 , \4072_b0 );
or ( \6607_b1 , \6605_b1 , w_21039 );
not ( w_21039 , w_21040 );
and ( \6607_b0 , \6605_b0 , w_21041 );
and ( w_21040 ,  , w_21041 );
buf ( w_21039 , \6606_b1 );
not ( w_21039 , w_21042 );
not (  , w_21043 );
and ( w_21042 , w_21043 , \6606_b0 );
buf ( \6608_b1 , \6607_b1 );
not ( \6608_b1 , w_21044 );
not ( \6608_b0 , w_21045 );
and ( w_21044 , w_21045 , \6607_b0 );
buf ( \6609_b1 , \4449_b1 );
not ( \6609_b1 , w_21046 );
not ( \6609_b0 , w_21047 );
and ( w_21046 , w_21047 , \4449_b0 );
or ( \6610_b1 , \6608_b1 , w_21048 );
or ( \6610_b0 , \6608_b0 , \6609_b0 );
not ( \6609_b0 , w_21049 );
and ( w_21049 , w_21048 , \6609_b1 );
or ( \6611_b1 , \6200_b1 , w_21051 );
not ( w_21051 , w_21052 );
and ( \6611_b0 , \6200_b0 , w_21053 );
and ( w_21052 ,  , w_21053 );
buf ( w_21051 , \4452_b1 );
not ( w_21051 , w_21054 );
not (  , w_21055 );
and ( w_21054 , w_21055 , \4452_b0 );
or ( \6612_b1 , \6610_b1 , w_21057 );
not ( w_21057 , w_21058 );
and ( \6612_b0 , \6610_b0 , w_21059 );
and ( w_21058 ,  , w_21059 );
buf ( w_21057 , \6611_b1 );
not ( w_21057 , w_21060 );
not (  , w_21061 );
and ( w_21060 , w_21061 , \6611_b0 );
buf ( \6613_b1 , \4093_b1 );
not ( \6613_b1 , w_21062 );
not ( \6613_b0 , w_21063 );
and ( w_21062 , w_21063 , \4093_b0 );
buf ( \6614_b1 , \5422_b1 );
not ( \6614_b1 , w_21064 );
not ( \6614_b0 , w_21065 );
and ( w_21064 , w_21065 , \5422_b0 );
or ( \6615_b1 , \6613_b1 , w_21066 );
or ( \6615_b0 , \6613_b0 , \6614_b0 );
not ( \6614_b0 , w_21067 );
and ( w_21067 , w_21066 , \6614_b1 );
or ( \6616_b1 , \5433_b1 , w_21069 );
not ( w_21069 , w_21070 );
and ( \6616_b0 , \5433_b0 , w_21071 );
and ( w_21070 ,  , w_21071 );
buf ( w_21069 , \4349_b1 );
not ( w_21069 , w_21072 );
not (  , w_21073 );
and ( w_21072 , w_21073 , \4349_b0 );
or ( \6617_b1 , \6615_b1 , w_21075 );
not ( w_21075 , w_21076 );
and ( \6617_b0 , \6615_b0 , w_21077 );
and ( w_21076 ,  , w_21077 );
buf ( w_21075 , \6616_b1 );
not ( w_21075 , w_21078 );
not (  , w_21079 );
and ( w_21078 , w_21079 , \6616_b0 );
buf ( \6618_b1 , \6617_b1 );
not ( \6618_b1 , w_21080 );
not ( \6618_b0 , w_21081 );
and ( w_21080 , w_21081 , \6617_b0 );
buf ( \6619_b1 , \6492_b1 );
not ( \6619_b1 , w_21082 );
not ( \6619_b0 , w_21083 );
and ( w_21082 , w_21083 , \6492_b0 );
or ( \6620_b1 , \6618_b1 , w_21084 );
or ( \6620_b0 , \6618_b0 , \6619_b0 );
not ( \6619_b0 , w_21085 );
and ( w_21085 , w_21084 , \6619_b1 );
or ( \6621_b1 , \6168_b1 , w_21087 );
not ( w_21087 , w_21088 );
and ( \6621_b0 , \6168_b0 , w_21089 );
and ( w_21088 ,  , w_21089 );
buf ( w_21087 , \5266_b1 );
not ( w_21087 , w_21090 );
not (  , w_21091 );
and ( w_21090 , w_21091 , \5266_b0 );
or ( \6622_b1 , \6620_b1 , w_21093 );
not ( w_21093 , w_21094 );
and ( \6622_b0 , \6620_b0 , w_21095 );
and ( w_21094 ,  , w_21095 );
buf ( w_21093 , \6621_b1 );
not ( w_21093 , w_21096 );
not (  , w_21097 );
and ( w_21096 , w_21097 , \6621_b0 );
or ( \6623_b1 , \6612_b1 , \6622_b1 );
xor ( \6623_b0 , \6612_b0 , w_21098 );
not ( w_21098 , w_21099 );
and ( w_21099 , \6622_b1 , \6622_b0 );
buf ( \6624_b1 , \4079_b1 );
not ( \6624_b1 , w_21100 );
not ( \6624_b0 , w_21101 );
and ( w_21100 , w_21101 , \4079_b0 );
buf ( \6625_b1 , \4493_b1 );
not ( \6625_b1 , w_21102 );
not ( \6625_b0 , w_21103 );
and ( w_21102 , w_21103 , \4493_b0 );
or ( \6626_b1 , \6624_b1 , w_21104 );
or ( \6626_b0 , \6624_b0 , \6625_b0 );
not ( \6625_b0 , w_21105 );
and ( w_21105 , w_21104 , \6625_b1 );
or ( \6627_b1 , \4283_b1 , w_21107 );
not ( w_21107 , w_21108 );
and ( \6627_b0 , \4283_b0 , w_21109 );
and ( w_21108 ,  , w_21109 );
buf ( w_21107 , \5535_b1 );
not ( w_21107 , w_21110 );
not (  , w_21111 );
and ( w_21110 , w_21111 , \5535_b0 );
or ( \6628_b1 , \6626_b1 , w_21113 );
not ( w_21113 , w_21114 );
and ( \6628_b0 , \6626_b0 , w_21115 );
and ( w_21114 ,  , w_21115 );
buf ( w_21113 , \6627_b1 );
not ( w_21113 , w_21116 );
not (  , w_21117 );
and ( w_21116 , w_21117 , \6627_b0 );
buf ( \6629_b1 , \6628_b1 );
not ( \6629_b1 , w_21118 );
not ( \6629_b0 , w_21119 );
and ( w_21118 , w_21119 , \6628_b0 );
buf ( \6630_b1 , \4338_b1 );
not ( \6630_b1 , w_21120 );
not ( \6630_b0 , w_21121 );
and ( w_21120 , w_21121 , \4338_b0 );
or ( \6631_b1 , \6629_b1 , w_21122 );
or ( \6631_b0 , \6629_b0 , \6630_b0 );
not ( \6630_b0 , w_21123 );
and ( w_21123 , w_21122 , \6630_b1 );
or ( \6632_b1 , \5160_b1 , w_21125 );
not ( w_21125 , w_21126 );
and ( \6632_b0 , \5160_b0 , w_21127 );
and ( w_21126 ,  , w_21127 );
buf ( w_21125 , \6224_b1 );
not ( w_21125 , w_21128 );
not (  , w_21129 );
and ( w_21128 , w_21129 , \6224_b0 );
or ( \6633_b1 , \6631_b1 , w_21131 );
not ( w_21131 , w_21132 );
and ( \6633_b0 , \6631_b0 , w_21133 );
and ( w_21132 ,  , w_21133 );
buf ( w_21131 , \6632_b1 );
not ( w_21131 , w_21134 );
not (  , w_21135 );
and ( w_21134 , w_21135 , \6632_b0 );
or ( \6634_b1 , \6623_b1 , \6633_b1 );
xor ( \6634_b0 , \6623_b0 , w_21136 );
not ( w_21136 , w_21137 );
and ( w_21137 , \6633_b1 , \6633_b0 );
buf ( \6635_b1 , \6634_b1 );
not ( \6635_b1 , w_21138 );
not ( \6635_b0 , w_21139 );
and ( w_21138 , w_21139 , \6634_b0 );
buf ( \6636_b1 , \4862_b1 );
not ( \6636_b1 , w_21140 );
not ( \6636_b0 , w_21141 );
and ( w_21140 , w_21141 , \4862_b0 );
or ( \6637_b1 , \4866_b1 , \4017_b1 );
not ( \4017_b1 , w_21142 );
and ( \6637_b0 , \4866_b0 , w_21143 );
and ( w_21142 , w_21143 , \4017_b0 );
or ( \6638_b1 , \4934_b1 , \4662_b1 );
not ( \4662_b1 , w_21144 );
and ( \6638_b0 , \4934_b0 , w_21145 );
and ( w_21144 , w_21145 , \4662_b0 );
or ( \6639_b1 , \6637_b1 , w_21147 );
not ( w_21147 , w_21148 );
and ( \6639_b0 , \6637_b0 , w_21149 );
and ( w_21148 ,  , w_21149 );
buf ( w_21147 , \6638_b1 );
not ( w_21147 , w_21150 );
not (  , w_21151 );
and ( w_21150 , w_21151 , \6638_b0 );
buf ( \6640_b1 , \6639_b1 );
not ( \6640_b1 , w_21152 );
not ( \6640_b0 , w_21153 );
and ( w_21152 , w_21153 , \6639_b0 );
or ( \6641_b1 , \6636_b1 , \6640_b1 );
not ( \6640_b1 , w_21154 );
and ( \6641_b0 , \6636_b0 , w_21155 );
and ( w_21154 , w_21155 , \6640_b0 );
buf ( \6642_b1 , \4021_b1 );
not ( \6642_b1 , w_21156 );
not ( \6642_b0 , w_21157 );
and ( w_21156 , w_21157 , \4021_b0 );
buf ( \6643_b1 , \4939_b1 );
not ( \6643_b1 , w_21158 );
not ( \6643_b0 , w_21159 );
and ( w_21158 , w_21159 , \4939_b0 );
or ( \6644_b1 , \6642_b1 , w_21160 );
or ( \6644_b0 , \6642_b0 , \6643_b0 );
not ( \6643_b0 , w_21161 );
and ( w_21161 , w_21160 , \6643_b1 );
or ( \6645_b1 , \4867_b1 , w_21163 );
not ( w_21163 , w_21164 );
and ( \6645_b0 , \4867_b0 , w_21165 );
and ( w_21164 ,  , w_21165 );
buf ( w_21163 , \4780_b1 );
not ( w_21163 , w_21166 );
not (  , w_21167 );
and ( w_21166 , w_21167 , \4780_b0 );
or ( \6646_b1 , \6644_b1 , w_21169 );
not ( w_21169 , w_21170 );
and ( \6646_b0 , \6644_b0 , w_21171 );
and ( w_21170 ,  , w_21171 );
buf ( w_21169 , \6645_b1 );
not ( w_21169 , w_21172 );
not (  , w_21173 );
and ( w_21172 , w_21173 , \6645_b0 );
or ( \6647_b1 , \6646_b1 , w_21175 );
not ( w_21175 , w_21176 );
and ( \6647_b0 , \6646_b0 , w_21177 );
and ( w_21176 ,  , w_21177 );
buf ( w_21175 , \4859_b1 );
not ( w_21175 , w_21178 );
not (  , w_21179 );
and ( w_21178 , w_21179 , \4859_b0 );
buf ( \6648_b1 , \6647_b1 );
not ( \6648_b1 , w_21180 );
not ( \6648_b0 , w_21181 );
and ( w_21180 , w_21181 , \6647_b0 );
or ( \6649_b1 , \6648_b1 , \4862_b1 );
not ( \4862_b1 , w_21182 );
and ( \6649_b0 , \6648_b0 , w_21183 );
and ( w_21182 , w_21183 , \4862_b0 );
or ( \6650_b1 , \6641_b1 , w_21185 );
not ( w_21185 , w_21186 );
and ( \6650_b0 , \6641_b0 , w_21187 );
and ( w_21186 ,  , w_21187 );
buf ( w_21185 , \6649_b1 );
not ( w_21185 , w_21188 );
not (  , w_21189 );
and ( w_21188 , w_21189 , \6649_b0 );
buf ( \6651_b1 , \5418_b1 );
not ( \6651_b1 , w_21190 );
not ( \6651_b0 , w_21191 );
and ( w_21190 , w_21191 , \5418_b0 );
buf ( \6652_b1 , \4270_b1 );
not ( \6652_b1 , w_21192 );
not ( \6652_b0 , w_21193 );
and ( w_21192 , w_21193 , \4270_b0 );
or ( \6653_b1 , \6651_b1 , w_21194 );
or ( \6653_b0 , \6651_b0 , \6652_b0 );
not ( \6652_b0 , w_21195 );
and ( w_21195 , w_21194 , \6652_b1 );
or ( \6654_b1 , \6653_b1 , w_21197 );
not ( w_21197 , w_21198 );
and ( \6654_b0 , \6653_b0 , w_21199 );
and ( w_21198 ,  , w_21199 );
buf ( w_21197 , \4917_b1 );
not ( w_21197 , w_21200 );
not (  , w_21201 );
and ( w_21200 , w_21201 , \4917_b0 );
or ( \6655_b1 , \4274_b1 , w_21203 );
not ( w_21203 , w_21204 );
and ( \6655_b0 , \4274_b0 , w_21205 );
and ( w_21204 ,  , w_21205 );
buf ( w_21203 , \4098_b1 );
not ( w_21203 , w_21206 );
not (  , w_21207 );
and ( w_21206 , w_21207 , \4098_b0 );
or ( \6657_b1 , \6650_b1 , w_21208 );
or ( \6657_b0 , \6650_b0 , \6656_b0 );
not ( \6656_b0 , w_21209 );
and ( w_21209 , w_21208 , \6656_b1 );
buf ( \6658_b1 , \6657_b1 );
not ( \6658_b1 , w_21210 );
not ( \6658_b0 , w_21211 );
and ( w_21210 , w_21211 , \6657_b0 );
or ( \6659_b1 , \4150_b1 , w_21213 );
not ( w_21213 , w_21214 );
and ( \6659_b0 , \4150_b0 , w_21215 );
and ( w_21214 ,  , w_21215 );
buf ( w_21213 , \4098_b1 );
not ( w_21213 , w_21216 );
not (  , w_21217 );
and ( w_21216 , w_21217 , \4098_b0 );
buf ( \6660_b1 , \6659_b1 );
not ( \6660_b1 , w_21218 );
not ( \6660_b0 , w_21219 );
and ( w_21218 , w_21219 , \6659_b0 );
buf ( \6661_b1 , \4095_b1 );
not ( \6661_b1 , w_21220 );
not ( \6661_b0 , w_21221 );
and ( w_21220 , w_21221 , \4095_b0 );
buf ( \6662_b1 , \5274_b1 );
not ( \6662_b1 , w_21222 );
not ( \6662_b0 , w_21223 );
and ( w_21222 , w_21223 , \5274_b0 );
or ( \6663_b1 , \6661_b1 , w_21224 );
or ( \6663_b0 , \6661_b0 , \6662_b0 );
not ( \6662_b0 , w_21225 );
and ( w_21225 , w_21224 , \6662_b1 );
or ( \6664_b1 , \5433_b1 , w_21227 );
not ( w_21227 , w_21228 );
and ( \6664_b0 , \5433_b0 , w_21229 );
and ( w_21228 ,  , w_21229 );
buf ( w_21227 , \4391_b1 );
not ( w_21227 , w_21230 );
not (  , w_21231 );
and ( w_21230 , w_21231 , \4391_b0 );
or ( \6665_b1 , \6663_b1 , w_21233 );
not ( w_21233 , w_21234 );
and ( \6665_b0 , \6663_b0 , w_21235 );
and ( w_21234 ,  , w_21235 );
buf ( w_21233 , \6664_b1 );
not ( w_21233 , w_21236 );
not (  , w_21237 );
and ( w_21236 , w_21237 , \6664_b0 );
buf ( \6666_b1 , \6665_b1 );
not ( \6666_b1 , w_21238 );
not ( \6666_b0 , w_21239 );
and ( w_21238 , w_21239 , \6665_b0 );
buf ( \6667_b1 , \5270_b1 );
not ( \6667_b1 , w_21240 );
not ( \6667_b0 , w_21241 );
and ( w_21240 , w_21241 , \5270_b0 );
or ( \6668_b1 , \6666_b1 , w_21242 );
or ( \6668_b0 , \6666_b0 , \6667_b0 );
not ( \6667_b0 , w_21243 );
and ( w_21243 , w_21242 , \6667_b1 );
or ( \6669_b1 , \6617_b1 , w_21245 );
not ( w_21245 , w_21246 );
and ( \6669_b0 , \6617_b0 , w_21247 );
and ( w_21246 ,  , w_21247 );
buf ( w_21245 , \5266_b1 );
not ( w_21245 , w_21248 );
not (  , w_21249 );
and ( w_21248 , w_21249 , \5266_b0 );
or ( \6670_b1 , \6668_b1 , w_21251 );
not ( w_21251 , w_21252 );
and ( \6670_b0 , \6668_b0 , w_21253 );
and ( w_21252 ,  , w_21253 );
buf ( w_21251 , \6669_b1 );
not ( w_21251 , w_21254 );
not (  , w_21255 );
and ( w_21254 , w_21255 , \6669_b0 );
or ( \6671_b1 , \6660_b1 , \6670_b1 );
not ( \6670_b1 , w_21256 );
and ( \6671_b0 , \6660_b0 , w_21257 );
and ( w_21256 , w_21257 , \6670_b0 );
buf ( \6672_b1 , \6660_b1 );
not ( \6672_b1 , w_21258 );
not ( \6672_b0 , w_21259 );
and ( w_21258 , w_21259 , \6660_b0 );
buf ( \6673_b1 , \6670_b1 );
not ( \6673_b1 , w_21260 );
not ( \6673_b0 , w_21261 );
and ( w_21260 , w_21261 , \6670_b0 );
or ( \6674_b1 , \6672_b1 , \6673_b1 );
not ( \6673_b1 , w_21262 );
and ( \6674_b0 , \6672_b0 , w_21263 );
and ( w_21262 , w_21263 , \6673_b0 );
or ( \6675_b1 , \6671_b1 , w_21265 );
not ( w_21265 , w_21266 );
and ( \6675_b0 , \6671_b0 , w_21267 );
and ( w_21266 ,  , w_21267 );
buf ( w_21265 , \6674_b1 );
not ( w_21265 , w_21268 );
not (  , w_21269 );
and ( w_21268 , w_21269 , \6674_b0 );
buf ( \6676_b1 , \6639_b1 );
not ( \6676_b1 , w_21270 );
not ( \6676_b0 , w_21271 );
and ( w_21270 , w_21271 , \6639_b0 );
buf ( \6677_b1 , \6676_b1 );
not ( \6677_b1 , w_21272 );
not ( \6677_b0 , w_21273 );
and ( w_21272 , w_21273 , \6676_b0 );
buf ( \6678_b1 , \4945_b1 );
not ( \6678_b1 , w_21274 );
not ( \6678_b0 , w_21275 );
and ( w_21274 , w_21275 , \4945_b0 );
or ( \6679_b1 , \6677_b1 , w_21276 );
or ( \6679_b0 , \6677_b0 , \6678_b0 );
not ( \6678_b0 , w_21277 );
and ( w_21277 , w_21276 , \6678_b1 );
buf ( \6680_b1 , \4066_b1 );
not ( \6680_b1 , w_21278 );
not ( \6680_b0 , w_21279 );
and ( w_21278 , w_21279 , \4066_b0 );
buf ( \6681_b1 , \5903_b1 );
not ( \6681_b1 , w_21280 );
not ( \6681_b0 , w_21281 );
and ( w_21280 , w_21281 , \5903_b0 );
or ( \6682_b1 , \6680_b1 , w_21282 );
or ( \6682_b0 , \6680_b0 , \6681_b0 );
not ( \6681_b0 , w_21283 );
and ( w_21283 , w_21282 , \6681_b1 );
or ( \6683_b1 , \5905_b1 , w_21285 );
not ( w_21285 , w_21286 );
and ( \6683_b0 , \5905_b0 , w_21287 );
and ( w_21286 ,  , w_21287 );
buf ( w_21285 , \4519_b1 );
not ( w_21285 , w_21288 );
not (  , w_21289 );
and ( w_21288 , w_21289 , \4519_b0 );
or ( \6684_b1 , \6682_b1 , w_21291 );
not ( w_21291 , w_21292 );
and ( \6684_b0 , \6682_b0 , w_21293 );
and ( w_21292 ,  , w_21293 );
buf ( w_21291 , \6683_b1 );
not ( w_21291 , w_21294 );
not (  , w_21295 );
and ( w_21294 , w_21295 , \6683_b0 );
or ( \6685_b1 , \4948_b1 , w_21297 );
not ( w_21297 , w_21298 );
and ( \6685_b0 , \4948_b0 , w_21299 );
and ( w_21298 ,  , w_21299 );
buf ( w_21297 , \6684_b1 );
not ( w_21297 , w_21300 );
not (  , w_21301 );
and ( w_21300 , w_21301 , \6684_b0 );
or ( \6686_b1 , \6679_b1 , w_21303 );
not ( w_21303 , w_21304 );
and ( \6686_b0 , \6679_b0 , w_21305 );
and ( w_21304 ,  , w_21305 );
buf ( w_21303 , \6685_b1 );
not ( w_21303 , w_21306 );
not (  , w_21307 );
and ( w_21306 , w_21307 , \6685_b0 );
buf ( \6687_b1 , \6686_b1 );
not ( \6687_b1 , w_21308 );
not ( \6687_b0 , w_21309 );
and ( w_21308 , w_21309 , \6686_b0 );
or ( \6688_b1 , \6675_b1 , \6687_b1 );
xor ( \6688_b0 , \6675_b0 , w_21310 );
not ( w_21310 , w_21311 );
and ( w_21311 , \6687_b1 , \6687_b0 );
buf ( \6689_b1 , \6688_b1 );
not ( \6689_b1 , w_21312 );
not ( \6689_b0 , w_21313 );
and ( w_21312 , w_21313 , \6688_b0 );
or ( \6690_b1 , \6658_b1 , w_21314 );
or ( \6690_b0 , \6658_b0 , \6689_b0 );
not ( \6689_b0 , w_21315 );
and ( w_21315 , w_21314 , \6689_b1 );
buf ( \6691_b1 , \6492_b1 );
not ( \6691_b1 , w_21316 );
not ( \6691_b0 , w_21317 );
and ( w_21316 , w_21317 , \6492_b0 );
buf ( \6692_b1 , \4066_b1 );
not ( \6692_b1 , w_21318 );
not ( \6692_b0 , w_21319 );
and ( w_21318 , w_21319 , \4066_b0 );
buf ( \6693_b1 , \6541_b1 );
not ( \6693_b1 , w_21320 );
not ( \6693_b0 , w_21321 );
and ( w_21320 , w_21321 , \6541_b0 );
or ( \6694_b1 , \6692_b1 , w_21322 );
or ( \6694_b0 , \6692_b0 , \6693_b0 );
not ( \6693_b0 , w_21323 );
and ( w_21323 , w_21322 , \6693_b1 );
or ( \6695_b1 , \5433_b1 , w_21325 );
not ( w_21325 , w_21326 );
and ( \6695_b0 , \5433_b0 , w_21327 );
and ( w_21326 ,  , w_21327 );
buf ( w_21325 , \4519_b1 );
not ( w_21325 , w_21328 );
not (  , w_21329 );
and ( w_21328 , w_21329 , \4519_b0 );
or ( \6696_b1 , \6694_b1 , w_21331 );
not ( w_21331 , w_21332 );
and ( \6696_b0 , \6694_b0 , w_21333 );
and ( w_21332 ,  , w_21333 );
buf ( w_21331 , \6695_b1 );
not ( w_21331 , w_21334 );
not (  , w_21335 );
and ( w_21334 , w_21335 , \6695_b0 );
buf ( \6697_b1 , \6696_b1 );
not ( \6697_b1 , w_21336 );
not ( \6697_b0 , w_21337 );
and ( w_21336 , w_21337 , \6696_b0 );
or ( \6698_b1 , \6691_b1 , w_21338 );
or ( \6698_b0 , \6691_b0 , \6697_b0 );
not ( \6697_b0 , w_21339 );
and ( w_21339 , w_21338 , \6697_b1 );
or ( \6699_b1 , \6665_b1 , w_21341 );
not ( w_21341 , w_21342 );
and ( \6699_b0 , \6665_b0 , w_21343 );
and ( w_21342 ,  , w_21343 );
buf ( w_21341 , \5266_b1 );
not ( w_21341 , w_21344 );
not (  , w_21345 );
and ( w_21344 , w_21345 , \5266_b0 );
or ( \6700_b1 , \6698_b1 , w_21347 );
not ( w_21347 , w_21348 );
and ( \6700_b0 , \6698_b0 , w_21349 );
and ( w_21348 ,  , w_21349 );
buf ( w_21347 , \6699_b1 );
not ( w_21347 , w_21350 );
not (  , w_21351 );
and ( w_21350 , w_21351 , \6699_b0 );
buf ( \6701_b1 , \6700_b1 );
not ( \6701_b1 , w_21352 );
not ( \6701_b0 , w_21353 );
and ( w_21352 , w_21353 , \6700_b0 );
or ( \6702_b1 , \4079_b1 , \4917_b1 );
not ( \4917_b1 , w_21354 );
and ( \6702_b0 , \4079_b0 , w_21355 );
and ( w_21354 , w_21355 , \4917_b0 );
buf ( \6703_b1 , \4079_b1 );
not ( \6703_b1 , w_21356 );
not ( \6703_b0 , w_21357 );
and ( w_21356 , w_21357 , \4079_b0 );
or ( \6704_b1 , \6703_b1 , \4732_b1 );
not ( \4732_b1 , w_21358 );
and ( \6704_b0 , \6703_b0 , w_21359 );
and ( w_21358 , w_21359 , \4732_b0 );
or ( \6705_b1 , \6702_b1 , w_21361 );
not ( w_21361 , w_21362 );
and ( \6705_b0 , \6702_b0 , w_21363 );
and ( w_21362 ,  , w_21363 );
buf ( w_21361 , \6704_b1 );
not ( w_21361 , w_21364 );
not (  , w_21365 );
and ( w_21364 , w_21365 , \6704_b0 );
buf ( \6706_b1 , \6705_b1 );
not ( \6706_b1 , w_21366 );
not ( \6706_b0 , w_21367 );
and ( w_21366 , w_21367 , \6705_b0 );
buf ( \6707_b1 , \4632_b1 );
not ( \6707_b1 , w_21368 );
not ( \6707_b0 , w_21369 );
and ( w_21368 , w_21369 , \4632_b0 );
or ( \6708_b1 , \6706_b1 , w_21370 );
or ( \6708_b0 , \6706_b0 , \6707_b0 );
not ( \6707_b0 , w_21371 );
and ( w_21371 , w_21370 , \6707_b1 );
buf ( \6709_b1 , \4076_b1 );
not ( \6709_b1 , w_21372 );
not ( \6709_b0 , w_21373 );
and ( w_21372 , w_21373 , \4076_b0 );
buf ( \6710_b1 , \4535_b1 );
not ( \6710_b1 , w_21374 );
not ( \6710_b0 , w_21375 );
and ( w_21374 , w_21375 , \4535_b0 );
or ( \6711_b1 , \6709_b1 , w_21376 );
or ( \6711_b0 , \6709_b0 , \6710_b0 );
not ( \6710_b0 , w_21377 );
and ( w_21377 , w_21376 , \6710_b1 );
or ( \6712_b1 , \4917_b1 , w_21379 );
not ( w_21379 , w_21380 );
and ( \6712_b0 , \4917_b0 , w_21381 );
and ( w_21380 ,  , w_21381 );
buf ( w_21379 , \5284_b1 );
not ( w_21379 , w_21382 );
not (  , w_21383 );
and ( w_21382 , w_21383 , \5284_b0 );
or ( \6713_b1 , \6711_b1 , w_21385 );
not ( w_21385 , w_21386 );
and ( \6713_b0 , \6711_b0 , w_21387 );
and ( w_21386 ,  , w_21387 );
buf ( w_21385 , \6712_b1 );
not ( w_21385 , w_21388 );
not (  , w_21389 );
and ( w_21388 , w_21389 , \6712_b0 );
or ( \6714_b1 , \4453_b1 , w_21391 );
not ( w_21391 , w_21392 );
and ( \6714_b0 , \4453_b0 , w_21393 );
and ( w_21392 ,  , w_21393 );
buf ( w_21391 , \6713_b1 );
not ( w_21391 , w_21394 );
not (  , w_21395 );
and ( w_21394 , w_21395 , \6713_b0 );
or ( \6715_b1 , \6708_b1 , w_21397 );
not ( w_21397 , w_21398 );
and ( \6715_b0 , \6708_b0 , w_21399 );
and ( w_21398 ,  , w_21399 );
buf ( w_21397 , \6714_b1 );
not ( w_21397 , w_21400 );
not (  , w_21401 );
and ( w_21400 , w_21401 , \6714_b0 );
buf ( \6716_b1 , \6715_b1 );
not ( \6716_b1 , w_21402 );
not ( \6716_b0 , w_21403 );
and ( w_21402 , w_21403 , \6715_b0 );
or ( \6717_b1 , \6701_b1 , w_21404 );
or ( \6717_b0 , \6701_b0 , \6716_b0 );
not ( \6716_b0 , w_21405 );
and ( w_21405 , w_21404 , \6716_b1 );
buf ( \6718_b1 , \6715_b1 );
not ( \6718_b1 , w_21406 );
not ( \6718_b0 , w_21407 );
and ( w_21406 , w_21407 , \6715_b0 );
buf ( \6719_b1 , \6718_b1 );
not ( \6719_b1 , w_21408 );
not ( \6719_b0 , w_21409 );
and ( w_21408 , w_21409 , \6718_b0 );
buf ( \6720_b1 , \6700_b1 );
not ( \6720_b1 , w_21410 );
not ( \6720_b0 , w_21411 );
and ( w_21410 , w_21411 , \6700_b0 );
buf ( \6721_b1 , \6720_b1 );
not ( \6721_b1 , w_21412 );
not ( \6721_b0 , w_21413 );
and ( w_21412 , w_21413 , \6720_b0 );
or ( \6722_b1 , \6719_b1 , w_21414 );
or ( \6722_b0 , \6719_b0 , \6721_b0 );
not ( \6721_b0 , w_21415 );
and ( w_21415 , w_21414 , \6721_b1 );
buf ( \6723_b1 , \4098_b1 );
not ( \6723_b1 , w_21416 );
not ( \6723_b0 , w_21417 );
and ( w_21416 , w_21417 , \4098_b0 );
buf ( \6724_b1 , \4493_b1 );
not ( \6724_b1 , w_21418 );
not ( \6724_b0 , w_21419 );
and ( w_21418 , w_21419 , \4493_b0 );
or ( \6725_b1 , \6723_b1 , w_21420 );
or ( \6725_b0 , \6723_b0 , \6724_b0 );
not ( \6724_b0 , w_21421 );
and ( w_21421 , w_21420 , \6724_b1 );
or ( \6726_b1 , \4285_b1 , w_21423 );
not ( w_21423 , w_21424 );
and ( \6726_b0 , \4285_b0 , w_21425 );
and ( w_21424 ,  , w_21425 );
buf ( w_21423 , \5418_b1 );
not ( w_21423 , w_21426 );
not (  , w_21427 );
and ( w_21426 , w_21427 , \5418_b0 );
or ( \6727_b1 , \6725_b1 , w_21429 );
not ( w_21429 , w_21430 );
and ( \6727_b0 , \6725_b0 , w_21431 );
and ( w_21430 ,  , w_21431 );
buf ( w_21429 , \6726_b1 );
not ( w_21429 , w_21432 );
not (  , w_21433 );
and ( w_21432 , w_21433 , \6726_b0 );
buf ( \6728_b1 , \6727_b1 );
not ( \6728_b1 , w_21434 );
not ( \6728_b0 , w_21435 );
and ( w_21434 , w_21435 , \6727_b0 );
buf ( \6729_b1 , \4430_b1 );
not ( \6729_b1 , w_21436 );
not ( \6729_b0 , w_21437 );
and ( w_21436 , w_21437 , \4430_b0 );
or ( \6730_b1 , \6728_b1 , w_21438 );
or ( \6730_b0 , \6728_b0 , \6729_b0 );
not ( \6729_b0 , w_21439 );
and ( w_21439 , w_21438 , \6729_b1 );
buf ( \6731_b1 , \4082_b1 );
not ( \6731_b1 , w_21440 );
not ( \6731_b0 , w_21441 );
and ( w_21440 , w_21441 , \4082_b0 );
buf ( \6732_b1 , \4493_b1 );
not ( \6732_b1 , w_21442 );
not ( \6732_b0 , w_21443 );
and ( w_21442 , w_21443 , \4493_b0 );
or ( \6733_b1 , \6731_b1 , w_21444 );
or ( \6733_b0 , \6731_b0 , \6732_b0 );
not ( \6732_b0 , w_21445 );
and ( w_21445 , w_21444 , \6732_b1 );
or ( \6734_b1 , \4283_b1 , w_21447 );
not ( w_21447 , w_21448 );
and ( \6734_b0 , \4283_b0 , w_21449 );
and ( w_21448 ,  , w_21449 );
buf ( w_21447 , \5526_b1 );
not ( w_21447 , w_21450 );
not (  , w_21451 );
and ( w_21450 , w_21451 , \5526_b0 );
or ( \6735_b1 , \6733_b1 , w_21453 );
not ( w_21453 , w_21454 );
and ( \6735_b0 , \6733_b0 , w_21455 );
and ( w_21454 ,  , w_21455 );
buf ( w_21453 , \6734_b1 );
not ( w_21453 , w_21456 );
not (  , w_21457 );
and ( w_21456 , w_21457 , \6734_b0 );
or ( \6736_b1 , \6735_b1 , w_21459 );
not ( w_21459 , w_21460 );
and ( \6736_b0 , \6735_b0 , w_21461 );
and ( w_21460 ,  , w_21461 );
buf ( w_21459 , \5160_b1 );
not ( w_21459 , w_21462 );
not (  , w_21463 );
and ( w_21462 , w_21463 , \5160_b0 );
or ( \6737_b1 , \6730_b1 , w_21465 );
not ( w_21465 , w_21466 );
and ( \6737_b0 , \6730_b0 , w_21467 );
and ( w_21466 ,  , w_21467 );
buf ( w_21465 , \6736_b1 );
not ( w_21465 , w_21468 );
not (  , w_21469 );
and ( w_21468 , w_21469 , \6736_b0 );
or ( \6738_b1 , \6722_b1 , w_21471 );
not ( w_21471 , w_21472 );
and ( \6738_b0 , \6722_b0 , w_21473 );
and ( w_21472 ,  , w_21473 );
buf ( w_21471 , \6737_b1 );
not ( w_21471 , w_21474 );
not (  , w_21475 );
and ( w_21474 , w_21475 , \6737_b0 );
or ( \6739_b1 , \6717_b1 , w_21477 );
not ( w_21477 , w_21478 );
and ( \6739_b0 , \6717_b0 , w_21479 );
and ( w_21478 ,  , w_21479 );
buf ( w_21477 , \6738_b1 );
not ( w_21477 , w_21480 );
not (  , w_21481 );
and ( w_21480 , w_21481 , \6738_b0 );
or ( \6740_b1 , \6690_b1 , w_21483 );
not ( w_21483 , w_21484 );
and ( \6740_b0 , \6690_b0 , w_21485 );
and ( w_21484 ,  , w_21485 );
buf ( w_21483 , \6739_b1 );
not ( w_21483 , w_21486 );
not (  , w_21487 );
and ( w_21486 , w_21487 , \6739_b0 );
buf ( \6741_b1 , \6688_b1 );
not ( \6741_b1 , w_21488 );
not ( \6741_b0 , w_21489 );
and ( w_21488 , w_21489 , \6688_b0 );
buf ( \6742_b1 , \6657_b1 );
not ( \6742_b1 , w_21490 );
not ( \6742_b0 , w_21491 );
and ( w_21490 , w_21491 , \6657_b0 );
or ( \6743_b1 , \6741_b1 , w_21493 );
not ( w_21493 , w_21494 );
and ( \6743_b0 , \6741_b0 , w_21495 );
and ( w_21494 ,  , w_21495 );
buf ( w_21493 , \6742_b1 );
not ( w_21493 , w_21496 );
not (  , w_21497 );
and ( w_21496 , w_21497 , \6742_b0 );
or ( \6744_b1 , \6740_b1 , w_21499 );
not ( w_21499 , w_21500 );
and ( \6744_b0 , \6740_b0 , w_21501 );
and ( w_21500 ,  , w_21501 );
buf ( w_21499 , \6743_b1 );
not ( w_21499 , w_21502 );
not (  , w_21503 );
and ( w_21502 , w_21503 , \6743_b0 );
buf ( \6745_b1 , \6744_b1 );
not ( \6745_b1 , w_21504 );
not ( \6745_b0 , w_21505 );
and ( w_21504 , w_21505 , \6744_b0 );
buf ( \6746_b1 , \6745_b1 );
not ( \6746_b1 , w_21506 );
not ( \6746_b0 , w_21507 );
and ( w_21506 , w_21507 , \6745_b0 );
or ( \6747_b1 , \6635_b1 , w_21508 );
or ( \6747_b0 , \6635_b0 , \6746_b0 );
not ( \6746_b0 , w_21509 );
and ( w_21509 , w_21508 , \6746_b1 );
buf ( \6748_b1 , \6634_b1 );
not ( \6748_b1 , w_21510 );
not ( \6748_b0 , w_21511 );
and ( w_21510 , w_21511 , \6634_b0 );
or ( \6749_b1 , \6748_b1 , w_21513 );
not ( w_21513 , w_21514 );
and ( \6749_b0 , \6748_b0 , w_21515 );
and ( w_21514 ,  , w_21515 );
buf ( w_21513 , \6744_b1 );
not ( w_21513 , w_21516 );
not (  , w_21517 );
and ( w_21516 , w_21517 , \6744_b0 );
or ( \6750_b1 , \6747_b1 , w_21519 );
not ( w_21519 , w_21520 );
and ( \6750_b0 , \6747_b0 , w_21521 );
and ( w_21520 ,  , w_21521 );
buf ( w_21519 , \6749_b1 );
not ( w_21519 , w_21522 );
not (  , w_21523 );
and ( w_21522 , w_21523 , \6749_b0 );
or ( \6751_b1 , \6673_b1 , w_21525 );
not ( w_21525 , w_21526 );
and ( \6751_b0 , \6673_b0 , w_21527 );
and ( w_21526 ,  , w_21527 );
buf ( w_21525 , \6659_b1 );
not ( w_21525 , w_21528 );
not (  , w_21529 );
and ( w_21528 , w_21529 , \6659_b0 );
buf ( \6752_b1 , \6751_b1 );
not ( \6752_b1 , w_21530 );
not ( \6752_b0 , w_21531 );
and ( w_21530 , w_21531 , \6751_b0 );
buf ( \6753_b1 , \6686_b1 );
not ( \6753_b1 , w_21532 );
not ( \6753_b0 , w_21533 );
and ( w_21532 , w_21533 , \6686_b0 );
or ( \6754_b1 , \6752_b1 , w_21534 );
or ( \6754_b0 , \6752_b0 , \6753_b0 );
not ( \6753_b0 , w_21535 );
and ( w_21535 , w_21534 , \6753_b1 );
or ( \6755_b1 , \6670_b1 , w_21537 );
not ( w_21537 , w_21538 );
and ( \6755_b0 , \6670_b0 , w_21539 );
and ( w_21538 ,  , w_21539 );
buf ( w_21537 , \6660_b1 );
not ( w_21537 , w_21540 );
not (  , w_21541 );
and ( w_21540 , w_21541 , \6660_b0 );
or ( \6756_b1 , \6754_b1 , w_21543 );
not ( w_21543 , w_21544 );
and ( \6756_b0 , \6754_b0 , w_21545 );
and ( w_21544 ,  , w_21545 );
buf ( w_21543 , \6755_b1 );
not ( w_21543 , w_21546 );
not (  , w_21547 );
and ( w_21546 , w_21547 , \6755_b0 );
buf ( \6757_b1 , \4026_b1 );
not ( \6757_b1 , w_21548 );
not ( \6757_b0 , w_21549 );
and ( w_21548 , w_21549 , \4026_b0 );
buf ( \6758_b1 , \5301_b1 );
not ( \6758_b1 , w_21550 );
not ( \6758_b0 , w_21551 );
and ( w_21550 , w_21551 , \5301_b0 );
or ( \6759_b1 , \6757_b1 , w_21552 );
or ( \6759_b0 , \6757_b0 , \6758_b0 );
not ( \6758_b0 , w_21553 );
and ( w_21553 , w_21552 , \6758_b1 );
or ( \6760_b1 , \4616_b1 , w_21555 );
not ( w_21555 , w_21556 );
and ( \6760_b0 , \4616_b0 , w_21557 );
and ( w_21556 ,  , w_21557 );
buf ( w_21555 , \4969_b1 );
not ( w_21555 , w_21558 );
not (  , w_21559 );
and ( w_21558 , w_21559 , \4969_b0 );
or ( \6761_b1 , \6759_b1 , w_21561 );
not ( w_21561 , w_21562 );
and ( \6761_b0 , \6759_b0 , w_21563 );
and ( w_21562 ,  , w_21563 );
buf ( w_21561 , \6760_b1 );
not ( w_21561 , w_21564 );
not (  , w_21565 );
and ( w_21564 , w_21565 , \6760_b0 );
buf ( \6762_b1 , \6761_b1 );
not ( \6762_b1 , w_21566 );
not ( \6762_b0 , w_21567 );
and ( w_21566 , w_21567 , \6761_b0 );
buf ( \6763_b1 , \4611_b1 );
not ( \6763_b1 , w_21568 );
not ( \6763_b0 , w_21569 );
and ( w_21568 , w_21569 , \4611_b0 );
or ( \6764_b1 , \6762_b1 , w_21570 );
or ( \6764_b0 , \6762_b0 , \6763_b0 );
not ( \6763_b0 , w_21571 );
and ( w_21571 , w_21570 , \6763_b1 );
buf ( \6765_b1 , \4021_b1 );
not ( \6765_b1 , w_21572 );
not ( \6765_b0 , w_21573 );
and ( w_21572 , w_21573 , \4021_b0 );
buf ( \6766_b1 , \5138_b1 );
not ( \6766_b1 , w_21574 );
not ( \6766_b0 , w_21575 );
and ( w_21574 , w_21575 , \5138_b0 );
or ( \6767_b1 , \6765_b1 , w_21576 );
or ( \6767_b0 , \6765_b0 , \6766_b0 );
not ( \6766_b0 , w_21577 );
and ( w_21577 , w_21576 , \6766_b1 );
or ( \6768_b1 , \4745_b1 , w_21579 );
not ( w_21579 , w_21580 );
and ( \6768_b0 , \4745_b0 , w_21581 );
and ( w_21580 ,  , w_21581 );
buf ( w_21579 , \4780_b1 );
not ( w_21579 , w_21582 );
not (  , w_21583 );
and ( w_21582 , w_21583 , \4780_b0 );
or ( \6769_b1 , \6767_b1 , w_21585 );
not ( w_21585 , w_21586 );
and ( \6769_b0 , \6767_b0 , w_21587 );
and ( w_21586 ,  , w_21587 );
buf ( w_21585 , \6768_b1 );
not ( w_21585 , w_21588 );
not (  , w_21589 );
and ( w_21588 , w_21589 , \6768_b0 );
or ( \6770_b1 , \4881_b1 , w_21591 );
not ( w_21591 , w_21592 );
and ( \6770_b0 , \4881_b0 , w_21593 );
and ( w_21592 ,  , w_21593 );
buf ( w_21591 , \6769_b1 );
not ( w_21591 , w_21594 );
not (  , w_21595 );
and ( w_21594 , w_21595 , \6769_b0 );
or ( \6771_b1 , \6764_b1 , w_21597 );
not ( w_21597 , w_21598 );
and ( \6771_b0 , \6764_b0 , w_21599 );
and ( w_21598 ,  , w_21599 );
buf ( w_21597 , \6770_b1 );
not ( w_21597 , w_21600 );
not (  , w_21601 );
and ( w_21600 , w_21601 , \6770_b0 );
buf ( \6772_b1 , \6771_b1 );
not ( \6772_b1 , w_21602 );
not ( \6772_b0 , w_21603 );
and ( w_21602 , w_21603 , \6771_b0 );
buf ( \6773_b1 , \6772_b1 );
not ( \6773_b1 , w_21604 );
not ( \6773_b0 , w_21605 );
and ( w_21604 , w_21605 , \6772_b0 );
or ( \6774_b1 , \4632_b1 , \6713_b1 );
not ( \6713_b1 , w_21606 );
and ( \6774_b0 , \4632_b0 , w_21607 );
and ( w_21606 , w_21607 , \6713_b0 );
or ( \6775_b1 , \4453_b1 , \6607_b1 );
not ( \6607_b1 , w_21608 );
and ( \6775_b0 , \4453_b0 , w_21609 );
and ( w_21608 , w_21609 , \6607_b0 );
or ( \6776_b1 , \6774_b1 , w_21611 );
not ( w_21611 , w_21612 );
and ( \6776_b0 , \6774_b0 , w_21613 );
and ( w_21612 ,  , w_21613 );
buf ( w_21611 , \6775_b1 );
not ( w_21611 , w_21614 );
not (  , w_21615 );
and ( w_21614 , w_21615 , \6775_b0 );
buf ( \6777_b1 , \6776_b1 );
not ( \6777_b1 , w_21616 );
not ( \6777_b0 , w_21617 );
and ( w_21616 , w_21617 , \6776_b0 );
or ( \6778_b1 , \6773_b1 , w_21618 );
or ( \6778_b0 , \6773_b0 , \6777_b0 );
not ( \6777_b0 , w_21619 );
and ( w_21619 , w_21618 , \6777_b1 );
buf ( \6779_b1 , \6735_b1 );
not ( \6779_b1 , w_21620 );
not ( \6779_b0 , w_21621 );
and ( w_21620 , w_21621 , \6735_b0 );
buf ( \6780_b1 , \4338_b1 );
not ( \6780_b1 , w_21622 );
not ( \6780_b0 , w_21623 );
and ( w_21622 , w_21623 , \4338_b0 );
or ( \6781_b1 , \6779_b1 , w_21624 );
or ( \6781_b0 , \6779_b0 , \6780_b0 );
not ( \6780_b0 , w_21625 );
and ( w_21625 , w_21624 , \6780_b1 );
or ( \6782_b1 , \6628_b1 , w_21627 );
not ( w_21627 , w_21628 );
and ( \6782_b0 , \6628_b0 , w_21629 );
and ( w_21628 ,  , w_21629 );
buf ( w_21627 , \4341_b1 );
not ( w_21627 , w_21630 );
not (  , w_21631 );
and ( w_21630 , w_21631 , \4341_b0 );
or ( \6783_b1 , \6781_b1 , w_21633 );
not ( w_21633 , w_21634 );
and ( \6783_b0 , \6781_b0 , w_21635 );
and ( w_21634 ,  , w_21635 );
buf ( w_21633 , \6782_b1 );
not ( w_21633 , w_21636 );
not (  , w_21637 );
and ( w_21636 , w_21637 , \6782_b0 );
or ( \6784_b1 , \6778_b1 , w_21639 );
not ( w_21639 , w_21640 );
and ( \6784_b0 , \6778_b0 , w_21641 );
and ( w_21640 ,  , w_21641 );
buf ( w_21639 , \6783_b1 );
not ( w_21639 , w_21642 );
not (  , w_21643 );
and ( w_21642 , w_21643 , \6783_b0 );
buf ( \6785_b1 , \6776_b1 );
not ( \6785_b1 , w_21644 );
not ( \6785_b0 , w_21645 );
and ( w_21644 , w_21645 , \6776_b0 );
or ( \6786_b1 , \6785_b1 , w_21647 );
not ( w_21647 , w_21648 );
and ( \6786_b0 , \6785_b0 , w_21649 );
and ( w_21648 ,  , w_21649 );
buf ( w_21647 , \6771_b1 );
not ( w_21647 , w_21650 );
not (  , w_21651 );
and ( w_21650 , w_21651 , \6771_b0 );
or ( \6787_b1 , \6784_b1 , w_21653 );
not ( w_21653 , w_21654 );
and ( \6787_b0 , \6784_b0 , w_21655 );
and ( w_21654 ,  , w_21655 );
buf ( w_21653 , \6786_b1 );
not ( w_21653 , w_21656 );
not (  , w_21657 );
and ( w_21656 , w_21657 , \6786_b0 );
or ( \6788_b1 , \6756_b1 , \6787_b1 );
xor ( \6788_b0 , \6756_b0 , w_21658 );
not ( w_21658 , w_21659 );
and ( w_21659 , \6787_b1 , \6787_b0 );
buf ( \6789_b1 , \6769_b1 );
not ( \6789_b1 , w_21660 );
not ( \6789_b0 , w_21661 );
and ( w_21660 , w_21661 , \6769_b0 );
buf ( \6790_b1 , \4610_b1 );
not ( \6790_b1 , w_21662 );
not ( \6790_b0 , w_21663 );
and ( w_21662 , w_21663 , \4610_b0 );
or ( \6791_b1 , \6789_b1 , w_21664 );
or ( \6791_b0 , \6789_b0 , \6790_b0 );
not ( \6790_b0 , w_21665 );
and ( w_21665 , w_21664 , \6790_b1 );
buf ( \6792_b1 , \4017_b1 );
not ( \6792_b1 , w_21666 );
not ( \6792_b0 , w_21667 );
and ( w_21666 , w_21667 , \4017_b0 );
buf ( \6793_b1 , \5138_b1 );
not ( \6793_b1 , w_21668 );
not ( \6793_b0 , w_21669 );
and ( w_21668 , w_21669 , \5138_b0 );
or ( \6794_b1 , \6792_b1 , w_21670 );
or ( \6794_b0 , \6792_b0 , \6793_b0 );
not ( \6793_b0 , w_21671 );
and ( w_21671 , w_21670 , \6793_b1 );
or ( \6795_b1 , \4745_b1 , w_21673 );
not ( w_21673 , w_21674 );
and ( \6795_b0 , \4745_b0 , w_21675 );
and ( w_21674 ,  , w_21675 );
buf ( w_21673 , \4662_b1 );
not ( w_21673 , w_21676 );
not (  , w_21677 );
and ( w_21676 , w_21677 , \4662_b0 );
or ( \6796_b1 , \6794_b1 , w_21679 );
not ( w_21679 , w_21680 );
and ( \6796_b0 , \6794_b0 , w_21681 );
and ( w_21680 ,  , w_21681 );
buf ( w_21679 , \6795_b1 );
not ( w_21679 , w_21682 );
not (  , w_21683 );
and ( w_21682 , w_21683 , \6795_b0 );
or ( \6797_b1 , \6796_b1 , w_21685 );
not ( w_21685 , w_21686 );
and ( \6797_b0 , \6796_b0 , w_21687 );
and ( w_21686 ,  , w_21687 );
buf ( w_21685 , \5146_b1 );
not ( w_21685 , w_21688 );
not (  , w_21689 );
and ( w_21688 , w_21689 , \5146_b0 );
or ( \6798_b1 , \6791_b1 , w_21691 );
not ( w_21691 , w_21692 );
and ( \6798_b0 , \6791_b0 , w_21693 );
and ( w_21692 ,  , w_21693 );
buf ( w_21691 , \6797_b1 );
not ( w_21691 , w_21694 );
not (  , w_21695 );
and ( w_21694 , w_21695 , \6797_b0 );
or ( \6799_b1 , \4098_b1 , w_21697 );
not ( w_21697 , w_21698 );
and ( \6799_b0 , \4098_b0 , w_21699 );
and ( w_21698 ,  , w_21699 );
buf ( w_21697 , \3573_b1 );
not ( w_21697 , w_21700 );
not (  , w_21701 );
and ( w_21700 , w_21701 , \3573_b0 );
buf ( \6800_b1 , \6799_b1 );
not ( \6800_b1 , w_21702 );
not ( \6800_b0 , w_21703 );
and ( w_21702 , w_21703 , \6799_b0 );
buf ( \6801_b1 , \4284_b1 );
not ( \6801_b1 , w_21704 );
not ( \6801_b0 , w_21705 );
and ( w_21704 , w_21705 , \4284_b0 );
or ( \6802_b1 , \6800_b1 , \6801_b1 );
not ( \6801_b1 , w_21706 );
and ( \6802_b0 , \6800_b0 , w_21707 );
and ( w_21706 , w_21707 , \6801_b0 );
buf ( \6803_b1 , \4098_b1 );
not ( \6803_b1 , w_21708 );
not ( \6803_b0 , w_21709 );
and ( w_21708 , w_21709 , \4098_b0 );
buf ( \6804_b1 , \3573_b1 );
not ( \6804_b1 , w_21710 );
not ( \6804_b0 , w_21711 );
and ( w_21710 , w_21711 , \3573_b0 );
or ( \6805_b1 , \6803_b1 , w_21712 );
or ( \6805_b0 , \6803_b0 , \6804_b0 );
not ( \6804_b0 , w_21713 );
and ( w_21713 , w_21712 , \6804_b1 );
or ( \6806_b1 , \6805_b1 , w_21715 );
not ( w_21715 , w_21716 );
and ( \6806_b0 , \6805_b0 , w_21717 );
and ( w_21716 ,  , w_21717 );
buf ( w_21715 , \4154_b1 );
not ( w_21715 , w_21718 );
not (  , w_21719 );
and ( w_21718 , w_21719 , \4154_b0 );
or ( \6807_b1 , \6802_b1 , w_21721 );
not ( w_21721 , w_21722 );
and ( \6807_b0 , \6802_b0 , w_21723 );
and ( w_21722 ,  , w_21723 );
buf ( w_21721 , \6806_b1 );
not ( w_21721 , w_21724 );
not (  , w_21725 );
and ( w_21724 , w_21725 , \6806_b0 );
buf ( \6808_b1 , \6807_b1 );
not ( \6808_b1 , w_21726 );
not ( \6808_b0 , w_21727 );
and ( w_21726 , w_21727 , \6807_b0 );
or ( \6809_b1 , \6180_b1 , w_21728 );
or ( \6809_b0 , \6180_b0 , \4862_b0 );
not ( \4862_b0 , w_21729 );
and ( w_21729 , w_21728 , \4862_b1 );
or ( \6811_b1 , \6809_b1 , w_21731 );
not ( w_21731 , w_21732 );
and ( \6811_b0 , \6809_b0 , w_21733 );
and ( w_21732 ,  , w_21733 );
buf ( w_21731 , \6810_b1 );
not ( w_21731 , w_21734 );
not (  , w_21735 );
and ( w_21734 , w_21735 , \6810_b0 );
buf ( \6812_b1 , \6811_b1 );
not ( \6812_b1 , w_21736 );
not ( \6812_b0 , w_21737 );
and ( w_21736 , w_21737 , \6811_b0 );
buf ( \6813_b1 , \6812_b1 );
not ( \6813_b1 , w_21738 );
not ( \6813_b0 , w_21739 );
and ( w_21738 , w_21739 , \6812_b0 );
or ( \6814_b1 , \6808_b1 , w_21740 );
or ( \6814_b0 , \6808_b0 , \6813_b0 );
not ( \6813_b0 , w_21741 );
and ( w_21741 , w_21740 , \6813_b1 );
or ( \6815_b1 , \6812_b1 , w_21742 );
or ( \6815_b0 , \6812_b0 , \6807_b0 );
not ( \6807_b0 , w_21743 );
and ( w_21743 , w_21742 , \6807_b1 );
or ( \6816_b1 , \6814_b1 , w_21745 );
not ( w_21745 , w_21746 );
and ( \6816_b0 , \6814_b0 , w_21747 );
and ( w_21746 ,  , w_21747 );
buf ( w_21745 , \6815_b1 );
not ( w_21745 , w_21748 );
not (  , w_21749 );
and ( w_21748 , w_21749 , \6815_b0 );
or ( \6817_b1 , \6798_b1 , \6816_b1 );
xor ( \6817_b0 , \6798_b0 , w_21750 );
not ( w_21750 , w_21751 );
and ( w_21751 , \6816_b1 , \6816_b0 );
buf ( \6818_b1 , \4098_b1 );
not ( \6818_b1 , w_21752 );
not ( \6818_b0 , w_21753 );
and ( w_21752 , w_21753 , \4098_b0 );
buf ( \6819_b1 , \4163_b1 );
not ( \6819_b1 , w_21754 );
not ( \6819_b0 , w_21755 );
and ( w_21754 , w_21755 , \4163_b0 );
or ( \6820_b1 , \6818_b1 , w_21756 );
or ( \6820_b0 , \6818_b0 , \6819_b0 );
not ( \6819_b0 , w_21757 );
and ( w_21757 , w_21756 , \6819_b1 );
or ( \6821_b1 , \4170_b1 , w_21759 );
not ( w_21759 , w_21760 );
and ( \6821_b0 , \4170_b0 , w_21761 );
and ( w_21760 ,  , w_21761 );
buf ( w_21759 , \5418_b1 );
not ( w_21759 , w_21762 );
not (  , w_21763 );
and ( w_21762 , w_21763 , \5418_b0 );
or ( \6822_b1 , \6820_b1 , w_21765 );
not ( w_21765 , w_21766 );
and ( \6822_b0 , \6820_b0 , w_21767 );
and ( w_21766 ,  , w_21767 );
buf ( w_21765 , \6821_b1 );
not ( w_21765 , w_21768 );
not (  , w_21769 );
and ( w_21768 , w_21769 , \6821_b0 );
buf ( \6823_b1 , \6822_b1 );
not ( \6823_b1 , w_21770 );
not ( \6823_b0 , w_21771 );
and ( w_21770 , w_21771 , \6822_b0 );
buf ( \6824_b1 , \4159_b1 );
not ( \6824_b1 , w_21772 );
not ( \6824_b0 , w_21773 );
and ( w_21772 , w_21773 , \4159_b0 );
or ( \6825_b1 , \6823_b1 , w_21774 );
or ( \6825_b0 , \6823_b0 , \6824_b0 );
not ( \6824_b0 , w_21775 );
and ( w_21775 , w_21774 , \6824_b1 );
or ( \6826_b1 , \4317_b1 , w_21777 );
not ( w_21777 , w_21778 );
and ( \6826_b0 , \4317_b0 , w_21779 );
and ( w_21778 ,  , w_21779 );
buf ( w_21777 , \6211_b1 );
not ( w_21777 , w_21780 );
not (  , w_21781 );
and ( w_21780 , w_21781 , \6211_b0 );
or ( \6827_b1 , \6825_b1 , w_21783 );
not ( w_21783 , w_21784 );
and ( \6827_b0 , \6825_b0 , w_21785 );
and ( w_21784 ,  , w_21785 );
buf ( w_21783 , \6826_b1 );
not ( w_21783 , w_21786 );
not (  , w_21787 );
and ( w_21786 , w_21787 , \6826_b0 );
or ( \6828_b1 , \6817_b1 , \6827_b1 );
xor ( \6828_b0 , \6817_b0 , w_21788 );
not ( w_21788 , w_21789 );
and ( w_21789 , \6827_b1 , \6827_b0 );
or ( \6829_b1 , \6788_b1 , \6828_b1 );
xor ( \6829_b0 , \6788_b0 , w_21790 );
not ( w_21790 , w_21791 );
and ( w_21791 , \6828_b1 , \6828_b0 );
buf ( \6830_b1 , \6829_b1 );
not ( \6830_b1 , w_21792 );
not ( \6830_b0 , w_21793 );
and ( w_21792 , w_21793 , \6829_b0 );
or ( \6831_b1 , \6750_b1 , \6830_b1 );
not ( \6830_b1 , w_21794 );
and ( \6831_b0 , \6750_b0 , w_21795 );
and ( w_21794 , w_21795 , \6830_b0 );
buf ( \6832_b1 , \6750_b1 );
not ( \6832_b1 , w_21796 );
not ( \6832_b0 , w_21797 );
and ( w_21796 , w_21797 , \6750_b0 );
or ( \6833_b1 , \6832_b1 , \6829_b1 );
not ( \6829_b1 , w_21798 );
and ( \6833_b0 , \6832_b0 , w_21799 );
and ( w_21798 , w_21799 , \6829_b0 );
or ( \6834_b1 , \6831_b1 , w_21801 );
not ( w_21801 , w_21802 );
and ( \6834_b0 , \6831_b0 , w_21803 );
and ( w_21802 ,  , w_21803 );
buf ( w_21801 , \6833_b1 );
not ( w_21801 , w_21804 );
not (  , w_21805 );
and ( w_21804 , w_21805 , \6833_b0 );
buf ( \6835_b1 , \4072_b1 );
not ( \6835_b1 , w_21806 );
not ( \6835_b0 , w_21807 );
and ( w_21806 , w_21807 , \4072_b0 );
buf ( \6836_b1 , \5138_b1 );
not ( \6836_b1 , w_21808 );
not ( \6836_b0 , w_21809 );
and ( w_21808 , w_21809 , \5138_b0 );
or ( \6837_b1 , \6835_b1 , w_21810 );
or ( \6837_b0 , \6835_b0 , \6836_b0 );
not ( \6836_b0 , w_21811 );
and ( w_21811 , w_21810 , \6836_b1 );
or ( \6838_b1 , \4616_b1 , w_21813 );
not ( w_21813 , w_21814 );
and ( \6838_b0 , \4616_b0 , w_21815 );
and ( w_21814 ,  , w_21815 );
buf ( w_21813 , \5089_b1 );
not ( w_21813 , w_21816 );
not (  , w_21817 );
and ( w_21816 , w_21817 , \5089_b0 );
or ( \6839_b1 , \6837_b1 , w_21819 );
not ( w_21819 , w_21820 );
and ( \6839_b0 , \6837_b0 , w_21821 );
and ( w_21820 ,  , w_21821 );
buf ( w_21819 , \6838_b1 );
not ( w_21819 , w_21822 );
not (  , w_21823 );
and ( w_21822 , w_21823 , \6838_b0 );
buf ( \6840_b1 , \6839_b1 );
not ( \6840_b1 , w_21824 );
not ( \6840_b0 , w_21825 );
and ( w_21824 , w_21825 , \6839_b0 );
buf ( \6841_b1 , \4611_b1 );
not ( \6841_b1 , w_21826 );
not ( \6841_b0 , w_21827 );
and ( w_21826 , w_21827 , \4611_b0 );
or ( \6842_b1 , \6840_b1 , w_21828 );
or ( \6842_b0 , \6840_b0 , \6841_b0 );
not ( \6841_b0 , w_21829 );
and ( w_21829 , w_21828 , \6841_b1 );
or ( \6843_b1 , \4754_b1 , w_21831 );
not ( w_21831 , w_21832 );
and ( \6843_b0 , \4754_b0 , w_21833 );
and ( w_21832 ,  , w_21833 );
buf ( w_21831 , \6761_b1 );
not ( w_21831 , w_21834 );
not (  , w_21835 );
and ( w_21834 , w_21835 , \6761_b0 );
or ( \6844_b1 , \6842_b1 , w_21837 );
not ( w_21837 , w_21838 );
and ( \6844_b0 , \6842_b0 , w_21839 );
and ( w_21838 ,  , w_21839 );
buf ( w_21837 , \6843_b1 );
not ( w_21837 , w_21840 );
not (  , w_21841 );
and ( w_21840 , w_21841 , \6843_b0 );
buf ( \6845_b1 , \6844_b1 );
buf ( \6845_b0 , \6844_b0 );
buf ( \6846_b1 , \6845_b1 );
not ( \6846_b1 , w_21842 );
not ( \6846_b0 , w_21843 );
and ( w_21842 , w_21843 , \6845_b0 );
buf ( \6847_b1 , \6656_b1 );
not ( \6847_b1 , w_21844 );
not ( \6847_b0 , w_21845 );
and ( w_21844 , w_21845 , \6656_b0 );
buf ( \6848_b1 , \6650_b1 );
not ( \6848_b1 , w_21846 );
not ( \6848_b0 , w_21847 );
and ( w_21846 , w_21847 , \6650_b0 );
buf ( \6849_b1 , \6848_b1 );
not ( \6849_b1 , w_21848 );
not ( \6849_b0 , w_21849 );
and ( w_21848 , w_21849 , \6848_b0 );
or ( \6850_b1 , \6847_b1 , w_21850 );
or ( \6850_b0 , \6847_b0 , \6849_b0 );
not ( \6849_b0 , w_21851 );
and ( w_21851 , w_21850 , \6849_b1 );
buf ( \6851_b1 , \6656_b1 );
not ( \6851_b1 , w_21852 );
not ( \6851_b0 , w_21853 );
and ( w_21852 , w_21853 , \6656_b0 );
or ( \6852_b1 , \6851_b1 , w_21855 );
not ( w_21855 , w_21856 );
and ( \6852_b0 , \6851_b0 , w_21857 );
and ( w_21856 ,  , w_21857 );
buf ( w_21855 , \6650_b1 );
not ( w_21855 , w_21858 );
not (  , w_21859 );
and ( w_21858 , w_21859 , \6650_b0 );
or ( \6853_b1 , \6850_b1 , w_21861 );
not ( w_21861 , w_21862 );
and ( \6853_b0 , \6850_b0 , w_21863 );
and ( w_21862 ,  , w_21863 );
buf ( w_21861 , \6852_b1 );
not ( w_21861 , w_21864 );
not (  , w_21865 );
and ( w_21864 , w_21865 , \6852_b0 );
buf ( \6854_b1 , \6853_b1 );
buf ( \6854_b0 , \6853_b0 );
buf ( \6855_b1 , \6854_b1 );
not ( \6855_b1 , w_21866 );
not ( \6855_b0 , w_21867 );
and ( w_21866 , w_21867 , \6854_b0 );
or ( \6856_b1 , \6846_b1 , w_21868 );
or ( \6856_b0 , \6846_b0 , \6855_b0 );
not ( \6855_b0 , w_21869 );
and ( w_21869 , w_21868 , \6855_b1 );
or ( \6857_b1 , \6854_b1 , w_21870 );
or ( \6857_b0 , \6854_b0 , \6845_b0 );
not ( \6845_b0 , w_21871 );
and ( w_21871 , w_21870 , \6845_b1 );
or ( \6858_b1 , \4800_b1 , w_21873 );
not ( w_21873 , w_21874 );
and ( \6858_b0 , \4800_b0 , w_21875 );
and ( w_21874 ,  , w_21875 );
buf ( w_21873 , \4098_b1 );
not ( w_21873 , w_21876 );
not (  , w_21877 );
and ( w_21876 , w_21877 , \4098_b0 );
buf ( \6859_b1 , \6858_b1 );
not ( \6859_b1 , w_21878 );
not ( \6859_b0 , w_21879 );
and ( w_21878 , w_21879 , \6858_b0 );
buf ( \6860_b1 , \6859_b1 );
not ( \6860_b1 , w_21880 );
not ( \6860_b0 , w_21881 );
and ( w_21880 , w_21881 , \6859_b0 );
or ( \6861_b1 , \6382_b1 , w_21883 );
not ( w_21883 , w_21884 );
and ( \6861_b0 , \6382_b0 , w_21885 );
and ( w_21884 ,  , w_21885 );
buf ( w_21883 , \4859_b1 );
not ( w_21883 , w_21886 );
not (  , w_21887 );
and ( w_21886 , w_21887 , \4859_b0 );
or ( \6862_b1 , \6861_b1 , w_21888 );
or ( \6862_b0 , \6861_b0 , \4948_b0 );
not ( \4948_b0 , w_21889 );
and ( w_21889 , w_21888 , \4948_b1 );
or ( \6863_b1 , \4863_b1 , w_21891 );
not ( w_21891 , w_21892 );
and ( \6863_b0 , \4863_b0 , w_21893 );
and ( w_21892 ,  , w_21893 );
buf ( w_21891 , \6646_b1 );
not ( w_21891 , w_21894 );
not (  , w_21895 );
and ( w_21894 , w_21895 , \6646_b0 );
or ( \6864_b1 , \6862_b1 , w_21897 );
not ( w_21897 , w_21898 );
and ( \6864_b0 , \6862_b0 , w_21899 );
and ( w_21898 ,  , w_21899 );
buf ( w_21897 , \6863_b1 );
not ( w_21897 , w_21900 );
not (  , w_21901 );
and ( w_21900 , w_21901 , \6863_b0 );
buf ( \6865_b1 , \6864_b1 );
not ( \6865_b1 , w_21902 );
not ( \6865_b0 , w_21903 );
and ( w_21902 , w_21903 , \6864_b0 );
or ( \6866_b1 , \6860_b1 , w_21904 );
or ( \6866_b0 , \6860_b0 , \6865_b0 );
not ( \6865_b0 , w_21905 );
and ( w_21905 , w_21904 , \6865_b1 );
or ( \6867_b1 , \6864_b1 , w_21906 );
or ( \6867_b0 , \6864_b0 , \6859_b0 );
not ( \6859_b0 , w_21907 );
and ( w_21907 , w_21906 , \6859_b1 );
buf ( \6868_b1 , \6423_b1 );
not ( \6868_b1 , w_21908 );
not ( \6868_b0 , w_21909 );
and ( w_21908 , w_21909 , \6423_b0 );
buf ( \6869_b1 , \4632_b1 );
not ( \6869_b1 , w_21910 );
not ( \6869_b0 , w_21911 );
and ( w_21910 , w_21911 , \4632_b0 );
or ( \6870_b1 , \6868_b1 , w_21912 );
or ( \6870_b0 , \6868_b0 , \6869_b0 );
not ( \6869_b0 , w_21913 );
and ( w_21913 , w_21912 , \6869_b1 );
or ( \6871_b1 , \4453_b1 , w_21915 );
not ( w_21915 , w_21916 );
and ( \6871_b0 , \4453_b0 , w_21917 );
and ( w_21916 ,  , w_21917 );
buf ( w_21915 , \6705_b1 );
not ( w_21915 , w_21918 );
not (  , w_21919 );
and ( w_21918 , w_21919 , \6705_b0 );
or ( \6872_b1 , \6870_b1 , w_21921 );
not ( w_21921 , w_21922 );
and ( \6872_b0 , \6870_b0 , w_21923 );
and ( w_21922 ,  , w_21923 );
buf ( w_21921 , \6871_b1 );
not ( w_21921 , w_21924 );
not (  , w_21925 );
and ( w_21924 , w_21925 , \6871_b0 );
or ( \6873_b1 , \6867_b1 , w_21927 );
not ( w_21927 , w_21928 );
and ( \6873_b0 , \6867_b0 , w_21929 );
and ( w_21928 ,  , w_21929 );
buf ( w_21927 , \6872_b1 );
not ( w_21927 , w_21930 );
not (  , w_21931 );
and ( w_21930 , w_21931 , \6872_b0 );
or ( \6874_b1 , \6866_b1 , w_21933 );
not ( w_21933 , w_21934 );
and ( \6874_b0 , \6866_b0 , w_21935 );
and ( w_21934 ,  , w_21935 );
buf ( w_21933 , \6873_b1 );
not ( w_21933 , w_21936 );
not (  , w_21937 );
and ( w_21936 , w_21937 , \6873_b0 );
or ( \6875_b1 , \6857_b1 , w_21939 );
not ( w_21939 , w_21940 );
and ( \6875_b0 , \6857_b0 , w_21941 );
and ( w_21940 ,  , w_21941 );
buf ( w_21939 , \6874_b1 );
not ( w_21939 , w_21942 );
not (  , w_21943 );
and ( w_21942 , w_21943 , \6874_b0 );
or ( \6876_b1 , \6856_b1 , w_21945 );
not ( w_21945 , w_21946 );
and ( \6876_b0 , \6856_b0 , w_21947 );
and ( w_21946 ,  , w_21947 );
buf ( w_21945 , \6875_b1 );
not ( w_21945 , w_21948 );
not (  , w_21949 );
and ( w_21948 , w_21949 , \6875_b0 );
buf ( \6877_b1 , \6876_b1 );
not ( \6877_b1 , w_21950 );
not ( \6877_b0 , w_21951 );
and ( w_21950 , w_21951 , \6876_b0 );
buf ( \6878_b1 , \6783_b1 );
not ( \6878_b1 , w_21952 );
not ( \6878_b0 , w_21953 );
and ( w_21952 , w_21953 , \6783_b0 );
buf ( \6879_b1 , \6772_b1 );
not ( \6879_b1 , w_21954 );
not ( \6879_b0 , w_21955 );
and ( w_21954 , w_21955 , \6772_b0 );
or ( \6880_b1 , \6878_b1 , w_21956 );
or ( \6880_b0 , \6878_b0 , \6879_b0 );
not ( \6879_b0 , w_21957 );
and ( w_21957 , w_21956 , \6879_b1 );
or ( \6881_b1 , \6783_b1 , w_21958 );
or ( \6881_b0 , \6783_b0 , \6772_b0 );
not ( \6772_b0 , w_21959 );
and ( w_21959 , w_21958 , \6772_b1 );
or ( \6882_b1 , \6880_b1 , w_21961 );
not ( w_21961 , w_21962 );
and ( \6882_b0 , \6880_b0 , w_21963 );
and ( w_21962 ,  , w_21963 );
buf ( w_21961 , \6881_b1 );
not ( w_21961 , w_21964 );
not (  , w_21965 );
and ( w_21964 , w_21965 , \6881_b0 );
buf ( \6883_b1 , \6776_b1 );
buf ( \6883_b0 , \6776_b0 );
buf ( \6884_b1 , \6883_b1 );
not ( \6884_b1 , w_21966 );
not ( \6884_b0 , w_21967 );
and ( w_21966 , w_21967 , \6883_b0 );
or ( \6885_b1 , \6882_b1 , \6884_b1 );
not ( \6884_b1 , w_21968 );
and ( \6885_b0 , \6882_b0 , w_21969 );
and ( w_21968 , w_21969 , \6884_b0 );
buf ( \6886_b1 , \6882_b1 );
not ( \6886_b1 , w_21970 );
not ( \6886_b0 , w_21971 );
and ( w_21970 , w_21971 , \6882_b0 );
or ( \6887_b1 , \6886_b1 , \6883_b1 );
not ( \6883_b1 , w_21972 );
and ( \6887_b0 , \6886_b0 , w_21973 );
and ( w_21972 , w_21973 , \6883_b0 );
or ( \6888_b1 , \6885_b1 , w_21975 );
not ( w_21975 , w_21976 );
and ( \6888_b0 , \6885_b0 , w_21977 );
and ( w_21976 ,  , w_21977 );
buf ( w_21975 , \6887_b1 );
not ( w_21975 , w_21978 );
not (  , w_21979 );
and ( w_21978 , w_21979 , \6887_b0 );
buf ( \6889_b1 , \6888_b1 );
not ( \6889_b1 , w_21980 );
not ( \6889_b0 , w_21981 );
and ( w_21980 , w_21981 , \6888_b0 );
or ( \6890_b1 , \6877_b1 , w_21983 );
not ( w_21983 , w_21984 );
and ( \6890_b0 , \6877_b0 , w_21985 );
and ( w_21984 ,  , w_21985 );
buf ( w_21983 , \6889_b1 );
not ( w_21983 , w_21986 );
not (  , w_21987 );
and ( w_21986 , w_21987 , \6889_b0 );
buf ( \6891_b1 , \6890_b1 );
not ( \6891_b1 , w_21988 );
not ( \6891_b0 , w_21989 );
and ( w_21988 , w_21989 , \6890_b0 );
buf ( \6892_b1 , \6742_b1 );
not ( \6892_b1 , w_21990 );
not ( \6892_b0 , w_21991 );
and ( w_21990 , w_21991 , \6742_b0 );
buf ( \6893_b1 , \6688_b1 );
not ( \6893_b1 , w_21992 );
not ( \6893_b0 , w_21993 );
and ( w_21992 , w_21993 , \6688_b0 );
or ( \6894_b1 , \6892_b1 , w_21994 );
or ( \6894_b0 , \6892_b0 , \6893_b0 );
not ( \6893_b0 , w_21995 );
and ( w_21995 , w_21994 , \6893_b1 );
or ( \6895_b1 , \6741_b1 , w_21997 );
not ( w_21997 , w_21998 );
and ( \6895_b0 , \6741_b0 , w_21999 );
and ( w_21998 ,  , w_21999 );
buf ( w_21997 , \6657_b1 );
not ( w_21997 , w_22000 );
not (  , w_22001 );
and ( w_22000 , w_22001 , \6657_b0 );
or ( \6896_b1 , \6894_b1 , w_22003 );
not ( w_22003 , w_22004 );
and ( \6896_b0 , \6894_b0 , w_22005 );
and ( w_22004 ,  , w_22005 );
buf ( w_22003 , \6895_b1 );
not ( w_22003 , w_22006 );
not (  , w_22007 );
and ( w_22006 , w_22007 , \6895_b0 );
or ( \6897_b1 , \6896_b1 , \6739_b1 );
not ( \6739_b1 , w_22008 );
and ( \6897_b0 , \6896_b0 , w_22009 );
and ( w_22008 , w_22009 , \6739_b0 );
buf ( \6898_b1 , \6896_b1 );
not ( \6898_b1 , w_22010 );
not ( \6898_b0 , w_22011 );
and ( w_22010 , w_22011 , \6896_b0 );
buf ( \6899_b1 , \6739_b1 );
not ( \6899_b1 , w_22012 );
not ( \6899_b0 , w_22013 );
and ( w_22012 , w_22013 , \6739_b0 );
or ( \6900_b1 , \6898_b1 , \6899_b1 );
not ( \6899_b1 , w_22014 );
and ( \6900_b0 , \6898_b0 , w_22015 );
and ( w_22014 , w_22015 , \6899_b0 );
or ( \6901_b1 , \6897_b1 , w_22017 );
not ( w_22017 , w_22018 );
and ( \6901_b0 , \6897_b0 , w_22019 );
and ( w_22018 ,  , w_22019 );
buf ( w_22017 , \6900_b1 );
not ( w_22017 , w_22020 );
not (  , w_22021 );
and ( w_22020 , w_22021 , \6900_b0 );
buf ( \6902_b1 , \6901_b1 );
not ( \6902_b1 , w_22022 );
not ( \6902_b0 , w_22023 );
and ( w_22022 , w_22023 , \6901_b0 );
or ( \6903_b1 , \6891_b1 , w_22024 );
or ( \6903_b0 , \6891_b0 , \6902_b0 );
not ( \6902_b0 , w_22025 );
and ( w_22025 , w_22024 , \6902_b1 );
buf ( \6904_b1 , \6877_b1 );
not ( \6904_b1 , w_22026 );
not ( \6904_b0 , w_22027 );
and ( w_22026 , w_22027 , \6877_b0 );
or ( \6905_b1 , \6904_b1 , w_22029 );
not ( w_22029 , w_22030 );
and ( \6905_b0 , \6904_b0 , w_22031 );
and ( w_22030 ,  , w_22031 );
buf ( w_22029 , \6888_b1 );
not ( w_22029 , w_22032 );
not (  , w_22033 );
and ( w_22032 , w_22033 , \6888_b0 );
or ( \6906_b1 , \6903_b1 , w_22035 );
not ( w_22035 , w_22036 );
and ( \6906_b0 , \6903_b0 , w_22037 );
and ( w_22036 ,  , w_22037 );
buf ( w_22035 , \6905_b1 );
not ( w_22035 , w_22038 );
not (  , w_22039 );
and ( w_22038 , w_22039 , \6905_b0 );
buf ( \6907_b1 , \6906_b1 );
not ( \6907_b1 , w_22040 );
not ( \6907_b0 , w_22041 );
and ( w_22040 , w_22041 , \6906_b0 );
or ( \6908_b1 , \6834_b1 , w_22043 );
not ( w_22043 , w_22044 );
and ( \6908_b0 , \6834_b0 , w_22045 );
and ( w_22044 ,  , w_22045 );
buf ( w_22043 , \6907_b1 );
not ( w_22043 , w_22046 );
not (  , w_22047 );
and ( w_22046 , w_22047 , \6907_b0 );
or ( \6909_b1 , \6700_b1 , \6737_b1 );
xor ( \6909_b0 , \6700_b0 , w_22048 );
not ( w_22048 , w_22049 );
and ( w_22049 , \6737_b1 , \6737_b0 );
or ( \6910_b1 , \6909_b1 , w_22050 );
xor ( \6910_b0 , \6909_b0 , w_22052 );
not ( w_22052 , w_22053 );
and ( w_22053 , w_22050 , w_22051 );
buf ( w_22050 , \6715_b1 );
not ( w_22050 , w_22054 );
not ( w_22051 , w_22055 );
and ( w_22054 , w_22055 , \6715_b0 );
or ( \6911_b1 , \6384_b1 , w_22057 );
not ( w_22057 , w_22058 );
and ( \6911_b0 , \6384_b0 , w_22059 );
and ( w_22058 ,  , w_22059 );
buf ( w_22057 , \6372_b1 );
not ( w_22057 , w_22060 );
not (  , w_22061 );
and ( w_22060 , w_22061 , \6372_b0 );
buf ( \6912_b1 , \6911_b1 );
not ( \6912_b1 , w_22062 );
not ( \6912_b0 , w_22063 );
and ( w_22062 , w_22063 , \6911_b0 );
buf ( \6913_b1 , \6410_b1 );
not ( \6913_b1 , w_22064 );
not ( \6913_b0 , w_22065 );
and ( w_22064 , w_22065 , \6410_b0 );
buf ( \6914_b1 , \4611_b1 );
not ( \6914_b1 , w_22066 );
not ( \6914_b0 , w_22067 );
and ( w_22066 , w_22067 , \4611_b0 );
or ( \6915_b1 , \6913_b1 , w_22068 );
or ( \6915_b0 , \6913_b0 , \6914_b0 );
not ( \6914_b0 , w_22069 );
and ( w_22069 , w_22068 , \6914_b1 );
or ( \6916_b1 , \6839_b1 , w_22071 );
not ( w_22071 , w_22072 );
and ( \6916_b0 , \6839_b0 , w_22073 );
and ( w_22072 ,  , w_22073 );
buf ( w_22071 , \4754_b1 );
not ( w_22071 , w_22074 );
not (  , w_22075 );
and ( w_22074 , w_22075 , \4754_b0 );
or ( \6917_b1 , \6915_b1 , w_22077 );
not ( w_22077 , w_22078 );
and ( \6917_b0 , \6915_b0 , w_22079 );
and ( w_22078 ,  , w_22079 );
buf ( w_22077 , \6916_b1 );
not ( w_22077 , w_22080 );
not (  , w_22081 );
and ( w_22080 , w_22081 , \6916_b0 );
buf ( \6918_b1 , \6401_b1 );
not ( \6918_b1 , w_22082 );
not ( \6918_b0 , w_22083 );
and ( w_22082 , w_22083 , \6401_b0 );
buf ( \6919_b1 , \6492_b1 );
not ( \6919_b1 , w_22084 );
not ( \6919_b0 , w_22085 );
and ( w_22084 , w_22085 , \6492_b0 );
or ( \6920_b1 , \6918_b1 , w_22086 );
or ( \6920_b0 , \6918_b0 , \6919_b0 );
not ( \6919_b0 , w_22087 );
and ( w_22087 , w_22086 , \6919_b1 );
or ( \6921_b1 , \6696_b1 , w_22089 );
not ( w_22089 , w_22090 );
and ( \6921_b0 , \6696_b0 , w_22091 );
and ( w_22090 ,  , w_22091 );
buf ( w_22089 , \5266_b1 );
not ( w_22089 , w_22092 );
not (  , w_22093 );
and ( w_22092 , w_22093 , \5266_b0 );
or ( \6922_b1 , \6920_b1 , w_22095 );
not ( w_22095 , w_22096 );
and ( \6922_b0 , \6920_b0 , w_22097 );
and ( w_22096 ,  , w_22097 );
buf ( w_22095 , \6921_b1 );
not ( w_22095 , w_22098 );
not (  , w_22099 );
and ( w_22098 , w_22099 , \6921_b0 );
or ( \6923_b1 , \6917_b1 , w_22100 );
or ( \6923_b0 , \6917_b0 , \6922_b0 );
not ( \6922_b0 , w_22101 );
and ( w_22101 , w_22100 , \6922_b1 );
or ( \6924_b1 , \6912_b1 , w_22103 );
not ( w_22103 , w_22104 );
and ( \6924_b0 , \6912_b0 , w_22105 );
and ( w_22104 ,  , w_22105 );
buf ( w_22103 , \6923_b1 );
not ( w_22103 , w_22106 );
not (  , w_22107 );
and ( w_22106 , w_22107 , \6923_b0 );
or ( \6925_b1 , \6917_b1 , w_22109 );
not ( w_22109 , w_22110 );
and ( \6925_b0 , \6917_b0 , w_22111 );
and ( w_22110 ,  , w_22111 );
buf ( w_22109 , \6922_b1 );
not ( w_22109 , w_22112 );
not (  , w_22113 );
and ( w_22112 , w_22113 , \6922_b0 );
or ( \6926_b1 , \6924_b1 , \6925_b1 );
not ( \6925_b1 , w_22114 );
and ( \6926_b0 , \6924_b0 , w_22115 );
and ( w_22114 , w_22115 , \6925_b0 );
or ( \6927_b1 , \6910_b1 , \6926_b1 );
xor ( \6927_b0 , \6910_b0 , w_22116 );
not ( w_22116 , w_22117 );
and ( w_22117 , \6926_b1 , \6926_b0 );
or ( \6928_b1 , \6844_b1 , \6853_b1 );
xor ( \6928_b0 , \6844_b0 , w_22118 );
not ( w_22118 , w_22119 );
and ( w_22119 , \6853_b1 , \6853_b0 );
or ( \6929_b1 , \6928_b1 , w_22120 );
xor ( \6929_b0 , \6928_b0 , w_22122 );
not ( w_22122 , w_22123 );
and ( w_22123 , w_22120 , w_22121 );
buf ( w_22120 , \6874_b1 );
not ( w_22120 , w_22124 );
not ( w_22121 , w_22125 );
and ( w_22124 , w_22125 , \6874_b0 );
or ( \6930_b1 , \6927_b1 , \6929_b1 );
xor ( \6930_b0 , \6927_b0 , w_22126 );
not ( w_22126 , w_22127 );
and ( w_22127 , \6929_b1 , \6929_b0 );
or ( \6931_b1 , \6858_b1 , \6864_b1 );
xor ( \6931_b0 , \6858_b0 , w_22128 );
not ( w_22128 , w_22129 );
and ( w_22129 , \6864_b1 , \6864_b0 );
or ( \6932_b1 , \6931_b1 , w_22130 );
xor ( \6932_b0 , \6931_b0 , w_22132 );
not ( w_22132 , w_22133 );
and ( w_22133 , w_22130 , w_22131 );
buf ( w_22130 , \6872_b1 );
not ( w_22130 , w_22134 );
not ( w_22131 , w_22135 );
and ( w_22134 , w_22135 , \6872_b0 );
or ( \6933_b1 , \6403_b1 , \6412_b1 );
xor ( \6933_b0 , \6403_b0 , w_22136 );
not ( w_22136 , w_22137 );
and ( w_22137 , \6412_b1 , \6412_b0 );
or ( \6934_b1 , \6933_b1 , \6426_b1 );
not ( \6426_b1 , w_22138 );
and ( \6934_b0 , \6933_b0 , w_22139 );
and ( w_22138 , w_22139 , \6426_b0 );
or ( \6935_b1 , \6403_b1 , \6412_b1 );
not ( \6412_b1 , w_22140 );
and ( \6935_b0 , \6403_b0 , w_22141 );
and ( w_22140 , w_22141 , \6412_b0 );
or ( \6936_b1 , \6934_b1 , w_22142 );
or ( \6936_b0 , \6934_b0 , \6935_b0 );
not ( \6935_b0 , w_22143 );
and ( w_22143 , w_22142 , \6935_b1 );
or ( \6937_b1 , \6932_b1 , \6936_b1 );
xor ( \6937_b0 , \6932_b0 , w_22144 );
not ( w_22144 , w_22145 );
and ( w_22145 , \6936_b1 , \6936_b0 );
or ( \6938_b1 , \6922_b1 , \6917_b1 );
xor ( \6938_b0 , \6922_b0 , w_22146 );
not ( w_22146 , w_22147 );
and ( w_22147 , \6917_b1 , \6917_b0 );
or ( \6939_b1 , \6938_b1 , w_22148 );
xor ( \6939_b0 , \6938_b0 , w_22150 );
not ( w_22150 , w_22151 );
and ( w_22151 , w_22148 , w_22149 );
buf ( w_22148 , \6911_b1 );
not ( w_22148 , w_22152 );
not ( w_22149 , w_22153 );
and ( w_22152 , w_22153 , \6911_b0 );
or ( \6940_b1 , \6937_b1 , \6939_b1 );
not ( \6939_b1 , w_22154 );
and ( \6940_b0 , \6937_b0 , w_22155 );
and ( w_22154 , w_22155 , \6939_b0 );
or ( \6941_b1 , \6932_b1 , \6936_b1 );
not ( \6936_b1 , w_22156 );
and ( \6941_b0 , \6932_b0 , w_22157 );
and ( w_22156 , w_22157 , \6936_b0 );
or ( \6942_b1 , \6940_b1 , w_22158 );
or ( \6942_b0 , \6940_b0 , \6941_b0 );
not ( \6941_b0 , w_22159 );
and ( w_22159 , w_22158 , \6941_b1 );
buf ( \6943_b1 , \6942_b1 );
not ( \6943_b1 , w_22160 );
not ( \6943_b0 , w_22161 );
and ( w_22160 , w_22161 , \6942_b0 );
or ( \6944_b1 , \6930_b1 , w_22163 );
not ( w_22163 , w_22164 );
and ( \6944_b0 , \6930_b0 , w_22165 );
and ( w_22164 ,  , w_22165 );
buf ( w_22163 , \6943_b1 );
not ( w_22163 , w_22166 );
not (  , w_22167 );
and ( w_22166 , w_22167 , \6943_b0 );
or ( \6945_b1 , \6932_b1 , \6936_b1 );
xor ( \6945_b0 , \6932_b0 , w_22168 );
not ( w_22168 , w_22169 );
and ( w_22169 , \6936_b1 , \6936_b0 );
or ( \6946_b1 , \6945_b1 , \6939_b1 );
xor ( \6946_b0 , \6945_b0 , w_22170 );
not ( w_22170 , w_22171 );
and ( w_22171 , \6939_b1 , \6939_b0 );
buf ( \6947_b1 , \6946_b1 );
not ( \6947_b1 , w_22172 );
not ( \6947_b0 , w_22173 );
and ( w_22172 , w_22173 , \6946_b0 );
or ( \6948_b1 , \6388_b1 , \6392_b1 );
xor ( \6948_b0 , \6388_b0 , w_22174 );
not ( w_22174 , w_22175 );
and ( w_22175 , \6392_b1 , \6392_b0 );
or ( \6949_b1 , \6948_b1 , \6427_b1 );
not ( \6427_b1 , w_22176 );
and ( \6949_b0 , \6948_b0 , w_22177 );
and ( w_22176 , w_22177 , \6427_b0 );
or ( \6950_b1 , \6388_b1 , \6392_b1 );
not ( \6392_b1 , w_22178 );
and ( \6950_b0 , \6388_b0 , w_22179 );
and ( w_22178 , w_22179 , \6392_b0 );
or ( \6951_b1 , \6949_b1 , w_22180 );
or ( \6951_b0 , \6949_b0 , \6950_b0 );
not ( \6950_b0 , w_22181 );
and ( w_22181 , w_22180 , \6950_b1 );
buf ( \6952_b1 , \6951_b1 );
not ( \6952_b1 , w_22182 );
not ( \6952_b0 , w_22183 );
and ( w_22182 , w_22183 , \6951_b0 );
or ( \6953_b1 , \6947_b1 , w_22185 );
not ( w_22185 , w_22186 );
and ( \6953_b0 , \6947_b0 , w_22187 );
and ( w_22186 ,  , w_22187 );
buf ( w_22185 , \6952_b1 );
not ( w_22185 , w_22188 );
not (  , w_22189 );
and ( w_22188 , w_22189 , \6952_b0 );
or ( \6954_b1 , \6944_b1 , \6953_b1 );
not ( \6953_b1 , w_22190 );
and ( \6954_b0 , \6944_b0 , w_22191 );
and ( w_22190 , w_22191 , \6953_b0 );
or ( \6955_b1 , \6876_b1 , \6888_b1 );
not ( \6888_b1 , w_22192 );
and ( \6955_b0 , \6876_b0 , w_22193 );
and ( w_22192 , w_22193 , \6888_b0 );
buf ( \6956_b1 , \6876_b1 );
not ( \6956_b1 , w_22194 );
not ( \6956_b0 , w_22195 );
and ( w_22194 , w_22195 , \6876_b0 );
or ( \6957_b1 , \6956_b1 , \6889_b1 );
not ( \6889_b1 , w_22196 );
and ( \6957_b0 , \6956_b0 , w_22197 );
and ( w_22196 , w_22197 , \6889_b0 );
or ( \6958_b1 , \6955_b1 , w_22199 );
not ( w_22199 , w_22200 );
and ( \6958_b0 , \6955_b0 , w_22201 );
and ( w_22200 ,  , w_22201 );
buf ( w_22199 , \6957_b1 );
not ( w_22199 , w_22202 );
not (  , w_22203 );
and ( w_22202 , w_22203 , \6957_b0 );
or ( \6959_b1 , \6958_b1 , w_22204 );
xor ( \6959_b0 , \6958_b0 , w_22206 );
not ( w_22206 , w_22207 );
and ( w_22207 , w_22204 , w_22205 );
buf ( w_22204 , \6901_b1 );
not ( w_22204 , w_22208 );
not ( w_22205 , w_22209 );
and ( w_22208 , w_22209 , \6901_b0 );
or ( \6960_b1 , \6910_b1 , \6926_b1 );
xor ( \6960_b0 , \6910_b0 , w_22210 );
not ( w_22210 , w_22211 );
and ( w_22211 , \6926_b1 , \6926_b0 );
or ( \6961_b1 , \6960_b1 , \6929_b1 );
not ( \6929_b1 , w_22212 );
and ( \6961_b0 , \6960_b0 , w_22213 );
and ( w_22212 , w_22213 , \6929_b0 );
or ( \6962_b1 , \6910_b1 , \6926_b1 );
not ( \6926_b1 , w_22214 );
and ( \6962_b0 , \6910_b0 , w_22215 );
and ( w_22214 , w_22215 , \6926_b0 );
or ( \6963_b1 , \6961_b1 , w_22216 );
or ( \6963_b0 , \6961_b0 , \6962_b0 );
not ( \6962_b0 , w_22217 );
and ( w_22217 , w_22216 , \6962_b1 );
or ( \6964_b1 , \6959_b1 , w_22219 );
not ( w_22219 , w_22220 );
and ( \6964_b0 , \6959_b0 , w_22221 );
and ( w_22220 ,  , w_22221 );
buf ( w_22219 , \6963_b1 );
not ( w_22219 , w_22222 );
not (  , w_22223 );
and ( w_22222 , w_22223 , \6963_b0 );
buf ( \6966_b1 , \6965_b1 );
not ( \6966_b1 , w_22224 );
not ( \6966_b0 , w_22225 );
and ( w_22224 , w_22225 , \6965_b0 );
buf ( \6967_b1 , \6966_b1 );
not ( \6967_b1 , w_22226 );
not ( \6967_b0 , w_22227 );
and ( w_22226 , w_22227 , \6966_b0 );
or ( \6968_b1 , \6602_b1 , w_22228 );
or ( \6968_b0 , \6602_b0 , \6967_b0 );
not ( \6967_b0 , w_22229 );
and ( w_22229 , w_22228 , \6967_b1 );
buf ( \6969_b1 , \6834_b1 );
not ( \6969_b1 , w_22230 );
not ( \6969_b0 , w_22231 );
and ( w_22230 , w_22231 , \6834_b0 );
or ( \6970_b1 , \6969_b1 , w_22233 );
not ( w_22233 , w_22234 );
and ( \6970_b0 , \6969_b0 , w_22235 );
and ( w_22234 ,  , w_22235 );
buf ( w_22233 , \6906_b1 );
not ( w_22233 , w_22236 );
not (  , w_22237 );
and ( w_22236 , w_22237 , \6906_b0 );
buf ( \6971_b1 , \6959_b1 );
not ( \6971_b1 , w_22238 );
not ( \6971_b0 , w_22239 );
and ( w_22238 , w_22239 , \6959_b0 );
buf ( \6972_b1 , \6963_b1 );
not ( \6972_b1 , w_22240 );
not ( \6972_b0 , w_22241 );
and ( w_22240 , w_22241 , \6963_b0 );
or ( \6973_b1 , \6971_b1 , w_22243 );
not ( w_22243 , w_22244 );
and ( \6973_b0 , \6971_b0 , w_22245 );
and ( w_22244 ,  , w_22245 );
buf ( w_22243 , \6972_b1 );
not ( w_22243 , w_22246 );
not (  , w_22247 );
and ( w_22246 , w_22247 , \6972_b0 );
or ( \6974_b1 , \6970_b1 , w_22249 );
not ( w_22249 , w_22250 );
and ( \6974_b0 , \6970_b0 , w_22251 );
and ( w_22250 ,  , w_22251 );
buf ( w_22249 , \6973_b1 );
not ( w_22249 , w_22252 );
not (  , w_22253 );
and ( w_22252 , w_22253 , \6973_b0 );
buf ( \6975_b1 , \6930_b1 );
not ( \6975_b1 , w_22254 );
not ( \6975_b0 , w_22255 );
and ( w_22254 , w_22255 , \6930_b0 );
or ( \6976_b1 , \6975_b1 , w_22257 );
not ( w_22257 , w_22258 );
and ( \6976_b0 , \6975_b0 , w_22259 );
and ( w_22258 ,  , w_22259 );
buf ( w_22257 , \6942_b1 );
not ( w_22257 , w_22260 );
not (  , w_22261 );
and ( w_22260 , w_22261 , \6942_b0 );
or ( \6977_b1 , \6946_b1 , w_22263 );
not ( w_22263 , w_22264 );
and ( \6977_b0 , \6946_b0 , w_22265 );
and ( w_22264 ,  , w_22265 );
buf ( w_22263 , \6951_b1 );
not ( w_22263 , w_22266 );
not (  , w_22267 );
and ( w_22266 , w_22267 , \6951_b0 );
or ( \6978_b1 , \6976_b1 , w_22269 );
not ( w_22269 , w_22270 );
and ( \6978_b0 , \6976_b0 , w_22271 );
and ( w_22270 ,  , w_22271 );
buf ( w_22269 , \6977_b1 );
not ( w_22269 , w_22272 );
not (  , w_22273 );
and ( w_22272 , w_22273 , \6977_b0 );
or ( \6980_b1 , \6974_b1 , w_22274 );
or ( \6980_b0 , \6974_b0 , \6979_b0 );
not ( \6979_b0 , w_22275 );
and ( w_22275 , w_22274 , \6979_b1 );
buf ( \6981_b1 , \6908_b1 );
buf ( \6981_b0 , \6908_b0 );
or ( \6982_b1 , \6980_b1 , w_22277 );
not ( w_22277 , w_22278 );
and ( \6982_b0 , \6980_b0 , w_22279 );
and ( w_22278 ,  , w_22279 );
buf ( w_22277 , \6981_b1 );
not ( w_22277 , w_22280 );
not (  , w_22281 );
and ( w_22280 , w_22281 , \6981_b0 );
or ( \6983_b1 , \6968_b1 , w_22283 );
not ( w_22283 , w_22284 );
and ( \6983_b0 , \6968_b0 , w_22285 );
and ( w_22284 ,  , w_22285 );
buf ( w_22283 , \6982_b1 );
not ( w_22283 , w_22286 );
not (  , w_22287 );
and ( w_22286 , w_22287 , \6982_b0 );
or ( \6984_b1 , \6062_b1 , \6088_b1 );
xor ( \6984_b0 , \6062_b0 , w_22288 );
not ( w_22288 , w_22289 );
and ( w_22289 , \6088_b1 , \6088_b0 );
or ( \6985_b1 , \6984_b1 , w_22290 );
xor ( \6985_b0 , \6984_b0 , w_22292 );
not ( w_22292 , w_22293 );
and ( w_22293 , w_22290 , w_22291 );
buf ( w_22290 , \6074_b1 );
not ( w_22290 , w_22294 );
not ( w_22291 , w_22295 );
and ( w_22294 , w_22295 , \6074_b0 );
buf ( \6986_b1 , \6622_b1 );
not ( \6986_b1 , w_22296 );
not ( \6986_b0 , w_22297 );
and ( w_22296 , w_22297 , \6622_b0 );
buf ( \6987_b1 , \6612_b1 );
not ( \6987_b1 , w_22298 );
not ( \6987_b0 , w_22299 );
and ( w_22298 , w_22299 , \6612_b0 );
or ( \6988_b1 , \6986_b1 , w_22300 );
or ( \6988_b0 , \6986_b0 , \6987_b0 );
not ( \6987_b0 , w_22301 );
and ( w_22301 , w_22300 , \6987_b1 );
or ( \6989_b1 , \6612_b1 , w_22302 );
or ( \6989_b0 , \6612_b0 , \6622_b0 );
not ( \6622_b0 , w_22303 );
and ( w_22303 , w_22302 , \6622_b1 );
or ( \6990_b1 , \6989_b1 , w_22305 );
not ( w_22305 , w_22306 );
and ( \6990_b0 , \6989_b0 , w_22307 );
and ( w_22306 ,  , w_22307 );
buf ( w_22305 , \6633_b1 );
not ( w_22305 , w_22308 );
not (  , w_22309 );
and ( w_22308 , w_22309 , \6633_b0 );
or ( \6991_b1 , \6988_b1 , w_22311 );
not ( w_22311 , w_22312 );
and ( \6991_b0 , \6988_b0 , w_22313 );
and ( w_22312 ,  , w_22313 );
buf ( w_22311 , \6990_b1 );
not ( w_22311 , w_22314 );
not (  , w_22315 );
and ( w_22314 , w_22315 , \6990_b0 );
buf ( \6992_b1 , \6796_b1 );
not ( \6992_b1 , w_22316 );
not ( \6992_b0 , w_22317 );
and ( w_22316 , w_22317 , \6796_b0 );
buf ( \6993_b1 , \4611_b1 );
not ( \6993_b1 , w_22318 );
not ( \6993_b0 , w_22319 );
and ( w_22318 , w_22319 , \4611_b0 );
or ( \6994_b1 , \6992_b1 , w_22320 );
or ( \6994_b0 , \6992_b0 , \6993_b0 );
not ( \6993_b0 , w_22321 );
and ( w_22321 , w_22320 , \6993_b1 );
or ( \6995_b1 , \4754_b1 , w_22323 );
not ( w_22323 , w_22324 );
and ( \6995_b0 , \4754_b0 , w_22325 );
and ( w_22324 ,  , w_22325 );
buf ( w_22323 , \6108_b1 );
not ( w_22323 , w_22326 );
not (  , w_22327 );
and ( w_22326 , w_22327 , \6108_b0 );
or ( \6996_b1 , \6994_b1 , w_22329 );
not ( w_22329 , w_22330 );
and ( \6996_b0 , \6994_b0 , w_22331 );
and ( w_22330 ,  , w_22331 );
buf ( w_22329 , \6995_b1 );
not ( w_22329 , w_22332 );
not (  , w_22333 );
and ( w_22332 , w_22333 , \6995_b0 );
buf ( \6997_b1 , \6996_b1 );
not ( \6997_b1 , w_22334 );
not ( \6997_b0 , w_22335 );
and ( w_22334 , w_22335 , \6996_b0 );
buf ( \6998_b1 , \6812_b1 );
not ( \6998_b1 , w_22336 );
not ( \6998_b0 , w_22337 );
and ( w_22336 , w_22337 , \6812_b0 );
or ( \6999_b1 , \6998_b1 , w_22339 );
not ( w_22339 , w_22340 );
and ( \6999_b0 , \6998_b0 , w_22341 );
and ( w_22340 ,  , w_22341 );
buf ( w_22339 , \6807_b1 );
not ( w_22339 , w_22342 );
not (  , w_22343 );
and ( w_22342 , w_22343 , \6807_b0 );
or ( \7000_b1 , \6997_b1 , w_22345 );
not ( w_22345 , w_22346 );
and ( \7000_b0 , \6997_b0 , w_22347 );
and ( w_22346 ,  , w_22347 );
buf ( w_22345 , \6999_b1 );
not ( w_22345 , w_22348 );
not (  , w_22349 );
and ( w_22348 , w_22349 , \6999_b0 );
or ( \7001_b1 , \6991_b1 , \7000_b1 );
not ( \7000_b1 , w_22350 );
and ( \7001_b0 , \6991_b0 , w_22351 );
and ( w_22350 , w_22351 , \7000_b0 );
or ( \7002_b1 , \6997_b1 , w_22353 );
not ( w_22353 , w_22354 );
and ( \7002_b0 , \6997_b0 , w_22355 );
and ( w_22354 ,  , w_22355 );
buf ( w_22353 , \6999_b1 );
not ( w_22353 , w_22356 );
not (  , w_22357 );
and ( w_22356 , w_22357 , \6999_b0 );
or ( \7003_b1 , \7001_b1 , w_22359 );
not ( w_22359 , w_22360 );
and ( \7003_b0 , \7001_b0 , w_22361 );
and ( w_22360 ,  , w_22361 );
buf ( w_22359 , \7002_b1 );
not ( w_22359 , w_22362 );
not (  , w_22363 );
and ( w_22362 , w_22363 , \7002_b0 );
or ( \7004_b1 , \6985_b1 , \7003_b1 );
xor ( \7004_b0 , \6985_b0 , w_22364 );
not ( w_22364 , w_22365 );
and ( w_22365 , \7003_b1 , \7003_b0 );
buf ( \7005_b1 , \6113_b1 );
not ( \7005_b1 , w_22366 );
not ( \7005_b0 , w_22367 );
and ( w_22366 , w_22367 , \6113_b0 );
or ( \7006_b1 , \6124_b1 , \7005_b1 );
xor ( \7006_b0 , \6124_b0 , w_22368 );
not ( w_22368 , w_22369 );
and ( w_22369 , \7005_b1 , \7005_b0 );
or ( \7007_b1 , \7006_b1 , \6103_b1 );
not ( \6103_b1 , w_22370 );
and ( \7007_b0 , \7006_b0 , w_22371 );
and ( w_22370 , w_22371 , \6103_b0 );
buf ( \7008_b1 , \7006_b1 );
not ( \7008_b1 , w_22372 );
not ( \7008_b0 , w_22373 );
and ( w_22372 , w_22373 , \7006_b0 );
buf ( \7009_b1 , \6103_b1 );
not ( \7009_b1 , w_22374 );
not ( \7009_b0 , w_22375 );
and ( w_22374 , w_22375 , \6103_b0 );
or ( \7010_b1 , \7008_b1 , \7009_b1 );
not ( \7009_b1 , w_22376 );
and ( \7010_b0 , \7008_b0 , w_22377 );
and ( w_22376 , w_22377 , \7009_b0 );
or ( \7011_b1 , \7007_b1 , w_22379 );
not ( w_22379 , w_22380 );
and ( \7011_b0 , \7007_b0 , w_22381 );
and ( w_22380 ,  , w_22381 );
buf ( w_22379 , \7010_b1 );
not ( w_22379 , w_22382 );
not (  , w_22383 );
and ( w_22382 , w_22383 , \7010_b0 );
or ( \7012_b1 , \7004_b1 , \7011_b1 );
xor ( \7012_b0 , \7004_b0 , w_22384 );
not ( w_22384 , w_22385 );
and ( w_22385 , \7011_b1 , \7011_b0 );
buf ( \7013_b1 , \7012_b1 );
not ( \7013_b1 , w_22386 );
not ( \7013_b0 , w_22387 );
and ( w_22386 , w_22387 , \7012_b0 );
buf ( \7014_b1 , \7013_b1 );
not ( \7014_b1 , w_22388 );
not ( \7014_b0 , w_22389 );
and ( w_22388 , w_22389 , \7013_b0 );
or ( \7015_b1 , \6162_b1 , \6192_b1 );
xor ( \7015_b0 , \6162_b0 , w_22390 );
not ( w_22390 , w_22391 );
and ( w_22391 , \6192_b1 , \6192_b0 );
or ( \7016_b1 , \7015_b1 , w_22392 );
xor ( \7016_b0 , \7015_b0 , w_22394 );
not ( w_22394 , w_22395 );
and ( w_22395 , w_22392 , w_22393 );
buf ( w_22392 , \6232_b1 );
not ( w_22392 , w_22396 );
not ( w_22393 , w_22397 );
and ( w_22396 , w_22397 , \6232_b0 );
buf ( \7017_b1 , \7016_b1 );
not ( \7017_b1 , w_22398 );
not ( \7017_b0 , w_22399 );
and ( w_22398 , w_22399 , \7016_b0 );
or ( \7018_b1 , \7014_b1 , w_22400 );
or ( \7018_b0 , \7014_b0 , \7017_b0 );
not ( \7017_b0 , w_22401 );
and ( w_22401 , w_22400 , \7017_b1 );
buf ( \7019_b1 , \7016_b1 );
not ( \7019_b1 , w_22402 );
not ( \7019_b0 , w_22403 );
and ( w_22402 , w_22403 , \7016_b0 );
buf ( \7020_b1 , \7019_b1 );
not ( \7020_b1 , w_22404 );
not ( \7020_b0 , w_22405 );
and ( w_22404 , w_22405 , \7019_b0 );
buf ( \7021_b1 , \7012_b1 );
not ( \7021_b1 , w_22406 );
not ( \7021_b0 , w_22407 );
and ( w_22406 , w_22407 , \7012_b0 );
or ( \7022_b1 , \7020_b1 , w_22408 );
or ( \7022_b0 , \7020_b0 , \7021_b0 );
not ( \7021_b0 , w_22409 );
and ( w_22409 , w_22408 , \7021_b1 );
or ( \7023_b1 , \6173_b1 , \6175_b1 );
xor ( \7023_b0 , \6173_b0 , w_22410 );
not ( w_22410 , w_22411 );
and ( w_22411 , \6175_b1 , \6175_b0 );
or ( \7024_b1 , \7023_b1 , \6186_b1 );
xor ( \7024_b0 , \7023_b0 , w_22412 );
not ( w_22412 , w_22413 );
and ( w_22413 , \6186_b1 , \6186_b0 );
buf ( \7025_b1 , \7024_b1 );
not ( \7025_b1 , w_22414 );
not ( \7025_b0 , w_22415 );
and ( w_22414 , w_22415 , \7024_b0 );
or ( \7026_b1 , \6798_b1 , \6816_b1 );
xor ( \7026_b0 , \6798_b0 , w_22416 );
not ( w_22416 , w_22417 );
and ( w_22417 , \6816_b1 , \6816_b0 );
or ( \7027_b1 , \7026_b1 , \6827_b1 );
not ( \6827_b1 , w_22418 );
and ( \7027_b0 , \7026_b0 , w_22419 );
and ( w_22418 , w_22419 , \6827_b0 );
or ( \7028_b1 , \6798_b1 , \6816_b1 );
not ( \6816_b1 , w_22420 );
and ( \7028_b0 , \6798_b0 , w_22421 );
and ( w_22420 , w_22421 , \6816_b0 );
or ( \7029_b1 , \7027_b1 , w_22422 );
or ( \7029_b0 , \7027_b0 , \7028_b0 );
not ( \7028_b0 , w_22423 );
and ( w_22423 , w_22422 , \7028_b1 );
buf ( \7030_b1 , \7029_b1 );
not ( \7030_b1 , w_22424 );
not ( \7030_b0 , w_22425 );
and ( w_22424 , w_22425 , \7029_b0 );
buf ( \7031_b1 , \7030_b1 );
not ( \7031_b1 , w_22426 );
not ( \7031_b0 , w_22427 );
and ( w_22426 , w_22427 , \7030_b0 );
or ( \7032_b1 , \7025_b1 , w_22428 );
or ( \7032_b0 , \7025_b0 , \7031_b0 );
not ( \7031_b0 , w_22429 );
and ( w_22429 , w_22428 , \7031_b1 );
buf ( \7033_b1 , \6229_b1 );
not ( \7033_b1 , w_22430 );
not ( \7033_b0 , w_22431 );
and ( w_22430 , w_22431 , \6229_b0 );
buf ( \7034_b1 , \6205_b1 );
not ( \7034_b1 , w_22432 );
not ( \7034_b0 , w_22433 );
and ( w_22432 , w_22433 , \6205_b0 );
or ( \7035_b1 , \7033_b1 , w_22434 );
or ( \7035_b0 , \7033_b0 , \7034_b0 );
not ( \7034_b0 , w_22435 );
and ( w_22435 , w_22434 , \7034_b1 );
or ( \7036_b1 , \6205_b1 , w_22436 );
or ( \7036_b0 , \6205_b0 , \6229_b0 );
not ( \6229_b0 , w_22437 );
and ( w_22437 , w_22436 , \6229_b1 );
or ( \7037_b1 , \7035_b1 , w_22439 );
not ( w_22439 , w_22440 );
and ( \7037_b0 , \7035_b0 , w_22441 );
and ( w_22440 ,  , w_22441 );
buf ( w_22439 , \7036_b1 );
not ( w_22439 , w_22442 );
not (  , w_22443 );
and ( w_22442 , w_22443 , \7036_b0 );
or ( \7038_b1 , \7037_b1 , \6216_b1 );
not ( \6216_b1 , w_22444 );
and ( \7038_b0 , \7037_b0 , w_22445 );
and ( w_22444 , w_22445 , \6216_b0 );
buf ( \7039_b1 , \7037_b1 );
not ( \7039_b1 , w_22446 );
not ( \7039_b0 , w_22447 );
and ( w_22446 , w_22447 , \7037_b0 );
or ( \7040_b1 , \7039_b1 , \6217_b1 );
not ( \6217_b1 , w_22448 );
and ( \7040_b0 , \7039_b0 , w_22449 );
and ( w_22448 , w_22449 , \6217_b0 );
or ( \7041_b1 , \7038_b1 , w_22451 );
not ( w_22451 , w_22452 );
and ( \7041_b0 , \7038_b0 , w_22453 );
and ( w_22452 ,  , w_22453 );
buf ( w_22451 , \7040_b1 );
not ( w_22451 , w_22454 );
not (  , w_22455 );
and ( w_22454 , w_22455 , \7040_b0 );
or ( \7042_b1 , \7032_b1 , w_22457 );
not ( w_22457 , w_22458 );
and ( \7042_b0 , \7032_b0 , w_22459 );
and ( w_22458 ,  , w_22459 );
buf ( w_22457 , \7041_b1 );
not ( w_22457 , w_22460 );
not (  , w_22461 );
and ( w_22460 , w_22461 , \7041_b0 );
buf ( \7043_b1 , \7024_b1 );
not ( \7043_b1 , w_22462 );
not ( \7043_b0 , w_22463 );
and ( w_22462 , w_22463 , \7024_b0 );
or ( \7044_b1 , \7043_b1 , w_22465 );
not ( w_22465 , w_22466 );
and ( \7044_b0 , \7043_b0 , w_22467 );
and ( w_22466 ,  , w_22467 );
buf ( w_22465 , \7029_b1 );
not ( w_22465 , w_22468 );
not (  , w_22469 );
and ( w_22468 , w_22469 , \7029_b0 );
or ( \7045_b1 , \7042_b1 , w_22471 );
not ( w_22471 , w_22472 );
and ( \7045_b0 , \7042_b0 , w_22473 );
and ( w_22472 ,  , w_22473 );
buf ( w_22471 , \7044_b1 );
not ( w_22471 , w_22474 );
not (  , w_22475 );
and ( w_22474 , w_22475 , \7044_b0 );
or ( \7046_b1 , \7022_b1 , w_22477 );
not ( w_22477 , w_22478 );
and ( \7046_b0 , \7022_b0 , w_22479 );
and ( w_22478 ,  , w_22479 );
buf ( w_22477 , \7045_b1 );
not ( w_22477 , w_22480 );
not (  , w_22481 );
and ( w_22480 , w_22481 , \7045_b0 );
or ( \7047_b1 , \7018_b1 , w_22483 );
not ( w_22483 , w_22484 );
and ( \7047_b0 , \7018_b0 , w_22485 );
and ( w_22484 ,  , w_22485 );
buf ( w_22483 , \7046_b1 );
not ( w_22483 , w_22486 );
not (  , w_22487 );
and ( w_22486 , w_22487 , \7046_b0 );
buf ( \7048_b1 , \7047_b1 );
not ( \7048_b1 , w_22488 );
not ( \7048_b0 , w_22489 );
and ( w_22488 , w_22489 , \7047_b0 );
or ( \7049_b1 , \6090_b1 , \6051_b1 );
xor ( \7049_b0 , \6090_b0 , w_22490 );
not ( w_22490 , w_22491 );
and ( w_22491 , \6051_b1 , \6051_b0 );
buf ( \7050_b1 , \6127_b1 );
not ( \7050_b1 , w_22492 );
not ( \7050_b0 , w_22493 );
and ( w_22492 , w_22493 , \6127_b0 );
or ( \7051_b1 , \7049_b1 , \7050_b1 );
not ( \7050_b1 , w_22494 );
and ( \7051_b0 , \7049_b0 , w_22495 );
and ( w_22494 , w_22495 , \7050_b0 );
buf ( \7052_b1 , \7049_b1 );
not ( \7052_b1 , w_22496 );
not ( \7052_b0 , w_22497 );
and ( w_22496 , w_22497 , \7049_b0 );
or ( \7053_b1 , \7052_b1 , \6127_b1 );
not ( \6127_b1 , w_22498 );
and ( \7053_b0 , \7052_b0 , w_22499 );
and ( w_22498 , w_22499 , \6127_b0 );
or ( \7054_b1 , \7051_b1 , w_22501 );
not ( w_22501 , w_22502 );
and ( \7054_b0 , \7051_b0 , w_22503 );
and ( w_22502 ,  , w_22503 );
buf ( w_22501 , \7053_b1 );
not ( w_22501 , w_22504 );
not (  , w_22505 );
and ( w_22504 , w_22505 , \7053_b0 );
or ( \7055_b1 , \6985_b1 , \7003_b1 );
xor ( \7055_b0 , \6985_b0 , w_22506 );
not ( w_22506 , w_22507 );
and ( w_22507 , \7003_b1 , \7003_b0 );
or ( \7056_b1 , \7055_b1 , \7011_b1 );
not ( \7011_b1 , w_22508 );
and ( \7056_b0 , \7055_b0 , w_22509 );
and ( w_22508 , w_22509 , \7011_b0 );
or ( \7057_b1 , \6985_b1 , \7003_b1 );
not ( \7003_b1 , w_22510 );
and ( \7057_b0 , \6985_b0 , w_22511 );
and ( w_22510 , w_22511 , \7003_b0 );
or ( \7058_b1 , \7056_b1 , w_22512 );
or ( \7058_b0 , \7056_b0 , \7057_b0 );
not ( \7057_b0 , w_22513 );
and ( w_22513 , w_22512 , \7057_b1 );
or ( \7059_b1 , \7054_b1 , \7058_b1 );
xor ( \7059_b0 , \7054_b0 , w_22514 );
not ( w_22514 , w_22515 );
and ( w_22515 , \7058_b1 , \7058_b0 );
or ( \7060_b1 , \6251_b1 , \6261_b1 );
not ( \6261_b1 , w_22516 );
and ( \7060_b0 , \6251_b0 , w_22517 );
and ( w_22516 , w_22517 , \6261_b0 );
buf ( \7061_b1 , \6251_b1 );
not ( \7061_b1 , w_22518 );
not ( \7061_b0 , w_22519 );
and ( w_22518 , w_22519 , \6251_b0 );
buf ( \7062_b1 , \6261_b1 );
not ( \7062_b1 , w_22520 );
not ( \7062_b0 , w_22521 );
and ( w_22520 , w_22521 , \6261_b0 );
or ( \7063_b1 , \7061_b1 , \7062_b1 );
not ( \7062_b1 , w_22522 );
and ( \7063_b0 , \7061_b0 , w_22523 );
and ( w_22522 , w_22523 , \7062_b0 );
or ( \7064_b1 , \7060_b1 , w_22525 );
not ( w_22525 , w_22526 );
and ( \7064_b0 , \7060_b0 , w_22527 );
and ( w_22526 ,  , w_22527 );
buf ( w_22525 , \7063_b1 );
not ( w_22525 , w_22528 );
not (  , w_22529 );
and ( w_22528 , w_22529 , \7063_b0 );
or ( \7065_b1 , \6236_b1 , \7064_b1 );
xor ( \7065_b0 , \6236_b0 , w_22530 );
not ( w_22530 , w_22531 );
and ( w_22531 , \7064_b1 , \7064_b0 );
or ( \7066_b1 , \7059_b1 , \7065_b1 );
xor ( \7066_b0 , \7059_b0 , w_22532 );
not ( w_22532 , w_22533 );
and ( w_22533 , \7065_b1 , \7065_b0 );
buf ( \7067_b1 , \7066_b1 );
buf ( \7067_b0 , \7066_b0 );
or ( \7068_b1 , \7048_b1 , w_22535 );
not ( w_22535 , w_22536 );
and ( \7068_b0 , \7048_b0 , w_22537 );
and ( w_22536 ,  , w_22537 );
buf ( w_22535 , \7067_b1 );
not ( w_22535 , w_22538 );
not (  , w_22539 );
and ( w_22538 , w_22539 , \7067_b0 );
or ( \7069_b1 , \6161_b1 , \6267_b1 );
xor ( \7069_b0 , \6161_b0 , w_22540 );
not ( w_22540 , w_22541 );
and ( w_22541 , \6267_b1 , \6267_b0 );
or ( \7070_b1 , \7069_b1 , \6270_b1 );
xor ( \7070_b0 , \7069_b0 , w_22542 );
not ( w_22542 , w_22543 );
and ( w_22543 , \6270_b1 , \6270_b0 );
buf ( \7071_b1 , \7070_b1 );
not ( \7071_b1 , w_22544 );
not ( \7071_b0 , w_22545 );
and ( w_22544 , w_22545 , \7070_b0 );
or ( \7072_b1 , \7054_b1 , \7058_b1 );
xor ( \7072_b0 , \7054_b0 , w_22546 );
not ( w_22546 , w_22547 );
and ( w_22547 , \7058_b1 , \7058_b0 );
or ( \7073_b1 , \7072_b1 , \7065_b1 );
not ( \7065_b1 , w_22548 );
and ( \7073_b0 , \7072_b0 , w_22549 );
and ( w_22548 , w_22549 , \7065_b0 );
or ( \7074_b1 , \7054_b1 , \7058_b1 );
not ( \7058_b1 , w_22550 );
and ( \7074_b0 , \7054_b0 , w_22551 );
and ( w_22550 , w_22551 , \7058_b0 );
or ( \7075_b1 , \7073_b1 , w_22552 );
or ( \7075_b0 , \7073_b0 , \7074_b0 );
not ( \7074_b0 , w_22553 );
and ( w_22553 , w_22552 , \7074_b1 );
or ( \7076_b1 , \7071_b1 , w_22555 );
not ( w_22555 , w_22556 );
and ( \7076_b0 , \7071_b0 , w_22557 );
and ( w_22556 ,  , w_22557 );
buf ( w_22555 , \7075_b1 );
not ( w_22555 , w_22558 );
not (  , w_22559 );
and ( w_22558 , w_22559 , \7075_b0 );
or ( \7077_b1 , \7016_b1 , \7045_b1 );
xor ( \7077_b0 , \7016_b0 , w_22560 );
not ( w_22560 , w_22561 );
and ( w_22561 , \7045_b1 , \7045_b0 );
or ( \7078_b1 , \7077_b1 , \7012_b1 );
not ( \7012_b1 , w_22562 );
and ( \7078_b0 , \7077_b0 , w_22563 );
and ( w_22562 , w_22563 , \7012_b0 );
buf ( \7079_b1 , \7077_b1 );
not ( \7079_b1 , w_22564 );
not ( \7079_b0 , w_22565 );
and ( w_22564 , w_22565 , \7077_b0 );
or ( \7080_b1 , \7079_b1 , \7013_b1 );
not ( \7013_b1 , w_22566 );
and ( \7080_b0 , \7079_b0 , w_22567 );
and ( w_22566 , w_22567 , \7013_b0 );
or ( \7081_b1 , \7078_b1 , w_22569 );
not ( w_22569 , w_22570 );
and ( \7081_b0 , \7078_b0 , w_22571 );
and ( w_22570 ,  , w_22571 );
buf ( w_22569 , \7080_b1 );
not ( w_22569 , w_22572 );
not (  , w_22573 );
and ( w_22572 , w_22573 , \7080_b0 );
buf ( \7082_b1 , \6999_b1 );
not ( \7082_b1 , w_22574 );
not ( \7082_b0 , w_22575 );
and ( w_22574 , w_22575 , \6999_b0 );
buf ( \7083_b1 , \7082_b1 );
not ( \7083_b1 , w_22576 );
not ( \7083_b0 , w_22577 );
and ( w_22576 , w_22577 , \7082_b0 );
buf ( \7084_b1 , \6997_b1 );
not ( \7084_b1 , w_22578 );
not ( \7084_b0 , w_22579 );
and ( w_22578 , w_22579 , \6997_b0 );
or ( \7085_b1 , \7083_b1 , w_22580 );
or ( \7085_b0 , \7083_b0 , \7084_b0 );
not ( \7084_b0 , w_22581 );
and ( w_22581 , w_22580 , \7084_b1 );
or ( \7086_b1 , \6997_b1 , w_22582 );
or ( \7086_b0 , \6997_b0 , \7082_b0 );
not ( \7082_b0 , w_22583 );
and ( w_22583 , w_22582 , \7082_b1 );
or ( \7087_b1 , \7085_b1 , w_22585 );
not ( w_22585 , w_22586 );
and ( \7087_b0 , \7085_b0 , w_22587 );
and ( w_22586 ,  , w_22587 );
buf ( w_22585 , \7086_b1 );
not ( w_22585 , w_22588 );
not (  , w_22589 );
and ( w_22588 , w_22589 , \7086_b0 );
or ( \7088_b1 , \6991_b1 , \7087_b1 );
xor ( \7088_b0 , \6991_b0 , w_22590 );
not ( w_22590 , w_22591 );
and ( w_22591 , \7087_b1 , \7087_b0 );
buf ( \7089_b1 , \7088_b1 );
buf ( \7089_b0 , \7088_b0 );
buf ( \7090_b1 , \7089_b1 );
not ( \7090_b1 , w_22592 );
not ( \7090_b0 , w_22593 );
and ( w_22592 , w_22593 , \7089_b0 );
or ( \7091_b1 , \7024_b1 , \7029_b1 );
xor ( \7091_b0 , \7024_b0 , w_22594 );
not ( w_22594 , w_22595 );
and ( w_22595 , \7029_b1 , \7029_b0 );
or ( \7092_b1 , \7091_b1 , w_22596 );
xor ( \7092_b0 , \7091_b0 , w_22598 );
not ( w_22598 , w_22599 );
and ( w_22599 , w_22596 , w_22597 );
buf ( w_22596 , \7041_b1 );
not ( w_22596 , w_22600 );
not ( w_22597 , w_22601 );
and ( w_22600 , w_22601 , \7041_b0 );
buf ( \7093_b1 , \7092_b1 );
not ( \7093_b1 , w_22602 );
not ( \7093_b0 , w_22603 );
and ( w_22602 , w_22603 , \7092_b0 );
or ( \7094_b1 , \7090_b1 , w_22605 );
not ( w_22605 , w_22606 );
and ( \7094_b0 , \7090_b0 , w_22607 );
and ( w_22606 ,  , w_22607 );
buf ( w_22605 , \7093_b1 );
not ( w_22605 , w_22608 );
not (  , w_22609 );
and ( w_22608 , w_22609 , \7093_b0 );
or ( \7095_b1 , \6756_b1 , \6787_b1 );
xor ( \7095_b0 , \6756_b0 , w_22610 );
not ( w_22610 , w_22611 );
and ( w_22611 , \6787_b1 , \6787_b0 );
or ( \7096_b1 , \7095_b1 , \6828_b1 );
not ( \6828_b1 , w_22612 );
and ( \7096_b0 , \7095_b0 , w_22613 );
and ( w_22612 , w_22613 , \6828_b0 );
or ( \7097_b1 , \6756_b1 , \6787_b1 );
not ( \6787_b1 , w_22614 );
and ( \7097_b0 , \6756_b0 , w_22615 );
and ( w_22614 , w_22615 , \6787_b0 );
or ( \7098_b1 , \7096_b1 , w_22616 );
or ( \7098_b0 , \7096_b0 , \7097_b0 );
not ( \7097_b0 , w_22617 );
and ( w_22617 , w_22616 , \7097_b1 );
buf ( \7099_b1 , \7098_b1 );
buf ( \7099_b0 , \7098_b0 );
or ( \7100_b1 , \7094_b1 , \7099_b1 );
not ( \7099_b1 , w_22618 );
and ( \7100_b0 , \7094_b0 , w_22619 );
and ( w_22618 , w_22619 , \7099_b0 );
or ( \7101_b1 , \7092_b1 , \7089_b1 );
not ( \7089_b1 , w_22620 );
and ( \7101_b0 , \7092_b0 , w_22621 );
and ( w_22620 , w_22621 , \7089_b0 );
or ( \7102_b1 , \7100_b1 , w_22623 );
not ( w_22623 , w_22624 );
and ( \7102_b0 , \7100_b0 , w_22625 );
and ( w_22624 ,  , w_22625 );
buf ( w_22623 , \7101_b1 );
not ( w_22623 , w_22626 );
not (  , w_22627 );
and ( w_22626 , w_22627 , \7101_b0 );
or ( \7103_b1 , \7081_b1 , w_22629 );
not ( w_22629 , w_22630 );
and ( \7103_b0 , \7081_b0 , w_22631 );
and ( w_22630 ,  , w_22631 );
buf ( w_22629 , \7102_b1 );
not ( w_22629 , w_22632 );
not (  , w_22633 );
and ( w_22632 , w_22633 , \7102_b0 );
buf ( \7104_b1 , \6829_b1 );
not ( \7104_b1 , w_22634 );
not ( \7104_b0 , w_22635 );
and ( w_22634 , w_22635 , \6829_b0 );
buf ( \7105_b1 , \6634_b1 );
not ( \7105_b1 , w_22636 );
not ( \7105_b0 , w_22637 );
and ( w_22636 , w_22637 , \6634_b0 );
or ( \7106_b1 , \7105_b1 , w_22639 );
not ( w_22639 , w_22640 );
and ( \7106_b0 , \7105_b0 , w_22641 );
and ( w_22640 ,  , w_22641 );
buf ( w_22639 , \6745_b1 );
not ( w_22639 , w_22642 );
not (  , w_22643 );
and ( w_22642 , w_22643 , \6745_b0 );
buf ( \7107_b1 , \7106_b1 );
not ( \7107_b1 , w_22644 );
not ( \7107_b0 , w_22645 );
and ( w_22644 , w_22645 , \7106_b0 );
or ( \7108_b1 , \7104_b1 , w_22646 );
or ( \7108_b0 , \7104_b0 , \7107_b0 );
not ( \7107_b0 , w_22647 );
and ( w_22647 , w_22646 , \7107_b1 );
or ( \7109_b1 , \6744_b1 , w_22649 );
not ( w_22649 , w_22650 );
and ( \7109_b0 , \6744_b0 , w_22651 );
and ( w_22650 ,  , w_22651 );
buf ( w_22649 , \6634_b1 );
not ( w_22649 , w_22652 );
not (  , w_22653 );
and ( w_22652 , w_22653 , \6634_b0 );
or ( \7110_b1 , \7108_b1 , w_22655 );
not ( w_22655 , w_22656 );
and ( \7110_b0 , \7108_b0 , w_22657 );
and ( w_22656 ,  , w_22657 );
buf ( w_22655 , \7109_b1 );
not ( w_22655 , w_22658 );
not (  , w_22659 );
and ( w_22658 , w_22659 , \7109_b0 );
buf ( \7111_b1 , \7110_b1 );
not ( \7111_b1 , w_22660 );
not ( \7111_b0 , w_22661 );
and ( w_22660 , w_22661 , \7110_b0 );
or ( \7112_b1 , \7088_b1 , \7098_b1 );
xor ( \7112_b0 , \7088_b0 , w_22662 );
not ( w_22662 , w_22663 );
and ( w_22663 , \7098_b1 , \7098_b0 );
or ( \7113_b1 , \7112_b1 , w_22664 );
xor ( \7113_b0 , \7112_b0 , w_22666 );
not ( w_22666 , w_22667 );
and ( w_22667 , w_22664 , w_22665 );
buf ( w_22664 , \7092_b1 );
not ( w_22664 , w_22668 );
not ( w_22665 , w_22669 );
and ( w_22668 , w_22669 , \7092_b0 );
or ( \7114_b1 , \7111_b1 , w_22671 );
not ( w_22671 , w_22672 );
and ( \7114_b0 , \7111_b0 , w_22673 );
and ( w_22672 ,  , w_22673 );
buf ( w_22671 , \7113_b1 );
not ( w_22671 , w_22674 );
not (  , w_22675 );
and ( w_22674 , w_22675 , \7113_b0 );
or ( \7115_b1 , \7103_b1 , \7114_b1 );
not ( \7114_b1 , w_22676 );
and ( \7115_b0 , \7103_b0 , w_22677 );
and ( w_22676 , w_22677 , \7114_b0 );
or ( \7117_b1 , \6983_b1 , w_22679 );
not ( w_22679 , w_22680 );
and ( \7117_b0 , \6983_b0 , w_22681 );
and ( w_22680 ,  , w_22681 );
buf ( w_22679 , \7116_b1 );
not ( w_22679 , w_22682 );
not (  , w_22683 );
and ( w_22682 , w_22683 , \7116_b0 );
buf ( \7118_b1 , \7075_b1 );
not ( \7118_b1 , w_22684 );
not ( \7118_b0 , w_22685 );
and ( w_22684 , w_22685 , \7075_b0 );
or ( \7119_b1 , \7118_b1 , w_22687 );
not ( w_22687 , w_22688 );
and ( \7119_b0 , \7118_b0 , w_22689 );
and ( w_22688 ,  , w_22689 );
buf ( w_22687 , \7070_b1 );
not ( w_22687 , w_22690 );
not (  , w_22691 );
and ( w_22690 , w_22691 , \7070_b0 );
buf ( \7120_b1 , \7119_b1 );
not ( \7120_b1 , w_22692 );
not ( \7120_b0 , w_22693 );
and ( w_22692 , w_22693 , \7119_b0 );
buf ( \7121_b1 , \7103_b1 );
not ( \7121_b1 , w_22694 );
not ( \7121_b0 , w_22695 );
and ( w_22694 , w_22695 , \7103_b0 );
buf ( \7122_b1 , \7113_b1 );
not ( \7122_b1 , w_22696 );
not ( \7122_b0 , w_22697 );
and ( w_22696 , w_22697 , \7113_b0 );
or ( \7123_b1 , \7122_b1 , w_22699 );
not ( w_22699 , w_22700 );
and ( \7123_b0 , \7122_b0 , w_22701 );
and ( w_22700 ,  , w_22701 );
buf ( w_22699 , \7110_b1 );
not ( w_22699 , w_22702 );
not (  , w_22703 );
and ( w_22702 , w_22703 , \7110_b0 );
or ( \7124_b1 , \7121_b1 , w_22705 );
not ( w_22705 , w_22706 );
and ( \7124_b0 , \7121_b0 , w_22707 );
and ( w_22706 ,  , w_22707 );
buf ( w_22705 , \7123_b1 );
not ( w_22705 , w_22708 );
not (  , w_22709 );
and ( w_22708 , w_22709 , \7123_b0 );
buf ( \7125_b1 , \7081_b1 );
not ( \7125_b1 , w_22710 );
not ( \7125_b0 , w_22711 );
and ( w_22710 , w_22711 , \7081_b0 );
buf ( \7126_b1 , \7102_b1 );
not ( \7126_b1 , w_22712 );
not ( \7126_b0 , w_22713 );
and ( w_22712 , w_22713 , \7102_b0 );
or ( \7127_b1 , \7125_b1 , w_22715 );
not ( w_22715 , w_22716 );
and ( \7127_b0 , \7125_b0 , w_22717 );
and ( w_22716 ,  , w_22717 );
buf ( w_22715 , \7126_b1 );
not ( w_22715 , w_22718 );
not (  , w_22719 );
and ( w_22718 , w_22719 , \7126_b0 );
buf ( \7128_b1 , \7066_b1 );
not ( \7128_b1 , w_22720 );
not ( \7128_b0 , w_22721 );
and ( w_22720 , w_22721 , \7066_b0 );
or ( \7129_b1 , \7128_b1 , w_22723 );
not ( w_22723 , w_22724 );
and ( \7129_b0 , \7128_b0 , w_22725 );
and ( w_22724 ,  , w_22725 );
buf ( w_22723 , \7047_b1 );
not ( w_22723 , w_22726 );
not (  , w_22727 );
and ( w_22726 , w_22727 , \7047_b0 );
or ( \7130_b1 , \7127_b1 , w_22729 );
not ( w_22729 , w_22730 );
and ( \7130_b0 , \7127_b0 , w_22731 );
and ( w_22730 ,  , w_22731 );
buf ( w_22729 , \7129_b1 );
not ( w_22729 , w_22732 );
not (  , w_22733 );
and ( w_22732 , w_22733 , \7129_b0 );
or ( \7131_b1 , \7124_b1 , w_22734 );
or ( \7131_b0 , \7124_b0 , \7130_b0 );
not ( \7130_b0 , w_22735 );
and ( w_22735 , w_22734 , \7130_b1 );
or ( \7132_b1 , \7131_b1 , w_22737 );
not ( w_22737 , w_22738 );
and ( \7132_b0 , \7131_b0 , w_22739 );
and ( w_22738 ,  , w_22739 );
buf ( w_22737 , \7068_b1 );
not ( w_22737 , w_22740 );
not (  , w_22741 );
and ( w_22740 , w_22741 , \7068_b0 );
buf ( \7133_b1 , \7132_b1 );
not ( \7133_b1 , w_22742 );
not ( \7133_b0 , w_22743 );
and ( w_22742 , w_22743 , \7132_b0 );
or ( \7134_b1 , \7120_b1 , w_22744 );
or ( \7134_b0 , \7120_b0 , \7133_b0 );
not ( \7133_b0 , w_22745 );
and ( w_22745 , w_22744 , \7133_b1 );
buf ( \7135_b1 , \7076_b1 );
buf ( \7135_b0 , \7076_b0 );
or ( \7136_b1 , \7134_b1 , w_22747 );
not ( w_22747 , w_22748 );
and ( \7136_b0 , \7134_b0 , w_22749 );
and ( w_22748 ,  , w_22749 );
buf ( w_22747 , \7135_b1 );
not ( w_22747 , w_22750 );
not (  , w_22751 );
and ( w_22750 , w_22751 , \7135_b0 );
or ( \7137_b1 , \7117_b1 , w_22753 );
not ( w_22753 , w_22754 );
and ( \7137_b0 , \7117_b0 , w_22755 );
and ( w_22754 ,  , w_22755 );
buf ( w_22753 , \7136_b1 );
not ( w_22753 , w_22756 );
not (  , w_22757 );
and ( w_22756 , w_22757 , \7136_b0 );
buf ( \7139_b1 , \6288_b1 );
not ( \7139_b1 , w_22758 );
not ( \7139_b0 , w_22759 );
and ( w_22758 , w_22759 , \6288_b0 );
or ( \7140_b1 , \6044_b1 , w_22761 );
not ( w_22761 , w_22762 );
and ( \7140_b0 , \6044_b0 , w_22763 );
and ( w_22762 ,  , w_22763 );
buf ( w_22761 , \6149_b1 );
not ( w_22761 , w_22764 );
not (  , w_22765 );
and ( w_22764 , w_22765 , \6149_b0 );
buf ( \7141_b1 , \7140_b1 );
not ( \7141_b1 , w_22766 );
not ( \7141_b0 , w_22767 );
and ( w_22766 , w_22767 , \7140_b0 );
or ( \7142_b1 , \6276_b1 , w_22769 );
not ( w_22769 , w_22770 );
and ( \7142_b0 , \6276_b0 , w_22771 );
and ( w_22770 ,  , w_22771 );
buf ( w_22769 , \6273_b1 );
not ( w_22769 , w_22772 );
not (  , w_22773 );
and ( w_22772 , w_22773 , \6273_b0 );
buf ( \7143_b1 , \7142_b1 );
not ( \7143_b1 , w_22774 );
not ( \7143_b0 , w_22775 );
and ( w_22774 , w_22775 , \7142_b0 );
or ( \7144_b1 , \7141_b1 , w_22776 );
or ( \7144_b0 , \7141_b0 , \7143_b0 );
not ( \7143_b0 , w_22777 );
and ( w_22777 , w_22776 , \7143_b1 );
or ( \7145_b1 , \7144_b1 , w_22779 );
not ( w_22779 , w_22780 );
and ( \7145_b0 , \7144_b0 , w_22781 );
and ( w_22780 ,  , w_22781 );
buf ( w_22779 , \6151_b1 );
not ( w_22779 , w_22782 );
not (  , w_22783 );
and ( w_22782 , w_22783 , \6151_b0 );
or ( \7146_b1 , \7145_b1 , w_22784 );
or ( \7146_b0 , \7145_b0 , \6033_b0 );
not ( \6033_b0 , w_22785 );
and ( w_22785 , w_22784 , \6033_b1 );
or ( \7147_b1 , \5849_b1 , w_22787 );
not ( w_22787 , w_22788 );
and ( \7147_b0 , \5849_b0 , w_22789 );
and ( w_22788 ,  , w_22789 );
buf ( w_22787 , \6032_b1 );
not ( w_22787 , w_22790 );
not (  , w_22791 );
and ( w_22790 , w_22791 , \6032_b0 );
or ( \7148_b1 , \7146_b1 , w_22793 );
not ( w_22793 , w_22794 );
and ( \7148_b0 , \7146_b0 , w_22795 );
and ( w_22794 ,  , w_22795 );
buf ( w_22793 , \7147_b1 );
not ( w_22793 , w_22796 );
not (  , w_22797 );
and ( w_22796 , w_22797 , \7147_b0 );
buf ( \7149_b1 , \7148_b1 );
not ( \7149_b1 , w_22798 );
not ( \7149_b0 , w_22799 );
and ( w_22798 , w_22799 , \7148_b0 );
or ( \7150_b1 , \7139_b1 , w_22800 );
or ( \7150_b0 , \7139_b0 , \7149_b0 );
not ( \7149_b0 , w_22801 );
and ( w_22801 , w_22800 , \7149_b1 );
buf ( \7151_b1 , \6287_b1 );
not ( \7151_b1 , w_22802 );
not ( \7151_b0 , w_22803 );
and ( w_22802 , w_22803 , \6287_b0 );
buf ( \7152_b1 , \6281_b1 );
not ( \7152_b1 , w_22804 );
not ( \7152_b0 , w_22805 );
and ( w_22804 , w_22805 , \6281_b0 );
or ( \7153_b1 , \7151_b1 , w_22807 );
not ( w_22807 , w_22808 );
and ( \7153_b0 , \7151_b0 , w_22809 );
and ( w_22808 ,  , w_22809 );
buf ( w_22807 , \7152_b1 );
not ( w_22807 , w_22810 );
not (  , w_22811 );
and ( w_22810 , w_22811 , \7152_b0 );
or ( \7154_b1 , \7150_b1 , w_22813 );
not ( w_22813 , w_22814 );
and ( \7154_b0 , \7150_b0 , w_22815 );
and ( w_22814 ,  , w_22815 );
buf ( w_22813 , \7153_b1 );
not ( w_22813 , w_22816 );
not (  , w_22817 );
and ( w_22816 , w_22817 , \7153_b0 );
or ( \7155_b1 , \7154_b1 , w_22819 );
not ( w_22819 , w_22820 );
and ( \7155_b0 , \7154_b0 , w_22821 );
and ( w_22820 ,  , w_22821 );
buf ( w_22819 , \5707_b1 );
not ( w_22819 , w_22822 );
not (  , w_22823 );
and ( w_22822 , w_22823 , \5707_b0 );
buf ( \7156_b1 , \5649_b1 );
buf ( \7156_b0 , \5649_b0 );
buf ( \7157_b1 , \5651_b1 );
not ( \7157_b1 , w_22824 );
not ( \7157_b0 , w_22825 );
and ( w_22824 , w_22825 , \5651_b0 );
buf ( \7158_b1 , \5705_b1 );
not ( \7158_b1 , w_22826 );
not ( \7158_b0 , w_22827 );
and ( w_22826 , w_22827 , \5705_b0 );
or ( \7159_b1 , \7157_b1 , w_22829 );
not ( w_22829 , w_22830 );
and ( \7159_b0 , \7157_b0 , w_22831 );
and ( w_22830 ,  , w_22831 );
buf ( w_22829 , \7158_b1 );
not ( w_22829 , w_22832 );
not (  , w_22833 );
and ( w_22832 , w_22833 , \7158_b0 );
or ( \7160_b1 , \5354_b1 , w_22834 );
or ( \7160_b0 , \5354_b0 , \5617_b0 );
not ( \5617_b0 , w_22835 );
and ( w_22835 , w_22834 , \5617_b1 );
or ( \7161_b1 , \7159_b1 , w_22837 );
not ( w_22837 , w_22838 );
and ( \7161_b0 , \7159_b0 , w_22839 );
and ( w_22838 ,  , w_22839 );
buf ( w_22837 , \7160_b1 );
not ( w_22837 , w_22840 );
not (  , w_22841 );
and ( w_22840 , w_22841 , \7160_b0 );
or ( \7162_b1 , \7156_b1 , \7161_b1 );
not ( \7161_b1 , w_22842 );
and ( \7162_b0 , \7156_b0 , w_22843 );
and ( w_22842 , w_22843 , \7161_b0 );
buf ( \7163_b1 , \5648_b1 );
buf ( \7163_b0 , \5648_b0 );
buf ( \7164_b1 , \7163_b1 );
not ( \7164_b1 , w_22844 );
not ( \7164_b0 , w_22845 );
and ( w_22844 , w_22845 , \7163_b0 );
or ( \7165_b1 , \5640_b1 , w_22846 );
or ( \7165_b0 , \5640_b0 , \5622_b0 );
not ( \5622_b0 , w_22847 );
and ( w_22847 , w_22846 , \5622_b1 );
or ( \7166_b1 , \7164_b1 , w_22848 );
or ( \7166_b0 , \7164_b0 , \7165_b0 );
not ( \7165_b0 , w_22849 );
and ( w_22849 , w_22848 , \7165_b1 );
or ( \7167_b1 , \5647_b1 , w_22850 );
or ( \7167_b0 , \5647_b0 , \5645_b0 );
not ( \5645_b0 , w_22851 );
and ( w_22851 , w_22850 , \5645_b1 );
or ( \7168_b1 , \7166_b1 , w_22853 );
not ( w_22853 , w_22854 );
and ( \7168_b0 , \7166_b0 , w_22855 );
and ( w_22854 ,  , w_22855 );
buf ( w_22853 , \7167_b1 );
not ( w_22853 , w_22856 );
not (  , w_22857 );
and ( w_22856 , w_22857 , \7167_b0 );
or ( \7169_b1 , \7162_b1 , w_22859 );
not ( w_22859 , w_22860 );
and ( \7169_b0 , \7162_b0 , w_22861 );
and ( w_22860 ,  , w_22861 );
buf ( w_22859 , \7168_b1 );
not ( w_22859 , w_22862 );
not (  , w_22863 );
and ( w_22862 , w_22863 , \7168_b0 );
buf ( \7171_b1 , \7170_b1 );
not ( \7171_b1 , w_22864 );
not ( \7171_b0 , w_22865 );
and ( w_22864 , w_22865 , \7170_b0 );
or ( \7172_b1 , \5071_b1 , w_22866 );
or ( \7172_b0 , \5071_b0 , \7171_b0 );
not ( \7171_b0 , w_22867 );
and ( w_22867 , w_22866 , \7171_b1 );
buf ( \7173_b1 , \5069_b1 );
not ( \7173_b1 , w_22868 );
not ( \7173_b0 , w_22869 );
and ( w_22868 , w_22869 , \5069_b0 );
buf ( \7174_b1 , \7173_b1 );
not ( \7174_b1 , w_22870 );
not ( \7174_b0 , w_22871 );
and ( w_22870 , w_22871 , \7173_b0 );
buf ( \7175_b1 , \5045_b1 );
not ( \7175_b1 , w_22872 );
not ( \7175_b0 , w_22873 );
and ( w_22872 , w_22873 , \5045_b0 );
buf ( \7176_b1 , \4370_b1 );
not ( \7176_b1 , w_22874 );
not ( \7176_b0 , w_22875 );
and ( w_22874 , w_22875 , \4370_b0 );
or ( \7177_b1 , \4828_b1 , w_22877 );
not ( w_22877 , w_22878 );
and ( \7177_b0 , \4828_b0 , w_22879 );
and ( w_22878 ,  , w_22879 );
buf ( w_22877 , \5003_b1 );
not ( w_22877 , w_22880 );
not (  , w_22881 );
and ( w_22880 , w_22881 , \5003_b0 );
or ( \7178_b1 , \4825_b1 , w_22883 );
not ( w_22883 , w_22884 );
and ( \7178_b0 , \4825_b0 , w_22885 );
and ( w_22884 ,  , w_22885 );
buf ( w_22883 , \7177_b1 );
not ( w_22883 , w_22886 );
not (  , w_22887 );
and ( w_22886 , w_22887 , \7177_b0 );
or ( \7179_b1 , \4822_b1 , \4824_b1 );
not ( \4824_b1 , w_22888 );
and ( \7179_b0 , \4822_b0 , w_22889 );
and ( w_22888 , w_22889 , \4824_b0 );
or ( \7180_b1 , \7178_b1 , w_22891 );
not ( w_22891 , w_22892 );
and ( \7180_b0 , \7178_b0 , w_22893 );
and ( w_22892 ,  , w_22893 );
buf ( w_22891 , \7179_b1 );
not ( w_22891 , w_22894 );
not (  , w_22895 );
and ( w_22894 , w_22895 , \7179_b0 );
or ( \7181_b1 , \5010_b1 , w_22897 );
not ( w_22897 , w_22898 );
and ( \7181_b0 , \5010_b0 , w_22899 );
and ( w_22898 ,  , w_22899 );
buf ( w_22897 , \5012_b1 );
not ( w_22897 , w_22900 );
not (  , w_22901 );
and ( w_22900 , w_22901 , \5012_b0 );
buf ( \7182_b1 , \7181_b1 );
not ( \7182_b1 , w_22902 );
not ( \7182_b0 , w_22903 );
and ( w_22902 , w_22903 , \7181_b0 );
or ( \7183_b1 , \4488_b1 , \4586_b1 );
not ( \4586_b1 , w_22904 );
and ( \7183_b0 , \4488_b0 , w_22905 );
and ( w_22904 , w_22905 , \4586_b0 );
or ( \7184_b1 , \7182_b1 , w_22907 );
not ( w_22907 , w_22908 );
and ( \7184_b0 , \7182_b0 , w_22909 );
and ( w_22908 ,  , w_22909 );
buf ( w_22907 , \7183_b1 );
not ( w_22907 , w_22910 );
not (  , w_22911 );
and ( w_22910 , w_22911 , \7183_b0 );
or ( \7185_b1 , \7180_b1 , \7184_b1 );
not ( \7184_b1 , w_22912 );
and ( \7185_b0 , \7180_b0 , w_22913 );
and ( w_22912 , w_22913 , \7184_b0 );
buf ( \7186_b1 , \4588_b1 );
not ( \7186_b1 , w_22914 );
not ( \7186_b0 , w_22915 );
and ( w_22914 , w_22915 , \4588_b0 );
buf ( \7187_b1 , \5013_b1 );
not ( \7187_b1 , w_22916 );
not ( \7187_b0 , w_22917 );
and ( w_22916 , w_22917 , \5013_b0 );
or ( \7188_b1 , \7186_b1 , w_22918 );
or ( \7188_b0 , \7186_b0 , \7187_b0 );
not ( \7187_b0 , w_22919 );
and ( w_22919 , w_22918 , \7187_b1 );
or ( \7189_b1 , \7188_b1 , w_22921 );
not ( w_22921 , w_22922 );
and ( \7189_b0 , \7188_b0 , w_22923 );
and ( w_22922 ,  , w_22923 );
buf ( w_22921 , \7181_b1 );
not ( w_22921 , w_22924 );
not (  , w_22925 );
and ( w_22924 , w_22925 , \7181_b0 );
buf ( \7190_b1 , \7189_b1 );
not ( \7190_b1 , w_22926 );
not ( \7190_b0 , w_22927 );
and ( w_22926 , w_22927 , \7189_b0 );
or ( \7191_b1 , \7185_b1 , w_22929 );
not ( w_22929 , w_22930 );
and ( \7191_b0 , \7185_b0 , w_22931 );
and ( w_22930 ,  , w_22931 );
buf ( w_22929 , \7190_b1 );
not ( w_22929 , w_22932 );
not (  , w_22933 );
and ( w_22932 , w_22933 , \7190_b0 );
buf ( \7192_b1 , \7191_b1 );
not ( \7192_b1 , w_22934 );
not ( \7192_b0 , w_22935 );
and ( w_22934 , w_22935 , \7191_b0 );
or ( \7193_b1 , \7176_b1 , w_22936 );
or ( \7193_b0 , \7176_b0 , \7192_b0 );
not ( \7192_b0 , w_22937 );
and ( w_22937 , w_22936 , \7192_b1 );
or ( \7194_b1 , \4369_b1 , w_22938 );
or ( \7194_b0 , \4369_b0 , \4293_b0 );
not ( \4293_b0 , w_22939 );
and ( w_22939 , w_22938 , \4293_b1 );
or ( \7195_b1 , \7193_b1 , w_22941 );
not ( w_22941 , w_22942 );
and ( \7195_b0 , \7193_b0 , w_22943 );
and ( w_22942 ,  , w_22943 );
buf ( w_22941 , \7194_b1 );
not ( w_22941 , w_22944 );
not (  , w_22945 );
and ( w_22944 , w_22945 , \7194_b0 );
buf ( \7196_b1 , \7195_b1 );
not ( \7196_b1 , w_22946 );
not ( \7196_b0 , w_22947 );
and ( w_22946 , w_22947 , \7195_b0 );
or ( \7197_b1 , \7175_b1 , w_22948 );
or ( \7197_b0 , \7175_b0 , \7196_b0 );
not ( \7196_b0 , w_22949 );
and ( w_22949 , w_22948 , \7196_b1 );
or ( \7198_b1 , \5019_b1 , w_22951 );
not ( w_22951 , w_22952 );
and ( \7198_b0 , \5019_b0 , w_22953 );
and ( w_22952 ,  , w_22953 );
buf ( w_22951 , \5044_b1 );
not ( w_22951 , w_22954 );
not (  , w_22955 );
and ( w_22954 , w_22955 , \5044_b0 );
or ( \7199_b1 , \7197_b1 , w_22957 );
not ( w_22957 , w_22958 );
and ( \7199_b0 , \7197_b0 , w_22959 );
and ( w_22958 ,  , w_22959 );
buf ( w_22957 , \7198_b1 );
not ( w_22957 , w_22960 );
not (  , w_22961 );
and ( w_22960 , w_22961 , \7198_b0 );
buf ( \7200_b1 , \7199_b1 );
not ( \7200_b1 , w_22962 );
not ( \7200_b0 , w_22963 );
and ( w_22962 , w_22963 , \7199_b0 );
or ( \7201_b1 , \7174_b1 , w_22964 );
or ( \7201_b0 , \7174_b0 , \7200_b0 );
not ( \7200_b0 , w_22965 );
and ( w_22965 , w_22964 , \7200_b1 );
or ( \7202_b1 , \5050_b1 , w_22967 );
not ( w_22967 , w_22968 );
and ( \7202_b0 , \5050_b0 , w_22969 );
and ( w_22968 ,  , w_22969 );
buf ( w_22967 , \5068_b1 );
not ( w_22967 , w_22970 );
not (  , w_22971 );
and ( w_22970 , w_22971 , \5068_b0 );
or ( \7203_b1 , \7201_b1 , w_22973 );
not ( w_22973 , w_22974 );
and ( \7203_b0 , \7201_b0 , w_22975 );
and ( w_22974 ,  , w_22975 );
buf ( w_22973 , \7202_b1 );
not ( w_22973 , w_22976 );
not (  , w_22977 );
and ( w_22976 , w_22977 , \7202_b0 );
buf ( \7204_b1 , \7203_b1 );
not ( \7204_b1 , w_22978 );
not ( \7204_b0 , w_22979 );
and ( w_22978 , w_22979 , \7203_b0 );
or ( \7205_b1 , \7172_b1 , w_22981 );
not ( w_22981 , w_22982 );
and ( \7205_b0 , \7172_b0 , w_22983 );
and ( w_22982 ,  , w_22983 );
buf ( w_22981 , \7204_b1 );
not ( w_22981 , w_22984 );
not (  , w_22985 );
and ( w_22984 , w_22985 , \7204_b0 );
buf ( \7206_b1 , \5064_b1 );
not ( \7206_b1 , w_22986 );
not ( \7206_b0 , w_22987 );
and ( w_22986 , w_22987 , \5064_b0 );
or ( \7207_b1 , \4195_b1 , \7206_b1 );
not ( \7206_b1 , w_22988 );
and ( \7207_b0 , \4195_b0 , w_22989 );
and ( w_22988 , w_22989 , \7206_b0 );
or ( \7208_b1 , \4200_b1 , \4253_b1 );
not ( \4253_b1 , w_22990 );
and ( \7208_b0 , \4200_b0 , w_22991 );
and ( w_22990 , w_22991 , \4253_b0 );
or ( \7209_b1 , \7207_b1 , w_22993 );
not ( w_22993 , w_22994 );
and ( \7209_b0 , \7207_b0 , w_22995 );
and ( w_22994 ,  , w_22995 );
buf ( w_22993 , \7208_b1 );
not ( w_22993 , w_22996 );
not (  , w_22997 );
and ( w_22996 , w_22997 , \7208_b0 );
buf ( \7210_b1 , \7209_b1 );
not ( \7210_b1 , w_22998 );
not ( \7210_b0 , w_22999 );
and ( w_22998 , w_22999 , \7209_b0 );
or ( \7211_b1 , \4253_b1 , w_23001 );
not ( w_23001 , w_23002 );
and ( \7211_b0 , \4253_b0 , w_23003 );
and ( w_23002 ,  , w_23003 );
buf ( w_23001 , \3997_b1 );
not ( w_23001 , w_23004 );
not (  , w_23005 );
and ( w_23004 , w_23005 , \3997_b0 );
buf ( \7212_b1 , \7211_b1 );
not ( \7212_b1 , w_23006 );
not ( \7212_b0 , w_23007 );
and ( w_23006 , w_23007 , \7211_b0 );
or ( \7213_b1 , \7210_b1 , \7212_b1 );
not ( \7212_b1 , w_23008 );
and ( \7213_b0 , \7210_b0 , w_23009 );
and ( w_23008 , w_23009 , \7212_b0 );
or ( \7214_b1 , \7209_b1 , \7211_b1 );
not ( \7211_b1 , w_23010 );
and ( \7214_b0 , \7209_b0 , w_23011 );
and ( w_23010 , w_23011 , \7211_b0 );
or ( \7215_b1 , \7213_b1 , w_23013 );
not ( w_23013 , w_23014 );
and ( \7215_b0 , \7213_b0 , w_23015 );
and ( w_23014 ,  , w_23015 );
buf ( w_23013 , \7214_b1 );
not ( w_23013 , w_23016 );
not (  , w_23017 );
and ( w_23016 , w_23017 , \7214_b0 );
buf ( \7216_b1 , \7215_b1 );
not ( \7216_b1 , w_23018 );
not ( \7216_b0 , w_23019 );
and ( w_23018 , w_23019 , \7215_b0 );
or ( \7217_b1 , \5057_b1 , \5059_b1 );
xor ( \7217_b0 , \5057_b0 , w_23020 );
not ( w_23020 , w_23021 );
and ( w_23021 , \5059_b1 , \5059_b0 );
or ( \7218_b1 , \7217_b1 , \5066_b1 );
not ( \5066_b1 , w_23022 );
and ( \7218_b0 , \7217_b0 , w_23023 );
and ( w_23022 , w_23023 , \5066_b0 );
or ( \7219_b1 , \5057_b1 , \5059_b1 );
not ( \5059_b1 , w_23024 );
and ( \7219_b0 , \5057_b0 , w_23025 );
and ( w_23024 , w_23025 , \5059_b0 );
or ( \7220_b1 , \7218_b1 , w_23026 );
or ( \7220_b0 , \7218_b0 , \7219_b0 );
not ( \7219_b0 , w_23027 );
and ( w_23027 , w_23026 , \7219_b1 );
buf ( \7221_b1 , \7220_b1 );
not ( \7221_b1 , w_23028 );
not ( \7221_b0 , w_23029 );
and ( w_23028 , w_23029 , \7220_b0 );
or ( \7222_b1 , \7216_b1 , w_23030 );
or ( \7222_b0 , \7216_b0 , \7221_b0 );
not ( \7221_b0 , w_23031 );
and ( w_23031 , w_23030 , \7221_b1 );
or ( \7223_b1 , \7220_b1 , w_23032 );
or ( \7223_b0 , \7220_b0 , \7215_b0 );
not ( \7215_b0 , w_23033 );
and ( w_23033 , w_23032 , \7215_b1 );
or ( \7224_b1 , \7222_b1 , w_23035 );
not ( w_23035 , w_23036 );
and ( \7224_b0 , \7222_b0 , w_23037 );
and ( w_23036 ,  , w_23037 );
buf ( w_23035 , \7223_b1 );
not ( w_23035 , w_23038 );
not (  , w_23039 );
and ( w_23038 , w_23039 , \7223_b0 );
buf ( \7225_b1 , \7224_b1 );
not ( \7225_b1 , w_23040 );
not ( \7225_b0 , w_23041 );
and ( w_23040 , w_23041 , \7224_b0 );
or ( \7226_b1 , \5051_b1 , \5055_b1 );
xor ( \7226_b0 , \5051_b0 , w_23042 );
not ( w_23042 , w_23043 );
and ( w_23043 , \5055_b1 , \5055_b0 );
or ( \7227_b1 , \7226_b1 , \5067_b1 );
not ( \5067_b1 , w_23044 );
and ( \7227_b0 , \7226_b0 , w_23045 );
and ( w_23044 , w_23045 , \5067_b0 );
or ( \7228_b1 , \5051_b1 , \5055_b1 );
not ( \5055_b1 , w_23046 );
and ( \7228_b0 , \5051_b0 , w_23047 );
and ( w_23046 , w_23047 , \5055_b0 );
or ( \7229_b1 , \7227_b1 , w_23048 );
or ( \7229_b0 , \7227_b0 , \7228_b0 );
not ( \7228_b0 , w_23049 );
and ( w_23049 , w_23048 , \7228_b1 );
buf ( \7230_b1 , \7229_b1 );
not ( \7230_b1 , w_23050 );
not ( \7230_b0 , w_23051 );
and ( w_23050 , w_23051 , \7229_b0 );
or ( \7231_b1 , \7225_b1 , w_23052 );
or ( \7231_b0 , \7225_b0 , \7230_b0 );
not ( \7230_b0 , w_23053 );
and ( w_23053 , w_23052 , \7230_b1 );
or ( \7232_b1 , \7229_b1 , w_23054 );
or ( \7232_b0 , \7229_b0 , \7224_b0 );
not ( \7224_b0 , w_23055 );
and ( w_23055 , w_23054 , \7224_b1 );
or ( \7233_b1 , \7231_b1 , w_23057 );
not ( w_23057 , w_23058 );
and ( \7233_b0 , \7231_b0 , w_23059 );
and ( w_23058 ,  , w_23059 );
buf ( w_23057 , \7232_b1 );
not ( w_23057 , w_23060 );
not (  , w_23061 );
and ( w_23060 , w_23061 , \7232_b0 );
buf ( \7234_b1 , \7233_b1 );
not ( \7234_b1 , w_23062 );
not ( \7234_b0 , w_23063 );
and ( w_23062 , w_23063 , \7233_b0 );
or ( \7235_b1 , \7205_b1 , \7234_b1 );
not ( \7234_b1 , w_23064 );
and ( \7235_b0 , \7205_b0 , w_23065 );
and ( w_23064 , w_23065 , \7234_b0 );
buf ( \7236_b1 , \7205_b1 );
not ( \7236_b1 , w_23066 );
not ( \7236_b0 , w_23067 );
and ( w_23066 , w_23067 , \7205_b0 );
or ( \7237_b1 , \7236_b1 , \7233_b1 );
not ( \7233_b1 , w_23068 );
and ( \7237_b0 , \7236_b0 , w_23069 );
and ( w_23068 , w_23069 , \7233_b0 );
or ( \7238_b1 , \7235_b1 , w_23071 );
not ( w_23071 , w_23072 );
and ( \7238_b0 , \7235_b0 , w_23073 );
and ( w_23072 ,  , w_23073 );
buf ( w_23071 , \7237_b1 );
not ( w_23071 , w_23074 );
not (  , w_23075 );
and ( w_23074 , w_23075 , \7237_b0 );
buf ( \7239_b1 , \5046_b1 );
not ( \7239_b1 , w_23076 );
not ( \7239_b0 , w_23077 );
and ( w_23076 , w_23077 , \5046_b0 );
buf ( \7240_b1 , \7239_b1 );
not ( \7240_b1 , w_23078 );
not ( \7240_b0 , w_23079 );
and ( w_23078 , w_23079 , \7239_b0 );
buf ( \7242_b1 , \7241_b1 );
not ( \7242_b1 , w_23080 );
not ( \7242_b0 , w_23081 );
and ( w_23080 , w_23081 , \7241_b0 );
or ( \7243_b1 , \7240_b1 , w_23082 );
or ( \7243_b0 , \7240_b0 , \7242_b0 );
not ( \7242_b0 , w_23083 );
and ( w_23083 , w_23082 , \7242_b1 );
buf ( \7244_b1 , \7199_b1 );
not ( \7244_b1 , w_23084 );
not ( \7244_b0 , w_23085 );
and ( w_23084 , w_23085 , \7199_b0 );
or ( \7245_b1 , \7243_b1 , w_23087 );
not ( w_23087 , w_23088 );
and ( \7245_b0 , \7243_b0 , w_23089 );
and ( w_23088 ,  , w_23089 );
buf ( w_23087 , \7244_b1 );
not ( w_23087 , w_23090 );
not (  , w_23091 );
and ( w_23090 , w_23091 , \7244_b0 );
or ( \7246_b1 , \7173_b1 , w_23093 );
not ( w_23093 , w_23094 );
and ( \7246_b0 , \7173_b0 , w_23095 );
and ( w_23094 ,  , w_23095 );
buf ( w_23093 , \7202_b1 );
not ( w_23093 , w_23096 );
not (  , w_23097 );
and ( w_23096 , w_23097 , \7202_b0 );
buf ( \7247_b1 , \7246_b1 );
not ( \7247_b1 , w_23098 );
not ( \7247_b0 , w_23099 );
and ( w_23098 , w_23099 , \7246_b0 );
or ( \7248_b1 , \7245_b1 , \7247_b1 );
not ( \7247_b1 , w_23100 );
and ( \7248_b0 , \7245_b0 , w_23101 );
and ( w_23100 , w_23101 , \7247_b0 );
buf ( \7249_b1 , \7245_b1 );
not ( \7249_b1 , w_23102 );
not ( \7249_b0 , w_23103 );
and ( w_23102 , w_23103 , \7245_b0 );
or ( \7250_b1 , \7249_b1 , \7246_b1 );
not ( \7246_b1 , w_23104 );
and ( \7250_b0 , \7249_b0 , w_23105 );
and ( w_23104 , w_23105 , \7246_b0 );
or ( \7251_b1 , \7248_b1 , w_23107 );
not ( w_23107 , w_23108 );
and ( \7251_b0 , \7248_b0 , w_23109 );
and ( w_23108 ,  , w_23109 );
buf ( w_23107 , \7250_b1 );
not ( w_23107 , w_23110 );
not (  , w_23111 );
and ( w_23110 , w_23111 , \7250_b0 );
buf ( \7252_b1 , \5015_b1 );
not ( \7252_b1 , w_23112 );
not ( \7252_b0 , w_23113 );
and ( w_23112 , w_23113 , \5015_b0 );
buf ( \7253_b1 , \7241_b1 );
not ( \7253_b1 , w_23114 );
not ( \7253_b0 , w_23115 );
and ( w_23114 , w_23115 , \7241_b0 );
or ( \7254_b1 , \7252_b1 , w_23116 );
or ( \7254_b0 , \7252_b0 , \7253_b0 );
not ( \7253_b0 , w_23117 );
and ( w_23117 , w_23116 , \7253_b1 );
buf ( \7255_b1 , \7195_b1 );
not ( \7255_b1 , w_23118 );
not ( \7255_b0 , w_23119 );
and ( w_23118 , w_23119 , \7195_b0 );
or ( \7256_b1 , \7254_b1 , w_23121 );
not ( w_23121 , w_23122 );
and ( \7256_b0 , \7254_b0 , w_23123 );
and ( w_23122 ,  , w_23123 );
buf ( w_23121 , \7255_b1 );
not ( w_23121 , w_23124 );
not (  , w_23125 );
and ( w_23124 , w_23125 , \7255_b0 );
or ( \7257_b1 , \5045_b1 , w_23127 );
not ( w_23127 , w_23128 );
and ( \7257_b0 , \5045_b0 , w_23129 );
and ( w_23128 ,  , w_23129 );
buf ( w_23127 , \7198_b1 );
not ( w_23127 , w_23130 );
not (  , w_23131 );
and ( w_23130 , w_23131 , \7198_b0 );
buf ( \7258_b1 , \7257_b1 );
not ( \7258_b1 , w_23132 );
not ( \7258_b0 , w_23133 );
and ( w_23132 , w_23133 , \7257_b0 );
or ( \7259_b1 , \7256_b1 , \7258_b1 );
not ( \7258_b1 , w_23134 );
and ( \7259_b0 , \7256_b0 , w_23135 );
and ( w_23134 , w_23135 , \7258_b0 );
buf ( \7260_b1 , \7256_b1 );
not ( \7260_b1 , w_23136 );
not ( \7260_b0 , w_23137 );
and ( w_23136 , w_23137 , \7256_b0 );
or ( \7261_b1 , \7260_b1 , \7257_b1 );
not ( \7257_b1 , w_23138 );
and ( \7261_b0 , \7260_b0 , w_23139 );
and ( w_23138 , w_23139 , \7257_b0 );
or ( \7262_b1 , \7259_b1 , w_23141 );
not ( w_23141 , w_23142 );
and ( \7262_b0 , \7259_b0 , w_23143 );
and ( w_23142 ,  , w_23143 );
buf ( w_23141 , \7261_b1 );
not ( w_23141 , w_23144 );
not (  , w_23145 );
and ( w_23144 , w_23145 , \7261_b0 );
buf ( \7263_b1 , \5014_b1 );
not ( \7263_b1 , w_23146 );
not ( \7263_b0 , w_23147 );
and ( w_23146 , w_23147 , \5014_b0 );
buf ( \7264_b1 , \7263_b1 );
not ( \7264_b1 , w_23148 );
not ( \7264_b0 , w_23149 );
and ( w_23148 , w_23149 , \7263_b0 );
buf ( \7265_b1 , \7170_b1 );
not ( \7265_b1 , w_23150 );
not ( \7265_b0 , w_23151 );
and ( w_23150 , w_23151 , \7170_b0 );
or ( \7266_b1 , \7264_b1 , w_23152 );
or ( \7266_b0 , \7264_b0 , \7265_b0 );
not ( \7265_b0 , w_23153 );
and ( w_23153 , w_23152 , \7265_b1 );
buf ( \7267_b1 , \7191_b1 );
not ( \7267_b1 , w_23154 );
not ( \7267_b0 , w_23155 );
and ( w_23154 , w_23155 , \7191_b0 );
or ( \7268_b1 , \7266_b1 , w_23157 );
not ( w_23157 , w_23158 );
and ( \7268_b0 , \7266_b0 , w_23159 );
and ( w_23158 ,  , w_23159 );
buf ( w_23157 , \7267_b1 );
not ( w_23157 , w_23160 );
not (  , w_23161 );
and ( w_23160 , w_23161 , \7267_b0 );
or ( \7269_b1 , \4370_b1 , w_23163 );
not ( w_23163 , w_23164 );
and ( \7269_b0 , \4370_b0 , w_23165 );
and ( w_23164 ,  , w_23165 );
buf ( w_23163 , \7194_b1 );
not ( w_23163 , w_23166 );
not (  , w_23167 );
and ( w_23166 , w_23167 , \7194_b0 );
buf ( \7270_b1 , \7269_b1 );
not ( \7270_b1 , w_23168 );
not ( \7270_b0 , w_23169 );
and ( w_23168 , w_23169 , \7269_b0 );
or ( \7271_b1 , \7268_b1 , \7270_b1 );
not ( \7270_b1 , w_23170 );
and ( \7271_b0 , \7268_b0 , w_23171 );
and ( w_23170 , w_23171 , \7270_b0 );
buf ( \7272_b1 , \7268_b1 );
not ( \7272_b1 , w_23172 );
not ( \7272_b0 , w_23173 );
and ( w_23172 , w_23173 , \7268_b0 );
or ( \7273_b1 , \7272_b1 , \7269_b1 );
not ( \7269_b1 , w_23174 );
and ( \7273_b0 , \7272_b0 , w_23175 );
and ( w_23174 , w_23175 , \7269_b0 );
or ( \7274_b1 , \7271_b1 , w_23177 );
not ( w_23177 , w_23178 );
and ( \7274_b0 , \7271_b0 , w_23179 );
and ( w_23178 ,  , w_23179 );
buf ( w_23177 , \7273_b1 );
not ( w_23177 , w_23180 );
not (  , w_23181 );
and ( w_23180 , w_23181 , \7273_b0 );
buf ( \7275_b1 , \5006_b1 );
not ( \7275_b1 , w_23182 );
not ( \7275_b0 , w_23183 );
and ( w_23182 , w_23183 , \5006_b0 );
buf ( \7276_b1 , \7170_b1 );
not ( \7276_b1 , w_23184 );
not ( \7276_b0 , w_23185 );
and ( w_23184 , w_23185 , \7170_b0 );
or ( \7277_b1 , \7275_b1 , w_23186 );
or ( \7277_b0 , \7275_b0 , \7276_b0 );
not ( \7276_b0 , w_23187 );
and ( w_23187 , w_23186 , \7276_b1 );
buf ( \7278_b1 , \7180_b1 );
buf ( \7278_b0 , \7180_b0 );
buf ( \7279_b1 , \7278_b1 );
not ( \7279_b1 , w_23188 );
not ( \7279_b0 , w_23189 );
and ( w_23188 , w_23189 , \7278_b0 );
or ( \7280_b1 , \7279_b1 , \4589_b1 );
not ( \4589_b1 , w_23190 );
and ( \7280_b0 , \7279_b0 , w_23191 );
and ( w_23190 , w_23191 , \4589_b0 );
or ( \7281_b1 , \7280_b1 , w_23193 );
not ( w_23193 , w_23194 );
and ( \7281_b0 , \7280_b0 , w_23195 );
and ( w_23194 ,  , w_23195 );
buf ( w_23193 , \7183_b1 );
not ( w_23193 , w_23196 );
not (  , w_23197 );
and ( w_23196 , w_23197 , \7183_b0 );
or ( \7282_b1 , \7277_b1 , w_23199 );
not ( w_23199 , w_23200 );
and ( \7282_b0 , \7277_b0 , w_23201 );
and ( w_23200 ,  , w_23201 );
buf ( w_23199 , \7281_b1 );
not ( w_23199 , w_23202 );
not (  , w_23203 );
and ( w_23202 , w_23203 , \7281_b0 );
or ( \7283_b1 , \5013_b1 , w_23205 );
not ( w_23205 , w_23206 );
and ( \7283_b0 , \5013_b0 , w_23207 );
and ( w_23206 ,  , w_23207 );
buf ( w_23205 , \7181_b1 );
not ( w_23205 , w_23208 );
not (  , w_23209 );
and ( w_23208 , w_23209 , \7181_b0 );
buf ( \7284_b1 , \7283_b1 );
not ( \7284_b1 , w_23210 );
not ( \7284_b0 , w_23211 );
and ( w_23210 , w_23211 , \7283_b0 );
or ( \7285_b1 , \7282_b1 , \7284_b1 );
not ( \7284_b1 , w_23212 );
and ( \7285_b0 , \7282_b0 , w_23213 );
and ( w_23212 , w_23213 , \7284_b0 );
buf ( \7286_b1 , \7282_b1 );
not ( \7286_b1 , w_23214 );
not ( \7286_b0 , w_23215 );
and ( w_23214 , w_23215 , \7282_b0 );
or ( \7287_b1 , \7286_b1 , \7283_b1 );
not ( \7283_b1 , w_23216 );
and ( \7287_b0 , \7286_b0 , w_23217 );
and ( w_23216 , w_23217 , \7283_b0 );
or ( \7288_b1 , \7285_b1 , w_23219 );
not ( w_23219 , w_23220 );
and ( \7288_b0 , \7285_b0 , w_23221 );
and ( w_23220 ,  , w_23221 );
buf ( w_23219 , \7287_b1 );
not ( w_23219 , w_23222 );
not (  , w_23223 );
and ( w_23222 , w_23223 , \7287_b0 );
buf ( \7289_b1 , \5005_b1 );
not ( \7289_b1 , w_23224 );
not ( \7289_b0 , w_23225 );
and ( w_23224 , w_23225 , \5005_b0 );
buf ( \7290_b1 , \7289_b1 );
not ( \7290_b1 , w_23226 );
not ( \7290_b0 , w_23227 );
and ( w_23226 , w_23227 , \7289_b0 );
buf ( \7291_b1 , \7170_b1 );
not ( \7291_b1 , w_23228 );
not ( \7291_b0 , w_23229 );
and ( w_23228 , w_23229 , \7170_b0 );
or ( \7292_b1 , \7290_b1 , w_23230 );
or ( \7292_b0 , \7290_b0 , \7291_b0 );
not ( \7291_b0 , w_23231 );
and ( w_23231 , w_23230 , \7291_b1 );
or ( \7293_b1 , \7292_b1 , w_23233 );
not ( w_23233 , w_23234 );
and ( \7293_b0 , \7292_b0 , w_23235 );
and ( w_23234 ,  , w_23235 );
buf ( w_23233 , \7278_b1 );
not ( w_23233 , w_23236 );
not (  , w_23237 );
and ( w_23236 , w_23237 , \7278_b0 );
buf ( \7294_b1 , \7183_b1 );
not ( \7294_b1 , w_23238 );
not ( \7294_b0 , w_23239 );
and ( w_23238 , w_23239 , \7183_b0 );
or ( \7295_b1 , \7294_b1 , w_23241 );
not ( w_23241 , w_23242 );
and ( \7295_b0 , \7294_b0 , w_23243 );
and ( w_23242 ,  , w_23243 );
buf ( w_23241 , \4589_b1 );
not ( w_23241 , w_23244 );
not (  , w_23245 );
and ( w_23244 , w_23245 , \4589_b0 );
buf ( \7296_b1 , \7295_b1 );
not ( \7296_b1 , w_23246 );
not ( \7296_b0 , w_23247 );
and ( w_23246 , w_23247 , \7295_b0 );
or ( \7297_b1 , \7293_b1 , \7296_b1 );
not ( \7296_b1 , w_23248 );
and ( \7297_b0 , \7293_b0 , w_23249 );
and ( w_23248 , w_23249 , \7296_b0 );
buf ( \7298_b1 , \7293_b1 );
not ( \7298_b1 , w_23250 );
not ( \7298_b0 , w_23251 );
and ( w_23250 , w_23251 , \7293_b0 );
or ( \7299_b1 , \7298_b1 , \7295_b1 );
not ( \7295_b1 , w_23252 );
and ( \7299_b0 , \7298_b0 , w_23253 );
and ( w_23252 , w_23253 , \7295_b0 );
or ( \7300_b1 , \7297_b1 , w_23255 );
not ( w_23255 , w_23256 );
and ( \7300_b0 , \7297_b0 , w_23257 );
and ( w_23256 ,  , w_23257 );
buf ( w_23255 , \7299_b1 );
not ( w_23255 , w_23258 );
not (  , w_23259 );
and ( w_23258 , w_23259 , \7299_b0 );
buf ( \7301_b1 , \5004_b1 );
not ( \7301_b1 , w_23260 );
not ( \7301_b0 , w_23261 );
and ( w_23260 , w_23261 , \5004_b0 );
buf ( \7302_b1 , \7241_b1 );
not ( \7302_b1 , w_23262 );
not ( \7302_b0 , w_23263 );
and ( w_23262 , w_23263 , \7241_b0 );
or ( \7303_b1 , \7301_b1 , w_23264 );
or ( \7303_b0 , \7301_b0 , \7302_b0 );
not ( \7302_b0 , w_23265 );
and ( w_23265 , w_23264 , \7302_b1 );
buf ( \7304_b1 , \7177_b1 );
buf ( \7304_b0 , \7177_b0 );
or ( \7305_b1 , \7303_b1 , w_23267 );
not ( w_23267 , w_23268 );
and ( \7305_b0 , \7303_b0 , w_23269 );
and ( w_23268 ,  , w_23269 );
buf ( w_23267 , \7304_b1 );
not ( w_23267 , w_23270 );
not (  , w_23271 );
and ( w_23270 , w_23271 , \7304_b0 );
or ( \7306_b1 , \4825_b1 , w_23272 );
or ( \7306_b0 , \4825_b0 , \7179_b0 );
not ( \7179_b0 , w_23273 );
and ( w_23273 , w_23272 , \7179_b1 );
buf ( \7307_b1 , \7306_b1 );
not ( \7307_b1 , w_23274 );
not ( \7307_b0 , w_23275 );
and ( w_23274 , w_23275 , \7306_b0 );
or ( \7308_b1 , \7305_b1 , \7307_b1 );
not ( \7307_b1 , w_23276 );
and ( \7308_b0 , \7305_b0 , w_23277 );
and ( w_23276 , w_23277 , \7307_b0 );
buf ( \7309_b1 , \7305_b1 );
not ( \7309_b1 , w_23278 );
not ( \7309_b0 , w_23279 );
and ( w_23278 , w_23279 , \7305_b0 );
or ( \7310_b1 , \7309_b1 , \7306_b1 );
not ( \7306_b1 , w_23280 );
and ( \7310_b0 , \7309_b0 , w_23281 );
and ( w_23280 , w_23281 , \7306_b0 );
or ( \7311_b1 , \7308_b1 , w_23283 );
not ( w_23283 , w_23284 );
and ( \7311_b0 , \7308_b0 , w_23285 );
and ( w_23284 ,  , w_23285 );
buf ( w_23283 , \7310_b1 );
not ( w_23283 , w_23286 );
not (  , w_23287 );
and ( w_23286 , w_23287 , \7310_b0 );
buf ( \7312_b1 , \5641_b1 );
buf ( \7312_b0 , \5641_b0 );
buf ( \7313_b1 , \7312_b1 );
not ( \7313_b1 , w_23288 );
not ( \7313_b0 , w_23289 );
and ( w_23288 , w_23289 , \7312_b0 );
buf ( \7314_b1 , \5706_b1 );
buf ( \7314_b0 , \5706_b0 );
buf ( \7315_b1 , \5618_b1 );
buf ( \7315_b0 , \5618_b0 );
or ( \7316_b1 , \7314_b1 , \7315_b1 );
not ( \7315_b1 , w_23290 );
and ( \7316_b0 , \7314_b0 , w_23291 );
and ( w_23290 , w_23291 , \7315_b0 );
buf ( \7317_b1 , \7316_b1 );
not ( \7317_b1 , w_23292 );
not ( \7317_b0 , w_23293 );
and ( w_23292 , w_23293 , \7316_b0 );
buf ( \7318_b1 , \7154_b1 );
not ( \7318_b1 , w_23294 );
not ( \7318_b0 , w_23295 );
and ( w_23294 , w_23295 , \7154_b0 );
or ( \7319_b1 , \6290_b1 , w_23297 );
not ( w_23297 , w_23298 );
and ( \7319_b0 , \6290_b0 , w_23299 );
and ( w_23298 ,  , w_23299 );
buf ( w_23297 , \7137_b1 );
not ( w_23297 , w_23300 );
not (  , w_23301 );
and ( w_23300 , w_23301 , \7137_b0 );
or ( \7320_b1 , \7318_b1 , w_23303 );
not ( w_23303 , w_23304 );
and ( \7320_b0 , \7318_b0 , w_23305 );
and ( w_23304 ,  , w_23305 );
buf ( w_23303 , \7319_b1 );
not ( w_23303 , w_23306 );
not (  , w_23307 );
and ( w_23306 , w_23307 , \7319_b0 );
buf ( \7321_b1 , \7320_b1 );
not ( \7321_b1 , w_23308 );
not ( \7321_b0 , w_23309 );
and ( w_23308 , w_23309 , \7320_b0 );
or ( \7322_b1 , \7317_b1 , w_23310 );
or ( \7322_b0 , \7317_b0 , \7321_b0 );
not ( \7321_b0 , w_23311 );
and ( w_23311 , w_23310 , \7321_b1 );
buf ( \7323_b1 , \7159_b1 );
buf ( \7323_b0 , \7159_b0 );
buf ( \7324_b1 , \7323_b1 );
not ( \7324_b1 , w_23312 );
not ( \7324_b0 , w_23313 );
and ( w_23312 , w_23313 , \7323_b0 );
or ( \7325_b1 , \7324_b1 , \7315_b1 );
not ( \7315_b1 , w_23314 );
and ( \7325_b0 , \7324_b0 , w_23315 );
and ( w_23314 , w_23315 , \7315_b0 );
buf ( \7326_b1 , \7160_b1 );
not ( \7326_b1 , w_23316 );
not ( \7326_b0 , w_23317 );
and ( w_23316 , w_23317 , \7160_b0 );
or ( \7327_b1 , \7325_b1 , w_23319 );
not ( w_23319 , w_23320 );
and ( \7327_b0 , \7325_b0 , w_23321 );
and ( w_23320 ,  , w_23321 );
buf ( w_23319 , \7326_b1 );
not ( w_23319 , w_23322 );
not (  , w_23323 );
and ( w_23322 , w_23323 , \7326_b0 );
or ( \7328_b1 , \7322_b1 , w_23325 );
not ( w_23325 , w_23326 );
and ( \7328_b0 , \7322_b0 , w_23327 );
and ( w_23326 ,  , w_23327 );
buf ( w_23325 , \7327_b1 );
not ( w_23325 , w_23328 );
not (  , w_23329 );
and ( w_23328 , w_23329 , \7327_b0 );
buf ( \7329_b1 , \7328_b1 );
not ( \7329_b1 , w_23330 );
not ( \7329_b0 , w_23331 );
and ( w_23330 , w_23331 , \7328_b0 );
or ( \7330_b1 , \7313_b1 , w_23332 );
or ( \7330_b0 , \7313_b0 , \7329_b0 );
not ( \7329_b0 , w_23333 );
and ( w_23333 , w_23332 , \7329_b1 );
or ( \7331_b1 , \7330_b1 , w_23335 );
not ( w_23335 , w_23336 );
and ( \7331_b0 , \7330_b0 , w_23337 );
and ( w_23336 ,  , w_23337 );
buf ( w_23335 , \7165_b1 );
not ( w_23335 , w_23338 );
not (  , w_23339 );
and ( w_23338 , w_23339 , \7165_b0 );
or ( \7332_b1 , \7163_b1 , w_23341 );
not ( w_23341 , w_23342 );
and ( \7332_b0 , \7163_b0 , w_23343 );
and ( w_23342 ,  , w_23343 );
buf ( w_23341 , \7167_b1 );
not ( w_23341 , w_23344 );
not (  , w_23345 );
and ( w_23344 , w_23345 , \7167_b0 );
buf ( \7333_b1 , \7332_b1 );
not ( \7333_b1 , w_23346 );
not ( \7333_b0 , w_23347 );
and ( w_23346 , w_23347 , \7332_b0 );
or ( \7334_b1 , \7331_b1 , \7333_b1 );
not ( \7333_b1 , w_23348 );
and ( \7334_b0 , \7331_b0 , w_23349 );
and ( w_23348 , w_23349 , \7333_b0 );
buf ( \7335_b1 , \7331_b1 );
not ( \7335_b1 , w_23350 );
not ( \7335_b0 , w_23351 );
and ( w_23350 , w_23351 , \7331_b0 );
or ( \7336_b1 , \7335_b1 , \7332_b1 );
not ( \7332_b1 , w_23352 );
and ( \7336_b0 , \7335_b0 , w_23353 );
and ( w_23352 , w_23353 , \7332_b0 );
or ( \7337_b1 , \7334_b1 , w_23355 );
not ( w_23355 , w_23356 );
and ( \7337_b0 , \7334_b0 , w_23357 );
and ( w_23356 ,  , w_23357 );
buf ( w_23355 , \7336_b1 );
not ( w_23355 , w_23358 );
not (  , w_23359 );
and ( w_23358 , w_23359 , \7336_b0 );
or ( \7338_b1 , \7304_b1 , w_23361 );
not ( w_23361 , w_23362 );
and ( \7338_b0 , \7304_b0 , w_23363 );
and ( w_23362 ,  , w_23363 );
buf ( w_23361 , \5004_b1 );
not ( w_23361 , w_23364 );
not (  , w_23365 );
and ( w_23364 , w_23365 , \5004_b0 );
buf ( \7339_b1 , \7338_b1 );
not ( \7339_b1 , w_23366 );
not ( \7339_b0 , w_23367 );
and ( w_23366 , w_23367 , \7338_b0 );
buf ( \7340_b1 , \7241_b1 );
not ( \7340_b1 , w_23368 );
not ( \7340_b0 , w_23369 );
and ( w_23368 , w_23369 , \7241_b0 );
or ( \7341_b1 , \7339_b1 , w_23370 );
or ( \7341_b0 , \7339_b0 , \7340_b0 );
not ( \7340_b0 , w_23371 );
and ( w_23371 , w_23370 , \7340_b1 );
or ( \7342_b1 , \7170_b1 , w_23372 );
or ( \7342_b0 , \7170_b0 , \7338_b0 );
not ( \7338_b0 , w_23373 );
and ( w_23373 , w_23372 , \7338_b1 );
or ( \7343_b1 , \7341_b1 , w_23375 );
not ( w_23375 , w_23376 );
and ( \7343_b0 , \7341_b0 , w_23377 );
and ( w_23376 ,  , w_23377 );
buf ( w_23375 , \7342_b1 );
not ( w_23375 , w_23378 );
not (  , w_23379 );
and ( w_23378 , w_23379 , \7342_b0 );
buf ( \7344_b1 , \7314_b1 );
not ( \7344_b1 , w_23380 );
not ( \7344_b0 , w_23381 );
and ( w_23380 , w_23381 , \7314_b0 );
buf ( \7345_b1 , \7320_b1 );
buf ( \7345_b0 , \7320_b0 );
buf ( \7346_b1 , \7345_b1 );
not ( \7346_b1 , w_23382 );
not ( \7346_b0 , w_23383 );
and ( w_23382 , w_23383 , \7345_b0 );
or ( \7347_b1 , \7344_b1 , w_23384 );
or ( \7347_b0 , \7344_b0 , \7346_b0 );
not ( \7346_b0 , w_23385 );
and ( w_23385 , w_23384 , \7346_b1 );
or ( \7348_b1 , \7347_b1 , w_23387 );
not ( w_23387 , w_23388 );
and ( \7348_b0 , \7347_b0 , w_23389 );
and ( w_23388 ,  , w_23389 );
buf ( w_23387 , \7323_b1 );
not ( w_23387 , w_23390 );
not (  , w_23391 );
and ( w_23390 , w_23391 , \7323_b0 );
or ( \7349_b1 , \7160_b1 , w_23393 );
not ( w_23393 , w_23394 );
and ( \7349_b0 , \7160_b0 , w_23395 );
and ( w_23394 ,  , w_23395 );
buf ( w_23393 , \7315_b1 );
not ( w_23393 , w_23396 );
not (  , w_23397 );
and ( w_23396 , w_23397 , \7315_b0 );
buf ( \7350_b1 , \7349_b1 );
not ( \7350_b1 , w_23398 );
not ( \7350_b0 , w_23399 );
and ( w_23398 , w_23399 , \7349_b0 );
or ( \7351_b1 , \7348_b1 , \7350_b1 );
not ( \7350_b1 , w_23400 );
and ( \7351_b0 , \7348_b0 , w_23401 );
and ( w_23400 , w_23401 , \7350_b0 );
buf ( \7352_b1 , \7348_b1 );
not ( \7352_b1 , w_23402 );
not ( \7352_b0 , w_23403 );
and ( w_23402 , w_23403 , \7348_b0 );
or ( \7353_b1 , \7352_b1 , \7349_b1 );
not ( \7349_b1 , w_23404 );
and ( \7353_b0 , \7352_b0 , w_23405 );
and ( w_23404 , w_23405 , \7349_b0 );
or ( \7354_b1 , \7351_b1 , w_23407 );
not ( w_23407 , w_23408 );
and ( \7354_b0 , \7351_b0 , w_23409 );
and ( w_23408 ,  , w_23409 );
buf ( w_23407 , \7353_b1 );
not ( w_23407 , w_23410 );
not (  , w_23411 );
and ( w_23410 , w_23411 , \7353_b0 );
or ( \7355_b1 , \7323_b1 , w_23413 );
not ( w_23413 , w_23414 );
and ( \7355_b0 , \7323_b0 , w_23415 );
and ( w_23414 ,  , w_23415 );
buf ( w_23413 , \7314_b1 );
not ( w_23413 , w_23416 );
not (  , w_23417 );
and ( w_23416 , w_23417 , \7314_b0 );
buf ( \7356_b1 , \7355_b1 );
not ( \7356_b1 , w_23418 );
not ( \7356_b0 , w_23419 );
and ( w_23418 , w_23419 , \7355_b0 );
or ( \7357_b1 , \7345_b1 , \7356_b1 );
not ( \7356_b1 , w_23420 );
and ( \7357_b0 , \7345_b0 , w_23421 );
and ( w_23420 , w_23421 , \7356_b0 );
buf ( \7358_b1 , \7345_b1 );
not ( \7358_b1 , w_23422 );
not ( \7358_b0 , w_23423 );
and ( w_23422 , w_23423 , \7345_b0 );
or ( \7359_b1 , \7358_b1 , \7355_b1 );
not ( \7355_b1 , w_23424 );
and ( \7359_b0 , \7358_b0 , w_23425 );
and ( w_23424 , w_23425 , \7355_b0 );
or ( \7360_b1 , \7357_b1 , w_23427 );
not ( w_23427 , w_23428 );
and ( \7360_b0 , \7357_b0 , w_23429 );
and ( w_23428 ,  , w_23429 );
buf ( w_23427 , \7359_b1 );
not ( w_23427 , w_23430 );
not (  , w_23431 );
and ( w_23430 , w_23431 , \7359_b0 );
buf ( \7361_b1 , \6034_b1 );
buf ( \7361_b0 , \6034_b0 );
buf ( \7362_b1 , \7361_b1 );
not ( \7362_b1 , w_23432 );
not ( \7362_b0 , w_23433 );
and ( w_23432 , w_23433 , \7361_b0 );
buf ( \7363_b1 , \6279_b1 );
not ( \7363_b1 , w_23434 );
not ( \7363_b0 , w_23435 );
and ( w_23434 , w_23435 , \6279_b0 );
buf ( \7364_b1 , \7137_b1 );
not ( \7364_b1 , w_23436 );
not ( \7364_b0 , w_23437 );
and ( w_23436 , w_23437 , \7137_b0 );
or ( \7365_b1 , \7363_b1 , w_23438 );
or ( \7365_b0 , \7363_b0 , \7364_b0 );
not ( \7364_b0 , w_23439 );
and ( w_23439 , w_23438 , \7364_b1 );
or ( \7366_b1 , \7365_b1 , w_23441 );
not ( w_23441 , w_23442 );
and ( \7366_b0 , \7365_b0 , w_23443 );
and ( w_23442 ,  , w_23443 );
buf ( w_23441 , \7145_b1 );
not ( w_23441 , w_23444 );
not (  , w_23445 );
and ( w_23444 , w_23445 , \7145_b0 );
buf ( \7367_b1 , \7366_b1 );
not ( \7367_b1 , w_23446 );
not ( \7367_b0 , w_23447 );
and ( w_23446 , w_23447 , \7366_b0 );
or ( \7368_b1 , \7362_b1 , w_23448 );
or ( \7368_b0 , \7362_b0 , \7367_b0 );
not ( \7367_b0 , w_23449 );
and ( w_23449 , w_23448 , \7367_b1 );
or ( \7369_b1 , \7368_b1 , w_23451 );
not ( w_23451 , w_23452 );
and ( \7369_b0 , \7368_b0 , w_23453 );
and ( w_23452 ,  , w_23453 );
buf ( w_23451 , \7147_b1 );
not ( w_23451 , w_23454 );
not (  , w_23455 );
and ( w_23454 , w_23455 , \7147_b0 );
or ( \7370_b1 , \6288_b1 , w_23457 );
not ( w_23457 , w_23458 );
and ( \7370_b0 , \6288_b0 , w_23459 );
and ( w_23458 ,  , w_23459 );
buf ( w_23457 , \7153_b1 );
not ( w_23457 , w_23460 );
not (  , w_23461 );
and ( w_23460 , w_23461 , \7153_b0 );
buf ( \7371_b1 , \7370_b1 );
not ( \7371_b1 , w_23462 );
not ( \7371_b0 , w_23463 );
and ( w_23462 , w_23463 , \7370_b0 );
or ( \7372_b1 , \7369_b1 , \7371_b1 );
not ( \7371_b1 , w_23464 );
and ( \7372_b0 , \7369_b0 , w_23465 );
and ( w_23464 , w_23465 , \7371_b0 );
buf ( \7373_b1 , \7369_b1 );
not ( \7373_b1 , w_23466 );
not ( \7373_b0 , w_23467 );
and ( w_23466 , w_23467 , \7369_b0 );
or ( \7374_b1 , \7373_b1 , \7370_b1 );
not ( \7370_b1 , w_23468 );
and ( \7374_b0 , \7373_b0 , w_23469 );
and ( w_23468 , w_23469 , \7370_b0 );
or ( \7375_b1 , \7372_b1 , w_23471 );
not ( w_23471 , w_23472 );
and ( \7375_b0 , \7372_b0 , w_23473 );
and ( w_23472 ,  , w_23473 );
buf ( w_23471 , \7374_b1 );
not ( w_23471 , w_23474 );
not (  , w_23475 );
and ( w_23474 , w_23475 , \7374_b0 );
or ( \7376_b1 , \7147_b1 , w_23477 );
not ( w_23477 , w_23478 );
and ( \7376_b0 , \7147_b0 , w_23479 );
and ( w_23478 ,  , w_23479 );
buf ( w_23477 , \7361_b1 );
not ( w_23477 , w_23480 );
not (  , w_23481 );
and ( w_23480 , w_23481 , \7361_b0 );
buf ( \7377_b1 , \7376_b1 );
not ( \7377_b1 , w_23482 );
not ( \7377_b0 , w_23483 );
and ( w_23482 , w_23483 , \7376_b0 );
or ( \7378_b1 , \7366_b1 , \7377_b1 );
not ( \7377_b1 , w_23484 );
and ( \7378_b0 , \7366_b0 , w_23485 );
and ( w_23484 , w_23485 , \7377_b0 );
buf ( \7379_b1 , \7366_b1 );
not ( \7379_b1 , w_23486 );
not ( \7379_b0 , w_23487 );
and ( w_23486 , w_23487 , \7366_b0 );
or ( \7380_b1 , \7379_b1 , \7376_b1 );
not ( \7376_b1 , w_23488 );
and ( \7380_b0 , \7379_b0 , w_23489 );
and ( w_23488 , w_23489 , \7376_b0 );
or ( \7381_b1 , \7378_b1 , w_23491 );
not ( w_23491 , w_23492 );
and ( \7381_b0 , \7378_b0 , w_23493 );
and ( w_23492 ,  , w_23493 );
buf ( w_23491 , \7380_b1 );
not ( w_23491 , w_23494 );
not (  , w_23495 );
and ( w_23494 , w_23495 , \7380_b0 );
buf ( \7382_b1 , \6278_b1 );
not ( \7382_b1 , w_23496 );
not ( \7382_b0 , w_23497 );
and ( w_23496 , w_23497 , \6278_b0 );
buf ( \7383_b1 , \7137_b1 );
buf ( \7383_b0 , \7137_b0 );
buf ( \7384_b1 , \7383_b1 );
not ( \7384_b1 , w_23498 );
not ( \7384_b0 , w_23499 );
and ( w_23498 , w_23499 , \7383_b0 );
or ( \7385_b1 , \7382_b1 , w_23500 );
or ( \7385_b0 , \7382_b0 , \7384_b0 );
not ( \7384_b0 , w_23501 );
and ( w_23501 , w_23500 , \7384_b1 );
or ( \7386_b1 , \7385_b1 , w_23503 );
not ( w_23503 , w_23504 );
and ( \7386_b0 , \7385_b0 , w_23505 );
and ( w_23504 ,  , w_23505 );
buf ( w_23503 , \7142_b1 );
not ( w_23503 , w_23506 );
not (  , w_23507 );
and ( w_23506 , w_23507 , \7142_b0 );
or ( \7387_b1 , \6151_b1 , w_23509 );
not ( w_23509 , w_23510 );
and ( \7387_b0 , \6151_b0 , w_23511 );
and ( w_23510 ,  , w_23511 );
buf ( w_23509 , \7140_b1 );
not ( w_23509 , w_23512 );
not (  , w_23513 );
and ( w_23512 , w_23513 , \7140_b0 );
buf ( \7388_b1 , \7387_b1 );
not ( \7388_b1 , w_23514 );
not ( \7388_b0 , w_23515 );
and ( w_23514 , w_23515 , \7387_b0 );
or ( \7389_b1 , \7386_b1 , \7388_b1 );
not ( \7388_b1 , w_23516 );
and ( \7389_b0 , \7386_b0 , w_23517 );
and ( w_23516 , w_23517 , \7388_b0 );
buf ( \7390_b1 , \7386_b1 );
not ( \7390_b1 , w_23518 );
not ( \7390_b0 , w_23519 );
and ( w_23518 , w_23519 , \7386_b0 );
or ( \7391_b1 , \7390_b1 , \7387_b1 );
not ( \7387_b1 , w_23520 );
and ( \7391_b0 , \7390_b0 , w_23521 );
and ( w_23520 , w_23521 , \7387_b0 );
or ( \7392_b1 , \7389_b1 , w_23523 );
not ( w_23523 , w_23524 );
and ( \7392_b0 , \7389_b0 , w_23525 );
and ( w_23524 ,  , w_23525 );
buf ( w_23523 , \7391_b1 );
not ( w_23523 , w_23526 );
not (  , w_23527 );
and ( w_23526 , w_23527 , \7391_b0 );
or ( \7393_b1 , \7142_b1 , w_23529 );
not ( w_23529 , w_23530 );
and ( \7393_b0 , \7142_b0 , w_23531 );
and ( w_23530 ,  , w_23531 );
buf ( w_23529 , \6278_b1 );
not ( w_23529 , w_23532 );
not (  , w_23533 );
and ( w_23532 , w_23533 , \6278_b0 );
buf ( \7394_b1 , \7393_b1 );
not ( \7394_b1 , w_23534 );
not ( \7394_b0 , w_23535 );
and ( w_23534 , w_23535 , \7393_b0 );
buf ( \7395_b1 , \7383_b1 );
not ( \7395_b1 , w_23536 );
not ( \7395_b0 , w_23537 );
and ( w_23536 , w_23537 , \7383_b0 );
or ( \7396_b1 , \7394_b1 , w_23538 );
or ( \7396_b0 , \7394_b0 , \7395_b0 );
not ( \7395_b0 , w_23539 );
and ( w_23539 , w_23538 , \7395_b1 );
or ( \7397_b1 , \7393_b1 , w_23540 );
or ( \7397_b0 , \7393_b0 , \7383_b0 );
not ( \7383_b0 , w_23541 );
and ( w_23541 , w_23540 , \7383_b1 );
or ( \7398_b1 , \7396_b1 , w_23543 );
not ( w_23543 , w_23544 );
and ( \7398_b0 , \7396_b0 , w_23545 );
and ( w_23544 ,  , w_23545 );
buf ( w_23543 , \7397_b1 );
not ( w_23543 , w_23546 );
not (  , w_23547 );
and ( w_23546 , w_23547 , \7397_b0 );
buf ( \7399_b1 , \7068_b1 );
buf ( \7399_b0 , \7068_b0 );
buf ( \7400_b1 , \7399_b1 );
not ( \7400_b1 , w_23548 );
not ( \7400_b0 , w_23549 );
and ( w_23548 , w_23549 , \7399_b0 );
buf ( \7401_b1 , \7115_b1 );
not ( \7401_b1 , w_23550 );
not ( \7401_b0 , w_23551 );
and ( w_23550 , w_23551 , \7115_b0 );
buf ( \7402_b1 , \6983_b1 );
not ( \7402_b1 , w_23552 );
not ( \7402_b0 , w_23553 );
and ( w_23552 , w_23553 , \6983_b0 );
or ( \7403_b1 , \7401_b1 , w_23554 );
or ( \7403_b0 , \7401_b0 , \7402_b0 );
not ( \7402_b0 , w_23555 );
and ( w_23555 , w_23554 , \7402_b1 );
buf ( \7404_b1 , \7127_b1 );
buf ( \7404_b0 , \7127_b0 );
buf ( \7405_b1 , \7404_b1 );
not ( \7405_b1 , w_23556 );
not ( \7405_b0 , w_23557 );
and ( w_23556 , w_23557 , \7404_b0 );
or ( \7406_b1 , \7405_b1 , w_23559 );
not ( w_23559 , w_23560 );
and ( \7406_b0 , \7405_b0 , w_23561 );
and ( w_23560 ,  , w_23561 );
buf ( w_23559 , \7124_b1 );
not ( w_23559 , w_23562 );
not (  , w_23563 );
and ( w_23562 , w_23563 , \7124_b0 );
or ( \7407_b1 , \7403_b1 , w_23565 );
not ( w_23565 , w_23566 );
and ( \7407_b0 , \7403_b0 , w_23567 );
and ( w_23566 ,  , w_23567 );
buf ( w_23565 , \7406_b1 );
not ( w_23565 , w_23568 );
not (  , w_23569 );
and ( w_23568 , w_23569 , \7406_b0 );
buf ( \7408_b1 , \7407_b1 );
not ( \7408_b1 , w_23570 );
not ( \7408_b0 , w_23571 );
and ( w_23570 , w_23571 , \7407_b0 );
or ( \7409_b1 , \7400_b1 , w_23572 );
or ( \7409_b0 , \7400_b0 , \7408_b0 );
not ( \7408_b0 , w_23573 );
and ( w_23573 , w_23572 , \7408_b1 );
buf ( \7410_b1 , \7129_b1 );
not ( \7410_b1 , w_23574 );
not ( \7410_b0 , w_23575 );
and ( w_23574 , w_23575 , \7129_b0 );
buf ( \7411_b1 , \7410_b1 );
not ( \7411_b1 , w_23576 );
not ( \7411_b0 , w_23577 );
and ( w_23576 , w_23577 , \7410_b0 );
or ( \7412_b1 , \7409_b1 , w_23579 );
not ( w_23579 , w_23580 );
and ( \7412_b0 , \7409_b0 , w_23581 );
and ( w_23580 ,  , w_23581 );
buf ( w_23579 , \7411_b1 );
not ( w_23579 , w_23582 );
not (  , w_23583 );
and ( w_23582 , w_23583 , \7411_b0 );
or ( \7413_b1 , \7119_b1 , w_23585 );
not ( w_23585 , w_23586 );
and ( \7413_b0 , \7119_b0 , w_23587 );
and ( w_23586 ,  , w_23587 );
buf ( w_23585 , \7135_b1 );
not ( w_23585 , w_23588 );
not (  , w_23589 );
and ( w_23588 , w_23589 , \7135_b0 );
buf ( \7414_b1 , \7413_b1 );
not ( \7414_b1 , w_23590 );
not ( \7414_b0 , w_23591 );
and ( w_23590 , w_23591 , \7413_b0 );
or ( \7415_b1 , \7412_b1 , \7414_b1 );
not ( \7414_b1 , w_23592 );
and ( \7415_b0 , \7412_b0 , w_23593 );
and ( w_23592 , w_23593 , \7414_b0 );
buf ( \7416_b1 , \7412_b1 );
not ( \7416_b1 , w_23594 );
not ( \7416_b0 , w_23595 );
and ( w_23594 , w_23595 , \7412_b0 );
or ( \7417_b1 , \7416_b1 , \7413_b1 );
not ( \7413_b1 , w_23596 );
and ( \7417_b0 , \7416_b0 , w_23597 );
and ( w_23596 , w_23597 , \7413_b0 );
or ( \7418_b1 , \7415_b1 , w_23599 );
not ( w_23599 , w_23600 );
and ( \7418_b0 , \7415_b0 , w_23601 );
and ( w_23600 ,  , w_23601 );
buf ( w_23599 , \7417_b1 );
not ( w_23599 , w_23602 );
not (  , w_23603 );
and ( w_23602 , w_23603 , \7417_b0 );
or ( \7419_b1 , \7165_b1 , w_23605 );
not ( w_23605 , w_23606 );
and ( \7419_b0 , \7165_b0 , w_23607 );
and ( w_23606 ,  , w_23607 );
buf ( w_23605 , \7312_b1 );
not ( w_23605 , w_23608 );
not (  , w_23609 );
and ( w_23608 , w_23609 , \7312_b0 );
buf ( \7420_b1 , \7410_b1 );
not ( \7420_b1 , w_23610 );
not ( \7420_b0 , w_23611 );
and ( w_23610 , w_23611 , \7410_b0 );
or ( \7421_b1 , \7420_b1 , w_23613 );
not ( w_23613 , w_23614 );
and ( \7421_b0 , \7420_b0 , w_23615 );
and ( w_23614 ,  , w_23615 );
buf ( w_23613 , \7399_b1 );
not ( w_23613 , w_23616 );
not (  , w_23617 );
and ( w_23616 , w_23617 , \7399_b0 );
buf ( \7422_b1 , \7421_b1 );
not ( \7422_b1 , w_23618 );
not ( \7422_b0 , w_23619 );
and ( w_23618 , w_23619 , \7421_b0 );
buf ( \7423_b1 , \7407_b1 );
not ( \7423_b1 , w_23620 );
not ( \7423_b0 , w_23621 );
and ( w_23620 , w_23621 , \7407_b0 );
or ( \7424_b1 , \7422_b1 , w_23622 );
or ( \7424_b0 , \7422_b0 , \7423_b0 );
not ( \7423_b0 , w_23623 );
and ( w_23623 , w_23622 , \7423_b1 );
or ( \7425_b1 , \7421_b1 , w_23624 );
or ( \7425_b0 , \7421_b0 , \7407_b0 );
not ( \7407_b0 , w_23625 );
and ( w_23625 , w_23624 , \7407_b1 );
or ( \7426_b1 , \7424_b1 , w_23627 );
not ( w_23627 , w_23628 );
and ( \7426_b0 , \7424_b0 , w_23629 );
and ( w_23628 ,  , w_23629 );
buf ( w_23627 , \7425_b1 );
not ( w_23627 , w_23630 );
not (  , w_23631 );
and ( w_23630 , w_23631 , \7425_b0 );
buf ( \7427_b1 , \7114_b1 );
not ( \7427_b1 , w_23632 );
not ( \7427_b0 , w_23633 );
and ( w_23632 , w_23633 , \7114_b0 );
buf ( \7428_b1 , \6983_b1 );
not ( \7428_b1 , w_23634 );
not ( \7428_b0 , w_23635 );
and ( w_23634 , w_23635 , \6983_b0 );
or ( \7429_b1 , \7427_b1 , w_23636 );
or ( \7429_b0 , \7427_b0 , \7428_b0 );
not ( \7428_b0 , w_23637 );
and ( w_23637 , w_23636 , \7428_b1 );
or ( \7430_b1 , \7429_b1 , w_23639 );
not ( w_23639 , w_23640 );
and ( \7430_b0 , \7429_b0 , w_23641 );
and ( w_23640 ,  , w_23641 );
buf ( w_23639 , \7123_b1 );
not ( w_23639 , w_23642 );
not (  , w_23643 );
and ( w_23642 , w_23643 , \7123_b0 );
or ( \7431_b1 , \7404_b1 , w_23645 );
not ( w_23645 , w_23646 );
and ( \7431_b0 , \7404_b0 , w_23647 );
and ( w_23646 ,  , w_23647 );
buf ( w_23645 , \7103_b1 );
not ( w_23645 , w_23648 );
not (  , w_23649 );
and ( w_23648 , w_23649 , \7103_b0 );
buf ( \7432_b1 , \7431_b1 );
not ( \7432_b1 , w_23650 );
not ( \7432_b0 , w_23651 );
and ( w_23650 , w_23651 , \7431_b0 );
or ( \7433_b1 , \7430_b1 , \7432_b1 );
not ( \7432_b1 , w_23652 );
and ( \7433_b0 , \7430_b0 , w_23653 );
and ( w_23652 , w_23653 , \7432_b0 );
buf ( \7434_b1 , \7430_b1 );
not ( \7434_b1 , w_23654 );
not ( \7434_b0 , w_23655 );
and ( w_23654 , w_23655 , \7430_b0 );
or ( \7435_b1 , \7434_b1 , \7431_b1 );
not ( \7431_b1 , w_23656 );
and ( \7435_b0 , \7434_b0 , w_23657 );
and ( w_23656 , w_23657 , \7431_b0 );
or ( \7436_b1 , \7433_b1 , w_23659 );
not ( w_23659 , w_23660 );
and ( \7436_b0 , \7433_b0 , w_23661 );
and ( w_23660 ,  , w_23661 );
buf ( w_23659 , \7435_b1 );
not ( w_23659 , w_23662 );
not (  , w_23663 );
and ( w_23662 , w_23663 , \7435_b0 );
buf ( \7437_b1 , \6964_b1 );
buf ( \7437_b0 , \6964_b0 );
buf ( \7438_b1 , \7437_b1 );
not ( \7438_b1 , w_23664 );
not ( \7438_b0 , w_23665 );
and ( w_23664 , w_23665 , \7437_b0 );
buf ( \7439_b1 , \6954_b1 );
not ( \7439_b1 , w_23666 );
not ( \7439_b0 , w_23667 );
and ( w_23666 , w_23667 , \6954_b0 );
buf ( \7440_b1 , \6601_b1 );
not ( \7440_b1 , w_23668 );
not ( \7440_b0 , w_23669 );
and ( w_23668 , w_23669 , \6601_b0 );
or ( \7441_b1 , \7439_b1 , w_23670 );
or ( \7441_b0 , \7439_b0 , \7440_b0 );
not ( \7440_b0 , w_23671 );
and ( w_23671 , w_23670 , \7440_b1 );
or ( \7442_b1 , \6978_b1 , w_23673 );
not ( w_23673 , w_23674 );
and ( \7442_b0 , \6978_b0 , w_23675 );
and ( w_23674 ,  , w_23675 );
buf ( w_23673 , \6944_b1 );
not ( w_23673 , w_23676 );
not (  , w_23677 );
and ( w_23676 , w_23677 , \6944_b0 );
or ( \7443_b1 , \7441_b1 , w_23679 );
not ( w_23679 , w_23680 );
and ( \7443_b0 , \7441_b0 , w_23681 );
and ( w_23680 ,  , w_23681 );
buf ( w_23679 , \7442_b1 );
not ( w_23679 , w_23682 );
not (  , w_23683 );
and ( w_23682 , w_23683 , \7442_b0 );
buf ( \7444_b1 , \7443_b1 );
not ( \7444_b1 , w_23684 );
not ( \7444_b0 , w_23685 );
and ( w_23684 , w_23685 , \7443_b0 );
or ( \7445_b1 , \7438_b1 , w_23686 );
or ( \7445_b0 , \7438_b0 , \7444_b0 );
not ( \7444_b0 , w_23687 );
and ( w_23687 , w_23686 , \7444_b1 );
or ( \7446_b1 , \7445_b1 , w_23689 );
not ( w_23689 , w_23690 );
and ( \7446_b0 , \7445_b0 , w_23691 );
and ( w_23690 ,  , w_23691 );
buf ( w_23689 , \6973_b1 );
not ( w_23689 , w_23692 );
not (  , w_23693 );
and ( w_23692 , w_23693 , \6973_b0 );
or ( \7447_b1 , \6981_b1 , w_23695 );
not ( w_23695 , w_23696 );
and ( \7447_b0 , \6981_b0 , w_23697 );
and ( w_23696 ,  , w_23697 );
buf ( w_23695 , \6970_b1 );
not ( w_23695 , w_23698 );
not (  , w_23699 );
and ( w_23698 , w_23699 , \6970_b0 );
buf ( \7448_b1 , \7447_b1 );
not ( \7448_b1 , w_23700 );
not ( \7448_b0 , w_23701 );
and ( w_23700 , w_23701 , \7447_b0 );
or ( \7449_b1 , \7446_b1 , \7448_b1 );
not ( \7448_b1 , w_23702 );
and ( \7449_b0 , \7446_b0 , w_23703 );
and ( w_23702 , w_23703 , \7448_b0 );
buf ( \7450_b1 , \7446_b1 );
not ( \7450_b1 , w_23704 );
not ( \7450_b0 , w_23705 );
and ( w_23704 , w_23705 , \7446_b0 );
or ( \7451_b1 , \7450_b1 , \7447_b1 );
not ( \7447_b1 , w_23706 );
and ( \7451_b0 , \7450_b0 , w_23707 );
and ( w_23706 , w_23707 , \7447_b0 );
or ( \7452_b1 , \7449_b1 , w_23709 );
not ( w_23709 , w_23710 );
and ( \7452_b0 , \7449_b0 , w_23711 );
and ( w_23710 ,  , w_23711 );
buf ( w_23709 , \7451_b1 );
not ( w_23709 , w_23712 );
not (  , w_23713 );
and ( w_23712 , w_23713 , \7451_b0 );
or ( \7453_b1 , \7114_b1 , w_23715 );
not ( w_23715 , w_23716 );
and ( \7453_b0 , \7114_b0 , w_23717 );
and ( w_23716 ,  , w_23717 );
buf ( w_23715 , \7123_b1 );
not ( w_23715 , w_23718 );
not (  , w_23719 );
and ( w_23718 , w_23719 , \7123_b0 );
buf ( \7454_b1 , \7453_b1 );
not ( \7454_b1 , w_23720 );
not ( \7454_b0 , w_23721 );
and ( w_23720 , w_23721 , \7453_b0 );
buf ( \7455_b1 , \6983_b1 );
not ( \7455_b1 , w_23722 );
not ( \7455_b0 , w_23723 );
and ( w_23722 , w_23723 , \6983_b0 );
or ( \7456_b1 , \7454_b1 , w_23724 );
or ( \7456_b0 , \7454_b0 , \7455_b0 );
not ( \7455_b0 , w_23725 );
and ( w_23725 , w_23724 , \7455_b1 );
or ( \7457_b1 , \7453_b1 , w_23726 );
or ( \7457_b0 , \7453_b0 , \6983_b0 );
not ( \6983_b0 , w_23727 );
and ( w_23727 , w_23726 , \6983_b1 );
or ( \7458_b1 , \7456_b1 , w_23729 );
not ( w_23729 , w_23730 );
and ( \7458_b0 , \7456_b0 , w_23731 );
and ( w_23730 ,  , w_23731 );
buf ( w_23729 , \7457_b1 );
not ( w_23729 , w_23732 );
not (  , w_23733 );
and ( w_23732 , w_23733 , \7457_b0 );
or ( \7459_b1 , \7437_b1 , w_23735 );
not ( w_23735 , w_23736 );
and ( \7459_b0 , \7437_b0 , w_23737 );
and ( w_23736 ,  , w_23737 );
buf ( w_23735 , \6973_b1 );
not ( w_23735 , w_23738 );
not (  , w_23739 );
and ( w_23738 , w_23739 , \6973_b0 );
buf ( \7460_b1 , \7459_b1 );
not ( \7460_b1 , w_23740 );
not ( \7460_b0 , w_23741 );
and ( w_23740 , w_23741 , \7459_b0 );
or ( \7461_b1 , \7443_b1 , \7460_b1 );
not ( \7460_b1 , w_23742 );
and ( \7461_b0 , \7443_b0 , w_23743 );
and ( w_23742 , w_23743 , \7460_b0 );
buf ( \7462_b1 , \7443_b1 );
not ( \7462_b1 , w_23744 );
not ( \7462_b0 , w_23745 );
and ( w_23744 , w_23745 , \7443_b0 );
or ( \7463_b1 , \7462_b1 , \7459_b1 );
not ( \7459_b1 , w_23746 );
and ( \7463_b0 , \7462_b0 , w_23747 );
and ( w_23746 , w_23747 , \7459_b0 );
or ( \7464_b1 , \7461_b1 , w_23749 );
not ( w_23749 , w_23750 );
and ( \7464_b0 , \7461_b0 , w_23751 );
and ( w_23750 ,  , w_23751 );
buf ( w_23749 , \7463_b1 );
not ( w_23749 , w_23752 );
not (  , w_23753 );
and ( w_23752 , w_23753 , \7463_b0 );
buf ( \7465_b1 , \6953_b1 );
not ( \7465_b1 , w_23754 );
not ( \7465_b0 , w_23755 );
and ( w_23754 , w_23755 , \6953_b0 );
buf ( \7466_b1 , \6601_b1 );
not ( \7466_b1 , w_23756 );
not ( \7466_b0 , w_23757 );
and ( w_23756 , w_23757 , \6601_b0 );
or ( \7467_b1 , \7465_b1 , w_23758 );
or ( \7467_b0 , \7465_b0 , \7466_b0 );
not ( \7466_b0 , w_23759 );
and ( w_23759 , w_23758 , \7466_b1 );
or ( \7468_b1 , \7467_b1 , w_23761 );
not ( w_23761 , w_23762 );
and ( \7468_b0 , \7467_b0 , w_23763 );
and ( w_23762 ,  , w_23763 );
buf ( w_23761 , \6977_b1 );
not ( w_23761 , w_23764 );
not (  , w_23765 );
and ( w_23764 , w_23765 , \6977_b0 );
or ( \7469_b1 , \6976_b1 , w_23767 );
not ( w_23767 , w_23768 );
and ( \7469_b0 , \6976_b0 , w_23769 );
and ( w_23768 ,  , w_23769 );
buf ( w_23767 , \6944_b1 );
not ( w_23767 , w_23770 );
not (  , w_23771 );
and ( w_23770 , w_23771 , \6944_b0 );
buf ( \7470_b1 , \7469_b1 );
not ( \7470_b1 , w_23772 );
not ( \7470_b0 , w_23773 );
and ( w_23772 , w_23773 , \7469_b0 );
or ( \7471_b1 , \7468_b1 , \7470_b1 );
not ( \7470_b1 , w_23774 );
and ( \7471_b0 , \7468_b0 , w_23775 );
and ( w_23774 , w_23775 , \7470_b0 );
buf ( \7472_b1 , \7468_b1 );
not ( \7472_b1 , w_23776 );
not ( \7472_b0 , w_23777 );
and ( w_23776 , w_23777 , \7468_b0 );
or ( \7473_b1 , \7472_b1 , \7469_b1 );
not ( \7469_b1 , w_23778 );
and ( \7473_b0 , \7472_b0 , w_23779 );
and ( w_23778 , w_23779 , \7469_b0 );
or ( \7474_b1 , \7471_b1 , w_23781 );
not ( w_23781 , w_23782 );
and ( \7474_b0 , \7471_b0 , w_23783 );
and ( w_23782 ,  , w_23783 );
buf ( w_23781 , \7473_b1 );
not ( w_23781 , w_23784 );
not (  , w_23785 );
and ( w_23784 , w_23785 , \7473_b0 );
or ( \7475_b1 , \6977_b1 , w_23787 );
not ( w_23787 , w_23788 );
and ( \7475_b0 , \6977_b0 , w_23789 );
and ( w_23788 ,  , w_23789 );
buf ( w_23787 , \6953_b1 );
not ( w_23787 , w_23790 );
not (  , w_23791 );
and ( w_23790 , w_23791 , \6953_b0 );
buf ( \7476_b1 , \7475_b1 );
not ( \7476_b1 , w_23792 );
not ( \7476_b0 , w_23793 );
and ( w_23792 , w_23793 , \7475_b0 );
buf ( \7477_b1 , \6601_b1 );
not ( \7477_b1 , w_23794 );
not ( \7477_b0 , w_23795 );
and ( w_23794 , w_23795 , \6601_b0 );
or ( \7478_b1 , \7476_b1 , w_23796 );
or ( \7478_b0 , \7476_b0 , \7477_b0 );
not ( \7477_b0 , w_23797 );
and ( w_23797 , w_23796 , \7477_b1 );
or ( \7479_b1 , \7475_b1 , w_23798 );
or ( \7479_b0 , \7475_b0 , \6601_b0 );
not ( \6601_b0 , w_23799 );
and ( w_23799 , w_23798 , \6601_b1 );
or ( \7480_b1 , \7478_b1 , w_23801 );
not ( w_23801 , w_23802 );
and ( \7480_b0 , \7478_b0 , w_23803 );
and ( w_23802 ,  , w_23803 );
buf ( w_23801 , \7479_b1 );
not ( w_23801 , w_23804 );
not (  , w_23805 );
and ( w_23804 , w_23805 , \7479_b0 );
or ( \7481_b1 , \6364_b1 , \6428_b1 );
xor ( \7481_b0 , \6364_b0 , w_23806 );
not ( w_23806 , w_23807 );
and ( w_23807 , \6428_b1 , \6428_b0 );
or ( \7482_b1 , \7481_b1 , \6598_b1 );
xor ( \7482_b0 , \7481_b0 , w_23808 );
not ( w_23808 , w_23809 );
and ( w_23809 , \6598_b1 , \6598_b0 );
or ( \7483_b1 , \6592_b1 , \6589_b1 );
not ( \6589_b1 , w_23810 );
and ( \7483_b0 , \6592_b0 , w_23811 );
and ( w_23810 , w_23811 , \6589_b0 );
or ( \7484_b1 , \7483_b1 , \6571_b1 );
not ( \6571_b1 , w_23812 );
and ( \7484_b0 , \7483_b0 , w_23813 );
and ( w_23812 , w_23813 , \6571_b0 );
buf ( \7485_b1 , \7483_b1 );
not ( \7485_b1 , w_23814 );
not ( \7485_b0 , w_23815 );
and ( w_23814 , w_23815 , \7483_b0 );
buf ( \7486_b1 , \6571_b1 );
not ( \7486_b1 , w_23816 );
not ( \7486_b0 , w_23817 );
and ( w_23816 , w_23817 , \6571_b0 );
or ( \7487_b1 , \7485_b1 , \7486_b1 );
not ( \7486_b1 , w_23818 );
and ( \7487_b0 , \7485_b0 , w_23819 );
and ( w_23818 , w_23819 , \7486_b0 );
or ( \7488_b1 , \7484_b1 , w_23821 );
not ( w_23821 , w_23822 );
and ( \7488_b0 , \7484_b0 , w_23823 );
and ( w_23822 ,  , w_23823 );
buf ( w_23821 , \7487_b1 );
not ( w_23821 , w_23824 );
not (  , w_23825 );
and ( w_23824 , w_23825 , \7487_b0 );
or ( \7489_b1 , \6597_b1 , w_23827 );
not ( w_23827 , w_23828 );
and ( \7489_b0 , \6597_b0 , w_23829 );
and ( w_23828 ,  , w_23829 );
buf ( w_23827 , \6471_b1 );
not ( w_23827 , w_23830 );
not (  , w_23831 );
and ( w_23830 , w_23831 , \6471_b0 );
buf ( \7490_b1 , \6567_b1 );
not ( \7490_b1 , w_23832 );
not ( \7490_b0 , w_23833 );
and ( w_23832 , w_23833 , \6567_b0 );
or ( \7491_b1 , \6570_b1 , w_23835 );
not ( w_23835 , w_23836 );
and ( \7491_b0 , \6570_b0 , w_23837 );
and ( w_23836 ,  , w_23837 );
buf ( w_23835 , \6515_b1 );
not ( w_23835 , w_23838 );
not (  , w_23839 );
and ( w_23838 , w_23839 , \6515_b0 );
buf ( \7492_b1 , \7491_b1 );
not ( \7492_b1 , w_23840 );
not ( \7492_b0 , w_23841 );
and ( w_23840 , w_23841 , \7491_b0 );
or ( \7493_b1 , \7490_b1 , w_23842 );
or ( \7493_b0 , \7490_b0 , \7492_b0 );
not ( \7492_b0 , w_23843 );
and ( w_23843 , w_23842 , \7492_b1 );
or ( \7494_b1 , \6567_b1 , w_23844 );
or ( \7494_b0 , \6567_b0 , \7491_b0 );
not ( \7491_b0 , w_23845 );
and ( w_23845 , w_23844 , \7491_b1 );
or ( \7495_b1 , \7493_b1 , w_23847 );
not ( w_23847 , w_23848 );
and ( \7495_b0 , \7493_b0 , w_23849 );
and ( w_23848 ,  , w_23849 );
buf ( w_23847 , \7494_b1 );
not ( w_23847 , w_23850 );
not (  , w_23851 );
and ( w_23850 , w_23851 , \7494_b0 );
or ( \7496_b1 , \6526_b1 , \6558_b1 );
xor ( \7496_b0 , \6526_b0 , w_23852 );
not ( w_23852 , w_23853 );
and ( w_23853 , \6558_b1 , \6558_b0 );
or ( \7497_b1 , \7496_b1 , \6564_b1 );
xor ( \7497_b0 , \7496_b0 , w_23854 );
not ( w_23854 , w_23855 );
and ( w_23855 , \6564_b1 , \6564_b0 );
or ( \7498_b1 , \6557_b1 , w_23857 );
not ( w_23857 , w_23858 );
and ( \7498_b0 , \6557_b0 , w_23859 );
and ( w_23858 ,  , w_23859 );
buf ( w_23857 , \6539_b1 );
not ( w_23857 , w_23860 );
not (  , w_23861 );
and ( w_23860 , w_23861 , \6539_b0 );
or ( \7499_b1 , \7498_b1 , \6552_b1 );
not ( \6552_b1 , w_23862 );
and ( \7499_b0 , \7498_b0 , w_23863 );
and ( w_23862 , w_23863 , \6552_b0 );
buf ( \7500_b1 , \7498_b1 );
not ( \7500_b1 , w_23864 );
not ( \7500_b0 , w_23865 );
and ( w_23864 , w_23865 , \7498_b0 );
or ( \7501_b1 , \7500_b1 , \6553_b1 );
not ( \6553_b1 , w_23866 );
and ( \7501_b0 , \7500_b0 , w_23867 );
and ( w_23866 , w_23867 , \6553_b0 );
or ( \7502_b1 , \7499_b1 , w_23869 );
not ( w_23869 , w_23870 );
and ( \7502_b0 , \7499_b0 , w_23871 );
and ( w_23870 ,  , w_23871 );
buf ( w_23869 , \7501_b1 );
not ( w_23869 , w_23872 );
not (  , w_23873 );
and ( w_23872 , w_23873 , \7501_b0 );
buf ( \7503_b1 , \6552_b1 );
not ( \7503_b1 , w_23874 );
not ( \7503_b0 , w_23875 );
and ( w_23874 , w_23875 , \6552_b0 );
or ( \7504_b1 , \6549_b1 , w_23877 );
not ( w_23877 , w_23878 );
and ( \7504_b0 , \6549_b0 , w_23879 );
and ( w_23878 ,  , w_23879 );
buf ( w_23877 , \6551_b1 );
not ( w_23877 , w_23880 );
not (  , w_23881 );
and ( w_23880 , w_23881 , \6551_b0 );
or ( \7505_b1 , \7503_b1 , w_23883 );
not ( w_23883 , w_23884 );
and ( \7505_b0 , \7503_b0 , w_23885 );
and ( w_23884 ,  , w_23885 );
buf ( w_23883 , \7504_b1 );
not ( w_23883 , w_23886 );
not (  , w_23887 );
and ( w_23886 , w_23887 , \7504_b0 );
buf ( \7506_b1 , \6550_b1 );
not ( \7506_b1 , w_23888 );
not ( \7506_b0 , w_23889 );
and ( w_23888 , w_23889 , \6550_b0 );
or ( \7507_b1 , \6593_b1 , w_23890 );
xor ( \7507_b0 , \6593_b0 , w_23892 );
not ( w_23892 , w_23893 );
and ( w_23893 , w_23890 , w_23891 );
buf ( w_23890 , \7489_b1 );
not ( w_23890 , w_23894 );
not ( w_23891 , w_23895 );
and ( w_23894 , w_23895 , \7489_b0 );
or ( \7508_b1 , \7328_b1 , w_23896 );
xor ( \7508_b0 , \7328_b0 , w_23898 );
not ( w_23898 , w_23899 );
and ( w_23899 , w_23896 , w_23897 );
buf ( w_23896 , \7419_b1 );
not ( w_23896 , w_23900 );
not ( w_23897 , w_23901 );
and ( w_23900 , w_23901 , \7419_b0 );
or ( \113_b1 , \111_b1 , w_23902 );
not ( w_23902 , w_23906 );
and ( \113_b0 , \111_b0 , w_23907 );
and ( w_23906 , w_23907 , w_23903 );
or ( w_23902 , \112_b1 , w_23904 );
not ( w_23904 , w_23908 );
and ( w_23903 , \112_b0 , w_23909 );
and ( w_23908 , w_23909 , w_23905 );
buf ( w_23904 , \b[5]_b1 );
not ( w_23904 , w_23910 );
not ( w_23905 , w_23911 );
and ( w_23910 , w_23911 , \b[5]_b0 );
or ( \159_b1 , \157_b1 , w_23912 );
not ( w_23912 , w_23916 );
and ( \159_b0 , \157_b0 , w_23917 );
and ( w_23916 , w_23917 , w_23913 );
or ( w_23912 , \158_b1 , w_23914 );
not ( w_23914 , w_23918 );
and ( w_23913 , \158_b0 , w_23919 );
and ( w_23918 , w_23919 , w_23915 );
buf ( w_23914 , \b[7]_b1 );
not ( w_23914 , w_23920 );
not ( w_23915 , w_23921 );
and ( w_23920 , w_23921 , \b[7]_b0 );
or ( \218_b1 , \216_b1 , w_23922 );
not ( w_23922 , w_23926 );
and ( \218_b0 , \216_b0 , w_23927 );
and ( w_23926 , w_23927 , w_23923 );
or ( w_23922 , \133_b1 , w_23924 );
not ( w_23924 , w_23928 );
and ( w_23923 , \133_b0 , w_23929 );
and ( w_23928 , w_23929 , w_23925 );
buf ( w_23924 , \217_b1 );
not ( w_23924 , w_23930 );
not ( w_23925 , w_23931 );
and ( w_23930 , w_23931 , \217_b0 );
or ( \220_b1 , \216_b1 , w_23932 );
not ( w_23932 , w_23936 );
and ( \220_b0 , \216_b0 , w_23937 );
and ( w_23936 , w_23937 , w_23933 );
or ( w_23932 , \133_b1 , w_23934 );
not ( w_23934 , w_23938 );
and ( w_23933 , \133_b0 , w_23939 );
and ( w_23938 , w_23939 , w_23935 );
buf ( w_23934 , \219_b1 );
not ( w_23934 , w_23940 );
not ( w_23935 , w_23941 );
and ( w_23940 , w_23941 , \219_b0 );
or ( \222_b1 , \218_b1 , w_23942 );
not ( w_23942 , w_23944 );
and ( \222_b0 , \218_b0 , w_23945 );
and ( w_23944 , w_23945 , w_23943 );
or ( w_23942 , \220_b1 , \221_b1 );
not ( \221_b1 , w_23946 );
and ( w_23943 , \220_b0 , w_23947 );
and ( w_23946 , w_23947 , \221_b0 );
or ( \282_b1 , \279_b1 , w_23948 );
not ( w_23948 , w_23952 );
and ( \282_b0 , \279_b0 , w_23953 );
and ( w_23952 , w_23953 , w_23949 );
or ( w_23948 , \b[3]_b1 , w_23950 );
not ( w_23950 , w_23954 );
and ( w_23949 , \b[3]_b0 , w_23955 );
and ( w_23954 , w_23955 , w_23951 );
buf ( w_23950 , \281_b1 );
not ( w_23950 , w_23956 );
not ( w_23951 , w_23957 );
and ( w_23956 , w_23957 , \281_b0 );
or ( \412_b1 , \410_b1 , w_23958 );
not ( w_23958 , w_23960 );
and ( \412_b0 , \410_b0 , w_23961 );
and ( w_23960 , w_23961 , w_23959 );
or ( w_23958 , \411_b1 , \b[9]_b1 );
not ( \b[9]_b1 , w_23962 );
and ( w_23959 , \411_b0 , w_23963 );
and ( w_23962 , w_23963 , \b[9]_b0 );
or ( \533_b1 , \347_b1 , w_23964 );
not ( w_23964 , w_23968 );
and ( \533_b0 , \347_b0 , w_23969 );
and ( w_23968 , w_23969 , w_23965 );
or ( w_23964 , \471_b1 , w_23966 );
not ( w_23966 , w_23970 );
and ( w_23965 , \471_b0 , w_23971 );
and ( w_23970 , w_23971 , w_23967 );
buf ( w_23966 , \532_b1 );
not ( w_23966 , w_23972 );
not ( w_23967 , w_23973 );
and ( w_23972 , w_23973 , \532_b0 );
or ( \543_b1 , \541_b1 , w_23974 );
not ( w_23974 , w_23978 );
and ( \543_b0 , \541_b0 , w_23979 );
and ( w_23978 , w_23979 , w_23975 );
or ( w_23974 , \542_b1 , w_23976 );
not ( w_23976 , w_23980 );
and ( w_23975 , \542_b0 , w_23981 );
and ( w_23980 , w_23981 , w_23977 );
buf ( w_23976 , \532_b1 );
not ( w_23976 , w_23982 );
not ( w_23977 , w_23983 );
and ( w_23982 , w_23983 , \532_b0 );
or ( \547_b1 , \533_b1 , w_23984 );
not ( w_23984 , w_23988 );
and ( \547_b0 , \533_b0 , w_23989 );
and ( w_23988 , w_23989 , w_23985 );
or ( w_23984 , \543_b1 , w_23986 );
not ( w_23986 , w_23990 );
and ( w_23985 , \543_b0 , w_23991 );
and ( w_23990 , w_23991 , w_23987 );
buf ( w_23986 , \546_b1 );
not ( w_23986 , w_23992 );
not ( w_23987 , w_23993 );
and ( w_23992 , w_23993 , \546_b0 );
or ( \566_b1 , \564_b1 , w_23994 );
not ( w_23994 , w_23998 );
and ( \566_b0 , \564_b0 , w_23999 );
and ( w_23998 , w_23999 , w_23995 );
or ( w_23994 , \565_b1 , w_23996 );
not ( w_23996 , w_24000 );
and ( w_23995 , \565_b0 , w_24001 );
and ( w_24000 , w_24001 , w_23997 );
buf ( w_23996 , \b[11]_b1 );
not ( w_23996 , w_24002 );
not ( w_23997 , w_24003 );
and ( w_24002 , w_24003 , \b[11]_b0 );
or ( \671_b1 , \a[8]_b1 , w_24010 );
or ( \671_b0 , \a[8]_b0 , w_24005 );
not ( w_24005 , w_24011 );
and ( w_24011 , w_24010 , w_24004 );
or ( w_24004 , \a[7]_b1 , w_24012 );
or ( w_24005 , \a[7]_b0 , w_24007 );
not ( w_24007 , w_24013 );
and ( w_24013 , w_24012 , w_24006 );
or ( w_24006 , \a[6]_b1 , w_24014 );
or ( w_24007 , \a[6]_b0 , w_24009 );
not ( w_24009 , w_24015 );
and ( w_24015 , w_24014 , w_24008 );
buf ( w_24008 , \a[5]_b1 );
not ( w_24008 , w_24016 );
not ( w_24009 , w_24017 );
and ( w_24016 , w_24017 , \a[5]_b0 );
or ( \675_b1 , \671_b1 , w_24018 );
not ( w_24018 , w_24024 );
and ( \675_b0 , \671_b0 , w_24025 );
and ( w_24024 , w_24025 , w_24019 );
or ( w_24018 , \672_b1 , w_24020 );
not ( w_24020 , w_24026 );
and ( w_24019 , \672_b0 , w_24027 );
and ( w_24026 , w_24027 , w_24021 );
or ( w_24020 , \673_b1 , w_24022 );
not ( w_24022 , w_24028 );
and ( w_24021 , \673_b0 , w_24029 );
and ( w_24028 , w_24029 , w_24023 );
buf ( w_24022 , \674_b1 );
not ( w_24022 , w_24030 );
not ( w_24023 , w_24031 );
and ( w_24030 , w_24031 , \674_b0 );
or ( \676_b1 , \a[15]_b1 , w_24036 );
or ( \676_b0 , \a[15]_b0 , w_24033 );
not ( w_24033 , w_24037 );
and ( w_24037 , w_24036 , w_24032 );
or ( w_24032 , \a[4]_b1 , w_24038 );
or ( w_24033 , \a[4]_b0 , w_24035 );
not ( w_24035 , w_24039 );
and ( w_24039 , w_24038 , w_24034 );
or ( w_24034 , \d[8]_b1 , w_24040 );
or ( w_24035 , \d[8]_b0 , \d[7]_b0 );
not ( \d[7]_b0 , w_24041 );
and ( w_24041 , w_24040 , \d[7]_b1 );
or ( \677_b1 , \d[6]_b1 , w_24046 );
or ( \677_b0 , \d[6]_b0 , w_24043 );
not ( w_24043 , w_24047 );
and ( w_24047 , w_24046 , w_24042 );
or ( w_24042 , \d[5]_b1 , w_24048 );
or ( w_24043 , \d[5]_b0 , w_24045 );
not ( w_24045 , w_24049 );
and ( w_24049 , w_24048 , w_24044 );
or ( w_24044 , \d[15]_b1 , w_24050 );
or ( w_24045 , \d[15]_b0 , \d[4]_b0 );
not ( \d[4]_b0 , w_24051 );
and ( w_24051 , w_24050 , \d[4]_b1 );
or ( \678_b1 , \675_b1 , w_24056 );
or ( \678_b0 , \675_b0 , w_24053 );
not ( w_24053 , w_24057 );
and ( w_24057 , w_24056 , w_24052 );
or ( w_24052 , \676_b1 , w_24058 );
or ( w_24053 , \676_b0 , w_24055 );
not ( w_24055 , w_24059 );
and ( w_24059 , w_24058 , w_24054 );
buf ( w_24054 , \677_b1 );
not ( w_24054 , w_24060 );
not ( w_24055 , w_24061 );
and ( w_24060 , w_24061 , \677_b0 );
or ( \682_b1 , \679_b1 , w_24066 );
or ( \682_b0 , \679_b0 , w_24063 );
not ( w_24063 , w_24067 );
and ( w_24067 , w_24066 , w_24062 );
or ( w_24062 , \680_b1 , w_24068 );
or ( w_24063 , \680_b0 , w_24065 );
not ( w_24065 , w_24069 );
and ( w_24069 , w_24068 , w_24064 );
buf ( w_24064 , \681_b1 );
not ( w_24064 , w_24070 );
not ( w_24065 , w_24071 );
and ( w_24070 , w_24071 , \681_b0 );
or ( \685_b1 , \678_b1 , w_24072 );
not ( w_24072 , w_24078 );
and ( \685_b0 , \678_b0 , w_24079 );
and ( w_24078 , w_24079 , w_24073 );
or ( w_24072 , \682_b1 , w_24074 );
not ( w_24074 , w_24080 );
and ( w_24073 , \682_b0 , w_24081 );
and ( w_24080 , w_24081 , w_24075 );
or ( w_24074 , \683_b1 , w_24076 );
not ( w_24076 , w_24082 );
and ( w_24075 , \683_b0 , w_24083 );
and ( w_24082 , w_24083 , w_24077 );
buf ( w_24076 , \684_b1 );
not ( w_24076 , w_24084 );
not ( w_24077 , w_24085 );
and ( w_24084 , w_24085 , \684_b0 );
or ( \690_b1 , \686_b1 , w_24088 );
or ( \690_b0 , \686_b0 , w_24087 );
not ( w_24087 , w_24089 );
and ( w_24089 , w_24088 , w_24086 );
or ( w_24086 , \689_b1 , w_24090 );
or ( w_24087 , \689_b0 , \d[13]_b0 );
not ( \d[13]_b0 , w_24091 );
and ( w_24091 , w_24090 , \d[13]_b1 );
or ( \691_b1 , \670_b1 , w_24098 );
or ( \691_b0 , \670_b0 , w_24093 );
not ( w_24093 , w_24099 );
and ( w_24099 , w_24098 , w_24092 );
or ( w_24092 , \685_b1 , w_24100 );
or ( w_24093 , \685_b0 , w_24095 );
not ( w_24095 , w_24101 );
and ( w_24101 , w_24100 , w_24094 );
or ( w_24094 , \690_b1 , w_24102 );
or ( w_24095 , \690_b0 , w_24097 );
not ( w_24097 , w_24103 );
and ( w_24103 , w_24102 , w_24096 );
buf ( w_24096 , \a[13]_b1 );
not ( w_24096 , w_24104 );
not ( w_24097 , w_24105 );
and ( w_24104 , w_24105 , \a[13]_b0 );
or ( \720_b1 , \716_b1 , w_24106 );
not ( w_24106 , w_24110 );
and ( \720_b0 , \716_b0 , w_24111 );
and ( w_24110 , w_24111 , w_24107 );
or ( w_24106 , \717_b1 , w_24108 );
not ( w_24108 , w_24112 );
and ( w_24107 , \717_b0 , w_24113 );
and ( w_24112 , w_24113 , w_24109 );
buf ( w_24108 , \719_b1 );
not ( w_24108 , w_24114 );
not ( w_24109 , w_24115 );
and ( w_24114 , w_24115 , \719_b0 );
or ( \723_b1 , \720_b1 , w_24116 );
not ( w_24116 , w_24120 );
and ( \723_b0 , \720_b0 , w_24121 );
and ( w_24120 , w_24121 , w_24117 );
or ( w_24116 , \721_b1 , w_24118 );
not ( w_24118 , w_24122 );
and ( w_24117 , \721_b0 , w_24123 );
and ( w_24122 , w_24123 , w_24119 );
buf ( w_24118 , \722_b1 );
not ( w_24118 , w_24124 );
not ( w_24119 , w_24125 );
and ( w_24124 , w_24125 , \722_b0 );
or ( \745_b1 , \741_b1 , w_24126 );
not ( w_24126 , w_24132 );
and ( \745_b0 , \741_b0 , w_24133 );
and ( w_24132 , w_24133 , w_24127 );
or ( w_24126 , \736_b1 , w_24128 );
not ( w_24128 , w_24134 );
and ( w_24127 , \736_b0 , w_24135 );
and ( w_24134 , w_24135 , w_24129 );
or ( w_24128 , \742_b1 , w_24130 );
not ( w_24130 , w_24136 );
and ( w_24129 , \742_b0 , w_24137 );
and ( w_24136 , w_24137 , w_24131 );
buf ( w_24130 , \744_b1 );
not ( w_24130 , w_24138 );
not ( w_24131 , w_24139 );
and ( w_24138 , w_24139 , \744_b0 );
or ( \762_b1 , \747_b1 , w_24140 );
not ( w_24140 , w_24142 );
and ( \762_b0 , \747_b0 , w_24143 );
and ( w_24142 , w_24143 , w_24141 );
or ( w_24140 , \754_b1 , \761_b1 );
not ( \761_b1 , w_24144 );
and ( w_24141 , \754_b0 , w_24145 );
and ( w_24144 , w_24145 , \761_b0 );
or ( \786_b1 , \778_b1 , w_24146 );
not ( w_24146 , w_24150 );
and ( \786_b0 , \778_b0 , w_24151 );
and ( w_24150 , w_24151 , w_24147 );
or ( w_24146 , \784_b1 , w_24148 );
not ( w_24148 , w_24152 );
and ( w_24147 , \784_b0 , w_24153 );
and ( w_24152 , w_24153 , w_24149 );
buf ( w_24148 , \785_b1 );
not ( w_24148 , w_24154 );
not ( w_24149 , w_24155 );
and ( w_24154 , w_24155 , \785_b0 );
or ( \805_b1 , \801_b1 , w_24156 );
not ( w_24156 , w_24160 );
and ( \805_b0 , \801_b0 , w_24161 );
and ( w_24160 , w_24161 , w_24157 );
or ( w_24156 , \802_b1 , w_24158 );
not ( w_24158 , w_24162 );
and ( w_24157 , \802_b0 , w_24163 );
and ( w_24162 , w_24163 , w_24159 );
buf ( w_24158 , \804_b1 );
not ( w_24158 , w_24164 );
not ( w_24159 , w_24165 );
and ( w_24164 , w_24165 , \804_b0 );
or ( \808_b1 , \805_b1 , w_24166 );
not ( w_24166 , w_24170 );
and ( \808_b0 , \805_b0 , w_24171 );
and ( w_24170 , w_24171 , w_24167 );
or ( w_24166 , \806_b1 , w_24168 );
not ( w_24168 , w_24172 );
and ( w_24167 , \806_b0 , w_24173 );
and ( w_24172 , w_24173 , w_24169 );
buf ( w_24168 , \807_b1 );
not ( w_24168 , w_24174 );
not ( w_24169 , w_24175 );
and ( w_24174 , w_24175 , \807_b0 );
or ( \830_b1 , \826_b1 , w_24176 );
not ( w_24176 , w_24182 );
and ( \830_b0 , \826_b0 , w_24183 );
and ( w_24182 , w_24183 , w_24177 );
or ( w_24176 , \821_b1 , w_24178 );
not ( w_24178 , w_24184 );
and ( w_24177 , \821_b0 , w_24185 );
and ( w_24184 , w_24185 , w_24179 );
or ( w_24178 , \827_b1 , w_24180 );
not ( w_24180 , w_24186 );
and ( w_24179 , \827_b0 , w_24187 );
and ( w_24186 , w_24187 , w_24181 );
buf ( w_24180 , \829_b1 );
not ( w_24180 , w_24188 );
not ( w_24181 , w_24189 );
and ( w_24188 , w_24189 , \829_b0 );
or ( \847_b1 , \832_b1 , w_24190 );
not ( w_24190 , w_24192 );
and ( \847_b0 , \832_b0 , w_24193 );
and ( w_24192 , w_24193 , w_24191 );
or ( w_24190 , \839_b1 , \846_b1 );
not ( \846_b1 , w_24194 );
and ( w_24191 , \839_b0 , w_24195 );
and ( w_24194 , w_24195 , \846_b0 );
or ( \871_b1 , \863_b1 , w_24196 );
not ( w_24196 , w_24200 );
and ( \871_b0 , \863_b0 , w_24201 );
and ( w_24200 , w_24201 , w_24197 );
or ( w_24196 , \869_b1 , w_24198 );
not ( w_24198 , w_24202 );
and ( w_24197 , \869_b0 , w_24203 );
and ( w_24202 , w_24203 , w_24199 );
buf ( w_24198 , \870_b1 );
not ( w_24198 , w_24204 );
not ( w_24199 , w_24205 );
and ( w_24204 , w_24205 , \870_b0 );
or ( \956_b1 , \954_b1 , w_24206 );
not ( w_24206 , w_24208 );
and ( \956_b0 , \954_b0 , w_24209 );
and ( w_24208 , w_24209 , w_24207 );
or ( w_24206 , \955_b1 , \d[11]_b1 );
not ( \d[11]_b1 , w_24210 );
and ( w_24207 , \955_b0 , w_24211 );
and ( w_24210 , w_24211 , \d[11]_b0 );
or ( \974_b1 , \972_b1 , w_24212 );
not ( w_24212 , w_24216 );
and ( \974_b0 , \972_b0 , w_24217 );
and ( w_24216 , w_24217 , w_24213 );
or ( w_24212 , \973_b1 , w_24214 );
not ( w_24214 , w_24218 );
and ( w_24213 , \973_b0 , w_24219 );
and ( w_24218 , w_24219 , w_24215 );
buf ( w_24214 , \d[9]_b1 );
not ( w_24214 , w_24220 );
not ( w_24215 , w_24221 );
and ( w_24220 , w_24221 , \d[9]_b0 );
or ( \1026_b1 , \1022_b1 , w_24222 );
not ( w_24222 , w_24224 );
and ( \1026_b0 , \1022_b0 , w_24225 );
and ( w_24224 , w_24225 , w_24223 );
or ( w_24222 , \1024_b1 , \1025_b1 );
not ( \1025_b1 , w_24226 );
and ( w_24223 , \1024_b0 , w_24227 );
and ( w_24226 , w_24227 , \1025_b0 );
or ( \1109_b1 , \1024_b1 , w_24228 );
not ( w_24228 , w_24230 );
and ( \1109_b0 , \1024_b0 , w_24231 );
and ( w_24230 , w_24231 , w_24229 );
or ( w_24228 , \1022_b1 , \1025_b1 );
not ( \1025_b1 , w_24232 );
and ( w_24229 , \1022_b0 , w_24233 );
and ( w_24232 , w_24233 , \1025_b0 );
or ( \1181_b1 , \1179_b1 , w_24234 );
not ( w_24234 , w_24236 );
and ( \1181_b0 , \1179_b0 , w_24237 );
and ( w_24236 , w_24237 , w_24235 );
or ( w_24234 , \1180_b1 , \d[7]_b1 );
not ( \d[7]_b1 , w_24238 );
and ( w_24235 , \1180_b0 , w_24239 );
and ( w_24238 , w_24239 , \d[7]_b0 );
or ( \1310_b1 , \1161_b1 , w_24240 );
not ( w_24240 , w_24242 );
and ( \1310_b0 , \1161_b0 , w_24243 );
and ( w_24242 , w_24243 , w_24241 );
or ( w_24240 , \1214_b1 , \1309_b1 );
not ( \1309_b1 , w_24244 );
and ( w_24241 , \1214_b0 , w_24245 );
and ( w_24244 , w_24245 , \1309_b0 );
or ( \1396_b1 , \1394_b1 , w_24246 );
not ( w_24246 , w_24250 );
and ( \1396_b0 , \1394_b0 , w_24251 );
and ( w_24250 , w_24251 , w_24247 );
or ( w_24246 , \1395_b1 , w_24248 );
not ( w_24248 , w_24252 );
and ( w_24247 , \1395_b0 , w_24253 );
and ( w_24252 , w_24253 , w_24249 );
buf ( w_24248 , \d[5]_b1 );
not ( w_24248 , w_24254 );
not ( w_24249 , w_24255 );
and ( w_24254 , w_24255 , \d[5]_b0 );
or ( \1474_b1 , \1472_b1 , w_24256 );
not ( w_24256 , w_24260 );
and ( \1474_b0 , \1472_b0 , w_24261 );
and ( w_24260 , w_24261 , w_24257 );
or ( w_24256 , \1473_b1 , w_24258 );
not ( w_24258 , w_24262 );
and ( w_24257 , \1473_b0 , w_24263 );
and ( w_24262 , w_24263 , w_24259 );
buf ( w_24258 , \d[3]_b1 );
not ( w_24258 , w_24264 );
not ( w_24259 , w_24265 );
and ( w_24264 , w_24265 , \d[3]_b0 );
or ( \1529_b1 , \1310_b1 , w_24266 );
not ( w_24266 , w_24270 );
and ( \1529_b0 , \1310_b0 , w_24271 );
and ( w_24270 , w_24271 , w_24267 );
or ( w_24266 , \1388_b1 , w_24268 );
not ( w_24268 , w_24272 );
and ( w_24267 , \1388_b0 , w_24273 );
and ( w_24272 , w_24273 , w_24269 );
buf ( w_24268 , \1528_b1 );
not ( w_24268 , w_24274 );
not ( w_24269 , w_24275 );
and ( w_24274 , w_24275 , \1528_b0 );
or ( \1542_b1 , \1540_b1 , w_24276 );
not ( w_24276 , w_24282 );
and ( \1542_b0 , \1540_b0 , w_24283 );
and ( w_24282 , w_24283 , w_24277 );
or ( w_24276 , \1541_b1 , w_24278 );
not ( w_24278 , w_24284 );
and ( w_24277 , \1541_b0 , w_24285 );
and ( w_24284 , w_24285 , w_24279 );
or ( w_24278 , \1214_b1 , w_24280 );
not ( w_24280 , w_24286 );
and ( w_24279 , \1214_b0 , w_24287 );
and ( w_24286 , w_24287 , w_24281 );
buf ( w_24280 , \1388_b1 );
not ( w_24280 , w_24288 );
not ( w_24281 , w_24289 );
and ( w_24288 , w_24289 , \1388_b0 );
or ( \1544_b1 , \1529_b1 , w_24290 );
not ( w_24290 , w_24296 );
and ( \1544_b0 , \1529_b0 , w_24297 );
and ( w_24296 , w_24297 , w_24291 );
or ( w_24290 , \1531_b1 , w_24292 );
not ( w_24292 , w_24298 );
and ( w_24291 , \1531_b0 , w_24299 );
and ( w_24298 , w_24299 , w_24293 );
or ( w_24292 , \1542_b1 , w_24294 );
not ( w_24294 , w_24300 );
and ( w_24293 , \1542_b0 , w_24301 );
and ( w_24300 , w_24301 , w_24295 );
buf ( w_24294 , \1543_b1 );
not ( w_24294 , w_24302 );
not ( w_24295 , w_24303 );
and ( w_24302 , w_24303 , \1543_b0 );
or ( \1555_b1 , \1553_b1 , w_24304 );
not ( w_24304 , w_24308 );
and ( \1555_b0 , \1553_b0 , w_24309 );
and ( w_24308 , w_24309 , w_24305 );
or ( w_24304 , \1554_b1 , w_24306 );
not ( w_24306 , w_24310 );
and ( w_24305 , \1554_b0 , w_24311 );
and ( w_24310 , w_24311 , w_24307 );
buf ( w_24306 , \d[13]_b1 );
not ( w_24306 , w_24312 );
not ( w_24307 , w_24313 );
and ( w_24312 , w_24313 , \d[13]_b0 );
or ( \1698_b1 , \1696_b1 , w_24314 );
not ( w_24314 , w_24316 );
and ( \1698_b0 , \1696_b0 , w_24317 );
and ( w_24316 , w_24317 , w_24315 );
or ( w_24314 , \1697_b1 , \c[11]_b1 );
not ( \c[11]_b1 , w_24318 );
and ( w_24315 , \1697_b0 , w_24319 );
and ( w_24318 , w_24319 , \c[11]_b0 );
or ( \1717_b1 , \1715_b1 , w_24320 );
not ( w_24320 , w_24324 );
and ( \1717_b0 , \1715_b0 , w_24325 );
and ( w_24324 , w_24325 , w_24321 );
or ( w_24320 , \1716_b1 , w_24322 );
not ( w_24322 , w_24326 );
and ( w_24321 , \1716_b0 , w_24327 );
and ( w_24326 , w_24327 , w_24323 );
buf ( w_24322 , \c[9]_b1 );
not ( w_24322 , w_24328 );
not ( w_24323 , w_24329 );
and ( w_24328 , w_24329 , \c[9]_b0 );
or ( \1770_b1 , \1767_b1 , w_24330 );
not ( w_24330 , w_24332 );
and ( \1770_b0 , \1767_b0 , w_24333 );
and ( w_24332 , w_24333 , w_24331 );
or ( w_24330 , \1768_b1 , \1769_b1 );
not ( \1769_b1 , w_24334 );
and ( w_24331 , \1768_b0 , w_24335 );
and ( w_24334 , w_24335 , \1769_b0 );
or ( \1921_b1 , \1919_b1 , w_24336 );
not ( w_24336 , w_24338 );
and ( \1921_b0 , \1919_b0 , w_24339 );
and ( w_24338 , w_24339 , w_24337 );
or ( w_24336 , \1920_b1 , \c[7]_b1 );
not ( \c[7]_b1 , w_24340 );
and ( w_24337 , \1920_b0 , w_24341 );
and ( w_24340 , w_24341 , \c[7]_b0 );
or ( \2050_b1 , \1901_b1 , w_24342 );
not ( w_24342 , w_24344 );
and ( \2050_b0 , \1901_b0 , w_24345 );
and ( w_24344 , w_24345 , w_24343 );
or ( w_24342 , \1954_b1 , \2049_b1 );
not ( \2049_b1 , w_24346 );
and ( w_24343 , \1954_b0 , w_24347 );
and ( w_24346 , w_24347 , \2049_b0 );
or ( \2137_b1 , \c[5]_b1 , w_24348 );
not ( w_24348 , w_24352 );
and ( \2137_b0 , \c[5]_b0 , w_24353 );
and ( w_24352 , w_24353 , w_24349 );
or ( w_24348 , \2134_b1 , w_24350 );
not ( w_24350 , w_24354 );
and ( w_24349 , \2134_b0 , w_24355 );
and ( w_24354 , w_24355 , w_24351 );
buf ( w_24350 , \2136_b1 );
not ( w_24350 , w_24356 );
not ( w_24351 , w_24357 );
and ( w_24356 , w_24357 , \2136_b0 );
or ( \2190_b1 , \2188_b1 , w_24358 );
not ( w_24358 , w_24362 );
and ( \2190_b0 , \2188_b0 , w_24363 );
and ( w_24362 , w_24363 , w_24359 );
or ( w_24358 , \2189_b1 , w_24360 );
not ( w_24360 , w_24364 );
and ( w_24359 , \2189_b0 , w_24365 );
and ( w_24364 , w_24365 , w_24361 );
buf ( w_24360 , \c[3]_b1 );
not ( w_24360 , w_24366 );
not ( w_24361 , w_24367 );
and ( w_24366 , w_24367 , \c[3]_b0 );
or ( \2272_b1 , \2050_b1 , w_24368 );
not ( w_24368 , w_24372 );
and ( \2272_b0 , \2050_b0 , w_24373 );
and ( w_24372 , w_24373 , w_24369 );
or ( w_24368 , \2129_b1 , w_24370 );
not ( w_24370 , w_24374 );
and ( w_24369 , \2129_b0 , w_24375 );
and ( w_24374 , w_24375 , w_24371 );
buf ( w_24370 , \2271_b1 );
not ( w_24370 , w_24376 );
not ( w_24371 , w_24377 );
and ( w_24376 , w_24377 , \2271_b0 );
or ( \2286_b1 , \2283_b1 , w_24378 );
not ( w_24378 , w_24384 );
and ( \2286_b0 , \2283_b0 , w_24385 );
and ( w_24384 , w_24385 , w_24379 );
or ( w_24378 , \2284_b1 , w_24380 );
not ( w_24380 , w_24386 );
and ( w_24379 , \2284_b0 , w_24387 );
and ( w_24386 , w_24387 , w_24381 );
or ( w_24380 , \2285_b1 , w_24382 );
not ( w_24382 , w_24388 );
and ( w_24381 , \2285_b0 , w_24389 );
and ( w_24388 , w_24389 , w_24383 );
buf ( w_24382 , \2129_b1 );
not ( w_24382 , w_24390 );
not ( w_24383 , w_24391 );
and ( w_24390 , w_24391 , \2129_b0 );
or ( \2289_b1 , \2272_b1 , w_24392 );
not ( w_24392 , w_24398 );
and ( \2289_b0 , \2272_b0 , w_24399 );
and ( w_24398 , w_24399 , w_24393 );
or ( w_24392 , \2274_b1 , w_24394 );
not ( w_24394 , w_24400 );
and ( w_24393 , \2274_b0 , w_24401 );
and ( w_24400 , w_24401 , w_24395 );
or ( w_24394 , \2286_b1 , w_24396 );
not ( w_24396 , w_24402 );
and ( w_24395 , \2286_b0 , w_24403 );
and ( w_24402 , w_24403 , w_24397 );
buf ( w_24396 , \2288_b1 );
not ( w_24396 , w_24404 );
not ( w_24397 , w_24405 );
and ( w_24404 , w_24405 , \2288_b0 );
or ( \2300_b1 , \2298_b1 , w_24406 );
not ( w_24406 , w_24410 );
and ( \2300_b0 , \2298_b0 , w_24411 );
and ( w_24410 , w_24411 , w_24407 );
or ( w_24406 , \2299_b1 , w_24408 );
not ( w_24408 , w_24412 );
and ( w_24407 , \2299_b0 , w_24413 );
and ( w_24412 , w_24413 , w_24409 );
buf ( w_24408 , \c[13]_b1 );
not ( w_24408 , w_24414 );
not ( w_24409 , w_24415 );
and ( w_24414 , w_24415 , \c[13]_b0 );
or ( \2433_b1 , \2432_b1 , w_24416 );
not ( w_24416 , w_24420 );
and ( \2433_b0 , \2432_b0 , w_24421 );
and ( w_24420 , w_24421 , w_24417 );
or ( w_24416 , \747_b1 , w_24418 );
not ( w_24418 , w_24422 );
and ( w_24417 , \747_b0 , w_24423 );
and ( w_24422 , w_24423 , w_24419 );
buf ( w_24418 , \754_b1 );
not ( w_24418 , w_24424 );
not ( w_24419 , w_24425 );
and ( w_24424 , w_24425 , \754_b0 );
or ( \2434_b1 , \2431_b1 , w_24426 );
not ( w_24426 , w_24430 );
and ( \2434_b0 , \2431_b0 , w_24431 );
and ( w_24430 , w_24431 , w_24427 );
or ( w_24426 , \2433_b1 , w_24428 );
not ( w_24428 , w_24432 );
and ( w_24427 , \2433_b0 , w_24433 );
and ( w_24432 , w_24433 , w_24429 );
buf ( w_24428 , \779_b1 );
not ( w_24428 , w_24434 );
not ( w_24429 , w_24435 );
and ( w_24434 , w_24435 , \779_b0 );
or ( \2447_b1 , \2446_b1 , w_24436 );
not ( w_24436 , w_24440 );
and ( \2447_b0 , \2446_b0 , w_24441 );
and ( w_24440 , w_24441 , w_24437 );
or ( w_24436 , \832_b1 , w_24438 );
not ( w_24438 , w_24442 );
and ( w_24437 , \832_b0 , w_24443 );
and ( w_24442 , w_24443 , w_24439 );
buf ( w_24438 , \839_b1 );
not ( w_24438 , w_24444 );
not ( w_24439 , w_24445 );
and ( w_24444 , w_24445 , \839_b0 );
or ( \2448_b1 , \2445_b1 , w_24446 );
not ( w_24446 , w_24450 );
and ( \2448_b0 , \2445_b0 , w_24451 );
and ( w_24450 , w_24451 , w_24447 );
or ( w_24446 , \2447_b1 , w_24448 );
not ( w_24448 , w_24452 );
and ( w_24447 , \2447_b0 , w_24453 );
and ( w_24452 , w_24453 , w_24449 );
buf ( w_24448 , \864_b1 );
not ( w_24448 , w_24454 );
not ( w_24449 , w_24455 );
and ( w_24454 , w_24455 , \864_b0 );
or ( \2477_b1 , \1669_b1 , w_24456 );
not ( w_24456 , w_24462 );
and ( \2477_b0 , \1669_b0 , w_24463 );
and ( w_24462 , w_24463 , w_24457 );
or ( w_24456 , \2414_b1 , w_24458 );
not ( w_24458 , w_24464 );
and ( w_24457 , \2414_b0 , w_24465 );
and ( w_24464 , w_24465 , w_24459 );
or ( w_24458 , \2465_b1 , w_24460 );
not ( w_24460 , w_24466 );
and ( w_24459 , \2465_b0 , w_24467 );
and ( w_24466 , w_24467 , w_24461 );
buf ( w_24460 , \2476_b1 );
not ( w_24460 , w_24468 );
not ( w_24461 , w_24469 );
and ( w_24468 , w_24469 , \2476_b0 );
or ( \2584_b1 , \2129_b1 , w_24470 );
not ( w_24470 , w_24472 );
and ( \2584_b0 , \2129_b0 , w_24473 );
and ( w_24472 , w_24473 , w_24471 );
or ( w_24470 , \2403_b1 , \1901_b1 );
not ( \1901_b1 , w_24474 );
and ( w_24471 , \2403_b0 , w_24475 );
and ( w_24474 , w_24475 , \1901_b0 );
or ( \2621_b1 , \747_b1 , w_24476 );
not ( w_24476 , w_24478 );
and ( \2621_b0 , \747_b0 , w_24479 );
and ( w_24478 , w_24479 , w_24477 );
or ( w_24476 , \754_b1 , \759_b1 );
not ( \759_b1 , w_24480 );
and ( w_24477 , \754_b0 , w_24481 );
and ( w_24480 , w_24481 , \759_b0 );
or ( \2636_b1 , \832_b1 , w_24482 );
not ( w_24482 , w_24484 );
and ( \2636_b0 , \832_b0 , w_24485 );
and ( w_24484 , w_24485 , w_24483 );
or ( w_24482 , \839_b1 , \844_b1 );
not ( \844_b1 , w_24486 );
and ( w_24483 , \839_b0 , w_24487 );
and ( w_24486 , w_24487 , \844_b0 );
or ( \2766_b1 , \1388_b1 , w_24488 );
not ( w_24488 , w_24490 );
and ( \2766_b0 , \1388_b0 , w_24491 );
and ( w_24490 , w_24491 , w_24489 );
or ( w_24488 , \1657_b1 , \1161_b1 );
not ( \1161_b1 , w_24492 );
and ( w_24489 , \1657_b0 , w_24493 );
and ( w_24492 , w_24493 , \1161_b0 );
or ( \2790_b1 , \2603_b1 , w_24494 );
not ( w_24494 , w_24500 );
and ( \2790_b0 , \2603_b0 , w_24501 );
and ( w_24500 , w_24501 , w_24495 );
or ( w_24494 , \2657_b1 , w_24496 );
not ( w_24496 , w_24502 );
and ( w_24495 , \2657_b0 , w_24503 );
and ( w_24502 , w_24503 , w_24497 );
or ( w_24496 , \2788_b1 , w_24498 );
not ( w_24498 , w_24504 );
and ( w_24497 , \2788_b0 , w_24505 );
and ( w_24504 , w_24505 , w_24499 );
buf ( w_24498 , \2789_b1 );
not ( w_24498 , w_24506 );
not ( w_24499 , w_24507 );
and ( w_24506 , w_24507 , \2789_b0 );
or ( \2803_b1 , \747_b1 , w_24508 );
not ( w_24508 , w_24510 );
and ( \2803_b0 , \747_b0 , w_24511 );
and ( w_24510 , w_24511 , w_24509 );
or ( w_24508 , \753_b1 , \2802_b1 );
not ( \2802_b1 , w_24512 );
and ( w_24509 , \753_b0 , w_24513 );
and ( w_24512 , w_24513 , \2802_b0 );
or ( \2819_b1 , \832_b1 , w_24514 );
not ( w_24514 , w_24516 );
and ( \2819_b0 , \832_b0 , w_24517 );
and ( w_24516 , w_24517 , w_24515 );
or ( w_24514 , \838_b1 , \2818_b1 );
not ( \2818_b1 , w_24518 );
and ( w_24515 , \838_b0 , w_24519 );
and ( w_24518 , w_24519 , \2818_b0 );
or ( \2876_b1 , \2841_b1 , w_24520 );
not ( w_24520 , w_24526 );
and ( \2876_b0 , \2841_b0 , w_24527 );
and ( w_24526 , w_24527 , w_24521 );
or ( w_24520 , \2856_b1 , w_24522 );
not ( w_24522 , w_24528 );
and ( w_24521 , \2856_b0 , w_24529 );
and ( w_24528 , w_24529 , w_24523 );
or ( w_24522 , \2860_b1 , w_24524 );
not ( w_24524 , w_24530 );
and ( w_24523 , \2860_b0 , w_24531 );
and ( w_24530 , w_24531 , w_24525 );
buf ( w_24524 , \2875_b1 );
not ( w_24524 , w_24532 );
not ( w_24525 , w_24533 );
and ( w_24532 , w_24533 , \2875_b0 );
or ( \2944_b1 , \2884_b1 , w_24534 );
not ( w_24534 , w_24538 );
and ( \2944_b0 , \2884_b0 , w_24539 );
and ( w_24538 , w_24539 , w_24535 );
or ( w_24534 , \2885_b1 , w_24536 );
not ( w_24536 , w_24540 );
and ( w_24535 , \2885_b0 , w_24541 );
and ( w_24540 , w_24541 , w_24537 );
buf ( w_24536 , \2943_b1 );
not ( w_24536 , w_24542 );
not ( w_24537 , w_24543 );
and ( w_24542 , w_24543 , \2943_b0 );
or ( \3016_b1 , \2948_b1 , w_24544 );
not ( w_24544 , w_24550 );
and ( \3016_b0 , \2948_b0 , w_24551 );
and ( w_24550 , w_24551 , w_24545 );
or ( w_24544 , \3011_b1 , w_24546 );
not ( w_24546 , w_24552 );
and ( w_24545 , \3011_b0 , w_24553 );
and ( w_24552 , w_24553 , w_24547 );
or ( w_24546 , \3013_b1 , w_24548 );
not ( w_24548 , w_24554 );
and ( w_24547 , \3013_b0 , w_24555 );
and ( w_24554 , w_24555 , w_24549 );
buf ( w_24548 , \3015_b1 );
not ( w_24548 , w_24556 );
not ( w_24549 , w_24557 );
and ( w_24556 , w_24557 , \3015_b0 );
or ( \3070_b1 , \3059_b1 , w_24558 );
not ( w_24558 , w_24564 );
and ( \3070_b0 , \3059_b0 , w_24565 );
and ( w_24564 , w_24565 , w_24559 );
or ( w_24558 , \3061_b1 , w_24560 );
not ( w_24560 , w_24566 );
and ( w_24559 , \3061_b0 , w_24567 );
and ( w_24566 , w_24567 , w_24561 );
or ( w_24560 , \3067_b1 , w_24562 );
not ( w_24562 , w_24568 );
and ( w_24561 , \3067_b0 , w_24569 );
and ( w_24568 , w_24569 , w_24563 );
buf ( w_24562 , \3069_b1 );
not ( w_24562 , w_24570 );
not ( w_24563 , w_24571 );
and ( w_24570 , w_24571 , \3069_b0 );
or ( \3109_b1 , \3106_b1 , w_24576 );
or ( \3109_b0 , \3106_b0 , w_24573 );
not ( w_24573 , w_24577 );
and ( w_24577 , w_24576 , w_24572 );
or ( w_24572 , \3107_b1 , w_24578 );
or ( w_24573 , \3107_b0 , w_24575 );
not ( w_24575 , w_24579 );
and ( w_24579 , w_24578 , w_24574 );
buf ( w_24574 , \3108_b1 );
not ( w_24574 , w_24580 );
not ( w_24575 , w_24581 );
and ( w_24580 , w_24581 , \3108_b0 );
or ( \3133_b1 , \3121_b1 , w_24582 );
not ( w_24582 , w_24584 );
and ( \3133_b0 , \3121_b0 , w_24585 );
and ( w_24584 , w_24585 , w_24583 );
or ( w_24582 , \3123_b1 , \3132_b1 );
not ( \3132_b1 , w_24586 );
and ( w_24583 , \3123_b0 , w_24587 );
and ( w_24586 , w_24587 , \3132_b0 );
or ( \3192_b1 , \3148_b1 , w_24588 );
not ( w_24588 , w_24592 );
and ( \3192_b0 , \3148_b0 , w_24593 );
and ( w_24592 , w_24593 , w_24589 );
or ( w_24588 , \3153_b1 , w_24590 );
not ( w_24590 , w_24594 );
and ( w_24589 , \3153_b0 , w_24595 );
and ( w_24594 , w_24595 , w_24591 );
buf ( w_24590 , \3191_b1 );
not ( w_24590 , w_24596 );
not ( w_24591 , w_24597 );
and ( w_24596 , w_24597 , \3191_b0 );
or ( \3282_b1 , \3279_b1 , w_24598 );
not ( w_24598 , w_24602 );
and ( \3282_b0 , \3279_b0 , w_24603 );
and ( w_24602 , w_24603 , w_24599 );
or ( w_24598 , \3281_b1 , w_24600 );
not ( w_24600 , w_24604 );
and ( w_24599 , \3281_b0 , w_24605 );
and ( w_24604 , w_24605 , w_24601 );
buf ( w_24600 , \741_b1 );
not ( w_24600 , w_24606 );
not ( w_24601 , w_24607 );
and ( w_24606 , w_24607 , \741_b0 );
or ( \3303_b1 , \3300_b1 , w_24608 );
not ( w_24608 , w_24612 );
and ( \3303_b0 , \3300_b0 , w_24613 );
and ( w_24612 , w_24613 , w_24609 );
or ( w_24608 , \3302_b1 , w_24610 );
not ( w_24610 , w_24614 );
and ( w_24609 , \3302_b0 , w_24615 );
and ( w_24614 , w_24615 , w_24611 );
buf ( w_24610 , \826_b1 );
not ( w_24610 , w_24616 );
not ( w_24611 , w_24617 );
and ( w_24616 , w_24617 , \826_b0 );
or ( \3567_b1 , \3530_b1 , w_24618 );
not ( w_24618 , w_24620 );
and ( \3567_b0 , \3530_b0 , w_24621 );
and ( w_24620 , w_24621 , w_24619 );
or ( w_24618 , \3532_b1 , \3566_b1 );
not ( \3566_b1 , w_24622 );
and ( w_24619 , \3532_b0 , w_24623 );
and ( w_24622 , w_24623 , \3566_b0 );
or ( \3573_b1 , \3567_b1 , w_24624 );
not ( w_24624 , w_24630 );
and ( \3573_b0 , \3567_b0 , w_24631 );
and ( w_24630 , w_24631 , w_24625 );
or ( w_24624 , \3569_b1 , w_24626 );
not ( w_24626 , w_24632 );
and ( w_24625 , \3569_b0 , w_24633 );
and ( w_24632 , w_24633 , w_24627 );
or ( w_24626 , \3570_b1 , w_24628 );
not ( w_24628 , w_24634 );
and ( w_24627 , \3570_b0 , w_24635 );
and ( w_24634 , w_24635 , w_24629 );
buf ( w_24628 , \3572_b1 );
not ( w_24628 , w_24636 );
not ( w_24629 , w_24637 );
and ( w_24636 , w_24637 , \3572_b0 );
or ( \3629_b1 , \3626_b1 , w_24642 );
or ( \3629_b0 , \3626_b0 , w_24639 );
not ( w_24639 , w_24643 );
and ( w_24643 , w_24642 , w_24638 );
or ( w_24638 , \3627_b1 , w_24644 );
or ( w_24639 , \3627_b0 , w_24641 );
not ( w_24641 , w_24645 );
and ( w_24645 , w_24644 , w_24640 );
buf ( w_24640 , \3628_b1 );
not ( w_24640 , w_24646 );
not ( w_24641 , w_24647 );
and ( w_24646 , w_24647 , \3628_b0 );
or ( \3632_b1 , \3599_b1 , w_24648 );
not ( w_24648 , w_24652 );
and ( \3632_b0 , \3599_b0 , w_24653 );
and ( w_24652 , w_24653 , w_24649 );
or ( w_24648 , \3601_b1 , w_24650 );
not ( w_24650 , w_24654 );
and ( w_24649 , \3601_b0 , w_24655 );
and ( w_24654 , w_24655 , w_24651 );
buf ( w_24650 , \3631_b1 );
not ( w_24650 , w_24656 );
not ( w_24651 , w_24657 );
and ( w_24656 , w_24657 , \3631_b0 );
or ( \3637_b1 , \3585_b1 , w_24658 );
not ( w_24658 , w_24664 );
and ( \3637_b0 , \3585_b0 , w_24665 );
and ( w_24664 , w_24665 , w_24659 );
or ( w_24658 , \3633_b1 , w_24660 );
not ( w_24660 , w_24666 );
and ( w_24659 , \3633_b0 , w_24667 );
and ( w_24666 , w_24667 , w_24661 );
or ( w_24660 , \3634_b1 , w_24662 );
not ( w_24662 , w_24668 );
and ( w_24661 , \3634_b0 , w_24669 );
and ( w_24668 , w_24669 , w_24663 );
buf ( w_24662 , \3636_b1 );
not ( w_24662 , w_24670 );
not ( w_24663 , w_24671 );
and ( w_24670 , w_24671 , \3636_b0 );
or ( \3657_b1 , \2763_b1 , w_24672 );
not ( w_24672 , w_24674 );
and ( \3657_b0 , \2763_b0 , w_24675 );
and ( w_24674 , w_24675 , w_24673 );
or ( w_24672 , \1657_b1 , \1541_b1 );
not ( \1541_b1 , w_24676 );
and ( w_24673 , \1657_b0 , w_24677 );
and ( w_24676 , w_24677 , \1541_b0 );
or ( \3761_b1 , \3759_b1 , w_24678 );
not ( w_24678 , w_24680 );
and ( \3761_b0 , \3759_b0 , w_24681 );
and ( w_24680 , w_24681 , w_24679 );
or ( w_24678 , \3760_b1 , \d[15]_b1 );
not ( \d[15]_b1 , w_24682 );
and ( w_24679 , \3760_b0 , w_24683 );
and ( w_24682 , w_24683 , \d[15]_b0 );
or ( \3833_b1 , \3831_b1 , w_24684 );
not ( w_24684 , w_24686 );
and ( \3833_b0 , \3831_b0 , w_24687 );
and ( w_24686 , w_24687 , w_24685 );
or ( w_24684 , \3832_b1 , \c[15]_b1 );
not ( \c[15]_b1 , w_24688 );
and ( w_24685 , \3832_b0 , w_24689 );
and ( w_24688 , w_24689 , \c[15]_b0 );
or ( \3936_b1 , \3933_b1 , w_24694 );
or ( \3936_b0 , \3933_b0 , w_24691 );
not ( w_24691 , w_24695 );
and ( w_24695 , w_24694 , w_24690 );
or ( w_24690 , \3934_b1 , w_24696 );
or ( w_24691 , \3934_b0 , w_24693 );
not ( w_24693 , w_24697 );
and ( w_24697 , w_24696 , w_24692 );
buf ( w_24692 , \3935_b1 );
not ( w_24692 , w_24698 );
not ( w_24693 , w_24699 );
and ( w_24698 , w_24699 , \3935_b0 );
or ( \3940_b1 , \3937_b1 , w_24700 );
not ( w_24700 , w_24704 );
and ( \3940_b0 , \3937_b0 , w_24705 );
and ( w_24704 , w_24705 , w_24701 );
or ( w_24700 , \3938_b1 , w_24702 );
not ( w_24702 , w_24706 );
and ( w_24701 , \3938_b0 , w_24707 );
and ( w_24706 , w_24707 , w_24703 );
buf ( w_24702 , \3939_b1 );
not ( w_24702 , w_24708 );
not ( w_24703 , w_24709 );
and ( w_24708 , w_24709 , \3939_b0 );
or ( \3949_b1 , \3940_b1 , w_24710 );
not ( w_24710 , w_24716 );
and ( \3949_b0 , \3940_b0 , w_24717 );
and ( w_24716 , w_24717 , w_24711 );
or ( w_24710 , \3943_b1 , w_24712 );
not ( w_24712 , w_24718 );
and ( w_24711 , \3943_b0 , w_24719 );
and ( w_24718 , w_24719 , w_24713 );
or ( w_24712 , \3946_b1 , w_24714 );
not ( w_24714 , w_24720 );
and ( w_24713 , \3946_b0 , w_24721 );
and ( w_24720 , w_24721 , w_24715 );
buf ( w_24714 , \3948_b1 );
not ( w_24714 , w_24722 );
not ( w_24715 , w_24723 );
and ( w_24722 , w_24723 , \3948_b0 );
or ( \3955_b1 , \3952_b1 , w_24724 );
not ( w_24724 , w_24728 );
and ( \3955_b0 , \3952_b0 , w_24729 );
and ( w_24728 , w_24729 , w_24725 );
or ( w_24724 , \3953_b1 , w_24726 );
not ( w_24726 , w_24730 );
and ( w_24725 , \3953_b0 , w_24731 );
and ( w_24730 , w_24731 , w_24727 );
buf ( w_24726 , \3954_b1 );
not ( w_24726 , w_24732 );
not ( w_24727 , w_24733 );
and ( w_24732 , w_24733 , \3954_b0 );
or ( \3976_b1 , \3960_b1 , w_24734 );
not ( w_24734 , w_24736 );
and ( \3976_b0 , \3960_b0 , w_24737 );
and ( w_24736 , w_24737 , w_24735 );
or ( w_24734 , \3968_b1 , \3975_b1 );
not ( \3975_b1 , w_24738 );
and ( w_24735 , \3968_b0 , w_24739 );
and ( w_24738 , w_24739 , \3975_b0 );
or ( \3995_b1 , \3987_b1 , w_24740 );
not ( w_24740 , w_24744 );
and ( \3995_b0 , \3987_b0 , w_24745 );
and ( w_24744 , w_24745 , w_24741 );
or ( w_24740 , \3993_b1 , w_24742 );
not ( w_24742 , w_24746 );
and ( w_24741 , \3993_b0 , w_24747 );
and ( w_24746 , w_24747 , w_24743 );
buf ( w_24742 , \3994_b1 );
not ( w_24742 , w_24748 );
not ( w_24743 , w_24749 );
and ( w_24748 , w_24749 , \3994_b0 );
or ( \4009_b1 , \4007_b1 , w_24750 );
not ( w_24750 , w_24752 );
and ( \4009_b0 , \4007_b0 , w_24753 );
and ( w_24752 , w_24753 , w_24751 );
or ( w_24750 , \3943_b1 , \4008_b1 );
not ( \4008_b1 , w_24754 );
and ( w_24751 , \3943_b0 , w_24755 );
and ( w_24754 , w_24755 , \4008_b0 );
or ( \4030_b1 , \3960_b1 , w_24756 );
not ( w_24756 , w_24758 );
and ( \4030_b0 , \3960_b0 , w_24759 );
and ( w_24758 , w_24759 , w_24757 );
or ( w_24756 , \3968_b1 , \4029_b1 );
not ( \4029_b1 , w_24760 );
and ( w_24757 , \3968_b0 , w_24761 );
and ( w_24760 , w_24761 , \4029_b0 );
or ( \4034_b1 , \3960_b1 , w_24762 );
not ( w_24762 , w_24764 );
and ( \4034_b0 , \3960_b0 , w_24765 );
and ( w_24764 , w_24765 , w_24763 );
or ( w_24762 , \3968_b1 , \3973_b1 );
not ( \3973_b1 , w_24766 );
and ( w_24763 , \3968_b0 , w_24767 );
and ( w_24766 , w_24767 , \3973_b0 );
or ( \4045_b1 , \4040_b1 , w_24770 );
or ( \4045_b0 , \4040_b0 , w_24769 );
not ( w_24769 , w_24771 );
and ( w_24771 , w_24770 , w_24768 );
or ( w_24768 , \3967_b1 , w_24772 );
or ( w_24769 , \3967_b0 , \4044_b0 );
not ( \4044_b0 , w_24773 );
and ( w_24773 , w_24772 , \4044_b1 );
or ( \4050_b1 , \4046_b1 , w_24778 );
or ( \4050_b0 , \4046_b0 , w_24775 );
not ( w_24775 , w_24779 );
and ( w_24779 , w_24778 , w_24774 );
or ( w_24774 , \4047_b1 , w_24780 );
or ( w_24775 , \4047_b0 , w_24777 );
not ( w_24777 , w_24781 );
and ( w_24781 , w_24780 , w_24776 );
buf ( w_24776 , \4049_b1 );
not ( w_24776 , w_24782 );
not ( w_24777 , w_24783 );
and ( w_24782 , w_24783 , \4049_b0 );
or ( \4053_b1 , \3960_b1 , w_24784 );
not ( w_24784 , w_24786 );
and ( \4053_b0 , \3960_b0 , w_24787 );
and ( w_24786 , w_24787 , w_24785 );
or ( w_24784 , \3966_b1 , \4052_b1 );
not ( \4052_b1 , w_24788 );
and ( w_24785 , \3966_b0 , w_24789 );
and ( w_24788 , w_24789 , \4052_b0 );
or ( \4099_b1 , \3926_b1 , w_24790 );
not ( w_24790 , w_24796 );
and ( \4099_b0 , \3926_b0 , w_24797 );
and ( w_24796 , w_24797 , w_24791 );
or ( w_24790 , \3788_b1 , w_24792 );
not ( w_24792 , w_24798 );
and ( w_24791 , \3788_b0 , w_24799 );
and ( w_24798 , w_24799 , w_24793 );
or ( w_24792 , \3517_b1 , w_24794 );
not ( w_24794 , w_24800 );
and ( w_24793 , \3517_b0 , w_24801 );
and ( w_24800 , w_24801 , w_24795 );
buf ( w_24794 , \927_b1 );
not ( w_24794 , w_24802 );
not ( w_24795 , w_24803 );
and ( w_24802 , w_24803 , \927_b0 );
or ( \4185_b1 , \3926_b1 , w_24804 );
not ( w_24804 , w_24808 );
and ( \4185_b0 , \3926_b0 , w_24809 );
and ( w_24808 , w_24809 , w_24805 );
or ( w_24804 , \3788_b1 , w_24806 );
not ( w_24806 , w_24810 );
and ( w_24805 , \3788_b0 , w_24811 );
and ( w_24810 , w_24811 , w_24807 );
or ( w_24806 , \3517_b1 , \927_b1 );
not ( \927_b1 , w_24812 );
and ( w_24807 , \3517_b0 , w_24813 );
and ( w_24812 , w_24813 , \927_b0 );
or ( \5649_b1 , \5618_b1 , w_24814 );
not ( w_24814 , w_24816 );
and ( \5649_b0 , \5618_b0 , w_24817 );
and ( w_24816 , w_24817 , w_24815 );
or ( w_24814 , \5641_b1 , \5648_b1 );
not ( \5648_b1 , w_24818 );
and ( w_24815 , \5641_b0 , w_24819 );
and ( w_24818 , w_24819 , \5648_b0 );
or ( \5732_b1 , \4102_b1 , w_24820 );
not ( w_24820 , w_24824 );
and ( \5732_b0 , \4102_b0 , w_24825 );
and ( w_24824 , w_24825 , w_24821 );
or ( w_24820 , \5729_b1 , w_24822 );
not ( w_24822 , w_24826 );
and ( w_24821 , \5729_b0 , w_24827 );
and ( w_24826 , w_24827 , w_24823 );
buf ( w_24822 , \5731_b1 );
not ( w_24822 , w_24828 );
not ( w_24823 , w_24829 );
and ( w_24828 , w_24829 , \5731_b0 );
or ( \5979_b1 , \4862_b1 , w_24830 );
not ( w_24830 , w_24834 );
and ( \5979_b0 , \4862_b0 , w_24835 );
and ( w_24834 , w_24835 , w_24831 );
or ( w_24830 , \5978_b1 , w_24832 );
not ( w_24832 , w_24836 );
and ( w_24831 , \5978_b0 , w_24837 );
and ( w_24836 , w_24837 , w_24833 );
buf ( w_24832 , \4858_b1 );
not ( w_24832 , w_24838 );
not ( w_24833 , w_24839 );
and ( w_24838 , w_24839 , \4858_b0 );
or ( \6289_b1 , \6034_b1 , w_24840 );
not ( w_24840 , w_24844 );
and ( \6289_b0 , \6034_b0 , w_24845 );
and ( w_24844 , w_24845 , w_24841 );
or ( w_24840 , \6279_b1 , w_24842 );
not ( w_24842 , w_24846 );
and ( w_24841 , \6279_b0 , w_24847 );
and ( w_24846 , w_24847 , w_24843 );
buf ( w_24842 , \6288_b1 );
not ( w_24842 , w_24848 );
not ( w_24843 , w_24849 );
and ( w_24848 , w_24849 , \6288_b0 );
or ( \6327_b1 , \6325_b1 , w_24850 );
not ( w_24850 , w_24852 );
and ( \6327_b0 , \6325_b0 , w_24853 );
and ( w_24852 , w_24853 , w_24851 );
or ( w_24850 , \4616_b1 , \6326_b1 );
not ( \6326_b1 , w_24854 );
and ( w_24851 , \4616_b0 , w_24855 );
and ( w_24854 , w_24855 , \6326_b0 );
or ( \6656_b1 , \6654_b1 , w_24856 );
not ( w_24856 , w_24860 );
and ( \6656_b0 , \6654_b0 , w_24861 );
and ( w_24860 , w_24861 , w_24857 );
or ( w_24856 , \4285_b1 , w_24858 );
not ( w_24858 , w_24862 );
and ( w_24857 , \4285_b0 , w_24863 );
and ( w_24862 , w_24863 , w_24859 );
buf ( w_24858 , \6655_b1 );
not ( w_24858 , w_24864 );
not ( w_24859 , w_24865 );
and ( w_24864 , w_24865 , \6655_b0 );
or ( \6810_b1 , \4862_b1 , w_24866 );
not ( w_24866 , w_24870 );
and ( \6810_b0 , \4862_b0 , w_24871 );
and ( w_24870 , w_24871 , w_24867 );
or ( w_24866 , \6684_b1 , w_24868 );
not ( w_24868 , w_24872 );
and ( w_24867 , \6684_b0 , w_24873 );
and ( w_24872 , w_24873 , w_24869 );
buf ( w_24868 , \4858_b1 );
not ( w_24868 , w_24874 );
not ( w_24869 , w_24875 );
and ( w_24874 , w_24875 , \4858_b0 );
or ( \6965_b1 , \6908_b1 , w_24876 );
not ( w_24876 , w_24880 );
and ( \6965_b0 , \6908_b0 , w_24881 );
and ( w_24880 , w_24881 , w_24877 );
or ( w_24876 , \6954_b1 , w_24878 );
not ( w_24878 , w_24882 );
and ( w_24877 , \6954_b0 , w_24883 );
and ( w_24882 , w_24883 , w_24879 );
buf ( w_24878 , \6964_b1 );
not ( w_24878 , w_24884 );
not ( w_24879 , w_24885 );
and ( w_24884 , w_24885 , \6964_b0 );
or ( \6979_b1 , \6964_b1 , w_24886 );
not ( w_24886 , w_24888 );
and ( \6979_b0 , \6964_b0 , w_24889 );
and ( w_24888 , w_24889 , w_24887 );
or ( w_24886 , \6978_b1 , \6944_b1 );
not ( \6944_b1 , w_24890 );
and ( w_24887 , \6978_b0 , w_24891 );
and ( w_24890 , w_24891 , \6944_b0 );
or ( \7116_b1 , \7068_b1 , w_24892 );
not ( w_24892 , w_24894 );
and ( \7116_b0 , \7068_b0 , w_24895 );
and ( w_24894 , w_24895 , w_24893 );
or ( w_24892 , \7076_b1 , \7115_b1 );
not ( \7115_b1 , w_24896 );
and ( w_24893 , \7076_b0 , w_24897 );
and ( w_24896 , w_24897 , \7115_b0 );
or ( \7138_b1 , \5707_b1 , w_24898 );
not ( w_24898 , w_24902 );
and ( \7138_b0 , \5707_b0 , w_24903 );
and ( w_24902 , w_24903 , w_24899 );
or ( w_24898 , \6290_b1 , w_24900 );
not ( w_24900 , w_24904 );
and ( w_24899 , \6290_b0 , w_24905 );
and ( w_24904 , w_24905 , w_24901 );
buf ( w_24900 , \7137_b1 );
not ( w_24900 , w_24906 );
not ( w_24901 , w_24907 );
and ( w_24906 , w_24907 , \7137_b0 );
or ( \7170_b1 , \7138_b1 , w_24908 );
not ( w_24908 , w_24912 );
and ( \7170_b0 , \7138_b0 , w_24913 );
and ( w_24912 , w_24913 , w_24909 );
or ( w_24908 , \7155_b1 , w_24910 );
not ( w_24910 , w_24914 );
and ( w_24909 , \7155_b0 , w_24915 );
and ( w_24914 , w_24915 , w_24911 );
buf ( w_24910 , \7169_b1 );
not ( w_24910 , w_24916 );
not ( w_24911 , w_24917 );
and ( w_24916 , w_24917 , \7169_b0 );
or ( \7241_b1 , \7138_b1 , w_24918 );
not ( w_24918 , w_24922 );
and ( \7241_b0 , \7138_b0 , w_24923 );
and ( w_24922 , w_24923 , w_24919 );
or ( w_24918 , \7155_b1 , w_24920 );
not ( w_24920 , w_24924 );
and ( w_24919 , \7155_b0 , w_24925 );
and ( w_24924 , w_24925 , w_24921 );
buf ( w_24920 , \7169_b1 );
not ( w_24920 , w_24926 );
not ( w_24921 , w_24927 );
and ( w_24926 , w_24927 , \7169_b0 );
endmodule

