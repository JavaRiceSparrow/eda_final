// ...
module top(\s[31]_b1 ,\s[31]_b0 ,\s[30]_b1 ,\s[30]_b0 ,\s[29]_b1 ,\s[29]_b0 ,\s[28]_b1 ,\s[28]_b0 ,\s[27]_b1 ,
		\s[27]_b0 ,\s[26]_b1 ,\s[26]_b0 ,\s[25]_b1 ,\s[25]_b0 ,\s[24]_b1 ,\s[24]_b0 ,\s[23]_b1 ,\s[23]_b0 ,
		\s[22]_b1 ,\s[22]_b0 ,\s[21]_b1 ,\s[21]_b0 ,\s[20]_b1 ,\s[20]_b0 ,\s[19]_b1 ,\s[19]_b0 ,\s[18]_b1 ,
		\s[18]_b0 ,\s[17]_b1 ,\s[17]_b0 ,\s[16]_b1 ,\s[16]_b0 ,\s[15]_b1 ,\s[15]_b0 ,\s[14]_b1 ,\s[14]_b0 ,
		\s[13]_b1 ,\s[13]_b0 ,\s[12]_b1 ,\s[12]_b0 ,\s[11]_b1 ,\s[11]_b0 ,\s[10]_b1 ,\s[10]_b0 ,\s[9]_b1 ,
		\s[9]_b0 ,\s[8]_b1 ,\s[8]_b0 ,\s[7]_b1 ,\s[7]_b0 ,\s[6]_b1 ,\s[6]_b0 ,\s[5]_b1 ,\s[5]_b0 ,
		\s[4]_b1 ,\s[4]_b0 ,\s[3]_b1 ,\s[3]_b0 ,\s[2]_b1 ,\s[2]_b0 ,\s[1]_b1 ,\s[1]_b0 ,\s[0]_b1 ,
		\s[0]_b0 ,\a[31]_b1 ,\a[31]_b0 ,\a[30]_b1 ,\a[30]_b0 ,\a[29]_b1 ,\a[29]_b0 ,\a[28]_b1 ,\a[28]_b0 ,
		\a[27]_b1 ,\a[27]_b0 ,\a[26]_b1 ,\a[26]_b0 ,\a[25]_b1 ,\a[25]_b0 ,\a[24]_b1 ,\a[24]_b0 ,\a[23]_b1 ,
		\a[23]_b0 ,\a[22]_b1 ,\a[22]_b0 ,\a[21]_b1 ,\a[21]_b0 ,\a[20]_b1 ,\a[20]_b0 ,\a[19]_b1 ,\a[19]_b0 ,
		\a[18]_b1 ,\a[18]_b0 ,\a[17]_b1 ,\a[17]_b0 ,\a[16]_b1 ,\a[16]_b0 ,\a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,
		\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,
		\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,
		\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,
		\a[0]_b1 ,\a[0]_b0 ,\b[31]_b1 ,\b[31]_b0 ,\b[30]_b1 ,\b[30]_b0 ,\b[29]_b1 ,\b[29]_b0 ,\b[28]_b1 ,
		\b[28]_b0 ,\b[27]_b1 ,\b[27]_b0 ,\b[26]_b1 ,\b[26]_b0 ,\b[25]_b1 ,\b[25]_b0 ,\b[24]_b1 ,\b[24]_b0 ,
		\b[23]_b1 ,\b[23]_b0 ,\b[22]_b1 ,\b[22]_b0 ,\b[21]_b1 ,\b[21]_b0 ,\b[20]_b1 ,\b[20]_b0 ,\b[19]_b1 ,
		\b[19]_b0 ,\b[18]_b1 ,\b[18]_b0 ,\b[17]_b1 ,\b[17]_b0 ,\b[16]_b1 ,\b[16]_b0 ,\b[15]_b1 ,\b[15]_b0 ,
		\b[14]_b1 ,\b[14]_b0 ,\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,
		\b[10]_b0 ,\b[9]_b1 ,\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,
		\b[5]_b1 ,\b[5]_b0 ,\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,
		\b[1]_b0 ,\b[0]_b1 ,\b[0]_b0 ,\c[31]_b1 ,\c[31]_b0 ,\c[30]_b1 ,\c[30]_b0 ,\c[29]_b1 ,\c[29]_b0 ,
		\c[28]_b1 ,\c[28]_b0 ,\c[27]_b1 ,\c[27]_b0 ,\c[26]_b1 ,\c[26]_b0 ,\c[25]_b1 ,\c[25]_b0 ,\c[24]_b1 ,
		\c[24]_b0 ,\c[23]_b1 ,\c[23]_b0 ,\c[22]_b1 ,\c[22]_b0 ,\c[21]_b1 ,\c[21]_b0 ,\c[20]_b1 ,\c[20]_b0 ,
		\c[19]_b1 ,\c[19]_b0 ,\c[18]_b1 ,\c[18]_b0 ,\c[17]_b1 ,\c[17]_b0 ,\c[16]_b1 ,\c[16]_b0 ,\c[15]_b1 ,
		\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,\c[11]_b1 ,\c[11]_b0 ,
		\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,\c[7]_b0 ,\c[6]_b1 ,
		\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,\c[2]_b1 ,\c[2]_b0 ,
		\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[31]_b1 ,\d[31]_b0 ,\d[30]_b1 ,\d[30]_b0 ,\d[29]_b1 ,
		\d[29]_b0 ,\d[28]_b1 ,\d[28]_b0 ,\d[27]_b1 ,\d[27]_b0 ,\d[26]_b1 ,\d[26]_b0 ,\d[25]_b1 ,\d[25]_b0 ,
		\d[24]_b1 ,\d[24]_b0 ,\d[23]_b1 ,\d[23]_b0 ,\d[22]_b1 ,\d[22]_b0 ,\d[21]_b1 ,\d[21]_b0 ,\d[20]_b1 ,
		\d[20]_b0 ,\d[19]_b1 ,\d[19]_b0 ,\d[18]_b1 ,\d[18]_b0 ,\d[17]_b1 ,\d[17]_b0 ,\d[16]_b1 ,\d[16]_b0 ,
		\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,
		\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,
		\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,
		\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,\d[0]_b1 ,\d[0]_b0 ,\o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,
		\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,\o[28]_b0 ,\o[27]_b1 ,\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,
		\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,\o[23]_b1 ,\o[23]_b0 ,\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,
		\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,\o[19]_b0 ,\o[18]_b1 ,\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,
		\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,\o[14]_b1 ,\o[14]_b0 ,\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,
		\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,\o[10]_b0 ,\o[9]_b1 ,\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,
		\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,\o[5]_b1 ,\o[5]_b0 ,\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,
		\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,\o[1]_b0 ,\o[0]_b1 ,\o[0]_b0 );
input \s[31]_b1 ,\s[31]_b0 ,\s[30]_b1 ,\s[30]_b0 ,\s[29]_b1 ,\s[29]_b0 ,\s[28]_b1 ,\s[28]_b0 ,\s[27]_b1 ,
		\s[27]_b0 ,\s[26]_b1 ,\s[26]_b0 ,\s[25]_b1 ,\s[25]_b0 ,\s[24]_b1 ,\s[24]_b0 ,\s[23]_b1 ,\s[23]_b0 ,
		\s[22]_b1 ,\s[22]_b0 ,\s[21]_b1 ,\s[21]_b0 ,\s[20]_b1 ,\s[20]_b0 ,\s[19]_b1 ,\s[19]_b0 ,\s[18]_b1 ,
		\s[18]_b0 ,\s[17]_b1 ,\s[17]_b0 ,\s[16]_b1 ,\s[16]_b0 ,\s[15]_b1 ,\s[15]_b0 ,\s[14]_b1 ,\s[14]_b0 ,
		\s[13]_b1 ,\s[13]_b0 ,\s[12]_b1 ,\s[12]_b0 ,\s[11]_b1 ,\s[11]_b0 ,\s[10]_b1 ,\s[10]_b0 ,\s[9]_b1 ,
		\s[9]_b0 ,\s[8]_b1 ,\s[8]_b0 ,\s[7]_b1 ,\s[7]_b0 ,\s[6]_b1 ,\s[6]_b0 ,\s[5]_b1 ,\s[5]_b0 ,
		\s[4]_b1 ,\s[4]_b0 ,\s[3]_b1 ,\s[3]_b0 ,\s[2]_b1 ,\s[2]_b0 ,\s[1]_b1 ,\s[1]_b0 ,\s[0]_b1 ,
		\s[0]_b0 ,\a[31]_b1 ,\a[31]_b0 ,\a[30]_b1 ,\a[30]_b0 ,\a[29]_b1 ,\a[29]_b0 ,\a[28]_b1 ,\a[28]_b0 ,
		\a[27]_b1 ,\a[27]_b0 ,\a[26]_b1 ,\a[26]_b0 ,\a[25]_b1 ,\a[25]_b0 ,\a[24]_b1 ,\a[24]_b0 ,\a[23]_b1 ,
		\a[23]_b0 ,\a[22]_b1 ,\a[22]_b0 ,\a[21]_b1 ,\a[21]_b0 ,\a[20]_b1 ,\a[20]_b0 ,\a[19]_b1 ,\a[19]_b0 ,
		\a[18]_b1 ,\a[18]_b0 ,\a[17]_b1 ,\a[17]_b0 ,\a[16]_b1 ,\a[16]_b0 ,\a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,
		\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,
		\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,
		\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,
		\a[0]_b1 ,\a[0]_b0 ,\b[31]_b1 ,\b[31]_b0 ,\b[30]_b1 ,\b[30]_b0 ,\b[29]_b1 ,\b[29]_b0 ,\b[28]_b1 ,
		\b[28]_b0 ,\b[27]_b1 ,\b[27]_b0 ,\b[26]_b1 ,\b[26]_b0 ,\b[25]_b1 ,\b[25]_b0 ,\b[24]_b1 ,\b[24]_b0 ,
		\b[23]_b1 ,\b[23]_b0 ,\b[22]_b1 ,\b[22]_b0 ,\b[21]_b1 ,\b[21]_b0 ,\b[20]_b1 ,\b[20]_b0 ,\b[19]_b1 ,
		\b[19]_b0 ,\b[18]_b1 ,\b[18]_b0 ,\b[17]_b1 ,\b[17]_b0 ,\b[16]_b1 ,\b[16]_b0 ,\b[15]_b1 ,\b[15]_b0 ,
		\b[14]_b1 ,\b[14]_b0 ,\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,
		\b[10]_b0 ,\b[9]_b1 ,\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,
		\b[5]_b1 ,\b[5]_b0 ,\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,
		\b[1]_b0 ,\b[0]_b1 ,\b[0]_b0 ,\c[31]_b1 ,\c[31]_b0 ,\c[30]_b1 ,\c[30]_b0 ,\c[29]_b1 ,\c[29]_b0 ,
		\c[28]_b1 ,\c[28]_b0 ,\c[27]_b1 ,\c[27]_b0 ,\c[26]_b1 ,\c[26]_b0 ,\c[25]_b1 ,\c[25]_b0 ,\c[24]_b1 ,
		\c[24]_b0 ,\c[23]_b1 ,\c[23]_b0 ,\c[22]_b1 ,\c[22]_b0 ,\c[21]_b1 ,\c[21]_b0 ,\c[20]_b1 ,\c[20]_b0 ,
		\c[19]_b1 ,\c[19]_b0 ,\c[18]_b1 ,\c[18]_b0 ,\c[17]_b1 ,\c[17]_b0 ,\c[16]_b1 ,\c[16]_b0 ,\c[15]_b1 ,
		\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,\c[11]_b1 ,\c[11]_b0 ,
		\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,\c[7]_b0 ,\c[6]_b1 ,
		\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,\c[2]_b1 ,\c[2]_b0 ,
		\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[31]_b1 ,\d[31]_b0 ,\d[30]_b1 ,\d[30]_b0 ,\d[29]_b1 ,
		\d[29]_b0 ,\d[28]_b1 ,\d[28]_b0 ,\d[27]_b1 ,\d[27]_b0 ,\d[26]_b1 ,\d[26]_b0 ,\d[25]_b1 ,\d[25]_b0 ,
		\d[24]_b1 ,\d[24]_b0 ,\d[23]_b1 ,\d[23]_b0 ,\d[22]_b1 ,\d[22]_b0 ,\d[21]_b1 ,\d[21]_b0 ,\d[20]_b1 ,
		\d[20]_b0 ,\d[19]_b1 ,\d[19]_b0 ,\d[18]_b1 ,\d[18]_b0 ,\d[17]_b1 ,\d[17]_b0 ,\d[16]_b1 ,\d[16]_b0 ,
		\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,
		\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,
		\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,
		\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,\d[0]_b1 ,\d[0]_b0 ;
output \o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,\o[28]_b0 ,\o[27]_b1 ,
		\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,\o[23]_b1 ,\o[23]_b0 ,
		\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,\o[19]_b0 ,\o[18]_b1 ,
		\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,\o[14]_b1 ,\o[14]_b0 ,
		\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,\o[10]_b0 ,\o[9]_b1 ,
		\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,\o[5]_b1 ,\o[5]_b0 ,
		\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,\o[1]_b0 ,\o[0]_b1 ,
		\o[0]_b0 ;

wire \193_ZERO_b1 , \193_ZERO_b0 , \194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , \197_b1 , \197_b0 , 
		\198_b1 , \198_b0 , \199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , \202_b1 , \202_b0 , 
		\203_b1 , \203_b0 , \204_ONE_b1 , \204_ONE_b0 , \205_n5[0]_b1 , \205_n5[0]_b0 , \206_b1 , \206_b0 , \207_A[0]_b1 , \207_A[0]_b0 , 
		\208_B[0]_b1 , \208_B[0]_b0 , \209_b1 , \209_b0 , \210_SUM[0]_b1 , \210_SUM[0]_b0 , \211_b1 , \211_b0 , \212_b1 , \212_b0 , 
		\213_b1 , \213_b0 , \214_b1 , \214_b0 , \215_b1 , \215_b0 , \216_b1 , \216_b0 , \217_b1 , \217_b0 , 
		\218_b1 , \218_b0 , \219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , \222_b1 , \222_b0 , 
		\223_b1 , \223_b0 , \224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , \227_b1 , \227_b0 , 
		\228_b1 , \228_b0 , \229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , \232_b1 , \232_b0 , 
		\233_b1 , \233_b0 , \234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , \237_b1 , \237_b0 , 
		\238_b1 , \238_b0 , \239_b1 , \239_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , \242_b1 , \242_b0 , 
		\243_A[0]_b1 , \243_A[0]_b0 , \244_B[0]_b1 , \244_B[0]_b0 , \245_b1 , \245_b0 , \246_SUM[0]_b1 , \246_SUM[0]_b0 , \247_b1 , \247_b0 , 
		\248_b1 , \248_b0 , \249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , \252_b1 , \252_b0 , 
		\253_b1 , \253_b0 , \254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , \257_b1 , \257_b0 , 
		\258_b1 , \258_b0 , \259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , \262_b1 , \262_b0 , 
		\263_b1 , \263_b0 , \264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , \267_b1 , \267_b0 , 
		\268_b1 , \268_b0 , \269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , \272_b1 , \272_b0 , 
		\273_b1 , \273_b0 , \274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_b1 , \276_b0 , \277_b1 , \277_b0 , 
		\278_b1 , \278_b0 , \279_n5[1]_b1 , \279_n5[1]_b0 , \280_b1 , \280_b0 , \281_A[1]_b1 , \281_A[1]_b0 , \282_B[1]_b1 , \282_B[1]_b0 , 
		\283_b1 , \283_b0 , \284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , \287_b1 , \287_b0 , 
		\288_SUM[1]_b1 , \288_SUM[1]_b0 , \289_b1 , \289_b0 , \290_A[1]_b1 , \290_A[1]_b0 , \291_B[1]_b1 , \291_B[1]_b0 , \292_b1 , \292_b0 , 
		\293_b1 , \293_b0 , \294_b1 , \294_b0 , \295_SUM[1]_b1 , \295_SUM[1]_b0 , \296_b1 , \296_b0 , \297_n5[2]_b1 , \297_n5[2]_b0 , 
		\298_b1 , \298_b0 , \299_A[2]_b1 , \299_A[2]_b0 , \300_B[2]_b1 , \300_B[2]_b0 , \301_b1 , \301_b0 , \302_b1 , \302_b0 , 
		\303_b1 , \303_b0 , \304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , \307_b1 , \307_b0 , 
		\308_SUM[2]_b1 , \308_SUM[2]_b0 , \309_b1 , \309_b0 , \310_A[2]_b1 , \310_A[2]_b0 , \311_B[2]_b1 , \311_B[2]_b0 , \312_b1 , \312_b0 , 
		\313_b1 , \313_b0 , \314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_b1 , \316_b0 , \317_b1 , \317_b0 , 
		\318_SUM[2]_b1 , \318_SUM[2]_b0 , \319_b1 , \319_b0 , \320_n5[3]_b1 , \320_n5[3]_b0 , \321_b1 , \321_b0 , \322_A[3]_b1 , \322_A[3]_b0 , 
		\323_B[3]_b1 , \323_B[3]_b0 , \324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , \327_b1 , \327_b0 , 
		\328_b1 , \328_b0 , \329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_SUM[3]_b1 , \331_SUM[3]_b0 , \332_b1 , \332_b0 , 
		\333_A[3]_b1 , \333_A[3]_b0 , \334_B[3]_b1 , \334_B[3]_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , \337_b1 , \337_b0 , 
		\338_b1 , \338_b0 , \339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_SUM[3]_b1 , \341_SUM[3]_b0 , \342_b1 , \342_b0 , 
		\343_n5[4]_b1 , \343_n5[4]_b0 , \344_b1 , \344_b0 , \345_A[4]_b1 , \345_A[4]_b0 , \346_B[4]_b1 , \346_B[4]_b0 , \347_b1 , \347_b0 , 
		\348_b1 , \348_b0 , \349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , \352_b1 , \352_b0 , 
		\353_b1 , \353_b0 , \354_SUM[4]_b1 , \354_SUM[4]_b0 , \355_b1 , \355_b0 , \356_A[4]_b1 , \356_A[4]_b0 , \357_B[4]_b1 , \357_B[4]_b0 , 
		\358_b1 , \358_b0 , \359_b1 , \359_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , \362_b1 , \362_b0 , 
		\363_b1 , \363_b0 , \364_SUM[4]_b1 , \364_SUM[4]_b0 , \365_b1 , \365_b0 , \366_n5[5]_b1 , \366_n5[5]_b0 , \367_b1 , \367_b0 , 
		\368_A[5]_b1 , \368_A[5]_b0 , \369_B[5]_b1 , \369_B[5]_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , \372_b1 , \372_b0 , 
		\373_b1 , \373_b0 , \374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , \377_SUM[5]_b1 , \377_SUM[5]_b0 , 
		\378_b1 , \378_b0 , \379_A[5]_b1 , \379_A[5]_b0 , \380_B[5]_b1 , \380_B[5]_b0 , \381_b1 , \381_b0 , \382_b1 , \382_b0 , 
		\383_b1 , \383_b0 , \384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , \387_SUM[5]_b1 , \387_SUM[5]_b0 , 
		\388_b1 , \388_b0 , \389_n5[6]_b1 , \389_n5[6]_b0 , \390_b1 , \390_b0 , \391_A[6]_b1 , \391_A[6]_b0 , \392_B[6]_b1 , \392_B[6]_b0 , 
		\393_b1 , \393_b0 , \394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , \397_b1 , \397_b0 , 
		\398_b1 , \398_b0 , \399_b1 , \399_b0 , \400_SUM[6]_b1 , \400_SUM[6]_b0 , \401_b1 , \401_b0 , \402_A[6]_b1 , \402_A[6]_b0 , 
		\403_B[6]_b1 , \403_B[6]_b0 , \404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , \407_b1 , \407_b0 , 
		\408_b1 , \408_b0 , \409_b1 , \409_b0 , \410_SUM[6]_b1 , \410_SUM[6]_b0 , \411_b1 , \411_b0 , \412_n5[7]_b1 , \412_n5[7]_b0 , 
		\413_b1 , \413_b0 , \414_A[7]_b1 , \414_A[7]_b0 , \415_B[7]_b1 , \415_B[7]_b0 , \416_b1 , \416_b0 , \417_b1 , \417_b0 , 
		\418_b1 , \418_b0 , \419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , \422_b1 , \422_b0 , 
		\423_SUM[7]_b1 , \423_SUM[7]_b0 , \424_b1 , \424_b0 , \425_A[7]_b1 , \425_A[7]_b0 , \426_B[7]_b1 , \426_B[7]_b0 , \427_b1 , \427_b0 , 
		\428_b1 , \428_b0 , \429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , \432_b1 , \432_b0 , 
		\433_SUM[7]_b1 , \433_SUM[7]_b0 , \434_b1 , \434_b0 , \435_n5[8]_b1 , \435_n5[8]_b0 , \436_b1 , \436_b0 , \437_A[8]_b1 , \437_A[8]_b0 , 
		\438_B[8]_b1 , \438_B[8]_b0 , \439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , \442_b1 , \442_b0 , 
		\443_b1 , \443_b0 , \444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_SUM[8]_b1 , \446_SUM[8]_b0 , \447_b1 , \447_b0 , 
		\448_A[8]_b1 , \448_A[8]_b0 , \449_B[8]_b1 , \449_B[8]_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , \452_b1 , \452_b0 , 
		\453_b1 , \453_b0 , \454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_SUM[8]_b1 , \456_SUM[8]_b0 , \457_b1 , \457_b0 , 
		\458_n5[9]_b1 , \458_n5[9]_b0 , \459_b1 , \459_b0 , \460_A[9]_b1 , \460_A[9]_b0 , \461_B[9]_b1 , \461_B[9]_b0 , \462_b1 , \462_b0 , 
		\463_b1 , \463_b0 , \464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , \467_b1 , \467_b0 , 
		\468_b1 , \468_b0 , \469_SUM[9]_b1 , \469_SUM[9]_b0 , \470_b1 , \470_b0 , \471_A[9]_b1 , \471_A[9]_b0 , \472_B[9]_b1 , \472_B[9]_b0 , 
		\473_b1 , \473_b0 , \474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , \477_b1 , \477_b0 , 
		\478_b1 , \478_b0 , \479_SUM[9]_b1 , \479_SUM[9]_b0 , \480_b1 , \480_b0 , \481_n5[10]_b1 , \481_n5[10]_b0 , \482_b1 , \482_b0 , 
		\483_A[10]_b1 , \483_A[10]_b0 , \484_B[10]_b1 , \484_B[10]_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , \487_b1 , \487_b0 , 
		\488_b1 , \488_b0 , \489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , \492_SUM[10]_b1 , \492_SUM[10]_b0 , 
		\493_b1 , \493_b0 , \494_A[10]_b1 , \494_A[10]_b0 , \495_B[10]_b1 , \495_B[10]_b0 , \496_b1 , \496_b0 , \497_b1 , \497_b0 , 
		\498_b1 , \498_b0 , \499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , \502_SUM[10]_b1 , \502_SUM[10]_b0 , 
		\503_b1 , \503_b0 , \504_n5[11]_b1 , \504_n5[11]_b0 , \505_b1 , \505_b0 , \506_A[11]_b1 , \506_A[11]_b0 , \507_B[11]_b1 , \507_B[11]_b0 , 
		\508_b1 , \508_b0 , \509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , \512_b1 , \512_b0 , 
		\513_b1 , \513_b0 , \514_b1 , \514_b0 , \515_SUM[11]_b1 , \515_SUM[11]_b0 , \516_b1 , \516_b0 , \517_A[11]_b1 , \517_A[11]_b0 , 
		\518_B[11]_b1 , \518_B[11]_b0 , \519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , \522_b1 , \522_b0 , 
		\523_b1 , \523_b0 , \524_b1 , \524_b0 , \525_SUM[11]_b1 , \525_SUM[11]_b0 , \526_b1 , \526_b0 , \527_n5[12]_b1 , \527_n5[12]_b0 , 
		\528_b1 , \528_b0 , \529_A[12]_b1 , \529_A[12]_b0 , \530_B[12]_b1 , \530_B[12]_b0 , \531_b1 , \531_b0 , \532_b1 , \532_b0 , 
		\533_b1 , \533_b0 , \534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_b1 , \536_b0 , \537_b1 , \537_b0 , 
		\538_SUM[12]_b1 , \538_SUM[12]_b0 , \539_b1 , \539_b0 , \540_A[12]_b1 , \540_A[12]_b0 , \541_B[12]_b1 , \541_B[12]_b0 , \542_b1 , \542_b0 , 
		\543_b1 , \543_b0 , \544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , \547_b1 , \547_b0 , 
		\548_SUM[12]_b1 , \548_SUM[12]_b0 , \549_b1 , \549_b0 , \550_n5[13]_b1 , \550_n5[13]_b0 , \551_b1 , \551_b0 , \552_A[13]_b1 , \552_A[13]_b0 , 
		\553_B[13]_b1 , \553_B[13]_b0 , \554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , \557_b1 , \557_b0 , 
		\558_b1 , \558_b0 , \559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_SUM[13]_b1 , \561_SUM[13]_b0 , \562_b1 , \562_b0 , 
		\563_A[13]_b1 , \563_A[13]_b0 , \564_B[13]_b1 , \564_B[13]_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , \567_b1 , \567_b0 , 
		\568_b1 , \568_b0 , \569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_SUM[13]_b1 , \571_SUM[13]_b0 , \572_b1 , \572_b0 , 
		\573_n5[14]_b1 , \573_n5[14]_b0 , \574_b1 , \574_b0 , \575_A[14]_b1 , \575_A[14]_b0 , \576_B[14]_b1 , \576_B[14]_b0 , \577_b1 , \577_b0 , 
		\578_b1 , \578_b0 , \579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , \582_b1 , \582_b0 , 
		\583_b1 , \583_b0 , \584_SUM[14]_b1 , \584_SUM[14]_b0 , \585_b1 , \585_b0 , \586_A[14]_b1 , \586_A[14]_b0 , \587_B[14]_b1 , \587_B[14]_b0 , 
		\588_b1 , \588_b0 , \589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , \592_b1 , \592_b0 , 
		\593_b1 , \593_b0 , \594_SUM[14]_b1 , \594_SUM[14]_b0 , \595_b1 , \595_b0 , \596_n5[15]_b1 , \596_n5[15]_b0 , \597_b1 , \597_b0 , 
		\598_A[15]_b1 , \598_A[15]_b0 , \599_B[15]_b1 , \599_B[15]_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , \602_b1 , \602_b0 , 
		\603_b1 , \603_b0 , \604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_b1 , \606_b0 , \607_SUM[15]_b1 , \607_SUM[15]_b0 , 
		\608_b1 , \608_b0 , \609_A[15]_b1 , \609_A[15]_b0 , \610_B[15]_b1 , \610_B[15]_b0 , \611_b1 , \611_b0 , \612_b1 , \612_b0 , 
		\613_b1 , \613_b0 , \614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , \617_SUM[15]_b1 , \617_SUM[15]_b0 , 
		\618_b1 , \618_b0 , \619_n5[16]_b1 , \619_n5[16]_b0 , \620_b1 , \620_b0 , \621_A[16]_b1 , \621_A[16]_b0 , \622_B[16]_b1 , \622_B[16]_b0 , 
		\623_b1 , \623_b0 , \624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , \627_b1 , \627_b0 , 
		\628_b1 , \628_b0 , \629_b1 , \629_b0 , \630_SUM[16]_b1 , \630_SUM[16]_b0 , \631_b1 , \631_b0 , \632_A[16]_b1 , \632_A[16]_b0 , 
		\633_B[16]_b1 , \633_B[16]_b0 , \634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , \637_b1 , \637_b0 , 
		\638_b1 , \638_b0 , \639_b1 , \639_b0 , \640_SUM[16]_b1 , \640_SUM[16]_b0 , \641_b1 , \641_b0 , \642_n5[17]_b1 , \642_n5[17]_b0 , 
		\643_b1 , \643_b0 , \644_A[17]_b1 , \644_A[17]_b0 , \645_B[17]_b1 , \645_B[17]_b0 , \646_b1 , \646_b0 , \647_b1 , \647_b0 , 
		\648_b1 , \648_b0 , \649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , \652_b1 , \652_b0 , 
		\653_SUM[17]_b1 , \653_SUM[17]_b0 , \654_b1 , \654_b0 , \655_A[17]_b1 , \655_A[17]_b0 , \656_B[17]_b1 , \656_B[17]_b0 , \657_b1 , \657_b0 , 
		\658_b1 , \658_b0 , \659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , \662_b1 , \662_b0 , 
		\663_SUM[17]_b1 , \663_SUM[17]_b0 , \664_b1 , \664_b0 , \665_n5[18]_b1 , \665_n5[18]_b0 , \666_b1 , \666_b0 , \667_A[18]_b1 , \667_A[18]_b0 , 
		\668_B[18]_b1 , \668_B[18]_b0 , \669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , \672_b1 , \672_b0 , 
		\673_b1 , \673_b0 , \674_b1 , \674_b0 , \675_b1 , \675_b0 , \676_SUM[18]_b1 , \676_SUM[18]_b0 , \677_b1 , \677_b0 , 
		\678_A[18]_b1 , \678_A[18]_b0 , \679_B[18]_b1 , \679_B[18]_b0 , \680_b1 , \680_b0 , \681_b1 , \681_b0 , \682_b1 , \682_b0 , 
		\683_b1 , \683_b0 , \684_b1 , \684_b0 , \685_b1 , \685_b0 , \686_SUM[18]_b1 , \686_SUM[18]_b0 , \687_b1 , \687_b0 , 
		\688_n5[19]_b1 , \688_n5[19]_b0 , \689_b1 , \689_b0 , \690_A[19]_b1 , \690_A[19]_b0 , \691_B[19]_b1 , \691_B[19]_b0 , \692_b1 , \692_b0 , 
		\693_b1 , \693_b0 , \694_b1 , \694_b0 , \695_b1 , \695_b0 , \696_b1 , \696_b0 , \697_b1 , \697_b0 , 
		\698_b1 , \698_b0 , \699_SUM[19]_b1 , \699_SUM[19]_b0 , \700_b1 , \700_b0 , \701_A[19]_b1 , \701_A[19]_b0 , \702_B[19]_b1 , \702_B[19]_b0 , 
		\703_b1 , \703_b0 , \704_b1 , \704_b0 , \705_b1 , \705_b0 , \706_b1 , \706_b0 , \707_b1 , \707_b0 , 
		\708_b1 , \708_b0 , \709_SUM[19]_b1 , \709_SUM[19]_b0 , \710_b1 , \710_b0 , \711_n5[20]_b1 , \711_n5[20]_b0 , \712_b1 , \712_b0 , 
		\713_A[20]_b1 , \713_A[20]_b0 , \714_B[20]_b1 , \714_B[20]_b0 , \715_b1 , \715_b0 , \716_b1 , \716_b0 , \717_b1 , \717_b0 , 
		\718_b1 , \718_b0 , \719_b1 , \719_b0 , \720_b1 , \720_b0 , \721_b1 , \721_b0 , \722_SUM[20]_b1 , \722_SUM[20]_b0 , 
		\723_b1 , \723_b0 , \724_A[20]_b1 , \724_A[20]_b0 , \725_B[20]_b1 , \725_B[20]_b0 , \726_b1 , \726_b0 , \727_b1 , \727_b0 , 
		\728_b1 , \728_b0 , \729_b1 , \729_b0 , \730_b1 , \730_b0 , \731_b1 , \731_b0 , \732_SUM[20]_b1 , \732_SUM[20]_b0 , 
		\733_b1 , \733_b0 , \734_n5[21]_b1 , \734_n5[21]_b0 , \735_b1 , \735_b0 , \736_A[21]_b1 , \736_A[21]_b0 , \737_B[21]_b1 , \737_B[21]_b0 , 
		\738_b1 , \738_b0 , \739_b1 , \739_b0 , \740_b1 , \740_b0 , \741_b1 , \741_b0 , \742_b1 , \742_b0 , 
		\743_b1 , \743_b0 , \744_b1 , \744_b0 , \745_SUM[21]_b1 , \745_SUM[21]_b0 , \746_b1 , \746_b0 , \747_A[21]_b1 , \747_A[21]_b0 , 
		\748_B[21]_b1 , \748_B[21]_b0 , \749_b1 , \749_b0 , \750_b1 , \750_b0 , \751_b1 , \751_b0 , \752_b1 , \752_b0 , 
		\753_b1 , \753_b0 , \754_b1 , \754_b0 , \755_SUM[21]_b1 , \755_SUM[21]_b0 , \756_b1 , \756_b0 , \757_n5[22]_b1 , \757_n5[22]_b0 , 
		\758_b1 , \758_b0 , \759_A[22]_b1 , \759_A[22]_b0 , \760_B[22]_b1 , \760_B[22]_b0 , \761_b1 , \761_b0 , \762_b1 , \762_b0 , 
		\763_b1 , \763_b0 , \764_b1 , \764_b0 , \765_b1 , \765_b0 , \766_b1 , \766_b0 , \767_b1 , \767_b0 , 
		\768_SUM[22]_b1 , \768_SUM[22]_b0 , \769_b1 , \769_b0 , \770_A[22]_b1 , \770_A[22]_b0 , \771_B[22]_b1 , \771_B[22]_b0 , \772_b1 , \772_b0 , 
		\773_b1 , \773_b0 , \774_b1 , \774_b0 , \775_b1 , \775_b0 , \776_b1 , \776_b0 , \777_b1 , \777_b0 , 
		\778_SUM[22]_b1 , \778_SUM[22]_b0 , \779_b1 , \779_b0 , \780_n5[23]_b1 , \780_n5[23]_b0 , \781_b1 , \781_b0 , \782_A[23]_b1 , \782_A[23]_b0 , 
		\783_B[23]_b1 , \783_B[23]_b0 , \784_b1 , \784_b0 , \785_b1 , \785_b0 , \786_b1 , \786_b0 , \787_b1 , \787_b0 , 
		\788_b1 , \788_b0 , \789_b1 , \789_b0 , \790_b1 , \790_b0 , \791_SUM[23]_b1 , \791_SUM[23]_b0 , \792_b1 , \792_b0 , 
		\793_A[23]_b1 , \793_A[23]_b0 , \794_B[23]_b1 , \794_B[23]_b0 , \795_b1 , \795_b0 , \796_b1 , \796_b0 , \797_b1 , \797_b0 , 
		\798_b1 , \798_b0 , \799_b1 , \799_b0 , \800_b1 , \800_b0 , \801_SUM[23]_b1 , \801_SUM[23]_b0 , \802_b1 , \802_b0 , 
		\803_n5[24]_b1 , \803_n5[24]_b0 , \804_b1 , \804_b0 , \805_A[24]_b1 , \805_A[24]_b0 , \806_B[24]_b1 , \806_B[24]_b0 , \807_b1 , \807_b0 , 
		\808_b1 , \808_b0 , \809_b1 , \809_b0 , \810_b1 , \810_b0 , \811_b1 , \811_b0 , \812_b1 , \812_b0 , 
		\813_b1 , \813_b0 , \814_SUM[24]_b1 , \814_SUM[24]_b0 , \815_b1 , \815_b0 , \816_A[24]_b1 , \816_A[24]_b0 , \817_B[24]_b1 , \817_B[24]_b0 , 
		\818_b1 , \818_b0 , \819_b1 , \819_b0 , \820_b1 , \820_b0 , \821_b1 , \821_b0 , \822_b1 , \822_b0 , 
		\823_b1 , \823_b0 , \824_SUM[24]_b1 , \824_SUM[24]_b0 , \825_b1 , \825_b0 , \826_n5[25]_b1 , \826_n5[25]_b0 , \827_b1 , \827_b0 , 
		\828_A[25]_b1 , \828_A[25]_b0 , \829_B[25]_b1 , \829_B[25]_b0 , \830_b1 , \830_b0 , \831_b1 , \831_b0 , \832_b1 , \832_b0 , 
		\833_b1 , \833_b0 , \834_b1 , \834_b0 , \835_b1 , \835_b0 , \836_b1 , \836_b0 , \837_SUM[25]_b1 , \837_SUM[25]_b0 , 
		\838_b1 , \838_b0 , \839_A[25]_b1 , \839_A[25]_b0 , \840_B[25]_b1 , \840_B[25]_b0 , \841_b1 , \841_b0 , \842_b1 , \842_b0 , 
		\843_b1 , \843_b0 , \844_b1 , \844_b0 , \845_b1 , \845_b0 , \846_b1 , \846_b0 , \847_SUM[25]_b1 , \847_SUM[25]_b0 , 
		\848_b1 , \848_b0 , \849_n5[26]_b1 , \849_n5[26]_b0 , \850_b1 , \850_b0 , \851_A[26]_b1 , \851_A[26]_b0 , \852_B[26]_b1 , \852_B[26]_b0 , 
		\853_b1 , \853_b0 , \854_b1 , \854_b0 , \855_b1 , \855_b0 , \856_b1 , \856_b0 , \857_b1 , \857_b0 , 
		\858_b1 , \858_b0 , \859_b1 , \859_b0 , \860_SUM[26]_b1 , \860_SUM[26]_b0 , \861_b1 , \861_b0 , \862_A[26]_b1 , \862_A[26]_b0 , 
		\863_B[26]_b1 , \863_B[26]_b0 , \864_b1 , \864_b0 , \865_b1 , \865_b0 , \866_b1 , \866_b0 , \867_b1 , \867_b0 , 
		\868_b1 , \868_b0 , \869_b1 , \869_b0 , \870_SUM[26]_b1 , \870_SUM[26]_b0 , \871_b1 , \871_b0 , \872_n5[27]_b1 , \872_n5[27]_b0 , 
		\873_b1 , \873_b0 , \874_A[27]_b1 , \874_A[27]_b0 , \875_B[27]_b1 , \875_B[27]_b0 , \876_b1 , \876_b0 , \877_b1 , \877_b0 , 
		\878_b1 , \878_b0 , \879_b1 , \879_b0 , \880_b1 , \880_b0 , \881_b1 , \881_b0 , \882_b1 , \882_b0 , 
		\883_SUM[27]_b1 , \883_SUM[27]_b0 , \884_b1 , \884_b0 , \885_A[27]_b1 , \885_A[27]_b0 , \886_B[27]_b1 , \886_B[27]_b0 , \887_b1 , \887_b0 , 
		\888_b1 , \888_b0 , \889_b1 , \889_b0 , \890_b1 , \890_b0 , \891_b1 , \891_b0 , \892_b1 , \892_b0 , 
		\893_SUM[27]_b1 , \893_SUM[27]_b0 , \894_b1 , \894_b0 , \895_n5[28]_b1 , \895_n5[28]_b0 , \896_b1 , \896_b0 , \897_A[28]_b1 , \897_A[28]_b0 , 
		\898_B[28]_b1 , \898_B[28]_b0 , \899_b1 , \899_b0 , \900_b1 , \900_b0 , \901_b1 , \901_b0 , \902_b1 , \902_b0 , 
		\903_b1 , \903_b0 , \904_b1 , \904_b0 , \905_b1 , \905_b0 , \906_SUM[28]_b1 , \906_SUM[28]_b0 , \907_b1 , \907_b0 , 
		\908_A[28]_b1 , \908_A[28]_b0 , \909_B[28]_b1 , \909_B[28]_b0 , \910_b1 , \910_b0 , \911_b1 , \911_b0 , \912_b1 , \912_b0 , 
		\913_b1 , \913_b0 , \914_b1 , \914_b0 , \915_b1 , \915_b0 , \916_SUM[28]_b1 , \916_SUM[28]_b0 , \917_b1 , \917_b0 , 
		\918_n5[29]_b1 , \918_n5[29]_b0 , \919_b1 , \919_b0 , \920_A[29]_b1 , \920_A[29]_b0 , \921_B[29]_b1 , \921_B[29]_b0 , \922_b1 , \922_b0 , 
		\923_b1 , \923_b0 , \924_b1 , \924_b0 , \925_b1 , \925_b0 , \926_b1 , \926_b0 , \927_b1 , \927_b0 , 
		\928_b1 , \928_b0 , \929_SUM[29]_b1 , \929_SUM[29]_b0 , \930_b1 , \930_b0 , \931_A[29]_b1 , \931_A[29]_b0 , \932_B[29]_b1 , \932_B[29]_b0 , 
		\933_b1 , \933_b0 , \934_b1 , \934_b0 , \935_b1 , \935_b0 , \936_b1 , \936_b0 , \937_b1 , \937_b0 , 
		\938_b1 , \938_b0 , \939_SUM[29]_b1 , \939_SUM[29]_b0 , \940_b1 , \940_b0 , \941_n5[30]_b1 , \941_n5[30]_b0 , \942_b1 , \942_b0 , 
		\943_A[30]_b1 , \943_A[30]_b0 , \944_B[30]_b1 , \944_B[30]_b0 , \945_b1 , \945_b0 , \946_b1 , \946_b0 , \947_b1 , \947_b0 , 
		\948_b1 , \948_b0 , \949_b1 , \949_b0 , \950_b1 , \950_b0 , \951_b1 , \951_b0 , \952_SUM[30]_b1 , \952_SUM[30]_b0 , 
		\953_b1 , \953_b0 , \954_A[30]_b1 , \954_A[30]_b0 , \955_B[30]_b1 , \955_B[30]_b0 , \956_b1 , \956_b0 , \957_b1 , \957_b0 , 
		\958_b1 , \958_b0 , \959_b1 , \959_b0 , \960_b1 , \960_b0 , \961_b1 , \961_b0 , \962_SUM[30]_b1 , \962_SUM[30]_b0 , 
		\963_b1 , \963_b0 , \964_n5[31]_b1 , \964_n5[31]_b0 , \965_b1 , \965_b0 , \966_A[31]_b1 , \966_A[31]_b0 , \967_B[31]_b1 , \967_B[31]_b0 , 
		\968_b1 , \968_b0 , \969_b1 , \969_b0 , \970_b1 , \970_b0 , \971_b1 , \971_b0 , \972_b1 , \972_b0 , 
		\973_b1 , \973_b0 , \974_b1 , \974_b0 , \975_SUM[31]_b1 , \975_SUM[31]_b0 , \976_b1 , \976_b0 , \977_A[31]_b1 , \977_A[31]_b0 , 
		\978_B[31]_b1 , \978_B[31]_b0 , \979_b1 , \979_b0 , \980_b1 , \980_b0 , \981_b1 , \981_b0 , \982_b1 , \982_b0 , 
		\983_b1 , \983_b0 , \984_b1 , \984_b0 , \985_SUM[31]_b1 , \985_SUM[31]_b0 , \986_b1 , \986_b0 , \987_A[31]_b1 , \987_A[31]_b0 , 
		\988_B[31]_b1 , \988_B[31]_b0 , \989_b1 , \989_b0 , \990_A[30]_b1 , \990_A[30]_b0 , \991_B[30]_b1 , \991_B[30]_b0 , \992_b1 , \992_b0 , 
		\993_A[29]_b1 , \993_A[29]_b0 , \994_B[29]_b1 , \994_B[29]_b0 , \995_b1 , \995_b0 , \996_A[28]_b1 , \996_A[28]_b0 , \997_B[28]_b1 , \997_B[28]_b0 , 
		\998_b1 , \998_b0 , \999_A[27]_b1 , \999_A[27]_b0 , \1000_B[27]_b1 , \1000_B[27]_b0 , \1001_b1 , \1001_b0 , \1002_A[26]_b1 , \1002_A[26]_b0 , 
		\1003_B[26]_b1 , \1003_B[26]_b0 , \1004_b1 , \1004_b0 , \1005_A[25]_b1 , \1005_A[25]_b0 , \1006_B[25]_b1 , \1006_B[25]_b0 , \1007_b1 , \1007_b0 , 
		\1008_A[24]_b1 , \1008_A[24]_b0 , \1009_B[24]_b1 , \1009_B[24]_b0 , \1010_b1 , \1010_b0 , \1011_A[23]_b1 , \1011_A[23]_b0 , \1012_B[23]_b1 , \1012_B[23]_b0 , 
		\1013_b1 , \1013_b0 , \1014_A[22]_b1 , \1014_A[22]_b0 , \1015_B[22]_b1 , \1015_B[22]_b0 , \1016_b1 , \1016_b0 , \1017_A[21]_b1 , \1017_A[21]_b0 , 
		\1018_B[21]_b1 , \1018_B[21]_b0 , \1019_b1 , \1019_b0 , \1020_A[20]_b1 , \1020_A[20]_b0 , \1021_B[20]_b1 , \1021_B[20]_b0 , \1022_b1 , \1022_b0 , 
		\1023_A[19]_b1 , \1023_A[19]_b0 , \1024_B[19]_b1 , \1024_B[19]_b0 , \1025_b1 , \1025_b0 , \1026_A[18]_b1 , \1026_A[18]_b0 , \1027_B[18]_b1 , \1027_B[18]_b0 , 
		\1028_b1 , \1028_b0 , \1029_A[17]_b1 , \1029_A[17]_b0 , \1030_B[17]_b1 , \1030_B[17]_b0 , \1031_b1 , \1031_b0 , \1032_A[16]_b1 , \1032_A[16]_b0 , 
		\1033_B[16]_b1 , \1033_B[16]_b0 , \1034_b1 , \1034_b0 , \1035_A[15]_b1 , \1035_A[15]_b0 , \1036_B[15]_b1 , \1036_B[15]_b0 , \1037_b1 , \1037_b0 , 
		\1038_A[14]_b1 , \1038_A[14]_b0 , \1039_B[14]_b1 , \1039_B[14]_b0 , \1040_b1 , \1040_b0 , \1041_A[13]_b1 , \1041_A[13]_b0 , \1042_B[13]_b1 , \1042_B[13]_b0 , 
		\1043_b1 , \1043_b0 , \1044_A[12]_b1 , \1044_A[12]_b0 , \1045_B[12]_b1 , \1045_B[12]_b0 , \1046_b1 , \1046_b0 , \1047_A[11]_b1 , \1047_A[11]_b0 , 
		\1048_B[11]_b1 , \1048_B[11]_b0 , \1049_b1 , \1049_b0 , \1050_A[10]_b1 , \1050_A[10]_b0 , \1051_B[10]_b1 , \1051_B[10]_b0 , \1052_b1 , \1052_b0 , 
		\1053_A[9]_b1 , \1053_A[9]_b0 , \1054_B[9]_b1 , \1054_B[9]_b0 , \1055_b1 , \1055_b0 , \1056_A[8]_b1 , \1056_A[8]_b0 , \1057_B[8]_b1 , \1057_B[8]_b0 , 
		\1058_b1 , \1058_b0 , \1059_A[7]_b1 , \1059_A[7]_b0 , \1060_B[7]_b1 , \1060_B[7]_b0 , \1061_b1 , \1061_b0 , \1062_A[6]_b1 , \1062_A[6]_b0 , 
		\1063_B[6]_b1 , \1063_B[6]_b0 , \1064_b1 , \1064_b0 , \1065_A[5]_b1 , \1065_A[5]_b0 , \1066_B[5]_b1 , \1066_B[5]_b0 , \1067_b1 , \1067_b0 , 
		\1068_A[4]_b1 , \1068_A[4]_b0 , \1069_B[4]_b1 , \1069_B[4]_b0 , \1070_b1 , \1070_b0 , \1071_A[3]_b1 , \1071_A[3]_b0 , \1072_B[3]_b1 , \1072_B[3]_b0 , 
		\1073_b1 , \1073_b0 , \1074_A[2]_b1 , \1074_A[2]_b0 , \1075_B[2]_b1 , \1075_B[2]_b0 , \1076_b1 , \1076_b0 , \1077_A[1]_b1 , \1077_A[1]_b0 , 
		\1078_B[1]_b1 , \1078_B[1]_b0 , \1079_b1 , \1079_b0 , \1080_A[0]_b1 , \1080_A[0]_b0 , \1081_B[0]_b1 , \1081_B[0]_b0 , \1082_b1 , \1082_b0 , 
		\1083_b1 , \1083_b0 , \1084_b1 , \1084_b0 , \1085_b1 , \1085_b0 , \1086_b1 , \1086_b0 , \1087_b1 , \1087_b0 , 
		\1088_b1 , \1088_b0 , \1089_b1 , \1089_b0 , \1090_b1 , \1090_b0 , \1091_b1 , \1091_b0 , \1092_b1 , \1092_b0 , 
		\1093_b1 , \1093_b0 , \1094_b1 , \1094_b0 , \1095_b1 , \1095_b0 , \1096_b1 , \1096_b0 , \1097_b1 , \1097_b0 , 
		\1098_b1 , \1098_b0 , \1099_b1 , \1099_b0 , \1100_b1 , \1100_b0 , \1101_b1 , \1101_b0 , \1102_b1 , \1102_b0 , 
		\1103_b1 , \1103_b0 , \1104_b1 , \1104_b0 , \1105_b1 , \1105_b0 , \1106_b1 , \1106_b0 , \1107_b1 , \1107_b0 , 
		\1108_b1 , \1108_b0 , \1109_b1 , \1109_b0 , \1110_b1 , \1110_b0 , \1111_b1 , \1111_b0 , \1112_b1 , \1112_b0 , 
		\1113_b1 , \1113_b0 , \1114_b1 , \1114_b0 , \1115_b1 , \1115_b0 , \1116_b1 , \1116_b0 , \1117_b1 , \1117_b0 , 
		\1118_b1 , \1118_b0 , \1119_b1 , \1119_b0 , \1120_b1 , \1120_b0 , \1121_b1 , \1121_b0 , \1122_b1 , \1122_b0 , 
		\1123_b1 , \1123_b0 , \1124_b1 , \1124_b0 , \1125_b1 , \1125_b0 , \1126_b1 , \1126_b0 , \1127_b1 , \1127_b0 , 
		\1128_b1 , \1128_b0 , \1129_b1 , \1129_b0 , \1130_b1 , \1130_b0 , \1131_b1 , \1131_b0 , \1132_b1 , \1132_b0 , 
		\1133_b1 , \1133_b0 , \1134_b1 , \1134_b0 , \1135_b1 , \1135_b0 , \1136_b1 , \1136_b0 , \1137_b1 , \1137_b0 , 
		\1138_b1 , \1138_b0 , \1139_b1 , \1139_b0 , \1140_b1 , \1140_b0 , \1141_b1 , \1141_b0 , \1142_b1 , \1142_b0 , 
		\1143_b1 , \1143_b0 , \1144_b1 , \1144_b0 , \1145_b1 , \1145_b0 , \1146_b1 , \1146_b0 , \1147_b1 , \1147_b0 , 
		\1148_b1 , \1148_b0 , \1149_b1 , \1149_b0 , \1150_b1 , \1150_b0 , \1151_b1 , \1151_b0 , \1152_b1 , \1152_b0 , 
		\1153_b1 , \1153_b0 , \1154_b1 , \1154_b0 , \1155_b1 , \1155_b0 , \1156_b1 , \1156_b0 , \1157_b1 , \1157_b0 , 
		\1158_b1 , \1158_b0 , \1159_b1 , \1159_b0 , \1160_b1 , \1160_b0 , \1161_b1 , \1161_b0 , \1162_b1 , \1162_b0 , 
		\1163_b1 , \1163_b0 , \1164_b1 , \1164_b0 , \1165_b1 , \1165_b0 , \1166_b1 , \1166_b0 , \1167_b1 , \1167_b0 , 
		\1168_b1 , \1168_b0 , \1169_b1 , \1169_b0 , \1170_b1 , \1170_b0 , \1171_b1 , \1171_b0 , \1172_b1 , \1172_b0 , 
		\1173_b1 , \1173_b0 , \1174_SUM[31]_b1 , \1174_SUM[31]_b0 , \1175_A[31]_b1 , \1175_A[31]_b0 , \1176_b1 , \1176_b0 , \1177_b1 , \1177_b0 , 
		\1178_SUM[30]_b1 , \1178_SUM[30]_b0 , \1179_A[30]_b1 , \1179_A[30]_b0 , \1180_b1 , \1180_b0 , \1181_b1 , \1181_b0 , \1182_SUM[29]_b1 , \1182_SUM[29]_b0 , 
		\1183_A[29]_b1 , \1183_A[29]_b0 , \1184_b1 , \1184_b0 , \1185_b1 , \1185_b0 , \1186_SUM[28]_b1 , \1186_SUM[28]_b0 , \1187_A[28]_b1 , \1187_A[28]_b0 , 
		\1188_b1 , \1188_b0 , \1189_b1 , \1189_b0 , \1190_SUM[27]_b1 , \1190_SUM[27]_b0 , \1191_A[27]_b1 , \1191_A[27]_b0 , \1192_b1 , \1192_b0 , 
		\1193_b1 , \1193_b0 , \1194_SUM[26]_b1 , \1194_SUM[26]_b0 , \1195_A[26]_b1 , \1195_A[26]_b0 , \1196_b1 , \1196_b0 , \1197_b1 , \1197_b0 , 
		\1198_SUM[25]_b1 , \1198_SUM[25]_b0 , \1199_A[25]_b1 , \1199_A[25]_b0 , \1200_b1 , \1200_b0 , \1201_b1 , \1201_b0 , \1202_SUM[24]_b1 , \1202_SUM[24]_b0 , 
		\1203_A[24]_b1 , \1203_A[24]_b0 , \1204_b1 , \1204_b0 , \1205_b1 , \1205_b0 , \1206_SUM[23]_b1 , \1206_SUM[23]_b0 , \1207_A[23]_b1 , \1207_A[23]_b0 , 
		\1208_b1 , \1208_b0 , \1209_b1 , \1209_b0 , \1210_SUM[22]_b1 , \1210_SUM[22]_b0 , \1211_A[22]_b1 , \1211_A[22]_b0 , \1212_b1 , \1212_b0 , 
		\1213_b1 , \1213_b0 , \1214_SUM[21]_b1 , \1214_SUM[21]_b0 , \1215_A[21]_b1 , \1215_A[21]_b0 , \1216_b1 , \1216_b0 , \1217_b1 , \1217_b0 , 
		\1218_SUM[20]_b1 , \1218_SUM[20]_b0 , \1219_A[20]_b1 , \1219_A[20]_b0 , \1220_b1 , \1220_b0 , \1221_b1 , \1221_b0 , \1222_SUM[19]_b1 , \1222_SUM[19]_b0 , 
		\1223_A[19]_b1 , \1223_A[19]_b0 , \1224_b1 , \1224_b0 , \1225_b1 , \1225_b0 , \1226_SUM[18]_b1 , \1226_SUM[18]_b0 , \1227_A[18]_b1 , \1227_A[18]_b0 , 
		\1228_b1 , \1228_b0 , \1229_b1 , \1229_b0 , \1230_SUM[17]_b1 , \1230_SUM[17]_b0 , \1231_A[17]_b1 , \1231_A[17]_b0 , \1232_b1 , \1232_b0 , 
		\1233_b1 , \1233_b0 , \1234_SUM[16]_b1 , \1234_SUM[16]_b0 , \1235_A[16]_b1 , \1235_A[16]_b0 , \1236_b1 , \1236_b0 , \1237_b1 , \1237_b0 , 
		\1238_SUM[15]_b1 , \1238_SUM[15]_b0 , \1239_A[15]_b1 , \1239_A[15]_b0 , \1240_b1 , \1240_b0 , \1241_b1 , \1241_b0 , \1242_SUM[14]_b1 , \1242_SUM[14]_b0 , 
		\1243_A[14]_b1 , \1243_A[14]_b0 , \1244_b1 , \1244_b0 , \1245_b1 , \1245_b0 , \1246_SUM[13]_b1 , \1246_SUM[13]_b0 , \1247_A[13]_b1 , \1247_A[13]_b0 , 
		\1248_b1 , \1248_b0 , \1249_b1 , \1249_b0 , \1250_SUM[12]_b1 , \1250_SUM[12]_b0 , \1251_A[12]_b1 , \1251_A[12]_b0 , \1252_b1 , \1252_b0 , 
		\1253_b1 , \1253_b0 , \1254_SUM[11]_b1 , \1254_SUM[11]_b0 , \1255_A[11]_b1 , \1255_A[11]_b0 , \1256_b1 , \1256_b0 , \1257_b1 , \1257_b0 , 
		\1258_SUM[10]_b1 , \1258_SUM[10]_b0 , \1259_A[10]_b1 , \1259_A[10]_b0 , \1260_b1 , \1260_b0 , \1261_b1 , \1261_b0 , \1262_SUM[9]_b1 , \1262_SUM[9]_b0 , 
		\1263_A[9]_b1 , \1263_A[9]_b0 , \1264_b1 , \1264_b0 , \1265_b1 , \1265_b0 , \1266_SUM[8]_b1 , \1266_SUM[8]_b0 , \1267_A[8]_b1 , \1267_A[8]_b0 , 
		\1268_b1 , \1268_b0 , \1269_b1 , \1269_b0 , \1270_SUM[7]_b1 , \1270_SUM[7]_b0 , \1271_A[7]_b1 , \1271_A[7]_b0 , \1272_b1 , \1272_b0 , 
		\1273_b1 , \1273_b0 , \1274_SUM[6]_b1 , \1274_SUM[6]_b0 , \1275_A[6]_b1 , \1275_A[6]_b0 , \1276_b1 , \1276_b0 , \1277_b1 , \1277_b0 , 
		\1278_SUM[5]_b1 , \1278_SUM[5]_b0 , \1279_A[5]_b1 , \1279_A[5]_b0 , \1280_b1 , \1280_b0 , \1281_b1 , \1281_b0 , \1282_SUM[4]_b1 , \1282_SUM[4]_b0 , 
		\1283_A[4]_b1 , \1283_A[4]_b0 , \1284_b1 , \1284_b0 , \1285_b1 , \1285_b0 , \1286_SUM[3]_b1 , \1286_SUM[3]_b0 , \1287_A[3]_b1 , \1287_A[3]_b0 , 
		\1288_b1 , \1288_b0 , \1289_b1 , \1289_b0 , \1290_SUM[2]_b1 , \1290_SUM[2]_b0 , \1291_A[2]_b1 , \1291_A[2]_b0 , \1292_b1 , \1292_b0 , 
		\1293_b1 , \1293_b0 , \1294_SUM[1]_b1 , \1294_SUM[1]_b0 , \1295_A[1]_b1 , \1295_A[1]_b0 , \1296_b1 , \1296_b0 , \1297_SUM[0]_b1 , \1297_SUM[0]_b0 , 
		\1298_A[0]_b1 , \1298_A[0]_b0 , \1299_B[31]_b1 , \1299_B[31]_b0 , \1300_B[30]_b1 , \1300_B[30]_b0 , \1301_B[29]_b1 , \1301_B[29]_b0 , \1302_B[28]_b1 , \1302_B[28]_b0 , 
		\1303_B[27]_b1 , \1303_B[27]_b0 , \1304_B[26]_b1 , \1304_B[26]_b0 , \1305_B[25]_b1 , \1305_B[25]_b0 , \1306_B[24]_b1 , \1306_B[24]_b0 , \1307_B[23]_b1 , \1307_B[23]_b0 , 
		\1308_B[22]_b1 , \1308_B[22]_b0 , \1309_B[21]_b1 , \1309_B[21]_b0 , \1310_B[20]_b1 , \1310_B[20]_b0 , \1311_B[19]_b1 , \1311_B[19]_b0 , \1312_B[18]_b1 , \1312_B[18]_b0 , 
		\1313_B[17]_b1 , \1313_B[17]_b0 , \1314_B[16]_b1 , \1314_B[16]_b0 , \1315_B[15]_b1 , \1315_B[15]_b0 , \1316_B[14]_b1 , \1316_B[14]_b0 , \1317_B[13]_b1 , \1317_B[13]_b0 , 
		\1318_B[12]_b1 , \1318_B[12]_b0 , \1319_B[11]_b1 , \1319_B[11]_b0 , \1320_B[10]_b1 , \1320_B[10]_b0 , \1321_B[9]_b1 , \1321_B[9]_b0 , \1322_B[8]_b1 , \1322_B[8]_b0 , 
		\1323_B[7]_b1 , \1323_B[7]_b0 , \1324_B[6]_b1 , \1324_B[6]_b0 , \1325_B[5]_b1 , \1325_B[5]_b0 , \1326_B[4]_b1 , \1326_B[4]_b0 , \1327_B[3]_b1 , \1327_B[3]_b0 , 
		\1328_B[2]_b1 , \1328_B[2]_b0 , \1329_B[1]_b1 , \1329_B[1]_b0 , \1330_B[0]_b1 , \1330_B[0]_b0 , \1331_b1 , \1331_b0 , \1332_b1 , \1332_b0 , 
		\1333_b1 , \1333_b0 , \1334_b1 , \1334_b0 , \1335_b1 , \1335_b0 , \1336_b1 , \1336_b0 , \1337_b1 , \1337_b0 , 
		\1338_b1 , \1338_b0 , \1339_b1 , \1339_b0 , \1340_b1 , \1340_b0 , \1341_b1 , \1341_b0 , \1342_b1 , \1342_b0 , 
		\1343_b1 , \1343_b0 , \1344_b1 , \1344_b0 , \1345_b1 , \1345_b0 , \1346_b1 , \1346_b0 , \1347_b1 , \1347_b0 , 
		\1348_b1 , \1348_b0 , \1349_b1 , \1349_b0 , \1350_b1 , \1350_b0 , \1351_b1 , \1351_b0 , \1352_b1 , \1352_b0 , 
		\1353_b1 , \1353_b0 , \1354_b1 , \1354_b0 , \1355_b1 , \1355_b0 , \1356_b1 , \1356_b0 , \1357_b1 , \1357_b0 , 
		\1358_b1 , \1358_b0 , \1359_b1 , \1359_b0 , \1360_b1 , \1360_b0 , \1361_b1 , \1361_b0 , \1362_b1 , \1362_b0 , 
		\1363_b1 , \1363_b0 , \1364_b1 , \1364_b0 , \1365_b1 , \1365_b0 , \1366_b1 , \1366_b0 , \1367_b1 , \1367_b0 , 
		\1368_b1 , \1368_b0 , \1369_b1 , \1369_b0 , \1370_b1 , \1370_b0 , \1371_b1 , \1371_b0 , \1372_b1 , \1372_b0 , 
		\1373_b1 , \1373_b0 , \1374_b1 , \1374_b0 , \1375_b1 , \1375_b0 , \1376_b1 , \1376_b0 , \1377_b1 , \1377_b0 , 
		\1378_b1 , \1378_b0 , \1379_b1 , \1379_b0 , \1380_b1 , \1380_b0 , \1381_b1 , \1381_b0 , \1382_b1 , \1382_b0 , 
		\1383_b1 , \1383_b0 , \1384_b1 , \1384_b0 , \1385_b1 , \1385_b0 , \1386_b1 , \1386_b0 , \1387_b1 , \1387_b0 , 
		\1388_b1 , \1388_b0 , \1389_b1 , \1389_b0 , \1390_b1 , \1390_b0 , \1391_b1 , \1391_b0 , \1392_b1 , \1392_b0 , 
		\1393_b1 , \1393_b0 , \1394_b1 , \1394_b0 , \1395_b1 , \1395_b0 , \1396_b1 , \1396_b0 , \1397_b1 , \1397_b0 , 
		\1398_b1 , \1398_b0 , \1399_b1 , \1399_b0 , \1400_b1 , \1400_b0 , \1401_b1 , \1401_b0 , \1402_b1 , \1402_b0 , 
		\1403_b1 , \1403_b0 , \1404_b1 , \1404_b0 , \1405_b1 , \1405_b0 , \1406_b1 , \1406_b0 , \1407_b1 , \1407_b0 , 
		\1408_b1 , \1408_b0 , \1409_b1 , \1409_b0 , \1410_b1 , \1410_b0 , \1411_b1 , \1411_b0 , \1412_b1 , \1412_b0 , 
		\1413_b1 , \1413_b0 , \1414_b1 , \1414_b0 , \1415_b1 , \1415_b0 , \1416_b1 , \1416_b0 , \1417_b1 , \1417_b0 , 
		\1418_b1 , \1418_b0 , \1419_b1 , \1419_b0 , \1420_b1 , \1420_b0 , \1421_b1 , \1421_b0 , \1422_b1 , \1422_b0 , 
		\1423_b1 , \1423_b0 , \1424_b1 , \1424_b0 , \1425_b1 , \1425_b0 , \1426_b1 , \1426_b0 , \1427_b1 , \1427_b0 , 
		\1428_b1 , \1428_b0 , \1429_b1 , \1429_b0 , \1430_b1 , \1430_b0 , \1431_b1 , \1431_b0 , \1432_b1 , \1432_b0 , 
		\1433_b1 , \1433_b0 , \1434_b1 , \1434_b0 , \1435_b1 , \1435_b0 , \1436_b1 , \1436_b0 , \1437_b1 , \1437_b0 , 
		\1438_b1 , \1438_b0 , \1439_b1 , \1439_b0 , \1440_b1 , \1440_b0 , \1441_b1 , \1441_b0 , \1442_b1 , \1442_b0 , 
		\1443_b1 , \1443_b0 , \1444_b1 , \1444_b0 , \1445_b1 , \1445_b0 , \1446_b1 , \1446_b0 , \1447_b1 , \1447_b0 , 
		\1448_b1 , \1448_b0 , \1449_b1 , \1449_b0 , \1450_b1 , \1450_b0 , \1451_b1 , \1451_b0 , \1452_b1 , \1452_b0 , 
		\1453_b1 , \1453_b0 , \1454_b1 , \1454_b0 , \1455_b1 , \1455_b0 , \1456_b1 , \1456_b0 , \1457_b1 , \1457_b0 , 
		\1458_b1 , \1458_b0 , \1459_b1 , \1459_b0 , \1460_b1 , \1460_b0 , \1461_b1 , \1461_b0 , \1462_b1 , \1462_b0 , 
		\1463_b1 , \1463_b0 , \1464_b1 , \1464_b0 , \1465_b1 , \1465_b0 , \1466_b1 , \1466_b0 , \1467_b1 , \1467_b0 , 
		\1468_b1 , \1468_b0 , \1469_b1 , \1469_b0 , \1470_b1 , \1470_b0 , \1471_b1 , \1471_b0 , \1472_b1 , \1472_b0 , 
		\1473_b1 , \1473_b0 , \1474_b1 , \1474_b0 , \1475_b1 , \1475_b0 , \1476_b1 , \1476_b0 , \1477_b1 , \1477_b0 , 
		\1478_b1 , \1478_b0 , \1479_b1 , \1479_b0 , \1480_b1 , \1480_b0 , \1481_b1 , \1481_b0 , \1482_b1 , \1482_b0 , 
		\1483_b1 , \1483_b0 , \1484_b1 , \1484_b0 , \1485_b1 , \1485_b0 , \1486_b1 , \1486_b0 , \1487_b1 , \1487_b0 , 
		\1488_b1 , \1488_b0 , \1489_b1 , \1489_b0 , \1490_b1 , \1490_b0 , \1491_b1 , \1491_b0 , \1492_b1 , \1492_b0 , 
		\1493_b1 , \1493_b0 , \1494_b1 , \1494_b0 , \1495_b1 , \1495_b0 , \1496_b1 , \1496_b0 , \1497_b1 , \1497_b0 , 
		\1498_b1 , \1498_b0 , \1499_b1 , \1499_b0 , \1500_b1 , \1500_b0 , \1501_b1 , \1501_b0 , \1502_b1 , \1502_b0 , 
		\1503_b1 , \1503_b0 , \1504_b1 , \1504_b0 , \1505_b1 , \1505_b0 , \1506_b1 , \1506_b0 , \1507_b1 , \1507_b0 , 
		\1508_b1 , \1508_b0 , \1509_b1 , \1509_b0 , \1510_b1 , \1510_b0 , \1511_b1 , \1511_b0 , \1512_b1 , \1512_b0 , 
		\1513_b1 , \1513_b0 , \1514_b1 , \1514_b0 , \1515_b1 , \1515_b0 , \1516_b1 , \1516_b0 , \1517_b1 , \1517_b0 , 
		\1518_b1 , \1518_b0 , \1519_b1 , \1519_b0 , \1520_b1 , \1520_b0 , \1521_b1 , \1521_b0 , \1522_b1 , \1522_b0 , 
		\1523_b1 , \1523_b0 , \1524_b1 , \1524_b0 , \1525_b1 , \1525_b0 , \1526_b1 , \1526_b0 , \1527_b1 , \1527_b0 , 
		\1528_b1 , \1528_b0 , \1529_b1 , \1529_b0 , \1530_b1 , \1530_b0 , \1531_b1 , \1531_b0 , \1532_b1 , \1532_b0 , 
		\1533_b1 , \1533_b0 , \1534_b1 , \1534_b0 , \1535_b1 , \1535_b0 , \1536_b1 , \1536_b0 , \1537_b1 , \1537_b0 , 
		\1538_b1 , \1538_b0 , \1539_b1 , \1539_b0 , \1540_b1 , \1540_b0 , \1541_b1 , \1541_b0 , \1542_b1 , \1542_b0 , 
		\1543_b1 , \1543_b0 , \1544_b1 , \1544_b0 , \1545_b1 , \1545_b0 , \1546_b1 , \1546_b0 , \1547_b1 , \1547_b0 , 
		\1548_b1 , \1548_b0 , \1549_b1 , \1549_b0 , \1550_b1 , \1550_b0 , \1551_b1 , \1551_b0 , \1552_b1 , \1552_b0 , 
		\1553_b1 , \1553_b0 , \1554_b1 , \1554_b0 , \1555_b1 , \1555_b0 , \1556_b1 , \1556_b0 , \1557_b1 , \1557_b0 , 
		\1558_b1 , \1558_b0 , \1559_b1 , \1559_b0 , \1560_b1 , \1560_b0 , \1561_b1 , \1561_b0 , \1562_b1 , \1562_b0 , 
		\1563_b1 , \1563_b0 , \1564_b1 , \1564_b0 , \1565_b1 , \1565_b0 , \1566_b1 , \1566_b0 , \1567_b1 , \1567_b0 , 
		\1568_b1 , \1568_b0 , \1569_b1 , \1569_b0 , \1570_b1 , \1570_b0 , \1571_b1 , \1571_b0 , \1572_b1 , \1572_b0 , 
		\1573_b1 , \1573_b0 , \1574_b1 , \1574_b0 , \1575_b1 , \1575_b0 , \1576_b1 , \1576_b0 , \1577_b1 , \1577_b0 , 
		\1578_b1 , \1578_b0 , \1579_b1 , \1579_b0 , \1580_b1 , \1580_b0 , \1581_b1 , \1581_b0 , \1582_b1 , \1582_b0 , 
		\1583_b1 , \1583_b0 , \1584_b1 , \1584_b0 , \1585_b1 , \1585_b0 , \1586_b1 , \1586_b0 , \1587_b1 , \1587_b0 , 
		\1588_b1 , \1588_b0 , \1589_b1 , \1589_b0 , \1590_b1 , \1590_b0 , \1591_b1 , \1591_b0 , \1592_b1 , \1592_b0 , 
		\1593_b1 , \1593_b0 , \1594_b1 , \1594_b0 , \1595_b1 , \1595_b0 , \1596_b1 , \1596_b0 , \1597_b1 , \1597_b0 , 
		\1598_b1 , \1598_b0 , \1599_b1 , \1599_b0 , \1600_b1 , \1600_b0 , \1601_b1 , \1601_b0 , \1602_b1 , \1602_b0 , 
		\1603_b1 , \1603_b0 , \1604_b1 , \1604_b0 , \1605_b1 , \1605_b0 , \1606_b1 , \1606_b0 , \1607_b1 , \1607_b0 , 
		\1608_b1 , \1608_b0 , \1609_b1 , \1609_b0 , \1610_b1 , \1610_b0 , \1611_b1 , \1611_b0 , \1612_b1 , \1612_b0 , 
		\1613_b1 , \1613_b0 , \1614_b1 , \1614_b0 , \1615_b1 , \1615_b0 , \1616_b1 , \1616_b0 , \1617_b1 , \1617_b0 , 
		\1618_b1 , \1618_b0 , \1619_b1 , \1619_b0 , \1620_b1 , \1620_b0 , \1621_b1 , \1621_b0 , \1622_b1 , \1622_b0 , 
		\1623_b1 , \1623_b0 , \1624_b1 , \1624_b0 , \1625_b1 , \1625_b0 , \1626_b1 , \1626_b0 , \1627_b1 , \1627_b0 , 
		\1628_b1 , \1628_b0 , \1629_b1 , \1629_b0 , \1630_b1 , \1630_b0 , \1631_b1 , \1631_b0 , \1632_b1 , \1632_b0 , 
		\1633_b1 , \1633_b0 , \1634_b1 , \1634_b0 , \1635_b1 , \1635_b0 , \1636_b1 , \1636_b0 , \1637_b1 , \1637_b0 , 
		\1638_b1 , \1638_b0 , \1639_b1 , \1639_b0 , \1640_b1 , \1640_b0 , \1641_b1 , \1641_b0 , \1642_b1 , \1642_b0 , 
		\1643_b1 , \1643_b0 , \1644_b1 , \1644_b0 , \1645_b1 , \1645_b0 , \1646_b1 , \1646_b0 , \1647_b1 , \1647_b0 , 
		\1648_b1 , \1648_b0 , \1649_b1 , \1649_b0 , \1650_b1 , \1650_b0 , \1651_b1 , \1651_b0 , \1652_b1 , \1652_b0 , 
		\1653_b1 , \1653_b0 , \1654_b1 , \1654_b0 , \1655_b1 , \1655_b0 , \1656_b1 , \1656_b0 , \1657_b1 , \1657_b0 , 
		\1658_b1 , \1658_b0 , \1659_b1 , \1659_b0 , \1660_b1 , \1660_b0 , \1661_b1 , \1661_b0 , \1662_b1 , \1662_b0 , 
		\1663_b1 , \1663_b0 , \1664_b1 , \1664_b0 , \1665_b1 , \1665_b0 , \1666_b1 , \1666_b0 , \1667_b1 , \1667_b0 , 
		\1668_b1 , \1668_b0 , \1669_b1 , \1669_b0 , \1670_b1 , \1670_b0 , \1671_b1 , \1671_b0 , \1672_b1 , \1672_b0 , 
		\1673_b1 , \1673_b0 , \1674_b1 , \1674_b0 , \1675_b1 , \1675_b0 , \1676_b1 , \1676_b0 , \1677_b1 , \1677_b0 , 
		\1678_b1 , \1678_b0 , \1679_b1 , \1679_b0 , \1680_b1 , \1680_b0 , \1681_b1 , \1681_b0 , \1682_b1 , \1682_b0 , 
		\1683_b1 , \1683_b0 , \1684_b1 , \1684_b0 , \1685_b1 , \1685_b0 , \1686_b1 , \1686_b0 , \1687_b1 , \1687_b0 , 
		\1688_b1 , \1688_b0 , \1689_b1 , \1689_b0 , \1690_b1 , \1690_b0 , \1691_b1 , \1691_b0 , \1692_b1 , \1692_b0 , 
		\1693_b1 , \1693_b0 , \1694_b1 , \1694_b0 , \1695_b1 , \1695_b0 , \1696_b1 , \1696_b0 , \1697_b1 , \1697_b0 , 
		\1698_b1 , \1698_b0 , \1699_b1 , \1699_b0 , \1700_b1 , \1700_b0 , \1701_b1 , \1701_b0 , \1702_b1 , \1702_b0 , 
		\1703_b1 , \1703_b0 , \1704_b1 , \1704_b0 , \1705_b1 , \1705_b0 , \1706_b1 , \1706_b0 , \1707_b1 , \1707_b0 , 
		\1708_b1 , \1708_b0 , \1709_b1 , \1709_b0 , \1710_b1 , \1710_b0 , \1711_b1 , \1711_b0 , \1712_b1 , \1712_b0 , 
		\1713_b1 , \1713_b0 , \1714_b1 , \1714_b0 , \1715_b1 , \1715_b0 , \1716_b1 , \1716_b0 , \1717_b1 , \1717_b0 , 
		\1718_b1 , \1718_b0 , \1719_b1 , \1719_b0 , \1720_b1 , \1720_b0 , \1721_b1 , \1721_b0 , \1722_b1 , \1722_b0 , 
		\1723_b1 , \1723_b0 , \1724_b1 , \1724_b0 , \1725_b1 , \1725_b0 , \1726_b1 , \1726_b0 , \1727_b1 , \1727_b0 , 
		\1728_b1 , \1728_b0 , \1729_b1 , \1729_b0 , \1730_b1 , \1730_b0 , \1731_b1 , \1731_b0 , \1732_b1 , \1732_b0 , 
		\1733_b1 , \1733_b0 , \1734_b1 , \1734_b0 , \1735_b1 , \1735_b0 , \1736_b1 , \1736_b0 , \1737_b1 , \1737_b0 , 
		\1738_b1 , \1738_b0 , \1739_b1 , \1739_b0 , \1740_b1 , \1740_b0 , \1741_b1 , \1741_b0 , \1742_b1 , \1742_b0 , 
		\1743_b1 , \1743_b0 , \1744_b1 , \1744_b0 , \1745_b1 , \1745_b0 , \1746_b1 , \1746_b0 , \1747_b1 , \1747_b0 , 
		\1748_b1 , \1748_b0 , \1749_b1 , \1749_b0 , \1750_b1 , \1750_b0 , \1751_b1 , \1751_b0 , \1752_b1 , \1752_b0 , 
		\1753_b1 , \1753_b0 , \1754_b1 , \1754_b0 , \1755_b1 , \1755_b0 , \1756_b1 , \1756_b0 , \1757_b1 , \1757_b0 , 
		\1758_b1 , \1758_b0 , \1759_b1 , \1759_b0 , \1760_b1 , \1760_b0 , \1761_b1 , \1761_b0 , \1762_b1 , \1762_b0 , 
		\1763_b1 , \1763_b0 , \1764_b1 , \1764_b0 , \1765_b1 , \1765_b0 , \1766_b1 , \1766_b0 , \1767_b1 , \1767_b0 , 
		\1768_b1 , \1768_b0 , \1769_b1 , \1769_b0 , \1770_b1 , \1770_b0 , \1771_b1 , \1771_b0 , \1772_b1 , \1772_b0 , 
		\1773_b1 , \1773_b0 , \1774_b1 , \1774_b0 , \1775_b1 , \1775_b0 , \1776_b1 , \1776_b0 , \1777_b1 , \1777_b0 , 
		\1778_b1 , \1778_b0 , \1779_b1 , \1779_b0 , \1780_b1 , \1780_b0 , \1781_b1 , \1781_b0 , \1782_b1 , \1782_b0 , 
		\1783_b1 , \1783_b0 , \1784_b1 , \1784_b0 , \1785_b1 , \1785_b0 , \1786_b1 , \1786_b0 , \1787_b1 , \1787_b0 , 
		\1788_b1 , \1788_b0 , \1789_b1 , \1789_b0 , \1790_b1 , \1790_b0 , \1791_b1 , \1791_b0 , \1792_b1 , \1792_b0 , 
		\1793_b1 , \1793_b0 , \1794_b1 , \1794_b0 , \1795_b1 , \1795_b0 , \1796_b1 , \1796_b0 , \1797_b1 , \1797_b0 , 
		\1798_b1 , \1798_b0 , \1799_b1 , \1799_b0 , \1800_b1 , \1800_b0 , \1801_b1 , \1801_b0 , \1802_b1 , \1802_b0 , 
		\1803_b1 , \1803_b0 , \1804_b1 , \1804_b0 , \1805_b1 , \1805_b0 , \1806_b1 , \1806_b0 , \1807_b1 , \1807_b0 , 
		\1808_b1 , \1808_b0 , \1809_b1 , \1809_b0 , \1810_b1 , \1810_b0 , \1811_b1 , \1811_b0 , \1812_b1 , \1812_b0 , 
		\1813_b1 , \1813_b0 , \1814_b1 , \1814_b0 , \1815_b1 , \1815_b0 , \1816_b1 , \1816_b0 , \1817_b1 , \1817_b0 , 
		\1818_b1 , \1818_b0 , \1819_b1 , \1819_b0 , \1820_b1 , \1820_b0 , \1821_b1 , \1821_b0 , \1822_b1 , \1822_b0 , 
		\1823_b1 , \1823_b0 , \1824_b1 , \1824_b0 , \1825_b1 , \1825_b0 , \1826_b1 , \1826_b0 , \1827_b1 , \1827_b0 , 
		\1828_b1 , \1828_b0 , \1829_b1 , \1829_b0 , \1830_b1 , \1830_b0 , \1831_b1 , \1831_b0 , \1832_b1 , \1832_b0 , 
		\1833_b1 , \1833_b0 , \1834_b1 , \1834_b0 , \1835_b1 , \1835_b0 , \1836_b1 , \1836_b0 , \1837_b1 , \1837_b0 , 
		\1838_b1 , \1838_b0 , \1839_b1 , \1839_b0 , \1840_b1 , \1840_b0 , \1841_b1 , \1841_b0 , \1842_b1 , \1842_b0 , 
		\1843_b1 , \1843_b0 , \1844_b1 , \1844_b0 , \1845_b1 , \1845_b0 , \1846_b1 , \1846_b0 , \1847_b1 , \1847_b0 , 
		\1848_b1 , \1848_b0 , \1849_b1 , \1849_b0 , \1850_b1 , \1850_b0 , \1851_b1 , \1851_b0 , \1852_b1 , \1852_b0 , 
		\1853_b1 , \1853_b0 , \1854_b1 , \1854_b0 , \1855_b1 , \1855_b0 , \1856_b1 , \1856_b0 , \1857_b1 , \1857_b0 , 
		\1858_b1 , \1858_b0 , \1859_b1 , \1859_b0 , \1860_b1 , \1860_b0 , \1861_b1 , \1861_b0 , \1862_b1 , \1862_b0 , 
		\1863_b1 , \1863_b0 , \1864_b1 , \1864_b0 , \1865_b1 , \1865_b0 , \1866_b1 , \1866_b0 , \1867_b1 , \1867_b0 , 
		\1868_b1 , \1868_b0 , \1869_b1 , \1869_b0 , \1870_b1 , \1870_b0 , \1871_b1 , \1871_b0 , \1872_b1 , \1872_b0 , 
		\1873_b1 , \1873_b0 , \1874_b1 , \1874_b0 , \1875_b1 , \1875_b0 , \1876_b1 , \1876_b0 , \1877_b1 , \1877_b0 , 
		\1878_b1 , \1878_b0 , \1879_b1 , \1879_b0 , \1880_b1 , \1880_b0 , \1881_b1 , \1881_b0 , \1882_b1 , \1882_b0 , 
		\1883_b1 , \1883_b0 , \1884_b1 , \1884_b0 , \1885_b1 , \1885_b0 , \1886_b1 , \1886_b0 , \1887_b1 , \1887_b0 , 
		\1888_b1 , \1888_b0 , \1889_b1 , \1889_b0 , \1890_b1 , \1890_b0 , \1891_b1 , \1891_b0 , \1892_b1 , \1892_b0 , 
		\1893_b1 , \1893_b0 , \1894_b1 , \1894_b0 , \1895_b1 , \1895_b0 , \1896_b1 , \1896_b0 , \1897_b1 , \1897_b0 , 
		\1898_b1 , \1898_b0 , \1899_b1 , \1899_b0 , \1900_b1 , \1900_b0 , \1901_b1 , \1901_b0 , \1902_b1 , \1902_b0 , 
		\1903_b1 , \1903_b0 , \1904_b1 , \1904_b0 , \1905_b1 , \1905_b0 , \1906_b1 , \1906_b0 , \1907_b1 , \1907_b0 , 
		\1908_b1 , \1908_b0 , \1909_b1 , \1909_b0 , \1910_b1 , \1910_b0 , \1911_b1 , \1911_b0 , \1912_b1 , \1912_b0 , 
		\1913_b1 , \1913_b0 , \1914_b1 , \1914_b0 , \1915_b1 , \1915_b0 , \1916_b1 , \1916_b0 , \1917_b1 , \1917_b0 , 
		\1918_b1 , \1918_b0 , \1919_b1 , \1919_b0 , \1920_b1 , \1920_b0 , \1921_b1 , \1921_b0 , \1922_b1 , \1922_b0 , 
		\1923_b1 , \1923_b0 , \1924_b1 , \1924_b0 , \1925_b1 , \1925_b0 , \1926_b1 , \1926_b0 , \1927_b1 , \1927_b0 , 
		\1928_b1 , \1928_b0 , \1929_b1 , \1929_b0 , \1930_b1 , \1930_b0 , \1931_b1 , \1931_b0 , \1932_b1 , \1932_b0 , 
		\1933_b1 , \1933_b0 , \1934_b1 , \1934_b0 , \1935_b1 , \1935_b0 , \1936_b1 , \1936_b0 , \1937_b1 , \1937_b0 , 
		\1938_b1 , \1938_b0 , \1939_b1 , \1939_b0 , \1940_b1 , \1940_b0 , \1941_b1 , \1941_b0 , \1942_b1 , \1942_b0 , 
		\1943_b1 , \1943_b0 , \1944_b1 , \1944_b0 , \1945_b1 , \1945_b0 , \1946_b1 , \1946_b0 , \1947_b1 , \1947_b0 , 
		\1948_b1 , \1948_b0 , \1949_b1 , \1949_b0 , \1950_b1 , \1950_b0 , \1951_b1 , \1951_b0 , \1952_b1 , \1952_b0 , 
		\1953_b1 , \1953_b0 , \1954_b1 , \1954_b0 , \1955_b1 , \1955_b0 , \1956_b1 , \1956_b0 , \1957_b1 , \1957_b0 , 
		\1958_b1 , \1958_b0 , \1959_b1 , \1959_b0 , \1960_b1 , \1960_b0 , \1961_b1 , \1961_b0 , \1962_b1 , \1962_b0 , 
		\1963_b1 , \1963_b0 , \1964_b1 , \1964_b0 , \1965_b1 , \1965_b0 , \1966_b1 , \1966_b0 , \1967_b1 , \1967_b0 , 
		\1968_b1 , \1968_b0 , \1969_b1 , \1969_b0 , \1970_b1 , \1970_b0 , \1971_b1 , \1971_b0 , \1972_b1 , \1972_b0 , 
		\1973_b1 , \1973_b0 , \1974_b1 , \1974_b0 , \1975_b1 , \1975_b0 , \1976_b1 , \1976_b0 , \1977_b1 , \1977_b0 , 
		\1978_b1 , \1978_b0 , \1979_b1 , \1979_b0 , \1980_b1 , \1980_b0 , \1981_b1 , \1981_b0 , \1982_b1 , \1982_b0 , 
		\1983_b1 , \1983_b0 , \1984_b1 , \1984_b0 , \1985_b1 , \1985_b0 , \1986_b1 , \1986_b0 , \1987_b1 , \1987_b0 , 
		\1988_b1 , \1988_b0 , \1989_b1 , \1989_b0 , \1990_b1 , \1990_b0 , \1991_b1 , \1991_b0 , \1992_b1 , \1992_b0 , 
		\1993_b1 , \1993_b0 , \1994_b1 , \1994_b0 , \1995_b1 , \1995_b0 , \1996_b1 , \1996_b0 , \1997_b1 , \1997_b0 , 
		\1998_b1 , \1998_b0 , \1999_b1 , \1999_b0 , \2000_b1 , \2000_b0 , \2001_b1 , \2001_b0 , \2002_b1 , \2002_b0 , 
		\2003_b1 , \2003_b0 , \2004_b1 , \2004_b0 , \2005_b1 , \2005_b0 , \2006_b1 , \2006_b0 , \2007_b1 , \2007_b0 , 
		\2008_b1 , \2008_b0 , \2009_b1 , \2009_b0 , \2010_b1 , \2010_b0 , \2011_b1 , \2011_b0 , \2012_b1 , \2012_b0 , 
		\2013_b1 , \2013_b0 , \2014_b1 , \2014_b0 , \2015_b1 , \2015_b0 , \2016_b1 , \2016_b0 , \2017_b1 , \2017_b0 , 
		\2018_b1 , \2018_b0 , \2019_b1 , \2019_b0 , \2020_b1 , \2020_b0 , \2021_b1 , \2021_b0 , \2022_b1 , \2022_b0 , 
		\2023_b1 , \2023_b0 , \2024_b1 , \2024_b0 , \2025_b1 , \2025_b0 , \2026_b1 , \2026_b0 , \2027_b1 , \2027_b0 , 
		\2028_b1 , \2028_b0 , \2029_b1 , \2029_b0 , \2030_b1 , \2030_b0 , \2031_b1 , \2031_b0 , \2032_b1 , \2032_b0 , 
		\2033_b1 , \2033_b0 , \2034_b1 , \2034_b0 , \2035_b1 , \2035_b0 , \2036_b1 , \2036_b0 , \2037_b1 , \2037_b0 , 
		\2038_b1 , \2038_b0 , \2039_b1 , \2039_b0 , \2040_b1 , \2040_b0 , \2041_b1 , \2041_b0 , \2042_b1 , \2042_b0 , 
		\2043_b1 , \2043_b0 , \2044_b1 , \2044_b0 , \2045_b1 , \2045_b0 , \2046_b1 , \2046_b0 , \2047_b1 , \2047_b0 , 
		\2048_b1 , \2048_b0 , \2049_b1 , \2049_b0 , \2050_b1 , \2050_b0 , \2051_b1 , \2051_b0 , \2052_b1 , \2052_b0 , 
		\2053_b1 , \2053_b0 , \2054_b1 , \2054_b0 , \2055_b1 , \2055_b0 , \2056_b1 , \2056_b0 , \2057_b1 , \2057_b0 , 
		\2058_b1 , \2058_b0 , \2059_b1 , \2059_b0 , \2060_b1 , \2060_b0 , \2061_b1 , \2061_b0 , \2062_b1 , \2062_b0 , 
		\2063_b1 , \2063_b0 , \2064_b1 , \2064_b0 , \2065_b1 , \2065_b0 , \2066_b1 , \2066_b0 , \2067_b1 , \2067_b0 , 
		\2068_b1 , \2068_b0 , \2069_b1 , \2069_b0 , \2070_b1 , \2070_b0 , \2071_b1 , \2071_b0 , \2072_b1 , \2072_b0 , 
		\2073_b1 , \2073_b0 , \2074_b1 , \2074_b0 , \2075_b1 , \2075_b0 , \2076_b1 , \2076_b0 , \2077_b1 , \2077_b0 , 
		\2078_b1 , \2078_b0 , \2079_b1 , \2079_b0 , \2080_b1 , \2080_b0 , \2081_b1 , \2081_b0 , \2082_b1 , \2082_b0 , 
		\2083_b1 , \2083_b0 , \2084_b1 , \2084_b0 , \2085_b1 , \2085_b0 , \2086_b1 , \2086_b0 , \2087_b1 , \2087_b0 , 
		\2088_b1 , \2088_b0 , \2089_b1 , \2089_b0 , \2090_b1 , \2090_b0 , \2091_b1 , \2091_b0 , \2092_b1 , \2092_b0 , 
		\2093_b1 , \2093_b0 , \2094_b1 , \2094_b0 , \2095_b1 , \2095_b0 , \2096_b1 , \2096_b0 , \2097_b1 , \2097_b0 , 
		\2098_b1 , \2098_b0 , \2099_b1 , \2099_b0 , \2100_b1 , \2100_b0 , \2101_b1 , \2101_b0 , \2102_b1 , \2102_b0 , 
		\2103_b1 , \2103_b0 , \2104_b1 , \2104_b0 , \2105_b1 , \2105_b0 , \2106_b1 , \2106_b0 , \2107_b1 , \2107_b0 , 
		\2108_b1 , \2108_b0 , \2109_b1 , \2109_b0 , \2110_b1 , \2110_b0 , \2111_b1 , \2111_b0 , \2112_b1 , \2112_b0 , 
		\2113_b1 , \2113_b0 , \2114_b1 , \2114_b0 , \2115_b1 , \2115_b0 , \2116_b1 , \2116_b0 , \2117_b1 , \2117_b0 , 
		\2118_b1 , \2118_b0 , \2119_b1 , \2119_b0 , \2120_b1 , \2120_b0 , \2121_b1 , \2121_b0 , \2122_b1 , \2122_b0 , 
		\2123_b1 , \2123_b0 , \2124_b1 , \2124_b0 , \2125_b1 , \2125_b0 , \2126_b1 , \2126_b0 , \2127_b1 , \2127_b0 , 
		\2128_b1 , \2128_b0 , \2129_b1 , \2129_b0 , \2130_b1 , \2130_b0 , \2131_b1 , \2131_b0 , \2132_b1 , \2132_b0 , 
		\2133_b1 , \2133_b0 , \2134_b1 , \2134_b0 , \2135_b1 , \2135_b0 , \2136_b1 , \2136_b0 , \2137_b1 , \2137_b0 , 
		\2138_b1 , \2138_b0 , \2139_b1 , \2139_b0 , \2140_b1 , \2140_b0 , \2141_b1 , \2141_b0 , \2142_b1 , \2142_b0 , 
		\2143_b1 , \2143_b0 , \2144_b1 , \2144_b0 , \2145_b1 , \2145_b0 , \2146_b1 , \2146_b0 , \2147_b1 , \2147_b0 , 
		\2148_b1 , \2148_b0 , \2149_b1 , \2149_b0 , \2150_b1 , \2150_b0 , \2151_b1 , \2151_b0 , \2152_b1 , \2152_b0 , 
		\2153_b1 , \2153_b0 , \2154_b1 , \2154_b0 , \2155_b1 , \2155_b0 , \2156_b1 , \2156_b0 , \2157_b1 , \2157_b0 , 
		\2158_b1 , \2158_b0 , \2159_b1 , \2159_b0 , \2160_b1 , \2160_b0 , \2161_b1 , \2161_b0 , \2162_b1 , \2162_b0 , 
		\2163_b1 , \2163_b0 , \2164_b1 , \2164_b0 , \2165_b1 , \2165_b0 , \2166_b1 , \2166_b0 , \2167_b1 , \2167_b0 , 
		\2168_b1 , \2168_b0 , \2169_b1 , \2169_b0 , \2170_b1 , \2170_b0 , \2171_b1 , \2171_b0 , \2172_b1 , \2172_b0 , 
		\2173_b1 , \2173_b0 , \2174_b1 , \2174_b0 , \2175_b1 , \2175_b0 , \2176_b1 , \2176_b0 , \2177_b1 , \2177_b0 , 
		\2178_b1 , \2178_b0 , \2179_b1 , \2179_b0 , \2180_b1 , \2180_b0 , \2181_b1 , \2181_b0 , \2182_b1 , \2182_b0 , 
		\2183_b1 , \2183_b0 , \2184_b1 , \2184_b0 , \2185_b1 , \2185_b0 , \2186_b1 , \2186_b0 , \2187_b1 , \2187_b0 , 
		\2188_b1 , \2188_b0 , \2189_b1 , \2189_b0 , \2190_b1 , \2190_b0 , \2191_b1 , \2191_b0 , \2192_b1 , \2192_b0 , 
		\2193_b1 , \2193_b0 , \2194_b1 , \2194_b0 , \2195_b1 , \2195_b0 , \2196_b1 , \2196_b0 , \2197_b1 , \2197_b0 , 
		\2198_b1 , \2198_b0 , \2199_b1 , \2199_b0 , \2200_b1 , \2200_b0 , \2201_b1 , \2201_b0 , \2202_b1 , \2202_b0 , 
		\2203_b1 , \2203_b0 , \2204_b1 , \2204_b0 , \2205_b1 , \2205_b0 , \2206_b1 , \2206_b0 , \2207_b1 , \2207_b0 , 
		\2208_b1 , \2208_b0 , \2209_b1 , \2209_b0 , \2210_b1 , \2210_b0 , \2211_b1 , \2211_b0 , \2212_b1 , \2212_b0 , 
		\2213_b1 , \2213_b0 , \2214_b1 , \2214_b0 , \2215_b1 , \2215_b0 , \2216_b1 , \2216_b0 , \2217_b1 , \2217_b0 , 
		\2218_b1 , \2218_b0 , \2219_b1 , \2219_b0 , \2220_b1 , \2220_b0 , \2221_b1 , \2221_b0 , \2222_b1 , \2222_b0 , 
		\2223_b1 , \2223_b0 , \2224_b1 , \2224_b0 , \2225_b1 , \2225_b0 , \2226_b1 , \2226_b0 , \2227_b1 , \2227_b0 , 
		\2228_b1 , \2228_b0 , \2229_b1 , \2229_b0 , \2230_b1 , \2230_b0 , \2231_b1 , \2231_b0 , \2232_b1 , \2232_b0 , 
		\2233_b1 , \2233_b0 , \2234_b1 , \2234_b0 , \2235_b1 , \2235_b0 , \2236_b1 , \2236_b0 , \2237_b1 , \2237_b0 , 
		\2238_b1 , \2238_b0 , \2239_b1 , \2239_b0 , \2240_b1 , \2240_b0 , \2241_b1 , \2241_b0 , \2242_b1 , \2242_b0 , 
		\2243_b1 , \2243_b0 , \2244_b1 , \2244_b0 , \2245_b1 , \2245_b0 , \2246_b1 , \2246_b0 , \2247_b1 , \2247_b0 , 
		\2248_b1 , \2248_b0 , \2249_b1 , \2249_b0 , \2250_b1 , \2250_b0 , \2251_b1 , \2251_b0 , \2252_b1 , \2252_b0 , 
		\2253_b1 , \2253_b0 , \2254_b1 , \2254_b0 , \2255_b1 , \2255_b0 , \2256_b1 , \2256_b0 , \2257_b1 , \2257_b0 , 
		\2258_b1 , \2258_b0 , \2259_b1 , \2259_b0 , \2260_b1 , \2260_b0 , \2261_b1 , \2261_b0 , \2262_b1 , \2262_b0 , 
		\2263_b1 , \2263_b0 , \2264_b1 , \2264_b0 , \2265_b1 , \2265_b0 , \2266_b1 , \2266_b0 , \2267_b1 , \2267_b0 , 
		\2268_b1 , \2268_b0 , \2269_b1 , \2269_b0 , \2270_b1 , \2270_b0 , \2271_b1 , \2271_b0 , \2272_b1 , \2272_b0 , 
		\2273_b1 , \2273_b0 , \2274_b1 , \2274_b0 , \2275_b1 , \2275_b0 , \2276_b1 , \2276_b0 , \2277_b1 , \2277_b0 , 
		\2278_b1 , \2278_b0 , \2279_b1 , \2279_b0 , \2280_b1 , \2280_b0 , \2281_b1 , \2281_b0 , \2282_b1 , \2282_b0 , 
		\2283_b1 , \2283_b0 , \2284_b1 , \2284_b0 , \2285_b1 , \2285_b0 , \2286_b1 , \2286_b0 , \2287_b1 , \2287_b0 , 
		\2288_b1 , \2288_b0 , \2289_b1 , \2289_b0 , \2290_b1 , \2290_b0 , \2291_b1 , \2291_b0 , \2292_b1 , \2292_b0 , 
		\2293_b1 , \2293_b0 , \2294_b1 , \2294_b0 , \2295_b1 , \2295_b0 , \2296_b1 , \2296_b0 , \2297_b1 , \2297_b0 , 
		\2298_b1 , \2298_b0 , \2299_b1 , \2299_b0 , \2300_b1 , \2300_b0 , \2301_b1 , \2301_b0 , \2302_b1 , \2302_b0 , 
		\2303_b1 , \2303_b0 , \2304_b1 , \2304_b0 , \2305_b1 , \2305_b0 , \2306_b1 , \2306_b0 , \2307_b1 , \2307_b0 , 
		\2308_b1 , \2308_b0 , \2309_b1 , \2309_b0 , \2310_b1 , \2310_b0 , \2311_b1 , \2311_b0 , \2312_b1 , \2312_b0 , 
		\2313_b1 , \2313_b0 , \2314_b1 , \2314_b0 , \2315_b1 , \2315_b0 , \2316_b1 , \2316_b0 , \2317_b1 , \2317_b0 , 
		\2318_b1 , \2318_b0 , \2319_b1 , \2319_b0 , \2320_b1 , \2320_b0 , \2321_b1 , \2321_b0 , \2322_b1 , \2322_b0 , 
		\2323_b1 , \2323_b0 , \2324_b1 , \2324_b0 , \2325_b1 , \2325_b0 , \2326_b1 , \2326_b0 , \2327_b1 , \2327_b0 , 
		\2328_b1 , \2328_b0 , \2329_b1 , \2329_b0 , \2330_b1 , \2330_b0 , \2331_b1 , \2331_b0 , \2332_b1 , \2332_b0 , 
		\2333_b1 , \2333_b0 , \2334_b1 , \2334_b0 , \2335_b1 , \2335_b0 , \2336_b1 , \2336_b0 , \2337_b1 , \2337_b0 , 
		\2338_b1 , \2338_b0 , \2339_b1 , \2339_b0 , \2340_b1 , \2340_b0 , \2341_b1 , \2341_b0 , \2342_b1 , \2342_b0 , 
		\2343_b1 , \2343_b0 , \2344_b1 , \2344_b0 , \2345_b1 , \2345_b0 , \2346_b1 , \2346_b0 , \2347_b1 , \2347_b0 , 
		\2348_b1 , \2348_b0 , \2349_b1 , \2349_b0 , \2350_b1 , \2350_b0 , \2351_b1 , \2351_b0 , \2352_b1 , \2352_b0 , 
		\2353_b1 , \2353_b0 , \2354_b1 , \2354_b0 , \2355_b1 , \2355_b0 , \2356_b1 , \2356_b0 , \2357_b1 , \2357_b0 , 
		\2358_b1 , \2358_b0 , \2359_b1 , \2359_b0 , \2360_b1 , \2360_b0 , \2361_b1 , \2361_b0 , \2362_b1 , \2362_b0 , 
		\2363_b1 , \2363_b0 , \2364_b1 , \2364_b0 , \2365_b1 , \2365_b0 , \2366_b1 , \2366_b0 , \2367_b1 , \2367_b0 , 
		\2368_b1 , \2368_b0 , \2369_b1 , \2369_b0 , \2370_b1 , \2370_b0 , \2371_b1 , \2371_b0 , \2372_b1 , \2372_b0 , 
		\2373_b1 , \2373_b0 , \2374_b1 , \2374_b0 , \2375_b1 , \2375_b0 , \2376_b1 , \2376_b0 , \2377_b1 , \2377_b0 , 
		\2378_b1 , \2378_b0 , \2379_b1 , \2379_b0 , \2380_b1 , \2380_b0 , \2381_b1 , \2381_b0 , \2382_b1 , \2382_b0 , 
		\2383_b1 , \2383_b0 , \2384_b1 , \2384_b0 , \2385_b1 , \2385_b0 , \2386_b1 , \2386_b0 , \2387_b1 , \2387_b0 , 
		\2388_b1 , \2388_b0 , \2389_b1 , \2389_b0 , \2390_b1 , \2390_b0 , \2391_b1 , \2391_b0 , \2392_b1 , \2392_b0 , 
		\2393_b1 , \2393_b0 , \2394_b1 , \2394_b0 , \2395_b1 , \2395_b0 , \2396_b1 , \2396_b0 , \2397_b1 , \2397_b0 , 
		\2398_b1 , \2398_b0 , \2399_b1 , \2399_b0 , \2400_b1 , \2400_b0 , \2401_b1 , \2401_b0 , \2402_b1 , \2402_b0 , 
		\2403_b1 , \2403_b0 , \2404_b1 , \2404_b0 , \2405_b1 , \2405_b0 , \2406_b1 , \2406_b0 , \2407_b1 , \2407_b0 , 
		\2408_b1 , \2408_b0 , \2409_b1 , \2409_b0 , \2410_b1 , \2410_b0 , \2411_b1 , \2411_b0 , \2412_b1 , \2412_b0 , 
		\2413_b1 , \2413_b0 , \2414_b1 , \2414_b0 , \2415_b1 , \2415_b0 , \2416_b1 , \2416_b0 , \2417_b1 , \2417_b0 , 
		\2418_b1 , \2418_b0 , \2419_b1 , \2419_b0 , \2420_b1 , \2420_b0 , \2421_b1 , \2421_b0 , \2422_b1 , \2422_b0 , 
		\2423_b1 , \2423_b0 , \2424_b1 , \2424_b0 , \2425_b1 , \2425_b0 , \2426_b1 , \2426_b0 , \2427_b1 , \2427_b0 , 
		\2428_b1 , \2428_b0 , \2429_b1 , \2429_b0 , \2430_b1 , \2430_b0 , \2431_b1 , \2431_b0 , \2432_b1 , \2432_b0 , 
		\2433_b1 , \2433_b0 , \2434_b1 , \2434_b0 , \2435_b1 , \2435_b0 , \2436_b1 , \2436_b0 , \2437_b1 , \2437_b0 , 
		\2438_b1 , \2438_b0 , \2439_b1 , \2439_b0 , \2440_b1 , \2440_b0 , \2441_b1 , \2441_b0 , \2442_b1 , \2442_b0 , 
		\2443_b1 , \2443_b0 , \2444_b1 , \2444_b0 , \2445_b1 , \2445_b0 , \2446_b1 , \2446_b0 , \2447_b1 , \2447_b0 , 
		\2448_b1 , \2448_b0 , \2449_b1 , \2449_b0 , \2450_b1 , \2450_b0 , \2451_b1 , \2451_b0 , \2452_b1 , \2452_b0 , 
		\2453_b1 , \2453_b0 , \2454_b1 , \2454_b0 , \2455_b1 , \2455_b0 , \2456_b1 , \2456_b0 , \2457_b1 , \2457_b0 , 
		\2458_b1 , \2458_b0 , \2459_b1 , \2459_b0 , \2460_b1 , \2460_b0 , \2461_b1 , \2461_b0 , \2462_b1 , \2462_b0 , 
		\2463_b1 , \2463_b0 , \2464_b1 , \2464_b0 , \2465_b1 , \2465_b0 , \2466_b1 , \2466_b0 , \2467_b1 , \2467_b0 , 
		\2468_b1 , \2468_b0 , \2469_b1 , \2469_b0 , \2470_b1 , \2470_b0 , \2471_b1 , \2471_b0 , \2472_b1 , \2472_b0 , 
		\2473_b1 , \2473_b0 , \2474_b1 , \2474_b0 , \2475_b1 , \2475_b0 , \2476_b1 , \2476_b0 , \2477_b1 , \2477_b0 , 
		\2478_b1 , \2478_b0 , \2479_b1 , \2479_b0 , \2480_b1 , \2480_b0 , \2481_b1 , \2481_b0 , \2482_b1 , \2482_b0 , 
		\2483_b1 , \2483_b0 , \2484_b1 , \2484_b0 , \2485_b1 , \2485_b0 , \2486_b1 , \2486_b0 , \2487_b1 , \2487_b0 , 
		\2488_b1 , \2488_b0 , \2489_b1 , \2489_b0 , \2490_b1 , \2490_b0 , \2491_b1 , \2491_b0 , \2492_b1 , \2492_b0 , 
		\2493_b1 , \2493_b0 , \2494_b1 , \2494_b0 , \2495_b1 , \2495_b0 , \2496_b1 , \2496_b0 , \2497_b1 , \2497_b0 , 
		\2498_b1 , \2498_b0 , \2499_b1 , \2499_b0 , \2500_b1 , \2500_b0 , \2501_b1 , \2501_b0 , \2502_b1 , \2502_b0 , 
		\2503_b1 , \2503_b0 , \2504_b1 , \2504_b0 , \2505_b1 , \2505_b0 , \2506_b1 , \2506_b0 , \2507_b1 , \2507_b0 , 
		\2508_b1 , \2508_b0 , \2509_b1 , \2509_b0 , \2510_b1 , \2510_b0 , \2511_b1 , \2511_b0 , \2512_b1 , \2512_b0 , 
		\2513_b1 , \2513_b0 , \2514_b1 , \2514_b0 , \2515_b1 , \2515_b0 , \2516_b1 , \2516_b0 , \2517_b1 , \2517_b0 , 
		\2518_b1 , \2518_b0 , \2519_b1 , \2519_b0 , \2520_b1 , \2520_b0 , \2521_b1 , \2521_b0 , \2522_b1 , \2522_b0 , 
		\2523_b1 , \2523_b0 , \2524_b1 , \2524_b0 , \2525_b1 , \2525_b0 , \2526_b1 , \2526_b0 , \2527_b1 , \2527_b0 , 
		\2528_b1 , \2528_b0 , \2529_b1 , \2529_b0 , \2530_b1 , \2530_b0 , \2531_b1 , \2531_b0 , \2532_b1 , \2532_b0 , 
		\2533_b1 , \2533_b0 , \2534_b1 , \2534_b0 , \2535_b1 , \2535_b0 , \2536_b1 , \2536_b0 , \2537_b1 , \2537_b0 , 
		\2538_b1 , \2538_b0 , \2539_b1 , \2539_b0 , \2540_b1 , \2540_b0 , \2541_b1 , \2541_b0 , \2542_b1 , \2542_b0 , 
		\2543_b1 , \2543_b0 , \2544_b1 , \2544_b0 , \2545_b1 , \2545_b0 , \2546_b1 , \2546_b0 , \2547_b1 , \2547_b0 , 
		\2548_b1 , \2548_b0 , \2549_b1 , \2549_b0 , \2550_b1 , \2550_b0 , \2551_b1 , \2551_b0 , \2552_b1 , \2552_b0 , 
		\2553_b1 , \2553_b0 , \2554_b1 , \2554_b0 , \2555_b1 , \2555_b0 , \2556_b1 , \2556_b0 , \2557_b1 , \2557_b0 , 
		\2558_b1 , \2558_b0 , \2559_b1 , \2559_b0 , \2560_b1 , \2560_b0 , \2561_b1 , \2561_b0 , \2562_b1 , \2562_b0 , 
		\2563_b1 , \2563_b0 , \2564_b1 , \2564_b0 , \2565_b1 , \2565_b0 , \2566_b1 , \2566_b0 , \2567_b1 , \2567_b0 , 
		\2568_b1 , \2568_b0 , \2569_b1 , \2569_b0 , \2570_b1 , \2570_b0 , \2571_b1 , \2571_b0 , \2572_b1 , \2572_b0 , 
		\2573_b1 , \2573_b0 , \2574_b1 , \2574_b0 , \2575_b1 , \2575_b0 , \2576_b1 , \2576_b0 , \2577_b1 , \2577_b0 , 
		\2578_b1 , \2578_b0 , \2579_b1 , \2579_b0 , \2580_b1 , \2580_b0 , \2581_b1 , \2581_b0 , \2582_b1 , \2582_b0 , 
		\2583_b1 , \2583_b0 , \2584_b1 , \2584_b0 , \2585_b1 , \2585_b0 , \2586_b1 , \2586_b0 , \2587_b1 , \2587_b0 , 
		\2588_b1 , \2588_b0 , \2589_b1 , \2589_b0 , \2590_b1 , \2590_b0 , \2591_b1 , \2591_b0 , \2592_b1 , \2592_b0 , 
		\2593_b1 , \2593_b0 , \2594_b1 , \2594_b0 , \2595_b1 , \2595_b0 , \2596_b1 , \2596_b0 , \2597_b1 , \2597_b0 , 
		\2598_b1 , \2598_b0 , \2599_b1 , \2599_b0 , \2600_b1 , \2600_b0 , \2601_b1 , \2601_b0 , \2602_b1 , \2602_b0 , 
		\2603_b1 , \2603_b0 , \2604_b1 , \2604_b0 , \2605_b1 , \2605_b0 , \2606_b1 , \2606_b0 , \2607_b1 , \2607_b0 , 
		\2608_b1 , \2608_b0 , \2609_b1 , \2609_b0 , \2610_b1 , \2610_b0 , \2611_b1 , \2611_b0 , \2612_b1 , \2612_b0 , 
		\2613_b1 , \2613_b0 , \2614_b1 , \2614_b0 , \2615_b1 , \2615_b0 , \2616_b1 , \2616_b0 , \2617_b1 , \2617_b0 , 
		\2618_b1 , \2618_b0 , \2619_b1 , \2619_b0 , \2620_b1 , \2620_b0 , \2621_b1 , \2621_b0 , \2622_b1 , \2622_b0 , 
		\2623_b1 , \2623_b0 , \2624_b1 , \2624_b0 , \2625_b1 , \2625_b0 , \2626_b1 , \2626_b0 , \2627_b1 , \2627_b0 , 
		\2628_b1 , \2628_b0 , \2629_b1 , \2629_b0 , \2630_b1 , \2630_b0 , \2631_b1 , \2631_b0 , \2632_b1 , \2632_b0 , 
		\2633_b1 , \2633_b0 , \2634_b1 , \2634_b0 , \2635_b1 , \2635_b0 , \2636_b1 , \2636_b0 , \2637_b1 , \2637_b0 , 
		\2638_b1 , \2638_b0 , \2639_b1 , \2639_b0 , \2640_b1 , \2640_b0 , \2641_b1 , \2641_b0 , \2642_b1 , \2642_b0 , 
		\2643_b1 , \2643_b0 , \2644_b1 , \2644_b0 , \2645_b1 , \2645_b0 , \2646_b1 , \2646_b0 , \2647_b1 , \2647_b0 , 
		\2648_b1 , \2648_b0 , \2649_b1 , \2649_b0 , \2650_b1 , \2650_b0 , \2651_b1 , \2651_b0 , \2652_b1 , \2652_b0 , 
		\2653_b1 , \2653_b0 , \2654_b1 , \2654_b0 , \2655_b1 , \2655_b0 , \2656_b1 , \2656_b0 , \2657_b1 , \2657_b0 , 
		\2658_b1 , \2658_b0 , \2659_b1 , \2659_b0 , \2660_b1 , \2660_b0 , \2661_b1 , \2661_b0 , \2662_b1 , \2662_b0 , 
		\2663_b1 , \2663_b0 , \2664_b1 , \2664_b0 , \2665_b1 , \2665_b0 , \2666_b1 , \2666_b0 , \2667_b1 , \2667_b0 , 
		\2668_b1 , \2668_b0 , \2669_b1 , \2669_b0 , \2670_b1 , \2670_b0 , \2671_b1 , \2671_b0 , \2672_b1 , \2672_b0 , 
		\2673_b1 , \2673_b0 , \2674_b1 , \2674_b0 , \2675_b1 , \2675_b0 , \2676_b1 , \2676_b0 , \2677_b1 , \2677_b0 , 
		\2678_b1 , \2678_b0 , \2679_b1 , \2679_b0 , \2680_b1 , \2680_b0 , \2681_b1 , \2681_b0 , \2682_b1 , \2682_b0 , 
		\2683_b1 , \2683_b0 , \2684_b1 , \2684_b0 , \2685_b1 , \2685_b0 , \2686_b1 , \2686_b0 , \2687_b1 , \2687_b0 , 
		\2688_b1 , \2688_b0 , \2689_b1 , \2689_b0 , \2690_b1 , \2690_b0 , \2691_b1 , \2691_b0 , \2692_b1 , \2692_b0 , 
		\2693_b1 , \2693_b0 , \2694_b1 , \2694_b0 , \2695_b1 , \2695_b0 , \2696_b1 , \2696_b0 , \2697_b1 , \2697_b0 , 
		\2698_b1 , \2698_b0 , \2699_b1 , \2699_b0 , \2700_b1 , \2700_b0 , \2701_b1 , \2701_b0 , \2702_b1 , \2702_b0 , 
		\2703_b1 , \2703_b0 , \2704_b1 , \2704_b0 , \2705_b1 , \2705_b0 , \2706_b1 , \2706_b0 , \2707_b1 , \2707_b0 , 
		\2708_b1 , \2708_b0 , \2709_b1 , \2709_b0 , \2710_b1 , \2710_b0 , \2711_b1 , \2711_b0 , \2712_b1 , \2712_b0 , 
		\2713_b1 , \2713_b0 , \2714_b1 , \2714_b0 , \2715_b1 , \2715_b0 , \2716_b1 , \2716_b0 , \2717_b1 , \2717_b0 , 
		\2718_b1 , \2718_b0 , \2719_b1 , \2719_b0 , \2720_b1 , \2720_b0 , \2721_b1 , \2721_b0 , \2722_b1 , \2722_b0 , 
		\2723_b1 , \2723_b0 , \2724_b1 , \2724_b0 , \2725_b1 , \2725_b0 , \2726_b1 , \2726_b0 , \2727_b1 , \2727_b0 , 
		\2728_b1 , \2728_b0 , \2729_b1 , \2729_b0 , \2730_b1 , \2730_b0 , \2731_b1 , \2731_b0 , \2732_b1 , \2732_b0 , 
		\2733_b1 , \2733_b0 , \2734_b1 , \2734_b0 , \2735_b1 , \2735_b0 , \2736_b1 , \2736_b0 , \2737_b1 , \2737_b0 , 
		\2738_b1 , \2738_b0 , \2739_b1 , \2739_b0 , \2740_b1 , \2740_b0 , \2741_b1 , \2741_b0 , \2742_b1 , \2742_b0 , 
		\2743_b1 , \2743_b0 , \2744_b1 , \2744_b0 , \2745_b1 , \2745_b0 , \2746_b1 , \2746_b0 , \2747_b1 , \2747_b0 , 
		\2748_b1 , \2748_b0 , \2749_b1 , \2749_b0 , \2750_b1 , \2750_b0 , \2751_b1 , \2751_b0 , \2752_b1 , \2752_b0 , 
		\2753_b1 , \2753_b0 , \2754_b1 , \2754_b0 , \2755_b1 , \2755_b0 , \2756_b1 , \2756_b0 , \2757_b1 , \2757_b0 , 
		\2758_b1 , \2758_b0 , \2759_b1 , \2759_b0 , \2760_b1 , \2760_b0 , \2761_b1 , \2761_b0 , \2762_b1 , \2762_b0 , 
		\2763_b1 , \2763_b0 , \2764_b1 , \2764_b0 , \2765_b1 , \2765_b0 , \2766_b1 , \2766_b0 , \2767_b1 , \2767_b0 , 
		\2768_b1 , \2768_b0 , \2769_b1 , \2769_b0 , \2770_b1 , \2770_b0 , \2771_b1 , \2771_b0 , \2772_b1 , \2772_b0 , 
		\2773_b1 , \2773_b0 , \2774_b1 , \2774_b0 , \2775_b1 , \2775_b0 , \2776_b1 , \2776_b0 , \2777_b1 , \2777_b0 , 
		\2778_b1 , \2778_b0 , \2779_b1 , \2779_b0 , \2780_b1 , \2780_b0 , \2781_b1 , \2781_b0 , \2782_b1 , \2782_b0 , 
		\2783_b1 , \2783_b0 , \2784_b1 , \2784_b0 , \2785_b1 , \2785_b0 , \2786_b1 , \2786_b0 , \2787_b1 , \2787_b0 , 
		\2788_b1 , \2788_b0 , \2789_b1 , \2789_b0 , \2790_b1 , \2790_b0 , \2791_b1 , \2791_b0 , \2792_b1 , \2792_b0 , 
		\2793_b1 , \2793_b0 , \2794_b1 , \2794_b0 , \2795_b1 , \2795_b0 , \2796_b1 , \2796_b0 , \2797_b1 , \2797_b0 , 
		\2798_b1 , \2798_b0 , \2799_b1 , \2799_b0 , \2800_b1 , \2800_b0 , \2801_b1 , \2801_b0 , \2802_b1 , \2802_b0 , 
		\2803_b1 , \2803_b0 , \2804_b1 , \2804_b0 , \2805_b1 , \2805_b0 , \2806_b1 , \2806_b0 , \2807_b1 , \2807_b0 , 
		\2808_b1 , \2808_b0 , \2809_b1 , \2809_b0 , \2810_b1 , \2810_b0 , \2811_b1 , \2811_b0 , \2812_b1 , \2812_b0 , 
		\2813_b1 , \2813_b0 , \2814_b1 , \2814_b0 , \2815_b1 , \2815_b0 , \2816_b1 , \2816_b0 , \2817_b1 , \2817_b0 , 
		\2818_b1 , \2818_b0 , \2819_b1 , \2819_b0 , \2820_b1 , \2820_b0 , \2821_b1 , \2821_b0 , \2822_b1 , \2822_b0 , 
		\2823_b1 , \2823_b0 , \2824_b1 , \2824_b0 , \2825_b1 , \2825_b0 , \2826_b1 , \2826_b0 , \2827_b1 , \2827_b0 , 
		\2828_b1 , \2828_b0 , \2829_b1 , \2829_b0 , \2830_b1 , \2830_b0 , \2831_b1 , \2831_b0 , \2832_b1 , \2832_b0 , 
		\2833_b1 , \2833_b0 , \2834_b1 , \2834_b0 , \2835_b1 , \2835_b0 , \2836_b1 , \2836_b0 , \2837_b1 , \2837_b0 , 
		\2838_b1 , \2838_b0 , \2839_b1 , \2839_b0 , \2840_b1 , \2840_b0 , \2841_b1 , \2841_b0 , \2842_b1 , \2842_b0 , 
		\2843_b1 , \2843_b0 , \2844_b1 , \2844_b0 , \2845_b1 , \2845_b0 , \2846_b1 , \2846_b0 , \2847_b1 , \2847_b0 , 
		\2848_b1 , \2848_b0 , \2849_b1 , \2849_b0 , \2850_b1 , \2850_b0 , \2851_b1 , \2851_b0 , \2852_b1 , \2852_b0 , 
		\2853_b1 , \2853_b0 , \2854_b1 , \2854_b0 , \2855_b1 , \2855_b0 , \2856_b1 , \2856_b0 , \2857_b1 , \2857_b0 , 
		\2858_b1 , \2858_b0 , \2859_b1 , \2859_b0 , \2860_b1 , \2860_b0 , \2861_b1 , \2861_b0 , \2862_b1 , \2862_b0 , 
		\2863_b1 , \2863_b0 , \2864_b1 , \2864_b0 , \2865_b1 , \2865_b0 , \2866_b1 , \2866_b0 , \2867_b1 , \2867_b0 , 
		\2868_b1 , \2868_b0 , \2869_b1 , \2869_b0 , \2870_b1 , \2870_b0 , \2871_b1 , \2871_b0 , \2872_b1 , \2872_b0 , 
		\2873_b1 , \2873_b0 , \2874_b1 , \2874_b0 , \2875_b1 , \2875_b0 , \2876_b1 , \2876_b0 , \2877_b1 , \2877_b0 , 
		\2878_b1 , \2878_b0 , \2879_b1 , \2879_b0 , \2880_b1 , \2880_b0 , \2881_b1 , \2881_b0 , \2882_b1 , \2882_b0 , 
		\2883_b1 , \2883_b0 , \2884_b1 , \2884_b0 , \2885_b1 , \2885_b0 , \2886_b1 , \2886_b0 , \2887_b1 , \2887_b0 , 
		\2888_b1 , \2888_b0 , \2889_b1 , \2889_b0 , \2890_b1 , \2890_b0 , \2891_b1 , \2891_b0 , \2892_b1 , \2892_b0 , 
		\2893_b1 , \2893_b0 , \2894_b1 , \2894_b0 , \2895_b1 , \2895_b0 , \2896_b1 , \2896_b0 , \2897_b1 , \2897_b0 , 
		\2898_b1 , \2898_b0 , \2899_b1 , \2899_b0 , \2900_b1 , \2900_b0 , \2901_b1 , \2901_b0 , \2902_b1 , \2902_b0 , 
		\2903_b1 , \2903_b0 , \2904_b1 , \2904_b0 , \2905_b1 , \2905_b0 , \2906_b1 , \2906_b0 , \2907_b1 , \2907_b0 , 
		\2908_b1 , \2908_b0 , \2909_b1 , \2909_b0 , \2910_b1 , \2910_b0 , \2911_b1 , \2911_b0 , \2912_b1 , \2912_b0 , 
		\2913_b1 , \2913_b0 , \2914_b1 , \2914_b0 , \2915_b1 , \2915_b0 , \2916_b1 , \2916_b0 , \2917_b1 , \2917_b0 , 
		\2918_b1 , \2918_b0 , \2919_b1 , \2919_b0 , \2920_b1 , \2920_b0 , \2921_b1 , \2921_b0 , \2922_b1 , \2922_b0 , 
		\2923_b1 , \2923_b0 , \2924_b1 , \2924_b0 , \2925_b1 , \2925_b0 , \2926_b1 , \2926_b0 , \2927_b1 , \2927_b0 , 
		\2928_b1 , \2928_b0 , \2929_b1 , \2929_b0 , \2930_b1 , \2930_b0 , \2931_b1 , \2931_b0 , \2932_b1 , \2932_b0 , 
		\2933_b1 , \2933_b0 , \2934_b1 , \2934_b0 , \2935_b1 , \2935_b0 , \2936_b1 , \2936_b0 , \2937_b1 , \2937_b0 , 
		\2938_b1 , \2938_b0 , \2939_b1 , \2939_b0 , \2940_b1 , \2940_b0 , \2941_b1 , \2941_b0 , \2942_b1 , \2942_b0 , 
		\2943_b1 , \2943_b0 , \2944_b1 , \2944_b0 , \2945_b1 , \2945_b0 , \2946_b1 , \2946_b0 , \2947_b1 , \2947_b0 , 
		\2948_b1 , \2948_b0 , \2949_b1 , \2949_b0 , \2950_b1 , \2950_b0 , \2951_b1 , \2951_b0 , \2952_b1 , \2952_b0 , 
		\2953_b1 , \2953_b0 , \2954_b1 , \2954_b0 , \2955_b1 , \2955_b0 , \2956_b1 , \2956_b0 , \2957_b1 , \2957_b0 , 
		\2958_b1 , \2958_b0 , \2959_b1 , \2959_b0 , \2960_b1 , \2960_b0 , \2961_b1 , \2961_b0 , \2962_b1 , \2962_b0 , 
		\2963_b1 , \2963_b0 , \2964_b1 , \2964_b0 , \2965_b1 , \2965_b0 , \2966_b1 , \2966_b0 , \2967_b1 , \2967_b0 , 
		\2968_b1 , \2968_b0 , \2969_b1 , \2969_b0 , \2970_b1 , \2970_b0 , \2971_b1 , \2971_b0 , \2972_b1 , \2972_b0 , 
		\2973_b1 , \2973_b0 , \2974_b1 , \2974_b0 , \2975_b1 , \2975_b0 , \2976_b1 , \2976_b0 , \2977_b1 , \2977_b0 , 
		\2978_b1 , \2978_b0 , \2979_b1 , \2979_b0 , \2980_b1 , \2980_b0 , \2981_b1 , \2981_b0 , \2982_b1 , \2982_b0 , 
		\2983_b1 , \2983_b0 , \2984_b1 , \2984_b0 , \2985_b1 , \2985_b0 , \2986_b1 , \2986_b0 , \2987_b1 , \2987_b0 , 
		\2988_b1 , \2988_b0 , \2989_b1 , \2989_b0 , \2990_b1 , \2990_b0 , \2991_b1 , \2991_b0 , \2992_b1 , \2992_b0 , 
		\2993_b1 , \2993_b0 , \2994_b1 , \2994_b0 , \2995_b1 , \2995_b0 , \2996_b1 , \2996_b0 , \2997_b1 , \2997_b0 , 
		\2998_b1 , \2998_b0 , \2999_b1 , \2999_b0 , \3000_b1 , \3000_b0 , \3001_b1 , \3001_b0 , \3002_b1 , \3002_b0 , 
		\3003_b1 , \3003_b0 , \3004_b1 , \3004_b0 , \3005_b1 , \3005_b0 , \3006_b1 , \3006_b0 , \3007_b1 , \3007_b0 , 
		\3008_b1 , \3008_b0 , \3009_b1 , \3009_b0 , \3010_b1 , \3010_b0 , \3011_b1 , \3011_b0 , \3012_b1 , \3012_b0 , 
		\3013_b1 , \3013_b0 , \3014_b1 , \3014_b0 , \3015_b1 , \3015_b0 , \3016_b1 , \3016_b0 , \3017_b1 , \3017_b0 , 
		\3018_b1 , \3018_b0 , \3019_b1 , \3019_b0 , \3020_b1 , \3020_b0 , \3021_b1 , \3021_b0 , \3022_b1 , \3022_b0 , 
		\3023_b1 , \3023_b0 , \3024_b1 , \3024_b0 , \3025_b1 , \3025_b0 , \3026_b1 , \3026_b0 , \3027_b1 , \3027_b0 , 
		\3028_b1 , \3028_b0 , \3029_b1 , \3029_b0 , \3030_b1 , \3030_b0 , \3031_b1 , \3031_b0 , \3032_b1 , \3032_b0 , 
		\3033_b1 , \3033_b0 , \3034_b1 , \3034_b0 , \3035_b1 , \3035_b0 , \3036_b1 , \3036_b0 , \3037_b1 , \3037_b0 , 
		\3038_b1 , \3038_b0 , \3039_b1 , \3039_b0 , \3040_b1 , \3040_b0 , \3041_b1 , \3041_b0 , \3042_b1 , \3042_b0 , 
		\3043_b1 , \3043_b0 , \3044_b1 , \3044_b0 , \3045_b1 , \3045_b0 , \3046_b1 , \3046_b0 , \3047_b1 , \3047_b0 , 
		\3048_b1 , \3048_b0 , \3049_b1 , \3049_b0 , \3050_b1 , \3050_b0 , \3051_b1 , \3051_b0 , \3052_b1 , \3052_b0 , 
		\3053_b1 , \3053_b0 , \3054_b1 , \3054_b0 , \3055_b1 , \3055_b0 , \3056_b1 , \3056_b0 , \3057_b1 , \3057_b0 , 
		\3058_b1 , \3058_b0 , \3059_b1 , \3059_b0 , \3060_b1 , \3060_b0 , \3061_b1 , \3061_b0 , \3062_b1 , \3062_b0 , 
		\3063_b1 , \3063_b0 , \3064_b1 , \3064_b0 , \3065_b1 , \3065_b0 , \3066_b1 , \3066_b0 , \3067_b1 , \3067_b0 , 
		\3068_b1 , \3068_b0 , \3069_b1 , \3069_b0 , \3070_b1 , \3070_b0 , \3071_b1 , \3071_b0 , \3072_b1 , \3072_b0 , 
		\3073_b1 , \3073_b0 , \3074_b1 , \3074_b0 , \3075_b1 , \3075_b0 , \3076_b1 , \3076_b0 , \3077_b1 , \3077_b0 , 
		\3078_b1 , \3078_b0 , \3079_b1 , \3079_b0 , \3080_b1 , \3080_b0 , \3081_b1 , \3081_b0 , \3082_b1 , \3082_b0 , 
		\3083_b1 , \3083_b0 , \3084_b1 , \3084_b0 , \3085_b1 , \3085_b0 , \3086_b1 , \3086_b0 , \3087_b1 , \3087_b0 , 
		\3088_b1 , \3088_b0 , \3089_b1 , \3089_b0 , \3090_b1 , \3090_b0 , \3091_b1 , \3091_b0 , \3092_b1 , \3092_b0 , 
		\3093_b1 , \3093_b0 , \3094_b1 , \3094_b0 , \3095_b1 , \3095_b0 , \3096_b1 , \3096_b0 , \3097_b1 , \3097_b0 , 
		\3098_b1 , \3098_b0 , \3099_b1 , \3099_b0 , \3100_b1 , \3100_b0 , \3101_b1 , \3101_b0 , \3102_b1 , \3102_b0 , 
		\3103_b1 , \3103_b0 , \3104_b1 , \3104_b0 , \3105_b1 , \3105_b0 , \3106_b1 , \3106_b0 , \3107_b1 , \3107_b0 , 
		\3108_b1 , \3108_b0 , \3109_b1 , \3109_b0 , \3110_b1 , \3110_b0 , \3111_b1 , \3111_b0 , \3112_b1 , \3112_b0 , 
		\3113_b1 , \3113_b0 , \3114_b1 , \3114_b0 , \3115_b1 , \3115_b0 , \3116_b1 , \3116_b0 , \3117_b1 , \3117_b0 , 
		\3118_b1 , \3118_b0 , \3119_b1 , \3119_b0 , \3120_b1 , \3120_b0 , \3121_b1 , \3121_b0 , \3122_b1 , \3122_b0 , 
		\3123_b1 , \3123_b0 , \3124_b1 , \3124_b0 , \3125_b1 , \3125_b0 , \3126_b1 , \3126_b0 , \3127_b1 , \3127_b0 , 
		\3128_b1 , \3128_b0 , \3129_b1 , \3129_b0 , \3130_b1 , \3130_b0 , \3131_b1 , \3131_b0 , \3132_b1 , \3132_b0 , 
		\3133_b1 , \3133_b0 , \3134_b1 , \3134_b0 , \3135_b1 , \3135_b0 , \3136_b1 , \3136_b0 , \3137_b1 , \3137_b0 , 
		\3138_b1 , \3138_b0 , \3139_b1 , \3139_b0 , \3140_b1 , \3140_b0 , \3141_b1 , \3141_b0 , \3142_b1 , \3142_b0 , 
		\3143_b1 , \3143_b0 , \3144_b1 , \3144_b0 , \3145_b1 , \3145_b0 , \3146_b1 , \3146_b0 , \3147_b1 , \3147_b0 , 
		\3148_b1 , \3148_b0 , \3149_b1 , \3149_b0 , \3150_b1 , \3150_b0 , \3151_b1 , \3151_b0 , \3152_b1 , \3152_b0 , 
		\3153_b1 , \3153_b0 , \3154_b1 , \3154_b0 , \3155_b1 , \3155_b0 , \3156_b1 , \3156_b0 , \3157_b1 , \3157_b0 , 
		\3158_b1 , \3158_b0 , \3159_b1 , \3159_b0 , \3160_b1 , \3160_b0 , \3161_b1 , \3161_b0 , \3162_b1 , \3162_b0 , 
		\3163_b1 , \3163_b0 , \3164_b1 , \3164_b0 , \3165_b1 , \3165_b0 , \3166_b1 , \3166_b0 , \3167_b1 , \3167_b0 , 
		\3168_b1 , \3168_b0 , \3169_b1 , \3169_b0 , \3170_b1 , \3170_b0 , \3171_b1 , \3171_b0 , \3172_b1 , \3172_b0 , 
		\3173_b1 , \3173_b0 , \3174_b1 , \3174_b0 , \3175_b1 , \3175_b0 , \3176_b1 , \3176_b0 , \3177_b1 , \3177_b0 , 
		\3178_b1 , \3178_b0 , \3179_b1 , \3179_b0 , \3180_b1 , \3180_b0 , \3181_b1 , \3181_b0 , \3182_b1 , \3182_b0 , 
		\3183_b1 , \3183_b0 , \3184_b1 , \3184_b0 , \3185_b1 , \3185_b0 , \3186_b1 , \3186_b0 , \3187_b1 , \3187_b0 , 
		\3188_b1 , \3188_b0 , \3189_b1 , \3189_b0 , \3190_b1 , \3190_b0 , \3191_b1 , \3191_b0 , \3192_b1 , \3192_b0 , 
		\3193_b1 , \3193_b0 , \3194_b1 , \3194_b0 , \3195_b1 , \3195_b0 , \3196_b1 , \3196_b0 , \3197_b1 , \3197_b0 , 
		\3198_b1 , \3198_b0 , \3199_b1 , \3199_b0 , \3200_b1 , \3200_b0 , \3201_b1 , \3201_b0 , \3202_b1 , \3202_b0 , 
		\3203_b1 , \3203_b0 , \3204_b1 , \3204_b0 , \3205_b1 , \3205_b0 , \3206_b1 , \3206_b0 , \3207_b1 , \3207_b0 , 
		\3208_b1 , \3208_b0 , \3209_b1 , \3209_b0 , \3210_b1 , \3210_b0 , \3211_b1 , \3211_b0 , \3212_b1 , \3212_b0 , 
		\3213_b1 , \3213_b0 , \3214_b1 , \3214_b0 , \3215_b1 , \3215_b0 , \3216_b1 , \3216_b0 , \3217_b1 , \3217_b0 , 
		\3218_b1 , \3218_b0 , \3219_b1 , \3219_b0 , \3220_b1 , \3220_b0 , \3221_b1 , \3221_b0 , \3222_b1 , \3222_b0 , 
		\3223_b1 , \3223_b0 , \3224_b1 , \3224_b0 , \3225_b1 , \3225_b0 , \3226_b1 , \3226_b0 , \3227_b1 , \3227_b0 , 
		\3228_b1 , \3228_b0 , \3229_b1 , \3229_b0 , \3230_b1 , \3230_b0 , \3231_b1 , \3231_b0 , \3232_b1 , \3232_b0 , 
		\3233_b1 , \3233_b0 , \3234_b1 , \3234_b0 , \3235_b1 , \3235_b0 , \3236_b1 , \3236_b0 , \3237_b1 , \3237_b0 , 
		\3238_b1 , \3238_b0 , \3239_b1 , \3239_b0 , \3240_b1 , \3240_b0 , \3241_b1 , \3241_b0 , \3242_b1 , \3242_b0 , 
		\3243_b1 , \3243_b0 , \3244_b1 , \3244_b0 , \3245_b1 , \3245_b0 , \3246_b1 , \3246_b0 , \3247_b1 , \3247_b0 , 
		\3248_b1 , \3248_b0 , \3249_b1 , \3249_b0 , \3250_b1 , \3250_b0 , \3251_b1 , \3251_b0 , \3252_b1 , \3252_b0 , 
		\3253_b1 , \3253_b0 , \3254_b1 , \3254_b0 , \3255_b1 , \3255_b0 , \3256_b1 , \3256_b0 , \3257_b1 , \3257_b0 , 
		\3258_b1 , \3258_b0 , \3259_b1 , \3259_b0 , \3260_b1 , \3260_b0 , \3261_b1 , \3261_b0 , \3262_b1 , \3262_b0 , 
		\3263_b1 , \3263_b0 , \3264_b1 , \3264_b0 , \3265_b1 , \3265_b0 , \3266_b1 , \3266_b0 , \3267_b1 , \3267_b0 , 
		\3268_b1 , \3268_b0 , \3269_b1 , \3269_b0 , \3270_b1 , \3270_b0 , \3271_b1 , \3271_b0 , \3272_b1 , \3272_b0 , 
		\3273_b1 , \3273_b0 , \3274_b1 , \3274_b0 , \3275_b1 , \3275_b0 , \3276_b1 , \3276_b0 , \3277_b1 , \3277_b0 , 
		\3278_b1 , \3278_b0 , \3279_b1 , \3279_b0 , \3280_b1 , \3280_b0 , \3281_b1 , \3281_b0 , \3282_b1 , \3282_b0 , 
		\3283_b1 , \3283_b0 , \3284_b1 , \3284_b0 , \3285_b1 , \3285_b0 , \3286_b1 , \3286_b0 , \3287_b1 , \3287_b0 , 
		\3288_b1 , \3288_b0 , \3289_b1 , \3289_b0 , \3290_b1 , \3290_b0 , \3291_b1 , \3291_b0 , \3292_b1 , \3292_b0 , 
		\3293_b1 , \3293_b0 , \3294_b1 , \3294_b0 , \3295_b1 , \3295_b0 , \3296_b1 , \3296_b0 , \3297_b1 , \3297_b0 , 
		\3298_b1 , \3298_b0 , \3299_b1 , \3299_b0 , \3300_b1 , \3300_b0 , \3301_b1 , \3301_b0 , \3302_b1 , \3302_b0 , 
		\3303_b1 , \3303_b0 , \3304_b1 , \3304_b0 , \3305_b1 , \3305_b0 , \3306_b1 , \3306_b0 , \3307_b1 , \3307_b0 , 
		\3308_b1 , \3308_b0 , \3309_b1 , \3309_b0 , \3310_b1 , \3310_b0 , \3311_b1 , \3311_b0 , \3312_b1 , \3312_b0 , 
		\3313_b1 , \3313_b0 , \3314_b1 , \3314_b0 , \3315_b1 , \3315_b0 , \3316_b1 , \3316_b0 , \3317_b1 , \3317_b0 , 
		\3318_b1 , \3318_b0 , \3319_b1 , \3319_b0 , \3320_b1 , \3320_b0 , \3321_b1 , \3321_b0 , \3322_b1 , \3322_b0 , 
		\3323_b1 , \3323_b0 , \3324_b1 , \3324_b0 , \3325_b1 , \3325_b0 , \3326_b1 , \3326_b0 , \3327_b1 , \3327_b0 , 
		\3328_b1 , \3328_b0 , \3329_b1 , \3329_b0 , \3330_b1 , \3330_b0 , \3331_b1 , \3331_b0 , \3332_b1 , \3332_b0 , 
		\3333_b1 , \3333_b0 , \3334_b1 , \3334_b0 , \3335_b1 , \3335_b0 , \3336_b1 , \3336_b0 , \3337_b1 , \3337_b0 , 
		\3338_b1 , \3338_b0 , \3339_b1 , \3339_b0 , \3340_b1 , \3340_b0 , \3341_b1 , \3341_b0 , \3342_b1 , \3342_b0 , 
		\3343_b1 , \3343_b0 , \3344_b1 , \3344_b0 , \3345_b1 , \3345_b0 , \3346_b1 , \3346_b0 , \3347_b1 , \3347_b0 , 
		\3348_b1 , \3348_b0 , \3349_b1 , \3349_b0 , \3350_b1 , \3350_b0 , \3351_b1 , \3351_b0 , \3352_b1 , \3352_b0 , 
		\3353_b1 , \3353_b0 , \3354_b1 , \3354_b0 , \3355_b1 , \3355_b0 , \3356_b1 , \3356_b0 , \3357_b1 , \3357_b0 , 
		\3358_b1 , \3358_b0 , \3359_b1 , \3359_b0 , \3360_b1 , \3360_b0 , \3361_b1 , \3361_b0 , \3362_b1 , \3362_b0 , 
		\3363_b1 , \3363_b0 , \3364_b1 , \3364_b0 , \3365_b1 , \3365_b0 , \3366_b1 , \3366_b0 , \3367_b1 , \3367_b0 , 
		\3368_b1 , \3368_b0 , \3369_b1 , \3369_b0 , \3370_b1 , \3370_b0 , \3371_b1 , \3371_b0 , \3372_b1 , \3372_b0 , 
		\3373_b1 , \3373_b0 , \3374_b1 , \3374_b0 , \3375_b1 , \3375_b0 , \3376_b1 , \3376_b0 , \3377_b1 , \3377_b0 , 
		\3378_b1 , \3378_b0 , \3379_b1 , \3379_b0 , \3380_b1 , \3380_b0 , \3381_b1 , \3381_b0 , \3382_b1 , \3382_b0 , 
		\3383_b1 , \3383_b0 , \3384_b1 , \3384_b0 , \3385_b1 , \3385_b0 , \3386_b1 , \3386_b0 , \3387_b1 , \3387_b0 , 
		\3388_b1 , \3388_b0 , \3389_b1 , \3389_b0 , \3390_b1 , \3390_b0 , \3391_b1 , \3391_b0 , \3392_b1 , \3392_b0 , 
		\3393_b1 , \3393_b0 , \3394_b1 , \3394_b0 , \3395_b1 , \3395_b0 , \3396_b1 , \3396_b0 , \3397_b1 , \3397_b0 , 
		\3398_b1 , \3398_b0 , \3399_b1 , \3399_b0 , \3400_b1 , \3400_b0 , \3401_b1 , \3401_b0 , \3402_b1 , \3402_b0 , 
		\3403_b1 , \3403_b0 , \3404_b1 , \3404_b0 , \3405_b1 , \3405_b0 , \3406_b1 , \3406_b0 , \3407_b1 , \3407_b0 , 
		\3408_b1 , \3408_b0 , \3409_b1 , \3409_b0 , \3410_b1 , \3410_b0 , \3411_b1 , \3411_b0 , \3412_b1 , \3412_b0 , 
		\3413_b1 , \3413_b0 , \3414_b1 , \3414_b0 , \3415_b1 , \3415_b0 , \3416_b1 , \3416_b0 , \3417_b1 , \3417_b0 , 
		\3418_b1 , \3418_b0 , \3419_b1 , \3419_b0 , \3420_b1 , \3420_b0 , \3421_b1 , \3421_b0 , \3422_b1 , \3422_b0 , 
		\3423_b1 , \3423_b0 , \3424_b1 , \3424_b0 , \3425_b1 , \3425_b0 , \3426_b1 , \3426_b0 , \3427_b1 , \3427_b0 , 
		\3428_b1 , \3428_b0 , \3429_b1 , \3429_b0 , \3430_b1 , \3430_b0 , \3431_b1 , \3431_b0 , \3432_b1 , \3432_b0 , 
		\3433_b1 , \3433_b0 , \3434_b1 , \3434_b0 , \3435_b1 , \3435_b0 , \3436_b1 , \3436_b0 , \3437_b1 , \3437_b0 , 
		\3438_b1 , \3438_b0 , \3439_b1 , \3439_b0 , \3440_b1 , \3440_b0 , \3441_b1 , \3441_b0 , \3442_b1 , \3442_b0 , 
		\3443_b1 , \3443_b0 , \3444_b1 , \3444_b0 , \3445_b1 , \3445_b0 , \3446_b1 , \3446_b0 , \3447_b1 , \3447_b0 , 
		\3448_b1 , \3448_b0 , \3449_b1 , \3449_b0 , \3450_b1 , \3450_b0 , \3451_b1 , \3451_b0 , \3452_b1 , \3452_b0 , 
		\3453_b1 , \3453_b0 , \3454_b1 , \3454_b0 , \3455_b1 , \3455_b0 , \3456_b1 , \3456_b0 , \3457_b1 , \3457_b0 , 
		\3458_b1 , \3458_b0 , \3459_b1 , \3459_b0 , \3460_b1 , \3460_b0 , \3461_b1 , \3461_b0 , \3462_b1 , \3462_b0 , 
		\3463_b1 , \3463_b0 , \3464_b1 , \3464_b0 , \3465_b1 , \3465_b0 , \3466_b1 , \3466_b0 , \3467_b1 , \3467_b0 , 
		\3468_b1 , \3468_b0 , \3469_b1 , \3469_b0 , \3470_b1 , \3470_b0 , \3471_b1 , \3471_b0 , \3472_b1 , \3472_b0 , 
		\3473_b1 , \3473_b0 , \3474_b1 , \3474_b0 , \3475_b1 , \3475_b0 , \3476_b1 , \3476_b0 , \3477_b1 , \3477_b0 , 
		\3478_b1 , \3478_b0 , \3479_b1 , \3479_b0 , \3480_b1 , \3480_b0 , \3481_b1 , \3481_b0 , \3482_b1 , \3482_b0 , 
		\3483_b1 , \3483_b0 , \3484_b1 , \3484_b0 , \3485_b1 , \3485_b0 , \3486_b1 , \3486_b0 , \3487_b1 , \3487_b0 , 
		\3488_b1 , \3488_b0 , \3489_b1 , \3489_b0 , \3490_b1 , \3490_b0 , \3491_b1 , \3491_b0 , \3492_b1 , \3492_b0 , 
		\3493_b1 , \3493_b0 , \3494_b1 , \3494_b0 , \3495_b1 , \3495_b0 , \3496_b1 , \3496_b0 , \3497_b1 , \3497_b0 , 
		\3498_b1 , \3498_b0 , \3499_b1 , \3499_b0 , \3500_b1 , \3500_b0 , \3501_b1 , \3501_b0 , \3502_b1 , \3502_b0 , 
		\3503_b1 , \3503_b0 , \3504_b1 , \3504_b0 , \3505_b1 , \3505_b0 , \3506_b1 , \3506_b0 , \3507_b1 , \3507_b0 , 
		\3508_b1 , \3508_b0 , \3509_b1 , \3509_b0 , \3510_b1 , \3510_b0 , \3511_b1 , \3511_b0 , \3512_b1 , \3512_b0 , 
		\3513_b1 , \3513_b0 , \3514_b1 , \3514_b0 , \3515_b1 , \3515_b0 , \3516_b1 , \3516_b0 , \3517_b1 , \3517_b0 , 
		\3518_b1 , \3518_b0 , \3519_b1 , \3519_b0 , \3520_b1 , \3520_b0 , \3521_b1 , \3521_b0 , \3522_b1 , \3522_b0 , 
		\3523_b1 , \3523_b0 , \3524_b1 , \3524_b0 , \3525_b1 , \3525_b0 , \3526_b1 , \3526_b0 , \3527_b1 , \3527_b0 , 
		\3528_b1 , \3528_b0 , \3529_b1 , \3529_b0 , \3530_b1 , \3530_b0 , \3531_b1 , \3531_b0 , \3532_b1 , \3532_b0 , 
		\3533_b1 , \3533_b0 , \3534_b1 , \3534_b0 , \3535_b1 , \3535_b0 , \3536_b1 , \3536_b0 , \3537_b1 , \3537_b0 , 
		\3538_b1 , \3538_b0 , \3539_b1 , \3539_b0 , \3540_b1 , \3540_b0 , \3541_b1 , \3541_b0 , \3542_b1 , \3542_b0 , 
		\3543_b1 , \3543_b0 , \3544_b1 , \3544_b0 , \3545_b1 , \3545_b0 , \3546_b1 , \3546_b0 , \3547_b1 , \3547_b0 , 
		\3548_b1 , \3548_b0 , \3549_b1 , \3549_b0 , \3550_b1 , \3550_b0 , \3551_b1 , \3551_b0 , \3552_b1 , \3552_b0 , 
		\3553_b1 , \3553_b0 , \3554_b1 , \3554_b0 , \3555_b1 , \3555_b0 , \3556_b1 , \3556_b0 , \3557_b1 , \3557_b0 , 
		\3558_b1 , \3558_b0 , \3559_b1 , \3559_b0 , \3560_b1 , \3560_b0 , \3561_b1 , \3561_b0 , \3562_b1 , \3562_b0 , 
		\3563_b1 , \3563_b0 , \3564_b1 , \3564_b0 , \3565_b1 , \3565_b0 , \3566_b1 , \3566_b0 , \3567_b1 , \3567_b0 , 
		\3568_b1 , \3568_b0 , \3569_b1 , \3569_b0 , \3570_b1 , \3570_b0 , \3571_b1 , \3571_b0 , \3572_b1 , \3572_b0 , 
		\3573_b1 , \3573_b0 , \3574_b1 , \3574_b0 , \3575_b1 , \3575_b0 , \3576_b1 , \3576_b0 , \3577_b1 , \3577_b0 , 
		\3578_b1 , \3578_b0 , \3579_b1 , \3579_b0 , \3580_b1 , \3580_b0 , \3581_b1 , \3581_b0 , \3582_b1 , \3582_b0 , 
		\3583_b1 , \3583_b0 , \3584_b1 , \3584_b0 , \3585_b1 , \3585_b0 , \3586_b1 , \3586_b0 , \3587_b1 , \3587_b0 , 
		\3588_b1 , \3588_b0 , \3589_b1 , \3589_b0 , \3590_b1 , \3590_b0 , \3591_b1 , \3591_b0 , \3592_b1 , \3592_b0 , 
		\3593_b1 , \3593_b0 , \3594_b1 , \3594_b0 , \3595_b1 , \3595_b0 , \3596_b1 , \3596_b0 , \3597_b1 , \3597_b0 , 
		\3598_b1 , \3598_b0 , \3599_b1 , \3599_b0 , \3600_b1 , \3600_b0 , \3601_b1 , \3601_b0 , \3602_b1 , \3602_b0 , 
		\3603_b1 , \3603_b0 , \3604_b1 , \3604_b0 , \3605_b1 , \3605_b0 , \3606_b1 , \3606_b0 , \3607_b1 , \3607_b0 , 
		\3608_b1 , \3608_b0 , \3609_b1 , \3609_b0 , \3610_b1 , \3610_b0 , \3611_b1 , \3611_b0 , \3612_b1 , \3612_b0 , 
		\3613_b1 , \3613_b0 , \3614_b1 , \3614_b0 , \3615_b1 , \3615_b0 , \3616_b1 , \3616_b0 , \3617_b1 , \3617_b0 , 
		\3618_b1 , \3618_b0 , \3619_b1 , \3619_b0 , \3620_b1 , \3620_b0 , \3621_b1 , \3621_b0 , \3622_b1 , \3622_b0 , 
		\3623_b1 , \3623_b0 , \3624_b1 , \3624_b0 , \3625_b1 , \3625_b0 , \3626_b1 , \3626_b0 , \3627_b1 , \3627_b0 , 
		\3628_b1 , \3628_b0 , \3629_b1 , \3629_b0 , \3630_b1 , \3630_b0 , \3631_b1 , \3631_b0 , \3632_b1 , \3632_b0 , 
		\3633_b1 , \3633_b0 , \3634_b1 , \3634_b0 , \3635_b1 , \3635_b0 , \3636_b1 , \3636_b0 , \3637_b1 , \3637_b0 , 
		\3638_b1 , \3638_b0 , \3639_b1 , \3639_b0 , \3640_b1 , \3640_b0 , \3641_b1 , \3641_b0 , \3642_b1 , \3642_b0 , 
		\3643_b1 , \3643_b0 , \3644_b1 , \3644_b0 , \3645_b1 , \3645_b0 , \3646_b1 , \3646_b0 , \3647_b1 , \3647_b0 , 
		\3648_b1 , \3648_b0 , \3649_b1 , \3649_b0 , \3650_b1 , \3650_b0 , \3651_b1 , \3651_b0 , \3652_b1 , \3652_b0 , 
		\3653_b1 , \3653_b0 , \3654_b1 , \3654_b0 , \3655_b1 , \3655_b0 , \3656_b1 , \3656_b0 , \3657_b1 , \3657_b0 , 
		\3658_b1 , \3658_b0 , \3659_b1 , \3659_b0 , \3660_b1 , \3660_b0 , \3661_b1 , \3661_b0 , \3662_b1 , \3662_b0 , 
		\3663_b1 , \3663_b0 , \3664_b1 , \3664_b0 , \3665_b1 , \3665_b0 , \3666_b1 , \3666_b0 , \3667_b1 , \3667_b0 , 
		\3668_b1 , \3668_b0 , \3669_b1 , \3669_b0 , \3670_b1 , \3670_b0 , \3671_b1 , \3671_b0 , \3672_b1 , \3672_b0 , 
		\3673_b1 , \3673_b0 , \3674_b1 , \3674_b0 , \3675_b1 , \3675_b0 , \3676_b1 , \3676_b0 , \3677_b1 , \3677_b0 , 
		\3678_b1 , \3678_b0 , \3679_b1 , \3679_b0 , \3680_b1 , \3680_b0 , \3681_b1 , \3681_b0 , \3682_b1 , \3682_b0 , 
		\3683_b1 , \3683_b0 , \3684_b1 , \3684_b0 , \3685_b1 , \3685_b0 , \3686_b1 , \3686_b0 , \3687_b1 , \3687_b0 , 
		\3688_b1 , \3688_b0 , \3689_b1 , \3689_b0 , \3690_b1 , \3690_b0 , \3691_b1 , \3691_b0 , \3692_b1 , \3692_b0 , 
		\3693_b1 , \3693_b0 , \3694_b1 , \3694_b0 , \3695_b1 , \3695_b0 , \3696_b1 , \3696_b0 , \3697_b1 , \3697_b0 , 
		\3698_b1 , \3698_b0 , \3699_b1 , \3699_b0 , \3700_b1 , \3700_b0 , \3701_b1 , \3701_b0 , \3702_b1 , \3702_b0 , 
		\3703_b1 , \3703_b0 , \3704_b1 , \3704_b0 , \3705_b1 , \3705_b0 , \3706_b1 , \3706_b0 , \3707_b1 , \3707_b0 , 
		\3708_b1 , \3708_b0 , \3709_b1 , \3709_b0 , \3710_b1 , \3710_b0 , \3711_b1 , \3711_b0 , \3712_b1 , \3712_b0 , 
		\3713_b1 , \3713_b0 , \3714_b1 , \3714_b0 , \3715_b1 , \3715_b0 , \3716_b1 , \3716_b0 , \3717_b1 , \3717_b0 , 
		\3718_b1 , \3718_b0 , \3719_b1 , \3719_b0 , \3720_b1 , \3720_b0 , \3721_b1 , \3721_b0 , \3722_b1 , \3722_b0 , 
		\3723_b1 , \3723_b0 , \3724_b1 , \3724_b0 , \3725_b1 , \3725_b0 , \3726_b1 , \3726_b0 , \3727_b1 , \3727_b0 , 
		\3728_b1 , \3728_b0 , \3729_b1 , \3729_b0 , \3730_b1 , \3730_b0 , \3731_b1 , \3731_b0 , \3732_b1 , \3732_b0 , 
		\3733_b1 , \3733_b0 , \3734_b1 , \3734_b0 , \3735_b1 , \3735_b0 , \3736_b1 , \3736_b0 , \3737_b1 , \3737_b0 , 
		\3738_b1 , \3738_b0 , \3739_b1 , \3739_b0 , \3740_b1 , \3740_b0 , \3741_b1 , \3741_b0 , \3742_b1 , \3742_b0 , 
		\3743_b1 , \3743_b0 , \3744_b1 , \3744_b0 , \3745_b1 , \3745_b0 , \3746_b1 , \3746_b0 , \3747_b1 , \3747_b0 , 
		\3748_b1 , \3748_b0 , \3749_b1 , \3749_b0 , \3750_b1 , \3750_b0 , \3751_b1 , \3751_b0 , \3752_b1 , \3752_b0 , 
		\3753_b1 , \3753_b0 , \3754_b1 , \3754_b0 , \3755_b1 , \3755_b0 , \3756_b1 , \3756_b0 , \3757_b1 , \3757_b0 , 
		\3758_b1 , \3758_b0 , \3759_b1 , \3759_b0 , \3760_b1 , \3760_b0 , \3761_b1 , \3761_b0 , \3762_b1 , \3762_b0 , 
		\3763_b1 , \3763_b0 , \3764_b1 , \3764_b0 , \3765_b1 , \3765_b0 , \3766_b1 , \3766_b0 , \3767_b1 , \3767_b0 , 
		\3768_b1 , \3768_b0 , \3769_b1 , \3769_b0 , \3770_b1 , \3770_b0 , \3771_b1 , \3771_b0 , \3772_b1 , \3772_b0 , 
		\3773_b1 , \3773_b0 , \3774_b1 , \3774_b0 , \3775_b1 , \3775_b0 , \3776_b1 , \3776_b0 , \3777_b1 , \3777_b0 , 
		\3778_b1 , \3778_b0 , \3779_b1 , \3779_b0 , \3780_b1 , \3780_b0 , \3781_b1 , \3781_b0 , \3782_b1 , \3782_b0 , 
		\3783_b1 , \3783_b0 , \3784_b1 , \3784_b0 , \3785_b1 , \3785_b0 , \3786_b1 , \3786_b0 , \3787_b1 , \3787_b0 , 
		\3788_b1 , \3788_b0 , \3789_b1 , \3789_b0 , \3790_b1 , \3790_b0 , \3791_b1 , \3791_b0 , \3792_b1 , \3792_b0 , 
		\3793_b1 , \3793_b0 , \3794_b1 , \3794_b0 , \3795_b1 , \3795_b0 , \3796_b1 , \3796_b0 , \3797_b1 , \3797_b0 , 
		\3798_b1 , \3798_b0 , \3799_b1 , \3799_b0 , \3800_b1 , \3800_b0 , \3801_b1 , \3801_b0 , \3802_b1 , \3802_b0 , 
		\3803_b1 , \3803_b0 , \3804_b1 , \3804_b0 , \3805_b1 , \3805_b0 , \3806_b1 , \3806_b0 , \3807_b1 , \3807_b0 , 
		\3808_b1 , \3808_b0 , \3809_b1 , \3809_b0 , \3810_b1 , \3810_b0 , \3811_b1 , \3811_b0 , \3812_b1 , \3812_b0 , 
		\3813_b1 , \3813_b0 , \3814_b1 , \3814_b0 , \3815_b1 , \3815_b0 , \3816_b1 , \3816_b0 , \3817_b1 , \3817_b0 , 
		\3818_b1 , \3818_b0 , \3819_b1 , \3819_b0 , \3820_b1 , \3820_b0 , \3821_b1 , \3821_b0 , \3822_b1 , \3822_b0 , 
		\3823_b1 , \3823_b0 , \3824_b1 , \3824_b0 , \3825_b1 , \3825_b0 , \3826_b1 , \3826_b0 , \3827_b1 , \3827_b0 , 
		\3828_b1 , \3828_b0 , \3829_b1 , \3829_b0 , \3830_b1 , \3830_b0 , \3831_b1 , \3831_b0 , \3832_b1 , \3832_b0 , 
		\3833_b1 , \3833_b0 , \3834_b1 , \3834_b0 , \3835_b1 , \3835_b0 , \3836_b1 , \3836_b0 , \3837_b1 , \3837_b0 , 
		\3838_b1 , \3838_b0 , \3839_b1 , \3839_b0 , \3840_b1 , \3840_b0 , \3841_b1 , \3841_b0 , \3842_b1 , \3842_b0 , 
		\3843_b1 , \3843_b0 , \3844_b1 , \3844_b0 , \3845_b1 , \3845_b0 , \3846_b1 , \3846_b0 , \3847_b1 , \3847_b0 , 
		\3848_b1 , \3848_b0 , \3849_b1 , \3849_b0 , \3850_b1 , \3850_b0 , \3851_b1 , \3851_b0 , \3852_b1 , \3852_b0 , 
		\3853_b1 , \3853_b0 , \3854_b1 , \3854_b0 , \3855_b1 , \3855_b0 , \3856_b1 , \3856_b0 , \3857_b1 , \3857_b0 , 
		\3858_b1 , \3858_b0 , \3859_b1 , \3859_b0 , \3860_b1 , \3860_b0 , \3861_b1 , \3861_b0 , \3862_b1 , \3862_b0 , 
		\3863_b1 , \3863_b0 , \3864_b1 , \3864_b0 , \3865_b1 , \3865_b0 , \3866_b1 , \3866_b0 , \3867_b1 , \3867_b0 , 
		\3868_b1 , \3868_b0 , \3869_b1 , \3869_b0 , \3870_b1 , \3870_b0 , \3871_b1 , \3871_b0 , \3872_b1 , \3872_b0 , 
		\3873_b1 , \3873_b0 , \3874_b1 , \3874_b0 , \3875_b1 , \3875_b0 , \3876_b1 , \3876_b0 , \3877_b1 , \3877_b0 , 
		\3878_b1 , \3878_b0 , \3879_b1 , \3879_b0 , \3880_b1 , \3880_b0 , \3881_b1 , \3881_b0 , \3882_b1 , \3882_b0 , 
		\3883_b1 , \3883_b0 , \3884_b1 , \3884_b0 , \3885_b1 , \3885_b0 , \3886_b1 , \3886_b0 , \3887_b1 , \3887_b0 , 
		\3888_b1 , \3888_b0 , \3889_b1 , \3889_b0 , \3890_b1 , \3890_b0 , \3891_b1 , \3891_b0 , \3892_b1 , \3892_b0 , 
		\3893_b1 , \3893_b0 , \3894_b1 , \3894_b0 , \3895_b1 , \3895_b0 , \3896_b1 , \3896_b0 , \3897_b1 , \3897_b0 , 
		\3898_b1 , \3898_b0 , \3899_b1 , \3899_b0 , \3900_b1 , \3900_b0 , \3901_b1 , \3901_b0 , \3902_b1 , \3902_b0 , 
		\3903_b1 , \3903_b0 , \3904_b1 , \3904_b0 , \3905_b1 , \3905_b0 , \3906_b1 , \3906_b0 , \3907_b1 , \3907_b0 , 
		\3908_b1 , \3908_b0 , \3909_b1 , \3909_b0 , \3910_b1 , \3910_b0 , \3911_b1 , \3911_b0 , \3912_b1 , \3912_b0 , 
		\3913_b1 , \3913_b0 , \3914_b1 , \3914_b0 , \3915_b1 , \3915_b0 , \3916_b1 , \3916_b0 , \3917_b1 , \3917_b0 , 
		\3918_b1 , \3918_b0 , \3919_b1 , \3919_b0 , \3920_b1 , \3920_b0 , \3921_b1 , \3921_b0 , \3922_b1 , \3922_b0 , 
		\3923_b1 , \3923_b0 , \3924_b1 , \3924_b0 , \3925_b1 , \3925_b0 , \3926_b1 , \3926_b0 , \3927_Z[31]_b1 , \3927_Z[31]_b0 , 
		\3928_b1 , \3928_b0 , \3929_Z[30]_b1 , \3929_Z[30]_b0 , \3930_b1 , \3930_b0 , \3931_Z[29]_b1 , \3931_Z[29]_b0 , \3932_b1 , \3932_b0 , 
		\3933_Z[28]_b1 , \3933_Z[28]_b0 , \3934_b1 , \3934_b0 , \3935_Z[27]_b1 , \3935_Z[27]_b0 , \3936_b1 , \3936_b0 , \3937_Z[26]_b1 , \3937_Z[26]_b0 , 
		\3938_b1 , \3938_b0 , \3939_Z[25]_b1 , \3939_Z[25]_b0 , \3940_b1 , \3940_b0 , \3941_Z[24]_b1 , \3941_Z[24]_b0 , \3942_b1 , \3942_b0 , 
		\3943_Z[23]_b1 , \3943_Z[23]_b0 , \3944_b1 , \3944_b0 , \3945_Z[22]_b1 , \3945_Z[22]_b0 , \3946_b1 , \3946_b0 , \3947_Z[21]_b1 , \3947_Z[21]_b0 , 
		\3948_b1 , \3948_b0 , \3949_Z[20]_b1 , \3949_Z[20]_b0 , \3950_b1 , \3950_b0 , \3951_Z[19]_b1 , \3951_Z[19]_b0 , \3952_b1 , \3952_b0 , 
		\3953_Z[18]_b1 , \3953_Z[18]_b0 , \3954_b1 , \3954_b0 , \3955_Z[17]_b1 , \3955_Z[17]_b0 , \3956_b1 , \3956_b0 , \3957_Z[16]_b1 , \3957_Z[16]_b0 , 
		\3958_b1 , \3958_b0 , \3959_Z[15]_b1 , \3959_Z[15]_b0 , \3960_b1 , \3960_b0 , \3961_Z[14]_b1 , \3961_Z[14]_b0 , \3962_b1 , \3962_b0 , 
		\3963_Z[13]_b1 , \3963_Z[13]_b0 , \3964_b1 , \3964_b0 , \3965_Z[12]_b1 , \3965_Z[12]_b0 , \3966_b1 , \3966_b0 , \3967_Z[11]_b1 , \3967_Z[11]_b0 , 
		\3968_b1 , \3968_b0 , \3969_Z[10]_b1 , \3969_Z[10]_b0 , \3970_b1 , \3970_b0 , \3971_Z[9]_b1 , \3971_Z[9]_b0 , \3972_b1 , \3972_b0 , 
		\3973_Z[8]_b1 , \3973_Z[8]_b0 , \3974_b1 , \3974_b0 , \3975_Z[7]_b1 , \3975_Z[7]_b0 , \3976_b1 , \3976_b0 , \3977_Z[6]_b1 , \3977_Z[6]_b0 , 
		\3978_b1 , \3978_b0 , \3979_Z[5]_b1 , \3979_Z[5]_b0 , \3980_b1 , \3980_b0 , \3981_Z[4]_b1 , \3981_Z[4]_b0 , \3982_b1 , \3982_b0 , 
		\3983_Z[3]_b1 , \3983_Z[3]_b0 , \3984_b1 , \3984_b0 , \3985_Z[2]_b1 , \3985_Z[2]_b0 , \3986_b1 , \3986_b0 , \3987_Z[1]_b1 , \3987_Z[1]_b0 , 
		\3988_b1 , \3988_b0 , \3989_Z[0]_b1 , \3989_Z[0]_b0 , w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , 
		w_6 , w_7 , w_8 , w_9 , w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , 
		w_16 , w_17 , w_18 , w_19 , w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , 
		w_26 , w_27 , w_28 , w_29 , w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , 
		w_36 , w_37 , w_38 , w_39 , w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , 
		w_46 , w_47 , w_48 , w_49 , w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , 
		w_56 , w_57 , w_58 , w_59 , w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , 
		w_66 , w_67 , w_68 , w_69 , w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , 
		w_76 , w_77 , w_78 , w_79 , w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , 
		w_86 , w_87 , w_88 , w_89 , w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , 
		w_96 , w_97 , w_98 , w_99 , w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , 
		w_106 , w_107 , w_108 , w_109 , w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , 
		w_116 , w_117 , w_118 , w_119 , w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , 
		w_126 , w_127 , w_128 , w_129 , w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , 
		w_136 , w_137 , w_138 , w_139 , w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , 
		w_146 , w_147 , w_148 , w_149 , w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , 
		w_156 , w_157 , w_158 , w_159 , w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , 
		w_166 , w_167 , w_168 , w_169 , w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , 
		w_176 , w_177 , w_178 , w_179 , w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , 
		w_186 , w_187 , w_188 , w_189 , w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , 
		w_196 , w_197 , w_198 , w_199 , w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , 
		w_206 , w_207 , w_208 , w_209 , w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , 
		w_216 , w_217 , w_218 , w_219 , w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , 
		w_226 , w_227 , w_228 , w_229 , w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , 
		w_236 , w_237 , w_238 , w_239 , w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , 
		w_246 , w_247 , w_248 , w_249 , w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , 
		w_256 , w_257 , w_258 , w_259 , w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , 
		w_266 , w_267 , w_268 , w_269 , w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , 
		w_276 , w_277 , w_278 , w_279 , w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , 
		w_286 , w_287 , w_288 , w_289 , w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , 
		w_296 , w_297 , w_298 , w_299 , w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , 
		w_306 , w_307 , w_308 , w_309 , w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , 
		w_316 , w_317 , w_318 , w_319 , w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , 
		w_326 , w_327 , w_328 , w_329 , w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , 
		w_336 , w_337 , w_338 , w_339 , w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , 
		w_346 , w_347 , w_348 , w_349 , w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , 
		w_356 , w_357 , w_358 , w_359 , w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , 
		w_366 , w_367 , w_368 , w_369 , w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , 
		w_376 , w_377 , w_378 , w_379 , w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , 
		w_386 , w_387 , w_388 , w_389 , w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , 
		w_396 , w_397 , w_398 , w_399 , w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , 
		w_406 , w_407 , w_408 , w_409 , w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , 
		w_416 , w_417 , w_418 , w_419 , w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , 
		w_426 , w_427 , w_428 , w_429 , w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , 
		w_436 , w_437 , w_438 , w_439 , w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , 
		w_446 , w_447 , w_448 , w_449 , w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , 
		w_456 , w_457 , w_458 , w_459 , w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , 
		w_466 , w_467 , w_468 , w_469 , w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , 
		w_476 , w_477 , w_478 , w_479 , w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , 
		w_486 , w_487 , w_488 , w_489 , w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , 
		w_496 , w_497 , w_498 , w_499 , w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , 
		w_506 , w_507 , w_508 , w_509 , w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , 
		w_516 , w_517 , w_518 , w_519 , w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , 
		w_526 , w_527 , w_528 , w_529 , w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , 
		w_536 , w_537 , w_538 , w_539 , w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , 
		w_546 , w_547 , w_548 , w_549 , w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , 
		w_556 , w_557 , w_558 , w_559 , w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , 
		w_566 , w_567 , w_568 , w_569 , w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , 
		w_576 , w_577 , w_578 , w_579 , w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , 
		w_586 , w_587 , w_588 , w_589 , w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , 
		w_596 , w_597 , w_598 , w_599 , w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , 
		w_606 , w_607 , w_608 , w_609 , w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , 
		w_616 , w_617 , w_618 , w_619 , w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , 
		w_626 , w_627 , w_628 , w_629 , w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , 
		w_636 , w_637 , w_638 , w_639 , w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , 
		w_646 , w_647 , w_648 , w_649 , w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , 
		w_656 , w_657 , w_658 , w_659 , w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , 
		w_666 , w_667 , w_668 , w_669 , w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , 
		w_676 , w_677 , w_678 , w_679 , w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , 
		w_686 , w_687 , w_688 , w_689 , w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , 
		w_696 , w_697 , w_698 , w_699 , w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , 
		w_706 , w_707 , w_708 , w_709 , w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , 
		w_716 , w_717 , w_718 , w_719 , w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , 
		w_726 , w_727 , w_728 , w_729 , w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , 
		w_736 , w_737 , w_738 , w_739 , w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , 
		w_746 , w_747 , w_748 , w_749 , w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , 
		w_756 , w_757 , w_758 , w_759 , w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , 
		w_766 , w_767 , w_768 , w_769 , w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , 
		w_776 , w_777 , w_778 , w_779 , w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , 
		w_786 , w_787 , w_788 , w_789 , w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , 
		w_796 , w_797 , w_798 , w_799 , w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , 
		w_806 , w_807 , w_808 , w_809 , w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , 
		w_816 , w_817 , w_818 , w_819 , w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , 
		w_826 , w_827 , w_828 , w_829 , w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , 
		w_836 , w_837 , w_838 , w_839 , w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , 
		w_846 , w_847 , w_848 , w_849 , w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , 
		w_856 , w_857 , w_858 , w_859 , w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , 
		w_866 , w_867 , w_868 , w_869 , w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , 
		w_876 , w_877 , w_878 , w_879 , w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , 
		w_886 , w_887 , w_888 , w_889 , w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , 
		w_896 , w_897 , w_898 , w_899 , w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , 
		w_906 , w_907 , w_908 , w_909 , w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , 
		w_916 , w_917 , w_918 , w_919 , w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , 
		w_926 , w_927 , w_928 , w_929 , w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , 
		w_936 , w_937 , w_938 , w_939 , w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , 
		w_946 , w_947 , w_948 , w_949 , w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , 
		w_956 , w_957 , w_958 , w_959 , w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , 
		w_966 , w_967 , w_968 , w_969 , w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , 
		w_976 , w_977 , w_978 , w_979 , w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , 
		w_986 , w_987 , w_988 , w_989 , w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , 
		w_996 , w_997 , w_998 , w_999 , w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , 
		w_1006 , w_1007 , w_1008 , w_1009 , w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , 
		w_1016 , w_1017 , w_1018 , w_1019 , w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , 
		w_1026 , w_1027 , w_1028 , w_1029 , w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , 
		w_1036 , w_1037 , w_1038 , w_1039 , w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , 
		w_1046 , w_1047 , w_1048 , w_1049 , w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , 
		w_1056 , w_1057 , w_1058 , w_1059 , w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , 
		w_1066 , w_1067 , w_1068 , w_1069 , w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , 
		w_1076 , w_1077 , w_1078 , w_1079 , w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , 
		w_1086 , w_1087 , w_1088 , w_1089 , w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , 
		w_1096 , w_1097 , w_1098 , w_1099 , w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , 
		w_1106 , w_1107 , w_1108 , w_1109 , w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , 
		w_1116 , w_1117 , w_1118 , w_1119 , w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , 
		w_1126 , w_1127 , w_1128 , w_1129 , w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , 
		w_1136 , w_1137 , w_1138 , w_1139 , w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , 
		w_1146 , w_1147 , w_1148 , w_1149 , w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , 
		w_1156 , w_1157 , w_1158 , w_1159 , w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , 
		w_1166 , w_1167 , w_1168 , w_1169 , w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , 
		w_1176 , w_1177 , w_1178 , w_1179 , w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , 
		w_1186 , w_1187 , w_1188 , w_1189 , w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , 
		w_1196 , w_1197 , w_1198 , w_1199 , w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , 
		w_1206 , w_1207 , w_1208 , w_1209 , w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , 
		w_1216 , w_1217 , w_1218 , w_1219 , w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , 
		w_1226 , w_1227 , w_1228 , w_1229 , w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , 
		w_1236 , w_1237 , w_1238 , w_1239 , w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , 
		w_1246 , w_1247 , w_1248 , w_1249 , w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , 
		w_1256 , w_1257 , w_1258 , w_1259 , w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , 
		w_1266 , w_1267 , w_1268 , w_1269 , w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , 
		w_1276 , w_1277 , w_1278 , w_1279 , w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , 
		w_1286 , w_1287 , w_1288 , w_1289 , w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , 
		w_1296 , w_1297 , w_1298 , w_1299 , w_1300 , w_1301 , w_1302 , w_1303 , w_1304 , w_1305 , 
		w_1306 , w_1307 , w_1308 , w_1309 , w_1310 , w_1311 , w_1312 , w_1313 , w_1314 , w_1315 , 
		w_1316 , w_1317 , w_1318 , w_1319 , w_1320 , w_1321 , w_1322 , w_1323 , w_1324 , w_1325 , 
		w_1326 , w_1327 , w_1328 , w_1329 , w_1330 , w_1331 , w_1332 , w_1333 , w_1334 , w_1335 , 
		w_1336 , w_1337 , w_1338 , w_1339 , w_1340 , w_1341 , w_1342 , w_1343 , w_1344 , w_1345 , 
		w_1346 , w_1347 , w_1348 , w_1349 , w_1350 , w_1351 , w_1352 , w_1353 , w_1354 , w_1355 , 
		w_1356 , w_1357 , w_1358 , w_1359 , w_1360 , w_1361 , w_1362 , w_1363 , w_1364 , w_1365 , 
		w_1366 , w_1367 , w_1368 , w_1369 , w_1370 , w_1371 , w_1372 , w_1373 , w_1374 , w_1375 , 
		w_1376 , w_1377 , w_1378 , w_1379 , w_1380 , w_1381 , w_1382 , w_1383 , w_1384 , w_1385 , 
		w_1386 , w_1387 , w_1388 , w_1389 , w_1390 , w_1391 , w_1392 , w_1393 , w_1394 , w_1395 , 
		w_1396 , w_1397 , w_1398 , w_1399 , w_1400 , w_1401 , w_1402 , w_1403 , w_1404 , w_1405 , 
		w_1406 , w_1407 , w_1408 , w_1409 , w_1410 , w_1411 , w_1412 , w_1413 , w_1414 , w_1415 , 
		w_1416 , w_1417 , w_1418 , w_1419 , w_1420 , w_1421 , w_1422 , w_1423 , w_1424 , w_1425 , 
		w_1426 , w_1427 , w_1428 , w_1429 , w_1430 , w_1431 , w_1432 , w_1433 , w_1434 , w_1435 , 
		w_1436 , w_1437 , w_1438 , w_1439 , w_1440 , w_1441 , w_1442 , w_1443 , w_1444 , w_1445 , 
		w_1446 , w_1447 , w_1448 , w_1449 , w_1450 , w_1451 , w_1452 , w_1453 , w_1454 , w_1455 , 
		w_1456 , w_1457 , w_1458 , w_1459 , w_1460 , w_1461 , w_1462 , w_1463 , w_1464 , w_1465 , 
		w_1466 , w_1467 , w_1468 , w_1469 , w_1470 , w_1471 , w_1472 , w_1473 , w_1474 , w_1475 , 
		w_1476 , w_1477 , w_1478 , w_1479 , w_1480 , w_1481 , w_1482 , w_1483 , w_1484 , w_1485 , 
		w_1486 , w_1487 , w_1488 , w_1489 , w_1490 , w_1491 , w_1492 , w_1493 , w_1494 , w_1495 , 
		w_1496 , w_1497 , w_1498 , w_1499 , w_1500 , w_1501 , w_1502 , w_1503 , w_1504 , w_1505 , 
		w_1506 , w_1507 , w_1508 , w_1509 , w_1510 , w_1511 , w_1512 , w_1513 , w_1514 , w_1515 , 
		w_1516 , w_1517 , w_1518 , w_1519 , w_1520 , w_1521 , w_1522 , w_1523 , w_1524 , w_1525 , 
		w_1526 , w_1527 , w_1528 , w_1529 , w_1530 , w_1531 , w_1532 , w_1533 , w_1534 , w_1535 , 
		w_1536 , w_1537 , w_1538 , w_1539 , w_1540 , w_1541 , w_1542 , w_1543 , w_1544 , w_1545 , 
		w_1546 , w_1547 , w_1548 , w_1549 , w_1550 , w_1551 , w_1552 , w_1553 , w_1554 , w_1555 , 
		w_1556 , w_1557 , w_1558 , w_1559 , w_1560 , w_1561 , w_1562 , w_1563 , w_1564 , w_1565 , 
		w_1566 , w_1567 , w_1568 , w_1569 , w_1570 , w_1571 , w_1572 , w_1573 , w_1574 , w_1575 , 
		w_1576 , w_1577 , w_1578 , w_1579 , w_1580 , w_1581 , w_1582 , w_1583 , w_1584 , w_1585 , 
		w_1586 , w_1587 , w_1588 , w_1589 , w_1590 , w_1591 , w_1592 , w_1593 , w_1594 , w_1595 , 
		w_1596 , w_1597 , w_1598 , w_1599 , w_1600 , w_1601 , w_1602 , w_1603 , w_1604 , w_1605 , 
		w_1606 , w_1607 , w_1608 , w_1609 , w_1610 , w_1611 , w_1612 , w_1613 , w_1614 , w_1615 , 
		w_1616 , w_1617 , w_1618 , w_1619 , w_1620 , w_1621 , w_1622 , w_1623 , w_1624 , w_1625 , 
		w_1626 , w_1627 , w_1628 , w_1629 , w_1630 , w_1631 , w_1632 , w_1633 , w_1634 , w_1635 , 
		w_1636 , w_1637 , w_1638 , w_1639 , w_1640 , w_1641 , w_1642 , w_1643 , w_1644 , w_1645 , 
		w_1646 , w_1647 , w_1648 , w_1649 , w_1650 , w_1651 , w_1652 , w_1653 , w_1654 , w_1655 , 
		w_1656 , w_1657 , w_1658 , w_1659 , w_1660 , w_1661 , w_1662 , w_1663 , w_1664 , w_1665 , 
		w_1666 , w_1667 , w_1668 , w_1669 , w_1670 , w_1671 , w_1672 , w_1673 , w_1674 , w_1675 , 
		w_1676 , w_1677 , w_1678 , w_1679 , w_1680 , w_1681 , w_1682 , w_1683 , w_1684 , w_1685 , 
		w_1686 , w_1687 , w_1688 , w_1689 , w_1690 , w_1691 , w_1692 , w_1693 , w_1694 , w_1695 , 
		w_1696 , w_1697 , w_1698 , w_1699 , w_1700 , w_1701 , w_1702 , w_1703 , w_1704 , w_1705 , 
		w_1706 , w_1707 , w_1708 , w_1709 , w_1710 , w_1711 , w_1712 , w_1713 , w_1714 , w_1715 , 
		w_1716 , w_1717 , w_1718 , w_1719 , w_1720 , w_1721 , w_1722 , w_1723 , w_1724 , w_1725 , 
		w_1726 , w_1727 , w_1728 , w_1729 , w_1730 , w_1731 , w_1732 , w_1733 , w_1734 , w_1735 , 
		w_1736 , w_1737 , w_1738 , w_1739 , w_1740 , w_1741 , w_1742 , w_1743 , w_1744 , w_1745 , 
		w_1746 , w_1747 , w_1748 , w_1749 , w_1750 , w_1751 , w_1752 , w_1753 , w_1754 , w_1755 , 
		w_1756 , w_1757 , w_1758 , w_1759 , w_1760 , w_1761 , w_1762 , w_1763 , w_1764 , w_1765 , 
		w_1766 , w_1767 , w_1768 , w_1769 , w_1770 , w_1771 , w_1772 , w_1773 , w_1774 , w_1775 , 
		w_1776 , w_1777 , w_1778 , w_1779 , w_1780 , w_1781 , w_1782 , w_1783 , w_1784 , w_1785 , 
		w_1786 , w_1787 , w_1788 , w_1789 , w_1790 , w_1791 , w_1792 , w_1793 , w_1794 , w_1795 , 
		w_1796 , w_1797 , w_1798 , w_1799 , w_1800 , w_1801 , w_1802 , w_1803 , w_1804 , w_1805 , 
		w_1806 , w_1807 , w_1808 , w_1809 , w_1810 , w_1811 , w_1812 , w_1813 , w_1814 , w_1815 , 
		w_1816 , w_1817 , w_1818 , w_1819 , w_1820 , w_1821 , w_1822 , w_1823 , w_1824 , w_1825 , 
		w_1826 , w_1827 , w_1828 , w_1829 , w_1830 , w_1831 , w_1832 , w_1833 , w_1834 , w_1835 , 
		w_1836 , w_1837 , w_1838 , w_1839 , w_1840 , w_1841 , w_1842 , w_1843 , w_1844 , w_1845 , 
		w_1846 , w_1847 , w_1848 , w_1849 , w_1850 , w_1851 , w_1852 , w_1853 , w_1854 , w_1855 , 
		w_1856 , w_1857 , w_1858 , w_1859 , w_1860 , w_1861 , w_1862 , w_1863 , w_1864 , w_1865 , 
		w_1866 , w_1867 , w_1868 , w_1869 , w_1870 , w_1871 , w_1872 , w_1873 , w_1874 , w_1875 , 
		w_1876 , w_1877 , w_1878 , w_1879 , w_1880 , w_1881 , w_1882 , w_1883 , w_1884 , w_1885 , 
		w_1886 , w_1887 , w_1888 , w_1889 , w_1890 , w_1891 , w_1892 , w_1893 , w_1894 , w_1895 , 
		w_1896 , w_1897 , w_1898 , w_1899 , w_1900 , w_1901 , w_1902 , w_1903 , w_1904 , w_1905 , 
		w_1906 , w_1907 , w_1908 , w_1909 , w_1910 , w_1911 , w_1912 , w_1913 , w_1914 , w_1915 , 
		w_1916 , w_1917 , w_1918 , w_1919 , w_1920 , w_1921 , w_1922 , w_1923 , w_1924 , w_1925 , 
		w_1926 , w_1927 , w_1928 , w_1929 , w_1930 , w_1931 , w_1932 , w_1933 , w_1934 , w_1935 , 
		w_1936 , w_1937 , w_1938 , w_1939 , w_1940 , w_1941 , w_1942 , w_1943 , w_1944 , w_1945 , 
		w_1946 , w_1947 , w_1948 , w_1949 , w_1950 , w_1951 , w_1952 , w_1953 , w_1954 , w_1955 , 
		w_1956 , w_1957 , w_1958 , w_1959 , w_1960 , w_1961 , w_1962 , w_1963 , w_1964 , w_1965 , 
		w_1966 , w_1967 , w_1968 , w_1969 , w_1970 , w_1971 , w_1972 , w_1973 , w_1974 , w_1975 , 
		w_1976 , w_1977 , w_1978 , w_1979 , w_1980 , w_1981 , w_1982 , w_1983 , w_1984 , w_1985 , 
		w_1986 , w_1987 , w_1988 , w_1989 , w_1990 , w_1991 , w_1992 , w_1993 , w_1994 , w_1995 , 
		w_1996 , w_1997 , w_1998 , w_1999 , w_2000 , w_2001 , w_2002 , w_2003 , w_2004 , w_2005 , 
		w_2006 , w_2007 , w_2008 , w_2009 , w_2010 , w_2011 , w_2012 , w_2013 , w_2014 , w_2015 , 
		w_2016 , w_2017 , w_2018 , w_2019 , w_2020 , w_2021 , w_2022 , w_2023 , w_2024 , w_2025 , 
		w_2026 , w_2027 , w_2028 , w_2029 , w_2030 , w_2031 , w_2032 , w_2033 , w_2034 , w_2035 , 
		w_2036 , w_2037 , w_2038 , w_2039 , w_2040 , w_2041 , w_2042 , w_2043 , w_2044 , w_2045 , 
		w_2046 , w_2047 , w_2048 , w_2049 , w_2050 , w_2051 , w_2052 , w_2053 , w_2054 , w_2055 , 
		w_2056 , w_2057 , w_2058 , w_2059 , w_2060 , w_2061 , w_2062 , w_2063 , w_2064 , w_2065 , 
		w_2066 , w_2067 , w_2068 , w_2069 , w_2070 , w_2071 , w_2072 , w_2073 , w_2074 , w_2075 , 
		w_2076 , w_2077 , w_2078 , w_2079 , w_2080 , w_2081 , w_2082 , w_2083 , w_2084 , w_2085 , 
		w_2086 , w_2087 , w_2088 , w_2089 , w_2090 , w_2091 , w_2092 , w_2093 , w_2094 , w_2095 , 
		w_2096 , w_2097 , w_2098 , w_2099 , w_2100 , w_2101 , w_2102 , w_2103 , w_2104 , w_2105 , 
		w_2106 , w_2107 , w_2108 , w_2109 , w_2110 , w_2111 , w_2112 , w_2113 , w_2114 , w_2115 , 
		w_2116 , w_2117 , w_2118 , w_2119 , w_2120 , w_2121 , w_2122 , w_2123 , w_2124 , w_2125 , 
		w_2126 , w_2127 , w_2128 , w_2129 , w_2130 , w_2131 , w_2132 , w_2133 , w_2134 , w_2135 , 
		w_2136 , w_2137 , w_2138 , w_2139 , w_2140 , w_2141 , w_2142 , w_2143 , w_2144 , w_2145 , 
		w_2146 , w_2147 , w_2148 , w_2149 , w_2150 , w_2151 , w_2152 , w_2153 , w_2154 , w_2155 , 
		w_2156 , w_2157 , w_2158 , w_2159 , w_2160 , w_2161 , w_2162 , w_2163 , w_2164 , w_2165 , 
		w_2166 , w_2167 , w_2168 , w_2169 , w_2170 , w_2171 , w_2172 , w_2173 , w_2174 , w_2175 , 
		w_2176 , w_2177 , w_2178 , w_2179 , w_2180 , w_2181 , w_2182 , w_2183 , w_2184 , w_2185 , 
		w_2186 , w_2187 , w_2188 , w_2189 , w_2190 , w_2191 , w_2192 , w_2193 , w_2194 , w_2195 , 
		w_2196 , w_2197 , w_2198 , w_2199 , w_2200 , w_2201 , w_2202 , w_2203 , w_2204 , w_2205 , 
		w_2206 , w_2207 , w_2208 , w_2209 , w_2210 , w_2211 , w_2212 , w_2213 , w_2214 , w_2215 , 
		w_2216 , w_2217 , w_2218 , w_2219 , w_2220 , w_2221 , w_2222 , w_2223 , w_2224 , w_2225 , 
		w_2226 , w_2227 , w_2228 , w_2229 , w_2230 , w_2231 , w_2232 , w_2233 , w_2234 , w_2235 , 
		w_2236 , w_2237 , w_2238 , w_2239 , w_2240 , w_2241 , w_2242 , w_2243 , w_2244 , w_2245 , 
		w_2246 , w_2247 , w_2248 , w_2249 , w_2250 , w_2251 , w_2252 , w_2253 , w_2254 , w_2255 , 
		w_2256 , w_2257 , w_2258 , w_2259 , w_2260 , w_2261 , w_2262 , w_2263 , w_2264 , w_2265 , 
		w_2266 , w_2267 , w_2268 , w_2269 , w_2270 , w_2271 , w_2272 , w_2273 , w_2274 , w_2275 , 
		w_2276 , w_2277 , w_2278 , w_2279 , w_2280 , w_2281 , w_2282 , w_2283 , w_2284 , w_2285 , 
		w_2286 , w_2287 , w_2288 , w_2289 , w_2290 , w_2291 , w_2292 , w_2293 , w_2294 , w_2295 , 
		w_2296 , w_2297 , w_2298 , w_2299 , w_2300 , w_2301 , w_2302 , w_2303 , w_2304 , w_2305 , 
		w_2306 , w_2307 , w_2308 , w_2309 , w_2310 , w_2311 , w_2312 , w_2313 , w_2314 , w_2315 , 
		w_2316 , w_2317 , w_2318 , w_2319 , w_2320 , w_2321 , w_2322 , w_2323 , w_2324 , w_2325 , 
		w_2326 , w_2327 , w_2328 , w_2329 , w_2330 , w_2331 , w_2332 , w_2333 , w_2334 , w_2335 , 
		w_2336 , w_2337 , w_2338 , w_2339 , w_2340 , w_2341 , w_2342 , w_2343 , w_2344 , w_2345 , 
		w_2346 , w_2347 , w_2348 , w_2349 , w_2350 , w_2351 , w_2352 , w_2353 , w_2354 , w_2355 , 
		w_2356 , w_2357 , w_2358 , w_2359 , w_2360 , w_2361 , w_2362 , w_2363 , w_2364 , w_2365 , 
		w_2366 , w_2367 , w_2368 , w_2369 , w_2370 , w_2371 , w_2372 , w_2373 , w_2374 , w_2375 , 
		w_2376 , w_2377 , w_2378 , w_2379 , w_2380 , w_2381 , w_2382 , w_2383 , w_2384 , w_2385 , 
		w_2386 , w_2387 , w_2388 , w_2389 , w_2390 , w_2391 , w_2392 , w_2393 , w_2394 , w_2395 , 
		w_2396 , w_2397 , w_2398 , w_2399 , w_2400 , w_2401 , w_2402 , w_2403 , w_2404 , w_2405 , 
		w_2406 , w_2407 , w_2408 , w_2409 , w_2410 , w_2411 , w_2412 , w_2413 , w_2414 , w_2415 , 
		w_2416 , w_2417 , w_2418 , w_2419 , w_2420 , w_2421 , w_2422 , w_2423 , w_2424 , w_2425 , 
		w_2426 , w_2427 , w_2428 , w_2429 , w_2430 , w_2431 , w_2432 , w_2433 , w_2434 , w_2435 , 
		w_2436 , w_2437 , w_2438 , w_2439 , w_2440 , w_2441 , w_2442 , w_2443 , w_2444 , w_2445 , 
		w_2446 , w_2447 , w_2448 , w_2449 , w_2450 , w_2451 , w_2452 , w_2453 , w_2454 , w_2455 , 
		w_2456 , w_2457 , w_2458 , w_2459 , w_2460 , w_2461 , w_2462 , w_2463 , w_2464 , w_2465 , 
		w_2466 , w_2467 , w_2468 , w_2469 , w_2470 , w_2471 , w_2472 , w_2473 , w_2474 , w_2475 , 
		w_2476 , w_2477 , w_2478 , w_2479 , w_2480 , w_2481 , w_2482 , w_2483 , w_2484 , w_2485 , 
		w_2486 , w_2487 , w_2488 , w_2489 , w_2490 , w_2491 , w_2492 , w_2493 , w_2494 , w_2495 , 
		w_2496 , w_2497 , w_2498 , w_2499 , w_2500 , w_2501 , w_2502 , w_2503 , w_2504 , w_2505 , 
		w_2506 , w_2507 , w_2508 , w_2509 , w_2510 , w_2511 , w_2512 , w_2513 , w_2514 , w_2515 , 
		w_2516 , w_2517 , w_2518 , w_2519 , w_2520 , w_2521 , w_2522 , w_2523 , w_2524 , w_2525 , 
		w_2526 , w_2527 , w_2528 , w_2529 , w_2530 , w_2531 , w_2532 , w_2533 , w_2534 , w_2535 , 
		w_2536 , w_2537 , w_2538 , w_2539 , w_2540 , w_2541 , w_2542 , w_2543 , w_2544 , w_2545 , 
		w_2546 , w_2547 , w_2548 , w_2549 , w_2550 , w_2551 , w_2552 , w_2553 , w_2554 , w_2555 , 
		w_2556 , w_2557 , w_2558 , w_2559 , w_2560 , w_2561 , w_2562 , w_2563 , w_2564 , w_2565 , 
		w_2566 , w_2567 , w_2568 , w_2569 , w_2570 , w_2571 , w_2572 , w_2573 , w_2574 , w_2575 , 
		w_2576 , w_2577 , w_2578 , w_2579 , w_2580 , w_2581 , w_2582 , w_2583 , w_2584 , w_2585 , 
		w_2586 , w_2587 , w_2588 , w_2589 , w_2590 , w_2591 , w_2592 , w_2593 , w_2594 , w_2595 , 
		w_2596 , w_2597 , w_2598 , w_2599 , w_2600 , w_2601 , w_2602 , w_2603 , w_2604 , w_2605 , 
		w_2606 , w_2607 , w_2608 , w_2609 , w_2610 , w_2611 , w_2612 , w_2613 , w_2614 , w_2615 , 
		w_2616 , w_2617 , w_2618 , w_2619 , w_2620 , w_2621 , w_2622 , w_2623 , w_2624 , w_2625 , 
		w_2626 , w_2627 , w_2628 , w_2629 , w_2630 , w_2631 , w_2632 , w_2633 , w_2634 , w_2635 , 
		w_2636 , w_2637 , w_2638 , w_2639 , w_2640 , w_2641 , w_2642 , w_2643 , w_2644 , w_2645 , 
		w_2646 , w_2647 , w_2648 , w_2649 , w_2650 , w_2651 , w_2652 , w_2653 , w_2654 , w_2655 , 
		w_2656 , w_2657 , w_2658 , w_2659 , w_2660 , w_2661 , w_2662 , w_2663 , w_2664 , w_2665 , 
		w_2666 , w_2667 , w_2668 , w_2669 , w_2670 , w_2671 , w_2672 , w_2673 , w_2674 , w_2675 , 
		w_2676 , w_2677 , w_2678 , w_2679 , w_2680 , w_2681 , w_2682 , w_2683 , w_2684 , w_2685 , 
		w_2686 , w_2687 , w_2688 , w_2689 , w_2690 , w_2691 , w_2692 , w_2693 , w_2694 , w_2695 , 
		w_2696 , w_2697 , w_2698 , w_2699 , w_2700 , w_2701 , w_2702 , w_2703 , w_2704 , w_2705 , 
		w_2706 , w_2707 , w_2708 , w_2709 , w_2710 , w_2711 , w_2712 , w_2713 , w_2714 , w_2715 , 
		w_2716 , w_2717 , w_2718 , w_2719 , w_2720 , w_2721 , w_2722 , w_2723 , w_2724 , w_2725 , 
		w_2726 , w_2727 , w_2728 , w_2729 , w_2730 , w_2731 , w_2732 , w_2733 , w_2734 , w_2735 , 
		w_2736 , w_2737 , w_2738 , w_2739 , w_2740 , w_2741 , w_2742 , w_2743 , w_2744 , w_2745 , 
		w_2746 , w_2747 , w_2748 , w_2749 , w_2750 , w_2751 , w_2752 , w_2753 , w_2754 , w_2755 , 
		w_2756 , w_2757 , w_2758 , w_2759 , w_2760 , w_2761 , w_2762 , w_2763 , w_2764 , w_2765 , 
		w_2766 , w_2767 , w_2768 , w_2769 , w_2770 , w_2771 , w_2772 , w_2773 , w_2774 , w_2775 , 
		w_2776 , w_2777 , w_2778 , w_2779 , w_2780 , w_2781 , w_2782 , w_2783 , w_2784 , w_2785 , 
		w_2786 , w_2787 , w_2788 , w_2789 , w_2790 , w_2791 , w_2792 , w_2793 , w_2794 , w_2795 , 
		w_2796 , w_2797 , w_2798 , w_2799 , w_2800 , w_2801 , w_2802 , w_2803 , w_2804 , w_2805 , 
		w_2806 , w_2807 , w_2808 , w_2809 , w_2810 , w_2811 , w_2812 , w_2813 , w_2814 , w_2815 , 
		w_2816 , w_2817 , w_2818 , w_2819 , w_2820 , w_2821 , w_2822 , w_2823 , w_2824 , w_2825 , 
		w_2826 , w_2827 , w_2828 , w_2829 , w_2830 , w_2831 , w_2832 , w_2833 , w_2834 , w_2835 , 
		w_2836 , w_2837 , w_2838 , w_2839 , w_2840 , w_2841 , w_2842 , w_2843 , w_2844 , w_2845 , 
		w_2846 , w_2847 , w_2848 , w_2849 , w_2850 , w_2851 , w_2852 , w_2853 , w_2854 , w_2855 , 
		w_2856 , w_2857 , w_2858 , w_2859 , w_2860 , w_2861 , w_2862 , w_2863 , w_2864 , w_2865 , 
		w_2866 , w_2867 , w_2868 , w_2869 , w_2870 , w_2871 , w_2872 , w_2873 , w_2874 , w_2875 , 
		w_2876 , w_2877 , w_2878 , w_2879 , w_2880 , w_2881 , w_2882 , w_2883 , w_2884 , w_2885 , 
		w_2886 , w_2887 , w_2888 , w_2889 , w_2890 , w_2891 , w_2892 , w_2893 , w_2894 , w_2895 , 
		w_2896 , w_2897 , w_2898 , w_2899 , w_2900 , w_2901 , w_2902 , w_2903 , w_2904 , w_2905 , 
		w_2906 , w_2907 , w_2908 , w_2909 , w_2910 , w_2911 , w_2912 , w_2913 , w_2914 , w_2915 , 
		w_2916 , w_2917 , w_2918 , w_2919 , w_2920 , w_2921 , w_2922 , w_2923 , w_2924 , w_2925 , 
		w_2926 , w_2927 , w_2928 , w_2929 , w_2930 , w_2931 , w_2932 , w_2933 , w_2934 , w_2935 , 
		w_2936 , w_2937 , w_2938 , w_2939 , w_2940 , w_2941 , w_2942 , w_2943 , w_2944 , w_2945 , 
		w_2946 , w_2947 , w_2948 , w_2949 , w_2950 , w_2951 , w_2952 , w_2953 , w_2954 , w_2955 , 
		w_2956 , w_2957 , w_2958 , w_2959 , w_2960 , w_2961 , w_2962 , w_2963 , w_2964 , w_2965 , 
		w_2966 , w_2967 , w_2968 , w_2969 , w_2970 , w_2971 , w_2972 , w_2973 , w_2974 , w_2975 , 
		w_2976 , w_2977 , w_2978 , w_2979 , w_2980 , w_2981 , w_2982 , w_2983 , w_2984 , w_2985 , 
		w_2986 , w_2987 , w_2988 , w_2989 , w_2990 , w_2991 , w_2992 , w_2993 , w_2994 , w_2995 , 
		w_2996 , w_2997 , w_2998 , w_2999 , w_3000 , w_3001 , w_3002 , w_3003 , w_3004 , w_3005 , 
		w_3006 , w_3007 , w_3008 , w_3009 , w_3010 , w_3011 , w_3012 , w_3013 , w_3014 , w_3015 , 
		w_3016 , w_3017 , w_3018 , w_3019 , w_3020 , w_3021 , w_3022 , w_3023 , w_3024 , w_3025 , 
		w_3026 , w_3027 , w_3028 , w_3029 , w_3030 , w_3031 , w_3032 , w_3033 , w_3034 , w_3035 , 
		w_3036 , w_3037 , w_3038 , w_3039 , w_3040 , w_3041 , w_3042 , w_3043 , w_3044 , w_3045 , 
		w_3046 , w_3047 , w_3048 , w_3049 , w_3050 , w_3051 , w_3052 , w_3053 , w_3054 , w_3055 , 
		w_3056 , w_3057 , w_3058 , w_3059 , w_3060 , w_3061 , w_3062 , w_3063 , w_3064 , w_3065 , 
		w_3066 , w_3067 , w_3068 , w_3069 , w_3070 , w_3071 , w_3072 , w_3073 , w_3074 , w_3075 , 
		w_3076 , w_3077 , w_3078 , w_3079 , w_3080 , w_3081 , w_3082 , w_3083 , w_3084 , w_3085 , 
		w_3086 , w_3087 , w_3088 , w_3089 , w_3090 , w_3091 , w_3092 , w_3093 , w_3094 , w_3095 , 
		w_3096 , w_3097 , w_3098 , w_3099 , w_3100 , w_3101 , w_3102 , w_3103 , w_3104 , w_3105 , 
		w_3106 , w_3107 , w_3108 , w_3109 , w_3110 , w_3111 , w_3112 , w_3113 , w_3114 , w_3115 , 
		w_3116 , w_3117 , w_3118 , w_3119 , w_3120 , w_3121 , w_3122 , w_3123 , w_3124 , w_3125 , 
		w_3126 , w_3127 , w_3128 , w_3129 , w_3130 , w_3131 , w_3132 , w_3133 , w_3134 , w_3135 , 
		w_3136 , w_3137 , w_3138 , w_3139 , w_3140 , w_3141 , w_3142 , w_3143 , w_3144 , w_3145 , 
		w_3146 , w_3147 , w_3148 , w_3149 , w_3150 , w_3151 , w_3152 , w_3153 , w_3154 , w_3155 , 
		w_3156 , w_3157 , w_3158 , w_3159 , w_3160 , w_3161 , w_3162 , w_3163 , w_3164 , w_3165 , 
		w_3166 , w_3167 , w_3168 , w_3169 , w_3170 , w_3171 , w_3172 , w_3173 , w_3174 , w_3175 , 
		w_3176 , w_3177 , w_3178 , w_3179 , w_3180 , w_3181 , w_3182 , w_3183 , w_3184 , w_3185 , 
		w_3186 , w_3187 , w_3188 , w_3189 , w_3190 , w_3191 , w_3192 , w_3193 , w_3194 , w_3195 , 
		w_3196 , w_3197 , w_3198 , w_3199 , w_3200 , w_3201 , w_3202 , w_3203 , w_3204 , w_3205 , 
		w_3206 , w_3207 , w_3208 , w_3209 , w_3210 , w_3211 , w_3212 , w_3213 , w_3214 , w_3215 , 
		w_3216 , w_3217 , w_3218 , w_3219 , w_3220 , w_3221 , w_3222 , w_3223 , w_3224 , w_3225 , 
		w_3226 , w_3227 , w_3228 , w_3229 , w_3230 , w_3231 , w_3232 , w_3233 , w_3234 , w_3235 , 
		w_3236 , w_3237 , w_3238 , w_3239 , w_3240 , w_3241 , w_3242 , w_3243 , w_3244 , w_3245 , 
		w_3246 , w_3247 , w_3248 , w_3249 , w_3250 , w_3251 , w_3252 , w_3253 , w_3254 , w_3255 , 
		w_3256 , w_3257 , w_3258 , w_3259 , w_3260 , w_3261 , w_3262 , w_3263 , w_3264 , w_3265 , 
		w_3266 , w_3267 , w_3268 , w_3269 , w_3270 , w_3271 , w_3272 , w_3273 , w_3274 , w_3275 , 
		w_3276 , w_3277 , w_3278 , w_3279 , w_3280 , w_3281 , w_3282 , w_3283 , w_3284 , w_3285 , 
		w_3286 , w_3287 , w_3288 , w_3289 , w_3290 , w_3291 , w_3292 , w_3293 , w_3294 , w_3295 , 
		w_3296 , w_3297 , w_3298 , w_3299 , w_3300 , w_3301 , w_3302 , w_3303 , w_3304 , w_3305 , 
		w_3306 , w_3307 , w_3308 , w_3309 , w_3310 , w_3311 , w_3312 , w_3313 , w_3314 , w_3315 , 
		w_3316 , w_3317 , w_3318 , w_3319 , w_3320 , w_3321 , w_3322 , w_3323 , w_3324 , w_3325 , 
		w_3326 , w_3327 , w_3328 , w_3329 , w_3330 , w_3331 , w_3332 , w_3333 , w_3334 , w_3335 , 
		w_3336 , w_3337 , w_3338 , w_3339 , w_3340 , w_3341 , w_3342 , w_3343 , w_3344 , w_3345 , 
		w_3346 , w_3347 , w_3348 , w_3349 , w_3350 , w_3351 , w_3352 , w_3353 , w_3354 , w_3355 , 
		w_3356 , w_3357 , w_3358 , w_3359 , w_3360 , w_3361 , w_3362 , w_3363 , w_3364 , w_3365 , 
		w_3366 , w_3367 , w_3368 , w_3369 , w_3370 , w_3371 , w_3372 , w_3373 , w_3374 , w_3375 , 
		w_3376 , w_3377 , w_3378 , w_3379 , w_3380 , w_3381 , w_3382 , w_3383 , w_3384 , w_3385 , 
		w_3386 , w_3387 , w_3388 , w_3389 , w_3390 , w_3391 , w_3392 , w_3393 , w_3394 , w_3395 , 
		w_3396 , w_3397 , w_3398 , w_3399 , w_3400 , w_3401 , w_3402 , w_3403 , w_3404 , w_3405 , 
		w_3406 , w_3407 , w_3408 , w_3409 , w_3410 , w_3411 , w_3412 , w_3413 , w_3414 , w_3415 , 
		w_3416 , w_3417 , w_3418 , w_3419 , w_3420 , w_3421 , w_3422 , w_3423 , w_3424 , w_3425 , 
		w_3426 , w_3427 , w_3428 , w_3429 , w_3430 , w_3431 , w_3432 , w_3433 , w_3434 , w_3435 , 
		w_3436 , w_3437 , w_3438 , w_3439 , w_3440 , w_3441 , w_3442 , w_3443 , w_3444 , w_3445 , 
		w_3446 , w_3447 , w_3448 , w_3449 , w_3450 , w_3451 , w_3452 , w_3453 , w_3454 , w_3455 , 
		w_3456 , w_3457 , w_3458 , w_3459 , w_3460 , w_3461 , w_3462 , w_3463 , w_3464 , w_3465 , 
		w_3466 , w_3467 , w_3468 , w_3469 , w_3470 , w_3471 , w_3472 , w_3473 , w_3474 , w_3475 , 
		w_3476 , w_3477 , w_3478 , w_3479 , w_3480 , w_3481 , w_3482 , w_3483 , w_3484 , w_3485 , 
		w_3486 , w_3487 , w_3488 , w_3489 , w_3490 , w_3491 , w_3492 , w_3493 , w_3494 , w_3495 , 
		w_3496 , w_3497 , w_3498 , w_3499 , w_3500 , w_3501 , w_3502 , w_3503 , w_3504 , w_3505 , 
		w_3506 , w_3507 , w_3508 , w_3509 , w_3510 , w_3511 , w_3512 , w_3513 , w_3514 , w_3515 , 
		w_3516 , w_3517 , w_3518 , w_3519 , w_3520 , w_3521 , w_3522 , w_3523 , w_3524 , w_3525 , 
		w_3526 , w_3527 , w_3528 , w_3529 , w_3530 , w_3531 , w_3532 , w_3533 , w_3534 , w_3535 , 
		w_3536 , w_3537 , w_3538 , w_3539 , w_3540 , w_3541 , w_3542 , w_3543 , w_3544 , w_3545 , 
		w_3546 , w_3547 , w_3548 , w_3549 , w_3550 , w_3551 , w_3552 , w_3553 , w_3554 , w_3555 , 
		w_3556 , w_3557 , w_3558 , w_3559 , w_3560 , w_3561 , w_3562 , w_3563 , w_3564 , w_3565 , 
		w_3566 , w_3567 , w_3568 , w_3569 , w_3570 , w_3571 , w_3572 , w_3573 , w_3574 , w_3575 , 
		w_3576 , w_3577 , w_3578 , w_3579 , w_3580 , w_3581 , w_3582 , w_3583 , w_3584 , w_3585 , 
		w_3586 , w_3587 , w_3588 , w_3589 , w_3590 , w_3591 , w_3592 , w_3593 , w_3594 , w_3595 , 
		w_3596 , w_3597 , w_3598 , w_3599 , w_3600 , w_3601 , w_3602 , w_3603 , w_3604 , w_3605 , 
		w_3606 , w_3607 , w_3608 , w_3609 , w_3610 , w_3611 , w_3612 , w_3613 , w_3614 , w_3615 , 
		w_3616 , w_3617 , w_3618 , w_3619 , w_3620 , w_3621 , w_3622 , w_3623 , w_3624 , w_3625 , 
		w_3626 , w_3627 , w_3628 , w_3629 , w_3630 , w_3631 , w_3632 , w_3633 , w_3634 , w_3635 , 
		w_3636 , w_3637 , w_3638 , w_3639 , w_3640 , w_3641 , w_3642 , w_3643 , w_3644 , w_3645 , 
		w_3646 , w_3647 , w_3648 , w_3649 , w_3650 , w_3651 , w_3652 , w_3653 , w_3654 , w_3655 , 
		w_3656 , w_3657 , w_3658 , w_3659 , w_3660 , w_3661 , w_3662 , w_3663 , w_3664 , w_3665 , 
		w_3666 , w_3667 , w_3668 , w_3669 , w_3670 , w_3671 , w_3672 , w_3673 , w_3674 , w_3675 , 
		w_3676 , w_3677 , w_3678 , w_3679 , w_3680 , w_3681 , w_3682 , w_3683 , w_3684 , w_3685 , 
		w_3686 , w_3687 , w_3688 , w_3689 , w_3690 , w_3691 , w_3692 , w_3693 , w_3694 , w_3695 , 
		w_3696 , w_3697 , w_3698 , w_3699 , w_3700 , w_3701 , w_3702 , w_3703 , w_3704 , w_3705 , 
		w_3706 , w_3707 , w_3708 , w_3709 , w_3710 , w_3711 , w_3712 , w_3713 , w_3714 , w_3715 , 
		w_3716 , w_3717 , w_3718 , w_3719 , w_3720 , w_3721 , w_3722 , w_3723 , w_3724 , w_3725 , 
		w_3726 , w_3727 , w_3728 , w_3729 , w_3730 , w_3731 , w_3732 , w_3733 , w_3734 , w_3735 , 
		w_3736 , w_3737 , w_3738 , w_3739 , w_3740 , w_3741 , w_3742 , w_3743 , w_3744 , w_3745 , 
		w_3746 , w_3747 , w_3748 , w_3749 , w_3750 , w_3751 , w_3752 , w_3753 , w_3754 , w_3755 , 
		w_3756 , w_3757 , w_3758 , w_3759 , w_3760 , w_3761 , w_3762 , w_3763 , w_3764 , w_3765 , 
		w_3766 , w_3767 , w_3768 , w_3769 , w_3770 , w_3771 , w_3772 , w_3773 , w_3774 , w_3775 , 
		w_3776 , w_3777 , w_3778 , w_3779 , w_3780 , w_3781 , w_3782 , w_3783 , w_3784 , w_3785 , 
		w_3786 , w_3787 , w_3788 , w_3789 , w_3790 , w_3791 , w_3792 , w_3793 , w_3794 , w_3795 , 
		w_3796 , w_3797 , w_3798 , w_3799 , w_3800 , w_3801 , w_3802 , w_3803 , w_3804 , w_3805 , 
		w_3806 , w_3807 , w_3808 , w_3809 , w_3810 , w_3811 , w_3812 , w_3813 , w_3814 , w_3815 , 
		w_3816 , w_3817 , w_3818 , w_3819 , w_3820 , w_3821 , w_3822 , w_3823 , w_3824 , w_3825 , 
		w_3826 , w_3827 , w_3828 , w_3829 , w_3830 , w_3831 , w_3832 , w_3833 , w_3834 , w_3835 , 
		w_3836 , w_3837 , w_3838 , w_3839 , w_3840 , w_3841 , w_3842 , w_3843 , w_3844 , w_3845 , 
		w_3846 , w_3847 , w_3848 , w_3849 , w_3850 , w_3851 , w_3852 , w_3853 , w_3854 , w_3855 , 
		w_3856 , w_3857 , w_3858 , w_3859 , w_3860 , w_3861 , w_3862 , w_3863 , w_3864 , w_3865 , 
		w_3866 , w_3867 , w_3868 , w_3869 , w_3870 , w_3871 , w_3872 , w_3873 , w_3874 , w_3875 , 
		w_3876 , w_3877 , w_3878 , w_3879 , w_3880 , w_3881 , w_3882 , w_3883 , w_3884 , w_3885 , 
		w_3886 , w_3887 , w_3888 , w_3889 , w_3890 , w_3891 , w_3892 , w_3893 , w_3894 , w_3895 , 
		w_3896 , w_3897 , w_3898 , w_3899 , w_3900 , w_3901 , w_3902 , w_3903 , w_3904 , w_3905 , 
		w_3906 , w_3907 , w_3908 , w_3909 , w_3910 , w_3911 , w_3912 , w_3913 , w_3914 , w_3915 , 
		w_3916 , w_3917 , w_3918 , w_3919 , w_3920 , w_3921 , w_3922 , w_3923 , w_3924 , w_3925 , 
		w_3926 , w_3927 , w_3928 , w_3929 , w_3930 , w_3931 , w_3932 , w_3933 , w_3934 , w_3935 , 
		w_3936 , w_3937 , w_3938 , w_3939 , w_3940 , w_3941 , w_3942 , w_3943 , w_3944 , w_3945 , 
		w_3946 , w_3947 , w_3948 , w_3949 , w_3950 , w_3951 , w_3952 , w_3953 , w_3954 , w_3955 , 
		w_3956 , w_3957 , w_3958 , w_3959 , w_3960 , w_3961 , w_3962 , w_3963 , w_3964 , w_3965 , 
		w_3966 , w_3967 , w_3968 , w_3969 , w_3970 , w_3971 , w_3972 , w_3973 , w_3974 , w_3975 , 
		w_3976 , w_3977 , w_3978 , w_3979 , w_3980 , w_3981 , w_3982 , w_3983 , w_3984 , w_3985 , 
		w_3986 , w_3987 , w_3988 , w_3989 , w_3990 , w_3991 , w_3992 , w_3993 , w_3994 , w_3995 , 
		w_3996 , w_3997 , w_3998 , w_3999 , w_4000 , w_4001 , w_4002 , w_4003 , w_4004 , w_4005 , 
		w_4006 , w_4007 , w_4008 , w_4009 , w_4010 , w_4011 , w_4012 , w_4013 , w_4014 , w_4015 , 
		w_4016 , w_4017 , w_4018 , w_4019 , w_4020 , w_4021 , w_4022 , w_4023 , w_4024 , w_4025 , 
		w_4026 , w_4027 , w_4028 , w_4029 , w_4030 , w_4031 , w_4032 , w_4033 , w_4034 , w_4035 , 
		w_4036 , w_4037 , w_4038 , w_4039 , w_4040 , w_4041 , w_4042 , w_4043 , w_4044 , w_4045 , 
		w_4046 , w_4047 , w_4048 , w_4049 , w_4050 , w_4051 , w_4052 , w_4053 , w_4054 , w_4055 , 
		w_4056 , w_4057 , w_4058 , w_4059 , w_4060 , w_4061 , w_4062 , w_4063 , w_4064 , w_4065 , 
		w_4066 , w_4067 , w_4068 , w_4069 , w_4070 , w_4071 , w_4072 , w_4073 , w_4074 , w_4075 , 
		w_4076 , w_4077 , w_4078 , w_4079 , w_4080 , w_4081 , w_4082 , w_4083 , w_4084 , w_4085 , 
		w_4086 , w_4087 , w_4088 , w_4089 , w_4090 , w_4091 , w_4092 , w_4093 , w_4094 , w_4095 , 
		w_4096 , w_4097 , w_4098 , w_4099 , w_4100 , w_4101 , w_4102 , w_4103 , w_4104 , w_4105 , 
		w_4106 , w_4107 , w_4108 , w_4109 , w_4110 , w_4111 , w_4112 , w_4113 , w_4114 , w_4115 , 
		w_4116 , w_4117 , w_4118 , w_4119 , w_4120 , w_4121 , w_4122 , w_4123 , w_4124 , w_4125 , 
		w_4126 , w_4127 , w_4128 , w_4129 , w_4130 , w_4131 , w_4132 , w_4133 , w_4134 , w_4135 , 
		w_4136 , w_4137 , w_4138 , w_4139 , w_4140 , w_4141 , w_4142 , w_4143 , w_4144 , w_4145 , 
		w_4146 , w_4147 , w_4148 , w_4149 , w_4150 , w_4151 , w_4152 , w_4153 , w_4154 , w_4155 , 
		w_4156 , w_4157 , w_4158 , w_4159 , w_4160 , w_4161 , w_4162 , w_4163 , w_4164 , w_4165 , 
		w_4166 , w_4167 , w_4168 , w_4169 , w_4170 , w_4171 , w_4172 , w_4173 , w_4174 , w_4175 , 
		w_4176 , w_4177 , w_4178 , w_4179 , w_4180 , w_4181 , w_4182 , w_4183 , w_4184 , w_4185 , 
		w_4186 , w_4187 , w_4188 , w_4189 , w_4190 , w_4191 , w_4192 , w_4193 , w_4194 , w_4195 , 
		w_4196 , w_4197 , w_4198 , w_4199 , w_4200 , w_4201 , w_4202 , w_4203 , w_4204 , w_4205 , 
		w_4206 , w_4207 , w_4208 , w_4209 , w_4210 , w_4211 , w_4212 , w_4213 , w_4214 , w_4215 , 
		w_4216 , w_4217 , w_4218 , w_4219 , w_4220 , w_4221 , w_4222 , w_4223 , w_4224 , w_4225 , 
		w_4226 , w_4227 , w_4228 , w_4229 , w_4230 , w_4231 , w_4232 , w_4233 , w_4234 , w_4235 , 
		w_4236 , w_4237 , w_4238 , w_4239 , w_4240 , w_4241 , w_4242 , w_4243 , w_4244 , w_4245 , 
		w_4246 , w_4247 , w_4248 , w_4249 , w_4250 , w_4251 , w_4252 , w_4253 , w_4254 , w_4255 , 
		w_4256 , w_4257 , w_4258 , w_4259 , w_4260 , w_4261 , w_4262 , w_4263 , w_4264 , w_4265 , 
		w_4266 , w_4267 , w_4268 , w_4269 , w_4270 , w_4271 , w_4272 , w_4273 , w_4274 , w_4275 , 
		w_4276 , w_4277 , w_4278 , w_4279 , w_4280 , w_4281 , w_4282 , w_4283 , w_4284 , w_4285 , 
		w_4286 , w_4287 , w_4288 , w_4289 , w_4290 , w_4291 , w_4292 , w_4293 , w_4294 , w_4295 , 
		w_4296 , w_4297 , w_4298 , w_4299 , w_4300 , w_4301 , w_4302 , w_4303 , w_4304 , w_4305 , 
		w_4306 , w_4307 , w_4308 , w_4309 , w_4310 , w_4311 , w_4312 , w_4313 , w_4314 , w_4315 , 
		w_4316 , w_4317 , w_4318 , w_4319 , w_4320 , w_4321 , w_4322 , w_4323 , w_4324 , w_4325 , 
		w_4326 , w_4327 , w_4328 , w_4329 , w_4330 , w_4331 , w_4332 , w_4333 , w_4334 , w_4335 , 
		w_4336 , w_4337 , w_4338 , w_4339 , w_4340 , w_4341 , w_4342 , w_4343 , w_4344 , w_4345 , 
		w_4346 , w_4347 , w_4348 , w_4349 , w_4350 , w_4351 , w_4352 , w_4353 , w_4354 , w_4355 , 
		w_4356 , w_4357 , w_4358 , w_4359 , w_4360 , w_4361 , w_4362 , w_4363 , w_4364 , w_4365 , 
		w_4366 , w_4367 , w_4368 , w_4369 , w_4370 , w_4371 , w_4372 , w_4373 , w_4374 , w_4375 , 
		w_4376 , w_4377 , w_4378 , w_4379 , w_4380 , w_4381 , w_4382 , w_4383 , w_4384 , w_4385 , 
		w_4386 , w_4387 , w_4388 , w_4389 , w_4390 , w_4391 , w_4392 , w_4393 , w_4394 , w_4395 , 
		w_4396 , w_4397 , w_4398 , w_4399 , w_4400 , w_4401 , w_4402 , w_4403 , w_4404 , w_4405 , 
		w_4406 , w_4407 , w_4408 , w_4409 , w_4410 , w_4411 , w_4412 , w_4413 , w_4414 , w_4415 , 
		w_4416 , w_4417 , w_4418 , w_4419 , w_4420 , w_4421 , w_4422 , w_4423 , w_4424 , w_4425 , 
		w_4426 , w_4427 , w_4428 , w_4429 , w_4430 , w_4431 , w_4432 , w_4433 , w_4434 , w_4435 , 
		w_4436 , w_4437 , w_4438 , w_4439 , w_4440 , w_4441 , w_4442 , w_4443 , w_4444 , w_4445 , 
		w_4446 , w_4447 , w_4448 , w_4449 , w_4450 , w_4451 , w_4452 , w_4453 , w_4454 , w_4455 , 
		w_4456 , w_4457 , w_4458 , w_4459 , w_4460 , w_4461 , w_4462 , w_4463 , w_4464 , w_4465 , 
		w_4466 , w_4467 , w_4468 , w_4469 , w_4470 , w_4471 , w_4472 , w_4473 , w_4474 , w_4475 , 
		w_4476 , w_4477 , w_4478 , w_4479 , w_4480 , w_4481 , w_4482 , w_4483 , w_4484 , w_4485 , 
		w_4486 , w_4487 , w_4488 , w_4489 , w_4490 , w_4491 , w_4492 , w_4493 , w_4494 , w_4495 , 
		w_4496 , w_4497 , w_4498 , w_4499 , w_4500 , w_4501 , w_4502 , w_4503 , w_4504 , w_4505 , 
		w_4506 , w_4507 , w_4508 , w_4509 , w_4510 , w_4511 , w_4512 , w_4513 , w_4514 , w_4515 , 
		w_4516 , w_4517 , w_4518 , w_4519 , w_4520 , w_4521 , w_4522 , w_4523 , w_4524 , w_4525 , 
		w_4526 , w_4527 , w_4528 , w_4529 , w_4530 , w_4531 , w_4532 , w_4533 , w_4534 , w_4535 , 
		w_4536 , w_4537 , w_4538 , w_4539 , w_4540 , w_4541 , w_4542 , w_4543 , w_4544 , w_4545 , 
		w_4546 , w_4547 , w_4548 , w_4549 , w_4550 , w_4551 , w_4552 , w_4553 , w_4554 , w_4555 , 
		w_4556 , w_4557 , w_4558 , w_4559 , w_4560 , w_4561 , w_4562 , w_4563 , w_4564 , w_4565 , 
		w_4566 , w_4567 , w_4568 , w_4569 , w_4570 , w_4571 , w_4572 , w_4573 , w_4574 , w_4575 , 
		w_4576 , w_4577 , w_4578 , w_4579 , w_4580 , w_4581 , w_4582 , w_4583 , w_4584 , w_4585 , 
		w_4586 , w_4587 , w_4588 , w_4589 , w_4590 , w_4591 , w_4592 , w_4593 , w_4594 , w_4595 , 
		w_4596 , w_4597 , w_4598 , w_4599 , w_4600 , w_4601 , w_4602 , w_4603 , w_4604 , w_4605 , 
		w_4606 , w_4607 , w_4608 , w_4609 , w_4610 , w_4611 , w_4612 , w_4613 , w_4614 , w_4615 , 
		w_4616 , w_4617 , w_4618 , w_4619 , w_4620 , w_4621 , w_4622 , w_4623 , w_4624 , w_4625 , 
		w_4626 , w_4627 , w_4628 , w_4629 , w_4630 , w_4631 , w_4632 , w_4633 , w_4634 , w_4635 , 
		w_4636 , w_4637 , w_4638 , w_4639 , w_4640 , w_4641 , w_4642 , w_4643 , w_4644 , w_4645 , 
		w_4646 , w_4647 , w_4648 , w_4649 , w_4650 , w_4651 , w_4652 , w_4653 , w_4654 , w_4655 , 
		w_4656 , w_4657 , w_4658 , w_4659 , w_4660 , w_4661 , w_4662 , w_4663 , w_4664 , w_4665 , 
		w_4666 , w_4667 , w_4668 , w_4669 , w_4670 , w_4671 , w_4672 , w_4673 , w_4674 , w_4675 , 
		w_4676 , w_4677 , w_4678 , w_4679 , w_4680 , w_4681 , w_4682 , w_4683 , w_4684 , w_4685 , 
		w_4686 , w_4687 , w_4688 , w_4689 , w_4690 , w_4691 , w_4692 , w_4693 , w_4694 , w_4695 , 
		w_4696 , w_4697 , w_4698 , w_4699 , w_4700 , w_4701 , w_4702 , w_4703 , w_4704 , w_4705 , 
		w_4706 , w_4707 , w_4708 , w_4709 , w_4710 , w_4711 , w_4712 , w_4713 , w_4714 , w_4715 , 
		w_4716 , w_4717 , w_4718 , w_4719 , w_4720 , w_4721 , w_4722 , w_4723 , w_4724 , w_4725 , 
		w_4726 , w_4727 , w_4728 , w_4729 , w_4730 , w_4731 , w_4732 , w_4733 , w_4734 , w_4735 , 
		w_4736 , w_4737 , w_4738 , w_4739 , w_4740 , w_4741 , w_4742 , w_4743 , w_4744 , w_4745 , 
		w_4746 , w_4747 , w_4748 , w_4749 , w_4750 , w_4751 , w_4752 , w_4753 , w_4754 , w_4755 , 
		w_4756 , w_4757 , w_4758 , w_4759 , w_4760 , w_4761 , w_4762 , w_4763 , w_4764 , w_4765 , 
		w_4766 , w_4767 , w_4768 , w_4769 , w_4770 , w_4771 , w_4772 , w_4773 , w_4774 , w_4775 , 
		w_4776 , w_4777 , w_4778 , w_4779 , w_4780 , w_4781 , w_4782 , w_4783 , w_4784 , w_4785 , 
		w_4786 , w_4787 , w_4788 , w_4789 , w_4790 , w_4791 , w_4792 , w_4793 , w_4794 , w_4795 , 
		w_4796 , w_4797 , w_4798 , w_4799 , w_4800 , w_4801 , w_4802 , w_4803 , w_4804 , w_4805 , 
		w_4806 , w_4807 , w_4808 , w_4809 , w_4810 , w_4811 , w_4812 , w_4813 , w_4814 , w_4815 , 
		w_4816 , w_4817 , w_4818 , w_4819 , w_4820 , w_4821 , w_4822 , w_4823 , w_4824 , w_4825 , 
		w_4826 , w_4827 , w_4828 , w_4829 , w_4830 , w_4831 , w_4832 , w_4833 , w_4834 , w_4835 , 
		w_4836 , w_4837 , w_4838 , w_4839 , w_4840 , w_4841 , w_4842 , w_4843 , w_4844 , w_4845 , 
		w_4846 , w_4847 , w_4848 , w_4849 , w_4850 , w_4851 , w_4852 , w_4853 , w_4854 , w_4855 , 
		w_4856 , w_4857 , w_4858 , w_4859 , w_4860 , w_4861 , w_4862 , w_4863 , w_4864 , w_4865 , 
		w_4866 , w_4867 , w_4868 , w_4869 , w_4870 , w_4871 , w_4872 , w_4873 , w_4874 , w_4875 , 
		w_4876 , w_4877 , w_4878 , w_4879 , w_4880 , w_4881 , w_4882 , w_4883 , w_4884 , w_4885 , 
		w_4886 , w_4887 , w_4888 , w_4889 , w_4890 , w_4891 , w_4892 , w_4893 , w_4894 , w_4895 , 
		w_4896 , w_4897 , w_4898 , w_4899 , w_4900 , w_4901 , w_4902 , w_4903 , w_4904 , w_4905 , 
		w_4906 , w_4907 , w_4908 , w_4909 , w_4910 , w_4911 , w_4912 , w_4913 , w_4914 , w_4915 , 
		w_4916 , w_4917 , w_4918 , w_4919 , w_4920 , w_4921 , w_4922 , w_4923 , w_4924 , w_4925 , 
		w_4926 , w_4927 , w_4928 , w_4929 , w_4930 , w_4931 , w_4932 , w_4933 , w_4934 , w_4935 , 
		w_4936 , w_4937 , w_4938 , w_4939 , w_4940 , w_4941 , w_4942 , w_4943 , w_4944 , w_4945 , 
		w_4946 , w_4947 , w_4948 , w_4949 , w_4950 , w_4951 , w_4952 , w_4953 , w_4954 , w_4955 , 
		w_4956 , w_4957 , w_4958 , w_4959 , w_4960 , w_4961 , w_4962 , w_4963 , w_4964 , w_4965 , 
		w_4966 , w_4967 , w_4968 , w_4969 , w_4970 , w_4971 , w_4972 , w_4973 , w_4974 , w_4975 , 
		w_4976 , w_4977 , w_4978 , w_4979 , w_4980 , w_4981 , w_4982 , w_4983 , w_4984 , w_4985 , 
		w_4986 , w_4987 , w_4988 , w_4989 , w_4990 , w_4991 , w_4992 , w_4993 , w_4994 , w_4995 , 
		w_4996 , w_4997 , w_4998 , w_4999 , w_5000 , w_5001 , w_5002 , w_5003 , w_5004 , w_5005 , 
		w_5006 , w_5007 , w_5008 , w_5009 , w_5010 , w_5011 , w_5012 , w_5013 , w_5014 , w_5015 , 
		w_5016 , w_5017 , w_5018 , w_5019 , w_5020 , w_5021 , w_5022 , w_5023 , w_5024 , w_5025 , 
		w_5026 , w_5027 , w_5028 , w_5029 , w_5030 , w_5031 , w_5032 , w_5033 , w_5034 , w_5035 , 
		w_5036 , w_5037 , w_5038 , w_5039 , w_5040 , w_5041 , w_5042 , w_5043 , w_5044 , w_5045 , 
		w_5046 , w_5047 , w_5048 , w_5049 , w_5050 , w_5051 , w_5052 , w_5053 , w_5054 , w_5055 , 
		w_5056 , w_5057 , w_5058 , w_5059 , w_5060 , w_5061 , w_5062 , w_5063 , w_5064 , w_5065 , 
		w_5066 , w_5067 , w_5068 , w_5069 , w_5070 , w_5071 , w_5072 , w_5073 , w_5074 , w_5075 , 
		w_5076 , w_5077 , w_5078 , w_5079 , w_5080 , w_5081 , w_5082 , w_5083 , w_5084 , w_5085 , 
		w_5086 , w_5087 , w_5088 , w_5089 , w_5090 , w_5091 , w_5092 , w_5093 , w_5094 , w_5095 , 
		w_5096 , w_5097 , w_5098 , w_5099 , w_5100 , w_5101 , w_5102 , w_5103 , w_5104 , w_5105 , 
		w_5106 , w_5107 , w_5108 , w_5109 , w_5110 , w_5111 , w_5112 , w_5113 , w_5114 , w_5115 , 
		w_5116 , w_5117 , w_5118 , w_5119 , w_5120 , w_5121 , w_5122 , w_5123 , w_5124 , w_5125 , 
		w_5126 , w_5127 , w_5128 , w_5129 , w_5130 , w_5131 , w_5132 , w_5133 , w_5134 , w_5135 , 
		w_5136 , w_5137 , w_5138 , w_5139 , w_5140 , w_5141 , w_5142 , w_5143 , w_5144 , w_5145 , 
		w_5146 , w_5147 , w_5148 , w_5149 , w_5150 , w_5151 , w_5152 , w_5153 , w_5154 , w_5155 , 
		w_5156 , w_5157 , w_5158 , w_5159 , w_5160 , w_5161 , w_5162 , w_5163 , w_5164 , w_5165 , 
		w_5166 , w_5167 , w_5168 , w_5169 , w_5170 , w_5171 , w_5172 , w_5173 , w_5174 , w_5175 , 
		w_5176 , w_5177 , w_5178 , w_5179 , w_5180 , w_5181 , w_5182 , w_5183 , w_5184 , w_5185 , 
		w_5186 , w_5187 , w_5188 , w_5189 , w_5190 , w_5191 , w_5192 , w_5193 , w_5194 , w_5195 , 
		w_5196 , w_5197 , w_5198 , w_5199 , w_5200 , w_5201 , w_5202 , w_5203 , w_5204 , w_5205 , 
		w_5206 , w_5207 , w_5208 , w_5209 , w_5210 , w_5211 , w_5212 , w_5213 , w_5214 , w_5215 , 
		w_5216 , w_5217 , w_5218 , w_5219 , w_5220 , w_5221 , w_5222 , w_5223 , w_5224 , w_5225 , 
		w_5226 , w_5227 , w_5228 , w_5229 , w_5230 , w_5231 , w_5232 , w_5233 , w_5234 , w_5235 , 
		w_5236 , w_5237 , w_5238 , w_5239 , w_5240 , w_5241 , w_5242 , w_5243 , w_5244 , w_5245 , 
		w_5246 , w_5247 , w_5248 , w_5249 , w_5250 , w_5251 , w_5252 , w_5253 , w_5254 , w_5255 , 
		w_5256 , w_5257 , w_5258 , w_5259 , w_5260 , w_5261 , w_5262 , w_5263 , w_5264 , w_5265 , 
		w_5266 , w_5267 , w_5268 , w_5269 , w_5270 , w_5271 , w_5272 , w_5273 , w_5274 , w_5275 , 
		w_5276 , w_5277 , w_5278 , w_5279 , w_5280 , w_5281 , w_5282 , w_5283 , w_5284 , w_5285 , 
		w_5286 , w_5287 , w_5288 , w_5289 , w_5290 , w_5291 , w_5292 , w_5293 , w_5294 , w_5295 , 
		w_5296 , w_5297 , w_5298 , w_5299 , w_5300 , w_5301 , w_5302 , w_5303 , w_5304 , w_5305 , 
		w_5306 , w_5307 , w_5308 , w_5309 , w_5310 , w_5311 , w_5312 , w_5313 , w_5314 , w_5315 , 
		w_5316 , w_5317 , w_5318 , w_5319 , w_5320 , w_5321 , w_5322 , w_5323 , w_5324 , w_5325 , 
		w_5326 , w_5327 , w_5328 , w_5329 , w_5330 , w_5331 , w_5332 , w_5333 , w_5334 , w_5335 , 
		w_5336 , w_5337 , w_5338 , w_5339 , w_5340 , w_5341 , w_5342 , w_5343 , w_5344 , w_5345 , 
		w_5346 , w_5347 , w_5348 , w_5349 , w_5350 , w_5351 , w_5352 , w_5353 , w_5354 , w_5355 , 
		w_5356 , w_5357 , w_5358 , w_5359 , w_5360 , w_5361 , w_5362 , w_5363 , w_5364 , w_5365 , 
		w_5366 , w_5367 , w_5368 , w_5369 , w_5370 , w_5371 , w_5372 , w_5373 , w_5374 , w_5375 , 
		w_5376 , w_5377 , w_5378 , w_5379 , w_5380 , w_5381 , w_5382 , w_5383 , w_5384 , w_5385 , 
		w_5386 , w_5387 , w_5388 , w_5389 , w_5390 , w_5391 , w_5392 , w_5393 , w_5394 , w_5395 , 
		w_5396 , w_5397 , w_5398 , w_5399 , w_5400 , w_5401 , w_5402 , w_5403 , w_5404 , w_5405 , 
		w_5406 , w_5407 , w_5408 , w_5409 , w_5410 , w_5411 , w_5412 , w_5413 , w_5414 , w_5415 , 
		w_5416 , w_5417 , w_5418 , w_5419 , w_5420 , w_5421 , w_5422 , w_5423 , w_5424 , w_5425 , 
		w_5426 , w_5427 , w_5428 , w_5429 , w_5430 , w_5431 , w_5432 , w_5433 , w_5434 , w_5435 , 
		w_5436 , w_5437 , w_5438 , w_5439 , w_5440 , w_5441 , w_5442 , w_5443 , w_5444 , w_5445 , 
		w_5446 , w_5447 , w_5448 , w_5449 , w_5450 , w_5451 , w_5452 , w_5453 , w_5454 , w_5455 , 
		w_5456 , w_5457 , w_5458 , w_5459 , w_5460 , w_5461 , w_5462 , w_5463 , w_5464 , w_5465 , 
		w_5466 , w_5467 , w_5468 , w_5469 , w_5470 , w_5471 , w_5472 , w_5473 , w_5474 , w_5475 , 
		w_5476 , w_5477 , w_5478 , w_5479 , w_5480 , w_5481 , w_5482 , w_5483 , w_5484 , w_5485 , 
		w_5486 , w_5487 , w_5488 , w_5489 , w_5490 , w_5491 , w_5492 , w_5493 , w_5494 , w_5495 , 
		w_5496 , w_5497 , w_5498 , w_5499 , w_5500 , w_5501 , w_5502 , w_5503 , w_5504 , w_5505 , 
		w_5506 , w_5507 , w_5508 , w_5509 , w_5510 , w_5511 , w_5512 , w_5513 , w_5514 , w_5515 , 
		w_5516 , w_5517 , w_5518 , w_5519 , w_5520 , w_5521 , w_5522 , w_5523 , w_5524 , w_5525 , 
		w_5526 , w_5527 , w_5528 , w_5529 , w_5530 , w_5531 , w_5532 , w_5533 , w_5534 , w_5535 , 
		w_5536 , w_5537 , w_5538 , w_5539 , w_5540 , w_5541 , w_5542 , w_5543 , w_5544 , w_5545 , 
		w_5546 , w_5547 , w_5548 , w_5549 , w_5550 , w_5551 , w_5552 , w_5553 , w_5554 , w_5555 , 
		w_5556 , w_5557 , w_5558 , w_5559 , w_5560 , w_5561 , w_5562 , w_5563 , w_5564 , w_5565 , 
		w_5566 , w_5567 , w_5568 , w_5569 , w_5570 , w_5571 , w_5572 , w_5573 , w_5574 , w_5575 , 
		w_5576 , w_5577 , w_5578 , w_5579 , w_5580 , w_5581 , w_5582 , w_5583 , w_5584 , w_5585 , 
		w_5586 , w_5587 , w_5588 , w_5589 , w_5590 , w_5591 , w_5592 , w_5593 , w_5594 , w_5595 , 
		w_5596 , w_5597 , w_5598 , w_5599 , w_5600 , w_5601 , w_5602 , w_5603 , w_5604 , w_5605 , 
		w_5606 , w_5607 , w_5608 , w_5609 , w_5610 , w_5611 , w_5612 , w_5613 , w_5614 , w_5615 , 
		w_5616 , w_5617 , w_5618 , w_5619 , w_5620 , w_5621 , w_5622 , w_5623 , w_5624 , w_5625 , 
		w_5626 , w_5627 , w_5628 , w_5629 , w_5630 , w_5631 , w_5632 , w_5633 , w_5634 , w_5635 , 
		w_5636 , w_5637 , w_5638 , w_5639 , w_5640 , w_5641 , w_5642 , w_5643 , w_5644 , w_5645 , 
		w_5646 , w_5647 , w_5648 , w_5649 , w_5650 , w_5651 , w_5652 , w_5653 , w_5654 , w_5655 , 
		w_5656 , w_5657 , w_5658 , w_5659 , w_5660 , w_5661 , w_5662 , w_5663 , w_5664 , w_5665 , 
		w_5666 , w_5667 , w_5668 , w_5669 , w_5670 , w_5671 , w_5672 , w_5673 , w_5674 , w_5675 , 
		w_5676 , w_5677 , w_5678 , w_5679 , w_5680 , w_5681 , w_5682 , w_5683 , w_5684 , w_5685 , 
		w_5686 , w_5687 , w_5688 , w_5689 , w_5690 , w_5691 , w_5692 , w_5693 , w_5694 , w_5695 , 
		w_5696 , w_5697 , w_5698 , w_5699 , w_5700 , w_5701 , w_5702 , w_5703 , w_5704 , w_5705 , 
		w_5706 , w_5707 , w_5708 , w_5709 , w_5710 , w_5711 , w_5712 , w_5713 , w_5714 , w_5715 , 
		w_5716 , w_5717 , w_5718 , w_5719 , w_5720 , w_5721 , w_5722 , w_5723 , w_5724 , w_5725 , 
		w_5726 , w_5727 , w_5728 , w_5729 , w_5730 , w_5731 , w_5732 , w_5733 , w_5734 , w_5735 , 
		w_5736 , w_5737 , w_5738 , w_5739 , w_5740 , w_5741 , w_5742 , w_5743 , w_5744 , w_5745 , 
		w_5746 , w_5747 , w_5748 , w_5749 , w_5750 , w_5751 , w_5752 , w_5753 , w_5754 , w_5755 , 
		w_5756 , w_5757 , w_5758 , w_5759 , w_5760 , w_5761 , w_5762 , w_5763 , w_5764 , w_5765 , 
		w_5766 , w_5767 , w_5768 , w_5769 , w_5770 , w_5771 , w_5772 , w_5773 , w_5774 , w_5775 , 
		w_5776 , w_5777 , w_5778 , w_5779 , w_5780 , w_5781 , w_5782 , w_5783 , w_5784 , w_5785 , 
		w_5786 , w_5787 , w_5788 , w_5789 , w_5790 , w_5791 , w_5792 , w_5793 , w_5794 , w_5795 , 
		w_5796 , w_5797 , w_5798 , w_5799 , w_5800 , w_5801 , w_5802 , w_5803 , w_5804 , w_5805 , 
		w_5806 , w_5807 , w_5808 , w_5809 , w_5810 , w_5811 , w_5812 , w_5813 , w_5814 , w_5815 , 
		w_5816 , w_5817 , w_5818 , w_5819 , w_5820 , w_5821 , w_5822 , w_5823 , w_5824 , w_5825 , 
		w_5826 , w_5827 , w_5828 , w_5829 , w_5830 , w_5831 , w_5832 , w_5833 , w_5834 , w_5835 , 
		w_5836 , w_5837 , w_5838 , w_5839 , w_5840 , w_5841 , w_5842 , w_5843 , w_5844 , w_5845 , 
		w_5846 , w_5847 , w_5848 , w_5849 , w_5850 , w_5851 , w_5852 , w_5853 , w_5854 , w_5855 , 
		w_5856 , w_5857 , w_5858 , w_5859 , w_5860 , w_5861 , w_5862 , w_5863 , w_5864 , w_5865 , 
		w_5866 , w_5867 , w_5868 , w_5869 , w_5870 , w_5871 , w_5872 , w_5873 , w_5874 , w_5875 , 
		w_5876 , w_5877 , w_5878 , w_5879 , w_5880 , w_5881 , w_5882 , w_5883 , w_5884 , w_5885 , 
		w_5886 , w_5887 , w_5888 , w_5889 , w_5890 , w_5891 , w_5892 , w_5893 , w_5894 , w_5895 , 
		w_5896 , w_5897 , w_5898 , w_5899 , w_5900 , w_5901 , w_5902 , w_5903 , w_5904 , w_5905 , 
		w_5906 , w_5907 , w_5908 , w_5909 , w_5910 , w_5911 , w_5912 , w_5913 , w_5914 , w_5915 , 
		w_5916 , w_5917 , w_5918 , w_5919 , w_5920 , w_5921 , w_5922 , w_5923 , w_5924 , w_5925 , 
		w_5926 , w_5927 , w_5928 , w_5929 , w_5930 , w_5931 , w_5932 , w_5933 , w_5934 , w_5935 , 
		w_5936 , w_5937 , w_5938 , w_5939 , w_5940 , w_5941 , w_5942 , w_5943 , w_5944 , w_5945 , 
		w_5946 , w_5947 , w_5948 , w_5949 , w_5950 , w_5951 , w_5952 , w_5953 , w_5954 , w_5955 , 
		w_5956 , w_5957 , w_5958 , w_5959 , w_5960 , w_5961 , w_5962 , w_5963 , w_5964 , w_5965 , 
		w_5966 , w_5967 , w_5968 , w_5969 , w_5970 , w_5971 , w_5972 , w_5973 , w_5974 , w_5975 , 
		w_5976 , w_5977 , w_5978 , w_5979 , w_5980 , w_5981 , w_5982 , w_5983 , w_5984 , w_5985 , 
		w_5986 , w_5987 , w_5988 , w_5989 , w_5990 , w_5991 , w_5992 , w_5993 , w_5994 , w_5995 , 
		w_5996 , w_5997 , w_5998 , w_5999 , w_6000 , w_6001 , w_6002 , w_6003 , w_6004 , w_6005 , 
		w_6006 , w_6007 , w_6008 , w_6009 , w_6010 , w_6011 , w_6012 , w_6013 , w_6014 , w_6015 , 
		w_6016 , w_6017 , w_6018 , w_6019 , w_6020 , w_6021 , w_6022 , w_6023 , w_6024 , w_6025 , 
		w_6026 , w_6027 , w_6028 , w_6029 , w_6030 , w_6031 , w_6032 , w_6033 , w_6034 , w_6035 , 
		w_6036 , w_6037 , w_6038 , w_6039 , w_6040 , w_6041 , w_6042 , w_6043 , w_6044 , w_6045 , 
		w_6046 , w_6047 , w_6048 , w_6049 , w_6050 , w_6051 , w_6052 , w_6053 , w_6054 , w_6055 , 
		w_6056 , w_6057 , w_6058 , w_6059 , w_6060 , w_6061 , w_6062 , w_6063 , w_6064 , w_6065 , 
		w_6066 , w_6067 , w_6068 , w_6069 , w_6070 , w_6071 , w_6072 , w_6073 , w_6074 , w_6075 , 
		w_6076 , w_6077 , w_6078 , w_6079 , w_6080 , w_6081 , w_6082 , w_6083 , w_6084 , w_6085 , 
		w_6086 , w_6087 , w_6088 , w_6089 , w_6090 , w_6091 , w_6092 , w_6093 , w_6094 , w_6095 , 
		w_6096 , w_6097 , w_6098 , w_6099 , w_6100 , w_6101 , w_6102 , w_6103 , w_6104 , w_6105 , 
		w_6106 , w_6107 , w_6108 , w_6109 , w_6110 , w_6111 , w_6112 , w_6113 , w_6114 , w_6115 , 
		w_6116 , w_6117 , w_6118 , w_6119 , w_6120 , w_6121 , w_6122 , w_6123 , w_6124 , w_6125 , 
		w_6126 , w_6127 , w_6128 , w_6129 , w_6130 , w_6131 , w_6132 , w_6133 , w_6134 , w_6135 , 
		w_6136 , w_6137 , w_6138 , w_6139 , w_6140 , w_6141 , w_6142 , w_6143 , w_6144 , w_6145 , 
		w_6146 , w_6147 , w_6148 , w_6149 , w_6150 , w_6151 , w_6152 , w_6153 , w_6154 , w_6155 , 
		w_6156 , w_6157 , w_6158 , w_6159 , w_6160 , w_6161 , w_6162 , w_6163 , w_6164 , w_6165 , 
		w_6166 , w_6167 , w_6168 , w_6169 , w_6170 , w_6171 , w_6172 , w_6173 , w_6174 , w_6175 , 
		w_6176 , w_6177 , w_6178 , w_6179 , w_6180 , w_6181 , w_6182 , w_6183 , w_6184 , w_6185 , 
		w_6186 , w_6187 , w_6188 , w_6189 , w_6190 , w_6191 , w_6192 , w_6193 , w_6194 , w_6195 , 
		w_6196 , w_6197 , w_6198 , w_6199 , w_6200 , w_6201 , w_6202 , w_6203 , w_6204 , w_6205 , 
		w_6206 , w_6207 , w_6208 , w_6209 , w_6210 , w_6211 , w_6212 , w_6213 , w_6214 , w_6215 , 
		w_6216 , w_6217 , w_6218 , w_6219 , w_6220 , w_6221 , w_6222 , w_6223 , w_6224 , w_6225 , 
		w_6226 , w_6227 , w_6228 , w_6229 , w_6230 , w_6231 , w_6232 , w_6233 , w_6234 , w_6235 , 
		w_6236 , w_6237 , w_6238 , w_6239 , w_6240 , w_6241 , w_6242 , w_6243 , w_6244 , w_6245 , 
		w_6246 , w_6247 , w_6248 , w_6249 , w_6250 , w_6251 , w_6252 , w_6253 , w_6254 , w_6255 , 
		w_6256 , w_6257 , w_6258 , w_6259 , w_6260 , w_6261 , w_6262 , w_6263 , w_6264 , w_6265 , 
		w_6266 , w_6267 , w_6268 , w_6269 , w_6270 , w_6271 , w_6272 , w_6273 , w_6274 , w_6275 , 
		w_6276 , w_6277 , w_6278 , w_6279 , w_6280 , w_6281 , w_6282 , w_6283 , w_6284 , w_6285 , 
		w_6286 , w_6287 , w_6288 , w_6289 , w_6290 , w_6291 , w_6292 , w_6293 , w_6294 , w_6295 , 
		w_6296 , w_6297 , w_6298 , w_6299 , w_6300 , w_6301 , w_6302 , w_6303 , w_6304 , w_6305 , 
		w_6306 , w_6307 , w_6308 , w_6309 , w_6310 , w_6311 , w_6312 , w_6313 , w_6314 , w_6315 , 
		w_6316 , w_6317 , w_6318 , w_6319 , w_6320 , w_6321 , w_6322 , w_6323 , w_6324 , w_6325 , 
		w_6326 , w_6327 , w_6328 , w_6329 , w_6330 , w_6331 , w_6332 , w_6333 , w_6334 , w_6335 , 
		w_6336 , w_6337 , w_6338 , w_6339 , w_6340 , w_6341 , w_6342 , w_6343 , w_6344 , w_6345 , 
		w_6346 , w_6347 , w_6348 , w_6349 , w_6350 , w_6351 , w_6352 , w_6353 , w_6354 , w_6355 , 
		w_6356 , w_6357 , w_6358 , w_6359 , w_6360 , w_6361 , w_6362 , w_6363 , w_6364 , w_6365 , 
		w_6366 , w_6367 , w_6368 , w_6369 , w_6370 , w_6371 , w_6372 , w_6373 , w_6374 , w_6375 , 
		w_6376 , w_6377 , w_6378 , w_6379 , w_6380 , w_6381 , w_6382 , w_6383 , w_6384 , w_6385 , 
		w_6386 , w_6387 , w_6388 , w_6389 , w_6390 , w_6391 , w_6392 , w_6393 , w_6394 , w_6395 , 
		w_6396 , w_6397 , w_6398 , w_6399 , w_6400 , w_6401 , w_6402 , w_6403 , w_6404 , w_6405 , 
		w_6406 , w_6407 , w_6408 , w_6409 , w_6410 , w_6411 , w_6412 , w_6413 , w_6414 , w_6415 , 
		w_6416 , w_6417 , w_6418 , w_6419 , w_6420 , w_6421 , w_6422 , w_6423 , w_6424 , w_6425 , 
		w_6426 , w_6427 , w_6428 , w_6429 , w_6430 , w_6431 , w_6432 , w_6433 , w_6434 , w_6435 , 
		w_6436 , w_6437 , w_6438 , w_6439 , w_6440 , w_6441 , w_6442 , w_6443 , w_6444 , w_6445 , 
		w_6446 , w_6447 , w_6448 , w_6449 , w_6450 , w_6451 , w_6452 , w_6453 , w_6454 , w_6455 , 
		w_6456 , w_6457 , w_6458 , w_6459 , w_6460 , w_6461 , w_6462 , w_6463 , w_6464 , w_6465 , 
		w_6466 , w_6467 , w_6468 , w_6469 , w_6470 , w_6471 , w_6472 , w_6473 , w_6474 , w_6475 , 
		w_6476 , w_6477 , w_6478 , w_6479 , w_6480 , w_6481 , w_6482 , w_6483 , w_6484 , w_6485 , 
		w_6486 , w_6487 , w_6488 , w_6489 , w_6490 , w_6491 , w_6492 , w_6493 , w_6494 , w_6495 , 
		w_6496 , w_6497 , w_6498 , w_6499 , w_6500 , w_6501 , w_6502 , w_6503 , w_6504 , w_6505 , 
		w_6506 , w_6507 , w_6508 , w_6509 , w_6510 , w_6511 , w_6512 , w_6513 , w_6514 , w_6515 , 
		w_6516 , w_6517 , w_6518 , w_6519 , w_6520 , w_6521 , w_6522 , w_6523 , w_6524 , w_6525 , 
		w_6526 , w_6527 , w_6528 , w_6529 , w_6530 , w_6531 , w_6532 , w_6533 , w_6534 , w_6535 , 
		w_6536 , w_6537 , w_6538 , w_6539 , w_6540 , w_6541 , w_6542 , w_6543 , w_6544 , w_6545 , 
		w_6546 , w_6547 , w_6548 , w_6549 , w_6550 , w_6551 , w_6552 , w_6553 , w_6554 , w_6555 , 
		w_6556 , w_6557 , w_6558 , w_6559 , w_6560 , w_6561 , w_6562 , w_6563 , w_6564 , w_6565 , 
		w_6566 , w_6567 , w_6568 , w_6569 , w_6570 , w_6571 , w_6572 , w_6573 , w_6574 , w_6575 , 
		w_6576 , w_6577 , w_6578 , w_6579 , w_6580 , w_6581 , w_6582 , w_6583 , w_6584 , w_6585 , 
		w_6586 , w_6587 , w_6588 , w_6589 , w_6590 , w_6591 , w_6592 , w_6593 , w_6594 , w_6595 , 
		w_6596 , w_6597 , w_6598 , w_6599 , w_6600 , w_6601 , w_6602 , w_6603 , w_6604 , w_6605 , 
		w_6606 , w_6607 , w_6608 , w_6609 , w_6610 , w_6611 , w_6612 , w_6613 , w_6614 , w_6615 , 
		w_6616 , w_6617 , w_6618 , w_6619 , w_6620 , w_6621 , w_6622 , w_6623 , w_6624 , w_6625 , 
		w_6626 , w_6627 , w_6628 , w_6629 , w_6630 , w_6631 , w_6632 , w_6633 , w_6634 , w_6635 , 
		w_6636 , w_6637 , w_6638 , w_6639 , w_6640 , w_6641 , w_6642 , w_6643 , w_6644 , w_6645 , 
		w_6646 , w_6647 , w_6648 , w_6649 , w_6650 , w_6651 , w_6652 , w_6653 , w_6654 , w_6655 , 
		w_6656 , w_6657 , w_6658 , w_6659 , w_6660 , w_6661 , w_6662 , w_6663 , w_6664 , w_6665 , 
		w_6666 , w_6667 , w_6668 , w_6669 , w_6670 , w_6671 , w_6672 , w_6673 , w_6674 , w_6675 , 
		w_6676 , w_6677 , w_6678 , w_6679 , w_6680 , w_6681 , w_6682 , w_6683 , w_6684 , w_6685 , 
		w_6686 , w_6687 , w_6688 , w_6689 , w_6690 , w_6691 , w_6692 , w_6693 , w_6694 , w_6695 , 
		w_6696 , w_6697 , w_6698 , w_6699 , w_6700 , w_6701 , w_6702 , w_6703 , w_6704 , w_6705 , 
		w_6706 , w_6707 , w_6708 , w_6709 , w_6710 , w_6711 , w_6712 , w_6713 , w_6714 , w_6715 , 
		w_6716 , w_6717 , w_6718 , w_6719 , w_6720 , w_6721 , w_6722 , w_6723 , w_6724 , w_6725 , 
		w_6726 , w_6727 , w_6728 , w_6729 , w_6730 , w_6731 , w_6732 , w_6733 , w_6734 , w_6735 , 
		w_6736 , w_6737 , w_6738 , w_6739 , w_6740 , w_6741 , w_6742 , w_6743 , w_6744 , w_6745 , 
		w_6746 , w_6747 , w_6748 , w_6749 , w_6750 , w_6751 , w_6752 , w_6753 , w_6754 , w_6755 , 
		w_6756 , w_6757 , w_6758 , w_6759 , w_6760 , w_6761 , w_6762 , w_6763 , w_6764 , w_6765 , 
		w_6766 , w_6767 , w_6768 , w_6769 , w_6770 , w_6771 , w_6772 , w_6773 , w_6774 , w_6775 , 
		w_6776 , w_6777 , w_6778 , w_6779 , w_6780 , w_6781 , w_6782 , w_6783 , w_6784 , w_6785 , 
		w_6786 , w_6787 , w_6788 , w_6789 , w_6790 , w_6791 , w_6792 , w_6793 , w_6794 , w_6795 , 
		w_6796 , w_6797 , w_6798 , w_6799 , w_6800 , w_6801 , w_6802 , w_6803 , w_6804 , w_6805 , 
		w_6806 , w_6807 , w_6808 , w_6809 , w_6810 , w_6811 , w_6812 , w_6813 , w_6814 , w_6815 , 
		w_6816 , w_6817 , w_6818 , w_6819 , w_6820 , w_6821 , w_6822 , w_6823 , w_6824 , w_6825 , 
		w_6826 , w_6827 , w_6828 , w_6829 , w_6830 , w_6831 , w_6832 , w_6833 , w_6834 , w_6835 , 
		w_6836 , w_6837 , w_6838 , w_6839 , w_6840 , w_6841 , w_6842 , w_6843 , w_6844 , w_6845 , 
		w_6846 , w_6847 , w_6848 , w_6849 , w_6850 , w_6851 , w_6852 , w_6853 , w_6854 , w_6855 , 
		w_6856 , w_6857 , w_6858 , w_6859 , w_6860 , w_6861 , w_6862 , w_6863 , w_6864 , w_6865 , 
		w_6866 , w_6867 , w_6868 , w_6869 , w_6870 , w_6871 , w_6872 , w_6873 , w_6874 , w_6875 , 
		w_6876 , w_6877 , w_6878 , w_6879 , w_6880 , w_6881 , w_6882 , w_6883 , w_6884 , w_6885 , 
		w_6886 , w_6887 , w_6888 , w_6889 , w_6890 , w_6891 , w_6892 , w_6893 , w_6894 , w_6895 , 
		w_6896 , w_6897 , w_6898 , w_6899 , w_6900 , w_6901 , w_6902 , w_6903 , w_6904 , w_6905 , 
		w_6906 , w_6907 , w_6908 , w_6909 , w_6910 , w_6911 , w_6912 , w_6913 , w_6914 , w_6915 , 
		w_6916 , w_6917 , w_6918 , w_6919 , w_6920 , w_6921 , w_6922 , w_6923 , w_6924 , w_6925 , 
		w_6926 , w_6927 , w_6928 , w_6929 , w_6930 , w_6931 , w_6932 , w_6933 , w_6934 , w_6935 , 
		w_6936 , w_6937 , w_6938 , w_6939 , w_6940 , w_6941 , w_6942 , w_6943 , w_6944 , w_6945 , 
		w_6946 , w_6947 , w_6948 , w_6949 , w_6950 , w_6951 , w_6952 , w_6953 , w_6954 , w_6955 , 
		w_6956 , w_6957 , w_6958 , w_6959 , w_6960 , w_6961 , w_6962 , w_6963 , w_6964 , w_6965 , 
		w_6966 , w_6967 , w_6968 , w_6969 , w_6970 , w_6971 , w_6972 , w_6973 , w_6974 , w_6975 , 
		w_6976 , w_6977 , w_6978 , w_6979 , w_6980 , w_6981 , w_6982 , w_6983 , w_6984 , w_6985 , 
		w_6986 , w_6987 , w_6988 , w_6989 , w_6990 , w_6991 , w_6992 , w_6993 , w_6994 , w_6995 , 
		w_6996 , w_6997 , w_6998 , w_6999 , w_7000 , w_7001 , w_7002 , w_7003 , w_7004 , w_7005 , 
		w_7006 , w_7007 , w_7008 , w_7009 , w_7010 , w_7011 , w_7012 , w_7013 , w_7014 , w_7015 , 
		w_7016 , w_7017 , w_7018 , w_7019 , w_7020 , w_7021 , w_7022 , w_7023 , w_7024 , w_7025 , 
		w_7026 , w_7027 , w_7028 , w_7029 , w_7030 , w_7031 , w_7032 , w_7033 , w_7034 , w_7035 , 
		w_7036 , w_7037 , w_7038 , w_7039 , w_7040 , w_7041 , w_7042 , w_7043 , w_7044 , w_7045 , 
		w_7046 , w_7047 , w_7048 , w_7049 , w_7050 , w_7051 , w_7052 , w_7053 , w_7054 , w_7055 , 
		w_7056 , w_7057 , w_7058 , w_7059 , w_7060 , w_7061 , w_7062 , w_7063 , w_7064 , w_7065 , 
		w_7066 , w_7067 , w_7068 , w_7069 , w_7070 , w_7071 , w_7072 , w_7073 , w_7074 , w_7075 , 
		w_7076 , w_7077 , w_7078 , w_7079 , w_7080 , w_7081 , w_7082 , w_7083 , w_7084 , w_7085 , 
		w_7086 , w_7087 , w_7088 , w_7089 , w_7090 , w_7091 , w_7092 , w_7093 , w_7094 , w_7095 , 
		w_7096 , w_7097 , w_7098 , w_7099 , w_7100 , w_7101 , w_7102 , w_7103 , w_7104 , w_7105 , 
		w_7106 , w_7107 , w_7108 , w_7109 , w_7110 , w_7111 , w_7112 , w_7113 , w_7114 , w_7115 , 
		w_7116 , w_7117 , w_7118 , w_7119 , w_7120 , w_7121 , w_7122 , w_7123 , w_7124 , w_7125 , 
		w_7126 , w_7127 , w_7128 , w_7129 , w_7130 , w_7131 , w_7132 , w_7133 , w_7134 , w_7135 , 
		w_7136 , w_7137 , w_7138 , w_7139 , w_7140 , w_7141 , w_7142 , w_7143 , w_7144 , w_7145 , 
		w_7146 , w_7147 , w_7148 , w_7149 , w_7150 , w_7151 , w_7152 , w_7153 , w_7154 , w_7155 , 
		w_7156 , w_7157 , w_7158 , w_7159 , w_7160 , w_7161 , w_7162 , w_7163 , w_7164 , w_7165 , 
		w_7166 , w_7167 , w_7168 , w_7169 , w_7170 , w_7171 , w_7172 , w_7173 , w_7174 , w_7175 , 
		w_7176 , w_7177 , w_7178 , w_7179 , w_7180 , w_7181 , w_7182 , w_7183 , w_7184 , w_7185 , 
		w_7186 , w_7187 , w_7188 , w_7189 , w_7190 , w_7191 , w_7192 , w_7193 , w_7194 , w_7195 , 
		w_7196 , w_7197 , w_7198 , w_7199 , w_7200 , w_7201 , w_7202 , w_7203 , w_7204 , w_7205 , 
		w_7206 , w_7207 , w_7208 , w_7209 , w_7210 , w_7211 , w_7212 , w_7213 , w_7214 , w_7215 , 
		w_7216 , w_7217 , w_7218 , w_7219 , w_7220 , w_7221 , w_7222 , w_7223 , w_7224 , w_7225 , 
		w_7226 , w_7227 , w_7228 , w_7229 , w_7230 , w_7231 , w_7232 , w_7233 , w_7234 , w_7235 , 
		w_7236 , w_7237 , w_7238 , w_7239 , w_7240 , w_7241 , w_7242 , w_7243 , w_7244 , w_7245 , 
		w_7246 , w_7247 , w_7248 , w_7249 , w_7250 , w_7251 , w_7252 , w_7253 , w_7254 , w_7255 , 
		w_7256 , w_7257 , w_7258 , w_7259 , w_7260 , w_7261 , w_7262 , w_7263 , w_7264 , w_7265 , 
		w_7266 , w_7267 , w_7268 , w_7269 , w_7270 , w_7271 , w_7272 , w_7273 , w_7274 , w_7275 , 
		w_7276 , w_7277 , w_7278 , w_7279 , w_7280 , w_7281 , w_7282 , w_7283 , w_7284 , w_7285 , 
		w_7286 , w_7287 , w_7288 , w_7289 , w_7290 , w_7291 , w_7292 , w_7293 , w_7294 , w_7295 , 
		w_7296 , w_7297 , w_7298 , w_7299 , w_7300 , w_7301 , w_7302 , w_7303 , w_7304 , w_7305 , 
		w_7306 , w_7307 , w_7308 , w_7309 , w_7310 , w_7311 , w_7312 , w_7313 , w_7314 , w_7315 , 
		w_7316 , w_7317 , w_7318 , w_7319 , w_7320 , w_7321 , w_7322 , w_7323 , w_7324 , w_7325 , 
		w_7326 , w_7327 , w_7328 , w_7329 , w_7330 , w_7331 , w_7332 , w_7333 , w_7334 , w_7335 , 
		w_7336 , w_7337 , w_7338 , w_7339 , w_7340 , w_7341 , w_7342 , w_7343 , w_7344 , w_7345 , 
		w_7346 , w_7347 , w_7348 , w_7349 , w_7350 , w_7351 , w_7352 , w_7353 , w_7354 , w_7355 , 
		w_7356 , w_7357 , w_7358 , w_7359 , w_7360 , w_7361 , w_7362 , w_7363 , w_7364 , w_7365 , 
		w_7366 , w_7367 , w_7368 , w_7369 , w_7370 , w_7371 , w_7372 , w_7373 , w_7374 , w_7375 , 
		w_7376 , w_7377 , w_7378 , w_7379 , w_7380 , w_7381 , w_7382 , w_7383 , w_7384 , w_7385 , 
		w_7386 , w_7387 , w_7388 , w_7389 , w_7390 , w_7391 , w_7392 , w_7393 , w_7394 , w_7395 , 
		w_7396 , w_7397 , w_7398 , w_7399 , w_7400 , w_7401 , w_7402 , w_7403 , w_7404 , w_7405 , 
		w_7406 , w_7407 , w_7408 , w_7409 , w_7410 , w_7411 , w_7412 , w_7413 , w_7414 , w_7415 , 
		w_7416 , w_7417 , w_7418 , w_7419 , w_7420 , w_7421 , w_7422 , w_7423 , w_7424 , w_7425 , 
		w_7426 , w_7427 , w_7428 , w_7429 , w_7430 , w_7431 , w_7432 , w_7433 , w_7434 , w_7435 , 
		w_7436 , w_7437 , w_7438 , w_7439 , w_7440 , w_7441 , w_7442 , w_7443 , w_7444 , w_7445 , 
		w_7446 , w_7447 , w_7448 , w_7449 , w_7450 , w_7451 , w_7452 , w_7453 , w_7454 , w_7455 , 
		w_7456 , w_7457 , w_7458 , w_7459 , w_7460 , w_7461 , w_7462 , w_7463 , w_7464 , w_7465 , 
		w_7466 , w_7467 , w_7468 , w_7469 , w_7470 , w_7471 , w_7472 , w_7473 , w_7474 , w_7475 , 
		w_7476 , w_7477 , w_7478 , w_7479 , w_7480 , w_7481 , w_7482 , w_7483 , w_7484 , w_7485 , 
		w_7486 , w_7487 , w_7488 , w_7489 , w_7490 , w_7491 , w_7492 , w_7493 , w_7494 , w_7495 , 
		w_7496 , w_7497 , w_7498 , w_7499 , w_7500 , w_7501 , w_7502 , w_7503 , w_7504 , w_7505 , 
		w_7506 , w_7507 , w_7508 , w_7509 , w_7510 , w_7511 , w_7512 , w_7513 , w_7514 , w_7515 , 
		w_7516 , w_7517 , w_7518 , w_7519 , w_7520 , w_7521 , w_7522 , w_7523 , w_7524 , w_7525 , 
		w_7526 , w_7527 , w_7528 , w_7529 , w_7530 , w_7531 , w_7532 , w_7533 , w_7534 , w_7535 , 
		w_7536 , w_7537 , w_7538 , w_7539 , w_7540 , w_7541 , w_7542 , w_7543 , w_7544 , w_7545 , 
		w_7546 , w_7547 , w_7548 , w_7549 , w_7550 , w_7551 , w_7552 , w_7553 , w_7554 , w_7555 , 
		w_7556 , w_7557 , w_7558 , w_7559 , w_7560 , w_7561 , w_7562 , w_7563 , w_7564 , w_7565 , 
		w_7566 , w_7567 , w_7568 , w_7569 , w_7570 , w_7571 , w_7572 , w_7573 , w_7574 , w_7575 , 
		w_7576 , w_7577 , w_7578 , w_7579 , w_7580 , w_7581 , w_7582 , w_7583 , w_7584 , w_7585 , 
		w_7586 , w_7587 , w_7588 , w_7589 , w_7590 , w_7591 , w_7592 , w_7593 , w_7594 , w_7595 , 
		w_7596 , w_7597 , w_7598 , w_7599 , w_7600 , w_7601 , w_7602 , w_7603 , w_7604 , w_7605 , 
		w_7606 , w_7607 , w_7608 , w_7609 , w_7610 , w_7611 , w_7612 , w_7613 , w_7614 , w_7615 , 
		w_7616 , w_7617 , w_7618 , w_7619 , w_7620 , w_7621 , w_7622 , w_7623 , w_7624 , w_7625 , 
		w_7626 , w_7627 , w_7628 , w_7629 , w_7630 , w_7631 , w_7632 , w_7633 , w_7634 , w_7635 , 
		w_7636 , w_7637 , w_7638 , w_7639 , w_7640 , w_7641 , w_7642 , w_7643 , w_7644 , w_7645 , 
		w_7646 , w_7647 , w_7648 , w_7649 , w_7650 , w_7651 , w_7652 , w_7653 , w_7654 , w_7655 , 
		w_7656 , w_7657 , w_7658 , w_7659 , w_7660 , w_7661 , w_7662 , w_7663 , w_7664 , w_7665 , 
		w_7666 , w_7667 , w_7668 , w_7669 , w_7670 , w_7671 , w_7672 , w_7673 , w_7674 , w_7675 , 
		w_7676 , w_7677 , w_7678 , w_7679 , w_7680 , w_7681 , w_7682 , w_7683 , w_7684 , w_7685 , 
		w_7686 , w_7687 , w_7688 , w_7689 , w_7690 , w_7691 , w_7692 , w_7693 , w_7694 , w_7695 , 
		w_7696 , w_7697 , w_7698 , w_7699 , w_7700 , w_7701 , w_7702 , w_7703 , w_7704 , w_7705 , 
		w_7706 , w_7707 , w_7708 , w_7709 , w_7710 , w_7711 , w_7712 , w_7713 , w_7714 , w_7715 , 
		w_7716 , w_7717 , w_7718 , w_7719 , w_7720 , w_7721 , w_7722 , w_7723 , w_7724 , w_7725 , 
		w_7726 , w_7727 , w_7728 , w_7729 , w_7730 , w_7731 , w_7732 , w_7733 , w_7734 , w_7735 , 
		w_7736 , w_7737 , w_7738 , w_7739 , w_7740 , w_7741 , w_7742 , w_7743 , w_7744 , w_7745 , 
		w_7746 , w_7747 , w_7748 , w_7749 , w_7750 , w_7751 , w_7752 , w_7753 , w_7754 , w_7755 , 
		w_7756 , w_7757 , w_7758 , w_7759 , w_7760 , w_7761 , w_7762 , w_7763 , w_7764 , w_7765 , 
		w_7766 , w_7767 , w_7768 , w_7769 , w_7770 , w_7771 , w_7772 , w_7773 , w_7774 , w_7775 , 
		w_7776 , w_7777 , w_7778 , w_7779 , w_7780 , w_7781 , w_7782 , w_7783 , w_7784 , w_7785 , 
		w_7786 , w_7787 , w_7788 , w_7789 , w_7790 , w_7791 , w_7792 , w_7793 , w_7794 , w_7795 , 
		w_7796 , w_7797 , w_7798 , w_7799 , w_7800 , w_7801 , w_7802 , w_7803 , w_7804 , w_7805 , 
		w_7806 , w_7807 , w_7808 , w_7809 , w_7810 , w_7811 , w_7812 , w_7813 , w_7814 , w_7815 , 
		w_7816 , w_7817 , w_7818 , w_7819 , w_7820 , w_7821 , w_7822 , w_7823 , w_7824 , w_7825 , 
		w_7826 , w_7827 , w_7828 , w_7829 , w_7830 , w_7831 , w_7832 , w_7833 , w_7834 , w_7835 , 
		w_7836 , w_7837 , w_7838 , w_7839 , w_7840 , w_7841 , w_7842 , w_7843 , w_7844 , w_7845 , 
		w_7846 , w_7847 , w_7848 , w_7849 , w_7850 , w_7851 , w_7852 , w_7853 , w_7854 , w_7855 , 
		w_7856 , w_7857 , w_7858 , w_7859 , w_7860 , w_7861 , w_7862 , w_7863 , w_7864 , w_7865 , 
		w_7866 , w_7867 , w_7868 , w_7869 , w_7870 , w_7871 , w_7872 , w_7873 , w_7874 , w_7875 , 
		w_7876 , w_7877 , w_7878 , w_7879 , w_7880 , w_7881 , w_7882 , w_7883 , w_7884 , w_7885 , 
		w_7886 , w_7887 , w_7888 , w_7889 , w_7890 , w_7891 , w_7892 , w_7893 , w_7894 , w_7895 , 
		w_7896 , w_7897 , w_7898 , w_7899 , w_7900 , w_7901 , w_7902 , w_7903 , w_7904 , w_7905 , 
		w_7906 , w_7907 , w_7908 , w_7909 , w_7910 , w_7911 , w_7912 , w_7913 , w_7914 , w_7915 , 
		w_7916 , w_7917 , w_7918 , w_7919 , w_7920 , w_7921 , w_7922 , w_7923 , w_7924 , w_7925 , 
		w_7926 , w_7927 , w_7928 , w_7929 , w_7930 , w_7931 , w_7932 , w_7933 , w_7934 , w_7935 , 
		w_7936 , w_7937 , w_7938 , w_7939 , w_7940 , w_7941 , w_7942 , w_7943 , w_7944 , w_7945 , 
		w_7946 , w_7947 , w_7948 , w_7949 , w_7950 , w_7951 , w_7952 , w_7953 , w_7954 , w_7955 , 
		w_7956 , w_7957 , w_7958 , w_7959 , w_7960 , w_7961 , w_7962 , w_7963 , w_7964 , w_7965 , 
		w_7966 , w_7967 , w_7968 , w_7969 , w_7970 , w_7971 , w_7972 , w_7973 , w_7974 , w_7975 , 
		w_7976 , w_7977 , w_7978 , w_7979 , w_7980 , w_7981 , w_7982 , w_7983 , w_7984 , w_7985 , 
		w_7986 , w_7987 , w_7988 , w_7989 , w_7990 , w_7991 , w_7992 , w_7993 , w_7994 , w_7995 , 
		w_7996 , w_7997 , w_7998 , w_7999 , w_8000 , w_8001 , w_8002 , w_8003 , w_8004 , w_8005 , 
		w_8006 , w_8007 , w_8008 , w_8009 , w_8010 , w_8011 , w_8012 , w_8013 , w_8014 , w_8015 , 
		w_8016 , w_8017 , w_8018 , w_8019 , w_8020 , w_8021 , w_8022 , w_8023 , w_8024 , w_8025 , 
		w_8026 , w_8027 , w_8028 , w_8029 , w_8030 , w_8031 , w_8032 , w_8033 , w_8034 , w_8035 , 
		w_8036 , w_8037 , w_8038 , w_8039 , w_8040 , w_8041 , w_8042 , w_8043 , w_8044 , w_8045 , 
		w_8046 , w_8047 , w_8048 , w_8049 , w_8050 , w_8051 , w_8052 , w_8053 , w_8054 , w_8055 , 
		w_8056 , w_8057 , w_8058 , w_8059 , w_8060 , w_8061 , w_8062 , w_8063 , w_8064 , w_8065 , 
		w_8066 , w_8067 , w_8068 , w_8069 , w_8070 , w_8071 , w_8072 , w_8073 , w_8074 , w_8075 , 
		w_8076 , w_8077 , w_8078 , w_8079 , w_8080 , w_8081 , w_8082 , w_8083 , w_8084 , w_8085 , 
		w_8086 , w_8087 , w_8088 , w_8089 , w_8090 , w_8091 , w_8092 , w_8093 , w_8094 , w_8095 , 
		w_8096 , w_8097 , w_8098 , w_8099 , w_8100 , w_8101 , w_8102 , w_8103 , w_8104 , w_8105 , 
		w_8106 , w_8107 , w_8108 , w_8109 , w_8110 , w_8111 , w_8112 , w_8113 , w_8114 , w_8115 , 
		w_8116 , w_8117 , w_8118 , w_8119 , w_8120 , w_8121 , w_8122 , w_8123 , w_8124 , w_8125 , 
		w_8126 , w_8127 , w_8128 , w_8129 , w_8130 , w_8131 , w_8132 , w_8133 , w_8134 , w_8135 , 
		w_8136 , w_8137 , w_8138 , w_8139 , w_8140 , w_8141 , w_8142 , w_8143 , w_8144 , w_8145 , 
		w_8146 , w_8147 , w_8148 , w_8149 , w_8150 , w_8151 , w_8152 , w_8153 , w_8154 , w_8155 , 
		w_8156 , w_8157 , w_8158 , w_8159 , w_8160 , w_8161 , w_8162 , w_8163 , w_8164 , w_8165 , 
		w_8166 , w_8167 , w_8168 , w_8169 , w_8170 , w_8171 , w_8172 , w_8173 , w_8174 , w_8175 , 
		w_8176 , w_8177 , w_8178 , w_8179 , w_8180 , w_8181 , w_8182 , w_8183 , w_8184 , w_8185 , 
		w_8186 , w_8187 , w_8188 , w_8189 , w_8190 , w_8191 , w_8192 , w_8193 , w_8194 , w_8195 , 
		w_8196 , w_8197 , w_8198 , w_8199 , w_8200 , w_8201 , w_8202 , w_8203 , w_8204 , w_8205 , 
		w_8206 , w_8207 , w_8208 , w_8209 , w_8210 , w_8211 , w_8212 , w_8213 , w_8214 , w_8215 , 
		w_8216 , w_8217 , w_8218 , w_8219 , w_8220 , w_8221 , w_8222 , w_8223 , w_8224 , w_8225 , 
		w_8226 , w_8227 , w_8228 , w_8229 , w_8230 , w_8231 , w_8232 , w_8233 , w_8234 , w_8235 , 
		w_8236 , w_8237 , w_8238 , w_8239 , w_8240 , w_8241 , w_8242 , w_8243 , w_8244 , w_8245 , 
		w_8246 , w_8247 , w_8248 , w_8249 , w_8250 , w_8251 , w_8252 , w_8253 , w_8254 , w_8255 , 
		w_8256 , w_8257 , w_8258 , w_8259 , w_8260 , w_8261 , w_8262 , w_8263 , w_8264 , w_8265 , 
		w_8266 , w_8267 , w_8268 , w_8269 , w_8270 , w_8271 , w_8272 , w_8273 , w_8274 , w_8275 , 
		w_8276 , w_8277 , w_8278 , w_8279 , w_8280 , w_8281 , w_8282 , w_8283 , w_8284 , w_8285 , 
		w_8286 , w_8287 , w_8288 , w_8289 , w_8290 , w_8291 , w_8292 , w_8293 , w_8294 , w_8295 , 
		w_8296 , w_8297 , w_8298 , w_8299 , w_8300 , w_8301 , w_8302 , w_8303 , w_8304 , w_8305 , 
		w_8306 , w_8307 , w_8308 , w_8309 , w_8310 , w_8311 , w_8312 , w_8313 , w_8314 , w_8315 , 
		w_8316 , w_8317 , w_8318 , w_8319 , w_8320 , w_8321 , w_8322 , w_8323 , w_8324 , w_8325 , 
		w_8326 , w_8327 , w_8328 , w_8329 , w_8330 , w_8331 , w_8332 , w_8333 , w_8334 , w_8335 , 
		w_8336 , w_8337 , w_8338 , w_8339 , w_8340 , w_8341 , w_8342 , w_8343 , w_8344 , w_8345 , 
		w_8346 , w_8347 , w_8348 , w_8349 , w_8350 , w_8351 , w_8352 , w_8353 , w_8354 , w_8355 , 
		w_8356 , w_8357 , w_8358 , w_8359 , w_8360 , w_8361 , w_8362 , w_8363 , w_8364 , w_8365 , 
		w_8366 , w_8367 , w_8368 , w_8369 , w_8370 , w_8371 , w_8372 , w_8373 , w_8374 , w_8375 , 
		w_8376 , w_8377 , w_8378 , w_8379 , w_8380 , w_8381 , w_8382 , w_8383 , w_8384 , w_8385 , 
		w_8386 , w_8387 , w_8388 , w_8389 , w_8390 , w_8391 , w_8392 , w_8393 , w_8394 , w_8395 , 
		w_8396 , w_8397 , w_8398 , w_8399 , w_8400 , w_8401 , w_8402 , w_8403 , w_8404 , w_8405 , 
		w_8406 , w_8407 , w_8408 , w_8409 , w_8410 , w_8411 , w_8412 , w_8413 , w_8414 , w_8415 , 
		w_8416 , w_8417 , w_8418 , w_8419 , w_8420 , w_8421 , w_8422 , w_8423 , w_8424 , w_8425 , 
		w_8426 , w_8427 , w_8428 , w_8429 , w_8430 , w_8431 , w_8432 , w_8433 , w_8434 , w_8435 , 
		w_8436 , w_8437 , w_8438 , w_8439 , w_8440 , w_8441 , w_8442 , w_8443 , w_8444 , w_8445 , 
		w_8446 , w_8447 , w_8448 , w_8449 , w_8450 , w_8451 , w_8452 , w_8453 , w_8454 , w_8455 , 
		w_8456 , w_8457 , w_8458 , w_8459 , w_8460 , w_8461 , w_8462 , w_8463 , w_8464 , w_8465 , 
		w_8466 , w_8467 , w_8468 , w_8469 , w_8470 , w_8471 , w_8472 , w_8473 , w_8474 , w_8475 , 
		w_8476 , w_8477 , w_8478 , w_8479 , w_8480 , w_8481 , w_8482 , w_8483 , w_8484 , w_8485 , 
		w_8486 , w_8487 , w_8488 , w_8489 , w_8490 , w_8491 , w_8492 , w_8493 , w_8494 , w_8495 , 
		w_8496 , w_8497 , w_8498 , w_8499 , w_8500 , w_8501 , w_8502 , w_8503 , w_8504 , w_8505 , 
		w_8506 , w_8507 , w_8508 , w_8509 , w_8510 , w_8511 , w_8512 , w_8513 , w_8514 , w_8515 , 
		w_8516 , w_8517 , w_8518 , w_8519 , w_8520 , w_8521 , w_8522 , w_8523 , w_8524 , w_8525 , 
		w_8526 , w_8527 , w_8528 , w_8529 , w_8530 , w_8531 , w_8532 , w_8533 , w_8534 , w_8535 , 
		w_8536 , w_8537 , w_8538 , w_8539 , w_8540 , w_8541 , w_8542 , w_8543 , w_8544 , w_8545 , 
		w_8546 , w_8547 , w_8548 , w_8549 , w_8550 , w_8551 , w_8552 , w_8553 , w_8554 , w_8555 , 
		w_8556 , w_8557 , w_8558 , w_8559 , w_8560 , w_8561 , w_8562 , w_8563 , w_8564 , w_8565 , 
		w_8566 , w_8567 , w_8568 , w_8569 , w_8570 , w_8571 , w_8572 , w_8573 , w_8574 , w_8575 , 
		w_8576 , w_8577 , w_8578 , w_8579 , w_8580 , w_8581 , w_8582 , w_8583 , w_8584 , w_8585 , 
		w_8586 , w_8587 , w_8588 , w_8589 , w_8590 , w_8591 , w_8592 , w_8593 , w_8594 , w_8595 , 
		w_8596 , w_8597 , w_8598 , w_8599 , w_8600 , w_8601 , w_8602 , w_8603 , w_8604 , w_8605 , 
		w_8606 , w_8607 , w_8608 , w_8609 , w_8610 , w_8611 , w_8612 , w_8613 , w_8614 , w_8615 , 
		w_8616 , w_8617 , w_8618 , w_8619 , w_8620 , w_8621 , w_8622 , w_8623 , w_8624 , w_8625 , 
		w_8626 , w_8627 , w_8628 , w_8629 , w_8630 , w_8631 , w_8632 , w_8633 , w_8634 , w_8635 , 
		w_8636 , w_8637 , w_8638 , w_8639 , w_8640 , w_8641 , w_8642 , w_8643 , w_8644 , w_8645 , 
		w_8646 , w_8647 , w_8648 , w_8649 , w_8650 , w_8651 , w_8652 , w_8653 , w_8654 , w_8655 , 
		w_8656 , w_8657 , w_8658 , w_8659 , w_8660 , w_8661 , w_8662 , w_8663 , w_8664 , w_8665 , 
		w_8666 , w_8667 , w_8668 , w_8669 , w_8670 , w_8671 , w_8672 , w_8673 , w_8674 , w_8675 , 
		w_8676 , w_8677 , w_8678 , w_8679 , w_8680 , w_8681 , w_8682 , w_8683 , w_8684 , w_8685 , 
		w_8686 , w_8687 , w_8688 , w_8689 , w_8690 , w_8691 , w_8692 , w_8693 , w_8694 , w_8695 , 
		w_8696 , w_8697 , w_8698 , w_8699 , w_8700 , w_8701 , w_8702 , w_8703 , w_8704 , w_8705 , 
		w_8706 , w_8707 , w_8708 , w_8709 , w_8710 , w_8711 , w_8712 , w_8713 , w_8714 , w_8715 , 
		w_8716 , w_8717 , w_8718 , w_8719 , w_8720 , w_8721 , w_8722 , w_8723 , w_8724 , w_8725 , 
		w_8726 , w_8727 , w_8728 , w_8729 , w_8730 , w_8731 , w_8732 , w_8733 , w_8734 , w_8735 , 
		w_8736 , w_8737 , w_8738 , w_8739 , w_8740 , w_8741 , w_8742 , w_8743 , w_8744 , w_8745 , 
		w_8746 , w_8747 , w_8748 , w_8749 , w_8750 , w_8751 , w_8752 , w_8753 , w_8754 , w_8755 , 
		w_8756 , w_8757 , w_8758 , w_8759 , w_8760 , w_8761 , w_8762 , w_8763 , w_8764 , w_8765 , 
		w_8766 , w_8767 , w_8768 , w_8769 , w_8770 , w_8771 , w_8772 , w_8773 , w_8774 , w_8775 , 
		w_8776 , w_8777 , w_8778 , w_8779 , w_8780 , w_8781 , w_8782 , w_8783 , w_8784 , w_8785 , 
		w_8786 , w_8787 , w_8788 , w_8789 , w_8790 , w_8791 , w_8792 , w_8793 , w_8794 , w_8795 , 
		w_8796 , w_8797 , w_8798 , w_8799 , w_8800 , w_8801 , w_8802 , w_8803 , w_8804 , w_8805 , 
		w_8806 , w_8807 , w_8808 , w_8809 , w_8810 , w_8811 , w_8812 , w_8813 , w_8814 , w_8815 , 
		w_8816 , w_8817 , w_8818 , w_8819 , w_8820 , w_8821 , w_8822 , w_8823 , w_8824 , w_8825 , 
		w_8826 , w_8827 , w_8828 , w_8829 , w_8830 , w_8831 , w_8832 , w_8833 , w_8834 , w_8835 , 
		w_8836 , w_8837 , w_8838 , w_8839 , w_8840 , w_8841 , w_8842 , w_8843 , w_8844 , w_8845 , 
		w_8846 , w_8847 , w_8848 , w_8849 , w_8850 , w_8851 , w_8852 , w_8853 , w_8854 , w_8855 , 
		w_8856 , w_8857 , w_8858 , w_8859 , w_8860 , w_8861 , w_8862 , w_8863 , w_8864 , w_8865 , 
		w_8866 , w_8867 , w_8868 , w_8869 , w_8870 , w_8871 , w_8872 , w_8873 , w_8874 , w_8875 , 
		w_8876 , w_8877 , w_8878 , w_8879 , w_8880 , w_8881 , w_8882 , w_8883 , w_8884 , w_8885 , 
		w_8886 , w_8887 , w_8888 , w_8889 , w_8890 , w_8891 , w_8892 , w_8893 , w_8894 , w_8895 , 
		w_8896 , w_8897 , w_8898 , w_8899 , w_8900 , w_8901 , w_8902 , w_8903 , w_8904 , w_8905 , 
		w_8906 , w_8907 , w_8908 , w_8909 , w_8910 , w_8911 , w_8912 , w_8913 , w_8914 , w_8915 , 
		w_8916 , w_8917 , w_8918 , w_8919 , w_8920 , w_8921 , w_8922 , w_8923 , w_8924 , w_8925 , 
		w_8926 , w_8927 , w_8928 , w_8929 , w_8930 , w_8931 , w_8932 , w_8933 , w_8934 , w_8935 , 
		w_8936 , w_8937 , w_8938 , w_8939 , w_8940 , w_8941 , w_8942 , w_8943 , w_8944 , w_8945 , 
		w_8946 , w_8947 , w_8948 , w_8949 , w_8950 , w_8951 , w_8952 , w_8953 , w_8954 , w_8955 , 
		w_8956 , w_8957 , w_8958 , w_8959 , w_8960 , w_8961 , w_8962 , w_8963 , w_8964 , w_8965 , 
		w_8966 , w_8967 , w_8968 , w_8969 , w_8970 , w_8971 , w_8972 , w_8973 , w_8974 , w_8975 , 
		w_8976 , w_8977 , w_8978 , w_8979 , w_8980 , w_8981 , w_8982 , w_8983 , w_8984 , w_8985 , 
		w_8986 , w_8987 , w_8988 , w_8989 , w_8990 , w_8991 , w_8992 , w_8993 , w_8994 , w_8995 , 
		w_8996 , w_8997 , w_8998 , w_8999 , w_9000 , w_9001 , w_9002 , w_9003 , w_9004 , w_9005 , 
		w_9006 , w_9007 , w_9008 , w_9009 , w_9010 , w_9011 , w_9012 , w_9013 , w_9014 , w_9015 , 
		w_9016 , w_9017 , w_9018 , w_9019 , w_9020 , w_9021 , w_9022 , w_9023 , w_9024 , w_9025 , 
		w_9026 , w_9027 , w_9028 , w_9029 , w_9030 , w_9031 , w_9032 , w_9033 , w_9034 , w_9035 , 
		w_9036 , w_9037 , w_9038 , w_9039 , w_9040 , w_9041 , w_9042 , w_9043 , w_9044 , w_9045 , 
		w_9046 , w_9047 , w_9048 , w_9049 , w_9050 , w_9051 , w_9052 , w_9053 , w_9054 , w_9055 , 
		w_9056 , w_9057 , w_9058 , w_9059 , w_9060 , w_9061 , w_9062 , w_9063 , w_9064 , w_9065 , 
		w_9066 , w_9067 , w_9068 , w_9069 , w_9070 , w_9071 , w_9072 , w_9073 , w_9074 , w_9075 , 
		w_9076 , w_9077 , w_9078 , w_9079 , w_9080 , w_9081 , w_9082 , w_9083 , w_9084 , w_9085 , 
		w_9086 , w_9087 , w_9088 , w_9089 , w_9090 , w_9091 , w_9092 , w_9093 , w_9094 , w_9095 , 
		w_9096 , w_9097 , w_9098 , w_9099 , w_9100 , w_9101 , w_9102 , w_9103 , w_9104 , w_9105 , 
		w_9106 , w_9107 , w_9108 , w_9109 , w_9110 , w_9111 , w_9112 , w_9113 , w_9114 , w_9115 , 
		w_9116 , w_9117 , w_9118 , w_9119 , w_9120 , w_9121 , w_9122 , w_9123 , w_9124 , w_9125 , 
		w_9126 , w_9127 , w_9128 , w_9129 , w_9130 , w_9131 , w_9132 , w_9133 , w_9134 , w_9135 , 
		w_9136 , w_9137 , w_9138 , w_9139 , w_9140 , w_9141 , w_9142 , w_9143 , w_9144 , w_9145 , 
		w_9146 , w_9147 , w_9148 , w_9149 , w_9150 , w_9151 , w_9152 , w_9153 , w_9154 , w_9155 , 
		w_9156 , w_9157 , w_9158 , w_9159 , w_9160 , w_9161 , w_9162 , w_9163 , w_9164 , w_9165 , 
		w_9166 , w_9167 , w_9168 , w_9169 , w_9170 , w_9171 , w_9172 , w_9173 , w_9174 , w_9175 , 
		w_9176 , w_9177 , w_9178 , w_9179 , w_9180 , w_9181 , w_9182 , w_9183 , w_9184 , w_9185 , 
		w_9186 , w_9187 , w_9188 , w_9189 , w_9190 , w_9191 , w_9192 , w_9193 , w_9194 , w_9195 , 
		w_9196 , w_9197 , w_9198 , w_9199 , w_9200 , w_9201 , w_9202 , w_9203 , w_9204 , w_9205 , 
		w_9206 , w_9207 , w_9208 , w_9209 , w_9210 , w_9211 , w_9212 , w_9213 , w_9214 , w_9215 , 
		w_9216 , w_9217 , w_9218 , w_9219 , w_9220 , w_9221 , w_9222 , w_9223 , w_9224 , w_9225 , 
		w_9226 , w_9227 , w_9228 , w_9229 , w_9230 , w_9231 , w_9232 , w_9233 , w_9234 , w_9235 , 
		w_9236 , w_9237 , w_9238 , w_9239 , w_9240 , w_9241 , w_9242 , w_9243 , w_9244 , w_9245 , 
		w_9246 , w_9247 , w_9248 , w_9249 , w_9250 , w_9251 , w_9252 , w_9253 , w_9254 , w_9255 , 
		w_9256 , w_9257 , w_9258 , w_9259 , w_9260 , w_9261 , w_9262 , w_9263 , w_9264 , w_9265 , 
		w_9266 , w_9267 , w_9268 , w_9269 , w_9270 , w_9271 , w_9272 , w_9273 , w_9274 , w_9275 , 
		w_9276 , w_9277 , w_9278 , w_9279 , w_9280 , w_9281 , w_9282 , w_9283 , w_9284 , w_9285 , 
		w_9286 , w_9287 , w_9288 , w_9289 , w_9290 , w_9291 , w_9292 , w_9293 , w_9294 , w_9295 , 
		w_9296 , w_9297 , w_9298 , w_9299 , w_9300 , w_9301 , w_9302 , w_9303 , w_9304 , w_9305 , 
		w_9306 , w_9307 , w_9308 , w_9309 , w_9310 , w_9311 , w_9312 , w_9313 , w_9314 , w_9315 , 
		w_9316 , w_9317 , w_9318 , w_9319 , w_9320 , w_9321 , w_9322 , w_9323 , w_9324 , w_9325 , 
		w_9326 , w_9327 , w_9328 , w_9329 , w_9330 , w_9331 , w_9332 , w_9333 , w_9334 , w_9335 , 
		w_9336 , w_9337 , w_9338 , w_9339 , w_9340 , w_9341 , w_9342 , w_9343 , w_9344 , w_9345 , 
		w_9346 , w_9347 , w_9348 , w_9349 , w_9350 , w_9351 , w_9352 , w_9353 , w_9354 , w_9355 , 
		w_9356 , w_9357 , w_9358 , w_9359 , w_9360 , w_9361 , w_9362 , w_9363 , w_9364 , w_9365 , 
		w_9366 , w_9367 , w_9368 , w_9369 , w_9370 , w_9371 , w_9372 , w_9373 , w_9374 , w_9375 , 
		w_9376 , w_9377 , w_9378 , w_9379 , w_9380 , w_9381 , w_9382 , w_9383 , w_9384 , w_9385 , 
		w_9386 , w_9387 , w_9388 , w_9389 , w_9390 , w_9391 , w_9392 , w_9393 , w_9394 , w_9395 , 
		w_9396 , w_9397 , w_9398 , w_9399 , w_9400 , w_9401 , w_9402 , w_9403 , w_9404 , w_9405 , 
		w_9406 , w_9407 , w_9408 , w_9409 , w_9410 , w_9411 , w_9412 , w_9413 , w_9414 , w_9415 , 
		w_9416 , w_9417 , w_9418 , w_9419 , w_9420 , w_9421 , w_9422 , w_9423 , w_9424 , w_9425 , 
		w_9426 , w_9427 , w_9428 , w_9429 , w_9430 , w_9431 , w_9432 , w_9433 , w_9434 , w_9435 , 
		w_9436 , w_9437 , w_9438 , w_9439 , w_9440 , w_9441 , w_9442 , w_9443 , w_9444 , w_9445 , 
		w_9446 , w_9447 , w_9448 , w_9449 , w_9450 , w_9451 , w_9452 , w_9453 , w_9454 , w_9455 , 
		w_9456 , w_9457 , w_9458 , w_9459 , w_9460 , w_9461 , w_9462 , w_9463 , w_9464 , w_9465 , 
		w_9466 , w_9467 , w_9468 , w_9469 , w_9470 , w_9471 , w_9472 , w_9473 , w_9474 , w_9475 , 
		w_9476 , w_9477 , w_9478 , w_9479 , w_9480 , w_9481 , w_9482 , w_9483 , w_9484 , w_9485 , 
		w_9486 , w_9487 , w_9488 , w_9489 , w_9490 , w_9491 , w_9492 , w_9493 , w_9494 , w_9495 , 
		w_9496 , w_9497 , w_9498 , w_9499 , w_9500 , w_9501 , w_9502 , w_9503 , w_9504 , w_9505 , 
		w_9506 , w_9507 , w_9508 , w_9509 , w_9510 , w_9511 , w_9512 , w_9513 , w_9514 , w_9515 , 
		w_9516 , w_9517 , w_9518 , w_9519 , w_9520 , w_9521 , w_9522 , w_9523 , w_9524 , w_9525 , 
		w_9526 , w_9527 , w_9528 , w_9529 , w_9530 , w_9531 , w_9532 , w_9533 , w_9534 , w_9535 , 
		w_9536 , w_9537 , w_9538 , w_9539 , w_9540 , w_9541 , w_9542 , w_9543 , w_9544 , w_9545 , 
		w_9546 , w_9547 , w_9548 , w_9549 , w_9550 , w_9551 , w_9552 , w_9553 , w_9554 , w_9555 , 
		w_9556 , w_9557 , w_9558 , w_9559 , w_9560 , w_9561 , w_9562 , w_9563 , w_9564 , w_9565 , 
		w_9566 , w_9567 , w_9568 , w_9569 , w_9570 , w_9571 , w_9572 , w_9573 , w_9574 , w_9575 , 
		w_9576 , w_9577 , w_9578 , w_9579 , w_9580 , w_9581 , w_9582 , w_9583 , w_9584 , w_9585 , 
		w_9586 , w_9587 , w_9588 , w_9589 , w_9590 , w_9591 , w_9592 , w_9593 , w_9594 , w_9595 , 
		w_9596 , w_9597 , w_9598 , w_9599 , w_9600 , w_9601 , w_9602 , w_9603 , w_9604 , w_9605 , 
		w_9606 , w_9607 , w_9608 , w_9609 , w_9610 , w_9611 , w_9612 , w_9613 , w_9614 , w_9615 , 
		w_9616 , w_9617 , w_9618 , w_9619 , w_9620 , w_9621 , w_9622 , w_9623 , w_9624 , w_9625 , 
		w_9626 , w_9627 , w_9628 , w_9629 , w_9630 , w_9631 , w_9632 , w_9633 , w_9634 , w_9635 , 
		w_9636 , w_9637 , w_9638 , w_9639 , w_9640 , w_9641 , w_9642 , w_9643 , w_9644 , w_9645 , 
		w_9646 , w_9647 , w_9648 , w_9649 , w_9650 , w_9651 , w_9652 , w_9653 , w_9654 , w_9655 , 
		w_9656 , w_9657 , w_9658 , w_9659 , w_9660 , w_9661 , w_9662 , w_9663 , w_9664 , w_9665 , 
		w_9666 , w_9667 , w_9668 , w_9669 , w_9670 , w_9671 , w_9672 , w_9673 , w_9674 , w_9675 , 
		w_9676 , w_9677 , w_9678 , w_9679 , w_9680 , w_9681 , w_9682 , w_9683 , w_9684 , w_9685 , 
		w_9686 , w_9687 , w_9688 , w_9689 , w_9690 , w_9691 , w_9692 , w_9693 , w_9694 , w_9695 , 
		w_9696 , w_9697 , w_9698 , w_9699 , w_9700 , w_9701 , w_9702 , w_9703 , w_9704 , w_9705 , 
		w_9706 , w_9707 , w_9708 , w_9709 , w_9710 , w_9711 , w_9712 , w_9713 , w_9714 , w_9715 , 
		w_9716 , w_9717 , w_9718 , w_9719 , w_9720 , w_9721 , w_9722 , w_9723 , w_9724 , w_9725 , 
		w_9726 , w_9727 , w_9728 , w_9729 , w_9730 , w_9731 , w_9732 , w_9733 , w_9734 , w_9735 , 
		w_9736 , w_9737 , w_9738 , w_9739 , w_9740 , w_9741 , w_9742 , w_9743 , w_9744 , w_9745 , 
		w_9746 , w_9747 , w_9748 , w_9749 , w_9750 , w_9751 , w_9752 , w_9753 , w_9754 , w_9755 , 
		w_9756 , w_9757 , w_9758 , w_9759 , w_9760 , w_9761 , w_9762 , w_9763 , w_9764 , w_9765 , 
		w_9766 , w_9767 , w_9768 , w_9769 , w_9770 , w_9771 , w_9772 , w_9773 , w_9774 , w_9775 , 
		w_9776 , w_9777 , w_9778 , w_9779 , w_9780 , w_9781 , w_9782 , w_9783 , w_9784 , w_9785 , 
		w_9786 , w_9787 , w_9788 , w_9789 , w_9790 , w_9791 , w_9792 , w_9793 , w_9794 , w_9795 , 
		w_9796 , w_9797 , w_9798 , w_9799 , w_9800 , w_9801 , w_9802 , w_9803 , w_9804 , w_9805 , 
		w_9806 , w_9807 , w_9808 , w_9809 , w_9810 , w_9811 , w_9812 , w_9813 , w_9814 , w_9815 , 
		w_9816 , w_9817 , w_9818 , w_9819 , w_9820 , w_9821 , w_9822 , w_9823 , w_9824 , w_9825 , 
		w_9826 , w_9827 , w_9828 , w_9829 , w_9830 , w_9831 , w_9832 , w_9833 , w_9834 , w_9835 , 
		w_9836 , w_9837 , w_9838 , w_9839 , w_9840 , w_9841 , w_9842 , w_9843 , w_9844 , w_9845 , 
		w_9846 , w_9847 , w_9848 , w_9849 , w_9850 , w_9851 , w_9852 , w_9853 , w_9854 , w_9855 , 
		w_9856 , w_9857 , w_9858 , w_9859 , w_9860 , w_9861 , w_9862 , w_9863 , w_9864 , w_9865 , 
		w_9866 , w_9867 , w_9868 , w_9869 , w_9870 , w_9871 , w_9872 , w_9873 , w_9874 , w_9875 , 
		w_9876 , w_9877 , w_9878 , w_9879 , w_9880 , w_9881 , w_9882 , w_9883 , w_9884 , w_9885 , 
		w_9886 , w_9887 , w_9888 , w_9889 , w_9890 , w_9891 , w_9892 , w_9893 , w_9894 , w_9895 , 
		w_9896 , w_9897 , w_9898 , w_9899 , w_9900 , w_9901 , w_9902 , w_9903 , w_9904 , w_9905 , 
		w_9906 , w_9907 , w_9908 , w_9909 , w_9910 , w_9911 , w_9912 , w_9913 , w_9914 , w_9915 , 
		w_9916 , w_9917 , w_9918 , w_9919 , w_9920 , w_9921 , w_9922 , w_9923 , w_9924 , w_9925 , 
		w_9926 , w_9927 , w_9928 , w_9929 , w_9930 , w_9931 , w_9932 , w_9933 , w_9934 , w_9935 , 
		w_9936 , w_9937 , w_9938 , w_9939 , w_9940 , w_9941 , w_9942 , w_9943 , w_9944 , w_9945 , 
		w_9946 , w_9947 , w_9948 , w_9949 , w_9950 , w_9951 , w_9952 , w_9953 , w_9954 , w_9955 , 
		w_9956 , w_9957 , w_9958 , w_9959 , w_9960 , w_9961 , w_9962 , w_9963 , w_9964 , w_9965 , 
		w_9966 , w_9967 , w_9968 , w_9969 , w_9970 , w_9971 , w_9972 , w_9973 , w_9974 , w_9975 , 
		w_9976 , w_9977 , w_9978 , w_9979 , w_9980 , w_9981 , w_9982 , w_9983 , w_9984 , w_9985 , 
		w_9986 , w_9987 , w_9988 , w_9989 , w_9990 , w_9991 , w_9992 , w_9993 , w_9994 , w_9995 , 
		w_9996 , w_9997 , w_9998 , w_9999 , w_10000 , w_10001 , w_10002 , w_10003 , w_10004 , w_10005 , 
		w_10006 , w_10007 , w_10008 , w_10009 , w_10010 , w_10011 , w_10012 , w_10013 , w_10014 , w_10015 , 
		w_10016 , w_10017 , w_10018 , w_10019 , w_10020 , w_10021 , w_10022 , w_10023 , w_10024 , w_10025 , 
		w_10026 , w_10027 , w_10028 , w_10029 , w_10030 , w_10031 , w_10032 , w_10033 , w_10034 , w_10035 , 
		w_10036 , w_10037 , w_10038 , w_10039 , w_10040 , w_10041 , w_10042 , w_10043 , w_10044 , w_10045 , 
		w_10046 , w_10047 , w_10048 , w_10049 , w_10050 , w_10051 , w_10052 , w_10053 , w_10054 , w_10055 , 
		w_10056 , w_10057 , w_10058 , w_10059 , w_10060 , w_10061 , w_10062 , w_10063 , w_10064 , w_10065 , 
		w_10066 , w_10067 , w_10068 , w_10069 , w_10070 , w_10071 , w_10072 , w_10073 , w_10074 , w_10075 , 
		w_10076 , w_10077 , w_10078 , w_10079 , w_10080 , w_10081 , w_10082 , w_10083 , w_10084 , w_10085 , 
		w_10086 , w_10087 , w_10088 , w_10089 , w_10090 , w_10091 , w_10092 , w_10093 , w_10094 , w_10095 , 
		w_10096 , w_10097 , w_10098 , w_10099 , w_10100 , w_10101 , w_10102 , w_10103 , w_10104 , w_10105 , 
		w_10106 , w_10107 , w_10108 , w_10109 , w_10110 , w_10111 , w_10112 , w_10113 , w_10114 , w_10115 , 
		w_10116 , w_10117 , w_10118 , w_10119 , w_10120 , w_10121 , w_10122 , w_10123 , w_10124 , w_10125 , 
		w_10126 , w_10127 , w_10128 , w_10129 , w_10130 , w_10131 , w_10132 , w_10133 , w_10134 , w_10135 , 
		w_10136 , w_10137 , w_10138 , w_10139 , w_10140 , w_10141 , w_10142 , w_10143 , w_10144 , w_10145 , 
		w_10146 , w_10147 , w_10148 , w_10149 , w_10150 , w_10151 , w_10152 , w_10153 , w_10154 , w_10155 , 
		w_10156 , w_10157 , w_10158 , w_10159 , w_10160 , w_10161 , w_10162 , w_10163 , w_10164 , w_10165 , 
		w_10166 , w_10167 , w_10168 , w_10169 , w_10170 , w_10171 , w_10172 , w_10173 , w_10174 , w_10175 , 
		w_10176 , w_10177 , w_10178 , w_10179 , w_10180 , w_10181 , w_10182 , w_10183 , w_10184 , w_10185 , 
		w_10186 , w_10187 , w_10188 , w_10189 , w_10190 , w_10191 , w_10192 , w_10193 , w_10194 , w_10195 , 
		w_10196 , w_10197 , w_10198 , w_10199 , w_10200 , w_10201 , w_10202 , w_10203 , w_10204 , w_10205 , 
		w_10206 , w_10207 , w_10208 , w_10209 , w_10210 , w_10211 , w_10212 , w_10213 , w_10214 , w_10215 , 
		w_10216 , w_10217 , w_10218 , w_10219 , w_10220 , w_10221 , w_10222 , w_10223 , w_10224 , w_10225 , 
		w_10226 , w_10227 , w_10228 , w_10229 , w_10230 , w_10231 , w_10232 , w_10233 , w_10234 , w_10235 , 
		w_10236 , w_10237 , w_10238 , w_10239 , w_10240 , w_10241 , w_10242 , w_10243 , w_10244 , w_10245 , 
		w_10246 , w_10247 , w_10248 , w_10249 , w_10250 , w_10251 , w_10252 , w_10253 , w_10254 , w_10255 , 
		w_10256 , w_10257 , w_10258 , w_10259 , w_10260 , w_10261 , w_10262 , w_10263 , w_10264 , w_10265 , 
		w_10266 , w_10267 , w_10268 , w_10269 , w_10270 , w_10271 , w_10272 , w_10273 , w_10274 , w_10275 , 
		w_10276 , w_10277 , w_10278 , w_10279 , w_10280 , w_10281 , w_10282 , w_10283 , w_10284 , w_10285 , 
		w_10286 , w_10287 , w_10288 , w_10289 , w_10290 , w_10291 , w_10292 , w_10293 , w_10294 , w_10295 , 
		w_10296 , w_10297 , w_10298 , w_10299 , w_10300 , w_10301 , w_10302 , w_10303 , w_10304 , w_10305 , 
		w_10306 , w_10307 , w_10308 , w_10309 , w_10310 , w_10311 , w_10312 , w_10313 , w_10314 , w_10315 , 
		w_10316 , w_10317 , w_10318 , w_10319 , w_10320 , w_10321 , w_10322 , w_10323 , w_10324 , w_10325 , 
		w_10326 , w_10327 , w_10328 , w_10329 , w_10330 , w_10331 , w_10332 , w_10333 , w_10334 , w_10335 , 
		w_10336 , w_10337 , w_10338 , w_10339 , w_10340 , w_10341 , w_10342 , w_10343 , w_10344 , w_10345 , 
		w_10346 , w_10347 , w_10348 , w_10349 , w_10350 , w_10351 , w_10352 , w_10353 , w_10354 , w_10355 , 
		w_10356 , w_10357 , w_10358 , w_10359 , w_10360 , w_10361 , w_10362 , w_10363 , w_10364 , w_10365 , 
		w_10366 , w_10367 , w_10368 , w_10369 , w_10370 , w_10371 , w_10372 , w_10373 , w_10374 , w_10375 , 
		w_10376 , w_10377 , w_10378 , w_10379 , w_10380 , w_10381 , w_10382 , w_10383 , w_10384 , w_10385 , 
		w_10386 , w_10387 , w_10388 , w_10389 , w_10390 , w_10391 , w_10392 , w_10393 , w_10394 , w_10395 , 
		w_10396 , w_10397 , w_10398 , w_10399 , w_10400 , w_10401 , w_10402 , w_10403 , w_10404 , w_10405 , 
		w_10406 , w_10407 , w_10408 , w_10409 , w_10410 , w_10411 , w_10412 , w_10413 , w_10414 , w_10415 , 
		w_10416 , w_10417 , w_10418 , w_10419 , w_10420 , w_10421 , w_10422 , w_10423 , w_10424 , w_10425 , 
		w_10426 , w_10427 , w_10428 , w_10429 , w_10430 , w_10431 , w_10432 , w_10433 , w_10434 , w_10435 , 
		w_10436 , w_10437 , w_10438 , w_10439 , w_10440 , w_10441 , w_10442 , w_10443 , w_10444 , w_10445 , 
		w_10446 , w_10447 , w_10448 , w_10449 , w_10450 , w_10451 , w_10452 , w_10453 , w_10454 , w_10455 , 
		w_10456 , w_10457 , w_10458 , w_10459 , w_10460 , w_10461 , w_10462 , w_10463 , w_10464 , w_10465 , 
		w_10466 , w_10467 , w_10468 , w_10469 , w_10470 , w_10471 , w_10472 , w_10473 , w_10474 , w_10475 , 
		w_10476 , w_10477 , w_10478 , w_10479 , w_10480 , w_10481 , w_10482 , w_10483 , w_10484 , w_10485 , 
		w_10486 , w_10487 , w_10488 , w_10489 , w_10490 , w_10491 , w_10492 , w_10493 , w_10494 , w_10495 , 
		w_10496 , w_10497 , w_10498 , w_10499 , w_10500 , w_10501 , w_10502 , w_10503 , w_10504 , w_10505 , 
		w_10506 , w_10507 , w_10508 , w_10509 , w_10510 , w_10511 , w_10512 , w_10513 , w_10514 , w_10515 , 
		w_10516 , w_10517 , w_10518 , w_10519 , w_10520 , w_10521 , w_10522 , w_10523 , w_10524 , w_10525 , 
		w_10526 , w_10527 , w_10528 , w_10529 , w_10530 , w_10531 , w_10532 , w_10533 , w_10534 , w_10535 , 
		w_10536 , w_10537 , w_10538 , w_10539 , w_10540 , w_10541 , w_10542 , w_10543 , w_10544 , w_10545 , 
		w_10546 , w_10547 , w_10548 , w_10549 , w_10550 , w_10551 , w_10552 , w_10553 , w_10554 , w_10555 , 
		w_10556 , w_10557 , w_10558 , w_10559 , w_10560 , w_10561 , w_10562 , w_10563 , w_10564 , w_10565 , 
		w_10566 , w_10567 , w_10568 , w_10569 , w_10570 , w_10571 , w_10572 , w_10573 , w_10574 , w_10575 , 
		w_10576 , w_10577 , w_10578 , w_10579 , w_10580 , w_10581 , w_10582 , w_10583 , w_10584 , w_10585 , 
		w_10586 , w_10587 , w_10588 , w_10589 , w_10590 , w_10591 , w_10592 , w_10593 , w_10594 , w_10595 , 
		w_10596 , w_10597 , w_10598 , w_10599 , w_10600 , w_10601 , w_10602 , w_10603 , w_10604 , w_10605 , 
		w_10606 , w_10607 , w_10608 , w_10609 , w_10610 , w_10611 , w_10612 , w_10613 , w_10614 , w_10615 , 
		w_10616 , w_10617 , w_10618 , w_10619 , w_10620 , w_10621 , w_10622 , w_10623 , w_10624 , w_10625 , 
		w_10626 , w_10627 , w_10628 , w_10629 , w_10630 , w_10631 , w_10632 , w_10633 , w_10634 , w_10635 , 
		w_10636 , w_10637 , w_10638 , w_10639 , w_10640 , w_10641 , w_10642 , w_10643 , w_10644 , w_10645 , 
		w_10646 , w_10647 , w_10648 , w_10649 , w_10650 , w_10651 , w_10652 , w_10653 , w_10654 , w_10655 , 
		w_10656 , w_10657 , w_10658 , w_10659 , w_10660 , w_10661 , w_10662 , w_10663 , w_10664 , w_10665 , 
		w_10666 , w_10667 , w_10668 , w_10669 , w_10670 , w_10671 , w_10672 , w_10673 , w_10674 , w_10675 , 
		w_10676 , w_10677 , w_10678 , w_10679 , w_10680 , w_10681 , w_10682 , w_10683 , w_10684 , w_10685 , 
		w_10686 , w_10687 , w_10688 , w_10689 , w_10690 , w_10691 , w_10692 , w_10693 , w_10694 , w_10695 , 
		w_10696 , w_10697 , w_10698 , w_10699 , w_10700 , w_10701 , w_10702 , w_10703 , w_10704 , w_10705 , 
		w_10706 , w_10707 , w_10708 , w_10709 , w_10710 , w_10711 , w_10712 , w_10713 , w_10714 , w_10715 , 
		w_10716 , w_10717 , w_10718 , w_10719 , w_10720 , w_10721 , w_10722 , w_10723 , w_10724 , w_10725 , 
		w_10726 , w_10727 , w_10728 , w_10729 , w_10730 , w_10731 , w_10732 , w_10733 , w_10734 , w_10735 , 
		w_10736 , w_10737 , w_10738 , w_10739 , w_10740 , w_10741 , w_10742 , w_10743 , w_10744 , w_10745 , 
		w_10746 , w_10747 , w_10748 , w_10749 , w_10750 , w_10751 , w_10752 , w_10753 , w_10754 , w_10755 , 
		w_10756 , w_10757 , w_10758 , w_10759 , w_10760 , w_10761 , w_10762 , w_10763 , w_10764 , w_10765 , 
		w_10766 , w_10767 , w_10768 , w_10769 , w_10770 , w_10771 , w_10772 , w_10773 , w_10774 , w_10775 , 
		w_10776 , w_10777 , w_10778 , w_10779 , w_10780 , w_10781 , w_10782 , w_10783 , w_10784 , w_10785 , 
		w_10786 , w_10787 , w_10788 , w_10789 , w_10790 , w_10791 , w_10792 , w_10793 , w_10794 , w_10795 , 
		w_10796 , w_10797 , w_10798 , w_10799 , w_10800 , w_10801 , w_10802 , w_10803 , w_10804 , w_10805 , 
		w_10806 , w_10807 , w_10808 , w_10809 , w_10810 , w_10811 , w_10812 , w_10813 , w_10814 , w_10815 , 
		w_10816 , w_10817 , w_10818 , w_10819 , w_10820 , w_10821 , w_10822 , w_10823 , w_10824 , w_10825 , 
		w_10826 , w_10827 , w_10828 , w_10829 , w_10830 , w_10831 , w_10832 , w_10833 , w_10834 , w_10835 , 
		w_10836 , w_10837 , w_10838 , w_10839 , w_10840 , w_10841 , w_10842 , w_10843 , w_10844 , w_10845 , 
		w_10846 , w_10847 , w_10848 , w_10849 , w_10850 , w_10851 , w_10852 , w_10853 , w_10854 , w_10855 , 
		w_10856 , w_10857 , w_10858 , w_10859 , w_10860 , w_10861 , w_10862 , w_10863 , w_10864 , w_10865 , 
		w_10866 , w_10867 , w_10868 , w_10869 , w_10870 , w_10871 , w_10872 , w_10873 , w_10874 , w_10875 , 
		w_10876 , w_10877 , w_10878 , w_10879 , w_10880 , w_10881 , w_10882 , w_10883 , w_10884 , w_10885 , 
		w_10886 , w_10887 ;
buf ( \o[31]_b1 , \3927_Z[31]_b1 );
buf ( \o[31]_b0 , \3927_Z[31]_b0 );
buf ( \o[30]_b1 , \3929_Z[30]_b1 );
buf ( \o[30]_b0 , \3929_Z[30]_b0 );
buf ( \o[29]_b1 , \3931_Z[29]_b1 );
buf ( \o[29]_b0 , \3931_Z[29]_b0 );
buf ( \o[28]_b1 , \3933_Z[28]_b1 );
buf ( \o[28]_b0 , \3933_Z[28]_b0 );
buf ( \o[27]_b1 , \3935_Z[27]_b1 );
buf ( \o[27]_b0 , \3935_Z[27]_b0 );
buf ( \o[26]_b1 , \3937_Z[26]_b1 );
buf ( \o[26]_b0 , \3937_Z[26]_b0 );
buf ( \o[25]_b1 , \3939_Z[25]_b1 );
buf ( \o[25]_b0 , \3939_Z[25]_b0 );
buf ( \o[24]_b1 , \3941_Z[24]_b1 );
buf ( \o[24]_b0 , \3941_Z[24]_b0 );
buf ( \o[23]_b1 , \3943_Z[23]_b1 );
buf ( \o[23]_b0 , \3943_Z[23]_b0 );
buf ( \o[22]_b1 , \3945_Z[22]_b1 );
buf ( \o[22]_b0 , \3945_Z[22]_b0 );
buf ( \o[21]_b1 , \3947_Z[21]_b1 );
buf ( \o[21]_b0 , \3947_Z[21]_b0 );
buf ( \o[20]_b1 , \3949_Z[20]_b1 );
buf ( \o[20]_b0 , \3949_Z[20]_b0 );
buf ( \o[19]_b1 , \3951_Z[19]_b1 );
buf ( \o[19]_b0 , \3951_Z[19]_b0 );
buf ( \o[18]_b1 , \3953_Z[18]_b1 );
buf ( \o[18]_b0 , \3953_Z[18]_b0 );
buf ( \o[17]_b1 , \3955_Z[17]_b1 );
buf ( \o[17]_b0 , \3955_Z[17]_b0 );
buf ( \o[16]_b1 , \3957_Z[16]_b1 );
buf ( \o[16]_b0 , \3957_Z[16]_b0 );
buf ( \o[15]_b1 , \3959_Z[15]_b1 );
buf ( \o[15]_b0 , \3959_Z[15]_b0 );
buf ( \o[14]_b1 , \3961_Z[14]_b1 );
buf ( \o[14]_b0 , \3961_Z[14]_b0 );
buf ( \o[13]_b1 , \3963_Z[13]_b1 );
buf ( \o[13]_b0 , \3963_Z[13]_b0 );
buf ( \o[12]_b1 , \3965_Z[12]_b1 );
buf ( \o[12]_b0 , \3965_Z[12]_b0 );
buf ( \o[11]_b1 , \3967_Z[11]_b1 );
buf ( \o[11]_b0 , \3967_Z[11]_b0 );
buf ( \o[10]_b1 , \3969_Z[10]_b1 );
buf ( \o[10]_b0 , \3969_Z[10]_b0 );
buf ( \o[9]_b1 , \3971_Z[9]_b1 );
buf ( \o[9]_b0 , \3971_Z[9]_b0 );
buf ( \o[8]_b1 , \3973_Z[8]_b1 );
buf ( \o[8]_b0 , \3973_Z[8]_b0 );
buf ( \o[7]_b1 , \3975_Z[7]_b1 );
buf ( \o[7]_b0 , \3975_Z[7]_b0 );
buf ( \o[6]_b1 , \3977_Z[6]_b1 );
buf ( \o[6]_b0 , \3977_Z[6]_b0 );
buf ( \o[5]_b1 , \3979_Z[5]_b1 );
buf ( \o[5]_b0 , \3979_Z[5]_b0 );
buf ( \o[4]_b1 , \3981_Z[4]_b1 );
buf ( \o[4]_b0 , \3981_Z[4]_b0 );
buf ( \o[3]_b1 , \3983_Z[3]_b1 );
buf ( \o[3]_b0 , \3983_Z[3]_b0 );
buf ( \o[2]_b1 , \3985_Z[2]_b1 );
buf ( \o[2]_b0 , \3985_Z[2]_b0 );
buf ( \o[1]_b1 , \3987_Z[1]_b1 );
buf ( \o[1]_b0 , \3987_Z[1]_b0 );
buf ( \o[0]_b1 , \3989_Z[0]_b1 );
buf ( \o[0]_b0 , \3989_Z[0]_b0 );
and ( \205_n5[0]_b1 , 1'b0_b1 , w_0 );
xor ( w_0 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1 );
and ( \205_n5[0]_b0 , w_1 , 1'b1_b0 );
or ( \206_b1 , \b[0]_b1 , w_2 );
or ( \206_b0 , \b[0]_b0 , \205_n5[0]_b0 );
not ( \205_n5[0]_b0 , w_3 );
and ( w_3 , w_2 , \205_n5[0]_b1 );
buf ( \207_A[0]_b1 , \c[0]_b1 );
buf ( \207_A[0]_b0 , \c[0]_b0 );
buf ( \208_B[0]_b1 , \d[0]_b1 );
buf ( \208_B[0]_b0 , \d[0]_b0 );
or ( \209_b1 , \207_A[0]_b1 , \208_B[0]_b1 );
xor ( \209_b0 , \207_A[0]_b0 , w_4 );
not ( w_4 , w_5 );
and ( w_5 , \208_B[0]_b1 , \208_B[0]_b0 );
buf ( \210_SUM[0]_b1 , \209_b1 );
buf ( \210_SUM[0]_b0 , \209_b0 );
or ( \211_b1 , \a[31]_b1 , \a[30]_b1 );
xor ( \211_b0 , \a[31]_b0 , w_6 );
not ( w_6 , w_7 );
and ( w_7 , \a[30]_b1 , \a[30]_b0 );
or ( \212_b1 , \a[29]_b1 , \a[28]_b1 );
xor ( \212_b0 , \a[29]_b0 , w_8 );
not ( w_8 , w_9 );
and ( w_9 , \a[28]_b1 , \a[28]_b0 );
or ( \213_b1 , \211_b1 , \212_b1 );
xor ( \213_b0 , \211_b0 , w_10 );
not ( w_10 , w_11 );
and ( w_11 , \212_b1 , \212_b0 );
or ( \214_b1 , \a[27]_b1 , \a[26]_b1 );
xor ( \214_b0 , \a[27]_b0 , w_12 );
not ( w_12 , w_13 );
and ( w_13 , \a[26]_b1 , \a[26]_b0 );
or ( \215_b1 , \a[25]_b1 , \a[24]_b1 );
xor ( \215_b0 , \a[25]_b0 , w_14 );
not ( w_14 , w_15 );
and ( w_15 , \a[24]_b1 , \a[24]_b0 );
or ( \216_b1 , \214_b1 , \215_b1 );
xor ( \216_b0 , \214_b0 , w_16 );
not ( w_16 , w_17 );
and ( w_17 , \215_b1 , \215_b0 );
or ( \217_b1 , \213_b1 , \216_b1 );
xor ( \217_b0 , \213_b0 , w_18 );
not ( w_18 , w_19 );
and ( w_19 , \216_b1 , \216_b0 );
or ( \218_b1 , \a[23]_b1 , \a[22]_b1 );
xor ( \218_b0 , \a[23]_b0 , w_20 );
not ( w_20 , w_21 );
and ( w_21 , \a[22]_b1 , \a[22]_b0 );
or ( \219_b1 , \a[21]_b1 , \a[20]_b1 );
xor ( \219_b0 , \a[21]_b0 , w_22 );
not ( w_22 , w_23 );
and ( w_23 , \a[20]_b1 , \a[20]_b0 );
or ( \220_b1 , \218_b1 , \219_b1 );
xor ( \220_b0 , \218_b0 , w_24 );
not ( w_24 , w_25 );
and ( w_25 , \219_b1 , \219_b0 );
or ( \221_b1 , \a[19]_b1 , \a[18]_b1 );
xor ( \221_b0 , \a[19]_b0 , w_26 );
not ( w_26 , w_27 );
and ( w_27 , \a[18]_b1 , \a[18]_b0 );
or ( \222_b1 , \a[17]_b1 , \a[16]_b1 );
xor ( \222_b0 , \a[17]_b0 , w_28 );
not ( w_28 , w_29 );
and ( w_29 , \a[16]_b1 , \a[16]_b0 );
or ( \223_b1 , \221_b1 , \222_b1 );
xor ( \223_b0 , \221_b0 , w_30 );
not ( w_30 , w_31 );
and ( w_31 , \222_b1 , \222_b0 );
or ( \224_b1 , \220_b1 , \223_b1 );
xor ( \224_b0 , \220_b0 , w_32 );
not ( w_32 , w_33 );
and ( w_33 , \223_b1 , \223_b0 );
or ( \225_b1 , \217_b1 , \224_b1 );
xor ( \225_b0 , \217_b0 , w_34 );
not ( w_34 , w_35 );
and ( w_35 , \224_b1 , \224_b0 );
or ( \226_b1 , \a[15]_b1 , \a[14]_b1 );
xor ( \226_b0 , \a[15]_b0 , w_36 );
not ( w_36 , w_37 );
and ( w_37 , \a[14]_b1 , \a[14]_b0 );
or ( \227_b1 , \a[13]_b1 , \a[12]_b1 );
xor ( \227_b0 , \a[13]_b0 , w_38 );
not ( w_38 , w_39 );
and ( w_39 , \a[12]_b1 , \a[12]_b0 );
or ( \228_b1 , \226_b1 , \227_b1 );
xor ( \228_b0 , \226_b0 , w_40 );
not ( w_40 , w_41 );
and ( w_41 , \227_b1 , \227_b0 );
or ( \229_b1 , \a[11]_b1 , \a[10]_b1 );
xor ( \229_b0 , \a[11]_b0 , w_42 );
not ( w_42 , w_43 );
and ( w_43 , \a[10]_b1 , \a[10]_b0 );
or ( \230_b1 , \a[9]_b1 , \a[8]_b1 );
xor ( \230_b0 , \a[9]_b0 , w_44 );
not ( w_44 , w_45 );
and ( w_45 , \a[8]_b1 , \a[8]_b0 );
or ( \231_b1 , \229_b1 , \230_b1 );
xor ( \231_b0 , \229_b0 , w_46 );
not ( w_46 , w_47 );
and ( w_47 , \230_b1 , \230_b0 );
or ( \232_b1 , \228_b1 , \231_b1 );
xor ( \232_b0 , \228_b0 , w_48 );
not ( w_48 , w_49 );
and ( w_49 , \231_b1 , \231_b0 );
or ( \233_b1 , \a[7]_b1 , \a[6]_b1 );
xor ( \233_b0 , \a[7]_b0 , w_50 );
not ( w_50 , w_51 );
and ( w_51 , \a[6]_b1 , \a[6]_b0 );
or ( \234_b1 , \a[5]_b1 , \a[4]_b1 );
xor ( \234_b0 , \a[5]_b0 , w_52 );
not ( w_52 , w_53 );
and ( w_53 , \a[4]_b1 , \a[4]_b0 );
or ( \235_b1 , \233_b1 , \234_b1 );
xor ( \235_b0 , \233_b0 , w_54 );
not ( w_54 , w_55 );
and ( w_55 , \234_b1 , \234_b0 );
or ( \236_b1 , \a[3]_b1 , \a[2]_b1 );
xor ( \236_b0 , \a[3]_b0 , w_56 );
not ( w_56 , w_57 );
and ( w_57 , \a[2]_b1 , \a[2]_b0 );
or ( \237_b1 , \a[1]_b1 , \a[0]_b1 );
xor ( \237_b0 , \a[1]_b0 , w_58 );
not ( w_58 , w_59 );
and ( w_59 , \a[0]_b1 , \a[0]_b0 );
or ( \238_b1 , \236_b1 , \237_b1 );
xor ( \238_b0 , \236_b0 , w_60 );
not ( w_60 , w_61 );
and ( w_61 , \237_b1 , \237_b0 );
or ( \239_b1 , \235_b1 , \238_b1 );
xor ( \239_b0 , \235_b0 , w_62 );
not ( w_62 , w_63 );
and ( w_63 , \238_b1 , \238_b0 );
or ( \240_b1 , \232_b1 , \239_b1 );
xor ( \240_b0 , \232_b0 , w_64 );
not ( w_64 , w_65 );
and ( w_65 , \239_b1 , \239_b0 );
or ( \241_b1 , \225_b1 , \240_b1 );
xor ( \241_b0 , \225_b0 , w_66 );
not ( w_66 , w_67 );
and ( w_67 , \240_b1 , \240_b0 );
and ( \242_b0 , \210_SUM[0]_b0 , w_68 );
and ( \242_b0 , \206_b0 , w_69 );
and ( w_82 , w_83 , w_70 );
and ( w_70 , \206_b0 , w_71 );
and ( w_83 , \206_b1 , w_72 );
and ( \242_b1 , \210_SUM[0]_b0 , w_73 );
and ( \210_SUM[0]_b1 , w_84 , w_74 );
and ( w_83 , \206_b0 , w_75 );
and ( \242_b1 , \242_b0 , w_76 );
and ( w_81 , w_85 , \241_b1 );
or ( w_68 , w_69 , w_77 );
or ( w_77 , w_71 , \241_b0 );
or ( w_72 , w_73 , w_78 );
or ( w_78 , w_74 , w_79 );
or ( w_79 , w_75 , w_80 );
or ( w_80 , w_76 , w_81 );
not ( \210_SUM[0]_b1 , w_82 );
not ( \210_SUM[0]_b0 , w_83 );
not ( \242_b1 , w_84 );
not ( \241_b0 , w_85 );
buf ( \243_A[0]_b1 , \c[0]_b1 );
buf ( \243_A[0]_b0 , \c[0]_b0 );
buf ( \244_B[0]_b1 , \d[0]_b1 );
buf ( \244_B[0]_b0 , \d[0]_b0 );
or ( \245_b1 , \243_A[0]_b1 , \244_B[0]_b1 );
xor ( \245_b0 , \243_A[0]_b0 , w_86 );
not ( w_86 , w_87 );
and ( w_87 , \244_B[0]_b1 , \244_B[0]_b0 );
buf ( \246_SUM[0]_b1 , \245_b1 );
buf ( \246_SUM[0]_b0 , \245_b0 );
or ( \247_b1 , \s[31]_b1 , \s[30]_b1 );
xor ( \247_b0 , \s[31]_b0 , w_88 );
not ( w_88 , w_89 );
and ( w_89 , \s[30]_b1 , \s[30]_b0 );
or ( \248_b1 , \s[29]_b1 , \s[28]_b1 );
xor ( \248_b0 , \s[29]_b0 , w_90 );
not ( w_90 , w_91 );
and ( w_91 , \s[28]_b1 , \s[28]_b0 );
or ( \249_b1 , \247_b1 , \248_b1 );
xor ( \249_b0 , \247_b0 , w_92 );
not ( w_92 , w_93 );
and ( w_93 , \248_b1 , \248_b0 );
or ( \250_b1 , \s[27]_b1 , \s[26]_b1 );
xor ( \250_b0 , \s[27]_b0 , w_94 );
not ( w_94 , w_95 );
and ( w_95 , \s[26]_b1 , \s[26]_b0 );
or ( \251_b1 , \s[25]_b1 , \s[24]_b1 );
xor ( \251_b0 , \s[25]_b0 , w_96 );
not ( w_96 , w_97 );
and ( w_97 , \s[24]_b1 , \s[24]_b0 );
or ( \252_b1 , \250_b1 , \251_b1 );
xor ( \252_b0 , \250_b0 , w_98 );
not ( w_98 , w_99 );
and ( w_99 , \251_b1 , \251_b0 );
or ( \253_b1 , \249_b1 , \252_b1 );
xor ( \253_b0 , \249_b0 , w_100 );
not ( w_100 , w_101 );
and ( w_101 , \252_b1 , \252_b0 );
or ( \254_b1 , \s[23]_b1 , \s[22]_b1 );
xor ( \254_b0 , \s[23]_b0 , w_102 );
not ( w_102 , w_103 );
and ( w_103 , \s[22]_b1 , \s[22]_b0 );
or ( \255_b1 , \s[21]_b1 , \s[20]_b1 );
xor ( \255_b0 , \s[21]_b0 , w_104 );
not ( w_104 , w_105 );
and ( w_105 , \s[20]_b1 , \s[20]_b0 );
or ( \256_b1 , \254_b1 , \255_b1 );
xor ( \256_b0 , \254_b0 , w_106 );
not ( w_106 , w_107 );
and ( w_107 , \255_b1 , \255_b0 );
or ( \257_b1 , \s[19]_b1 , \s[18]_b1 );
xor ( \257_b0 , \s[19]_b0 , w_108 );
not ( w_108 , w_109 );
and ( w_109 , \s[18]_b1 , \s[18]_b0 );
or ( \258_b1 , \s[17]_b1 , \s[16]_b1 );
xor ( \258_b0 , \s[17]_b0 , w_110 );
not ( w_110 , w_111 );
and ( w_111 , \s[16]_b1 , \s[16]_b0 );
or ( \259_b1 , \257_b1 , \258_b1 );
xor ( \259_b0 , \257_b0 , w_112 );
not ( w_112 , w_113 );
and ( w_113 , \258_b1 , \258_b0 );
or ( \260_b1 , \256_b1 , \259_b1 );
xor ( \260_b0 , \256_b0 , w_114 );
not ( w_114 , w_115 );
and ( w_115 , \259_b1 , \259_b0 );
or ( \261_b1 , \253_b1 , \260_b1 );
xor ( \261_b0 , \253_b0 , w_116 );
not ( w_116 , w_117 );
and ( w_117 , \260_b1 , \260_b0 );
or ( \262_b1 , \s[15]_b1 , \s[14]_b1 );
xor ( \262_b0 , \s[15]_b0 , w_118 );
not ( w_118 , w_119 );
and ( w_119 , \s[14]_b1 , \s[14]_b0 );
or ( \263_b1 , \s[13]_b1 , \s[12]_b1 );
xor ( \263_b0 , \s[13]_b0 , w_120 );
not ( w_120 , w_121 );
and ( w_121 , \s[12]_b1 , \s[12]_b0 );
or ( \264_b1 , \262_b1 , \263_b1 );
xor ( \264_b0 , \262_b0 , w_122 );
not ( w_122 , w_123 );
and ( w_123 , \263_b1 , \263_b0 );
or ( \265_b1 , \s[11]_b1 , \s[10]_b1 );
xor ( \265_b0 , \s[11]_b0 , w_124 );
not ( w_124 , w_125 );
and ( w_125 , \s[10]_b1 , \s[10]_b0 );
or ( \266_b1 , \s[9]_b1 , \s[8]_b1 );
xor ( \266_b0 , \s[9]_b0 , w_126 );
not ( w_126 , w_127 );
and ( w_127 , \s[8]_b1 , \s[8]_b0 );
or ( \267_b1 , \265_b1 , \266_b1 );
xor ( \267_b0 , \265_b0 , w_128 );
not ( w_128 , w_129 );
and ( w_129 , \266_b1 , \266_b0 );
or ( \268_b1 , \264_b1 , \267_b1 );
xor ( \268_b0 , \264_b0 , w_130 );
not ( w_130 , w_131 );
and ( w_131 , \267_b1 , \267_b0 );
or ( \269_b1 , \s[7]_b1 , \s[6]_b1 );
xor ( \269_b0 , \s[7]_b0 , w_132 );
not ( w_132 , w_133 );
and ( w_133 , \s[6]_b1 , \s[6]_b0 );
or ( \270_b1 , \s[5]_b1 , \s[4]_b1 );
xor ( \270_b0 , \s[5]_b0 , w_134 );
not ( w_134 , w_135 );
and ( w_135 , \s[4]_b1 , \s[4]_b0 );
or ( \271_b1 , \269_b1 , \270_b1 );
xor ( \271_b0 , \269_b0 , w_136 );
not ( w_136 , w_137 );
and ( w_137 , \270_b1 , \270_b0 );
or ( \272_b1 , \s[3]_b1 , \s[2]_b1 );
xor ( \272_b0 , \s[3]_b0 , w_138 );
not ( w_138 , w_139 );
and ( w_139 , \s[2]_b1 , \s[2]_b0 );
or ( \273_b1 , \s[1]_b1 , \s[0]_b1 );
xor ( \273_b0 , \s[1]_b0 , w_140 );
not ( w_140 , w_141 );
and ( w_141 , \s[0]_b1 , \s[0]_b0 );
or ( \274_b1 , \272_b1 , \273_b1 );
xor ( \274_b0 , \272_b0 , w_142 );
not ( w_142 , w_143 );
and ( w_143 , \273_b1 , \273_b0 );
or ( \275_b1 , \271_b1 , \274_b1 );
xor ( \275_b0 , \271_b0 , w_144 );
not ( w_144 , w_145 );
and ( w_145 , \274_b1 , \274_b0 );
or ( \276_b1 , \268_b1 , \275_b1 );
xor ( \276_b0 , \268_b0 , w_146 );
not ( w_146 , w_147 );
and ( w_147 , \275_b1 , \275_b0 );
or ( \277_b1 , \261_b1 , \276_b1 );
xor ( \277_b0 , \261_b0 , w_148 );
not ( w_148 , w_149 );
and ( w_149 , \276_b1 , \276_b0 );
and ( \278_b0 , \246_SUM[0]_b0 , w_150 );
and ( \278_b0 , \242_b0 , w_151 );
and ( w_164 , w_165 , w_152 );
and ( w_152 , \242_b0 , w_153 );
and ( w_165 , \242_b1 , w_154 );
and ( \278_b1 , \246_SUM[0]_b0 , w_155 );
and ( \246_SUM[0]_b1 , w_166 , w_156 );
and ( w_165 , \242_b0 , w_157 );
and ( \278_b1 , \278_b0 , w_158 );
and ( w_163 , w_167 , \277_b1 );
or ( w_150 , w_151 , w_159 );
or ( w_159 , w_153 , \277_b0 );
or ( w_154 , w_155 , w_160 );
or ( w_160 , w_156 , w_161 );
or ( w_161 , w_157 , w_162 );
or ( w_162 , w_158 , w_163 );
not ( \246_SUM[0]_b1 , w_164 );
not ( \246_SUM[0]_b0 , w_165 );
not ( \278_b1 , w_166 );
not ( \277_b0 , w_167 );
and ( \279_n5[1]_b1 , 1'b0_b1 , w_168 );
xor ( w_168 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_169 );
and ( \279_n5[1]_b0 , w_169 , 1'b1_b0 );
or ( \280_b1 , \b[1]_b1 , w_170 );
or ( \280_b0 , \b[1]_b0 , \279_n5[1]_b0 );
not ( \279_n5[1]_b0 , w_171 );
and ( w_171 , w_170 , \279_n5[1]_b1 );
buf ( \281_A[1]_b1 , \c[1]_b1 );
buf ( \281_A[1]_b0 , \c[1]_b0 );
buf ( \282_B[1]_b1 , \d[1]_b1 );
buf ( \282_B[1]_b0 , \d[1]_b0 );
buf ( \283_b1 , \282_B[1]_b1 );
not ( \283_b1 , w_172 );
not ( \283_b0 , w_173 );
and ( w_172 , w_173 , \282_B[1]_b0 );
or ( \284_b1 , \281_A[1]_b1 , \283_b1 );
xor ( \284_b0 , \281_A[1]_b0 , w_174 );
not ( w_174 , w_175 );
and ( w_175 , \283_b1 , \283_b0 );
buf ( \285_b1 , \208_B[0]_b1 );
not ( \285_b1 , w_176 );
not ( \285_b0 , w_177 );
and ( w_176 , w_177 , \208_B[0]_b0 );
or ( \286_b1 , \207_A[0]_b1 , w_178 );
or ( \286_b0 , \207_A[0]_b0 , \285_b0 );
not ( \285_b0 , w_179 );
and ( w_179 , w_178 , \285_b1 );
or ( \287_b1 , \284_b1 , \286_b1 );
xor ( \287_b0 , \284_b0 , w_180 );
not ( w_180 , w_181 );
and ( w_181 , \286_b1 , \286_b0 );
buf ( \288_SUM[1]_b1 , \287_b1 );
buf ( \288_SUM[1]_b0 , \287_b0 );
and ( \289_b0 , \288_SUM[1]_b0 , w_182 );
and ( \289_b0 , \280_b0 , w_183 );
and ( w_196 , w_197 , w_184 );
and ( w_184 , \280_b0 , w_185 );
and ( w_197 , \280_b1 , w_186 );
and ( \289_b1 , \288_SUM[1]_b0 , w_187 );
and ( \288_SUM[1]_b1 , w_198 , w_188 );
and ( w_197 , \280_b0 , w_189 );
and ( \289_b1 , \289_b0 , w_190 );
and ( w_195 , w_199 , \241_b1 );
or ( w_182 , w_183 , w_191 );
or ( w_191 , w_185 , \241_b0 );
or ( w_186 , w_187 , w_192 );
or ( w_192 , w_188 , w_193 );
or ( w_193 , w_189 , w_194 );
or ( w_194 , w_190 , w_195 );
not ( \288_SUM[1]_b1 , w_196 );
not ( \288_SUM[1]_b0 , w_197 );
not ( \289_b1 , w_198 );
not ( \241_b0 , w_199 );
buf ( \290_A[1]_b1 , \c[1]_b1 );
buf ( \290_A[1]_b0 , \c[1]_b0 );
buf ( \291_B[1]_b1 , \d[1]_b1 );
buf ( \291_B[1]_b0 , \d[1]_b0 );
or ( \292_b1 , \290_A[1]_b1 , \291_B[1]_b1 );
xor ( \292_b0 , \290_A[1]_b0 , w_200 );
not ( w_200 , w_201 );
and ( w_201 , \291_B[1]_b1 , \291_B[1]_b0 );
or ( \293_b1 , \243_A[0]_b1 , \244_B[0]_b1 );
not ( \244_B[0]_b1 , w_202 );
and ( \293_b0 , \243_A[0]_b0 , w_203 );
and ( w_202 , w_203 , \244_B[0]_b0 );
or ( \294_b1 , \292_b1 , \293_b1 );
xor ( \294_b0 , \292_b0 , w_204 );
not ( w_204 , w_205 );
and ( w_205 , \293_b1 , \293_b0 );
buf ( \295_SUM[1]_b1 , \294_b1 );
buf ( \295_SUM[1]_b0 , \294_b0 );
and ( \296_b0 , \295_SUM[1]_b0 , w_206 );
and ( \296_b0 , \289_b0 , w_207 );
and ( w_220 , w_221 , w_208 );
and ( w_208 , \289_b0 , w_209 );
and ( w_221 , \289_b1 , w_210 );
and ( \296_b1 , \295_SUM[1]_b0 , w_211 );
and ( \295_SUM[1]_b1 , w_222 , w_212 );
and ( w_221 , \289_b0 , w_213 );
and ( \296_b1 , \296_b0 , w_214 );
and ( w_219 , w_223 , \277_b1 );
or ( w_206 , w_207 , w_215 );
or ( w_215 , w_209 , \277_b0 );
or ( w_210 , w_211 , w_216 );
or ( w_216 , w_212 , w_217 );
or ( w_217 , w_213 , w_218 );
or ( w_218 , w_214 , w_219 );
not ( \295_SUM[1]_b1 , w_220 );
not ( \295_SUM[1]_b0 , w_221 );
not ( \296_b1 , w_222 );
not ( \277_b0 , w_223 );
and ( \297_n5[2]_b1 , 1'b0_b1 , w_224 );
xor ( w_224 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_225 );
and ( \297_n5[2]_b0 , w_225 , 1'b1_b0 );
or ( \298_b1 , \b[2]_b1 , w_226 );
or ( \298_b0 , \b[2]_b0 , \297_n5[2]_b0 );
not ( \297_n5[2]_b0 , w_227 );
and ( w_227 , w_226 , \297_n5[2]_b1 );
buf ( \299_A[2]_b1 , \c[2]_b1 );
buf ( \299_A[2]_b0 , \c[2]_b0 );
buf ( \300_B[2]_b1 , \d[2]_b1 );
buf ( \300_B[2]_b0 , \d[2]_b0 );
buf ( \301_b1 , \300_B[2]_b1 );
not ( \301_b1 , w_228 );
not ( \301_b0 , w_229 );
and ( w_228 , w_229 , \300_B[2]_b0 );
or ( \302_b1 , \299_A[2]_b1 , \301_b1 );
xor ( \302_b0 , \299_A[2]_b0 , w_230 );
not ( w_230 , w_231 );
and ( w_231 , \301_b1 , \301_b0 );
or ( \303_b1 , \281_A[1]_b1 , \283_b1 );
not ( \283_b1 , w_232 );
and ( \303_b0 , \281_A[1]_b0 , w_233 );
and ( w_232 , w_233 , \283_b0 );
or ( \304_b1 , \283_b1 , \286_b1 );
not ( \286_b1 , w_234 );
and ( \304_b0 , \283_b0 , w_235 );
and ( w_234 , w_235 , \286_b0 );
or ( \305_b1 , \281_A[1]_b1 , \286_b1 );
not ( \286_b1 , w_236 );
and ( \305_b0 , \281_A[1]_b0 , w_237 );
and ( w_236 , w_237 , \286_b0 );
or ( \307_b1 , \302_b1 , \306_b1 );
xor ( \307_b0 , \302_b0 , w_238 );
not ( w_238 , w_239 );
and ( w_239 , \306_b1 , \306_b0 );
buf ( \308_SUM[2]_b1 , \307_b1 );
buf ( \308_SUM[2]_b0 , \307_b0 );
and ( \309_b0 , \308_SUM[2]_b0 , w_240 );
and ( \309_b0 , \298_b0 , w_241 );
and ( w_254 , w_255 , w_242 );
and ( w_242 , \298_b0 , w_243 );
and ( w_255 , \298_b1 , w_244 );
and ( \309_b1 , \308_SUM[2]_b0 , w_245 );
and ( \308_SUM[2]_b1 , w_256 , w_246 );
and ( w_255 , \298_b0 , w_247 );
and ( \309_b1 , \309_b0 , w_248 );
and ( w_253 , w_257 , \241_b1 );
or ( w_240 , w_241 , w_249 );
or ( w_249 , w_243 , \241_b0 );
or ( w_244 , w_245 , w_250 );
or ( w_250 , w_246 , w_251 );
or ( w_251 , w_247 , w_252 );
or ( w_252 , w_248 , w_253 );
not ( \308_SUM[2]_b1 , w_254 );
not ( \308_SUM[2]_b0 , w_255 );
not ( \309_b1 , w_256 );
not ( \241_b0 , w_257 );
buf ( \310_A[2]_b1 , \c[2]_b1 );
buf ( \310_A[2]_b0 , \c[2]_b0 );
buf ( \311_B[2]_b1 , \d[2]_b1 );
buf ( \311_B[2]_b0 , \d[2]_b0 );
or ( \312_b1 , \310_A[2]_b1 , \311_B[2]_b1 );
xor ( \312_b0 , \310_A[2]_b0 , w_258 );
not ( w_258 , w_259 );
and ( w_259 , \311_B[2]_b1 , \311_B[2]_b0 );
or ( \313_b1 , \290_A[1]_b1 , \291_B[1]_b1 );
not ( \291_B[1]_b1 , w_260 );
and ( \313_b0 , \290_A[1]_b0 , w_261 );
and ( w_260 , w_261 , \291_B[1]_b0 );
or ( \314_b1 , \291_B[1]_b1 , \293_b1 );
not ( \293_b1 , w_262 );
and ( \314_b0 , \291_B[1]_b0 , w_263 );
and ( w_262 , w_263 , \293_b0 );
or ( \315_b1 , \290_A[1]_b1 , \293_b1 );
not ( \293_b1 , w_264 );
and ( \315_b0 , \290_A[1]_b0 , w_265 );
and ( w_264 , w_265 , \293_b0 );
or ( \317_b1 , \312_b1 , \316_b1 );
xor ( \317_b0 , \312_b0 , w_266 );
not ( w_266 , w_267 );
and ( w_267 , \316_b1 , \316_b0 );
buf ( \318_SUM[2]_b1 , \317_b1 );
buf ( \318_SUM[2]_b0 , \317_b0 );
and ( \319_b0 , \318_SUM[2]_b0 , w_268 );
and ( \319_b0 , \309_b0 , w_269 );
and ( w_282 , w_283 , w_270 );
and ( w_270 , \309_b0 , w_271 );
and ( w_283 , \309_b1 , w_272 );
and ( \319_b1 , \318_SUM[2]_b0 , w_273 );
and ( \318_SUM[2]_b1 , w_284 , w_274 );
and ( w_283 , \309_b0 , w_275 );
and ( \319_b1 , \319_b0 , w_276 );
and ( w_281 , w_285 , \277_b1 );
or ( w_268 , w_269 , w_277 );
or ( w_277 , w_271 , \277_b0 );
or ( w_272 , w_273 , w_278 );
or ( w_278 , w_274 , w_279 );
or ( w_279 , w_275 , w_280 );
or ( w_280 , w_276 , w_281 );
not ( \318_SUM[2]_b1 , w_282 );
not ( \318_SUM[2]_b0 , w_283 );
not ( \319_b1 , w_284 );
not ( \277_b0 , w_285 );
and ( \320_n5[3]_b1 , 1'b0_b1 , w_286 );
xor ( w_286 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_287 );
and ( \320_n5[3]_b0 , w_287 , 1'b1_b0 );
or ( \321_b1 , \b[3]_b1 , w_288 );
or ( \321_b0 , \b[3]_b0 , \320_n5[3]_b0 );
not ( \320_n5[3]_b0 , w_289 );
and ( w_289 , w_288 , \320_n5[3]_b1 );
buf ( \322_A[3]_b1 , \c[3]_b1 );
buf ( \322_A[3]_b0 , \c[3]_b0 );
buf ( \323_B[3]_b1 , \d[3]_b1 );
buf ( \323_B[3]_b0 , \d[3]_b0 );
buf ( \324_b1 , \323_B[3]_b1 );
not ( \324_b1 , w_290 );
not ( \324_b0 , w_291 );
and ( w_290 , w_291 , \323_B[3]_b0 );
or ( \325_b1 , \322_A[3]_b1 , \324_b1 );
xor ( \325_b0 , \322_A[3]_b0 , w_292 );
not ( w_292 , w_293 );
and ( w_293 , \324_b1 , \324_b0 );
or ( \326_b1 , \299_A[2]_b1 , \301_b1 );
not ( \301_b1 , w_294 );
and ( \326_b0 , \299_A[2]_b0 , w_295 );
and ( w_294 , w_295 , \301_b0 );
or ( \327_b1 , \301_b1 , \306_b1 );
not ( \306_b1 , w_296 );
and ( \327_b0 , \301_b0 , w_297 );
and ( w_296 , w_297 , \306_b0 );
or ( \328_b1 , \299_A[2]_b1 , \306_b1 );
not ( \306_b1 , w_298 );
and ( \328_b0 , \299_A[2]_b0 , w_299 );
and ( w_298 , w_299 , \306_b0 );
or ( \330_b1 , \325_b1 , \329_b1 );
xor ( \330_b0 , \325_b0 , w_300 );
not ( w_300 , w_301 );
and ( w_301 , \329_b1 , \329_b0 );
buf ( \331_SUM[3]_b1 , \330_b1 );
buf ( \331_SUM[3]_b0 , \330_b0 );
and ( \332_b0 , \331_SUM[3]_b0 , w_302 );
and ( \332_b0 , \321_b0 , w_303 );
and ( w_316 , w_317 , w_304 );
and ( w_304 , \321_b0 , w_305 );
and ( w_317 , \321_b1 , w_306 );
and ( \332_b1 , \331_SUM[3]_b0 , w_307 );
and ( \331_SUM[3]_b1 , w_318 , w_308 );
and ( w_317 , \321_b0 , w_309 );
and ( \332_b1 , \332_b0 , w_310 );
and ( w_315 , w_319 , \241_b1 );
or ( w_302 , w_303 , w_311 );
or ( w_311 , w_305 , \241_b0 );
or ( w_306 , w_307 , w_312 );
or ( w_312 , w_308 , w_313 );
or ( w_313 , w_309 , w_314 );
or ( w_314 , w_310 , w_315 );
not ( \331_SUM[3]_b1 , w_316 );
not ( \331_SUM[3]_b0 , w_317 );
not ( \332_b1 , w_318 );
not ( \241_b0 , w_319 );
buf ( \333_A[3]_b1 , \c[3]_b1 );
buf ( \333_A[3]_b0 , \c[3]_b0 );
buf ( \334_B[3]_b1 , \d[3]_b1 );
buf ( \334_B[3]_b0 , \d[3]_b0 );
or ( \335_b1 , \333_A[3]_b1 , \334_B[3]_b1 );
xor ( \335_b0 , \333_A[3]_b0 , w_320 );
not ( w_320 , w_321 );
and ( w_321 , \334_B[3]_b1 , \334_B[3]_b0 );
or ( \336_b1 , \310_A[2]_b1 , \311_B[2]_b1 );
not ( \311_B[2]_b1 , w_322 );
and ( \336_b0 , \310_A[2]_b0 , w_323 );
and ( w_322 , w_323 , \311_B[2]_b0 );
or ( \337_b1 , \311_B[2]_b1 , \316_b1 );
not ( \316_b1 , w_324 );
and ( \337_b0 , \311_B[2]_b0 , w_325 );
and ( w_324 , w_325 , \316_b0 );
or ( \338_b1 , \310_A[2]_b1 , \316_b1 );
not ( \316_b1 , w_326 );
and ( \338_b0 , \310_A[2]_b0 , w_327 );
and ( w_326 , w_327 , \316_b0 );
or ( \340_b1 , \335_b1 , \339_b1 );
xor ( \340_b0 , \335_b0 , w_328 );
not ( w_328 , w_329 );
and ( w_329 , \339_b1 , \339_b0 );
buf ( \341_SUM[3]_b1 , \340_b1 );
buf ( \341_SUM[3]_b0 , \340_b0 );
and ( \342_b0 , \341_SUM[3]_b0 , w_330 );
and ( \342_b0 , \332_b0 , w_331 );
and ( w_344 , w_345 , w_332 );
and ( w_332 , \332_b0 , w_333 );
and ( w_345 , \332_b1 , w_334 );
and ( \342_b1 , \341_SUM[3]_b0 , w_335 );
and ( \341_SUM[3]_b1 , w_346 , w_336 );
and ( w_345 , \332_b0 , w_337 );
and ( \342_b1 , \342_b0 , w_338 );
and ( w_343 , w_347 , \277_b1 );
or ( w_330 , w_331 , w_339 );
or ( w_339 , w_333 , \277_b0 );
or ( w_334 , w_335 , w_340 );
or ( w_340 , w_336 , w_341 );
or ( w_341 , w_337 , w_342 );
or ( w_342 , w_338 , w_343 );
not ( \341_SUM[3]_b1 , w_344 );
not ( \341_SUM[3]_b0 , w_345 );
not ( \342_b1 , w_346 );
not ( \277_b0 , w_347 );
and ( \343_n5[4]_b1 , 1'b0_b1 , w_348 );
xor ( w_348 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_349 );
and ( \343_n5[4]_b0 , w_349 , 1'b1_b0 );
or ( \344_b1 , \b[4]_b1 , w_350 );
or ( \344_b0 , \b[4]_b0 , \343_n5[4]_b0 );
not ( \343_n5[4]_b0 , w_351 );
and ( w_351 , w_350 , \343_n5[4]_b1 );
buf ( \345_A[4]_b1 , \c[4]_b1 );
buf ( \345_A[4]_b0 , \c[4]_b0 );
buf ( \346_B[4]_b1 , \d[4]_b1 );
buf ( \346_B[4]_b0 , \d[4]_b0 );
buf ( \347_b1 , \346_B[4]_b1 );
not ( \347_b1 , w_352 );
not ( \347_b0 , w_353 );
and ( w_352 , w_353 , \346_B[4]_b0 );
or ( \348_b1 , \345_A[4]_b1 , \347_b1 );
xor ( \348_b0 , \345_A[4]_b0 , w_354 );
not ( w_354 , w_355 );
and ( w_355 , \347_b1 , \347_b0 );
or ( \349_b1 , \322_A[3]_b1 , \324_b1 );
not ( \324_b1 , w_356 );
and ( \349_b0 , \322_A[3]_b0 , w_357 );
and ( w_356 , w_357 , \324_b0 );
or ( \350_b1 , \324_b1 , \329_b1 );
not ( \329_b1 , w_358 );
and ( \350_b0 , \324_b0 , w_359 );
and ( w_358 , w_359 , \329_b0 );
or ( \351_b1 , \322_A[3]_b1 , \329_b1 );
not ( \329_b1 , w_360 );
and ( \351_b0 , \322_A[3]_b0 , w_361 );
and ( w_360 , w_361 , \329_b0 );
or ( \353_b1 , \348_b1 , \352_b1 );
xor ( \353_b0 , \348_b0 , w_362 );
not ( w_362 , w_363 );
and ( w_363 , \352_b1 , \352_b0 );
buf ( \354_SUM[4]_b1 , \353_b1 );
buf ( \354_SUM[4]_b0 , \353_b0 );
and ( \355_b0 , \354_SUM[4]_b0 , w_364 );
and ( \355_b0 , \344_b0 , w_365 );
and ( w_378 , w_379 , w_366 );
and ( w_366 , \344_b0 , w_367 );
and ( w_379 , \344_b1 , w_368 );
and ( \355_b1 , \354_SUM[4]_b0 , w_369 );
and ( \354_SUM[4]_b1 , w_380 , w_370 );
and ( w_379 , \344_b0 , w_371 );
and ( \355_b1 , \355_b0 , w_372 );
and ( w_377 , w_381 , \241_b1 );
or ( w_364 , w_365 , w_373 );
or ( w_373 , w_367 , \241_b0 );
or ( w_368 , w_369 , w_374 );
or ( w_374 , w_370 , w_375 );
or ( w_375 , w_371 , w_376 );
or ( w_376 , w_372 , w_377 );
not ( \354_SUM[4]_b1 , w_378 );
not ( \354_SUM[4]_b0 , w_379 );
not ( \355_b1 , w_380 );
not ( \241_b0 , w_381 );
buf ( \356_A[4]_b1 , \c[4]_b1 );
buf ( \356_A[4]_b0 , \c[4]_b0 );
buf ( \357_B[4]_b1 , \d[4]_b1 );
buf ( \357_B[4]_b0 , \d[4]_b0 );
or ( \358_b1 , \356_A[4]_b1 , \357_B[4]_b1 );
xor ( \358_b0 , \356_A[4]_b0 , w_382 );
not ( w_382 , w_383 );
and ( w_383 , \357_B[4]_b1 , \357_B[4]_b0 );
or ( \359_b1 , \333_A[3]_b1 , \334_B[3]_b1 );
not ( \334_B[3]_b1 , w_384 );
and ( \359_b0 , \333_A[3]_b0 , w_385 );
and ( w_384 , w_385 , \334_B[3]_b0 );
or ( \360_b1 , \334_B[3]_b1 , \339_b1 );
not ( \339_b1 , w_386 );
and ( \360_b0 , \334_B[3]_b0 , w_387 );
and ( w_386 , w_387 , \339_b0 );
or ( \361_b1 , \333_A[3]_b1 , \339_b1 );
not ( \339_b1 , w_388 );
and ( \361_b0 , \333_A[3]_b0 , w_389 );
and ( w_388 , w_389 , \339_b0 );
or ( \363_b1 , \358_b1 , \362_b1 );
xor ( \363_b0 , \358_b0 , w_390 );
not ( w_390 , w_391 );
and ( w_391 , \362_b1 , \362_b0 );
buf ( \364_SUM[4]_b1 , \363_b1 );
buf ( \364_SUM[4]_b0 , \363_b0 );
and ( \365_b0 , \364_SUM[4]_b0 , w_392 );
and ( \365_b0 , \355_b0 , w_393 );
and ( w_406 , w_407 , w_394 );
and ( w_394 , \355_b0 , w_395 );
and ( w_407 , \355_b1 , w_396 );
and ( \365_b1 , \364_SUM[4]_b0 , w_397 );
and ( \364_SUM[4]_b1 , w_408 , w_398 );
and ( w_407 , \355_b0 , w_399 );
and ( \365_b1 , \365_b0 , w_400 );
and ( w_405 , w_409 , \277_b1 );
or ( w_392 , w_393 , w_401 );
or ( w_401 , w_395 , \277_b0 );
or ( w_396 , w_397 , w_402 );
or ( w_402 , w_398 , w_403 );
or ( w_403 , w_399 , w_404 );
or ( w_404 , w_400 , w_405 );
not ( \364_SUM[4]_b1 , w_406 );
not ( \364_SUM[4]_b0 , w_407 );
not ( \365_b1 , w_408 );
not ( \277_b0 , w_409 );
and ( \366_n5[5]_b1 , 1'b0_b1 , w_410 );
xor ( w_410 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_411 );
and ( \366_n5[5]_b0 , w_411 , 1'b1_b0 );
or ( \367_b1 , \b[5]_b1 , w_412 );
or ( \367_b0 , \b[5]_b0 , \366_n5[5]_b0 );
not ( \366_n5[5]_b0 , w_413 );
and ( w_413 , w_412 , \366_n5[5]_b1 );
buf ( \368_A[5]_b1 , \c[5]_b1 );
buf ( \368_A[5]_b0 , \c[5]_b0 );
buf ( \369_B[5]_b1 , \d[5]_b1 );
buf ( \369_B[5]_b0 , \d[5]_b0 );
buf ( \370_b1 , \369_B[5]_b1 );
not ( \370_b1 , w_414 );
not ( \370_b0 , w_415 );
and ( w_414 , w_415 , \369_B[5]_b0 );
or ( \371_b1 , \368_A[5]_b1 , \370_b1 );
xor ( \371_b0 , \368_A[5]_b0 , w_416 );
not ( w_416 , w_417 );
and ( w_417 , \370_b1 , \370_b0 );
or ( \372_b1 , \345_A[4]_b1 , \347_b1 );
not ( \347_b1 , w_418 );
and ( \372_b0 , \345_A[4]_b0 , w_419 );
and ( w_418 , w_419 , \347_b0 );
or ( \373_b1 , \347_b1 , \352_b1 );
not ( \352_b1 , w_420 );
and ( \373_b0 , \347_b0 , w_421 );
and ( w_420 , w_421 , \352_b0 );
or ( \374_b1 , \345_A[4]_b1 , \352_b1 );
not ( \352_b1 , w_422 );
and ( \374_b0 , \345_A[4]_b0 , w_423 );
and ( w_422 , w_423 , \352_b0 );
or ( \376_b1 , \371_b1 , \375_b1 );
xor ( \376_b0 , \371_b0 , w_424 );
not ( w_424 , w_425 );
and ( w_425 , \375_b1 , \375_b0 );
buf ( \377_SUM[5]_b1 , \376_b1 );
buf ( \377_SUM[5]_b0 , \376_b0 );
and ( \378_b0 , \377_SUM[5]_b0 , w_426 );
and ( \378_b0 , \367_b0 , w_427 );
and ( w_440 , w_441 , w_428 );
and ( w_428 , \367_b0 , w_429 );
and ( w_441 , \367_b1 , w_430 );
and ( \378_b1 , \377_SUM[5]_b0 , w_431 );
and ( \377_SUM[5]_b1 , w_442 , w_432 );
and ( w_441 , \367_b0 , w_433 );
and ( \378_b1 , \378_b0 , w_434 );
and ( w_439 , w_443 , \241_b1 );
or ( w_426 , w_427 , w_435 );
or ( w_435 , w_429 , \241_b0 );
or ( w_430 , w_431 , w_436 );
or ( w_436 , w_432 , w_437 );
or ( w_437 , w_433 , w_438 );
or ( w_438 , w_434 , w_439 );
not ( \377_SUM[5]_b1 , w_440 );
not ( \377_SUM[5]_b0 , w_441 );
not ( \378_b1 , w_442 );
not ( \241_b0 , w_443 );
buf ( \379_A[5]_b1 , \c[5]_b1 );
buf ( \379_A[5]_b0 , \c[5]_b0 );
buf ( \380_B[5]_b1 , \d[5]_b1 );
buf ( \380_B[5]_b0 , \d[5]_b0 );
or ( \381_b1 , \379_A[5]_b1 , \380_B[5]_b1 );
xor ( \381_b0 , \379_A[5]_b0 , w_444 );
not ( w_444 , w_445 );
and ( w_445 , \380_B[5]_b1 , \380_B[5]_b0 );
or ( \382_b1 , \356_A[4]_b1 , \357_B[4]_b1 );
not ( \357_B[4]_b1 , w_446 );
and ( \382_b0 , \356_A[4]_b0 , w_447 );
and ( w_446 , w_447 , \357_B[4]_b0 );
or ( \383_b1 , \357_B[4]_b1 , \362_b1 );
not ( \362_b1 , w_448 );
and ( \383_b0 , \357_B[4]_b0 , w_449 );
and ( w_448 , w_449 , \362_b0 );
or ( \384_b1 , \356_A[4]_b1 , \362_b1 );
not ( \362_b1 , w_450 );
and ( \384_b0 , \356_A[4]_b0 , w_451 );
and ( w_450 , w_451 , \362_b0 );
or ( \386_b1 , \381_b1 , \385_b1 );
xor ( \386_b0 , \381_b0 , w_452 );
not ( w_452 , w_453 );
and ( w_453 , \385_b1 , \385_b0 );
buf ( \387_SUM[5]_b1 , \386_b1 );
buf ( \387_SUM[5]_b0 , \386_b0 );
and ( \388_b0 , \387_SUM[5]_b0 , w_454 );
and ( \388_b0 , \378_b0 , w_455 );
and ( w_468 , w_469 , w_456 );
and ( w_456 , \378_b0 , w_457 );
and ( w_469 , \378_b1 , w_458 );
and ( \388_b1 , \387_SUM[5]_b0 , w_459 );
and ( \387_SUM[5]_b1 , w_470 , w_460 );
and ( w_469 , \378_b0 , w_461 );
and ( \388_b1 , \388_b0 , w_462 );
and ( w_467 , w_471 , \277_b1 );
or ( w_454 , w_455 , w_463 );
or ( w_463 , w_457 , \277_b0 );
or ( w_458 , w_459 , w_464 );
or ( w_464 , w_460 , w_465 );
or ( w_465 , w_461 , w_466 );
or ( w_466 , w_462 , w_467 );
not ( \387_SUM[5]_b1 , w_468 );
not ( \387_SUM[5]_b0 , w_469 );
not ( \388_b1 , w_470 );
not ( \277_b0 , w_471 );
and ( \389_n5[6]_b1 , 1'b0_b1 , w_472 );
xor ( w_472 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_473 );
and ( \389_n5[6]_b0 , w_473 , 1'b1_b0 );
or ( \390_b1 , \b[6]_b1 , w_474 );
or ( \390_b0 , \b[6]_b0 , \389_n5[6]_b0 );
not ( \389_n5[6]_b0 , w_475 );
and ( w_475 , w_474 , \389_n5[6]_b1 );
buf ( \391_A[6]_b1 , \c[6]_b1 );
buf ( \391_A[6]_b0 , \c[6]_b0 );
buf ( \392_B[6]_b1 , \d[6]_b1 );
buf ( \392_B[6]_b0 , \d[6]_b0 );
buf ( \393_b1 , \392_B[6]_b1 );
not ( \393_b1 , w_476 );
not ( \393_b0 , w_477 );
and ( w_476 , w_477 , \392_B[6]_b0 );
or ( \394_b1 , \391_A[6]_b1 , \393_b1 );
xor ( \394_b0 , \391_A[6]_b0 , w_478 );
not ( w_478 , w_479 );
and ( w_479 , \393_b1 , \393_b0 );
or ( \395_b1 , \368_A[5]_b1 , \370_b1 );
not ( \370_b1 , w_480 );
and ( \395_b0 , \368_A[5]_b0 , w_481 );
and ( w_480 , w_481 , \370_b0 );
or ( \396_b1 , \370_b1 , \375_b1 );
not ( \375_b1 , w_482 );
and ( \396_b0 , \370_b0 , w_483 );
and ( w_482 , w_483 , \375_b0 );
or ( \397_b1 , \368_A[5]_b1 , \375_b1 );
not ( \375_b1 , w_484 );
and ( \397_b0 , \368_A[5]_b0 , w_485 );
and ( w_484 , w_485 , \375_b0 );
or ( \399_b1 , \394_b1 , \398_b1 );
xor ( \399_b0 , \394_b0 , w_486 );
not ( w_486 , w_487 );
and ( w_487 , \398_b1 , \398_b0 );
buf ( \400_SUM[6]_b1 , \399_b1 );
buf ( \400_SUM[6]_b0 , \399_b0 );
and ( \401_b0 , \400_SUM[6]_b0 , w_488 );
and ( \401_b0 , \390_b0 , w_489 );
and ( w_502 , w_503 , w_490 );
and ( w_490 , \390_b0 , w_491 );
and ( w_503 , \390_b1 , w_492 );
and ( \401_b1 , \400_SUM[6]_b0 , w_493 );
and ( \400_SUM[6]_b1 , w_504 , w_494 );
and ( w_503 , \390_b0 , w_495 );
and ( \401_b1 , \401_b0 , w_496 );
and ( w_501 , w_505 , \241_b1 );
or ( w_488 , w_489 , w_497 );
or ( w_497 , w_491 , \241_b0 );
or ( w_492 , w_493 , w_498 );
or ( w_498 , w_494 , w_499 );
or ( w_499 , w_495 , w_500 );
or ( w_500 , w_496 , w_501 );
not ( \400_SUM[6]_b1 , w_502 );
not ( \400_SUM[6]_b0 , w_503 );
not ( \401_b1 , w_504 );
not ( \241_b0 , w_505 );
buf ( \402_A[6]_b1 , \c[6]_b1 );
buf ( \402_A[6]_b0 , \c[6]_b0 );
buf ( \403_B[6]_b1 , \d[6]_b1 );
buf ( \403_B[6]_b0 , \d[6]_b0 );
or ( \404_b1 , \402_A[6]_b1 , \403_B[6]_b1 );
xor ( \404_b0 , \402_A[6]_b0 , w_506 );
not ( w_506 , w_507 );
and ( w_507 , \403_B[6]_b1 , \403_B[6]_b0 );
or ( \405_b1 , \379_A[5]_b1 , \380_B[5]_b1 );
not ( \380_B[5]_b1 , w_508 );
and ( \405_b0 , \379_A[5]_b0 , w_509 );
and ( w_508 , w_509 , \380_B[5]_b0 );
or ( \406_b1 , \380_B[5]_b1 , \385_b1 );
not ( \385_b1 , w_510 );
and ( \406_b0 , \380_B[5]_b0 , w_511 );
and ( w_510 , w_511 , \385_b0 );
or ( \407_b1 , \379_A[5]_b1 , \385_b1 );
not ( \385_b1 , w_512 );
and ( \407_b0 , \379_A[5]_b0 , w_513 );
and ( w_512 , w_513 , \385_b0 );
or ( \409_b1 , \404_b1 , \408_b1 );
xor ( \409_b0 , \404_b0 , w_514 );
not ( w_514 , w_515 );
and ( w_515 , \408_b1 , \408_b0 );
buf ( \410_SUM[6]_b1 , \409_b1 );
buf ( \410_SUM[6]_b0 , \409_b0 );
and ( \411_b0 , \410_SUM[6]_b0 , w_516 );
and ( \411_b0 , \401_b0 , w_517 );
and ( w_530 , w_531 , w_518 );
and ( w_518 , \401_b0 , w_519 );
and ( w_531 , \401_b1 , w_520 );
and ( \411_b1 , \410_SUM[6]_b0 , w_521 );
and ( \410_SUM[6]_b1 , w_532 , w_522 );
and ( w_531 , \401_b0 , w_523 );
and ( \411_b1 , \411_b0 , w_524 );
and ( w_529 , w_533 , \277_b1 );
or ( w_516 , w_517 , w_525 );
or ( w_525 , w_519 , \277_b0 );
or ( w_520 , w_521 , w_526 );
or ( w_526 , w_522 , w_527 );
or ( w_527 , w_523 , w_528 );
or ( w_528 , w_524 , w_529 );
not ( \410_SUM[6]_b1 , w_530 );
not ( \410_SUM[6]_b0 , w_531 );
not ( \411_b1 , w_532 );
not ( \277_b0 , w_533 );
and ( \412_n5[7]_b1 , 1'b0_b1 , w_534 );
xor ( w_534 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_535 );
and ( \412_n5[7]_b0 , w_535 , 1'b1_b0 );
or ( \413_b1 , \b[7]_b1 , w_536 );
or ( \413_b0 , \b[7]_b0 , \412_n5[7]_b0 );
not ( \412_n5[7]_b0 , w_537 );
and ( w_537 , w_536 , \412_n5[7]_b1 );
buf ( \414_A[7]_b1 , \c[7]_b1 );
buf ( \414_A[7]_b0 , \c[7]_b0 );
buf ( \415_B[7]_b1 , \d[7]_b1 );
buf ( \415_B[7]_b0 , \d[7]_b0 );
buf ( \416_b1 , \415_B[7]_b1 );
not ( \416_b1 , w_538 );
not ( \416_b0 , w_539 );
and ( w_538 , w_539 , \415_B[7]_b0 );
or ( \417_b1 , \414_A[7]_b1 , \416_b1 );
xor ( \417_b0 , \414_A[7]_b0 , w_540 );
not ( w_540 , w_541 );
and ( w_541 , \416_b1 , \416_b0 );
or ( \418_b1 , \391_A[6]_b1 , \393_b1 );
not ( \393_b1 , w_542 );
and ( \418_b0 , \391_A[6]_b0 , w_543 );
and ( w_542 , w_543 , \393_b0 );
or ( \419_b1 , \393_b1 , \398_b1 );
not ( \398_b1 , w_544 );
and ( \419_b0 , \393_b0 , w_545 );
and ( w_544 , w_545 , \398_b0 );
or ( \420_b1 , \391_A[6]_b1 , \398_b1 );
not ( \398_b1 , w_546 );
and ( \420_b0 , \391_A[6]_b0 , w_547 );
and ( w_546 , w_547 , \398_b0 );
or ( \422_b1 , \417_b1 , \421_b1 );
xor ( \422_b0 , \417_b0 , w_548 );
not ( w_548 , w_549 );
and ( w_549 , \421_b1 , \421_b0 );
buf ( \423_SUM[7]_b1 , \422_b1 );
buf ( \423_SUM[7]_b0 , \422_b0 );
and ( \424_b0 , \423_SUM[7]_b0 , w_550 );
and ( \424_b0 , \413_b0 , w_551 );
and ( w_564 , w_565 , w_552 );
and ( w_552 , \413_b0 , w_553 );
and ( w_565 , \413_b1 , w_554 );
and ( \424_b1 , \423_SUM[7]_b0 , w_555 );
and ( \423_SUM[7]_b1 , w_566 , w_556 );
and ( w_565 , \413_b0 , w_557 );
and ( \424_b1 , \424_b0 , w_558 );
and ( w_563 , w_567 , \241_b1 );
or ( w_550 , w_551 , w_559 );
or ( w_559 , w_553 , \241_b0 );
or ( w_554 , w_555 , w_560 );
or ( w_560 , w_556 , w_561 );
or ( w_561 , w_557 , w_562 );
or ( w_562 , w_558 , w_563 );
not ( \423_SUM[7]_b1 , w_564 );
not ( \423_SUM[7]_b0 , w_565 );
not ( \424_b1 , w_566 );
not ( \241_b0 , w_567 );
buf ( \425_A[7]_b1 , \c[7]_b1 );
buf ( \425_A[7]_b0 , \c[7]_b0 );
buf ( \426_B[7]_b1 , \d[7]_b1 );
buf ( \426_B[7]_b0 , \d[7]_b0 );
or ( \427_b1 , \425_A[7]_b1 , \426_B[7]_b1 );
xor ( \427_b0 , \425_A[7]_b0 , w_568 );
not ( w_568 , w_569 );
and ( w_569 , \426_B[7]_b1 , \426_B[7]_b0 );
or ( \428_b1 , \402_A[6]_b1 , \403_B[6]_b1 );
not ( \403_B[6]_b1 , w_570 );
and ( \428_b0 , \402_A[6]_b0 , w_571 );
and ( w_570 , w_571 , \403_B[6]_b0 );
or ( \429_b1 , \403_B[6]_b1 , \408_b1 );
not ( \408_b1 , w_572 );
and ( \429_b0 , \403_B[6]_b0 , w_573 );
and ( w_572 , w_573 , \408_b0 );
or ( \430_b1 , \402_A[6]_b1 , \408_b1 );
not ( \408_b1 , w_574 );
and ( \430_b0 , \402_A[6]_b0 , w_575 );
and ( w_574 , w_575 , \408_b0 );
or ( \432_b1 , \427_b1 , \431_b1 );
xor ( \432_b0 , \427_b0 , w_576 );
not ( w_576 , w_577 );
and ( w_577 , \431_b1 , \431_b0 );
buf ( \433_SUM[7]_b1 , \432_b1 );
buf ( \433_SUM[7]_b0 , \432_b0 );
and ( \434_b0 , \433_SUM[7]_b0 , w_578 );
and ( \434_b0 , \424_b0 , w_579 );
and ( w_592 , w_593 , w_580 );
and ( w_580 , \424_b0 , w_581 );
and ( w_593 , \424_b1 , w_582 );
and ( \434_b1 , \433_SUM[7]_b0 , w_583 );
and ( \433_SUM[7]_b1 , w_594 , w_584 );
and ( w_593 , \424_b0 , w_585 );
and ( \434_b1 , \434_b0 , w_586 );
and ( w_591 , w_595 , \277_b1 );
or ( w_578 , w_579 , w_587 );
or ( w_587 , w_581 , \277_b0 );
or ( w_582 , w_583 , w_588 );
or ( w_588 , w_584 , w_589 );
or ( w_589 , w_585 , w_590 );
or ( w_590 , w_586 , w_591 );
not ( \433_SUM[7]_b1 , w_592 );
not ( \433_SUM[7]_b0 , w_593 );
not ( \434_b1 , w_594 );
not ( \277_b0 , w_595 );
and ( \435_n5[8]_b1 , 1'b0_b1 , w_596 );
xor ( w_596 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_597 );
and ( \435_n5[8]_b0 , w_597 , 1'b1_b0 );
or ( \436_b1 , \b[8]_b1 , w_598 );
or ( \436_b0 , \b[8]_b0 , \435_n5[8]_b0 );
not ( \435_n5[8]_b0 , w_599 );
and ( w_599 , w_598 , \435_n5[8]_b1 );
buf ( \437_A[8]_b1 , \c[8]_b1 );
buf ( \437_A[8]_b0 , \c[8]_b0 );
buf ( \438_B[8]_b1 , \d[8]_b1 );
buf ( \438_B[8]_b0 , \d[8]_b0 );
buf ( \439_b1 , \438_B[8]_b1 );
not ( \439_b1 , w_600 );
not ( \439_b0 , w_601 );
and ( w_600 , w_601 , \438_B[8]_b0 );
or ( \440_b1 , \437_A[8]_b1 , \439_b1 );
xor ( \440_b0 , \437_A[8]_b0 , w_602 );
not ( w_602 , w_603 );
and ( w_603 , \439_b1 , \439_b0 );
or ( \441_b1 , \414_A[7]_b1 , \416_b1 );
not ( \416_b1 , w_604 );
and ( \441_b0 , \414_A[7]_b0 , w_605 );
and ( w_604 , w_605 , \416_b0 );
or ( \442_b1 , \416_b1 , \421_b1 );
not ( \421_b1 , w_606 );
and ( \442_b0 , \416_b0 , w_607 );
and ( w_606 , w_607 , \421_b0 );
or ( \443_b1 , \414_A[7]_b1 , \421_b1 );
not ( \421_b1 , w_608 );
and ( \443_b0 , \414_A[7]_b0 , w_609 );
and ( w_608 , w_609 , \421_b0 );
or ( \445_b1 , \440_b1 , \444_b1 );
xor ( \445_b0 , \440_b0 , w_610 );
not ( w_610 , w_611 );
and ( w_611 , \444_b1 , \444_b0 );
buf ( \446_SUM[8]_b1 , \445_b1 );
buf ( \446_SUM[8]_b0 , \445_b0 );
and ( \447_b0 , \446_SUM[8]_b0 , w_612 );
and ( \447_b0 , \436_b0 , w_613 );
and ( w_626 , w_627 , w_614 );
and ( w_614 , \436_b0 , w_615 );
and ( w_627 , \436_b1 , w_616 );
and ( \447_b1 , \446_SUM[8]_b0 , w_617 );
and ( \446_SUM[8]_b1 , w_628 , w_618 );
and ( w_627 , \436_b0 , w_619 );
and ( \447_b1 , \447_b0 , w_620 );
and ( w_625 , w_629 , \241_b1 );
or ( w_612 , w_613 , w_621 );
or ( w_621 , w_615 , \241_b0 );
or ( w_616 , w_617 , w_622 );
or ( w_622 , w_618 , w_623 );
or ( w_623 , w_619 , w_624 );
or ( w_624 , w_620 , w_625 );
not ( \446_SUM[8]_b1 , w_626 );
not ( \446_SUM[8]_b0 , w_627 );
not ( \447_b1 , w_628 );
not ( \241_b0 , w_629 );
buf ( \448_A[8]_b1 , \c[8]_b1 );
buf ( \448_A[8]_b0 , \c[8]_b0 );
buf ( \449_B[8]_b1 , \d[8]_b1 );
buf ( \449_B[8]_b0 , \d[8]_b0 );
or ( \450_b1 , \448_A[8]_b1 , \449_B[8]_b1 );
xor ( \450_b0 , \448_A[8]_b0 , w_630 );
not ( w_630 , w_631 );
and ( w_631 , \449_B[8]_b1 , \449_B[8]_b0 );
or ( \451_b1 , \425_A[7]_b1 , \426_B[7]_b1 );
not ( \426_B[7]_b1 , w_632 );
and ( \451_b0 , \425_A[7]_b0 , w_633 );
and ( w_632 , w_633 , \426_B[7]_b0 );
or ( \452_b1 , \426_B[7]_b1 , \431_b1 );
not ( \431_b1 , w_634 );
and ( \452_b0 , \426_B[7]_b0 , w_635 );
and ( w_634 , w_635 , \431_b0 );
or ( \453_b1 , \425_A[7]_b1 , \431_b1 );
not ( \431_b1 , w_636 );
and ( \453_b0 , \425_A[7]_b0 , w_637 );
and ( w_636 , w_637 , \431_b0 );
or ( \455_b1 , \450_b1 , \454_b1 );
xor ( \455_b0 , \450_b0 , w_638 );
not ( w_638 , w_639 );
and ( w_639 , \454_b1 , \454_b0 );
buf ( \456_SUM[8]_b1 , \455_b1 );
buf ( \456_SUM[8]_b0 , \455_b0 );
and ( \457_b0 , \456_SUM[8]_b0 , w_640 );
and ( \457_b0 , \447_b0 , w_641 );
and ( w_654 , w_655 , w_642 );
and ( w_642 , \447_b0 , w_643 );
and ( w_655 , \447_b1 , w_644 );
and ( \457_b1 , \456_SUM[8]_b0 , w_645 );
and ( \456_SUM[8]_b1 , w_656 , w_646 );
and ( w_655 , \447_b0 , w_647 );
and ( \457_b1 , \457_b0 , w_648 );
and ( w_653 , w_657 , \277_b1 );
or ( w_640 , w_641 , w_649 );
or ( w_649 , w_643 , \277_b0 );
or ( w_644 , w_645 , w_650 );
or ( w_650 , w_646 , w_651 );
or ( w_651 , w_647 , w_652 );
or ( w_652 , w_648 , w_653 );
not ( \456_SUM[8]_b1 , w_654 );
not ( \456_SUM[8]_b0 , w_655 );
not ( \457_b1 , w_656 );
not ( \277_b0 , w_657 );
and ( \458_n5[9]_b1 , 1'b0_b1 , w_658 );
xor ( w_658 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_659 );
and ( \458_n5[9]_b0 , w_659 , 1'b1_b0 );
or ( \459_b1 , \b[9]_b1 , w_660 );
or ( \459_b0 , \b[9]_b0 , \458_n5[9]_b0 );
not ( \458_n5[9]_b0 , w_661 );
and ( w_661 , w_660 , \458_n5[9]_b1 );
buf ( \460_A[9]_b1 , \c[9]_b1 );
buf ( \460_A[9]_b0 , \c[9]_b0 );
buf ( \461_B[9]_b1 , \d[9]_b1 );
buf ( \461_B[9]_b0 , \d[9]_b0 );
buf ( \462_b1 , \461_B[9]_b1 );
not ( \462_b1 , w_662 );
not ( \462_b0 , w_663 );
and ( w_662 , w_663 , \461_B[9]_b0 );
or ( \463_b1 , \460_A[9]_b1 , \462_b1 );
xor ( \463_b0 , \460_A[9]_b0 , w_664 );
not ( w_664 , w_665 );
and ( w_665 , \462_b1 , \462_b0 );
or ( \464_b1 , \437_A[8]_b1 , \439_b1 );
not ( \439_b1 , w_666 );
and ( \464_b0 , \437_A[8]_b0 , w_667 );
and ( w_666 , w_667 , \439_b0 );
or ( \465_b1 , \439_b1 , \444_b1 );
not ( \444_b1 , w_668 );
and ( \465_b0 , \439_b0 , w_669 );
and ( w_668 , w_669 , \444_b0 );
or ( \466_b1 , \437_A[8]_b1 , \444_b1 );
not ( \444_b1 , w_670 );
and ( \466_b0 , \437_A[8]_b0 , w_671 );
and ( w_670 , w_671 , \444_b0 );
or ( \468_b1 , \463_b1 , \467_b1 );
xor ( \468_b0 , \463_b0 , w_672 );
not ( w_672 , w_673 );
and ( w_673 , \467_b1 , \467_b0 );
buf ( \469_SUM[9]_b1 , \468_b1 );
buf ( \469_SUM[9]_b0 , \468_b0 );
and ( \470_b0 , \469_SUM[9]_b0 , w_674 );
and ( \470_b0 , \459_b0 , w_675 );
and ( w_688 , w_689 , w_676 );
and ( w_676 , \459_b0 , w_677 );
and ( w_689 , \459_b1 , w_678 );
and ( \470_b1 , \469_SUM[9]_b0 , w_679 );
and ( \469_SUM[9]_b1 , w_690 , w_680 );
and ( w_689 , \459_b0 , w_681 );
and ( \470_b1 , \470_b0 , w_682 );
and ( w_687 , w_691 , \241_b1 );
or ( w_674 , w_675 , w_683 );
or ( w_683 , w_677 , \241_b0 );
or ( w_678 , w_679 , w_684 );
or ( w_684 , w_680 , w_685 );
or ( w_685 , w_681 , w_686 );
or ( w_686 , w_682 , w_687 );
not ( \469_SUM[9]_b1 , w_688 );
not ( \469_SUM[9]_b0 , w_689 );
not ( \470_b1 , w_690 );
not ( \241_b0 , w_691 );
buf ( \471_A[9]_b1 , \c[9]_b1 );
buf ( \471_A[9]_b0 , \c[9]_b0 );
buf ( \472_B[9]_b1 , \d[9]_b1 );
buf ( \472_B[9]_b0 , \d[9]_b0 );
or ( \473_b1 , \471_A[9]_b1 , \472_B[9]_b1 );
xor ( \473_b0 , \471_A[9]_b0 , w_692 );
not ( w_692 , w_693 );
and ( w_693 , \472_B[9]_b1 , \472_B[9]_b0 );
or ( \474_b1 , \448_A[8]_b1 , \449_B[8]_b1 );
not ( \449_B[8]_b1 , w_694 );
and ( \474_b0 , \448_A[8]_b0 , w_695 );
and ( w_694 , w_695 , \449_B[8]_b0 );
or ( \475_b1 , \449_B[8]_b1 , \454_b1 );
not ( \454_b1 , w_696 );
and ( \475_b0 , \449_B[8]_b0 , w_697 );
and ( w_696 , w_697 , \454_b0 );
or ( \476_b1 , \448_A[8]_b1 , \454_b1 );
not ( \454_b1 , w_698 );
and ( \476_b0 , \448_A[8]_b0 , w_699 );
and ( w_698 , w_699 , \454_b0 );
or ( \478_b1 , \473_b1 , \477_b1 );
xor ( \478_b0 , \473_b0 , w_700 );
not ( w_700 , w_701 );
and ( w_701 , \477_b1 , \477_b0 );
buf ( \479_SUM[9]_b1 , \478_b1 );
buf ( \479_SUM[9]_b0 , \478_b0 );
and ( \480_b0 , \479_SUM[9]_b0 , w_702 );
and ( \480_b0 , \470_b0 , w_703 );
and ( w_716 , w_717 , w_704 );
and ( w_704 , \470_b0 , w_705 );
and ( w_717 , \470_b1 , w_706 );
and ( \480_b1 , \479_SUM[9]_b0 , w_707 );
and ( \479_SUM[9]_b1 , w_718 , w_708 );
and ( w_717 , \470_b0 , w_709 );
and ( \480_b1 , \480_b0 , w_710 );
and ( w_715 , w_719 , \277_b1 );
or ( w_702 , w_703 , w_711 );
or ( w_711 , w_705 , \277_b0 );
or ( w_706 , w_707 , w_712 );
or ( w_712 , w_708 , w_713 );
or ( w_713 , w_709 , w_714 );
or ( w_714 , w_710 , w_715 );
not ( \479_SUM[9]_b1 , w_716 );
not ( \479_SUM[9]_b0 , w_717 );
not ( \480_b1 , w_718 );
not ( \277_b0 , w_719 );
and ( \481_n5[10]_b1 , 1'b0_b1 , w_720 );
xor ( w_720 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_721 );
and ( \481_n5[10]_b0 , w_721 , 1'b1_b0 );
or ( \482_b1 , \b[10]_b1 , w_722 );
or ( \482_b0 , \b[10]_b0 , \481_n5[10]_b0 );
not ( \481_n5[10]_b0 , w_723 );
and ( w_723 , w_722 , \481_n5[10]_b1 );
buf ( \483_A[10]_b1 , \c[10]_b1 );
buf ( \483_A[10]_b0 , \c[10]_b0 );
buf ( \484_B[10]_b1 , \d[10]_b1 );
buf ( \484_B[10]_b0 , \d[10]_b0 );
buf ( \485_b1 , \484_B[10]_b1 );
not ( \485_b1 , w_724 );
not ( \485_b0 , w_725 );
and ( w_724 , w_725 , \484_B[10]_b0 );
or ( \486_b1 , \483_A[10]_b1 , \485_b1 );
xor ( \486_b0 , \483_A[10]_b0 , w_726 );
not ( w_726 , w_727 );
and ( w_727 , \485_b1 , \485_b0 );
or ( \487_b1 , \460_A[9]_b1 , \462_b1 );
not ( \462_b1 , w_728 );
and ( \487_b0 , \460_A[9]_b0 , w_729 );
and ( w_728 , w_729 , \462_b0 );
or ( \488_b1 , \462_b1 , \467_b1 );
not ( \467_b1 , w_730 );
and ( \488_b0 , \462_b0 , w_731 );
and ( w_730 , w_731 , \467_b0 );
or ( \489_b1 , \460_A[9]_b1 , \467_b1 );
not ( \467_b1 , w_732 );
and ( \489_b0 , \460_A[9]_b0 , w_733 );
and ( w_732 , w_733 , \467_b0 );
or ( \491_b1 , \486_b1 , \490_b1 );
xor ( \491_b0 , \486_b0 , w_734 );
not ( w_734 , w_735 );
and ( w_735 , \490_b1 , \490_b0 );
buf ( \492_SUM[10]_b1 , \491_b1 );
buf ( \492_SUM[10]_b0 , \491_b0 );
and ( \493_b0 , \492_SUM[10]_b0 , w_736 );
and ( \493_b0 , \482_b0 , w_737 );
and ( w_750 , w_751 , w_738 );
and ( w_738 , \482_b0 , w_739 );
and ( w_751 , \482_b1 , w_740 );
and ( \493_b1 , \492_SUM[10]_b0 , w_741 );
and ( \492_SUM[10]_b1 , w_752 , w_742 );
and ( w_751 , \482_b0 , w_743 );
and ( \493_b1 , \493_b0 , w_744 );
and ( w_749 , w_753 , \241_b1 );
or ( w_736 , w_737 , w_745 );
or ( w_745 , w_739 , \241_b0 );
or ( w_740 , w_741 , w_746 );
or ( w_746 , w_742 , w_747 );
or ( w_747 , w_743 , w_748 );
or ( w_748 , w_744 , w_749 );
not ( \492_SUM[10]_b1 , w_750 );
not ( \492_SUM[10]_b0 , w_751 );
not ( \493_b1 , w_752 );
not ( \241_b0 , w_753 );
buf ( \494_A[10]_b1 , \c[10]_b1 );
buf ( \494_A[10]_b0 , \c[10]_b0 );
buf ( \495_B[10]_b1 , \d[10]_b1 );
buf ( \495_B[10]_b0 , \d[10]_b0 );
or ( \496_b1 , \494_A[10]_b1 , \495_B[10]_b1 );
xor ( \496_b0 , \494_A[10]_b0 , w_754 );
not ( w_754 , w_755 );
and ( w_755 , \495_B[10]_b1 , \495_B[10]_b0 );
or ( \497_b1 , \471_A[9]_b1 , \472_B[9]_b1 );
not ( \472_B[9]_b1 , w_756 );
and ( \497_b0 , \471_A[9]_b0 , w_757 );
and ( w_756 , w_757 , \472_B[9]_b0 );
or ( \498_b1 , \472_B[9]_b1 , \477_b1 );
not ( \477_b1 , w_758 );
and ( \498_b0 , \472_B[9]_b0 , w_759 );
and ( w_758 , w_759 , \477_b0 );
or ( \499_b1 , \471_A[9]_b1 , \477_b1 );
not ( \477_b1 , w_760 );
and ( \499_b0 , \471_A[9]_b0 , w_761 );
and ( w_760 , w_761 , \477_b0 );
or ( \501_b1 , \496_b1 , \500_b1 );
xor ( \501_b0 , \496_b0 , w_762 );
not ( w_762 , w_763 );
and ( w_763 , \500_b1 , \500_b0 );
buf ( \502_SUM[10]_b1 , \501_b1 );
buf ( \502_SUM[10]_b0 , \501_b0 );
and ( \503_b0 , \502_SUM[10]_b0 , w_764 );
and ( \503_b0 , \493_b0 , w_765 );
and ( w_778 , w_779 , w_766 );
and ( w_766 , \493_b0 , w_767 );
and ( w_779 , \493_b1 , w_768 );
and ( \503_b1 , \502_SUM[10]_b0 , w_769 );
and ( \502_SUM[10]_b1 , w_780 , w_770 );
and ( w_779 , \493_b0 , w_771 );
and ( \503_b1 , \503_b0 , w_772 );
and ( w_777 , w_781 , \277_b1 );
or ( w_764 , w_765 , w_773 );
or ( w_773 , w_767 , \277_b0 );
or ( w_768 , w_769 , w_774 );
or ( w_774 , w_770 , w_775 );
or ( w_775 , w_771 , w_776 );
or ( w_776 , w_772 , w_777 );
not ( \502_SUM[10]_b1 , w_778 );
not ( \502_SUM[10]_b0 , w_779 );
not ( \503_b1 , w_780 );
not ( \277_b0 , w_781 );
and ( \504_n5[11]_b1 , 1'b0_b1 , w_782 );
xor ( w_782 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_783 );
and ( \504_n5[11]_b0 , w_783 , 1'b1_b0 );
or ( \505_b1 , \b[11]_b1 , w_784 );
or ( \505_b0 , \b[11]_b0 , \504_n5[11]_b0 );
not ( \504_n5[11]_b0 , w_785 );
and ( w_785 , w_784 , \504_n5[11]_b1 );
buf ( \506_A[11]_b1 , \c[11]_b1 );
buf ( \506_A[11]_b0 , \c[11]_b0 );
buf ( \507_B[11]_b1 , \d[11]_b1 );
buf ( \507_B[11]_b0 , \d[11]_b0 );
buf ( \508_b1 , \507_B[11]_b1 );
not ( \508_b1 , w_786 );
not ( \508_b0 , w_787 );
and ( w_786 , w_787 , \507_B[11]_b0 );
or ( \509_b1 , \506_A[11]_b1 , \508_b1 );
xor ( \509_b0 , \506_A[11]_b0 , w_788 );
not ( w_788 , w_789 );
and ( w_789 , \508_b1 , \508_b0 );
or ( \510_b1 , \483_A[10]_b1 , \485_b1 );
not ( \485_b1 , w_790 );
and ( \510_b0 , \483_A[10]_b0 , w_791 );
and ( w_790 , w_791 , \485_b0 );
or ( \511_b1 , \485_b1 , \490_b1 );
not ( \490_b1 , w_792 );
and ( \511_b0 , \485_b0 , w_793 );
and ( w_792 , w_793 , \490_b0 );
or ( \512_b1 , \483_A[10]_b1 , \490_b1 );
not ( \490_b1 , w_794 );
and ( \512_b0 , \483_A[10]_b0 , w_795 );
and ( w_794 , w_795 , \490_b0 );
or ( \514_b1 , \509_b1 , \513_b1 );
xor ( \514_b0 , \509_b0 , w_796 );
not ( w_796 , w_797 );
and ( w_797 , \513_b1 , \513_b0 );
buf ( \515_SUM[11]_b1 , \514_b1 );
buf ( \515_SUM[11]_b0 , \514_b0 );
and ( \516_b0 , \515_SUM[11]_b0 , w_798 );
and ( \516_b0 , \505_b0 , w_799 );
and ( w_812 , w_813 , w_800 );
and ( w_800 , \505_b0 , w_801 );
and ( w_813 , \505_b1 , w_802 );
and ( \516_b1 , \515_SUM[11]_b0 , w_803 );
and ( \515_SUM[11]_b1 , w_814 , w_804 );
and ( w_813 , \505_b0 , w_805 );
and ( \516_b1 , \516_b0 , w_806 );
and ( w_811 , w_815 , \241_b1 );
or ( w_798 , w_799 , w_807 );
or ( w_807 , w_801 , \241_b0 );
or ( w_802 , w_803 , w_808 );
or ( w_808 , w_804 , w_809 );
or ( w_809 , w_805 , w_810 );
or ( w_810 , w_806 , w_811 );
not ( \515_SUM[11]_b1 , w_812 );
not ( \515_SUM[11]_b0 , w_813 );
not ( \516_b1 , w_814 );
not ( \241_b0 , w_815 );
buf ( \517_A[11]_b1 , \c[11]_b1 );
buf ( \517_A[11]_b0 , \c[11]_b0 );
buf ( \518_B[11]_b1 , \d[11]_b1 );
buf ( \518_B[11]_b0 , \d[11]_b0 );
or ( \519_b1 , \517_A[11]_b1 , \518_B[11]_b1 );
xor ( \519_b0 , \517_A[11]_b0 , w_816 );
not ( w_816 , w_817 );
and ( w_817 , \518_B[11]_b1 , \518_B[11]_b0 );
or ( \520_b1 , \494_A[10]_b1 , \495_B[10]_b1 );
not ( \495_B[10]_b1 , w_818 );
and ( \520_b0 , \494_A[10]_b0 , w_819 );
and ( w_818 , w_819 , \495_B[10]_b0 );
or ( \521_b1 , \495_B[10]_b1 , \500_b1 );
not ( \500_b1 , w_820 );
and ( \521_b0 , \495_B[10]_b0 , w_821 );
and ( w_820 , w_821 , \500_b0 );
or ( \522_b1 , \494_A[10]_b1 , \500_b1 );
not ( \500_b1 , w_822 );
and ( \522_b0 , \494_A[10]_b0 , w_823 );
and ( w_822 , w_823 , \500_b0 );
or ( \524_b1 , \519_b1 , \523_b1 );
xor ( \524_b0 , \519_b0 , w_824 );
not ( w_824 , w_825 );
and ( w_825 , \523_b1 , \523_b0 );
buf ( \525_SUM[11]_b1 , \524_b1 );
buf ( \525_SUM[11]_b0 , \524_b0 );
and ( \526_b0 , \525_SUM[11]_b0 , w_826 );
and ( \526_b0 , \516_b0 , w_827 );
and ( w_840 , w_841 , w_828 );
and ( w_828 , \516_b0 , w_829 );
and ( w_841 , \516_b1 , w_830 );
and ( \526_b1 , \525_SUM[11]_b0 , w_831 );
and ( \525_SUM[11]_b1 , w_842 , w_832 );
and ( w_841 , \516_b0 , w_833 );
and ( \526_b1 , \526_b0 , w_834 );
and ( w_839 , w_843 , \277_b1 );
or ( w_826 , w_827 , w_835 );
or ( w_835 , w_829 , \277_b0 );
or ( w_830 , w_831 , w_836 );
or ( w_836 , w_832 , w_837 );
or ( w_837 , w_833 , w_838 );
or ( w_838 , w_834 , w_839 );
not ( \525_SUM[11]_b1 , w_840 );
not ( \525_SUM[11]_b0 , w_841 );
not ( \526_b1 , w_842 );
not ( \277_b0 , w_843 );
and ( \527_n5[12]_b1 , 1'b0_b1 , w_844 );
xor ( w_844 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_845 );
and ( \527_n5[12]_b0 , w_845 , 1'b1_b0 );
or ( \528_b1 , \b[12]_b1 , w_846 );
or ( \528_b0 , \b[12]_b0 , \527_n5[12]_b0 );
not ( \527_n5[12]_b0 , w_847 );
and ( w_847 , w_846 , \527_n5[12]_b1 );
buf ( \529_A[12]_b1 , \c[12]_b1 );
buf ( \529_A[12]_b0 , \c[12]_b0 );
buf ( \530_B[12]_b1 , \d[12]_b1 );
buf ( \530_B[12]_b0 , \d[12]_b0 );
buf ( \531_b1 , \530_B[12]_b1 );
not ( \531_b1 , w_848 );
not ( \531_b0 , w_849 );
and ( w_848 , w_849 , \530_B[12]_b0 );
or ( \532_b1 , \529_A[12]_b1 , \531_b1 );
xor ( \532_b0 , \529_A[12]_b0 , w_850 );
not ( w_850 , w_851 );
and ( w_851 , \531_b1 , \531_b0 );
or ( \533_b1 , \506_A[11]_b1 , \508_b1 );
not ( \508_b1 , w_852 );
and ( \533_b0 , \506_A[11]_b0 , w_853 );
and ( w_852 , w_853 , \508_b0 );
or ( \534_b1 , \508_b1 , \513_b1 );
not ( \513_b1 , w_854 );
and ( \534_b0 , \508_b0 , w_855 );
and ( w_854 , w_855 , \513_b0 );
or ( \535_b1 , \506_A[11]_b1 , \513_b1 );
not ( \513_b1 , w_856 );
and ( \535_b0 , \506_A[11]_b0 , w_857 );
and ( w_856 , w_857 , \513_b0 );
or ( \537_b1 , \532_b1 , \536_b1 );
xor ( \537_b0 , \532_b0 , w_858 );
not ( w_858 , w_859 );
and ( w_859 , \536_b1 , \536_b0 );
buf ( \538_SUM[12]_b1 , \537_b1 );
buf ( \538_SUM[12]_b0 , \537_b0 );
and ( \539_b0 , \538_SUM[12]_b0 , w_860 );
and ( \539_b0 , \528_b0 , w_861 );
and ( w_874 , w_875 , w_862 );
and ( w_862 , \528_b0 , w_863 );
and ( w_875 , \528_b1 , w_864 );
and ( \539_b1 , \538_SUM[12]_b0 , w_865 );
and ( \538_SUM[12]_b1 , w_876 , w_866 );
and ( w_875 , \528_b0 , w_867 );
and ( \539_b1 , \539_b0 , w_868 );
and ( w_873 , w_877 , \241_b1 );
or ( w_860 , w_861 , w_869 );
or ( w_869 , w_863 , \241_b0 );
or ( w_864 , w_865 , w_870 );
or ( w_870 , w_866 , w_871 );
or ( w_871 , w_867 , w_872 );
or ( w_872 , w_868 , w_873 );
not ( \538_SUM[12]_b1 , w_874 );
not ( \538_SUM[12]_b0 , w_875 );
not ( \539_b1 , w_876 );
not ( \241_b0 , w_877 );
buf ( \540_A[12]_b1 , \c[12]_b1 );
buf ( \540_A[12]_b0 , \c[12]_b0 );
buf ( \541_B[12]_b1 , \d[12]_b1 );
buf ( \541_B[12]_b0 , \d[12]_b0 );
or ( \542_b1 , \540_A[12]_b1 , \541_B[12]_b1 );
xor ( \542_b0 , \540_A[12]_b0 , w_878 );
not ( w_878 , w_879 );
and ( w_879 , \541_B[12]_b1 , \541_B[12]_b0 );
or ( \543_b1 , \517_A[11]_b1 , \518_B[11]_b1 );
not ( \518_B[11]_b1 , w_880 );
and ( \543_b0 , \517_A[11]_b0 , w_881 );
and ( w_880 , w_881 , \518_B[11]_b0 );
or ( \544_b1 , \518_B[11]_b1 , \523_b1 );
not ( \523_b1 , w_882 );
and ( \544_b0 , \518_B[11]_b0 , w_883 );
and ( w_882 , w_883 , \523_b0 );
or ( \545_b1 , \517_A[11]_b1 , \523_b1 );
not ( \523_b1 , w_884 );
and ( \545_b0 , \517_A[11]_b0 , w_885 );
and ( w_884 , w_885 , \523_b0 );
or ( \547_b1 , \542_b1 , \546_b1 );
xor ( \547_b0 , \542_b0 , w_886 );
not ( w_886 , w_887 );
and ( w_887 , \546_b1 , \546_b0 );
buf ( \548_SUM[12]_b1 , \547_b1 );
buf ( \548_SUM[12]_b0 , \547_b0 );
and ( \549_b0 , \548_SUM[12]_b0 , w_888 );
and ( \549_b0 , \539_b0 , w_889 );
and ( w_902 , w_903 , w_890 );
and ( w_890 , \539_b0 , w_891 );
and ( w_903 , \539_b1 , w_892 );
and ( \549_b1 , \548_SUM[12]_b0 , w_893 );
and ( \548_SUM[12]_b1 , w_904 , w_894 );
and ( w_903 , \539_b0 , w_895 );
and ( \549_b1 , \549_b0 , w_896 );
and ( w_901 , w_905 , \277_b1 );
or ( w_888 , w_889 , w_897 );
or ( w_897 , w_891 , \277_b0 );
or ( w_892 , w_893 , w_898 );
or ( w_898 , w_894 , w_899 );
or ( w_899 , w_895 , w_900 );
or ( w_900 , w_896 , w_901 );
not ( \548_SUM[12]_b1 , w_902 );
not ( \548_SUM[12]_b0 , w_903 );
not ( \549_b1 , w_904 );
not ( \277_b0 , w_905 );
and ( \550_n5[13]_b1 , 1'b0_b1 , w_906 );
xor ( w_906 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_907 );
and ( \550_n5[13]_b0 , w_907 , 1'b1_b0 );
or ( \551_b1 , \b[13]_b1 , w_908 );
or ( \551_b0 , \b[13]_b0 , \550_n5[13]_b0 );
not ( \550_n5[13]_b0 , w_909 );
and ( w_909 , w_908 , \550_n5[13]_b1 );
buf ( \552_A[13]_b1 , \c[13]_b1 );
buf ( \552_A[13]_b0 , \c[13]_b0 );
buf ( \553_B[13]_b1 , \d[13]_b1 );
buf ( \553_B[13]_b0 , \d[13]_b0 );
buf ( \554_b1 , \553_B[13]_b1 );
not ( \554_b1 , w_910 );
not ( \554_b0 , w_911 );
and ( w_910 , w_911 , \553_B[13]_b0 );
or ( \555_b1 , \552_A[13]_b1 , \554_b1 );
xor ( \555_b0 , \552_A[13]_b0 , w_912 );
not ( w_912 , w_913 );
and ( w_913 , \554_b1 , \554_b0 );
or ( \556_b1 , \529_A[12]_b1 , \531_b1 );
not ( \531_b1 , w_914 );
and ( \556_b0 , \529_A[12]_b0 , w_915 );
and ( w_914 , w_915 , \531_b0 );
or ( \557_b1 , \531_b1 , \536_b1 );
not ( \536_b1 , w_916 );
and ( \557_b0 , \531_b0 , w_917 );
and ( w_916 , w_917 , \536_b0 );
or ( \558_b1 , \529_A[12]_b1 , \536_b1 );
not ( \536_b1 , w_918 );
and ( \558_b0 , \529_A[12]_b0 , w_919 );
and ( w_918 , w_919 , \536_b0 );
or ( \560_b1 , \555_b1 , \559_b1 );
xor ( \560_b0 , \555_b0 , w_920 );
not ( w_920 , w_921 );
and ( w_921 , \559_b1 , \559_b0 );
buf ( \561_SUM[13]_b1 , \560_b1 );
buf ( \561_SUM[13]_b0 , \560_b0 );
and ( \562_b0 , \561_SUM[13]_b0 , w_922 );
and ( \562_b0 , \551_b0 , w_923 );
and ( w_936 , w_937 , w_924 );
and ( w_924 , \551_b0 , w_925 );
and ( w_937 , \551_b1 , w_926 );
and ( \562_b1 , \561_SUM[13]_b0 , w_927 );
and ( \561_SUM[13]_b1 , w_938 , w_928 );
and ( w_937 , \551_b0 , w_929 );
and ( \562_b1 , \562_b0 , w_930 );
and ( w_935 , w_939 , \241_b1 );
or ( w_922 , w_923 , w_931 );
or ( w_931 , w_925 , \241_b0 );
or ( w_926 , w_927 , w_932 );
or ( w_932 , w_928 , w_933 );
or ( w_933 , w_929 , w_934 );
or ( w_934 , w_930 , w_935 );
not ( \561_SUM[13]_b1 , w_936 );
not ( \561_SUM[13]_b0 , w_937 );
not ( \562_b1 , w_938 );
not ( \241_b0 , w_939 );
buf ( \563_A[13]_b1 , \c[13]_b1 );
buf ( \563_A[13]_b0 , \c[13]_b0 );
buf ( \564_B[13]_b1 , \d[13]_b1 );
buf ( \564_B[13]_b0 , \d[13]_b0 );
or ( \565_b1 , \563_A[13]_b1 , \564_B[13]_b1 );
xor ( \565_b0 , \563_A[13]_b0 , w_940 );
not ( w_940 , w_941 );
and ( w_941 , \564_B[13]_b1 , \564_B[13]_b0 );
or ( \566_b1 , \540_A[12]_b1 , \541_B[12]_b1 );
not ( \541_B[12]_b1 , w_942 );
and ( \566_b0 , \540_A[12]_b0 , w_943 );
and ( w_942 , w_943 , \541_B[12]_b0 );
or ( \567_b1 , \541_B[12]_b1 , \546_b1 );
not ( \546_b1 , w_944 );
and ( \567_b0 , \541_B[12]_b0 , w_945 );
and ( w_944 , w_945 , \546_b0 );
or ( \568_b1 , \540_A[12]_b1 , \546_b1 );
not ( \546_b1 , w_946 );
and ( \568_b0 , \540_A[12]_b0 , w_947 );
and ( w_946 , w_947 , \546_b0 );
or ( \570_b1 , \565_b1 , \569_b1 );
xor ( \570_b0 , \565_b0 , w_948 );
not ( w_948 , w_949 );
and ( w_949 , \569_b1 , \569_b0 );
buf ( \571_SUM[13]_b1 , \570_b1 );
buf ( \571_SUM[13]_b0 , \570_b0 );
and ( \572_b0 , \571_SUM[13]_b0 , w_950 );
and ( \572_b0 , \562_b0 , w_951 );
and ( w_964 , w_965 , w_952 );
and ( w_952 , \562_b0 , w_953 );
and ( w_965 , \562_b1 , w_954 );
and ( \572_b1 , \571_SUM[13]_b0 , w_955 );
and ( \571_SUM[13]_b1 , w_966 , w_956 );
and ( w_965 , \562_b0 , w_957 );
and ( \572_b1 , \572_b0 , w_958 );
and ( w_963 , w_967 , \277_b1 );
or ( w_950 , w_951 , w_959 );
or ( w_959 , w_953 , \277_b0 );
or ( w_954 , w_955 , w_960 );
or ( w_960 , w_956 , w_961 );
or ( w_961 , w_957 , w_962 );
or ( w_962 , w_958 , w_963 );
not ( \571_SUM[13]_b1 , w_964 );
not ( \571_SUM[13]_b0 , w_965 );
not ( \572_b1 , w_966 );
not ( \277_b0 , w_967 );
and ( \573_n5[14]_b1 , 1'b0_b1 , w_968 );
xor ( w_968 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_969 );
and ( \573_n5[14]_b0 , w_969 , 1'b1_b0 );
or ( \574_b1 , \b[14]_b1 , w_970 );
or ( \574_b0 , \b[14]_b0 , \573_n5[14]_b0 );
not ( \573_n5[14]_b0 , w_971 );
and ( w_971 , w_970 , \573_n5[14]_b1 );
buf ( \575_A[14]_b1 , \c[14]_b1 );
buf ( \575_A[14]_b0 , \c[14]_b0 );
buf ( \576_B[14]_b1 , \d[14]_b1 );
buf ( \576_B[14]_b0 , \d[14]_b0 );
buf ( \577_b1 , \576_B[14]_b1 );
not ( \577_b1 , w_972 );
not ( \577_b0 , w_973 );
and ( w_972 , w_973 , \576_B[14]_b0 );
or ( \578_b1 , \575_A[14]_b1 , \577_b1 );
xor ( \578_b0 , \575_A[14]_b0 , w_974 );
not ( w_974 , w_975 );
and ( w_975 , \577_b1 , \577_b0 );
or ( \579_b1 , \552_A[13]_b1 , \554_b1 );
not ( \554_b1 , w_976 );
and ( \579_b0 , \552_A[13]_b0 , w_977 );
and ( w_976 , w_977 , \554_b0 );
or ( \580_b1 , \554_b1 , \559_b1 );
not ( \559_b1 , w_978 );
and ( \580_b0 , \554_b0 , w_979 );
and ( w_978 , w_979 , \559_b0 );
or ( \581_b1 , \552_A[13]_b1 , \559_b1 );
not ( \559_b1 , w_980 );
and ( \581_b0 , \552_A[13]_b0 , w_981 );
and ( w_980 , w_981 , \559_b0 );
or ( \583_b1 , \578_b1 , \582_b1 );
xor ( \583_b0 , \578_b0 , w_982 );
not ( w_982 , w_983 );
and ( w_983 , \582_b1 , \582_b0 );
buf ( \584_SUM[14]_b1 , \583_b1 );
buf ( \584_SUM[14]_b0 , \583_b0 );
and ( \585_b0 , \584_SUM[14]_b0 , w_984 );
and ( \585_b0 , \574_b0 , w_985 );
and ( w_998 , w_999 , w_986 );
and ( w_986 , \574_b0 , w_987 );
and ( w_999 , \574_b1 , w_988 );
and ( \585_b1 , \584_SUM[14]_b0 , w_989 );
and ( \584_SUM[14]_b1 , w_1000 , w_990 );
and ( w_999 , \574_b0 , w_991 );
and ( \585_b1 , \585_b0 , w_992 );
and ( w_997 , w_1001 , \241_b1 );
or ( w_984 , w_985 , w_993 );
or ( w_993 , w_987 , \241_b0 );
or ( w_988 , w_989 , w_994 );
or ( w_994 , w_990 , w_995 );
or ( w_995 , w_991 , w_996 );
or ( w_996 , w_992 , w_997 );
not ( \584_SUM[14]_b1 , w_998 );
not ( \584_SUM[14]_b0 , w_999 );
not ( \585_b1 , w_1000 );
not ( \241_b0 , w_1001 );
buf ( \586_A[14]_b1 , \c[14]_b1 );
buf ( \586_A[14]_b0 , \c[14]_b0 );
buf ( \587_B[14]_b1 , \d[14]_b1 );
buf ( \587_B[14]_b0 , \d[14]_b0 );
or ( \588_b1 , \586_A[14]_b1 , \587_B[14]_b1 );
xor ( \588_b0 , \586_A[14]_b0 , w_1002 );
not ( w_1002 , w_1003 );
and ( w_1003 , \587_B[14]_b1 , \587_B[14]_b0 );
or ( \589_b1 , \563_A[13]_b1 , \564_B[13]_b1 );
not ( \564_B[13]_b1 , w_1004 );
and ( \589_b0 , \563_A[13]_b0 , w_1005 );
and ( w_1004 , w_1005 , \564_B[13]_b0 );
or ( \590_b1 , \564_B[13]_b1 , \569_b1 );
not ( \569_b1 , w_1006 );
and ( \590_b0 , \564_B[13]_b0 , w_1007 );
and ( w_1006 , w_1007 , \569_b0 );
or ( \591_b1 , \563_A[13]_b1 , \569_b1 );
not ( \569_b1 , w_1008 );
and ( \591_b0 , \563_A[13]_b0 , w_1009 );
and ( w_1008 , w_1009 , \569_b0 );
or ( \593_b1 , \588_b1 , \592_b1 );
xor ( \593_b0 , \588_b0 , w_1010 );
not ( w_1010 , w_1011 );
and ( w_1011 , \592_b1 , \592_b0 );
buf ( \594_SUM[14]_b1 , \593_b1 );
buf ( \594_SUM[14]_b0 , \593_b0 );
and ( \595_b0 , \594_SUM[14]_b0 , w_1012 );
and ( \595_b0 , \585_b0 , w_1013 );
and ( w_1026 , w_1027 , w_1014 );
and ( w_1014 , \585_b0 , w_1015 );
and ( w_1027 , \585_b1 , w_1016 );
and ( \595_b1 , \594_SUM[14]_b0 , w_1017 );
and ( \594_SUM[14]_b1 , w_1028 , w_1018 );
and ( w_1027 , \585_b0 , w_1019 );
and ( \595_b1 , \595_b0 , w_1020 );
and ( w_1025 , w_1029 , \277_b1 );
or ( w_1012 , w_1013 , w_1021 );
or ( w_1021 , w_1015 , \277_b0 );
or ( w_1016 , w_1017 , w_1022 );
or ( w_1022 , w_1018 , w_1023 );
or ( w_1023 , w_1019 , w_1024 );
or ( w_1024 , w_1020 , w_1025 );
not ( \594_SUM[14]_b1 , w_1026 );
not ( \594_SUM[14]_b0 , w_1027 );
not ( \595_b1 , w_1028 );
not ( \277_b0 , w_1029 );
and ( \596_n5[15]_b1 , 1'b0_b1 , w_1030 );
xor ( w_1030 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1031 );
and ( \596_n5[15]_b0 , w_1031 , 1'b1_b0 );
or ( \597_b1 , \b[15]_b1 , w_1032 );
or ( \597_b0 , \b[15]_b0 , \596_n5[15]_b0 );
not ( \596_n5[15]_b0 , w_1033 );
and ( w_1033 , w_1032 , \596_n5[15]_b1 );
buf ( \598_A[15]_b1 , \c[15]_b1 );
buf ( \598_A[15]_b0 , \c[15]_b0 );
buf ( \599_B[15]_b1 , \d[15]_b1 );
buf ( \599_B[15]_b0 , \d[15]_b0 );
buf ( \600_b1 , \599_B[15]_b1 );
not ( \600_b1 , w_1034 );
not ( \600_b0 , w_1035 );
and ( w_1034 , w_1035 , \599_B[15]_b0 );
or ( \601_b1 , \598_A[15]_b1 , \600_b1 );
xor ( \601_b0 , \598_A[15]_b0 , w_1036 );
not ( w_1036 , w_1037 );
and ( w_1037 , \600_b1 , \600_b0 );
or ( \602_b1 , \575_A[14]_b1 , \577_b1 );
not ( \577_b1 , w_1038 );
and ( \602_b0 , \575_A[14]_b0 , w_1039 );
and ( w_1038 , w_1039 , \577_b0 );
or ( \603_b1 , \577_b1 , \582_b1 );
not ( \582_b1 , w_1040 );
and ( \603_b0 , \577_b0 , w_1041 );
and ( w_1040 , w_1041 , \582_b0 );
or ( \604_b1 , \575_A[14]_b1 , \582_b1 );
not ( \582_b1 , w_1042 );
and ( \604_b0 , \575_A[14]_b0 , w_1043 );
and ( w_1042 , w_1043 , \582_b0 );
or ( \606_b1 , \601_b1 , \605_b1 );
xor ( \606_b0 , \601_b0 , w_1044 );
not ( w_1044 , w_1045 );
and ( w_1045 , \605_b1 , \605_b0 );
buf ( \607_SUM[15]_b1 , \606_b1 );
buf ( \607_SUM[15]_b0 , \606_b0 );
and ( \608_b0 , \607_SUM[15]_b0 , w_1046 );
and ( \608_b0 , \597_b0 , w_1047 );
and ( w_1060 , w_1061 , w_1048 );
and ( w_1048 , \597_b0 , w_1049 );
and ( w_1061 , \597_b1 , w_1050 );
and ( \608_b1 , \607_SUM[15]_b0 , w_1051 );
and ( \607_SUM[15]_b1 , w_1062 , w_1052 );
and ( w_1061 , \597_b0 , w_1053 );
and ( \608_b1 , \608_b0 , w_1054 );
and ( w_1059 , w_1063 , \241_b1 );
or ( w_1046 , w_1047 , w_1055 );
or ( w_1055 , w_1049 , \241_b0 );
or ( w_1050 , w_1051 , w_1056 );
or ( w_1056 , w_1052 , w_1057 );
or ( w_1057 , w_1053 , w_1058 );
or ( w_1058 , w_1054 , w_1059 );
not ( \607_SUM[15]_b1 , w_1060 );
not ( \607_SUM[15]_b0 , w_1061 );
not ( \608_b1 , w_1062 );
not ( \241_b0 , w_1063 );
buf ( \609_A[15]_b1 , \c[15]_b1 );
buf ( \609_A[15]_b0 , \c[15]_b0 );
buf ( \610_B[15]_b1 , \d[15]_b1 );
buf ( \610_B[15]_b0 , \d[15]_b0 );
or ( \611_b1 , \609_A[15]_b1 , \610_B[15]_b1 );
xor ( \611_b0 , \609_A[15]_b0 , w_1064 );
not ( w_1064 , w_1065 );
and ( w_1065 , \610_B[15]_b1 , \610_B[15]_b0 );
or ( \612_b1 , \586_A[14]_b1 , \587_B[14]_b1 );
not ( \587_B[14]_b1 , w_1066 );
and ( \612_b0 , \586_A[14]_b0 , w_1067 );
and ( w_1066 , w_1067 , \587_B[14]_b0 );
or ( \613_b1 , \587_B[14]_b1 , \592_b1 );
not ( \592_b1 , w_1068 );
and ( \613_b0 , \587_B[14]_b0 , w_1069 );
and ( w_1068 , w_1069 , \592_b0 );
or ( \614_b1 , \586_A[14]_b1 , \592_b1 );
not ( \592_b1 , w_1070 );
and ( \614_b0 , \586_A[14]_b0 , w_1071 );
and ( w_1070 , w_1071 , \592_b0 );
or ( \616_b1 , \611_b1 , \615_b1 );
xor ( \616_b0 , \611_b0 , w_1072 );
not ( w_1072 , w_1073 );
and ( w_1073 , \615_b1 , \615_b0 );
buf ( \617_SUM[15]_b1 , \616_b1 );
buf ( \617_SUM[15]_b0 , \616_b0 );
and ( \618_b0 , \617_SUM[15]_b0 , w_1074 );
and ( \618_b0 , \608_b0 , w_1075 );
and ( w_1088 , w_1089 , w_1076 );
and ( w_1076 , \608_b0 , w_1077 );
and ( w_1089 , \608_b1 , w_1078 );
and ( \618_b1 , \617_SUM[15]_b0 , w_1079 );
and ( \617_SUM[15]_b1 , w_1090 , w_1080 );
and ( w_1089 , \608_b0 , w_1081 );
and ( \618_b1 , \618_b0 , w_1082 );
and ( w_1087 , w_1091 , \277_b1 );
or ( w_1074 , w_1075 , w_1083 );
or ( w_1083 , w_1077 , \277_b0 );
or ( w_1078 , w_1079 , w_1084 );
or ( w_1084 , w_1080 , w_1085 );
or ( w_1085 , w_1081 , w_1086 );
or ( w_1086 , w_1082 , w_1087 );
not ( \617_SUM[15]_b1 , w_1088 );
not ( \617_SUM[15]_b0 , w_1089 );
not ( \618_b1 , w_1090 );
not ( \277_b0 , w_1091 );
and ( \619_n5[16]_b1 , 1'b0_b1 , w_1092 );
xor ( w_1092 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1093 );
and ( \619_n5[16]_b0 , w_1093 , 1'b1_b0 );
or ( \620_b1 , \b[16]_b1 , w_1094 );
or ( \620_b0 , \b[16]_b0 , \619_n5[16]_b0 );
not ( \619_n5[16]_b0 , w_1095 );
and ( w_1095 , w_1094 , \619_n5[16]_b1 );
buf ( \621_A[16]_b1 , \c[16]_b1 );
buf ( \621_A[16]_b0 , \c[16]_b0 );
buf ( \622_B[16]_b1 , \d[16]_b1 );
buf ( \622_B[16]_b0 , \d[16]_b0 );
buf ( \623_b1 , \622_B[16]_b1 );
not ( \623_b1 , w_1096 );
not ( \623_b0 , w_1097 );
and ( w_1096 , w_1097 , \622_B[16]_b0 );
or ( \624_b1 , \621_A[16]_b1 , \623_b1 );
xor ( \624_b0 , \621_A[16]_b0 , w_1098 );
not ( w_1098 , w_1099 );
and ( w_1099 , \623_b1 , \623_b0 );
or ( \625_b1 , \598_A[15]_b1 , \600_b1 );
not ( \600_b1 , w_1100 );
and ( \625_b0 , \598_A[15]_b0 , w_1101 );
and ( w_1100 , w_1101 , \600_b0 );
or ( \626_b1 , \600_b1 , \605_b1 );
not ( \605_b1 , w_1102 );
and ( \626_b0 , \600_b0 , w_1103 );
and ( w_1102 , w_1103 , \605_b0 );
or ( \627_b1 , \598_A[15]_b1 , \605_b1 );
not ( \605_b1 , w_1104 );
and ( \627_b0 , \598_A[15]_b0 , w_1105 );
and ( w_1104 , w_1105 , \605_b0 );
or ( \629_b1 , \624_b1 , \628_b1 );
xor ( \629_b0 , \624_b0 , w_1106 );
not ( w_1106 , w_1107 );
and ( w_1107 , \628_b1 , \628_b0 );
buf ( \630_SUM[16]_b1 , \629_b1 );
buf ( \630_SUM[16]_b0 , \629_b0 );
and ( \631_b0 , \630_SUM[16]_b0 , w_1108 );
and ( \631_b0 , \620_b0 , w_1109 );
and ( w_1122 , w_1123 , w_1110 );
and ( w_1110 , \620_b0 , w_1111 );
and ( w_1123 , \620_b1 , w_1112 );
and ( \631_b1 , \630_SUM[16]_b0 , w_1113 );
and ( \630_SUM[16]_b1 , w_1124 , w_1114 );
and ( w_1123 , \620_b0 , w_1115 );
and ( \631_b1 , \631_b0 , w_1116 );
and ( w_1121 , w_1125 , \241_b1 );
or ( w_1108 , w_1109 , w_1117 );
or ( w_1117 , w_1111 , \241_b0 );
or ( w_1112 , w_1113 , w_1118 );
or ( w_1118 , w_1114 , w_1119 );
or ( w_1119 , w_1115 , w_1120 );
or ( w_1120 , w_1116 , w_1121 );
not ( \630_SUM[16]_b1 , w_1122 );
not ( \630_SUM[16]_b0 , w_1123 );
not ( \631_b1 , w_1124 );
not ( \241_b0 , w_1125 );
buf ( \632_A[16]_b1 , \c[16]_b1 );
buf ( \632_A[16]_b0 , \c[16]_b0 );
buf ( \633_B[16]_b1 , \d[16]_b1 );
buf ( \633_B[16]_b0 , \d[16]_b0 );
or ( \634_b1 , \632_A[16]_b1 , \633_B[16]_b1 );
xor ( \634_b0 , \632_A[16]_b0 , w_1126 );
not ( w_1126 , w_1127 );
and ( w_1127 , \633_B[16]_b1 , \633_B[16]_b0 );
or ( \635_b1 , \609_A[15]_b1 , \610_B[15]_b1 );
not ( \610_B[15]_b1 , w_1128 );
and ( \635_b0 , \609_A[15]_b0 , w_1129 );
and ( w_1128 , w_1129 , \610_B[15]_b0 );
or ( \636_b1 , \610_B[15]_b1 , \615_b1 );
not ( \615_b1 , w_1130 );
and ( \636_b0 , \610_B[15]_b0 , w_1131 );
and ( w_1130 , w_1131 , \615_b0 );
or ( \637_b1 , \609_A[15]_b1 , \615_b1 );
not ( \615_b1 , w_1132 );
and ( \637_b0 , \609_A[15]_b0 , w_1133 );
and ( w_1132 , w_1133 , \615_b0 );
or ( \639_b1 , \634_b1 , \638_b1 );
xor ( \639_b0 , \634_b0 , w_1134 );
not ( w_1134 , w_1135 );
and ( w_1135 , \638_b1 , \638_b0 );
buf ( \640_SUM[16]_b1 , \639_b1 );
buf ( \640_SUM[16]_b0 , \639_b0 );
and ( \641_b0 , \640_SUM[16]_b0 , w_1136 );
and ( \641_b0 , \631_b0 , w_1137 );
and ( w_1150 , w_1151 , w_1138 );
and ( w_1138 , \631_b0 , w_1139 );
and ( w_1151 , \631_b1 , w_1140 );
and ( \641_b1 , \640_SUM[16]_b0 , w_1141 );
and ( \640_SUM[16]_b1 , w_1152 , w_1142 );
and ( w_1151 , \631_b0 , w_1143 );
and ( \641_b1 , \641_b0 , w_1144 );
and ( w_1149 , w_1153 , \277_b1 );
or ( w_1136 , w_1137 , w_1145 );
or ( w_1145 , w_1139 , \277_b0 );
or ( w_1140 , w_1141 , w_1146 );
or ( w_1146 , w_1142 , w_1147 );
or ( w_1147 , w_1143 , w_1148 );
or ( w_1148 , w_1144 , w_1149 );
not ( \640_SUM[16]_b1 , w_1150 );
not ( \640_SUM[16]_b0 , w_1151 );
not ( \641_b1 , w_1152 );
not ( \277_b0 , w_1153 );
and ( \642_n5[17]_b1 , 1'b0_b1 , w_1154 );
xor ( w_1154 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1155 );
and ( \642_n5[17]_b0 , w_1155 , 1'b1_b0 );
or ( \643_b1 , \b[17]_b1 , w_1156 );
or ( \643_b0 , \b[17]_b0 , \642_n5[17]_b0 );
not ( \642_n5[17]_b0 , w_1157 );
and ( w_1157 , w_1156 , \642_n5[17]_b1 );
buf ( \644_A[17]_b1 , \c[17]_b1 );
buf ( \644_A[17]_b0 , \c[17]_b0 );
buf ( \645_B[17]_b1 , \d[17]_b1 );
buf ( \645_B[17]_b0 , \d[17]_b0 );
buf ( \646_b1 , \645_B[17]_b1 );
not ( \646_b1 , w_1158 );
not ( \646_b0 , w_1159 );
and ( w_1158 , w_1159 , \645_B[17]_b0 );
or ( \647_b1 , \644_A[17]_b1 , \646_b1 );
xor ( \647_b0 , \644_A[17]_b0 , w_1160 );
not ( w_1160 , w_1161 );
and ( w_1161 , \646_b1 , \646_b0 );
or ( \648_b1 , \621_A[16]_b1 , \623_b1 );
not ( \623_b1 , w_1162 );
and ( \648_b0 , \621_A[16]_b0 , w_1163 );
and ( w_1162 , w_1163 , \623_b0 );
or ( \649_b1 , \623_b1 , \628_b1 );
not ( \628_b1 , w_1164 );
and ( \649_b0 , \623_b0 , w_1165 );
and ( w_1164 , w_1165 , \628_b0 );
or ( \650_b1 , \621_A[16]_b1 , \628_b1 );
not ( \628_b1 , w_1166 );
and ( \650_b0 , \621_A[16]_b0 , w_1167 );
and ( w_1166 , w_1167 , \628_b0 );
or ( \652_b1 , \647_b1 , \651_b1 );
xor ( \652_b0 , \647_b0 , w_1168 );
not ( w_1168 , w_1169 );
and ( w_1169 , \651_b1 , \651_b0 );
buf ( \653_SUM[17]_b1 , \652_b1 );
buf ( \653_SUM[17]_b0 , \652_b0 );
and ( \654_b0 , \653_SUM[17]_b0 , w_1170 );
and ( \654_b0 , \643_b0 , w_1171 );
and ( w_1184 , w_1185 , w_1172 );
and ( w_1172 , \643_b0 , w_1173 );
and ( w_1185 , \643_b1 , w_1174 );
and ( \654_b1 , \653_SUM[17]_b0 , w_1175 );
and ( \653_SUM[17]_b1 , w_1186 , w_1176 );
and ( w_1185 , \643_b0 , w_1177 );
and ( \654_b1 , \654_b0 , w_1178 );
and ( w_1183 , w_1187 , \241_b1 );
or ( w_1170 , w_1171 , w_1179 );
or ( w_1179 , w_1173 , \241_b0 );
or ( w_1174 , w_1175 , w_1180 );
or ( w_1180 , w_1176 , w_1181 );
or ( w_1181 , w_1177 , w_1182 );
or ( w_1182 , w_1178 , w_1183 );
not ( \653_SUM[17]_b1 , w_1184 );
not ( \653_SUM[17]_b0 , w_1185 );
not ( \654_b1 , w_1186 );
not ( \241_b0 , w_1187 );
buf ( \655_A[17]_b1 , \c[17]_b1 );
buf ( \655_A[17]_b0 , \c[17]_b0 );
buf ( \656_B[17]_b1 , \d[17]_b1 );
buf ( \656_B[17]_b0 , \d[17]_b0 );
or ( \657_b1 , \655_A[17]_b1 , \656_B[17]_b1 );
xor ( \657_b0 , \655_A[17]_b0 , w_1188 );
not ( w_1188 , w_1189 );
and ( w_1189 , \656_B[17]_b1 , \656_B[17]_b0 );
or ( \658_b1 , \632_A[16]_b1 , \633_B[16]_b1 );
not ( \633_B[16]_b1 , w_1190 );
and ( \658_b0 , \632_A[16]_b0 , w_1191 );
and ( w_1190 , w_1191 , \633_B[16]_b0 );
or ( \659_b1 , \633_B[16]_b1 , \638_b1 );
not ( \638_b1 , w_1192 );
and ( \659_b0 , \633_B[16]_b0 , w_1193 );
and ( w_1192 , w_1193 , \638_b0 );
or ( \660_b1 , \632_A[16]_b1 , \638_b1 );
not ( \638_b1 , w_1194 );
and ( \660_b0 , \632_A[16]_b0 , w_1195 );
and ( w_1194 , w_1195 , \638_b0 );
or ( \662_b1 , \657_b1 , \661_b1 );
xor ( \662_b0 , \657_b0 , w_1196 );
not ( w_1196 , w_1197 );
and ( w_1197 , \661_b1 , \661_b0 );
buf ( \663_SUM[17]_b1 , \662_b1 );
buf ( \663_SUM[17]_b0 , \662_b0 );
and ( \664_b0 , \663_SUM[17]_b0 , w_1198 );
and ( \664_b0 , \654_b0 , w_1199 );
and ( w_1212 , w_1213 , w_1200 );
and ( w_1200 , \654_b0 , w_1201 );
and ( w_1213 , \654_b1 , w_1202 );
and ( \664_b1 , \663_SUM[17]_b0 , w_1203 );
and ( \663_SUM[17]_b1 , w_1214 , w_1204 );
and ( w_1213 , \654_b0 , w_1205 );
and ( \664_b1 , \664_b0 , w_1206 );
and ( w_1211 , w_1215 , \277_b1 );
or ( w_1198 , w_1199 , w_1207 );
or ( w_1207 , w_1201 , \277_b0 );
or ( w_1202 , w_1203 , w_1208 );
or ( w_1208 , w_1204 , w_1209 );
or ( w_1209 , w_1205 , w_1210 );
or ( w_1210 , w_1206 , w_1211 );
not ( \663_SUM[17]_b1 , w_1212 );
not ( \663_SUM[17]_b0 , w_1213 );
not ( \664_b1 , w_1214 );
not ( \277_b0 , w_1215 );
and ( \665_n5[18]_b1 , 1'b0_b1 , w_1216 );
xor ( w_1216 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1217 );
and ( \665_n5[18]_b0 , w_1217 , 1'b1_b0 );
or ( \666_b1 , \b[18]_b1 , w_1218 );
or ( \666_b0 , \b[18]_b0 , \665_n5[18]_b0 );
not ( \665_n5[18]_b0 , w_1219 );
and ( w_1219 , w_1218 , \665_n5[18]_b1 );
buf ( \667_A[18]_b1 , \c[18]_b1 );
buf ( \667_A[18]_b0 , \c[18]_b0 );
buf ( \668_B[18]_b1 , \d[18]_b1 );
buf ( \668_B[18]_b0 , \d[18]_b0 );
buf ( \669_b1 , \668_B[18]_b1 );
not ( \669_b1 , w_1220 );
not ( \669_b0 , w_1221 );
and ( w_1220 , w_1221 , \668_B[18]_b0 );
or ( \670_b1 , \667_A[18]_b1 , \669_b1 );
xor ( \670_b0 , \667_A[18]_b0 , w_1222 );
not ( w_1222 , w_1223 );
and ( w_1223 , \669_b1 , \669_b0 );
or ( \671_b1 , \644_A[17]_b1 , \646_b1 );
not ( \646_b1 , w_1224 );
and ( \671_b0 , \644_A[17]_b0 , w_1225 );
and ( w_1224 , w_1225 , \646_b0 );
or ( \672_b1 , \646_b1 , \651_b1 );
not ( \651_b1 , w_1226 );
and ( \672_b0 , \646_b0 , w_1227 );
and ( w_1226 , w_1227 , \651_b0 );
or ( \673_b1 , \644_A[17]_b1 , \651_b1 );
not ( \651_b1 , w_1228 );
and ( \673_b0 , \644_A[17]_b0 , w_1229 );
and ( w_1228 , w_1229 , \651_b0 );
or ( \675_b1 , \670_b1 , \674_b1 );
xor ( \675_b0 , \670_b0 , w_1230 );
not ( w_1230 , w_1231 );
and ( w_1231 , \674_b1 , \674_b0 );
buf ( \676_SUM[18]_b1 , \675_b1 );
buf ( \676_SUM[18]_b0 , \675_b0 );
and ( \677_b0 , \676_SUM[18]_b0 , w_1232 );
and ( \677_b0 , \666_b0 , w_1233 );
and ( w_1246 , w_1247 , w_1234 );
and ( w_1234 , \666_b0 , w_1235 );
and ( w_1247 , \666_b1 , w_1236 );
and ( \677_b1 , \676_SUM[18]_b0 , w_1237 );
and ( \676_SUM[18]_b1 , w_1248 , w_1238 );
and ( w_1247 , \666_b0 , w_1239 );
and ( \677_b1 , \677_b0 , w_1240 );
and ( w_1245 , w_1249 , \241_b1 );
or ( w_1232 , w_1233 , w_1241 );
or ( w_1241 , w_1235 , \241_b0 );
or ( w_1236 , w_1237 , w_1242 );
or ( w_1242 , w_1238 , w_1243 );
or ( w_1243 , w_1239 , w_1244 );
or ( w_1244 , w_1240 , w_1245 );
not ( \676_SUM[18]_b1 , w_1246 );
not ( \676_SUM[18]_b0 , w_1247 );
not ( \677_b1 , w_1248 );
not ( \241_b0 , w_1249 );
buf ( \678_A[18]_b1 , \c[18]_b1 );
buf ( \678_A[18]_b0 , \c[18]_b0 );
buf ( \679_B[18]_b1 , \d[18]_b1 );
buf ( \679_B[18]_b0 , \d[18]_b0 );
or ( \680_b1 , \678_A[18]_b1 , \679_B[18]_b1 );
xor ( \680_b0 , \678_A[18]_b0 , w_1250 );
not ( w_1250 , w_1251 );
and ( w_1251 , \679_B[18]_b1 , \679_B[18]_b0 );
or ( \681_b1 , \655_A[17]_b1 , \656_B[17]_b1 );
not ( \656_B[17]_b1 , w_1252 );
and ( \681_b0 , \655_A[17]_b0 , w_1253 );
and ( w_1252 , w_1253 , \656_B[17]_b0 );
or ( \682_b1 , \656_B[17]_b1 , \661_b1 );
not ( \661_b1 , w_1254 );
and ( \682_b0 , \656_B[17]_b0 , w_1255 );
and ( w_1254 , w_1255 , \661_b0 );
or ( \683_b1 , \655_A[17]_b1 , \661_b1 );
not ( \661_b1 , w_1256 );
and ( \683_b0 , \655_A[17]_b0 , w_1257 );
and ( w_1256 , w_1257 , \661_b0 );
or ( \685_b1 , \680_b1 , \684_b1 );
xor ( \685_b0 , \680_b0 , w_1258 );
not ( w_1258 , w_1259 );
and ( w_1259 , \684_b1 , \684_b0 );
buf ( \686_SUM[18]_b1 , \685_b1 );
buf ( \686_SUM[18]_b0 , \685_b0 );
and ( \687_b0 , \686_SUM[18]_b0 , w_1260 );
and ( \687_b0 , \677_b0 , w_1261 );
and ( w_1274 , w_1275 , w_1262 );
and ( w_1262 , \677_b0 , w_1263 );
and ( w_1275 , \677_b1 , w_1264 );
and ( \687_b1 , \686_SUM[18]_b0 , w_1265 );
and ( \686_SUM[18]_b1 , w_1276 , w_1266 );
and ( w_1275 , \677_b0 , w_1267 );
and ( \687_b1 , \687_b0 , w_1268 );
and ( w_1273 , w_1277 , \277_b1 );
or ( w_1260 , w_1261 , w_1269 );
or ( w_1269 , w_1263 , \277_b0 );
or ( w_1264 , w_1265 , w_1270 );
or ( w_1270 , w_1266 , w_1271 );
or ( w_1271 , w_1267 , w_1272 );
or ( w_1272 , w_1268 , w_1273 );
not ( \686_SUM[18]_b1 , w_1274 );
not ( \686_SUM[18]_b0 , w_1275 );
not ( \687_b1 , w_1276 );
not ( \277_b0 , w_1277 );
and ( \688_n5[19]_b1 , 1'b0_b1 , w_1278 );
xor ( w_1278 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1279 );
and ( \688_n5[19]_b0 , w_1279 , 1'b1_b0 );
or ( \689_b1 , \b[19]_b1 , w_1280 );
or ( \689_b0 , \b[19]_b0 , \688_n5[19]_b0 );
not ( \688_n5[19]_b0 , w_1281 );
and ( w_1281 , w_1280 , \688_n5[19]_b1 );
buf ( \690_A[19]_b1 , \c[19]_b1 );
buf ( \690_A[19]_b0 , \c[19]_b0 );
buf ( \691_B[19]_b1 , \d[19]_b1 );
buf ( \691_B[19]_b0 , \d[19]_b0 );
buf ( \692_b1 , \691_B[19]_b1 );
not ( \692_b1 , w_1282 );
not ( \692_b0 , w_1283 );
and ( w_1282 , w_1283 , \691_B[19]_b0 );
or ( \693_b1 , \690_A[19]_b1 , \692_b1 );
xor ( \693_b0 , \690_A[19]_b0 , w_1284 );
not ( w_1284 , w_1285 );
and ( w_1285 , \692_b1 , \692_b0 );
or ( \694_b1 , \667_A[18]_b1 , \669_b1 );
not ( \669_b1 , w_1286 );
and ( \694_b0 , \667_A[18]_b0 , w_1287 );
and ( w_1286 , w_1287 , \669_b0 );
or ( \695_b1 , \669_b1 , \674_b1 );
not ( \674_b1 , w_1288 );
and ( \695_b0 , \669_b0 , w_1289 );
and ( w_1288 , w_1289 , \674_b0 );
or ( \696_b1 , \667_A[18]_b1 , \674_b1 );
not ( \674_b1 , w_1290 );
and ( \696_b0 , \667_A[18]_b0 , w_1291 );
and ( w_1290 , w_1291 , \674_b0 );
or ( \698_b1 , \693_b1 , \697_b1 );
xor ( \698_b0 , \693_b0 , w_1292 );
not ( w_1292 , w_1293 );
and ( w_1293 , \697_b1 , \697_b0 );
buf ( \699_SUM[19]_b1 , \698_b1 );
buf ( \699_SUM[19]_b0 , \698_b0 );
and ( \700_b0 , \699_SUM[19]_b0 , w_1294 );
and ( \700_b0 , \689_b0 , w_1295 );
and ( w_1308 , w_1309 , w_1296 );
and ( w_1296 , \689_b0 , w_1297 );
and ( w_1309 , \689_b1 , w_1298 );
and ( \700_b1 , \699_SUM[19]_b0 , w_1299 );
and ( \699_SUM[19]_b1 , w_1310 , w_1300 );
and ( w_1309 , \689_b0 , w_1301 );
and ( \700_b1 , \700_b0 , w_1302 );
and ( w_1307 , w_1311 , \241_b1 );
or ( w_1294 , w_1295 , w_1303 );
or ( w_1303 , w_1297 , \241_b0 );
or ( w_1298 , w_1299 , w_1304 );
or ( w_1304 , w_1300 , w_1305 );
or ( w_1305 , w_1301 , w_1306 );
or ( w_1306 , w_1302 , w_1307 );
not ( \699_SUM[19]_b1 , w_1308 );
not ( \699_SUM[19]_b0 , w_1309 );
not ( \700_b1 , w_1310 );
not ( \241_b0 , w_1311 );
buf ( \701_A[19]_b1 , \c[19]_b1 );
buf ( \701_A[19]_b0 , \c[19]_b0 );
buf ( \702_B[19]_b1 , \d[19]_b1 );
buf ( \702_B[19]_b0 , \d[19]_b0 );
or ( \703_b1 , \701_A[19]_b1 , \702_B[19]_b1 );
xor ( \703_b0 , \701_A[19]_b0 , w_1312 );
not ( w_1312 , w_1313 );
and ( w_1313 , \702_B[19]_b1 , \702_B[19]_b0 );
or ( \704_b1 , \678_A[18]_b1 , \679_B[18]_b1 );
not ( \679_B[18]_b1 , w_1314 );
and ( \704_b0 , \678_A[18]_b0 , w_1315 );
and ( w_1314 , w_1315 , \679_B[18]_b0 );
or ( \705_b1 , \679_B[18]_b1 , \684_b1 );
not ( \684_b1 , w_1316 );
and ( \705_b0 , \679_B[18]_b0 , w_1317 );
and ( w_1316 , w_1317 , \684_b0 );
or ( \706_b1 , \678_A[18]_b1 , \684_b1 );
not ( \684_b1 , w_1318 );
and ( \706_b0 , \678_A[18]_b0 , w_1319 );
and ( w_1318 , w_1319 , \684_b0 );
or ( \708_b1 , \703_b1 , \707_b1 );
xor ( \708_b0 , \703_b0 , w_1320 );
not ( w_1320 , w_1321 );
and ( w_1321 , \707_b1 , \707_b0 );
buf ( \709_SUM[19]_b1 , \708_b1 );
buf ( \709_SUM[19]_b0 , \708_b0 );
and ( \710_b0 , \709_SUM[19]_b0 , w_1322 );
and ( \710_b0 , \700_b0 , w_1323 );
and ( w_1336 , w_1337 , w_1324 );
and ( w_1324 , \700_b0 , w_1325 );
and ( w_1337 , \700_b1 , w_1326 );
and ( \710_b1 , \709_SUM[19]_b0 , w_1327 );
and ( \709_SUM[19]_b1 , w_1338 , w_1328 );
and ( w_1337 , \700_b0 , w_1329 );
and ( \710_b1 , \710_b0 , w_1330 );
and ( w_1335 , w_1339 , \277_b1 );
or ( w_1322 , w_1323 , w_1331 );
or ( w_1331 , w_1325 , \277_b0 );
or ( w_1326 , w_1327 , w_1332 );
or ( w_1332 , w_1328 , w_1333 );
or ( w_1333 , w_1329 , w_1334 );
or ( w_1334 , w_1330 , w_1335 );
not ( \709_SUM[19]_b1 , w_1336 );
not ( \709_SUM[19]_b0 , w_1337 );
not ( \710_b1 , w_1338 );
not ( \277_b0 , w_1339 );
and ( \711_n5[20]_b1 , 1'b0_b1 , w_1340 );
xor ( w_1340 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1341 );
and ( \711_n5[20]_b0 , w_1341 , 1'b1_b0 );
or ( \712_b1 , \b[20]_b1 , w_1342 );
or ( \712_b0 , \b[20]_b0 , \711_n5[20]_b0 );
not ( \711_n5[20]_b0 , w_1343 );
and ( w_1343 , w_1342 , \711_n5[20]_b1 );
buf ( \713_A[20]_b1 , \c[20]_b1 );
buf ( \713_A[20]_b0 , \c[20]_b0 );
buf ( \714_B[20]_b1 , \d[20]_b1 );
buf ( \714_B[20]_b0 , \d[20]_b0 );
buf ( \715_b1 , \714_B[20]_b1 );
not ( \715_b1 , w_1344 );
not ( \715_b0 , w_1345 );
and ( w_1344 , w_1345 , \714_B[20]_b0 );
or ( \716_b1 , \713_A[20]_b1 , \715_b1 );
xor ( \716_b0 , \713_A[20]_b0 , w_1346 );
not ( w_1346 , w_1347 );
and ( w_1347 , \715_b1 , \715_b0 );
or ( \717_b1 , \690_A[19]_b1 , \692_b1 );
not ( \692_b1 , w_1348 );
and ( \717_b0 , \690_A[19]_b0 , w_1349 );
and ( w_1348 , w_1349 , \692_b0 );
or ( \718_b1 , \692_b1 , \697_b1 );
not ( \697_b1 , w_1350 );
and ( \718_b0 , \692_b0 , w_1351 );
and ( w_1350 , w_1351 , \697_b0 );
or ( \719_b1 , \690_A[19]_b1 , \697_b1 );
not ( \697_b1 , w_1352 );
and ( \719_b0 , \690_A[19]_b0 , w_1353 );
and ( w_1352 , w_1353 , \697_b0 );
or ( \721_b1 , \716_b1 , \720_b1 );
xor ( \721_b0 , \716_b0 , w_1354 );
not ( w_1354 , w_1355 );
and ( w_1355 , \720_b1 , \720_b0 );
buf ( \722_SUM[20]_b1 , \721_b1 );
buf ( \722_SUM[20]_b0 , \721_b0 );
and ( \723_b0 , \722_SUM[20]_b0 , w_1356 );
and ( \723_b0 , \712_b0 , w_1357 );
and ( w_1370 , w_1371 , w_1358 );
and ( w_1358 , \712_b0 , w_1359 );
and ( w_1371 , \712_b1 , w_1360 );
and ( \723_b1 , \722_SUM[20]_b0 , w_1361 );
and ( \722_SUM[20]_b1 , w_1372 , w_1362 );
and ( w_1371 , \712_b0 , w_1363 );
and ( \723_b1 , \723_b0 , w_1364 );
and ( w_1369 , w_1373 , \241_b1 );
or ( w_1356 , w_1357 , w_1365 );
or ( w_1365 , w_1359 , \241_b0 );
or ( w_1360 , w_1361 , w_1366 );
or ( w_1366 , w_1362 , w_1367 );
or ( w_1367 , w_1363 , w_1368 );
or ( w_1368 , w_1364 , w_1369 );
not ( \722_SUM[20]_b1 , w_1370 );
not ( \722_SUM[20]_b0 , w_1371 );
not ( \723_b1 , w_1372 );
not ( \241_b0 , w_1373 );
buf ( \724_A[20]_b1 , \c[20]_b1 );
buf ( \724_A[20]_b0 , \c[20]_b0 );
buf ( \725_B[20]_b1 , \d[20]_b1 );
buf ( \725_B[20]_b0 , \d[20]_b0 );
or ( \726_b1 , \724_A[20]_b1 , \725_B[20]_b1 );
xor ( \726_b0 , \724_A[20]_b0 , w_1374 );
not ( w_1374 , w_1375 );
and ( w_1375 , \725_B[20]_b1 , \725_B[20]_b0 );
or ( \727_b1 , \701_A[19]_b1 , \702_B[19]_b1 );
not ( \702_B[19]_b1 , w_1376 );
and ( \727_b0 , \701_A[19]_b0 , w_1377 );
and ( w_1376 , w_1377 , \702_B[19]_b0 );
or ( \728_b1 , \702_B[19]_b1 , \707_b1 );
not ( \707_b1 , w_1378 );
and ( \728_b0 , \702_B[19]_b0 , w_1379 );
and ( w_1378 , w_1379 , \707_b0 );
or ( \729_b1 , \701_A[19]_b1 , \707_b1 );
not ( \707_b1 , w_1380 );
and ( \729_b0 , \701_A[19]_b0 , w_1381 );
and ( w_1380 , w_1381 , \707_b0 );
or ( \731_b1 , \726_b1 , \730_b1 );
xor ( \731_b0 , \726_b0 , w_1382 );
not ( w_1382 , w_1383 );
and ( w_1383 , \730_b1 , \730_b0 );
buf ( \732_SUM[20]_b1 , \731_b1 );
buf ( \732_SUM[20]_b0 , \731_b0 );
and ( \733_b0 , \732_SUM[20]_b0 , w_1384 );
and ( \733_b0 , \723_b0 , w_1385 );
and ( w_1398 , w_1399 , w_1386 );
and ( w_1386 , \723_b0 , w_1387 );
and ( w_1399 , \723_b1 , w_1388 );
and ( \733_b1 , \732_SUM[20]_b0 , w_1389 );
and ( \732_SUM[20]_b1 , w_1400 , w_1390 );
and ( w_1399 , \723_b0 , w_1391 );
and ( \733_b1 , \733_b0 , w_1392 );
and ( w_1397 , w_1401 , \277_b1 );
or ( w_1384 , w_1385 , w_1393 );
or ( w_1393 , w_1387 , \277_b0 );
or ( w_1388 , w_1389 , w_1394 );
or ( w_1394 , w_1390 , w_1395 );
or ( w_1395 , w_1391 , w_1396 );
or ( w_1396 , w_1392 , w_1397 );
not ( \732_SUM[20]_b1 , w_1398 );
not ( \732_SUM[20]_b0 , w_1399 );
not ( \733_b1 , w_1400 );
not ( \277_b0 , w_1401 );
and ( \734_n5[21]_b1 , 1'b0_b1 , w_1402 );
xor ( w_1402 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1403 );
and ( \734_n5[21]_b0 , w_1403 , 1'b1_b0 );
or ( \735_b1 , \b[21]_b1 , w_1404 );
or ( \735_b0 , \b[21]_b0 , \734_n5[21]_b0 );
not ( \734_n5[21]_b0 , w_1405 );
and ( w_1405 , w_1404 , \734_n5[21]_b1 );
buf ( \736_A[21]_b1 , \c[21]_b1 );
buf ( \736_A[21]_b0 , \c[21]_b0 );
buf ( \737_B[21]_b1 , \d[21]_b1 );
buf ( \737_B[21]_b0 , \d[21]_b0 );
buf ( \738_b1 , \737_B[21]_b1 );
not ( \738_b1 , w_1406 );
not ( \738_b0 , w_1407 );
and ( w_1406 , w_1407 , \737_B[21]_b0 );
or ( \739_b1 , \736_A[21]_b1 , \738_b1 );
xor ( \739_b0 , \736_A[21]_b0 , w_1408 );
not ( w_1408 , w_1409 );
and ( w_1409 , \738_b1 , \738_b0 );
or ( \740_b1 , \713_A[20]_b1 , \715_b1 );
not ( \715_b1 , w_1410 );
and ( \740_b0 , \713_A[20]_b0 , w_1411 );
and ( w_1410 , w_1411 , \715_b0 );
or ( \741_b1 , \715_b1 , \720_b1 );
not ( \720_b1 , w_1412 );
and ( \741_b0 , \715_b0 , w_1413 );
and ( w_1412 , w_1413 , \720_b0 );
or ( \742_b1 , \713_A[20]_b1 , \720_b1 );
not ( \720_b1 , w_1414 );
and ( \742_b0 , \713_A[20]_b0 , w_1415 );
and ( w_1414 , w_1415 , \720_b0 );
or ( \744_b1 , \739_b1 , \743_b1 );
xor ( \744_b0 , \739_b0 , w_1416 );
not ( w_1416 , w_1417 );
and ( w_1417 , \743_b1 , \743_b0 );
buf ( \745_SUM[21]_b1 , \744_b1 );
buf ( \745_SUM[21]_b0 , \744_b0 );
and ( \746_b0 , \745_SUM[21]_b0 , w_1418 );
and ( \746_b0 , \735_b0 , w_1419 );
and ( w_1432 , w_1433 , w_1420 );
and ( w_1420 , \735_b0 , w_1421 );
and ( w_1433 , \735_b1 , w_1422 );
and ( \746_b1 , \745_SUM[21]_b0 , w_1423 );
and ( \745_SUM[21]_b1 , w_1434 , w_1424 );
and ( w_1433 , \735_b0 , w_1425 );
and ( \746_b1 , \746_b0 , w_1426 );
and ( w_1431 , w_1435 , \241_b1 );
or ( w_1418 , w_1419 , w_1427 );
or ( w_1427 , w_1421 , \241_b0 );
or ( w_1422 , w_1423 , w_1428 );
or ( w_1428 , w_1424 , w_1429 );
or ( w_1429 , w_1425 , w_1430 );
or ( w_1430 , w_1426 , w_1431 );
not ( \745_SUM[21]_b1 , w_1432 );
not ( \745_SUM[21]_b0 , w_1433 );
not ( \746_b1 , w_1434 );
not ( \241_b0 , w_1435 );
buf ( \747_A[21]_b1 , \c[21]_b1 );
buf ( \747_A[21]_b0 , \c[21]_b0 );
buf ( \748_B[21]_b1 , \d[21]_b1 );
buf ( \748_B[21]_b0 , \d[21]_b0 );
or ( \749_b1 , \747_A[21]_b1 , \748_B[21]_b1 );
xor ( \749_b0 , \747_A[21]_b0 , w_1436 );
not ( w_1436 , w_1437 );
and ( w_1437 , \748_B[21]_b1 , \748_B[21]_b0 );
or ( \750_b1 , \724_A[20]_b1 , \725_B[20]_b1 );
not ( \725_B[20]_b1 , w_1438 );
and ( \750_b0 , \724_A[20]_b0 , w_1439 );
and ( w_1438 , w_1439 , \725_B[20]_b0 );
or ( \751_b1 , \725_B[20]_b1 , \730_b1 );
not ( \730_b1 , w_1440 );
and ( \751_b0 , \725_B[20]_b0 , w_1441 );
and ( w_1440 , w_1441 , \730_b0 );
or ( \752_b1 , \724_A[20]_b1 , \730_b1 );
not ( \730_b1 , w_1442 );
and ( \752_b0 , \724_A[20]_b0 , w_1443 );
and ( w_1442 , w_1443 , \730_b0 );
or ( \754_b1 , \749_b1 , \753_b1 );
xor ( \754_b0 , \749_b0 , w_1444 );
not ( w_1444 , w_1445 );
and ( w_1445 , \753_b1 , \753_b0 );
buf ( \755_SUM[21]_b1 , \754_b1 );
buf ( \755_SUM[21]_b0 , \754_b0 );
and ( \756_b0 , \755_SUM[21]_b0 , w_1446 );
and ( \756_b0 , \746_b0 , w_1447 );
and ( w_1460 , w_1461 , w_1448 );
and ( w_1448 , \746_b0 , w_1449 );
and ( w_1461 , \746_b1 , w_1450 );
and ( \756_b1 , \755_SUM[21]_b0 , w_1451 );
and ( \755_SUM[21]_b1 , w_1462 , w_1452 );
and ( w_1461 , \746_b0 , w_1453 );
and ( \756_b1 , \756_b0 , w_1454 );
and ( w_1459 , w_1463 , \277_b1 );
or ( w_1446 , w_1447 , w_1455 );
or ( w_1455 , w_1449 , \277_b0 );
or ( w_1450 , w_1451 , w_1456 );
or ( w_1456 , w_1452 , w_1457 );
or ( w_1457 , w_1453 , w_1458 );
or ( w_1458 , w_1454 , w_1459 );
not ( \755_SUM[21]_b1 , w_1460 );
not ( \755_SUM[21]_b0 , w_1461 );
not ( \756_b1 , w_1462 );
not ( \277_b0 , w_1463 );
and ( \757_n5[22]_b1 , 1'b0_b1 , w_1464 );
xor ( w_1464 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1465 );
and ( \757_n5[22]_b0 , w_1465 , 1'b1_b0 );
or ( \758_b1 , \b[22]_b1 , w_1466 );
or ( \758_b0 , \b[22]_b0 , \757_n5[22]_b0 );
not ( \757_n5[22]_b0 , w_1467 );
and ( w_1467 , w_1466 , \757_n5[22]_b1 );
buf ( \759_A[22]_b1 , \c[22]_b1 );
buf ( \759_A[22]_b0 , \c[22]_b0 );
buf ( \760_B[22]_b1 , \d[22]_b1 );
buf ( \760_B[22]_b0 , \d[22]_b0 );
buf ( \761_b1 , \760_B[22]_b1 );
not ( \761_b1 , w_1468 );
not ( \761_b0 , w_1469 );
and ( w_1468 , w_1469 , \760_B[22]_b0 );
or ( \762_b1 , \759_A[22]_b1 , \761_b1 );
xor ( \762_b0 , \759_A[22]_b0 , w_1470 );
not ( w_1470 , w_1471 );
and ( w_1471 , \761_b1 , \761_b0 );
or ( \763_b1 , \736_A[21]_b1 , \738_b1 );
not ( \738_b1 , w_1472 );
and ( \763_b0 , \736_A[21]_b0 , w_1473 );
and ( w_1472 , w_1473 , \738_b0 );
or ( \764_b1 , \738_b1 , \743_b1 );
not ( \743_b1 , w_1474 );
and ( \764_b0 , \738_b0 , w_1475 );
and ( w_1474 , w_1475 , \743_b0 );
or ( \765_b1 , \736_A[21]_b1 , \743_b1 );
not ( \743_b1 , w_1476 );
and ( \765_b0 , \736_A[21]_b0 , w_1477 );
and ( w_1476 , w_1477 , \743_b0 );
or ( \767_b1 , \762_b1 , \766_b1 );
xor ( \767_b0 , \762_b0 , w_1478 );
not ( w_1478 , w_1479 );
and ( w_1479 , \766_b1 , \766_b0 );
buf ( \768_SUM[22]_b1 , \767_b1 );
buf ( \768_SUM[22]_b0 , \767_b0 );
and ( \769_b0 , \768_SUM[22]_b0 , w_1480 );
and ( \769_b0 , \758_b0 , w_1481 );
and ( w_1494 , w_1495 , w_1482 );
and ( w_1482 , \758_b0 , w_1483 );
and ( w_1495 , \758_b1 , w_1484 );
and ( \769_b1 , \768_SUM[22]_b0 , w_1485 );
and ( \768_SUM[22]_b1 , w_1496 , w_1486 );
and ( w_1495 , \758_b0 , w_1487 );
and ( \769_b1 , \769_b0 , w_1488 );
and ( w_1493 , w_1497 , \241_b1 );
or ( w_1480 , w_1481 , w_1489 );
or ( w_1489 , w_1483 , \241_b0 );
or ( w_1484 , w_1485 , w_1490 );
or ( w_1490 , w_1486 , w_1491 );
or ( w_1491 , w_1487 , w_1492 );
or ( w_1492 , w_1488 , w_1493 );
not ( \768_SUM[22]_b1 , w_1494 );
not ( \768_SUM[22]_b0 , w_1495 );
not ( \769_b1 , w_1496 );
not ( \241_b0 , w_1497 );
buf ( \770_A[22]_b1 , \c[22]_b1 );
buf ( \770_A[22]_b0 , \c[22]_b0 );
buf ( \771_B[22]_b1 , \d[22]_b1 );
buf ( \771_B[22]_b0 , \d[22]_b0 );
or ( \772_b1 , \770_A[22]_b1 , \771_B[22]_b1 );
xor ( \772_b0 , \770_A[22]_b0 , w_1498 );
not ( w_1498 , w_1499 );
and ( w_1499 , \771_B[22]_b1 , \771_B[22]_b0 );
or ( \773_b1 , \747_A[21]_b1 , \748_B[21]_b1 );
not ( \748_B[21]_b1 , w_1500 );
and ( \773_b0 , \747_A[21]_b0 , w_1501 );
and ( w_1500 , w_1501 , \748_B[21]_b0 );
or ( \774_b1 , \748_B[21]_b1 , \753_b1 );
not ( \753_b1 , w_1502 );
and ( \774_b0 , \748_B[21]_b0 , w_1503 );
and ( w_1502 , w_1503 , \753_b0 );
or ( \775_b1 , \747_A[21]_b1 , \753_b1 );
not ( \753_b1 , w_1504 );
and ( \775_b0 , \747_A[21]_b0 , w_1505 );
and ( w_1504 , w_1505 , \753_b0 );
or ( \777_b1 , \772_b1 , \776_b1 );
xor ( \777_b0 , \772_b0 , w_1506 );
not ( w_1506 , w_1507 );
and ( w_1507 , \776_b1 , \776_b0 );
buf ( \778_SUM[22]_b1 , \777_b1 );
buf ( \778_SUM[22]_b0 , \777_b0 );
and ( \779_b0 , \778_SUM[22]_b0 , w_1508 );
and ( \779_b0 , \769_b0 , w_1509 );
and ( w_1522 , w_1523 , w_1510 );
and ( w_1510 , \769_b0 , w_1511 );
and ( w_1523 , \769_b1 , w_1512 );
and ( \779_b1 , \778_SUM[22]_b0 , w_1513 );
and ( \778_SUM[22]_b1 , w_1524 , w_1514 );
and ( w_1523 , \769_b0 , w_1515 );
and ( \779_b1 , \779_b0 , w_1516 );
and ( w_1521 , w_1525 , \277_b1 );
or ( w_1508 , w_1509 , w_1517 );
or ( w_1517 , w_1511 , \277_b0 );
or ( w_1512 , w_1513 , w_1518 );
or ( w_1518 , w_1514 , w_1519 );
or ( w_1519 , w_1515 , w_1520 );
or ( w_1520 , w_1516 , w_1521 );
not ( \778_SUM[22]_b1 , w_1522 );
not ( \778_SUM[22]_b0 , w_1523 );
not ( \779_b1 , w_1524 );
not ( \277_b0 , w_1525 );
and ( \780_n5[23]_b1 , 1'b0_b1 , w_1526 );
xor ( w_1526 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1527 );
and ( \780_n5[23]_b0 , w_1527 , 1'b1_b0 );
or ( \781_b1 , \b[23]_b1 , w_1528 );
or ( \781_b0 , \b[23]_b0 , \780_n5[23]_b0 );
not ( \780_n5[23]_b0 , w_1529 );
and ( w_1529 , w_1528 , \780_n5[23]_b1 );
buf ( \782_A[23]_b1 , \c[23]_b1 );
buf ( \782_A[23]_b0 , \c[23]_b0 );
buf ( \783_B[23]_b1 , \d[23]_b1 );
buf ( \783_B[23]_b0 , \d[23]_b0 );
buf ( \784_b1 , \783_B[23]_b1 );
not ( \784_b1 , w_1530 );
not ( \784_b0 , w_1531 );
and ( w_1530 , w_1531 , \783_B[23]_b0 );
or ( \785_b1 , \782_A[23]_b1 , \784_b1 );
xor ( \785_b0 , \782_A[23]_b0 , w_1532 );
not ( w_1532 , w_1533 );
and ( w_1533 , \784_b1 , \784_b0 );
or ( \786_b1 , \759_A[22]_b1 , \761_b1 );
not ( \761_b1 , w_1534 );
and ( \786_b0 , \759_A[22]_b0 , w_1535 );
and ( w_1534 , w_1535 , \761_b0 );
or ( \787_b1 , \761_b1 , \766_b1 );
not ( \766_b1 , w_1536 );
and ( \787_b0 , \761_b0 , w_1537 );
and ( w_1536 , w_1537 , \766_b0 );
or ( \788_b1 , \759_A[22]_b1 , \766_b1 );
not ( \766_b1 , w_1538 );
and ( \788_b0 , \759_A[22]_b0 , w_1539 );
and ( w_1538 , w_1539 , \766_b0 );
or ( \790_b1 , \785_b1 , \789_b1 );
xor ( \790_b0 , \785_b0 , w_1540 );
not ( w_1540 , w_1541 );
and ( w_1541 , \789_b1 , \789_b0 );
buf ( \791_SUM[23]_b1 , \790_b1 );
buf ( \791_SUM[23]_b0 , \790_b0 );
and ( \792_b0 , \791_SUM[23]_b0 , w_1542 );
and ( \792_b0 , \781_b0 , w_1543 );
and ( w_1556 , w_1557 , w_1544 );
and ( w_1544 , \781_b0 , w_1545 );
and ( w_1557 , \781_b1 , w_1546 );
and ( \792_b1 , \791_SUM[23]_b0 , w_1547 );
and ( \791_SUM[23]_b1 , w_1558 , w_1548 );
and ( w_1557 , \781_b0 , w_1549 );
and ( \792_b1 , \792_b0 , w_1550 );
and ( w_1555 , w_1559 , \241_b1 );
or ( w_1542 , w_1543 , w_1551 );
or ( w_1551 , w_1545 , \241_b0 );
or ( w_1546 , w_1547 , w_1552 );
or ( w_1552 , w_1548 , w_1553 );
or ( w_1553 , w_1549 , w_1554 );
or ( w_1554 , w_1550 , w_1555 );
not ( \791_SUM[23]_b1 , w_1556 );
not ( \791_SUM[23]_b0 , w_1557 );
not ( \792_b1 , w_1558 );
not ( \241_b0 , w_1559 );
buf ( \793_A[23]_b1 , \c[23]_b1 );
buf ( \793_A[23]_b0 , \c[23]_b0 );
buf ( \794_B[23]_b1 , \d[23]_b1 );
buf ( \794_B[23]_b0 , \d[23]_b0 );
or ( \795_b1 , \793_A[23]_b1 , \794_B[23]_b1 );
xor ( \795_b0 , \793_A[23]_b0 , w_1560 );
not ( w_1560 , w_1561 );
and ( w_1561 , \794_B[23]_b1 , \794_B[23]_b0 );
or ( \796_b1 , \770_A[22]_b1 , \771_B[22]_b1 );
not ( \771_B[22]_b1 , w_1562 );
and ( \796_b0 , \770_A[22]_b0 , w_1563 );
and ( w_1562 , w_1563 , \771_B[22]_b0 );
or ( \797_b1 , \771_B[22]_b1 , \776_b1 );
not ( \776_b1 , w_1564 );
and ( \797_b0 , \771_B[22]_b0 , w_1565 );
and ( w_1564 , w_1565 , \776_b0 );
or ( \798_b1 , \770_A[22]_b1 , \776_b1 );
not ( \776_b1 , w_1566 );
and ( \798_b0 , \770_A[22]_b0 , w_1567 );
and ( w_1566 , w_1567 , \776_b0 );
or ( \800_b1 , \795_b1 , \799_b1 );
xor ( \800_b0 , \795_b0 , w_1568 );
not ( w_1568 , w_1569 );
and ( w_1569 , \799_b1 , \799_b0 );
buf ( \801_SUM[23]_b1 , \800_b1 );
buf ( \801_SUM[23]_b0 , \800_b0 );
and ( \802_b0 , \801_SUM[23]_b0 , w_1570 );
and ( \802_b0 , \792_b0 , w_1571 );
and ( w_1584 , w_1585 , w_1572 );
and ( w_1572 , \792_b0 , w_1573 );
and ( w_1585 , \792_b1 , w_1574 );
and ( \802_b1 , \801_SUM[23]_b0 , w_1575 );
and ( \801_SUM[23]_b1 , w_1586 , w_1576 );
and ( w_1585 , \792_b0 , w_1577 );
and ( \802_b1 , \802_b0 , w_1578 );
and ( w_1583 , w_1587 , \277_b1 );
or ( w_1570 , w_1571 , w_1579 );
or ( w_1579 , w_1573 , \277_b0 );
or ( w_1574 , w_1575 , w_1580 );
or ( w_1580 , w_1576 , w_1581 );
or ( w_1581 , w_1577 , w_1582 );
or ( w_1582 , w_1578 , w_1583 );
not ( \801_SUM[23]_b1 , w_1584 );
not ( \801_SUM[23]_b0 , w_1585 );
not ( \802_b1 , w_1586 );
not ( \277_b0 , w_1587 );
and ( \803_n5[24]_b1 , 1'b0_b1 , w_1588 );
xor ( w_1588 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1589 );
and ( \803_n5[24]_b0 , w_1589 , 1'b1_b0 );
or ( \804_b1 , \b[24]_b1 , w_1590 );
or ( \804_b0 , \b[24]_b0 , \803_n5[24]_b0 );
not ( \803_n5[24]_b0 , w_1591 );
and ( w_1591 , w_1590 , \803_n5[24]_b1 );
buf ( \805_A[24]_b1 , \c[24]_b1 );
buf ( \805_A[24]_b0 , \c[24]_b0 );
buf ( \806_B[24]_b1 , \d[24]_b1 );
buf ( \806_B[24]_b0 , \d[24]_b0 );
buf ( \807_b1 , \806_B[24]_b1 );
not ( \807_b1 , w_1592 );
not ( \807_b0 , w_1593 );
and ( w_1592 , w_1593 , \806_B[24]_b0 );
or ( \808_b1 , \805_A[24]_b1 , \807_b1 );
xor ( \808_b0 , \805_A[24]_b0 , w_1594 );
not ( w_1594 , w_1595 );
and ( w_1595 , \807_b1 , \807_b0 );
or ( \809_b1 , \782_A[23]_b1 , \784_b1 );
not ( \784_b1 , w_1596 );
and ( \809_b0 , \782_A[23]_b0 , w_1597 );
and ( w_1596 , w_1597 , \784_b0 );
or ( \810_b1 , \784_b1 , \789_b1 );
not ( \789_b1 , w_1598 );
and ( \810_b0 , \784_b0 , w_1599 );
and ( w_1598 , w_1599 , \789_b0 );
or ( \811_b1 , \782_A[23]_b1 , \789_b1 );
not ( \789_b1 , w_1600 );
and ( \811_b0 , \782_A[23]_b0 , w_1601 );
and ( w_1600 , w_1601 , \789_b0 );
or ( \813_b1 , \808_b1 , \812_b1 );
xor ( \813_b0 , \808_b0 , w_1602 );
not ( w_1602 , w_1603 );
and ( w_1603 , \812_b1 , \812_b0 );
buf ( \814_SUM[24]_b1 , \813_b1 );
buf ( \814_SUM[24]_b0 , \813_b0 );
and ( \815_b0 , \814_SUM[24]_b0 , w_1604 );
and ( \815_b0 , \804_b0 , w_1605 );
and ( w_1618 , w_1619 , w_1606 );
and ( w_1606 , \804_b0 , w_1607 );
and ( w_1619 , \804_b1 , w_1608 );
and ( \815_b1 , \814_SUM[24]_b0 , w_1609 );
and ( \814_SUM[24]_b1 , w_1620 , w_1610 );
and ( w_1619 , \804_b0 , w_1611 );
and ( \815_b1 , \815_b0 , w_1612 );
and ( w_1617 , w_1621 , \241_b1 );
or ( w_1604 , w_1605 , w_1613 );
or ( w_1613 , w_1607 , \241_b0 );
or ( w_1608 , w_1609 , w_1614 );
or ( w_1614 , w_1610 , w_1615 );
or ( w_1615 , w_1611 , w_1616 );
or ( w_1616 , w_1612 , w_1617 );
not ( \814_SUM[24]_b1 , w_1618 );
not ( \814_SUM[24]_b0 , w_1619 );
not ( \815_b1 , w_1620 );
not ( \241_b0 , w_1621 );
buf ( \816_A[24]_b1 , \c[24]_b1 );
buf ( \816_A[24]_b0 , \c[24]_b0 );
buf ( \817_B[24]_b1 , \d[24]_b1 );
buf ( \817_B[24]_b0 , \d[24]_b0 );
or ( \818_b1 , \816_A[24]_b1 , \817_B[24]_b1 );
xor ( \818_b0 , \816_A[24]_b0 , w_1622 );
not ( w_1622 , w_1623 );
and ( w_1623 , \817_B[24]_b1 , \817_B[24]_b0 );
or ( \819_b1 , \793_A[23]_b1 , \794_B[23]_b1 );
not ( \794_B[23]_b1 , w_1624 );
and ( \819_b0 , \793_A[23]_b0 , w_1625 );
and ( w_1624 , w_1625 , \794_B[23]_b0 );
or ( \820_b1 , \794_B[23]_b1 , \799_b1 );
not ( \799_b1 , w_1626 );
and ( \820_b0 , \794_B[23]_b0 , w_1627 );
and ( w_1626 , w_1627 , \799_b0 );
or ( \821_b1 , \793_A[23]_b1 , \799_b1 );
not ( \799_b1 , w_1628 );
and ( \821_b0 , \793_A[23]_b0 , w_1629 );
and ( w_1628 , w_1629 , \799_b0 );
or ( \823_b1 , \818_b1 , \822_b1 );
xor ( \823_b0 , \818_b0 , w_1630 );
not ( w_1630 , w_1631 );
and ( w_1631 , \822_b1 , \822_b0 );
buf ( \824_SUM[24]_b1 , \823_b1 );
buf ( \824_SUM[24]_b0 , \823_b0 );
and ( \825_b0 , \824_SUM[24]_b0 , w_1632 );
and ( \825_b0 , \815_b0 , w_1633 );
and ( w_1646 , w_1647 , w_1634 );
and ( w_1634 , \815_b0 , w_1635 );
and ( w_1647 , \815_b1 , w_1636 );
and ( \825_b1 , \824_SUM[24]_b0 , w_1637 );
and ( \824_SUM[24]_b1 , w_1648 , w_1638 );
and ( w_1647 , \815_b0 , w_1639 );
and ( \825_b1 , \825_b0 , w_1640 );
and ( w_1645 , w_1649 , \277_b1 );
or ( w_1632 , w_1633 , w_1641 );
or ( w_1641 , w_1635 , \277_b0 );
or ( w_1636 , w_1637 , w_1642 );
or ( w_1642 , w_1638 , w_1643 );
or ( w_1643 , w_1639 , w_1644 );
or ( w_1644 , w_1640 , w_1645 );
not ( \824_SUM[24]_b1 , w_1646 );
not ( \824_SUM[24]_b0 , w_1647 );
not ( \825_b1 , w_1648 );
not ( \277_b0 , w_1649 );
and ( \826_n5[25]_b1 , 1'b0_b1 , w_1650 );
xor ( w_1650 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1651 );
and ( \826_n5[25]_b0 , w_1651 , 1'b1_b0 );
or ( \827_b1 , \b[25]_b1 , w_1652 );
or ( \827_b0 , \b[25]_b0 , \826_n5[25]_b0 );
not ( \826_n5[25]_b0 , w_1653 );
and ( w_1653 , w_1652 , \826_n5[25]_b1 );
buf ( \828_A[25]_b1 , \c[25]_b1 );
buf ( \828_A[25]_b0 , \c[25]_b0 );
buf ( \829_B[25]_b1 , \d[25]_b1 );
buf ( \829_B[25]_b0 , \d[25]_b0 );
buf ( \830_b1 , \829_B[25]_b1 );
not ( \830_b1 , w_1654 );
not ( \830_b0 , w_1655 );
and ( w_1654 , w_1655 , \829_B[25]_b0 );
or ( \831_b1 , \828_A[25]_b1 , \830_b1 );
xor ( \831_b0 , \828_A[25]_b0 , w_1656 );
not ( w_1656 , w_1657 );
and ( w_1657 , \830_b1 , \830_b0 );
or ( \832_b1 , \805_A[24]_b1 , \807_b1 );
not ( \807_b1 , w_1658 );
and ( \832_b0 , \805_A[24]_b0 , w_1659 );
and ( w_1658 , w_1659 , \807_b0 );
or ( \833_b1 , \807_b1 , \812_b1 );
not ( \812_b1 , w_1660 );
and ( \833_b0 , \807_b0 , w_1661 );
and ( w_1660 , w_1661 , \812_b0 );
or ( \834_b1 , \805_A[24]_b1 , \812_b1 );
not ( \812_b1 , w_1662 );
and ( \834_b0 , \805_A[24]_b0 , w_1663 );
and ( w_1662 , w_1663 , \812_b0 );
or ( \836_b1 , \831_b1 , \835_b1 );
xor ( \836_b0 , \831_b0 , w_1664 );
not ( w_1664 , w_1665 );
and ( w_1665 , \835_b1 , \835_b0 );
buf ( \837_SUM[25]_b1 , \836_b1 );
buf ( \837_SUM[25]_b0 , \836_b0 );
and ( \838_b0 , \837_SUM[25]_b0 , w_1666 );
and ( \838_b0 , \827_b0 , w_1667 );
and ( w_1680 , w_1681 , w_1668 );
and ( w_1668 , \827_b0 , w_1669 );
and ( w_1681 , \827_b1 , w_1670 );
and ( \838_b1 , \837_SUM[25]_b0 , w_1671 );
and ( \837_SUM[25]_b1 , w_1682 , w_1672 );
and ( w_1681 , \827_b0 , w_1673 );
and ( \838_b1 , \838_b0 , w_1674 );
and ( w_1679 , w_1683 , \241_b1 );
or ( w_1666 , w_1667 , w_1675 );
or ( w_1675 , w_1669 , \241_b0 );
or ( w_1670 , w_1671 , w_1676 );
or ( w_1676 , w_1672 , w_1677 );
or ( w_1677 , w_1673 , w_1678 );
or ( w_1678 , w_1674 , w_1679 );
not ( \837_SUM[25]_b1 , w_1680 );
not ( \837_SUM[25]_b0 , w_1681 );
not ( \838_b1 , w_1682 );
not ( \241_b0 , w_1683 );
buf ( \839_A[25]_b1 , \c[25]_b1 );
buf ( \839_A[25]_b0 , \c[25]_b0 );
buf ( \840_B[25]_b1 , \d[25]_b1 );
buf ( \840_B[25]_b0 , \d[25]_b0 );
or ( \841_b1 , \839_A[25]_b1 , \840_B[25]_b1 );
xor ( \841_b0 , \839_A[25]_b0 , w_1684 );
not ( w_1684 , w_1685 );
and ( w_1685 , \840_B[25]_b1 , \840_B[25]_b0 );
or ( \842_b1 , \816_A[24]_b1 , \817_B[24]_b1 );
not ( \817_B[24]_b1 , w_1686 );
and ( \842_b0 , \816_A[24]_b0 , w_1687 );
and ( w_1686 , w_1687 , \817_B[24]_b0 );
or ( \843_b1 , \817_B[24]_b1 , \822_b1 );
not ( \822_b1 , w_1688 );
and ( \843_b0 , \817_B[24]_b0 , w_1689 );
and ( w_1688 , w_1689 , \822_b0 );
or ( \844_b1 , \816_A[24]_b1 , \822_b1 );
not ( \822_b1 , w_1690 );
and ( \844_b0 , \816_A[24]_b0 , w_1691 );
and ( w_1690 , w_1691 , \822_b0 );
or ( \846_b1 , \841_b1 , \845_b1 );
xor ( \846_b0 , \841_b0 , w_1692 );
not ( w_1692 , w_1693 );
and ( w_1693 , \845_b1 , \845_b0 );
buf ( \847_SUM[25]_b1 , \846_b1 );
buf ( \847_SUM[25]_b0 , \846_b0 );
and ( \848_b0 , \847_SUM[25]_b0 , w_1694 );
and ( \848_b0 , \838_b0 , w_1695 );
and ( w_1708 , w_1709 , w_1696 );
and ( w_1696 , \838_b0 , w_1697 );
and ( w_1709 , \838_b1 , w_1698 );
and ( \848_b1 , \847_SUM[25]_b0 , w_1699 );
and ( \847_SUM[25]_b1 , w_1710 , w_1700 );
and ( w_1709 , \838_b0 , w_1701 );
and ( \848_b1 , \848_b0 , w_1702 );
and ( w_1707 , w_1711 , \277_b1 );
or ( w_1694 , w_1695 , w_1703 );
or ( w_1703 , w_1697 , \277_b0 );
or ( w_1698 , w_1699 , w_1704 );
or ( w_1704 , w_1700 , w_1705 );
or ( w_1705 , w_1701 , w_1706 );
or ( w_1706 , w_1702 , w_1707 );
not ( \847_SUM[25]_b1 , w_1708 );
not ( \847_SUM[25]_b0 , w_1709 );
not ( \848_b1 , w_1710 );
not ( \277_b0 , w_1711 );
and ( \849_n5[26]_b1 , 1'b0_b1 , w_1712 );
xor ( w_1712 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1713 );
and ( \849_n5[26]_b0 , w_1713 , 1'b1_b0 );
or ( \850_b1 , \b[26]_b1 , w_1714 );
or ( \850_b0 , \b[26]_b0 , \849_n5[26]_b0 );
not ( \849_n5[26]_b0 , w_1715 );
and ( w_1715 , w_1714 , \849_n5[26]_b1 );
buf ( \851_A[26]_b1 , \c[26]_b1 );
buf ( \851_A[26]_b0 , \c[26]_b0 );
buf ( \852_B[26]_b1 , \d[26]_b1 );
buf ( \852_B[26]_b0 , \d[26]_b0 );
buf ( \853_b1 , \852_B[26]_b1 );
not ( \853_b1 , w_1716 );
not ( \853_b0 , w_1717 );
and ( w_1716 , w_1717 , \852_B[26]_b0 );
or ( \854_b1 , \851_A[26]_b1 , \853_b1 );
xor ( \854_b0 , \851_A[26]_b0 , w_1718 );
not ( w_1718 , w_1719 );
and ( w_1719 , \853_b1 , \853_b0 );
or ( \855_b1 , \828_A[25]_b1 , \830_b1 );
not ( \830_b1 , w_1720 );
and ( \855_b0 , \828_A[25]_b0 , w_1721 );
and ( w_1720 , w_1721 , \830_b0 );
or ( \856_b1 , \830_b1 , \835_b1 );
not ( \835_b1 , w_1722 );
and ( \856_b0 , \830_b0 , w_1723 );
and ( w_1722 , w_1723 , \835_b0 );
or ( \857_b1 , \828_A[25]_b1 , \835_b1 );
not ( \835_b1 , w_1724 );
and ( \857_b0 , \828_A[25]_b0 , w_1725 );
and ( w_1724 , w_1725 , \835_b0 );
or ( \859_b1 , \854_b1 , \858_b1 );
xor ( \859_b0 , \854_b0 , w_1726 );
not ( w_1726 , w_1727 );
and ( w_1727 , \858_b1 , \858_b0 );
buf ( \860_SUM[26]_b1 , \859_b1 );
buf ( \860_SUM[26]_b0 , \859_b0 );
and ( \861_b0 , \860_SUM[26]_b0 , w_1728 );
and ( \861_b0 , \850_b0 , w_1729 );
and ( w_1742 , w_1743 , w_1730 );
and ( w_1730 , \850_b0 , w_1731 );
and ( w_1743 , \850_b1 , w_1732 );
and ( \861_b1 , \860_SUM[26]_b0 , w_1733 );
and ( \860_SUM[26]_b1 , w_1744 , w_1734 );
and ( w_1743 , \850_b0 , w_1735 );
and ( \861_b1 , \861_b0 , w_1736 );
and ( w_1741 , w_1745 , \241_b1 );
or ( w_1728 , w_1729 , w_1737 );
or ( w_1737 , w_1731 , \241_b0 );
or ( w_1732 , w_1733 , w_1738 );
or ( w_1738 , w_1734 , w_1739 );
or ( w_1739 , w_1735 , w_1740 );
or ( w_1740 , w_1736 , w_1741 );
not ( \860_SUM[26]_b1 , w_1742 );
not ( \860_SUM[26]_b0 , w_1743 );
not ( \861_b1 , w_1744 );
not ( \241_b0 , w_1745 );
buf ( \862_A[26]_b1 , \c[26]_b1 );
buf ( \862_A[26]_b0 , \c[26]_b0 );
buf ( \863_B[26]_b1 , \d[26]_b1 );
buf ( \863_B[26]_b0 , \d[26]_b0 );
or ( \864_b1 , \862_A[26]_b1 , \863_B[26]_b1 );
xor ( \864_b0 , \862_A[26]_b0 , w_1746 );
not ( w_1746 , w_1747 );
and ( w_1747 , \863_B[26]_b1 , \863_B[26]_b0 );
or ( \865_b1 , \839_A[25]_b1 , \840_B[25]_b1 );
not ( \840_B[25]_b1 , w_1748 );
and ( \865_b0 , \839_A[25]_b0 , w_1749 );
and ( w_1748 , w_1749 , \840_B[25]_b0 );
or ( \866_b1 , \840_B[25]_b1 , \845_b1 );
not ( \845_b1 , w_1750 );
and ( \866_b0 , \840_B[25]_b0 , w_1751 );
and ( w_1750 , w_1751 , \845_b0 );
or ( \867_b1 , \839_A[25]_b1 , \845_b1 );
not ( \845_b1 , w_1752 );
and ( \867_b0 , \839_A[25]_b0 , w_1753 );
and ( w_1752 , w_1753 , \845_b0 );
or ( \869_b1 , \864_b1 , \868_b1 );
xor ( \869_b0 , \864_b0 , w_1754 );
not ( w_1754 , w_1755 );
and ( w_1755 , \868_b1 , \868_b0 );
buf ( \870_SUM[26]_b1 , \869_b1 );
buf ( \870_SUM[26]_b0 , \869_b0 );
and ( \871_b0 , \870_SUM[26]_b0 , w_1756 );
and ( \871_b0 , \861_b0 , w_1757 );
and ( w_1770 , w_1771 , w_1758 );
and ( w_1758 , \861_b0 , w_1759 );
and ( w_1771 , \861_b1 , w_1760 );
and ( \871_b1 , \870_SUM[26]_b0 , w_1761 );
and ( \870_SUM[26]_b1 , w_1772 , w_1762 );
and ( w_1771 , \861_b0 , w_1763 );
and ( \871_b1 , \871_b0 , w_1764 );
and ( w_1769 , w_1773 , \277_b1 );
or ( w_1756 , w_1757 , w_1765 );
or ( w_1765 , w_1759 , \277_b0 );
or ( w_1760 , w_1761 , w_1766 );
or ( w_1766 , w_1762 , w_1767 );
or ( w_1767 , w_1763 , w_1768 );
or ( w_1768 , w_1764 , w_1769 );
not ( \870_SUM[26]_b1 , w_1770 );
not ( \870_SUM[26]_b0 , w_1771 );
not ( \871_b1 , w_1772 );
not ( \277_b0 , w_1773 );
and ( \872_n5[27]_b1 , 1'b0_b1 , w_1774 );
xor ( w_1774 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1775 );
and ( \872_n5[27]_b0 , w_1775 , 1'b1_b0 );
or ( \873_b1 , \b[27]_b1 , w_1776 );
or ( \873_b0 , \b[27]_b0 , \872_n5[27]_b0 );
not ( \872_n5[27]_b0 , w_1777 );
and ( w_1777 , w_1776 , \872_n5[27]_b1 );
buf ( \874_A[27]_b1 , \c[27]_b1 );
buf ( \874_A[27]_b0 , \c[27]_b0 );
buf ( \875_B[27]_b1 , \d[27]_b1 );
buf ( \875_B[27]_b0 , \d[27]_b0 );
buf ( \876_b1 , \875_B[27]_b1 );
not ( \876_b1 , w_1778 );
not ( \876_b0 , w_1779 );
and ( w_1778 , w_1779 , \875_B[27]_b0 );
or ( \877_b1 , \874_A[27]_b1 , \876_b1 );
xor ( \877_b0 , \874_A[27]_b0 , w_1780 );
not ( w_1780 , w_1781 );
and ( w_1781 , \876_b1 , \876_b0 );
or ( \878_b1 , \851_A[26]_b1 , \853_b1 );
not ( \853_b1 , w_1782 );
and ( \878_b0 , \851_A[26]_b0 , w_1783 );
and ( w_1782 , w_1783 , \853_b0 );
or ( \879_b1 , \853_b1 , \858_b1 );
not ( \858_b1 , w_1784 );
and ( \879_b0 , \853_b0 , w_1785 );
and ( w_1784 , w_1785 , \858_b0 );
or ( \880_b1 , \851_A[26]_b1 , \858_b1 );
not ( \858_b1 , w_1786 );
and ( \880_b0 , \851_A[26]_b0 , w_1787 );
and ( w_1786 , w_1787 , \858_b0 );
or ( \882_b1 , \877_b1 , \881_b1 );
xor ( \882_b0 , \877_b0 , w_1788 );
not ( w_1788 , w_1789 );
and ( w_1789 , \881_b1 , \881_b0 );
buf ( \883_SUM[27]_b1 , \882_b1 );
buf ( \883_SUM[27]_b0 , \882_b0 );
and ( \884_b0 , \883_SUM[27]_b0 , w_1790 );
and ( \884_b0 , \873_b0 , w_1791 );
and ( w_1804 , w_1805 , w_1792 );
and ( w_1792 , \873_b0 , w_1793 );
and ( w_1805 , \873_b1 , w_1794 );
and ( \884_b1 , \883_SUM[27]_b0 , w_1795 );
and ( \883_SUM[27]_b1 , w_1806 , w_1796 );
and ( w_1805 , \873_b0 , w_1797 );
and ( \884_b1 , \884_b0 , w_1798 );
and ( w_1803 , w_1807 , \241_b1 );
or ( w_1790 , w_1791 , w_1799 );
or ( w_1799 , w_1793 , \241_b0 );
or ( w_1794 , w_1795 , w_1800 );
or ( w_1800 , w_1796 , w_1801 );
or ( w_1801 , w_1797 , w_1802 );
or ( w_1802 , w_1798 , w_1803 );
not ( \883_SUM[27]_b1 , w_1804 );
not ( \883_SUM[27]_b0 , w_1805 );
not ( \884_b1 , w_1806 );
not ( \241_b0 , w_1807 );
buf ( \885_A[27]_b1 , \c[27]_b1 );
buf ( \885_A[27]_b0 , \c[27]_b0 );
buf ( \886_B[27]_b1 , \d[27]_b1 );
buf ( \886_B[27]_b0 , \d[27]_b0 );
or ( \887_b1 , \885_A[27]_b1 , \886_B[27]_b1 );
xor ( \887_b0 , \885_A[27]_b0 , w_1808 );
not ( w_1808 , w_1809 );
and ( w_1809 , \886_B[27]_b1 , \886_B[27]_b0 );
or ( \888_b1 , \862_A[26]_b1 , \863_B[26]_b1 );
not ( \863_B[26]_b1 , w_1810 );
and ( \888_b0 , \862_A[26]_b0 , w_1811 );
and ( w_1810 , w_1811 , \863_B[26]_b0 );
or ( \889_b1 , \863_B[26]_b1 , \868_b1 );
not ( \868_b1 , w_1812 );
and ( \889_b0 , \863_B[26]_b0 , w_1813 );
and ( w_1812 , w_1813 , \868_b0 );
or ( \890_b1 , \862_A[26]_b1 , \868_b1 );
not ( \868_b1 , w_1814 );
and ( \890_b0 , \862_A[26]_b0 , w_1815 );
and ( w_1814 , w_1815 , \868_b0 );
or ( \892_b1 , \887_b1 , \891_b1 );
xor ( \892_b0 , \887_b0 , w_1816 );
not ( w_1816 , w_1817 );
and ( w_1817 , \891_b1 , \891_b0 );
buf ( \893_SUM[27]_b1 , \892_b1 );
buf ( \893_SUM[27]_b0 , \892_b0 );
and ( \894_b0 , \893_SUM[27]_b0 , w_1818 );
and ( \894_b0 , \884_b0 , w_1819 );
and ( w_1832 , w_1833 , w_1820 );
and ( w_1820 , \884_b0 , w_1821 );
and ( w_1833 , \884_b1 , w_1822 );
and ( \894_b1 , \893_SUM[27]_b0 , w_1823 );
and ( \893_SUM[27]_b1 , w_1834 , w_1824 );
and ( w_1833 , \884_b0 , w_1825 );
and ( \894_b1 , \894_b0 , w_1826 );
and ( w_1831 , w_1835 , \277_b1 );
or ( w_1818 , w_1819 , w_1827 );
or ( w_1827 , w_1821 , \277_b0 );
or ( w_1822 , w_1823 , w_1828 );
or ( w_1828 , w_1824 , w_1829 );
or ( w_1829 , w_1825 , w_1830 );
or ( w_1830 , w_1826 , w_1831 );
not ( \893_SUM[27]_b1 , w_1832 );
not ( \893_SUM[27]_b0 , w_1833 );
not ( \894_b1 , w_1834 );
not ( \277_b0 , w_1835 );
and ( \895_n5[28]_b1 , 1'b0_b1 , w_1836 );
xor ( w_1836 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1837 );
and ( \895_n5[28]_b0 , w_1837 , 1'b1_b0 );
or ( \896_b1 , \b[28]_b1 , w_1838 );
or ( \896_b0 , \b[28]_b0 , \895_n5[28]_b0 );
not ( \895_n5[28]_b0 , w_1839 );
and ( w_1839 , w_1838 , \895_n5[28]_b1 );
buf ( \897_A[28]_b1 , \c[28]_b1 );
buf ( \897_A[28]_b0 , \c[28]_b0 );
buf ( \898_B[28]_b1 , \d[28]_b1 );
buf ( \898_B[28]_b0 , \d[28]_b0 );
buf ( \899_b1 , \898_B[28]_b1 );
not ( \899_b1 , w_1840 );
not ( \899_b0 , w_1841 );
and ( w_1840 , w_1841 , \898_B[28]_b0 );
or ( \900_b1 , \897_A[28]_b1 , \899_b1 );
xor ( \900_b0 , \897_A[28]_b0 , w_1842 );
not ( w_1842 , w_1843 );
and ( w_1843 , \899_b1 , \899_b0 );
or ( \901_b1 , \874_A[27]_b1 , \876_b1 );
not ( \876_b1 , w_1844 );
and ( \901_b0 , \874_A[27]_b0 , w_1845 );
and ( w_1844 , w_1845 , \876_b0 );
or ( \902_b1 , \876_b1 , \881_b1 );
not ( \881_b1 , w_1846 );
and ( \902_b0 , \876_b0 , w_1847 );
and ( w_1846 , w_1847 , \881_b0 );
or ( \903_b1 , \874_A[27]_b1 , \881_b1 );
not ( \881_b1 , w_1848 );
and ( \903_b0 , \874_A[27]_b0 , w_1849 );
and ( w_1848 , w_1849 , \881_b0 );
or ( \905_b1 , \900_b1 , \904_b1 );
xor ( \905_b0 , \900_b0 , w_1850 );
not ( w_1850 , w_1851 );
and ( w_1851 , \904_b1 , \904_b0 );
buf ( \906_SUM[28]_b1 , \905_b1 );
buf ( \906_SUM[28]_b0 , \905_b0 );
and ( \907_b0 , \906_SUM[28]_b0 , w_1852 );
and ( \907_b0 , \896_b0 , w_1853 );
and ( w_1866 , w_1867 , w_1854 );
and ( w_1854 , \896_b0 , w_1855 );
and ( w_1867 , \896_b1 , w_1856 );
and ( \907_b1 , \906_SUM[28]_b0 , w_1857 );
and ( \906_SUM[28]_b1 , w_1868 , w_1858 );
and ( w_1867 , \896_b0 , w_1859 );
and ( \907_b1 , \907_b0 , w_1860 );
and ( w_1865 , w_1869 , \241_b1 );
or ( w_1852 , w_1853 , w_1861 );
or ( w_1861 , w_1855 , \241_b0 );
or ( w_1856 , w_1857 , w_1862 );
or ( w_1862 , w_1858 , w_1863 );
or ( w_1863 , w_1859 , w_1864 );
or ( w_1864 , w_1860 , w_1865 );
not ( \906_SUM[28]_b1 , w_1866 );
not ( \906_SUM[28]_b0 , w_1867 );
not ( \907_b1 , w_1868 );
not ( \241_b0 , w_1869 );
buf ( \908_A[28]_b1 , \c[28]_b1 );
buf ( \908_A[28]_b0 , \c[28]_b0 );
buf ( \909_B[28]_b1 , \d[28]_b1 );
buf ( \909_B[28]_b0 , \d[28]_b0 );
or ( \910_b1 , \908_A[28]_b1 , \909_B[28]_b1 );
xor ( \910_b0 , \908_A[28]_b0 , w_1870 );
not ( w_1870 , w_1871 );
and ( w_1871 , \909_B[28]_b1 , \909_B[28]_b0 );
or ( \911_b1 , \885_A[27]_b1 , \886_B[27]_b1 );
not ( \886_B[27]_b1 , w_1872 );
and ( \911_b0 , \885_A[27]_b0 , w_1873 );
and ( w_1872 , w_1873 , \886_B[27]_b0 );
or ( \912_b1 , \886_B[27]_b1 , \891_b1 );
not ( \891_b1 , w_1874 );
and ( \912_b0 , \886_B[27]_b0 , w_1875 );
and ( w_1874 , w_1875 , \891_b0 );
or ( \913_b1 , \885_A[27]_b1 , \891_b1 );
not ( \891_b1 , w_1876 );
and ( \913_b0 , \885_A[27]_b0 , w_1877 );
and ( w_1876 , w_1877 , \891_b0 );
or ( \915_b1 , \910_b1 , \914_b1 );
xor ( \915_b0 , \910_b0 , w_1878 );
not ( w_1878 , w_1879 );
and ( w_1879 , \914_b1 , \914_b0 );
buf ( \916_SUM[28]_b1 , \915_b1 );
buf ( \916_SUM[28]_b0 , \915_b0 );
and ( \917_b0 , \916_SUM[28]_b0 , w_1880 );
and ( \917_b0 , \907_b0 , w_1881 );
and ( w_1894 , w_1895 , w_1882 );
and ( w_1882 , \907_b0 , w_1883 );
and ( w_1895 , \907_b1 , w_1884 );
and ( \917_b1 , \916_SUM[28]_b0 , w_1885 );
and ( \916_SUM[28]_b1 , w_1896 , w_1886 );
and ( w_1895 , \907_b0 , w_1887 );
and ( \917_b1 , \917_b0 , w_1888 );
and ( w_1893 , w_1897 , \277_b1 );
or ( w_1880 , w_1881 , w_1889 );
or ( w_1889 , w_1883 , \277_b0 );
or ( w_1884 , w_1885 , w_1890 );
or ( w_1890 , w_1886 , w_1891 );
or ( w_1891 , w_1887 , w_1892 );
or ( w_1892 , w_1888 , w_1893 );
not ( \916_SUM[28]_b1 , w_1894 );
not ( \916_SUM[28]_b0 , w_1895 );
not ( \917_b1 , w_1896 );
not ( \277_b0 , w_1897 );
and ( \918_n5[29]_b1 , 1'b0_b1 , w_1898 );
xor ( w_1898 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1899 );
and ( \918_n5[29]_b0 , w_1899 , 1'b1_b0 );
or ( \919_b1 , \b[29]_b1 , w_1900 );
or ( \919_b0 , \b[29]_b0 , \918_n5[29]_b0 );
not ( \918_n5[29]_b0 , w_1901 );
and ( w_1901 , w_1900 , \918_n5[29]_b1 );
buf ( \920_A[29]_b1 , \c[29]_b1 );
buf ( \920_A[29]_b0 , \c[29]_b0 );
buf ( \921_B[29]_b1 , \d[29]_b1 );
buf ( \921_B[29]_b0 , \d[29]_b0 );
buf ( \922_b1 , \921_B[29]_b1 );
not ( \922_b1 , w_1902 );
not ( \922_b0 , w_1903 );
and ( w_1902 , w_1903 , \921_B[29]_b0 );
or ( \923_b1 , \920_A[29]_b1 , \922_b1 );
xor ( \923_b0 , \920_A[29]_b0 , w_1904 );
not ( w_1904 , w_1905 );
and ( w_1905 , \922_b1 , \922_b0 );
or ( \924_b1 , \897_A[28]_b1 , \899_b1 );
not ( \899_b1 , w_1906 );
and ( \924_b0 , \897_A[28]_b0 , w_1907 );
and ( w_1906 , w_1907 , \899_b0 );
or ( \925_b1 , \899_b1 , \904_b1 );
not ( \904_b1 , w_1908 );
and ( \925_b0 , \899_b0 , w_1909 );
and ( w_1908 , w_1909 , \904_b0 );
or ( \926_b1 , \897_A[28]_b1 , \904_b1 );
not ( \904_b1 , w_1910 );
and ( \926_b0 , \897_A[28]_b0 , w_1911 );
and ( w_1910 , w_1911 , \904_b0 );
or ( \928_b1 , \923_b1 , \927_b1 );
xor ( \928_b0 , \923_b0 , w_1912 );
not ( w_1912 , w_1913 );
and ( w_1913 , \927_b1 , \927_b0 );
buf ( \929_SUM[29]_b1 , \928_b1 );
buf ( \929_SUM[29]_b0 , \928_b0 );
and ( \930_b0 , \929_SUM[29]_b0 , w_1914 );
and ( \930_b0 , \919_b0 , w_1915 );
and ( w_1928 , w_1929 , w_1916 );
and ( w_1916 , \919_b0 , w_1917 );
and ( w_1929 , \919_b1 , w_1918 );
and ( \930_b1 , \929_SUM[29]_b0 , w_1919 );
and ( \929_SUM[29]_b1 , w_1930 , w_1920 );
and ( w_1929 , \919_b0 , w_1921 );
and ( \930_b1 , \930_b0 , w_1922 );
and ( w_1927 , w_1931 , \241_b1 );
or ( w_1914 , w_1915 , w_1923 );
or ( w_1923 , w_1917 , \241_b0 );
or ( w_1918 , w_1919 , w_1924 );
or ( w_1924 , w_1920 , w_1925 );
or ( w_1925 , w_1921 , w_1926 );
or ( w_1926 , w_1922 , w_1927 );
not ( \929_SUM[29]_b1 , w_1928 );
not ( \929_SUM[29]_b0 , w_1929 );
not ( \930_b1 , w_1930 );
not ( \241_b0 , w_1931 );
buf ( \931_A[29]_b1 , \c[29]_b1 );
buf ( \931_A[29]_b0 , \c[29]_b0 );
buf ( \932_B[29]_b1 , \d[29]_b1 );
buf ( \932_B[29]_b0 , \d[29]_b0 );
or ( \933_b1 , \931_A[29]_b1 , \932_B[29]_b1 );
xor ( \933_b0 , \931_A[29]_b0 , w_1932 );
not ( w_1932 , w_1933 );
and ( w_1933 , \932_B[29]_b1 , \932_B[29]_b0 );
or ( \934_b1 , \908_A[28]_b1 , \909_B[28]_b1 );
not ( \909_B[28]_b1 , w_1934 );
and ( \934_b0 , \908_A[28]_b0 , w_1935 );
and ( w_1934 , w_1935 , \909_B[28]_b0 );
or ( \935_b1 , \909_B[28]_b1 , \914_b1 );
not ( \914_b1 , w_1936 );
and ( \935_b0 , \909_B[28]_b0 , w_1937 );
and ( w_1936 , w_1937 , \914_b0 );
or ( \936_b1 , \908_A[28]_b1 , \914_b1 );
not ( \914_b1 , w_1938 );
and ( \936_b0 , \908_A[28]_b0 , w_1939 );
and ( w_1938 , w_1939 , \914_b0 );
or ( \938_b1 , \933_b1 , \937_b1 );
xor ( \938_b0 , \933_b0 , w_1940 );
not ( w_1940 , w_1941 );
and ( w_1941 , \937_b1 , \937_b0 );
buf ( \939_SUM[29]_b1 , \938_b1 );
buf ( \939_SUM[29]_b0 , \938_b0 );
and ( \940_b0 , \939_SUM[29]_b0 , w_1942 );
and ( \940_b0 , \930_b0 , w_1943 );
and ( w_1956 , w_1957 , w_1944 );
and ( w_1944 , \930_b0 , w_1945 );
and ( w_1957 , \930_b1 , w_1946 );
and ( \940_b1 , \939_SUM[29]_b0 , w_1947 );
and ( \939_SUM[29]_b1 , w_1958 , w_1948 );
and ( w_1957 , \930_b0 , w_1949 );
and ( \940_b1 , \940_b0 , w_1950 );
and ( w_1955 , w_1959 , \277_b1 );
or ( w_1942 , w_1943 , w_1951 );
or ( w_1951 , w_1945 , \277_b0 );
or ( w_1946 , w_1947 , w_1952 );
or ( w_1952 , w_1948 , w_1953 );
or ( w_1953 , w_1949 , w_1954 );
or ( w_1954 , w_1950 , w_1955 );
not ( \939_SUM[29]_b1 , w_1956 );
not ( \939_SUM[29]_b0 , w_1957 );
not ( \940_b1 , w_1958 );
not ( \277_b0 , w_1959 );
and ( \941_n5[30]_b1 , 1'b0_b1 , w_1960 );
xor ( w_1960 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_1961 );
and ( \941_n5[30]_b0 , w_1961 , 1'b1_b0 );
or ( \942_b1 , \b[30]_b1 , w_1962 );
or ( \942_b0 , \b[30]_b0 , \941_n5[30]_b0 );
not ( \941_n5[30]_b0 , w_1963 );
and ( w_1963 , w_1962 , \941_n5[30]_b1 );
buf ( \943_A[30]_b1 , \c[30]_b1 );
buf ( \943_A[30]_b0 , \c[30]_b0 );
buf ( \944_B[30]_b1 , \d[30]_b1 );
buf ( \944_B[30]_b0 , \d[30]_b0 );
buf ( \945_b1 , \944_B[30]_b1 );
not ( \945_b1 , w_1964 );
not ( \945_b0 , w_1965 );
and ( w_1964 , w_1965 , \944_B[30]_b0 );
or ( \946_b1 , \943_A[30]_b1 , \945_b1 );
xor ( \946_b0 , \943_A[30]_b0 , w_1966 );
not ( w_1966 , w_1967 );
and ( w_1967 , \945_b1 , \945_b0 );
or ( \947_b1 , \920_A[29]_b1 , \922_b1 );
not ( \922_b1 , w_1968 );
and ( \947_b0 , \920_A[29]_b0 , w_1969 );
and ( w_1968 , w_1969 , \922_b0 );
or ( \948_b1 , \922_b1 , \927_b1 );
not ( \927_b1 , w_1970 );
and ( \948_b0 , \922_b0 , w_1971 );
and ( w_1970 , w_1971 , \927_b0 );
or ( \949_b1 , \920_A[29]_b1 , \927_b1 );
not ( \927_b1 , w_1972 );
and ( \949_b0 , \920_A[29]_b0 , w_1973 );
and ( w_1972 , w_1973 , \927_b0 );
or ( \951_b1 , \946_b1 , \950_b1 );
xor ( \951_b0 , \946_b0 , w_1974 );
not ( w_1974 , w_1975 );
and ( w_1975 , \950_b1 , \950_b0 );
buf ( \952_SUM[30]_b1 , \951_b1 );
buf ( \952_SUM[30]_b0 , \951_b0 );
and ( \953_b0 , \952_SUM[30]_b0 , w_1976 );
and ( \953_b0 , \942_b0 , w_1977 );
and ( w_1990 , w_1991 , w_1978 );
and ( w_1978 , \942_b0 , w_1979 );
and ( w_1991 , \942_b1 , w_1980 );
and ( \953_b1 , \952_SUM[30]_b0 , w_1981 );
and ( \952_SUM[30]_b1 , w_1992 , w_1982 );
and ( w_1991 , \942_b0 , w_1983 );
and ( \953_b1 , \953_b0 , w_1984 );
and ( w_1989 , w_1993 , \241_b1 );
or ( w_1976 , w_1977 , w_1985 );
or ( w_1985 , w_1979 , \241_b0 );
or ( w_1980 , w_1981 , w_1986 );
or ( w_1986 , w_1982 , w_1987 );
or ( w_1987 , w_1983 , w_1988 );
or ( w_1988 , w_1984 , w_1989 );
not ( \952_SUM[30]_b1 , w_1990 );
not ( \952_SUM[30]_b0 , w_1991 );
not ( \953_b1 , w_1992 );
not ( \241_b0 , w_1993 );
buf ( \954_A[30]_b1 , \c[30]_b1 );
buf ( \954_A[30]_b0 , \c[30]_b0 );
buf ( \955_B[30]_b1 , \d[30]_b1 );
buf ( \955_B[30]_b0 , \d[30]_b0 );
or ( \956_b1 , \954_A[30]_b1 , \955_B[30]_b1 );
xor ( \956_b0 , \954_A[30]_b0 , w_1994 );
not ( w_1994 , w_1995 );
and ( w_1995 , \955_B[30]_b1 , \955_B[30]_b0 );
or ( \957_b1 , \931_A[29]_b1 , \932_B[29]_b1 );
not ( \932_B[29]_b1 , w_1996 );
and ( \957_b0 , \931_A[29]_b0 , w_1997 );
and ( w_1996 , w_1997 , \932_B[29]_b0 );
or ( \958_b1 , \932_B[29]_b1 , \937_b1 );
not ( \937_b1 , w_1998 );
and ( \958_b0 , \932_B[29]_b0 , w_1999 );
and ( w_1998 , w_1999 , \937_b0 );
or ( \959_b1 , \931_A[29]_b1 , \937_b1 );
not ( \937_b1 , w_2000 );
and ( \959_b0 , \931_A[29]_b0 , w_2001 );
and ( w_2000 , w_2001 , \937_b0 );
or ( \961_b1 , \956_b1 , \960_b1 );
xor ( \961_b0 , \956_b0 , w_2002 );
not ( w_2002 , w_2003 );
and ( w_2003 , \960_b1 , \960_b0 );
buf ( \962_SUM[30]_b1 , \961_b1 );
buf ( \962_SUM[30]_b0 , \961_b0 );
and ( \963_b0 , \962_SUM[30]_b0 , w_2004 );
and ( \963_b0 , \953_b0 , w_2005 );
and ( w_2018 , w_2019 , w_2006 );
and ( w_2006 , \953_b0 , w_2007 );
and ( w_2019 , \953_b1 , w_2008 );
and ( \963_b1 , \962_SUM[30]_b0 , w_2009 );
and ( \962_SUM[30]_b1 , w_2020 , w_2010 );
and ( w_2019 , \953_b0 , w_2011 );
and ( \963_b1 , \963_b0 , w_2012 );
and ( w_2017 , w_2021 , \277_b1 );
or ( w_2004 , w_2005 , w_2013 );
or ( w_2013 , w_2007 , \277_b0 );
or ( w_2008 , w_2009 , w_2014 );
or ( w_2014 , w_2010 , w_2015 );
or ( w_2015 , w_2011 , w_2016 );
or ( w_2016 , w_2012 , w_2017 );
not ( \962_SUM[30]_b1 , w_2018 );
not ( \962_SUM[30]_b0 , w_2019 );
not ( \963_b1 , w_2020 );
not ( \277_b0 , w_2021 );
and ( \964_n5[31]_b1 , 1'b0_b1 , w_2022 );
xor ( w_2022 , 1'b0_b0 , 1'b1_b1 );
not ( 1'b1_b1 , w_2023 );
and ( \964_n5[31]_b0 , w_2023 , 1'b1_b0 );
or ( \965_b1 , \b[31]_b1 , w_2024 );
or ( \965_b0 , \b[31]_b0 , \964_n5[31]_b0 );
not ( \964_n5[31]_b0 , w_2025 );
and ( w_2025 , w_2024 , \964_n5[31]_b1 );
buf ( \966_A[31]_b1 , \c[31]_b1 );
buf ( \966_A[31]_b0 , \c[31]_b0 );
buf ( \967_B[31]_b1 , \d[31]_b1 );
buf ( \967_B[31]_b0 , \d[31]_b0 );
buf ( \968_b1 , \967_B[31]_b1 );
not ( \968_b1 , w_2026 );
not ( \968_b0 , w_2027 );
and ( w_2026 , w_2027 , \967_B[31]_b0 );
or ( \969_b1 , \966_A[31]_b1 , \968_b1 );
xor ( \969_b0 , \966_A[31]_b0 , w_2028 );
not ( w_2028 , w_2029 );
and ( w_2029 , \968_b1 , \968_b0 );
or ( \970_b1 , \943_A[30]_b1 , \945_b1 );
not ( \945_b1 , w_2030 );
and ( \970_b0 , \943_A[30]_b0 , w_2031 );
and ( w_2030 , w_2031 , \945_b0 );
or ( \971_b1 , \945_b1 , \950_b1 );
not ( \950_b1 , w_2032 );
and ( \971_b0 , \945_b0 , w_2033 );
and ( w_2032 , w_2033 , \950_b0 );
or ( \972_b1 , \943_A[30]_b1 , \950_b1 );
not ( \950_b1 , w_2034 );
and ( \972_b0 , \943_A[30]_b0 , w_2035 );
and ( w_2034 , w_2035 , \950_b0 );
or ( \974_b1 , \969_b1 , \973_b1 );
xor ( \974_b0 , \969_b0 , w_2036 );
not ( w_2036 , w_2037 );
and ( w_2037 , \973_b1 , \973_b0 );
buf ( \975_SUM[31]_b1 , \974_b1 );
buf ( \975_SUM[31]_b0 , \974_b0 );
and ( \976_b0 , \975_SUM[31]_b0 , w_2038 );
and ( \976_b0 , \965_b0 , w_2039 );
and ( w_2052 , w_2053 , w_2040 );
and ( w_2040 , \965_b0 , w_2041 );
and ( w_2053 , \965_b1 , w_2042 );
and ( \976_b1 , \975_SUM[31]_b0 , w_2043 );
and ( \975_SUM[31]_b1 , w_2054 , w_2044 );
and ( w_2053 , \965_b0 , w_2045 );
and ( \976_b1 , \976_b0 , w_2046 );
and ( w_2051 , w_2055 , \241_b1 );
or ( w_2038 , w_2039 , w_2047 );
or ( w_2047 , w_2041 , \241_b0 );
or ( w_2042 , w_2043 , w_2048 );
or ( w_2048 , w_2044 , w_2049 );
or ( w_2049 , w_2045 , w_2050 );
or ( w_2050 , w_2046 , w_2051 );
not ( \975_SUM[31]_b1 , w_2052 );
not ( \975_SUM[31]_b0 , w_2053 );
not ( \976_b1 , w_2054 );
not ( \241_b0 , w_2055 );
buf ( \977_A[31]_b1 , \c[31]_b1 );
buf ( \977_A[31]_b0 , \c[31]_b0 );
buf ( \978_B[31]_b1 , \d[31]_b1 );
buf ( \978_B[31]_b0 , \d[31]_b0 );
or ( \979_b1 , \977_A[31]_b1 , \978_B[31]_b1 );
xor ( \979_b0 , \977_A[31]_b0 , w_2056 );
not ( w_2056 , w_2057 );
and ( w_2057 , \978_B[31]_b1 , \978_B[31]_b0 );
or ( \980_b1 , \954_A[30]_b1 , \955_B[30]_b1 );
not ( \955_B[30]_b1 , w_2058 );
and ( \980_b0 , \954_A[30]_b0 , w_2059 );
and ( w_2058 , w_2059 , \955_B[30]_b0 );
or ( \981_b1 , \955_B[30]_b1 , \960_b1 );
not ( \960_b1 , w_2060 );
and ( \981_b0 , \955_B[30]_b0 , w_2061 );
and ( w_2060 , w_2061 , \960_b0 );
or ( \982_b1 , \954_A[30]_b1 , \960_b1 );
not ( \960_b1 , w_2062 );
and ( \982_b0 , \954_A[30]_b0 , w_2063 );
and ( w_2062 , w_2063 , \960_b0 );
or ( \984_b1 , \979_b1 , \983_b1 );
xor ( \984_b0 , \979_b0 , w_2064 );
not ( w_2064 , w_2065 );
and ( w_2065 , \983_b1 , \983_b0 );
buf ( \985_SUM[31]_b1 , \984_b1 );
buf ( \985_SUM[31]_b0 , \984_b0 );
and ( \986_b0 , \985_SUM[31]_b0 , w_2066 );
and ( \986_b0 , \976_b0 , w_2067 );
and ( w_2080 , w_2081 , w_2068 );
and ( w_2068 , \976_b0 , w_2069 );
and ( w_2081 , \976_b1 , w_2070 );
and ( \986_b1 , \985_SUM[31]_b0 , w_2071 );
and ( \985_SUM[31]_b1 , w_2082 , w_2072 );
and ( w_2081 , \976_b0 , w_2073 );
and ( \986_b1 , \986_b0 , w_2074 );
and ( w_2079 , w_2083 , \277_b1 );
or ( w_2066 , w_2067 , w_2075 );
or ( w_2075 , w_2069 , \277_b0 );
or ( w_2070 , w_2071 , w_2076 );
or ( w_2076 , w_2072 , w_2077 );
or ( w_2077 , w_2073 , w_2078 );
or ( w_2078 , w_2074 , w_2079 );
not ( \985_SUM[31]_b1 , w_2080 );
not ( \985_SUM[31]_b0 , w_2081 );
not ( \986_b1 , w_2082 );
not ( \277_b0 , w_2083 );
buf ( \987_A[31]_b1 , \a[31]_b1 );
buf ( \987_A[31]_b0 , \a[31]_b0 );
buf ( \988_B[31]_b1 , \b[31]_b1 );
buf ( \988_B[31]_b0 , \b[31]_b0 );
or ( \989_b1 , \987_A[31]_b1 , \988_B[31]_b1 );
xor ( \989_b0 , \987_A[31]_b0 , w_2084 );
not ( w_2084 , w_2085 );
and ( w_2085 , \988_B[31]_b1 , \988_B[31]_b0 );
buf ( \990_A[30]_b1 , \a[30]_b1 );
buf ( \990_A[30]_b0 , \a[30]_b0 );
buf ( \991_B[30]_b1 , \b[30]_b1 );
buf ( \991_B[30]_b0 , \b[30]_b0 );
or ( \992_b1 , \990_A[30]_b1 , \991_B[30]_b1 );
not ( \991_B[30]_b1 , w_2086 );
and ( \992_b0 , \990_A[30]_b0 , w_2087 );
and ( w_2086 , w_2087 , \991_B[30]_b0 );
buf ( \993_A[29]_b1 , \a[29]_b1 );
buf ( \993_A[29]_b0 , \a[29]_b0 );
buf ( \994_B[29]_b1 , \b[29]_b1 );
buf ( \994_B[29]_b0 , \b[29]_b0 );
or ( \995_b1 , \993_A[29]_b1 , \994_B[29]_b1 );
not ( \994_B[29]_b1 , w_2088 );
and ( \995_b0 , \993_A[29]_b0 , w_2089 );
and ( w_2088 , w_2089 , \994_B[29]_b0 );
buf ( \996_A[28]_b1 , \a[28]_b1 );
buf ( \996_A[28]_b0 , \a[28]_b0 );
buf ( \997_B[28]_b1 , \b[28]_b1 );
buf ( \997_B[28]_b0 , \b[28]_b0 );
or ( \998_b1 , \996_A[28]_b1 , \997_B[28]_b1 );
not ( \997_B[28]_b1 , w_2090 );
and ( \998_b0 , \996_A[28]_b0 , w_2091 );
and ( w_2090 , w_2091 , \997_B[28]_b0 );
buf ( \999_A[27]_b1 , \a[27]_b1 );
buf ( \999_A[27]_b0 , \a[27]_b0 );
buf ( \1000_B[27]_b1 , \b[27]_b1 );
buf ( \1000_B[27]_b0 , \b[27]_b0 );
or ( \1001_b1 , \999_A[27]_b1 , \1000_B[27]_b1 );
not ( \1000_B[27]_b1 , w_2092 );
and ( \1001_b0 , \999_A[27]_b0 , w_2093 );
and ( w_2092 , w_2093 , \1000_B[27]_b0 );
buf ( \1002_A[26]_b1 , \a[26]_b1 );
buf ( \1002_A[26]_b0 , \a[26]_b0 );
buf ( \1003_B[26]_b1 , \b[26]_b1 );
buf ( \1003_B[26]_b0 , \b[26]_b0 );
or ( \1004_b1 , \1002_A[26]_b1 , \1003_B[26]_b1 );
not ( \1003_B[26]_b1 , w_2094 );
and ( \1004_b0 , \1002_A[26]_b0 , w_2095 );
and ( w_2094 , w_2095 , \1003_B[26]_b0 );
buf ( \1005_A[25]_b1 , \a[25]_b1 );
buf ( \1005_A[25]_b0 , \a[25]_b0 );
buf ( \1006_B[25]_b1 , \b[25]_b1 );
buf ( \1006_B[25]_b0 , \b[25]_b0 );
or ( \1007_b1 , \1005_A[25]_b1 , \1006_B[25]_b1 );
not ( \1006_B[25]_b1 , w_2096 );
and ( \1007_b0 , \1005_A[25]_b0 , w_2097 );
and ( w_2096 , w_2097 , \1006_B[25]_b0 );
buf ( \1008_A[24]_b1 , \a[24]_b1 );
buf ( \1008_A[24]_b0 , \a[24]_b0 );
buf ( \1009_B[24]_b1 , \b[24]_b1 );
buf ( \1009_B[24]_b0 , \b[24]_b0 );
or ( \1010_b1 , \1008_A[24]_b1 , \1009_B[24]_b1 );
not ( \1009_B[24]_b1 , w_2098 );
and ( \1010_b0 , \1008_A[24]_b0 , w_2099 );
and ( w_2098 , w_2099 , \1009_B[24]_b0 );
buf ( \1011_A[23]_b1 , \a[23]_b1 );
buf ( \1011_A[23]_b0 , \a[23]_b0 );
buf ( \1012_B[23]_b1 , \b[23]_b1 );
buf ( \1012_B[23]_b0 , \b[23]_b0 );
or ( \1013_b1 , \1011_A[23]_b1 , \1012_B[23]_b1 );
not ( \1012_B[23]_b1 , w_2100 );
and ( \1013_b0 , \1011_A[23]_b0 , w_2101 );
and ( w_2100 , w_2101 , \1012_B[23]_b0 );
buf ( \1014_A[22]_b1 , \a[22]_b1 );
buf ( \1014_A[22]_b0 , \a[22]_b0 );
buf ( \1015_B[22]_b1 , \b[22]_b1 );
buf ( \1015_B[22]_b0 , \b[22]_b0 );
or ( \1016_b1 , \1014_A[22]_b1 , \1015_B[22]_b1 );
not ( \1015_B[22]_b1 , w_2102 );
and ( \1016_b0 , \1014_A[22]_b0 , w_2103 );
and ( w_2102 , w_2103 , \1015_B[22]_b0 );
buf ( \1017_A[21]_b1 , \a[21]_b1 );
buf ( \1017_A[21]_b0 , \a[21]_b0 );
buf ( \1018_B[21]_b1 , \b[21]_b1 );
buf ( \1018_B[21]_b0 , \b[21]_b0 );
or ( \1019_b1 , \1017_A[21]_b1 , \1018_B[21]_b1 );
not ( \1018_B[21]_b1 , w_2104 );
and ( \1019_b0 , \1017_A[21]_b0 , w_2105 );
and ( w_2104 , w_2105 , \1018_B[21]_b0 );
buf ( \1020_A[20]_b1 , \a[20]_b1 );
buf ( \1020_A[20]_b0 , \a[20]_b0 );
buf ( \1021_B[20]_b1 , \b[20]_b1 );
buf ( \1021_B[20]_b0 , \b[20]_b0 );
or ( \1022_b1 , \1020_A[20]_b1 , \1021_B[20]_b1 );
not ( \1021_B[20]_b1 , w_2106 );
and ( \1022_b0 , \1020_A[20]_b0 , w_2107 );
and ( w_2106 , w_2107 , \1021_B[20]_b0 );
buf ( \1023_A[19]_b1 , \a[19]_b1 );
buf ( \1023_A[19]_b0 , \a[19]_b0 );
buf ( \1024_B[19]_b1 , \b[19]_b1 );
buf ( \1024_B[19]_b0 , \b[19]_b0 );
or ( \1025_b1 , \1023_A[19]_b1 , \1024_B[19]_b1 );
not ( \1024_B[19]_b1 , w_2108 );
and ( \1025_b0 , \1023_A[19]_b0 , w_2109 );
and ( w_2108 , w_2109 , \1024_B[19]_b0 );
buf ( \1026_A[18]_b1 , \a[18]_b1 );
buf ( \1026_A[18]_b0 , \a[18]_b0 );
buf ( \1027_B[18]_b1 , \b[18]_b1 );
buf ( \1027_B[18]_b0 , \b[18]_b0 );
or ( \1028_b1 , \1026_A[18]_b1 , \1027_B[18]_b1 );
not ( \1027_B[18]_b1 , w_2110 );
and ( \1028_b0 , \1026_A[18]_b0 , w_2111 );
and ( w_2110 , w_2111 , \1027_B[18]_b0 );
buf ( \1029_A[17]_b1 , \a[17]_b1 );
buf ( \1029_A[17]_b0 , \a[17]_b0 );
buf ( \1030_B[17]_b1 , \b[17]_b1 );
buf ( \1030_B[17]_b0 , \b[17]_b0 );
or ( \1031_b1 , \1029_A[17]_b1 , \1030_B[17]_b1 );
not ( \1030_B[17]_b1 , w_2112 );
and ( \1031_b0 , \1029_A[17]_b0 , w_2113 );
and ( w_2112 , w_2113 , \1030_B[17]_b0 );
buf ( \1032_A[16]_b1 , \a[16]_b1 );
buf ( \1032_A[16]_b0 , \a[16]_b0 );
buf ( \1033_B[16]_b1 , \b[16]_b1 );
buf ( \1033_B[16]_b0 , \b[16]_b0 );
or ( \1034_b1 , \1032_A[16]_b1 , \1033_B[16]_b1 );
not ( \1033_B[16]_b1 , w_2114 );
and ( \1034_b0 , \1032_A[16]_b0 , w_2115 );
and ( w_2114 , w_2115 , \1033_B[16]_b0 );
buf ( \1035_A[15]_b1 , \a[15]_b1 );
buf ( \1035_A[15]_b0 , \a[15]_b0 );
buf ( \1036_B[15]_b1 , \b[15]_b1 );
buf ( \1036_B[15]_b0 , \b[15]_b0 );
or ( \1037_b1 , \1035_A[15]_b1 , \1036_B[15]_b1 );
not ( \1036_B[15]_b1 , w_2116 );
and ( \1037_b0 , \1035_A[15]_b0 , w_2117 );
and ( w_2116 , w_2117 , \1036_B[15]_b0 );
buf ( \1038_A[14]_b1 , \a[14]_b1 );
buf ( \1038_A[14]_b0 , \a[14]_b0 );
buf ( \1039_B[14]_b1 , \b[14]_b1 );
buf ( \1039_B[14]_b0 , \b[14]_b0 );
or ( \1040_b1 , \1038_A[14]_b1 , \1039_B[14]_b1 );
not ( \1039_B[14]_b1 , w_2118 );
and ( \1040_b0 , \1038_A[14]_b0 , w_2119 );
and ( w_2118 , w_2119 , \1039_B[14]_b0 );
buf ( \1041_A[13]_b1 , \a[13]_b1 );
buf ( \1041_A[13]_b0 , \a[13]_b0 );
buf ( \1042_B[13]_b1 , \b[13]_b1 );
buf ( \1042_B[13]_b0 , \b[13]_b0 );
or ( \1043_b1 , \1041_A[13]_b1 , \1042_B[13]_b1 );
not ( \1042_B[13]_b1 , w_2120 );
and ( \1043_b0 , \1041_A[13]_b0 , w_2121 );
and ( w_2120 , w_2121 , \1042_B[13]_b0 );
buf ( \1044_A[12]_b1 , \a[12]_b1 );
buf ( \1044_A[12]_b0 , \a[12]_b0 );
buf ( \1045_B[12]_b1 , \b[12]_b1 );
buf ( \1045_B[12]_b0 , \b[12]_b0 );
or ( \1046_b1 , \1044_A[12]_b1 , \1045_B[12]_b1 );
not ( \1045_B[12]_b1 , w_2122 );
and ( \1046_b0 , \1044_A[12]_b0 , w_2123 );
and ( w_2122 , w_2123 , \1045_B[12]_b0 );
buf ( \1047_A[11]_b1 , \a[11]_b1 );
buf ( \1047_A[11]_b0 , \a[11]_b0 );
buf ( \1048_B[11]_b1 , \b[11]_b1 );
buf ( \1048_B[11]_b0 , \b[11]_b0 );
or ( \1049_b1 , \1047_A[11]_b1 , \1048_B[11]_b1 );
not ( \1048_B[11]_b1 , w_2124 );
and ( \1049_b0 , \1047_A[11]_b0 , w_2125 );
and ( w_2124 , w_2125 , \1048_B[11]_b0 );
buf ( \1050_A[10]_b1 , \a[10]_b1 );
buf ( \1050_A[10]_b0 , \a[10]_b0 );
buf ( \1051_B[10]_b1 , \b[10]_b1 );
buf ( \1051_B[10]_b0 , \b[10]_b0 );
or ( \1052_b1 , \1050_A[10]_b1 , \1051_B[10]_b1 );
not ( \1051_B[10]_b1 , w_2126 );
and ( \1052_b0 , \1050_A[10]_b0 , w_2127 );
and ( w_2126 , w_2127 , \1051_B[10]_b0 );
buf ( \1053_A[9]_b1 , \a[9]_b1 );
buf ( \1053_A[9]_b0 , \a[9]_b0 );
buf ( \1054_B[9]_b1 , \b[9]_b1 );
buf ( \1054_B[9]_b0 , \b[9]_b0 );
or ( \1055_b1 , \1053_A[9]_b1 , \1054_B[9]_b1 );
not ( \1054_B[9]_b1 , w_2128 );
and ( \1055_b0 , \1053_A[9]_b0 , w_2129 );
and ( w_2128 , w_2129 , \1054_B[9]_b0 );
buf ( \1056_A[8]_b1 , \a[8]_b1 );
buf ( \1056_A[8]_b0 , \a[8]_b0 );
buf ( \1057_B[8]_b1 , \b[8]_b1 );
buf ( \1057_B[8]_b0 , \b[8]_b0 );
or ( \1058_b1 , \1056_A[8]_b1 , \1057_B[8]_b1 );
not ( \1057_B[8]_b1 , w_2130 );
and ( \1058_b0 , \1056_A[8]_b0 , w_2131 );
and ( w_2130 , w_2131 , \1057_B[8]_b0 );
buf ( \1059_A[7]_b1 , \a[7]_b1 );
buf ( \1059_A[7]_b0 , \a[7]_b0 );
buf ( \1060_B[7]_b1 , \b[7]_b1 );
buf ( \1060_B[7]_b0 , \b[7]_b0 );
or ( \1061_b1 , \1059_A[7]_b1 , \1060_B[7]_b1 );
not ( \1060_B[7]_b1 , w_2132 );
and ( \1061_b0 , \1059_A[7]_b0 , w_2133 );
and ( w_2132 , w_2133 , \1060_B[7]_b0 );
buf ( \1062_A[6]_b1 , \a[6]_b1 );
buf ( \1062_A[6]_b0 , \a[6]_b0 );
buf ( \1063_B[6]_b1 , \b[6]_b1 );
buf ( \1063_B[6]_b0 , \b[6]_b0 );
or ( \1064_b1 , \1062_A[6]_b1 , \1063_B[6]_b1 );
not ( \1063_B[6]_b1 , w_2134 );
and ( \1064_b0 , \1062_A[6]_b0 , w_2135 );
and ( w_2134 , w_2135 , \1063_B[6]_b0 );
buf ( \1065_A[5]_b1 , \a[5]_b1 );
buf ( \1065_A[5]_b0 , \a[5]_b0 );
buf ( \1066_B[5]_b1 , \b[5]_b1 );
buf ( \1066_B[5]_b0 , \b[5]_b0 );
or ( \1067_b1 , \1065_A[5]_b1 , \1066_B[5]_b1 );
not ( \1066_B[5]_b1 , w_2136 );
and ( \1067_b0 , \1065_A[5]_b0 , w_2137 );
and ( w_2136 , w_2137 , \1066_B[5]_b0 );
buf ( \1068_A[4]_b1 , \a[4]_b1 );
buf ( \1068_A[4]_b0 , \a[4]_b0 );
buf ( \1069_B[4]_b1 , \b[4]_b1 );
buf ( \1069_B[4]_b0 , \b[4]_b0 );
or ( \1070_b1 , \1068_A[4]_b1 , \1069_B[4]_b1 );
not ( \1069_B[4]_b1 , w_2138 );
and ( \1070_b0 , \1068_A[4]_b0 , w_2139 );
and ( w_2138 , w_2139 , \1069_B[4]_b0 );
buf ( \1071_A[3]_b1 , \a[3]_b1 );
buf ( \1071_A[3]_b0 , \a[3]_b0 );
buf ( \1072_B[3]_b1 , \b[3]_b1 );
buf ( \1072_B[3]_b0 , \b[3]_b0 );
or ( \1073_b1 , \1071_A[3]_b1 , \1072_B[3]_b1 );
not ( \1072_B[3]_b1 , w_2140 );
and ( \1073_b0 , \1071_A[3]_b0 , w_2141 );
and ( w_2140 , w_2141 , \1072_B[3]_b0 );
buf ( \1074_A[2]_b1 , \a[2]_b1 );
buf ( \1074_A[2]_b0 , \a[2]_b0 );
buf ( \1075_B[2]_b1 , \b[2]_b1 );
buf ( \1075_B[2]_b0 , \b[2]_b0 );
or ( \1076_b1 , \1074_A[2]_b1 , \1075_B[2]_b1 );
not ( \1075_B[2]_b1 , w_2142 );
and ( \1076_b0 , \1074_A[2]_b0 , w_2143 );
and ( w_2142 , w_2143 , \1075_B[2]_b0 );
buf ( \1077_A[1]_b1 , \a[1]_b1 );
buf ( \1077_A[1]_b0 , \a[1]_b0 );
buf ( \1078_B[1]_b1 , \b[1]_b1 );
buf ( \1078_B[1]_b0 , \b[1]_b0 );
or ( \1079_b1 , \1077_A[1]_b1 , \1078_B[1]_b1 );
not ( \1078_B[1]_b1 , w_2144 );
and ( \1079_b0 , \1077_A[1]_b0 , w_2145 );
and ( w_2144 , w_2145 , \1078_B[1]_b0 );
buf ( \1080_A[0]_b1 , \a[0]_b1 );
buf ( \1080_A[0]_b0 , \a[0]_b0 );
buf ( \1081_B[0]_b1 , \b[0]_b1 );
buf ( \1081_B[0]_b0 , \b[0]_b0 );
or ( \1082_b1 , \1080_A[0]_b1 , \1081_B[0]_b1 );
not ( \1081_B[0]_b1 , w_2146 );
and ( \1082_b0 , \1080_A[0]_b0 , w_2147 );
and ( w_2146 , w_2147 , \1081_B[0]_b0 );
or ( \1083_b1 , \1078_B[1]_b1 , \1082_b1 );
not ( \1082_b1 , w_2148 );
and ( \1083_b0 , \1078_B[1]_b0 , w_2149 );
and ( w_2148 , w_2149 , \1082_b0 );
or ( \1084_b1 , \1077_A[1]_b1 , \1082_b1 );
not ( \1082_b1 , w_2150 );
and ( \1084_b0 , \1077_A[1]_b0 , w_2151 );
and ( w_2150 , w_2151 , \1082_b0 );
or ( \1086_b1 , \1075_B[2]_b1 , \1085_b1 );
not ( \1085_b1 , w_2152 );
and ( \1086_b0 , \1075_B[2]_b0 , w_2153 );
and ( w_2152 , w_2153 , \1085_b0 );
or ( \1087_b1 , \1074_A[2]_b1 , \1085_b1 );
not ( \1085_b1 , w_2154 );
and ( \1087_b0 , \1074_A[2]_b0 , w_2155 );
and ( w_2154 , w_2155 , \1085_b0 );
or ( \1089_b1 , \1072_B[3]_b1 , \1088_b1 );
not ( \1088_b1 , w_2156 );
and ( \1089_b0 , \1072_B[3]_b0 , w_2157 );
and ( w_2156 , w_2157 , \1088_b0 );
or ( \1090_b1 , \1071_A[3]_b1 , \1088_b1 );
not ( \1088_b1 , w_2158 );
and ( \1090_b0 , \1071_A[3]_b0 , w_2159 );
and ( w_2158 , w_2159 , \1088_b0 );
or ( \1092_b1 , \1069_B[4]_b1 , \1091_b1 );
not ( \1091_b1 , w_2160 );
and ( \1092_b0 , \1069_B[4]_b0 , w_2161 );
and ( w_2160 , w_2161 , \1091_b0 );
or ( \1093_b1 , \1068_A[4]_b1 , \1091_b1 );
not ( \1091_b1 , w_2162 );
and ( \1093_b0 , \1068_A[4]_b0 , w_2163 );
and ( w_2162 , w_2163 , \1091_b0 );
or ( \1095_b1 , \1066_B[5]_b1 , \1094_b1 );
not ( \1094_b1 , w_2164 );
and ( \1095_b0 , \1066_B[5]_b0 , w_2165 );
and ( w_2164 , w_2165 , \1094_b0 );
or ( \1096_b1 , \1065_A[5]_b1 , \1094_b1 );
not ( \1094_b1 , w_2166 );
and ( \1096_b0 , \1065_A[5]_b0 , w_2167 );
and ( w_2166 , w_2167 , \1094_b0 );
or ( \1098_b1 , \1063_B[6]_b1 , \1097_b1 );
not ( \1097_b1 , w_2168 );
and ( \1098_b0 , \1063_B[6]_b0 , w_2169 );
and ( w_2168 , w_2169 , \1097_b0 );
or ( \1099_b1 , \1062_A[6]_b1 , \1097_b1 );
not ( \1097_b1 , w_2170 );
and ( \1099_b0 , \1062_A[6]_b0 , w_2171 );
and ( w_2170 , w_2171 , \1097_b0 );
or ( \1101_b1 , \1060_B[7]_b1 , \1100_b1 );
not ( \1100_b1 , w_2172 );
and ( \1101_b0 , \1060_B[7]_b0 , w_2173 );
and ( w_2172 , w_2173 , \1100_b0 );
or ( \1102_b1 , \1059_A[7]_b1 , \1100_b1 );
not ( \1100_b1 , w_2174 );
and ( \1102_b0 , \1059_A[7]_b0 , w_2175 );
and ( w_2174 , w_2175 , \1100_b0 );
or ( \1104_b1 , \1057_B[8]_b1 , \1103_b1 );
not ( \1103_b1 , w_2176 );
and ( \1104_b0 , \1057_B[8]_b0 , w_2177 );
and ( w_2176 , w_2177 , \1103_b0 );
or ( \1105_b1 , \1056_A[8]_b1 , \1103_b1 );
not ( \1103_b1 , w_2178 );
and ( \1105_b0 , \1056_A[8]_b0 , w_2179 );
and ( w_2178 , w_2179 , \1103_b0 );
or ( \1107_b1 , \1054_B[9]_b1 , \1106_b1 );
not ( \1106_b1 , w_2180 );
and ( \1107_b0 , \1054_B[9]_b0 , w_2181 );
and ( w_2180 , w_2181 , \1106_b0 );
or ( \1108_b1 , \1053_A[9]_b1 , \1106_b1 );
not ( \1106_b1 , w_2182 );
and ( \1108_b0 , \1053_A[9]_b0 , w_2183 );
and ( w_2182 , w_2183 , \1106_b0 );
or ( \1110_b1 , \1051_B[10]_b1 , \1109_b1 );
not ( \1109_b1 , w_2184 );
and ( \1110_b0 , \1051_B[10]_b0 , w_2185 );
and ( w_2184 , w_2185 , \1109_b0 );
or ( \1111_b1 , \1050_A[10]_b1 , \1109_b1 );
not ( \1109_b1 , w_2186 );
and ( \1111_b0 , \1050_A[10]_b0 , w_2187 );
and ( w_2186 , w_2187 , \1109_b0 );
or ( \1113_b1 , \1048_B[11]_b1 , \1112_b1 );
not ( \1112_b1 , w_2188 );
and ( \1113_b0 , \1048_B[11]_b0 , w_2189 );
and ( w_2188 , w_2189 , \1112_b0 );
or ( \1114_b1 , \1047_A[11]_b1 , \1112_b1 );
not ( \1112_b1 , w_2190 );
and ( \1114_b0 , \1047_A[11]_b0 , w_2191 );
and ( w_2190 , w_2191 , \1112_b0 );
or ( \1116_b1 , \1045_B[12]_b1 , \1115_b1 );
not ( \1115_b1 , w_2192 );
and ( \1116_b0 , \1045_B[12]_b0 , w_2193 );
and ( w_2192 , w_2193 , \1115_b0 );
or ( \1117_b1 , \1044_A[12]_b1 , \1115_b1 );
not ( \1115_b1 , w_2194 );
and ( \1117_b0 , \1044_A[12]_b0 , w_2195 );
and ( w_2194 , w_2195 , \1115_b0 );
or ( \1119_b1 , \1042_B[13]_b1 , \1118_b1 );
not ( \1118_b1 , w_2196 );
and ( \1119_b0 , \1042_B[13]_b0 , w_2197 );
and ( w_2196 , w_2197 , \1118_b0 );
or ( \1120_b1 , \1041_A[13]_b1 , \1118_b1 );
not ( \1118_b1 , w_2198 );
and ( \1120_b0 , \1041_A[13]_b0 , w_2199 );
and ( w_2198 , w_2199 , \1118_b0 );
or ( \1122_b1 , \1039_B[14]_b1 , \1121_b1 );
not ( \1121_b1 , w_2200 );
and ( \1122_b0 , \1039_B[14]_b0 , w_2201 );
and ( w_2200 , w_2201 , \1121_b0 );
or ( \1123_b1 , \1038_A[14]_b1 , \1121_b1 );
not ( \1121_b1 , w_2202 );
and ( \1123_b0 , \1038_A[14]_b0 , w_2203 );
and ( w_2202 , w_2203 , \1121_b0 );
or ( \1125_b1 , \1036_B[15]_b1 , \1124_b1 );
not ( \1124_b1 , w_2204 );
and ( \1125_b0 , \1036_B[15]_b0 , w_2205 );
and ( w_2204 , w_2205 , \1124_b0 );
or ( \1126_b1 , \1035_A[15]_b1 , \1124_b1 );
not ( \1124_b1 , w_2206 );
and ( \1126_b0 , \1035_A[15]_b0 , w_2207 );
and ( w_2206 , w_2207 , \1124_b0 );
or ( \1128_b1 , \1033_B[16]_b1 , \1127_b1 );
not ( \1127_b1 , w_2208 );
and ( \1128_b0 , \1033_B[16]_b0 , w_2209 );
and ( w_2208 , w_2209 , \1127_b0 );
or ( \1129_b1 , \1032_A[16]_b1 , \1127_b1 );
not ( \1127_b1 , w_2210 );
and ( \1129_b0 , \1032_A[16]_b0 , w_2211 );
and ( w_2210 , w_2211 , \1127_b0 );
or ( \1131_b1 , \1030_B[17]_b1 , \1130_b1 );
not ( \1130_b1 , w_2212 );
and ( \1131_b0 , \1030_B[17]_b0 , w_2213 );
and ( w_2212 , w_2213 , \1130_b0 );
or ( \1132_b1 , \1029_A[17]_b1 , \1130_b1 );
not ( \1130_b1 , w_2214 );
and ( \1132_b0 , \1029_A[17]_b0 , w_2215 );
and ( w_2214 , w_2215 , \1130_b0 );
or ( \1134_b1 , \1027_B[18]_b1 , \1133_b1 );
not ( \1133_b1 , w_2216 );
and ( \1134_b0 , \1027_B[18]_b0 , w_2217 );
and ( w_2216 , w_2217 , \1133_b0 );
or ( \1135_b1 , \1026_A[18]_b1 , \1133_b1 );
not ( \1133_b1 , w_2218 );
and ( \1135_b0 , \1026_A[18]_b0 , w_2219 );
and ( w_2218 , w_2219 , \1133_b0 );
or ( \1137_b1 , \1024_B[19]_b1 , \1136_b1 );
not ( \1136_b1 , w_2220 );
and ( \1137_b0 , \1024_B[19]_b0 , w_2221 );
and ( w_2220 , w_2221 , \1136_b0 );
or ( \1138_b1 , \1023_A[19]_b1 , \1136_b1 );
not ( \1136_b1 , w_2222 );
and ( \1138_b0 , \1023_A[19]_b0 , w_2223 );
and ( w_2222 , w_2223 , \1136_b0 );
or ( \1140_b1 , \1021_B[20]_b1 , \1139_b1 );
not ( \1139_b1 , w_2224 );
and ( \1140_b0 , \1021_B[20]_b0 , w_2225 );
and ( w_2224 , w_2225 , \1139_b0 );
or ( \1141_b1 , \1020_A[20]_b1 , \1139_b1 );
not ( \1139_b1 , w_2226 );
and ( \1141_b0 , \1020_A[20]_b0 , w_2227 );
and ( w_2226 , w_2227 , \1139_b0 );
or ( \1143_b1 , \1018_B[21]_b1 , \1142_b1 );
not ( \1142_b1 , w_2228 );
and ( \1143_b0 , \1018_B[21]_b0 , w_2229 );
and ( w_2228 , w_2229 , \1142_b0 );
or ( \1144_b1 , \1017_A[21]_b1 , \1142_b1 );
not ( \1142_b1 , w_2230 );
and ( \1144_b0 , \1017_A[21]_b0 , w_2231 );
and ( w_2230 , w_2231 , \1142_b0 );
or ( \1146_b1 , \1015_B[22]_b1 , \1145_b1 );
not ( \1145_b1 , w_2232 );
and ( \1146_b0 , \1015_B[22]_b0 , w_2233 );
and ( w_2232 , w_2233 , \1145_b0 );
or ( \1147_b1 , \1014_A[22]_b1 , \1145_b1 );
not ( \1145_b1 , w_2234 );
and ( \1147_b0 , \1014_A[22]_b0 , w_2235 );
and ( w_2234 , w_2235 , \1145_b0 );
or ( \1149_b1 , \1012_B[23]_b1 , \1148_b1 );
not ( \1148_b1 , w_2236 );
and ( \1149_b0 , \1012_B[23]_b0 , w_2237 );
and ( w_2236 , w_2237 , \1148_b0 );
or ( \1150_b1 , \1011_A[23]_b1 , \1148_b1 );
not ( \1148_b1 , w_2238 );
and ( \1150_b0 , \1011_A[23]_b0 , w_2239 );
and ( w_2238 , w_2239 , \1148_b0 );
or ( \1152_b1 , \1009_B[24]_b1 , \1151_b1 );
not ( \1151_b1 , w_2240 );
and ( \1152_b0 , \1009_B[24]_b0 , w_2241 );
and ( w_2240 , w_2241 , \1151_b0 );
or ( \1153_b1 , \1008_A[24]_b1 , \1151_b1 );
not ( \1151_b1 , w_2242 );
and ( \1153_b0 , \1008_A[24]_b0 , w_2243 );
and ( w_2242 , w_2243 , \1151_b0 );
or ( \1155_b1 , \1006_B[25]_b1 , \1154_b1 );
not ( \1154_b1 , w_2244 );
and ( \1155_b0 , \1006_B[25]_b0 , w_2245 );
and ( w_2244 , w_2245 , \1154_b0 );
or ( \1156_b1 , \1005_A[25]_b1 , \1154_b1 );
not ( \1154_b1 , w_2246 );
and ( \1156_b0 , \1005_A[25]_b0 , w_2247 );
and ( w_2246 , w_2247 , \1154_b0 );
or ( \1158_b1 , \1003_B[26]_b1 , \1157_b1 );
not ( \1157_b1 , w_2248 );
and ( \1158_b0 , \1003_B[26]_b0 , w_2249 );
and ( w_2248 , w_2249 , \1157_b0 );
or ( \1159_b1 , \1002_A[26]_b1 , \1157_b1 );
not ( \1157_b1 , w_2250 );
and ( \1159_b0 , \1002_A[26]_b0 , w_2251 );
and ( w_2250 , w_2251 , \1157_b0 );
or ( \1161_b1 , \1000_B[27]_b1 , \1160_b1 );
not ( \1160_b1 , w_2252 );
and ( \1161_b0 , \1000_B[27]_b0 , w_2253 );
and ( w_2252 , w_2253 , \1160_b0 );
or ( \1162_b1 , \999_A[27]_b1 , \1160_b1 );
not ( \1160_b1 , w_2254 );
and ( \1162_b0 , \999_A[27]_b0 , w_2255 );
and ( w_2254 , w_2255 , \1160_b0 );
or ( \1164_b1 , \997_B[28]_b1 , \1163_b1 );
not ( \1163_b1 , w_2256 );
and ( \1164_b0 , \997_B[28]_b0 , w_2257 );
and ( w_2256 , w_2257 , \1163_b0 );
or ( \1165_b1 , \996_A[28]_b1 , \1163_b1 );
not ( \1163_b1 , w_2258 );
and ( \1165_b0 , \996_A[28]_b0 , w_2259 );
and ( w_2258 , w_2259 , \1163_b0 );
or ( \1167_b1 , \994_B[29]_b1 , \1166_b1 );
not ( \1166_b1 , w_2260 );
and ( \1167_b0 , \994_B[29]_b0 , w_2261 );
and ( w_2260 , w_2261 , \1166_b0 );
or ( \1168_b1 , \993_A[29]_b1 , \1166_b1 );
not ( \1166_b1 , w_2262 );
and ( \1168_b0 , \993_A[29]_b0 , w_2263 );
and ( w_2262 , w_2263 , \1166_b0 );
or ( \1170_b1 , \991_B[30]_b1 , \1169_b1 );
not ( \1169_b1 , w_2264 );
and ( \1170_b0 , \991_B[30]_b0 , w_2265 );
and ( w_2264 , w_2265 , \1169_b0 );
or ( \1171_b1 , \990_A[30]_b1 , \1169_b1 );
not ( \1169_b1 , w_2266 );
and ( \1171_b0 , \990_A[30]_b0 , w_2267 );
and ( w_2266 , w_2267 , \1169_b0 );
or ( \1173_b1 , \989_b1 , \1172_b1 );
xor ( \1173_b0 , \989_b0 , w_2268 );
not ( w_2268 , w_2269 );
and ( w_2269 , \1172_b1 , \1172_b0 );
buf ( \1174_SUM[31]_b1 , \1173_b1 );
buf ( \1174_SUM[31]_b0 , \1173_b0 );
buf ( \1175_A[31]_b1 , \1174_SUM[31]_b1 );
buf ( \1175_A[31]_b0 , \1174_SUM[31]_b0 );
or ( \1176_b1 , \990_A[30]_b1 , \991_B[30]_b1 );
xor ( \1176_b0 , \990_A[30]_b0 , w_2270 );
not ( w_2270 , w_2271 );
and ( w_2271 , \991_B[30]_b1 , \991_B[30]_b0 );
or ( \1177_b1 , \1176_b1 , \1169_b1 );
xor ( \1177_b0 , \1176_b0 , w_2272 );
not ( w_2272 , w_2273 );
and ( w_2273 , \1169_b1 , \1169_b0 );
buf ( \1178_SUM[30]_b1 , \1177_b1 );
buf ( \1178_SUM[30]_b0 , \1177_b0 );
buf ( \1179_A[30]_b1 , \1178_SUM[30]_b1 );
buf ( \1179_A[30]_b0 , \1178_SUM[30]_b0 );
or ( \1180_b1 , \993_A[29]_b1 , \994_B[29]_b1 );
xor ( \1180_b0 , \993_A[29]_b0 , w_2274 );
not ( w_2274 , w_2275 );
and ( w_2275 , \994_B[29]_b1 , \994_B[29]_b0 );
or ( \1181_b1 , \1180_b1 , \1166_b1 );
xor ( \1181_b0 , \1180_b0 , w_2276 );
not ( w_2276 , w_2277 );
and ( w_2277 , \1166_b1 , \1166_b0 );
buf ( \1182_SUM[29]_b1 , \1181_b1 );
buf ( \1182_SUM[29]_b0 , \1181_b0 );
buf ( \1183_A[29]_b1 , \1182_SUM[29]_b1 );
buf ( \1183_A[29]_b0 , \1182_SUM[29]_b0 );
or ( \1184_b1 , \996_A[28]_b1 , \997_B[28]_b1 );
xor ( \1184_b0 , \996_A[28]_b0 , w_2278 );
not ( w_2278 , w_2279 );
and ( w_2279 , \997_B[28]_b1 , \997_B[28]_b0 );
or ( \1185_b1 , \1184_b1 , \1163_b1 );
xor ( \1185_b0 , \1184_b0 , w_2280 );
not ( w_2280 , w_2281 );
and ( w_2281 , \1163_b1 , \1163_b0 );
buf ( \1186_SUM[28]_b1 , \1185_b1 );
buf ( \1186_SUM[28]_b0 , \1185_b0 );
buf ( \1187_A[28]_b1 , \1186_SUM[28]_b1 );
buf ( \1187_A[28]_b0 , \1186_SUM[28]_b0 );
or ( \1188_b1 , \999_A[27]_b1 , \1000_B[27]_b1 );
xor ( \1188_b0 , \999_A[27]_b0 , w_2282 );
not ( w_2282 , w_2283 );
and ( w_2283 , \1000_B[27]_b1 , \1000_B[27]_b0 );
or ( \1189_b1 , \1188_b1 , \1160_b1 );
xor ( \1189_b0 , \1188_b0 , w_2284 );
not ( w_2284 , w_2285 );
and ( w_2285 , \1160_b1 , \1160_b0 );
buf ( \1190_SUM[27]_b1 , \1189_b1 );
buf ( \1190_SUM[27]_b0 , \1189_b0 );
buf ( \1191_A[27]_b1 , \1190_SUM[27]_b1 );
buf ( \1191_A[27]_b0 , \1190_SUM[27]_b0 );
or ( \1192_b1 , \1002_A[26]_b1 , \1003_B[26]_b1 );
xor ( \1192_b0 , \1002_A[26]_b0 , w_2286 );
not ( w_2286 , w_2287 );
and ( w_2287 , \1003_B[26]_b1 , \1003_B[26]_b0 );
or ( \1193_b1 , \1192_b1 , \1157_b1 );
xor ( \1193_b0 , \1192_b0 , w_2288 );
not ( w_2288 , w_2289 );
and ( w_2289 , \1157_b1 , \1157_b0 );
buf ( \1194_SUM[26]_b1 , \1193_b1 );
buf ( \1194_SUM[26]_b0 , \1193_b0 );
buf ( \1195_A[26]_b1 , \1194_SUM[26]_b1 );
buf ( \1195_A[26]_b0 , \1194_SUM[26]_b0 );
or ( \1196_b1 , \1005_A[25]_b1 , \1006_B[25]_b1 );
xor ( \1196_b0 , \1005_A[25]_b0 , w_2290 );
not ( w_2290 , w_2291 );
and ( w_2291 , \1006_B[25]_b1 , \1006_B[25]_b0 );
or ( \1197_b1 , \1196_b1 , \1154_b1 );
xor ( \1197_b0 , \1196_b0 , w_2292 );
not ( w_2292 , w_2293 );
and ( w_2293 , \1154_b1 , \1154_b0 );
buf ( \1198_SUM[25]_b1 , \1197_b1 );
buf ( \1198_SUM[25]_b0 , \1197_b0 );
buf ( \1199_A[25]_b1 , \1198_SUM[25]_b1 );
buf ( \1199_A[25]_b0 , \1198_SUM[25]_b0 );
or ( \1200_b1 , \1008_A[24]_b1 , \1009_B[24]_b1 );
xor ( \1200_b0 , \1008_A[24]_b0 , w_2294 );
not ( w_2294 , w_2295 );
and ( w_2295 , \1009_B[24]_b1 , \1009_B[24]_b0 );
or ( \1201_b1 , \1200_b1 , \1151_b1 );
xor ( \1201_b0 , \1200_b0 , w_2296 );
not ( w_2296 , w_2297 );
and ( w_2297 , \1151_b1 , \1151_b0 );
buf ( \1202_SUM[24]_b1 , \1201_b1 );
buf ( \1202_SUM[24]_b0 , \1201_b0 );
buf ( \1203_A[24]_b1 , \1202_SUM[24]_b1 );
buf ( \1203_A[24]_b0 , \1202_SUM[24]_b0 );
or ( \1204_b1 , \1011_A[23]_b1 , \1012_B[23]_b1 );
xor ( \1204_b0 , \1011_A[23]_b0 , w_2298 );
not ( w_2298 , w_2299 );
and ( w_2299 , \1012_B[23]_b1 , \1012_B[23]_b0 );
or ( \1205_b1 , \1204_b1 , \1148_b1 );
xor ( \1205_b0 , \1204_b0 , w_2300 );
not ( w_2300 , w_2301 );
and ( w_2301 , \1148_b1 , \1148_b0 );
buf ( \1206_SUM[23]_b1 , \1205_b1 );
buf ( \1206_SUM[23]_b0 , \1205_b0 );
buf ( \1207_A[23]_b1 , \1206_SUM[23]_b1 );
buf ( \1207_A[23]_b0 , \1206_SUM[23]_b0 );
or ( \1208_b1 , \1014_A[22]_b1 , \1015_B[22]_b1 );
xor ( \1208_b0 , \1014_A[22]_b0 , w_2302 );
not ( w_2302 , w_2303 );
and ( w_2303 , \1015_B[22]_b1 , \1015_B[22]_b0 );
or ( \1209_b1 , \1208_b1 , \1145_b1 );
xor ( \1209_b0 , \1208_b0 , w_2304 );
not ( w_2304 , w_2305 );
and ( w_2305 , \1145_b1 , \1145_b0 );
buf ( \1210_SUM[22]_b1 , \1209_b1 );
buf ( \1210_SUM[22]_b0 , \1209_b0 );
buf ( \1211_A[22]_b1 , \1210_SUM[22]_b1 );
buf ( \1211_A[22]_b0 , \1210_SUM[22]_b0 );
or ( \1212_b1 , \1017_A[21]_b1 , \1018_B[21]_b1 );
xor ( \1212_b0 , \1017_A[21]_b0 , w_2306 );
not ( w_2306 , w_2307 );
and ( w_2307 , \1018_B[21]_b1 , \1018_B[21]_b0 );
or ( \1213_b1 , \1212_b1 , \1142_b1 );
xor ( \1213_b0 , \1212_b0 , w_2308 );
not ( w_2308 , w_2309 );
and ( w_2309 , \1142_b1 , \1142_b0 );
buf ( \1214_SUM[21]_b1 , \1213_b1 );
buf ( \1214_SUM[21]_b0 , \1213_b0 );
buf ( \1215_A[21]_b1 , \1214_SUM[21]_b1 );
buf ( \1215_A[21]_b0 , \1214_SUM[21]_b0 );
or ( \1216_b1 , \1020_A[20]_b1 , \1021_B[20]_b1 );
xor ( \1216_b0 , \1020_A[20]_b0 , w_2310 );
not ( w_2310 , w_2311 );
and ( w_2311 , \1021_B[20]_b1 , \1021_B[20]_b0 );
or ( \1217_b1 , \1216_b1 , \1139_b1 );
xor ( \1217_b0 , \1216_b0 , w_2312 );
not ( w_2312 , w_2313 );
and ( w_2313 , \1139_b1 , \1139_b0 );
buf ( \1218_SUM[20]_b1 , \1217_b1 );
buf ( \1218_SUM[20]_b0 , \1217_b0 );
buf ( \1219_A[20]_b1 , \1218_SUM[20]_b1 );
buf ( \1219_A[20]_b0 , \1218_SUM[20]_b0 );
or ( \1220_b1 , \1023_A[19]_b1 , \1024_B[19]_b1 );
xor ( \1220_b0 , \1023_A[19]_b0 , w_2314 );
not ( w_2314 , w_2315 );
and ( w_2315 , \1024_B[19]_b1 , \1024_B[19]_b0 );
or ( \1221_b1 , \1220_b1 , \1136_b1 );
xor ( \1221_b0 , \1220_b0 , w_2316 );
not ( w_2316 , w_2317 );
and ( w_2317 , \1136_b1 , \1136_b0 );
buf ( \1222_SUM[19]_b1 , \1221_b1 );
buf ( \1222_SUM[19]_b0 , \1221_b0 );
buf ( \1223_A[19]_b1 , \1222_SUM[19]_b1 );
buf ( \1223_A[19]_b0 , \1222_SUM[19]_b0 );
or ( \1224_b1 , \1026_A[18]_b1 , \1027_B[18]_b1 );
xor ( \1224_b0 , \1026_A[18]_b0 , w_2318 );
not ( w_2318 , w_2319 );
and ( w_2319 , \1027_B[18]_b1 , \1027_B[18]_b0 );
or ( \1225_b1 , \1224_b1 , \1133_b1 );
xor ( \1225_b0 , \1224_b0 , w_2320 );
not ( w_2320 , w_2321 );
and ( w_2321 , \1133_b1 , \1133_b0 );
buf ( \1226_SUM[18]_b1 , \1225_b1 );
buf ( \1226_SUM[18]_b0 , \1225_b0 );
buf ( \1227_A[18]_b1 , \1226_SUM[18]_b1 );
buf ( \1227_A[18]_b0 , \1226_SUM[18]_b0 );
or ( \1228_b1 , \1029_A[17]_b1 , \1030_B[17]_b1 );
xor ( \1228_b0 , \1029_A[17]_b0 , w_2322 );
not ( w_2322 , w_2323 );
and ( w_2323 , \1030_B[17]_b1 , \1030_B[17]_b0 );
or ( \1229_b1 , \1228_b1 , \1130_b1 );
xor ( \1229_b0 , \1228_b0 , w_2324 );
not ( w_2324 , w_2325 );
and ( w_2325 , \1130_b1 , \1130_b0 );
buf ( \1230_SUM[17]_b1 , \1229_b1 );
buf ( \1230_SUM[17]_b0 , \1229_b0 );
buf ( \1231_A[17]_b1 , \1230_SUM[17]_b1 );
buf ( \1231_A[17]_b0 , \1230_SUM[17]_b0 );
or ( \1232_b1 , \1032_A[16]_b1 , \1033_B[16]_b1 );
xor ( \1232_b0 , \1032_A[16]_b0 , w_2326 );
not ( w_2326 , w_2327 );
and ( w_2327 , \1033_B[16]_b1 , \1033_B[16]_b0 );
or ( \1233_b1 , \1232_b1 , \1127_b1 );
xor ( \1233_b0 , \1232_b0 , w_2328 );
not ( w_2328 , w_2329 );
and ( w_2329 , \1127_b1 , \1127_b0 );
buf ( \1234_SUM[16]_b1 , \1233_b1 );
buf ( \1234_SUM[16]_b0 , \1233_b0 );
buf ( \1235_A[16]_b1 , \1234_SUM[16]_b1 );
buf ( \1235_A[16]_b0 , \1234_SUM[16]_b0 );
or ( \1236_b1 , \1035_A[15]_b1 , \1036_B[15]_b1 );
xor ( \1236_b0 , \1035_A[15]_b0 , w_2330 );
not ( w_2330 , w_2331 );
and ( w_2331 , \1036_B[15]_b1 , \1036_B[15]_b0 );
or ( \1237_b1 , \1236_b1 , \1124_b1 );
xor ( \1237_b0 , \1236_b0 , w_2332 );
not ( w_2332 , w_2333 );
and ( w_2333 , \1124_b1 , \1124_b0 );
buf ( \1238_SUM[15]_b1 , \1237_b1 );
buf ( \1238_SUM[15]_b0 , \1237_b0 );
buf ( \1239_A[15]_b1 , \1238_SUM[15]_b1 );
buf ( \1239_A[15]_b0 , \1238_SUM[15]_b0 );
or ( \1240_b1 , \1038_A[14]_b1 , \1039_B[14]_b1 );
xor ( \1240_b0 , \1038_A[14]_b0 , w_2334 );
not ( w_2334 , w_2335 );
and ( w_2335 , \1039_B[14]_b1 , \1039_B[14]_b0 );
or ( \1241_b1 , \1240_b1 , \1121_b1 );
xor ( \1241_b0 , \1240_b0 , w_2336 );
not ( w_2336 , w_2337 );
and ( w_2337 , \1121_b1 , \1121_b0 );
buf ( \1242_SUM[14]_b1 , \1241_b1 );
buf ( \1242_SUM[14]_b0 , \1241_b0 );
buf ( \1243_A[14]_b1 , \1242_SUM[14]_b1 );
buf ( \1243_A[14]_b0 , \1242_SUM[14]_b0 );
or ( \1244_b1 , \1041_A[13]_b1 , \1042_B[13]_b1 );
xor ( \1244_b0 , \1041_A[13]_b0 , w_2338 );
not ( w_2338 , w_2339 );
and ( w_2339 , \1042_B[13]_b1 , \1042_B[13]_b0 );
or ( \1245_b1 , \1244_b1 , \1118_b1 );
xor ( \1245_b0 , \1244_b0 , w_2340 );
not ( w_2340 , w_2341 );
and ( w_2341 , \1118_b1 , \1118_b0 );
buf ( \1246_SUM[13]_b1 , \1245_b1 );
buf ( \1246_SUM[13]_b0 , \1245_b0 );
buf ( \1247_A[13]_b1 , \1246_SUM[13]_b1 );
buf ( \1247_A[13]_b0 , \1246_SUM[13]_b0 );
or ( \1248_b1 , \1044_A[12]_b1 , \1045_B[12]_b1 );
xor ( \1248_b0 , \1044_A[12]_b0 , w_2342 );
not ( w_2342 , w_2343 );
and ( w_2343 , \1045_B[12]_b1 , \1045_B[12]_b0 );
or ( \1249_b1 , \1248_b1 , \1115_b1 );
xor ( \1249_b0 , \1248_b0 , w_2344 );
not ( w_2344 , w_2345 );
and ( w_2345 , \1115_b1 , \1115_b0 );
buf ( \1250_SUM[12]_b1 , \1249_b1 );
buf ( \1250_SUM[12]_b0 , \1249_b0 );
buf ( \1251_A[12]_b1 , \1250_SUM[12]_b1 );
buf ( \1251_A[12]_b0 , \1250_SUM[12]_b0 );
or ( \1252_b1 , \1047_A[11]_b1 , \1048_B[11]_b1 );
xor ( \1252_b0 , \1047_A[11]_b0 , w_2346 );
not ( w_2346 , w_2347 );
and ( w_2347 , \1048_B[11]_b1 , \1048_B[11]_b0 );
or ( \1253_b1 , \1252_b1 , \1112_b1 );
xor ( \1253_b0 , \1252_b0 , w_2348 );
not ( w_2348 , w_2349 );
and ( w_2349 , \1112_b1 , \1112_b0 );
buf ( \1254_SUM[11]_b1 , \1253_b1 );
buf ( \1254_SUM[11]_b0 , \1253_b0 );
buf ( \1255_A[11]_b1 , \1254_SUM[11]_b1 );
buf ( \1255_A[11]_b0 , \1254_SUM[11]_b0 );
or ( \1256_b1 , \1050_A[10]_b1 , \1051_B[10]_b1 );
xor ( \1256_b0 , \1050_A[10]_b0 , w_2350 );
not ( w_2350 , w_2351 );
and ( w_2351 , \1051_B[10]_b1 , \1051_B[10]_b0 );
or ( \1257_b1 , \1256_b1 , \1109_b1 );
xor ( \1257_b0 , \1256_b0 , w_2352 );
not ( w_2352 , w_2353 );
and ( w_2353 , \1109_b1 , \1109_b0 );
buf ( \1258_SUM[10]_b1 , \1257_b1 );
buf ( \1258_SUM[10]_b0 , \1257_b0 );
buf ( \1259_A[10]_b1 , \1258_SUM[10]_b1 );
buf ( \1259_A[10]_b0 , \1258_SUM[10]_b0 );
or ( \1260_b1 , \1053_A[9]_b1 , \1054_B[9]_b1 );
xor ( \1260_b0 , \1053_A[9]_b0 , w_2354 );
not ( w_2354 , w_2355 );
and ( w_2355 , \1054_B[9]_b1 , \1054_B[9]_b0 );
or ( \1261_b1 , \1260_b1 , \1106_b1 );
xor ( \1261_b0 , \1260_b0 , w_2356 );
not ( w_2356 , w_2357 );
and ( w_2357 , \1106_b1 , \1106_b0 );
buf ( \1262_SUM[9]_b1 , \1261_b1 );
buf ( \1262_SUM[9]_b0 , \1261_b0 );
buf ( \1263_A[9]_b1 , \1262_SUM[9]_b1 );
buf ( \1263_A[9]_b0 , \1262_SUM[9]_b0 );
or ( \1264_b1 , \1056_A[8]_b1 , \1057_B[8]_b1 );
xor ( \1264_b0 , \1056_A[8]_b0 , w_2358 );
not ( w_2358 , w_2359 );
and ( w_2359 , \1057_B[8]_b1 , \1057_B[8]_b0 );
or ( \1265_b1 , \1264_b1 , \1103_b1 );
xor ( \1265_b0 , \1264_b0 , w_2360 );
not ( w_2360 , w_2361 );
and ( w_2361 , \1103_b1 , \1103_b0 );
buf ( \1266_SUM[8]_b1 , \1265_b1 );
buf ( \1266_SUM[8]_b0 , \1265_b0 );
buf ( \1267_A[8]_b1 , \1266_SUM[8]_b1 );
buf ( \1267_A[8]_b0 , \1266_SUM[8]_b0 );
or ( \1268_b1 , \1059_A[7]_b1 , \1060_B[7]_b1 );
xor ( \1268_b0 , \1059_A[7]_b0 , w_2362 );
not ( w_2362 , w_2363 );
and ( w_2363 , \1060_B[7]_b1 , \1060_B[7]_b0 );
or ( \1269_b1 , \1268_b1 , \1100_b1 );
xor ( \1269_b0 , \1268_b0 , w_2364 );
not ( w_2364 , w_2365 );
and ( w_2365 , \1100_b1 , \1100_b0 );
buf ( \1270_SUM[7]_b1 , \1269_b1 );
buf ( \1270_SUM[7]_b0 , \1269_b0 );
buf ( \1271_A[7]_b1 , \1270_SUM[7]_b1 );
buf ( \1271_A[7]_b0 , \1270_SUM[7]_b0 );
or ( \1272_b1 , \1062_A[6]_b1 , \1063_B[6]_b1 );
xor ( \1272_b0 , \1062_A[6]_b0 , w_2366 );
not ( w_2366 , w_2367 );
and ( w_2367 , \1063_B[6]_b1 , \1063_B[6]_b0 );
or ( \1273_b1 , \1272_b1 , \1097_b1 );
xor ( \1273_b0 , \1272_b0 , w_2368 );
not ( w_2368 , w_2369 );
and ( w_2369 , \1097_b1 , \1097_b0 );
buf ( \1274_SUM[6]_b1 , \1273_b1 );
buf ( \1274_SUM[6]_b0 , \1273_b0 );
buf ( \1275_A[6]_b1 , \1274_SUM[6]_b1 );
buf ( \1275_A[6]_b0 , \1274_SUM[6]_b0 );
or ( \1276_b1 , \1065_A[5]_b1 , \1066_B[5]_b1 );
xor ( \1276_b0 , \1065_A[5]_b0 , w_2370 );
not ( w_2370 , w_2371 );
and ( w_2371 , \1066_B[5]_b1 , \1066_B[5]_b0 );
or ( \1277_b1 , \1276_b1 , \1094_b1 );
xor ( \1277_b0 , \1276_b0 , w_2372 );
not ( w_2372 , w_2373 );
and ( w_2373 , \1094_b1 , \1094_b0 );
buf ( \1278_SUM[5]_b1 , \1277_b1 );
buf ( \1278_SUM[5]_b0 , \1277_b0 );
buf ( \1279_A[5]_b1 , \1278_SUM[5]_b1 );
buf ( \1279_A[5]_b0 , \1278_SUM[5]_b0 );
or ( \1280_b1 , \1068_A[4]_b1 , \1069_B[4]_b1 );
xor ( \1280_b0 , \1068_A[4]_b0 , w_2374 );
not ( w_2374 , w_2375 );
and ( w_2375 , \1069_B[4]_b1 , \1069_B[4]_b0 );
or ( \1281_b1 , \1280_b1 , \1091_b1 );
xor ( \1281_b0 , \1280_b0 , w_2376 );
not ( w_2376 , w_2377 );
and ( w_2377 , \1091_b1 , \1091_b0 );
buf ( \1282_SUM[4]_b1 , \1281_b1 );
buf ( \1282_SUM[4]_b0 , \1281_b0 );
buf ( \1283_A[4]_b1 , \1282_SUM[4]_b1 );
buf ( \1283_A[4]_b0 , \1282_SUM[4]_b0 );
or ( \1284_b1 , \1071_A[3]_b1 , \1072_B[3]_b1 );
xor ( \1284_b0 , \1071_A[3]_b0 , w_2378 );
not ( w_2378 , w_2379 );
and ( w_2379 , \1072_B[3]_b1 , \1072_B[3]_b0 );
or ( \1285_b1 , \1284_b1 , \1088_b1 );
xor ( \1285_b0 , \1284_b0 , w_2380 );
not ( w_2380 , w_2381 );
and ( w_2381 , \1088_b1 , \1088_b0 );
buf ( \1286_SUM[3]_b1 , \1285_b1 );
buf ( \1286_SUM[3]_b0 , \1285_b0 );
buf ( \1287_A[3]_b1 , \1286_SUM[3]_b1 );
buf ( \1287_A[3]_b0 , \1286_SUM[3]_b0 );
or ( \1288_b1 , \1074_A[2]_b1 , \1075_B[2]_b1 );
xor ( \1288_b0 , \1074_A[2]_b0 , w_2382 );
not ( w_2382 , w_2383 );
and ( w_2383 , \1075_B[2]_b1 , \1075_B[2]_b0 );
or ( \1289_b1 , \1288_b1 , \1085_b1 );
xor ( \1289_b0 , \1288_b0 , w_2384 );
not ( w_2384 , w_2385 );
and ( w_2385 , \1085_b1 , \1085_b0 );
buf ( \1290_SUM[2]_b1 , \1289_b1 );
buf ( \1290_SUM[2]_b0 , \1289_b0 );
buf ( \1291_A[2]_b1 , \1290_SUM[2]_b1 );
buf ( \1291_A[2]_b0 , \1290_SUM[2]_b0 );
or ( \1292_b1 , \1077_A[1]_b1 , \1078_B[1]_b1 );
xor ( \1292_b0 , \1077_A[1]_b0 , w_2386 );
not ( w_2386 , w_2387 );
and ( w_2387 , \1078_B[1]_b1 , \1078_B[1]_b0 );
or ( \1293_b1 , \1292_b1 , \1082_b1 );
xor ( \1293_b0 , \1292_b0 , w_2388 );
not ( w_2388 , w_2389 );
and ( w_2389 , \1082_b1 , \1082_b0 );
buf ( \1294_SUM[1]_b1 , \1293_b1 );
buf ( \1294_SUM[1]_b0 , \1293_b0 );
buf ( \1295_A[1]_b1 , \1294_SUM[1]_b1 );
buf ( \1295_A[1]_b0 , \1294_SUM[1]_b0 );
or ( \1296_b1 , \1080_A[0]_b1 , \1081_B[0]_b1 );
xor ( \1296_b0 , \1080_A[0]_b0 , w_2390 );
not ( w_2390 , w_2391 );
and ( w_2391 , \1081_B[0]_b1 , \1081_B[0]_b0 );
buf ( \1297_SUM[0]_b1 , \1296_b1 );
buf ( \1297_SUM[0]_b0 , \1296_b0 );
buf ( \1298_A[0]_b1 , \1297_SUM[0]_b1 );
buf ( \1298_A[0]_b0 , \1297_SUM[0]_b0 );
buf ( \1299_B[31]_b1 , \986_b1 );
buf ( \1299_B[31]_b0 , \986_b0 );
buf ( \1300_B[30]_b1 , \963_b1 );
buf ( \1300_B[30]_b0 , \963_b0 );
buf ( \1301_B[29]_b1 , \940_b1 );
buf ( \1301_B[29]_b0 , \940_b0 );
buf ( \1302_B[28]_b1 , \917_b1 );
buf ( \1302_B[28]_b0 , \917_b0 );
buf ( \1303_B[27]_b1 , \894_b1 );
buf ( \1303_B[27]_b0 , \894_b0 );
buf ( \1304_B[26]_b1 , \871_b1 );
buf ( \1304_B[26]_b0 , \871_b0 );
buf ( \1305_B[25]_b1 , \848_b1 );
buf ( \1305_B[25]_b0 , \848_b0 );
buf ( \1306_B[24]_b1 , \825_b1 );
buf ( \1306_B[24]_b0 , \825_b0 );
buf ( \1307_B[23]_b1 , \802_b1 );
buf ( \1307_B[23]_b0 , \802_b0 );
buf ( \1308_B[22]_b1 , \779_b1 );
buf ( \1308_B[22]_b0 , \779_b0 );
buf ( \1309_B[21]_b1 , \756_b1 );
buf ( \1309_B[21]_b0 , \756_b0 );
buf ( \1310_B[20]_b1 , \733_b1 );
buf ( \1310_B[20]_b0 , \733_b0 );
buf ( \1311_B[19]_b1 , \710_b1 );
buf ( \1311_B[19]_b0 , \710_b0 );
buf ( \1312_B[18]_b1 , \687_b1 );
buf ( \1312_B[18]_b0 , \687_b0 );
buf ( \1313_B[17]_b1 , \664_b1 );
buf ( \1313_B[17]_b0 , \664_b0 );
buf ( \1314_B[16]_b1 , \641_b1 );
buf ( \1314_B[16]_b0 , \641_b0 );
buf ( \1315_B[15]_b1 , \618_b1 );
buf ( \1315_B[15]_b0 , \618_b0 );
buf ( \1316_B[14]_b1 , \595_b1 );
buf ( \1316_B[14]_b0 , \595_b0 );
buf ( \1317_B[13]_b1 , \572_b1 );
buf ( \1317_B[13]_b0 , \572_b0 );
buf ( \1318_B[12]_b1 , \549_b1 );
buf ( \1318_B[12]_b0 , \549_b0 );
buf ( \1319_B[11]_b1 , \526_b1 );
buf ( \1319_B[11]_b0 , \526_b0 );
buf ( \1320_B[10]_b1 , \503_b1 );
buf ( \1320_B[10]_b0 , \503_b0 );
buf ( \1321_B[9]_b1 , \480_b1 );
buf ( \1321_B[9]_b0 , \480_b0 );
buf ( \1322_B[8]_b1 , \457_b1 );
buf ( \1322_B[8]_b0 , \457_b0 );
buf ( \1323_B[7]_b1 , \434_b1 );
buf ( \1323_B[7]_b0 , \434_b0 );
buf ( \1324_B[6]_b1 , \411_b1 );
buf ( \1324_B[6]_b0 , \411_b0 );
buf ( \1325_B[5]_b1 , \388_b1 );
buf ( \1325_B[5]_b0 , \388_b0 );
buf ( \1326_B[4]_b1 , \365_b1 );
buf ( \1326_B[4]_b0 , \365_b0 );
buf ( \1327_B[3]_b1 , \342_b1 );
buf ( \1327_B[3]_b0 , \342_b0 );
buf ( \1328_B[2]_b1 , \319_b1 );
buf ( \1328_B[2]_b0 , \319_b0 );
buf ( \1329_B[1]_b1 , \296_b1 );
buf ( \1329_B[1]_b0 , \296_b0 );
buf ( \1330_B[0]_b1 , \278_b1 );
buf ( \1330_B[0]_b0 , \278_b0 );
buf ( \1331_b1 , \1191_A[27]_b1 );
buf ( \1331_b0 , \1191_A[27]_b0 );
buf ( \1332_b1 , \1329_B[1]_b1 );
buf ( \1332_b0 , \1329_B[1]_b0 );
buf ( \1333_b1 , \1330_B[0]_b1 );
buf ( \1333_b0 , \1330_B[0]_b0 );
or ( \1334_b1 , \1332_b1 , \1333_b1 );
xor ( \1334_b0 , \1332_b0 , w_2392 );
not ( w_2392 , w_2393 );
and ( w_2393 , \1333_b1 , \1333_b0 );
buf ( \1335_b1 , \1333_b1 );
not ( \1335_b1 , w_2394 );
not ( \1335_b0 , w_2395 );
and ( w_2394 , w_2395 , \1333_b0 );
or ( \1336_b1 , \1334_b1 , \1335_b1 );
not ( \1335_b1 , w_2396 );
and ( \1336_b0 , \1334_b0 , w_2397 );
and ( w_2396 , w_2397 , \1335_b0 );
or ( \1337_b1 , \1331_b1 , \1336_b1 );
not ( \1336_b1 , w_2398 );
and ( \1337_b0 , \1331_b0 , w_2399 );
and ( w_2398 , w_2399 , \1336_b0 );
buf ( \1338_b1 , \1187_A[28]_b1 );
buf ( \1338_b0 , \1187_A[28]_b0 );
or ( \1339_b1 , \1338_b1 , \1333_b1 );
not ( \1333_b1 , w_2400 );
and ( \1339_b0 , \1338_b0 , w_2401 );
and ( w_2400 , w_2401 , \1333_b0 );
or ( \1340_b1 , \1337_b1 , w_2403 );
not ( w_2403 , w_2404 );
and ( \1340_b0 , \1337_b0 , w_2405 );
and ( w_2404 ,  , w_2405 );
buf ( w_2403 , \1339_b1 );
not ( w_2403 , w_2406 );
not (  , w_2407 );
and ( w_2406 , w_2407 , \1339_b0 );
or ( \1341_b1 , \1340_b1 , w_2408 );
xor ( \1341_b0 , \1340_b0 , w_2410 );
not ( w_2410 , w_2411 );
and ( w_2411 , w_2408 , w_2409 );
buf ( w_2408 , \1332_b1 );
not ( w_2408 , w_2412 );
not ( w_2409 , w_2413 );
and ( w_2412 , w_2413 , \1332_b0 );
buf ( \1342_b1 , \1215_A[21]_b1 );
buf ( \1342_b0 , \1215_A[21]_b0 );
buf ( \1343_b1 , \1323_B[7]_b1 );
buf ( \1343_b0 , \1323_B[7]_b0 );
buf ( \1344_b1 , \1324_B[6]_b1 );
buf ( \1344_b0 , \1324_B[6]_b0 );
or ( \1345_b1 , \1343_b1 , \1344_b1 );
xor ( \1345_b0 , \1343_b0 , w_2414 );
not ( w_2414 , w_2415 );
and ( w_2415 , \1344_b1 , \1344_b0 );
buf ( \1346_b1 , \1325_B[5]_b1 );
buf ( \1346_b0 , \1325_B[5]_b0 );
or ( \1347_b1 , \1344_b1 , \1346_b1 );
xor ( \1347_b0 , \1344_b0 , w_2416 );
not ( w_2416 , w_2417 );
and ( w_2417 , \1346_b1 , \1346_b0 );
buf ( \1348_b1 , \1347_b1 );
not ( \1348_b1 , w_2418 );
not ( \1348_b0 , w_2419 );
and ( w_2418 , w_2419 , \1347_b0 );
or ( \1349_b1 , \1345_b1 , \1348_b1 );
not ( \1348_b1 , w_2420 );
and ( \1349_b0 , \1345_b0 , w_2421 );
and ( w_2420 , w_2421 , \1348_b0 );
or ( \1350_b1 , \1342_b1 , \1349_b1 );
not ( \1349_b1 , w_2422 );
and ( \1350_b0 , \1342_b0 , w_2423 );
and ( w_2422 , w_2423 , \1349_b0 );
buf ( \1351_b1 , \1211_A[22]_b1 );
buf ( \1351_b0 , \1211_A[22]_b0 );
or ( \1352_b1 , \1351_b1 , \1347_b1 );
not ( \1347_b1 , w_2424 );
and ( \1352_b0 , \1351_b0 , w_2425 );
and ( w_2424 , w_2425 , \1347_b0 );
or ( \1353_b1 , \1350_b1 , w_2427 );
not ( w_2427 , w_2428 );
and ( \1353_b0 , \1350_b0 , w_2429 );
and ( w_2428 ,  , w_2429 );
buf ( w_2427 , \1352_b1 );
not ( w_2427 , w_2430 );
not (  , w_2431 );
and ( w_2430 , w_2431 , \1352_b0 );
or ( \1354_b1 , \1344_b1 , \1346_b1 );
not ( \1346_b1 , w_2432 );
and ( \1354_b0 , \1344_b0 , w_2433 );
and ( w_2432 , w_2433 , \1346_b0 );
buf ( \1355_b1 , \1354_b1 );
not ( \1355_b1 , w_2434 );
not ( \1355_b0 , w_2435 );
and ( w_2434 , w_2435 , \1354_b0 );
or ( \1356_b1 , \1343_b1 , \1355_b1 );
not ( \1355_b1 , w_2436 );
and ( \1356_b0 , \1343_b0 , w_2437 );
and ( w_2436 , w_2437 , \1355_b0 );
or ( \1357_b1 , \1353_b1 , w_2438 );
xor ( \1357_b0 , \1353_b0 , w_2440 );
not ( w_2440 , w_2441 );
and ( w_2441 , w_2438 , w_2439 );
buf ( w_2438 , \1356_b1 );
not ( w_2438 , w_2442 );
not ( w_2439 , w_2443 );
and ( w_2442 , w_2443 , \1356_b0 );
or ( \1358_b1 , \1341_b1 , \1357_b1 );
xor ( \1358_b0 , \1341_b0 , w_2444 );
not ( w_2444 , w_2445 );
and ( w_2445 , \1357_b1 , \1357_b0 );
buf ( \1359_b1 , \1247_A[13]_b1 );
buf ( \1359_b0 , \1247_A[13]_b0 );
buf ( \1360_b1 , \1315_B[15]_b1 );
buf ( \1360_b0 , \1315_B[15]_b0 );
buf ( \1361_b1 , \1316_B[14]_b1 );
buf ( \1361_b0 , \1316_B[14]_b0 );
or ( \1362_b1 , \1360_b1 , \1361_b1 );
xor ( \1362_b0 , \1360_b0 , w_2446 );
not ( w_2446 , w_2447 );
and ( w_2447 , \1361_b1 , \1361_b0 );
buf ( \1363_b1 , \1317_B[13]_b1 );
buf ( \1363_b0 , \1317_B[13]_b0 );
or ( \1364_b1 , \1361_b1 , \1363_b1 );
xor ( \1364_b0 , \1361_b0 , w_2448 );
not ( w_2448 , w_2449 );
and ( w_2449 , \1363_b1 , \1363_b0 );
buf ( \1365_b1 , \1364_b1 );
not ( \1365_b1 , w_2450 );
not ( \1365_b0 , w_2451 );
and ( w_2450 , w_2451 , \1364_b0 );
or ( \1366_b1 , \1362_b1 , \1365_b1 );
not ( \1365_b1 , w_2452 );
and ( \1366_b0 , \1362_b0 , w_2453 );
and ( w_2452 , w_2453 , \1365_b0 );
or ( \1367_b1 , \1359_b1 , \1366_b1 );
not ( \1366_b1 , w_2454 );
and ( \1367_b0 , \1359_b0 , w_2455 );
and ( w_2454 , w_2455 , \1366_b0 );
buf ( \1368_b1 , \1243_A[14]_b1 );
buf ( \1368_b0 , \1243_A[14]_b0 );
or ( \1369_b1 , \1368_b1 , \1364_b1 );
not ( \1364_b1 , w_2456 );
and ( \1369_b0 , \1368_b0 , w_2457 );
and ( w_2456 , w_2457 , \1364_b0 );
or ( \1370_b1 , \1367_b1 , w_2459 );
not ( w_2459 , w_2460 );
and ( \1370_b0 , \1367_b0 , w_2461 );
and ( w_2460 ,  , w_2461 );
buf ( w_2459 , \1369_b1 );
not ( w_2459 , w_2462 );
not (  , w_2463 );
and ( w_2462 , w_2463 , \1369_b0 );
or ( \1371_b1 , \1361_b1 , \1363_b1 );
not ( \1363_b1 , w_2464 );
and ( \1371_b0 , \1361_b0 , w_2465 );
and ( w_2464 , w_2465 , \1363_b0 );
buf ( \1372_b1 , \1371_b1 );
not ( \1372_b1 , w_2466 );
not ( \1372_b0 , w_2467 );
and ( w_2466 , w_2467 , \1371_b0 );
or ( \1373_b1 , \1360_b1 , \1372_b1 );
not ( \1372_b1 , w_2468 );
and ( \1373_b0 , \1360_b0 , w_2469 );
and ( w_2468 , w_2469 , \1372_b0 );
or ( \1374_b1 , \1370_b1 , w_2470 );
xor ( \1374_b0 , \1370_b0 , w_2472 );
not ( w_2472 , w_2473 );
and ( w_2473 , w_2470 , w_2471 );
buf ( w_2470 , \1373_b1 );
not ( w_2470 , w_2474 );
not ( w_2471 , w_2475 );
and ( w_2474 , w_2475 , \1373_b0 );
or ( \1375_b1 , \1358_b1 , \1374_b1 );
xor ( \1375_b0 , \1358_b0 , w_2476 );
not ( w_2476 , w_2477 );
and ( w_2477 , \1374_b1 , \1374_b0 );
buf ( \1376_b1 , \1223_A[19]_b1 );
buf ( \1376_b0 , \1223_A[19]_b0 );
buf ( \1377_b1 , \1321_B[9]_b1 );
buf ( \1377_b0 , \1321_B[9]_b0 );
buf ( \1378_b1 , \1322_B[8]_b1 );
buf ( \1378_b0 , \1322_B[8]_b0 );
or ( \1379_b1 , \1377_b1 , \1378_b1 );
xor ( \1379_b0 , \1377_b0 , w_2478 );
not ( w_2478 , w_2479 );
and ( w_2479 , \1378_b1 , \1378_b0 );
or ( \1380_b1 , \1378_b1 , \1343_b1 );
xor ( \1380_b0 , \1378_b0 , w_2480 );
not ( w_2480 , w_2481 );
and ( w_2481 , \1343_b1 , \1343_b0 );
buf ( \1381_b1 , \1380_b1 );
not ( \1381_b1 , w_2482 );
not ( \1381_b0 , w_2483 );
and ( w_2482 , w_2483 , \1380_b0 );
or ( \1382_b1 , \1379_b1 , \1381_b1 );
not ( \1381_b1 , w_2484 );
and ( \1382_b0 , \1379_b0 , w_2485 );
and ( w_2484 , w_2485 , \1381_b0 );
or ( \1383_b1 , \1376_b1 , \1382_b1 );
not ( \1382_b1 , w_2486 );
and ( \1383_b0 , \1376_b0 , w_2487 );
and ( w_2486 , w_2487 , \1382_b0 );
buf ( \1384_b1 , \1219_A[20]_b1 );
buf ( \1384_b0 , \1219_A[20]_b0 );
or ( \1385_b1 , \1384_b1 , \1380_b1 );
not ( \1380_b1 , w_2488 );
and ( \1385_b0 , \1384_b0 , w_2489 );
and ( w_2488 , w_2489 , \1380_b0 );
or ( \1386_b1 , \1383_b1 , w_2491 );
not ( w_2491 , w_2492 );
and ( \1386_b0 , \1383_b0 , w_2493 );
and ( w_2492 ,  , w_2493 );
buf ( w_2491 , \1385_b1 );
not ( w_2491 , w_2494 );
not (  , w_2495 );
and ( w_2494 , w_2495 , \1385_b0 );
or ( \1387_b1 , \1378_b1 , \1343_b1 );
not ( \1343_b1 , w_2496 );
and ( \1387_b0 , \1378_b0 , w_2497 );
and ( w_2496 , w_2497 , \1343_b0 );
buf ( \1388_b1 , \1387_b1 );
not ( \1388_b1 , w_2498 );
not ( \1388_b0 , w_2499 );
and ( w_2498 , w_2499 , \1387_b0 );
or ( \1389_b1 , \1377_b1 , \1388_b1 );
not ( \1388_b1 , w_2500 );
and ( \1389_b0 , \1377_b0 , w_2501 );
and ( w_2500 , w_2501 , \1388_b0 );
or ( \1390_b1 , \1386_b1 , w_2502 );
xor ( \1390_b0 , \1386_b0 , w_2504 );
not ( w_2504 , w_2505 );
and ( w_2505 , w_2502 , w_2503 );
buf ( w_2502 , \1389_b1 );
not ( w_2502 , w_2506 );
not ( w_2503 , w_2507 );
and ( w_2506 , w_2507 , \1389_b0 );
buf ( \1391_b1 , \1255_A[11]_b1 );
buf ( \1391_b0 , \1255_A[11]_b0 );
buf ( \1392_b1 , \1313_B[17]_b1 );
buf ( \1392_b0 , \1313_B[17]_b0 );
buf ( \1393_b1 , \1314_B[16]_b1 );
buf ( \1393_b0 , \1314_B[16]_b0 );
or ( \1394_b1 , \1392_b1 , \1393_b1 );
xor ( \1394_b0 , \1392_b0 , w_2508 );
not ( w_2508 , w_2509 );
and ( w_2509 , \1393_b1 , \1393_b0 );
or ( \1395_b1 , \1393_b1 , \1360_b1 );
xor ( \1395_b0 , \1393_b0 , w_2510 );
not ( w_2510 , w_2511 );
and ( w_2511 , \1360_b1 , \1360_b0 );
buf ( \1396_b1 , \1395_b1 );
not ( \1396_b1 , w_2512 );
not ( \1396_b0 , w_2513 );
and ( w_2512 , w_2513 , \1395_b0 );
or ( \1397_b1 , \1394_b1 , \1396_b1 );
not ( \1396_b1 , w_2514 );
and ( \1397_b0 , \1394_b0 , w_2515 );
and ( w_2514 , w_2515 , \1396_b0 );
or ( \1398_b1 , \1391_b1 , \1397_b1 );
not ( \1397_b1 , w_2516 );
and ( \1398_b0 , \1391_b0 , w_2517 );
and ( w_2516 , w_2517 , \1397_b0 );
buf ( \1399_b1 , \1251_A[12]_b1 );
buf ( \1399_b0 , \1251_A[12]_b0 );
or ( \1400_b1 , \1399_b1 , \1395_b1 );
not ( \1395_b1 , w_2518 );
and ( \1400_b0 , \1399_b0 , w_2519 );
and ( w_2518 , w_2519 , \1395_b0 );
or ( \1401_b1 , \1398_b1 , w_2521 );
not ( w_2521 , w_2522 );
and ( \1401_b0 , \1398_b0 , w_2523 );
and ( w_2522 ,  , w_2523 );
buf ( w_2521 , \1400_b1 );
not ( w_2521 , w_2524 );
not (  , w_2525 );
and ( w_2524 , w_2525 , \1400_b0 );
or ( \1402_b1 , \1393_b1 , \1360_b1 );
not ( \1360_b1 , w_2526 );
and ( \1402_b0 , \1393_b0 , w_2527 );
and ( w_2526 , w_2527 , \1360_b0 );
buf ( \1403_b1 , \1402_b1 );
not ( \1403_b1 , w_2528 );
not ( \1403_b0 , w_2529 );
and ( w_2528 , w_2529 , \1402_b0 );
or ( \1404_b1 , \1392_b1 , \1403_b1 );
not ( \1403_b1 , w_2530 );
and ( \1404_b0 , \1392_b0 , w_2531 );
and ( w_2530 , w_2531 , \1403_b0 );
or ( \1405_b1 , \1401_b1 , w_2532 );
xor ( \1405_b0 , \1401_b0 , w_2534 );
not ( w_2534 , w_2535 );
and ( w_2535 , w_2532 , w_2533 );
buf ( w_2532 , \1404_b1 );
not ( w_2532 , w_2536 );
not ( w_2533 , w_2537 );
and ( w_2536 , w_2537 , \1404_b0 );
or ( \1406_b1 , \1390_b1 , \1405_b1 );
xor ( \1406_b0 , \1390_b0 , w_2538 );
not ( w_2538 , w_2539 );
and ( w_2539 , \1405_b1 , \1405_b0 );
buf ( \1407_b1 , \1271_A[7]_b1 );
buf ( \1407_b0 , \1271_A[7]_b0 );
buf ( \1408_b1 , \1309_B[21]_b1 );
buf ( \1408_b0 , \1309_B[21]_b0 );
buf ( \1409_b1 , \1310_B[20]_b1 );
buf ( \1409_b0 , \1310_B[20]_b0 );
or ( \1410_b1 , \1408_b1 , \1409_b1 );
xor ( \1410_b0 , \1408_b0 , w_2540 );
not ( w_2540 , w_2541 );
and ( w_2541 , \1409_b1 , \1409_b0 );
buf ( \1411_b1 , \1311_B[19]_b1 );
buf ( \1411_b0 , \1311_B[19]_b0 );
or ( \1412_b1 , \1409_b1 , \1411_b1 );
xor ( \1412_b0 , \1409_b0 , w_2542 );
not ( w_2542 , w_2543 );
and ( w_2543 , \1411_b1 , \1411_b0 );
buf ( \1413_b1 , \1412_b1 );
not ( \1413_b1 , w_2544 );
not ( \1413_b0 , w_2545 );
and ( w_2544 , w_2545 , \1412_b0 );
or ( \1414_b1 , \1410_b1 , \1413_b1 );
not ( \1413_b1 , w_2546 );
and ( \1414_b0 , \1410_b0 , w_2547 );
and ( w_2546 , w_2547 , \1413_b0 );
or ( \1415_b1 , \1407_b1 , \1414_b1 );
not ( \1414_b1 , w_2548 );
and ( \1415_b0 , \1407_b0 , w_2549 );
and ( w_2548 , w_2549 , \1414_b0 );
buf ( \1416_b1 , \1267_A[8]_b1 );
buf ( \1416_b0 , \1267_A[8]_b0 );
or ( \1417_b1 , \1416_b1 , \1412_b1 );
not ( \1412_b1 , w_2550 );
and ( \1417_b0 , \1416_b0 , w_2551 );
and ( w_2550 , w_2551 , \1412_b0 );
or ( \1418_b1 , \1415_b1 , w_2553 );
not ( w_2553 , w_2554 );
and ( \1418_b0 , \1415_b0 , w_2555 );
and ( w_2554 ,  , w_2555 );
buf ( w_2553 , \1417_b1 );
not ( w_2553 , w_2556 );
not (  , w_2557 );
and ( w_2556 , w_2557 , \1417_b0 );
or ( \1419_b1 , \1409_b1 , \1411_b1 );
not ( \1411_b1 , w_2558 );
and ( \1419_b0 , \1409_b0 , w_2559 );
and ( w_2558 , w_2559 , \1411_b0 );
buf ( \1420_b1 , \1419_b1 );
not ( \1420_b1 , w_2560 );
not ( \1420_b0 , w_2561 );
and ( w_2560 , w_2561 , \1419_b0 );
or ( \1421_b1 , \1408_b1 , \1420_b1 );
not ( \1420_b1 , w_2562 );
and ( \1421_b0 , \1408_b0 , w_2563 );
and ( w_2562 , w_2563 , \1420_b0 );
or ( \1422_b1 , \1418_b1 , w_2564 );
xor ( \1422_b0 , \1418_b0 , w_2566 );
not ( w_2566 , w_2567 );
and ( w_2567 , w_2564 , w_2565 );
buf ( w_2564 , \1421_b1 );
not ( w_2564 , w_2568 );
not ( w_2565 , w_2569 );
and ( w_2568 , w_2569 , \1421_b0 );
or ( \1423_b1 , \1406_b1 , \1422_b1 );
xor ( \1423_b0 , \1406_b0 , w_2570 );
not ( w_2570 , w_2571 );
and ( w_2571 , \1422_b1 , \1422_b0 );
or ( \1424_b1 , \1375_b1 , \1423_b1 );
not ( \1423_b1 , w_2572 );
and ( \1424_b0 , \1375_b0 , w_2573 );
and ( w_2572 , w_2573 , \1423_b0 );
buf ( \1425_b1 , \1203_A[24]_b1 );
buf ( \1425_b0 , \1203_A[24]_b0 );
buf ( \1426_b1 , \1327_B[3]_b1 );
buf ( \1426_b0 , \1327_B[3]_b0 );
buf ( \1427_b1 , \1328_B[2]_b1 );
buf ( \1427_b0 , \1328_B[2]_b0 );
or ( \1428_b1 , \1426_b1 , \1427_b1 );
xor ( \1428_b0 , \1426_b0 , w_2574 );
not ( w_2574 , w_2575 );
and ( w_2575 , \1427_b1 , \1427_b0 );
or ( \1429_b1 , \1427_b1 , \1332_b1 );
xor ( \1429_b0 , \1427_b0 , w_2576 );
not ( w_2576 , w_2577 );
and ( w_2577 , \1332_b1 , \1332_b0 );
buf ( \1430_b1 , \1429_b1 );
not ( \1430_b1 , w_2578 );
not ( \1430_b0 , w_2579 );
and ( w_2578 , w_2579 , \1429_b0 );
or ( \1431_b1 , \1428_b1 , \1430_b1 );
not ( \1430_b1 , w_2580 );
and ( \1431_b0 , \1428_b0 , w_2581 );
and ( w_2580 , w_2581 , \1430_b0 );
or ( \1432_b1 , \1425_b1 , \1431_b1 );
not ( \1431_b1 , w_2582 );
and ( \1432_b0 , \1425_b0 , w_2583 );
and ( w_2582 , w_2583 , \1431_b0 );
buf ( \1433_b1 , \1199_A[25]_b1 );
buf ( \1433_b0 , \1199_A[25]_b0 );
or ( \1434_b1 , \1433_b1 , \1429_b1 );
not ( \1429_b1 , w_2584 );
and ( \1434_b0 , \1433_b0 , w_2585 );
and ( w_2584 , w_2585 , \1429_b0 );
or ( \1435_b1 , \1432_b1 , w_2587 );
not ( w_2587 , w_2588 );
and ( \1435_b0 , \1432_b0 , w_2589 );
and ( w_2588 ,  , w_2589 );
buf ( w_2587 , \1434_b1 );
not ( w_2587 , w_2590 );
not (  , w_2591 );
and ( w_2590 , w_2591 , \1434_b0 );
or ( \1436_b1 , \1427_b1 , \1332_b1 );
not ( \1332_b1 , w_2592 );
and ( \1436_b0 , \1427_b0 , w_2593 );
and ( w_2592 , w_2593 , \1332_b0 );
buf ( \1437_b1 , \1436_b1 );
not ( \1437_b1 , w_2594 );
not ( \1437_b0 , w_2595 );
and ( w_2594 , w_2595 , \1436_b0 );
or ( \1438_b1 , \1426_b1 , \1437_b1 );
not ( \1437_b1 , w_2596 );
and ( \1438_b0 , \1426_b0 , w_2597 );
and ( w_2596 , w_2597 , \1437_b0 );
or ( \1439_b1 , \1435_b1 , w_2598 );
xor ( \1439_b0 , \1435_b0 , w_2600 );
not ( w_2600 , w_2601 );
and ( w_2601 , w_2598 , w_2599 );
buf ( w_2598 , \1438_b1 );
not ( w_2598 , w_2602 );
not ( w_2599 , w_2603 );
and ( w_2602 , w_2603 , \1438_b0 );
buf ( \1440_b1 , \1326_B[4]_b1 );
buf ( \1440_b0 , \1326_B[4]_b0 );
or ( \1441_b1 , \1346_b1 , \1440_b1 );
xor ( \1441_b0 , \1346_b0 , w_2604 );
not ( w_2604 , w_2605 );
and ( w_2605 , \1440_b1 , \1440_b0 );
or ( \1442_b1 , \1440_b1 , \1426_b1 );
xor ( \1442_b0 , \1440_b0 , w_2606 );
not ( w_2606 , w_2607 );
and ( w_2607 , \1426_b1 , \1426_b0 );
buf ( \1443_b1 , \1442_b1 );
not ( \1443_b1 , w_2608 );
not ( \1443_b0 , w_2609 );
and ( w_2608 , w_2609 , \1442_b0 );
or ( \1444_b1 , \1441_b1 , \1443_b1 );
not ( \1443_b1 , w_2610 );
and ( \1444_b0 , \1441_b0 , w_2611 );
and ( w_2610 , w_2611 , \1443_b0 );
or ( \1445_b1 , \1351_b1 , \1444_b1 );
not ( \1444_b1 , w_2612 );
and ( \1445_b0 , \1351_b0 , w_2613 );
and ( w_2612 , w_2613 , \1444_b0 );
buf ( \1446_b1 , \1207_A[23]_b1 );
buf ( \1446_b0 , \1207_A[23]_b0 );
or ( \1447_b1 , \1446_b1 , \1442_b1 );
not ( \1442_b1 , w_2614 );
and ( \1447_b0 , \1446_b0 , w_2615 );
and ( w_2614 , w_2615 , \1442_b0 );
or ( \1448_b1 , \1445_b1 , w_2617 );
not ( w_2617 , w_2618 );
and ( \1448_b0 , \1445_b0 , w_2619 );
and ( w_2618 ,  , w_2619 );
buf ( w_2617 , \1447_b1 );
not ( w_2617 , w_2620 );
not (  , w_2621 );
and ( w_2620 , w_2621 , \1447_b0 );
or ( \1449_b1 , \1440_b1 , \1426_b1 );
not ( \1426_b1 , w_2622 );
and ( \1449_b0 , \1440_b0 , w_2623 );
and ( w_2622 , w_2623 , \1426_b0 );
buf ( \1450_b1 , \1449_b1 );
not ( \1450_b1 , w_2624 );
not ( \1450_b0 , w_2625 );
and ( w_2624 , w_2625 , \1449_b0 );
or ( \1451_b1 , \1346_b1 , \1450_b1 );
not ( \1450_b1 , w_2626 );
and ( \1451_b0 , \1346_b0 , w_2627 );
and ( w_2626 , w_2627 , \1450_b0 );
or ( \1452_b1 , \1448_b1 , w_2628 );
xor ( \1452_b0 , \1448_b0 , w_2630 );
not ( w_2630 , w_2631 );
and ( w_2631 , w_2628 , w_2629 );
buf ( w_2628 , \1451_b1 );
not ( w_2628 , w_2632 );
not ( w_2629 , w_2633 );
and ( w_2632 , w_2633 , \1451_b0 );
or ( \1453_b1 , \1439_b1 , \1452_b1 );
not ( \1452_b1 , w_2634 );
and ( \1453_b0 , \1439_b0 , w_2635 );
and ( w_2634 , w_2635 , \1452_b0 );
buf ( \1454_b1 , \1231_A[17]_b1 );
buf ( \1454_b0 , \1231_A[17]_b0 );
buf ( \1455_b1 , \1319_B[11]_b1 );
buf ( \1455_b0 , \1319_B[11]_b0 );
buf ( \1456_b1 , \1320_B[10]_b1 );
buf ( \1456_b0 , \1320_B[10]_b0 );
or ( \1457_b1 , \1455_b1 , \1456_b1 );
xor ( \1457_b0 , \1455_b0 , w_2636 );
not ( w_2636 , w_2637 );
and ( w_2637 , \1456_b1 , \1456_b0 );
or ( \1458_b1 , \1456_b1 , \1377_b1 );
xor ( \1458_b0 , \1456_b0 , w_2638 );
not ( w_2638 , w_2639 );
and ( w_2639 , \1377_b1 , \1377_b0 );
buf ( \1459_b1 , \1458_b1 );
not ( \1459_b1 , w_2640 );
not ( \1459_b0 , w_2641 );
and ( w_2640 , w_2641 , \1458_b0 );
or ( \1460_b1 , \1457_b1 , \1459_b1 );
not ( \1459_b1 , w_2642 );
and ( \1460_b0 , \1457_b0 , w_2643 );
and ( w_2642 , w_2643 , \1459_b0 );
or ( \1461_b1 , \1454_b1 , \1460_b1 );
not ( \1460_b1 , w_2644 );
and ( \1461_b0 , \1454_b0 , w_2645 );
and ( w_2644 , w_2645 , \1460_b0 );
buf ( \1462_b1 , \1227_A[18]_b1 );
buf ( \1462_b0 , \1227_A[18]_b0 );
or ( \1463_b1 , \1462_b1 , \1458_b1 );
not ( \1458_b1 , w_2646 );
and ( \1463_b0 , \1462_b0 , w_2647 );
and ( w_2646 , w_2647 , \1458_b0 );
or ( \1464_b1 , \1461_b1 , w_2649 );
not ( w_2649 , w_2650 );
and ( \1464_b0 , \1461_b0 , w_2651 );
and ( w_2650 ,  , w_2651 );
buf ( w_2649 , \1463_b1 );
not ( w_2649 , w_2652 );
not (  , w_2653 );
and ( w_2652 , w_2653 , \1463_b0 );
or ( \1465_b1 , \1456_b1 , \1377_b1 );
not ( \1377_b1 , w_2654 );
and ( \1465_b0 , \1456_b0 , w_2655 );
and ( w_2654 , w_2655 , \1377_b0 );
buf ( \1466_b1 , \1465_b1 );
not ( \1466_b1 , w_2656 );
not ( \1466_b0 , w_2657 );
and ( w_2656 , w_2657 , \1465_b0 );
or ( \1467_b1 , \1455_b1 , \1466_b1 );
not ( \1466_b1 , w_2658 );
and ( \1467_b0 , \1455_b0 , w_2659 );
and ( w_2658 , w_2659 , \1466_b0 );
or ( \1468_b1 , \1464_b1 , w_2660 );
xor ( \1468_b0 , \1464_b0 , w_2662 );
not ( w_2662 , w_2663 );
and ( w_2663 , w_2660 , w_2661 );
buf ( w_2660 , \1467_b1 );
not ( w_2660 , w_2664 );
not ( w_2661 , w_2665 );
and ( w_2664 , w_2665 , \1467_b0 );
or ( \1469_b1 , \1453_b1 , \1468_b1 );
xor ( \1469_b0 , \1453_b0 , w_2666 );
not ( w_2666 , w_2667 );
and ( w_2667 , \1468_b1 , \1468_b0 );
buf ( \1470_b1 , \1239_A[15]_b1 );
buf ( \1470_b0 , \1239_A[15]_b0 );
buf ( \1471_b1 , \1318_B[12]_b1 );
buf ( \1471_b0 , \1318_B[12]_b0 );
or ( \1472_b1 , \1363_b1 , \1471_b1 );
xor ( \1472_b0 , \1363_b0 , w_2668 );
not ( w_2668 , w_2669 );
and ( w_2669 , \1471_b1 , \1471_b0 );
or ( \1473_b1 , \1471_b1 , \1455_b1 );
xor ( \1473_b0 , \1471_b0 , w_2670 );
not ( w_2670 , w_2671 );
and ( w_2671 , \1455_b1 , \1455_b0 );
buf ( \1474_b1 , \1473_b1 );
not ( \1474_b1 , w_2672 );
not ( \1474_b0 , w_2673 );
and ( w_2672 , w_2673 , \1473_b0 );
or ( \1475_b1 , \1472_b1 , \1474_b1 );
not ( \1474_b1 , w_2674 );
and ( \1475_b0 , \1472_b0 , w_2675 );
and ( w_2674 , w_2675 , \1474_b0 );
or ( \1476_b1 , \1470_b1 , \1475_b1 );
not ( \1475_b1 , w_2676 );
and ( \1476_b0 , \1470_b0 , w_2677 );
and ( w_2676 , w_2677 , \1475_b0 );
buf ( \1477_b1 , \1235_A[16]_b1 );
buf ( \1477_b0 , \1235_A[16]_b0 );
or ( \1478_b1 , \1477_b1 , \1473_b1 );
not ( \1473_b1 , w_2678 );
and ( \1478_b0 , \1477_b0 , w_2679 );
and ( w_2678 , w_2679 , \1473_b0 );
or ( \1479_b1 , \1476_b1 , w_2681 );
not ( w_2681 , w_2682 );
and ( \1479_b0 , \1476_b0 , w_2683 );
and ( w_2682 ,  , w_2683 );
buf ( w_2681 , \1478_b1 );
not ( w_2681 , w_2684 );
not (  , w_2685 );
and ( w_2684 , w_2685 , \1478_b0 );
or ( \1480_b1 , \1471_b1 , \1455_b1 );
not ( \1455_b1 , w_2686 );
and ( \1480_b0 , \1471_b0 , w_2687 );
and ( w_2686 , w_2687 , \1455_b0 );
buf ( \1481_b1 , \1480_b1 );
not ( \1481_b1 , w_2688 );
not ( \1481_b0 , w_2689 );
and ( w_2688 , w_2689 , \1480_b0 );
or ( \1482_b1 , \1363_b1 , \1481_b1 );
not ( \1481_b1 , w_2690 );
and ( \1482_b0 , \1363_b0 , w_2691 );
and ( w_2690 , w_2691 , \1481_b0 );
or ( \1483_b1 , \1479_b1 , w_2692 );
xor ( \1483_b0 , \1479_b0 , w_2694 );
not ( w_2694 , w_2695 );
and ( w_2695 , w_2692 , w_2693 );
buf ( w_2692 , \1482_b1 );
not ( w_2692 , w_2696 );
not ( w_2693 , w_2697 );
and ( w_2696 , w_2697 , \1482_b0 );
or ( \1484_b1 , \1469_b1 , \1483_b1 );
xor ( \1484_b0 , \1469_b0 , w_2698 );
not ( w_2698 , w_2699 );
and ( w_2699 , \1483_b1 , \1483_b0 );
or ( \1485_b1 , \1423_b1 , \1484_b1 );
not ( \1484_b1 , w_2700 );
and ( \1485_b0 , \1423_b0 , w_2701 );
and ( w_2700 , w_2701 , \1484_b0 );
or ( \1486_b1 , \1375_b1 , \1484_b1 );
not ( \1484_b1 , w_2702 );
and ( \1486_b0 , \1375_b0 , w_2703 );
and ( w_2702 , w_2703 , \1484_b0 );
or ( \1488_b1 , \1433_b1 , \1431_b1 );
not ( \1431_b1 , w_2704 );
and ( \1488_b0 , \1433_b0 , w_2705 );
and ( w_2704 , w_2705 , \1431_b0 );
buf ( \1489_b1 , \1195_A[26]_b1 );
buf ( \1489_b0 , \1195_A[26]_b0 );
or ( \1490_b1 , \1489_b1 , \1429_b1 );
not ( \1429_b1 , w_2706 );
and ( \1490_b0 , \1489_b0 , w_2707 );
and ( w_2706 , w_2707 , \1429_b0 );
or ( \1491_b1 , \1488_b1 , w_2709 );
not ( w_2709 , w_2710 );
and ( \1491_b0 , \1488_b0 , w_2711 );
and ( w_2710 ,  , w_2711 );
buf ( w_2709 , \1490_b1 );
not ( w_2709 , w_2712 );
not (  , w_2713 );
and ( w_2712 , w_2713 , \1490_b0 );
or ( \1492_b1 , \1491_b1 , w_2714 );
xor ( \1492_b0 , \1491_b0 , w_2716 );
not ( w_2716 , w_2717 );
and ( w_2717 , w_2714 , w_2715 );
buf ( w_2714 , \1438_b1 );
not ( w_2714 , w_2718 );
not ( w_2715 , w_2719 );
and ( w_2718 , w_2719 , \1438_b0 );
or ( \1493_b1 , \1446_b1 , \1444_b1 );
not ( \1444_b1 , w_2720 );
and ( \1493_b0 , \1446_b0 , w_2721 );
and ( w_2720 , w_2721 , \1444_b0 );
or ( \1494_b1 , \1425_b1 , \1442_b1 );
not ( \1442_b1 , w_2722 );
and ( \1494_b0 , \1425_b0 , w_2723 );
and ( w_2722 , w_2723 , \1442_b0 );
or ( \1495_b1 , \1493_b1 , w_2725 );
not ( w_2725 , w_2726 );
and ( \1495_b0 , \1493_b0 , w_2727 );
and ( w_2726 ,  , w_2727 );
buf ( w_2725 , \1494_b1 );
not ( w_2725 , w_2728 );
not (  , w_2729 );
and ( w_2728 , w_2729 , \1494_b0 );
or ( \1496_b1 , \1495_b1 , w_2730 );
xor ( \1496_b0 , \1495_b0 , w_2732 );
not ( w_2732 , w_2733 );
and ( w_2733 , w_2730 , w_2731 );
buf ( w_2730 , \1451_b1 );
not ( w_2730 , w_2734 );
not ( w_2731 , w_2735 );
and ( w_2734 , w_2735 , \1451_b0 );
or ( \1497_b1 , \1492_b1 , \1496_b1 );
not ( \1496_b1 , w_2736 );
and ( \1497_b0 , \1492_b0 , w_2737 );
and ( w_2736 , w_2737 , \1496_b0 );
buf ( \1498_b1 , \1298_A[0]_b1 );
buf ( \1498_b0 , \1298_A[0]_b0 );
buf ( \1499_b1 , \1302_B[28]_b1 );
buf ( \1499_b0 , \1302_B[28]_b0 );
buf ( \1500_b1 , \1303_B[27]_b1 );
buf ( \1500_b0 , \1303_B[27]_b0 );
or ( \1501_b1 , \1499_b1 , \1500_b1 );
xor ( \1501_b0 , \1499_b0 , w_2738 );
not ( w_2738 , w_2739 );
and ( w_2739 , \1500_b1 , \1500_b0 );
or ( \1502_b1 , \1498_b1 , \1501_b1 );
not ( \1501_b1 , w_2740 );
and ( \1502_b0 , \1498_b0 , w_2741 );
and ( w_2740 , w_2741 , \1501_b0 );
or ( \1503_b1 , \1496_b1 , \1502_b1 );
not ( \1502_b1 , w_2742 );
and ( \1503_b0 , \1496_b0 , w_2743 );
and ( w_2742 , w_2743 , \1502_b0 );
or ( \1504_b1 , \1492_b1 , \1502_b1 );
not ( \1502_b1 , w_2744 );
and ( \1504_b0 , \1492_b0 , w_2745 );
and ( w_2744 , w_2745 , \1502_b0 );
or ( \1506_b1 , \1341_b1 , \1357_b1 );
not ( \1357_b1 , w_2746 );
and ( \1506_b0 , \1341_b0 , w_2747 );
and ( w_2746 , w_2747 , \1357_b0 );
or ( \1507_b1 , \1357_b1 , \1374_b1 );
not ( \1374_b1 , w_2748 );
and ( \1507_b0 , \1357_b0 , w_2749 );
and ( w_2748 , w_2749 , \1374_b0 );
or ( \1508_b1 , \1341_b1 , \1374_b1 );
not ( \1374_b1 , w_2750 );
and ( \1508_b0 , \1341_b0 , w_2751 );
and ( w_2750 , w_2751 , \1374_b0 );
or ( \1510_b1 , \1505_b1 , \1509_b1 );
xor ( \1510_b0 , \1505_b0 , w_2752 );
not ( w_2752 , w_2753 );
and ( w_2753 , \1509_b1 , \1509_b0 );
or ( \1511_b1 , \1390_b1 , \1405_b1 );
not ( \1405_b1 , w_2754 );
and ( \1511_b0 , \1390_b0 , w_2755 );
and ( w_2754 , w_2755 , \1405_b0 );
or ( \1512_b1 , \1405_b1 , \1422_b1 );
not ( \1422_b1 , w_2756 );
and ( \1512_b0 , \1405_b0 , w_2757 );
and ( w_2756 , w_2757 , \1422_b0 );
or ( \1513_b1 , \1390_b1 , \1422_b1 );
not ( \1422_b1 , w_2758 );
and ( \1513_b0 , \1390_b0 , w_2759 );
and ( w_2758 , w_2759 , \1422_b0 );
or ( \1515_b1 , \1510_b1 , \1514_b1 );
xor ( \1515_b0 , \1510_b0 , w_2760 );
not ( w_2760 , w_2761 );
and ( w_2761 , \1514_b1 , \1514_b0 );
or ( \1516_b1 , \1487_b1 , \1515_b1 );
not ( \1515_b1 , w_2762 );
and ( \1516_b0 , \1487_b0 , w_2763 );
and ( w_2762 , w_2763 , \1515_b0 );
buf ( \1517_b1 , \1283_A[4]_b1 );
buf ( \1517_b0 , \1283_A[4]_b0 );
buf ( \1518_b1 , \1305_B[25]_b1 );
buf ( \1518_b0 , \1305_B[25]_b0 );
buf ( \1519_b1 , \1306_B[24]_b1 );
buf ( \1519_b0 , \1306_B[24]_b0 );
or ( \1520_b1 , \1518_b1 , \1519_b1 );
xor ( \1520_b0 , \1518_b0 , w_2764 );
not ( w_2764 , w_2765 );
and ( w_2765 , \1519_b1 , \1519_b0 );
buf ( \1521_b1 , \1307_B[23]_b1 );
buf ( \1521_b0 , \1307_B[23]_b0 );
or ( \1522_b1 , \1519_b1 , \1521_b1 );
xor ( \1522_b0 , \1519_b0 , w_2766 );
not ( w_2766 , w_2767 );
and ( w_2767 , \1521_b1 , \1521_b0 );
buf ( \1523_b1 , \1522_b1 );
not ( \1523_b1 , w_2768 );
not ( \1523_b0 , w_2769 );
and ( w_2768 , w_2769 , \1522_b0 );
or ( \1524_b1 , \1520_b1 , \1523_b1 );
not ( \1523_b1 , w_2770 );
and ( \1524_b0 , \1520_b0 , w_2771 );
and ( w_2770 , w_2771 , \1523_b0 );
or ( \1525_b1 , \1517_b1 , \1524_b1 );
not ( \1524_b1 , w_2772 );
and ( \1525_b0 , \1517_b0 , w_2773 );
and ( w_2772 , w_2773 , \1524_b0 );
buf ( \1526_b1 , \1279_A[5]_b1 );
buf ( \1526_b0 , \1279_A[5]_b0 );
or ( \1527_b1 , \1526_b1 , \1522_b1 );
not ( \1522_b1 , w_2774 );
and ( \1527_b0 , \1526_b0 , w_2775 );
and ( w_2774 , w_2775 , \1522_b0 );
or ( \1528_b1 , \1525_b1 , w_2777 );
not ( w_2777 , w_2778 );
and ( \1528_b0 , \1525_b0 , w_2779 );
and ( w_2778 ,  , w_2779 );
buf ( w_2777 , \1527_b1 );
not ( w_2777 , w_2780 );
not (  , w_2781 );
and ( w_2780 , w_2781 , \1527_b0 );
or ( \1529_b1 , \1519_b1 , \1521_b1 );
not ( \1521_b1 , w_2782 );
and ( \1529_b0 , \1519_b0 , w_2783 );
and ( w_2782 , w_2783 , \1521_b0 );
buf ( \1530_b1 , \1529_b1 );
not ( \1530_b1 , w_2784 );
not ( \1530_b0 , w_2785 );
and ( w_2784 , w_2785 , \1529_b0 );
or ( \1531_b1 , \1518_b1 , \1530_b1 );
not ( \1530_b1 , w_2786 );
and ( \1531_b0 , \1518_b0 , w_2787 );
and ( w_2786 , w_2787 , \1530_b0 );
or ( \1532_b1 , \1528_b1 , w_2788 );
xor ( \1532_b0 , \1528_b0 , w_2790 );
not ( w_2790 , w_2791 );
and ( w_2791 , w_2788 , w_2789 );
buf ( w_2788 , \1531_b1 );
not ( w_2788 , w_2792 );
not ( w_2789 , w_2793 );
and ( w_2792 , w_2793 , \1531_b0 );
buf ( \1533_b1 , \1291_A[2]_b1 );
buf ( \1533_b0 , \1291_A[2]_b0 );
buf ( \1534_b1 , \1304_B[26]_b1 );
buf ( \1534_b0 , \1304_B[26]_b0 );
or ( \1535_b1 , \1500_b1 , \1534_b1 );
xor ( \1535_b0 , \1500_b0 , w_2794 );
not ( w_2794 , w_2795 );
and ( w_2795 , \1534_b1 , \1534_b0 );
or ( \1536_b1 , \1534_b1 , \1518_b1 );
xor ( \1536_b0 , \1534_b0 , w_2796 );
not ( w_2796 , w_2797 );
and ( w_2797 , \1518_b1 , \1518_b0 );
buf ( \1537_b1 , \1536_b1 );
not ( \1537_b1 , w_2798 );
not ( \1537_b0 , w_2799 );
and ( w_2798 , w_2799 , \1536_b0 );
or ( \1538_b1 , \1535_b1 , \1537_b1 );
not ( \1537_b1 , w_2800 );
and ( \1538_b0 , \1535_b0 , w_2801 );
and ( w_2800 , w_2801 , \1537_b0 );
or ( \1539_b1 , \1533_b1 , \1538_b1 );
not ( \1538_b1 , w_2802 );
and ( \1539_b0 , \1533_b0 , w_2803 );
and ( w_2802 , w_2803 , \1538_b0 );
buf ( \1540_b1 , \1287_A[3]_b1 );
buf ( \1540_b0 , \1287_A[3]_b0 );
or ( \1541_b1 , \1540_b1 , \1536_b1 );
not ( \1536_b1 , w_2804 );
and ( \1541_b0 , \1540_b0 , w_2805 );
and ( w_2804 , w_2805 , \1536_b0 );
or ( \1542_b1 , \1539_b1 , w_2807 );
not ( w_2807 , w_2808 );
and ( \1542_b0 , \1539_b0 , w_2809 );
and ( w_2808 ,  , w_2809 );
buf ( w_2807 , \1541_b1 );
not ( w_2807 , w_2810 );
not (  , w_2811 );
and ( w_2810 , w_2811 , \1541_b0 );
or ( \1543_b1 , \1534_b1 , \1518_b1 );
not ( \1518_b1 , w_2812 );
and ( \1543_b0 , \1534_b0 , w_2813 );
and ( w_2812 , w_2813 , \1518_b0 );
buf ( \1544_b1 , \1543_b1 );
not ( \1544_b1 , w_2814 );
not ( \1544_b0 , w_2815 );
and ( w_2814 , w_2815 , \1543_b0 );
or ( \1545_b1 , \1500_b1 , \1544_b1 );
not ( \1544_b1 , w_2816 );
and ( \1545_b0 , \1500_b0 , w_2817 );
and ( w_2816 , w_2817 , \1544_b0 );
or ( \1546_b1 , \1542_b1 , w_2818 );
xor ( \1546_b0 , \1542_b0 , w_2820 );
not ( w_2820 , w_2821 );
and ( w_2821 , w_2818 , w_2819 );
buf ( w_2818 , \1545_b1 );
not ( w_2818 , w_2822 );
not ( w_2819 , w_2823 );
and ( w_2822 , w_2823 , \1545_b0 );
or ( \1547_b1 , \1532_b1 , \1546_b1 );
xor ( \1547_b0 , \1532_b0 , w_2824 );
not ( w_2824 , w_2825 );
and ( w_2825 , \1546_b1 , \1546_b0 );
buf ( \1548_b1 , \1301_B[29]_b1 );
buf ( \1548_b0 , \1301_B[29]_b0 );
or ( \1549_b1 , \1548_b1 , \1499_b1 );
xor ( \1549_b0 , \1548_b0 , w_2826 );
not ( w_2826 , w_2827 );
and ( w_2827 , \1499_b1 , \1499_b0 );
buf ( \1550_b1 , \1501_b1 );
not ( \1550_b1 , w_2828 );
not ( \1550_b0 , w_2829 );
and ( w_2828 , w_2829 , \1501_b0 );
or ( \1551_b1 , \1549_b1 , \1550_b1 );
not ( \1550_b1 , w_2830 );
and ( \1551_b0 , \1549_b0 , w_2831 );
and ( w_2830 , w_2831 , \1550_b0 );
or ( \1552_b1 , \1498_b1 , \1551_b1 );
not ( \1551_b1 , w_2832 );
and ( \1552_b0 , \1498_b0 , w_2833 );
and ( w_2832 , w_2833 , \1551_b0 );
buf ( \1553_b1 , \1295_A[1]_b1 );
buf ( \1553_b0 , \1295_A[1]_b0 );
or ( \1554_b1 , \1553_b1 , \1501_b1 );
not ( \1501_b1 , w_2834 );
and ( \1554_b0 , \1553_b0 , w_2835 );
and ( w_2834 , w_2835 , \1501_b0 );
or ( \1555_b1 , \1552_b1 , w_2837 );
not ( w_2837 , w_2838 );
and ( \1555_b0 , \1552_b0 , w_2839 );
and ( w_2838 ,  , w_2839 );
buf ( w_2837 , \1554_b1 );
not ( w_2837 , w_2840 );
not (  , w_2841 );
and ( w_2840 , w_2841 , \1554_b0 );
or ( \1556_b1 , \1499_b1 , \1500_b1 );
not ( \1500_b1 , w_2842 );
and ( \1556_b0 , \1499_b0 , w_2843 );
and ( w_2842 , w_2843 , \1500_b0 );
buf ( \1557_b1 , \1556_b1 );
not ( \1557_b1 , w_2844 );
not ( \1557_b0 , w_2845 );
and ( w_2844 , w_2845 , \1556_b0 );
or ( \1558_b1 , \1548_b1 , \1557_b1 );
not ( \1557_b1 , w_2846 );
and ( \1558_b0 , \1548_b0 , w_2847 );
and ( w_2846 , w_2847 , \1557_b0 );
or ( \1559_b1 , \1555_b1 , w_2848 );
xor ( \1559_b0 , \1555_b0 , w_2850 );
not ( w_2850 , w_2851 );
and ( w_2851 , w_2848 , w_2849 );
buf ( w_2848 , \1558_b1 );
not ( w_2848 , w_2852 );
not ( w_2849 , w_2853 );
and ( w_2852 , w_2853 , \1558_b0 );
or ( \1560_b1 , \1547_b1 , \1559_b1 );
xor ( \1560_b0 , \1547_b0 , w_2854 );
not ( w_2854 , w_2855 );
and ( w_2855 , \1559_b1 , \1559_b0 );
or ( \1561_b1 , \1384_b1 , \1382_b1 );
not ( \1382_b1 , w_2856 );
and ( \1561_b0 , \1384_b0 , w_2857 );
and ( w_2856 , w_2857 , \1382_b0 );
or ( \1562_b1 , \1342_b1 , \1380_b1 );
not ( \1380_b1 , w_2858 );
and ( \1562_b0 , \1342_b0 , w_2859 );
and ( w_2858 , w_2859 , \1380_b0 );
or ( \1563_b1 , \1561_b1 , w_2861 );
not ( w_2861 , w_2862 );
and ( \1563_b0 , \1561_b0 , w_2863 );
and ( w_2862 ,  , w_2863 );
buf ( w_2861 , \1562_b1 );
not ( w_2861 , w_2864 );
not (  , w_2865 );
and ( w_2864 , w_2865 , \1562_b0 );
or ( \1564_b1 , \1563_b1 , w_2866 );
xor ( \1564_b0 , \1563_b0 , w_2868 );
not ( w_2868 , w_2869 );
and ( w_2869 , w_2866 , w_2867 );
buf ( w_2866 , \1389_b1 );
not ( w_2866 , w_2870 );
not ( w_2867 , w_2871 );
and ( w_2870 , w_2871 , \1389_b0 );
or ( \1565_b1 , \1368_b1 , \1366_b1 );
not ( \1366_b1 , w_2872 );
and ( \1565_b0 , \1368_b0 , w_2873 );
and ( w_2872 , w_2873 , \1366_b0 );
or ( \1566_b1 , \1470_b1 , \1364_b1 );
not ( \1364_b1 , w_2874 );
and ( \1566_b0 , \1470_b0 , w_2875 );
and ( w_2874 , w_2875 , \1364_b0 );
or ( \1567_b1 , \1565_b1 , w_2877 );
not ( w_2877 , w_2878 );
and ( \1567_b0 , \1565_b0 , w_2879 );
and ( w_2878 ,  , w_2879 );
buf ( w_2877 , \1566_b1 );
not ( w_2877 , w_2880 );
not (  , w_2881 );
and ( w_2880 , w_2881 , \1566_b0 );
or ( \1568_b1 , \1567_b1 , w_2882 );
xor ( \1568_b0 , \1567_b0 , w_2884 );
not ( w_2884 , w_2885 );
and ( w_2885 , w_2882 , w_2883 );
buf ( w_2882 , \1373_b1 );
not ( w_2882 , w_2886 );
not ( w_2883 , w_2887 );
and ( w_2886 , w_2887 , \1373_b0 );
or ( \1569_b1 , \1564_b1 , \1568_b1 );
xor ( \1569_b0 , \1564_b0 , w_2888 );
not ( w_2888 , w_2889 );
and ( w_2889 , \1568_b1 , \1568_b0 );
or ( \1570_b1 , \1399_b1 , \1397_b1 );
not ( \1397_b1 , w_2890 );
and ( \1570_b0 , \1399_b0 , w_2891 );
and ( w_2890 , w_2891 , \1397_b0 );
or ( \1571_b1 , \1359_b1 , \1395_b1 );
not ( \1395_b1 , w_2892 );
and ( \1571_b0 , \1359_b0 , w_2893 );
and ( w_2892 , w_2893 , \1395_b0 );
or ( \1572_b1 , \1570_b1 , w_2895 );
not ( w_2895 , w_2896 );
and ( \1572_b0 , \1570_b0 , w_2897 );
and ( w_2896 ,  , w_2897 );
buf ( w_2895 , \1571_b1 );
not ( w_2895 , w_2898 );
not (  , w_2899 );
and ( w_2898 , w_2899 , \1571_b0 );
or ( \1573_b1 , \1572_b1 , w_2900 );
xor ( \1573_b0 , \1572_b0 , w_2902 );
not ( w_2902 , w_2903 );
and ( w_2903 , w_2900 , w_2901 );
buf ( w_2900 , \1404_b1 );
not ( w_2900 , w_2904 );
not ( w_2901 , w_2905 );
and ( w_2904 , w_2905 , \1404_b0 );
or ( \1574_b1 , \1569_b1 , \1573_b1 );
xor ( \1574_b0 , \1569_b0 , w_2906 );
not ( w_2906 , w_2907 );
and ( w_2907 , \1573_b1 , \1573_b0 );
or ( \1575_b1 , \1560_b1 , \1574_b1 );
xor ( \1575_b0 , \1560_b0 , w_2908 );
not ( w_2908 , w_2909 );
and ( w_2909 , \1574_b1 , \1574_b0 );
or ( \1576_b1 , \1462_b1 , \1460_b1 );
not ( \1460_b1 , w_2910 );
and ( \1576_b0 , \1462_b0 , w_2911 );
and ( w_2910 , w_2911 , \1460_b0 );
or ( \1577_b1 , \1376_b1 , \1458_b1 );
not ( \1458_b1 , w_2912 );
and ( \1577_b0 , \1376_b0 , w_2913 );
and ( w_2912 , w_2913 , \1458_b0 );
or ( \1578_b1 , \1576_b1 , w_2915 );
not ( w_2915 , w_2916 );
and ( \1578_b0 , \1576_b0 , w_2917 );
and ( w_2916 ,  , w_2917 );
buf ( w_2915 , \1577_b1 );
not ( w_2915 , w_2918 );
not (  , w_2919 );
and ( w_2918 , w_2919 , \1577_b0 );
or ( \1579_b1 , \1578_b1 , w_2920 );
xor ( \1579_b0 , \1578_b0 , w_2922 );
not ( w_2922 , w_2923 );
and ( w_2923 , w_2920 , w_2921 );
buf ( w_2920 , \1467_b1 );
not ( w_2920 , w_2924 );
not ( w_2921 , w_2925 );
and ( w_2924 , w_2925 , \1467_b0 );
or ( \1580_b1 , \1477_b1 , \1475_b1 );
not ( \1475_b1 , w_2926 );
and ( \1580_b0 , \1477_b0 , w_2927 );
and ( w_2926 , w_2927 , \1475_b0 );
or ( \1581_b1 , \1454_b1 , \1473_b1 );
not ( \1473_b1 , w_2928 );
and ( \1581_b0 , \1454_b0 , w_2929 );
and ( w_2928 , w_2929 , \1473_b0 );
or ( \1582_b1 , \1580_b1 , w_2931 );
not ( w_2931 , w_2932 );
and ( \1582_b0 , \1580_b0 , w_2933 );
and ( w_2932 ,  , w_2933 );
buf ( w_2931 , \1581_b1 );
not ( w_2931 , w_2934 );
not (  , w_2935 );
and ( w_2934 , w_2935 , \1581_b0 );
or ( \1583_b1 , \1582_b1 , w_2936 );
xor ( \1583_b0 , \1582_b0 , w_2938 );
not ( w_2938 , w_2939 );
and ( w_2939 , w_2936 , w_2937 );
buf ( w_2936 , \1482_b1 );
not ( w_2936 , w_2940 );
not ( w_2937 , w_2941 );
and ( w_2940 , w_2941 , \1482_b0 );
or ( \1584_b1 , \1579_b1 , \1583_b1 );
xor ( \1584_b0 , \1579_b0 , w_2942 );
not ( w_2942 , w_2943 );
and ( w_2943 , \1583_b1 , \1583_b0 );
or ( \1585_b1 , \1416_b1 , \1414_b1 );
not ( \1414_b1 , w_2944 );
and ( \1585_b0 , \1416_b0 , w_2945 );
and ( w_2944 , w_2945 , \1414_b0 );
buf ( \1586_b1 , \1263_A[9]_b1 );
buf ( \1586_b0 , \1263_A[9]_b0 );
or ( \1587_b1 , \1586_b1 , \1412_b1 );
not ( \1412_b1 , w_2946 );
and ( \1587_b0 , \1586_b0 , w_2947 );
and ( w_2946 , w_2947 , \1412_b0 );
or ( \1588_b1 , \1585_b1 , w_2949 );
not ( w_2949 , w_2950 );
and ( \1588_b0 , \1585_b0 , w_2951 );
and ( w_2950 ,  , w_2951 );
buf ( w_2949 , \1587_b1 );
not ( w_2949 , w_2952 );
not (  , w_2953 );
and ( w_2952 , w_2953 , \1587_b0 );
or ( \1589_b1 , \1588_b1 , w_2954 );
xor ( \1589_b0 , \1588_b0 , w_2956 );
not ( w_2956 , w_2957 );
and ( w_2957 , w_2954 , w_2955 );
buf ( w_2954 , \1421_b1 );
not ( w_2954 , w_2958 );
not ( w_2955 , w_2959 );
and ( w_2958 , w_2959 , \1421_b0 );
or ( \1590_b1 , \1584_b1 , \1589_b1 );
xor ( \1590_b0 , \1584_b0 , w_2960 );
not ( w_2960 , w_2961 );
and ( w_2961 , \1589_b1 , \1589_b0 );
or ( \1591_b1 , \1575_b1 , \1590_b1 );
xor ( \1591_b0 , \1575_b0 , w_2962 );
not ( w_2962 , w_2963 );
and ( w_2963 , \1590_b1 , \1590_b0 );
or ( \1592_b1 , \1515_b1 , \1591_b1 );
not ( \1591_b1 , w_2964 );
and ( \1592_b0 , \1515_b0 , w_2965 );
and ( w_2964 , w_2965 , \1591_b0 );
or ( \1593_b1 , \1487_b1 , \1591_b1 );
not ( \1591_b1 , w_2966 );
and ( \1593_b0 , \1487_b0 , w_2967 );
and ( w_2966 , w_2967 , \1591_b0 );
or ( \1595_b1 , \1433_b1 , \1336_b1 );
not ( \1336_b1 , w_2968 );
and ( \1595_b0 , \1433_b0 , w_2969 );
and ( w_2968 , w_2969 , \1336_b0 );
or ( \1596_b1 , \1489_b1 , \1333_b1 );
not ( \1333_b1 , w_2970 );
and ( \1596_b0 , \1489_b0 , w_2971 );
and ( w_2970 , w_2971 , \1333_b0 );
or ( \1597_b1 , \1595_b1 , w_2973 );
not ( w_2973 , w_2974 );
and ( \1597_b0 , \1595_b0 , w_2975 );
and ( w_2974 ,  , w_2975 );
buf ( w_2973 , \1596_b1 );
not ( w_2973 , w_2976 );
not (  , w_2977 );
and ( w_2976 , w_2977 , \1596_b0 );
or ( \1598_b1 , \1597_b1 , w_2978 );
xor ( \1598_b0 , \1597_b0 , w_2980 );
not ( w_2980 , w_2981 );
and ( w_2981 , w_2978 , w_2979 );
buf ( w_2978 , \1332_b1 );
not ( w_2978 , w_2982 );
not ( w_2979 , w_2983 );
and ( w_2982 , w_2983 , \1332_b0 );
or ( \1599_b1 , \1376_b1 , \1349_b1 );
not ( \1349_b1 , w_2984 );
and ( \1599_b0 , \1376_b0 , w_2985 );
and ( w_2984 , w_2985 , \1349_b0 );
or ( \1600_b1 , \1384_b1 , \1347_b1 );
not ( \1347_b1 , w_2986 );
and ( \1600_b0 , \1384_b0 , w_2987 );
and ( w_2986 , w_2987 , \1347_b0 );
or ( \1601_b1 , \1599_b1 , w_2989 );
not ( w_2989 , w_2990 );
and ( \1601_b0 , \1599_b0 , w_2991 );
and ( w_2990 ,  , w_2991 );
buf ( w_2989 , \1600_b1 );
not ( w_2989 , w_2992 );
not (  , w_2993 );
and ( w_2992 , w_2993 , \1600_b0 );
or ( \1602_b1 , \1601_b1 , w_2994 );
xor ( \1602_b0 , \1601_b0 , w_2996 );
not ( w_2996 , w_2997 );
and ( w_2997 , w_2994 , w_2995 );
buf ( w_2994 , \1356_b1 );
not ( w_2994 , w_2998 );
not ( w_2995 , w_2999 );
and ( w_2998 , w_2999 , \1356_b0 );
or ( \1603_b1 , \1598_b1 , \1602_b1 );
not ( \1602_b1 , w_3000 );
and ( \1603_b0 , \1598_b0 , w_3001 );
and ( w_3000 , w_3001 , \1602_b0 );
or ( \1604_b1 , \1391_b1 , \1366_b1 );
not ( \1366_b1 , w_3002 );
and ( \1604_b0 , \1391_b0 , w_3003 );
and ( w_3002 , w_3003 , \1366_b0 );
or ( \1605_b1 , \1399_b1 , \1364_b1 );
not ( \1364_b1 , w_3004 );
and ( \1605_b0 , \1399_b0 , w_3005 );
and ( w_3004 , w_3005 , \1364_b0 );
or ( \1606_b1 , \1604_b1 , w_3007 );
not ( w_3007 , w_3008 );
and ( \1606_b0 , \1604_b0 , w_3009 );
and ( w_3008 ,  , w_3009 );
buf ( w_3007 , \1605_b1 );
not ( w_3007 , w_3010 );
not (  , w_3011 );
and ( w_3010 , w_3011 , \1605_b0 );
or ( \1607_b1 , \1606_b1 , w_3012 );
xor ( \1607_b0 , \1606_b0 , w_3014 );
not ( w_3014 , w_3015 );
and ( w_3015 , w_3012 , w_3013 );
buf ( w_3012 , \1373_b1 );
not ( w_3012 , w_3016 );
not ( w_3013 , w_3017 );
and ( w_3016 , w_3017 , \1373_b0 );
or ( \1608_b1 , \1602_b1 , \1607_b1 );
not ( \1607_b1 , w_3018 );
and ( \1608_b0 , \1602_b0 , w_3019 );
and ( w_3018 , w_3019 , \1607_b0 );
or ( \1609_b1 , \1598_b1 , \1607_b1 );
not ( \1607_b1 , w_3020 );
and ( \1609_b0 , \1598_b0 , w_3021 );
and ( w_3020 , w_3021 , \1607_b0 );
or ( \1611_b1 , \1454_b1 , \1382_b1 );
not ( \1382_b1 , w_3022 );
and ( \1611_b0 , \1454_b0 , w_3023 );
and ( w_3022 , w_3023 , \1382_b0 );
or ( \1612_b1 , \1462_b1 , \1380_b1 );
not ( \1380_b1 , w_3024 );
and ( \1612_b0 , \1462_b0 , w_3025 );
and ( w_3024 , w_3025 , \1380_b0 );
or ( \1613_b1 , \1611_b1 , w_3027 );
not ( w_3027 , w_3028 );
and ( \1613_b0 , \1611_b0 , w_3029 );
and ( w_3028 ,  , w_3029 );
buf ( w_3027 , \1612_b1 );
not ( w_3027 , w_3030 );
not (  , w_3031 );
and ( w_3030 , w_3031 , \1612_b0 );
or ( \1614_b1 , \1613_b1 , w_3032 );
xor ( \1614_b0 , \1613_b0 , w_3034 );
not ( w_3034 , w_3035 );
and ( w_3035 , w_3032 , w_3033 );
buf ( w_3032 , \1389_b1 );
not ( w_3032 , w_3036 );
not ( w_3033 , w_3037 );
and ( w_3036 , w_3037 , \1389_b0 );
or ( \1615_b1 , \1586_b1 , \1397_b1 );
not ( \1397_b1 , w_3038 );
and ( \1615_b0 , \1586_b0 , w_3039 );
and ( w_3038 , w_3039 , \1397_b0 );
buf ( \1616_b1 , \1259_A[10]_b1 );
buf ( \1616_b0 , \1259_A[10]_b0 );
or ( \1617_b1 , \1616_b1 , \1395_b1 );
not ( \1395_b1 , w_3040 );
and ( \1617_b0 , \1616_b0 , w_3041 );
and ( w_3040 , w_3041 , \1395_b0 );
or ( \1618_b1 , \1615_b1 , w_3043 );
not ( w_3043 , w_3044 );
and ( \1618_b0 , \1615_b0 , w_3045 );
and ( w_3044 ,  , w_3045 );
buf ( w_3043 , \1617_b1 );
not ( w_3043 , w_3046 );
not (  , w_3047 );
and ( w_3046 , w_3047 , \1617_b0 );
or ( \1619_b1 , \1618_b1 , w_3048 );
xor ( \1619_b0 , \1618_b0 , w_3050 );
not ( w_3050 , w_3051 );
and ( w_3051 , w_3048 , w_3049 );
buf ( w_3048 , \1404_b1 );
not ( w_3048 , w_3052 );
not ( w_3049 , w_3053 );
and ( w_3052 , w_3053 , \1404_b0 );
or ( \1620_b1 , \1614_b1 , \1619_b1 );
not ( \1619_b1 , w_3054 );
and ( \1620_b0 , \1614_b0 , w_3055 );
and ( w_3054 , w_3055 , \1619_b0 );
or ( \1621_b1 , \1526_b1 , \1414_b1 );
not ( \1414_b1 , w_3056 );
and ( \1621_b0 , \1526_b0 , w_3057 );
and ( w_3056 , w_3057 , \1414_b0 );
buf ( \1622_b1 , \1275_A[6]_b1 );
buf ( \1622_b0 , \1275_A[6]_b0 );
or ( \1623_b1 , \1622_b1 , \1412_b1 );
not ( \1412_b1 , w_3058 );
and ( \1623_b0 , \1622_b0 , w_3059 );
and ( w_3058 , w_3059 , \1412_b0 );
or ( \1624_b1 , \1621_b1 , w_3061 );
not ( w_3061 , w_3062 );
and ( \1624_b0 , \1621_b0 , w_3063 );
and ( w_3062 ,  , w_3063 );
buf ( w_3061 , \1623_b1 );
not ( w_3061 , w_3064 );
not (  , w_3065 );
and ( w_3064 , w_3065 , \1623_b0 );
or ( \1625_b1 , \1624_b1 , w_3066 );
xor ( \1625_b0 , \1624_b0 , w_3068 );
not ( w_3068 , w_3069 );
and ( w_3069 , w_3066 , w_3067 );
buf ( w_3066 , \1421_b1 );
not ( w_3066 , w_3070 );
not ( w_3067 , w_3071 );
and ( w_3070 , w_3071 , \1421_b0 );
or ( \1626_b1 , \1619_b1 , \1625_b1 );
not ( \1625_b1 , w_3072 );
and ( \1626_b0 , \1619_b0 , w_3073 );
and ( w_3072 , w_3073 , \1625_b0 );
or ( \1627_b1 , \1614_b1 , \1625_b1 );
not ( \1625_b1 , w_3074 );
and ( \1627_b0 , \1614_b0 , w_3075 );
and ( w_3074 , w_3075 , \1625_b0 );
or ( \1629_b1 , \1610_b1 , \1628_b1 );
not ( \1628_b1 , w_3076 );
and ( \1629_b0 , \1610_b0 , w_3077 );
and ( w_3076 , w_3077 , \1628_b0 );
or ( \1630_b1 , \1351_b1 , \1431_b1 );
not ( \1431_b1 , w_3078 );
and ( \1630_b0 , \1351_b0 , w_3079 );
and ( w_3078 , w_3079 , \1431_b0 );
or ( \1631_b1 , \1446_b1 , \1429_b1 );
not ( \1429_b1 , w_3080 );
and ( \1631_b0 , \1446_b0 , w_3081 );
and ( w_3080 , w_3081 , \1429_b0 );
or ( \1632_b1 , \1630_b1 , w_3083 );
not ( w_3083 , w_3084 );
and ( \1632_b0 , \1630_b0 , w_3085 );
and ( w_3084 ,  , w_3085 );
buf ( w_3083 , \1631_b1 );
not ( w_3083 , w_3086 );
not (  , w_3087 );
and ( w_3086 , w_3087 , \1631_b0 );
or ( \1633_b1 , \1632_b1 , w_3088 );
xor ( \1633_b0 , \1632_b0 , w_3090 );
not ( w_3090 , w_3091 );
and ( w_3091 , w_3088 , w_3089 );
buf ( w_3088 , \1438_b1 );
not ( w_3088 , w_3092 );
not ( w_3089 , w_3093 );
and ( w_3092 , w_3093 , \1438_b0 );
or ( \1634_b1 , \1384_b1 , \1444_b1 );
not ( \1444_b1 , w_3094 );
and ( \1634_b0 , \1384_b0 , w_3095 );
and ( w_3094 , w_3095 , \1444_b0 );
or ( \1635_b1 , \1342_b1 , \1442_b1 );
not ( \1442_b1 , w_3096 );
and ( \1635_b0 , \1342_b0 , w_3097 );
and ( w_3096 , w_3097 , \1442_b0 );
or ( \1636_b1 , \1634_b1 , w_3099 );
not ( w_3099 , w_3100 );
and ( \1636_b0 , \1634_b0 , w_3101 );
and ( w_3100 ,  , w_3101 );
buf ( w_3099 , \1635_b1 );
not ( w_3099 , w_3102 );
not (  , w_3103 );
and ( w_3102 , w_3103 , \1635_b0 );
or ( \1637_b1 , \1636_b1 , w_3104 );
xor ( \1637_b0 , \1636_b0 , w_3106 );
not ( w_3106 , w_3107 );
and ( w_3107 , w_3104 , w_3105 );
buf ( w_3104 , \1451_b1 );
not ( w_3104 , w_3108 );
not ( w_3105 , w_3109 );
and ( w_3108 , w_3109 , \1451_b0 );
or ( \1638_b1 , \1633_b1 , \1637_b1 );
not ( \1637_b1 , w_3110 );
and ( \1638_b0 , \1633_b0 , w_3111 );
and ( w_3110 , w_3111 , \1637_b0 );
buf ( \1639_b1 , \1308_B[22]_b1 );
buf ( \1639_b0 , \1308_B[22]_b0 );
or ( \1640_b1 , \1521_b1 , \1639_b1 );
xor ( \1640_b0 , \1521_b0 , w_3112 );
not ( w_3112 , w_3113 );
and ( w_3113 , \1639_b1 , \1639_b0 );
or ( \1641_b1 , \1639_b1 , \1408_b1 );
xor ( \1641_b0 , \1639_b0 , w_3114 );
not ( w_3114 , w_3115 );
and ( w_3115 , \1408_b1 , \1408_b0 );
buf ( \1642_b1 , \1641_b1 );
not ( \1642_b1 , w_3116 );
not ( \1642_b0 , w_3117 );
and ( w_3116 , w_3117 , \1641_b0 );
or ( \1643_b1 , \1640_b1 , \1642_b1 );
not ( \1642_b1 , w_3118 );
and ( \1643_b0 , \1640_b0 , w_3119 );
and ( w_3118 , w_3119 , \1642_b0 );
or ( \1644_b1 , \1540_b1 , \1643_b1 );
not ( \1643_b1 , w_3120 );
and ( \1644_b0 , \1540_b0 , w_3121 );
and ( w_3120 , w_3121 , \1643_b0 );
or ( \1645_b1 , \1517_b1 , \1641_b1 );
not ( \1641_b1 , w_3122 );
and ( \1645_b0 , \1517_b0 , w_3123 );
and ( w_3122 , w_3123 , \1641_b0 );
or ( \1646_b1 , \1644_b1 , w_3125 );
not ( w_3125 , w_3126 );
and ( \1646_b0 , \1644_b0 , w_3127 );
and ( w_3126 ,  , w_3127 );
buf ( w_3125 , \1645_b1 );
not ( w_3125 , w_3128 );
not (  , w_3129 );
and ( w_3128 , w_3129 , \1645_b0 );
or ( \1647_b1 , \1639_b1 , \1408_b1 );
not ( \1408_b1 , w_3130 );
and ( \1647_b0 , \1639_b0 , w_3131 );
and ( w_3130 , w_3131 , \1408_b0 );
buf ( \1648_b1 , \1647_b1 );
not ( \1648_b1 , w_3132 );
not ( \1648_b0 , w_3133 );
and ( w_3132 , w_3133 , \1647_b0 );
or ( \1649_b1 , \1521_b1 , \1648_b1 );
not ( \1648_b1 , w_3134 );
and ( \1649_b0 , \1521_b0 , w_3135 );
and ( w_3134 , w_3135 , \1648_b0 );
or ( \1650_b1 , \1646_b1 , w_3136 );
xor ( \1650_b0 , \1646_b0 , w_3138 );
not ( w_3138 , w_3139 );
and ( w_3139 , w_3136 , w_3137 );
buf ( w_3136 , \1649_b1 );
not ( w_3136 , w_3140 );
not ( w_3137 , w_3141 );
and ( w_3140 , w_3141 , \1649_b0 );
or ( \1651_b1 , \1638_b1 , \1650_b1 );
not ( \1650_b1 , w_3142 );
and ( \1651_b0 , \1638_b0 , w_3143 );
and ( w_3142 , w_3143 , \1650_b0 );
or ( \1652_b1 , \1553_b1 , \1524_b1 );
not ( \1524_b1 , w_3144 );
and ( \1652_b0 , \1553_b0 , w_3145 );
and ( w_3144 , w_3145 , \1524_b0 );
or ( \1653_b1 , \1533_b1 , \1522_b1 );
not ( \1522_b1 , w_3146 );
and ( \1653_b0 , \1533_b0 , w_3147 );
and ( w_3146 , w_3147 , \1522_b0 );
or ( \1654_b1 , \1652_b1 , w_3149 );
not ( w_3149 , w_3150 );
and ( \1654_b0 , \1652_b0 , w_3151 );
and ( w_3150 ,  , w_3151 );
buf ( w_3149 , \1653_b1 );
not ( w_3149 , w_3152 );
not (  , w_3153 );
and ( w_3152 , w_3153 , \1653_b0 );
or ( \1655_b1 , \1654_b1 , w_3154 );
xor ( \1655_b0 , \1654_b0 , w_3156 );
not ( w_3156 , w_3157 );
and ( w_3157 , w_3154 , w_3155 );
buf ( w_3154 , \1531_b1 );
not ( w_3154 , w_3158 );
not ( w_3155 , w_3159 );
and ( w_3158 , w_3159 , \1531_b0 );
or ( \1656_b1 , \1650_b1 , \1655_b1 );
not ( \1655_b1 , w_3160 );
and ( \1656_b0 , \1650_b0 , w_3161 );
and ( w_3160 , w_3161 , \1655_b0 );
or ( \1657_b1 , \1638_b1 , \1655_b1 );
not ( \1655_b1 , w_3162 );
and ( \1657_b0 , \1638_b0 , w_3163 );
and ( w_3162 , w_3163 , \1655_b0 );
or ( \1659_b1 , \1628_b1 , \1658_b1 );
not ( \1658_b1 , w_3164 );
and ( \1659_b0 , \1628_b0 , w_3165 );
and ( w_3164 , w_3165 , \1658_b0 );
or ( \1660_b1 , \1610_b1 , \1658_b1 );
not ( \1658_b1 , w_3166 );
and ( \1660_b0 , \1610_b0 , w_3167 );
and ( w_3166 , w_3167 , \1658_b0 );
or ( \1662_b1 , \1470_b1 , \1460_b1 );
not ( \1460_b1 , w_3168 );
and ( \1662_b0 , \1470_b0 , w_3169 );
and ( w_3168 , w_3169 , \1460_b0 );
or ( \1663_b1 , \1477_b1 , \1458_b1 );
not ( \1458_b1 , w_3170 );
and ( \1663_b0 , \1477_b0 , w_3171 );
and ( w_3170 , w_3171 , \1458_b0 );
or ( \1664_b1 , \1662_b1 , w_3173 );
not ( w_3173 , w_3174 );
and ( \1664_b0 , \1662_b0 , w_3175 );
and ( w_3174 ,  , w_3175 );
buf ( w_3173 , \1663_b1 );
not ( w_3173 , w_3176 );
not (  , w_3177 );
and ( w_3176 , w_3177 , \1663_b0 );
or ( \1665_b1 , \1664_b1 , w_3178 );
xor ( \1665_b0 , \1664_b0 , w_3180 );
not ( w_3180 , w_3181 );
and ( w_3181 , w_3178 , w_3179 );
buf ( w_3178 , \1467_b1 );
not ( w_3178 , w_3182 );
not ( w_3179 , w_3183 );
and ( w_3182 , w_3183 , \1467_b0 );
or ( \1666_b1 , \1359_b1 , \1475_b1 );
not ( \1475_b1 , w_3184 );
and ( \1666_b0 , \1359_b0 , w_3185 );
and ( w_3184 , w_3185 , \1475_b0 );
or ( \1667_b1 , \1368_b1 , \1473_b1 );
not ( \1473_b1 , w_3186 );
and ( \1667_b0 , \1368_b0 , w_3187 );
and ( w_3186 , w_3187 , \1473_b0 );
or ( \1668_b1 , \1666_b1 , w_3189 );
not ( w_3189 , w_3190 );
and ( \1668_b0 , \1666_b0 , w_3191 );
and ( w_3190 ,  , w_3191 );
buf ( w_3189 , \1667_b1 );
not ( w_3189 , w_3192 );
not (  , w_3193 );
and ( w_3192 , w_3193 , \1667_b0 );
or ( \1669_b1 , \1668_b1 , w_3194 );
xor ( \1669_b0 , \1668_b0 , w_3196 );
not ( w_3196 , w_3197 );
and ( w_3197 , w_3194 , w_3195 );
buf ( w_3194 , \1482_b1 );
not ( w_3194 , w_3198 );
not ( w_3195 , w_3199 );
and ( w_3198 , w_3199 , \1482_b0 );
or ( \1670_b1 , \1665_b1 , \1669_b1 );
not ( \1669_b1 , w_3200 );
and ( \1670_b0 , \1665_b0 , w_3201 );
and ( w_3200 , w_3201 , \1669_b0 );
buf ( \1671_b1 , \1312_B[18]_b1 );
buf ( \1671_b0 , \1312_B[18]_b0 );
or ( \1672_b1 , \1411_b1 , \1671_b1 );
xor ( \1672_b0 , \1411_b0 , w_3202 );
not ( w_3202 , w_3203 );
and ( w_3203 , \1671_b1 , \1671_b0 );
or ( \1673_b1 , \1671_b1 , \1392_b1 );
xor ( \1673_b0 , \1671_b0 , w_3204 );
not ( w_3204 , w_3205 );
and ( w_3205 , \1392_b1 , \1392_b0 );
buf ( \1674_b1 , \1673_b1 );
not ( \1674_b1 , w_3206 );
not ( \1674_b0 , w_3207 );
and ( w_3206 , w_3207 , \1673_b0 );
or ( \1675_b1 , \1672_b1 , \1674_b1 );
not ( \1674_b1 , w_3208 );
and ( \1675_b0 , \1672_b0 , w_3209 );
and ( w_3208 , w_3209 , \1674_b0 );
or ( \1676_b1 , \1407_b1 , \1675_b1 );
not ( \1675_b1 , w_3210 );
and ( \1676_b0 , \1407_b0 , w_3211 );
and ( w_3210 , w_3211 , \1675_b0 );
or ( \1677_b1 , \1416_b1 , \1673_b1 );
not ( \1673_b1 , w_3212 );
and ( \1677_b0 , \1416_b0 , w_3213 );
and ( w_3212 , w_3213 , \1673_b0 );
or ( \1678_b1 , \1676_b1 , w_3215 );
not ( w_3215 , w_3216 );
and ( \1678_b0 , \1676_b0 , w_3217 );
and ( w_3216 ,  , w_3217 );
buf ( w_3215 , \1677_b1 );
not ( w_3215 , w_3218 );
not (  , w_3219 );
and ( w_3218 , w_3219 , \1677_b0 );
or ( \1679_b1 , \1671_b1 , \1392_b1 );
not ( \1392_b1 , w_3220 );
and ( \1679_b0 , \1671_b0 , w_3221 );
and ( w_3220 , w_3221 , \1392_b0 );
buf ( \1680_b1 , \1679_b1 );
not ( \1680_b1 , w_3222 );
not ( \1680_b0 , w_3223 );
and ( w_3222 , w_3223 , \1679_b0 );
or ( \1681_b1 , \1411_b1 , \1680_b1 );
not ( \1680_b1 , w_3224 );
and ( \1681_b0 , \1411_b0 , w_3225 );
and ( w_3224 , w_3225 , \1680_b0 );
or ( \1682_b1 , \1678_b1 , w_3226 );
xor ( \1682_b0 , \1678_b0 , w_3228 );
not ( w_3228 , w_3229 );
and ( w_3229 , w_3226 , w_3227 );
buf ( w_3226 , \1681_b1 );
not ( w_3226 , w_3230 );
not ( w_3227 , w_3231 );
and ( w_3230 , w_3231 , \1681_b0 );
or ( \1683_b1 , \1669_b1 , \1682_b1 );
not ( \1682_b1 , w_3232 );
and ( \1683_b0 , \1669_b0 , w_3233 );
and ( w_3232 , w_3233 , \1682_b0 );
or ( \1684_b1 , \1665_b1 , \1682_b1 );
not ( \1682_b1 , w_3234 );
and ( \1684_b0 , \1665_b0 , w_3235 );
and ( w_3234 , w_3235 , \1682_b0 );
or ( \1686_b1 , \1462_b1 , \1382_b1 );
not ( \1382_b1 , w_3236 );
and ( \1686_b0 , \1462_b0 , w_3237 );
and ( w_3236 , w_3237 , \1382_b0 );
or ( \1687_b1 , \1376_b1 , \1380_b1 );
not ( \1380_b1 , w_3238 );
and ( \1687_b0 , \1376_b0 , w_3239 );
and ( w_3238 , w_3239 , \1380_b0 );
or ( \1688_b1 , \1686_b1 , w_3241 );
not ( w_3241 , w_3242 );
and ( \1688_b0 , \1686_b0 , w_3243 );
and ( w_3242 ,  , w_3243 );
buf ( w_3241 , \1687_b1 );
not ( w_3241 , w_3244 );
not (  , w_3245 );
and ( w_3244 , w_3245 , \1687_b0 );
or ( \1689_b1 , \1688_b1 , w_3246 );
xor ( \1689_b0 , \1688_b0 , w_3248 );
not ( w_3248 , w_3249 );
and ( w_3249 , w_3246 , w_3247 );
buf ( w_3246 , \1389_b1 );
not ( w_3246 , w_3250 );
not ( w_3247 , w_3251 );
and ( w_3250 , w_3251 , \1389_b0 );
or ( \1690_b1 , \1399_b1 , \1366_b1 );
not ( \1366_b1 , w_3252 );
and ( \1690_b0 , \1399_b0 , w_3253 );
and ( w_3252 , w_3253 , \1366_b0 );
or ( \1691_b1 , \1359_b1 , \1364_b1 );
not ( \1364_b1 , w_3254 );
and ( \1691_b0 , \1359_b0 , w_3255 );
and ( w_3254 , w_3255 , \1364_b0 );
or ( \1692_b1 , \1690_b1 , w_3257 );
not ( w_3257 , w_3258 );
and ( \1692_b0 , \1690_b0 , w_3259 );
and ( w_3258 ,  , w_3259 );
buf ( w_3257 , \1691_b1 );
not ( w_3257 , w_3260 );
not (  , w_3261 );
and ( w_3260 , w_3261 , \1691_b0 );
or ( \1693_b1 , \1692_b1 , w_3262 );
xor ( \1693_b0 , \1692_b0 , w_3264 );
not ( w_3264 , w_3265 );
and ( w_3265 , w_3262 , w_3263 );
buf ( w_3262 , \1373_b1 );
not ( w_3262 , w_3266 );
not ( w_3263 , w_3267 );
and ( w_3266 , w_3267 , \1373_b0 );
or ( \1694_b1 , \1689_b1 , \1693_b1 );
xor ( \1694_b0 , \1689_b0 , w_3268 );
not ( w_3268 , w_3269 );
and ( w_3269 , \1693_b1 , \1693_b0 );
or ( \1695_b1 , \1616_b1 , \1397_b1 );
not ( \1397_b1 , w_3270 );
and ( \1695_b0 , \1616_b0 , w_3271 );
and ( w_3270 , w_3271 , \1397_b0 );
or ( \1696_b1 , \1391_b1 , \1395_b1 );
not ( \1395_b1 , w_3272 );
and ( \1696_b0 , \1391_b0 , w_3273 );
and ( w_3272 , w_3273 , \1395_b0 );
or ( \1697_b1 , \1695_b1 , w_3275 );
not ( w_3275 , w_3276 );
and ( \1697_b0 , \1695_b0 , w_3277 );
and ( w_3276 ,  , w_3277 );
buf ( w_3275 , \1696_b1 );
not ( w_3275 , w_3278 );
not (  , w_3279 );
and ( w_3278 , w_3279 , \1696_b0 );
or ( \1698_b1 , \1697_b1 , w_3280 );
xor ( \1698_b0 , \1697_b0 , w_3282 );
not ( w_3282 , w_3283 );
and ( w_3283 , w_3280 , w_3281 );
buf ( w_3280 , \1404_b1 );
not ( w_3280 , w_3284 );
not ( w_3281 , w_3285 );
and ( w_3284 , w_3285 , \1404_b0 );
or ( \1699_b1 , \1694_b1 , \1698_b1 );
xor ( \1699_b0 , \1694_b0 , w_3286 );
not ( w_3286 , w_3287 );
and ( w_3287 , \1698_b1 , \1698_b0 );
or ( \1700_b1 , \1685_b1 , \1699_b1 );
not ( \1699_b1 , w_3288 );
and ( \1700_b0 , \1685_b0 , w_3289 );
and ( w_3288 , w_3289 , \1699_b0 );
or ( \1701_b1 , \1477_b1 , \1460_b1 );
not ( \1460_b1 , w_3290 );
and ( \1701_b0 , \1477_b0 , w_3291 );
and ( w_3290 , w_3291 , \1460_b0 );
or ( \1702_b1 , \1454_b1 , \1458_b1 );
not ( \1458_b1 , w_3292 );
and ( \1702_b0 , \1454_b0 , w_3293 );
and ( w_3292 , w_3293 , \1458_b0 );
or ( \1703_b1 , \1701_b1 , w_3295 );
not ( w_3295 , w_3296 );
and ( \1703_b0 , \1701_b0 , w_3297 );
and ( w_3296 ,  , w_3297 );
buf ( w_3295 , \1702_b1 );
not ( w_3295 , w_3298 );
not (  , w_3299 );
and ( w_3298 , w_3299 , \1702_b0 );
or ( \1704_b1 , \1703_b1 , w_3300 );
xor ( \1704_b0 , \1703_b0 , w_3302 );
not ( w_3302 , w_3303 );
and ( w_3303 , w_3300 , w_3301 );
buf ( w_3300 , \1467_b1 );
not ( w_3300 , w_3304 );
not ( w_3301 , w_3305 );
and ( w_3304 , w_3305 , \1467_b0 );
or ( \1705_b1 , \1368_b1 , \1475_b1 );
not ( \1475_b1 , w_3306 );
and ( \1705_b0 , \1368_b0 , w_3307 );
and ( w_3306 , w_3307 , \1475_b0 );
or ( \1706_b1 , \1470_b1 , \1473_b1 );
not ( \1473_b1 , w_3308 );
and ( \1706_b0 , \1470_b0 , w_3309 );
and ( w_3308 , w_3309 , \1473_b0 );
or ( \1707_b1 , \1705_b1 , w_3311 );
not ( w_3311 , w_3312 );
and ( \1707_b0 , \1705_b0 , w_3313 );
and ( w_3312 ,  , w_3313 );
buf ( w_3311 , \1706_b1 );
not ( w_3311 , w_3314 );
not (  , w_3315 );
and ( w_3314 , w_3315 , \1706_b0 );
or ( \1708_b1 , \1707_b1 , w_3316 );
xor ( \1708_b0 , \1707_b0 , w_3318 );
not ( w_3318 , w_3319 );
and ( w_3319 , w_3316 , w_3317 );
buf ( w_3316 , \1482_b1 );
not ( w_3316 , w_3320 );
not ( w_3317 , w_3321 );
and ( w_3320 , w_3321 , \1482_b0 );
or ( \1709_b1 , \1704_b1 , \1708_b1 );
xor ( \1709_b0 , \1704_b0 , w_3322 );
not ( w_3322 , w_3323 );
and ( w_3323 , \1708_b1 , \1708_b0 );
or ( \1710_b1 , \1622_b1 , \1414_b1 );
not ( \1414_b1 , w_3324 );
and ( \1710_b0 , \1622_b0 , w_3325 );
and ( w_3324 , w_3325 , \1414_b0 );
or ( \1711_b1 , \1407_b1 , \1412_b1 );
not ( \1412_b1 , w_3326 );
and ( \1711_b0 , \1407_b0 , w_3327 );
and ( w_3326 , w_3327 , \1412_b0 );
or ( \1712_b1 , \1710_b1 , w_3329 );
not ( w_3329 , w_3330 );
and ( \1712_b0 , \1710_b0 , w_3331 );
and ( w_3330 ,  , w_3331 );
buf ( w_3329 , \1711_b1 );
not ( w_3329 , w_3332 );
not (  , w_3333 );
and ( w_3332 , w_3333 , \1711_b0 );
or ( \1713_b1 , \1712_b1 , w_3334 );
xor ( \1713_b0 , \1712_b0 , w_3336 );
not ( w_3336 , w_3337 );
and ( w_3337 , w_3334 , w_3335 );
buf ( w_3334 , \1421_b1 );
not ( w_3334 , w_3338 );
not ( w_3335 , w_3339 );
and ( w_3338 , w_3339 , \1421_b0 );
or ( \1714_b1 , \1709_b1 , \1713_b1 );
xor ( \1714_b0 , \1709_b0 , w_3340 );
not ( w_3340 , w_3341 );
and ( w_3341 , \1713_b1 , \1713_b0 );
or ( \1715_b1 , \1699_b1 , \1714_b1 );
not ( \1714_b1 , w_3342 );
and ( \1715_b0 , \1699_b0 , w_3343 );
and ( w_3342 , w_3343 , \1714_b0 );
or ( \1716_b1 , \1685_b1 , \1714_b1 );
not ( \1714_b1 , w_3344 );
and ( \1716_b0 , \1685_b0 , w_3345 );
and ( w_3344 , w_3345 , \1714_b0 );
or ( \1718_b1 , \1661_b1 , \1717_b1 );
not ( \1717_b1 , w_3346 );
and ( \1718_b0 , \1661_b0 , w_3347 );
and ( w_3346 , w_3347 , \1717_b0 );
or ( \1719_b1 , \1689_b1 , \1693_b1 );
not ( \1693_b1 , w_3348 );
and ( \1719_b0 , \1689_b0 , w_3349 );
and ( w_3348 , w_3349 , \1693_b0 );
or ( \1720_b1 , \1693_b1 , \1698_b1 );
not ( \1698_b1 , w_3350 );
and ( \1720_b0 , \1693_b0 , w_3351 );
and ( w_3350 , w_3351 , \1698_b0 );
or ( \1721_b1 , \1689_b1 , \1698_b1 );
not ( \1698_b1 , w_3352 );
and ( \1721_b0 , \1689_b0 , w_3353 );
and ( w_3352 , w_3353 , \1698_b0 );
or ( \1723_b1 , \1704_b1 , \1708_b1 );
not ( \1708_b1 , w_3354 );
and ( \1723_b0 , \1704_b0 , w_3355 );
and ( w_3354 , w_3355 , \1708_b0 );
or ( \1724_b1 , \1708_b1 , \1713_b1 );
not ( \1713_b1 , w_3356 );
and ( \1724_b0 , \1708_b0 , w_3357 );
and ( w_3356 , w_3357 , \1713_b0 );
or ( \1725_b1 , \1704_b1 , \1713_b1 );
not ( \1713_b1 , w_3358 );
and ( \1725_b0 , \1704_b0 , w_3359 );
and ( w_3358 , w_3359 , \1713_b0 );
or ( \1727_b1 , \1722_b1 , \1726_b1 );
xor ( \1727_b0 , \1722_b0 , w_3360 );
not ( w_3360 , w_3361 );
and ( w_3361 , \1726_b1 , \1726_b0 );
or ( \1728_b1 , \1439_b1 , \1452_b1 );
xor ( \1728_b0 , \1439_b0 , w_3362 );
not ( w_3362 , w_3363 );
and ( w_3363 , \1452_b1 , \1452_b0 );
or ( \1729_b1 , \1416_b1 , \1675_b1 );
not ( \1675_b1 , w_3364 );
and ( \1729_b0 , \1416_b0 , w_3365 );
and ( w_3364 , w_3365 , \1675_b0 );
or ( \1730_b1 , \1586_b1 , \1673_b1 );
not ( \1673_b1 , w_3366 );
and ( \1730_b0 , \1586_b0 , w_3367 );
and ( w_3366 , w_3367 , \1673_b0 );
or ( \1731_b1 , \1729_b1 , w_3369 );
not ( w_3369 , w_3370 );
and ( \1731_b0 , \1729_b0 , w_3371 );
and ( w_3370 ,  , w_3371 );
buf ( w_3369 , \1730_b1 );
not ( w_3369 , w_3372 );
not (  , w_3373 );
and ( w_3372 , w_3373 , \1730_b0 );
or ( \1732_b1 , \1731_b1 , w_3374 );
xor ( \1732_b0 , \1731_b0 , w_3376 );
not ( w_3376 , w_3377 );
and ( w_3377 , w_3374 , w_3375 );
buf ( w_3374 , \1681_b1 );
not ( w_3374 , w_3378 );
not ( w_3375 , w_3379 );
and ( w_3378 , w_3379 , \1681_b0 );
or ( \1733_b1 , \1728_b1 , \1732_b1 );
not ( \1732_b1 , w_3380 );
and ( \1733_b0 , \1728_b0 , w_3381 );
and ( w_3380 , w_3381 , \1732_b0 );
or ( \1734_b1 , \1517_b1 , \1643_b1 );
not ( \1643_b1 , w_3382 );
and ( \1734_b0 , \1517_b0 , w_3383 );
and ( w_3382 , w_3383 , \1643_b0 );
or ( \1735_b1 , \1526_b1 , \1641_b1 );
not ( \1641_b1 , w_3384 );
and ( \1735_b0 , \1526_b0 , w_3385 );
and ( w_3384 , w_3385 , \1641_b0 );
or ( \1736_b1 , \1734_b1 , w_3387 );
not ( w_3387 , w_3388 );
and ( \1736_b0 , \1734_b0 , w_3389 );
and ( w_3388 ,  , w_3389 );
buf ( w_3387 , \1735_b1 );
not ( w_3387 , w_3390 );
not (  , w_3391 );
and ( w_3390 , w_3391 , \1735_b0 );
or ( \1737_b1 , \1736_b1 , w_3392 );
xor ( \1737_b0 , \1736_b0 , w_3394 );
not ( w_3394 , w_3395 );
and ( w_3395 , w_3392 , w_3393 );
buf ( w_3392 , \1649_b1 );
not ( w_3392 , w_3396 );
not ( w_3393 , w_3397 );
and ( w_3396 , w_3397 , \1649_b0 );
or ( \1738_b1 , \1732_b1 , \1737_b1 );
not ( \1737_b1 , w_3398 );
and ( \1738_b0 , \1732_b0 , w_3399 );
and ( w_3398 , w_3399 , \1737_b0 );
or ( \1739_b1 , \1728_b1 , \1737_b1 );
not ( \1737_b1 , w_3400 );
and ( \1739_b0 , \1728_b0 , w_3401 );
and ( w_3400 , w_3401 , \1737_b0 );
or ( \1741_b1 , \1727_b1 , \1740_b1 );
xor ( \1741_b0 , \1727_b0 , w_3402 );
not ( w_3402 , w_3403 );
and ( w_3403 , \1740_b1 , \1740_b0 );
or ( \1742_b1 , \1717_b1 , \1741_b1 );
not ( \1741_b1 , w_3404 );
and ( \1742_b0 , \1717_b0 , w_3405 );
and ( w_3404 , w_3405 , \1741_b0 );
or ( \1743_b1 , \1661_b1 , \1741_b1 );
not ( \1741_b1 , w_3406 );
and ( \1743_b0 , \1661_b0 , w_3407 );
and ( w_3406 , w_3407 , \1741_b0 );
or ( \1745_b1 , \1446_b1 , \1431_b1 );
not ( \1431_b1 , w_3408 );
and ( \1745_b0 , \1446_b0 , w_3409 );
and ( w_3408 , w_3409 , \1431_b0 );
or ( \1746_b1 , \1425_b1 , \1429_b1 );
not ( \1429_b1 , w_3410 );
and ( \1746_b0 , \1425_b0 , w_3411 );
and ( w_3410 , w_3411 , \1429_b0 );
or ( \1747_b1 , \1745_b1 , w_3413 );
not ( w_3413 , w_3414 );
and ( \1747_b0 , \1745_b0 , w_3415 );
and ( w_3414 ,  , w_3415 );
buf ( w_3413 , \1746_b1 );
not ( w_3413 , w_3416 );
not (  , w_3417 );
and ( w_3416 , w_3417 , \1746_b0 );
or ( \1748_b1 , \1747_b1 , w_3418 );
xor ( \1748_b0 , \1747_b0 , w_3420 );
not ( w_3420 , w_3421 );
and ( w_3421 , w_3418 , w_3419 );
buf ( w_3418 , \1438_b1 );
not ( w_3418 , w_3422 );
not ( w_3419 , w_3423 );
and ( w_3422 , w_3423 , \1438_b0 );
or ( \1749_b1 , \1342_b1 , \1444_b1 );
not ( \1444_b1 , w_3424 );
and ( \1749_b0 , \1342_b0 , w_3425 );
and ( w_3424 , w_3425 , \1444_b0 );
or ( \1750_b1 , \1351_b1 , \1442_b1 );
not ( \1442_b1 , w_3426 );
and ( \1750_b0 , \1351_b0 , w_3427 );
and ( w_3426 , w_3427 , \1442_b0 );
or ( \1751_b1 , \1749_b1 , w_3429 );
not ( w_3429 , w_3430 );
and ( \1751_b0 , \1749_b0 , w_3431 );
and ( w_3430 ,  , w_3431 );
buf ( w_3429 , \1750_b1 );
not ( w_3429 , w_3432 );
not (  , w_3433 );
and ( w_3432 , w_3433 , \1750_b0 );
or ( \1752_b1 , \1751_b1 , w_3434 );
xor ( \1752_b0 , \1751_b0 , w_3436 );
not ( w_3436 , w_3437 );
and ( w_3437 , w_3434 , w_3435 );
buf ( w_3434 , \1451_b1 );
not ( w_3434 , w_3438 );
not ( w_3435 , w_3439 );
and ( w_3438 , w_3439 , \1451_b0 );
or ( \1753_b1 , \1748_b1 , \1752_b1 );
not ( \1752_b1 , w_3440 );
and ( \1753_b0 , \1748_b0 , w_3441 );
and ( w_3440 , w_3441 , \1752_b0 );
or ( \1754_b1 , \1498_b1 , \1536_b1 );
not ( \1536_b1 , w_3442 );
and ( \1754_b0 , \1498_b0 , w_3443 );
and ( w_3442 , w_3443 , \1536_b0 );
or ( \1755_b1 , \1752_b1 , \1754_b1 );
not ( \1754_b1 , w_3444 );
and ( \1755_b0 , \1752_b0 , w_3445 );
and ( w_3444 , w_3445 , \1754_b0 );
or ( \1756_b1 , \1748_b1 , \1754_b1 );
not ( \1754_b1 , w_3446 );
and ( \1756_b0 , \1748_b0 , w_3447 );
and ( w_3446 , w_3447 , \1754_b0 );
or ( \1758_b1 , \1533_b1 , \1524_b1 );
not ( \1524_b1 , w_3448 );
and ( \1758_b0 , \1533_b0 , w_3449 );
and ( w_3448 , w_3449 , \1524_b0 );
or ( \1759_b1 , \1540_b1 , \1522_b1 );
not ( \1522_b1 , w_3450 );
and ( \1759_b0 , \1540_b0 , w_3451 );
and ( w_3450 , w_3451 , \1522_b0 );
or ( \1760_b1 , \1758_b1 , w_3453 );
not ( w_3453 , w_3454 );
and ( \1760_b0 , \1758_b0 , w_3455 );
and ( w_3454 ,  , w_3455 );
buf ( w_3453 , \1759_b1 );
not ( w_3453 , w_3456 );
not (  , w_3457 );
and ( w_3456 , w_3457 , \1759_b0 );
or ( \1761_b1 , \1760_b1 , w_3458 );
xor ( \1761_b0 , \1760_b0 , w_3460 );
not ( w_3460 , w_3461 );
and ( w_3461 , w_3458 , w_3459 );
buf ( w_3458 , \1531_b1 );
not ( w_3458 , w_3462 );
not ( w_3459 , w_3463 );
and ( w_3462 , w_3463 , \1531_b0 );
or ( \1762_b1 , \1757_b1 , \1761_b1 );
not ( \1761_b1 , w_3464 );
and ( \1762_b0 , \1757_b0 , w_3465 );
and ( w_3464 , w_3465 , \1761_b0 );
or ( \1763_b1 , \1498_b1 , \1538_b1 );
not ( \1538_b1 , w_3466 );
and ( \1763_b0 , \1498_b0 , w_3467 );
and ( w_3466 , w_3467 , \1538_b0 );
or ( \1764_b1 , \1553_b1 , \1536_b1 );
not ( \1536_b1 , w_3468 );
and ( \1764_b0 , \1553_b0 , w_3469 );
and ( w_3468 , w_3469 , \1536_b0 );
or ( \1765_b1 , \1763_b1 , w_3471 );
not ( w_3471 , w_3472 );
and ( \1765_b0 , \1763_b0 , w_3473 );
and ( w_3472 ,  , w_3473 );
buf ( w_3471 , \1764_b1 );
not ( w_3471 , w_3474 );
not (  , w_3475 );
and ( w_3474 , w_3475 , \1764_b0 );
or ( \1766_b1 , \1765_b1 , w_3476 );
xor ( \1766_b0 , \1765_b0 , w_3478 );
not ( w_3478 , w_3479 );
and ( w_3479 , w_3476 , w_3477 );
buf ( w_3476 , \1545_b1 );
not ( w_3476 , w_3480 );
not ( w_3477 , w_3481 );
and ( w_3480 , w_3481 , \1545_b0 );
or ( \1767_b1 , \1761_b1 , \1766_b1 );
not ( \1766_b1 , w_3482 );
and ( \1767_b0 , \1761_b0 , w_3483 );
and ( w_3482 , w_3483 , \1766_b0 );
or ( \1768_b1 , \1757_b1 , \1766_b1 );
not ( \1766_b1 , w_3484 );
and ( \1768_b0 , \1757_b0 , w_3485 );
and ( w_3484 , w_3485 , \1766_b0 );
or ( \1770_b1 , \1586_b1 , \1675_b1 );
not ( \1675_b1 , w_3486 );
and ( \1770_b0 , \1586_b0 , w_3487 );
and ( w_3486 , w_3487 , \1675_b0 );
or ( \1771_b1 , \1616_b1 , \1673_b1 );
not ( \1673_b1 , w_3488 );
and ( \1771_b0 , \1616_b0 , w_3489 );
and ( w_3488 , w_3489 , \1673_b0 );
or ( \1772_b1 , \1770_b1 , w_3491 );
not ( w_3491 , w_3492 );
and ( \1772_b0 , \1770_b0 , w_3493 );
and ( w_3492 ,  , w_3493 );
buf ( w_3491 , \1771_b1 );
not ( w_3491 , w_3494 );
not (  , w_3495 );
and ( w_3494 , w_3495 , \1771_b0 );
or ( \1773_b1 , \1772_b1 , w_3496 );
xor ( \1773_b0 , \1772_b0 , w_3498 );
not ( w_3498 , w_3499 );
and ( w_3499 , w_3496 , w_3497 );
buf ( w_3496 , \1681_b1 );
not ( w_3496 , w_3500 );
not ( w_3497 , w_3501 );
and ( w_3500 , w_3501 , \1681_b0 );
or ( \1774_b1 , \1526_b1 , \1643_b1 );
not ( \1643_b1 , w_3502 );
and ( \1774_b0 , \1526_b0 , w_3503 );
and ( w_3502 , w_3503 , \1643_b0 );
or ( \1775_b1 , \1622_b1 , \1641_b1 );
not ( \1641_b1 , w_3504 );
and ( \1775_b0 , \1622_b0 , w_3505 );
and ( w_3504 , w_3505 , \1641_b0 );
or ( \1776_b1 , \1774_b1 , w_3507 );
not ( w_3507 , w_3508 );
and ( \1776_b0 , \1774_b0 , w_3509 );
and ( w_3508 ,  , w_3509 );
buf ( w_3507 , \1775_b1 );
not ( w_3507 , w_3510 );
not (  , w_3511 );
and ( w_3510 , w_3511 , \1775_b0 );
or ( \1777_b1 , \1776_b1 , w_3512 );
xor ( \1777_b0 , \1776_b0 , w_3514 );
not ( w_3514 , w_3515 );
and ( w_3515 , w_3512 , w_3513 );
buf ( w_3512 , \1649_b1 );
not ( w_3512 , w_3516 );
not ( w_3513 , w_3517 );
and ( w_3516 , w_3517 , \1649_b0 );
or ( \1778_b1 , \1773_b1 , \1777_b1 );
xor ( \1778_b0 , \1773_b0 , w_3518 );
not ( w_3518 , w_3519 );
and ( w_3519 , \1777_b1 , \1777_b0 );
or ( \1779_b1 , \1540_b1 , \1524_b1 );
not ( \1524_b1 , w_3520 );
and ( \1779_b0 , \1540_b0 , w_3521 );
and ( w_3520 , w_3521 , \1524_b0 );
or ( \1780_b1 , \1517_b1 , \1522_b1 );
not ( \1522_b1 , w_3522 );
and ( \1780_b0 , \1517_b0 , w_3523 );
and ( w_3522 , w_3523 , \1522_b0 );
or ( \1781_b1 , \1779_b1 , w_3525 );
not ( w_3525 , w_3526 );
and ( \1781_b0 , \1779_b0 , w_3527 );
and ( w_3526 ,  , w_3527 );
buf ( w_3525 , \1780_b1 );
not ( w_3525 , w_3528 );
not (  , w_3529 );
and ( w_3528 , w_3529 , \1780_b0 );
or ( \1782_b1 , \1781_b1 , w_3530 );
xor ( \1782_b0 , \1781_b0 , w_3532 );
not ( w_3532 , w_3533 );
and ( w_3533 , w_3530 , w_3531 );
buf ( w_3530 , \1531_b1 );
not ( w_3530 , w_3534 );
not ( w_3531 , w_3535 );
and ( w_3534 , w_3535 , \1531_b0 );
or ( \1783_b1 , \1778_b1 , \1782_b1 );
xor ( \1783_b0 , \1778_b0 , w_3536 );
not ( w_3536 , w_3537 );
and ( w_3537 , \1782_b1 , \1782_b0 );
or ( \1784_b1 , \1769_b1 , \1783_b1 );
not ( \1783_b1 , w_3538 );
and ( \1784_b0 , \1769_b0 , w_3539 );
and ( w_3538 , w_3539 , \1783_b0 );
or ( \1785_b1 , \1489_b1 , \1336_b1 );
not ( \1336_b1 , w_3540 );
and ( \1785_b0 , \1489_b0 , w_3541 );
and ( w_3540 , w_3541 , \1336_b0 );
or ( \1786_b1 , \1331_b1 , \1333_b1 );
not ( \1333_b1 , w_3542 );
and ( \1786_b0 , \1331_b0 , w_3543 );
and ( w_3542 , w_3543 , \1333_b0 );
or ( \1787_b1 , \1785_b1 , w_3545 );
not ( w_3545 , w_3546 );
and ( \1787_b0 , \1785_b0 , w_3547 );
and ( w_3546 ,  , w_3547 );
buf ( w_3545 , \1786_b1 );
not ( w_3545 , w_3548 );
not (  , w_3549 );
and ( w_3548 , w_3549 , \1786_b0 );
or ( \1788_b1 , \1787_b1 , w_3550 );
xor ( \1788_b0 , \1787_b0 , w_3552 );
not ( w_3552 , w_3553 );
and ( w_3553 , w_3550 , w_3551 );
buf ( w_3550 , \1332_b1 );
not ( w_3550 , w_3554 );
not ( w_3551 , w_3555 );
and ( w_3554 , w_3555 , \1332_b0 );
or ( \1789_b1 , \1384_b1 , \1349_b1 );
not ( \1349_b1 , w_3556 );
and ( \1789_b0 , \1384_b0 , w_3557 );
and ( w_3556 , w_3557 , \1349_b0 );
or ( \1790_b1 , \1342_b1 , \1347_b1 );
not ( \1347_b1 , w_3558 );
and ( \1790_b0 , \1342_b0 , w_3559 );
and ( w_3558 , w_3559 , \1347_b0 );
or ( \1791_b1 , \1789_b1 , w_3561 );
not ( w_3561 , w_3562 );
and ( \1791_b0 , \1789_b0 , w_3563 );
and ( w_3562 ,  , w_3563 );
buf ( w_3561 , \1790_b1 );
not ( w_3561 , w_3564 );
not (  , w_3565 );
and ( w_3564 , w_3565 , \1790_b0 );
or ( \1792_b1 , \1791_b1 , w_3566 );
xor ( \1792_b0 , \1791_b0 , w_3568 );
not ( w_3568 , w_3569 );
and ( w_3569 , w_3566 , w_3567 );
buf ( w_3566 , \1356_b1 );
not ( w_3566 , w_3570 );
not ( w_3567 , w_3571 );
and ( w_3570 , w_3571 , \1356_b0 );
or ( \1793_b1 , \1788_b1 , \1792_b1 );
not ( \1792_b1 , w_3572 );
and ( \1793_b0 , \1788_b0 , w_3573 );
and ( w_3572 , w_3573 , \1792_b0 );
buf ( \1794_b1 , \1754_b1 );
not ( \1794_b1 , w_3574 );
not ( \1794_b0 , w_3575 );
and ( w_3574 , w_3575 , \1754_b0 );
or ( \1795_b1 , \1794_b1 , \1545_b1 );
not ( \1545_b1 , w_3576 );
and ( \1795_b0 , \1794_b0 , w_3577 );
and ( w_3576 , w_3577 , \1545_b0 );
or ( \1796_b1 , \1792_b1 , \1795_b1 );
not ( \1795_b1 , w_3578 );
and ( \1796_b0 , \1792_b0 , w_3579 );
and ( w_3578 , w_3579 , \1795_b0 );
or ( \1797_b1 , \1788_b1 , \1795_b1 );
not ( \1795_b1 , w_3580 );
and ( \1797_b0 , \1788_b0 , w_3581 );
and ( w_3580 , w_3581 , \1795_b0 );
or ( \1799_b1 , \1553_b1 , \1538_b1 );
not ( \1538_b1 , w_3582 );
and ( \1799_b0 , \1553_b0 , w_3583 );
and ( w_3582 , w_3583 , \1538_b0 );
or ( \1800_b1 , \1533_b1 , \1536_b1 );
not ( \1536_b1 , w_3584 );
and ( \1800_b0 , \1533_b0 , w_3585 );
and ( w_3584 , w_3585 , \1536_b0 );
or ( \1801_b1 , \1799_b1 , w_3587 );
not ( w_3587 , w_3588 );
and ( \1801_b0 , \1799_b0 , w_3589 );
and ( w_3588 ,  , w_3589 );
buf ( w_3587 , \1800_b1 );
not ( w_3587 , w_3590 );
not (  , w_3591 );
and ( w_3590 , w_3591 , \1800_b0 );
or ( \1802_b1 , \1801_b1 , w_3592 );
xor ( \1802_b0 , \1801_b0 , w_3594 );
not ( w_3594 , w_3595 );
and ( w_3595 , w_3592 , w_3593 );
buf ( w_3592 , \1545_b1 );
not ( w_3592 , w_3596 );
not ( w_3593 , w_3597 );
and ( w_3596 , w_3597 , \1545_b0 );
or ( \1803_b1 , \1798_b1 , \1802_b1 );
xor ( \1803_b0 , \1798_b0 , w_3598 );
not ( w_3598 , w_3599 );
and ( w_3599 , \1802_b1 , \1802_b0 );
or ( \1804_b1 , \1492_b1 , \1496_b1 );
xor ( \1804_b0 , \1492_b0 , w_3600 );
not ( w_3600 , w_3601 );
and ( w_3601 , \1496_b1 , \1496_b0 );
or ( \1805_b1 , \1804_b1 , \1502_b1 );
xor ( \1805_b0 , \1804_b0 , w_3602 );
not ( w_3602 , w_3603 );
and ( w_3603 , \1502_b1 , \1502_b0 );
or ( \1806_b1 , \1803_b1 , \1805_b1 );
xor ( \1806_b0 , \1803_b0 , w_3604 );
not ( w_3604 , w_3605 );
and ( w_3605 , \1805_b1 , \1805_b0 );
or ( \1807_b1 , \1783_b1 , \1806_b1 );
not ( \1806_b1 , w_3606 );
and ( \1807_b0 , \1783_b0 , w_3607 );
and ( w_3606 , w_3607 , \1806_b0 );
or ( \1808_b1 , \1769_b1 , \1806_b1 );
not ( \1806_b1 , w_3608 );
and ( \1808_b0 , \1769_b0 , w_3609 );
and ( w_3608 , w_3609 , \1806_b0 );
or ( \1810_b1 , \1744_b1 , \1809_b1 );
not ( \1809_b1 , w_3610 );
and ( \1810_b0 , \1744_b0 , w_3611 );
and ( w_3610 , w_3611 , \1809_b0 );
or ( \1811_b1 , \1773_b1 , \1777_b1 );
not ( \1777_b1 , w_3612 );
and ( \1811_b0 , \1773_b0 , w_3613 );
and ( w_3612 , w_3613 , \1777_b0 );
or ( \1812_b1 , \1777_b1 , \1782_b1 );
not ( \1782_b1 , w_3614 );
and ( \1812_b0 , \1777_b0 , w_3615 );
and ( w_3614 , w_3615 , \1782_b0 );
or ( \1813_b1 , \1773_b1 , \1782_b1 );
not ( \1782_b1 , w_3616 );
and ( \1813_b0 , \1773_b0 , w_3617 );
and ( w_3616 , w_3617 , \1782_b0 );
or ( \1815_b1 , \1453_b1 , \1468_b1 );
not ( \1468_b1 , w_3618 );
and ( \1815_b0 , \1453_b0 , w_3619 );
and ( w_3618 , w_3619 , \1468_b0 );
or ( \1816_b1 , \1468_b1 , \1483_b1 );
not ( \1483_b1 , w_3620 );
and ( \1816_b0 , \1468_b0 , w_3621 );
and ( w_3620 , w_3621 , \1483_b0 );
or ( \1817_b1 , \1453_b1 , \1483_b1 );
not ( \1483_b1 , w_3622 );
and ( \1817_b0 , \1453_b0 , w_3623 );
and ( w_3622 , w_3623 , \1483_b0 );
or ( \1819_b1 , \1814_b1 , \1818_b1 );
xor ( \1819_b0 , \1814_b0 , w_3624 );
not ( w_3624 , w_3625 );
and ( w_3625 , \1818_b1 , \1818_b0 );
or ( \1820_b1 , \1338_b1 , \1336_b1 );
not ( \1336_b1 , w_3626 );
and ( \1820_b0 , \1338_b0 , w_3627 );
and ( w_3626 , w_3627 , \1336_b0 );
buf ( \1821_b1 , \1183_A[29]_b1 );
buf ( \1821_b0 , \1183_A[29]_b0 );
or ( \1822_b1 , \1821_b1 , \1333_b1 );
not ( \1333_b1 , w_3628 );
and ( \1822_b0 , \1821_b0 , w_3629 );
and ( w_3628 , w_3629 , \1333_b0 );
or ( \1823_b1 , \1820_b1 , w_3631 );
not ( w_3631 , w_3632 );
and ( \1823_b0 , \1820_b0 , w_3633 );
and ( w_3632 ,  , w_3633 );
buf ( w_3631 , \1822_b1 );
not ( w_3631 , w_3634 );
not (  , w_3635 );
and ( w_3634 , w_3635 , \1822_b0 );
or ( \1824_b1 , \1823_b1 , w_3636 );
xor ( \1824_b0 , \1823_b0 , w_3638 );
not ( w_3638 , w_3639 );
and ( w_3639 , w_3636 , w_3637 );
buf ( w_3636 , \1332_b1 );
not ( w_3636 , w_3640 );
not ( w_3637 , w_3641 );
and ( w_3640 , w_3641 , \1332_b0 );
or ( \1825_b1 , \1425_b1 , \1444_b1 );
not ( \1444_b1 , w_3642 );
and ( \1825_b0 , \1425_b0 , w_3643 );
and ( w_3642 , w_3643 , \1444_b0 );
or ( \1826_b1 , \1433_b1 , \1442_b1 );
not ( \1442_b1 , w_3644 );
and ( \1826_b0 , \1433_b0 , w_3645 );
and ( w_3644 , w_3645 , \1442_b0 );
or ( \1827_b1 , \1825_b1 , w_3647 );
not ( w_3647 , w_3648 );
and ( \1827_b0 , \1825_b0 , w_3649 );
and ( w_3648 ,  , w_3649 );
buf ( w_3647 , \1826_b1 );
not ( w_3647 , w_3650 );
not (  , w_3651 );
and ( w_3650 , w_3651 , \1826_b0 );
or ( \1828_b1 , \1827_b1 , w_3652 );
xor ( \1828_b0 , \1827_b0 , w_3654 );
not ( w_3654 , w_3655 );
and ( w_3655 , w_3652 , w_3653 );
buf ( w_3652 , \1451_b1 );
not ( w_3652 , w_3656 );
not ( w_3653 , w_3657 );
and ( w_3656 , w_3657 , \1451_b0 );
or ( \1829_b1 , \1824_b1 , \1828_b1 );
xor ( \1829_b0 , \1824_b0 , w_3658 );
not ( w_3658 , w_3659 );
and ( w_3659 , \1828_b1 , \1828_b0 );
or ( \1830_b1 , \1351_b1 , \1349_b1 );
not ( \1349_b1 , w_3660 );
and ( \1830_b0 , \1351_b0 , w_3661 );
and ( w_3660 , w_3661 , \1349_b0 );
or ( \1831_b1 , \1446_b1 , \1347_b1 );
not ( \1347_b1 , w_3662 );
and ( \1831_b0 , \1446_b0 , w_3663 );
and ( w_3662 , w_3663 , \1347_b0 );
or ( \1832_b1 , \1830_b1 , w_3665 );
not ( w_3665 , w_3666 );
and ( \1832_b0 , \1830_b0 , w_3667 );
and ( w_3666 ,  , w_3667 );
buf ( w_3665 , \1831_b1 );
not ( w_3665 , w_3668 );
not (  , w_3669 );
and ( w_3668 , w_3669 , \1831_b0 );
or ( \1833_b1 , \1832_b1 , w_3670 );
xor ( \1833_b0 , \1832_b0 , w_3672 );
not ( w_3672 , w_3673 );
and ( w_3673 , w_3670 , w_3671 );
buf ( w_3670 , \1356_b1 );
not ( w_3670 , w_3674 );
not ( w_3671 , w_3675 );
and ( w_3674 , w_3675 , \1356_b0 );
or ( \1834_b1 , \1829_b1 , \1833_b1 );
xor ( \1834_b0 , \1829_b0 , w_3676 );
not ( w_3676 , w_3677 );
and ( w_3677 , \1833_b1 , \1833_b0 );
or ( \1835_b1 , \1819_b1 , \1834_b1 );
xor ( \1835_b0 , \1819_b0 , w_3678 );
not ( w_3678 , w_3679 );
and ( w_3679 , \1834_b1 , \1834_b0 );
or ( \1836_b1 , \1809_b1 , \1835_b1 );
not ( \1835_b1 , w_3680 );
and ( \1836_b0 , \1809_b0 , w_3681 );
and ( w_3680 , w_3681 , \1835_b0 );
or ( \1837_b1 , \1744_b1 , \1835_b1 );
not ( \1835_b1 , w_3682 );
and ( \1837_b0 , \1744_b0 , w_3683 );
and ( w_3682 , w_3683 , \1835_b0 );
or ( \1839_b1 , \1594_b1 , \1838_b1 );
not ( \1838_b1 , w_3684 );
and ( \1839_b0 , \1594_b0 , w_3685 );
and ( w_3684 , w_3685 , \1838_b0 );
or ( \1840_b1 , \1560_b1 , \1574_b1 );
not ( \1574_b1 , w_3686 );
and ( \1840_b0 , \1560_b0 , w_3687 );
and ( w_3686 , w_3687 , \1574_b0 );
or ( \1841_b1 , \1574_b1 , \1590_b1 );
not ( \1590_b1 , w_3688 );
and ( \1841_b0 , \1574_b0 , w_3689 );
and ( w_3688 , w_3689 , \1590_b0 );
or ( \1842_b1 , \1560_b1 , \1590_b1 );
not ( \1590_b1 , w_3690 );
and ( \1842_b0 , \1560_b0 , w_3691 );
and ( w_3690 , w_3691 , \1590_b0 );
or ( \1844_b1 , \1814_b1 , \1818_b1 );
not ( \1818_b1 , w_3692 );
and ( \1844_b0 , \1814_b0 , w_3693 );
and ( w_3692 , w_3693 , \1818_b0 );
or ( \1845_b1 , \1818_b1 , \1834_b1 );
not ( \1834_b1 , w_3694 );
and ( \1845_b0 , \1818_b0 , w_3695 );
and ( w_3694 , w_3695 , \1834_b0 );
or ( \1846_b1 , \1814_b1 , \1834_b1 );
not ( \1834_b1 , w_3696 );
and ( \1846_b0 , \1814_b0 , w_3697 );
and ( w_3696 , w_3697 , \1834_b0 );
or ( \1848_b1 , \1843_b1 , \1847_b1 );
xor ( \1848_b0 , \1843_b0 , w_3698 );
not ( w_3698 , w_3699 );
and ( w_3699 , \1847_b1 , \1847_b0 );
or ( \1849_b1 , \1489_b1 , \1431_b1 );
not ( \1431_b1 , w_3700 );
and ( \1849_b0 , \1489_b0 , w_3701 );
and ( w_3700 , w_3701 , \1431_b0 );
or ( \1850_b1 , \1331_b1 , \1429_b1 );
not ( \1429_b1 , w_3702 );
and ( \1850_b0 , \1331_b0 , w_3703 );
and ( w_3702 , w_3703 , \1429_b0 );
or ( \1851_b1 , \1849_b1 , w_3705 );
not ( w_3705 , w_3706 );
and ( \1851_b0 , \1849_b0 , w_3707 );
and ( w_3706 ,  , w_3707 );
buf ( w_3705 , \1850_b1 );
not ( w_3705 , w_3708 );
not (  , w_3709 );
and ( w_3708 , w_3709 , \1850_b0 );
or ( \1852_b1 , \1851_b1 , w_3710 );
xor ( \1852_b0 , \1851_b0 , w_3712 );
not ( w_3712 , w_3713 );
and ( w_3713 , w_3710 , w_3711 );
buf ( w_3710 , \1438_b1 );
not ( w_3710 , w_3714 );
not ( w_3711 , w_3715 );
and ( w_3714 , w_3715 , \1438_b0 );
buf ( \1853_b1 , \1502_b1 );
not ( \1853_b1 , w_3716 );
not ( \1853_b0 , w_3717 );
and ( w_3716 , w_3717 , \1502_b0 );
or ( \1854_b1 , \1853_b1 , \1558_b1 );
not ( \1558_b1 , w_3718 );
and ( \1854_b0 , \1853_b0 , w_3719 );
and ( w_3718 , w_3719 , \1558_b0 );
or ( \1855_b1 , \1852_b1 , \1854_b1 );
xor ( \1855_b0 , \1852_b0 , w_3720 );
not ( w_3720 , w_3721 );
and ( w_3721 , \1854_b1 , \1854_b0 );
or ( \1856_b1 , \1616_b1 , \1675_b1 );
not ( \1675_b1 , w_3722 );
and ( \1856_b0 , \1616_b0 , w_3723 );
and ( w_3722 , w_3723 , \1675_b0 );
or ( \1857_b1 , \1391_b1 , \1673_b1 );
not ( \1673_b1 , w_3724 );
and ( \1857_b0 , \1391_b0 , w_3725 );
and ( w_3724 , w_3725 , \1673_b0 );
or ( \1858_b1 , \1856_b1 , w_3727 );
not ( w_3727 , w_3728 );
and ( \1858_b0 , \1856_b0 , w_3729 );
and ( w_3728 ,  , w_3729 );
buf ( w_3727 , \1857_b1 );
not ( w_3727 , w_3730 );
not (  , w_3731 );
and ( w_3730 , w_3731 , \1857_b0 );
or ( \1859_b1 , \1858_b1 , w_3732 );
xor ( \1859_b0 , \1858_b0 , w_3734 );
not ( w_3734 , w_3735 );
and ( w_3735 , w_3732 , w_3733 );
buf ( w_3732 , \1681_b1 );
not ( w_3732 , w_3736 );
not ( w_3733 , w_3737 );
and ( w_3736 , w_3737 , \1681_b0 );
or ( \1860_b1 , \1855_b1 , \1859_b1 );
not ( \1859_b1 , w_3738 );
and ( \1860_b0 , \1855_b0 , w_3739 );
and ( w_3738 , w_3739 , \1859_b0 );
or ( \1861_b1 , \1622_b1 , \1643_b1 );
not ( \1643_b1 , w_3740 );
and ( \1861_b0 , \1622_b0 , w_3741 );
and ( w_3740 , w_3741 , \1643_b0 );
or ( \1862_b1 , \1407_b1 , \1641_b1 );
not ( \1641_b1 , w_3742 );
and ( \1862_b0 , \1407_b0 , w_3743 );
and ( w_3742 , w_3743 , \1641_b0 );
or ( \1863_b1 , \1861_b1 , w_3745 );
not ( w_3745 , w_3746 );
and ( \1863_b0 , \1861_b0 , w_3747 );
and ( w_3746 ,  , w_3747 );
buf ( w_3745 , \1862_b1 );
not ( w_3745 , w_3748 );
not (  , w_3749 );
and ( w_3748 , w_3749 , \1862_b0 );
or ( \1864_b1 , \1863_b1 , w_3750 );
xor ( \1864_b0 , \1863_b0 , w_3752 );
not ( w_3752 , w_3753 );
and ( w_3753 , w_3750 , w_3751 );
buf ( w_3750 , \1649_b1 );
not ( w_3750 , w_3754 );
not ( w_3751 , w_3755 );
and ( w_3754 , w_3755 , \1649_b0 );
or ( \1865_b1 , \1859_b1 , \1864_b1 );
not ( \1864_b1 , w_3756 );
and ( \1865_b0 , \1859_b0 , w_3757 );
and ( w_3756 , w_3757 , \1864_b0 );
or ( \1866_b1 , \1855_b1 , \1864_b1 );
not ( \1864_b1 , w_3758 );
and ( \1866_b0 , \1855_b0 , w_3759 );
and ( w_3758 , w_3759 , \1864_b0 );
or ( \1868_b1 , \1342_b1 , \1382_b1 );
not ( \1382_b1 , w_3760 );
and ( \1868_b0 , \1342_b0 , w_3761 );
and ( w_3760 , w_3761 , \1382_b0 );
or ( \1869_b1 , \1351_b1 , \1380_b1 );
not ( \1380_b1 , w_3762 );
and ( \1869_b0 , \1351_b0 , w_3763 );
and ( w_3762 , w_3763 , \1380_b0 );
or ( \1870_b1 , \1868_b1 , w_3765 );
not ( w_3765 , w_3766 );
and ( \1870_b0 , \1868_b0 , w_3767 );
and ( w_3766 ,  , w_3767 );
buf ( w_3765 , \1869_b1 );
not ( w_3765 , w_3768 );
not (  , w_3769 );
and ( w_3768 , w_3769 , \1869_b0 );
or ( \1871_b1 , \1870_b1 , w_3770 );
xor ( \1871_b0 , \1870_b0 , w_3772 );
not ( w_3772 , w_3773 );
and ( w_3773 , w_3770 , w_3771 );
buf ( w_3770 , \1389_b1 );
not ( w_3770 , w_3774 );
not ( w_3771 , w_3775 );
and ( w_3774 , w_3775 , \1389_b0 );
or ( \1872_b1 , \1359_b1 , \1397_b1 );
not ( \1397_b1 , w_3776 );
and ( \1872_b0 , \1359_b0 , w_3777 );
and ( w_3776 , w_3777 , \1397_b0 );
or ( \1873_b1 , \1368_b1 , \1395_b1 );
not ( \1395_b1 , w_3778 );
and ( \1873_b0 , \1368_b0 , w_3779 );
and ( w_3778 , w_3779 , \1395_b0 );
or ( \1874_b1 , \1872_b1 , w_3781 );
not ( w_3781 , w_3782 );
and ( \1874_b0 , \1872_b0 , w_3783 );
and ( w_3782 ,  , w_3783 );
buf ( w_3781 , \1873_b1 );
not ( w_3781 , w_3784 );
not (  , w_3785 );
and ( w_3784 , w_3785 , \1873_b0 );
or ( \1875_b1 , \1874_b1 , w_3786 );
xor ( \1875_b0 , \1874_b0 , w_3788 );
not ( w_3788 , w_3789 );
and ( w_3789 , w_3786 , w_3787 );
buf ( w_3786 , \1404_b1 );
not ( w_3786 , w_3790 );
not ( w_3787 , w_3791 );
and ( w_3790 , w_3791 , \1404_b0 );
or ( \1876_b1 , \1871_b1 , \1875_b1 );
xor ( \1876_b0 , \1871_b0 , w_3792 );
not ( w_3792 , w_3793 );
and ( w_3793 , \1875_b1 , \1875_b0 );
or ( \1877_b1 , \1586_b1 , \1414_b1 );
not ( \1414_b1 , w_3794 );
and ( \1877_b0 , \1586_b0 , w_3795 );
and ( w_3794 , w_3795 , \1414_b0 );
or ( \1878_b1 , \1616_b1 , \1412_b1 );
not ( \1412_b1 , w_3796 );
and ( \1878_b0 , \1616_b0 , w_3797 );
and ( w_3796 , w_3797 , \1412_b0 );
or ( \1879_b1 , \1877_b1 , w_3799 );
not ( w_3799 , w_3800 );
and ( \1879_b0 , \1877_b0 , w_3801 );
and ( w_3800 ,  , w_3801 );
buf ( w_3799 , \1878_b1 );
not ( w_3799 , w_3802 );
not (  , w_3803 );
and ( w_3802 , w_3803 , \1878_b0 );
or ( \1880_b1 , \1879_b1 , w_3804 );
xor ( \1880_b0 , \1879_b0 , w_3806 );
not ( w_3806 , w_3807 );
and ( w_3807 , w_3804 , w_3805 );
buf ( w_3804 , \1421_b1 );
not ( w_3804 , w_3808 );
not ( w_3805 , w_3809 );
and ( w_3808 , w_3809 , \1421_b0 );
or ( \1881_b1 , \1876_b1 , \1880_b1 );
xor ( \1881_b0 , \1876_b0 , w_3810 );
not ( w_3810 , w_3811 );
and ( w_3811 , \1880_b1 , \1880_b0 );
or ( \1882_b1 , \1867_b1 , \1881_b1 );
xor ( \1882_b0 , \1867_b0 , w_3812 );
not ( w_3812 , w_3813 );
and ( w_3813 , \1881_b1 , \1881_b0 );
or ( \1883_b1 , \1391_b1 , \1675_b1 );
not ( \1675_b1 , w_3814 );
and ( \1883_b0 , \1391_b0 , w_3815 );
and ( w_3814 , w_3815 , \1675_b0 );
or ( \1884_b1 , \1399_b1 , \1673_b1 );
not ( \1673_b1 , w_3816 );
and ( \1884_b0 , \1399_b0 , w_3817 );
and ( w_3816 , w_3817 , \1673_b0 );
or ( \1885_b1 , \1883_b1 , w_3819 );
not ( w_3819 , w_3820 );
and ( \1885_b0 , \1883_b0 , w_3821 );
and ( w_3820 ,  , w_3821 );
buf ( w_3819 , \1884_b1 );
not ( w_3819 , w_3822 );
not (  , w_3823 );
and ( w_3822 , w_3823 , \1884_b0 );
or ( \1886_b1 , \1885_b1 , w_3824 );
xor ( \1886_b0 , \1885_b0 , w_3826 );
not ( w_3826 , w_3827 );
and ( w_3827 , w_3824 , w_3825 );
buf ( w_3824 , \1681_b1 );
not ( w_3824 , w_3828 );
not ( w_3825 , w_3829 );
and ( w_3828 , w_3829 , \1681_b0 );
or ( \1887_b1 , \1407_b1 , \1643_b1 );
not ( \1643_b1 , w_3830 );
and ( \1887_b0 , \1407_b0 , w_3831 );
and ( w_3830 , w_3831 , \1643_b0 );
or ( \1888_b1 , \1416_b1 , \1641_b1 );
not ( \1641_b1 , w_3832 );
and ( \1888_b0 , \1416_b0 , w_3833 );
and ( w_3832 , w_3833 , \1641_b0 );
or ( \1889_b1 , \1887_b1 , w_3835 );
not ( w_3835 , w_3836 );
and ( \1889_b0 , \1887_b0 , w_3837 );
and ( w_3836 ,  , w_3837 );
buf ( w_3835 , \1888_b1 );
not ( w_3835 , w_3838 );
not (  , w_3839 );
and ( w_3838 , w_3839 , \1888_b0 );
or ( \1890_b1 , \1889_b1 , w_3840 );
xor ( \1890_b0 , \1889_b0 , w_3842 );
not ( w_3842 , w_3843 );
and ( w_3843 , w_3840 , w_3841 );
buf ( w_3840 , \1649_b1 );
not ( w_3840 , w_3844 );
not ( w_3841 , w_3845 );
and ( w_3844 , w_3845 , \1649_b0 );
or ( \1891_b1 , \1886_b1 , \1890_b1 );
xor ( \1891_b0 , \1886_b0 , w_3846 );
not ( w_3846 , w_3847 );
and ( w_3847 , \1890_b1 , \1890_b0 );
or ( \1892_b1 , \1526_b1 , \1524_b1 );
not ( \1524_b1 , w_3848 );
and ( \1892_b0 , \1526_b0 , w_3849 );
and ( w_3848 , w_3849 , \1524_b0 );
or ( \1893_b1 , \1622_b1 , \1522_b1 );
not ( \1522_b1 , w_3850 );
and ( \1893_b0 , \1622_b0 , w_3851 );
and ( w_3850 , w_3851 , \1522_b0 );
or ( \1894_b1 , \1892_b1 , w_3853 );
not ( w_3853 , w_3854 );
and ( \1894_b0 , \1892_b0 , w_3855 );
and ( w_3854 ,  , w_3855 );
buf ( w_3853 , \1893_b1 );
not ( w_3853 , w_3856 );
not (  , w_3857 );
and ( w_3856 , w_3857 , \1893_b0 );
or ( \1895_b1 , \1894_b1 , w_3858 );
xor ( \1895_b0 , \1894_b0 , w_3860 );
not ( w_3860 , w_3861 );
and ( w_3861 , w_3858 , w_3859 );
buf ( w_3858 , \1531_b1 );
not ( w_3858 , w_3862 );
not ( w_3859 , w_3863 );
and ( w_3862 , w_3863 , \1531_b0 );
or ( \1896_b1 , \1891_b1 , \1895_b1 );
xor ( \1896_b0 , \1891_b0 , w_3864 );
not ( w_3864 , w_3865 );
and ( w_3865 , \1895_b1 , \1895_b0 );
or ( \1897_b1 , \1882_b1 , \1896_b1 );
xor ( \1897_b0 , \1882_b0 , w_3866 );
not ( w_3866 , w_3867 );
and ( w_3867 , \1896_b1 , \1896_b0 );
or ( \1898_b1 , \1848_b1 , \1897_b1 );
xor ( \1898_b0 , \1848_b0 , w_3868 );
not ( w_3868 , w_3869 );
and ( w_3869 , \1897_b1 , \1897_b0 );
or ( \1899_b1 , \1838_b1 , \1898_b1 );
not ( \1898_b1 , w_3870 );
and ( \1899_b0 , \1838_b0 , w_3871 );
and ( w_3870 , w_3871 , \1898_b0 );
or ( \1900_b1 , \1594_b1 , \1898_b1 );
not ( \1898_b1 , w_3872 );
and ( \1900_b0 , \1594_b0 , w_3873 );
and ( w_3872 , w_3873 , \1898_b0 );
or ( \1902_b1 , \1788_b1 , \1792_b1 );
xor ( \1902_b0 , \1788_b0 , w_3874 );
not ( w_3874 , w_3875 );
and ( w_3875 , \1792_b1 , \1792_b0 );
or ( \1903_b1 , \1902_b1 , \1795_b1 );
xor ( \1903_b0 , \1902_b0 , w_3876 );
not ( w_3876 , w_3877 );
and ( w_3877 , \1795_b1 , \1795_b0 );
or ( \1904_b1 , \1757_b1 , \1761_b1 );
xor ( \1904_b0 , \1757_b0 , w_3878 );
not ( w_3878 , w_3879 );
and ( w_3879 , \1761_b1 , \1761_b0 );
or ( \1905_b1 , \1904_b1 , \1766_b1 );
xor ( \1905_b0 , \1904_b0 , w_3880 );
not ( w_3880 , w_3881 );
and ( w_3881 , \1766_b1 , \1766_b0 );
or ( \1906_b1 , \1903_b1 , \1905_b1 );
not ( \1905_b1 , w_3882 );
and ( \1906_b0 , \1903_b0 , w_3883 );
and ( w_3882 , w_3883 , \1905_b0 );
or ( \1907_b1 , \1728_b1 , \1732_b1 );
xor ( \1907_b0 , \1728_b0 , w_3884 );
not ( w_3884 , w_3885 );
and ( w_3885 , \1732_b1 , \1732_b0 );
or ( \1908_b1 , \1907_b1 , \1737_b1 );
xor ( \1908_b0 , \1907_b0 , w_3886 );
not ( w_3886 , w_3887 );
and ( w_3887 , \1737_b1 , \1737_b0 );
or ( \1909_b1 , \1905_b1 , \1908_b1 );
not ( \1908_b1 , w_3888 );
and ( \1909_b0 , \1905_b0 , w_3889 );
and ( w_3888 , w_3889 , \1908_b0 );
or ( \1910_b1 , \1903_b1 , \1908_b1 );
not ( \1908_b1 , w_3890 );
and ( \1910_b0 , \1903_b0 , w_3891 );
and ( w_3890 , w_3891 , \1908_b0 );
or ( \1912_b1 , \1425_b1 , \1336_b1 );
not ( \1336_b1 , w_3892 );
and ( \1912_b0 , \1425_b0 , w_3893 );
and ( w_3892 , w_3893 , \1336_b0 );
or ( \1913_b1 , \1433_b1 , \1333_b1 );
not ( \1333_b1 , w_3894 );
and ( \1913_b0 , \1433_b0 , w_3895 );
and ( w_3894 , w_3895 , \1333_b0 );
or ( \1914_b1 , \1912_b1 , w_3897 );
not ( w_3897 , w_3898 );
and ( \1914_b0 , \1912_b0 , w_3899 );
and ( w_3898 ,  , w_3899 );
buf ( w_3897 , \1913_b1 );
not ( w_3897 , w_3900 );
not (  , w_3901 );
and ( w_3900 , w_3901 , \1913_b0 );
or ( \1915_b1 , \1914_b1 , w_3902 );
xor ( \1915_b0 , \1914_b0 , w_3904 );
not ( w_3904 , w_3905 );
and ( w_3905 , w_3902 , w_3903 );
buf ( w_3902 , \1332_b1 );
not ( w_3902 , w_3906 );
not ( w_3903 , w_3907 );
and ( w_3906 , w_3907 , \1332_b0 );
or ( \1916_b1 , \1462_b1 , \1349_b1 );
not ( \1349_b1 , w_3908 );
and ( \1916_b0 , \1462_b0 , w_3909 );
and ( w_3908 , w_3909 , \1349_b0 );
or ( \1917_b1 , \1376_b1 , \1347_b1 );
not ( \1347_b1 , w_3910 );
and ( \1917_b0 , \1376_b0 , w_3911 );
and ( w_3910 , w_3911 , \1347_b0 );
or ( \1918_b1 , \1916_b1 , w_3913 );
not ( w_3913 , w_3914 );
and ( \1918_b0 , \1916_b0 , w_3915 );
and ( w_3914 ,  , w_3915 );
buf ( w_3913 , \1917_b1 );
not ( w_3913 , w_3916 );
not (  , w_3917 );
and ( w_3916 , w_3917 , \1917_b0 );
or ( \1919_b1 , \1918_b1 , w_3918 );
xor ( \1919_b0 , \1918_b0 , w_3920 );
not ( w_3920 , w_3921 );
and ( w_3921 , w_3918 , w_3919 );
buf ( w_3918 , \1356_b1 );
not ( w_3918 , w_3922 );
not ( w_3919 , w_3923 );
and ( w_3922 , w_3923 , \1356_b0 );
or ( \1920_b1 , \1915_b1 , \1919_b1 );
not ( \1919_b1 , w_3924 );
and ( \1920_b0 , \1915_b0 , w_3925 );
and ( w_3924 , w_3925 , \1919_b0 );
or ( \1921_b1 , \1498_b1 , \1522_b1 );
not ( \1522_b1 , w_3926 );
and ( \1921_b0 , \1498_b0 , w_3927 );
and ( w_3926 , w_3927 , \1522_b0 );
buf ( \1922_b1 , \1921_b1 );
not ( \1922_b1 , w_3928 );
not ( \1922_b0 , w_3929 );
and ( w_3928 , w_3929 , \1921_b0 );
or ( \1923_b1 , \1922_b1 , \1531_b1 );
not ( \1531_b1 , w_3930 );
and ( \1923_b0 , \1922_b0 , w_3931 );
and ( w_3930 , w_3931 , \1531_b0 );
or ( \1924_b1 , \1919_b1 , \1923_b1 );
not ( \1923_b1 , w_3932 );
and ( \1924_b0 , \1919_b0 , w_3933 );
and ( w_3932 , w_3933 , \1923_b0 );
or ( \1925_b1 , \1915_b1 , \1923_b1 );
not ( \1923_b1 , w_3934 );
and ( \1925_b0 , \1915_b0 , w_3935 );
and ( w_3934 , w_3935 , \1923_b0 );
or ( \1927_b1 , \1368_b1 , \1460_b1 );
not ( \1460_b1 , w_3936 );
and ( \1927_b0 , \1368_b0 , w_3937 );
and ( w_3936 , w_3937 , \1460_b0 );
or ( \1928_b1 , \1470_b1 , \1458_b1 );
not ( \1458_b1 , w_3938 );
and ( \1928_b0 , \1470_b0 , w_3939 );
and ( w_3938 , w_3939 , \1458_b0 );
or ( \1929_b1 , \1927_b1 , w_3941 );
not ( w_3941 , w_3942 );
and ( \1929_b0 , \1927_b0 , w_3943 );
and ( w_3942 ,  , w_3943 );
buf ( w_3941 , \1928_b1 );
not ( w_3941 , w_3944 );
not (  , w_3945 );
and ( w_3944 , w_3945 , \1928_b0 );
or ( \1930_b1 , \1929_b1 , w_3946 );
xor ( \1930_b0 , \1929_b0 , w_3948 );
not ( w_3948 , w_3949 );
and ( w_3949 , w_3946 , w_3947 );
buf ( w_3946 , \1467_b1 );
not ( w_3946 , w_3950 );
not ( w_3947 , w_3951 );
and ( w_3950 , w_3951 , \1467_b0 );
or ( \1931_b1 , \1399_b1 , \1475_b1 );
not ( \1475_b1 , w_3952 );
and ( \1931_b0 , \1399_b0 , w_3953 );
and ( w_3952 , w_3953 , \1475_b0 );
or ( \1932_b1 , \1359_b1 , \1473_b1 );
not ( \1473_b1 , w_3954 );
and ( \1932_b0 , \1359_b0 , w_3955 );
and ( w_3954 , w_3955 , \1473_b0 );
or ( \1933_b1 , \1931_b1 , w_3957 );
not ( w_3957 , w_3958 );
and ( \1933_b0 , \1931_b0 , w_3959 );
and ( w_3958 ,  , w_3959 );
buf ( w_3957 , \1932_b1 );
not ( w_3957 , w_3960 );
not (  , w_3961 );
and ( w_3960 , w_3961 , \1932_b0 );
or ( \1934_b1 , \1933_b1 , w_3962 );
xor ( \1934_b0 , \1933_b0 , w_3964 );
not ( w_3964 , w_3965 );
and ( w_3965 , w_3962 , w_3963 );
buf ( w_3962 , \1482_b1 );
not ( w_3962 , w_3966 );
not ( w_3963 , w_3967 );
and ( w_3966 , w_3967 , \1482_b0 );
or ( \1935_b1 , \1930_b1 , \1934_b1 );
not ( \1934_b1 , w_3968 );
and ( \1935_b0 , \1930_b0 , w_3969 );
and ( w_3968 , w_3969 , \1934_b0 );
or ( \1936_b1 , \1517_b1 , \1414_b1 );
not ( \1414_b1 , w_3970 );
and ( \1936_b0 , \1517_b0 , w_3971 );
and ( w_3970 , w_3971 , \1414_b0 );
or ( \1937_b1 , \1526_b1 , \1412_b1 );
not ( \1412_b1 , w_3972 );
and ( \1937_b0 , \1526_b0 , w_3973 );
and ( w_3972 , w_3973 , \1412_b0 );
or ( \1938_b1 , \1936_b1 , w_3975 );
not ( w_3975 , w_3976 );
and ( \1938_b0 , \1936_b0 , w_3977 );
and ( w_3976 ,  , w_3977 );
buf ( w_3975 , \1937_b1 );
not ( w_3975 , w_3978 );
not (  , w_3979 );
and ( w_3978 , w_3979 , \1937_b0 );
or ( \1939_b1 , \1938_b1 , w_3980 );
xor ( \1939_b0 , \1938_b0 , w_3982 );
not ( w_3982 , w_3983 );
and ( w_3983 , w_3980 , w_3981 );
buf ( w_3980 , \1421_b1 );
not ( w_3980 , w_3984 );
not ( w_3981 , w_3985 );
and ( w_3984 , w_3985 , \1421_b0 );
or ( \1940_b1 , \1934_b1 , \1939_b1 );
not ( \1939_b1 , w_3986 );
and ( \1940_b0 , \1934_b0 , w_3987 );
and ( w_3986 , w_3987 , \1939_b0 );
or ( \1941_b1 , \1930_b1 , \1939_b1 );
not ( \1939_b1 , w_3988 );
and ( \1941_b0 , \1930_b0 , w_3989 );
and ( w_3988 , w_3989 , \1939_b0 );
or ( \1943_b1 , \1926_b1 , \1942_b1 );
not ( \1942_b1 , w_3990 );
and ( \1943_b0 , \1926_b0 , w_3991 );
and ( w_3990 , w_3991 , \1942_b0 );
or ( \1944_b1 , \1477_b1 , \1382_b1 );
not ( \1382_b1 , w_3992 );
and ( \1944_b0 , \1477_b0 , w_3993 );
and ( w_3992 , w_3993 , \1382_b0 );
or ( \1945_b1 , \1454_b1 , \1380_b1 );
not ( \1380_b1 , w_3994 );
and ( \1945_b0 , \1454_b0 , w_3995 );
and ( w_3994 , w_3995 , \1380_b0 );
or ( \1946_b1 , \1944_b1 , w_3997 );
not ( w_3997 , w_3998 );
and ( \1946_b0 , \1944_b0 , w_3999 );
and ( w_3998 ,  , w_3999 );
buf ( w_3997 , \1945_b1 );
not ( w_3997 , w_4000 );
not (  , w_4001 );
and ( w_4000 , w_4001 , \1945_b0 );
or ( \1947_b1 , \1946_b1 , w_4002 );
xor ( \1947_b0 , \1946_b0 , w_4004 );
not ( w_4004 , w_4005 );
and ( w_4005 , w_4002 , w_4003 );
buf ( w_4002 , \1389_b1 );
not ( w_4002 , w_4006 );
not ( w_4003 , w_4007 );
and ( w_4006 , w_4007 , \1389_b0 );
or ( \1948_b1 , \1616_b1 , \1366_b1 );
not ( \1366_b1 , w_4008 );
and ( \1948_b0 , \1616_b0 , w_4009 );
and ( w_4008 , w_4009 , \1366_b0 );
or ( \1949_b1 , \1391_b1 , \1364_b1 );
not ( \1364_b1 , w_4010 );
and ( \1949_b0 , \1391_b0 , w_4011 );
and ( w_4010 , w_4011 , \1364_b0 );
or ( \1950_b1 , \1948_b1 , w_4013 );
not ( w_4013 , w_4014 );
and ( \1950_b0 , \1948_b0 , w_4015 );
and ( w_4014 ,  , w_4015 );
buf ( w_4013 , \1949_b1 );
not ( w_4013 , w_4016 );
not (  , w_4017 );
and ( w_4016 , w_4017 , \1949_b0 );
or ( \1951_b1 , \1950_b1 , w_4018 );
xor ( \1951_b0 , \1950_b0 , w_4020 );
not ( w_4020 , w_4021 );
and ( w_4021 , w_4018 , w_4019 );
buf ( w_4018 , \1373_b1 );
not ( w_4018 , w_4022 );
not ( w_4019 , w_4023 );
and ( w_4022 , w_4023 , \1373_b0 );
or ( \1952_b1 , \1947_b1 , \1951_b1 );
not ( \1951_b1 , w_4024 );
and ( \1952_b0 , \1947_b0 , w_4025 );
and ( w_4024 , w_4025 , \1951_b0 );
or ( \1953_b1 , \1416_b1 , \1397_b1 );
not ( \1397_b1 , w_4026 );
and ( \1953_b0 , \1416_b0 , w_4027 );
and ( w_4026 , w_4027 , \1397_b0 );
or ( \1954_b1 , \1586_b1 , \1395_b1 );
not ( \1395_b1 , w_4028 );
and ( \1954_b0 , \1586_b0 , w_4029 );
and ( w_4028 , w_4029 , \1395_b0 );
or ( \1955_b1 , \1953_b1 , w_4031 );
not ( w_4031 , w_4032 );
and ( \1955_b0 , \1953_b0 , w_4033 );
and ( w_4032 ,  , w_4033 );
buf ( w_4031 , \1954_b1 );
not ( w_4031 , w_4034 );
not (  , w_4035 );
and ( w_4034 , w_4035 , \1954_b0 );
or ( \1956_b1 , \1955_b1 , w_4036 );
xor ( \1956_b0 , \1955_b0 , w_4038 );
not ( w_4038 , w_4039 );
and ( w_4039 , w_4036 , w_4037 );
buf ( w_4036 , \1404_b1 );
not ( w_4036 , w_4040 );
not ( w_4037 , w_4041 );
and ( w_4040 , w_4041 , \1404_b0 );
or ( \1957_b1 , \1951_b1 , \1956_b1 );
not ( \1956_b1 , w_4042 );
and ( \1957_b0 , \1951_b0 , w_4043 );
and ( w_4042 , w_4043 , \1956_b0 );
or ( \1958_b1 , \1947_b1 , \1956_b1 );
not ( \1956_b1 , w_4044 );
and ( \1958_b0 , \1947_b0 , w_4045 );
and ( w_4044 , w_4045 , \1956_b0 );
or ( \1960_b1 , \1942_b1 , \1959_b1 );
not ( \1959_b1 , w_4046 );
and ( \1960_b0 , \1942_b0 , w_4047 );
and ( w_4046 , w_4047 , \1959_b0 );
or ( \1961_b1 , \1926_b1 , \1959_b1 );
not ( \1959_b1 , w_4048 );
and ( \1961_b0 , \1926_b0 , w_4049 );
and ( w_4048 , w_4049 , \1959_b0 );
or ( \1963_b1 , \1633_b1 , \1637_b1 );
xor ( \1963_b0 , \1633_b0 , w_4050 );
not ( w_4050 , w_4051 );
and ( w_4051 , \1637_b1 , \1637_b0 );
or ( \1964_b1 , \1622_b1 , \1675_b1 );
not ( \1675_b1 , w_4052 );
and ( \1964_b0 , \1622_b0 , w_4053 );
and ( w_4052 , w_4053 , \1675_b0 );
or ( \1965_b1 , \1407_b1 , \1673_b1 );
not ( \1673_b1 , w_4054 );
and ( \1965_b0 , \1407_b0 , w_4055 );
and ( w_4054 , w_4055 , \1673_b0 );
or ( \1966_b1 , \1964_b1 , w_4057 );
not ( w_4057 , w_4058 );
and ( \1966_b0 , \1964_b0 , w_4059 );
and ( w_4058 ,  , w_4059 );
buf ( w_4057 , \1965_b1 );
not ( w_4057 , w_4060 );
not (  , w_4061 );
and ( w_4060 , w_4061 , \1965_b0 );
or ( \1967_b1 , \1966_b1 , w_4062 );
xor ( \1967_b0 , \1966_b0 , w_4064 );
not ( w_4064 , w_4065 );
and ( w_4065 , w_4062 , w_4063 );
buf ( w_4062 , \1681_b1 );
not ( w_4062 , w_4066 );
not ( w_4063 , w_4067 );
and ( w_4066 , w_4067 , \1681_b0 );
or ( \1968_b1 , \1963_b1 , \1967_b1 );
not ( \1967_b1 , w_4068 );
and ( \1968_b0 , \1963_b0 , w_4069 );
and ( w_4068 , w_4069 , \1967_b0 );
or ( \1969_b1 , \1533_b1 , \1643_b1 );
not ( \1643_b1 , w_4070 );
and ( \1969_b0 , \1533_b0 , w_4071 );
and ( w_4070 , w_4071 , \1643_b0 );
or ( \1970_b1 , \1540_b1 , \1641_b1 );
not ( \1641_b1 , w_4072 );
and ( \1970_b0 , \1540_b0 , w_4073 );
and ( w_4072 , w_4073 , \1641_b0 );
or ( \1971_b1 , \1969_b1 , w_4075 );
not ( w_4075 , w_4076 );
and ( \1971_b0 , \1969_b0 , w_4077 );
and ( w_4076 ,  , w_4077 );
buf ( w_4075 , \1970_b1 );
not ( w_4075 , w_4078 );
not (  , w_4079 );
and ( w_4078 , w_4079 , \1970_b0 );
or ( \1972_b1 , \1971_b1 , w_4080 );
xor ( \1972_b0 , \1971_b0 , w_4082 );
not ( w_4082 , w_4083 );
and ( w_4083 , w_4080 , w_4081 );
buf ( w_4080 , \1649_b1 );
not ( w_4080 , w_4084 );
not ( w_4081 , w_4085 );
and ( w_4084 , w_4085 , \1649_b0 );
or ( \1973_b1 , \1967_b1 , \1972_b1 );
not ( \1972_b1 , w_4086 );
and ( \1973_b0 , \1967_b0 , w_4087 );
and ( w_4086 , w_4087 , \1972_b0 );
or ( \1974_b1 , \1963_b1 , \1972_b1 );
not ( \1972_b1 , w_4088 );
and ( \1974_b0 , \1963_b0 , w_4089 );
and ( w_4088 , w_4089 , \1972_b0 );
or ( \1976_b1 , \1748_b1 , \1752_b1 );
xor ( \1976_b0 , \1748_b0 , w_4090 );
not ( w_4090 , w_4091 );
and ( w_4091 , \1752_b1 , \1752_b0 );
or ( \1977_b1 , \1976_b1 , \1754_b1 );
xor ( \1977_b0 , \1976_b0 , w_4092 );
not ( w_4092 , w_4093 );
and ( w_4093 , \1754_b1 , \1754_b0 );
or ( \1978_b1 , \1975_b1 , \1977_b1 );
not ( \1977_b1 , w_4094 );
and ( \1978_b0 , \1975_b0 , w_4095 );
and ( w_4094 , w_4095 , \1977_b0 );
or ( \1979_b1 , \1598_b1 , \1602_b1 );
xor ( \1979_b0 , \1598_b0 , w_4096 );
not ( w_4096 , w_4097 );
and ( w_4097 , \1602_b1 , \1602_b0 );
or ( \1980_b1 , \1979_b1 , \1607_b1 );
xor ( \1980_b0 , \1979_b0 , w_4098 );
not ( w_4098 , w_4099 );
and ( w_4099 , \1607_b1 , \1607_b0 );
or ( \1981_b1 , \1977_b1 , \1980_b1 );
not ( \1980_b1 , w_4100 );
and ( \1981_b0 , \1977_b0 , w_4101 );
and ( w_4100 , w_4101 , \1980_b0 );
or ( \1982_b1 , \1975_b1 , \1980_b1 );
not ( \1980_b1 , w_4102 );
and ( \1982_b0 , \1975_b0 , w_4103 );
and ( w_4102 , w_4103 , \1980_b0 );
or ( \1984_b1 , \1962_b1 , \1983_b1 );
not ( \1983_b1 , w_4104 );
and ( \1984_b0 , \1962_b0 , w_4105 );
and ( w_4104 , w_4105 , \1983_b0 );
or ( \1985_b1 , \1610_b1 , \1628_b1 );
xor ( \1985_b0 , \1610_b0 , w_4106 );
not ( w_4106 , w_4107 );
and ( w_4107 , \1628_b1 , \1628_b0 );
or ( \1986_b1 , \1985_b1 , \1658_b1 );
xor ( \1986_b0 , \1985_b0 , w_4108 );
not ( w_4108 , w_4109 );
and ( w_4109 , \1658_b1 , \1658_b0 );
or ( \1987_b1 , \1983_b1 , \1986_b1 );
not ( \1986_b1 , w_4110 );
and ( \1987_b0 , \1983_b0 , w_4111 );
and ( w_4110 , w_4111 , \1986_b0 );
or ( \1988_b1 , \1962_b1 , \1986_b1 );
not ( \1986_b1 , w_4112 );
and ( \1988_b0 , \1962_b0 , w_4113 );
and ( w_4112 , w_4113 , \1986_b0 );
or ( \1990_b1 , \1911_b1 , \1989_b1 );
not ( \1989_b1 , w_4114 );
and ( \1990_b0 , \1911_b0 , w_4115 );
and ( w_4114 , w_4115 , \1989_b0 );
or ( \1991_b1 , \1375_b1 , \1423_b1 );
xor ( \1991_b0 , \1375_b0 , w_4116 );
not ( w_4116 , w_4117 );
and ( w_4117 , \1423_b1 , \1423_b0 );
or ( \1992_b1 , \1991_b1 , \1484_b1 );
xor ( \1992_b0 , \1991_b0 , w_4118 );
not ( w_4118 , w_4119 );
and ( w_4119 , \1484_b1 , \1484_b0 );
or ( \1993_b1 , \1989_b1 , \1992_b1 );
not ( \1992_b1 , w_4120 );
and ( \1993_b0 , \1989_b0 , w_4121 );
and ( w_4120 , w_4121 , \1992_b0 );
or ( \1994_b1 , \1911_b1 , \1992_b1 );
not ( \1992_b1 , w_4122 );
and ( \1994_b0 , \1911_b0 , w_4123 );
and ( w_4122 , w_4123 , \1992_b0 );
or ( \1996_b1 , \1722_b1 , \1726_b1 );
not ( \1726_b1 , w_4124 );
and ( \1996_b0 , \1722_b0 , w_4125 );
and ( w_4124 , w_4125 , \1726_b0 );
or ( \1997_b1 , \1726_b1 , \1740_b1 );
not ( \1740_b1 , w_4126 );
and ( \1997_b0 , \1726_b0 , w_4127 );
and ( w_4126 , w_4127 , \1740_b0 );
or ( \1998_b1 , \1722_b1 , \1740_b1 );
not ( \1740_b1 , w_4128 );
and ( \1998_b0 , \1722_b0 , w_4129 );
and ( w_4128 , w_4129 , \1740_b0 );
or ( \2000_b1 , \1798_b1 , \1802_b1 );
not ( \1802_b1 , w_4130 );
and ( \2000_b0 , \1798_b0 , w_4131 );
and ( w_4130 , w_4131 , \1802_b0 );
or ( \2001_b1 , \1802_b1 , \1805_b1 );
not ( \1805_b1 , w_4132 );
and ( \2001_b0 , \1802_b0 , w_4133 );
and ( w_4132 , w_4133 , \1805_b0 );
or ( \2002_b1 , \1798_b1 , \1805_b1 );
not ( \1805_b1 , w_4134 );
and ( \2002_b0 , \1798_b0 , w_4135 );
and ( w_4134 , w_4135 , \1805_b0 );
or ( \2004_b1 , \1999_b1 , \2003_b1 );
xor ( \2004_b0 , \1999_b0 , w_4136 );
not ( w_4136 , w_4137 );
and ( w_4137 , \2003_b1 , \2003_b0 );
or ( \2005_b1 , \1855_b1 , \1859_b1 );
xor ( \2005_b0 , \1855_b0 , w_4138 );
not ( w_4138 , w_4139 );
and ( w_4139 , \1859_b1 , \1859_b0 );
or ( \2006_b1 , \2005_b1 , \1864_b1 );
xor ( \2006_b0 , \2005_b0 , w_4140 );
not ( w_4140 , w_4141 );
and ( w_4141 , \1864_b1 , \1864_b0 );
or ( \2007_b1 , \2004_b1 , \2006_b1 );
xor ( \2007_b0 , \2004_b0 , w_4142 );
not ( w_4142 , w_4143 );
and ( w_4143 , \2006_b1 , \2006_b0 );
or ( \2008_b1 , \1995_b1 , \2007_b1 );
not ( \2007_b1 , w_4144 );
and ( \2008_b0 , \1995_b0 , w_4145 );
and ( w_4144 , w_4145 , \2007_b0 );
or ( \2009_b1 , \1487_b1 , \1515_b1 );
xor ( \2009_b0 , \1487_b0 , w_4146 );
not ( w_4146 , w_4147 );
and ( w_4147 , \1515_b1 , \1515_b0 );
or ( \2010_b1 , \2009_b1 , \1591_b1 );
xor ( \2010_b0 , \2009_b0 , w_4148 );
not ( w_4148 , w_4149 );
and ( w_4149 , \1591_b1 , \1591_b0 );
or ( \2011_b1 , \2007_b1 , \2010_b1 );
not ( \2010_b1 , w_4150 );
and ( \2011_b0 , \2007_b0 , w_4151 );
and ( w_4150 , w_4151 , \2010_b0 );
or ( \2012_b1 , \1995_b1 , \2010_b1 );
not ( \2010_b1 , w_4152 );
and ( \2012_b0 , \1995_b0 , w_4153 );
and ( w_4152 , w_4153 , \2010_b0 );
or ( \2014_b1 , \1999_b1 , \2003_b1 );
not ( \2003_b1 , w_4154 );
and ( \2014_b0 , \1999_b0 , w_4155 );
and ( w_4154 , w_4155 , \2003_b0 );
or ( \2015_b1 , \2003_b1 , \2006_b1 );
not ( \2006_b1 , w_4156 );
and ( \2015_b0 , \2003_b0 , w_4157 );
and ( w_4156 , w_4157 , \2006_b0 );
or ( \2016_b1 , \1999_b1 , \2006_b1 );
not ( \2006_b1 , w_4158 );
and ( \2016_b0 , \1999_b0 , w_4159 );
and ( w_4158 , w_4159 , \2006_b0 );
or ( \2018_b1 , \1532_b1 , \1546_b1 );
not ( \1546_b1 , w_4160 );
and ( \2018_b0 , \1532_b0 , w_4161 );
and ( w_4160 , w_4161 , \1546_b0 );
or ( \2019_b1 , \1546_b1 , \1559_b1 );
not ( \1559_b1 , w_4162 );
and ( \2019_b0 , \1546_b0 , w_4163 );
and ( w_4162 , w_4163 , \1559_b0 );
or ( \2020_b1 , \1532_b1 , \1559_b1 );
not ( \1559_b1 , w_4164 );
and ( \2020_b0 , \1532_b0 , w_4165 );
and ( w_4164 , w_4165 , \1559_b0 );
or ( \2022_b1 , \1821_b1 , \1336_b1 );
not ( \1336_b1 , w_4166 );
and ( \2022_b0 , \1821_b0 , w_4167 );
and ( w_4166 , w_4167 , \1336_b0 );
buf ( \2023_b1 , \1179_A[30]_b1 );
buf ( \2023_b0 , \1179_A[30]_b0 );
or ( \2024_b1 , \2023_b1 , \1333_b1 );
not ( \1333_b1 , w_4168 );
and ( \2024_b0 , \2023_b0 , w_4169 );
and ( w_4168 , w_4169 , \1333_b0 );
or ( \2025_b1 , \2022_b1 , w_4171 );
not ( w_4171 , w_4172 );
and ( \2025_b0 , \2022_b0 , w_4173 );
and ( w_4172 ,  , w_4173 );
buf ( w_4171 , \2024_b1 );
not ( w_4171 , w_4174 );
not (  , w_4175 );
and ( w_4174 , w_4175 , \2024_b0 );
or ( \2026_b1 , \2025_b1 , w_4176 );
xor ( \2026_b0 , \2025_b0 , w_4178 );
not ( w_4178 , w_4179 );
and ( w_4179 , w_4176 , w_4177 );
buf ( w_4176 , \1332_b1 );
not ( w_4176 , w_4180 );
not ( w_4177 , w_4181 );
and ( w_4180 , w_4181 , \1332_b0 );
or ( \2027_b1 , \1446_b1 , \1349_b1 );
not ( \1349_b1 , w_4182 );
and ( \2027_b0 , \1446_b0 , w_4183 );
and ( w_4182 , w_4183 , \1349_b0 );
or ( \2028_b1 , \1425_b1 , \1347_b1 );
not ( \1347_b1 , w_4184 );
and ( \2028_b0 , \1425_b0 , w_4185 );
and ( w_4184 , w_4185 , \1347_b0 );
or ( \2029_b1 , \2027_b1 , w_4187 );
not ( w_4187 , w_4188 );
and ( \2029_b0 , \2027_b0 , w_4189 );
and ( w_4188 ,  , w_4189 );
buf ( w_4187 , \2028_b1 );
not ( w_4187 , w_4190 );
not (  , w_4191 );
and ( w_4190 , w_4191 , \2028_b0 );
or ( \2030_b1 , \2029_b1 , w_4192 );
xor ( \2030_b0 , \2029_b0 , w_4194 );
not ( w_4194 , w_4195 );
and ( w_4195 , w_4192 , w_4193 );
buf ( w_4192 , \1356_b1 );
not ( w_4192 , w_4196 );
not ( w_4193 , w_4197 );
and ( w_4196 , w_4197 , \1356_b0 );
or ( \2031_b1 , \2026_b1 , \2030_b1 );
xor ( \2031_b0 , \2026_b0 , w_4198 );
not ( w_4198 , w_4199 );
and ( w_4199 , \2030_b1 , \2030_b0 );
or ( \2032_b1 , \1470_b1 , \1366_b1 );
not ( \1366_b1 , w_4200 );
and ( \2032_b0 , \1470_b0 , w_4201 );
and ( w_4200 , w_4201 , \1366_b0 );
or ( \2033_b1 , \1477_b1 , \1364_b1 );
not ( \1364_b1 , w_4202 );
and ( \2033_b0 , \1477_b0 , w_4203 );
and ( w_4202 , w_4203 , \1364_b0 );
or ( \2034_b1 , \2032_b1 , w_4205 );
not ( w_4205 , w_4206 );
and ( \2034_b0 , \2032_b0 , w_4207 );
and ( w_4206 ,  , w_4207 );
buf ( w_4205 , \2033_b1 );
not ( w_4205 , w_4208 );
not (  , w_4209 );
and ( w_4208 , w_4209 , \2033_b0 );
or ( \2035_b1 , \2034_b1 , w_4210 );
xor ( \2035_b0 , \2034_b0 , w_4212 );
not ( w_4212 , w_4213 );
and ( w_4213 , w_4210 , w_4211 );
buf ( w_4210 , \1373_b1 );
not ( w_4210 , w_4214 );
not ( w_4211 , w_4215 );
and ( w_4214 , w_4215 , \1373_b0 );
or ( \2036_b1 , \2031_b1 , \2035_b1 );
xor ( \2036_b0 , \2031_b0 , w_4216 );
not ( w_4216 , w_4217 );
and ( w_4217 , \2035_b1 , \2035_b0 );
or ( \2037_b1 , \2021_b1 , \2036_b1 );
xor ( \2037_b0 , \2021_b0 , w_4218 );
not ( w_4218 , w_4219 );
and ( w_4219 , \2036_b1 , \2036_b0 );
or ( \2038_b1 , \1852_b1 , \1854_b1 );
not ( \1854_b1 , w_4220 );
and ( \2038_b0 , \1852_b0 , w_4221 );
and ( w_4220 , w_4221 , \1854_b0 );
or ( \2039_b1 , \1376_b1 , \1460_b1 );
not ( \1460_b1 , w_4222 );
and ( \2039_b0 , \1376_b0 , w_4223 );
and ( w_4222 , w_4223 , \1460_b0 );
or ( \2040_b1 , \1384_b1 , \1458_b1 );
not ( \1458_b1 , w_4224 );
and ( \2040_b0 , \1384_b0 , w_4225 );
and ( w_4224 , w_4225 , \1458_b0 );
or ( \2041_b1 , \2039_b1 , w_4227 );
not ( w_4227 , w_4228 );
and ( \2041_b0 , \2039_b0 , w_4229 );
and ( w_4228 ,  , w_4229 );
buf ( w_4227 , \2040_b1 );
not ( w_4227 , w_4230 );
not (  , w_4231 );
and ( w_4230 , w_4231 , \2040_b0 );
or ( \2042_b1 , \2041_b1 , w_4232 );
xor ( \2042_b0 , \2041_b0 , w_4234 );
not ( w_4234 , w_4235 );
and ( w_4235 , w_4232 , w_4233 );
buf ( w_4232 , \1467_b1 );
not ( w_4232 , w_4236 );
not ( w_4233 , w_4237 );
and ( w_4236 , w_4237 , \1467_b0 );
or ( \2043_b1 , \2038_b1 , \2042_b1 );
xor ( \2043_b0 , \2038_b0 , w_4238 );
not ( w_4238 , w_4239 );
and ( w_4239 , \2042_b1 , \2042_b0 );
or ( \2044_b1 , \1454_b1 , \1475_b1 );
not ( \1475_b1 , w_4240 );
and ( \2044_b0 , \1454_b0 , w_4241 );
and ( w_4240 , w_4241 , \1475_b0 );
or ( \2045_b1 , \1462_b1 , \1473_b1 );
not ( \1473_b1 , w_4242 );
and ( \2045_b0 , \1462_b0 , w_4243 );
and ( w_4242 , w_4243 , \1473_b0 );
or ( \2046_b1 , \2044_b1 , w_4245 );
not ( w_4245 , w_4246 );
and ( \2046_b0 , \2044_b0 , w_4247 );
and ( w_4246 ,  , w_4247 );
buf ( w_4245 , \2045_b1 );
not ( w_4245 , w_4248 );
not (  , w_4249 );
and ( w_4248 , w_4249 , \2045_b0 );
or ( \2047_b1 , \2046_b1 , w_4250 );
xor ( \2047_b0 , \2046_b0 , w_4252 );
not ( w_4252 , w_4253 );
and ( w_4253 , w_4250 , w_4251 );
buf ( w_4250 , \1482_b1 );
not ( w_4250 , w_4254 );
not ( w_4251 , w_4255 );
and ( w_4254 , w_4255 , \1482_b0 );
or ( \2048_b1 , \2043_b1 , \2047_b1 );
xor ( \2048_b0 , \2043_b0 , w_4256 );
not ( w_4256 , w_4257 );
and ( w_4257 , \2047_b1 , \2047_b0 );
or ( \2049_b1 , \2037_b1 , \2048_b1 );
xor ( \2049_b0 , \2037_b0 , w_4258 );
not ( w_4258 , w_4259 );
and ( w_4259 , \2048_b1 , \2048_b0 );
or ( \2050_b1 , \2017_b1 , \2049_b1 );
xor ( \2050_b0 , \2017_b0 , w_4260 );
not ( w_4260 , w_4261 );
and ( w_4261 , \2049_b1 , \2049_b0 );
or ( \2051_b1 , \1505_b1 , \1509_b1 );
not ( \1509_b1 , w_4262 );
and ( \2051_b0 , \1505_b0 , w_4263 );
and ( w_4262 , w_4263 , \1509_b0 );
or ( \2052_b1 , \1509_b1 , \1514_b1 );
not ( \1514_b1 , w_4264 );
and ( \2052_b0 , \1509_b0 , w_4265 );
and ( w_4264 , w_4265 , \1514_b0 );
or ( \2053_b1 , \1505_b1 , \1514_b1 );
not ( \1514_b1 , w_4266 );
and ( \2053_b0 , \1505_b0 , w_4267 );
and ( w_4266 , w_4267 , \1514_b0 );
or ( \2055_b1 , \1564_b1 , \1568_b1 );
not ( \1568_b1 , w_4268 );
and ( \2055_b0 , \1564_b0 , w_4269 );
and ( w_4268 , w_4269 , \1568_b0 );
or ( \2056_b1 , \1568_b1 , \1573_b1 );
not ( \1573_b1 , w_4270 );
and ( \2056_b0 , \1568_b0 , w_4271 );
and ( w_4270 , w_4271 , \1573_b0 );
or ( \2057_b1 , \1564_b1 , \1573_b1 );
not ( \1573_b1 , w_4272 );
and ( \2057_b0 , \1564_b0 , w_4273 );
and ( w_4272 , w_4273 , \1573_b0 );
or ( \2059_b1 , \1579_b1 , \1583_b1 );
not ( \1583_b1 , w_4274 );
and ( \2059_b0 , \1579_b0 , w_4275 );
and ( w_4274 , w_4275 , \1583_b0 );
or ( \2060_b1 , \1583_b1 , \1589_b1 );
not ( \1589_b1 , w_4276 );
and ( \2060_b0 , \1583_b0 , w_4277 );
and ( w_4276 , w_4277 , \1589_b0 );
or ( \2061_b1 , \1579_b1 , \1589_b1 );
not ( \1589_b1 , w_4278 );
and ( \2061_b0 , \1579_b0 , w_4279 );
and ( w_4278 , w_4279 , \1589_b0 );
or ( \2063_b1 , \2058_b1 , \2062_b1 );
xor ( \2063_b0 , \2058_b0 , w_4280 );
not ( w_4280 , w_4281 );
and ( w_4281 , \2062_b1 , \2062_b0 );
or ( \2064_b1 , \1824_b1 , \1828_b1 );
not ( \1828_b1 , w_4282 );
and ( \2064_b0 , \1824_b0 , w_4283 );
and ( w_4282 , w_4283 , \1828_b0 );
or ( \2065_b1 , \1828_b1 , \1833_b1 );
not ( \1833_b1 , w_4284 );
and ( \2065_b0 , \1828_b0 , w_4285 );
and ( w_4284 , w_4285 , \1833_b0 );
or ( \2066_b1 , \1824_b1 , \1833_b1 );
not ( \1833_b1 , w_4286 );
and ( \2066_b0 , \1824_b0 , w_4287 );
and ( w_4286 , w_4287 , \1833_b0 );
or ( \2068_b1 , \2063_b1 , \2067_b1 );
xor ( \2068_b0 , \2063_b0 , w_4288 );
not ( w_4288 , w_4289 );
and ( w_4289 , \2067_b1 , \2067_b0 );
or ( \2069_b1 , \2054_b1 , \2068_b1 );
xor ( \2069_b0 , \2054_b0 , w_4290 );
not ( w_4290 , w_4291 );
and ( w_4291 , \2068_b1 , \2068_b0 );
or ( \2070_b1 , \1540_b1 , \1538_b1 );
not ( \1538_b1 , w_4292 );
and ( \2070_b0 , \1540_b0 , w_4293 );
and ( w_4292 , w_4293 , \1538_b0 );
or ( \2071_b1 , \1517_b1 , \1536_b1 );
not ( \1536_b1 , w_4294 );
and ( \2071_b0 , \1517_b0 , w_4295 );
and ( w_4294 , w_4295 , \1536_b0 );
or ( \2072_b1 , \2070_b1 , w_4297 );
not ( w_4297 , w_4298 );
and ( \2072_b0 , \2070_b0 , w_4299 );
and ( w_4298 ,  , w_4299 );
buf ( w_4297 , \2071_b1 );
not ( w_4297 , w_4300 );
not (  , w_4301 );
and ( w_4300 , w_4301 , \2071_b0 );
or ( \2073_b1 , \2072_b1 , w_4302 );
xor ( \2073_b0 , \2072_b0 , w_4304 );
not ( w_4304 , w_4305 );
and ( w_4305 , w_4302 , w_4303 );
buf ( w_4302 , \1545_b1 );
not ( w_4302 , w_4306 );
not ( w_4303 , w_4307 );
and ( w_4306 , w_4307 , \1545_b0 );
or ( \2074_b1 , \1553_b1 , \1551_b1 );
not ( \1551_b1 , w_4308 );
and ( \2074_b0 , \1553_b0 , w_4309 );
and ( w_4308 , w_4309 , \1551_b0 );
or ( \2075_b1 , \1533_b1 , \1501_b1 );
not ( \1501_b1 , w_4310 );
and ( \2075_b0 , \1533_b0 , w_4311 );
and ( w_4310 , w_4311 , \1501_b0 );
or ( \2076_b1 , \2074_b1 , w_4313 );
not ( w_4313 , w_4314 );
and ( \2076_b0 , \2074_b0 , w_4315 );
and ( w_4314 ,  , w_4315 );
buf ( w_4313 , \2075_b1 );
not ( w_4313 , w_4316 );
not (  , w_4317 );
and ( w_4316 , w_4317 , \2075_b0 );
or ( \2077_b1 , \2076_b1 , w_4318 );
xor ( \2077_b0 , \2076_b0 , w_4320 );
not ( w_4320 , w_4321 );
and ( w_4321 , w_4318 , w_4319 );
buf ( w_4318 , \1558_b1 );
not ( w_4318 , w_4322 );
not ( w_4319 , w_4323 );
and ( w_4322 , w_4323 , \1558_b0 );
or ( \2078_b1 , \2073_b1 , \2077_b1 );
xor ( \2078_b0 , \2073_b0 , w_4324 );
not ( w_4324 , w_4325 );
and ( w_4325 , \2077_b1 , \2077_b0 );
or ( \2079_b1 , \1331_b1 , \1431_b1 );
not ( \1431_b1 , w_4326 );
and ( \2079_b0 , \1331_b0 , w_4327 );
and ( w_4326 , w_4327 , \1431_b0 );
or ( \2080_b1 , \1338_b1 , \1429_b1 );
not ( \1429_b1 , w_4328 );
and ( \2080_b0 , \1338_b0 , w_4329 );
and ( w_4328 , w_4329 , \1429_b0 );
or ( \2081_b1 , \2079_b1 , w_4331 );
not ( w_4331 , w_4332 );
and ( \2081_b0 , \2079_b0 , w_4333 );
and ( w_4332 ,  , w_4333 );
buf ( w_4331 , \2080_b1 );
not ( w_4331 , w_4334 );
not (  , w_4335 );
and ( w_4334 , w_4335 , \2080_b0 );
or ( \2082_b1 , \2081_b1 , w_4336 );
xor ( \2082_b0 , \2081_b0 , w_4338 );
not ( w_4338 , w_4339 );
and ( w_4339 , w_4336 , w_4337 );
buf ( w_4336 , \1438_b1 );
not ( w_4336 , w_4340 );
not ( w_4337 , w_4341 );
and ( w_4340 , w_4341 , \1438_b0 );
or ( \2083_b1 , \1433_b1 , \1444_b1 );
not ( \1444_b1 , w_4342 );
and ( \2083_b0 , \1433_b0 , w_4343 );
and ( w_4342 , w_4343 , \1444_b0 );
or ( \2084_b1 , \1489_b1 , \1442_b1 );
not ( \1442_b1 , w_4344 );
and ( \2084_b0 , \1489_b0 , w_4345 );
and ( w_4344 , w_4345 , \1442_b0 );
or ( \2085_b1 , \2083_b1 , w_4347 );
not ( w_4347 , w_4348 );
and ( \2085_b0 , \2083_b0 , w_4349 );
and ( w_4348 ,  , w_4349 );
buf ( w_4347 , \2084_b1 );
not ( w_4347 , w_4350 );
not (  , w_4351 );
and ( w_4350 , w_4351 , \2084_b0 );
or ( \2086_b1 , \2085_b1 , w_4352 );
xor ( \2086_b0 , \2085_b0 , w_4354 );
not ( w_4354 , w_4355 );
and ( w_4355 , w_4352 , w_4353 );
buf ( w_4352 , \1451_b1 );
not ( w_4352 , w_4356 );
not ( w_4353 , w_4357 );
and ( w_4356 , w_4357 , \1451_b0 );
or ( \2087_b1 , \2082_b1 , \2086_b1 );
xor ( \2087_b0 , \2082_b0 , w_4358 );
not ( w_4358 , w_4359 );
and ( w_4359 , \2086_b1 , \2086_b0 );
buf ( \2088_b1 , \1300_B[30]_b1 );
buf ( \2088_b0 , \1300_B[30]_b0 );
or ( \2089_b1 , \2088_b1 , \1548_b1 );
xor ( \2089_b0 , \2088_b0 , w_4360 );
not ( w_4360 , w_4361 );
and ( w_4361 , \1548_b1 , \1548_b0 );
or ( \2090_b1 , \1498_b1 , \2089_b1 );
not ( \2089_b1 , w_4362 );
and ( \2090_b0 , \1498_b0 , w_4363 );
and ( w_4362 , w_4363 , \2089_b0 );
or ( \2091_b1 , \2087_b1 , \2090_b1 );
xor ( \2091_b0 , \2087_b0 , w_4364 );
not ( w_4364 , w_4365 );
and ( w_4365 , \2090_b1 , \2090_b0 );
or ( \2092_b1 , \2078_b1 , \2091_b1 );
xor ( \2092_b0 , \2078_b0 , w_4366 );
not ( w_4366 , w_4367 );
and ( w_4367 , \2091_b1 , \2091_b0 );
or ( \2093_b1 , \2069_b1 , \2092_b1 );
xor ( \2093_b0 , \2069_b0 , w_4368 );
not ( w_4368 , w_4369 );
and ( w_4369 , \2092_b1 , \2092_b0 );
or ( \2094_b1 , \2050_b1 , \2093_b1 );
xor ( \2094_b0 , \2050_b0 , w_4370 );
not ( w_4370 , w_4371 );
and ( w_4371 , \2093_b1 , \2093_b0 );
or ( \2095_b1 , \2013_b1 , \2094_b1 );
not ( \2094_b1 , w_4372 );
and ( \2095_b0 , \2013_b0 , w_4373 );
and ( w_4372 , w_4373 , \2094_b0 );
or ( \2096_b1 , \1594_b1 , \1838_b1 );
xor ( \2096_b0 , \1594_b0 , w_4374 );
not ( w_4374 , w_4375 );
and ( w_4375 , \1838_b1 , \1838_b0 );
or ( \2097_b1 , \2096_b1 , \1898_b1 );
xor ( \2097_b0 , \2096_b0 , w_4376 );
not ( w_4376 , w_4377 );
and ( w_4377 , \1898_b1 , \1898_b0 );
or ( \2098_b1 , \2094_b1 , \2097_b1 );
not ( \2097_b1 , w_4378 );
and ( \2098_b0 , \2094_b0 , w_4379 );
and ( w_4378 , w_4379 , \2097_b0 );
or ( \2099_b1 , \2013_b1 , \2097_b1 );
not ( \2097_b1 , w_4380 );
and ( \2099_b0 , \2013_b0 , w_4381 );
and ( w_4380 , w_4381 , \2097_b0 );
or ( \2101_b1 , \1901_b1 , \2100_b1 );
xor ( \2101_b0 , \1901_b0 , w_4382 );
not ( w_4382 , w_4383 );
and ( w_4383 , \2100_b1 , \2100_b0 );
or ( \2102_b1 , \2017_b1 , \2049_b1 );
not ( \2049_b1 , w_4384 );
and ( \2102_b0 , \2017_b0 , w_4385 );
and ( w_4384 , w_4385 , \2049_b0 );
or ( \2103_b1 , \2049_b1 , \2093_b1 );
not ( \2093_b1 , w_4386 );
and ( \2103_b0 , \2049_b0 , w_4387 );
and ( w_4386 , w_4387 , \2093_b0 );
or ( \2104_b1 , \2017_b1 , \2093_b1 );
not ( \2093_b1 , w_4388 );
and ( \2104_b0 , \2017_b0 , w_4389 );
and ( w_4388 , w_4389 , \2093_b0 );
or ( \2106_b1 , \2054_b1 , \2068_b1 );
not ( \2068_b1 , w_4390 );
and ( \2106_b0 , \2054_b0 , w_4391 );
and ( w_4390 , w_4391 , \2068_b0 );
or ( \2107_b1 , \2068_b1 , \2092_b1 );
not ( \2092_b1 , w_4392 );
and ( \2107_b0 , \2068_b0 , w_4393 );
and ( w_4392 , w_4393 , \2092_b0 );
or ( \2108_b1 , \2054_b1 , \2092_b1 );
not ( \2092_b1 , w_4394 );
and ( \2108_b0 , \2054_b0 , w_4395 );
and ( w_4394 , w_4395 , \2092_b0 );
or ( \2110_b1 , \1871_b1 , \1875_b1 );
not ( \1875_b1 , w_4396 );
and ( \2110_b0 , \1871_b0 , w_4397 );
and ( w_4396 , w_4397 , \1875_b0 );
or ( \2111_b1 , \1875_b1 , \1880_b1 );
not ( \1880_b1 , w_4398 );
and ( \2111_b0 , \1875_b0 , w_4399 );
and ( w_4398 , w_4399 , \1880_b0 );
or ( \2112_b1 , \1871_b1 , \1880_b1 );
not ( \1880_b1 , w_4400 );
and ( \2112_b0 , \1871_b0 , w_4401 );
and ( w_4400 , w_4401 , \1880_b0 );
or ( \2114_b1 , \2073_b1 , \2077_b1 );
not ( \2077_b1 , w_4402 );
and ( \2114_b0 , \2073_b0 , w_4403 );
and ( w_4402 , w_4403 , \2077_b0 );
or ( \2115_b1 , \2077_b1 , \2091_b1 );
not ( \2091_b1 , w_4404 );
and ( \2115_b0 , \2077_b0 , w_4405 );
and ( w_4404 , w_4405 , \2091_b0 );
or ( \2116_b1 , \2073_b1 , \2091_b1 );
not ( \2091_b1 , w_4406 );
and ( \2116_b0 , \2073_b0 , w_4407 );
and ( w_4406 , w_4407 , \2091_b0 );
or ( \2118_b1 , \2113_b1 , \2117_b1 );
xor ( \2118_b0 , \2113_b0 , w_4408 );
not ( w_4408 , w_4409 );
and ( w_4409 , \2117_b1 , \2117_b0 );
or ( \2119_b1 , \1399_b1 , \1675_b1 );
not ( \1675_b1 , w_4410 );
and ( \2119_b0 , \1399_b0 , w_4411 );
and ( w_4410 , w_4411 , \1675_b0 );
or ( \2120_b1 , \1359_b1 , \1673_b1 );
not ( \1673_b1 , w_4412 );
and ( \2120_b0 , \1359_b0 , w_4413 );
and ( w_4412 , w_4413 , \1673_b0 );
or ( \2121_b1 , \2119_b1 , w_4415 );
not ( w_4415 , w_4416 );
and ( \2121_b0 , \2119_b0 , w_4417 );
and ( w_4416 ,  , w_4417 );
buf ( w_4415 , \2120_b1 );
not ( w_4415 , w_4418 );
not (  , w_4419 );
and ( w_4418 , w_4419 , \2120_b0 );
or ( \2122_b1 , \2121_b1 , w_4420 );
xor ( \2122_b0 , \2121_b0 , w_4422 );
not ( w_4422 , w_4423 );
and ( w_4423 , w_4420 , w_4421 );
buf ( w_4420 , \1681_b1 );
not ( w_4420 , w_4424 );
not ( w_4421 , w_4425 );
and ( w_4424 , w_4425 , \1681_b0 );
or ( \2123_b1 , \1517_b1 , \1538_b1 );
not ( \1538_b1 , w_4426 );
and ( \2123_b0 , \1517_b0 , w_4427 );
and ( w_4426 , w_4427 , \1538_b0 );
or ( \2124_b1 , \1526_b1 , \1536_b1 );
not ( \1536_b1 , w_4428 );
and ( \2124_b0 , \1526_b0 , w_4429 );
and ( w_4428 , w_4429 , \1536_b0 );
or ( \2125_b1 , \2123_b1 , w_4431 );
not ( w_4431 , w_4432 );
and ( \2125_b0 , \2123_b0 , w_4433 );
and ( w_4432 ,  , w_4433 );
buf ( w_4431 , \2124_b1 );
not ( w_4431 , w_4434 );
not (  , w_4435 );
and ( w_4434 , w_4435 , \2124_b0 );
or ( \2126_b1 , \2125_b1 , w_4436 );
xor ( \2126_b0 , \2125_b0 , w_4438 );
not ( w_4438 , w_4439 );
and ( w_4439 , w_4436 , w_4437 );
buf ( w_4436 , \1545_b1 );
not ( w_4436 , w_4440 );
not ( w_4437 , w_4441 );
and ( w_4440 , w_4441 , \1545_b0 );
or ( \2127_b1 , \2122_b1 , \2126_b1 );
xor ( \2127_b0 , \2122_b0 , w_4442 );
not ( w_4442 , w_4443 );
and ( w_4443 , \2126_b1 , \2126_b0 );
or ( \2128_b1 , \1533_b1 , \1551_b1 );
not ( \1551_b1 , w_4444 );
and ( \2128_b0 , \1533_b0 , w_4445 );
and ( w_4444 , w_4445 , \1551_b0 );
or ( \2129_b1 , \1540_b1 , \1501_b1 );
not ( \1501_b1 , w_4446 );
and ( \2129_b0 , \1540_b0 , w_4447 );
and ( w_4446 , w_4447 , \1501_b0 );
or ( \2130_b1 , \2128_b1 , w_4449 );
not ( w_4449 , w_4450 );
and ( \2130_b0 , \2128_b0 , w_4451 );
and ( w_4450 ,  , w_4451 );
buf ( w_4449 , \2129_b1 );
not ( w_4449 , w_4452 );
not (  , w_4453 );
and ( w_4452 , w_4453 , \2129_b0 );
or ( \2131_b1 , \2130_b1 , w_4454 );
xor ( \2131_b0 , \2130_b0 , w_4456 );
not ( w_4456 , w_4457 );
and ( w_4457 , w_4454 , w_4455 );
buf ( w_4454 , \1558_b1 );
not ( w_4454 , w_4458 );
not ( w_4455 , w_4459 );
and ( w_4458 , w_4459 , \1558_b0 );
or ( \2132_b1 , \2127_b1 , \2131_b1 );
xor ( \2132_b0 , \2127_b0 , w_4460 );
not ( w_4460 , w_4461 );
and ( w_4461 , \2131_b1 , \2131_b0 );
or ( \2133_b1 , \2118_b1 , \2132_b1 );
xor ( \2133_b0 , \2118_b0 , w_4462 );
not ( w_4462 , w_4463 );
and ( w_4463 , \2132_b1 , \2132_b0 );
or ( \2134_b1 , \2109_b1 , \2133_b1 );
xor ( \2134_b0 , \2109_b0 , w_4464 );
not ( w_4464 , w_4465 );
and ( w_4465 , \2133_b1 , \2133_b0 );
or ( \2135_b1 , \1886_b1 , \1890_b1 );
not ( \1890_b1 , w_4466 );
and ( \2135_b0 , \1886_b0 , w_4467 );
and ( w_4466 , w_4467 , \1890_b0 );
or ( \2136_b1 , \1890_b1 , \1895_b1 );
not ( \1895_b1 , w_4468 );
and ( \2136_b0 , \1890_b0 , w_4469 );
and ( w_4468 , w_4469 , \1895_b0 );
or ( \2137_b1 , \1886_b1 , \1895_b1 );
not ( \1895_b1 , w_4470 );
and ( \2137_b0 , \1886_b0 , w_4471 );
and ( w_4470 , w_4471 , \1895_b0 );
or ( \2139_b1 , \2038_b1 , \2042_b1 );
not ( \2042_b1 , w_4472 );
and ( \2139_b0 , \2038_b0 , w_4473 );
and ( w_4472 , w_4473 , \2042_b0 );
or ( \2140_b1 , \2042_b1 , \2047_b1 );
not ( \2047_b1 , w_4474 );
and ( \2140_b0 , \2042_b0 , w_4475 );
and ( w_4474 , w_4475 , \2047_b0 );
or ( \2141_b1 , \2038_b1 , \2047_b1 );
not ( \2047_b1 , w_4476 );
and ( \2141_b0 , \2038_b0 , w_4477 );
and ( w_4476 , w_4477 , \2047_b0 );
or ( \2143_b1 , \2138_b1 , \2142_b1 );
xor ( \2143_b0 , \2138_b0 , w_4478 );
not ( w_4478 , w_4479 );
and ( w_4479 , \2142_b1 , \2142_b0 );
or ( \2144_b1 , \1338_b1 , \1431_b1 );
not ( \1431_b1 , w_4480 );
and ( \2144_b0 , \1338_b0 , w_4481 );
and ( w_4480 , w_4481 , \1431_b0 );
or ( \2145_b1 , \1821_b1 , \1429_b1 );
not ( \1429_b1 , w_4482 );
and ( \2145_b0 , \1821_b0 , w_4483 );
and ( w_4482 , w_4483 , \1429_b0 );
or ( \2146_b1 , \2144_b1 , w_4485 );
not ( w_4485 , w_4486 );
and ( \2146_b0 , \2144_b0 , w_4487 );
and ( w_4486 ,  , w_4487 );
buf ( w_4485 , \2145_b1 );
not ( w_4485 , w_4488 );
not (  , w_4489 );
and ( w_4488 , w_4489 , \2145_b0 );
or ( \2147_b1 , \2146_b1 , w_4490 );
xor ( \2147_b0 , \2146_b0 , w_4492 );
not ( w_4492 , w_4493 );
and ( w_4493 , w_4490 , w_4491 );
buf ( w_4490 , \1438_b1 );
not ( w_4490 , w_4494 );
not ( w_4491 , w_4495 );
and ( w_4494 , w_4495 , \1438_b0 );
or ( \2148_b1 , \1489_b1 , \1444_b1 );
not ( \1444_b1 , w_4496 );
and ( \2148_b0 , \1489_b0 , w_4497 );
and ( w_4496 , w_4497 , \1444_b0 );
or ( \2149_b1 , \1331_b1 , \1442_b1 );
not ( \1442_b1 , w_4498 );
and ( \2149_b0 , \1331_b0 , w_4499 );
and ( w_4498 , w_4499 , \1442_b0 );
or ( \2150_b1 , \2148_b1 , w_4501 );
not ( w_4501 , w_4502 );
and ( \2150_b0 , \2148_b0 , w_4503 );
and ( w_4502 ,  , w_4503 );
buf ( w_4501 , \2149_b1 );
not ( w_4501 , w_4504 );
not (  , w_4505 );
and ( w_4504 , w_4505 , \2149_b0 );
or ( \2151_b1 , \2150_b1 , w_4506 );
xor ( \2151_b0 , \2150_b0 , w_4508 );
not ( w_4508 , w_4509 );
and ( w_4509 , w_4506 , w_4507 );
buf ( w_4506 , \1451_b1 );
not ( w_4506 , w_4510 );
not ( w_4507 , w_4511 );
and ( w_4510 , w_4511 , \1451_b0 );
or ( \2152_b1 , \2147_b1 , \2151_b1 );
xor ( \2152_b0 , \2147_b0 , w_4512 );
not ( w_4512 , w_4513 );
and ( w_4513 , \2151_b1 , \2151_b0 );
or ( \2153_b1 , \1616_b1 , \1414_b1 );
not ( \1414_b1 , w_4514 );
and ( \2153_b0 , \1616_b0 , w_4515 );
and ( w_4514 , w_4515 , \1414_b0 );
or ( \2154_b1 , \1391_b1 , \1412_b1 );
not ( \1412_b1 , w_4516 );
and ( \2154_b0 , \1391_b0 , w_4517 );
and ( w_4516 , w_4517 , \1412_b0 );
or ( \2155_b1 , \2153_b1 , w_4519 );
not ( w_4519 , w_4520 );
and ( \2155_b0 , \2153_b0 , w_4521 );
and ( w_4520 ,  , w_4521 );
buf ( w_4519 , \2154_b1 );
not ( w_4519 , w_4522 );
not (  , w_4523 );
and ( w_4522 , w_4523 , \2154_b0 );
or ( \2156_b1 , \2155_b1 , w_4524 );
xor ( \2156_b0 , \2155_b0 , w_4526 );
not ( w_4526 , w_4527 );
and ( w_4527 , w_4524 , w_4525 );
buf ( w_4524 , \1421_b1 );
not ( w_4524 , w_4528 );
not ( w_4525 , w_4529 );
and ( w_4528 , w_4529 , \1421_b0 );
or ( \2157_b1 , \2152_b1 , \2156_b1 );
xor ( \2157_b0 , \2152_b0 , w_4530 );
not ( w_4530 , w_4531 );
and ( w_4531 , \2156_b1 , \2156_b0 );
or ( \2158_b1 , \1622_b1 , \1524_b1 );
not ( \1524_b1 , w_4532 );
and ( \2158_b0 , \1622_b0 , w_4533 );
and ( w_4532 , w_4533 , \1524_b0 );
or ( \2159_b1 , \1407_b1 , \1522_b1 );
not ( \1522_b1 , w_4534 );
and ( \2159_b0 , \1407_b0 , w_4535 );
and ( w_4534 , w_4535 , \1522_b0 );
or ( \2160_b1 , \2158_b1 , w_4537 );
not ( w_4537 , w_4538 );
and ( \2160_b0 , \2158_b0 , w_4539 );
and ( w_4538 ,  , w_4539 );
buf ( w_4537 , \2159_b1 );
not ( w_4537 , w_4540 );
not (  , w_4541 );
and ( w_4540 , w_4541 , \2159_b0 );
or ( \2161_b1 , \2160_b1 , w_4542 );
xor ( \2161_b0 , \2160_b0 , w_4544 );
not ( w_4544 , w_4545 );
and ( w_4545 , w_4542 , w_4543 );
buf ( w_4542 , \1531_b1 );
not ( w_4542 , w_4546 );
not ( w_4543 , w_4547 );
and ( w_4546 , w_4547 , \1531_b0 );
or ( \2162_b1 , \2157_b1 , \2161_b1 );
xor ( \2162_b0 , \2157_b0 , w_4548 );
not ( w_4548 , w_4549 );
and ( w_4549 , \2161_b1 , \2161_b0 );
or ( \2163_b1 , \2143_b1 , \2162_b1 );
xor ( \2163_b0 , \2143_b0 , w_4550 );
not ( w_4550 , w_4551 );
and ( w_4551 , \2162_b1 , \2162_b0 );
or ( \2164_b1 , \1425_b1 , \1349_b1 );
not ( \1349_b1 , w_4552 );
and ( \2164_b0 , \1425_b0 , w_4553 );
and ( w_4552 , w_4553 , \1349_b0 );
or ( \2165_b1 , \1433_b1 , \1347_b1 );
not ( \1347_b1 , w_4554 );
and ( \2165_b0 , \1433_b0 , w_4555 );
and ( w_4554 , w_4555 , \1347_b0 );
or ( \2166_b1 , \2164_b1 , w_4557 );
not ( w_4557 , w_4558 );
and ( \2166_b0 , \2164_b0 , w_4559 );
and ( w_4558 ,  , w_4559 );
buf ( w_4557 , \2165_b1 );
not ( w_4557 , w_4560 );
not (  , w_4561 );
and ( w_4560 , w_4561 , \2165_b0 );
or ( \2167_b1 , \2166_b1 , w_4562 );
xor ( \2167_b0 , \2166_b0 , w_4564 );
not ( w_4564 , w_4565 );
and ( w_4565 , w_4562 , w_4563 );
buf ( w_4562 , \1356_b1 );
not ( w_4562 , w_4566 );
not ( w_4563 , w_4567 );
and ( w_4566 , w_4567 , \1356_b0 );
or ( \2168_b1 , \1462_b1 , \1475_b1 );
not ( \1475_b1 , w_4568 );
and ( \2168_b0 , \1462_b0 , w_4569 );
and ( w_4568 , w_4569 , \1475_b0 );
or ( \2169_b1 , \1376_b1 , \1473_b1 );
not ( \1473_b1 , w_4570 );
and ( \2169_b0 , \1376_b0 , w_4571 );
and ( w_4570 , w_4571 , \1473_b0 );
or ( \2170_b1 , \2168_b1 , w_4573 );
not ( w_4573 , w_4574 );
and ( \2170_b0 , \2168_b0 , w_4575 );
and ( w_4574 ,  , w_4575 );
buf ( w_4573 , \2169_b1 );
not ( w_4573 , w_4576 );
not (  , w_4577 );
and ( w_4576 , w_4577 , \2169_b0 );
or ( \2171_b1 , \2170_b1 , w_4578 );
xor ( \2171_b0 , \2170_b0 , w_4580 );
not ( w_4580 , w_4581 );
and ( w_4581 , w_4578 , w_4579 );
buf ( w_4578 , \1482_b1 );
not ( w_4578 , w_4582 );
not ( w_4579 , w_4583 );
and ( w_4582 , w_4583 , \1482_b0 );
or ( \2172_b1 , \2167_b1 , \2171_b1 );
xor ( \2172_b0 , \2167_b0 , w_4584 );
not ( w_4584 , w_4585 );
and ( w_4585 , \2171_b1 , \2171_b0 );
or ( \2173_b1 , \1477_b1 , \1366_b1 );
not ( \1366_b1 , w_4586 );
and ( \2173_b0 , \1477_b0 , w_4587 );
and ( w_4586 , w_4587 , \1366_b0 );
or ( \2174_b1 , \1454_b1 , \1364_b1 );
not ( \1364_b1 , w_4588 );
and ( \2174_b0 , \1454_b0 , w_4589 );
and ( w_4588 , w_4589 , \1364_b0 );
or ( \2175_b1 , \2173_b1 , w_4591 );
not ( w_4591 , w_4592 );
and ( \2175_b0 , \2173_b0 , w_4593 );
and ( w_4592 ,  , w_4593 );
buf ( w_4591 , \2174_b1 );
not ( w_4591 , w_4594 );
not (  , w_4595 );
and ( w_4594 , w_4595 , \2174_b0 );
or ( \2176_b1 , \2175_b1 , w_4596 );
xor ( \2176_b0 , \2175_b0 , w_4598 );
not ( w_4598 , w_4599 );
and ( w_4599 , w_4596 , w_4597 );
buf ( w_4596 , \1373_b1 );
not ( w_4596 , w_4600 );
not ( w_4597 , w_4601 );
and ( w_4600 , w_4601 , \1373_b0 );
or ( \2177_b1 , \2172_b1 , \2176_b1 );
xor ( \2177_b0 , \2172_b0 , w_4602 );
not ( w_4602 , w_4603 );
and ( w_4603 , \2176_b1 , \2176_b0 );
or ( \2178_b1 , \1368_b1 , \1397_b1 );
not ( \1397_b1 , w_4604 );
and ( \2178_b0 , \1368_b0 , w_4605 );
and ( w_4604 , w_4605 , \1397_b0 );
or ( \2179_b1 , \1470_b1 , \1395_b1 );
not ( \1395_b1 , w_4606 );
and ( \2179_b0 , \1470_b0 , w_4607 );
and ( w_4606 , w_4607 , \1395_b0 );
or ( \2180_b1 , \2178_b1 , w_4609 );
not ( w_4609 , w_4610 );
and ( \2180_b0 , \2178_b0 , w_4611 );
and ( w_4610 ,  , w_4611 );
buf ( w_4609 , \2179_b1 );
not ( w_4609 , w_4612 );
not (  , w_4613 );
and ( w_4612 , w_4613 , \2179_b0 );
or ( \2181_b1 , \2180_b1 , w_4614 );
xor ( \2181_b0 , \2180_b0 , w_4616 );
not ( w_4616 , w_4617 );
and ( w_4617 , w_4614 , w_4615 );
buf ( w_4614 , \1404_b1 );
not ( w_4614 , w_4618 );
not ( w_4615 , w_4619 );
and ( w_4618 , w_4619 , \1404_b0 );
or ( \2182_b1 , \2177_b1 , \2181_b1 );
xor ( \2182_b0 , \2177_b0 , w_4620 );
not ( w_4620 , w_4621 );
and ( w_4621 , \2181_b1 , \2181_b0 );
or ( \2183_b1 , \2163_b1 , \2182_b1 );
xor ( \2183_b0 , \2163_b0 , w_4622 );
not ( w_4622 , w_4623 );
and ( w_4623 , \2182_b1 , \2182_b0 );
or ( \2184_b1 , \2134_b1 , \2183_b1 );
xor ( \2184_b0 , \2134_b0 , w_4624 );
not ( w_4624 , w_4625 );
and ( w_4625 , \2183_b1 , \2183_b0 );
or ( \2185_b1 , \2105_b1 , \2184_b1 );
xor ( \2185_b0 , \2105_b0 , w_4626 );
not ( w_4626 , w_4627 );
and ( w_4627 , \2184_b1 , \2184_b0 );
or ( \2186_b1 , \2058_b1 , \2062_b1 );
not ( \2062_b1 , w_4628 );
and ( \2186_b0 , \2058_b0 , w_4629 );
and ( w_4628 , w_4629 , \2062_b0 );
or ( \2187_b1 , \2062_b1 , \2067_b1 );
not ( \2067_b1 , w_4630 );
and ( \2187_b0 , \2062_b0 , w_4631 );
and ( w_4630 , w_4631 , \2067_b0 );
or ( \2188_b1 , \2058_b1 , \2067_b1 );
not ( \2067_b1 , w_4632 );
and ( \2188_b0 , \2058_b0 , w_4633 );
and ( w_4632 , w_4633 , \2067_b0 );
or ( \2190_b1 , \2021_b1 , \2036_b1 );
not ( \2036_b1 , w_4634 );
and ( \2190_b0 , \2021_b0 , w_4635 );
and ( w_4634 , w_4635 , \2036_b0 );
or ( \2191_b1 , \2036_b1 , \2048_b1 );
not ( \2048_b1 , w_4636 );
and ( \2191_b0 , \2036_b0 , w_4637 );
and ( w_4636 , w_4637 , \2048_b0 );
or ( \2192_b1 , \2021_b1 , \2048_b1 );
not ( \2048_b1 , w_4638 );
and ( \2192_b0 , \2021_b0 , w_4639 );
and ( w_4638 , w_4639 , \2048_b0 );
or ( \2194_b1 , \2189_b1 , \2193_b1 );
xor ( \2194_b0 , \2189_b0 , w_4640 );
not ( w_4640 , w_4641 );
and ( w_4641 , \2193_b1 , \2193_b0 );
or ( \2195_b1 , \1867_b1 , \1881_b1 );
not ( \1881_b1 , w_4642 );
and ( \2195_b0 , \1867_b0 , w_4643 );
and ( w_4642 , w_4643 , \1881_b0 );
or ( \2196_b1 , \1881_b1 , \1896_b1 );
not ( \1896_b1 , w_4644 );
and ( \2196_b0 , \1881_b0 , w_4645 );
and ( w_4644 , w_4645 , \1896_b0 );
or ( \2197_b1 , \1867_b1 , \1896_b1 );
not ( \1896_b1 , w_4646 );
and ( \2197_b0 , \1867_b0 , w_4647 );
and ( w_4646 , w_4647 , \1896_b0 );
or ( \2199_b1 , \1843_b1 , \1847_b1 );
not ( \1847_b1 , w_4648 );
and ( \2199_b0 , \1843_b0 , w_4649 );
and ( w_4648 , w_4649 , \1847_b0 );
or ( \2200_b1 , \1847_b1 , \1897_b1 );
not ( \1897_b1 , w_4650 );
and ( \2200_b0 , \1847_b0 , w_4651 );
and ( w_4650 , w_4651 , \1897_b0 );
or ( \2201_b1 , \1843_b1 , \1897_b1 );
not ( \1897_b1 , w_4652 );
and ( \2201_b0 , \1843_b0 , w_4653 );
and ( w_4652 , w_4653 , \1897_b0 );
or ( \2203_b1 , \2198_b1 , \2202_b1 );
xor ( \2203_b0 , \2198_b0 , w_4654 );
not ( w_4654 , w_4655 );
and ( w_4655 , \2202_b1 , \2202_b0 );
or ( \2204_b1 , \2026_b1 , \2030_b1 );
not ( \2030_b1 , w_4656 );
and ( \2204_b0 , \2026_b0 , w_4657 );
and ( w_4656 , w_4657 , \2030_b0 );
or ( \2205_b1 , \2030_b1 , \2035_b1 );
not ( \2035_b1 , w_4658 );
and ( \2205_b0 , \2030_b0 , w_4659 );
and ( w_4658 , w_4659 , \2035_b0 );
or ( \2206_b1 , \2026_b1 , \2035_b1 );
not ( \2035_b1 , w_4660 );
and ( \2206_b0 , \2026_b0 , w_4661 );
and ( w_4660 , w_4661 , \2035_b0 );
or ( \2208_b1 , \2082_b1 , \2086_b1 );
not ( \2086_b1 , w_4662 );
and ( \2208_b0 , \2082_b0 , w_4663 );
and ( w_4662 , w_4663 , \2086_b0 );
or ( \2209_b1 , \2086_b1 , \2090_b1 );
not ( \2090_b1 , w_4664 );
and ( \2209_b0 , \2086_b0 , w_4665 );
and ( w_4664 , w_4665 , \2090_b0 );
or ( \2210_b1 , \2082_b1 , \2090_b1 );
not ( \2090_b1 , w_4666 );
and ( \2210_b0 , \2082_b0 , w_4667 );
and ( w_4666 , w_4667 , \2090_b0 );
or ( \2212_b1 , \2207_b1 , \2211_b1 );
xor ( \2212_b0 , \2207_b0 , w_4668 );
not ( w_4668 , w_4669 );
and ( w_4669 , \2211_b1 , \2211_b0 );
or ( \2213_b1 , \1351_b1 , \1382_b1 );
not ( \1382_b1 , w_4670 );
and ( \2213_b0 , \1351_b0 , w_4671 );
and ( w_4670 , w_4671 , \1382_b0 );
or ( \2214_b1 , \1446_b1 , \1380_b1 );
not ( \1380_b1 , w_4672 );
and ( \2214_b0 , \1446_b0 , w_4673 );
and ( w_4672 , w_4673 , \1380_b0 );
or ( \2215_b1 , \2213_b1 , w_4675 );
not ( w_4675 , w_4676 );
and ( \2215_b0 , \2213_b0 , w_4677 );
and ( w_4676 ,  , w_4677 );
buf ( w_4675 , \2214_b1 );
not ( w_4675 , w_4678 );
not (  , w_4679 );
and ( w_4678 , w_4679 , \2214_b0 );
or ( \2216_b1 , \2215_b1 , w_4680 );
xor ( \2216_b0 , \2215_b0 , w_4682 );
not ( w_4682 , w_4683 );
and ( w_4683 , w_4680 , w_4681 );
buf ( w_4680 , \1389_b1 );
not ( w_4680 , w_4684 );
not ( w_4681 , w_4685 );
and ( w_4684 , w_4685 , \1389_b0 );
or ( \2217_b1 , \1384_b1 , \1460_b1 );
not ( \1460_b1 , w_4686 );
and ( \2217_b0 , \1384_b0 , w_4687 );
and ( w_4686 , w_4687 , \1460_b0 );
or ( \2218_b1 , \1342_b1 , \1458_b1 );
not ( \1458_b1 , w_4688 );
and ( \2218_b0 , \1342_b0 , w_4689 );
and ( w_4688 , w_4689 , \1458_b0 );
or ( \2219_b1 , \2217_b1 , w_4691 );
not ( w_4691 , w_4692 );
and ( \2219_b0 , \2217_b0 , w_4693 );
and ( w_4692 ,  , w_4693 );
buf ( w_4691 , \2218_b1 );
not ( w_4691 , w_4694 );
not (  , w_4695 );
and ( w_4694 , w_4695 , \2218_b0 );
or ( \2220_b1 , \2219_b1 , w_4696 );
xor ( \2220_b0 , \2219_b0 , w_4698 );
not ( w_4698 , w_4699 );
and ( w_4699 , w_4696 , w_4697 );
buf ( w_4696 , \1467_b1 );
not ( w_4696 , w_4700 );
not ( w_4697 , w_4701 );
and ( w_4700 , w_4701 , \1467_b0 );
or ( \2221_b1 , \2216_b1 , \2220_b1 );
xor ( \2221_b0 , \2216_b0 , w_4702 );
not ( w_4702 , w_4703 );
and ( w_4703 , \2220_b1 , \2220_b0 );
or ( \2222_b1 , \1416_b1 , \1643_b1 );
not ( \1643_b1 , w_4704 );
and ( \2222_b0 , \1416_b0 , w_4705 );
and ( w_4704 , w_4705 , \1643_b0 );
or ( \2223_b1 , \1586_b1 , \1641_b1 );
not ( \1641_b1 , w_4706 );
and ( \2223_b0 , \1586_b0 , w_4707 );
and ( w_4706 , w_4707 , \1641_b0 );
or ( \2224_b1 , \2222_b1 , w_4709 );
not ( w_4709 , w_4710 );
and ( \2224_b0 , \2222_b0 , w_4711 );
and ( w_4710 ,  , w_4711 );
buf ( w_4709 , \2223_b1 );
not ( w_4709 , w_4712 );
not (  , w_4713 );
and ( w_4712 , w_4713 , \2223_b0 );
or ( \2225_b1 , \2224_b1 , w_4714 );
xor ( \2225_b0 , \2224_b0 , w_4716 );
not ( w_4716 , w_4717 );
and ( w_4717 , w_4714 , w_4715 );
buf ( w_4714 , \1649_b1 );
not ( w_4714 , w_4718 );
not ( w_4715 , w_4719 );
and ( w_4718 , w_4719 , \1649_b0 );
or ( \2226_b1 , \2221_b1 , \2225_b1 );
xor ( \2226_b0 , \2221_b0 , w_4720 );
not ( w_4720 , w_4721 );
and ( w_4721 , \2225_b1 , \2225_b0 );
or ( \2227_b1 , \2023_b1 , \1336_b1 );
not ( \1336_b1 , w_4722 );
and ( \2227_b0 , \2023_b0 , w_4723 );
and ( w_4722 , w_4723 , \1336_b0 );
buf ( \2228_b1 , \1175_A[31]_b1 );
buf ( \2228_b0 , \1175_A[31]_b0 );
or ( \2229_b1 , \2228_b1 , \1333_b1 );
not ( \1333_b1 , w_4724 );
and ( \2229_b0 , \2228_b0 , w_4725 );
and ( w_4724 , w_4725 , \1333_b0 );
or ( \2230_b1 , \2227_b1 , w_4727 );
not ( w_4727 , w_4728 );
and ( \2230_b0 , \2227_b0 , w_4729 );
and ( w_4728 ,  , w_4729 );
buf ( w_4727 , \2229_b1 );
not ( w_4727 , w_4730 );
not (  , w_4731 );
and ( w_4730 , w_4731 , \2229_b0 );
or ( \2231_b1 , \2230_b1 , w_4732 );
xor ( \2231_b0 , \2230_b0 , w_4734 );
not ( w_4734 , w_4735 );
and ( w_4735 , w_4732 , w_4733 );
buf ( w_4732 , \1332_b1 );
not ( w_4732 , w_4736 );
not ( w_4733 , w_4737 );
and ( w_4736 , w_4737 , \1332_b0 );
buf ( \2232_b1 , \2090_b1 );
not ( \2232_b1 , w_4738 );
not ( \2232_b0 , w_4739 );
and ( w_4738 , w_4739 , \2090_b0 );
buf ( \2233_b1 , \1299_B[31]_b1 );
buf ( \2233_b0 , \1299_B[31]_b0 );
or ( \2234_b1 , \2088_b1 , \1548_b1 );
not ( \1548_b1 , w_4740 );
and ( \2234_b0 , \2088_b0 , w_4741 );
and ( w_4740 , w_4741 , \1548_b0 );
buf ( \2235_b1 , \2234_b1 );
not ( \2235_b1 , w_4742 );
not ( \2235_b0 , w_4743 );
and ( w_4742 , w_4743 , \2234_b0 );
or ( \2236_b1 , \2233_b1 , \2235_b1 );
not ( \2235_b1 , w_4744 );
and ( \2236_b0 , \2233_b0 , w_4745 );
and ( w_4744 , w_4745 , \2235_b0 );
or ( \2237_b1 , \2232_b1 , \2236_b1 );
not ( \2236_b1 , w_4746 );
and ( \2237_b0 , \2232_b0 , w_4747 );
and ( w_4746 , w_4747 , \2236_b0 );
or ( \2238_b1 , \2231_b1 , \2237_b1 );
xor ( \2238_b0 , \2231_b0 , w_4748 );
not ( w_4748 , w_4749 );
and ( w_4749 , \2237_b1 , \2237_b0 );
or ( \2239_b1 , \2233_b1 , \2088_b1 );
xor ( \2239_b0 , \2233_b0 , w_4750 );
not ( w_4750 , w_4751 );
and ( w_4751 , \2088_b1 , \2088_b0 );
buf ( \2240_b1 , \2089_b1 );
not ( \2240_b1 , w_4752 );
not ( \2240_b0 , w_4753 );
and ( w_4752 , w_4753 , \2089_b0 );
or ( \2241_b1 , \2239_b1 , \2240_b1 );
not ( \2240_b1 , w_4754 );
and ( \2241_b0 , \2239_b0 , w_4755 );
and ( w_4754 , w_4755 , \2240_b0 );
or ( \2242_b1 , \1498_b1 , \2241_b1 );
not ( \2241_b1 , w_4756 );
and ( \2242_b0 , \1498_b0 , w_4757 );
and ( w_4756 , w_4757 , \2241_b0 );
or ( \2243_b1 , \1553_b1 , \2089_b1 );
not ( \2089_b1 , w_4758 );
and ( \2243_b0 , \1553_b0 , w_4759 );
and ( w_4758 , w_4759 , \2089_b0 );
or ( \2244_b1 , \2242_b1 , w_4761 );
not ( w_4761 , w_4762 );
and ( \2244_b0 , \2242_b0 , w_4763 );
and ( w_4762 ,  , w_4763 );
buf ( w_4761 , \2243_b1 );
not ( w_4761 , w_4764 );
not (  , w_4765 );
and ( w_4764 , w_4765 , \2243_b0 );
or ( \2245_b1 , \2244_b1 , w_4766 );
xor ( \2245_b0 , \2244_b0 , w_4768 );
not ( w_4768 , w_4769 );
and ( w_4769 , w_4766 , w_4767 );
buf ( w_4766 , \2236_b1 );
not ( w_4766 , w_4770 );
not ( w_4767 , w_4771 );
and ( w_4770 , w_4771 , \2236_b0 );
or ( \2246_b1 , \2238_b1 , \2245_b1 );
xor ( \2246_b0 , \2238_b0 , w_4772 );
not ( w_4772 , w_4773 );
and ( w_4773 , \2245_b1 , \2245_b0 );
or ( \2247_b1 , \2226_b1 , \2246_b1 );
xor ( \2247_b0 , \2226_b0 , w_4774 );
not ( w_4774 , w_4775 );
and ( w_4775 , \2246_b1 , \2246_b0 );
or ( \2248_b1 , \2212_b1 , \2247_b1 );
xor ( \2248_b0 , \2212_b0 , w_4776 );
not ( w_4776 , w_4777 );
and ( w_4777 , \2247_b1 , \2247_b0 );
or ( \2249_b1 , \2203_b1 , \2248_b1 );
xor ( \2249_b0 , \2203_b0 , w_4778 );
not ( w_4778 , w_4779 );
and ( w_4779 , \2248_b1 , \2248_b0 );
or ( \2250_b1 , \2194_b1 , \2249_b1 );
xor ( \2250_b0 , \2194_b0 , w_4780 );
not ( w_4780 , w_4781 );
and ( w_4781 , \2249_b1 , \2249_b0 );
or ( \2251_b1 , \2185_b1 , \2250_b1 );
xor ( \2251_b0 , \2185_b0 , w_4782 );
not ( w_4782 , w_4783 );
and ( w_4783 , \2250_b1 , \2250_b0 );
or ( \2252_b1 , \2101_b1 , \2251_b1 );
xor ( \2252_b0 , \2101_b0 , w_4784 );
not ( w_4784 , w_4785 );
and ( w_4785 , \2251_b1 , \2251_b0 );
or ( \2253_b1 , \2013_b1 , \2094_b1 );
xor ( \2253_b0 , \2013_b0 , w_4786 );
not ( w_4786 , w_4787 );
and ( w_4787 , \2094_b1 , \2094_b0 );
or ( \2254_b1 , \2253_b1 , \2097_b1 );
xor ( \2254_b0 , \2253_b0 , w_4788 );
not ( w_4788 , w_4789 );
and ( w_4789 , \2097_b1 , \2097_b0 );
or ( \2255_b1 , \1665_b1 , \1669_b1 );
xor ( \2255_b0 , \1665_b0 , w_4790 );
not ( w_4790 , w_4791 );
and ( w_4791 , \1669_b1 , \1669_b0 );
or ( \2256_b1 , \2255_b1 , \1682_b1 );
xor ( \2256_b0 , \2255_b0 , w_4792 );
not ( w_4792 , w_4793 );
and ( w_4793 , \1682_b1 , \1682_b0 );
or ( \2257_b1 , \1614_b1 , \1619_b1 );
xor ( \2257_b0 , \1614_b0 , w_4794 );
not ( w_4794 , w_4795 );
and ( w_4795 , \1619_b1 , \1619_b0 );
or ( \2258_b1 , \2257_b1 , \1625_b1 );
xor ( \2258_b0 , \2257_b0 , w_4796 );
not ( w_4796 , w_4797 );
and ( w_4797 , \1625_b1 , \1625_b0 );
or ( \2259_b1 , \2256_b1 , \2258_b1 );
not ( \2258_b1 , w_4798 );
and ( \2259_b0 , \2256_b0 , w_4799 );
and ( w_4798 , w_4799 , \2258_b0 );
or ( \2260_b1 , \1638_b1 , \1650_b1 );
xor ( \2260_b0 , \1638_b0 , w_4800 );
not ( w_4800 , w_4801 );
and ( w_4801 , \1650_b1 , \1650_b0 );
or ( \2261_b1 , \2260_b1 , \1655_b1 );
xor ( \2261_b0 , \2260_b0 , w_4802 );
not ( w_4802 , w_4803 );
and ( w_4803 , \1655_b1 , \1655_b0 );
or ( \2262_b1 , \2258_b1 , \2261_b1 );
not ( \2261_b1 , w_4804 );
and ( \2262_b0 , \2258_b0 , w_4805 );
and ( w_4804 , w_4805 , \2261_b0 );
or ( \2263_b1 , \2256_b1 , \2261_b1 );
not ( \2261_b1 , w_4806 );
and ( \2263_b0 , \2256_b0 , w_4807 );
and ( w_4806 , w_4807 , \2261_b0 );
or ( \2265_b1 , \1685_b1 , \1699_b1 );
xor ( \2265_b0 , \1685_b0 , w_4808 );
not ( w_4808 , w_4809 );
and ( w_4809 , \1699_b1 , \1699_b0 );
or ( \2266_b1 , \2265_b1 , \1714_b1 );
xor ( \2266_b0 , \2265_b0 , w_4810 );
not ( w_4810 , w_4811 );
and ( w_4811 , \1714_b1 , \1714_b0 );
or ( \2267_b1 , \2264_b1 , \2266_b1 );
not ( \2266_b1 , w_4812 );
and ( \2267_b0 , \2264_b0 , w_4813 );
and ( w_4812 , w_4813 , \2266_b0 );
or ( \2268_b1 , \1903_b1 , \1905_b1 );
xor ( \2268_b0 , \1903_b0 , w_4814 );
not ( w_4814 , w_4815 );
and ( w_4815 , \1905_b1 , \1905_b0 );
or ( \2269_b1 , \2268_b1 , \1908_b1 );
xor ( \2269_b0 , \2268_b0 , w_4816 );
not ( w_4816 , w_4817 );
and ( w_4817 , \1908_b1 , \1908_b0 );
or ( \2270_b1 , \2266_b1 , \2269_b1 );
not ( \2269_b1 , w_4818 );
and ( \2270_b0 , \2266_b0 , w_4819 );
and ( w_4818 , w_4819 , \2269_b0 );
or ( \2271_b1 , \2264_b1 , \2269_b1 );
not ( \2269_b1 , w_4820 );
and ( \2271_b0 , \2264_b0 , w_4821 );
and ( w_4820 , w_4821 , \2269_b0 );
or ( \2273_b1 , \1661_b1 , \1717_b1 );
xor ( \2273_b0 , \1661_b0 , w_4822 );
not ( w_4822 , w_4823 );
and ( w_4823 , \1717_b1 , \1717_b0 );
or ( \2274_b1 , \2273_b1 , \1741_b1 );
xor ( \2274_b0 , \2273_b0 , w_4824 );
not ( w_4824 , w_4825 );
and ( w_4825 , \1741_b1 , \1741_b0 );
or ( \2275_b1 , \2272_b1 , \2274_b1 );
not ( \2274_b1 , w_4826 );
and ( \2275_b0 , \2272_b0 , w_4827 );
and ( w_4826 , w_4827 , \2274_b0 );
or ( \2276_b1 , \1769_b1 , \1783_b1 );
xor ( \2276_b0 , \1769_b0 , w_4828 );
not ( w_4828 , w_4829 );
and ( w_4829 , \1783_b1 , \1783_b0 );
or ( \2277_b1 , \2276_b1 , \1806_b1 );
xor ( \2277_b0 , \2276_b0 , w_4830 );
not ( w_4830 , w_4831 );
and ( w_4831 , \1806_b1 , \1806_b0 );
or ( \2278_b1 , \2274_b1 , \2277_b1 );
not ( \2277_b1 , w_4832 );
and ( \2278_b0 , \2274_b0 , w_4833 );
and ( w_4832 , w_4833 , \2277_b0 );
or ( \2279_b1 , \2272_b1 , \2277_b1 );
not ( \2277_b1 , w_4834 );
and ( \2279_b0 , \2272_b0 , w_4835 );
and ( w_4834 , w_4835 , \2277_b0 );
or ( \2281_b1 , \1744_b1 , \1809_b1 );
xor ( \2281_b0 , \1744_b0 , w_4836 );
not ( w_4836 , w_4837 );
and ( w_4837 , \1809_b1 , \1809_b0 );
or ( \2282_b1 , \2281_b1 , \1835_b1 );
xor ( \2282_b0 , \2281_b0 , w_4838 );
not ( w_4838 , w_4839 );
and ( w_4839 , \1835_b1 , \1835_b0 );
or ( \2283_b1 , \2280_b1 , \2282_b1 );
not ( \2282_b1 , w_4840 );
and ( \2283_b0 , \2280_b0 , w_4841 );
and ( w_4840 , w_4841 , \2282_b0 );
or ( \2284_b1 , \1995_b1 , \2007_b1 );
xor ( \2284_b0 , \1995_b0 , w_4842 );
not ( w_4842 , w_4843 );
and ( w_4843 , \2007_b1 , \2007_b0 );
or ( \2285_b1 , \2284_b1 , \2010_b1 );
xor ( \2285_b0 , \2284_b0 , w_4844 );
not ( w_4844 , w_4845 );
and ( w_4845 , \2010_b1 , \2010_b0 );
or ( \2286_b1 , \2282_b1 , \2285_b1 );
not ( \2285_b1 , w_4846 );
and ( \2286_b0 , \2282_b0 , w_4847 );
and ( w_4846 , w_4847 , \2285_b0 );
or ( \2287_b1 , \2280_b1 , \2285_b1 );
not ( \2285_b1 , w_4848 );
and ( \2287_b0 , \2280_b0 , w_4849 );
and ( w_4848 , w_4849 , \2285_b0 );
or ( \2289_b1 , \2254_b1 , \2288_b1 );
not ( \2288_b1 , w_4850 );
and ( \2289_b0 , \2254_b0 , w_4851 );
and ( w_4850 , w_4851 , \2288_b0 );
or ( \2290_b1 , \2254_b1 , \2288_b1 );
xor ( \2290_b0 , \2254_b0 , w_4852 );
not ( w_4852 , w_4853 );
and ( w_4853 , \2288_b1 , \2288_b0 );
or ( \2291_b1 , \1342_b1 , \1431_b1 );
not ( \1431_b1 , w_4854 );
and ( \2291_b0 , \1342_b0 , w_4855 );
and ( w_4854 , w_4855 , \1431_b0 );
or ( \2292_b1 , \1351_b1 , \1429_b1 );
not ( \1429_b1 , w_4856 );
and ( \2292_b0 , \1351_b0 , w_4857 );
and ( w_4856 , w_4857 , \1429_b0 );
or ( \2293_b1 , \2291_b1 , w_4859 );
not ( w_4859 , w_4860 );
and ( \2293_b0 , \2291_b0 , w_4861 );
and ( w_4860 ,  , w_4861 );
buf ( w_4859 , \2292_b1 );
not ( w_4859 , w_4862 );
not (  , w_4863 );
and ( w_4862 , w_4863 , \2292_b0 );
or ( \2294_b1 , \2293_b1 , w_4864 );
xor ( \2294_b0 , \2293_b0 , w_4866 );
not ( w_4866 , w_4867 );
and ( w_4867 , w_4864 , w_4865 );
buf ( w_4864 , \1438_b1 );
not ( w_4864 , w_4868 );
not ( w_4865 , w_4869 );
and ( w_4868 , w_4869 , \1438_b0 );
or ( \2295_b1 , \1376_b1 , \1444_b1 );
not ( \1444_b1 , w_4870 );
and ( \2295_b0 , \1376_b0 , w_4871 );
and ( w_4870 , w_4871 , \1444_b0 );
or ( \2296_b1 , \1384_b1 , \1442_b1 );
not ( \1442_b1 , w_4872 );
and ( \2296_b0 , \1384_b0 , w_4873 );
and ( w_4872 , w_4873 , \1442_b0 );
or ( \2297_b1 , \2295_b1 , w_4875 );
not ( w_4875 , w_4876 );
and ( \2297_b0 , \2295_b0 , w_4877 );
and ( w_4876 ,  , w_4877 );
buf ( w_4875 , \2296_b1 );
not ( w_4875 , w_4878 );
not (  , w_4879 );
and ( w_4878 , w_4879 , \2296_b0 );
or ( \2298_b1 , \2297_b1 , w_4880 );
xor ( \2298_b0 , \2297_b0 , w_4882 );
not ( w_4882 , w_4883 );
and ( w_4883 , w_4880 , w_4881 );
buf ( w_4880 , \1451_b1 );
not ( w_4880 , w_4884 );
not ( w_4881 , w_4885 );
and ( w_4884 , w_4885 , \1451_b0 );
or ( \2299_b1 , \2294_b1 , \2298_b1 );
not ( \2298_b1 , w_4886 );
and ( \2299_b0 , \2294_b0 , w_4887 );
and ( w_4886 , w_4887 , \2298_b0 );
or ( \2300_b1 , \2298_b1 , \1921_b1 );
not ( \1921_b1 , w_4888 );
and ( \2300_b0 , \2298_b0 , w_4889 );
and ( w_4888 , w_4889 , \1921_b0 );
or ( \2301_b1 , \2294_b1 , \1921_b1 );
not ( \1921_b1 , w_4890 );
and ( \2301_b0 , \2294_b0 , w_4891 );
and ( w_4890 , w_4891 , \1921_b0 );
or ( \2303_b1 , \1446_b1 , \1336_b1 );
not ( \1336_b1 , w_4892 );
and ( \2303_b0 , \1446_b0 , w_4893 );
and ( w_4892 , w_4893 , \1336_b0 );
or ( \2304_b1 , \1425_b1 , \1333_b1 );
not ( \1333_b1 , w_4894 );
and ( \2304_b0 , \1425_b0 , w_4895 );
and ( w_4894 , w_4895 , \1333_b0 );
or ( \2305_b1 , \2303_b1 , w_4897 );
not ( w_4897 , w_4898 );
and ( \2305_b0 , \2303_b0 , w_4899 );
and ( w_4898 ,  , w_4899 );
buf ( w_4897 , \2304_b1 );
not ( w_4897 , w_4900 );
not (  , w_4901 );
and ( w_4900 , w_4901 , \2304_b0 );
or ( \2306_b1 , \2305_b1 , w_4902 );
xor ( \2306_b0 , \2305_b0 , w_4904 );
not ( w_4904 , w_4905 );
and ( w_4905 , w_4902 , w_4903 );
buf ( w_4902 , \1332_b1 );
not ( w_4902 , w_4906 );
not ( w_4903 , w_4907 );
and ( w_4906 , w_4907 , \1332_b0 );
or ( \2307_b1 , \1454_b1 , \1349_b1 );
not ( \1349_b1 , w_4908 );
and ( \2307_b0 , \1454_b0 , w_4909 );
and ( w_4908 , w_4909 , \1349_b0 );
or ( \2308_b1 , \1462_b1 , \1347_b1 );
not ( \1347_b1 , w_4910 );
and ( \2308_b0 , \1462_b0 , w_4911 );
and ( w_4910 , w_4911 , \1347_b0 );
or ( \2309_b1 , \2307_b1 , w_4913 );
not ( w_4913 , w_4914 );
and ( \2309_b0 , \2307_b0 , w_4915 );
and ( w_4914 ,  , w_4915 );
buf ( w_4913 , \2308_b1 );
not ( w_4913 , w_4916 );
not (  , w_4917 );
and ( w_4916 , w_4917 , \2308_b0 );
or ( \2310_b1 , \2309_b1 , w_4918 );
xor ( \2310_b0 , \2309_b0 , w_4920 );
not ( w_4920 , w_4921 );
and ( w_4921 , w_4918 , w_4919 );
buf ( w_4918 , \1356_b1 );
not ( w_4918 , w_4922 );
not ( w_4919 , w_4923 );
and ( w_4922 , w_4923 , \1356_b0 );
or ( \2311_b1 , \2306_b1 , \2310_b1 );
not ( \2310_b1 , w_4924 );
and ( \2311_b0 , \2306_b0 , w_4925 );
and ( w_4924 , w_4925 , \2310_b0 );
or ( \2312_b1 , \1586_b1 , \1366_b1 );
not ( \1366_b1 , w_4926 );
and ( \2312_b0 , \1586_b0 , w_4927 );
and ( w_4926 , w_4927 , \1366_b0 );
or ( \2313_b1 , \1616_b1 , \1364_b1 );
not ( \1364_b1 , w_4928 );
and ( \2313_b0 , \1616_b0 , w_4929 );
and ( w_4928 , w_4929 , \1364_b0 );
or ( \2314_b1 , \2312_b1 , w_4931 );
not ( w_4931 , w_4932 );
and ( \2314_b0 , \2312_b0 , w_4933 );
and ( w_4932 ,  , w_4933 );
buf ( w_4931 , \2313_b1 );
not ( w_4931 , w_4934 );
not (  , w_4935 );
and ( w_4934 , w_4935 , \2313_b0 );
or ( \2315_b1 , \2314_b1 , w_4936 );
xor ( \2315_b0 , \2314_b0 , w_4938 );
not ( w_4938 , w_4939 );
and ( w_4939 , w_4936 , w_4937 );
buf ( w_4936 , \1373_b1 );
not ( w_4936 , w_4940 );
not ( w_4937 , w_4941 );
and ( w_4940 , w_4941 , \1373_b0 );
or ( \2316_b1 , \2310_b1 , \2315_b1 );
not ( \2315_b1 , w_4942 );
and ( \2316_b0 , \2310_b0 , w_4943 );
and ( w_4942 , w_4943 , \2315_b0 );
or ( \2317_b1 , \2306_b1 , \2315_b1 );
not ( \2315_b1 , w_4944 );
and ( \2317_b0 , \2306_b0 , w_4945 );
and ( w_4944 , w_4945 , \2315_b0 );
or ( \2319_b1 , \2302_b1 , \2318_b1 );
not ( \2318_b1 , w_4946 );
and ( \2319_b0 , \2302_b0 , w_4947 );
and ( w_4946 , w_4947 , \2318_b0 );
or ( \2320_b1 , \1498_b1 , \1524_b1 );
not ( \1524_b1 , w_4948 );
and ( \2320_b0 , \1498_b0 , w_4949 );
and ( w_4948 , w_4949 , \1524_b0 );
or ( \2321_b1 , \1553_b1 , \1522_b1 );
not ( \1522_b1 , w_4950 );
and ( \2321_b0 , \1553_b0 , w_4951 );
and ( w_4950 , w_4951 , \1522_b0 );
or ( \2322_b1 , \2320_b1 , w_4953 );
not ( w_4953 , w_4954 );
and ( \2322_b0 , \2320_b0 , w_4955 );
and ( w_4954 ,  , w_4955 );
buf ( w_4953 , \2321_b1 );
not ( w_4953 , w_4956 );
not (  , w_4957 );
and ( w_4956 , w_4957 , \2321_b0 );
or ( \2323_b1 , \2322_b1 , w_4958 );
xor ( \2323_b0 , \2322_b0 , w_4960 );
not ( w_4960 , w_4961 );
and ( w_4961 , w_4958 , w_4959 );
buf ( w_4958 , \1531_b1 );
not ( w_4958 , w_4962 );
not ( w_4959 , w_4963 );
and ( w_4962 , w_4963 , \1531_b0 );
or ( \2324_b1 , \2318_b1 , \2323_b1 );
not ( \2323_b1 , w_4964 );
and ( \2324_b0 , \2318_b0 , w_4965 );
and ( w_4964 , w_4965 , \2323_b0 );
or ( \2325_b1 , \2302_b1 , \2323_b1 );
not ( \2323_b1 , w_4966 );
and ( \2325_b0 , \2302_b0 , w_4967 );
and ( w_4966 , w_4967 , \2323_b0 );
or ( \2327_b1 , \1470_b1 , \1382_b1 );
not ( \1382_b1 , w_4968 );
and ( \2327_b0 , \1470_b0 , w_4969 );
and ( w_4968 , w_4969 , \1382_b0 );
or ( \2328_b1 , \1477_b1 , \1380_b1 );
not ( \1380_b1 , w_4970 );
and ( \2328_b0 , \1477_b0 , w_4971 );
and ( w_4970 , w_4971 , \1380_b0 );
or ( \2329_b1 , \2327_b1 , w_4973 );
not ( w_4973 , w_4974 );
and ( \2329_b0 , \2327_b0 , w_4975 );
and ( w_4974 ,  , w_4975 );
buf ( w_4973 , \2328_b1 );
not ( w_4973 , w_4976 );
not (  , w_4977 );
and ( w_4976 , w_4977 , \2328_b0 );
or ( \2330_b1 , \2329_b1 , w_4978 );
xor ( \2330_b0 , \2329_b0 , w_4980 );
not ( w_4980 , w_4981 );
and ( w_4981 , w_4978 , w_4979 );
buf ( w_4978 , \1389_b1 );
not ( w_4978 , w_4982 );
not ( w_4979 , w_4983 );
and ( w_4982 , w_4983 , \1389_b0 );
or ( \2331_b1 , \1407_b1 , \1397_b1 );
not ( \1397_b1 , w_4984 );
and ( \2331_b0 , \1407_b0 , w_4985 );
and ( w_4984 , w_4985 , \1397_b0 );
or ( \2332_b1 , \1416_b1 , \1395_b1 );
not ( \1395_b1 , w_4986 );
and ( \2332_b0 , \1416_b0 , w_4987 );
and ( w_4986 , w_4987 , \1395_b0 );
or ( \2333_b1 , \2331_b1 , w_4989 );
not ( w_4989 , w_4990 );
and ( \2333_b0 , \2331_b0 , w_4991 );
and ( w_4990 ,  , w_4991 );
buf ( w_4989 , \2332_b1 );
not ( w_4989 , w_4992 );
not (  , w_4993 );
and ( w_4992 , w_4993 , \2332_b0 );
or ( \2334_b1 , \2333_b1 , w_4994 );
xor ( \2334_b0 , \2333_b0 , w_4996 );
not ( w_4996 , w_4997 );
and ( w_4997 , w_4994 , w_4995 );
buf ( w_4994 , \1404_b1 );
not ( w_4994 , w_4998 );
not ( w_4995 , w_4999 );
and ( w_4998 , w_4999 , \1404_b0 );
or ( \2335_b1 , \2330_b1 , \2334_b1 );
not ( \2334_b1 , w_5000 );
and ( \2335_b0 , \2330_b0 , w_5001 );
and ( w_5000 , w_5001 , \2334_b0 );
or ( \2336_b1 , \1540_b1 , \1414_b1 );
not ( \1414_b1 , w_5002 );
and ( \2336_b0 , \1540_b0 , w_5003 );
and ( w_5002 , w_5003 , \1414_b0 );
or ( \2337_b1 , \1517_b1 , \1412_b1 );
not ( \1412_b1 , w_5004 );
and ( \2337_b0 , \1517_b0 , w_5005 );
and ( w_5004 , w_5005 , \1412_b0 );
or ( \2338_b1 , \2336_b1 , w_5007 );
not ( w_5007 , w_5008 );
and ( \2338_b0 , \2336_b0 , w_5009 );
and ( w_5008 ,  , w_5009 );
buf ( w_5007 , \2337_b1 );
not ( w_5007 , w_5010 );
not (  , w_5011 );
and ( w_5010 , w_5011 , \2337_b0 );
or ( \2339_b1 , \2338_b1 , w_5012 );
xor ( \2339_b0 , \2338_b0 , w_5014 );
not ( w_5014 , w_5015 );
and ( w_5015 , w_5012 , w_5013 );
buf ( w_5012 , \1421_b1 );
not ( w_5012 , w_5016 );
not ( w_5013 , w_5017 );
and ( w_5016 , w_5017 , \1421_b0 );
or ( \2340_b1 , \2334_b1 , \2339_b1 );
not ( \2339_b1 , w_5018 );
and ( \2340_b0 , \2334_b0 , w_5019 );
and ( w_5018 , w_5019 , \2339_b0 );
or ( \2341_b1 , \2330_b1 , \2339_b1 );
not ( \2339_b1 , w_5020 );
and ( \2341_b0 , \2330_b0 , w_5021 );
and ( w_5020 , w_5021 , \2339_b0 );
or ( \2343_b1 , \1359_b1 , \1460_b1 );
not ( \1460_b1 , w_5022 );
and ( \2343_b0 , \1359_b0 , w_5023 );
and ( w_5022 , w_5023 , \1460_b0 );
or ( \2344_b1 , \1368_b1 , \1458_b1 );
not ( \1458_b1 , w_5024 );
and ( \2344_b0 , \1368_b0 , w_5025 );
and ( w_5024 , w_5025 , \1458_b0 );
or ( \2345_b1 , \2343_b1 , w_5027 );
not ( w_5027 , w_5028 );
and ( \2345_b0 , \2343_b0 , w_5029 );
and ( w_5028 ,  , w_5029 );
buf ( w_5027 , \2344_b1 );
not ( w_5027 , w_5030 );
not (  , w_5031 );
and ( w_5030 , w_5031 , \2344_b0 );
or ( \2346_b1 , \2345_b1 , w_5032 );
xor ( \2346_b0 , \2345_b0 , w_5034 );
not ( w_5034 , w_5035 );
and ( w_5035 , w_5032 , w_5033 );
buf ( w_5032 , \1467_b1 );
not ( w_5032 , w_5036 );
not ( w_5033 , w_5037 );
and ( w_5036 , w_5037 , \1467_b0 );
or ( \2347_b1 , \1391_b1 , \1475_b1 );
not ( \1475_b1 , w_5038 );
and ( \2347_b0 , \1391_b0 , w_5039 );
and ( w_5038 , w_5039 , \1475_b0 );
or ( \2348_b1 , \1399_b1 , \1473_b1 );
not ( \1473_b1 , w_5040 );
and ( \2348_b0 , \1399_b0 , w_5041 );
and ( w_5040 , w_5041 , \1473_b0 );
or ( \2349_b1 , \2347_b1 , w_5043 );
not ( w_5043 , w_5044 );
and ( \2349_b0 , \2347_b0 , w_5045 );
and ( w_5044 ,  , w_5045 );
buf ( w_5043 , \2348_b1 );
not ( w_5043 , w_5046 );
not (  , w_5047 );
and ( w_5046 , w_5047 , \2348_b0 );
or ( \2350_b1 , \2349_b1 , w_5048 );
xor ( \2350_b0 , \2349_b0 , w_5050 );
not ( w_5050 , w_5051 );
and ( w_5051 , w_5048 , w_5049 );
buf ( w_5048 , \1482_b1 );
not ( w_5048 , w_5052 );
not ( w_5049 , w_5053 );
and ( w_5052 , w_5053 , \1482_b0 );
or ( \2351_b1 , \2346_b1 , \2350_b1 );
not ( \2350_b1 , w_5054 );
and ( \2351_b0 , \2346_b0 , w_5055 );
and ( w_5054 , w_5055 , \2350_b0 );
or ( \2352_b1 , \1526_b1 , \1675_b1 );
not ( \1675_b1 , w_5056 );
and ( \2352_b0 , \1526_b0 , w_5057 );
and ( w_5056 , w_5057 , \1675_b0 );
or ( \2353_b1 , \1622_b1 , \1673_b1 );
not ( \1673_b1 , w_5058 );
and ( \2353_b0 , \1622_b0 , w_5059 );
and ( w_5058 , w_5059 , \1673_b0 );
or ( \2354_b1 , \2352_b1 , w_5061 );
not ( w_5061 , w_5062 );
and ( \2354_b0 , \2352_b0 , w_5063 );
and ( w_5062 ,  , w_5063 );
buf ( w_5061 , \2353_b1 );
not ( w_5061 , w_5064 );
not (  , w_5065 );
and ( w_5064 , w_5065 , \2353_b0 );
or ( \2355_b1 , \2354_b1 , w_5066 );
xor ( \2355_b0 , \2354_b0 , w_5068 );
not ( w_5068 , w_5069 );
and ( w_5069 , w_5066 , w_5067 );
buf ( w_5066 , \1681_b1 );
not ( w_5066 , w_5070 );
not ( w_5067 , w_5071 );
and ( w_5070 , w_5071 , \1681_b0 );
or ( \2356_b1 , \2350_b1 , \2355_b1 );
not ( \2355_b1 , w_5072 );
and ( \2356_b0 , \2350_b0 , w_5073 );
and ( w_5072 , w_5073 , \2355_b0 );
or ( \2357_b1 , \2346_b1 , \2355_b1 );
not ( \2355_b1 , w_5074 );
and ( \2357_b0 , \2346_b0 , w_5075 );
and ( w_5074 , w_5075 , \2355_b0 );
or ( \2359_b1 , \2342_b1 , \2358_b1 );
not ( \2358_b1 , w_5076 );
and ( \2359_b0 , \2342_b0 , w_5077 );
and ( w_5076 , w_5077 , \2358_b0 );
or ( \2360_b1 , \1915_b1 , \1919_b1 );
xor ( \2360_b0 , \1915_b0 , w_5078 );
not ( w_5078 , w_5079 );
and ( w_5079 , \1919_b1 , \1919_b0 );
or ( \2361_b1 , \2360_b1 , \1923_b1 );
xor ( \2361_b0 , \2360_b0 , w_5080 );
not ( w_5080 , w_5081 );
and ( w_5081 , \1923_b1 , \1923_b0 );
or ( \2362_b1 , \2358_b1 , \2361_b1 );
not ( \2361_b1 , w_5082 );
and ( \2362_b0 , \2358_b0 , w_5083 );
and ( w_5082 , w_5083 , \2361_b0 );
or ( \2363_b1 , \2342_b1 , \2361_b1 );
not ( \2361_b1 , w_5084 );
and ( \2363_b0 , \2342_b0 , w_5085 );
and ( w_5084 , w_5085 , \2361_b0 );
or ( \2365_b1 , \2326_b1 , \2364_b1 );
not ( \2364_b1 , w_5086 );
and ( \2365_b0 , \2326_b0 , w_5087 );
and ( w_5086 , w_5087 , \2364_b0 );
or ( \2366_b1 , \1926_b1 , \1942_b1 );
xor ( \2366_b0 , \1926_b0 , w_5088 );
not ( w_5088 , w_5089 );
and ( w_5089 , \1942_b1 , \1942_b0 );
or ( \2367_b1 , \2366_b1 , \1959_b1 );
xor ( \2367_b0 , \2366_b0 , w_5090 );
not ( w_5090 , w_5091 );
and ( w_5091 , \1959_b1 , \1959_b0 );
or ( \2368_b1 , \2364_b1 , \2367_b1 );
not ( \2367_b1 , w_5092 );
and ( \2368_b0 , \2364_b0 , w_5093 );
and ( w_5092 , w_5093 , \2367_b0 );
or ( \2369_b1 , \2326_b1 , \2367_b1 );
not ( \2367_b1 , w_5094 );
and ( \2369_b0 , \2326_b0 , w_5095 );
and ( w_5094 , w_5095 , \2367_b0 );
or ( \2371_b1 , \1930_b1 , \1934_b1 );
xor ( \2371_b0 , \1930_b0 , w_5096 );
not ( w_5096 , w_5097 );
and ( w_5097 , \1934_b1 , \1934_b0 );
or ( \2372_b1 , \2371_b1 , \1939_b1 );
xor ( \2372_b0 , \2371_b0 , w_5098 );
not ( w_5098 , w_5099 );
and ( w_5099 , \1939_b1 , \1939_b0 );
or ( \2373_b1 , \1947_b1 , \1951_b1 );
xor ( \2373_b0 , \1947_b0 , w_5100 );
not ( w_5100 , w_5101 );
and ( w_5101 , \1951_b1 , \1951_b0 );
or ( \2374_b1 , \2373_b1 , \1956_b1 );
xor ( \2374_b0 , \2373_b0 , w_5102 );
not ( w_5102 , w_5103 );
and ( w_5103 , \1956_b1 , \1956_b0 );
or ( \2375_b1 , \2372_b1 , \2374_b1 );
not ( \2374_b1 , w_5104 );
and ( \2375_b0 , \2372_b0 , w_5105 );
and ( w_5104 , w_5105 , \2374_b0 );
or ( \2376_b1 , \1963_b1 , \1967_b1 );
xor ( \2376_b0 , \1963_b0 , w_5106 );
not ( w_5106 , w_5107 );
and ( w_5107 , \1967_b1 , \1967_b0 );
or ( \2377_b1 , \2376_b1 , \1972_b1 );
xor ( \2377_b0 , \2376_b0 , w_5108 );
not ( w_5108 , w_5109 );
and ( w_5109 , \1972_b1 , \1972_b0 );
or ( \2378_b1 , \2374_b1 , \2377_b1 );
not ( \2377_b1 , w_5110 );
and ( \2378_b0 , \2374_b0 , w_5111 );
and ( w_5110 , w_5111 , \2377_b0 );
or ( \2379_b1 , \2372_b1 , \2377_b1 );
not ( \2377_b1 , w_5112 );
and ( \2379_b0 , \2372_b0 , w_5113 );
and ( w_5112 , w_5113 , \2377_b0 );
or ( \2381_b1 , \2256_b1 , \2258_b1 );
xor ( \2381_b0 , \2256_b0 , w_5114 );
not ( w_5114 , w_5115 );
and ( w_5115 , \2258_b1 , \2258_b0 );
or ( \2382_b1 , \2381_b1 , \2261_b1 );
xor ( \2382_b0 , \2381_b0 , w_5116 );
not ( w_5116 , w_5117 );
and ( w_5117 , \2261_b1 , \2261_b0 );
or ( \2383_b1 , \2380_b1 , \2382_b1 );
not ( \2382_b1 , w_5118 );
and ( \2383_b0 , \2380_b0 , w_5119 );
and ( w_5118 , w_5119 , \2382_b0 );
or ( \2384_b1 , \1975_b1 , \1977_b1 );
xor ( \2384_b0 , \1975_b0 , w_5120 );
not ( w_5120 , w_5121 );
and ( w_5121 , \1977_b1 , \1977_b0 );
or ( \2385_b1 , \2384_b1 , \1980_b1 );
xor ( \2385_b0 , \2384_b0 , w_5122 );
not ( w_5122 , w_5123 );
and ( w_5123 , \1980_b1 , \1980_b0 );
or ( \2386_b1 , \2382_b1 , \2385_b1 );
not ( \2385_b1 , w_5124 );
and ( \2386_b0 , \2382_b0 , w_5125 );
and ( w_5124 , w_5125 , \2385_b0 );
or ( \2387_b1 , \2380_b1 , \2385_b1 );
not ( \2385_b1 , w_5126 );
and ( \2387_b0 , \2380_b0 , w_5127 );
and ( w_5126 , w_5127 , \2385_b0 );
or ( \2389_b1 , \2370_b1 , \2388_b1 );
not ( \2388_b1 , w_5128 );
and ( \2389_b0 , \2370_b0 , w_5129 );
and ( w_5128 , w_5129 , \2388_b0 );
or ( \2390_b1 , \1962_b1 , \1983_b1 );
xor ( \2390_b0 , \1962_b0 , w_5130 );
not ( w_5130 , w_5131 );
and ( w_5131 , \1983_b1 , \1983_b0 );
or ( \2391_b1 , \2390_b1 , \1986_b1 );
xor ( \2391_b0 , \2390_b0 , w_5132 );
not ( w_5132 , w_5133 );
and ( w_5133 , \1986_b1 , \1986_b0 );
or ( \2392_b1 , \2388_b1 , \2391_b1 );
not ( \2391_b1 , w_5134 );
and ( \2392_b0 , \2388_b0 , w_5135 );
and ( w_5134 , w_5135 , \2391_b0 );
or ( \2393_b1 , \2370_b1 , \2391_b1 );
not ( \2391_b1 , w_5136 );
and ( \2393_b0 , \2370_b0 , w_5137 );
and ( w_5136 , w_5137 , \2391_b0 );
or ( \2395_b1 , \1911_b1 , \1989_b1 );
xor ( \2395_b0 , \1911_b0 , w_5138 );
not ( w_5138 , w_5139 );
and ( w_5139 , \1989_b1 , \1989_b0 );
or ( \2396_b1 , \2395_b1 , \1992_b1 );
xor ( \2396_b0 , \2395_b0 , w_5140 );
not ( w_5140 , w_5141 );
and ( w_5141 , \1992_b1 , \1992_b0 );
or ( \2397_b1 , \2394_b1 , \2396_b1 );
not ( \2396_b1 , w_5142 );
and ( \2397_b0 , \2394_b0 , w_5143 );
and ( w_5142 , w_5143 , \2396_b0 );
or ( \2398_b1 , \2272_b1 , \2274_b1 );
xor ( \2398_b0 , \2272_b0 , w_5144 );
not ( w_5144 , w_5145 );
and ( w_5145 , \2274_b1 , \2274_b0 );
or ( \2399_b1 , \2398_b1 , \2277_b1 );
xor ( \2399_b0 , \2398_b0 , w_5146 );
not ( w_5146 , w_5147 );
and ( w_5147 , \2277_b1 , \2277_b0 );
or ( \2400_b1 , \2396_b1 , \2399_b1 );
not ( \2399_b1 , w_5148 );
and ( \2400_b0 , \2396_b0 , w_5149 );
and ( w_5148 , w_5149 , \2399_b0 );
or ( \2401_b1 , \2394_b1 , \2399_b1 );
not ( \2399_b1 , w_5150 );
and ( \2401_b0 , \2394_b0 , w_5151 );
and ( w_5150 , w_5151 , \2399_b0 );
or ( \2403_b1 , \2280_b1 , \2282_b1 );
xor ( \2403_b0 , \2280_b0 , w_5152 );
not ( w_5152 , w_5153 );
and ( w_5153 , \2282_b1 , \2282_b0 );
or ( \2404_b1 , \2403_b1 , \2285_b1 );
xor ( \2404_b0 , \2403_b0 , w_5154 );
not ( w_5154 , w_5155 );
and ( w_5155 , \2285_b1 , \2285_b0 );
or ( \2405_b1 , \2402_b1 , \2404_b1 );
not ( \2404_b1 , w_5156 );
and ( \2405_b0 , \2402_b0 , w_5157 );
and ( w_5156 , w_5157 , \2404_b0 );
or ( \2406_b1 , \2402_b1 , \2404_b1 );
xor ( \2406_b0 , \2402_b0 , w_5158 );
not ( w_5158 , w_5159 );
and ( w_5159 , \2404_b1 , \2404_b0 );
or ( \2407_b1 , \2394_b1 , \2396_b1 );
xor ( \2407_b0 , \2394_b0 , w_5160 );
not ( w_5160 , w_5161 );
and ( w_5161 , \2396_b1 , \2396_b0 );
or ( \2408_b1 , \2407_b1 , \2399_b1 );
xor ( \2408_b0 , \2407_b0 , w_5162 );
not ( w_5162 , w_5163 );
and ( w_5163 , \2399_b1 , \2399_b0 );
or ( \2409_b1 , \1368_b1 , \1382_b1 );
not ( \1382_b1 , w_5164 );
and ( \2409_b0 , \1368_b0 , w_5165 );
and ( w_5164 , w_5165 , \1382_b0 );
or ( \2410_b1 , \1470_b1 , \1380_b1 );
not ( \1380_b1 , w_5166 );
and ( \2410_b0 , \1470_b0 , w_5167 );
and ( w_5166 , w_5167 , \1380_b0 );
or ( \2411_b1 , \2409_b1 , w_5169 );
not ( w_5169 , w_5170 );
and ( \2411_b0 , \2409_b0 , w_5171 );
and ( w_5170 ,  , w_5171 );
buf ( w_5169 , \2410_b1 );
not ( w_5169 , w_5172 );
not (  , w_5173 );
and ( w_5172 , w_5173 , \2410_b0 );
or ( \2412_b1 , \2411_b1 , w_5174 );
xor ( \2412_b0 , \2411_b0 , w_5176 );
not ( w_5176 , w_5177 );
and ( w_5177 , w_5174 , w_5175 );
buf ( w_5174 , \1389_b1 );
not ( w_5174 , w_5178 );
not ( w_5175 , w_5179 );
and ( w_5178 , w_5179 , \1389_b0 );
or ( \2413_b1 , \1416_b1 , \1366_b1 );
not ( \1366_b1 , w_5180 );
and ( \2413_b0 , \1416_b0 , w_5181 );
and ( w_5180 , w_5181 , \1366_b0 );
or ( \2414_b1 , \1586_b1 , \1364_b1 );
not ( \1364_b1 , w_5182 );
and ( \2414_b0 , \1586_b0 , w_5183 );
and ( w_5182 , w_5183 , \1364_b0 );
or ( \2415_b1 , \2413_b1 , w_5185 );
not ( w_5185 , w_5186 );
and ( \2415_b0 , \2413_b0 , w_5187 );
and ( w_5186 ,  , w_5187 );
buf ( w_5185 , \2414_b1 );
not ( w_5185 , w_5188 );
not (  , w_5189 );
and ( w_5188 , w_5189 , \2414_b0 );
or ( \2416_b1 , \2415_b1 , w_5190 );
xor ( \2416_b0 , \2415_b0 , w_5192 );
not ( w_5192 , w_5193 );
and ( w_5193 , w_5190 , w_5191 );
buf ( w_5190 , \1373_b1 );
not ( w_5190 , w_5194 );
not ( w_5191 , w_5195 );
and ( w_5194 , w_5195 , \1373_b0 );
or ( \2417_b1 , \2412_b1 , \2416_b1 );
not ( \2416_b1 , w_5196 );
and ( \2417_b0 , \2412_b0 , w_5197 );
and ( w_5196 , w_5197 , \2416_b0 );
or ( \2418_b1 , \1622_b1 , \1397_b1 );
not ( \1397_b1 , w_5198 );
and ( \2418_b0 , \1622_b0 , w_5199 );
and ( w_5198 , w_5199 , \1397_b0 );
or ( \2419_b1 , \1407_b1 , \1395_b1 );
not ( \1395_b1 , w_5200 );
and ( \2419_b0 , \1407_b0 , w_5201 );
and ( w_5200 , w_5201 , \1395_b0 );
or ( \2420_b1 , \2418_b1 , w_5203 );
not ( w_5203 , w_5204 );
and ( \2420_b0 , \2418_b0 , w_5205 );
and ( w_5204 ,  , w_5205 );
buf ( w_5203 , \2419_b1 );
not ( w_5203 , w_5206 );
not (  , w_5207 );
and ( w_5206 , w_5207 , \2419_b0 );
or ( \2421_b1 , \2420_b1 , w_5208 );
xor ( \2421_b0 , \2420_b0 , w_5210 );
not ( w_5210 , w_5211 );
and ( w_5211 , w_5208 , w_5209 );
buf ( w_5208 , \1404_b1 );
not ( w_5208 , w_5212 );
not ( w_5209 , w_5213 );
and ( w_5212 , w_5213 , \1404_b0 );
or ( \2422_b1 , \2416_b1 , \2421_b1 );
not ( \2421_b1 , w_5214 );
and ( \2422_b0 , \2416_b0 , w_5215 );
and ( w_5214 , w_5215 , \2421_b0 );
or ( \2423_b1 , \2412_b1 , \2421_b1 );
not ( \2421_b1 , w_5216 );
and ( \2423_b0 , \2412_b0 , w_5217 );
and ( w_5216 , w_5217 , \2421_b0 );
or ( \2425_b1 , \1384_b1 , \1431_b1 );
not ( \1431_b1 , w_5218 );
and ( \2425_b0 , \1384_b0 , w_5219 );
and ( w_5218 , w_5219 , \1431_b0 );
or ( \2426_b1 , \1342_b1 , \1429_b1 );
not ( \1429_b1 , w_5220 );
and ( \2426_b0 , \1342_b0 , w_5221 );
and ( w_5220 , w_5221 , \1429_b0 );
or ( \2427_b1 , \2425_b1 , w_5223 );
not ( w_5223 , w_5224 );
and ( \2427_b0 , \2425_b0 , w_5225 );
and ( w_5224 ,  , w_5225 );
buf ( w_5223 , \2426_b1 );
not ( w_5223 , w_5226 );
not (  , w_5227 );
and ( w_5226 , w_5227 , \2426_b0 );
or ( \2428_b1 , \2427_b1 , w_5228 );
xor ( \2428_b0 , \2427_b0 , w_5230 );
not ( w_5230 , w_5231 );
and ( w_5231 , w_5228 , w_5229 );
buf ( w_5228 , \1438_b1 );
not ( w_5228 , w_5232 );
not ( w_5229 , w_5233 );
and ( w_5232 , w_5233 , \1438_b0 );
or ( \2429_b1 , \1462_b1 , \1444_b1 );
not ( \1444_b1 , w_5234 );
and ( \2429_b0 , \1462_b0 , w_5235 );
and ( w_5234 , w_5235 , \1444_b0 );
or ( \2430_b1 , \1376_b1 , \1442_b1 );
not ( \1442_b1 , w_5236 );
and ( \2430_b0 , \1376_b0 , w_5237 );
and ( w_5236 , w_5237 , \1442_b0 );
or ( \2431_b1 , \2429_b1 , w_5239 );
not ( w_5239 , w_5240 );
and ( \2431_b0 , \2429_b0 , w_5241 );
and ( w_5240 ,  , w_5241 );
buf ( w_5239 , \2430_b1 );
not ( w_5239 , w_5242 );
not (  , w_5243 );
and ( w_5242 , w_5243 , \2430_b0 );
or ( \2432_b1 , \2431_b1 , w_5244 );
xor ( \2432_b0 , \2431_b0 , w_5246 );
not ( w_5246 , w_5247 );
and ( w_5247 , w_5244 , w_5245 );
buf ( w_5244 , \1451_b1 );
not ( w_5244 , w_5248 );
not ( w_5245 , w_5249 );
and ( w_5248 , w_5249 , \1451_b0 );
or ( \2433_b1 , \2428_b1 , \2432_b1 );
not ( \2432_b1 , w_5250 );
and ( \2433_b0 , \2428_b0 , w_5251 );
and ( w_5250 , w_5251 , \2432_b0 );
or ( \2434_b1 , \2424_b1 , \2433_b1 );
not ( \2433_b1 , w_5252 );
and ( \2434_b0 , \2424_b0 , w_5253 );
and ( w_5252 , w_5253 , \2433_b0 );
or ( \2435_b1 , \1553_b1 , \1643_b1 );
not ( \1643_b1 , w_5254 );
and ( \2435_b0 , \1553_b0 , w_5255 );
and ( w_5254 , w_5255 , \1643_b0 );
or ( \2436_b1 , \1533_b1 , \1641_b1 );
not ( \1641_b1 , w_5256 );
and ( \2436_b0 , \1533_b0 , w_5257 );
and ( w_5256 , w_5257 , \1641_b0 );
or ( \2437_b1 , \2435_b1 , w_5259 );
not ( w_5259 , w_5260 );
and ( \2437_b0 , \2435_b0 , w_5261 );
and ( w_5260 ,  , w_5261 );
buf ( w_5259 , \2436_b1 );
not ( w_5259 , w_5262 );
not (  , w_5263 );
and ( w_5262 , w_5263 , \2436_b0 );
or ( \2438_b1 , \2437_b1 , w_5264 );
xor ( \2438_b0 , \2437_b0 , w_5266 );
not ( w_5266 , w_5267 );
and ( w_5267 , w_5264 , w_5265 );
buf ( w_5264 , \1649_b1 );
not ( w_5264 , w_5268 );
not ( w_5265 , w_5269 );
and ( w_5268 , w_5269 , \1649_b0 );
or ( \2439_b1 , \2433_b1 , \2438_b1 );
not ( \2438_b1 , w_5270 );
and ( \2439_b0 , \2433_b0 , w_5271 );
and ( w_5270 , w_5271 , \2438_b0 );
or ( \2440_b1 , \2424_b1 , \2438_b1 );
not ( \2438_b1 , w_5272 );
and ( \2440_b0 , \2424_b0 , w_5273 );
and ( w_5272 , w_5273 , \2438_b0 );
or ( \2442_b1 , \1399_b1 , \1460_b1 );
not ( \1460_b1 , w_5274 );
and ( \2442_b0 , \1399_b0 , w_5275 );
and ( w_5274 , w_5275 , \1460_b0 );
or ( \2443_b1 , \1359_b1 , \1458_b1 );
not ( \1458_b1 , w_5276 );
and ( \2443_b0 , \1359_b0 , w_5277 );
and ( w_5276 , w_5277 , \1458_b0 );
or ( \2444_b1 , \2442_b1 , w_5279 );
not ( w_5279 , w_5280 );
and ( \2444_b0 , \2442_b0 , w_5281 );
and ( w_5280 ,  , w_5281 );
buf ( w_5279 , \2443_b1 );
not ( w_5279 , w_5282 );
not (  , w_5283 );
and ( w_5282 , w_5283 , \2443_b0 );
or ( \2445_b1 , \2444_b1 , w_5284 );
xor ( \2445_b0 , \2444_b0 , w_5286 );
not ( w_5286 , w_5287 );
and ( w_5287 , w_5284 , w_5285 );
buf ( w_5284 , \1467_b1 );
not ( w_5284 , w_5288 );
not ( w_5285 , w_5289 );
and ( w_5288 , w_5289 , \1467_b0 );
or ( \2446_b1 , \1616_b1 , \1475_b1 );
not ( \1475_b1 , w_5290 );
and ( \2446_b0 , \1616_b0 , w_5291 );
and ( w_5290 , w_5291 , \1475_b0 );
or ( \2447_b1 , \1391_b1 , \1473_b1 );
not ( \1473_b1 , w_5292 );
and ( \2447_b0 , \1391_b0 , w_5293 );
and ( w_5292 , w_5293 , \1473_b0 );
or ( \2448_b1 , \2446_b1 , w_5295 );
not ( w_5295 , w_5296 );
and ( \2448_b0 , \2446_b0 , w_5297 );
and ( w_5296 ,  , w_5297 );
buf ( w_5295 , \2447_b1 );
not ( w_5295 , w_5298 );
not (  , w_5299 );
and ( w_5298 , w_5299 , \2447_b0 );
or ( \2449_b1 , \2448_b1 , w_5300 );
xor ( \2449_b0 , \2448_b0 , w_5302 );
not ( w_5302 , w_5303 );
and ( w_5303 , w_5300 , w_5301 );
buf ( w_5300 , \1482_b1 );
not ( w_5300 , w_5304 );
not ( w_5301 , w_5305 );
and ( w_5304 , w_5305 , \1482_b0 );
or ( \2450_b1 , \2445_b1 , \2449_b1 );
not ( \2449_b1 , w_5306 );
and ( \2450_b0 , \2445_b0 , w_5307 );
and ( w_5306 , w_5307 , \2449_b0 );
or ( \2451_b1 , \1533_b1 , \1414_b1 );
not ( \1414_b1 , w_5308 );
and ( \2451_b0 , \1533_b0 , w_5309 );
and ( w_5308 , w_5309 , \1414_b0 );
or ( \2452_b1 , \1540_b1 , \1412_b1 );
not ( \1412_b1 , w_5310 );
and ( \2452_b0 , \1540_b0 , w_5311 );
and ( w_5310 , w_5311 , \1412_b0 );
or ( \2453_b1 , \2451_b1 , w_5313 );
not ( w_5313 , w_5314 );
and ( \2453_b0 , \2451_b0 , w_5315 );
and ( w_5314 ,  , w_5315 );
buf ( w_5313 , \2452_b1 );
not ( w_5313 , w_5316 );
not (  , w_5317 );
and ( w_5316 , w_5317 , \2452_b0 );
or ( \2454_b1 , \2453_b1 , w_5318 );
xor ( \2454_b0 , \2453_b0 , w_5320 );
not ( w_5320 , w_5321 );
and ( w_5321 , w_5318 , w_5319 );
buf ( w_5318 , \1421_b1 );
not ( w_5318 , w_5322 );
not ( w_5319 , w_5323 );
and ( w_5322 , w_5323 , \1421_b0 );
or ( \2455_b1 , \2449_b1 , \2454_b1 );
not ( \2454_b1 , w_5324 );
and ( \2455_b0 , \2449_b0 , w_5325 );
and ( w_5324 , w_5325 , \2454_b0 );
or ( \2456_b1 , \2445_b1 , \2454_b1 );
not ( \2454_b1 , w_5326 );
and ( \2456_b0 , \2445_b0 , w_5327 );
and ( w_5326 , w_5327 , \2454_b0 );
or ( \2458_b1 , \1351_b1 , \1336_b1 );
not ( \1336_b1 , w_5328 );
and ( \2458_b0 , \1351_b0 , w_5329 );
and ( w_5328 , w_5329 , \1336_b0 );
or ( \2459_b1 , \1446_b1 , \1333_b1 );
not ( \1333_b1 , w_5330 );
and ( \2459_b0 , \1446_b0 , w_5331 );
and ( w_5330 , w_5331 , \1333_b0 );
or ( \2460_b1 , \2458_b1 , w_5333 );
not ( w_5333 , w_5334 );
and ( \2460_b0 , \2458_b0 , w_5335 );
and ( w_5334 ,  , w_5335 );
buf ( w_5333 , \2459_b1 );
not ( w_5333 , w_5336 );
not (  , w_5337 );
and ( w_5336 , w_5337 , \2459_b0 );
or ( \2461_b1 , \2460_b1 , w_5338 );
xor ( \2461_b0 , \2460_b0 , w_5340 );
not ( w_5340 , w_5341 );
and ( w_5341 , w_5338 , w_5339 );
buf ( w_5338 , \1332_b1 );
not ( w_5338 , w_5342 );
not ( w_5339 , w_5343 );
and ( w_5342 , w_5343 , \1332_b0 );
or ( \2462_b1 , \1477_b1 , \1349_b1 );
not ( \1349_b1 , w_5344 );
and ( \2462_b0 , \1477_b0 , w_5345 );
and ( w_5344 , w_5345 , \1349_b0 );
or ( \2463_b1 , \1454_b1 , \1347_b1 );
not ( \1347_b1 , w_5346 );
and ( \2463_b0 , \1454_b0 , w_5347 );
and ( w_5346 , w_5347 , \1347_b0 );
or ( \2464_b1 , \2462_b1 , w_5349 );
not ( w_5349 , w_5350 );
and ( \2464_b0 , \2462_b0 , w_5351 );
and ( w_5350 ,  , w_5351 );
buf ( w_5349 , \2463_b1 );
not ( w_5349 , w_5352 );
not (  , w_5353 );
and ( w_5352 , w_5353 , \2463_b0 );
or ( \2465_b1 , \2464_b1 , w_5354 );
xor ( \2465_b0 , \2464_b0 , w_5356 );
not ( w_5356 , w_5357 );
and ( w_5357 , w_5354 , w_5355 );
buf ( w_5354 , \1356_b1 );
not ( w_5354 , w_5358 );
not ( w_5355 , w_5359 );
and ( w_5358 , w_5359 , \1356_b0 );
or ( \2466_b1 , \2461_b1 , \2465_b1 );
not ( \2465_b1 , w_5360 );
and ( \2466_b0 , \2461_b0 , w_5361 );
and ( w_5360 , w_5361 , \2465_b0 );
or ( \2467_b1 , \1498_b1 , \1641_b1 );
not ( \1641_b1 , w_5362 );
and ( \2467_b0 , \1498_b0 , w_5363 );
and ( w_5362 , w_5363 , \1641_b0 );
buf ( \2468_b1 , \2467_b1 );
not ( \2468_b1 , w_5364 );
not ( \2468_b0 , w_5365 );
and ( w_5364 , w_5365 , \2467_b0 );
or ( \2469_b1 , \2468_b1 , \1649_b1 );
not ( \1649_b1 , w_5366 );
and ( \2469_b0 , \2468_b0 , w_5367 );
and ( w_5366 , w_5367 , \1649_b0 );
or ( \2470_b1 , \2465_b1 , \2469_b1 );
not ( \2469_b1 , w_5368 );
and ( \2470_b0 , \2465_b0 , w_5369 );
and ( w_5368 , w_5369 , \2469_b0 );
or ( \2471_b1 , \2461_b1 , \2469_b1 );
not ( \2469_b1 , w_5370 );
and ( \2471_b0 , \2461_b0 , w_5371 );
and ( w_5370 , w_5371 , \2469_b0 );
or ( \2473_b1 , \2457_b1 , \2472_b1 );
not ( \2472_b1 , w_5372 );
and ( \2473_b0 , \2457_b0 , w_5373 );
and ( w_5372 , w_5373 , \2472_b0 );
or ( \2474_b1 , \2294_b1 , \2298_b1 );
xor ( \2474_b0 , \2294_b0 , w_5374 );
not ( w_5374 , w_5375 );
and ( w_5375 , \2298_b1 , \2298_b0 );
or ( \2475_b1 , \2474_b1 , \1921_b1 );
xor ( \2475_b0 , \2474_b0 , w_5376 );
not ( w_5376 , w_5377 );
and ( w_5377 , \1921_b1 , \1921_b0 );
or ( \2476_b1 , \2472_b1 , \2475_b1 );
not ( \2475_b1 , w_5378 );
and ( \2476_b0 , \2472_b0 , w_5379 );
and ( w_5378 , w_5379 , \2475_b0 );
or ( \2477_b1 , \2457_b1 , \2475_b1 );
not ( \2475_b1 , w_5380 );
and ( \2477_b0 , \2457_b0 , w_5381 );
and ( w_5380 , w_5381 , \2475_b0 );
or ( \2479_b1 , \2441_b1 , \2478_b1 );
not ( \2478_b1 , w_5382 );
and ( \2479_b0 , \2441_b0 , w_5383 );
and ( w_5382 , w_5383 , \2478_b0 );
or ( \2480_b1 , \2302_b1 , \2318_b1 );
xor ( \2480_b0 , \2302_b0 , w_5384 );
not ( w_5384 , w_5385 );
and ( w_5385 , \2318_b1 , \2318_b0 );
or ( \2481_b1 , \2480_b1 , \2323_b1 );
xor ( \2481_b0 , \2480_b0 , w_5386 );
not ( w_5386 , w_5387 );
and ( w_5387 , \2323_b1 , \2323_b0 );
or ( \2482_b1 , \2478_b1 , \2481_b1 );
not ( \2481_b1 , w_5388 );
and ( \2482_b0 , \2478_b0 , w_5389 );
and ( w_5388 , w_5389 , \2481_b0 );
or ( \2483_b1 , \2441_b1 , \2481_b1 );
not ( \2481_b1 , w_5390 );
and ( \2483_b0 , \2441_b0 , w_5391 );
and ( w_5390 , w_5391 , \2481_b0 );
or ( \2485_b1 , \2306_b1 , \2310_b1 );
xor ( \2485_b0 , \2306_b0 , w_5392 );
not ( w_5392 , w_5393 );
and ( w_5393 , \2310_b1 , \2310_b0 );
or ( \2486_b1 , \2485_b1 , \2315_b1 );
xor ( \2486_b0 , \2485_b0 , w_5394 );
not ( w_5394 , w_5395 );
and ( w_5395 , \2315_b1 , \2315_b0 );
or ( \2487_b1 , \2330_b1 , \2334_b1 );
xor ( \2487_b0 , \2330_b0 , w_5396 );
not ( w_5396 , w_5397 );
and ( w_5397 , \2334_b1 , \2334_b0 );
or ( \2488_b1 , \2487_b1 , \2339_b1 );
xor ( \2488_b0 , \2487_b0 , w_5398 );
not ( w_5398 , w_5399 );
and ( w_5399 , \2339_b1 , \2339_b0 );
or ( \2489_b1 , \2486_b1 , \2488_b1 );
not ( \2488_b1 , w_5400 );
and ( \2489_b0 , \2486_b0 , w_5401 );
and ( w_5400 , w_5401 , \2488_b0 );
or ( \2490_b1 , \2346_b1 , \2350_b1 );
xor ( \2490_b0 , \2346_b0 , w_5402 );
not ( w_5402 , w_5403 );
and ( w_5403 , \2350_b1 , \2350_b0 );
or ( \2491_b1 , \2490_b1 , \2355_b1 );
xor ( \2491_b0 , \2490_b0 , w_5404 );
not ( w_5404 , w_5405 );
and ( w_5405 , \2355_b1 , \2355_b0 );
or ( \2492_b1 , \2488_b1 , \2491_b1 );
not ( \2491_b1 , w_5406 );
and ( \2492_b0 , \2488_b0 , w_5407 );
and ( w_5406 , w_5407 , \2491_b0 );
or ( \2493_b1 , \2486_b1 , \2491_b1 );
not ( \2491_b1 , w_5408 );
and ( \2493_b0 , \2486_b0 , w_5409 );
and ( w_5408 , w_5409 , \2491_b0 );
or ( \2495_b1 , \2342_b1 , \2358_b1 );
xor ( \2495_b0 , \2342_b0 , w_5410 );
not ( w_5410 , w_5411 );
and ( w_5411 , \2358_b1 , \2358_b0 );
or ( \2496_b1 , \2495_b1 , \2361_b1 );
xor ( \2496_b0 , \2495_b0 , w_5412 );
not ( w_5412 , w_5413 );
and ( w_5413 , \2361_b1 , \2361_b0 );
or ( \2497_b1 , \2494_b1 , \2496_b1 );
not ( \2496_b1 , w_5414 );
and ( \2497_b0 , \2494_b0 , w_5415 );
and ( w_5414 , w_5415 , \2496_b0 );
or ( \2498_b1 , \2372_b1 , \2374_b1 );
xor ( \2498_b0 , \2372_b0 , w_5416 );
not ( w_5416 , w_5417 );
and ( w_5417 , \2374_b1 , \2374_b0 );
or ( \2499_b1 , \2498_b1 , \2377_b1 );
xor ( \2499_b0 , \2498_b0 , w_5418 );
not ( w_5418 , w_5419 );
and ( w_5419 , \2377_b1 , \2377_b0 );
or ( \2500_b1 , \2496_b1 , \2499_b1 );
not ( \2499_b1 , w_5420 );
and ( \2500_b0 , \2496_b0 , w_5421 );
and ( w_5420 , w_5421 , \2499_b0 );
or ( \2501_b1 , \2494_b1 , \2499_b1 );
not ( \2499_b1 , w_5422 );
and ( \2501_b0 , \2494_b0 , w_5423 );
and ( w_5422 , w_5423 , \2499_b0 );
or ( \2503_b1 , \2484_b1 , \2502_b1 );
not ( \2502_b1 , w_5424 );
and ( \2503_b0 , \2484_b0 , w_5425 );
and ( w_5424 , w_5425 , \2502_b0 );
or ( \2504_b1 , \2326_b1 , \2364_b1 );
xor ( \2504_b0 , \2326_b0 , w_5426 );
not ( w_5426 , w_5427 );
and ( w_5427 , \2364_b1 , \2364_b0 );
or ( \2505_b1 , \2504_b1 , \2367_b1 );
xor ( \2505_b0 , \2504_b0 , w_5428 );
not ( w_5428 , w_5429 );
and ( w_5429 , \2367_b1 , \2367_b0 );
or ( \2506_b1 , \2502_b1 , \2505_b1 );
not ( \2505_b1 , w_5430 );
and ( \2506_b0 , \2502_b0 , w_5431 );
and ( w_5430 , w_5431 , \2505_b0 );
or ( \2507_b1 , \2484_b1 , \2505_b1 );
not ( \2505_b1 , w_5432 );
and ( \2507_b0 , \2484_b0 , w_5433 );
and ( w_5432 , w_5433 , \2505_b0 );
or ( \2509_b1 , \2264_b1 , \2266_b1 );
xor ( \2509_b0 , \2264_b0 , w_5434 );
not ( w_5434 , w_5435 );
and ( w_5435 , \2266_b1 , \2266_b0 );
or ( \2510_b1 , \2509_b1 , \2269_b1 );
xor ( \2510_b0 , \2509_b0 , w_5436 );
not ( w_5436 , w_5437 );
and ( w_5437 , \2269_b1 , \2269_b0 );
or ( \2511_b1 , \2508_b1 , \2510_b1 );
not ( \2510_b1 , w_5438 );
and ( \2511_b0 , \2508_b0 , w_5439 );
and ( w_5438 , w_5439 , \2510_b0 );
or ( \2512_b1 , \2370_b1 , \2388_b1 );
xor ( \2512_b0 , \2370_b0 , w_5440 );
not ( w_5440 , w_5441 );
and ( w_5441 , \2388_b1 , \2388_b0 );
or ( \2513_b1 , \2512_b1 , \2391_b1 );
xor ( \2513_b0 , \2512_b0 , w_5442 );
not ( w_5442 , w_5443 );
and ( w_5443 , \2391_b1 , \2391_b0 );
or ( \2514_b1 , \2510_b1 , \2513_b1 );
not ( \2513_b1 , w_5444 );
and ( \2514_b0 , \2510_b0 , w_5445 );
and ( w_5444 , w_5445 , \2513_b0 );
or ( \2515_b1 , \2508_b1 , \2513_b1 );
not ( \2513_b1 , w_5446 );
and ( \2515_b0 , \2508_b0 , w_5447 );
and ( w_5446 , w_5447 , \2513_b0 );
or ( \2517_b1 , \2408_b1 , \2516_b1 );
not ( \2516_b1 , w_5448 );
and ( \2517_b0 , \2408_b0 , w_5449 );
and ( w_5448 , w_5449 , \2516_b0 );
or ( \2518_b1 , \2408_b1 , \2516_b1 );
xor ( \2518_b0 , \2408_b0 , w_5450 );
not ( w_5450 , w_5451 );
and ( w_5451 , \2516_b1 , \2516_b0 );
or ( \2519_b1 , \2508_b1 , \2510_b1 );
xor ( \2519_b0 , \2508_b0 , w_5452 );
not ( w_5452 , w_5453 );
and ( w_5453 , \2510_b1 , \2510_b0 );
or ( \2520_b1 , \2519_b1 , \2513_b1 );
xor ( \2520_b0 , \2519_b0 , w_5454 );
not ( w_5454 , w_5455 );
and ( w_5455 , \2513_b1 , \2513_b0 );
or ( \2521_b1 , \1376_b1 , \1431_b1 );
not ( \1431_b1 , w_5456 );
and ( \2521_b0 , \1376_b0 , w_5457 );
and ( w_5456 , w_5457 , \1431_b0 );
or ( \2522_b1 , \1384_b1 , \1429_b1 );
not ( \1429_b1 , w_5458 );
and ( \2522_b0 , \1384_b0 , w_5459 );
and ( w_5458 , w_5459 , \1429_b0 );
or ( \2523_b1 , \2521_b1 , w_5461 );
not ( w_5461 , w_5462 );
and ( \2523_b0 , \2521_b0 , w_5463 );
and ( w_5462 ,  , w_5463 );
buf ( w_5461 , \2522_b1 );
not ( w_5461 , w_5464 );
not (  , w_5465 );
and ( w_5464 , w_5465 , \2522_b0 );
or ( \2524_b1 , \2523_b1 , w_5466 );
xor ( \2524_b0 , \2523_b0 , w_5468 );
not ( w_5468 , w_5469 );
and ( w_5469 , w_5466 , w_5467 );
buf ( w_5466 , \1438_b1 );
not ( w_5466 , w_5470 );
not ( w_5467 , w_5471 );
and ( w_5470 , w_5471 , \1438_b0 );
or ( \2525_b1 , \1454_b1 , \1444_b1 );
not ( \1444_b1 , w_5472 );
and ( \2525_b0 , \1454_b0 , w_5473 );
and ( w_5472 , w_5473 , \1444_b0 );
or ( \2526_b1 , \1462_b1 , \1442_b1 );
not ( \1442_b1 , w_5474 );
and ( \2526_b0 , \1462_b0 , w_5475 );
and ( w_5474 , w_5475 , \1442_b0 );
or ( \2527_b1 , \2525_b1 , w_5477 );
not ( w_5477 , w_5478 );
and ( \2527_b0 , \2525_b0 , w_5479 );
and ( w_5478 ,  , w_5479 );
buf ( w_5477 , \2526_b1 );
not ( w_5477 , w_5480 );
not (  , w_5481 );
and ( w_5480 , w_5481 , \2526_b0 );
or ( \2528_b1 , \2527_b1 , w_5482 );
xor ( \2528_b0 , \2527_b0 , w_5484 );
not ( w_5484 , w_5485 );
and ( w_5485 , w_5482 , w_5483 );
buf ( w_5482 , \1451_b1 );
not ( w_5482 , w_5486 );
not ( w_5483 , w_5487 );
and ( w_5486 , w_5487 , \1451_b0 );
or ( \2529_b1 , \2524_b1 , \2528_b1 );
not ( \2528_b1 , w_5488 );
and ( \2529_b0 , \2524_b0 , w_5489 );
and ( w_5488 , w_5489 , \2528_b0 );
or ( \2530_b1 , \2528_b1 , \2467_b1 );
not ( \2467_b1 , w_5490 );
and ( \2530_b0 , \2528_b0 , w_5491 );
and ( w_5490 , w_5491 , \2467_b0 );
or ( \2531_b1 , \2524_b1 , \2467_b1 );
not ( \2467_b1 , w_5492 );
and ( \2531_b0 , \2524_b0 , w_5493 );
and ( w_5492 , w_5493 , \2467_b0 );
or ( \2533_b1 , \1359_b1 , \1382_b1 );
not ( \1382_b1 , w_5494 );
and ( \2533_b0 , \1359_b0 , w_5495 );
and ( w_5494 , w_5495 , \1382_b0 );
or ( \2534_b1 , \1368_b1 , \1380_b1 );
not ( \1380_b1 , w_5496 );
and ( \2534_b0 , \1368_b0 , w_5497 );
and ( w_5496 , w_5497 , \1380_b0 );
or ( \2535_b1 , \2533_b1 , w_5499 );
not ( w_5499 , w_5500 );
and ( \2535_b0 , \2533_b0 , w_5501 );
and ( w_5500 ,  , w_5501 );
buf ( w_5499 , \2534_b1 );
not ( w_5499 , w_5502 );
not (  , w_5503 );
and ( w_5502 , w_5503 , \2534_b0 );
or ( \2536_b1 , \2535_b1 , w_5504 );
xor ( \2536_b0 , \2535_b0 , w_5506 );
not ( w_5506 , w_5507 );
and ( w_5507 , w_5504 , w_5505 );
buf ( w_5504 , \1389_b1 );
not ( w_5504 , w_5508 );
not ( w_5505 , w_5509 );
and ( w_5508 , w_5509 , \1389_b0 );
or ( \2537_b1 , \1526_b1 , \1397_b1 );
not ( \1397_b1 , w_5510 );
and ( \2537_b0 , \1526_b0 , w_5511 );
and ( w_5510 , w_5511 , \1397_b0 );
or ( \2538_b1 , \1622_b1 , \1395_b1 );
not ( \1395_b1 , w_5512 );
and ( \2538_b0 , \1622_b0 , w_5513 );
and ( w_5512 , w_5513 , \1395_b0 );
or ( \2539_b1 , \2537_b1 , w_5515 );
not ( w_5515 , w_5516 );
and ( \2539_b0 , \2537_b0 , w_5517 );
and ( w_5516 ,  , w_5517 );
buf ( w_5515 , \2538_b1 );
not ( w_5515 , w_5518 );
not (  , w_5519 );
and ( w_5518 , w_5519 , \2538_b0 );
or ( \2540_b1 , \2539_b1 , w_5520 );
xor ( \2540_b0 , \2539_b0 , w_5522 );
not ( w_5522 , w_5523 );
and ( w_5523 , w_5520 , w_5521 );
buf ( w_5520 , \1404_b1 );
not ( w_5520 , w_5524 );
not ( w_5521 , w_5525 );
and ( w_5524 , w_5525 , \1404_b0 );
or ( \2541_b1 , \2536_b1 , \2540_b1 );
not ( \2540_b1 , w_5526 );
and ( \2541_b0 , \2536_b0 , w_5527 );
and ( w_5526 , w_5527 , \2540_b0 );
or ( \2542_b1 , \1553_b1 , \1414_b1 );
not ( \1414_b1 , w_5528 );
and ( \2542_b0 , \1553_b0 , w_5529 );
and ( w_5528 , w_5529 , \1414_b0 );
or ( \2543_b1 , \1533_b1 , \1412_b1 );
not ( \1412_b1 , w_5530 );
and ( \2543_b0 , \1533_b0 , w_5531 );
and ( w_5530 , w_5531 , \1412_b0 );
or ( \2544_b1 , \2542_b1 , w_5533 );
not ( w_5533 , w_5534 );
and ( \2544_b0 , \2542_b0 , w_5535 );
and ( w_5534 ,  , w_5535 );
buf ( w_5533 , \2543_b1 );
not ( w_5533 , w_5536 );
not (  , w_5537 );
and ( w_5536 , w_5537 , \2543_b0 );
or ( \2545_b1 , \2544_b1 , w_5538 );
xor ( \2545_b0 , \2544_b0 , w_5540 );
not ( w_5540 , w_5541 );
and ( w_5541 , w_5538 , w_5539 );
buf ( w_5538 , \1421_b1 );
not ( w_5538 , w_5542 );
not ( w_5539 , w_5543 );
and ( w_5542 , w_5543 , \1421_b0 );
or ( \2546_b1 , \2540_b1 , \2545_b1 );
not ( \2545_b1 , w_5544 );
and ( \2546_b0 , \2540_b0 , w_5545 );
and ( w_5544 , w_5545 , \2545_b0 );
or ( \2547_b1 , \2536_b1 , \2545_b1 );
not ( \2545_b1 , w_5546 );
and ( \2547_b0 , \2536_b0 , w_5547 );
and ( w_5546 , w_5547 , \2545_b0 );
or ( \2549_b1 , \2532_b1 , \2548_b1 );
not ( \2548_b1 , w_5548 );
and ( \2549_b0 , \2532_b0 , w_5549 );
and ( w_5548 , w_5549 , \2548_b0 );
or ( \2550_b1 , \1342_b1 , \1336_b1 );
not ( \1336_b1 , w_5550 );
and ( \2550_b0 , \1342_b0 , w_5551 );
and ( w_5550 , w_5551 , \1336_b0 );
or ( \2551_b1 , \1351_b1 , \1333_b1 );
not ( \1333_b1 , w_5552 );
and ( \2551_b0 , \1351_b0 , w_5553 );
and ( w_5552 , w_5553 , \1333_b0 );
or ( \2552_b1 , \2550_b1 , w_5555 );
not ( w_5555 , w_5556 );
and ( \2552_b0 , \2550_b0 , w_5557 );
and ( w_5556 ,  , w_5557 );
buf ( w_5555 , \2551_b1 );
not ( w_5555 , w_5558 );
not (  , w_5559 );
and ( w_5558 , w_5559 , \2551_b0 );
or ( \2553_b1 , \2552_b1 , w_5560 );
xor ( \2553_b0 , \2552_b0 , w_5562 );
not ( w_5562 , w_5563 );
and ( w_5563 , w_5560 , w_5561 );
buf ( w_5560 , \1332_b1 );
not ( w_5560 , w_5564 );
not ( w_5561 , w_5565 );
and ( w_5564 , w_5565 , \1332_b0 );
or ( \2554_b1 , \1470_b1 , \1349_b1 );
not ( \1349_b1 , w_5566 );
and ( \2554_b0 , \1470_b0 , w_5567 );
and ( w_5566 , w_5567 , \1349_b0 );
or ( \2555_b1 , \1477_b1 , \1347_b1 );
not ( \1347_b1 , w_5568 );
and ( \2555_b0 , \1477_b0 , w_5569 );
and ( w_5568 , w_5569 , \1347_b0 );
or ( \2556_b1 , \2554_b1 , w_5571 );
not ( w_5571 , w_5572 );
and ( \2556_b0 , \2554_b0 , w_5573 );
and ( w_5572 ,  , w_5573 );
buf ( w_5571 , \2555_b1 );
not ( w_5571 , w_5574 );
not (  , w_5575 );
and ( w_5574 , w_5575 , \2555_b0 );
or ( \2557_b1 , \2556_b1 , w_5576 );
xor ( \2557_b0 , \2556_b0 , w_5578 );
not ( w_5578 , w_5579 );
and ( w_5579 , w_5576 , w_5577 );
buf ( w_5576 , \1356_b1 );
not ( w_5576 , w_5580 );
not ( w_5577 , w_5581 );
and ( w_5580 , w_5581 , \1356_b0 );
or ( \2558_b1 , \2553_b1 , \2557_b1 );
not ( \2557_b1 , w_5582 );
and ( \2558_b0 , \2553_b0 , w_5583 );
and ( w_5582 , w_5583 , \2557_b0 );
or ( \2559_b1 , \1407_b1 , \1366_b1 );
not ( \1366_b1 , w_5584 );
and ( \2559_b0 , \1407_b0 , w_5585 );
and ( w_5584 , w_5585 , \1366_b0 );
or ( \2560_b1 , \1416_b1 , \1364_b1 );
not ( \1364_b1 , w_5586 );
and ( \2560_b0 , \1416_b0 , w_5587 );
and ( w_5586 , w_5587 , \1364_b0 );
or ( \2561_b1 , \2559_b1 , w_5589 );
not ( w_5589 , w_5590 );
and ( \2561_b0 , \2559_b0 , w_5591 );
and ( w_5590 ,  , w_5591 );
buf ( w_5589 , \2560_b1 );
not ( w_5589 , w_5592 );
not (  , w_5593 );
and ( w_5592 , w_5593 , \2560_b0 );
or ( \2562_b1 , \2561_b1 , w_5594 );
xor ( \2562_b0 , \2561_b0 , w_5596 );
not ( w_5596 , w_5597 );
and ( w_5597 , w_5594 , w_5595 );
buf ( w_5594 , \1373_b1 );
not ( w_5594 , w_5598 );
not ( w_5595 , w_5599 );
and ( w_5598 , w_5599 , \1373_b0 );
or ( \2563_b1 , \2557_b1 , \2562_b1 );
not ( \2562_b1 , w_5600 );
and ( \2563_b0 , \2557_b0 , w_5601 );
and ( w_5600 , w_5601 , \2562_b0 );
or ( \2564_b1 , \2553_b1 , \2562_b1 );
not ( \2562_b1 , w_5602 );
and ( \2564_b0 , \2553_b0 , w_5603 );
and ( w_5602 , w_5603 , \2562_b0 );
or ( \2566_b1 , \2548_b1 , \2565_b1 );
not ( \2565_b1 , w_5604 );
and ( \2566_b0 , \2548_b0 , w_5605 );
and ( w_5604 , w_5605 , \2565_b0 );
or ( \2567_b1 , \2532_b1 , \2565_b1 );
not ( \2565_b1 , w_5606 );
and ( \2567_b0 , \2532_b0 , w_5607 );
and ( w_5606 , w_5607 , \2565_b0 );
or ( \2569_b1 , \2428_b1 , \2432_b1 );
xor ( \2569_b0 , \2428_b0 , w_5608 );
not ( w_5608 , w_5609 );
and ( w_5609 , \2432_b1 , \2432_b0 );
or ( \2570_b1 , \1517_b1 , \1675_b1 );
not ( \1675_b1 , w_5610 );
and ( \2570_b0 , \1517_b0 , w_5611 );
and ( w_5610 , w_5611 , \1675_b0 );
or ( \2571_b1 , \1526_b1 , \1673_b1 );
not ( \1673_b1 , w_5612 );
and ( \2571_b0 , \1526_b0 , w_5613 );
and ( w_5612 , w_5613 , \1673_b0 );
or ( \2572_b1 , \2570_b1 , w_5615 );
not ( w_5615 , w_5616 );
and ( \2572_b0 , \2570_b0 , w_5617 );
and ( w_5616 ,  , w_5617 );
buf ( w_5615 , \2571_b1 );
not ( w_5615 , w_5618 );
not (  , w_5619 );
and ( w_5618 , w_5619 , \2571_b0 );
or ( \2573_b1 , \2572_b1 , w_5620 );
xor ( \2573_b0 , \2572_b0 , w_5622 );
not ( w_5622 , w_5623 );
and ( w_5623 , w_5620 , w_5621 );
buf ( w_5620 , \1681_b1 );
not ( w_5620 , w_5624 );
not ( w_5621 , w_5625 );
and ( w_5624 , w_5625 , \1681_b0 );
or ( \2574_b1 , \2569_b1 , \2573_b1 );
not ( \2573_b1 , w_5626 );
and ( \2574_b0 , \2569_b0 , w_5627 );
and ( w_5626 , w_5627 , \2573_b0 );
or ( \2575_b1 , \1498_b1 , \1643_b1 );
not ( \1643_b1 , w_5628 );
and ( \2575_b0 , \1498_b0 , w_5629 );
and ( w_5628 , w_5629 , \1643_b0 );
or ( \2576_b1 , \1553_b1 , \1641_b1 );
not ( \1641_b1 , w_5630 );
and ( \2576_b0 , \1553_b0 , w_5631 );
and ( w_5630 , w_5631 , \1641_b0 );
or ( \2577_b1 , \2575_b1 , w_5633 );
not ( w_5633 , w_5634 );
and ( \2577_b0 , \2575_b0 , w_5635 );
and ( w_5634 ,  , w_5635 );
buf ( w_5633 , \2576_b1 );
not ( w_5633 , w_5636 );
not (  , w_5637 );
and ( w_5636 , w_5637 , \2576_b0 );
or ( \2578_b1 , \2577_b1 , w_5638 );
xor ( \2578_b0 , \2577_b0 , w_5640 );
not ( w_5640 , w_5641 );
and ( w_5641 , w_5638 , w_5639 );
buf ( w_5638 , \1649_b1 );
not ( w_5638 , w_5642 );
not ( w_5639 , w_5643 );
and ( w_5642 , w_5643 , \1649_b0 );
or ( \2579_b1 , \2573_b1 , \2578_b1 );
not ( \2578_b1 , w_5644 );
and ( \2579_b0 , \2573_b0 , w_5645 );
and ( w_5644 , w_5645 , \2578_b0 );
or ( \2580_b1 , \2569_b1 , \2578_b1 );
not ( \2578_b1 , w_5646 );
and ( \2580_b0 , \2569_b0 , w_5647 );
and ( w_5646 , w_5647 , \2578_b0 );
or ( \2582_b1 , \2568_b1 , \2581_b1 );
not ( \2581_b1 , w_5648 );
and ( \2582_b0 , \2568_b0 , w_5649 );
and ( w_5648 , w_5649 , \2581_b0 );
or ( \2583_b1 , \2424_b1 , \2433_b1 );
xor ( \2583_b0 , \2424_b0 , w_5650 );
not ( w_5650 , w_5651 );
and ( w_5651 , \2433_b1 , \2433_b0 );
or ( \2584_b1 , \2583_b1 , \2438_b1 );
xor ( \2584_b0 , \2583_b0 , w_5652 );
not ( w_5652 , w_5653 );
and ( w_5653 , \2438_b1 , \2438_b0 );
or ( \2585_b1 , \2581_b1 , \2584_b1 );
not ( \2584_b1 , w_5654 );
and ( \2585_b0 , \2581_b0 , w_5655 );
and ( w_5654 , w_5655 , \2584_b0 );
or ( \2586_b1 , \2568_b1 , \2584_b1 );
not ( \2584_b1 , w_5656 );
and ( \2586_b0 , \2568_b0 , w_5657 );
and ( w_5656 , w_5657 , \2584_b0 );
or ( \2588_b1 , \1391_b1 , \1460_b1 );
not ( \1460_b1 , w_5658 );
and ( \2588_b0 , \1391_b0 , w_5659 );
and ( w_5658 , w_5659 , \1460_b0 );
or ( \2589_b1 , \1399_b1 , \1458_b1 );
not ( \1458_b1 , w_5660 );
and ( \2589_b0 , \1399_b0 , w_5661 );
and ( w_5660 , w_5661 , \1458_b0 );
or ( \2590_b1 , \2588_b1 , w_5663 );
not ( w_5663 , w_5664 );
and ( \2590_b0 , \2588_b0 , w_5665 );
and ( w_5664 ,  , w_5665 );
buf ( w_5663 , \2589_b1 );
not ( w_5663 , w_5666 );
not (  , w_5667 );
and ( w_5666 , w_5667 , \2589_b0 );
or ( \2591_b1 , \2590_b1 , w_5668 );
xor ( \2591_b0 , \2590_b0 , w_5670 );
not ( w_5670 , w_5671 );
and ( w_5671 , w_5668 , w_5669 );
buf ( w_5668 , \1467_b1 );
not ( w_5668 , w_5672 );
not ( w_5669 , w_5673 );
and ( w_5672 , w_5673 , \1467_b0 );
or ( \2592_b1 , \1586_b1 , \1475_b1 );
not ( \1475_b1 , w_5674 );
and ( \2592_b0 , \1586_b0 , w_5675 );
and ( w_5674 , w_5675 , \1475_b0 );
or ( \2593_b1 , \1616_b1 , \1473_b1 );
not ( \1473_b1 , w_5676 );
and ( \2593_b0 , \1616_b0 , w_5677 );
and ( w_5676 , w_5677 , \1473_b0 );
or ( \2594_b1 , \2592_b1 , w_5679 );
not ( w_5679 , w_5680 );
and ( \2594_b0 , \2592_b0 , w_5681 );
and ( w_5680 ,  , w_5681 );
buf ( w_5679 , \2593_b1 );
not ( w_5679 , w_5682 );
not (  , w_5683 );
and ( w_5682 , w_5683 , \2593_b0 );
or ( \2595_b1 , \2594_b1 , w_5684 );
xor ( \2595_b0 , \2594_b0 , w_5686 );
not ( w_5686 , w_5687 );
and ( w_5687 , w_5684 , w_5685 );
buf ( w_5684 , \1482_b1 );
not ( w_5684 , w_5688 );
not ( w_5685 , w_5689 );
and ( w_5688 , w_5689 , \1482_b0 );
or ( \2596_b1 , \2591_b1 , \2595_b1 );
not ( \2595_b1 , w_5690 );
and ( \2596_b0 , \2591_b0 , w_5691 );
and ( w_5690 , w_5691 , \2595_b0 );
or ( \2597_b1 , \1540_b1 , \1675_b1 );
not ( \1675_b1 , w_5692 );
and ( \2597_b0 , \1540_b0 , w_5693 );
and ( w_5692 , w_5693 , \1675_b0 );
or ( \2598_b1 , \1517_b1 , \1673_b1 );
not ( \1673_b1 , w_5694 );
and ( \2598_b0 , \1517_b0 , w_5695 );
and ( w_5694 , w_5695 , \1673_b0 );
or ( \2599_b1 , \2597_b1 , w_5697 );
not ( w_5697 , w_5698 );
and ( \2599_b0 , \2597_b0 , w_5699 );
and ( w_5698 ,  , w_5699 );
buf ( w_5697 , \2598_b1 );
not ( w_5697 , w_5700 );
not (  , w_5701 );
and ( w_5700 , w_5701 , \2598_b0 );
or ( \2600_b1 , \2599_b1 , w_5702 );
xor ( \2600_b0 , \2599_b0 , w_5704 );
not ( w_5704 , w_5705 );
and ( w_5705 , w_5702 , w_5703 );
buf ( w_5702 , \1681_b1 );
not ( w_5702 , w_5706 );
not ( w_5703 , w_5707 );
and ( w_5706 , w_5707 , \1681_b0 );
or ( \2601_b1 , \2595_b1 , \2600_b1 );
not ( \2600_b1 , w_5708 );
and ( \2601_b0 , \2595_b0 , w_5709 );
and ( w_5708 , w_5709 , \2600_b0 );
or ( \2602_b1 , \2591_b1 , \2600_b1 );
not ( \2600_b1 , w_5710 );
and ( \2602_b0 , \2591_b0 , w_5711 );
and ( w_5710 , w_5711 , \2600_b0 );
or ( \2604_b1 , \2412_b1 , \2416_b1 );
xor ( \2604_b0 , \2412_b0 , w_5712 );
not ( w_5712 , w_5713 );
and ( w_5713 , \2416_b1 , \2416_b0 );
or ( \2605_b1 , \2604_b1 , \2421_b1 );
xor ( \2605_b0 , \2604_b0 , w_5714 );
not ( w_5714 , w_5715 );
and ( w_5715 , \2421_b1 , \2421_b0 );
or ( \2606_b1 , \2603_b1 , \2605_b1 );
not ( \2605_b1 , w_5716 );
and ( \2606_b0 , \2603_b0 , w_5717 );
and ( w_5716 , w_5717 , \2605_b0 );
or ( \2607_b1 , \2445_b1 , \2449_b1 );
xor ( \2607_b0 , \2445_b0 , w_5718 );
not ( w_5718 , w_5719 );
and ( w_5719 , \2449_b1 , \2449_b0 );
or ( \2608_b1 , \2607_b1 , \2454_b1 );
xor ( \2608_b0 , \2607_b0 , w_5720 );
not ( w_5720 , w_5721 );
and ( w_5721 , \2454_b1 , \2454_b0 );
or ( \2609_b1 , \2605_b1 , \2608_b1 );
not ( \2608_b1 , w_5722 );
and ( \2609_b0 , \2605_b0 , w_5723 );
and ( w_5722 , w_5723 , \2608_b0 );
or ( \2610_b1 , \2603_b1 , \2608_b1 );
not ( \2608_b1 , w_5724 );
and ( \2610_b0 , \2603_b0 , w_5725 );
and ( w_5724 , w_5725 , \2608_b0 );
or ( \2612_b1 , \2457_b1 , \2472_b1 );
xor ( \2612_b0 , \2457_b0 , w_5726 );
not ( w_5726 , w_5727 );
and ( w_5727 , \2472_b1 , \2472_b0 );
or ( \2613_b1 , \2612_b1 , \2475_b1 );
xor ( \2613_b0 , \2612_b0 , w_5728 );
not ( w_5728 , w_5729 );
and ( w_5729 , \2475_b1 , \2475_b0 );
or ( \2614_b1 , \2611_b1 , \2613_b1 );
not ( \2613_b1 , w_5730 );
and ( \2614_b0 , \2611_b0 , w_5731 );
and ( w_5730 , w_5731 , \2613_b0 );
or ( \2615_b1 , \2486_b1 , \2488_b1 );
xor ( \2615_b0 , \2486_b0 , w_5732 );
not ( w_5732 , w_5733 );
and ( w_5733 , \2488_b1 , \2488_b0 );
or ( \2616_b1 , \2615_b1 , \2491_b1 );
xor ( \2616_b0 , \2615_b0 , w_5734 );
not ( w_5734 , w_5735 );
and ( w_5735 , \2491_b1 , \2491_b0 );
or ( \2617_b1 , \2613_b1 , \2616_b1 );
not ( \2616_b1 , w_5736 );
and ( \2617_b0 , \2613_b0 , w_5737 );
and ( w_5736 , w_5737 , \2616_b0 );
or ( \2618_b1 , \2611_b1 , \2616_b1 );
not ( \2616_b1 , w_5738 );
and ( \2618_b0 , \2611_b0 , w_5739 );
and ( w_5738 , w_5739 , \2616_b0 );
or ( \2620_b1 , \2587_b1 , \2619_b1 );
not ( \2619_b1 , w_5740 );
and ( \2620_b0 , \2587_b0 , w_5741 );
and ( w_5740 , w_5741 , \2619_b0 );
or ( \2621_b1 , \2441_b1 , \2478_b1 );
xor ( \2621_b0 , \2441_b0 , w_5742 );
not ( w_5742 , w_5743 );
and ( w_5743 , \2478_b1 , \2478_b0 );
or ( \2622_b1 , \2621_b1 , \2481_b1 );
xor ( \2622_b0 , \2621_b0 , w_5744 );
not ( w_5744 , w_5745 );
and ( w_5745 , \2481_b1 , \2481_b0 );
or ( \2623_b1 , \2619_b1 , \2622_b1 );
not ( \2622_b1 , w_5746 );
and ( \2623_b0 , \2619_b0 , w_5747 );
and ( w_5746 , w_5747 , \2622_b0 );
or ( \2624_b1 , \2587_b1 , \2622_b1 );
not ( \2622_b1 , w_5748 );
and ( \2624_b0 , \2587_b0 , w_5749 );
and ( w_5748 , w_5749 , \2622_b0 );
or ( \2626_b1 , \2380_b1 , \2382_b1 );
xor ( \2626_b0 , \2380_b0 , w_5750 );
not ( w_5750 , w_5751 );
and ( w_5751 , \2382_b1 , \2382_b0 );
or ( \2627_b1 , \2626_b1 , \2385_b1 );
xor ( \2627_b0 , \2626_b0 , w_5752 );
not ( w_5752 , w_5753 );
and ( w_5753 , \2385_b1 , \2385_b0 );
or ( \2628_b1 , \2625_b1 , \2627_b1 );
not ( \2627_b1 , w_5754 );
and ( \2628_b0 , \2625_b0 , w_5755 );
and ( w_5754 , w_5755 , \2627_b0 );
or ( \2629_b1 , \2484_b1 , \2502_b1 );
xor ( \2629_b0 , \2484_b0 , w_5756 );
not ( w_5756 , w_5757 );
and ( w_5757 , \2502_b1 , \2502_b0 );
or ( \2630_b1 , \2629_b1 , \2505_b1 );
xor ( \2630_b0 , \2629_b0 , w_5758 );
not ( w_5758 , w_5759 );
and ( w_5759 , \2505_b1 , \2505_b0 );
or ( \2631_b1 , \2627_b1 , \2630_b1 );
not ( \2630_b1 , w_5760 );
and ( \2631_b0 , \2627_b0 , w_5761 );
and ( w_5760 , w_5761 , \2630_b0 );
or ( \2632_b1 , \2625_b1 , \2630_b1 );
not ( \2630_b1 , w_5762 );
and ( \2632_b0 , \2625_b0 , w_5763 );
and ( w_5762 , w_5763 , \2630_b0 );
or ( \2634_b1 , \2520_b1 , \2633_b1 );
not ( \2633_b1 , w_5764 );
and ( \2634_b0 , \2520_b0 , w_5765 );
and ( w_5764 , w_5765 , \2633_b0 );
or ( \2635_b1 , \2520_b1 , \2633_b1 );
xor ( \2635_b0 , \2520_b0 , w_5766 );
not ( w_5766 , w_5767 );
and ( w_5767 , \2633_b1 , \2633_b0 );
or ( \2636_b1 , \2625_b1 , \2627_b1 );
xor ( \2636_b0 , \2625_b0 , w_5768 );
not ( w_5768 , w_5769 );
and ( w_5769 , \2627_b1 , \2627_b0 );
or ( \2637_b1 , \2636_b1 , \2630_b1 );
xor ( \2637_b0 , \2636_b0 , w_5770 );
not ( w_5770 , w_5771 );
and ( w_5771 , \2630_b1 , \2630_b0 );
or ( \2638_b1 , \1616_b1 , \1460_b1 );
not ( \1460_b1 , w_5772 );
and ( \2638_b0 , \1616_b0 , w_5773 );
and ( w_5772 , w_5773 , \1460_b0 );
or ( \2639_b1 , \1391_b1 , \1458_b1 );
not ( \1458_b1 , w_5774 );
and ( \2639_b0 , \1391_b0 , w_5775 );
and ( w_5774 , w_5775 , \1458_b0 );
or ( \2640_b1 , \2638_b1 , w_5777 );
not ( w_5777 , w_5778 );
and ( \2640_b0 , \2638_b0 , w_5779 );
and ( w_5778 ,  , w_5779 );
buf ( w_5777 , \2639_b1 );
not ( w_5777 , w_5780 );
not (  , w_5781 );
and ( w_5780 , w_5781 , \2639_b0 );
or ( \2641_b1 , \2640_b1 , w_5782 );
xor ( \2641_b0 , \2640_b0 , w_5784 );
not ( w_5784 , w_5785 );
and ( w_5785 , w_5782 , w_5783 );
buf ( w_5782 , \1467_b1 );
not ( w_5782 , w_5786 );
not ( w_5783 , w_5787 );
and ( w_5786 , w_5787 , \1467_b0 );
or ( \2642_b1 , \1416_b1 , \1475_b1 );
not ( \1475_b1 , w_5788 );
and ( \2642_b0 , \1416_b0 , w_5789 );
and ( w_5788 , w_5789 , \1475_b0 );
or ( \2643_b1 , \1586_b1 , \1473_b1 );
not ( \1473_b1 , w_5790 );
and ( \2643_b0 , \1586_b0 , w_5791 );
and ( w_5790 , w_5791 , \1473_b0 );
or ( \2644_b1 , \2642_b1 , w_5793 );
not ( w_5793 , w_5794 );
and ( \2644_b0 , \2642_b0 , w_5795 );
and ( w_5794 ,  , w_5795 );
buf ( w_5793 , \2643_b1 );
not ( w_5793 , w_5796 );
not (  , w_5797 );
and ( w_5796 , w_5797 , \2643_b0 );
or ( \2645_b1 , \2644_b1 , w_5798 );
xor ( \2645_b0 , \2644_b0 , w_5800 );
not ( w_5800 , w_5801 );
and ( w_5801 , w_5798 , w_5799 );
buf ( w_5798 , \1482_b1 );
not ( w_5798 , w_5802 );
not ( w_5799 , w_5803 );
and ( w_5802 , w_5803 , \1482_b0 );
or ( \2646_b1 , \2641_b1 , \2645_b1 );
not ( \2645_b1 , w_5804 );
and ( \2646_b0 , \2641_b0 , w_5805 );
and ( w_5804 , w_5805 , \2645_b0 );
or ( \2647_b1 , \1498_b1 , \1414_b1 );
not ( \1414_b1 , w_5806 );
and ( \2647_b0 , \1498_b0 , w_5807 );
and ( w_5806 , w_5807 , \1414_b0 );
or ( \2648_b1 , \1553_b1 , \1412_b1 );
not ( \1412_b1 , w_5808 );
and ( \2648_b0 , \1553_b0 , w_5809 );
and ( w_5808 , w_5809 , \1412_b0 );
or ( \2649_b1 , \2647_b1 , w_5811 );
not ( w_5811 , w_5812 );
and ( \2649_b0 , \2647_b0 , w_5813 );
and ( w_5812 ,  , w_5813 );
buf ( w_5811 , \2648_b1 );
not ( w_5811 , w_5814 );
not (  , w_5815 );
and ( w_5814 , w_5815 , \2648_b0 );
or ( \2650_b1 , \2649_b1 , w_5816 );
xor ( \2650_b0 , \2649_b0 , w_5818 );
not ( w_5818 , w_5819 );
and ( w_5819 , w_5816 , w_5817 );
buf ( w_5816 , \1421_b1 );
not ( w_5816 , w_5820 );
not ( w_5817 , w_5821 );
and ( w_5820 , w_5821 , \1421_b0 );
or ( \2651_b1 , \2645_b1 , \2650_b1 );
not ( \2650_b1 , w_5822 );
and ( \2651_b0 , \2645_b0 , w_5823 );
and ( w_5822 , w_5823 , \2650_b0 );
or ( \2652_b1 , \2641_b1 , \2650_b1 );
not ( \2650_b1 , w_5824 );
and ( \2652_b0 , \2641_b0 , w_5825 );
and ( w_5824 , w_5825 , \2650_b0 );
or ( \2654_b1 , \1399_b1 , \1382_b1 );
not ( \1382_b1 , w_5826 );
and ( \2654_b0 , \1399_b0 , w_5827 );
and ( w_5826 , w_5827 , \1382_b0 );
or ( \2655_b1 , \1359_b1 , \1380_b1 );
not ( \1380_b1 , w_5828 );
and ( \2655_b0 , \1359_b0 , w_5829 );
and ( w_5828 , w_5829 , \1380_b0 );
or ( \2656_b1 , \2654_b1 , w_5831 );
not ( w_5831 , w_5832 );
and ( \2656_b0 , \2654_b0 , w_5833 );
and ( w_5832 ,  , w_5833 );
buf ( w_5831 , \2655_b1 );
not ( w_5831 , w_5834 );
not (  , w_5835 );
and ( w_5834 , w_5835 , \2655_b0 );
or ( \2657_b1 , \2656_b1 , w_5836 );
xor ( \2657_b0 , \2656_b0 , w_5838 );
not ( w_5838 , w_5839 );
and ( w_5839 , w_5836 , w_5837 );
buf ( w_5836 , \1389_b1 );
not ( w_5836 , w_5840 );
not ( w_5837 , w_5841 );
and ( w_5840 , w_5841 , \1389_b0 );
or ( \2658_b1 , \1622_b1 , \1366_b1 );
not ( \1366_b1 , w_5842 );
and ( \2658_b0 , \1622_b0 , w_5843 );
and ( w_5842 , w_5843 , \1366_b0 );
or ( \2659_b1 , \1407_b1 , \1364_b1 );
not ( \1364_b1 , w_5844 );
and ( \2659_b0 , \1407_b0 , w_5845 );
and ( w_5844 , w_5845 , \1364_b0 );
or ( \2660_b1 , \2658_b1 , w_5847 );
not ( w_5847 , w_5848 );
and ( \2660_b0 , \2658_b0 , w_5849 );
and ( w_5848 ,  , w_5849 );
buf ( w_5847 , \2659_b1 );
not ( w_5847 , w_5850 );
not (  , w_5851 );
and ( w_5850 , w_5851 , \2659_b0 );
or ( \2661_b1 , \2660_b1 , w_5852 );
xor ( \2661_b0 , \2660_b0 , w_5854 );
not ( w_5854 , w_5855 );
and ( w_5855 , w_5852 , w_5853 );
buf ( w_5852 , \1373_b1 );
not ( w_5852 , w_5856 );
not ( w_5853 , w_5857 );
and ( w_5856 , w_5857 , \1373_b0 );
or ( \2662_b1 , \2657_b1 , \2661_b1 );
not ( \2661_b1 , w_5858 );
and ( \2662_b0 , \2657_b0 , w_5859 );
and ( w_5858 , w_5859 , \2661_b0 );
or ( \2663_b1 , \1517_b1 , \1397_b1 );
not ( \1397_b1 , w_5860 );
and ( \2663_b0 , \1517_b0 , w_5861 );
and ( w_5860 , w_5861 , \1397_b0 );
or ( \2664_b1 , \1526_b1 , \1395_b1 );
not ( \1395_b1 , w_5862 );
and ( \2664_b0 , \1526_b0 , w_5863 );
and ( w_5862 , w_5863 , \1395_b0 );
or ( \2665_b1 , \2663_b1 , w_5865 );
not ( w_5865 , w_5866 );
and ( \2665_b0 , \2663_b0 , w_5867 );
and ( w_5866 ,  , w_5867 );
buf ( w_5865 , \2664_b1 );
not ( w_5865 , w_5868 );
not (  , w_5869 );
and ( w_5868 , w_5869 , \2664_b0 );
or ( \2666_b1 , \2665_b1 , w_5870 );
xor ( \2666_b0 , \2665_b0 , w_5872 );
not ( w_5872 , w_5873 );
and ( w_5873 , w_5870 , w_5871 );
buf ( w_5870 , \1404_b1 );
not ( w_5870 , w_5874 );
not ( w_5871 , w_5875 );
and ( w_5874 , w_5875 , \1404_b0 );
or ( \2667_b1 , \2661_b1 , \2666_b1 );
not ( \2666_b1 , w_5876 );
and ( \2667_b0 , \2661_b0 , w_5877 );
and ( w_5876 , w_5877 , \2666_b0 );
or ( \2668_b1 , \2657_b1 , \2666_b1 );
not ( \2666_b1 , w_5878 );
and ( \2668_b0 , \2657_b0 , w_5879 );
and ( w_5878 , w_5879 , \2666_b0 );
or ( \2670_b1 , \2653_b1 , \2669_b1 );
not ( \2669_b1 , w_5880 );
and ( \2670_b0 , \2653_b0 , w_5881 );
and ( w_5880 , w_5881 , \2669_b0 );
or ( \2671_b1 , \1462_b1 , \1431_b1 );
not ( \1431_b1 , w_5882 );
and ( \2671_b0 , \1462_b0 , w_5883 );
and ( w_5882 , w_5883 , \1431_b0 );
or ( \2672_b1 , \1376_b1 , \1429_b1 );
not ( \1429_b1 , w_5884 );
and ( \2672_b0 , \1376_b0 , w_5885 );
and ( w_5884 , w_5885 , \1429_b0 );
or ( \2673_b1 , \2671_b1 , w_5887 );
not ( w_5887 , w_5888 );
and ( \2673_b0 , \2671_b0 , w_5889 );
and ( w_5888 ,  , w_5889 );
buf ( w_5887 , \2672_b1 );
not ( w_5887 , w_5890 );
not (  , w_5891 );
and ( w_5890 , w_5891 , \2672_b0 );
or ( \2674_b1 , \2673_b1 , w_5892 );
xor ( \2674_b0 , \2673_b0 , w_5894 );
not ( w_5894 , w_5895 );
and ( w_5895 , w_5892 , w_5893 );
buf ( w_5892 , \1438_b1 );
not ( w_5892 , w_5896 );
not ( w_5893 , w_5897 );
and ( w_5896 , w_5897 , \1438_b0 );
or ( \2675_b1 , \1498_b1 , \1412_b1 );
not ( \1412_b1 , w_5898 );
and ( \2675_b0 , \1498_b0 , w_5899 );
and ( w_5898 , w_5899 , \1412_b0 );
buf ( \2676_b1 , \2675_b1 );
not ( \2676_b1 , w_5900 );
not ( \2676_b0 , w_5901 );
and ( w_5900 , w_5901 , \2675_b0 );
or ( \2677_b1 , \2676_b1 , \1421_b1 );
not ( \1421_b1 , w_5902 );
and ( \2677_b0 , \2676_b0 , w_5903 );
and ( w_5902 , w_5903 , \1421_b0 );
or ( \2678_b1 , \2674_b1 , \2677_b1 );
not ( \2677_b1 , w_5904 );
and ( \2678_b0 , \2674_b0 , w_5905 );
and ( w_5904 , w_5905 , \2677_b0 );
or ( \2679_b1 , \2669_b1 , \2678_b1 );
not ( \2678_b1 , w_5906 );
and ( \2679_b0 , \2669_b0 , w_5907 );
and ( w_5906 , w_5907 , \2678_b0 );
or ( \2680_b1 , \2653_b1 , \2678_b1 );
not ( \2678_b1 , w_5908 );
and ( \2680_b0 , \2653_b0 , w_5909 );
and ( w_5908 , w_5909 , \2678_b0 );
or ( \2682_b1 , \2461_b1 , \2465_b1 );
xor ( \2682_b0 , \2461_b0 , w_5910 );
not ( w_5910 , w_5911 );
and ( w_5911 , \2465_b1 , \2465_b0 );
or ( \2683_b1 , \2682_b1 , \2469_b1 );
xor ( \2683_b0 , \2682_b0 , w_5912 );
not ( w_5912 , w_5913 );
and ( w_5913 , \2469_b1 , \2469_b0 );
or ( \2684_b1 , \2681_b1 , \2683_b1 );
not ( \2683_b1 , w_5914 );
and ( \2684_b0 , \2681_b0 , w_5915 );
and ( w_5914 , w_5915 , \2683_b0 );
or ( \2685_b1 , \2569_b1 , \2573_b1 );
xor ( \2685_b0 , \2569_b0 , w_5916 );
not ( w_5916 , w_5917 );
and ( w_5917 , \2573_b1 , \2573_b0 );
or ( \2686_b1 , \2685_b1 , \2578_b1 );
xor ( \2686_b0 , \2685_b0 , w_5918 );
not ( w_5918 , w_5919 );
and ( w_5919 , \2578_b1 , \2578_b0 );
or ( \2687_b1 , \2683_b1 , \2686_b1 );
not ( \2686_b1 , w_5920 );
and ( \2687_b0 , \2683_b0 , w_5921 );
and ( w_5920 , w_5921 , \2686_b0 );
or ( \2688_b1 , \2681_b1 , \2686_b1 );
not ( \2686_b1 , w_5922 );
and ( \2688_b0 , \2681_b0 , w_5923 );
and ( w_5922 , w_5923 , \2686_b0 );
or ( \2690_b1 , \1384_b1 , \1336_b1 );
not ( \1336_b1 , w_5924 );
and ( \2690_b0 , \1384_b0 , w_5925 );
and ( w_5924 , w_5925 , \1336_b0 );
or ( \2691_b1 , \1342_b1 , \1333_b1 );
not ( \1333_b1 , w_5926 );
and ( \2691_b0 , \1342_b0 , w_5927 );
and ( w_5926 , w_5927 , \1333_b0 );
or ( \2692_b1 , \2690_b1 , w_5929 );
not ( w_5929 , w_5930 );
and ( \2692_b0 , \2690_b0 , w_5931 );
and ( w_5930 ,  , w_5931 );
buf ( w_5929 , \2691_b1 );
not ( w_5929 , w_5932 );
not (  , w_5933 );
and ( w_5932 , w_5933 , \2691_b0 );
or ( \2693_b1 , \2692_b1 , w_5934 );
xor ( \2693_b0 , \2692_b0 , w_5936 );
not ( w_5936 , w_5937 );
and ( w_5937 , w_5934 , w_5935 );
buf ( w_5934 , \1332_b1 );
not ( w_5934 , w_5938 );
not ( w_5935 , w_5939 );
and ( w_5938 , w_5939 , \1332_b0 );
or ( \2694_b1 , \1477_b1 , \1444_b1 );
not ( \1444_b1 , w_5940 );
and ( \2694_b0 , \1477_b0 , w_5941 );
and ( w_5940 , w_5941 , \1444_b0 );
or ( \2695_b1 , \1454_b1 , \1442_b1 );
not ( \1442_b1 , w_5942 );
and ( \2695_b0 , \1454_b0 , w_5943 );
and ( w_5942 , w_5943 , \1442_b0 );
or ( \2696_b1 , \2694_b1 , w_5945 );
not ( w_5945 , w_5946 );
and ( \2696_b0 , \2694_b0 , w_5947 );
and ( w_5946 ,  , w_5947 );
buf ( w_5945 , \2695_b1 );
not ( w_5945 , w_5948 );
not (  , w_5949 );
and ( w_5948 , w_5949 , \2695_b0 );
or ( \2697_b1 , \2696_b1 , w_5950 );
xor ( \2697_b0 , \2696_b0 , w_5952 );
not ( w_5952 , w_5953 );
and ( w_5953 , w_5950 , w_5951 );
buf ( w_5950 , \1451_b1 );
not ( w_5950 , w_5954 );
not ( w_5951 , w_5955 );
and ( w_5954 , w_5955 , \1451_b0 );
or ( \2698_b1 , \2693_b1 , \2697_b1 );
not ( \2697_b1 , w_5956 );
and ( \2698_b0 , \2693_b0 , w_5957 );
and ( w_5956 , w_5957 , \2697_b0 );
or ( \2699_b1 , \1368_b1 , \1349_b1 );
not ( \1349_b1 , w_5958 );
and ( \2699_b0 , \1368_b0 , w_5959 );
and ( w_5958 , w_5959 , \1349_b0 );
or ( \2700_b1 , \1470_b1 , \1347_b1 );
not ( \1347_b1 , w_5960 );
and ( \2700_b0 , \1470_b0 , w_5961 );
and ( w_5960 , w_5961 , \1347_b0 );
or ( \2701_b1 , \2699_b1 , w_5963 );
not ( w_5963 , w_5964 );
and ( \2701_b0 , \2699_b0 , w_5965 );
and ( w_5964 ,  , w_5965 );
buf ( w_5963 , \2700_b1 );
not ( w_5963 , w_5966 );
not (  , w_5967 );
and ( w_5966 , w_5967 , \2700_b0 );
or ( \2702_b1 , \2701_b1 , w_5968 );
xor ( \2702_b0 , \2701_b0 , w_5970 );
not ( w_5970 , w_5971 );
and ( w_5971 , w_5968 , w_5969 );
buf ( w_5968 , \1356_b1 );
not ( w_5968 , w_5972 );
not ( w_5969 , w_5973 );
and ( w_5972 , w_5973 , \1356_b0 );
or ( \2703_b1 , \2697_b1 , \2702_b1 );
not ( \2702_b1 , w_5974 );
and ( \2703_b0 , \2697_b0 , w_5975 );
and ( w_5974 , w_5975 , \2702_b0 );
or ( \2704_b1 , \2693_b1 , \2702_b1 );
not ( \2702_b1 , w_5976 );
and ( \2704_b0 , \2693_b0 , w_5977 );
and ( w_5976 , w_5977 , \2702_b0 );
or ( \2706_b1 , \2524_b1 , \2528_b1 );
xor ( \2706_b0 , \2524_b0 , w_5978 );
not ( w_5978 , w_5979 );
and ( w_5979 , \2528_b1 , \2528_b0 );
or ( \2707_b1 , \2706_b1 , \2467_b1 );
xor ( \2707_b0 , \2706_b0 , w_5980 );
not ( w_5980 , w_5981 );
and ( w_5981 , \2467_b1 , \2467_b0 );
or ( \2708_b1 , \2705_b1 , \2707_b1 );
not ( \2707_b1 , w_5982 );
and ( \2708_b0 , \2705_b0 , w_5983 );
and ( w_5982 , w_5983 , \2707_b0 );
or ( \2709_b1 , \2536_b1 , \2540_b1 );
xor ( \2709_b0 , \2536_b0 , w_5984 );
not ( w_5984 , w_5985 );
and ( w_5985 , \2540_b1 , \2540_b0 );
or ( \2710_b1 , \2709_b1 , \2545_b1 );
xor ( \2710_b0 , \2709_b0 , w_5986 );
not ( w_5986 , w_5987 );
and ( w_5987 , \2545_b1 , \2545_b0 );
or ( \2711_b1 , \2707_b1 , \2710_b1 );
not ( \2710_b1 , w_5988 );
and ( \2711_b0 , \2707_b0 , w_5989 );
and ( w_5988 , w_5989 , \2710_b0 );
or ( \2712_b1 , \2705_b1 , \2710_b1 );
not ( \2710_b1 , w_5990 );
and ( \2712_b0 , \2705_b0 , w_5991 );
and ( w_5990 , w_5991 , \2710_b0 );
or ( \2714_b1 , \2674_b1 , \2677_b1 );
xor ( \2714_b0 , \2674_b0 , w_5992 );
not ( w_5992 , w_5993 );
and ( w_5993 , \2677_b1 , \2677_b0 );
or ( \2715_b1 , \1454_b1 , \1431_b1 );
not ( \1431_b1 , w_5994 );
and ( \2715_b0 , \1454_b0 , w_5995 );
and ( w_5994 , w_5995 , \1431_b0 );
or ( \2716_b1 , \1462_b1 , \1429_b1 );
not ( \1429_b1 , w_5996 );
and ( \2716_b0 , \1462_b0 , w_5997 );
and ( w_5996 , w_5997 , \1429_b0 );
or ( \2717_b1 , \2715_b1 , w_5999 );
not ( w_5999 , w_6000 );
and ( \2717_b0 , \2715_b0 , w_6001 );
and ( w_6000 ,  , w_6001 );
buf ( w_5999 , \2716_b1 );
not ( w_5999 , w_6002 );
not (  , w_6003 );
and ( w_6002 , w_6003 , \2716_b0 );
or ( \2718_b1 , \2717_b1 , w_6004 );
xor ( \2718_b0 , \2717_b0 , w_6006 );
not ( w_6006 , w_6007 );
and ( w_6007 , w_6004 , w_6005 );
buf ( w_6004 , \1438_b1 );
not ( w_6004 , w_6008 );
not ( w_6005 , w_6009 );
and ( w_6008 , w_6009 , \1438_b0 );
or ( \2719_b1 , \1470_b1 , \1444_b1 );
not ( \1444_b1 , w_6010 );
and ( \2719_b0 , \1470_b0 , w_6011 );
and ( w_6010 , w_6011 , \1444_b0 );
or ( \2720_b1 , \1477_b1 , \1442_b1 );
not ( \1442_b1 , w_6012 );
and ( \2720_b0 , \1477_b0 , w_6013 );
and ( w_6012 , w_6013 , \1442_b0 );
or ( \2721_b1 , \2719_b1 , w_6015 );
not ( w_6015 , w_6016 );
and ( \2721_b0 , \2719_b0 , w_6017 );
and ( w_6016 ,  , w_6017 );
buf ( w_6015 , \2720_b1 );
not ( w_6015 , w_6018 );
not (  , w_6019 );
and ( w_6018 , w_6019 , \2720_b0 );
or ( \2722_b1 , \2721_b1 , w_6020 );
xor ( \2722_b0 , \2721_b0 , w_6022 );
not ( w_6022 , w_6023 );
and ( w_6023 , w_6020 , w_6021 );
buf ( w_6020 , \1451_b1 );
not ( w_6020 , w_6024 );
not ( w_6021 , w_6025 );
and ( w_6024 , w_6025 , \1451_b0 );
or ( \2723_b1 , \2718_b1 , \2722_b1 );
not ( \2722_b1 , w_6026 );
and ( \2723_b0 , \2718_b0 , w_6027 );
and ( w_6026 , w_6027 , \2722_b0 );
or ( \2724_b1 , \2722_b1 , \2675_b1 );
not ( \2675_b1 , w_6028 );
and ( \2724_b0 , \2722_b0 , w_6029 );
and ( w_6028 , w_6029 , \2675_b0 );
or ( \2725_b1 , \2718_b1 , \2675_b1 );
not ( \2675_b1 , w_6030 );
and ( \2725_b0 , \2718_b0 , w_6031 );
and ( w_6030 , w_6031 , \2675_b0 );
or ( \2727_b1 , \2714_b1 , \2726_b1 );
not ( \2726_b1 , w_6032 );
and ( \2727_b0 , \2714_b0 , w_6033 );
and ( w_6032 , w_6033 , \2726_b0 );
or ( \2728_b1 , \1533_b1 , \1675_b1 );
not ( \1675_b1 , w_6034 );
and ( \2728_b0 , \1533_b0 , w_6035 );
and ( w_6034 , w_6035 , \1675_b0 );
or ( \2729_b1 , \1540_b1 , \1673_b1 );
not ( \1673_b1 , w_6036 );
and ( \2729_b0 , \1540_b0 , w_6037 );
and ( w_6036 , w_6037 , \1673_b0 );
or ( \2730_b1 , \2728_b1 , w_6039 );
not ( w_6039 , w_6040 );
and ( \2730_b0 , \2728_b0 , w_6041 );
and ( w_6040 ,  , w_6041 );
buf ( w_6039 , \2729_b1 );
not ( w_6039 , w_6042 );
not (  , w_6043 );
and ( w_6042 , w_6043 , \2729_b0 );
or ( \2731_b1 , \2730_b1 , w_6044 );
xor ( \2731_b0 , \2730_b0 , w_6046 );
not ( w_6046 , w_6047 );
and ( w_6047 , w_6044 , w_6045 );
buf ( w_6044 , \1681_b1 );
not ( w_6044 , w_6048 );
not ( w_6045 , w_6049 );
and ( w_6048 , w_6049 , \1681_b0 );
or ( \2732_b1 , \2726_b1 , \2731_b1 );
not ( \2731_b1 , w_6050 );
and ( \2732_b0 , \2726_b0 , w_6051 );
and ( w_6050 , w_6051 , \2731_b0 );
or ( \2733_b1 , \2714_b1 , \2731_b1 );
not ( \2731_b1 , w_6052 );
and ( \2733_b0 , \2714_b0 , w_6053 );
and ( w_6052 , w_6053 , \2731_b0 );
or ( \2735_b1 , \2591_b1 , \2595_b1 );
xor ( \2735_b0 , \2591_b0 , w_6054 );
not ( w_6054 , w_6055 );
and ( w_6055 , \2595_b1 , \2595_b0 );
or ( \2736_b1 , \2735_b1 , \2600_b1 );
xor ( \2736_b0 , \2735_b0 , w_6056 );
not ( w_6056 , w_6057 );
and ( w_6057 , \2600_b1 , \2600_b0 );
or ( \2737_b1 , \2734_b1 , \2736_b1 );
not ( \2736_b1 , w_6058 );
and ( \2737_b0 , \2734_b0 , w_6059 );
and ( w_6058 , w_6059 , \2736_b0 );
or ( \2738_b1 , \2553_b1 , \2557_b1 );
xor ( \2738_b0 , \2553_b0 , w_6060 );
not ( w_6060 , w_6061 );
and ( w_6061 , \2557_b1 , \2557_b0 );
or ( \2739_b1 , \2738_b1 , \2562_b1 );
xor ( \2739_b0 , \2738_b0 , w_6062 );
not ( w_6062 , w_6063 );
and ( w_6063 , \2562_b1 , \2562_b0 );
or ( \2740_b1 , \2736_b1 , \2739_b1 );
not ( \2739_b1 , w_6064 );
and ( \2740_b0 , \2736_b0 , w_6065 );
and ( w_6064 , w_6065 , \2739_b0 );
or ( \2741_b1 , \2734_b1 , \2739_b1 );
not ( \2739_b1 , w_6066 );
and ( \2741_b0 , \2734_b0 , w_6067 );
and ( w_6066 , w_6067 , \2739_b0 );
or ( \2743_b1 , \2713_b1 , \2742_b1 );
not ( \2742_b1 , w_6068 );
and ( \2743_b0 , \2713_b0 , w_6069 );
and ( w_6068 , w_6069 , \2742_b0 );
or ( \2744_b1 , \2532_b1 , \2548_b1 );
xor ( \2744_b0 , \2532_b0 , w_6070 );
not ( w_6070 , w_6071 );
and ( w_6071 , \2548_b1 , \2548_b0 );
or ( \2745_b1 , \2744_b1 , \2565_b1 );
xor ( \2745_b0 , \2744_b0 , w_6072 );
not ( w_6072 , w_6073 );
and ( w_6073 , \2565_b1 , \2565_b0 );
or ( \2746_b1 , \2742_b1 , \2745_b1 );
not ( \2745_b1 , w_6074 );
and ( \2746_b0 , \2742_b0 , w_6075 );
and ( w_6074 , w_6075 , \2745_b0 );
or ( \2747_b1 , \2713_b1 , \2745_b1 );
not ( \2745_b1 , w_6076 );
and ( \2747_b0 , \2713_b0 , w_6077 );
and ( w_6076 , w_6077 , \2745_b0 );
or ( \2749_b1 , \2689_b1 , \2748_b1 );
not ( \2748_b1 , w_6078 );
and ( \2749_b0 , \2689_b0 , w_6079 );
and ( w_6078 , w_6079 , \2748_b0 );
or ( \2750_b1 , \2568_b1 , \2581_b1 );
xor ( \2750_b0 , \2568_b0 , w_6080 );
not ( w_6080 , w_6081 );
and ( w_6081 , \2581_b1 , \2581_b0 );
or ( \2751_b1 , \2750_b1 , \2584_b1 );
xor ( \2751_b0 , \2750_b0 , w_6082 );
not ( w_6082 , w_6083 );
and ( w_6083 , \2584_b1 , \2584_b0 );
or ( \2752_b1 , \2748_b1 , \2751_b1 );
not ( \2751_b1 , w_6084 );
and ( \2752_b0 , \2748_b0 , w_6085 );
and ( w_6084 , w_6085 , \2751_b0 );
or ( \2753_b1 , \2689_b1 , \2751_b1 );
not ( \2751_b1 , w_6086 );
and ( \2753_b0 , \2689_b0 , w_6087 );
and ( w_6086 , w_6087 , \2751_b0 );
or ( \2755_b1 , \2494_b1 , \2496_b1 );
xor ( \2755_b0 , \2494_b0 , w_6088 );
not ( w_6088 , w_6089 );
and ( w_6089 , \2496_b1 , \2496_b0 );
or ( \2756_b1 , \2755_b1 , \2499_b1 );
xor ( \2756_b0 , \2755_b0 , w_6090 );
not ( w_6090 , w_6091 );
and ( w_6091 , \2499_b1 , \2499_b0 );
or ( \2757_b1 , \2754_b1 , \2756_b1 );
not ( \2756_b1 , w_6092 );
and ( \2757_b0 , \2754_b0 , w_6093 );
and ( w_6092 , w_6093 , \2756_b0 );
or ( \2758_b1 , \2587_b1 , \2619_b1 );
xor ( \2758_b0 , \2587_b0 , w_6094 );
not ( w_6094 , w_6095 );
and ( w_6095 , \2619_b1 , \2619_b0 );
or ( \2759_b1 , \2758_b1 , \2622_b1 );
xor ( \2759_b0 , \2758_b0 , w_6096 );
not ( w_6096 , w_6097 );
and ( w_6097 , \2622_b1 , \2622_b0 );
or ( \2760_b1 , \2756_b1 , \2759_b1 );
not ( \2759_b1 , w_6098 );
and ( \2760_b0 , \2756_b0 , w_6099 );
and ( w_6098 , w_6099 , \2759_b0 );
or ( \2761_b1 , \2754_b1 , \2759_b1 );
not ( \2759_b1 , w_6100 );
and ( \2761_b0 , \2754_b0 , w_6101 );
and ( w_6100 , w_6101 , \2759_b0 );
or ( \2763_b1 , \2637_b1 , \2762_b1 );
not ( \2762_b1 , w_6102 );
and ( \2763_b0 , \2637_b0 , w_6103 );
and ( w_6102 , w_6103 , \2762_b0 );
or ( \2764_b1 , \2637_b1 , \2762_b1 );
xor ( \2764_b0 , \2637_b0 , w_6104 );
not ( w_6104 , w_6105 );
and ( w_6105 , \2762_b1 , \2762_b0 );
or ( \2765_b1 , \2754_b1 , \2756_b1 );
xor ( \2765_b0 , \2754_b0 , w_6106 );
not ( w_6106 , w_6107 );
and ( w_6107 , \2756_b1 , \2756_b0 );
or ( \2766_b1 , \2765_b1 , \2759_b1 );
xor ( \2766_b0 , \2765_b0 , w_6108 );
not ( w_6108 , w_6109 );
and ( w_6109 , \2759_b1 , \2759_b0 );
or ( \2767_b1 , \1376_b1 , \1336_b1 );
not ( \1336_b1 , w_6110 );
and ( \2767_b0 , \1376_b0 , w_6111 );
and ( w_6110 , w_6111 , \1336_b0 );
or ( \2768_b1 , \1384_b1 , \1333_b1 );
not ( \1333_b1 , w_6112 );
and ( \2768_b0 , \1384_b0 , w_6113 );
and ( w_6112 , w_6113 , \1333_b0 );
or ( \2769_b1 , \2767_b1 , w_6115 );
not ( w_6115 , w_6116 );
and ( \2769_b0 , \2767_b0 , w_6117 );
and ( w_6116 ,  , w_6117 );
buf ( w_6115 , \2768_b1 );
not ( w_6115 , w_6118 );
not (  , w_6119 );
and ( w_6118 , w_6119 , \2768_b0 );
or ( \2770_b1 , \2769_b1 , w_6120 );
xor ( \2770_b0 , \2769_b0 , w_6122 );
not ( w_6122 , w_6123 );
and ( w_6123 , w_6120 , w_6121 );
buf ( w_6120 , \1332_b1 );
not ( w_6120 , w_6124 );
not ( w_6121 , w_6125 );
and ( w_6124 , w_6125 , \1332_b0 );
or ( \2771_b1 , \1391_b1 , \1382_b1 );
not ( \1382_b1 , w_6126 );
and ( \2771_b0 , \1391_b0 , w_6127 );
and ( w_6126 , w_6127 , \1382_b0 );
or ( \2772_b1 , \1399_b1 , \1380_b1 );
not ( \1380_b1 , w_6128 );
and ( \2772_b0 , \1399_b0 , w_6129 );
and ( w_6128 , w_6129 , \1380_b0 );
or ( \2773_b1 , \2771_b1 , w_6131 );
not ( w_6131 , w_6132 );
and ( \2773_b0 , \2771_b0 , w_6133 );
and ( w_6132 ,  , w_6133 );
buf ( w_6131 , \2772_b1 );
not ( w_6131 , w_6134 );
not (  , w_6135 );
and ( w_6134 , w_6135 , \2772_b0 );
or ( \2774_b1 , \2773_b1 , w_6136 );
xor ( \2774_b0 , \2773_b0 , w_6138 );
not ( w_6138 , w_6139 );
and ( w_6139 , w_6136 , w_6137 );
buf ( w_6136 , \1389_b1 );
not ( w_6136 , w_6140 );
not ( w_6137 , w_6141 );
and ( w_6140 , w_6141 , \1389_b0 );
or ( \2775_b1 , \2770_b1 , \2774_b1 );
not ( \2774_b1 , w_6142 );
and ( \2775_b0 , \2770_b0 , w_6143 );
and ( w_6142 , w_6143 , \2774_b0 );
or ( \2776_b1 , \1586_b1 , \1460_b1 );
not ( \1460_b1 , w_6144 );
and ( \2776_b0 , \1586_b0 , w_6145 );
and ( w_6144 , w_6145 , \1460_b0 );
or ( \2777_b1 , \1616_b1 , \1458_b1 );
not ( \1458_b1 , w_6146 );
and ( \2777_b0 , \1616_b0 , w_6147 );
and ( w_6146 , w_6147 , \1458_b0 );
or ( \2778_b1 , \2776_b1 , w_6149 );
not ( w_6149 , w_6150 );
and ( \2778_b0 , \2776_b0 , w_6151 );
and ( w_6150 ,  , w_6151 );
buf ( w_6149 , \2777_b1 );
not ( w_6149 , w_6152 );
not (  , w_6153 );
and ( w_6152 , w_6153 , \2777_b0 );
or ( \2779_b1 , \2778_b1 , w_6154 );
xor ( \2779_b0 , \2778_b0 , w_6156 );
not ( w_6156 , w_6157 );
and ( w_6157 , w_6154 , w_6155 );
buf ( w_6154 , \1467_b1 );
not ( w_6154 , w_6158 );
not ( w_6155 , w_6159 );
and ( w_6158 , w_6159 , \1467_b0 );
or ( \2780_b1 , \2774_b1 , \2779_b1 );
not ( \2779_b1 , w_6160 );
and ( \2780_b0 , \2774_b0 , w_6161 );
and ( w_6160 , w_6161 , \2779_b0 );
or ( \2781_b1 , \2770_b1 , \2779_b1 );
not ( \2779_b1 , w_6162 );
and ( \2781_b0 , \2770_b0 , w_6163 );
and ( w_6162 , w_6163 , \2779_b0 );
or ( \2783_b1 , \1359_b1 , \1349_b1 );
not ( \1349_b1 , w_6164 );
and ( \2783_b0 , \1359_b0 , w_6165 );
and ( w_6164 , w_6165 , \1349_b0 );
or ( \2784_b1 , \1368_b1 , \1347_b1 );
not ( \1347_b1 , w_6166 );
and ( \2784_b0 , \1368_b0 , w_6167 );
and ( w_6166 , w_6167 , \1347_b0 );
or ( \2785_b1 , \2783_b1 , w_6169 );
not ( w_6169 , w_6170 );
and ( \2785_b0 , \2783_b0 , w_6171 );
and ( w_6170 ,  , w_6171 );
buf ( w_6169 , \2784_b1 );
not ( w_6169 , w_6172 );
not (  , w_6173 );
and ( w_6172 , w_6173 , \2784_b0 );
or ( \2786_b1 , \2785_b1 , w_6174 );
xor ( \2786_b0 , \2785_b0 , w_6176 );
not ( w_6176 , w_6177 );
and ( w_6177 , w_6174 , w_6175 );
buf ( w_6174 , \1356_b1 );
not ( w_6174 , w_6178 );
not ( w_6175 , w_6179 );
and ( w_6178 , w_6179 , \1356_b0 );
or ( \2787_b1 , \1526_b1 , \1366_b1 );
not ( \1366_b1 , w_6180 );
and ( \2787_b0 , \1526_b0 , w_6181 );
and ( w_6180 , w_6181 , \1366_b0 );
or ( \2788_b1 , \1622_b1 , \1364_b1 );
not ( \1364_b1 , w_6182 );
and ( \2788_b0 , \1622_b0 , w_6183 );
and ( w_6182 , w_6183 , \1364_b0 );
or ( \2789_b1 , \2787_b1 , w_6185 );
not ( w_6185 , w_6186 );
and ( \2789_b0 , \2787_b0 , w_6187 );
and ( w_6186 ,  , w_6187 );
buf ( w_6185 , \2788_b1 );
not ( w_6185 , w_6188 );
not (  , w_6189 );
and ( w_6188 , w_6189 , \2788_b0 );
or ( \2790_b1 , \2789_b1 , w_6190 );
xor ( \2790_b0 , \2789_b0 , w_6192 );
not ( w_6192 , w_6193 );
and ( w_6193 , w_6190 , w_6191 );
buf ( w_6190 , \1373_b1 );
not ( w_6190 , w_6194 );
not ( w_6191 , w_6195 );
and ( w_6194 , w_6195 , \1373_b0 );
or ( \2791_b1 , \2786_b1 , \2790_b1 );
not ( \2790_b1 , w_6196 );
and ( \2791_b0 , \2786_b0 , w_6197 );
and ( w_6196 , w_6197 , \2790_b0 );
or ( \2792_b1 , \1540_b1 , \1397_b1 );
not ( \1397_b1 , w_6198 );
and ( \2792_b0 , \1540_b0 , w_6199 );
and ( w_6198 , w_6199 , \1397_b0 );
or ( \2793_b1 , \1517_b1 , \1395_b1 );
not ( \1395_b1 , w_6200 );
and ( \2793_b0 , \1517_b0 , w_6201 );
and ( w_6200 , w_6201 , \1395_b0 );
or ( \2794_b1 , \2792_b1 , w_6203 );
not ( w_6203 , w_6204 );
and ( \2794_b0 , \2792_b0 , w_6205 );
and ( w_6204 ,  , w_6205 );
buf ( w_6203 , \2793_b1 );
not ( w_6203 , w_6206 );
not (  , w_6207 );
and ( w_6206 , w_6207 , \2793_b0 );
or ( \2795_b1 , \2794_b1 , w_6208 );
xor ( \2795_b0 , \2794_b0 , w_6210 );
not ( w_6210 , w_6211 );
and ( w_6211 , w_6208 , w_6209 );
buf ( w_6208 , \1404_b1 );
not ( w_6208 , w_6212 );
not ( w_6209 , w_6213 );
and ( w_6212 , w_6213 , \1404_b0 );
or ( \2796_b1 , \2790_b1 , \2795_b1 );
not ( \2795_b1 , w_6214 );
and ( \2796_b0 , \2790_b0 , w_6215 );
and ( w_6214 , w_6215 , \2795_b0 );
or ( \2797_b1 , \2786_b1 , \2795_b1 );
not ( \2795_b1 , w_6216 );
and ( \2797_b0 , \2786_b0 , w_6217 );
and ( w_6216 , w_6217 , \2795_b0 );
or ( \2799_b1 , \2782_b1 , \2798_b1 );
not ( \2798_b1 , w_6218 );
and ( \2799_b0 , \2782_b0 , w_6219 );
and ( w_6218 , w_6219 , \2798_b0 );
or ( \2800_b1 , \2641_b1 , \2645_b1 );
xor ( \2800_b0 , \2641_b0 , w_6220 );
not ( w_6220 , w_6221 );
and ( w_6221 , \2645_b1 , \2645_b0 );
or ( \2801_b1 , \2800_b1 , \2650_b1 );
xor ( \2801_b0 , \2800_b0 , w_6222 );
not ( w_6222 , w_6223 );
and ( w_6223 , \2650_b1 , \2650_b0 );
or ( \2802_b1 , \2798_b1 , \2801_b1 );
not ( \2801_b1 , w_6224 );
and ( \2802_b0 , \2798_b0 , w_6225 );
and ( w_6224 , w_6225 , \2801_b0 );
or ( \2803_b1 , \2782_b1 , \2801_b1 );
not ( \2801_b1 , w_6226 );
and ( \2803_b0 , \2782_b0 , w_6227 );
and ( w_6226 , w_6227 , \2801_b0 );
or ( \2805_b1 , \1477_b1 , \1431_b1 );
not ( \1431_b1 , w_6228 );
and ( \2805_b0 , \1477_b0 , w_6229 );
and ( w_6228 , w_6229 , \1431_b0 );
or ( \2806_b1 , \1454_b1 , \1429_b1 );
not ( \1429_b1 , w_6230 );
and ( \2806_b0 , \1454_b0 , w_6231 );
and ( w_6230 , w_6231 , \1429_b0 );
or ( \2807_b1 , \2805_b1 , w_6233 );
not ( w_6233 , w_6234 );
and ( \2807_b0 , \2805_b0 , w_6235 );
and ( w_6234 ,  , w_6235 );
buf ( w_6233 , \2806_b1 );
not ( w_6233 , w_6236 );
not (  , w_6237 );
and ( w_6236 , w_6237 , \2806_b0 );
or ( \2808_b1 , \2807_b1 , w_6238 );
xor ( \2808_b0 , \2807_b0 , w_6240 );
not ( w_6240 , w_6241 );
and ( w_6241 , w_6238 , w_6239 );
buf ( w_6238 , \1438_b1 );
not ( w_6238 , w_6242 );
not ( w_6239 , w_6243 );
and ( w_6242 , w_6243 , \1438_b0 );
or ( \2809_b1 , \1498_b1 , \1673_b1 );
not ( \1673_b1 , w_6244 );
and ( \2809_b0 , \1498_b0 , w_6245 );
and ( w_6244 , w_6245 , \1673_b0 );
buf ( \2810_b1 , \2809_b1 );
not ( \2810_b1 , w_6246 );
not ( \2810_b0 , w_6247 );
and ( w_6246 , w_6247 , \2809_b0 );
or ( \2811_b1 , \2810_b1 , \1681_b1 );
not ( \1681_b1 , w_6248 );
and ( \2811_b0 , \2810_b0 , w_6249 );
and ( w_6248 , w_6249 , \1681_b0 );
or ( \2812_b1 , \2808_b1 , \2811_b1 );
not ( \2811_b1 , w_6250 );
and ( \2812_b0 , \2808_b0 , w_6251 );
and ( w_6250 , w_6251 , \2811_b0 );
or ( \2813_b1 , \1407_b1 , \1475_b1 );
not ( \1475_b1 , w_6252 );
and ( \2813_b0 , \1407_b0 , w_6253 );
and ( w_6252 , w_6253 , \1475_b0 );
or ( \2814_b1 , \1416_b1 , \1473_b1 );
not ( \1473_b1 , w_6254 );
and ( \2814_b0 , \1416_b0 , w_6255 );
and ( w_6254 , w_6255 , \1473_b0 );
or ( \2815_b1 , \2813_b1 , w_6257 );
not ( w_6257 , w_6258 );
and ( \2815_b0 , \2813_b0 , w_6259 );
and ( w_6258 ,  , w_6259 );
buf ( w_6257 , \2814_b1 );
not ( w_6257 , w_6260 );
not (  , w_6261 );
and ( w_6260 , w_6261 , \2814_b0 );
or ( \2816_b1 , \2815_b1 , w_6262 );
xor ( \2816_b0 , \2815_b0 , w_6264 );
not ( w_6264 , w_6265 );
and ( w_6265 , w_6262 , w_6263 );
buf ( w_6262 , \1482_b1 );
not ( w_6262 , w_6266 );
not ( w_6263 , w_6267 );
and ( w_6266 , w_6267 , \1482_b0 );
or ( \2817_b1 , \2812_b1 , \2816_b1 );
not ( \2816_b1 , w_6268 );
and ( \2817_b0 , \2812_b0 , w_6269 );
and ( w_6268 , w_6269 , \2816_b0 );
or ( \2818_b1 , \1553_b1 , \1675_b1 );
not ( \1675_b1 , w_6270 );
and ( \2818_b0 , \1553_b0 , w_6271 );
and ( w_6270 , w_6271 , \1675_b0 );
or ( \2819_b1 , \1533_b1 , \1673_b1 );
not ( \1673_b1 , w_6272 );
and ( \2819_b0 , \1533_b0 , w_6273 );
and ( w_6272 , w_6273 , \1673_b0 );
or ( \2820_b1 , \2818_b1 , w_6275 );
not ( w_6275 , w_6276 );
and ( \2820_b0 , \2818_b0 , w_6277 );
and ( w_6276 ,  , w_6277 );
buf ( w_6275 , \2819_b1 );
not ( w_6275 , w_6278 );
not (  , w_6279 );
and ( w_6278 , w_6279 , \2819_b0 );
or ( \2821_b1 , \2820_b1 , w_6280 );
xor ( \2821_b0 , \2820_b0 , w_6282 );
not ( w_6282 , w_6283 );
and ( w_6283 , w_6280 , w_6281 );
buf ( w_6280 , \1681_b1 );
not ( w_6280 , w_6284 );
not ( w_6281 , w_6285 );
and ( w_6284 , w_6285 , \1681_b0 );
or ( \2822_b1 , \2816_b1 , \2821_b1 );
not ( \2821_b1 , w_6286 );
and ( \2822_b0 , \2816_b0 , w_6287 );
and ( w_6286 , w_6287 , \2821_b0 );
or ( \2823_b1 , \2812_b1 , \2821_b1 );
not ( \2821_b1 , w_6288 );
and ( \2823_b0 , \2812_b0 , w_6289 );
and ( w_6288 , w_6289 , \2821_b0 );
or ( \2825_b1 , \2693_b1 , \2697_b1 );
xor ( \2825_b0 , \2693_b0 , w_6290 );
not ( w_6290 , w_6291 );
and ( w_6291 , \2697_b1 , \2697_b0 );
or ( \2826_b1 , \2825_b1 , \2702_b1 );
xor ( \2826_b0 , \2825_b0 , w_6292 );
not ( w_6292 , w_6293 );
and ( w_6293 , \2702_b1 , \2702_b0 );
or ( \2827_b1 , \2824_b1 , \2826_b1 );
not ( \2826_b1 , w_6294 );
and ( \2827_b0 , \2824_b0 , w_6295 );
and ( w_6294 , w_6295 , \2826_b0 );
or ( \2828_b1 , \2657_b1 , \2661_b1 );
xor ( \2828_b0 , \2657_b0 , w_6296 );
not ( w_6296 , w_6297 );
and ( w_6297 , \2661_b1 , \2661_b0 );
or ( \2829_b1 , \2828_b1 , \2666_b1 );
xor ( \2829_b0 , \2828_b0 , w_6298 );
not ( w_6298 , w_6299 );
and ( w_6299 , \2666_b1 , \2666_b0 );
or ( \2830_b1 , \2826_b1 , \2829_b1 );
not ( \2829_b1 , w_6300 );
and ( \2830_b0 , \2826_b0 , w_6301 );
and ( w_6300 , w_6301 , \2829_b0 );
or ( \2831_b1 , \2824_b1 , \2829_b1 );
not ( \2829_b1 , w_6302 );
and ( \2831_b0 , \2824_b0 , w_6303 );
and ( w_6302 , w_6303 , \2829_b0 );
or ( \2833_b1 , \2804_b1 , \2832_b1 );
not ( \2832_b1 , w_6304 );
and ( \2833_b0 , \2804_b0 , w_6305 );
and ( w_6304 , w_6305 , \2832_b0 );
or ( \2834_b1 , \2653_b1 , \2669_b1 );
xor ( \2834_b0 , \2653_b0 , w_6306 );
not ( w_6306 , w_6307 );
and ( w_6307 , \2669_b1 , \2669_b0 );
or ( \2835_b1 , \2834_b1 , \2678_b1 );
xor ( \2835_b0 , \2834_b0 , w_6308 );
not ( w_6308 , w_6309 );
and ( w_6309 , \2678_b1 , \2678_b0 );
or ( \2836_b1 , \2832_b1 , \2835_b1 );
not ( \2835_b1 , w_6310 );
and ( \2836_b0 , \2832_b0 , w_6311 );
and ( w_6310 , w_6311 , \2835_b0 );
or ( \2837_b1 , \2804_b1 , \2835_b1 );
not ( \2835_b1 , w_6312 );
and ( \2837_b0 , \2804_b0 , w_6313 );
and ( w_6312 , w_6313 , \2835_b0 );
or ( \2839_b1 , \2603_b1 , \2605_b1 );
xor ( \2839_b0 , \2603_b0 , w_6314 );
not ( w_6314 , w_6315 );
and ( w_6315 , \2605_b1 , \2605_b0 );
or ( \2840_b1 , \2839_b1 , \2608_b1 );
xor ( \2840_b0 , \2839_b0 , w_6316 );
not ( w_6316 , w_6317 );
and ( w_6317 , \2608_b1 , \2608_b0 );
or ( \2841_b1 , \2838_b1 , \2840_b1 );
not ( \2840_b1 , w_6318 );
and ( \2841_b0 , \2838_b0 , w_6319 );
and ( w_6318 , w_6319 , \2840_b0 );
or ( \2842_b1 , \2681_b1 , \2683_b1 );
xor ( \2842_b0 , \2681_b0 , w_6320 );
not ( w_6320 , w_6321 );
and ( w_6321 , \2683_b1 , \2683_b0 );
or ( \2843_b1 , \2842_b1 , \2686_b1 );
xor ( \2843_b0 , \2842_b0 , w_6322 );
not ( w_6322 , w_6323 );
and ( w_6323 , \2686_b1 , \2686_b0 );
or ( \2844_b1 , \2840_b1 , \2843_b1 );
not ( \2843_b1 , w_6324 );
and ( \2844_b0 , \2840_b0 , w_6325 );
and ( w_6324 , w_6325 , \2843_b0 );
or ( \2845_b1 , \2838_b1 , \2843_b1 );
not ( \2843_b1 , w_6326 );
and ( \2845_b0 , \2838_b0 , w_6327 );
and ( w_6326 , w_6327 , \2843_b0 );
or ( \2847_b1 , \2611_b1 , \2613_b1 );
xor ( \2847_b0 , \2611_b0 , w_6328 );
not ( w_6328 , w_6329 );
and ( w_6329 , \2613_b1 , \2613_b0 );
or ( \2848_b1 , \2847_b1 , \2616_b1 );
xor ( \2848_b0 , \2847_b0 , w_6330 );
not ( w_6330 , w_6331 );
and ( w_6331 , \2616_b1 , \2616_b0 );
or ( \2849_b1 , \2846_b1 , \2848_b1 );
not ( \2848_b1 , w_6332 );
and ( \2849_b0 , \2846_b0 , w_6333 );
and ( w_6332 , w_6333 , \2848_b0 );
or ( \2850_b1 , \2689_b1 , \2748_b1 );
xor ( \2850_b0 , \2689_b0 , w_6334 );
not ( w_6334 , w_6335 );
and ( w_6335 , \2748_b1 , \2748_b0 );
or ( \2851_b1 , \2850_b1 , \2751_b1 );
xor ( \2851_b0 , \2850_b0 , w_6336 );
not ( w_6336 , w_6337 );
and ( w_6337 , \2751_b1 , \2751_b0 );
or ( \2852_b1 , \2848_b1 , \2851_b1 );
not ( \2851_b1 , w_6338 );
and ( \2852_b0 , \2848_b0 , w_6339 );
and ( w_6338 , w_6339 , \2851_b0 );
or ( \2853_b1 , \2846_b1 , \2851_b1 );
not ( \2851_b1 , w_6340 );
and ( \2853_b0 , \2846_b0 , w_6341 );
and ( w_6340 , w_6341 , \2851_b0 );
or ( \2855_b1 , \2766_b1 , \2854_b1 );
not ( \2854_b1 , w_6342 );
and ( \2855_b0 , \2766_b0 , w_6343 );
and ( w_6342 , w_6343 , \2854_b0 );
or ( \2856_b1 , \2766_b1 , \2854_b1 );
xor ( \2856_b0 , \2766_b0 , w_6344 );
not ( w_6344 , w_6345 );
and ( w_6345 , \2854_b1 , \2854_b0 );
or ( \2857_b1 , \2846_b1 , \2848_b1 );
xor ( \2857_b0 , \2846_b0 , w_6346 );
not ( w_6346 , w_6347 );
and ( w_6347 , \2848_b1 , \2848_b0 );
or ( \2858_b1 , \2857_b1 , \2851_b1 );
xor ( \2858_b0 , \2857_b0 , w_6348 );
not ( w_6348 , w_6349 );
and ( w_6349 , \2851_b1 , \2851_b0 );
or ( \2859_b1 , \1462_b1 , \1336_b1 );
not ( \1336_b1 , w_6350 );
and ( \2859_b0 , \1462_b0 , w_6351 );
and ( w_6350 , w_6351 , \1336_b0 );
or ( \2860_b1 , \1376_b1 , \1333_b1 );
not ( \1333_b1 , w_6352 );
and ( \2860_b0 , \1376_b0 , w_6353 );
and ( w_6352 , w_6353 , \1333_b0 );
or ( \2861_b1 , \2859_b1 , w_6355 );
not ( w_6355 , w_6356 );
and ( \2861_b0 , \2859_b0 , w_6357 );
and ( w_6356 ,  , w_6357 );
buf ( w_6355 , \2860_b1 );
not ( w_6355 , w_6358 );
not (  , w_6359 );
and ( w_6358 , w_6359 , \2860_b0 );
or ( \2862_b1 , \2861_b1 , w_6360 );
xor ( \2862_b0 , \2861_b0 , w_6362 );
not ( w_6362 , w_6363 );
and ( w_6363 , w_6360 , w_6361 );
buf ( w_6360 , \1332_b1 );
not ( w_6360 , w_6364 );
not ( w_6361 , w_6365 );
and ( w_6364 , w_6365 , \1332_b0 );
or ( \2863_b1 , \1616_b1 , \1382_b1 );
not ( \1382_b1 , w_6366 );
and ( \2863_b0 , \1616_b0 , w_6367 );
and ( w_6366 , w_6367 , \1382_b0 );
or ( \2864_b1 , \1391_b1 , \1380_b1 );
not ( \1380_b1 , w_6368 );
and ( \2864_b0 , \1391_b0 , w_6369 );
and ( w_6368 , w_6369 , \1380_b0 );
or ( \2865_b1 , \2863_b1 , w_6371 );
not ( w_6371 , w_6372 );
and ( \2865_b0 , \2863_b0 , w_6373 );
and ( w_6372 ,  , w_6373 );
buf ( w_6371 , \2864_b1 );
not ( w_6371 , w_6374 );
not (  , w_6375 );
and ( w_6374 , w_6375 , \2864_b0 );
or ( \2866_b1 , \2865_b1 , w_6376 );
xor ( \2866_b0 , \2865_b0 , w_6378 );
not ( w_6378 , w_6379 );
and ( w_6379 , w_6376 , w_6377 );
buf ( w_6376 , \1389_b1 );
not ( w_6376 , w_6380 );
not ( w_6377 , w_6381 );
and ( w_6380 , w_6381 , \1389_b0 );
or ( \2867_b1 , \2862_b1 , \2866_b1 );
not ( \2866_b1 , w_6382 );
and ( \2867_b0 , \2862_b0 , w_6383 );
and ( w_6382 , w_6383 , \2866_b0 );
or ( \2868_b1 , \1533_b1 , \1397_b1 );
not ( \1397_b1 , w_6384 );
and ( \2868_b0 , \1533_b0 , w_6385 );
and ( w_6384 , w_6385 , \1397_b0 );
or ( \2869_b1 , \1540_b1 , \1395_b1 );
not ( \1395_b1 , w_6386 );
and ( \2869_b0 , \1540_b0 , w_6387 );
and ( w_6386 , w_6387 , \1395_b0 );
or ( \2870_b1 , \2868_b1 , w_6389 );
not ( w_6389 , w_6390 );
and ( \2870_b0 , \2868_b0 , w_6391 );
and ( w_6390 ,  , w_6391 );
buf ( w_6389 , \2869_b1 );
not ( w_6389 , w_6392 );
not (  , w_6393 );
and ( w_6392 , w_6393 , \2869_b0 );
or ( \2871_b1 , \2870_b1 , w_6394 );
xor ( \2871_b0 , \2870_b0 , w_6396 );
not ( w_6396 , w_6397 );
and ( w_6397 , w_6394 , w_6395 );
buf ( w_6394 , \1404_b1 );
not ( w_6394 , w_6398 );
not ( w_6395 , w_6399 );
and ( w_6398 , w_6399 , \1404_b0 );
or ( \2872_b1 , \2866_b1 , \2871_b1 );
not ( \2871_b1 , w_6400 );
and ( \2872_b0 , \2866_b0 , w_6401 );
and ( w_6400 , w_6401 , \2871_b0 );
or ( \2873_b1 , \2862_b1 , \2871_b1 );
not ( \2871_b1 , w_6402 );
and ( \2873_b0 , \2862_b0 , w_6403 );
and ( w_6402 , w_6403 , \2871_b0 );
or ( \2875_b1 , \1368_b1 , \1444_b1 );
not ( \1444_b1 , w_6404 );
and ( \2875_b0 , \1368_b0 , w_6405 );
and ( w_6404 , w_6405 , \1444_b0 );
or ( \2876_b1 , \1470_b1 , \1442_b1 );
not ( \1442_b1 , w_6406 );
and ( \2876_b0 , \1470_b0 , w_6407 );
and ( w_6406 , w_6407 , \1442_b0 );
or ( \2877_b1 , \2875_b1 , w_6409 );
not ( w_6409 , w_6410 );
and ( \2877_b0 , \2875_b0 , w_6411 );
and ( w_6410 ,  , w_6411 );
buf ( w_6409 , \2876_b1 );
not ( w_6409 , w_6412 );
not (  , w_6413 );
and ( w_6412 , w_6413 , \2876_b0 );
or ( \2878_b1 , \2877_b1 , w_6414 );
xor ( \2878_b0 , \2877_b0 , w_6416 );
not ( w_6416 , w_6417 );
and ( w_6417 , w_6414 , w_6415 );
buf ( w_6414 , \1451_b1 );
not ( w_6414 , w_6418 );
not ( w_6415 , w_6419 );
and ( w_6418 , w_6419 , \1451_b0 );
or ( \2879_b1 , \1399_b1 , \1349_b1 );
not ( \1349_b1 , w_6420 );
and ( \2879_b0 , \1399_b0 , w_6421 );
and ( w_6420 , w_6421 , \1349_b0 );
or ( \2880_b1 , \1359_b1 , \1347_b1 );
not ( \1347_b1 , w_6422 );
and ( \2880_b0 , \1359_b0 , w_6423 );
and ( w_6422 , w_6423 , \1347_b0 );
or ( \2881_b1 , \2879_b1 , w_6425 );
not ( w_6425 , w_6426 );
and ( \2881_b0 , \2879_b0 , w_6427 );
and ( w_6426 ,  , w_6427 );
buf ( w_6425 , \2880_b1 );
not ( w_6425 , w_6428 );
not (  , w_6429 );
and ( w_6428 , w_6429 , \2880_b0 );
or ( \2882_b1 , \2881_b1 , w_6430 );
xor ( \2882_b0 , \2881_b0 , w_6432 );
not ( w_6432 , w_6433 );
and ( w_6433 , w_6430 , w_6431 );
buf ( w_6430 , \1356_b1 );
not ( w_6430 , w_6434 );
not ( w_6431 , w_6435 );
and ( w_6434 , w_6435 , \1356_b0 );
or ( \2883_b1 , \2878_b1 , \2882_b1 );
not ( \2882_b1 , w_6436 );
and ( \2883_b0 , \2878_b0 , w_6437 );
and ( w_6436 , w_6437 , \2882_b0 );
or ( \2884_b1 , \1517_b1 , \1366_b1 );
not ( \1366_b1 , w_6438 );
and ( \2884_b0 , \1517_b0 , w_6439 );
and ( w_6438 , w_6439 , \1366_b0 );
or ( \2885_b1 , \1526_b1 , \1364_b1 );
not ( \1364_b1 , w_6440 );
and ( \2885_b0 , \1526_b0 , w_6441 );
and ( w_6440 , w_6441 , \1364_b0 );
or ( \2886_b1 , \2884_b1 , w_6443 );
not ( w_6443 , w_6444 );
and ( \2886_b0 , \2884_b0 , w_6445 );
and ( w_6444 ,  , w_6445 );
buf ( w_6443 , \2885_b1 );
not ( w_6443 , w_6446 );
not (  , w_6447 );
and ( w_6446 , w_6447 , \2885_b0 );
or ( \2887_b1 , \2886_b1 , w_6448 );
xor ( \2887_b0 , \2886_b0 , w_6450 );
not ( w_6450 , w_6451 );
and ( w_6451 , w_6448 , w_6449 );
buf ( w_6448 , \1373_b1 );
not ( w_6448 , w_6452 );
not ( w_6449 , w_6453 );
and ( w_6452 , w_6453 , \1373_b0 );
or ( \2888_b1 , \2882_b1 , \2887_b1 );
not ( \2887_b1 , w_6454 );
and ( \2888_b0 , \2882_b0 , w_6455 );
and ( w_6454 , w_6455 , \2887_b0 );
or ( \2889_b1 , \2878_b1 , \2887_b1 );
not ( \2887_b1 , w_6456 );
and ( \2889_b0 , \2878_b0 , w_6457 );
and ( w_6456 , w_6457 , \2887_b0 );
or ( \2891_b1 , \2874_b1 , \2890_b1 );
not ( \2890_b1 , w_6458 );
and ( \2891_b0 , \2874_b0 , w_6459 );
and ( w_6458 , w_6459 , \2890_b0 );
or ( \2892_b1 , \2718_b1 , \2722_b1 );
xor ( \2892_b0 , \2718_b0 , w_6460 );
not ( w_6460 , w_6461 );
and ( w_6461 , \2722_b1 , \2722_b0 );
or ( \2893_b1 , \2892_b1 , \2675_b1 );
xor ( \2893_b0 , \2892_b0 , w_6462 );
not ( w_6462 , w_6463 );
and ( w_6463 , \2675_b1 , \2675_b0 );
or ( \2894_b1 , \2890_b1 , \2893_b1 );
not ( \2893_b1 , w_6464 );
and ( \2894_b0 , \2890_b0 , w_6465 );
and ( w_6464 , w_6465 , \2893_b0 );
or ( \2895_b1 , \2874_b1 , \2893_b1 );
not ( \2893_b1 , w_6466 );
and ( \2895_b0 , \2874_b0 , w_6467 );
and ( w_6466 , w_6467 , \2893_b0 );
or ( \2897_b1 , \2714_b1 , \2726_b1 );
xor ( \2897_b0 , \2714_b0 , w_6468 );
not ( w_6468 , w_6469 );
and ( w_6469 , \2726_b1 , \2726_b0 );
or ( \2898_b1 , \2897_b1 , \2731_b1 );
xor ( \2898_b0 , \2897_b0 , w_6470 );
not ( w_6470 , w_6471 );
and ( w_6471 , \2731_b1 , \2731_b0 );
or ( \2899_b1 , \2896_b1 , \2898_b1 );
not ( \2898_b1 , w_6472 );
and ( \2899_b0 , \2896_b0 , w_6473 );
and ( w_6472 , w_6473 , \2898_b0 );
or ( \2900_b1 , \2782_b1 , \2798_b1 );
xor ( \2900_b0 , \2782_b0 , w_6474 );
not ( w_6474 , w_6475 );
and ( w_6475 , \2798_b1 , \2798_b0 );
or ( \2901_b1 , \2900_b1 , \2801_b1 );
xor ( \2901_b0 , \2900_b0 , w_6476 );
not ( w_6476 , w_6477 );
and ( w_6477 , \2801_b1 , \2801_b0 );
or ( \2902_b1 , \2898_b1 , \2901_b1 );
not ( \2901_b1 , w_6478 );
and ( \2902_b0 , \2898_b0 , w_6479 );
and ( w_6478 , w_6479 , \2901_b0 );
or ( \2903_b1 , \2896_b1 , \2901_b1 );
not ( \2901_b1 , w_6480 );
and ( \2903_b0 , \2896_b0 , w_6481 );
and ( w_6480 , w_6481 , \2901_b0 );
or ( \2905_b1 , \2705_b1 , \2707_b1 );
xor ( \2905_b0 , \2705_b0 , w_6482 );
not ( w_6482 , w_6483 );
and ( w_6483 , \2707_b1 , \2707_b0 );
or ( \2906_b1 , \2905_b1 , \2710_b1 );
xor ( \2906_b0 , \2905_b0 , w_6484 );
not ( w_6484 , w_6485 );
and ( w_6485 , \2710_b1 , \2710_b0 );
or ( \2907_b1 , \2904_b1 , \2906_b1 );
not ( \2906_b1 , w_6486 );
and ( \2907_b0 , \2904_b0 , w_6487 );
and ( w_6486 , w_6487 , \2906_b0 );
or ( \2908_b1 , \2734_b1 , \2736_b1 );
xor ( \2908_b0 , \2734_b0 , w_6488 );
not ( w_6488 , w_6489 );
and ( w_6489 , \2736_b1 , \2736_b0 );
or ( \2909_b1 , \2908_b1 , \2739_b1 );
xor ( \2909_b0 , \2908_b0 , w_6490 );
not ( w_6490 , w_6491 );
and ( w_6491 , \2739_b1 , \2739_b0 );
or ( \2910_b1 , \2906_b1 , \2909_b1 );
not ( \2909_b1 , w_6492 );
and ( \2910_b0 , \2906_b0 , w_6493 );
and ( w_6492 , w_6493 , \2909_b0 );
or ( \2911_b1 , \2904_b1 , \2909_b1 );
not ( \2909_b1 , w_6494 );
and ( \2911_b0 , \2904_b0 , w_6495 );
and ( w_6494 , w_6495 , \2909_b0 );
or ( \2913_b1 , \2713_b1 , \2742_b1 );
xor ( \2913_b0 , \2713_b0 , w_6496 );
not ( w_6496 , w_6497 );
and ( w_6497 , \2742_b1 , \2742_b0 );
or ( \2914_b1 , \2913_b1 , \2745_b1 );
xor ( \2914_b0 , \2913_b0 , w_6498 );
not ( w_6498 , w_6499 );
and ( w_6499 , \2745_b1 , \2745_b0 );
or ( \2915_b1 , \2912_b1 , \2914_b1 );
not ( \2914_b1 , w_6500 );
and ( \2915_b0 , \2912_b0 , w_6501 );
and ( w_6500 , w_6501 , \2914_b0 );
or ( \2916_b1 , \2838_b1 , \2840_b1 );
xor ( \2916_b0 , \2838_b0 , w_6502 );
not ( w_6502 , w_6503 );
and ( w_6503 , \2840_b1 , \2840_b0 );
or ( \2917_b1 , \2916_b1 , \2843_b1 );
xor ( \2917_b0 , \2916_b0 , w_6504 );
not ( w_6504 , w_6505 );
and ( w_6505 , \2843_b1 , \2843_b0 );
or ( \2918_b1 , \2914_b1 , \2917_b1 );
not ( \2917_b1 , w_6506 );
and ( \2918_b0 , \2914_b0 , w_6507 );
and ( w_6506 , w_6507 , \2917_b0 );
or ( \2919_b1 , \2912_b1 , \2917_b1 );
not ( \2917_b1 , w_6508 );
and ( \2919_b0 , \2912_b0 , w_6509 );
and ( w_6508 , w_6509 , \2917_b0 );
or ( \2921_b1 , \2858_b1 , \2920_b1 );
not ( \2920_b1 , w_6510 );
and ( \2921_b0 , \2858_b0 , w_6511 );
and ( w_6510 , w_6511 , \2920_b0 );
or ( \2922_b1 , \2858_b1 , \2920_b1 );
xor ( \2922_b0 , \2858_b0 , w_6512 );
not ( w_6512 , w_6513 );
and ( w_6513 , \2920_b1 , \2920_b0 );
or ( \2923_b1 , \2808_b1 , \2811_b1 );
xor ( \2923_b0 , \2808_b0 , w_6514 );
not ( w_6514 , w_6515 );
and ( w_6515 , \2811_b1 , \2811_b0 );
or ( \2924_b1 , \1416_b1 , \1460_b1 );
not ( \1460_b1 , w_6516 );
and ( \2924_b0 , \1416_b0 , w_6517 );
and ( w_6516 , w_6517 , \1460_b0 );
or ( \2925_b1 , \1586_b1 , \1458_b1 );
not ( \1458_b1 , w_6518 );
and ( \2925_b0 , \1586_b0 , w_6519 );
and ( w_6518 , w_6519 , \1458_b0 );
or ( \2926_b1 , \2924_b1 , w_6521 );
not ( w_6521 , w_6522 );
and ( \2926_b0 , \2924_b0 , w_6523 );
and ( w_6522 ,  , w_6523 );
buf ( w_6521 , \2925_b1 );
not ( w_6521 , w_6524 );
not (  , w_6525 );
and ( w_6524 , w_6525 , \2925_b0 );
or ( \2927_b1 , \2926_b1 , w_6526 );
xor ( \2927_b0 , \2926_b0 , w_6528 );
not ( w_6528 , w_6529 );
and ( w_6529 , w_6526 , w_6527 );
buf ( w_6526 , \1467_b1 );
not ( w_6526 , w_6530 );
not ( w_6527 , w_6531 );
and ( w_6530 , w_6531 , \1467_b0 );
or ( \2928_b1 , \2923_b1 , \2927_b1 );
not ( \2927_b1 , w_6532 );
and ( \2928_b0 , \2923_b0 , w_6533 );
and ( w_6532 , w_6533 , \2927_b0 );
or ( \2929_b1 , \1622_b1 , \1475_b1 );
not ( \1475_b1 , w_6534 );
and ( \2929_b0 , \1622_b0 , w_6535 );
and ( w_6534 , w_6535 , \1475_b0 );
or ( \2930_b1 , \1407_b1 , \1473_b1 );
not ( \1473_b1 , w_6536 );
and ( \2930_b0 , \1407_b0 , w_6537 );
and ( w_6536 , w_6537 , \1473_b0 );
or ( \2931_b1 , \2929_b1 , w_6539 );
not ( w_6539 , w_6540 );
and ( \2931_b0 , \2929_b0 , w_6541 );
and ( w_6540 ,  , w_6541 );
buf ( w_6539 , \2930_b1 );
not ( w_6539 , w_6542 );
not (  , w_6543 );
and ( w_6542 , w_6543 , \2930_b0 );
or ( \2932_b1 , \2931_b1 , w_6544 );
xor ( \2932_b0 , \2931_b0 , w_6546 );
not ( w_6546 , w_6547 );
and ( w_6547 , w_6544 , w_6545 );
buf ( w_6544 , \1482_b1 );
not ( w_6544 , w_6548 );
not ( w_6545 , w_6549 );
and ( w_6548 , w_6549 , \1482_b0 );
or ( \2933_b1 , \2927_b1 , \2932_b1 );
not ( \2932_b1 , w_6550 );
and ( \2933_b0 , \2927_b0 , w_6551 );
and ( w_6550 , w_6551 , \2932_b0 );
or ( \2934_b1 , \2923_b1 , \2932_b1 );
not ( \2932_b1 , w_6552 );
and ( \2934_b0 , \2923_b0 , w_6553 );
and ( w_6552 , w_6553 , \2932_b0 );
or ( \2936_b1 , \2770_b1 , \2774_b1 );
xor ( \2936_b0 , \2770_b0 , w_6554 );
not ( w_6554 , w_6555 );
and ( w_6555 , \2774_b1 , \2774_b0 );
or ( \2937_b1 , \2936_b1 , \2779_b1 );
xor ( \2937_b0 , \2936_b0 , w_6556 );
not ( w_6556 , w_6557 );
and ( w_6557 , \2779_b1 , \2779_b0 );
or ( \2938_b1 , \2935_b1 , \2937_b1 );
not ( \2937_b1 , w_6558 );
and ( \2938_b0 , \2935_b0 , w_6559 );
and ( w_6558 , w_6559 , \2937_b0 );
or ( \2939_b1 , \2786_b1 , \2790_b1 );
xor ( \2939_b0 , \2786_b0 , w_6560 );
not ( w_6560 , w_6561 );
and ( w_6561 , \2790_b1 , \2790_b0 );
or ( \2940_b1 , \2939_b1 , \2795_b1 );
xor ( \2940_b0 , \2939_b0 , w_6562 );
not ( w_6562 , w_6563 );
and ( w_6563 , \2795_b1 , \2795_b0 );
or ( \2941_b1 , \2937_b1 , \2940_b1 );
not ( \2940_b1 , w_6564 );
and ( \2941_b0 , \2937_b0 , w_6565 );
and ( w_6564 , w_6565 , \2940_b0 );
or ( \2942_b1 , \2935_b1 , \2940_b1 );
not ( \2940_b1 , w_6566 );
and ( \2942_b0 , \2935_b0 , w_6567 );
and ( w_6566 , w_6567 , \2940_b0 );
or ( \2944_b1 , \1470_b1 , \1431_b1 );
not ( \1431_b1 , w_6568 );
and ( \2944_b0 , \1470_b0 , w_6569 );
and ( w_6568 , w_6569 , \1431_b0 );
or ( \2945_b1 , \1477_b1 , \1429_b1 );
not ( \1429_b1 , w_6570 );
and ( \2945_b0 , \1477_b0 , w_6571 );
and ( w_6570 , w_6571 , \1429_b0 );
or ( \2946_b1 , \2944_b1 , w_6573 );
not ( w_6573 , w_6574 );
and ( \2946_b0 , \2944_b0 , w_6575 );
and ( w_6574 ,  , w_6575 );
buf ( w_6573 , \2945_b1 );
not ( w_6573 , w_6576 );
not (  , w_6577 );
and ( w_6576 , w_6577 , \2945_b0 );
or ( \2947_b1 , \2946_b1 , w_6578 );
xor ( \2947_b0 , \2946_b0 , w_6580 );
not ( w_6580 , w_6581 );
and ( w_6581 , w_6578 , w_6579 );
buf ( w_6578 , \1438_b1 );
not ( w_6578 , w_6582 );
not ( w_6579 , w_6583 );
and ( w_6582 , w_6583 , \1438_b0 );
or ( \2948_b1 , \1359_b1 , \1444_b1 );
not ( \1444_b1 , w_6584 );
and ( \2948_b0 , \1359_b0 , w_6585 );
and ( w_6584 , w_6585 , \1444_b0 );
or ( \2949_b1 , \1368_b1 , \1442_b1 );
not ( \1442_b1 , w_6586 );
and ( \2949_b0 , \1368_b0 , w_6587 );
and ( w_6586 , w_6587 , \1442_b0 );
or ( \2950_b1 , \2948_b1 , w_6589 );
not ( w_6589 , w_6590 );
and ( \2950_b0 , \2948_b0 , w_6591 );
and ( w_6590 ,  , w_6591 );
buf ( w_6589 , \2949_b1 );
not ( w_6589 , w_6592 );
not (  , w_6593 );
and ( w_6592 , w_6593 , \2949_b0 );
or ( \2951_b1 , \2950_b1 , w_6594 );
xor ( \2951_b0 , \2950_b0 , w_6596 );
not ( w_6596 , w_6597 );
and ( w_6597 , w_6594 , w_6595 );
buf ( w_6594 , \1451_b1 );
not ( w_6594 , w_6598 );
not ( w_6595 , w_6599 );
and ( w_6598 , w_6599 , \1451_b0 );
or ( \2952_b1 , \2947_b1 , \2951_b1 );
not ( \2951_b1 , w_6600 );
and ( \2952_b0 , \2947_b0 , w_6601 );
and ( w_6600 , w_6601 , \2951_b0 );
or ( \2953_b1 , \2951_b1 , \2809_b1 );
not ( \2809_b1 , w_6602 );
and ( \2953_b0 , \2951_b0 , w_6603 );
and ( w_6602 , w_6603 , \2809_b0 );
or ( \2954_b1 , \2947_b1 , \2809_b1 );
not ( \2809_b1 , w_6604 );
and ( \2954_b0 , \2947_b0 , w_6605 );
and ( w_6604 , w_6605 , \2809_b0 );
or ( \2956_b1 , \1391_b1 , \1349_b1 );
not ( \1349_b1 , w_6606 );
and ( \2956_b0 , \1391_b0 , w_6607 );
and ( w_6606 , w_6607 , \1349_b0 );
or ( \2957_b1 , \1399_b1 , \1347_b1 );
not ( \1347_b1 , w_6608 );
and ( \2957_b0 , \1399_b0 , w_6609 );
and ( w_6608 , w_6609 , \1347_b0 );
or ( \2958_b1 , \2956_b1 , w_6611 );
not ( w_6611 , w_6612 );
and ( \2958_b0 , \2956_b0 , w_6613 );
and ( w_6612 ,  , w_6613 );
buf ( w_6611 , \2957_b1 );
not ( w_6611 , w_6614 );
not (  , w_6615 );
and ( w_6614 , w_6615 , \2957_b0 );
or ( \2959_b1 , \2958_b1 , w_6616 );
xor ( \2959_b0 , \2958_b0 , w_6618 );
not ( w_6618 , w_6619 );
and ( w_6619 , w_6616 , w_6617 );
buf ( w_6616 , \1356_b1 );
not ( w_6616 , w_6620 );
not ( w_6617 , w_6621 );
and ( w_6620 , w_6621 , \1356_b0 );
or ( \2960_b1 , \1540_b1 , \1366_b1 );
not ( \1366_b1 , w_6622 );
and ( \2960_b0 , \1540_b0 , w_6623 );
and ( w_6622 , w_6623 , \1366_b0 );
or ( \2961_b1 , \1517_b1 , \1364_b1 );
not ( \1364_b1 , w_6624 );
and ( \2961_b0 , \1517_b0 , w_6625 );
and ( w_6624 , w_6625 , \1364_b0 );
or ( \2962_b1 , \2960_b1 , w_6627 );
not ( w_6627 , w_6628 );
and ( \2962_b0 , \2960_b0 , w_6629 );
and ( w_6628 ,  , w_6629 );
buf ( w_6627 , \2961_b1 );
not ( w_6627 , w_6630 );
not (  , w_6631 );
and ( w_6630 , w_6631 , \2961_b0 );
or ( \2963_b1 , \2962_b1 , w_6632 );
xor ( \2963_b0 , \2962_b0 , w_6634 );
not ( w_6634 , w_6635 );
and ( w_6635 , w_6632 , w_6633 );
buf ( w_6632 , \1373_b1 );
not ( w_6632 , w_6636 );
not ( w_6633 , w_6637 );
and ( w_6636 , w_6637 , \1373_b0 );
or ( \2964_b1 , \2959_b1 , \2963_b1 );
not ( \2963_b1 , w_6638 );
and ( \2964_b0 , \2959_b0 , w_6639 );
and ( w_6638 , w_6639 , \2963_b0 );
or ( \2965_b1 , \1553_b1 , \1397_b1 );
not ( \1397_b1 , w_6640 );
and ( \2965_b0 , \1553_b0 , w_6641 );
and ( w_6640 , w_6641 , \1397_b0 );
or ( \2966_b1 , \1533_b1 , \1395_b1 );
not ( \1395_b1 , w_6642 );
and ( \2966_b0 , \1533_b0 , w_6643 );
and ( w_6642 , w_6643 , \1395_b0 );
or ( \2967_b1 , \2965_b1 , w_6645 );
not ( w_6645 , w_6646 );
and ( \2967_b0 , \2965_b0 , w_6647 );
and ( w_6646 ,  , w_6647 );
buf ( w_6645 , \2966_b1 );
not ( w_6645 , w_6648 );
not (  , w_6649 );
and ( w_6648 , w_6649 , \2966_b0 );
or ( \2968_b1 , \2967_b1 , w_6650 );
xor ( \2968_b0 , \2967_b0 , w_6652 );
not ( w_6652 , w_6653 );
and ( w_6653 , w_6650 , w_6651 );
buf ( w_6650 , \1404_b1 );
not ( w_6650 , w_6654 );
not ( w_6651 , w_6655 );
and ( w_6654 , w_6655 , \1404_b0 );
or ( \2969_b1 , \2963_b1 , \2968_b1 );
not ( \2968_b1 , w_6656 );
and ( \2969_b0 , \2963_b0 , w_6657 );
and ( w_6656 , w_6657 , \2968_b0 );
or ( \2970_b1 , \2959_b1 , \2968_b1 );
not ( \2968_b1 , w_6658 );
and ( \2970_b0 , \2959_b0 , w_6659 );
and ( w_6658 , w_6659 , \2968_b0 );
or ( \2972_b1 , \2955_b1 , \2971_b1 );
not ( \2971_b1 , w_6660 );
and ( \2972_b0 , \2955_b0 , w_6661 );
and ( w_6660 , w_6661 , \2971_b0 );
or ( \2973_b1 , \1498_b1 , \1675_b1 );
not ( \1675_b1 , w_6662 );
and ( \2973_b0 , \1498_b0 , w_6663 );
and ( w_6662 , w_6663 , \1675_b0 );
or ( \2974_b1 , \1553_b1 , \1673_b1 );
not ( \1673_b1 , w_6664 );
and ( \2974_b0 , \1553_b0 , w_6665 );
and ( w_6664 , w_6665 , \1673_b0 );
or ( \2975_b1 , \2973_b1 , w_6667 );
not ( w_6667 , w_6668 );
and ( \2975_b0 , \2973_b0 , w_6669 );
and ( w_6668 ,  , w_6669 );
buf ( w_6667 , \2974_b1 );
not ( w_6667 , w_6670 );
not (  , w_6671 );
and ( w_6670 , w_6671 , \2974_b0 );
or ( \2976_b1 , \2975_b1 , w_6672 );
xor ( \2976_b0 , \2975_b0 , w_6674 );
not ( w_6674 , w_6675 );
and ( w_6675 , w_6672 , w_6673 );
buf ( w_6672 , \1681_b1 );
not ( w_6672 , w_6676 );
not ( w_6673 , w_6677 );
and ( w_6676 , w_6677 , \1681_b0 );
or ( \2977_b1 , \2971_b1 , \2976_b1 );
not ( \2976_b1 , w_6678 );
and ( \2977_b0 , \2971_b0 , w_6679 );
and ( w_6678 , w_6679 , \2976_b0 );
or ( \2978_b1 , \2955_b1 , \2976_b1 );
not ( \2976_b1 , w_6680 );
and ( \2978_b0 , \2955_b0 , w_6681 );
and ( w_6680 , w_6681 , \2976_b0 );
or ( \2980_b1 , \2812_b1 , \2816_b1 );
xor ( \2980_b0 , \2812_b0 , w_6682 );
not ( w_6682 , w_6683 );
and ( w_6683 , \2816_b1 , \2816_b0 );
or ( \2981_b1 , \2980_b1 , \2821_b1 );
xor ( \2981_b0 , \2980_b0 , w_6684 );
not ( w_6684 , w_6685 );
and ( w_6685 , \2821_b1 , \2821_b0 );
or ( \2982_b1 , \2979_b1 , \2981_b1 );
not ( \2981_b1 , w_6686 );
and ( \2982_b0 , \2979_b0 , w_6687 );
and ( w_6686 , w_6687 , \2981_b0 );
or ( \2983_b1 , \2874_b1 , \2890_b1 );
xor ( \2983_b0 , \2874_b0 , w_6688 );
not ( w_6688 , w_6689 );
and ( w_6689 , \2890_b1 , \2890_b0 );
or ( \2984_b1 , \2983_b1 , \2893_b1 );
xor ( \2984_b0 , \2983_b0 , w_6690 );
not ( w_6690 , w_6691 );
and ( w_6691 , \2893_b1 , \2893_b0 );
or ( \2985_b1 , \2981_b1 , \2984_b1 );
not ( \2984_b1 , w_6692 );
and ( \2985_b0 , \2981_b0 , w_6693 );
and ( w_6692 , w_6693 , \2984_b0 );
or ( \2986_b1 , \2979_b1 , \2984_b1 );
not ( \2984_b1 , w_6694 );
and ( \2986_b0 , \2979_b0 , w_6695 );
and ( w_6694 , w_6695 , \2984_b0 );
or ( \2988_b1 , \2943_b1 , \2987_b1 );
not ( \2987_b1 , w_6696 );
and ( \2988_b0 , \2943_b0 , w_6697 );
and ( w_6696 , w_6697 , \2987_b0 );
or ( \2989_b1 , \2824_b1 , \2826_b1 );
xor ( \2989_b0 , \2824_b0 , w_6698 );
not ( w_6698 , w_6699 );
and ( w_6699 , \2826_b1 , \2826_b0 );
or ( \2990_b1 , \2989_b1 , \2829_b1 );
xor ( \2990_b0 , \2989_b0 , w_6700 );
not ( w_6700 , w_6701 );
and ( w_6701 , \2829_b1 , \2829_b0 );
or ( \2991_b1 , \2987_b1 , \2990_b1 );
not ( \2990_b1 , w_6702 );
and ( \2991_b0 , \2987_b0 , w_6703 );
and ( w_6702 , w_6703 , \2990_b0 );
or ( \2992_b1 , \2943_b1 , \2990_b1 );
not ( \2990_b1 , w_6704 );
and ( \2992_b0 , \2943_b0 , w_6705 );
and ( w_6704 , w_6705 , \2990_b0 );
or ( \2994_b1 , \2804_b1 , \2832_b1 );
xor ( \2994_b0 , \2804_b0 , w_6706 );
not ( w_6706 , w_6707 );
and ( w_6707 , \2832_b1 , \2832_b0 );
or ( \2995_b1 , \2994_b1 , \2835_b1 );
xor ( \2995_b0 , \2994_b0 , w_6708 );
not ( w_6708 , w_6709 );
and ( w_6709 , \2835_b1 , \2835_b0 );
or ( \2996_b1 , \2993_b1 , \2995_b1 );
not ( \2995_b1 , w_6710 );
and ( \2996_b0 , \2993_b0 , w_6711 );
and ( w_6710 , w_6711 , \2995_b0 );
or ( \2997_b1 , \2904_b1 , \2906_b1 );
xor ( \2997_b0 , \2904_b0 , w_6712 );
not ( w_6712 , w_6713 );
and ( w_6713 , \2906_b1 , \2906_b0 );
or ( \2998_b1 , \2997_b1 , \2909_b1 );
xor ( \2998_b0 , \2997_b0 , w_6714 );
not ( w_6714 , w_6715 );
and ( w_6715 , \2909_b1 , \2909_b0 );
or ( \2999_b1 , \2995_b1 , \2998_b1 );
not ( \2998_b1 , w_6716 );
and ( \2999_b0 , \2995_b0 , w_6717 );
and ( w_6716 , w_6717 , \2998_b0 );
or ( \3000_b1 , \2993_b1 , \2998_b1 );
not ( \2998_b1 , w_6718 );
and ( \3000_b0 , \2993_b0 , w_6719 );
and ( w_6718 , w_6719 , \2998_b0 );
or ( \3002_b1 , \2912_b1 , \2914_b1 );
xor ( \3002_b0 , \2912_b0 , w_6720 );
not ( w_6720 , w_6721 );
and ( w_6721 , \2914_b1 , \2914_b0 );
or ( \3003_b1 , \3002_b1 , \2917_b1 );
xor ( \3003_b0 , \3002_b0 , w_6722 );
not ( w_6722 , w_6723 );
and ( w_6723 , \2917_b1 , \2917_b0 );
or ( \3004_b1 , \3001_b1 , \3003_b1 );
not ( \3003_b1 , w_6724 );
and ( \3004_b0 , \3001_b0 , w_6725 );
and ( w_6724 , w_6725 , \3003_b0 );
or ( \3005_b1 , \3001_b1 , \3003_b1 );
xor ( \3005_b0 , \3001_b0 , w_6726 );
not ( w_6726 , w_6727 );
and ( w_6727 , \3003_b1 , \3003_b0 );
or ( \3006_b1 , \2993_b1 , \2995_b1 );
xor ( \3006_b0 , \2993_b0 , w_6728 );
not ( w_6728 , w_6729 );
and ( w_6729 , \2995_b1 , \2995_b0 );
or ( \3007_b1 , \3006_b1 , \2998_b1 );
xor ( \3007_b0 , \3006_b0 , w_6730 );
not ( w_6730 , w_6731 );
and ( w_6731 , \2998_b1 , \2998_b0 );
or ( \3008_b1 , \1454_b1 , \1336_b1 );
not ( \1336_b1 , w_6732 );
and ( \3008_b0 , \1454_b0 , w_6733 );
and ( w_6732 , w_6733 , \1336_b0 );
or ( \3009_b1 , \1462_b1 , \1333_b1 );
not ( \1333_b1 , w_6734 );
and ( \3009_b0 , \1462_b0 , w_6735 );
and ( w_6734 , w_6735 , \1333_b0 );
or ( \3010_b1 , \3008_b1 , w_6737 );
not ( w_6737 , w_6738 );
and ( \3010_b0 , \3008_b0 , w_6739 );
and ( w_6738 ,  , w_6739 );
buf ( w_6737 , \3009_b1 );
not ( w_6737 , w_6740 );
not (  , w_6741 );
and ( w_6740 , w_6741 , \3009_b0 );
or ( \3011_b1 , \3010_b1 , w_6742 );
xor ( \3011_b0 , \3010_b0 , w_6744 );
not ( w_6744 , w_6745 );
and ( w_6745 , w_6742 , w_6743 );
buf ( w_6742 , \1332_b1 );
not ( w_6742 , w_6746 );
not ( w_6743 , w_6747 );
and ( w_6746 , w_6747 , \1332_b0 );
or ( \3012_b1 , \1586_b1 , \1382_b1 );
not ( \1382_b1 , w_6748 );
and ( \3012_b0 , \1586_b0 , w_6749 );
and ( w_6748 , w_6749 , \1382_b0 );
or ( \3013_b1 , \1616_b1 , \1380_b1 );
not ( \1380_b1 , w_6750 );
and ( \3013_b0 , \1616_b0 , w_6751 );
and ( w_6750 , w_6751 , \1380_b0 );
or ( \3014_b1 , \3012_b1 , w_6753 );
not ( w_6753 , w_6754 );
and ( \3014_b0 , \3012_b0 , w_6755 );
and ( w_6754 ,  , w_6755 );
buf ( w_6753 , \3013_b1 );
not ( w_6753 , w_6756 );
not (  , w_6757 );
and ( w_6756 , w_6757 , \3013_b0 );
or ( \3015_b1 , \3014_b1 , w_6758 );
xor ( \3015_b0 , \3014_b0 , w_6760 );
not ( w_6760 , w_6761 );
and ( w_6761 , w_6758 , w_6759 );
buf ( w_6758 , \1389_b1 );
not ( w_6758 , w_6762 );
not ( w_6759 , w_6763 );
and ( w_6762 , w_6763 , \1389_b0 );
or ( \3016_b1 , \3011_b1 , \3015_b1 );
not ( \3015_b1 , w_6764 );
and ( \3016_b0 , \3011_b0 , w_6765 );
and ( w_6764 , w_6765 , \3015_b0 );
or ( \3017_b1 , \1407_b1 , \1460_b1 );
not ( \1460_b1 , w_6766 );
and ( \3017_b0 , \1407_b0 , w_6767 );
and ( w_6766 , w_6767 , \1460_b0 );
or ( \3018_b1 , \1416_b1 , \1458_b1 );
not ( \1458_b1 , w_6768 );
and ( \3018_b0 , \1416_b0 , w_6769 );
and ( w_6768 , w_6769 , \1458_b0 );
or ( \3019_b1 , \3017_b1 , w_6771 );
not ( w_6771 , w_6772 );
and ( \3019_b0 , \3017_b0 , w_6773 );
and ( w_6772 ,  , w_6773 );
buf ( w_6771 , \3018_b1 );
not ( w_6771 , w_6774 );
not (  , w_6775 );
and ( w_6774 , w_6775 , \3018_b0 );
or ( \3020_b1 , \3019_b1 , w_6776 );
xor ( \3020_b0 , \3019_b0 , w_6778 );
not ( w_6778 , w_6779 );
and ( w_6779 , w_6776 , w_6777 );
buf ( w_6776 , \1467_b1 );
not ( w_6776 , w_6780 );
not ( w_6777 , w_6781 );
and ( w_6780 , w_6781 , \1467_b0 );
or ( \3021_b1 , \3015_b1 , \3020_b1 );
not ( \3020_b1 , w_6782 );
and ( \3021_b0 , \3015_b0 , w_6783 );
and ( w_6782 , w_6783 , \3020_b0 );
or ( \3022_b1 , \3011_b1 , \3020_b1 );
not ( \3020_b1 , w_6784 );
and ( \3022_b0 , \3011_b0 , w_6785 );
and ( w_6784 , w_6785 , \3020_b0 );
or ( \3024_b1 , \2862_b1 , \2866_b1 );
xor ( \3024_b0 , \2862_b0 , w_6786 );
not ( w_6786 , w_6787 );
and ( w_6787 , \2866_b1 , \2866_b0 );
or ( \3025_b1 , \3024_b1 , \2871_b1 );
xor ( \3025_b0 , \3024_b0 , w_6788 );
not ( w_6788 , w_6789 );
and ( w_6789 , \2871_b1 , \2871_b0 );
or ( \3026_b1 , \3023_b1 , \3025_b1 );
not ( \3025_b1 , w_6790 );
and ( \3026_b0 , \3023_b0 , w_6791 );
and ( w_6790 , w_6791 , \3025_b0 );
or ( \3027_b1 , \2878_b1 , \2882_b1 );
xor ( \3027_b0 , \2878_b0 , w_6792 );
not ( w_6792 , w_6793 );
and ( w_6793 , \2882_b1 , \2882_b0 );
or ( \3028_b1 , \3027_b1 , \2887_b1 );
xor ( \3028_b0 , \3027_b0 , w_6794 );
not ( w_6794 , w_6795 );
and ( w_6795 , \2887_b1 , \2887_b0 );
or ( \3029_b1 , \3025_b1 , \3028_b1 );
not ( \3028_b1 , w_6796 );
and ( \3029_b0 , \3025_b0 , w_6797 );
and ( w_6796 , w_6797 , \3028_b0 );
or ( \3030_b1 , \3023_b1 , \3028_b1 );
not ( \3028_b1 , w_6798 );
and ( \3030_b0 , \3023_b0 , w_6799 );
and ( w_6798 , w_6799 , \3028_b0 );
or ( \3032_b1 , \1368_b1 , \1431_b1 );
not ( \1431_b1 , w_6800 );
and ( \3032_b0 , \1368_b0 , w_6801 );
and ( w_6800 , w_6801 , \1431_b0 );
or ( \3033_b1 , \1470_b1 , \1429_b1 );
not ( \1429_b1 , w_6802 );
and ( \3033_b0 , \1470_b0 , w_6803 );
and ( w_6802 , w_6803 , \1429_b0 );
or ( \3034_b1 , \3032_b1 , w_6805 );
not ( w_6805 , w_6806 );
and ( \3034_b0 , \3032_b0 , w_6807 );
and ( w_6806 ,  , w_6807 );
buf ( w_6805 , \3033_b1 );
not ( w_6805 , w_6808 );
not (  , w_6809 );
and ( w_6808 , w_6809 , \3033_b0 );
or ( \3035_b1 , \3034_b1 , w_6810 );
xor ( \3035_b0 , \3034_b0 , w_6812 );
not ( w_6812 , w_6813 );
and ( w_6813 , w_6810 , w_6811 );
buf ( w_6810 , \1438_b1 );
not ( w_6810 , w_6814 );
not ( w_6811 , w_6815 );
and ( w_6814 , w_6815 , \1438_b0 );
or ( \3036_b1 , \1498_b1 , \1395_b1 );
not ( \1395_b1 , w_6816 );
and ( \3036_b0 , \1498_b0 , w_6817 );
and ( w_6816 , w_6817 , \1395_b0 );
buf ( \3037_b1 , \3036_b1 );
not ( \3037_b1 , w_6818 );
not ( \3037_b0 , w_6819 );
and ( w_6818 , w_6819 , \3036_b0 );
or ( \3038_b1 , \3037_b1 , \1404_b1 );
not ( \1404_b1 , w_6820 );
and ( \3038_b0 , \3037_b0 , w_6821 );
and ( w_6820 , w_6821 , \1404_b0 );
or ( \3039_b1 , \3035_b1 , \3038_b1 );
not ( \3038_b1 , w_6822 );
and ( \3039_b0 , \3035_b0 , w_6823 );
and ( w_6822 , w_6823 , \3038_b0 );
or ( \3040_b1 , \1526_b1 , \1475_b1 );
not ( \1475_b1 , w_6824 );
and ( \3040_b0 , \1526_b0 , w_6825 );
and ( w_6824 , w_6825 , \1475_b0 );
or ( \3041_b1 , \1622_b1 , \1473_b1 );
not ( \1473_b1 , w_6826 );
and ( \3041_b0 , \1622_b0 , w_6827 );
and ( w_6826 , w_6827 , \1473_b0 );
or ( \3042_b1 , \3040_b1 , w_6829 );
not ( w_6829 , w_6830 );
and ( \3042_b0 , \3040_b0 , w_6831 );
and ( w_6830 ,  , w_6831 );
buf ( w_6829 , \3041_b1 );
not ( w_6829 , w_6832 );
not (  , w_6833 );
and ( w_6832 , w_6833 , \3041_b0 );
or ( \3043_b1 , \3042_b1 , w_6834 );
xor ( \3043_b0 , \3042_b0 , w_6836 );
not ( w_6836 , w_6837 );
and ( w_6837 , w_6834 , w_6835 );
buf ( w_6834 , \1482_b1 );
not ( w_6834 , w_6838 );
not ( w_6835 , w_6839 );
and ( w_6838 , w_6839 , \1482_b0 );
or ( \3044_b1 , \3039_b1 , \3043_b1 );
not ( \3043_b1 , w_6840 );
and ( \3044_b0 , \3039_b0 , w_6841 );
and ( w_6840 , w_6841 , \3043_b0 );
or ( \3045_b1 , \2947_b1 , \2951_b1 );
xor ( \3045_b0 , \2947_b0 , w_6842 );
not ( w_6842 , w_6843 );
and ( w_6843 , \2951_b1 , \2951_b0 );
or ( \3046_b1 , \3045_b1 , \2809_b1 );
xor ( \3046_b0 , \3045_b0 , w_6844 );
not ( w_6844 , w_6845 );
and ( w_6845 , \2809_b1 , \2809_b0 );
or ( \3047_b1 , \3043_b1 , \3046_b1 );
not ( \3046_b1 , w_6846 );
and ( \3047_b0 , \3043_b0 , w_6847 );
and ( w_6846 , w_6847 , \3046_b0 );
or ( \3048_b1 , \3039_b1 , \3046_b1 );
not ( \3046_b1 , w_6848 );
and ( \3048_b0 , \3039_b0 , w_6849 );
and ( w_6848 , w_6849 , \3046_b0 );
or ( \3050_b1 , \2955_b1 , \2971_b1 );
xor ( \3050_b0 , \2955_b0 , w_6850 );
not ( w_6850 , w_6851 );
and ( w_6851 , \2971_b1 , \2971_b0 );
or ( \3051_b1 , \3050_b1 , \2976_b1 );
xor ( \3051_b0 , \3050_b0 , w_6852 );
not ( w_6852 , w_6853 );
and ( w_6853 , \2976_b1 , \2976_b0 );
or ( \3052_b1 , \3049_b1 , \3051_b1 );
not ( \3051_b1 , w_6854 );
and ( \3052_b0 , \3049_b0 , w_6855 );
and ( w_6854 , w_6855 , \3051_b0 );
or ( \3053_b1 , \2923_b1 , \2927_b1 );
xor ( \3053_b0 , \2923_b0 , w_6856 );
not ( w_6856 , w_6857 );
and ( w_6857 , \2927_b1 , \2927_b0 );
or ( \3054_b1 , \3053_b1 , \2932_b1 );
xor ( \3054_b0 , \3053_b0 , w_6858 );
not ( w_6858 , w_6859 );
and ( w_6859 , \2932_b1 , \2932_b0 );
or ( \3055_b1 , \3051_b1 , \3054_b1 );
not ( \3054_b1 , w_6860 );
and ( \3055_b0 , \3051_b0 , w_6861 );
and ( w_6860 , w_6861 , \3054_b0 );
or ( \3056_b1 , \3049_b1 , \3054_b1 );
not ( \3054_b1 , w_6862 );
and ( \3056_b0 , \3049_b0 , w_6863 );
and ( w_6862 , w_6863 , \3054_b0 );
or ( \3058_b1 , \3031_b1 , \3057_b1 );
not ( \3057_b1 , w_6864 );
and ( \3058_b0 , \3031_b0 , w_6865 );
and ( w_6864 , w_6865 , \3057_b0 );
or ( \3059_b1 , \2935_b1 , \2937_b1 );
xor ( \3059_b0 , \2935_b0 , w_6866 );
not ( w_6866 , w_6867 );
and ( w_6867 , \2937_b1 , \2937_b0 );
or ( \3060_b1 , \3059_b1 , \2940_b1 );
xor ( \3060_b0 , \3059_b0 , w_6868 );
not ( w_6868 , w_6869 );
and ( w_6869 , \2940_b1 , \2940_b0 );
or ( \3061_b1 , \3057_b1 , \3060_b1 );
not ( \3060_b1 , w_6870 );
and ( \3061_b0 , \3057_b0 , w_6871 );
and ( w_6870 , w_6871 , \3060_b0 );
or ( \3062_b1 , \3031_b1 , \3060_b1 );
not ( \3060_b1 , w_6872 );
and ( \3062_b0 , \3031_b0 , w_6873 );
and ( w_6872 , w_6873 , \3060_b0 );
or ( \3064_b1 , \2896_b1 , \2898_b1 );
xor ( \3064_b0 , \2896_b0 , w_6874 );
not ( w_6874 , w_6875 );
and ( w_6875 , \2898_b1 , \2898_b0 );
or ( \3065_b1 , \3064_b1 , \2901_b1 );
xor ( \3065_b0 , \3064_b0 , w_6876 );
not ( w_6876 , w_6877 );
and ( w_6877 , \2901_b1 , \2901_b0 );
or ( \3066_b1 , \3063_b1 , \3065_b1 );
not ( \3065_b1 , w_6878 );
and ( \3066_b0 , \3063_b0 , w_6879 );
and ( w_6878 , w_6879 , \3065_b0 );
or ( \3067_b1 , \2943_b1 , \2987_b1 );
xor ( \3067_b0 , \2943_b0 , w_6880 );
not ( w_6880 , w_6881 );
and ( w_6881 , \2987_b1 , \2987_b0 );
or ( \3068_b1 , \3067_b1 , \2990_b1 );
xor ( \3068_b0 , \3067_b0 , w_6882 );
not ( w_6882 , w_6883 );
and ( w_6883 , \2990_b1 , \2990_b0 );
or ( \3069_b1 , \3065_b1 , \3068_b1 );
not ( \3068_b1 , w_6884 );
and ( \3069_b0 , \3065_b0 , w_6885 );
and ( w_6884 , w_6885 , \3068_b0 );
or ( \3070_b1 , \3063_b1 , \3068_b1 );
not ( \3068_b1 , w_6886 );
and ( \3070_b0 , \3063_b0 , w_6887 );
and ( w_6886 , w_6887 , \3068_b0 );
or ( \3072_b1 , \3007_b1 , \3071_b1 );
not ( \3071_b1 , w_6888 );
and ( \3072_b0 , \3007_b0 , w_6889 );
and ( w_6888 , w_6889 , \3071_b0 );
or ( \3073_b1 , \3007_b1 , \3071_b1 );
xor ( \3073_b0 , \3007_b0 , w_6890 );
not ( w_6890 , w_6891 );
and ( w_6891 , \3071_b1 , \3071_b0 );
or ( \3074_b1 , \3063_b1 , \3065_b1 );
xor ( \3074_b0 , \3063_b0 , w_6892 );
not ( w_6892 , w_6893 );
and ( w_6893 , \3065_b1 , \3065_b0 );
or ( \3075_b1 , \3074_b1 , \3068_b1 );
xor ( \3075_b0 , \3074_b0 , w_6894 );
not ( w_6894 , w_6895 );
and ( w_6895 , \3068_b1 , \3068_b0 );
or ( \3076_b1 , \1477_b1 , \1336_b1 );
not ( \1336_b1 , w_6896 );
and ( \3076_b0 , \1477_b0 , w_6897 );
and ( w_6896 , w_6897 , \1336_b0 );
or ( \3077_b1 , \1454_b1 , \1333_b1 );
not ( \1333_b1 , w_6898 );
and ( \3077_b0 , \1454_b0 , w_6899 );
and ( w_6898 , w_6899 , \1333_b0 );
or ( \3078_b1 , \3076_b1 , w_6901 );
not ( w_6901 , w_6902 );
and ( \3078_b0 , \3076_b0 , w_6903 );
and ( w_6902 ,  , w_6903 );
buf ( w_6901 , \3077_b1 );
not ( w_6901 , w_6904 );
not (  , w_6905 );
and ( w_6904 , w_6905 , \3077_b0 );
or ( \3079_b1 , \3078_b1 , w_6906 );
xor ( \3079_b0 , \3078_b0 , w_6908 );
not ( w_6908 , w_6909 );
and ( w_6909 , w_6906 , w_6907 );
buf ( w_6906 , \1332_b1 );
not ( w_6906 , w_6910 );
not ( w_6907 , w_6911 );
and ( w_6910 , w_6911 , \1332_b0 );
or ( \3080_b1 , \1416_b1 , \1382_b1 );
not ( \1382_b1 , w_6912 );
and ( \3080_b0 , \1416_b0 , w_6913 );
and ( w_6912 , w_6913 , \1382_b0 );
or ( \3081_b1 , \1586_b1 , \1380_b1 );
not ( \1380_b1 , w_6914 );
and ( \3081_b0 , \1586_b0 , w_6915 );
and ( w_6914 , w_6915 , \1380_b0 );
or ( \3082_b1 , \3080_b1 , w_6917 );
not ( w_6917 , w_6918 );
and ( \3082_b0 , \3080_b0 , w_6919 );
and ( w_6918 ,  , w_6919 );
buf ( w_6917 , \3081_b1 );
not ( w_6917 , w_6920 );
not (  , w_6921 );
and ( w_6920 , w_6921 , \3081_b0 );
or ( \3083_b1 , \3082_b1 , w_6922 );
xor ( \3083_b0 , \3082_b0 , w_6924 );
not ( w_6924 , w_6925 );
and ( w_6925 , w_6922 , w_6923 );
buf ( w_6922 , \1389_b1 );
not ( w_6922 , w_6926 );
not ( w_6923 , w_6927 );
and ( w_6926 , w_6927 , \1389_b0 );
or ( \3084_b1 , \3079_b1 , \3083_b1 );
not ( \3083_b1 , w_6928 );
and ( \3084_b0 , \3079_b0 , w_6929 );
and ( w_6928 , w_6929 , \3083_b0 );
or ( \3085_b1 , \1498_b1 , \1397_b1 );
not ( \1397_b1 , w_6930 );
and ( \3085_b0 , \1498_b0 , w_6931 );
and ( w_6930 , w_6931 , \1397_b0 );
or ( \3086_b1 , \1553_b1 , \1395_b1 );
not ( \1395_b1 , w_6932 );
and ( \3086_b0 , \1553_b0 , w_6933 );
and ( w_6932 , w_6933 , \1395_b0 );
or ( \3087_b1 , \3085_b1 , w_6935 );
not ( w_6935 , w_6936 );
and ( \3087_b0 , \3085_b0 , w_6937 );
and ( w_6936 ,  , w_6937 );
buf ( w_6935 , \3086_b1 );
not ( w_6935 , w_6938 );
not (  , w_6939 );
and ( w_6938 , w_6939 , \3086_b0 );
or ( \3088_b1 , \3087_b1 , w_6940 );
xor ( \3088_b0 , \3087_b0 , w_6942 );
not ( w_6942 , w_6943 );
and ( w_6943 , w_6940 , w_6941 );
buf ( w_6940 , \1404_b1 );
not ( w_6940 , w_6944 );
not ( w_6941 , w_6945 );
and ( w_6944 , w_6945 , \1404_b0 );
or ( \3089_b1 , \3083_b1 , \3088_b1 );
not ( \3088_b1 , w_6946 );
and ( \3089_b0 , \3083_b0 , w_6947 );
and ( w_6946 , w_6947 , \3088_b0 );
or ( \3090_b1 , \3079_b1 , \3088_b1 );
not ( \3088_b1 , w_6948 );
and ( \3090_b0 , \3079_b0 , w_6949 );
and ( w_6948 , w_6949 , \3088_b0 );
or ( \3092_b1 , \1399_b1 , \1444_b1 );
not ( \1444_b1 , w_6950 );
and ( \3092_b0 , \1399_b0 , w_6951 );
and ( w_6950 , w_6951 , \1444_b0 );
or ( \3093_b1 , \1359_b1 , \1442_b1 );
not ( \1442_b1 , w_6952 );
and ( \3093_b0 , \1359_b0 , w_6953 );
and ( w_6952 , w_6953 , \1442_b0 );
or ( \3094_b1 , \3092_b1 , w_6955 );
not ( w_6955 , w_6956 );
and ( \3094_b0 , \3092_b0 , w_6957 );
and ( w_6956 ,  , w_6957 );
buf ( w_6955 , \3093_b1 );
not ( w_6955 , w_6958 );
not (  , w_6959 );
and ( w_6958 , w_6959 , \3093_b0 );
or ( \3095_b1 , \3094_b1 , w_6960 );
xor ( \3095_b0 , \3094_b0 , w_6962 );
not ( w_6962 , w_6963 );
and ( w_6963 , w_6960 , w_6961 );
buf ( w_6960 , \1451_b1 );
not ( w_6960 , w_6964 );
not ( w_6961 , w_6965 );
and ( w_6964 , w_6965 , \1451_b0 );
or ( \3096_b1 , \1616_b1 , \1349_b1 );
not ( \1349_b1 , w_6966 );
and ( \3096_b0 , \1616_b0 , w_6967 );
and ( w_6966 , w_6967 , \1349_b0 );
or ( \3097_b1 , \1391_b1 , \1347_b1 );
not ( \1347_b1 , w_6968 );
and ( \3097_b0 , \1391_b0 , w_6969 );
and ( w_6968 , w_6969 , \1347_b0 );
or ( \3098_b1 , \3096_b1 , w_6971 );
not ( w_6971 , w_6972 );
and ( \3098_b0 , \3096_b0 , w_6973 );
and ( w_6972 ,  , w_6973 );
buf ( w_6971 , \3097_b1 );
not ( w_6971 , w_6974 );
not (  , w_6975 );
and ( w_6974 , w_6975 , \3097_b0 );
or ( \3099_b1 , \3098_b1 , w_6976 );
xor ( \3099_b0 , \3098_b0 , w_6978 );
not ( w_6978 , w_6979 );
and ( w_6979 , w_6976 , w_6977 );
buf ( w_6976 , \1356_b1 );
not ( w_6976 , w_6980 );
not ( w_6977 , w_6981 );
and ( w_6980 , w_6981 , \1356_b0 );
or ( \3100_b1 , \3095_b1 , \3099_b1 );
not ( \3099_b1 , w_6982 );
and ( \3100_b0 , \3095_b0 , w_6983 );
and ( w_6982 , w_6983 , \3099_b0 );
or ( \3101_b1 , \1533_b1 , \1366_b1 );
not ( \1366_b1 , w_6984 );
and ( \3101_b0 , \1533_b0 , w_6985 );
and ( w_6984 , w_6985 , \1366_b0 );
or ( \3102_b1 , \1540_b1 , \1364_b1 );
not ( \1364_b1 , w_6986 );
and ( \3102_b0 , \1540_b0 , w_6987 );
and ( w_6986 , w_6987 , \1364_b0 );
or ( \3103_b1 , \3101_b1 , w_6989 );
not ( w_6989 , w_6990 );
and ( \3103_b0 , \3101_b0 , w_6991 );
and ( w_6990 ,  , w_6991 );
buf ( w_6989 , \3102_b1 );
not ( w_6989 , w_6992 );
not (  , w_6993 );
and ( w_6992 , w_6993 , \3102_b0 );
or ( \3104_b1 , \3103_b1 , w_6994 );
xor ( \3104_b0 , \3103_b0 , w_6996 );
not ( w_6996 , w_6997 );
and ( w_6997 , w_6994 , w_6995 );
buf ( w_6994 , \1373_b1 );
not ( w_6994 , w_6998 );
not ( w_6995 , w_6999 );
and ( w_6998 , w_6999 , \1373_b0 );
or ( \3105_b1 , \3099_b1 , \3104_b1 );
not ( \3104_b1 , w_7000 );
and ( \3105_b0 , \3099_b0 , w_7001 );
and ( w_7000 , w_7001 , \3104_b0 );
or ( \3106_b1 , \3095_b1 , \3104_b1 );
not ( \3104_b1 , w_7002 );
and ( \3106_b0 , \3095_b0 , w_7003 );
and ( w_7002 , w_7003 , \3104_b0 );
or ( \3108_b1 , \3091_b1 , \3107_b1 );
not ( \3107_b1 , w_7004 );
and ( \3108_b0 , \3091_b0 , w_7005 );
and ( w_7004 , w_7005 , \3107_b0 );
or ( \3109_b1 , \3035_b1 , \3038_b1 );
xor ( \3109_b0 , \3035_b0 , w_7006 );
not ( w_7006 , w_7007 );
and ( w_7007 , \3038_b1 , \3038_b0 );
or ( \3110_b1 , \1622_b1 , \1460_b1 );
not ( \1460_b1 , w_7008 );
and ( \3110_b0 , \1622_b0 , w_7009 );
and ( w_7008 , w_7009 , \1460_b0 );
or ( \3111_b1 , \1407_b1 , \1458_b1 );
not ( \1458_b1 , w_7010 );
and ( \3111_b0 , \1407_b0 , w_7011 );
and ( w_7010 , w_7011 , \1458_b0 );
or ( \3112_b1 , \3110_b1 , w_7013 );
not ( w_7013 , w_7014 );
and ( \3112_b0 , \3110_b0 , w_7015 );
and ( w_7014 ,  , w_7015 );
buf ( w_7013 , \3111_b1 );
not ( w_7013 , w_7016 );
not (  , w_7017 );
and ( w_7016 , w_7017 , \3111_b0 );
or ( \3113_b1 , \3112_b1 , w_7018 );
xor ( \3113_b0 , \3112_b0 , w_7020 );
not ( w_7020 , w_7021 );
and ( w_7021 , w_7018 , w_7019 );
buf ( w_7018 , \1467_b1 );
not ( w_7018 , w_7022 );
not ( w_7019 , w_7023 );
and ( w_7022 , w_7023 , \1467_b0 );
or ( \3114_b1 , \3109_b1 , \3113_b1 );
not ( \3113_b1 , w_7024 );
and ( \3114_b0 , \3109_b0 , w_7025 );
and ( w_7024 , w_7025 , \3113_b0 );
or ( \3115_b1 , \1517_b1 , \1475_b1 );
not ( \1475_b1 , w_7026 );
and ( \3115_b0 , \1517_b0 , w_7027 );
and ( w_7026 , w_7027 , \1475_b0 );
or ( \3116_b1 , \1526_b1 , \1473_b1 );
not ( \1473_b1 , w_7028 );
and ( \3116_b0 , \1526_b0 , w_7029 );
and ( w_7028 , w_7029 , \1473_b0 );
or ( \3117_b1 , \3115_b1 , w_7031 );
not ( w_7031 , w_7032 );
and ( \3117_b0 , \3115_b0 , w_7033 );
and ( w_7032 ,  , w_7033 );
buf ( w_7031 , \3116_b1 );
not ( w_7031 , w_7034 );
not (  , w_7035 );
and ( w_7034 , w_7035 , \3116_b0 );
or ( \3118_b1 , \3117_b1 , w_7036 );
xor ( \3118_b0 , \3117_b0 , w_7038 );
not ( w_7038 , w_7039 );
and ( w_7039 , w_7036 , w_7037 );
buf ( w_7036 , \1482_b1 );
not ( w_7036 , w_7040 );
not ( w_7037 , w_7041 );
and ( w_7040 , w_7041 , \1482_b0 );
or ( \3119_b1 , \3113_b1 , \3118_b1 );
not ( \3118_b1 , w_7042 );
and ( \3119_b0 , \3113_b0 , w_7043 );
and ( w_7042 , w_7043 , \3118_b0 );
or ( \3120_b1 , \3109_b1 , \3118_b1 );
not ( \3118_b1 , w_7044 );
and ( \3120_b0 , \3109_b0 , w_7045 );
and ( w_7044 , w_7045 , \3118_b0 );
or ( \3122_b1 , \3107_b1 , \3121_b1 );
not ( \3121_b1 , w_7046 );
and ( \3122_b0 , \3107_b0 , w_7047 );
and ( w_7046 , w_7047 , \3121_b0 );
or ( \3123_b1 , \3091_b1 , \3121_b1 );
not ( \3121_b1 , w_7048 );
and ( \3123_b0 , \3091_b0 , w_7049 );
and ( w_7048 , w_7049 , \3121_b0 );
or ( \3125_b1 , \1407_b1 , \1382_b1 );
not ( \1382_b1 , w_7050 );
and ( \3125_b0 , \1407_b0 , w_7051 );
and ( w_7050 , w_7051 , \1382_b0 );
or ( \3126_b1 , \1416_b1 , \1380_b1 );
not ( \1380_b1 , w_7052 );
and ( \3126_b0 , \1416_b0 , w_7053 );
and ( w_7052 , w_7053 , \1380_b0 );
or ( \3127_b1 , \3125_b1 , w_7055 );
not ( w_7055 , w_7056 );
and ( \3127_b0 , \3125_b0 , w_7057 );
and ( w_7056 ,  , w_7057 );
buf ( w_7055 , \3126_b1 );
not ( w_7055 , w_7058 );
not (  , w_7059 );
and ( w_7058 , w_7059 , \3126_b0 );
or ( \3128_b1 , \3127_b1 , w_7060 );
xor ( \3128_b0 , \3127_b0 , w_7062 );
not ( w_7062 , w_7063 );
and ( w_7063 , w_7060 , w_7061 );
buf ( w_7060 , \1389_b1 );
not ( w_7060 , w_7064 );
not ( w_7061 , w_7065 );
and ( w_7064 , w_7065 , \1389_b0 );
or ( \3129_b1 , \1526_b1 , \1460_b1 );
not ( \1460_b1 , w_7066 );
and ( \3129_b0 , \1526_b0 , w_7067 );
and ( w_7066 , w_7067 , \1460_b0 );
or ( \3130_b1 , \1622_b1 , \1458_b1 );
not ( \1458_b1 , w_7068 );
and ( \3130_b0 , \1622_b0 , w_7069 );
and ( w_7068 , w_7069 , \1458_b0 );
or ( \3131_b1 , \3129_b1 , w_7071 );
not ( w_7071 , w_7072 );
and ( \3131_b0 , \3129_b0 , w_7073 );
and ( w_7072 ,  , w_7073 );
buf ( w_7071 , \3130_b1 );
not ( w_7071 , w_7074 );
not (  , w_7075 );
and ( w_7074 , w_7075 , \3130_b0 );
or ( \3132_b1 , \3131_b1 , w_7076 );
xor ( \3132_b0 , \3131_b0 , w_7078 );
not ( w_7078 , w_7079 );
and ( w_7079 , w_7076 , w_7077 );
buf ( w_7076 , \1467_b1 );
not ( w_7076 , w_7080 );
not ( w_7077 , w_7081 );
and ( w_7080 , w_7081 , \1467_b0 );
or ( \3133_b1 , \3128_b1 , \3132_b1 );
not ( \3132_b1 , w_7082 );
and ( \3133_b0 , \3128_b0 , w_7083 );
and ( w_7082 , w_7083 , \3132_b0 );
or ( \3134_b1 , \1540_b1 , \1475_b1 );
not ( \1475_b1 , w_7084 );
and ( \3134_b0 , \1540_b0 , w_7085 );
and ( w_7084 , w_7085 , \1475_b0 );
or ( \3135_b1 , \1517_b1 , \1473_b1 );
not ( \1473_b1 , w_7086 );
and ( \3135_b0 , \1517_b0 , w_7087 );
and ( w_7086 , w_7087 , \1473_b0 );
or ( \3136_b1 , \3134_b1 , w_7089 );
not ( w_7089 , w_7090 );
and ( \3136_b0 , \3134_b0 , w_7091 );
and ( w_7090 ,  , w_7091 );
buf ( w_7089 , \3135_b1 );
not ( w_7089 , w_7092 );
not (  , w_7093 );
and ( w_7092 , w_7093 , \3135_b0 );
or ( \3137_b1 , \3136_b1 , w_7094 );
xor ( \3137_b0 , \3136_b0 , w_7096 );
not ( w_7096 , w_7097 );
and ( w_7097 , w_7094 , w_7095 );
buf ( w_7094 , \1482_b1 );
not ( w_7094 , w_7098 );
not ( w_7095 , w_7099 );
and ( w_7098 , w_7099 , \1482_b0 );
or ( \3138_b1 , \3132_b1 , \3137_b1 );
not ( \3137_b1 , w_7100 );
and ( \3138_b0 , \3132_b0 , w_7101 );
and ( w_7100 , w_7101 , \3137_b0 );
or ( \3139_b1 , \3128_b1 , \3137_b1 );
not ( \3137_b1 , w_7102 );
and ( \3139_b0 , \3128_b0 , w_7103 );
and ( w_7102 , w_7103 , \3137_b0 );
or ( \3141_b1 , \1470_b1 , \1336_b1 );
not ( \1336_b1 , w_7104 );
and ( \3141_b0 , \1470_b0 , w_7105 );
and ( w_7104 , w_7105 , \1336_b0 );
or ( \3142_b1 , \1477_b1 , \1333_b1 );
not ( \1333_b1 , w_7106 );
and ( \3142_b0 , \1477_b0 , w_7107 );
and ( w_7106 , w_7107 , \1333_b0 );
or ( \3143_b1 , \3141_b1 , w_7109 );
not ( w_7109 , w_7110 );
and ( \3143_b0 , \3141_b0 , w_7111 );
and ( w_7110 ,  , w_7111 );
buf ( w_7109 , \3142_b1 );
not ( w_7109 , w_7112 );
not (  , w_7113 );
and ( w_7112 , w_7113 , \3142_b0 );
or ( \3144_b1 , \3143_b1 , w_7114 );
xor ( \3144_b0 , \3143_b0 , w_7116 );
not ( w_7116 , w_7117 );
and ( w_7117 , w_7114 , w_7115 );
buf ( w_7114 , \1332_b1 );
not ( w_7114 , w_7118 );
not ( w_7115 , w_7119 );
and ( w_7118 , w_7119 , \1332_b0 );
or ( \3145_b1 , \1586_b1 , \1349_b1 );
not ( \1349_b1 , w_7120 );
and ( \3145_b0 , \1586_b0 , w_7121 );
and ( w_7120 , w_7121 , \1349_b0 );
or ( \3146_b1 , \1616_b1 , \1347_b1 );
not ( \1347_b1 , w_7122 );
and ( \3146_b0 , \1616_b0 , w_7123 );
and ( w_7122 , w_7123 , \1347_b0 );
or ( \3147_b1 , \3145_b1 , w_7125 );
not ( w_7125 , w_7126 );
and ( \3147_b0 , \3145_b0 , w_7127 );
and ( w_7126 ,  , w_7127 );
buf ( w_7125 , \3146_b1 );
not ( w_7125 , w_7128 );
not (  , w_7129 );
and ( w_7128 , w_7129 , \3146_b0 );
or ( \3148_b1 , \3147_b1 , w_7130 );
xor ( \3148_b0 , \3147_b0 , w_7132 );
not ( w_7132 , w_7133 );
and ( w_7133 , w_7130 , w_7131 );
buf ( w_7130 , \1356_b1 );
not ( w_7130 , w_7134 );
not ( w_7131 , w_7135 );
and ( w_7134 , w_7135 , \1356_b0 );
or ( \3149_b1 , \3144_b1 , \3148_b1 );
not ( \3148_b1 , w_7136 );
and ( \3149_b0 , \3144_b0 , w_7137 );
and ( w_7136 , w_7137 , \3148_b0 );
or ( \3150_b1 , \1553_b1 , \1366_b1 );
not ( \1366_b1 , w_7138 );
and ( \3150_b0 , \1553_b0 , w_7139 );
and ( w_7138 , w_7139 , \1366_b0 );
or ( \3151_b1 , \1533_b1 , \1364_b1 );
not ( \1364_b1 , w_7140 );
and ( \3151_b0 , \1533_b0 , w_7141 );
and ( w_7140 , w_7141 , \1364_b0 );
or ( \3152_b1 , \3150_b1 , w_7143 );
not ( w_7143 , w_7144 );
and ( \3152_b0 , \3150_b0 , w_7145 );
and ( w_7144 ,  , w_7145 );
buf ( w_7143 , \3151_b1 );
not ( w_7143 , w_7146 );
not (  , w_7147 );
and ( w_7146 , w_7147 , \3151_b0 );
or ( \3153_b1 , \3152_b1 , w_7148 );
xor ( \3153_b0 , \3152_b0 , w_7150 );
not ( w_7150 , w_7151 );
and ( w_7151 , w_7148 , w_7149 );
buf ( w_7148 , \1373_b1 );
not ( w_7148 , w_7152 );
not ( w_7149 , w_7153 );
and ( w_7152 , w_7153 , \1373_b0 );
or ( \3154_b1 , \3148_b1 , \3153_b1 );
not ( \3153_b1 , w_7154 );
and ( \3154_b0 , \3148_b0 , w_7155 );
and ( w_7154 , w_7155 , \3153_b0 );
or ( \3155_b1 , \3144_b1 , \3153_b1 );
not ( \3153_b1 , w_7156 );
and ( \3155_b0 , \3144_b0 , w_7157 );
and ( w_7156 , w_7157 , \3153_b0 );
or ( \3157_b1 , \3140_b1 , \3156_b1 );
not ( \3156_b1 , w_7158 );
and ( \3157_b0 , \3140_b0 , w_7159 );
and ( w_7158 , w_7159 , \3156_b0 );
or ( \3158_b1 , \1359_b1 , \1431_b1 );
not ( \1431_b1 , w_7160 );
and ( \3158_b0 , \1359_b0 , w_7161 );
and ( w_7160 , w_7161 , \1431_b0 );
or ( \3159_b1 , \1368_b1 , \1429_b1 );
not ( \1429_b1 , w_7162 );
and ( \3159_b0 , \1368_b0 , w_7163 );
and ( w_7162 , w_7163 , \1429_b0 );
or ( \3160_b1 , \3158_b1 , w_7165 );
not ( w_7165 , w_7166 );
and ( \3160_b0 , \3158_b0 , w_7167 );
and ( w_7166 ,  , w_7167 );
buf ( w_7165 , \3159_b1 );
not ( w_7165 , w_7168 );
not (  , w_7169 );
and ( w_7168 , w_7169 , \3159_b0 );
or ( \3161_b1 , \3160_b1 , w_7170 );
xor ( \3161_b0 , \3160_b0 , w_7172 );
not ( w_7172 , w_7173 );
and ( w_7173 , w_7170 , w_7171 );
buf ( w_7170 , \1438_b1 );
not ( w_7170 , w_7174 );
not ( w_7171 , w_7175 );
and ( w_7174 , w_7175 , \1438_b0 );
or ( \3162_b1 , \1391_b1 , \1444_b1 );
not ( \1444_b1 , w_7176 );
and ( \3162_b0 , \1391_b0 , w_7177 );
and ( w_7176 , w_7177 , \1444_b0 );
or ( \3163_b1 , \1399_b1 , \1442_b1 );
not ( \1442_b1 , w_7178 );
and ( \3163_b0 , \1399_b0 , w_7179 );
and ( w_7178 , w_7179 , \1442_b0 );
or ( \3164_b1 , \3162_b1 , w_7181 );
not ( w_7181 , w_7182 );
and ( \3164_b0 , \3162_b0 , w_7183 );
and ( w_7182 ,  , w_7183 );
buf ( w_7181 , \3163_b1 );
not ( w_7181 , w_7184 );
not (  , w_7185 );
and ( w_7184 , w_7185 , \3163_b0 );
or ( \3165_b1 , \3164_b1 , w_7186 );
xor ( \3165_b0 , \3164_b0 , w_7188 );
not ( w_7188 , w_7189 );
and ( w_7189 , w_7186 , w_7187 );
buf ( w_7186 , \1451_b1 );
not ( w_7186 , w_7190 );
not ( w_7187 , w_7191 );
and ( w_7190 , w_7191 , \1451_b0 );
or ( \3166_b1 , \3161_b1 , \3165_b1 );
not ( \3165_b1 , w_7192 );
and ( \3166_b0 , \3161_b0 , w_7193 );
and ( w_7192 , w_7193 , \3165_b0 );
or ( \3167_b1 , \3165_b1 , \3036_b1 );
not ( \3036_b1 , w_7194 );
and ( \3167_b0 , \3165_b0 , w_7195 );
and ( w_7194 , w_7195 , \3036_b0 );
or ( \3168_b1 , \3161_b1 , \3036_b1 );
not ( \3036_b1 , w_7196 );
and ( \3168_b0 , \3161_b0 , w_7197 );
and ( w_7196 , w_7197 , \3036_b0 );
or ( \3170_b1 , \3156_b1 , \3169_b1 );
not ( \3169_b1 , w_7198 );
and ( \3170_b0 , \3156_b0 , w_7199 );
and ( w_7198 , w_7199 , \3169_b0 );
or ( \3171_b1 , \3140_b1 , \3169_b1 );
not ( \3169_b1 , w_7200 );
and ( \3171_b0 , \3140_b0 , w_7201 );
and ( w_7200 , w_7201 , \3169_b0 );
or ( \3173_b1 , \3011_b1 , \3015_b1 );
xor ( \3173_b0 , \3011_b0 , w_7202 );
not ( w_7202 , w_7203 );
and ( w_7203 , \3015_b1 , \3015_b0 );
or ( \3174_b1 , \3173_b1 , \3020_b1 );
xor ( \3174_b0 , \3173_b0 , w_7204 );
not ( w_7204 , w_7205 );
and ( w_7205 , \3020_b1 , \3020_b0 );
or ( \3175_b1 , \3172_b1 , \3174_b1 );
not ( \3174_b1 , w_7206 );
and ( \3175_b0 , \3172_b0 , w_7207 );
and ( w_7206 , w_7207 , \3174_b0 );
or ( \3176_b1 , \2959_b1 , \2963_b1 );
xor ( \3176_b0 , \2959_b0 , w_7208 );
not ( w_7208 , w_7209 );
and ( w_7209 , \2963_b1 , \2963_b0 );
or ( \3177_b1 , \3176_b1 , \2968_b1 );
xor ( \3177_b0 , \3176_b0 , w_7210 );
not ( w_7210 , w_7211 );
and ( w_7211 , \2968_b1 , \2968_b0 );
or ( \3178_b1 , \3174_b1 , \3177_b1 );
not ( \3177_b1 , w_7212 );
and ( \3178_b0 , \3174_b0 , w_7213 );
and ( w_7212 , w_7213 , \3177_b0 );
or ( \3179_b1 , \3172_b1 , \3177_b1 );
not ( \3177_b1 , w_7214 );
and ( \3179_b0 , \3172_b0 , w_7215 );
and ( w_7214 , w_7215 , \3177_b0 );
or ( \3181_b1 , \3124_b1 , \3180_b1 );
not ( \3180_b1 , w_7216 );
and ( \3181_b0 , \3124_b0 , w_7217 );
and ( w_7216 , w_7217 , \3180_b0 );
or ( \3182_b1 , \3023_b1 , \3025_b1 );
xor ( \3182_b0 , \3023_b0 , w_7218 );
not ( w_7218 , w_7219 );
and ( w_7219 , \3025_b1 , \3025_b0 );
or ( \3183_b1 , \3182_b1 , \3028_b1 );
xor ( \3183_b0 , \3182_b0 , w_7220 );
not ( w_7220 , w_7221 );
and ( w_7221 , \3028_b1 , \3028_b0 );
or ( \3184_b1 , \3180_b1 , \3183_b1 );
not ( \3183_b1 , w_7222 );
and ( \3184_b0 , \3180_b0 , w_7223 );
and ( w_7222 , w_7223 , \3183_b0 );
or ( \3185_b1 , \3124_b1 , \3183_b1 );
not ( \3183_b1 , w_7224 );
and ( \3185_b0 , \3124_b0 , w_7225 );
and ( w_7224 , w_7225 , \3183_b0 );
or ( \3187_b1 , \2979_b1 , \2981_b1 );
xor ( \3187_b0 , \2979_b0 , w_7226 );
not ( w_7226 , w_7227 );
and ( w_7227 , \2981_b1 , \2981_b0 );
or ( \3188_b1 , \3187_b1 , \2984_b1 );
xor ( \3188_b0 , \3187_b0 , w_7228 );
not ( w_7228 , w_7229 );
and ( w_7229 , \2984_b1 , \2984_b0 );
or ( \3189_b1 , \3186_b1 , \3188_b1 );
not ( \3188_b1 , w_7230 );
and ( \3189_b0 , \3186_b0 , w_7231 );
and ( w_7230 , w_7231 , \3188_b0 );
or ( \3190_b1 , \3031_b1 , \3057_b1 );
xor ( \3190_b0 , \3031_b0 , w_7232 );
not ( w_7232 , w_7233 );
and ( w_7233 , \3057_b1 , \3057_b0 );
or ( \3191_b1 , \3190_b1 , \3060_b1 );
xor ( \3191_b0 , \3190_b0 , w_7234 );
not ( w_7234 , w_7235 );
and ( w_7235 , \3060_b1 , \3060_b0 );
or ( \3192_b1 , \3188_b1 , \3191_b1 );
not ( \3191_b1 , w_7236 );
and ( \3192_b0 , \3188_b0 , w_7237 );
and ( w_7236 , w_7237 , \3191_b0 );
or ( \3193_b1 , \3186_b1 , \3191_b1 );
not ( \3191_b1 , w_7238 );
and ( \3193_b0 , \3186_b0 , w_7239 );
and ( w_7238 , w_7239 , \3191_b0 );
or ( \3195_b1 , \3075_b1 , \3194_b1 );
not ( \3194_b1 , w_7240 );
and ( \3195_b0 , \3075_b0 , w_7241 );
and ( w_7240 , w_7241 , \3194_b0 );
or ( \3196_b1 , \3075_b1 , \3194_b1 );
xor ( \3196_b0 , \3075_b0 , w_7242 );
not ( w_7242 , w_7243 );
and ( w_7243 , \3194_b1 , \3194_b0 );
or ( \3197_b1 , \3186_b1 , \3188_b1 );
xor ( \3197_b0 , \3186_b0 , w_7244 );
not ( w_7244 , w_7245 );
and ( w_7245 , \3188_b1 , \3188_b0 );
or ( \3198_b1 , \3197_b1 , \3191_b1 );
xor ( \3198_b0 , \3197_b0 , w_7246 );
not ( w_7246 , w_7247 );
and ( w_7247 , \3191_b1 , \3191_b0 );
or ( \3199_b1 , \3079_b1 , \3083_b1 );
xor ( \3199_b0 , \3079_b0 , w_7248 );
not ( w_7248 , w_7249 );
and ( w_7249 , \3083_b1 , \3083_b0 );
or ( \3200_b1 , \3199_b1 , \3088_b1 );
xor ( \3200_b0 , \3199_b0 , w_7250 );
not ( w_7250 , w_7251 );
and ( w_7251 , \3088_b1 , \3088_b0 );
or ( \3201_b1 , \3095_b1 , \3099_b1 );
xor ( \3201_b0 , \3095_b0 , w_7252 );
not ( w_7252 , w_7253 );
and ( w_7253 , \3099_b1 , \3099_b0 );
or ( \3202_b1 , \3201_b1 , \3104_b1 );
xor ( \3202_b0 , \3201_b0 , w_7254 );
not ( w_7254 , w_7255 );
and ( w_7255 , \3104_b1 , \3104_b0 );
or ( \3203_b1 , \3200_b1 , \3202_b1 );
not ( \3202_b1 , w_7256 );
and ( \3203_b0 , \3200_b0 , w_7257 );
and ( w_7256 , w_7257 , \3202_b0 );
or ( \3204_b1 , \3109_b1 , \3113_b1 );
xor ( \3204_b0 , \3109_b0 , w_7258 );
not ( w_7258 , w_7259 );
and ( w_7259 , \3113_b1 , \3113_b0 );
or ( \3205_b1 , \3204_b1 , \3118_b1 );
xor ( \3205_b0 , \3204_b0 , w_7260 );
not ( w_7260 , w_7261 );
and ( w_7261 , \3118_b1 , \3118_b0 );
or ( \3206_b1 , \3202_b1 , \3205_b1 );
not ( \3205_b1 , w_7262 );
and ( \3206_b0 , \3202_b0 , w_7263 );
and ( w_7262 , w_7263 , \3205_b0 );
or ( \3207_b1 , \3200_b1 , \3205_b1 );
not ( \3205_b1 , w_7264 );
and ( \3207_b0 , \3200_b0 , w_7265 );
and ( w_7264 , w_7265 , \3205_b0 );
or ( \3209_b1 , \3091_b1 , \3107_b1 );
xor ( \3209_b0 , \3091_b0 , w_7266 );
not ( w_7266 , w_7267 );
and ( w_7267 , \3107_b1 , \3107_b0 );
or ( \3210_b1 , \3209_b1 , \3121_b1 );
xor ( \3210_b0 , \3209_b0 , w_7268 );
not ( w_7268 , w_7269 );
and ( w_7269 , \3121_b1 , \3121_b0 );
or ( \3211_b1 , \3208_b1 , \3210_b1 );
not ( \3210_b1 , w_7270 );
and ( \3211_b0 , \3208_b0 , w_7271 );
and ( w_7270 , w_7271 , \3210_b0 );
or ( \3212_b1 , \3039_b1 , \3043_b1 );
xor ( \3212_b0 , \3039_b0 , w_7272 );
not ( w_7272 , w_7273 );
and ( w_7273 , \3043_b1 , \3043_b0 );
or ( \3213_b1 , \3212_b1 , \3046_b1 );
xor ( \3213_b0 , \3212_b0 , w_7274 );
not ( w_7274 , w_7275 );
and ( w_7275 , \3046_b1 , \3046_b0 );
or ( \3214_b1 , \3210_b1 , \3213_b1 );
not ( \3213_b1 , w_7276 );
and ( \3214_b0 , \3210_b0 , w_7277 );
and ( w_7276 , w_7277 , \3213_b0 );
or ( \3215_b1 , \3208_b1 , \3213_b1 );
not ( \3213_b1 , w_7278 );
and ( \3215_b0 , \3208_b0 , w_7279 );
and ( w_7278 , w_7279 , \3213_b0 );
or ( \3217_b1 , \3049_b1 , \3051_b1 );
xor ( \3217_b0 , \3049_b0 , w_7280 );
not ( w_7280 , w_7281 );
and ( w_7281 , \3051_b1 , \3051_b0 );
or ( \3218_b1 , \3217_b1 , \3054_b1 );
xor ( \3218_b0 , \3217_b0 , w_7282 );
not ( w_7282 , w_7283 );
and ( w_7283 , \3054_b1 , \3054_b0 );
or ( \3219_b1 , \3216_b1 , \3218_b1 );
not ( \3218_b1 , w_7284 );
and ( \3219_b0 , \3216_b0 , w_7285 );
and ( w_7284 , w_7285 , \3218_b0 );
or ( \3220_b1 , \3124_b1 , \3180_b1 );
xor ( \3220_b0 , \3124_b0 , w_7286 );
not ( w_7286 , w_7287 );
and ( w_7287 , \3180_b1 , \3180_b0 );
or ( \3221_b1 , \3220_b1 , \3183_b1 );
xor ( \3221_b0 , \3220_b0 , w_7288 );
not ( w_7288 , w_7289 );
and ( w_7289 , \3183_b1 , \3183_b0 );
or ( \3222_b1 , \3218_b1 , \3221_b1 );
not ( \3221_b1 , w_7290 );
and ( \3222_b0 , \3218_b0 , w_7291 );
and ( w_7290 , w_7291 , \3221_b0 );
or ( \3223_b1 , \3216_b1 , \3221_b1 );
not ( \3221_b1 , w_7292 );
and ( \3223_b0 , \3216_b0 , w_7293 );
and ( w_7292 , w_7293 , \3221_b0 );
or ( \3225_b1 , \3198_b1 , \3224_b1 );
not ( \3224_b1 , w_7294 );
and ( \3225_b0 , \3198_b0 , w_7295 );
and ( w_7294 , w_7295 , \3224_b0 );
or ( \3226_b1 , \3198_b1 , \3224_b1 );
xor ( \3226_b0 , \3198_b0 , w_7296 );
not ( w_7296 , w_7297 );
and ( w_7297 , \3224_b1 , \3224_b0 );
or ( \3227_b1 , \3216_b1 , \3218_b1 );
xor ( \3227_b0 , \3216_b0 , w_7298 );
not ( w_7298 , w_7299 );
and ( w_7299 , \3218_b1 , \3218_b0 );
or ( \3228_b1 , \3227_b1 , \3221_b1 );
xor ( \3228_b0 , \3227_b0 , w_7300 );
not ( w_7300 , w_7301 );
and ( w_7301 , \3221_b1 , \3221_b0 );
or ( \3229_b1 , \1416_b1 , \1349_b1 );
not ( \1349_b1 , w_7302 );
and ( \3229_b0 , \1416_b0 , w_7303 );
and ( w_7302 , w_7303 , \1349_b0 );
or ( \3230_b1 , \1586_b1 , \1347_b1 );
not ( \1347_b1 , w_7304 );
and ( \3230_b0 , \1586_b0 , w_7305 );
and ( w_7304 , w_7305 , \1347_b0 );
or ( \3231_b1 , \3229_b1 , w_7307 );
not ( w_7307 , w_7308 );
and ( \3231_b0 , \3229_b0 , w_7309 );
and ( w_7308 ,  , w_7309 );
buf ( w_7307 , \3230_b1 );
not ( w_7307 , w_7310 );
not (  , w_7311 );
and ( w_7310 , w_7311 , \3230_b0 );
or ( \3232_b1 , \3231_b1 , w_7312 );
xor ( \3232_b0 , \3231_b0 , w_7314 );
not ( w_7314 , w_7315 );
and ( w_7315 , w_7312 , w_7313 );
buf ( w_7312 , \1356_b1 );
not ( w_7312 , w_7316 );
not ( w_7313 , w_7317 );
and ( w_7316 , w_7317 , \1356_b0 );
or ( \3233_b1 , \1622_b1 , \1382_b1 );
not ( \1382_b1 , w_7318 );
and ( \3233_b0 , \1622_b0 , w_7319 );
and ( w_7318 , w_7319 , \1382_b0 );
or ( \3234_b1 , \1407_b1 , \1380_b1 );
not ( \1380_b1 , w_7320 );
and ( \3234_b0 , \1407_b0 , w_7321 );
and ( w_7320 , w_7321 , \1380_b0 );
or ( \3235_b1 , \3233_b1 , w_7323 );
not ( w_7323 , w_7324 );
and ( \3235_b0 , \3233_b0 , w_7325 );
and ( w_7324 ,  , w_7325 );
buf ( w_7323 , \3234_b1 );
not ( w_7323 , w_7326 );
not (  , w_7327 );
and ( w_7326 , w_7327 , \3234_b0 );
or ( \3236_b1 , \3235_b1 , w_7328 );
xor ( \3236_b0 , \3235_b0 , w_7330 );
not ( w_7330 , w_7331 );
and ( w_7331 , w_7328 , w_7329 );
buf ( w_7328 , \1389_b1 );
not ( w_7328 , w_7332 );
not ( w_7329 , w_7333 );
and ( w_7332 , w_7333 , \1389_b0 );
or ( \3237_b1 , \3232_b1 , \3236_b1 );
not ( \3236_b1 , w_7334 );
and ( \3237_b0 , \3232_b0 , w_7335 );
and ( w_7334 , w_7335 , \3236_b0 );
or ( \3238_b1 , \1517_b1 , \1460_b1 );
not ( \1460_b1 , w_7336 );
and ( \3238_b0 , \1517_b0 , w_7337 );
and ( w_7336 , w_7337 , \1460_b0 );
or ( \3239_b1 , \1526_b1 , \1458_b1 );
not ( \1458_b1 , w_7338 );
and ( \3239_b0 , \1526_b0 , w_7339 );
and ( w_7338 , w_7339 , \1458_b0 );
or ( \3240_b1 , \3238_b1 , w_7341 );
not ( w_7341 , w_7342 );
and ( \3240_b0 , \3238_b0 , w_7343 );
and ( w_7342 ,  , w_7343 );
buf ( w_7341 , \3239_b1 );
not ( w_7341 , w_7344 );
not (  , w_7345 );
and ( w_7344 , w_7345 , \3239_b0 );
or ( \3241_b1 , \3240_b1 , w_7346 );
xor ( \3241_b0 , \3240_b0 , w_7348 );
not ( w_7348 , w_7349 );
and ( w_7349 , w_7346 , w_7347 );
buf ( w_7346 , \1467_b1 );
not ( w_7346 , w_7350 );
not ( w_7347 , w_7351 );
and ( w_7350 , w_7351 , \1467_b0 );
or ( \3242_b1 , \3236_b1 , \3241_b1 );
not ( \3241_b1 , w_7352 );
and ( \3242_b0 , \3236_b0 , w_7353 );
and ( w_7352 , w_7353 , \3241_b0 );
or ( \3243_b1 , \3232_b1 , \3241_b1 );
not ( \3241_b1 , w_7354 );
and ( \3243_b0 , \3232_b0 , w_7355 );
and ( w_7354 , w_7355 , \3241_b0 );
or ( \3245_b1 , \3128_b1 , \3132_b1 );
xor ( \3245_b0 , \3128_b0 , w_7356 );
not ( w_7356 , w_7357 );
and ( w_7357 , \3132_b1 , \3132_b0 );
or ( \3246_b1 , \3245_b1 , \3137_b1 );
xor ( \3246_b0 , \3245_b0 , w_7358 );
not ( w_7358 , w_7359 );
and ( w_7359 , \3137_b1 , \3137_b0 );
or ( \3247_b1 , \3244_b1 , \3246_b1 );
not ( \3246_b1 , w_7360 );
and ( \3247_b0 , \3244_b0 , w_7361 );
and ( w_7360 , w_7361 , \3246_b0 );
or ( \3248_b1 , \3144_b1 , \3148_b1 );
xor ( \3248_b0 , \3144_b0 , w_7362 );
not ( w_7362 , w_7363 );
and ( w_7363 , \3148_b1 , \3148_b0 );
or ( \3249_b1 , \3248_b1 , \3153_b1 );
xor ( \3249_b0 , \3248_b0 , w_7364 );
not ( w_7364 , w_7365 );
and ( w_7365 , \3153_b1 , \3153_b0 );
or ( \3250_b1 , \3246_b1 , \3249_b1 );
not ( \3249_b1 , w_7366 );
and ( \3250_b0 , \3246_b0 , w_7367 );
and ( w_7366 , w_7367 , \3249_b0 );
or ( \3251_b1 , \3244_b1 , \3249_b1 );
not ( \3249_b1 , w_7368 );
and ( \3251_b0 , \3244_b0 , w_7369 );
and ( w_7368 , w_7369 , \3249_b0 );
or ( \3253_b1 , \1368_b1 , \1336_b1 );
not ( \1336_b1 , w_7370 );
and ( \3253_b0 , \1368_b0 , w_7371 );
and ( w_7370 , w_7371 , \1336_b0 );
or ( \3254_b1 , \1470_b1 , \1333_b1 );
not ( \1333_b1 , w_7372 );
and ( \3254_b0 , \1470_b0 , w_7373 );
and ( w_7372 , w_7373 , \1333_b0 );
or ( \3255_b1 , \3253_b1 , w_7375 );
not ( w_7375 , w_7376 );
and ( \3255_b0 , \3253_b0 , w_7377 );
and ( w_7376 ,  , w_7377 );
buf ( w_7375 , \3254_b1 );
not ( w_7375 , w_7378 );
not (  , w_7379 );
and ( w_7378 , w_7379 , \3254_b0 );
or ( \3256_b1 , \3255_b1 , w_7380 );
xor ( \3256_b0 , \3255_b0 , w_7382 );
not ( w_7382 , w_7383 );
and ( w_7383 , w_7380 , w_7381 );
buf ( w_7380 , \1332_b1 );
not ( w_7380 , w_7384 );
not ( w_7381 , w_7385 );
and ( w_7384 , w_7385 , \1332_b0 );
or ( \3257_b1 , \1616_b1 , \1444_b1 );
not ( \1444_b1 , w_7386 );
and ( \3257_b0 , \1616_b0 , w_7387 );
and ( w_7386 , w_7387 , \1444_b0 );
or ( \3258_b1 , \1391_b1 , \1442_b1 );
not ( \1442_b1 , w_7388 );
and ( \3258_b0 , \1391_b0 , w_7389 );
and ( w_7388 , w_7389 , \1442_b0 );
or ( \3259_b1 , \3257_b1 , w_7391 );
not ( w_7391 , w_7392 );
and ( \3259_b0 , \3257_b0 , w_7393 );
and ( w_7392 ,  , w_7393 );
buf ( w_7391 , \3258_b1 );
not ( w_7391 , w_7394 );
not (  , w_7395 );
and ( w_7394 , w_7395 , \3258_b0 );
or ( \3260_b1 , \3259_b1 , w_7396 );
xor ( \3260_b0 , \3259_b0 , w_7398 );
not ( w_7398 , w_7399 );
and ( w_7399 , w_7396 , w_7397 );
buf ( w_7396 , \1451_b1 );
not ( w_7396 , w_7400 );
not ( w_7397 , w_7401 );
and ( w_7400 , w_7401 , \1451_b0 );
or ( \3261_b1 , \3256_b1 , \3260_b1 );
not ( \3260_b1 , w_7402 );
and ( \3261_b0 , \3256_b0 , w_7403 );
and ( w_7402 , w_7403 , \3260_b0 );
or ( \3262_b1 , \1498_b1 , \1366_b1 );
not ( \1366_b1 , w_7404 );
and ( \3262_b0 , \1498_b0 , w_7405 );
and ( w_7404 , w_7405 , \1366_b0 );
or ( \3263_b1 , \1553_b1 , \1364_b1 );
not ( \1364_b1 , w_7406 );
and ( \3263_b0 , \1553_b0 , w_7407 );
and ( w_7406 , w_7407 , \1364_b0 );
or ( \3264_b1 , \3262_b1 , w_7409 );
not ( w_7409 , w_7410 );
and ( \3264_b0 , \3262_b0 , w_7411 );
and ( w_7410 ,  , w_7411 );
buf ( w_7409 , \3263_b1 );
not ( w_7409 , w_7412 );
not (  , w_7413 );
and ( w_7412 , w_7413 , \3263_b0 );
or ( \3265_b1 , \3264_b1 , w_7414 );
xor ( \3265_b0 , \3264_b0 , w_7416 );
not ( w_7416 , w_7417 );
and ( w_7417 , w_7414 , w_7415 );
buf ( w_7414 , \1373_b1 );
not ( w_7414 , w_7418 );
not ( w_7415 , w_7419 );
and ( w_7418 , w_7419 , \1373_b0 );
or ( \3266_b1 , \3260_b1 , \3265_b1 );
not ( \3265_b1 , w_7420 );
and ( \3266_b0 , \3260_b0 , w_7421 );
and ( w_7420 , w_7421 , \3265_b0 );
or ( \3267_b1 , \3256_b1 , \3265_b1 );
not ( \3265_b1 , w_7422 );
and ( \3267_b0 , \3256_b0 , w_7423 );
and ( w_7422 , w_7423 , \3265_b0 );
or ( \3269_b1 , \1399_b1 , \1431_b1 );
not ( \1431_b1 , w_7424 );
and ( \3269_b0 , \1399_b0 , w_7425 );
and ( w_7424 , w_7425 , \1431_b0 );
or ( \3270_b1 , \1359_b1 , \1429_b1 );
not ( \1429_b1 , w_7426 );
and ( \3270_b0 , \1359_b0 , w_7427 );
and ( w_7426 , w_7427 , \1429_b0 );
or ( \3271_b1 , \3269_b1 , w_7429 );
not ( w_7429 , w_7430 );
and ( \3271_b0 , \3269_b0 , w_7431 );
and ( w_7430 ,  , w_7431 );
buf ( w_7429 , \3270_b1 );
not ( w_7429 , w_7432 );
not (  , w_7433 );
and ( w_7432 , w_7433 , \3270_b0 );
or ( \3272_b1 , \3271_b1 , w_7434 );
xor ( \3272_b0 , \3271_b0 , w_7436 );
not ( w_7436 , w_7437 );
and ( w_7437 , w_7434 , w_7435 );
buf ( w_7434 , \1438_b1 );
not ( w_7434 , w_7438 );
not ( w_7435 , w_7439 );
and ( w_7438 , w_7439 , \1438_b0 );
or ( \3273_b1 , \1498_b1 , \1364_b1 );
not ( \1364_b1 , w_7440 );
and ( \3273_b0 , \1498_b0 , w_7441 );
and ( w_7440 , w_7441 , \1364_b0 );
buf ( \3274_b1 , \3273_b1 );
not ( \3274_b1 , w_7442 );
not ( \3274_b0 , w_7443 );
and ( w_7442 , w_7443 , \3273_b0 );
or ( \3275_b1 , \3274_b1 , \1373_b1 );
not ( \1373_b1 , w_7444 );
and ( \3275_b0 , \3274_b0 , w_7445 );
and ( w_7444 , w_7445 , \1373_b0 );
or ( \3276_b1 , \3272_b1 , \3275_b1 );
not ( \3275_b1 , w_7446 );
and ( \3276_b0 , \3272_b0 , w_7447 );
and ( w_7446 , w_7447 , \3275_b0 );
or ( \3277_b1 , \3268_b1 , \3276_b1 );
not ( \3276_b1 , w_7448 );
and ( \3277_b0 , \3268_b0 , w_7449 );
and ( w_7448 , w_7449 , \3276_b0 );
or ( \3278_b1 , \3161_b1 , \3165_b1 );
xor ( \3278_b0 , \3161_b0 , w_7450 );
not ( w_7450 , w_7451 );
and ( w_7451 , \3165_b1 , \3165_b0 );
or ( \3279_b1 , \3278_b1 , \3036_b1 );
xor ( \3279_b0 , \3278_b0 , w_7452 );
not ( w_7452 , w_7453 );
and ( w_7453 , \3036_b1 , \3036_b0 );
or ( \3280_b1 , \3276_b1 , \3279_b1 );
not ( \3279_b1 , w_7454 );
and ( \3280_b0 , \3276_b0 , w_7455 );
and ( w_7454 , w_7455 , \3279_b0 );
or ( \3281_b1 , \3268_b1 , \3279_b1 );
not ( \3279_b1 , w_7456 );
and ( \3281_b0 , \3268_b0 , w_7457 );
and ( w_7456 , w_7457 , \3279_b0 );
or ( \3283_b1 , \3252_b1 , \3282_b1 );
not ( \3282_b1 , w_7458 );
and ( \3283_b0 , \3252_b0 , w_7459 );
and ( w_7458 , w_7459 , \3282_b0 );
or ( \3284_b1 , \3140_b1 , \3156_b1 );
xor ( \3284_b0 , \3140_b0 , w_7460 );
not ( w_7460 , w_7461 );
and ( w_7461 , \3156_b1 , \3156_b0 );
or ( \3285_b1 , \3284_b1 , \3169_b1 );
xor ( \3285_b0 , \3284_b0 , w_7462 );
not ( w_7462 , w_7463 );
and ( w_7463 , \3169_b1 , \3169_b0 );
or ( \3286_b1 , \3282_b1 , \3285_b1 );
not ( \3285_b1 , w_7464 );
and ( \3286_b0 , \3282_b0 , w_7465 );
and ( w_7464 , w_7465 , \3285_b0 );
or ( \3287_b1 , \3252_b1 , \3285_b1 );
not ( \3285_b1 , w_7466 );
and ( \3287_b0 , \3252_b0 , w_7467 );
and ( w_7466 , w_7467 , \3285_b0 );
or ( \3289_b1 , \3172_b1 , \3174_b1 );
xor ( \3289_b0 , \3172_b0 , w_7468 );
not ( w_7468 , w_7469 );
and ( w_7469 , \3174_b1 , \3174_b0 );
or ( \3290_b1 , \3289_b1 , \3177_b1 );
xor ( \3290_b0 , \3289_b0 , w_7470 );
not ( w_7470 , w_7471 );
and ( w_7471 , \3177_b1 , \3177_b0 );
or ( \3291_b1 , \3288_b1 , \3290_b1 );
not ( \3290_b1 , w_7472 );
and ( \3291_b0 , \3288_b0 , w_7473 );
and ( w_7472 , w_7473 , \3290_b0 );
or ( \3292_b1 , \3208_b1 , \3210_b1 );
xor ( \3292_b0 , \3208_b0 , w_7474 );
not ( w_7474 , w_7475 );
and ( w_7475 , \3210_b1 , \3210_b0 );
or ( \3293_b1 , \3292_b1 , \3213_b1 );
xor ( \3293_b0 , \3292_b0 , w_7476 );
not ( w_7476 , w_7477 );
and ( w_7477 , \3213_b1 , \3213_b0 );
or ( \3294_b1 , \3290_b1 , \3293_b1 );
not ( \3293_b1 , w_7478 );
and ( \3294_b0 , \3290_b0 , w_7479 );
and ( w_7478 , w_7479 , \3293_b0 );
or ( \3295_b1 , \3288_b1 , \3293_b1 );
not ( \3293_b1 , w_7480 );
and ( \3295_b0 , \3288_b0 , w_7481 );
and ( w_7480 , w_7481 , \3293_b0 );
or ( \3297_b1 , \3228_b1 , \3296_b1 );
not ( \3296_b1 , w_7482 );
and ( \3297_b0 , \3228_b0 , w_7483 );
and ( w_7482 , w_7483 , \3296_b0 );
or ( \3298_b1 , \3228_b1 , \3296_b1 );
xor ( \3298_b0 , \3228_b0 , w_7484 );
not ( w_7484 , w_7485 );
and ( w_7485 , \3296_b1 , \3296_b0 );
or ( \3299_b1 , \3272_b1 , \3275_b1 );
xor ( \3299_b0 , \3272_b0 , w_7486 );
not ( w_7486 , w_7487 );
and ( w_7487 , \3275_b1 , \3275_b0 );
or ( \3300_b1 , \1391_b1 , \1431_b1 );
not ( \1431_b1 , w_7488 );
and ( \3300_b0 , \1391_b0 , w_7489 );
and ( w_7488 , w_7489 , \1431_b0 );
or ( \3301_b1 , \1399_b1 , \1429_b1 );
not ( \1429_b1 , w_7490 );
and ( \3301_b0 , \1399_b0 , w_7491 );
and ( w_7490 , w_7491 , \1429_b0 );
or ( \3302_b1 , \3300_b1 , w_7493 );
not ( w_7493 , w_7494 );
and ( \3302_b0 , \3300_b0 , w_7495 );
and ( w_7494 ,  , w_7495 );
buf ( w_7493 , \3301_b1 );
not ( w_7493 , w_7496 );
not (  , w_7497 );
and ( w_7496 , w_7497 , \3301_b0 );
or ( \3303_b1 , \3302_b1 , w_7498 );
xor ( \3303_b0 , \3302_b0 , w_7500 );
not ( w_7500 , w_7501 );
and ( w_7501 , w_7498 , w_7499 );
buf ( w_7498 , \1438_b1 );
not ( w_7498 , w_7502 );
not ( w_7499 , w_7503 );
and ( w_7502 , w_7503 , \1438_b0 );
or ( \3304_b1 , \1586_b1 , \1444_b1 );
not ( \1444_b1 , w_7504 );
and ( \3304_b0 , \1586_b0 , w_7505 );
and ( w_7504 , w_7505 , \1444_b0 );
or ( \3305_b1 , \1616_b1 , \1442_b1 );
not ( \1442_b1 , w_7506 );
and ( \3305_b0 , \1616_b0 , w_7507 );
and ( w_7506 , w_7507 , \1442_b0 );
or ( \3306_b1 , \3304_b1 , w_7509 );
not ( w_7509 , w_7510 );
and ( \3306_b0 , \3304_b0 , w_7511 );
and ( w_7510 ,  , w_7511 );
buf ( w_7509 , \3305_b1 );
not ( w_7509 , w_7512 );
not (  , w_7513 );
and ( w_7512 , w_7513 , \3305_b0 );
or ( \3307_b1 , \3306_b1 , w_7514 );
xor ( \3307_b0 , \3306_b0 , w_7516 );
not ( w_7516 , w_7517 );
and ( w_7517 , w_7514 , w_7515 );
buf ( w_7514 , \1451_b1 );
not ( w_7514 , w_7518 );
not ( w_7515 , w_7519 );
and ( w_7518 , w_7519 , \1451_b0 );
or ( \3308_b1 , \3303_b1 , \3307_b1 );
not ( \3307_b1 , w_7520 );
and ( \3308_b0 , \3303_b0 , w_7521 );
and ( w_7520 , w_7521 , \3307_b0 );
or ( \3309_b1 , \3307_b1 , \3273_b1 );
not ( \3273_b1 , w_7522 );
and ( \3309_b0 , \3307_b0 , w_7523 );
and ( w_7522 , w_7523 , \3273_b0 );
or ( \3310_b1 , \3303_b1 , \3273_b1 );
not ( \3273_b1 , w_7524 );
and ( \3310_b0 , \3303_b0 , w_7525 );
and ( w_7524 , w_7525 , \3273_b0 );
or ( \3312_b1 , \3299_b1 , \3311_b1 );
not ( \3311_b1 , w_7526 );
and ( \3312_b0 , \3299_b0 , w_7527 );
and ( w_7526 , w_7527 , \3311_b0 );
or ( \3313_b1 , \1533_b1 , \1475_b1 );
not ( \1475_b1 , w_7528 );
and ( \3313_b0 , \1533_b0 , w_7529 );
and ( w_7528 , w_7529 , \1475_b0 );
or ( \3314_b1 , \1540_b1 , \1473_b1 );
not ( \1473_b1 , w_7530 );
and ( \3314_b0 , \1540_b0 , w_7531 );
and ( w_7530 , w_7531 , \1473_b0 );
or ( \3315_b1 , \3313_b1 , w_7533 );
not ( w_7533 , w_7534 );
and ( \3315_b0 , \3313_b0 , w_7535 );
and ( w_7534 ,  , w_7535 );
buf ( w_7533 , \3314_b1 );
not ( w_7533 , w_7536 );
not (  , w_7537 );
and ( w_7536 , w_7537 , \3314_b0 );
or ( \3316_b1 , \3315_b1 , w_7538 );
xor ( \3316_b0 , \3315_b0 , w_7540 );
not ( w_7540 , w_7541 );
and ( w_7541 , w_7538 , w_7539 );
buf ( w_7538 , \1482_b1 );
not ( w_7538 , w_7542 );
not ( w_7539 , w_7543 );
and ( w_7542 , w_7543 , \1482_b0 );
or ( \3317_b1 , \3311_b1 , \3316_b1 );
not ( \3316_b1 , w_7544 );
and ( \3317_b0 , \3311_b0 , w_7545 );
and ( w_7544 , w_7545 , \3316_b0 );
or ( \3318_b1 , \3299_b1 , \3316_b1 );
not ( \3316_b1 , w_7546 );
and ( \3318_b0 , \3299_b0 , w_7547 );
and ( w_7546 , w_7547 , \3316_b0 );
or ( \3320_b1 , \1359_b1 , \1336_b1 );
not ( \1336_b1 , w_7548 );
and ( \3320_b0 , \1359_b0 , w_7549 );
and ( w_7548 , w_7549 , \1336_b0 );
or ( \3321_b1 , \1368_b1 , \1333_b1 );
not ( \1333_b1 , w_7550 );
and ( \3321_b0 , \1368_b0 , w_7551 );
and ( w_7550 , w_7551 , \1333_b0 );
or ( \3322_b1 , \3320_b1 , w_7553 );
not ( w_7553 , w_7554 );
and ( \3322_b0 , \3320_b0 , w_7555 );
and ( w_7554 ,  , w_7555 );
buf ( w_7553 , \3321_b1 );
not ( w_7553 , w_7556 );
not (  , w_7557 );
and ( w_7556 , w_7557 , \3321_b0 );
or ( \3323_b1 , \3322_b1 , w_7558 );
xor ( \3323_b0 , \3322_b0 , w_7560 );
not ( w_7560 , w_7561 );
and ( w_7561 , w_7558 , w_7559 );
buf ( w_7558 , \1332_b1 );
not ( w_7558 , w_7562 );
not ( w_7559 , w_7563 );
and ( w_7562 , w_7563 , \1332_b0 );
or ( \3324_b1 , \1407_b1 , \1349_b1 );
not ( \1349_b1 , w_7564 );
and ( \3324_b0 , \1407_b0 , w_7565 );
and ( w_7564 , w_7565 , \1349_b0 );
or ( \3325_b1 , \1416_b1 , \1347_b1 );
not ( \1347_b1 , w_7566 );
and ( \3325_b0 , \1416_b0 , w_7567 );
and ( w_7566 , w_7567 , \1347_b0 );
or ( \3326_b1 , \3324_b1 , w_7569 );
not ( w_7569 , w_7570 );
and ( \3326_b0 , \3324_b0 , w_7571 );
and ( w_7570 ,  , w_7571 );
buf ( w_7569 , \3325_b1 );
not ( w_7569 , w_7572 );
not (  , w_7573 );
and ( w_7572 , w_7573 , \3325_b0 );
or ( \3327_b1 , \3326_b1 , w_7574 );
xor ( \3327_b0 , \3326_b0 , w_7576 );
not ( w_7576 , w_7577 );
and ( w_7577 , w_7574 , w_7575 );
buf ( w_7574 , \1356_b1 );
not ( w_7574 , w_7578 );
not ( w_7575 , w_7579 );
and ( w_7578 , w_7579 , \1356_b0 );
or ( \3328_b1 , \3323_b1 , \3327_b1 );
not ( \3327_b1 , w_7580 );
and ( \3328_b0 , \3323_b0 , w_7581 );
and ( w_7580 , w_7581 , \3327_b0 );
or ( \3329_b1 , \1526_b1 , \1382_b1 );
not ( \1382_b1 , w_7582 );
and ( \3329_b0 , \1526_b0 , w_7583 );
and ( w_7582 , w_7583 , \1382_b0 );
or ( \3330_b1 , \1622_b1 , \1380_b1 );
not ( \1380_b1 , w_7584 );
and ( \3330_b0 , \1622_b0 , w_7585 );
and ( w_7584 , w_7585 , \1380_b0 );
or ( \3331_b1 , \3329_b1 , w_7587 );
not ( w_7587 , w_7588 );
and ( \3331_b0 , \3329_b0 , w_7589 );
and ( w_7588 ,  , w_7589 );
buf ( w_7587 , \3330_b1 );
not ( w_7587 , w_7590 );
not (  , w_7591 );
and ( w_7590 , w_7591 , \3330_b0 );
or ( \3332_b1 , \3331_b1 , w_7592 );
xor ( \3332_b0 , \3331_b0 , w_7594 );
not ( w_7594 , w_7595 );
and ( w_7595 , w_7592 , w_7593 );
buf ( w_7592 , \1389_b1 );
not ( w_7592 , w_7596 );
not ( w_7593 , w_7597 );
and ( w_7596 , w_7597 , \1389_b0 );
or ( \3333_b1 , \3327_b1 , \3332_b1 );
not ( \3332_b1 , w_7598 );
and ( \3333_b0 , \3327_b0 , w_7599 );
and ( w_7598 , w_7599 , \3332_b0 );
or ( \3334_b1 , \3323_b1 , \3332_b1 );
not ( \3332_b1 , w_7600 );
and ( \3334_b0 , \3323_b0 , w_7601 );
and ( w_7600 , w_7601 , \3332_b0 );
or ( \3336_b1 , \3232_b1 , \3236_b1 );
xor ( \3336_b0 , \3232_b0 , w_7602 );
not ( w_7602 , w_7603 );
and ( w_7603 , \3236_b1 , \3236_b0 );
or ( \3337_b1 , \3336_b1 , \3241_b1 );
xor ( \3337_b0 , \3336_b0 , w_7604 );
not ( w_7604 , w_7605 );
and ( w_7605 , \3241_b1 , \3241_b0 );
or ( \3338_b1 , \3335_b1 , \3337_b1 );
not ( \3337_b1 , w_7606 );
and ( \3338_b0 , \3335_b0 , w_7607 );
and ( w_7606 , w_7607 , \3337_b0 );
or ( \3339_b1 , \3256_b1 , \3260_b1 );
xor ( \3339_b0 , \3256_b0 , w_7608 );
not ( w_7608 , w_7609 );
and ( w_7609 , \3260_b1 , \3260_b0 );
or ( \3340_b1 , \3339_b1 , \3265_b1 );
xor ( \3340_b0 , \3339_b0 , w_7610 );
not ( w_7610 , w_7611 );
and ( w_7611 , \3265_b1 , \3265_b0 );
or ( \3341_b1 , \3337_b1 , \3340_b1 );
not ( \3340_b1 , w_7612 );
and ( \3341_b0 , \3337_b0 , w_7613 );
and ( w_7612 , w_7613 , \3340_b0 );
or ( \3342_b1 , \3335_b1 , \3340_b1 );
not ( \3340_b1 , w_7614 );
and ( \3342_b0 , \3335_b0 , w_7615 );
and ( w_7614 , w_7615 , \3340_b0 );
or ( \3344_b1 , \3319_b1 , \3343_b1 );
not ( \3343_b1 , w_7616 );
and ( \3344_b0 , \3319_b0 , w_7617 );
and ( w_7616 , w_7617 , \3343_b0 );
or ( \3345_b1 , \3268_b1 , \3276_b1 );
xor ( \3345_b0 , \3268_b0 , w_7618 );
not ( w_7618 , w_7619 );
and ( w_7619 , \3276_b1 , \3276_b0 );
or ( \3346_b1 , \3345_b1 , \3279_b1 );
xor ( \3346_b0 , \3345_b0 , w_7620 );
not ( w_7620 , w_7621 );
and ( w_7621 , \3279_b1 , \3279_b0 );
or ( \3347_b1 , \3343_b1 , \3346_b1 );
not ( \3346_b1 , w_7622 );
and ( \3347_b0 , \3343_b0 , w_7623 );
and ( w_7622 , w_7623 , \3346_b0 );
or ( \3348_b1 , \3319_b1 , \3346_b1 );
not ( \3346_b1 , w_7624 );
and ( \3348_b0 , \3319_b0 , w_7625 );
and ( w_7624 , w_7625 , \3346_b0 );
or ( \3350_b1 , \3200_b1 , \3202_b1 );
xor ( \3350_b0 , \3200_b0 , w_7626 );
not ( w_7626 , w_7627 );
and ( w_7627 , \3202_b1 , \3202_b0 );
or ( \3351_b1 , \3350_b1 , \3205_b1 );
xor ( \3351_b0 , \3350_b0 , w_7628 );
not ( w_7628 , w_7629 );
and ( w_7629 , \3205_b1 , \3205_b0 );
or ( \3352_b1 , \3349_b1 , \3351_b1 );
not ( \3351_b1 , w_7630 );
and ( \3352_b0 , \3349_b0 , w_7631 );
and ( w_7630 , w_7631 , \3351_b0 );
or ( \3353_b1 , \3252_b1 , \3282_b1 );
xor ( \3353_b0 , \3252_b0 , w_7632 );
not ( w_7632 , w_7633 );
and ( w_7633 , \3282_b1 , \3282_b0 );
or ( \3354_b1 , \3353_b1 , \3285_b1 );
xor ( \3354_b0 , \3353_b0 , w_7634 );
not ( w_7634 , w_7635 );
and ( w_7635 , \3285_b1 , \3285_b0 );
or ( \3355_b1 , \3351_b1 , \3354_b1 );
not ( \3354_b1 , w_7636 );
and ( \3355_b0 , \3351_b0 , w_7637 );
and ( w_7636 , w_7637 , \3354_b0 );
or ( \3356_b1 , \3349_b1 , \3354_b1 );
not ( \3354_b1 , w_7638 );
and ( \3356_b0 , \3349_b0 , w_7639 );
and ( w_7638 , w_7639 , \3354_b0 );
or ( \3358_b1 , \3288_b1 , \3290_b1 );
xor ( \3358_b0 , \3288_b0 , w_7640 );
not ( w_7640 , w_7641 );
and ( w_7641 , \3290_b1 , \3290_b0 );
or ( \3359_b1 , \3358_b1 , \3293_b1 );
xor ( \3359_b0 , \3358_b0 , w_7642 );
not ( w_7642 , w_7643 );
and ( w_7643 , \3293_b1 , \3293_b0 );
or ( \3360_b1 , \3357_b1 , \3359_b1 );
not ( \3359_b1 , w_7644 );
and ( \3360_b0 , \3357_b0 , w_7645 );
and ( w_7644 , w_7645 , \3359_b0 );
or ( \3361_b1 , \3357_b1 , \3359_b1 );
xor ( \3361_b0 , \3357_b0 , w_7646 );
not ( w_7646 , w_7647 );
and ( w_7647 , \3359_b1 , \3359_b0 );
or ( \3362_b1 , \3349_b1 , \3351_b1 );
xor ( \3362_b0 , \3349_b0 , w_7648 );
not ( w_7648 , w_7649 );
and ( w_7649 , \3351_b1 , \3351_b0 );
or ( \3363_b1 , \3362_b1 , \3354_b1 );
xor ( \3363_b0 , \3362_b0 , w_7650 );
not ( w_7650 , w_7651 );
and ( w_7651 , \3354_b1 , \3354_b0 );
or ( \3364_b1 , \1616_b1 , \1431_b1 );
not ( \1431_b1 , w_7652 );
and ( \3364_b0 , \1616_b0 , w_7653 );
and ( w_7652 , w_7653 , \1431_b0 );
or ( \3365_b1 , \1391_b1 , \1429_b1 );
not ( \1429_b1 , w_7654 );
and ( \3365_b0 , \1391_b0 , w_7655 );
and ( w_7654 , w_7655 , \1429_b0 );
or ( \3366_b1 , \3364_b1 , w_7657 );
not ( w_7657 , w_7658 );
and ( \3366_b0 , \3364_b0 , w_7659 );
and ( w_7658 ,  , w_7659 );
buf ( w_7657 , \3365_b1 );
not ( w_7657 , w_7660 );
not (  , w_7661 );
and ( w_7660 , w_7661 , \3365_b0 );
or ( \3367_b1 , \3366_b1 , w_7662 );
xor ( \3367_b0 , \3366_b0 , w_7664 );
not ( w_7664 , w_7665 );
and ( w_7665 , w_7662 , w_7663 );
buf ( w_7662 , \1438_b1 );
not ( w_7662 , w_7666 );
not ( w_7663 , w_7667 );
and ( w_7666 , w_7667 , \1438_b0 );
or ( \3368_b1 , \1498_b1 , \1473_b1 );
not ( \1473_b1 , w_7668 );
and ( \3368_b0 , \1498_b0 , w_7669 );
and ( w_7668 , w_7669 , \1473_b0 );
buf ( \3369_b1 , \3368_b1 );
not ( \3369_b1 , w_7670 );
not ( \3369_b0 , w_7671 );
and ( w_7670 , w_7671 , \3368_b0 );
or ( \3370_b1 , \3369_b1 , \1482_b1 );
not ( \1482_b1 , w_7672 );
and ( \3370_b0 , \3369_b0 , w_7673 );
and ( w_7672 , w_7673 , \1482_b0 );
or ( \3371_b1 , \3367_b1 , \3370_b1 );
not ( \3370_b1 , w_7674 );
and ( \3371_b0 , \3367_b0 , w_7675 );
and ( w_7674 , w_7675 , \3370_b0 );
or ( \3372_b1 , \1540_b1 , \1460_b1 );
not ( \1460_b1 , w_7676 );
and ( \3372_b0 , \1540_b0 , w_7677 );
and ( w_7676 , w_7677 , \1460_b0 );
or ( \3373_b1 , \1517_b1 , \1458_b1 );
not ( \1458_b1 , w_7678 );
and ( \3373_b0 , \1517_b0 , w_7679 );
and ( w_7678 , w_7679 , \1458_b0 );
or ( \3374_b1 , \3372_b1 , w_7681 );
not ( w_7681 , w_7682 );
and ( \3374_b0 , \3372_b0 , w_7683 );
and ( w_7682 ,  , w_7683 );
buf ( w_7681 , \3373_b1 );
not ( w_7681 , w_7684 );
not (  , w_7685 );
and ( w_7684 , w_7685 , \3373_b0 );
or ( \3375_b1 , \3374_b1 , w_7686 );
xor ( \3375_b0 , \3374_b0 , w_7688 );
not ( w_7688 , w_7689 );
and ( w_7689 , w_7686 , w_7687 );
buf ( w_7686 , \1467_b1 );
not ( w_7686 , w_7690 );
not ( w_7687 , w_7691 );
and ( w_7690 , w_7691 , \1467_b0 );
or ( \3376_b1 , \3371_b1 , \3375_b1 );
not ( \3375_b1 , w_7692 );
and ( \3376_b0 , \3371_b0 , w_7693 );
and ( w_7692 , w_7693 , \3375_b0 );
or ( \3377_b1 , \1553_b1 , \1475_b1 );
not ( \1475_b1 , w_7694 );
and ( \3377_b0 , \1553_b0 , w_7695 );
and ( w_7694 , w_7695 , \1475_b0 );
or ( \3378_b1 , \1533_b1 , \1473_b1 );
not ( \1473_b1 , w_7696 );
and ( \3378_b0 , \1533_b0 , w_7697 );
and ( w_7696 , w_7697 , \1473_b0 );
or ( \3379_b1 , \3377_b1 , w_7699 );
not ( w_7699 , w_7700 );
and ( \3379_b0 , \3377_b0 , w_7701 );
and ( w_7700 ,  , w_7701 );
buf ( w_7699 , \3378_b1 );
not ( w_7699 , w_7702 );
not (  , w_7703 );
and ( w_7702 , w_7703 , \3378_b0 );
or ( \3380_b1 , \3379_b1 , w_7704 );
xor ( \3380_b0 , \3379_b0 , w_7706 );
not ( w_7706 , w_7707 );
and ( w_7707 , w_7704 , w_7705 );
buf ( w_7704 , \1482_b1 );
not ( w_7704 , w_7708 );
not ( w_7705 , w_7709 );
and ( w_7708 , w_7709 , \1482_b0 );
or ( \3381_b1 , \3375_b1 , \3380_b1 );
not ( \3380_b1 , w_7710 );
and ( \3381_b0 , \3375_b0 , w_7711 );
and ( w_7710 , w_7711 , \3380_b0 );
or ( \3382_b1 , \3371_b1 , \3380_b1 );
not ( \3380_b1 , w_7712 );
and ( \3382_b0 , \3371_b0 , w_7713 );
and ( w_7712 , w_7713 , \3380_b0 );
or ( \3384_b1 , \1399_b1 , \1336_b1 );
not ( \1336_b1 , w_7714 );
and ( \3384_b0 , \1399_b0 , w_7715 );
and ( w_7714 , w_7715 , \1336_b0 );
or ( \3385_b1 , \1359_b1 , \1333_b1 );
not ( \1333_b1 , w_7716 );
and ( \3385_b0 , \1359_b0 , w_7717 );
and ( w_7716 , w_7717 , \1333_b0 );
or ( \3386_b1 , \3384_b1 , w_7719 );
not ( w_7719 , w_7720 );
and ( \3386_b0 , \3384_b0 , w_7721 );
and ( w_7720 ,  , w_7721 );
buf ( w_7719 , \3385_b1 );
not ( w_7719 , w_7722 );
not (  , w_7723 );
and ( w_7722 , w_7723 , \3385_b0 );
or ( \3387_b1 , \3386_b1 , w_7724 );
xor ( \3387_b0 , \3386_b0 , w_7726 );
not ( w_7726 , w_7727 );
and ( w_7727 , w_7724 , w_7725 );
buf ( w_7724 , \1332_b1 );
not ( w_7724 , w_7728 );
not ( w_7725 , w_7729 );
and ( w_7728 , w_7729 , \1332_b0 );
or ( \3388_b1 , \1416_b1 , \1444_b1 );
not ( \1444_b1 , w_7730 );
and ( \3388_b0 , \1416_b0 , w_7731 );
and ( w_7730 , w_7731 , \1444_b0 );
or ( \3389_b1 , \1586_b1 , \1442_b1 );
not ( \1442_b1 , w_7732 );
and ( \3389_b0 , \1586_b0 , w_7733 );
and ( w_7732 , w_7733 , \1442_b0 );
or ( \3390_b1 , \3388_b1 , w_7735 );
not ( w_7735 , w_7736 );
and ( \3390_b0 , \3388_b0 , w_7737 );
and ( w_7736 ,  , w_7737 );
buf ( w_7735 , \3389_b1 );
not ( w_7735 , w_7738 );
not (  , w_7739 );
and ( w_7738 , w_7739 , \3389_b0 );
or ( \3391_b1 , \3390_b1 , w_7740 );
xor ( \3391_b0 , \3390_b0 , w_7742 );
not ( w_7742 , w_7743 );
and ( w_7743 , w_7740 , w_7741 );
buf ( w_7740 , \1451_b1 );
not ( w_7740 , w_7744 );
not ( w_7741 , w_7745 );
and ( w_7744 , w_7745 , \1451_b0 );
or ( \3392_b1 , \3387_b1 , \3391_b1 );
not ( \3391_b1 , w_7746 );
and ( \3392_b0 , \3387_b0 , w_7747 );
and ( w_7746 , w_7747 , \3391_b0 );
or ( \3393_b1 , \1622_b1 , \1349_b1 );
not ( \1349_b1 , w_7748 );
and ( \3393_b0 , \1622_b0 , w_7749 );
and ( w_7748 , w_7749 , \1349_b0 );
or ( \3394_b1 , \1407_b1 , \1347_b1 );
not ( \1347_b1 , w_7750 );
and ( \3394_b0 , \1407_b0 , w_7751 );
and ( w_7750 , w_7751 , \1347_b0 );
or ( \3395_b1 , \3393_b1 , w_7753 );
not ( w_7753 , w_7754 );
and ( \3395_b0 , \3393_b0 , w_7755 );
and ( w_7754 ,  , w_7755 );
buf ( w_7753 , \3394_b1 );
not ( w_7753 , w_7756 );
not (  , w_7757 );
and ( w_7756 , w_7757 , \3394_b0 );
or ( \3396_b1 , \3395_b1 , w_7758 );
xor ( \3396_b0 , \3395_b0 , w_7760 );
not ( w_7760 , w_7761 );
and ( w_7761 , w_7758 , w_7759 );
buf ( w_7758 , \1356_b1 );
not ( w_7758 , w_7762 );
not ( w_7759 , w_7763 );
and ( w_7762 , w_7763 , \1356_b0 );
or ( \3397_b1 , \3391_b1 , \3396_b1 );
not ( \3396_b1 , w_7764 );
and ( \3397_b0 , \3391_b0 , w_7765 );
and ( w_7764 , w_7765 , \3396_b0 );
or ( \3398_b1 , \3387_b1 , \3396_b1 );
not ( \3396_b1 , w_7766 );
and ( \3398_b0 , \3387_b0 , w_7767 );
and ( w_7766 , w_7767 , \3396_b0 );
or ( \3400_b1 , \1517_b1 , \1382_b1 );
not ( \1382_b1 , w_7768 );
and ( \3400_b0 , \1517_b0 , w_7769 );
and ( w_7768 , w_7769 , \1382_b0 );
or ( \3401_b1 , \1526_b1 , \1380_b1 );
not ( \1380_b1 , w_7770 );
and ( \3401_b0 , \1526_b0 , w_7771 );
and ( w_7770 , w_7771 , \1380_b0 );
or ( \3402_b1 , \3400_b1 , w_7773 );
not ( w_7773 , w_7774 );
and ( \3402_b0 , \3400_b0 , w_7775 );
and ( w_7774 ,  , w_7775 );
buf ( w_7773 , \3401_b1 );
not ( w_7773 , w_7776 );
not (  , w_7777 );
and ( w_7776 , w_7777 , \3401_b0 );
or ( \3403_b1 , \3402_b1 , w_7778 );
xor ( \3403_b0 , \3402_b0 , w_7780 );
not ( w_7780 , w_7781 );
and ( w_7781 , w_7778 , w_7779 );
buf ( w_7778 , \1389_b1 );
not ( w_7778 , w_7782 );
not ( w_7779 , w_7783 );
and ( w_7782 , w_7783 , \1389_b0 );
or ( \3404_b1 , \1533_b1 , \1460_b1 );
not ( \1460_b1 , w_7784 );
and ( \3404_b0 , \1533_b0 , w_7785 );
and ( w_7784 , w_7785 , \1460_b0 );
or ( \3405_b1 , \1540_b1 , \1458_b1 );
not ( \1458_b1 , w_7786 );
and ( \3405_b0 , \1540_b0 , w_7787 );
and ( w_7786 , w_7787 , \1458_b0 );
or ( \3406_b1 , \3404_b1 , w_7789 );
not ( w_7789 , w_7790 );
and ( \3406_b0 , \3404_b0 , w_7791 );
and ( w_7790 ,  , w_7791 );
buf ( w_7789 , \3405_b1 );
not ( w_7789 , w_7792 );
not (  , w_7793 );
and ( w_7792 , w_7793 , \3405_b0 );
or ( \3407_b1 , \3406_b1 , w_7794 );
xor ( \3407_b0 , \3406_b0 , w_7796 );
not ( w_7796 , w_7797 );
and ( w_7797 , w_7794 , w_7795 );
buf ( w_7794 , \1467_b1 );
not ( w_7794 , w_7798 );
not ( w_7795 , w_7799 );
and ( w_7798 , w_7799 , \1467_b0 );
or ( \3408_b1 , \3403_b1 , \3407_b1 );
not ( \3407_b1 , w_7800 );
and ( \3408_b0 , \3403_b0 , w_7801 );
and ( w_7800 , w_7801 , \3407_b0 );
or ( \3409_b1 , \1498_b1 , \1475_b1 );
not ( \1475_b1 , w_7802 );
and ( \3409_b0 , \1498_b0 , w_7803 );
and ( w_7802 , w_7803 , \1475_b0 );
or ( \3410_b1 , \1553_b1 , \1473_b1 );
not ( \1473_b1 , w_7804 );
and ( \3410_b0 , \1553_b0 , w_7805 );
and ( w_7804 , w_7805 , \1473_b0 );
or ( \3411_b1 , \3409_b1 , w_7807 );
not ( w_7807 , w_7808 );
and ( \3411_b0 , \3409_b0 , w_7809 );
and ( w_7808 ,  , w_7809 );
buf ( w_7807 , \3410_b1 );
not ( w_7807 , w_7810 );
not (  , w_7811 );
and ( w_7810 , w_7811 , \3410_b0 );
or ( \3412_b1 , \3411_b1 , w_7812 );
xor ( \3412_b0 , \3411_b0 , w_7814 );
not ( w_7814 , w_7815 );
and ( w_7815 , w_7812 , w_7813 );
buf ( w_7812 , \1482_b1 );
not ( w_7812 , w_7816 );
not ( w_7813 , w_7817 );
and ( w_7816 , w_7817 , \1482_b0 );
or ( \3413_b1 , \3407_b1 , \3412_b1 );
not ( \3412_b1 , w_7818 );
and ( \3413_b0 , \3407_b0 , w_7819 );
and ( w_7818 , w_7819 , \3412_b0 );
or ( \3414_b1 , \3403_b1 , \3412_b1 );
not ( \3412_b1 , w_7820 );
and ( \3414_b0 , \3403_b0 , w_7821 );
and ( w_7820 , w_7821 , \3412_b0 );
or ( \3416_b1 , \3399_b1 , \3415_b1 );
not ( \3415_b1 , w_7822 );
and ( \3416_b0 , \3399_b0 , w_7823 );
and ( w_7822 , w_7823 , \3415_b0 );
or ( \3417_b1 , \3303_b1 , \3307_b1 );
xor ( \3417_b0 , \3303_b0 , w_7824 );
not ( w_7824 , w_7825 );
and ( w_7825 , \3307_b1 , \3307_b0 );
or ( \3418_b1 , \3417_b1 , \3273_b1 );
xor ( \3418_b0 , \3417_b0 , w_7826 );
not ( w_7826 , w_7827 );
and ( w_7827 , \3273_b1 , \3273_b0 );
or ( \3419_b1 , \3415_b1 , \3418_b1 );
not ( \3418_b1 , w_7828 );
and ( \3419_b0 , \3415_b0 , w_7829 );
and ( w_7828 , w_7829 , \3418_b0 );
or ( \3420_b1 , \3399_b1 , \3418_b1 );
not ( \3418_b1 , w_7830 );
and ( \3420_b0 , \3399_b0 , w_7831 );
and ( w_7830 , w_7831 , \3418_b0 );
or ( \3422_b1 , \3383_b1 , \3421_b1 );
not ( \3421_b1 , w_7832 );
and ( \3422_b0 , \3383_b0 , w_7833 );
and ( w_7832 , w_7833 , \3421_b0 );
or ( \3423_b1 , \3299_b1 , \3311_b1 );
xor ( \3423_b0 , \3299_b0 , w_7834 );
not ( w_7834 , w_7835 );
and ( w_7835 , \3311_b1 , \3311_b0 );
or ( \3424_b1 , \3423_b1 , \3316_b1 );
xor ( \3424_b0 , \3423_b0 , w_7836 );
not ( w_7836 , w_7837 );
and ( w_7837 , \3316_b1 , \3316_b0 );
or ( \3425_b1 , \3421_b1 , \3424_b1 );
not ( \3424_b1 , w_7838 );
and ( \3425_b0 , \3421_b0 , w_7839 );
and ( w_7838 , w_7839 , \3424_b0 );
or ( \3426_b1 , \3383_b1 , \3424_b1 );
not ( \3424_b1 , w_7840 );
and ( \3426_b0 , \3383_b0 , w_7841 );
and ( w_7840 , w_7841 , \3424_b0 );
or ( \3428_b1 , \3244_b1 , \3246_b1 );
xor ( \3428_b0 , \3244_b0 , w_7842 );
not ( w_7842 , w_7843 );
and ( w_7843 , \3246_b1 , \3246_b0 );
or ( \3429_b1 , \3428_b1 , \3249_b1 );
xor ( \3429_b0 , \3428_b0 , w_7844 );
not ( w_7844 , w_7845 );
and ( w_7845 , \3249_b1 , \3249_b0 );
or ( \3430_b1 , \3427_b1 , \3429_b1 );
not ( \3429_b1 , w_7846 );
and ( \3430_b0 , \3427_b0 , w_7847 );
and ( w_7846 , w_7847 , \3429_b0 );
or ( \3431_b1 , \3319_b1 , \3343_b1 );
xor ( \3431_b0 , \3319_b0 , w_7848 );
not ( w_7848 , w_7849 );
and ( w_7849 , \3343_b1 , \3343_b0 );
or ( \3432_b1 , \3431_b1 , \3346_b1 );
xor ( \3432_b0 , \3431_b0 , w_7850 );
not ( w_7850 , w_7851 );
and ( w_7851 , \3346_b1 , \3346_b0 );
or ( \3433_b1 , \3429_b1 , \3432_b1 );
not ( \3432_b1 , w_7852 );
and ( \3433_b0 , \3429_b0 , w_7853 );
and ( w_7852 , w_7853 , \3432_b0 );
or ( \3434_b1 , \3427_b1 , \3432_b1 );
not ( \3432_b1 , w_7854 );
and ( \3434_b0 , \3427_b0 , w_7855 );
and ( w_7854 , w_7855 , \3432_b0 );
or ( \3436_b1 , \3363_b1 , \3435_b1 );
not ( \3435_b1 , w_7856 );
and ( \3436_b0 , \3363_b0 , w_7857 );
and ( w_7856 , w_7857 , \3435_b0 );
or ( \3437_b1 , \3363_b1 , \3435_b1 );
xor ( \3437_b0 , \3363_b0 , w_7858 );
not ( w_7858 , w_7859 );
and ( w_7859 , \3435_b1 , \3435_b0 );
or ( \3438_b1 , \3427_b1 , \3429_b1 );
xor ( \3438_b0 , \3427_b0 , w_7860 );
not ( w_7860 , w_7861 );
and ( w_7861 , \3429_b1 , \3429_b0 );
or ( \3439_b1 , \3438_b1 , \3432_b1 );
xor ( \3439_b0 , \3438_b0 , w_7862 );
not ( w_7862 , w_7863 );
and ( w_7863 , \3432_b1 , \3432_b0 );
or ( \3440_b1 , \3367_b1 , \3370_b1 );
xor ( \3440_b0 , \3367_b0 , w_7864 );
not ( w_7864 , w_7865 );
and ( w_7865 , \3370_b1 , \3370_b0 );
or ( \3441_b1 , \1586_b1 , \1431_b1 );
not ( \1431_b1 , w_7866 );
and ( \3441_b0 , \1586_b0 , w_7867 );
and ( w_7866 , w_7867 , \1431_b0 );
or ( \3442_b1 , \1616_b1 , \1429_b1 );
not ( \1429_b1 , w_7868 );
and ( \3442_b0 , \1616_b0 , w_7869 );
and ( w_7868 , w_7869 , \1429_b0 );
or ( \3443_b1 , \3441_b1 , w_7871 );
not ( w_7871 , w_7872 );
and ( \3443_b0 , \3441_b0 , w_7873 );
and ( w_7872 ,  , w_7873 );
buf ( w_7871 , \3442_b1 );
not ( w_7871 , w_7874 );
not (  , w_7875 );
and ( w_7874 , w_7875 , \3442_b0 );
or ( \3444_b1 , \3443_b1 , w_7876 );
xor ( \3444_b0 , \3443_b0 , w_7878 );
not ( w_7878 , w_7879 );
and ( w_7879 , w_7876 , w_7877 );
buf ( w_7876 , \1438_b1 );
not ( w_7876 , w_7880 );
not ( w_7877 , w_7881 );
and ( w_7880 , w_7881 , \1438_b0 );
or ( \3445_b1 , \1407_b1 , \1444_b1 );
not ( \1444_b1 , w_7882 );
and ( \3445_b0 , \1407_b0 , w_7883 );
and ( w_7882 , w_7883 , \1444_b0 );
or ( \3446_b1 , \1416_b1 , \1442_b1 );
not ( \1442_b1 , w_7884 );
and ( \3446_b0 , \1416_b0 , w_7885 );
and ( w_7884 , w_7885 , \1442_b0 );
or ( \3447_b1 , \3445_b1 , w_7887 );
not ( w_7887 , w_7888 );
and ( \3447_b0 , \3445_b0 , w_7889 );
and ( w_7888 ,  , w_7889 );
buf ( w_7887 , \3446_b1 );
not ( w_7887 , w_7890 );
not (  , w_7891 );
and ( w_7890 , w_7891 , \3446_b0 );
or ( \3448_b1 , \3447_b1 , w_7892 );
xor ( \3448_b0 , \3447_b0 , w_7894 );
not ( w_7894 , w_7895 );
and ( w_7895 , w_7892 , w_7893 );
buf ( w_7892 , \1451_b1 );
not ( w_7892 , w_7896 );
not ( w_7893 , w_7897 );
and ( w_7896 , w_7897 , \1451_b0 );
or ( \3449_b1 , \3444_b1 , \3448_b1 );
not ( \3448_b1 , w_7898 );
and ( \3449_b0 , \3444_b0 , w_7899 );
and ( w_7898 , w_7899 , \3448_b0 );
or ( \3450_b1 , \3448_b1 , \3368_b1 );
not ( \3368_b1 , w_7900 );
and ( \3450_b0 , \3448_b0 , w_7901 );
and ( w_7900 , w_7901 , \3368_b0 );
or ( \3451_b1 , \3444_b1 , \3368_b1 );
not ( \3368_b1 , w_7902 );
and ( \3451_b0 , \3444_b0 , w_7903 );
and ( w_7902 , w_7903 , \3368_b0 );
or ( \3453_b1 , \3440_b1 , \3452_b1 );
not ( \3452_b1 , w_7904 );
and ( \3453_b0 , \3440_b0 , w_7905 );
and ( w_7904 , w_7905 , \3452_b0 );
or ( \3454_b1 , \1391_b1 , \1336_b1 );
not ( \1336_b1 , w_7906 );
and ( \3454_b0 , \1391_b0 , w_7907 );
and ( w_7906 , w_7907 , \1336_b0 );
or ( \3455_b1 , \1399_b1 , \1333_b1 );
not ( \1333_b1 , w_7908 );
and ( \3455_b0 , \1399_b0 , w_7909 );
and ( w_7908 , w_7909 , \1333_b0 );
or ( \3456_b1 , \3454_b1 , w_7911 );
not ( w_7911 , w_7912 );
and ( \3456_b0 , \3454_b0 , w_7913 );
and ( w_7912 ,  , w_7913 );
buf ( w_7911 , \3455_b1 );
not ( w_7911 , w_7914 );
not (  , w_7915 );
and ( w_7914 , w_7915 , \3455_b0 );
or ( \3457_b1 , \3456_b1 , w_7916 );
xor ( \3457_b0 , \3456_b0 , w_7918 );
not ( w_7918 , w_7919 );
and ( w_7919 , w_7916 , w_7917 );
buf ( w_7916 , \1332_b1 );
not ( w_7916 , w_7920 );
not ( w_7917 , w_7921 );
and ( w_7920 , w_7921 , \1332_b0 );
or ( \3458_b1 , \1526_b1 , \1349_b1 );
not ( \1349_b1 , w_7922 );
and ( \3458_b0 , \1526_b0 , w_7923 );
and ( w_7922 , w_7923 , \1349_b0 );
or ( \3459_b1 , \1622_b1 , \1347_b1 );
not ( \1347_b1 , w_7924 );
and ( \3459_b0 , \1622_b0 , w_7925 );
and ( w_7924 , w_7925 , \1347_b0 );
or ( \3460_b1 , \3458_b1 , w_7927 );
not ( w_7927 , w_7928 );
and ( \3460_b0 , \3458_b0 , w_7929 );
and ( w_7928 ,  , w_7929 );
buf ( w_7927 , \3459_b1 );
not ( w_7927 , w_7930 );
not (  , w_7931 );
and ( w_7930 , w_7931 , \3459_b0 );
or ( \3461_b1 , \3460_b1 , w_7932 );
xor ( \3461_b0 , \3460_b0 , w_7934 );
not ( w_7934 , w_7935 );
and ( w_7935 , w_7932 , w_7933 );
buf ( w_7932 , \1356_b1 );
not ( w_7932 , w_7936 );
not ( w_7933 , w_7937 );
and ( w_7936 , w_7937 , \1356_b0 );
or ( \3462_b1 , \3457_b1 , \3461_b1 );
not ( \3461_b1 , w_7938 );
and ( \3462_b0 , \3457_b0 , w_7939 );
and ( w_7938 , w_7939 , \3461_b0 );
or ( \3463_b1 , \1540_b1 , \1382_b1 );
not ( \1382_b1 , w_7940 );
and ( \3463_b0 , \1540_b0 , w_7941 );
and ( w_7940 , w_7941 , \1382_b0 );
or ( \3464_b1 , \1517_b1 , \1380_b1 );
not ( \1380_b1 , w_7942 );
and ( \3464_b0 , \1517_b0 , w_7943 );
and ( w_7942 , w_7943 , \1380_b0 );
or ( \3465_b1 , \3463_b1 , w_7945 );
not ( w_7945 , w_7946 );
and ( \3465_b0 , \3463_b0 , w_7947 );
and ( w_7946 ,  , w_7947 );
buf ( w_7945 , \3464_b1 );
not ( w_7945 , w_7948 );
not (  , w_7949 );
and ( w_7948 , w_7949 , \3464_b0 );
or ( \3466_b1 , \3465_b1 , w_7950 );
xor ( \3466_b0 , \3465_b0 , w_7952 );
not ( w_7952 , w_7953 );
and ( w_7953 , w_7950 , w_7951 );
buf ( w_7950 , \1389_b1 );
not ( w_7950 , w_7954 );
not ( w_7951 , w_7955 );
and ( w_7954 , w_7955 , \1389_b0 );
or ( \3467_b1 , \3461_b1 , \3466_b1 );
not ( \3466_b1 , w_7956 );
and ( \3467_b0 , \3461_b0 , w_7957 );
and ( w_7956 , w_7957 , \3466_b0 );
or ( \3468_b1 , \3457_b1 , \3466_b1 );
not ( \3466_b1 , w_7958 );
and ( \3468_b0 , \3457_b0 , w_7959 );
and ( w_7958 , w_7959 , \3466_b0 );
or ( \3470_b1 , \3452_b1 , \3469_b1 );
not ( \3469_b1 , w_7960 );
and ( \3470_b0 , \3452_b0 , w_7961 );
and ( w_7960 , w_7961 , \3469_b0 );
or ( \3471_b1 , \3440_b1 , \3469_b1 );
not ( \3469_b1 , w_7962 );
and ( \3471_b0 , \3440_b0 , w_7963 );
and ( w_7962 , w_7963 , \3469_b0 );
or ( \3473_b1 , \3323_b1 , \3327_b1 );
xor ( \3473_b0 , \3323_b0 , w_7964 );
not ( w_7964 , w_7965 );
and ( w_7965 , \3327_b1 , \3327_b0 );
or ( \3474_b1 , \3473_b1 , \3332_b1 );
xor ( \3474_b0 , \3473_b0 , w_7966 );
not ( w_7966 , w_7967 );
and ( w_7967 , \3332_b1 , \3332_b0 );
or ( \3475_b1 , \3472_b1 , \3474_b1 );
not ( \3474_b1 , w_7968 );
and ( \3475_b0 , \3472_b0 , w_7969 );
and ( w_7968 , w_7969 , \3474_b0 );
or ( \3476_b1 , \3371_b1 , \3375_b1 );
xor ( \3476_b0 , \3371_b0 , w_7970 );
not ( w_7970 , w_7971 );
and ( w_7971 , \3375_b1 , \3375_b0 );
or ( \3477_b1 , \3476_b1 , \3380_b1 );
xor ( \3477_b0 , \3476_b0 , w_7972 );
not ( w_7972 , w_7973 );
and ( w_7973 , \3380_b1 , \3380_b0 );
or ( \3478_b1 , \3474_b1 , \3477_b1 );
not ( \3477_b1 , w_7974 );
and ( \3478_b0 , \3474_b0 , w_7975 );
and ( w_7974 , w_7975 , \3477_b0 );
or ( \3479_b1 , \3472_b1 , \3477_b1 );
not ( \3477_b1 , w_7976 );
and ( \3479_b0 , \3472_b0 , w_7977 );
and ( w_7976 , w_7977 , \3477_b0 );
or ( \3481_b1 , \3335_b1 , \3337_b1 );
xor ( \3481_b0 , \3335_b0 , w_7978 );
not ( w_7978 , w_7979 );
and ( w_7979 , \3337_b1 , \3337_b0 );
or ( \3482_b1 , \3481_b1 , \3340_b1 );
xor ( \3482_b0 , \3481_b0 , w_7980 );
not ( w_7980 , w_7981 );
and ( w_7981 , \3340_b1 , \3340_b0 );
or ( \3483_b1 , \3480_b1 , \3482_b1 );
not ( \3482_b1 , w_7982 );
and ( \3483_b0 , \3480_b0 , w_7983 );
and ( w_7982 , w_7983 , \3482_b0 );
or ( \3484_b1 , \3383_b1 , \3421_b1 );
xor ( \3484_b0 , \3383_b0 , w_7984 );
not ( w_7984 , w_7985 );
and ( w_7985 , \3421_b1 , \3421_b0 );
or ( \3485_b1 , \3484_b1 , \3424_b1 );
xor ( \3485_b0 , \3484_b0 , w_7986 );
not ( w_7986 , w_7987 );
and ( w_7987 , \3424_b1 , \3424_b0 );
or ( \3486_b1 , \3482_b1 , \3485_b1 );
not ( \3485_b1 , w_7988 );
and ( \3486_b0 , \3482_b0 , w_7989 );
and ( w_7988 , w_7989 , \3485_b0 );
or ( \3487_b1 , \3480_b1 , \3485_b1 );
not ( \3485_b1 , w_7990 );
and ( \3487_b0 , \3480_b0 , w_7991 );
and ( w_7990 , w_7991 , \3485_b0 );
or ( \3489_b1 , \3439_b1 , \3488_b1 );
not ( \3488_b1 , w_7992 );
and ( \3489_b0 , \3439_b0 , w_7993 );
and ( w_7992 , w_7993 , \3488_b0 );
or ( \3490_b1 , \3439_b1 , \3488_b1 );
xor ( \3490_b0 , \3439_b0 , w_7994 );
not ( w_7994 , w_7995 );
and ( w_7995 , \3488_b1 , \3488_b0 );
or ( \3491_b1 , \3480_b1 , \3482_b1 );
xor ( \3491_b0 , \3480_b0 , w_7996 );
not ( w_7996 , w_7997 );
and ( w_7997 , \3482_b1 , \3482_b0 );
or ( \3492_b1 , \3491_b1 , \3485_b1 );
xor ( \3492_b0 , \3491_b0 , w_7998 );
not ( w_7998 , w_7999 );
and ( w_7999 , \3485_b1 , \3485_b0 );
or ( \3493_b1 , \1616_b1 , \1336_b1 );
not ( \1336_b1 , w_8000 );
and ( \3493_b0 , \1616_b0 , w_8001 );
and ( w_8000 , w_8001 , \1336_b0 );
or ( \3494_b1 , \1391_b1 , \1333_b1 );
not ( \1333_b1 , w_8002 );
and ( \3494_b0 , \1391_b0 , w_8003 );
and ( w_8002 , w_8003 , \1333_b0 );
or ( \3495_b1 , \3493_b1 , w_8005 );
not ( w_8005 , w_8006 );
and ( \3495_b0 , \3493_b0 , w_8007 );
and ( w_8006 ,  , w_8007 );
buf ( w_8005 , \3494_b1 );
not ( w_8005 , w_8008 );
not (  , w_8009 );
and ( w_8008 , w_8009 , \3494_b0 );
or ( \3496_b1 , \3495_b1 , w_8010 );
xor ( \3496_b0 , \3495_b0 , w_8012 );
not ( w_8012 , w_8013 );
and ( w_8013 , w_8010 , w_8011 );
buf ( w_8010 , \1332_b1 );
not ( w_8010 , w_8014 );
not ( w_8011 , w_8015 );
and ( w_8014 , w_8015 , \1332_b0 );
or ( \3497_b1 , \1622_b1 , \1444_b1 );
not ( \1444_b1 , w_8016 );
and ( \3497_b0 , \1622_b0 , w_8017 );
and ( w_8016 , w_8017 , \1444_b0 );
or ( \3498_b1 , \1407_b1 , \1442_b1 );
not ( \1442_b1 , w_8018 );
and ( \3498_b0 , \1407_b0 , w_8019 );
and ( w_8018 , w_8019 , \1442_b0 );
or ( \3499_b1 , \3497_b1 , w_8021 );
not ( w_8021 , w_8022 );
and ( \3499_b0 , \3497_b0 , w_8023 );
and ( w_8022 ,  , w_8023 );
buf ( w_8021 , \3498_b1 );
not ( w_8021 , w_8024 );
not (  , w_8025 );
and ( w_8024 , w_8025 , \3498_b0 );
or ( \3500_b1 , \3499_b1 , w_8026 );
xor ( \3500_b0 , \3499_b0 , w_8028 );
not ( w_8028 , w_8029 );
and ( w_8029 , w_8026 , w_8027 );
buf ( w_8026 , \1451_b1 );
not ( w_8026 , w_8030 );
not ( w_8027 , w_8031 );
and ( w_8030 , w_8031 , \1451_b0 );
or ( \3501_b1 , \3496_b1 , \3500_b1 );
not ( \3500_b1 , w_8032 );
and ( \3501_b0 , \3496_b0 , w_8033 );
and ( w_8032 , w_8033 , \3500_b0 );
or ( \3502_b1 , \1517_b1 , \1349_b1 );
not ( \1349_b1 , w_8034 );
and ( \3502_b0 , \1517_b0 , w_8035 );
and ( w_8034 , w_8035 , \1349_b0 );
or ( \3503_b1 , \1526_b1 , \1347_b1 );
not ( \1347_b1 , w_8036 );
and ( \3503_b0 , \1526_b0 , w_8037 );
and ( w_8036 , w_8037 , \1347_b0 );
or ( \3504_b1 , \3502_b1 , w_8039 );
not ( w_8039 , w_8040 );
and ( \3504_b0 , \3502_b0 , w_8041 );
and ( w_8040 ,  , w_8041 );
buf ( w_8039 , \3503_b1 );
not ( w_8039 , w_8042 );
not (  , w_8043 );
and ( w_8042 , w_8043 , \3503_b0 );
or ( \3505_b1 , \3504_b1 , w_8044 );
xor ( \3505_b0 , \3504_b0 , w_8046 );
not ( w_8046 , w_8047 );
and ( w_8047 , w_8044 , w_8045 );
buf ( w_8044 , \1356_b1 );
not ( w_8044 , w_8048 );
not ( w_8045 , w_8049 );
and ( w_8048 , w_8049 , \1356_b0 );
or ( \3506_b1 , \3500_b1 , \3505_b1 );
not ( \3505_b1 , w_8050 );
and ( \3506_b0 , \3500_b0 , w_8051 );
and ( w_8050 , w_8051 , \3505_b0 );
or ( \3507_b1 , \3496_b1 , \3505_b1 );
not ( \3505_b1 , w_8052 );
and ( \3507_b0 , \3496_b0 , w_8053 );
and ( w_8052 , w_8053 , \3505_b0 );
or ( \3509_b1 , \1416_b1 , \1431_b1 );
not ( \1431_b1 , w_8054 );
and ( \3509_b0 , \1416_b0 , w_8055 );
and ( w_8054 , w_8055 , \1431_b0 );
or ( \3510_b1 , \1586_b1 , \1429_b1 );
not ( \1429_b1 , w_8056 );
and ( \3510_b0 , \1586_b0 , w_8057 );
and ( w_8056 , w_8057 , \1429_b0 );
or ( \3511_b1 , \3509_b1 , w_8059 );
not ( w_8059 , w_8060 );
and ( \3511_b0 , \3509_b0 , w_8061 );
and ( w_8060 ,  , w_8061 );
buf ( w_8059 , \3510_b1 );
not ( w_8059 , w_8062 );
not (  , w_8063 );
and ( w_8062 , w_8063 , \3510_b0 );
or ( \3512_b1 , \3511_b1 , w_8064 );
xor ( \3512_b0 , \3511_b0 , w_8066 );
not ( w_8066 , w_8067 );
and ( w_8067 , w_8064 , w_8065 );
buf ( w_8064 , \1438_b1 );
not ( w_8064 , w_8068 );
not ( w_8065 , w_8069 );
and ( w_8068 , w_8069 , \1438_b0 );
or ( \3513_b1 , \1498_b1 , \1458_b1 );
not ( \1458_b1 , w_8070 );
and ( \3513_b0 , \1498_b0 , w_8071 );
and ( w_8070 , w_8071 , \1458_b0 );
buf ( \3514_b1 , \3513_b1 );
not ( \3514_b1 , w_8072 );
not ( \3514_b0 , w_8073 );
and ( w_8072 , w_8073 , \3513_b0 );
or ( \3515_b1 , \3514_b1 , \1467_b1 );
not ( \1467_b1 , w_8074 );
and ( \3515_b0 , \3514_b0 , w_8075 );
and ( w_8074 , w_8075 , \1467_b0 );
or ( \3516_b1 , \3512_b1 , \3515_b1 );
not ( \3515_b1 , w_8076 );
and ( \3516_b0 , \3512_b0 , w_8077 );
and ( w_8076 , w_8077 , \3515_b0 );
or ( \3517_b1 , \3508_b1 , \3516_b1 );
not ( \3516_b1 , w_8078 );
and ( \3517_b0 , \3508_b0 , w_8079 );
and ( w_8078 , w_8079 , \3516_b0 );
or ( \3518_b1 , \1553_b1 , \1460_b1 );
not ( \1460_b1 , w_8080 );
and ( \3518_b0 , \1553_b0 , w_8081 );
and ( w_8080 , w_8081 , \1460_b0 );
or ( \3519_b1 , \1533_b1 , \1458_b1 );
not ( \1458_b1 , w_8082 );
and ( \3519_b0 , \1533_b0 , w_8083 );
and ( w_8082 , w_8083 , \1458_b0 );
or ( \3520_b1 , \3518_b1 , w_8085 );
not ( w_8085 , w_8086 );
and ( \3520_b0 , \3518_b0 , w_8087 );
and ( w_8086 ,  , w_8087 );
buf ( w_8085 , \3519_b1 );
not ( w_8085 , w_8088 );
not (  , w_8089 );
and ( w_8088 , w_8089 , \3519_b0 );
or ( \3521_b1 , \3520_b1 , w_8090 );
xor ( \3521_b0 , \3520_b0 , w_8092 );
not ( w_8092 , w_8093 );
and ( w_8093 , w_8090 , w_8091 );
buf ( w_8090 , \1467_b1 );
not ( w_8090 , w_8094 );
not ( w_8091 , w_8095 );
and ( w_8094 , w_8095 , \1467_b0 );
or ( \3522_b1 , \3516_b1 , \3521_b1 );
not ( \3521_b1 , w_8096 );
and ( \3522_b0 , \3516_b0 , w_8097 );
and ( w_8096 , w_8097 , \3521_b0 );
or ( \3523_b1 , \3508_b1 , \3521_b1 );
not ( \3521_b1 , w_8098 );
and ( \3523_b0 , \3508_b0 , w_8099 );
and ( w_8098 , w_8099 , \3521_b0 );
or ( \3525_b1 , \3387_b1 , \3391_b1 );
xor ( \3525_b0 , \3387_b0 , w_8100 );
not ( w_8100 , w_8101 );
and ( w_8101 , \3391_b1 , \3391_b0 );
or ( \3526_b1 , \3525_b1 , \3396_b1 );
xor ( \3526_b0 , \3525_b0 , w_8102 );
not ( w_8102 , w_8103 );
and ( w_8103 , \3396_b1 , \3396_b0 );
or ( \3527_b1 , \3524_b1 , \3526_b1 );
not ( \3526_b1 , w_8104 );
and ( \3527_b0 , \3524_b0 , w_8105 );
and ( w_8104 , w_8105 , \3526_b0 );
or ( \3528_b1 , \3403_b1 , \3407_b1 );
xor ( \3528_b0 , \3403_b0 , w_8106 );
not ( w_8106 , w_8107 );
and ( w_8107 , \3407_b1 , \3407_b0 );
or ( \3529_b1 , \3528_b1 , \3412_b1 );
xor ( \3529_b0 , \3528_b0 , w_8108 );
not ( w_8108 , w_8109 );
and ( w_8109 , \3412_b1 , \3412_b0 );
or ( \3530_b1 , \3526_b1 , \3529_b1 );
not ( \3529_b1 , w_8110 );
and ( \3530_b0 , \3526_b0 , w_8111 );
and ( w_8110 , w_8111 , \3529_b0 );
or ( \3531_b1 , \3524_b1 , \3529_b1 );
not ( \3529_b1 , w_8112 );
and ( \3531_b0 , \3524_b0 , w_8113 );
and ( w_8112 , w_8113 , \3529_b0 );
or ( \3533_b1 , \3399_b1 , \3415_b1 );
xor ( \3533_b0 , \3399_b0 , w_8114 );
not ( w_8114 , w_8115 );
and ( w_8115 , \3415_b1 , \3415_b0 );
or ( \3534_b1 , \3533_b1 , \3418_b1 );
xor ( \3534_b0 , \3533_b0 , w_8116 );
not ( w_8116 , w_8117 );
and ( w_8117 , \3418_b1 , \3418_b0 );
or ( \3535_b1 , \3532_b1 , \3534_b1 );
not ( \3534_b1 , w_8118 );
and ( \3535_b0 , \3532_b0 , w_8119 );
and ( w_8118 , w_8119 , \3534_b0 );
or ( \3536_b1 , \3472_b1 , \3474_b1 );
xor ( \3536_b0 , \3472_b0 , w_8120 );
not ( w_8120 , w_8121 );
and ( w_8121 , \3474_b1 , \3474_b0 );
or ( \3537_b1 , \3536_b1 , \3477_b1 );
xor ( \3537_b0 , \3536_b0 , w_8122 );
not ( w_8122 , w_8123 );
and ( w_8123 , \3477_b1 , \3477_b0 );
or ( \3538_b1 , \3534_b1 , \3537_b1 );
not ( \3537_b1 , w_8124 );
and ( \3538_b0 , \3534_b0 , w_8125 );
and ( w_8124 , w_8125 , \3537_b0 );
or ( \3539_b1 , \3532_b1 , \3537_b1 );
not ( \3537_b1 , w_8126 );
and ( \3539_b0 , \3532_b0 , w_8127 );
and ( w_8126 , w_8127 , \3537_b0 );
or ( \3541_b1 , \3492_b1 , \3540_b1 );
not ( \3540_b1 , w_8128 );
and ( \3541_b0 , \3492_b0 , w_8129 );
and ( w_8128 , w_8129 , \3540_b0 );
or ( \3542_b1 , \3492_b1 , \3540_b1 );
xor ( \3542_b0 , \3492_b0 , w_8130 );
not ( w_8130 , w_8131 );
and ( w_8131 , \3540_b1 , \3540_b0 );
or ( \3543_b1 , \3532_b1 , \3534_b1 );
xor ( \3543_b0 , \3532_b0 , w_8132 );
not ( w_8132 , w_8133 );
and ( w_8133 , \3534_b1 , \3534_b0 );
or ( \3544_b1 , \3543_b1 , \3537_b1 );
xor ( \3544_b0 , \3543_b0 , w_8134 );
not ( w_8134 , w_8135 );
and ( w_8135 , \3537_b1 , \3537_b0 );
or ( \3545_b1 , \3512_b1 , \3515_b1 );
xor ( \3545_b0 , \3512_b0 , w_8136 );
not ( w_8136 , w_8137 );
and ( w_8137 , \3515_b1 , \3515_b0 );
or ( \3546_b1 , \1533_b1 , \1382_b1 );
not ( \1382_b1 , w_8138 );
and ( \3546_b0 , \1533_b0 , w_8139 );
and ( w_8138 , w_8139 , \1382_b0 );
or ( \3547_b1 , \1540_b1 , \1380_b1 );
not ( \1380_b1 , w_8140 );
and ( \3547_b0 , \1540_b0 , w_8141 );
and ( w_8140 , w_8141 , \1380_b0 );
or ( \3548_b1 , \3546_b1 , w_8143 );
not ( w_8143 , w_8144 );
and ( \3548_b0 , \3546_b0 , w_8145 );
and ( w_8144 ,  , w_8145 );
buf ( w_8143 , \3547_b1 );
not ( w_8143 , w_8146 );
not (  , w_8147 );
and ( w_8146 , w_8147 , \3547_b0 );
or ( \3549_b1 , \3548_b1 , w_8148 );
xor ( \3549_b0 , \3548_b0 , w_8150 );
not ( w_8150 , w_8151 );
and ( w_8151 , w_8148 , w_8149 );
buf ( w_8148 , \1389_b1 );
not ( w_8148 , w_8152 );
not ( w_8149 , w_8153 );
and ( w_8152 , w_8153 , \1389_b0 );
or ( \3550_b1 , \3545_b1 , \3549_b1 );
not ( \3549_b1 , w_8154 );
and ( \3550_b0 , \3545_b0 , w_8155 );
and ( w_8154 , w_8155 , \3549_b0 );
or ( \3551_b1 , \1498_b1 , \1460_b1 );
not ( \1460_b1 , w_8156 );
and ( \3551_b0 , \1498_b0 , w_8157 );
and ( w_8156 , w_8157 , \1460_b0 );
or ( \3552_b1 , \1553_b1 , \1458_b1 );
not ( \1458_b1 , w_8158 );
and ( \3552_b0 , \1553_b0 , w_8159 );
and ( w_8158 , w_8159 , \1458_b0 );
or ( \3553_b1 , \3551_b1 , w_8161 );
not ( w_8161 , w_8162 );
and ( \3553_b0 , \3551_b0 , w_8163 );
and ( w_8162 ,  , w_8163 );
buf ( w_8161 , \3552_b1 );
not ( w_8161 , w_8164 );
not (  , w_8165 );
and ( w_8164 , w_8165 , \3552_b0 );
or ( \3554_b1 , \3553_b1 , w_8166 );
xor ( \3554_b0 , \3553_b0 , w_8168 );
not ( w_8168 , w_8169 );
and ( w_8169 , w_8166 , w_8167 );
buf ( w_8166 , \1467_b1 );
not ( w_8166 , w_8170 );
not ( w_8167 , w_8171 );
and ( w_8170 , w_8171 , \1467_b0 );
or ( \3555_b1 , \3549_b1 , \3554_b1 );
not ( \3554_b1 , w_8172 );
and ( \3555_b0 , \3549_b0 , w_8173 );
and ( w_8172 , w_8173 , \3554_b0 );
or ( \3556_b1 , \3545_b1 , \3554_b1 );
not ( \3554_b1 , w_8174 );
and ( \3556_b0 , \3545_b0 , w_8175 );
and ( w_8174 , w_8175 , \3554_b0 );
or ( \3558_b1 , \3444_b1 , \3448_b1 );
xor ( \3558_b0 , \3444_b0 , w_8176 );
not ( w_8176 , w_8177 );
and ( w_8177 , \3448_b1 , \3448_b0 );
or ( \3559_b1 , \3558_b1 , \3368_b1 );
xor ( \3559_b0 , \3558_b0 , w_8178 );
not ( w_8178 , w_8179 );
and ( w_8179 , \3368_b1 , \3368_b0 );
or ( \3560_b1 , \3557_b1 , \3559_b1 );
not ( \3559_b1 , w_8180 );
and ( \3560_b0 , \3557_b0 , w_8181 );
and ( w_8180 , w_8181 , \3559_b0 );
or ( \3561_b1 , \3457_b1 , \3461_b1 );
xor ( \3561_b0 , \3457_b0 , w_8182 );
not ( w_8182 , w_8183 );
and ( w_8183 , \3461_b1 , \3461_b0 );
or ( \3562_b1 , \3561_b1 , \3466_b1 );
xor ( \3562_b0 , \3561_b0 , w_8184 );
not ( w_8184 , w_8185 );
and ( w_8185 , \3466_b1 , \3466_b0 );
or ( \3563_b1 , \3559_b1 , \3562_b1 );
not ( \3562_b1 , w_8186 );
and ( \3563_b0 , \3559_b0 , w_8187 );
and ( w_8186 , w_8187 , \3562_b0 );
or ( \3564_b1 , \3557_b1 , \3562_b1 );
not ( \3562_b1 , w_8188 );
and ( \3564_b0 , \3557_b0 , w_8189 );
and ( w_8188 , w_8189 , \3562_b0 );
or ( \3566_b1 , \3440_b1 , \3452_b1 );
xor ( \3566_b0 , \3440_b0 , w_8190 );
not ( w_8190 , w_8191 );
and ( w_8191 , \3452_b1 , \3452_b0 );
or ( \3567_b1 , \3566_b1 , \3469_b1 );
xor ( \3567_b0 , \3566_b0 , w_8192 );
not ( w_8192 , w_8193 );
and ( w_8193 , \3469_b1 , \3469_b0 );
or ( \3568_b1 , \3565_b1 , \3567_b1 );
not ( \3567_b1 , w_8194 );
and ( \3568_b0 , \3565_b0 , w_8195 );
and ( w_8194 , w_8195 , \3567_b0 );
or ( \3569_b1 , \3524_b1 , \3526_b1 );
xor ( \3569_b0 , \3524_b0 , w_8196 );
not ( w_8196 , w_8197 );
and ( w_8197 , \3526_b1 , \3526_b0 );
or ( \3570_b1 , \3569_b1 , \3529_b1 );
xor ( \3570_b0 , \3569_b0 , w_8198 );
not ( w_8198 , w_8199 );
and ( w_8199 , \3529_b1 , \3529_b0 );
or ( \3571_b1 , \3567_b1 , \3570_b1 );
not ( \3570_b1 , w_8200 );
and ( \3571_b0 , \3567_b0 , w_8201 );
and ( w_8200 , w_8201 , \3570_b0 );
or ( \3572_b1 , \3565_b1 , \3570_b1 );
not ( \3570_b1 , w_8202 );
and ( \3572_b0 , \3565_b0 , w_8203 );
and ( w_8202 , w_8203 , \3570_b0 );
or ( \3574_b1 , \3544_b1 , \3573_b1 );
not ( \3573_b1 , w_8204 );
and ( \3574_b0 , \3544_b0 , w_8205 );
and ( w_8204 , w_8205 , \3573_b0 );
or ( \3575_b1 , \3544_b1 , \3573_b1 );
xor ( \3575_b0 , \3544_b0 , w_8206 );
not ( w_8206 , w_8207 );
and ( w_8207 , \3573_b1 , \3573_b0 );
or ( \3576_b1 , \3565_b1 , \3567_b1 );
xor ( \3576_b0 , \3565_b0 , w_8208 );
not ( w_8208 , w_8209 );
and ( w_8209 , \3567_b1 , \3567_b0 );
or ( \3577_b1 , \3576_b1 , \3570_b1 );
xor ( \3577_b0 , \3576_b0 , w_8210 );
not ( w_8210 , w_8211 );
and ( w_8211 , \3570_b1 , \3570_b0 );
or ( \3578_b1 , \1407_b1 , \1431_b1 );
not ( \1431_b1 , w_8212 );
and ( \3578_b0 , \1407_b0 , w_8213 );
and ( w_8212 , w_8213 , \1431_b0 );
or ( \3579_b1 , \1416_b1 , \1429_b1 );
not ( \1429_b1 , w_8214 );
and ( \3579_b0 , \1416_b0 , w_8215 );
and ( w_8214 , w_8215 , \1429_b0 );
or ( \3580_b1 , \3578_b1 , w_8217 );
not ( w_8217 , w_8218 );
and ( \3580_b0 , \3578_b0 , w_8219 );
and ( w_8218 ,  , w_8219 );
buf ( w_8217 , \3579_b1 );
not ( w_8217 , w_8220 );
not (  , w_8221 );
and ( w_8220 , w_8221 , \3579_b0 );
or ( \3581_b1 , \3580_b1 , w_8222 );
xor ( \3581_b0 , \3580_b0 , w_8224 );
not ( w_8224 , w_8225 );
and ( w_8225 , w_8222 , w_8223 );
buf ( w_8222 , \1438_b1 );
not ( w_8222 , w_8226 );
not ( w_8223 , w_8227 );
and ( w_8226 , w_8227 , \1438_b0 );
or ( \3582_b1 , \1526_b1 , \1444_b1 );
not ( \1444_b1 , w_8228 );
and ( \3582_b0 , \1526_b0 , w_8229 );
and ( w_8228 , w_8229 , \1444_b0 );
or ( \3583_b1 , \1622_b1 , \1442_b1 );
not ( \1442_b1 , w_8230 );
and ( \3583_b0 , \1622_b0 , w_8231 );
and ( w_8230 , w_8231 , \1442_b0 );
or ( \3584_b1 , \3582_b1 , w_8233 );
not ( w_8233 , w_8234 );
and ( \3584_b0 , \3582_b0 , w_8235 );
and ( w_8234 ,  , w_8235 );
buf ( w_8233 , \3583_b1 );
not ( w_8233 , w_8236 );
not (  , w_8237 );
and ( w_8236 , w_8237 , \3583_b0 );
or ( \3585_b1 , \3584_b1 , w_8238 );
xor ( \3585_b0 , \3584_b0 , w_8240 );
not ( w_8240 , w_8241 );
and ( w_8241 , w_8238 , w_8239 );
buf ( w_8238 , \1451_b1 );
not ( w_8238 , w_8242 );
not ( w_8239 , w_8243 );
and ( w_8242 , w_8243 , \1451_b0 );
or ( \3586_b1 , \3581_b1 , \3585_b1 );
not ( \3585_b1 , w_8244 );
and ( \3586_b0 , \3581_b0 , w_8245 );
and ( w_8244 , w_8245 , \3585_b0 );
or ( \3587_b1 , \3585_b1 , \3513_b1 );
not ( \3513_b1 , w_8246 );
and ( \3587_b0 , \3585_b0 , w_8247 );
and ( w_8246 , w_8247 , \3513_b0 );
or ( \3588_b1 , \3581_b1 , \3513_b1 );
not ( \3513_b1 , w_8248 );
and ( \3588_b0 , \3581_b0 , w_8249 );
and ( w_8248 , w_8249 , \3513_b0 );
or ( \3590_b1 , \1586_b1 , \1336_b1 );
not ( \1336_b1 , w_8250 );
and ( \3590_b0 , \1586_b0 , w_8251 );
and ( w_8250 , w_8251 , \1336_b0 );
or ( \3591_b1 , \1616_b1 , \1333_b1 );
not ( \1333_b1 , w_8252 );
and ( \3591_b0 , \1616_b0 , w_8253 );
and ( w_8252 , w_8253 , \1333_b0 );
or ( \3592_b1 , \3590_b1 , w_8255 );
not ( w_8255 , w_8256 );
and ( \3592_b0 , \3590_b0 , w_8257 );
and ( w_8256 ,  , w_8257 );
buf ( w_8255 , \3591_b1 );
not ( w_8255 , w_8258 );
not (  , w_8259 );
and ( w_8258 , w_8259 , \3591_b0 );
or ( \3593_b1 , \3592_b1 , w_8260 );
xor ( \3593_b0 , \3592_b0 , w_8262 );
not ( w_8262 , w_8263 );
and ( w_8263 , w_8260 , w_8261 );
buf ( w_8260 , \1332_b1 );
not ( w_8260 , w_8264 );
not ( w_8261 , w_8265 );
and ( w_8264 , w_8265 , \1332_b0 );
or ( \3594_b1 , \1540_b1 , \1349_b1 );
not ( \1349_b1 , w_8266 );
and ( \3594_b0 , \1540_b0 , w_8267 );
and ( w_8266 , w_8267 , \1349_b0 );
or ( \3595_b1 , \1517_b1 , \1347_b1 );
not ( \1347_b1 , w_8268 );
and ( \3595_b0 , \1517_b0 , w_8269 );
and ( w_8268 , w_8269 , \1347_b0 );
or ( \3596_b1 , \3594_b1 , w_8271 );
not ( w_8271 , w_8272 );
and ( \3596_b0 , \3594_b0 , w_8273 );
and ( w_8272 ,  , w_8273 );
buf ( w_8271 , \3595_b1 );
not ( w_8271 , w_8274 );
not (  , w_8275 );
and ( w_8274 , w_8275 , \3595_b0 );
or ( \3597_b1 , \3596_b1 , w_8276 );
xor ( \3597_b0 , \3596_b0 , w_8278 );
not ( w_8278 , w_8279 );
and ( w_8279 , w_8276 , w_8277 );
buf ( w_8276 , \1356_b1 );
not ( w_8276 , w_8280 );
not ( w_8277 , w_8281 );
and ( w_8280 , w_8281 , \1356_b0 );
or ( \3598_b1 , \3593_b1 , \3597_b1 );
not ( \3597_b1 , w_8282 );
and ( \3598_b0 , \3593_b0 , w_8283 );
and ( w_8282 , w_8283 , \3597_b0 );
or ( \3599_b1 , \1553_b1 , \1382_b1 );
not ( \1382_b1 , w_8284 );
and ( \3599_b0 , \1553_b0 , w_8285 );
and ( w_8284 , w_8285 , \1382_b0 );
or ( \3600_b1 , \1533_b1 , \1380_b1 );
not ( \1380_b1 , w_8286 );
and ( \3600_b0 , \1533_b0 , w_8287 );
and ( w_8286 , w_8287 , \1380_b0 );
or ( \3601_b1 , \3599_b1 , w_8289 );
not ( w_8289 , w_8290 );
and ( \3601_b0 , \3599_b0 , w_8291 );
and ( w_8290 ,  , w_8291 );
buf ( w_8289 , \3600_b1 );
not ( w_8289 , w_8292 );
not (  , w_8293 );
and ( w_8292 , w_8293 , \3600_b0 );
or ( \3602_b1 , \3601_b1 , w_8294 );
xor ( \3602_b0 , \3601_b0 , w_8296 );
not ( w_8296 , w_8297 );
and ( w_8297 , w_8294 , w_8295 );
buf ( w_8294 , \1389_b1 );
not ( w_8294 , w_8298 );
not ( w_8295 , w_8299 );
and ( w_8298 , w_8299 , \1389_b0 );
or ( \3603_b1 , \3597_b1 , \3602_b1 );
not ( \3602_b1 , w_8300 );
and ( \3603_b0 , \3597_b0 , w_8301 );
and ( w_8300 , w_8301 , \3602_b0 );
or ( \3604_b1 , \3593_b1 , \3602_b1 );
not ( \3602_b1 , w_8302 );
and ( \3604_b0 , \3593_b0 , w_8303 );
and ( w_8302 , w_8303 , \3602_b0 );
or ( \3606_b1 , \3589_b1 , \3605_b1 );
not ( \3605_b1 , w_8304 );
and ( \3606_b0 , \3589_b0 , w_8305 );
and ( w_8304 , w_8305 , \3605_b0 );
or ( \3607_b1 , \3545_b1 , \3549_b1 );
xor ( \3607_b0 , \3545_b0 , w_8306 );
not ( w_8306 , w_8307 );
and ( w_8307 , \3549_b1 , \3549_b0 );
or ( \3608_b1 , \3607_b1 , \3554_b1 );
xor ( \3608_b0 , \3607_b0 , w_8308 );
not ( w_8308 , w_8309 );
and ( w_8309 , \3554_b1 , \3554_b0 );
or ( \3609_b1 , \3605_b1 , \3608_b1 );
not ( \3608_b1 , w_8310 );
and ( \3609_b0 , \3605_b0 , w_8311 );
and ( w_8310 , w_8311 , \3608_b0 );
or ( \3610_b1 , \3589_b1 , \3608_b1 );
not ( \3608_b1 , w_8312 );
and ( \3610_b0 , \3589_b0 , w_8313 );
and ( w_8312 , w_8313 , \3608_b0 );
or ( \3612_b1 , \3508_b1 , \3516_b1 );
xor ( \3612_b0 , \3508_b0 , w_8314 );
not ( w_8314 , w_8315 );
and ( w_8315 , \3516_b1 , \3516_b0 );
or ( \3613_b1 , \3612_b1 , \3521_b1 );
xor ( \3613_b0 , \3612_b0 , w_8316 );
not ( w_8316 , w_8317 );
and ( w_8317 , \3521_b1 , \3521_b0 );
or ( \3614_b1 , \3611_b1 , \3613_b1 );
not ( \3613_b1 , w_8318 );
and ( \3614_b0 , \3611_b0 , w_8319 );
and ( w_8318 , w_8319 , \3613_b0 );
or ( \3615_b1 , \3557_b1 , \3559_b1 );
xor ( \3615_b0 , \3557_b0 , w_8320 );
not ( w_8320 , w_8321 );
and ( w_8321 , \3559_b1 , \3559_b0 );
or ( \3616_b1 , \3615_b1 , \3562_b1 );
xor ( \3616_b0 , \3615_b0 , w_8322 );
not ( w_8322 , w_8323 );
and ( w_8323 , \3562_b1 , \3562_b0 );
or ( \3617_b1 , \3613_b1 , \3616_b1 );
not ( \3616_b1 , w_8324 );
and ( \3617_b0 , \3613_b0 , w_8325 );
and ( w_8324 , w_8325 , \3616_b0 );
or ( \3618_b1 , \3611_b1 , \3616_b1 );
not ( \3616_b1 , w_8326 );
and ( \3618_b0 , \3611_b0 , w_8327 );
and ( w_8326 , w_8327 , \3616_b0 );
or ( \3620_b1 , \3577_b1 , \3619_b1 );
not ( \3619_b1 , w_8328 );
and ( \3620_b0 , \3577_b0 , w_8329 );
and ( w_8328 , w_8329 , \3619_b0 );
or ( \3621_b1 , \3577_b1 , \3619_b1 );
xor ( \3621_b0 , \3577_b0 , w_8330 );
not ( w_8330 , w_8331 );
and ( w_8331 , \3619_b1 , \3619_b0 );
or ( \3622_b1 , \3611_b1 , \3613_b1 );
xor ( \3622_b0 , \3611_b0 , w_8332 );
not ( w_8332 , w_8333 );
and ( w_8333 , \3613_b1 , \3613_b0 );
or ( \3623_b1 , \3622_b1 , \3616_b1 );
xor ( \3623_b0 , \3622_b0 , w_8334 );
not ( w_8334 , w_8335 );
and ( w_8335 , \3616_b1 , \3616_b0 );
or ( \3624_b1 , \1416_b1 , \1336_b1 );
not ( \1336_b1 , w_8336 );
and ( \3624_b0 , \1416_b0 , w_8337 );
and ( w_8336 , w_8337 , \1336_b0 );
or ( \3625_b1 , \1586_b1 , \1333_b1 );
not ( \1333_b1 , w_8338 );
and ( \3625_b0 , \1586_b0 , w_8339 );
and ( w_8338 , w_8339 , \1333_b0 );
or ( \3626_b1 , \3624_b1 , w_8341 );
not ( w_8341 , w_8342 );
and ( \3626_b0 , \3624_b0 , w_8343 );
and ( w_8342 ,  , w_8343 );
buf ( w_8341 , \3625_b1 );
not ( w_8341 , w_8344 );
not (  , w_8345 );
and ( w_8344 , w_8345 , \3625_b0 );
or ( \3627_b1 , \3626_b1 , w_8346 );
xor ( \3627_b0 , \3626_b0 , w_8348 );
not ( w_8348 , w_8349 );
and ( w_8349 , w_8346 , w_8347 );
buf ( w_8346 , \1332_b1 );
not ( w_8346 , w_8350 );
not ( w_8347 , w_8351 );
and ( w_8350 , w_8351 , \1332_b0 );
or ( \3628_b1 , \1517_b1 , \1444_b1 );
not ( \1444_b1 , w_8352 );
and ( \3628_b0 , \1517_b0 , w_8353 );
and ( w_8352 , w_8353 , \1444_b0 );
or ( \3629_b1 , \1526_b1 , \1442_b1 );
not ( \1442_b1 , w_8354 );
and ( \3629_b0 , \1526_b0 , w_8355 );
and ( w_8354 , w_8355 , \1442_b0 );
or ( \3630_b1 , \3628_b1 , w_8357 );
not ( w_8357 , w_8358 );
and ( \3630_b0 , \3628_b0 , w_8359 );
and ( w_8358 ,  , w_8359 );
buf ( w_8357 , \3629_b1 );
not ( w_8357 , w_8360 );
not (  , w_8361 );
and ( w_8360 , w_8361 , \3629_b0 );
or ( \3631_b1 , \3630_b1 , w_8362 );
xor ( \3631_b0 , \3630_b0 , w_8364 );
not ( w_8364 , w_8365 );
and ( w_8365 , w_8362 , w_8363 );
buf ( w_8362 , \1451_b1 );
not ( w_8362 , w_8366 );
not ( w_8363 , w_8367 );
and ( w_8366 , w_8367 , \1451_b0 );
or ( \3632_b1 , \3627_b1 , \3631_b1 );
not ( \3631_b1 , w_8368 );
and ( \3632_b0 , \3627_b0 , w_8369 );
and ( w_8368 , w_8369 , \3631_b0 );
or ( \3633_b1 , \1533_b1 , \1349_b1 );
not ( \1349_b1 , w_8370 );
and ( \3633_b0 , \1533_b0 , w_8371 );
and ( w_8370 , w_8371 , \1349_b0 );
or ( \3634_b1 , \1540_b1 , \1347_b1 );
not ( \1347_b1 , w_8372 );
and ( \3634_b0 , \1540_b0 , w_8373 );
and ( w_8372 , w_8373 , \1347_b0 );
or ( \3635_b1 , \3633_b1 , w_8375 );
not ( w_8375 , w_8376 );
and ( \3635_b0 , \3633_b0 , w_8377 );
and ( w_8376 ,  , w_8377 );
buf ( w_8375 , \3634_b1 );
not ( w_8375 , w_8378 );
not (  , w_8379 );
and ( w_8378 , w_8379 , \3634_b0 );
or ( \3636_b1 , \3635_b1 , w_8380 );
xor ( \3636_b0 , \3635_b0 , w_8382 );
not ( w_8382 , w_8383 );
and ( w_8383 , w_8380 , w_8381 );
buf ( w_8380 , \1356_b1 );
not ( w_8380 , w_8384 );
not ( w_8381 , w_8385 );
and ( w_8384 , w_8385 , \1356_b0 );
or ( \3637_b1 , \3631_b1 , \3636_b1 );
not ( \3636_b1 , w_8386 );
and ( \3637_b0 , \3631_b0 , w_8387 );
and ( w_8386 , w_8387 , \3636_b0 );
or ( \3638_b1 , \3627_b1 , \3636_b1 );
not ( \3636_b1 , w_8388 );
and ( \3638_b0 , \3627_b0 , w_8389 );
and ( w_8388 , w_8389 , \3636_b0 );
or ( \3640_b1 , \1622_b1 , \1431_b1 );
not ( \1431_b1 , w_8390 );
and ( \3640_b0 , \1622_b0 , w_8391 );
and ( w_8390 , w_8391 , \1431_b0 );
or ( \3641_b1 , \1407_b1 , \1429_b1 );
not ( \1429_b1 , w_8392 );
and ( \3641_b0 , \1407_b0 , w_8393 );
and ( w_8392 , w_8393 , \1429_b0 );
or ( \3642_b1 , \3640_b1 , w_8395 );
not ( w_8395 , w_8396 );
and ( \3642_b0 , \3640_b0 , w_8397 );
and ( w_8396 ,  , w_8397 );
buf ( w_8395 , \3641_b1 );
not ( w_8395 , w_8398 );
not (  , w_8399 );
and ( w_8398 , w_8399 , \3641_b0 );
or ( \3643_b1 , \3642_b1 , w_8400 );
xor ( \3643_b0 , \3642_b0 , w_8402 );
not ( w_8402 , w_8403 );
and ( w_8403 , w_8400 , w_8401 );
buf ( w_8400 , \1438_b1 );
not ( w_8400 , w_8404 );
not ( w_8401 , w_8405 );
and ( w_8404 , w_8405 , \1438_b0 );
or ( \3644_b1 , \1498_b1 , \1380_b1 );
not ( \1380_b1 , w_8406 );
and ( \3644_b0 , \1498_b0 , w_8407 );
and ( w_8406 , w_8407 , \1380_b0 );
buf ( \3645_b1 , \3644_b1 );
not ( \3645_b1 , w_8408 );
not ( \3645_b0 , w_8409 );
and ( w_8408 , w_8409 , \3644_b0 );
or ( \3646_b1 , \3645_b1 , \1389_b1 );
not ( \1389_b1 , w_8410 );
and ( \3646_b0 , \3645_b0 , w_8411 );
and ( w_8410 , w_8411 , \1389_b0 );
or ( \3647_b1 , \3643_b1 , \3646_b1 );
not ( \3646_b1 , w_8412 );
and ( \3647_b0 , \3643_b0 , w_8413 );
and ( w_8412 , w_8413 , \3646_b0 );
or ( \3648_b1 , \3639_b1 , \3647_b1 );
not ( \3647_b1 , w_8414 );
and ( \3648_b0 , \3639_b0 , w_8415 );
and ( w_8414 , w_8415 , \3647_b0 );
or ( \3649_b1 , \3581_b1 , \3585_b1 );
xor ( \3649_b0 , \3581_b0 , w_8416 );
not ( w_8416 , w_8417 );
and ( w_8417 , \3585_b1 , \3585_b0 );
or ( \3650_b1 , \3649_b1 , \3513_b1 );
xor ( \3650_b0 , \3649_b0 , w_8418 );
not ( w_8418 , w_8419 );
and ( w_8419 , \3513_b1 , \3513_b0 );
or ( \3651_b1 , \3647_b1 , \3650_b1 );
not ( \3650_b1 , w_8420 );
and ( \3651_b0 , \3647_b0 , w_8421 );
and ( w_8420 , w_8421 , \3650_b0 );
or ( \3652_b1 , \3639_b1 , \3650_b1 );
not ( \3650_b1 , w_8422 );
and ( \3652_b0 , \3639_b0 , w_8423 );
and ( w_8422 , w_8423 , \3650_b0 );
or ( \3654_b1 , \3496_b1 , \3500_b1 );
xor ( \3654_b0 , \3496_b0 , w_8424 );
not ( w_8424 , w_8425 );
and ( w_8425 , \3500_b1 , \3500_b0 );
or ( \3655_b1 , \3654_b1 , \3505_b1 );
xor ( \3655_b0 , \3654_b0 , w_8426 );
not ( w_8426 , w_8427 );
and ( w_8427 , \3505_b1 , \3505_b0 );
or ( \3656_b1 , \3653_b1 , \3655_b1 );
not ( \3655_b1 , w_8428 );
and ( \3656_b0 , \3653_b0 , w_8429 );
and ( w_8428 , w_8429 , \3655_b0 );
or ( \3657_b1 , \3589_b1 , \3605_b1 );
xor ( \3657_b0 , \3589_b0 , w_8430 );
not ( w_8430 , w_8431 );
and ( w_8431 , \3605_b1 , \3605_b0 );
or ( \3658_b1 , \3657_b1 , \3608_b1 );
xor ( \3658_b0 , \3657_b0 , w_8432 );
not ( w_8432 , w_8433 );
and ( w_8433 , \3608_b1 , \3608_b0 );
or ( \3659_b1 , \3655_b1 , \3658_b1 );
not ( \3658_b1 , w_8434 );
and ( \3659_b0 , \3655_b0 , w_8435 );
and ( w_8434 , w_8435 , \3658_b0 );
or ( \3660_b1 , \3653_b1 , \3658_b1 );
not ( \3658_b1 , w_8436 );
and ( \3660_b0 , \3653_b0 , w_8437 );
and ( w_8436 , w_8437 , \3658_b0 );
or ( \3662_b1 , \3623_b1 , \3661_b1 );
not ( \3661_b1 , w_8438 );
and ( \3662_b0 , \3623_b0 , w_8439 );
and ( w_8438 , w_8439 , \3661_b0 );
or ( \3663_b1 , \3623_b1 , \3661_b1 );
xor ( \3663_b0 , \3623_b0 , w_8440 );
not ( w_8440 , w_8441 );
and ( w_8441 , \3661_b1 , \3661_b0 );
or ( \3664_b1 , \3643_b1 , \3646_b1 );
xor ( \3664_b0 , \3643_b0 , w_8442 );
not ( w_8442 , w_8443 );
and ( w_8443 , \3646_b1 , \3646_b0 );
or ( \3665_b1 , \1526_b1 , \1431_b1 );
not ( \1431_b1 , w_8444 );
and ( \3665_b0 , \1526_b0 , w_8445 );
and ( w_8444 , w_8445 , \1431_b0 );
or ( \3666_b1 , \1622_b1 , \1429_b1 );
not ( \1429_b1 , w_8446 );
and ( \3666_b0 , \1622_b0 , w_8447 );
and ( w_8446 , w_8447 , \1429_b0 );
or ( \3667_b1 , \3665_b1 , w_8449 );
not ( w_8449 , w_8450 );
and ( \3667_b0 , \3665_b0 , w_8451 );
and ( w_8450 ,  , w_8451 );
buf ( w_8449 , \3666_b1 );
not ( w_8449 , w_8452 );
not (  , w_8453 );
and ( w_8452 , w_8453 , \3666_b0 );
or ( \3668_b1 , \3667_b1 , w_8454 );
xor ( \3668_b0 , \3667_b0 , w_8456 );
not ( w_8456 , w_8457 );
and ( w_8457 , w_8454 , w_8455 );
buf ( w_8454 , \1438_b1 );
not ( w_8454 , w_8458 );
not ( w_8455 , w_8459 );
and ( w_8458 , w_8459 , \1438_b0 );
or ( \3669_b1 , \1540_b1 , \1444_b1 );
not ( \1444_b1 , w_8460 );
and ( \3669_b0 , \1540_b0 , w_8461 );
and ( w_8460 , w_8461 , \1444_b0 );
or ( \3670_b1 , \1517_b1 , \1442_b1 );
not ( \1442_b1 , w_8462 );
and ( \3670_b0 , \1517_b0 , w_8463 );
and ( w_8462 , w_8463 , \1442_b0 );
or ( \3671_b1 , \3669_b1 , w_8465 );
not ( w_8465 , w_8466 );
and ( \3671_b0 , \3669_b0 , w_8467 );
and ( w_8466 ,  , w_8467 );
buf ( w_8465 , \3670_b1 );
not ( w_8465 , w_8468 );
not (  , w_8469 );
and ( w_8468 , w_8469 , \3670_b0 );
or ( \3672_b1 , \3671_b1 , w_8470 );
xor ( \3672_b0 , \3671_b0 , w_8472 );
not ( w_8472 , w_8473 );
and ( w_8473 , w_8470 , w_8471 );
buf ( w_8470 , \1451_b1 );
not ( w_8470 , w_8474 );
not ( w_8471 , w_8475 );
and ( w_8474 , w_8475 , \1451_b0 );
or ( \3673_b1 , \3668_b1 , \3672_b1 );
not ( \3672_b1 , w_8476 );
and ( \3673_b0 , \3668_b0 , w_8477 );
and ( w_8476 , w_8477 , \3672_b0 );
or ( \3674_b1 , \3672_b1 , \3644_b1 );
not ( \3644_b1 , w_8478 );
and ( \3674_b0 , \3672_b0 , w_8479 );
and ( w_8478 , w_8479 , \3644_b0 );
or ( \3675_b1 , \3668_b1 , \3644_b1 );
not ( \3644_b1 , w_8480 );
and ( \3675_b0 , \3668_b0 , w_8481 );
and ( w_8480 , w_8481 , \3644_b0 );
or ( \3677_b1 , \3664_b1 , \3676_b1 );
not ( \3676_b1 , w_8482 );
and ( \3677_b0 , \3664_b0 , w_8483 );
and ( w_8482 , w_8483 , \3676_b0 );
or ( \3678_b1 , \1498_b1 , \1382_b1 );
not ( \1382_b1 , w_8484 );
and ( \3678_b0 , \1498_b0 , w_8485 );
and ( w_8484 , w_8485 , \1382_b0 );
or ( \3679_b1 , \1553_b1 , \1380_b1 );
not ( \1380_b1 , w_8486 );
and ( \3679_b0 , \1553_b0 , w_8487 );
and ( w_8486 , w_8487 , \1380_b0 );
or ( \3680_b1 , \3678_b1 , w_8489 );
not ( w_8489 , w_8490 );
and ( \3680_b0 , \3678_b0 , w_8491 );
and ( w_8490 ,  , w_8491 );
buf ( w_8489 , \3679_b1 );
not ( w_8489 , w_8492 );
not (  , w_8493 );
and ( w_8492 , w_8493 , \3679_b0 );
or ( \3681_b1 , \3680_b1 , w_8494 );
xor ( \3681_b0 , \3680_b0 , w_8496 );
not ( w_8496 , w_8497 );
and ( w_8497 , w_8494 , w_8495 );
buf ( w_8494 , \1389_b1 );
not ( w_8494 , w_8498 );
not ( w_8495 , w_8499 );
and ( w_8498 , w_8499 , \1389_b0 );
or ( \3682_b1 , \3676_b1 , \3681_b1 );
not ( \3681_b1 , w_8500 );
and ( \3682_b0 , \3676_b0 , w_8501 );
and ( w_8500 , w_8501 , \3681_b0 );
or ( \3683_b1 , \3664_b1 , \3681_b1 );
not ( \3681_b1 , w_8502 );
and ( \3683_b0 , \3664_b0 , w_8503 );
and ( w_8502 , w_8503 , \3681_b0 );
or ( \3685_b1 , \3593_b1 , \3597_b1 );
xor ( \3685_b0 , \3593_b0 , w_8504 );
not ( w_8504 , w_8505 );
and ( w_8505 , \3597_b1 , \3597_b0 );
or ( \3686_b1 , \3685_b1 , \3602_b1 );
xor ( \3686_b0 , \3685_b0 , w_8506 );
not ( w_8506 , w_8507 );
and ( w_8507 , \3602_b1 , \3602_b0 );
or ( \3687_b1 , \3684_b1 , \3686_b1 );
not ( \3686_b1 , w_8508 );
and ( \3687_b0 , \3684_b0 , w_8509 );
and ( w_8508 , w_8509 , \3686_b0 );
or ( \3688_b1 , \3639_b1 , \3647_b1 );
xor ( \3688_b0 , \3639_b0 , w_8510 );
not ( w_8510 , w_8511 );
and ( w_8511 , \3647_b1 , \3647_b0 );
or ( \3689_b1 , \3688_b1 , \3650_b1 );
xor ( \3689_b0 , \3688_b0 , w_8512 );
not ( w_8512 , w_8513 );
and ( w_8513 , \3650_b1 , \3650_b0 );
or ( \3690_b1 , \3686_b1 , \3689_b1 );
not ( \3689_b1 , w_8514 );
and ( \3690_b0 , \3686_b0 , w_8515 );
and ( w_8514 , w_8515 , \3689_b0 );
or ( \3691_b1 , \3684_b1 , \3689_b1 );
not ( \3689_b1 , w_8516 );
and ( \3691_b0 , \3684_b0 , w_8517 );
and ( w_8516 , w_8517 , \3689_b0 );
or ( \3693_b1 , \3653_b1 , \3655_b1 );
xor ( \3693_b0 , \3653_b0 , w_8518 );
not ( w_8518 , w_8519 );
and ( w_8519 , \3655_b1 , \3655_b0 );
or ( \3694_b1 , \3693_b1 , \3658_b1 );
xor ( \3694_b0 , \3693_b0 , w_8520 );
not ( w_8520 , w_8521 );
and ( w_8521 , \3658_b1 , \3658_b0 );
or ( \3695_b1 , \3692_b1 , \3694_b1 );
not ( \3694_b1 , w_8522 );
and ( \3695_b0 , \3692_b0 , w_8523 );
and ( w_8522 , w_8523 , \3694_b0 );
or ( \3696_b1 , \3692_b1 , \3694_b1 );
xor ( \3696_b0 , \3692_b0 , w_8524 );
not ( w_8524 , w_8525 );
and ( w_8525 , \3694_b1 , \3694_b0 );
or ( \3697_b1 , \3684_b1 , \3686_b1 );
xor ( \3697_b0 , \3684_b0 , w_8526 );
not ( w_8526 , w_8527 );
and ( w_8527 , \3686_b1 , \3686_b0 );
or ( \3698_b1 , \3697_b1 , \3689_b1 );
xor ( \3698_b0 , \3697_b0 , w_8528 );
not ( w_8528 , w_8529 );
and ( w_8529 , \3689_b1 , \3689_b0 );
or ( \3699_b1 , \1517_b1 , \1431_b1 );
not ( \1431_b1 , w_8530 );
and ( \3699_b0 , \1517_b0 , w_8531 );
and ( w_8530 , w_8531 , \1431_b0 );
or ( \3700_b1 , \1526_b1 , \1429_b1 );
not ( \1429_b1 , w_8532 );
and ( \3700_b0 , \1526_b0 , w_8533 );
and ( w_8532 , w_8533 , \1429_b0 );
or ( \3701_b1 , \3699_b1 , w_8535 );
not ( w_8535 , w_8536 );
and ( \3701_b0 , \3699_b0 , w_8537 );
and ( w_8536 ,  , w_8537 );
buf ( w_8535 , \3700_b1 );
not ( w_8535 , w_8538 );
not (  , w_8539 );
and ( w_8538 , w_8539 , \3700_b0 );
or ( \3702_b1 , \3701_b1 , w_8540 );
xor ( \3702_b0 , \3701_b0 , w_8542 );
not ( w_8542 , w_8543 );
and ( w_8543 , w_8540 , w_8541 );
buf ( w_8540 , \1438_b1 );
not ( w_8540 , w_8544 );
not ( w_8541 , w_8545 );
and ( w_8544 , w_8545 , \1438_b0 );
or ( \3703_b1 , \1498_b1 , \1347_b1 );
not ( \1347_b1 , w_8546 );
and ( \3703_b0 , \1498_b0 , w_8547 );
and ( w_8546 , w_8547 , \1347_b0 );
buf ( \3704_b1 , \3703_b1 );
not ( \3704_b1 , w_8548 );
not ( \3704_b0 , w_8549 );
and ( w_8548 , w_8549 , \3703_b0 );
or ( \3705_b1 , \3704_b1 , \1356_b1 );
not ( \1356_b1 , w_8550 );
and ( \3705_b0 , \3704_b0 , w_8551 );
and ( w_8550 , w_8551 , \1356_b0 );
or ( \3706_b1 , \3702_b1 , \3705_b1 );
not ( \3705_b1 , w_8552 );
and ( \3706_b0 , \3702_b0 , w_8553 );
and ( w_8552 , w_8553 , \3705_b0 );
or ( \3707_b1 , \1407_b1 , \1336_b1 );
not ( \1336_b1 , w_8554 );
and ( \3707_b0 , \1407_b0 , w_8555 );
and ( w_8554 , w_8555 , \1336_b0 );
or ( \3708_b1 , \1416_b1 , \1333_b1 );
not ( \1333_b1 , w_8556 );
and ( \3708_b0 , \1416_b0 , w_8557 );
and ( w_8556 , w_8557 , \1333_b0 );
or ( \3709_b1 , \3707_b1 , w_8559 );
not ( w_8559 , w_8560 );
and ( \3709_b0 , \3707_b0 , w_8561 );
and ( w_8560 ,  , w_8561 );
buf ( w_8559 , \3708_b1 );
not ( w_8559 , w_8562 );
not (  , w_8563 );
and ( w_8562 , w_8563 , \3708_b0 );
or ( \3710_b1 , \3709_b1 , w_8564 );
xor ( \3710_b0 , \3709_b0 , w_8566 );
not ( w_8566 , w_8567 );
and ( w_8567 , w_8564 , w_8565 );
buf ( w_8564 , \1332_b1 );
not ( w_8564 , w_8568 );
not ( w_8565 , w_8569 );
and ( w_8568 , w_8569 , \1332_b0 );
or ( \3711_b1 , \3706_b1 , \3710_b1 );
not ( \3710_b1 , w_8570 );
and ( \3711_b0 , \3706_b0 , w_8571 );
and ( w_8570 , w_8571 , \3710_b0 );
or ( \3712_b1 , \1553_b1 , \1349_b1 );
not ( \1349_b1 , w_8572 );
and ( \3712_b0 , \1553_b0 , w_8573 );
and ( w_8572 , w_8573 , \1349_b0 );
or ( \3713_b1 , \1533_b1 , \1347_b1 );
not ( \1347_b1 , w_8574 );
and ( \3713_b0 , \1533_b0 , w_8575 );
and ( w_8574 , w_8575 , \1347_b0 );
or ( \3714_b1 , \3712_b1 , w_8577 );
not ( w_8577 , w_8578 );
and ( \3714_b0 , \3712_b0 , w_8579 );
and ( w_8578 ,  , w_8579 );
buf ( w_8577 , \3713_b1 );
not ( w_8577 , w_8580 );
not (  , w_8581 );
and ( w_8580 , w_8581 , \3713_b0 );
or ( \3715_b1 , \3714_b1 , w_8582 );
xor ( \3715_b0 , \3714_b0 , w_8584 );
not ( w_8584 , w_8585 );
and ( w_8585 , w_8582 , w_8583 );
buf ( w_8582 , \1356_b1 );
not ( w_8582 , w_8586 );
not ( w_8583 , w_8587 );
and ( w_8586 , w_8587 , \1356_b0 );
or ( \3716_b1 , \3710_b1 , \3715_b1 );
not ( \3715_b1 , w_8588 );
and ( \3716_b0 , \3710_b0 , w_8589 );
and ( w_8588 , w_8589 , \3715_b0 );
or ( \3717_b1 , \3706_b1 , \3715_b1 );
not ( \3715_b1 , w_8590 );
and ( \3717_b0 , \3706_b0 , w_8591 );
and ( w_8590 , w_8591 , \3715_b0 );
or ( \3719_b1 , \3627_b1 , \3631_b1 );
xor ( \3719_b0 , \3627_b0 , w_8592 );
not ( w_8592 , w_8593 );
and ( w_8593 , \3631_b1 , \3631_b0 );
or ( \3720_b1 , \3719_b1 , \3636_b1 );
xor ( \3720_b0 , \3719_b0 , w_8594 );
not ( w_8594 , w_8595 );
and ( w_8595 , \3636_b1 , \3636_b0 );
or ( \3721_b1 , \3718_b1 , \3720_b1 );
not ( \3720_b1 , w_8596 );
and ( \3721_b0 , \3718_b0 , w_8597 );
and ( w_8596 , w_8597 , \3720_b0 );
or ( \3722_b1 , \3664_b1 , \3676_b1 );
xor ( \3722_b0 , \3664_b0 , w_8598 );
not ( w_8598 , w_8599 );
and ( w_8599 , \3676_b1 , \3676_b0 );
or ( \3723_b1 , \3722_b1 , \3681_b1 );
xor ( \3723_b0 , \3722_b0 , w_8600 );
not ( w_8600 , w_8601 );
and ( w_8601 , \3681_b1 , \3681_b0 );
or ( \3724_b1 , \3720_b1 , \3723_b1 );
not ( \3723_b1 , w_8602 );
and ( \3724_b0 , \3720_b0 , w_8603 );
and ( w_8602 , w_8603 , \3723_b0 );
or ( \3725_b1 , \3718_b1 , \3723_b1 );
not ( \3723_b1 , w_8604 );
and ( \3725_b0 , \3718_b0 , w_8605 );
and ( w_8604 , w_8605 , \3723_b0 );
or ( \3727_b1 , \3698_b1 , \3726_b1 );
not ( \3726_b1 , w_8606 );
and ( \3727_b0 , \3698_b0 , w_8607 );
and ( w_8606 , w_8607 , \3726_b0 );
or ( \3728_b1 , \3698_b1 , \3726_b1 );
xor ( \3728_b0 , \3698_b0 , w_8608 );
not ( w_8608 , w_8609 );
and ( w_8609 , \3726_b1 , \3726_b0 );
or ( \3729_b1 , \3718_b1 , \3720_b1 );
xor ( \3729_b0 , \3718_b0 , w_8610 );
not ( w_8610 , w_8611 );
and ( w_8611 , \3720_b1 , \3720_b0 );
or ( \3730_b1 , \3729_b1 , \3723_b1 );
xor ( \3730_b0 , \3729_b0 , w_8612 );
not ( w_8612 , w_8613 );
and ( w_8613 , \3723_b1 , \3723_b0 );
or ( \3731_b1 , \1622_b1 , \1336_b1 );
not ( \1336_b1 , w_8614 );
and ( \3731_b0 , \1622_b0 , w_8615 );
and ( w_8614 , w_8615 , \1336_b0 );
or ( \3732_b1 , \1407_b1 , \1333_b1 );
not ( \1333_b1 , w_8616 );
and ( \3732_b0 , \1407_b0 , w_8617 );
and ( w_8616 , w_8617 , \1333_b0 );
or ( \3733_b1 , \3731_b1 , w_8619 );
not ( w_8619 , w_8620 );
and ( \3733_b0 , \3731_b0 , w_8621 );
and ( w_8620 ,  , w_8621 );
buf ( w_8619 , \3732_b1 );
not ( w_8619 , w_8622 );
not (  , w_8623 );
and ( w_8622 , w_8623 , \3732_b0 );
or ( \3734_b1 , \3733_b1 , w_8624 );
xor ( \3734_b0 , \3733_b0 , w_8626 );
not ( w_8626 , w_8627 );
and ( w_8627 , w_8624 , w_8625 );
buf ( w_8624 , \1332_b1 );
not ( w_8624 , w_8628 );
not ( w_8625 , w_8629 );
and ( w_8628 , w_8629 , \1332_b0 );
or ( \3735_b1 , \1533_b1 , \1444_b1 );
not ( \1444_b1 , w_8630 );
and ( \3735_b0 , \1533_b0 , w_8631 );
and ( w_8630 , w_8631 , \1444_b0 );
or ( \3736_b1 , \1540_b1 , \1442_b1 );
not ( \1442_b1 , w_8632 );
and ( \3736_b0 , \1540_b0 , w_8633 );
and ( w_8632 , w_8633 , \1442_b0 );
or ( \3737_b1 , \3735_b1 , w_8635 );
not ( w_8635 , w_8636 );
and ( \3737_b0 , \3735_b0 , w_8637 );
and ( w_8636 ,  , w_8637 );
buf ( w_8635 , \3736_b1 );
not ( w_8635 , w_8638 );
not (  , w_8639 );
and ( w_8638 , w_8639 , \3736_b0 );
or ( \3738_b1 , \3737_b1 , w_8640 );
xor ( \3738_b0 , \3737_b0 , w_8642 );
not ( w_8642 , w_8643 );
and ( w_8643 , w_8640 , w_8641 );
buf ( w_8640 , \1451_b1 );
not ( w_8640 , w_8644 );
not ( w_8641 , w_8645 );
and ( w_8644 , w_8645 , \1451_b0 );
or ( \3739_b1 , \3734_b1 , \3738_b1 );
not ( \3738_b1 , w_8646 );
and ( \3739_b0 , \3734_b0 , w_8647 );
and ( w_8646 , w_8647 , \3738_b0 );
or ( \3740_b1 , \1498_b1 , \1349_b1 );
not ( \1349_b1 , w_8648 );
and ( \3740_b0 , \1498_b0 , w_8649 );
and ( w_8648 , w_8649 , \1349_b0 );
or ( \3741_b1 , \1553_b1 , \1347_b1 );
not ( \1347_b1 , w_8650 );
and ( \3741_b0 , \1553_b0 , w_8651 );
and ( w_8650 , w_8651 , \1347_b0 );
or ( \3742_b1 , \3740_b1 , w_8653 );
not ( w_8653 , w_8654 );
and ( \3742_b0 , \3740_b0 , w_8655 );
and ( w_8654 ,  , w_8655 );
buf ( w_8653 , \3741_b1 );
not ( w_8653 , w_8656 );
not (  , w_8657 );
and ( w_8656 , w_8657 , \3741_b0 );
or ( \3743_b1 , \3742_b1 , w_8658 );
xor ( \3743_b0 , \3742_b0 , w_8660 );
not ( w_8660 , w_8661 );
and ( w_8661 , w_8658 , w_8659 );
buf ( w_8658 , \1356_b1 );
not ( w_8658 , w_8662 );
not ( w_8659 , w_8663 );
and ( w_8662 , w_8663 , \1356_b0 );
or ( \3744_b1 , \3738_b1 , \3743_b1 );
not ( \3743_b1 , w_8664 );
and ( \3744_b0 , \3738_b0 , w_8665 );
and ( w_8664 , w_8665 , \3743_b0 );
or ( \3745_b1 , \3734_b1 , \3743_b1 );
not ( \3743_b1 , w_8666 );
and ( \3745_b0 , \3734_b0 , w_8667 );
and ( w_8666 , w_8667 , \3743_b0 );
or ( \3747_b1 , \3668_b1 , \3672_b1 );
xor ( \3747_b0 , \3668_b0 , w_8668 );
not ( w_8668 , w_8669 );
and ( w_8669 , \3672_b1 , \3672_b0 );
or ( \3748_b1 , \3747_b1 , \3644_b1 );
xor ( \3748_b0 , \3747_b0 , w_8670 );
not ( w_8670 , w_8671 );
and ( w_8671 , \3644_b1 , \3644_b0 );
or ( \3749_b1 , \3746_b1 , \3748_b1 );
not ( \3748_b1 , w_8672 );
and ( \3749_b0 , \3746_b0 , w_8673 );
and ( w_8672 , w_8673 , \3748_b0 );
or ( \3750_b1 , \3706_b1 , \3710_b1 );
xor ( \3750_b0 , \3706_b0 , w_8674 );
not ( w_8674 , w_8675 );
and ( w_8675 , \3710_b1 , \3710_b0 );
or ( \3751_b1 , \3750_b1 , \3715_b1 );
xor ( \3751_b0 , \3750_b0 , w_8676 );
not ( w_8676 , w_8677 );
and ( w_8677 , \3715_b1 , \3715_b0 );
or ( \3752_b1 , \3748_b1 , \3751_b1 );
not ( \3751_b1 , w_8678 );
and ( \3752_b0 , \3748_b0 , w_8679 );
and ( w_8678 , w_8679 , \3751_b0 );
or ( \3753_b1 , \3746_b1 , \3751_b1 );
not ( \3751_b1 , w_8680 );
and ( \3753_b0 , \3746_b0 , w_8681 );
and ( w_8680 , w_8681 , \3751_b0 );
or ( \3755_b1 , \3730_b1 , \3754_b1 );
not ( \3754_b1 , w_8682 );
and ( \3755_b0 , \3730_b0 , w_8683 );
and ( w_8682 , w_8683 , \3754_b0 );
or ( \3756_b1 , \3730_b1 , \3754_b1 );
xor ( \3756_b0 , \3730_b0 , w_8684 );
not ( w_8684 , w_8685 );
and ( w_8685 , \3754_b1 , \3754_b0 );
or ( \3757_b1 , \3702_b1 , \3705_b1 );
xor ( \3757_b0 , \3702_b0 , w_8686 );
not ( w_8686 , w_8687 );
and ( w_8687 , \3705_b1 , \3705_b0 );
or ( \3758_b1 , \1540_b1 , \1431_b1 );
not ( \1431_b1 , w_8688 );
and ( \3758_b0 , \1540_b0 , w_8689 );
and ( w_8688 , w_8689 , \1431_b0 );
or ( \3759_b1 , \1517_b1 , \1429_b1 );
not ( \1429_b1 , w_8690 );
and ( \3759_b0 , \1517_b0 , w_8691 );
and ( w_8690 , w_8691 , \1429_b0 );
or ( \3760_b1 , \3758_b1 , w_8693 );
not ( w_8693 , w_8694 );
and ( \3760_b0 , \3758_b0 , w_8695 );
and ( w_8694 ,  , w_8695 );
buf ( w_8693 , \3759_b1 );
not ( w_8693 , w_8696 );
not (  , w_8697 );
and ( w_8696 , w_8697 , \3759_b0 );
or ( \3761_b1 , \3760_b1 , w_8698 );
xor ( \3761_b0 , \3760_b0 , w_8700 );
not ( w_8700 , w_8701 );
and ( w_8701 , w_8698 , w_8699 );
buf ( w_8698 , \1438_b1 );
not ( w_8698 , w_8702 );
not ( w_8699 , w_8703 );
and ( w_8702 , w_8703 , \1438_b0 );
or ( \3762_b1 , \1553_b1 , \1444_b1 );
not ( \1444_b1 , w_8704 );
and ( \3762_b0 , \1553_b0 , w_8705 );
and ( w_8704 , w_8705 , \1444_b0 );
or ( \3763_b1 , \1533_b1 , \1442_b1 );
not ( \1442_b1 , w_8706 );
and ( \3763_b0 , \1533_b0 , w_8707 );
and ( w_8706 , w_8707 , \1442_b0 );
or ( \3764_b1 , \3762_b1 , w_8709 );
not ( w_8709 , w_8710 );
and ( \3764_b0 , \3762_b0 , w_8711 );
and ( w_8710 ,  , w_8711 );
buf ( w_8709 , \3763_b1 );
not ( w_8709 , w_8712 );
not (  , w_8713 );
and ( w_8712 , w_8713 , \3763_b0 );
or ( \3765_b1 , \3764_b1 , w_8714 );
xor ( \3765_b0 , \3764_b0 , w_8716 );
not ( w_8716 , w_8717 );
and ( w_8717 , w_8714 , w_8715 );
buf ( w_8714 , \1451_b1 );
not ( w_8714 , w_8718 );
not ( w_8715 , w_8719 );
and ( w_8718 , w_8719 , \1451_b0 );
or ( \3766_b1 , \3761_b1 , \3765_b1 );
not ( \3765_b1 , w_8720 );
and ( \3766_b0 , \3761_b0 , w_8721 );
and ( w_8720 , w_8721 , \3765_b0 );
or ( \3767_b1 , \3765_b1 , \3703_b1 );
not ( \3703_b1 , w_8722 );
and ( \3767_b0 , \3765_b0 , w_8723 );
and ( w_8722 , w_8723 , \3703_b0 );
or ( \3768_b1 , \3761_b1 , \3703_b1 );
not ( \3703_b1 , w_8724 );
and ( \3768_b0 , \3761_b0 , w_8725 );
and ( w_8724 , w_8725 , \3703_b0 );
or ( \3770_b1 , \3757_b1 , \3769_b1 );
not ( \3769_b1 , w_8726 );
and ( \3770_b0 , \3757_b0 , w_8727 );
and ( w_8726 , w_8727 , \3769_b0 );
or ( \3771_b1 , \3734_b1 , \3738_b1 );
xor ( \3771_b0 , \3734_b0 , w_8728 );
not ( w_8728 , w_8729 );
and ( w_8729 , \3738_b1 , \3738_b0 );
or ( \3772_b1 , \3771_b1 , \3743_b1 );
xor ( \3772_b0 , \3771_b0 , w_8730 );
not ( w_8730 , w_8731 );
and ( w_8731 , \3743_b1 , \3743_b0 );
or ( \3773_b1 , \3769_b1 , \3772_b1 );
not ( \3772_b1 , w_8732 );
and ( \3773_b0 , \3769_b0 , w_8733 );
and ( w_8732 , w_8733 , \3772_b0 );
or ( \3774_b1 , \3757_b1 , \3772_b1 );
not ( \3772_b1 , w_8734 );
and ( \3774_b0 , \3757_b0 , w_8735 );
and ( w_8734 , w_8735 , \3772_b0 );
or ( \3776_b1 , \3746_b1 , \3748_b1 );
xor ( \3776_b0 , \3746_b0 , w_8736 );
not ( w_8736 , w_8737 );
and ( w_8737 , \3748_b1 , \3748_b0 );
or ( \3777_b1 , \3776_b1 , \3751_b1 );
xor ( \3777_b0 , \3776_b0 , w_8738 );
not ( w_8738 , w_8739 );
and ( w_8739 , \3751_b1 , \3751_b0 );
or ( \3778_b1 , \3775_b1 , \3777_b1 );
not ( \3777_b1 , w_8740 );
and ( \3778_b0 , \3775_b0 , w_8741 );
and ( w_8740 , w_8741 , \3777_b0 );
or ( \3779_b1 , \3775_b1 , \3777_b1 );
xor ( \3779_b0 , \3775_b0 , w_8742 );
not ( w_8742 , w_8743 );
and ( w_8743 , \3777_b1 , \3777_b0 );
or ( \3780_b1 , \3757_b1 , \3769_b1 );
xor ( \3780_b0 , \3757_b0 , w_8744 );
not ( w_8744 , w_8745 );
and ( w_8745 , \3769_b1 , \3769_b0 );
or ( \3781_b1 , \3780_b1 , \3772_b1 );
xor ( \3781_b0 , \3780_b0 , w_8746 );
not ( w_8746 , w_8747 );
and ( w_8747 , \3772_b1 , \3772_b0 );
or ( \3782_b1 , \1533_b1 , \1431_b1 );
not ( \1431_b1 , w_8748 );
and ( \3782_b0 , \1533_b0 , w_8749 );
and ( w_8748 , w_8749 , \1431_b0 );
or ( \3783_b1 , \1540_b1 , \1429_b1 );
not ( \1429_b1 , w_8750 );
and ( \3783_b0 , \1540_b0 , w_8751 );
and ( w_8750 , w_8751 , \1429_b0 );
or ( \3784_b1 , \3782_b1 , w_8753 );
not ( w_8753 , w_8754 );
and ( \3784_b0 , \3782_b0 , w_8755 );
and ( w_8754 ,  , w_8755 );
buf ( w_8753 , \3783_b1 );
not ( w_8753 , w_8756 );
not (  , w_8757 );
and ( w_8756 , w_8757 , \3783_b0 );
or ( \3785_b1 , \3784_b1 , w_8758 );
xor ( \3785_b0 , \3784_b0 , w_8760 );
not ( w_8760 , w_8761 );
and ( w_8761 , w_8758 , w_8759 );
buf ( w_8758 , \1438_b1 );
not ( w_8758 , w_8762 );
not ( w_8759 , w_8763 );
and ( w_8762 , w_8763 , \1438_b0 );
or ( \3786_b1 , \1498_b1 , \1442_b1 );
not ( \1442_b1 , w_8764 );
and ( \3786_b0 , \1498_b0 , w_8765 );
and ( w_8764 , w_8765 , \1442_b0 );
buf ( \3787_b1 , \3786_b1 );
not ( \3787_b1 , w_8766 );
not ( \3787_b0 , w_8767 );
and ( w_8766 , w_8767 , \3786_b0 );
or ( \3788_b1 , \3787_b1 , \1451_b1 );
not ( \1451_b1 , w_8768 );
and ( \3788_b0 , \3787_b0 , w_8769 );
and ( w_8768 , w_8769 , \1451_b0 );
or ( \3789_b1 , \3785_b1 , \3788_b1 );
not ( \3788_b1 , w_8770 );
and ( \3789_b0 , \3785_b0 , w_8771 );
and ( w_8770 , w_8771 , \3788_b0 );
or ( \3790_b1 , \1526_b1 , \1336_b1 );
not ( \1336_b1 , w_8772 );
and ( \3790_b0 , \1526_b0 , w_8773 );
and ( w_8772 , w_8773 , \1336_b0 );
or ( \3791_b1 , \1622_b1 , \1333_b1 );
not ( \1333_b1 , w_8774 );
and ( \3791_b0 , \1622_b0 , w_8775 );
and ( w_8774 , w_8775 , \1333_b0 );
or ( \3792_b1 , \3790_b1 , w_8777 );
not ( w_8777 , w_8778 );
and ( \3792_b0 , \3790_b0 , w_8779 );
and ( w_8778 ,  , w_8779 );
buf ( w_8777 , \3791_b1 );
not ( w_8777 , w_8780 );
not (  , w_8781 );
and ( w_8780 , w_8781 , \3791_b0 );
or ( \3793_b1 , \3792_b1 , w_8782 );
xor ( \3793_b0 , \3792_b0 , w_8784 );
not ( w_8784 , w_8785 );
and ( w_8785 , w_8782 , w_8783 );
buf ( w_8782 , \1332_b1 );
not ( w_8782 , w_8786 );
not ( w_8783 , w_8787 );
and ( w_8786 , w_8787 , \1332_b0 );
or ( \3794_b1 , \3789_b1 , \3793_b1 );
not ( \3793_b1 , w_8788 );
and ( \3794_b0 , \3789_b0 , w_8789 );
and ( w_8788 , w_8789 , \3793_b0 );
or ( \3795_b1 , \3761_b1 , \3765_b1 );
xor ( \3795_b0 , \3761_b0 , w_8790 );
not ( w_8790 , w_8791 );
and ( w_8791 , \3765_b1 , \3765_b0 );
or ( \3796_b1 , \3795_b1 , \3703_b1 );
xor ( \3796_b0 , \3795_b0 , w_8792 );
not ( w_8792 , w_8793 );
and ( w_8793 , \3703_b1 , \3703_b0 );
or ( \3797_b1 , \3793_b1 , \3796_b1 );
not ( \3796_b1 , w_8794 );
and ( \3797_b0 , \3793_b0 , w_8795 );
and ( w_8794 , w_8795 , \3796_b0 );
or ( \3798_b1 , \3789_b1 , \3796_b1 );
not ( \3796_b1 , w_8796 );
and ( \3798_b0 , \3789_b0 , w_8797 );
and ( w_8796 , w_8797 , \3796_b0 );
or ( \3800_b1 , \3781_b1 , \3799_b1 );
not ( \3799_b1 , w_8798 );
and ( \3800_b0 , \3781_b0 , w_8799 );
and ( w_8798 , w_8799 , \3799_b0 );
or ( \3801_b1 , \3781_b1 , \3799_b1 );
xor ( \3801_b0 , \3781_b0 , w_8800 );
not ( w_8800 , w_8801 );
and ( w_8801 , \3799_b1 , \3799_b0 );
or ( \3802_b1 , \3789_b1 , \3793_b1 );
xor ( \3802_b0 , \3789_b0 , w_8802 );
not ( w_8802 , w_8803 );
and ( w_8803 , \3793_b1 , \3793_b0 );
or ( \3803_b1 , \3802_b1 , \3796_b1 );
xor ( \3803_b0 , \3802_b0 , w_8804 );
not ( w_8804 , w_8805 );
and ( w_8805 , \3796_b1 , \3796_b0 );
or ( \3804_b1 , \3785_b1 , \3788_b1 );
xor ( \3804_b0 , \3785_b0 , w_8806 );
not ( w_8806 , w_8807 );
and ( w_8807 , \3788_b1 , \3788_b0 );
or ( \3805_b1 , \1517_b1 , \1336_b1 );
not ( \1336_b1 , w_8808 );
and ( \3805_b0 , \1517_b0 , w_8809 );
and ( w_8808 , w_8809 , \1336_b0 );
or ( \3806_b1 , \1526_b1 , \1333_b1 );
not ( \1333_b1 , w_8810 );
and ( \3806_b0 , \1526_b0 , w_8811 );
and ( w_8810 , w_8811 , \1333_b0 );
or ( \3807_b1 , \3805_b1 , w_8813 );
not ( w_8813 , w_8814 );
and ( \3807_b0 , \3805_b0 , w_8815 );
and ( w_8814 ,  , w_8815 );
buf ( w_8813 , \3806_b1 );
not ( w_8813 , w_8816 );
not (  , w_8817 );
and ( w_8816 , w_8817 , \3806_b0 );
or ( \3808_b1 , \3807_b1 , w_8818 );
xor ( \3808_b0 , \3807_b0 , w_8820 );
not ( w_8820 , w_8821 );
and ( w_8821 , w_8818 , w_8819 );
buf ( w_8818 , \1332_b1 );
not ( w_8818 , w_8822 );
not ( w_8819 , w_8823 );
and ( w_8822 , w_8823 , \1332_b0 );
or ( \3809_b1 , \3804_b1 , \3808_b1 );
not ( \3808_b1 , w_8824 );
and ( \3809_b0 , \3804_b0 , w_8825 );
and ( w_8824 , w_8825 , \3808_b0 );
or ( \3810_b1 , \1498_b1 , \1444_b1 );
not ( \1444_b1 , w_8826 );
and ( \3810_b0 , \1498_b0 , w_8827 );
and ( w_8826 , w_8827 , \1444_b0 );
or ( \3811_b1 , \1553_b1 , \1442_b1 );
not ( \1442_b1 , w_8828 );
and ( \3811_b0 , \1553_b0 , w_8829 );
and ( w_8828 , w_8829 , \1442_b0 );
or ( \3812_b1 , \3810_b1 , w_8831 );
not ( w_8831 , w_8832 );
and ( \3812_b0 , \3810_b0 , w_8833 );
and ( w_8832 ,  , w_8833 );
buf ( w_8831 , \3811_b1 );
not ( w_8831 , w_8834 );
not (  , w_8835 );
and ( w_8834 , w_8835 , \3811_b0 );
or ( \3813_b1 , \3812_b1 , w_8836 );
xor ( \3813_b0 , \3812_b0 , w_8838 );
not ( w_8838 , w_8839 );
and ( w_8839 , w_8836 , w_8837 );
buf ( w_8836 , \1451_b1 );
not ( w_8836 , w_8840 );
not ( w_8837 , w_8841 );
and ( w_8840 , w_8841 , \1451_b0 );
or ( \3814_b1 , \3808_b1 , \3813_b1 );
not ( \3813_b1 , w_8842 );
and ( \3814_b0 , \3808_b0 , w_8843 );
and ( w_8842 , w_8843 , \3813_b0 );
or ( \3815_b1 , \3804_b1 , \3813_b1 );
not ( \3813_b1 , w_8844 );
and ( \3815_b0 , \3804_b0 , w_8845 );
and ( w_8844 , w_8845 , \3813_b0 );
or ( \3817_b1 , \3803_b1 , \3816_b1 );
not ( \3816_b1 , w_8846 );
and ( \3817_b0 , \3803_b0 , w_8847 );
and ( w_8846 , w_8847 , \3816_b0 );
or ( \3818_b1 , \3803_b1 , \3816_b1 );
xor ( \3818_b0 , \3803_b0 , w_8848 );
not ( w_8848 , w_8849 );
and ( w_8849 , \3816_b1 , \3816_b0 );
or ( \3819_b1 , \1540_b1 , \1336_b1 );
not ( \1336_b1 , w_8850 );
and ( \3819_b0 , \1540_b0 , w_8851 );
and ( w_8850 , w_8851 , \1336_b0 );
or ( \3820_b1 , \1517_b1 , \1333_b1 );
not ( \1333_b1 , w_8852 );
and ( \3820_b0 , \1517_b0 , w_8853 );
and ( w_8852 , w_8853 , \1333_b0 );
or ( \3821_b1 , \3819_b1 , w_8855 );
not ( w_8855 , w_8856 );
and ( \3821_b0 , \3819_b0 , w_8857 );
and ( w_8856 ,  , w_8857 );
buf ( w_8855 , \3820_b1 );
not ( w_8855 , w_8858 );
not (  , w_8859 );
and ( w_8858 , w_8859 , \3820_b0 );
or ( \3822_b1 , \3821_b1 , w_8860 );
xor ( \3822_b0 , \3821_b0 , w_8862 );
not ( w_8862 , w_8863 );
and ( w_8863 , w_8860 , w_8861 );
buf ( w_8860 , \1332_b1 );
not ( w_8860 , w_8864 );
not ( w_8861 , w_8865 );
and ( w_8864 , w_8865 , \1332_b0 );
or ( \3823_b1 , \1553_b1 , \1431_b1 );
not ( \1431_b1 , w_8866 );
and ( \3823_b0 , \1553_b0 , w_8867 );
and ( w_8866 , w_8867 , \1431_b0 );
or ( \3824_b1 , \1533_b1 , \1429_b1 );
not ( \1429_b1 , w_8868 );
and ( \3824_b0 , \1533_b0 , w_8869 );
and ( w_8868 , w_8869 , \1429_b0 );
or ( \3825_b1 , \3823_b1 , w_8871 );
not ( w_8871 , w_8872 );
and ( \3825_b0 , \3823_b0 , w_8873 );
and ( w_8872 ,  , w_8873 );
buf ( w_8871 , \3824_b1 );
not ( w_8871 , w_8874 );
not (  , w_8875 );
and ( w_8874 , w_8875 , \3824_b0 );
or ( \3826_b1 , \3825_b1 , w_8876 );
xor ( \3826_b0 , \3825_b0 , w_8878 );
not ( w_8878 , w_8879 );
and ( w_8879 , w_8876 , w_8877 );
buf ( w_8876 , \1438_b1 );
not ( w_8876 , w_8880 );
not ( w_8877 , w_8881 );
and ( w_8880 , w_8881 , \1438_b0 );
or ( \3827_b1 , \3822_b1 , \3826_b1 );
not ( \3826_b1 , w_8882 );
and ( \3827_b0 , \3822_b0 , w_8883 );
and ( w_8882 , w_8883 , \3826_b0 );
or ( \3828_b1 , \3826_b1 , \3786_b1 );
not ( \3786_b1 , w_8884 );
and ( \3828_b0 , \3826_b0 , w_8885 );
and ( w_8884 , w_8885 , \3786_b0 );
or ( \3829_b1 , \3822_b1 , \3786_b1 );
not ( \3786_b1 , w_8886 );
and ( \3829_b0 , \3822_b0 , w_8887 );
and ( w_8886 , w_8887 , \3786_b0 );
or ( \3831_b1 , \3804_b1 , \3808_b1 );
xor ( \3831_b0 , \3804_b0 , w_8888 );
not ( w_8888 , w_8889 );
and ( w_8889 , \3808_b1 , \3808_b0 );
or ( \3832_b1 , \3831_b1 , \3813_b1 );
xor ( \3832_b0 , \3831_b0 , w_8890 );
not ( w_8890 , w_8891 );
and ( w_8891 , \3813_b1 , \3813_b0 );
or ( \3833_b1 , \3830_b1 , \3832_b1 );
not ( \3832_b1 , w_8892 );
and ( \3833_b0 , \3830_b0 , w_8893 );
and ( w_8892 , w_8893 , \3832_b0 );
or ( \3834_b1 , \3830_b1 , \3832_b1 );
xor ( \3834_b0 , \3830_b0 , w_8894 );
not ( w_8894 , w_8895 );
and ( w_8895 , \3832_b1 , \3832_b0 );
or ( \3835_b1 , \3822_b1 , \3826_b1 );
xor ( \3835_b0 , \3822_b0 , w_8896 );
not ( w_8896 , w_8897 );
and ( w_8897 , \3826_b1 , \3826_b0 );
or ( \3836_b1 , \3835_b1 , \3786_b1 );
xor ( \3836_b0 , \3835_b0 , w_8898 );
not ( w_8898 , w_8899 );
and ( w_8899 , \3786_b1 , \3786_b0 );
or ( \3837_b1 , \1498_b1 , \1429_b1 );
not ( \1429_b1 , w_8900 );
and ( \3837_b0 , \1498_b0 , w_8901 );
and ( w_8900 , w_8901 , \1429_b0 );
buf ( \3838_b1 , \3837_b1 );
not ( \3838_b1 , w_8902 );
not ( \3838_b0 , w_8903 );
and ( w_8902 , w_8903 , \3837_b0 );
or ( \3839_b1 , \3838_b1 , \1438_b1 );
not ( \1438_b1 , w_8904 );
and ( \3839_b0 , \3838_b0 , w_8905 );
and ( w_8904 , w_8905 , \1438_b0 );
or ( \3840_b1 , \1498_b1 , \1431_b1 );
not ( \1431_b1 , w_8906 );
and ( \3840_b0 , \1498_b0 , w_8907 );
and ( w_8906 , w_8907 , \1431_b0 );
or ( \3841_b1 , \1553_b1 , \1429_b1 );
not ( \1429_b1 , w_8908 );
and ( \3841_b0 , \1553_b0 , w_8909 );
and ( w_8908 , w_8909 , \1429_b0 );
or ( \3842_b1 , \3840_b1 , w_8911 );
not ( w_8911 , w_8912 );
and ( \3842_b0 , \3840_b0 , w_8913 );
and ( w_8912 ,  , w_8913 );
buf ( w_8911 , \3841_b1 );
not ( w_8911 , w_8914 );
not (  , w_8915 );
and ( w_8914 , w_8915 , \3841_b0 );
or ( \3843_b1 , \3842_b1 , w_8916 );
xor ( \3843_b0 , \3842_b0 , w_8918 );
not ( w_8918 , w_8919 );
and ( w_8919 , w_8916 , w_8917 );
buf ( w_8916 , \1438_b1 );
not ( w_8916 , w_8920 );
not ( w_8917 , w_8921 );
and ( w_8920 , w_8921 , \1438_b0 );
or ( \3844_b1 , \3839_b1 , \3843_b1 );
not ( \3843_b1 , w_8922 );
and ( \3844_b0 , \3839_b0 , w_8923 );
and ( w_8922 , w_8923 , \3843_b0 );
or ( \3845_b1 , \3836_b1 , \3844_b1 );
not ( \3844_b1 , w_8924 );
and ( \3845_b0 , \3836_b0 , w_8925 );
and ( w_8924 , w_8925 , \3844_b0 );
or ( \3846_b1 , \3836_b1 , \3844_b1 );
xor ( \3846_b0 , \3836_b0 , w_8926 );
not ( w_8926 , w_8927 );
and ( w_8927 , \3844_b1 , \3844_b0 );
or ( \3847_b1 , \1533_b1 , \1336_b1 );
not ( \1336_b1 , w_8928 );
and ( \3847_b0 , \1533_b0 , w_8929 );
and ( w_8928 , w_8929 , \1336_b0 );
or ( \3848_b1 , \1540_b1 , \1333_b1 );
not ( \1333_b1 , w_8930 );
and ( \3848_b0 , \1540_b0 , w_8931 );
and ( w_8930 , w_8931 , \1333_b0 );
or ( \3849_b1 , \3847_b1 , w_8933 );
not ( w_8933 , w_8934 );
and ( \3849_b0 , \3847_b0 , w_8935 );
and ( w_8934 ,  , w_8935 );
buf ( w_8933 , \3848_b1 );
not ( w_8933 , w_8936 );
not (  , w_8937 );
and ( w_8936 , w_8937 , \3848_b0 );
or ( \3850_b1 , \3849_b1 , w_8938 );
xor ( \3850_b0 , \3849_b0 , w_8940 );
not ( w_8940 , w_8941 );
and ( w_8941 , w_8938 , w_8939 );
buf ( w_8938 , \1332_b1 );
not ( w_8938 , w_8942 );
not ( w_8939 , w_8943 );
and ( w_8942 , w_8943 , \1332_b0 );
or ( \3851_b1 , \3839_b1 , \3843_b1 );
xor ( \3851_b0 , \3839_b0 , w_8944 );
not ( w_8944 , w_8945 );
and ( w_8945 , \3843_b1 , \3843_b0 );
or ( \3852_b1 , \3850_b1 , \3851_b1 );
not ( \3851_b1 , w_8946 );
and ( \3852_b0 , \3850_b0 , w_8947 );
and ( w_8946 , w_8947 , \3851_b0 );
or ( \3853_b1 , \3850_b1 , \3851_b1 );
xor ( \3853_b0 , \3850_b0 , w_8948 );
not ( w_8948 , w_8949 );
and ( w_8949 , \3851_b1 , \3851_b0 );
or ( \3854_b1 , \1553_b1 , \1336_b1 );
not ( \1336_b1 , w_8950 );
and ( \3854_b0 , \1553_b0 , w_8951 );
and ( w_8950 , w_8951 , \1336_b0 );
or ( \3855_b1 , \1533_b1 , \1333_b1 );
not ( \1333_b1 , w_8952 );
and ( \3855_b0 , \1533_b0 , w_8953 );
and ( w_8952 , w_8953 , \1333_b0 );
or ( \3856_b1 , \3854_b1 , w_8955 );
not ( w_8955 , w_8956 );
and ( \3856_b0 , \3854_b0 , w_8957 );
and ( w_8956 ,  , w_8957 );
buf ( w_8955 , \3855_b1 );
not ( w_8955 , w_8958 );
not (  , w_8959 );
and ( w_8958 , w_8959 , \3855_b0 );
or ( \3857_b1 , \3856_b1 , w_8960 );
xor ( \3857_b0 , \3856_b0 , w_8962 );
not ( w_8962 , w_8963 );
and ( w_8963 , w_8960 , w_8961 );
buf ( w_8960 , \1332_b1 );
not ( w_8960 , w_8964 );
not ( w_8961 , w_8965 );
and ( w_8964 , w_8965 , \1332_b0 );
or ( \3858_b1 , \3857_b1 , \3837_b1 );
not ( \3837_b1 , w_8966 );
and ( \3858_b0 , \3857_b0 , w_8967 );
and ( w_8966 , w_8967 , \3837_b0 );
or ( \3859_b1 , \3857_b1 , \3837_b1 );
xor ( \3859_b0 , \3857_b0 , w_8968 );
not ( w_8968 , w_8969 );
and ( w_8969 , \3837_b1 , \3837_b0 );
or ( \3860_b1 , \1498_b1 , \1336_b1 );
not ( \1336_b1 , w_8970 );
and ( \3860_b0 , \1498_b0 , w_8971 );
and ( w_8970 , w_8971 , \1336_b0 );
or ( \3861_b1 , \1553_b1 , \1333_b1 );
not ( \1333_b1 , w_8972 );
and ( \3861_b0 , \1553_b0 , w_8973 );
and ( w_8972 , w_8973 , \1333_b0 );
or ( \3862_b1 , \3860_b1 , w_8975 );
not ( w_8975 , w_8976 );
and ( \3862_b0 , \3860_b0 , w_8977 );
and ( w_8976 ,  , w_8977 );
buf ( w_8975 , \3861_b1 );
not ( w_8975 , w_8978 );
not (  , w_8979 );
and ( w_8978 , w_8979 , \3861_b0 );
or ( \3863_b1 , \3862_b1 , w_8980 );
xor ( \3863_b0 , \3862_b0 , w_8982 );
not ( w_8982 , w_8983 );
and ( w_8983 , w_8980 , w_8981 );
buf ( w_8980 , \1332_b1 );
not ( w_8980 , w_8984 );
not ( w_8981 , w_8985 );
and ( w_8984 , w_8985 , \1332_b0 );
or ( \3864_b1 , \1498_b1 , \1333_b1 );
not ( \1333_b1 , w_8986 );
and ( \3864_b0 , \1498_b0 , w_8987 );
and ( w_8986 , w_8987 , \1333_b0 );
buf ( \3865_b1 , \3864_b1 );
not ( \3865_b1 , w_8988 );
not ( \3865_b0 , w_8989 );
and ( w_8988 , w_8989 , \3864_b0 );
or ( \3866_b1 , \3865_b1 , \1332_b1 );
not ( \1332_b1 , w_8990 );
and ( \3866_b0 , \3865_b0 , w_8991 );
and ( w_8990 , w_8991 , \1332_b0 );
or ( \3867_b1 , \3863_b1 , \3866_b1 );
not ( \3866_b1 , w_8992 );
and ( \3867_b0 , \3863_b0 , w_8993 );
and ( w_8992 , w_8993 , \3866_b0 );
or ( \3868_b1 , \3859_b1 , \3867_b1 );
not ( \3867_b1 , w_8994 );
and ( \3868_b0 , \3859_b0 , w_8995 );
and ( w_8994 , w_8995 , \3867_b0 );
or ( \3869_b1 , \3858_b1 , w_8996 );
or ( \3869_b0 , \3858_b0 , \3868_b0 );
not ( \3868_b0 , w_8997 );
and ( w_8997 , w_8996 , \3868_b1 );
or ( \3870_b1 , \3853_b1 , \3869_b1 );
not ( \3869_b1 , w_8998 );
and ( \3870_b0 , \3853_b0 , w_8999 );
and ( w_8998 , w_8999 , \3869_b0 );
or ( \3871_b1 , \3852_b1 , w_9000 );
or ( \3871_b0 , \3852_b0 , \3870_b0 );
not ( \3870_b0 , w_9001 );
and ( w_9001 , w_9000 , \3870_b1 );
or ( \3872_b1 , \3846_b1 , \3871_b1 );
not ( \3871_b1 , w_9002 );
and ( \3872_b0 , \3846_b0 , w_9003 );
and ( w_9002 , w_9003 , \3871_b0 );
or ( \3873_b1 , \3845_b1 , w_9004 );
or ( \3873_b0 , \3845_b0 , \3872_b0 );
not ( \3872_b0 , w_9005 );
and ( w_9005 , w_9004 , \3872_b1 );
or ( \3874_b1 , \3834_b1 , \3873_b1 );
not ( \3873_b1 , w_9006 );
and ( \3874_b0 , \3834_b0 , w_9007 );
and ( w_9006 , w_9007 , \3873_b0 );
or ( \3875_b1 , \3833_b1 , w_9008 );
or ( \3875_b0 , \3833_b0 , \3874_b0 );
not ( \3874_b0 , w_9009 );
and ( w_9009 , w_9008 , \3874_b1 );
or ( \3876_b1 , \3818_b1 , \3875_b1 );
not ( \3875_b1 , w_9010 );
and ( \3876_b0 , \3818_b0 , w_9011 );
and ( w_9010 , w_9011 , \3875_b0 );
or ( \3877_b1 , \3817_b1 , w_9012 );
or ( \3877_b0 , \3817_b0 , \3876_b0 );
not ( \3876_b0 , w_9013 );
and ( w_9013 , w_9012 , \3876_b1 );
or ( \3878_b1 , \3801_b1 , \3877_b1 );
not ( \3877_b1 , w_9014 );
and ( \3878_b0 , \3801_b0 , w_9015 );
and ( w_9014 , w_9015 , \3877_b0 );
or ( \3879_b1 , \3800_b1 , w_9016 );
or ( \3879_b0 , \3800_b0 , \3878_b0 );
not ( \3878_b0 , w_9017 );
and ( w_9017 , w_9016 , \3878_b1 );
or ( \3880_b1 , \3779_b1 , \3879_b1 );
not ( \3879_b1 , w_9018 );
and ( \3880_b0 , \3779_b0 , w_9019 );
and ( w_9018 , w_9019 , \3879_b0 );
or ( \3881_b1 , \3778_b1 , w_9020 );
or ( \3881_b0 , \3778_b0 , \3880_b0 );
not ( \3880_b0 , w_9021 );
and ( w_9021 , w_9020 , \3880_b1 );
or ( \3882_b1 , \3756_b1 , \3881_b1 );
not ( \3881_b1 , w_9022 );
and ( \3882_b0 , \3756_b0 , w_9023 );
and ( w_9022 , w_9023 , \3881_b0 );
or ( \3883_b1 , \3755_b1 , w_9024 );
or ( \3883_b0 , \3755_b0 , \3882_b0 );
not ( \3882_b0 , w_9025 );
and ( w_9025 , w_9024 , \3882_b1 );
or ( \3884_b1 , \3728_b1 , \3883_b1 );
not ( \3883_b1 , w_9026 );
and ( \3884_b0 , \3728_b0 , w_9027 );
and ( w_9026 , w_9027 , \3883_b0 );
or ( \3885_b1 , \3727_b1 , w_9028 );
or ( \3885_b0 , \3727_b0 , \3884_b0 );
not ( \3884_b0 , w_9029 );
and ( w_9029 , w_9028 , \3884_b1 );
or ( \3886_b1 , \3696_b1 , \3885_b1 );
not ( \3885_b1 , w_9030 );
and ( \3886_b0 , \3696_b0 , w_9031 );
and ( w_9030 , w_9031 , \3885_b0 );
or ( \3887_b1 , \3695_b1 , w_9032 );
or ( \3887_b0 , \3695_b0 , \3886_b0 );
not ( \3886_b0 , w_9033 );
and ( w_9033 , w_9032 , \3886_b1 );
or ( \3888_b1 , \3663_b1 , \3887_b1 );
not ( \3887_b1 , w_9034 );
and ( \3888_b0 , \3663_b0 , w_9035 );
and ( w_9034 , w_9035 , \3887_b0 );
or ( \3889_b1 , \3662_b1 , w_9036 );
or ( \3889_b0 , \3662_b0 , \3888_b0 );
not ( \3888_b0 , w_9037 );
and ( w_9037 , w_9036 , \3888_b1 );
or ( \3890_b1 , \3621_b1 , \3889_b1 );
not ( \3889_b1 , w_9038 );
and ( \3890_b0 , \3621_b0 , w_9039 );
and ( w_9038 , w_9039 , \3889_b0 );
or ( \3891_b1 , \3620_b1 , w_9040 );
or ( \3891_b0 , \3620_b0 , \3890_b0 );
not ( \3890_b0 , w_9041 );
and ( w_9041 , w_9040 , \3890_b1 );
or ( \3892_b1 , \3575_b1 , \3891_b1 );
not ( \3891_b1 , w_9042 );
and ( \3892_b0 , \3575_b0 , w_9043 );
and ( w_9042 , w_9043 , \3891_b0 );
or ( \3893_b1 , \3574_b1 , w_9044 );
or ( \3893_b0 , \3574_b0 , \3892_b0 );
not ( \3892_b0 , w_9045 );
and ( w_9045 , w_9044 , \3892_b1 );
or ( \3894_b1 , \3542_b1 , \3893_b1 );
not ( \3893_b1 , w_9046 );
and ( \3894_b0 , \3542_b0 , w_9047 );
and ( w_9046 , w_9047 , \3893_b0 );
or ( \3895_b1 , \3541_b1 , w_9048 );
or ( \3895_b0 , \3541_b0 , \3894_b0 );
not ( \3894_b0 , w_9049 );
and ( w_9049 , w_9048 , \3894_b1 );
or ( \3896_b1 , \3490_b1 , \3895_b1 );
not ( \3895_b1 , w_9050 );
and ( \3896_b0 , \3490_b0 , w_9051 );
and ( w_9050 , w_9051 , \3895_b0 );
or ( \3897_b1 , \3489_b1 , w_9052 );
or ( \3897_b0 , \3489_b0 , \3896_b0 );
not ( \3896_b0 , w_9053 );
and ( w_9053 , w_9052 , \3896_b1 );
or ( \3898_b1 , \3437_b1 , \3897_b1 );
not ( \3897_b1 , w_9054 );
and ( \3898_b0 , \3437_b0 , w_9055 );
and ( w_9054 , w_9055 , \3897_b0 );
or ( \3899_b1 , \3436_b1 , w_9056 );
or ( \3899_b0 , \3436_b0 , \3898_b0 );
not ( \3898_b0 , w_9057 );
and ( w_9057 , w_9056 , \3898_b1 );
or ( \3900_b1 , \3361_b1 , \3899_b1 );
not ( \3899_b1 , w_9058 );
and ( \3900_b0 , \3361_b0 , w_9059 );
and ( w_9058 , w_9059 , \3899_b0 );
or ( \3901_b1 , \3360_b1 , w_9060 );
or ( \3901_b0 , \3360_b0 , \3900_b0 );
not ( \3900_b0 , w_9061 );
and ( w_9061 , w_9060 , \3900_b1 );
or ( \3902_b1 , \3298_b1 , \3901_b1 );
not ( \3901_b1 , w_9062 );
and ( \3902_b0 , \3298_b0 , w_9063 );
and ( w_9062 , w_9063 , \3901_b0 );
or ( \3903_b1 , \3297_b1 , w_9064 );
or ( \3903_b0 , \3297_b0 , \3902_b0 );
not ( \3902_b0 , w_9065 );
and ( w_9065 , w_9064 , \3902_b1 );
or ( \3904_b1 , \3226_b1 , \3903_b1 );
not ( \3903_b1 , w_9066 );
and ( \3904_b0 , \3226_b0 , w_9067 );
and ( w_9066 , w_9067 , \3903_b0 );
or ( \3905_b1 , \3225_b1 , w_9068 );
or ( \3905_b0 , \3225_b0 , \3904_b0 );
not ( \3904_b0 , w_9069 );
and ( w_9069 , w_9068 , \3904_b1 );
or ( \3906_b1 , \3196_b1 , \3905_b1 );
not ( \3905_b1 , w_9070 );
and ( \3906_b0 , \3196_b0 , w_9071 );
and ( w_9070 , w_9071 , \3905_b0 );
or ( \3907_b1 , \3195_b1 , w_9072 );
or ( \3907_b0 , \3195_b0 , \3906_b0 );
not ( \3906_b0 , w_9073 );
and ( w_9073 , w_9072 , \3906_b1 );
or ( \3908_b1 , \3073_b1 , \3907_b1 );
not ( \3907_b1 , w_9074 );
and ( \3908_b0 , \3073_b0 , w_9075 );
and ( w_9074 , w_9075 , \3907_b0 );
or ( \3909_b1 , \3072_b1 , w_9076 );
or ( \3909_b0 , \3072_b0 , \3908_b0 );
not ( \3908_b0 , w_9077 );
and ( w_9077 , w_9076 , \3908_b1 );
or ( \3910_b1 , \3005_b1 , \3909_b1 );
not ( \3909_b1 , w_9078 );
and ( \3910_b0 , \3005_b0 , w_9079 );
and ( w_9078 , w_9079 , \3909_b0 );
or ( \3911_b1 , \3004_b1 , w_9080 );
or ( \3911_b0 , \3004_b0 , \3910_b0 );
not ( \3910_b0 , w_9081 );
and ( w_9081 , w_9080 , \3910_b1 );
or ( \3912_b1 , \2922_b1 , \3911_b1 );
not ( \3911_b1 , w_9082 );
and ( \3912_b0 , \2922_b0 , w_9083 );
and ( w_9082 , w_9083 , \3911_b0 );
or ( \3913_b1 , \2921_b1 , w_9084 );
or ( \3913_b0 , \2921_b0 , \3912_b0 );
not ( \3912_b0 , w_9085 );
and ( w_9085 , w_9084 , \3912_b1 );
or ( \3914_b1 , \2856_b1 , \3913_b1 );
not ( \3913_b1 , w_9086 );
and ( \3914_b0 , \2856_b0 , w_9087 );
and ( w_9086 , w_9087 , \3913_b0 );
or ( \3915_b1 , \2855_b1 , w_9088 );
or ( \3915_b0 , \2855_b0 , \3914_b0 );
not ( \3914_b0 , w_9089 );
and ( w_9089 , w_9088 , \3914_b1 );
or ( \3916_b1 , \2764_b1 , \3915_b1 );
not ( \3915_b1 , w_9090 );
and ( \3916_b0 , \2764_b0 , w_9091 );
and ( w_9090 , w_9091 , \3915_b0 );
or ( \3917_b1 , \2763_b1 , w_9092 );
or ( \3917_b0 , \2763_b0 , \3916_b0 );
not ( \3916_b0 , w_9093 );
and ( w_9093 , w_9092 , \3916_b1 );
or ( \3918_b1 , \2635_b1 , \3917_b1 );
not ( \3917_b1 , w_9094 );
and ( \3918_b0 , \2635_b0 , w_9095 );
and ( w_9094 , w_9095 , \3917_b0 );
or ( \3919_b1 , \2634_b1 , w_9096 );
or ( \3919_b0 , \2634_b0 , \3918_b0 );
not ( \3918_b0 , w_9097 );
and ( w_9097 , w_9096 , \3918_b1 );
or ( \3920_b1 , \2518_b1 , \3919_b1 );
not ( \3919_b1 , w_9098 );
and ( \3920_b0 , \2518_b0 , w_9099 );
and ( w_9098 , w_9099 , \3919_b0 );
or ( \3921_b1 , \2517_b1 , w_9100 );
or ( \3921_b0 , \2517_b0 , \3920_b0 );
not ( \3920_b0 , w_9101 );
and ( w_9101 , w_9100 , \3920_b1 );
or ( \3922_b1 , \2406_b1 , \3921_b1 );
not ( \3921_b1 , w_9102 );
and ( \3922_b0 , \2406_b0 , w_9103 );
and ( w_9102 , w_9103 , \3921_b0 );
or ( \3923_b1 , \2405_b1 , w_9104 );
or ( \3923_b0 , \2405_b0 , \3922_b0 );
not ( \3922_b0 , w_9105 );
and ( w_9105 , w_9104 , \3922_b1 );
or ( \3924_b1 , \2290_b1 , \3923_b1 );
not ( \3923_b1 , w_9106 );
and ( \3924_b0 , \2290_b0 , w_9107 );
and ( w_9106 , w_9107 , \3923_b0 );
or ( \3925_b1 , \2289_b1 , w_9108 );
or ( \3925_b0 , \2289_b0 , \3924_b0 );
not ( \3924_b0 , w_9109 );
and ( w_9109 , w_9108 , \3924_b1 );
or ( \3926_b1 , \2252_b1 , \3925_b1 );
xor ( \3926_b0 , \2252_b0 , w_9110 );
not ( w_9110 , w_9111 );
and ( w_9111 , \3925_b1 , \3925_b0 );
buf ( \3927_Z[31]_b1 , \3926_b1 );
buf ( \3927_Z[31]_b0 , \3926_b0 );
or ( \3928_b1 , \2290_b1 , \3923_b1 );
xor ( \3928_b0 , \2290_b0 , w_9112 );
not ( w_9112 , w_9113 );
and ( w_9113 , \3923_b1 , \3923_b0 );
buf ( \3929_Z[30]_b1 , \3928_b1 );
buf ( \3929_Z[30]_b0 , \3928_b0 );
or ( \3930_b1 , \2406_b1 , \3921_b1 );
xor ( \3930_b0 , \2406_b0 , w_9114 );
not ( w_9114 , w_9115 );
and ( w_9115 , \3921_b1 , \3921_b0 );
buf ( \3931_Z[29]_b1 , \3930_b1 );
buf ( \3931_Z[29]_b0 , \3930_b0 );
or ( \3932_b1 , \2518_b1 , \3919_b1 );
xor ( \3932_b0 , \2518_b0 , w_9116 );
not ( w_9116 , w_9117 );
and ( w_9117 , \3919_b1 , \3919_b0 );
buf ( \3933_Z[28]_b1 , \3932_b1 );
buf ( \3933_Z[28]_b0 , \3932_b0 );
or ( \3934_b1 , \2635_b1 , \3917_b1 );
xor ( \3934_b0 , \2635_b0 , w_9118 );
not ( w_9118 , w_9119 );
and ( w_9119 , \3917_b1 , \3917_b0 );
buf ( \3935_Z[27]_b1 , \3934_b1 );
buf ( \3935_Z[27]_b0 , \3934_b0 );
or ( \3936_b1 , \2764_b1 , \3915_b1 );
xor ( \3936_b0 , \2764_b0 , w_9120 );
not ( w_9120 , w_9121 );
and ( w_9121 , \3915_b1 , \3915_b0 );
buf ( \3937_Z[26]_b1 , \3936_b1 );
buf ( \3937_Z[26]_b0 , \3936_b0 );
or ( \3938_b1 , \2856_b1 , \3913_b1 );
xor ( \3938_b0 , \2856_b0 , w_9122 );
not ( w_9122 , w_9123 );
and ( w_9123 , \3913_b1 , \3913_b0 );
buf ( \3939_Z[25]_b1 , \3938_b1 );
buf ( \3939_Z[25]_b0 , \3938_b0 );
or ( \3940_b1 , \2922_b1 , \3911_b1 );
xor ( \3940_b0 , \2922_b0 , w_9124 );
not ( w_9124 , w_9125 );
and ( w_9125 , \3911_b1 , \3911_b0 );
buf ( \3941_Z[24]_b1 , \3940_b1 );
buf ( \3941_Z[24]_b0 , \3940_b0 );
or ( \3942_b1 , \3005_b1 , \3909_b1 );
xor ( \3942_b0 , \3005_b0 , w_9126 );
not ( w_9126 , w_9127 );
and ( w_9127 , \3909_b1 , \3909_b0 );
buf ( \3943_Z[23]_b1 , \3942_b1 );
buf ( \3943_Z[23]_b0 , \3942_b0 );
or ( \3944_b1 , \3073_b1 , \3907_b1 );
xor ( \3944_b0 , \3073_b0 , w_9128 );
not ( w_9128 , w_9129 );
and ( w_9129 , \3907_b1 , \3907_b0 );
buf ( \3945_Z[22]_b1 , \3944_b1 );
buf ( \3945_Z[22]_b0 , \3944_b0 );
or ( \3946_b1 , \3196_b1 , \3905_b1 );
xor ( \3946_b0 , \3196_b0 , w_9130 );
not ( w_9130 , w_9131 );
and ( w_9131 , \3905_b1 , \3905_b0 );
buf ( \3947_Z[21]_b1 , \3946_b1 );
buf ( \3947_Z[21]_b0 , \3946_b0 );
or ( \3948_b1 , \3226_b1 , \3903_b1 );
xor ( \3948_b0 , \3226_b0 , w_9132 );
not ( w_9132 , w_9133 );
and ( w_9133 , \3903_b1 , \3903_b0 );
buf ( \3949_Z[20]_b1 , \3948_b1 );
buf ( \3949_Z[20]_b0 , \3948_b0 );
or ( \3950_b1 , \3298_b1 , \3901_b1 );
xor ( \3950_b0 , \3298_b0 , w_9134 );
not ( w_9134 , w_9135 );
and ( w_9135 , \3901_b1 , \3901_b0 );
buf ( \3951_Z[19]_b1 , \3950_b1 );
buf ( \3951_Z[19]_b0 , \3950_b0 );
or ( \3952_b1 , \3361_b1 , \3899_b1 );
xor ( \3952_b0 , \3361_b0 , w_9136 );
not ( w_9136 , w_9137 );
and ( w_9137 , \3899_b1 , \3899_b0 );
buf ( \3953_Z[18]_b1 , \3952_b1 );
buf ( \3953_Z[18]_b0 , \3952_b0 );
or ( \3954_b1 , \3437_b1 , \3897_b1 );
xor ( \3954_b0 , \3437_b0 , w_9138 );
not ( w_9138 , w_9139 );
and ( w_9139 , \3897_b1 , \3897_b0 );
buf ( \3955_Z[17]_b1 , \3954_b1 );
buf ( \3955_Z[17]_b0 , \3954_b0 );
or ( \3956_b1 , \3490_b1 , \3895_b1 );
xor ( \3956_b0 , \3490_b0 , w_9140 );
not ( w_9140 , w_9141 );
and ( w_9141 , \3895_b1 , \3895_b0 );
buf ( \3957_Z[16]_b1 , \3956_b1 );
buf ( \3957_Z[16]_b0 , \3956_b0 );
or ( \3958_b1 , \3542_b1 , \3893_b1 );
xor ( \3958_b0 , \3542_b0 , w_9142 );
not ( w_9142 , w_9143 );
and ( w_9143 , \3893_b1 , \3893_b0 );
buf ( \3959_Z[15]_b1 , \3958_b1 );
buf ( \3959_Z[15]_b0 , \3958_b0 );
or ( \3960_b1 , \3575_b1 , \3891_b1 );
xor ( \3960_b0 , \3575_b0 , w_9144 );
not ( w_9144 , w_9145 );
and ( w_9145 , \3891_b1 , \3891_b0 );
buf ( \3961_Z[14]_b1 , \3960_b1 );
buf ( \3961_Z[14]_b0 , \3960_b0 );
or ( \3962_b1 , \3621_b1 , \3889_b1 );
xor ( \3962_b0 , \3621_b0 , w_9146 );
not ( w_9146 , w_9147 );
and ( w_9147 , \3889_b1 , \3889_b0 );
buf ( \3963_Z[13]_b1 , \3962_b1 );
buf ( \3963_Z[13]_b0 , \3962_b0 );
or ( \3964_b1 , \3663_b1 , \3887_b1 );
xor ( \3964_b0 , \3663_b0 , w_9148 );
not ( w_9148 , w_9149 );
and ( w_9149 , \3887_b1 , \3887_b0 );
buf ( \3965_Z[12]_b1 , \3964_b1 );
buf ( \3965_Z[12]_b0 , \3964_b0 );
or ( \3966_b1 , \3696_b1 , \3885_b1 );
xor ( \3966_b0 , \3696_b0 , w_9150 );
not ( w_9150 , w_9151 );
and ( w_9151 , \3885_b1 , \3885_b0 );
buf ( \3967_Z[11]_b1 , \3966_b1 );
buf ( \3967_Z[11]_b0 , \3966_b0 );
or ( \3968_b1 , \3728_b1 , \3883_b1 );
xor ( \3968_b0 , \3728_b0 , w_9152 );
not ( w_9152 , w_9153 );
and ( w_9153 , \3883_b1 , \3883_b0 );
buf ( \3969_Z[10]_b1 , \3968_b1 );
buf ( \3969_Z[10]_b0 , \3968_b0 );
or ( \3970_b1 , \3756_b1 , \3881_b1 );
xor ( \3970_b0 , \3756_b0 , w_9154 );
not ( w_9154 , w_9155 );
and ( w_9155 , \3881_b1 , \3881_b0 );
buf ( \3971_Z[9]_b1 , \3970_b1 );
buf ( \3971_Z[9]_b0 , \3970_b0 );
or ( \3972_b1 , \3779_b1 , \3879_b1 );
xor ( \3972_b0 , \3779_b0 , w_9156 );
not ( w_9156 , w_9157 );
and ( w_9157 , \3879_b1 , \3879_b0 );
buf ( \3973_Z[8]_b1 , \3972_b1 );
buf ( \3973_Z[8]_b0 , \3972_b0 );
or ( \3974_b1 , \3801_b1 , \3877_b1 );
xor ( \3974_b0 , \3801_b0 , w_9158 );
not ( w_9158 , w_9159 );
and ( w_9159 , \3877_b1 , \3877_b0 );
buf ( \3975_Z[7]_b1 , \3974_b1 );
buf ( \3975_Z[7]_b0 , \3974_b0 );
or ( \3976_b1 , \3818_b1 , \3875_b1 );
xor ( \3976_b0 , \3818_b0 , w_9160 );
not ( w_9160 , w_9161 );
and ( w_9161 , \3875_b1 , \3875_b0 );
buf ( \3977_Z[6]_b1 , \3976_b1 );
buf ( \3977_Z[6]_b0 , \3976_b0 );
or ( \3978_b1 , \3834_b1 , \3873_b1 );
xor ( \3978_b0 , \3834_b0 , w_9162 );
not ( w_9162 , w_9163 );
and ( w_9163 , \3873_b1 , \3873_b0 );
buf ( \3979_Z[5]_b1 , \3978_b1 );
buf ( \3979_Z[5]_b0 , \3978_b0 );
or ( \3980_b1 , \3846_b1 , \3871_b1 );
xor ( \3980_b0 , \3846_b0 , w_9164 );
not ( w_9164 , w_9165 );
and ( w_9165 , \3871_b1 , \3871_b0 );
buf ( \3981_Z[4]_b1 , \3980_b1 );
buf ( \3981_Z[4]_b0 , \3980_b0 );
or ( \3982_b1 , \3853_b1 , \3869_b1 );
xor ( \3982_b0 , \3853_b0 , w_9166 );
not ( w_9166 , w_9167 );
and ( w_9167 , \3869_b1 , \3869_b0 );
buf ( \3983_Z[3]_b1 , \3982_b1 );
buf ( \3983_Z[3]_b0 , \3982_b0 );
or ( \3984_b1 , \3859_b1 , \3867_b1 );
xor ( \3984_b0 , \3859_b0 , w_9168 );
not ( w_9168 , w_9169 );
and ( w_9169 , \3867_b1 , \3867_b0 );
buf ( \3985_Z[2]_b1 , \3984_b1 );
buf ( \3985_Z[2]_b0 , \3984_b0 );
or ( \3986_b1 , \3863_b1 , \3866_b1 );
xor ( \3986_b0 , \3863_b0 , w_9170 );
not ( w_9170 , w_9171 );
and ( w_9171 , \3866_b1 , \3866_b0 );
buf ( \3987_Z[1]_b1 , \3986_b1 );
buf ( \3987_Z[1]_b0 , \3986_b0 );
buf ( \3988_b1 , \3864_b1 );
buf ( \3988_b0 , \3864_b0 );
buf ( \3989_Z[0]_b1 , \3988_b1 );
buf ( \3989_Z[0]_b0 , \3988_b0 );
or ( \306_b1 , \303_b1 , w_9174 );
or ( \306_b0 , \303_b0 , w_9173 );
not ( w_9173 , w_9175 );
and ( w_9175 , w_9174 , w_9172 );
or ( w_9172 , \304_b1 , w_9176 );
or ( w_9173 , \304_b0 , \305_b0 );
not ( \305_b0 , w_9177 );
and ( w_9177 , w_9176 , \305_b1 );
or ( \316_b1 , \313_b1 , w_9180 );
or ( \316_b0 , \313_b0 , w_9179 );
not ( w_9179 , w_9181 );
and ( w_9181 , w_9180 , w_9178 );
or ( w_9178 , \314_b1 , w_9182 );
or ( w_9179 , \314_b0 , \315_b0 );
not ( \315_b0 , w_9183 );
and ( w_9183 , w_9182 , \315_b1 );
or ( \329_b1 , \326_b1 , w_9186 );
or ( \329_b0 , \326_b0 , w_9185 );
not ( w_9185 , w_9187 );
and ( w_9187 , w_9186 , w_9184 );
or ( w_9184 , \327_b1 , w_9188 );
or ( w_9185 , \327_b0 , \328_b0 );
not ( \328_b0 , w_9189 );
and ( w_9189 , w_9188 , \328_b1 );
or ( \339_b1 , \336_b1 , w_9192 );
or ( \339_b0 , \336_b0 , w_9191 );
not ( w_9191 , w_9193 );
and ( w_9193 , w_9192 , w_9190 );
or ( w_9190 , \337_b1 , w_9194 );
or ( w_9191 , \337_b0 , \338_b0 );
not ( \338_b0 , w_9195 );
and ( w_9195 , w_9194 , \338_b1 );
or ( \352_b1 , \349_b1 , w_9198 );
or ( \352_b0 , \349_b0 , w_9197 );
not ( w_9197 , w_9199 );
and ( w_9199 , w_9198 , w_9196 );
or ( w_9196 , \350_b1 , w_9200 );
or ( w_9197 , \350_b0 , \351_b0 );
not ( \351_b0 , w_9201 );
and ( w_9201 , w_9200 , \351_b1 );
or ( \362_b1 , \359_b1 , w_9204 );
or ( \362_b0 , \359_b0 , w_9203 );
not ( w_9203 , w_9205 );
and ( w_9205 , w_9204 , w_9202 );
or ( w_9202 , \360_b1 , w_9206 );
or ( w_9203 , \360_b0 , \361_b0 );
not ( \361_b0 , w_9207 );
and ( w_9207 , w_9206 , \361_b1 );
or ( \375_b1 , \372_b1 , w_9210 );
or ( \375_b0 , \372_b0 , w_9209 );
not ( w_9209 , w_9211 );
and ( w_9211 , w_9210 , w_9208 );
or ( w_9208 , \373_b1 , w_9212 );
or ( w_9209 , \373_b0 , \374_b0 );
not ( \374_b0 , w_9213 );
and ( w_9213 , w_9212 , \374_b1 );
or ( \385_b1 , \382_b1 , w_9216 );
or ( \385_b0 , \382_b0 , w_9215 );
not ( w_9215 , w_9217 );
and ( w_9217 , w_9216 , w_9214 );
or ( w_9214 , \383_b1 , w_9218 );
or ( w_9215 , \383_b0 , \384_b0 );
not ( \384_b0 , w_9219 );
and ( w_9219 , w_9218 , \384_b1 );
or ( \398_b1 , \395_b1 , w_9222 );
or ( \398_b0 , \395_b0 , w_9221 );
not ( w_9221 , w_9223 );
and ( w_9223 , w_9222 , w_9220 );
or ( w_9220 , \396_b1 , w_9224 );
or ( w_9221 , \396_b0 , \397_b0 );
not ( \397_b0 , w_9225 );
and ( w_9225 , w_9224 , \397_b1 );
or ( \408_b1 , \405_b1 , w_9228 );
or ( \408_b0 , \405_b0 , w_9227 );
not ( w_9227 , w_9229 );
and ( w_9229 , w_9228 , w_9226 );
or ( w_9226 , \406_b1 , w_9230 );
or ( w_9227 , \406_b0 , \407_b0 );
not ( \407_b0 , w_9231 );
and ( w_9231 , w_9230 , \407_b1 );
or ( \421_b1 , \418_b1 , w_9234 );
or ( \421_b0 , \418_b0 , w_9233 );
not ( w_9233 , w_9235 );
and ( w_9235 , w_9234 , w_9232 );
or ( w_9232 , \419_b1 , w_9236 );
or ( w_9233 , \419_b0 , \420_b0 );
not ( \420_b0 , w_9237 );
and ( w_9237 , w_9236 , \420_b1 );
or ( \431_b1 , \428_b1 , w_9240 );
or ( \431_b0 , \428_b0 , w_9239 );
not ( w_9239 , w_9241 );
and ( w_9241 , w_9240 , w_9238 );
or ( w_9238 , \429_b1 , w_9242 );
or ( w_9239 , \429_b0 , \430_b0 );
not ( \430_b0 , w_9243 );
and ( w_9243 , w_9242 , \430_b1 );
or ( \444_b1 , \441_b1 , w_9246 );
or ( \444_b0 , \441_b0 , w_9245 );
not ( w_9245 , w_9247 );
and ( w_9247 , w_9246 , w_9244 );
or ( w_9244 , \442_b1 , w_9248 );
or ( w_9245 , \442_b0 , \443_b0 );
not ( \443_b0 , w_9249 );
and ( w_9249 , w_9248 , \443_b1 );
or ( \454_b1 , \451_b1 , w_9252 );
or ( \454_b0 , \451_b0 , w_9251 );
not ( w_9251 , w_9253 );
and ( w_9253 , w_9252 , w_9250 );
or ( w_9250 , \452_b1 , w_9254 );
or ( w_9251 , \452_b0 , \453_b0 );
not ( \453_b0 , w_9255 );
and ( w_9255 , w_9254 , \453_b1 );
or ( \467_b1 , \464_b1 , w_9258 );
or ( \467_b0 , \464_b0 , w_9257 );
not ( w_9257 , w_9259 );
and ( w_9259 , w_9258 , w_9256 );
or ( w_9256 , \465_b1 , w_9260 );
or ( w_9257 , \465_b0 , \466_b0 );
not ( \466_b0 , w_9261 );
and ( w_9261 , w_9260 , \466_b1 );
or ( \477_b1 , \474_b1 , w_9264 );
or ( \477_b0 , \474_b0 , w_9263 );
not ( w_9263 , w_9265 );
and ( w_9265 , w_9264 , w_9262 );
or ( w_9262 , \475_b1 , w_9266 );
or ( w_9263 , \475_b0 , \476_b0 );
not ( \476_b0 , w_9267 );
and ( w_9267 , w_9266 , \476_b1 );
or ( \490_b1 , \487_b1 , w_9270 );
or ( \490_b0 , \487_b0 , w_9269 );
not ( w_9269 , w_9271 );
and ( w_9271 , w_9270 , w_9268 );
or ( w_9268 , \488_b1 , w_9272 );
or ( w_9269 , \488_b0 , \489_b0 );
not ( \489_b0 , w_9273 );
and ( w_9273 , w_9272 , \489_b1 );
or ( \500_b1 , \497_b1 , w_9276 );
or ( \500_b0 , \497_b0 , w_9275 );
not ( w_9275 , w_9277 );
and ( w_9277 , w_9276 , w_9274 );
or ( w_9274 , \498_b1 , w_9278 );
or ( w_9275 , \498_b0 , \499_b0 );
not ( \499_b0 , w_9279 );
and ( w_9279 , w_9278 , \499_b1 );
or ( \513_b1 , \510_b1 , w_9282 );
or ( \513_b0 , \510_b0 , w_9281 );
not ( w_9281 , w_9283 );
and ( w_9283 , w_9282 , w_9280 );
or ( w_9280 , \511_b1 , w_9284 );
or ( w_9281 , \511_b0 , \512_b0 );
not ( \512_b0 , w_9285 );
and ( w_9285 , w_9284 , \512_b1 );
or ( \523_b1 , \520_b1 , w_9288 );
or ( \523_b0 , \520_b0 , w_9287 );
not ( w_9287 , w_9289 );
and ( w_9289 , w_9288 , w_9286 );
or ( w_9286 , \521_b1 , w_9290 );
or ( w_9287 , \521_b0 , \522_b0 );
not ( \522_b0 , w_9291 );
and ( w_9291 , w_9290 , \522_b1 );
or ( \536_b1 , \533_b1 , w_9294 );
or ( \536_b0 , \533_b0 , w_9293 );
not ( w_9293 , w_9295 );
and ( w_9295 , w_9294 , w_9292 );
or ( w_9292 , \534_b1 , w_9296 );
or ( w_9293 , \534_b0 , \535_b0 );
not ( \535_b0 , w_9297 );
and ( w_9297 , w_9296 , \535_b1 );
or ( \546_b1 , \543_b1 , w_9300 );
or ( \546_b0 , \543_b0 , w_9299 );
not ( w_9299 , w_9301 );
and ( w_9301 , w_9300 , w_9298 );
or ( w_9298 , \544_b1 , w_9302 );
or ( w_9299 , \544_b0 , \545_b0 );
not ( \545_b0 , w_9303 );
and ( w_9303 , w_9302 , \545_b1 );
or ( \559_b1 , \556_b1 , w_9306 );
or ( \559_b0 , \556_b0 , w_9305 );
not ( w_9305 , w_9307 );
and ( w_9307 , w_9306 , w_9304 );
or ( w_9304 , \557_b1 , w_9308 );
or ( w_9305 , \557_b0 , \558_b0 );
not ( \558_b0 , w_9309 );
and ( w_9309 , w_9308 , \558_b1 );
or ( \569_b1 , \566_b1 , w_9312 );
or ( \569_b0 , \566_b0 , w_9311 );
not ( w_9311 , w_9313 );
and ( w_9313 , w_9312 , w_9310 );
or ( w_9310 , \567_b1 , w_9314 );
or ( w_9311 , \567_b0 , \568_b0 );
not ( \568_b0 , w_9315 );
and ( w_9315 , w_9314 , \568_b1 );
or ( \582_b1 , \579_b1 , w_9318 );
or ( \582_b0 , \579_b0 , w_9317 );
not ( w_9317 , w_9319 );
and ( w_9319 , w_9318 , w_9316 );
or ( w_9316 , \580_b1 , w_9320 );
or ( w_9317 , \580_b0 , \581_b0 );
not ( \581_b0 , w_9321 );
and ( w_9321 , w_9320 , \581_b1 );
or ( \592_b1 , \589_b1 , w_9324 );
or ( \592_b0 , \589_b0 , w_9323 );
not ( w_9323 , w_9325 );
and ( w_9325 , w_9324 , w_9322 );
or ( w_9322 , \590_b1 , w_9326 );
or ( w_9323 , \590_b0 , \591_b0 );
not ( \591_b0 , w_9327 );
and ( w_9327 , w_9326 , \591_b1 );
or ( \605_b1 , \602_b1 , w_9330 );
or ( \605_b0 , \602_b0 , w_9329 );
not ( w_9329 , w_9331 );
and ( w_9331 , w_9330 , w_9328 );
or ( w_9328 , \603_b1 , w_9332 );
or ( w_9329 , \603_b0 , \604_b0 );
not ( \604_b0 , w_9333 );
and ( w_9333 , w_9332 , \604_b1 );
or ( \615_b1 , \612_b1 , w_9336 );
or ( \615_b0 , \612_b0 , w_9335 );
not ( w_9335 , w_9337 );
and ( w_9337 , w_9336 , w_9334 );
or ( w_9334 , \613_b1 , w_9338 );
or ( w_9335 , \613_b0 , \614_b0 );
not ( \614_b0 , w_9339 );
and ( w_9339 , w_9338 , \614_b1 );
or ( \628_b1 , \625_b1 , w_9342 );
or ( \628_b0 , \625_b0 , w_9341 );
not ( w_9341 , w_9343 );
and ( w_9343 , w_9342 , w_9340 );
or ( w_9340 , \626_b1 , w_9344 );
or ( w_9341 , \626_b0 , \627_b0 );
not ( \627_b0 , w_9345 );
and ( w_9345 , w_9344 , \627_b1 );
or ( \638_b1 , \635_b1 , w_9348 );
or ( \638_b0 , \635_b0 , w_9347 );
not ( w_9347 , w_9349 );
and ( w_9349 , w_9348 , w_9346 );
or ( w_9346 , \636_b1 , w_9350 );
or ( w_9347 , \636_b0 , \637_b0 );
not ( \637_b0 , w_9351 );
and ( w_9351 , w_9350 , \637_b1 );
or ( \651_b1 , \648_b1 , w_9354 );
or ( \651_b0 , \648_b0 , w_9353 );
not ( w_9353 , w_9355 );
and ( w_9355 , w_9354 , w_9352 );
or ( w_9352 , \649_b1 , w_9356 );
or ( w_9353 , \649_b0 , \650_b0 );
not ( \650_b0 , w_9357 );
and ( w_9357 , w_9356 , \650_b1 );
or ( \661_b1 , \658_b1 , w_9360 );
or ( \661_b0 , \658_b0 , w_9359 );
not ( w_9359 , w_9361 );
and ( w_9361 , w_9360 , w_9358 );
or ( w_9358 , \659_b1 , w_9362 );
or ( w_9359 , \659_b0 , \660_b0 );
not ( \660_b0 , w_9363 );
and ( w_9363 , w_9362 , \660_b1 );
or ( \674_b1 , \671_b1 , w_9366 );
or ( \674_b0 , \671_b0 , w_9365 );
not ( w_9365 , w_9367 );
and ( w_9367 , w_9366 , w_9364 );
or ( w_9364 , \672_b1 , w_9368 );
or ( w_9365 , \672_b0 , \673_b0 );
not ( \673_b0 , w_9369 );
and ( w_9369 , w_9368 , \673_b1 );
or ( \684_b1 , \681_b1 , w_9372 );
or ( \684_b0 , \681_b0 , w_9371 );
not ( w_9371 , w_9373 );
and ( w_9373 , w_9372 , w_9370 );
or ( w_9370 , \682_b1 , w_9374 );
or ( w_9371 , \682_b0 , \683_b0 );
not ( \683_b0 , w_9375 );
and ( w_9375 , w_9374 , \683_b1 );
or ( \697_b1 , \694_b1 , w_9378 );
or ( \697_b0 , \694_b0 , w_9377 );
not ( w_9377 , w_9379 );
and ( w_9379 , w_9378 , w_9376 );
or ( w_9376 , \695_b1 , w_9380 );
or ( w_9377 , \695_b0 , \696_b0 );
not ( \696_b0 , w_9381 );
and ( w_9381 , w_9380 , \696_b1 );
or ( \707_b1 , \704_b1 , w_9384 );
or ( \707_b0 , \704_b0 , w_9383 );
not ( w_9383 , w_9385 );
and ( w_9385 , w_9384 , w_9382 );
or ( w_9382 , \705_b1 , w_9386 );
or ( w_9383 , \705_b0 , \706_b0 );
not ( \706_b0 , w_9387 );
and ( w_9387 , w_9386 , \706_b1 );
or ( \720_b1 , \717_b1 , w_9390 );
or ( \720_b0 , \717_b0 , w_9389 );
not ( w_9389 , w_9391 );
and ( w_9391 , w_9390 , w_9388 );
or ( w_9388 , \718_b1 , w_9392 );
or ( w_9389 , \718_b0 , \719_b0 );
not ( \719_b0 , w_9393 );
and ( w_9393 , w_9392 , \719_b1 );
or ( \730_b1 , \727_b1 , w_9396 );
or ( \730_b0 , \727_b0 , w_9395 );
not ( w_9395 , w_9397 );
and ( w_9397 , w_9396 , w_9394 );
or ( w_9394 , \728_b1 , w_9398 );
or ( w_9395 , \728_b0 , \729_b0 );
not ( \729_b0 , w_9399 );
and ( w_9399 , w_9398 , \729_b1 );
or ( \743_b1 , \740_b1 , w_9402 );
or ( \743_b0 , \740_b0 , w_9401 );
not ( w_9401 , w_9403 );
and ( w_9403 , w_9402 , w_9400 );
or ( w_9400 , \741_b1 , w_9404 );
or ( w_9401 , \741_b0 , \742_b0 );
not ( \742_b0 , w_9405 );
and ( w_9405 , w_9404 , \742_b1 );
or ( \753_b1 , \750_b1 , w_9408 );
or ( \753_b0 , \750_b0 , w_9407 );
not ( w_9407 , w_9409 );
and ( w_9409 , w_9408 , w_9406 );
or ( w_9406 , \751_b1 , w_9410 );
or ( w_9407 , \751_b0 , \752_b0 );
not ( \752_b0 , w_9411 );
and ( w_9411 , w_9410 , \752_b1 );
or ( \766_b1 , \763_b1 , w_9414 );
or ( \766_b0 , \763_b0 , w_9413 );
not ( w_9413 , w_9415 );
and ( w_9415 , w_9414 , w_9412 );
or ( w_9412 , \764_b1 , w_9416 );
or ( w_9413 , \764_b0 , \765_b0 );
not ( \765_b0 , w_9417 );
and ( w_9417 , w_9416 , \765_b1 );
or ( \776_b1 , \773_b1 , w_9420 );
or ( \776_b0 , \773_b0 , w_9419 );
not ( w_9419 , w_9421 );
and ( w_9421 , w_9420 , w_9418 );
or ( w_9418 , \774_b1 , w_9422 );
or ( w_9419 , \774_b0 , \775_b0 );
not ( \775_b0 , w_9423 );
and ( w_9423 , w_9422 , \775_b1 );
or ( \789_b1 , \786_b1 , w_9426 );
or ( \789_b0 , \786_b0 , w_9425 );
not ( w_9425 , w_9427 );
and ( w_9427 , w_9426 , w_9424 );
or ( w_9424 , \787_b1 , w_9428 );
or ( w_9425 , \787_b0 , \788_b0 );
not ( \788_b0 , w_9429 );
and ( w_9429 , w_9428 , \788_b1 );
or ( \799_b1 , \796_b1 , w_9432 );
or ( \799_b0 , \796_b0 , w_9431 );
not ( w_9431 , w_9433 );
and ( w_9433 , w_9432 , w_9430 );
or ( w_9430 , \797_b1 , w_9434 );
or ( w_9431 , \797_b0 , \798_b0 );
not ( \798_b0 , w_9435 );
and ( w_9435 , w_9434 , \798_b1 );
or ( \812_b1 , \809_b1 , w_9438 );
or ( \812_b0 , \809_b0 , w_9437 );
not ( w_9437 , w_9439 );
and ( w_9439 , w_9438 , w_9436 );
or ( w_9436 , \810_b1 , w_9440 );
or ( w_9437 , \810_b0 , \811_b0 );
not ( \811_b0 , w_9441 );
and ( w_9441 , w_9440 , \811_b1 );
or ( \822_b1 , \819_b1 , w_9444 );
or ( \822_b0 , \819_b0 , w_9443 );
not ( w_9443 , w_9445 );
and ( w_9445 , w_9444 , w_9442 );
or ( w_9442 , \820_b1 , w_9446 );
or ( w_9443 , \820_b0 , \821_b0 );
not ( \821_b0 , w_9447 );
and ( w_9447 , w_9446 , \821_b1 );
or ( \835_b1 , \832_b1 , w_9450 );
or ( \835_b0 , \832_b0 , w_9449 );
not ( w_9449 , w_9451 );
and ( w_9451 , w_9450 , w_9448 );
or ( w_9448 , \833_b1 , w_9452 );
or ( w_9449 , \833_b0 , \834_b0 );
not ( \834_b0 , w_9453 );
and ( w_9453 , w_9452 , \834_b1 );
or ( \845_b1 , \842_b1 , w_9456 );
or ( \845_b0 , \842_b0 , w_9455 );
not ( w_9455 , w_9457 );
and ( w_9457 , w_9456 , w_9454 );
or ( w_9454 , \843_b1 , w_9458 );
or ( w_9455 , \843_b0 , \844_b0 );
not ( \844_b0 , w_9459 );
and ( w_9459 , w_9458 , \844_b1 );
or ( \858_b1 , \855_b1 , w_9462 );
or ( \858_b0 , \855_b0 , w_9461 );
not ( w_9461 , w_9463 );
and ( w_9463 , w_9462 , w_9460 );
or ( w_9460 , \856_b1 , w_9464 );
or ( w_9461 , \856_b0 , \857_b0 );
not ( \857_b0 , w_9465 );
and ( w_9465 , w_9464 , \857_b1 );
or ( \868_b1 , \865_b1 , w_9468 );
or ( \868_b0 , \865_b0 , w_9467 );
not ( w_9467 , w_9469 );
and ( w_9469 , w_9468 , w_9466 );
or ( w_9466 , \866_b1 , w_9470 );
or ( w_9467 , \866_b0 , \867_b0 );
not ( \867_b0 , w_9471 );
and ( w_9471 , w_9470 , \867_b1 );
or ( \881_b1 , \878_b1 , w_9474 );
or ( \881_b0 , \878_b0 , w_9473 );
not ( w_9473 , w_9475 );
and ( w_9475 , w_9474 , w_9472 );
or ( w_9472 , \879_b1 , w_9476 );
or ( w_9473 , \879_b0 , \880_b0 );
not ( \880_b0 , w_9477 );
and ( w_9477 , w_9476 , \880_b1 );
or ( \891_b1 , \888_b1 , w_9480 );
or ( \891_b0 , \888_b0 , w_9479 );
not ( w_9479 , w_9481 );
and ( w_9481 , w_9480 , w_9478 );
or ( w_9478 , \889_b1 , w_9482 );
or ( w_9479 , \889_b0 , \890_b0 );
not ( \890_b0 , w_9483 );
and ( w_9483 , w_9482 , \890_b1 );
or ( \904_b1 , \901_b1 , w_9486 );
or ( \904_b0 , \901_b0 , w_9485 );
not ( w_9485 , w_9487 );
and ( w_9487 , w_9486 , w_9484 );
or ( w_9484 , \902_b1 , w_9488 );
or ( w_9485 , \902_b0 , \903_b0 );
not ( \903_b0 , w_9489 );
and ( w_9489 , w_9488 , \903_b1 );
or ( \914_b1 , \911_b1 , w_9492 );
or ( \914_b0 , \911_b0 , w_9491 );
not ( w_9491 , w_9493 );
and ( w_9493 , w_9492 , w_9490 );
or ( w_9490 , \912_b1 , w_9494 );
or ( w_9491 , \912_b0 , \913_b0 );
not ( \913_b0 , w_9495 );
and ( w_9495 , w_9494 , \913_b1 );
or ( \927_b1 , \924_b1 , w_9498 );
or ( \927_b0 , \924_b0 , w_9497 );
not ( w_9497 , w_9499 );
and ( w_9499 , w_9498 , w_9496 );
or ( w_9496 , \925_b1 , w_9500 );
or ( w_9497 , \925_b0 , \926_b0 );
not ( \926_b0 , w_9501 );
and ( w_9501 , w_9500 , \926_b1 );
or ( \937_b1 , \934_b1 , w_9504 );
or ( \937_b0 , \934_b0 , w_9503 );
not ( w_9503 , w_9505 );
and ( w_9505 , w_9504 , w_9502 );
or ( w_9502 , \935_b1 , w_9506 );
or ( w_9503 , \935_b0 , \936_b0 );
not ( \936_b0 , w_9507 );
and ( w_9507 , w_9506 , \936_b1 );
or ( \950_b1 , \947_b1 , w_9510 );
or ( \950_b0 , \947_b0 , w_9509 );
not ( w_9509 , w_9511 );
and ( w_9511 , w_9510 , w_9508 );
or ( w_9508 , \948_b1 , w_9512 );
or ( w_9509 , \948_b0 , \949_b0 );
not ( \949_b0 , w_9513 );
and ( w_9513 , w_9512 , \949_b1 );
or ( \960_b1 , \957_b1 , w_9516 );
or ( \960_b0 , \957_b0 , w_9515 );
not ( w_9515 , w_9517 );
and ( w_9517 , w_9516 , w_9514 );
or ( w_9514 , \958_b1 , w_9518 );
or ( w_9515 , \958_b0 , \959_b0 );
not ( \959_b0 , w_9519 );
and ( w_9519 , w_9518 , \959_b1 );
or ( \973_b1 , \970_b1 , w_9522 );
or ( \973_b0 , \970_b0 , w_9521 );
not ( w_9521 , w_9523 );
and ( w_9523 , w_9522 , w_9520 );
or ( w_9520 , \971_b1 , w_9524 );
or ( w_9521 , \971_b0 , \972_b0 );
not ( \972_b0 , w_9525 );
and ( w_9525 , w_9524 , \972_b1 );
or ( \983_b1 , \980_b1 , w_9528 );
or ( \983_b0 , \980_b0 , w_9527 );
not ( w_9527 , w_9529 );
and ( w_9529 , w_9528 , w_9526 );
or ( w_9526 , \981_b1 , w_9530 );
or ( w_9527 , \981_b0 , \982_b0 );
not ( \982_b0 , w_9531 );
and ( w_9531 , w_9530 , \982_b1 );
or ( \1085_b1 , \1079_b1 , w_9534 );
or ( \1085_b0 , \1079_b0 , w_9533 );
not ( w_9533 , w_9535 );
and ( w_9535 , w_9534 , w_9532 );
or ( w_9532 , \1083_b1 , w_9536 );
or ( w_9533 , \1083_b0 , \1084_b0 );
not ( \1084_b0 , w_9537 );
and ( w_9537 , w_9536 , \1084_b1 );
or ( \1088_b1 , \1076_b1 , w_9540 );
or ( \1088_b0 , \1076_b0 , w_9539 );
not ( w_9539 , w_9541 );
and ( w_9541 , w_9540 , w_9538 );
or ( w_9538 , \1086_b1 , w_9542 );
or ( w_9539 , \1086_b0 , \1087_b0 );
not ( \1087_b0 , w_9543 );
and ( w_9543 , w_9542 , \1087_b1 );
or ( \1091_b1 , \1073_b1 , w_9546 );
or ( \1091_b0 , \1073_b0 , w_9545 );
not ( w_9545 , w_9547 );
and ( w_9547 , w_9546 , w_9544 );
or ( w_9544 , \1089_b1 , w_9548 );
or ( w_9545 , \1089_b0 , \1090_b0 );
not ( \1090_b0 , w_9549 );
and ( w_9549 , w_9548 , \1090_b1 );
or ( \1094_b1 , \1070_b1 , w_9552 );
or ( \1094_b0 , \1070_b0 , w_9551 );
not ( w_9551 , w_9553 );
and ( w_9553 , w_9552 , w_9550 );
or ( w_9550 , \1092_b1 , w_9554 );
or ( w_9551 , \1092_b0 , \1093_b0 );
not ( \1093_b0 , w_9555 );
and ( w_9555 , w_9554 , \1093_b1 );
or ( \1097_b1 , \1067_b1 , w_9558 );
or ( \1097_b0 , \1067_b0 , w_9557 );
not ( w_9557 , w_9559 );
and ( w_9559 , w_9558 , w_9556 );
or ( w_9556 , \1095_b1 , w_9560 );
or ( w_9557 , \1095_b0 , \1096_b0 );
not ( \1096_b0 , w_9561 );
and ( w_9561 , w_9560 , \1096_b1 );
or ( \1100_b1 , \1064_b1 , w_9564 );
or ( \1100_b0 , \1064_b0 , w_9563 );
not ( w_9563 , w_9565 );
and ( w_9565 , w_9564 , w_9562 );
or ( w_9562 , \1098_b1 , w_9566 );
or ( w_9563 , \1098_b0 , \1099_b0 );
not ( \1099_b0 , w_9567 );
and ( w_9567 , w_9566 , \1099_b1 );
or ( \1103_b1 , \1061_b1 , w_9570 );
or ( \1103_b0 , \1061_b0 , w_9569 );
not ( w_9569 , w_9571 );
and ( w_9571 , w_9570 , w_9568 );
or ( w_9568 , \1101_b1 , w_9572 );
or ( w_9569 , \1101_b0 , \1102_b0 );
not ( \1102_b0 , w_9573 );
and ( w_9573 , w_9572 , \1102_b1 );
or ( \1106_b1 , \1058_b1 , w_9576 );
or ( \1106_b0 , \1058_b0 , w_9575 );
not ( w_9575 , w_9577 );
and ( w_9577 , w_9576 , w_9574 );
or ( w_9574 , \1104_b1 , w_9578 );
or ( w_9575 , \1104_b0 , \1105_b0 );
not ( \1105_b0 , w_9579 );
and ( w_9579 , w_9578 , \1105_b1 );
or ( \1109_b1 , \1055_b1 , w_9582 );
or ( \1109_b0 , \1055_b0 , w_9581 );
not ( w_9581 , w_9583 );
and ( w_9583 , w_9582 , w_9580 );
or ( w_9580 , \1107_b1 , w_9584 );
or ( w_9581 , \1107_b0 , \1108_b0 );
not ( \1108_b0 , w_9585 );
and ( w_9585 , w_9584 , \1108_b1 );
or ( \1112_b1 , \1052_b1 , w_9588 );
or ( \1112_b0 , \1052_b0 , w_9587 );
not ( w_9587 , w_9589 );
and ( w_9589 , w_9588 , w_9586 );
or ( w_9586 , \1110_b1 , w_9590 );
or ( w_9587 , \1110_b0 , \1111_b0 );
not ( \1111_b0 , w_9591 );
and ( w_9591 , w_9590 , \1111_b1 );
or ( \1115_b1 , \1049_b1 , w_9594 );
or ( \1115_b0 , \1049_b0 , w_9593 );
not ( w_9593 , w_9595 );
and ( w_9595 , w_9594 , w_9592 );
or ( w_9592 , \1113_b1 , w_9596 );
or ( w_9593 , \1113_b0 , \1114_b0 );
not ( \1114_b0 , w_9597 );
and ( w_9597 , w_9596 , \1114_b1 );
or ( \1118_b1 , \1046_b1 , w_9600 );
or ( \1118_b0 , \1046_b0 , w_9599 );
not ( w_9599 , w_9601 );
and ( w_9601 , w_9600 , w_9598 );
or ( w_9598 , \1116_b1 , w_9602 );
or ( w_9599 , \1116_b0 , \1117_b0 );
not ( \1117_b0 , w_9603 );
and ( w_9603 , w_9602 , \1117_b1 );
or ( \1121_b1 , \1043_b1 , w_9606 );
or ( \1121_b0 , \1043_b0 , w_9605 );
not ( w_9605 , w_9607 );
and ( w_9607 , w_9606 , w_9604 );
or ( w_9604 , \1119_b1 , w_9608 );
or ( w_9605 , \1119_b0 , \1120_b0 );
not ( \1120_b0 , w_9609 );
and ( w_9609 , w_9608 , \1120_b1 );
or ( \1124_b1 , \1040_b1 , w_9612 );
or ( \1124_b0 , \1040_b0 , w_9611 );
not ( w_9611 , w_9613 );
and ( w_9613 , w_9612 , w_9610 );
or ( w_9610 , \1122_b1 , w_9614 );
or ( w_9611 , \1122_b0 , \1123_b0 );
not ( \1123_b0 , w_9615 );
and ( w_9615 , w_9614 , \1123_b1 );
or ( \1127_b1 , \1037_b1 , w_9618 );
or ( \1127_b0 , \1037_b0 , w_9617 );
not ( w_9617 , w_9619 );
and ( w_9619 , w_9618 , w_9616 );
or ( w_9616 , \1125_b1 , w_9620 );
or ( w_9617 , \1125_b0 , \1126_b0 );
not ( \1126_b0 , w_9621 );
and ( w_9621 , w_9620 , \1126_b1 );
or ( \1130_b1 , \1034_b1 , w_9624 );
or ( \1130_b0 , \1034_b0 , w_9623 );
not ( w_9623 , w_9625 );
and ( w_9625 , w_9624 , w_9622 );
or ( w_9622 , \1128_b1 , w_9626 );
or ( w_9623 , \1128_b0 , \1129_b0 );
not ( \1129_b0 , w_9627 );
and ( w_9627 , w_9626 , \1129_b1 );
or ( \1133_b1 , \1031_b1 , w_9630 );
or ( \1133_b0 , \1031_b0 , w_9629 );
not ( w_9629 , w_9631 );
and ( w_9631 , w_9630 , w_9628 );
or ( w_9628 , \1131_b1 , w_9632 );
or ( w_9629 , \1131_b0 , \1132_b0 );
not ( \1132_b0 , w_9633 );
and ( w_9633 , w_9632 , \1132_b1 );
or ( \1136_b1 , \1028_b1 , w_9636 );
or ( \1136_b0 , \1028_b0 , w_9635 );
not ( w_9635 , w_9637 );
and ( w_9637 , w_9636 , w_9634 );
or ( w_9634 , \1134_b1 , w_9638 );
or ( w_9635 , \1134_b0 , \1135_b0 );
not ( \1135_b0 , w_9639 );
and ( w_9639 , w_9638 , \1135_b1 );
or ( \1139_b1 , \1025_b1 , w_9642 );
or ( \1139_b0 , \1025_b0 , w_9641 );
not ( w_9641 , w_9643 );
and ( w_9643 , w_9642 , w_9640 );
or ( w_9640 , \1137_b1 , w_9644 );
or ( w_9641 , \1137_b0 , \1138_b0 );
not ( \1138_b0 , w_9645 );
and ( w_9645 , w_9644 , \1138_b1 );
or ( \1142_b1 , \1022_b1 , w_9648 );
or ( \1142_b0 , \1022_b0 , w_9647 );
not ( w_9647 , w_9649 );
and ( w_9649 , w_9648 , w_9646 );
or ( w_9646 , \1140_b1 , w_9650 );
or ( w_9647 , \1140_b0 , \1141_b0 );
not ( \1141_b0 , w_9651 );
and ( w_9651 , w_9650 , \1141_b1 );
or ( \1145_b1 , \1019_b1 , w_9654 );
or ( \1145_b0 , \1019_b0 , w_9653 );
not ( w_9653 , w_9655 );
and ( w_9655 , w_9654 , w_9652 );
or ( w_9652 , \1143_b1 , w_9656 );
or ( w_9653 , \1143_b0 , \1144_b0 );
not ( \1144_b0 , w_9657 );
and ( w_9657 , w_9656 , \1144_b1 );
or ( \1148_b1 , \1016_b1 , w_9660 );
or ( \1148_b0 , \1016_b0 , w_9659 );
not ( w_9659 , w_9661 );
and ( w_9661 , w_9660 , w_9658 );
or ( w_9658 , \1146_b1 , w_9662 );
or ( w_9659 , \1146_b0 , \1147_b0 );
not ( \1147_b0 , w_9663 );
and ( w_9663 , w_9662 , \1147_b1 );
or ( \1151_b1 , \1013_b1 , w_9666 );
or ( \1151_b0 , \1013_b0 , w_9665 );
not ( w_9665 , w_9667 );
and ( w_9667 , w_9666 , w_9664 );
or ( w_9664 , \1149_b1 , w_9668 );
or ( w_9665 , \1149_b0 , \1150_b0 );
not ( \1150_b0 , w_9669 );
and ( w_9669 , w_9668 , \1150_b1 );
or ( \1154_b1 , \1010_b1 , w_9672 );
or ( \1154_b0 , \1010_b0 , w_9671 );
not ( w_9671 , w_9673 );
and ( w_9673 , w_9672 , w_9670 );
or ( w_9670 , \1152_b1 , w_9674 );
or ( w_9671 , \1152_b0 , \1153_b0 );
not ( \1153_b0 , w_9675 );
and ( w_9675 , w_9674 , \1153_b1 );
or ( \1157_b1 , \1007_b1 , w_9678 );
or ( \1157_b0 , \1007_b0 , w_9677 );
not ( w_9677 , w_9679 );
and ( w_9679 , w_9678 , w_9676 );
or ( w_9676 , \1155_b1 , w_9680 );
or ( w_9677 , \1155_b0 , \1156_b0 );
not ( \1156_b0 , w_9681 );
and ( w_9681 , w_9680 , \1156_b1 );
or ( \1160_b1 , \1004_b1 , w_9684 );
or ( \1160_b0 , \1004_b0 , w_9683 );
not ( w_9683 , w_9685 );
and ( w_9685 , w_9684 , w_9682 );
or ( w_9682 , \1158_b1 , w_9686 );
or ( w_9683 , \1158_b0 , \1159_b0 );
not ( \1159_b0 , w_9687 );
and ( w_9687 , w_9686 , \1159_b1 );
or ( \1163_b1 , \1001_b1 , w_9690 );
or ( \1163_b0 , \1001_b0 , w_9689 );
not ( w_9689 , w_9691 );
and ( w_9691 , w_9690 , w_9688 );
or ( w_9688 , \1161_b1 , w_9692 );
or ( w_9689 , \1161_b0 , \1162_b0 );
not ( \1162_b0 , w_9693 );
and ( w_9693 , w_9692 , \1162_b1 );
or ( \1166_b1 , \998_b1 , w_9696 );
or ( \1166_b0 , \998_b0 , w_9695 );
not ( w_9695 , w_9697 );
and ( w_9697 , w_9696 , w_9694 );
or ( w_9694 , \1164_b1 , w_9698 );
or ( w_9695 , \1164_b0 , \1165_b0 );
not ( \1165_b0 , w_9699 );
and ( w_9699 , w_9698 , \1165_b1 );
or ( \1169_b1 , \995_b1 , w_9702 );
or ( \1169_b0 , \995_b0 , w_9701 );
not ( w_9701 , w_9703 );
and ( w_9703 , w_9702 , w_9700 );
or ( w_9700 , \1167_b1 , w_9704 );
or ( w_9701 , \1167_b0 , \1168_b0 );
not ( \1168_b0 , w_9705 );
and ( w_9705 , w_9704 , \1168_b1 );
or ( \1172_b1 , \992_b1 , w_9708 );
or ( \1172_b0 , \992_b0 , w_9707 );
not ( w_9707 , w_9709 );
and ( w_9709 , w_9708 , w_9706 );
or ( w_9706 , \1170_b1 , w_9710 );
or ( w_9707 , \1170_b0 , \1171_b0 );
not ( \1171_b0 , w_9711 );
and ( w_9711 , w_9710 , \1171_b1 );
or ( \1487_b1 , \1424_b1 , w_9714 );
or ( \1487_b0 , \1424_b0 , w_9713 );
not ( w_9713 , w_9715 );
and ( w_9715 , w_9714 , w_9712 );
or ( w_9712 , \1485_b1 , w_9716 );
or ( w_9713 , \1485_b0 , \1486_b0 );
not ( \1486_b0 , w_9717 );
and ( w_9717 , w_9716 , \1486_b1 );
or ( \1505_b1 , \1497_b1 , w_9720 );
or ( \1505_b0 , \1497_b0 , w_9719 );
not ( w_9719 , w_9721 );
and ( w_9721 , w_9720 , w_9718 );
or ( w_9718 , \1503_b1 , w_9722 );
or ( w_9719 , \1503_b0 , \1504_b0 );
not ( \1504_b0 , w_9723 );
and ( w_9723 , w_9722 , \1504_b1 );
or ( \1509_b1 , \1506_b1 , w_9726 );
or ( \1509_b0 , \1506_b0 , w_9725 );
not ( w_9725 , w_9727 );
and ( w_9727 , w_9726 , w_9724 );
or ( w_9724 , \1507_b1 , w_9728 );
or ( w_9725 , \1507_b0 , \1508_b0 );
not ( \1508_b0 , w_9729 );
and ( w_9729 , w_9728 , \1508_b1 );
or ( \1514_b1 , \1511_b1 , w_9732 );
or ( \1514_b0 , \1511_b0 , w_9731 );
not ( w_9731 , w_9733 );
and ( w_9733 , w_9732 , w_9730 );
or ( w_9730 , \1512_b1 , w_9734 );
or ( w_9731 , \1512_b0 , \1513_b0 );
not ( \1513_b0 , w_9735 );
and ( w_9735 , w_9734 , \1513_b1 );
or ( \1594_b1 , \1516_b1 , w_9738 );
or ( \1594_b0 , \1516_b0 , w_9737 );
not ( w_9737 , w_9739 );
and ( w_9739 , w_9738 , w_9736 );
or ( w_9736 , \1592_b1 , w_9740 );
or ( w_9737 , \1592_b0 , \1593_b0 );
not ( \1593_b0 , w_9741 );
and ( w_9741 , w_9740 , \1593_b1 );
or ( \1610_b1 , \1603_b1 , w_9744 );
or ( \1610_b0 , \1603_b0 , w_9743 );
not ( w_9743 , w_9745 );
and ( w_9745 , w_9744 , w_9742 );
or ( w_9742 , \1608_b1 , w_9746 );
or ( w_9743 , \1608_b0 , \1609_b0 );
not ( \1609_b0 , w_9747 );
and ( w_9747 , w_9746 , \1609_b1 );
or ( \1628_b1 , \1620_b1 , w_9750 );
or ( \1628_b0 , \1620_b0 , w_9749 );
not ( w_9749 , w_9751 );
and ( w_9751 , w_9750 , w_9748 );
or ( w_9748 , \1626_b1 , w_9752 );
or ( w_9749 , \1626_b0 , \1627_b0 );
not ( \1627_b0 , w_9753 );
and ( w_9753 , w_9752 , \1627_b1 );
or ( \1658_b1 , \1651_b1 , w_9756 );
or ( \1658_b0 , \1651_b0 , w_9755 );
not ( w_9755 , w_9757 );
and ( w_9757 , w_9756 , w_9754 );
or ( w_9754 , \1656_b1 , w_9758 );
or ( w_9755 , \1656_b0 , \1657_b0 );
not ( \1657_b0 , w_9759 );
and ( w_9759 , w_9758 , \1657_b1 );
or ( \1661_b1 , \1629_b1 , w_9762 );
or ( \1661_b0 , \1629_b0 , w_9761 );
not ( w_9761 , w_9763 );
and ( w_9763 , w_9762 , w_9760 );
or ( w_9760 , \1659_b1 , w_9764 );
or ( w_9761 , \1659_b0 , \1660_b0 );
not ( \1660_b0 , w_9765 );
and ( w_9765 , w_9764 , \1660_b1 );
or ( \1685_b1 , \1670_b1 , w_9768 );
or ( \1685_b0 , \1670_b0 , w_9767 );
not ( w_9767 , w_9769 );
and ( w_9769 , w_9768 , w_9766 );
or ( w_9766 , \1683_b1 , w_9770 );
or ( w_9767 , \1683_b0 , \1684_b0 );
not ( \1684_b0 , w_9771 );
and ( w_9771 , w_9770 , \1684_b1 );
or ( \1717_b1 , \1700_b1 , w_9774 );
or ( \1717_b0 , \1700_b0 , w_9773 );
not ( w_9773 , w_9775 );
and ( w_9775 , w_9774 , w_9772 );
or ( w_9772 , \1715_b1 , w_9776 );
or ( w_9773 , \1715_b0 , \1716_b0 );
not ( \1716_b0 , w_9777 );
and ( w_9777 , w_9776 , \1716_b1 );
or ( \1722_b1 , \1719_b1 , w_9780 );
or ( \1722_b0 , \1719_b0 , w_9779 );
not ( w_9779 , w_9781 );
and ( w_9781 , w_9780 , w_9778 );
or ( w_9778 , \1720_b1 , w_9782 );
or ( w_9779 , \1720_b0 , \1721_b0 );
not ( \1721_b0 , w_9783 );
and ( w_9783 , w_9782 , \1721_b1 );
or ( \1726_b1 , \1723_b1 , w_9786 );
or ( \1726_b0 , \1723_b0 , w_9785 );
not ( w_9785 , w_9787 );
and ( w_9787 , w_9786 , w_9784 );
or ( w_9784 , \1724_b1 , w_9788 );
or ( w_9785 , \1724_b0 , \1725_b0 );
not ( \1725_b0 , w_9789 );
and ( w_9789 , w_9788 , \1725_b1 );
or ( \1740_b1 , \1733_b1 , w_9792 );
or ( \1740_b0 , \1733_b0 , w_9791 );
not ( w_9791 , w_9793 );
and ( w_9793 , w_9792 , w_9790 );
or ( w_9790 , \1738_b1 , w_9794 );
or ( w_9791 , \1738_b0 , \1739_b0 );
not ( \1739_b0 , w_9795 );
and ( w_9795 , w_9794 , \1739_b1 );
or ( \1744_b1 , \1718_b1 , w_9798 );
or ( \1744_b0 , \1718_b0 , w_9797 );
not ( w_9797 , w_9799 );
and ( w_9799 , w_9798 , w_9796 );
or ( w_9796 , \1742_b1 , w_9800 );
or ( w_9797 , \1742_b0 , \1743_b0 );
not ( \1743_b0 , w_9801 );
and ( w_9801 , w_9800 , \1743_b1 );
or ( \1757_b1 , \1753_b1 , w_9804 );
or ( \1757_b0 , \1753_b0 , w_9803 );
not ( w_9803 , w_9805 );
and ( w_9805 , w_9804 , w_9802 );
or ( w_9802 , \1755_b1 , w_9806 );
or ( w_9803 , \1755_b0 , \1756_b0 );
not ( \1756_b0 , w_9807 );
and ( w_9807 , w_9806 , \1756_b1 );
or ( \1769_b1 , \1762_b1 , w_9810 );
or ( \1769_b0 , \1762_b0 , w_9809 );
not ( w_9809 , w_9811 );
and ( w_9811 , w_9810 , w_9808 );
or ( w_9808 , \1767_b1 , w_9812 );
or ( w_9809 , \1767_b0 , \1768_b0 );
not ( \1768_b0 , w_9813 );
and ( w_9813 , w_9812 , \1768_b1 );
or ( \1798_b1 , \1793_b1 , w_9816 );
or ( \1798_b0 , \1793_b0 , w_9815 );
not ( w_9815 , w_9817 );
and ( w_9817 , w_9816 , w_9814 );
or ( w_9814 , \1796_b1 , w_9818 );
or ( w_9815 , \1796_b0 , \1797_b0 );
not ( \1797_b0 , w_9819 );
and ( w_9819 , w_9818 , \1797_b1 );
or ( \1809_b1 , \1784_b1 , w_9822 );
or ( \1809_b0 , \1784_b0 , w_9821 );
not ( w_9821 , w_9823 );
and ( w_9823 , w_9822 , w_9820 );
or ( w_9820 , \1807_b1 , w_9824 );
or ( w_9821 , \1807_b0 , \1808_b0 );
not ( \1808_b0 , w_9825 );
and ( w_9825 , w_9824 , \1808_b1 );
or ( \1814_b1 , \1811_b1 , w_9828 );
or ( \1814_b0 , \1811_b0 , w_9827 );
not ( w_9827 , w_9829 );
and ( w_9829 , w_9828 , w_9826 );
or ( w_9826 , \1812_b1 , w_9830 );
or ( w_9827 , \1812_b0 , \1813_b0 );
not ( \1813_b0 , w_9831 );
and ( w_9831 , w_9830 , \1813_b1 );
or ( \1818_b1 , \1815_b1 , w_9834 );
or ( \1818_b0 , \1815_b0 , w_9833 );
not ( w_9833 , w_9835 );
and ( w_9835 , w_9834 , w_9832 );
or ( w_9832 , \1816_b1 , w_9836 );
or ( w_9833 , \1816_b0 , \1817_b0 );
not ( \1817_b0 , w_9837 );
and ( w_9837 , w_9836 , \1817_b1 );
or ( \1838_b1 , \1810_b1 , w_9840 );
or ( \1838_b0 , \1810_b0 , w_9839 );
not ( w_9839 , w_9841 );
and ( w_9841 , w_9840 , w_9838 );
or ( w_9838 , \1836_b1 , w_9842 );
or ( w_9839 , \1836_b0 , \1837_b0 );
not ( \1837_b0 , w_9843 );
and ( w_9843 , w_9842 , \1837_b1 );
or ( \1843_b1 , \1840_b1 , w_9846 );
or ( \1843_b0 , \1840_b0 , w_9845 );
not ( w_9845 , w_9847 );
and ( w_9847 , w_9846 , w_9844 );
or ( w_9844 , \1841_b1 , w_9848 );
or ( w_9845 , \1841_b0 , \1842_b0 );
not ( \1842_b0 , w_9849 );
and ( w_9849 , w_9848 , \1842_b1 );
or ( \1847_b1 , \1844_b1 , w_9852 );
or ( \1847_b0 , \1844_b0 , w_9851 );
not ( w_9851 , w_9853 );
and ( w_9853 , w_9852 , w_9850 );
or ( w_9850 , \1845_b1 , w_9854 );
or ( w_9851 , \1845_b0 , \1846_b0 );
not ( \1846_b0 , w_9855 );
and ( w_9855 , w_9854 , \1846_b1 );
or ( \1867_b1 , \1860_b1 , w_9858 );
or ( \1867_b0 , \1860_b0 , w_9857 );
not ( w_9857 , w_9859 );
and ( w_9859 , w_9858 , w_9856 );
or ( w_9856 , \1865_b1 , w_9860 );
or ( w_9857 , \1865_b0 , \1866_b0 );
not ( \1866_b0 , w_9861 );
and ( w_9861 , w_9860 , \1866_b1 );
or ( \1901_b1 , \1839_b1 , w_9864 );
or ( \1901_b0 , \1839_b0 , w_9863 );
not ( w_9863 , w_9865 );
and ( w_9865 , w_9864 , w_9862 );
or ( w_9862 , \1899_b1 , w_9866 );
or ( w_9863 , \1899_b0 , \1900_b0 );
not ( \1900_b0 , w_9867 );
and ( w_9867 , w_9866 , \1900_b1 );
or ( \1911_b1 , \1906_b1 , w_9870 );
or ( \1911_b0 , \1906_b0 , w_9869 );
not ( w_9869 , w_9871 );
and ( w_9871 , w_9870 , w_9868 );
or ( w_9868 , \1909_b1 , w_9872 );
or ( w_9869 , \1909_b0 , \1910_b0 );
not ( \1910_b0 , w_9873 );
and ( w_9873 , w_9872 , \1910_b1 );
or ( \1926_b1 , \1920_b1 , w_9876 );
or ( \1926_b0 , \1920_b0 , w_9875 );
not ( w_9875 , w_9877 );
and ( w_9877 , w_9876 , w_9874 );
or ( w_9874 , \1924_b1 , w_9878 );
or ( w_9875 , \1924_b0 , \1925_b0 );
not ( \1925_b0 , w_9879 );
and ( w_9879 , w_9878 , \1925_b1 );
or ( \1942_b1 , \1935_b1 , w_9882 );
or ( \1942_b0 , \1935_b0 , w_9881 );
not ( w_9881 , w_9883 );
and ( w_9883 , w_9882 , w_9880 );
or ( w_9880 , \1940_b1 , w_9884 );
or ( w_9881 , \1940_b0 , \1941_b0 );
not ( \1941_b0 , w_9885 );
and ( w_9885 , w_9884 , \1941_b1 );
or ( \1959_b1 , \1952_b1 , w_9888 );
or ( \1959_b0 , \1952_b0 , w_9887 );
not ( w_9887 , w_9889 );
and ( w_9889 , w_9888 , w_9886 );
or ( w_9886 , \1957_b1 , w_9890 );
or ( w_9887 , \1957_b0 , \1958_b0 );
not ( \1958_b0 , w_9891 );
and ( w_9891 , w_9890 , \1958_b1 );
or ( \1962_b1 , \1943_b1 , w_9894 );
or ( \1962_b0 , \1943_b0 , w_9893 );
not ( w_9893 , w_9895 );
and ( w_9895 , w_9894 , w_9892 );
or ( w_9892 , \1960_b1 , w_9896 );
or ( w_9893 , \1960_b0 , \1961_b0 );
not ( \1961_b0 , w_9897 );
and ( w_9897 , w_9896 , \1961_b1 );
or ( \1975_b1 , \1968_b1 , w_9900 );
or ( \1975_b0 , \1968_b0 , w_9899 );
not ( w_9899 , w_9901 );
and ( w_9901 , w_9900 , w_9898 );
or ( w_9898 , \1973_b1 , w_9902 );
or ( w_9899 , \1973_b0 , \1974_b0 );
not ( \1974_b0 , w_9903 );
and ( w_9903 , w_9902 , \1974_b1 );
or ( \1983_b1 , \1978_b1 , w_9906 );
or ( \1983_b0 , \1978_b0 , w_9905 );
not ( w_9905 , w_9907 );
and ( w_9907 , w_9906 , w_9904 );
or ( w_9904 , \1981_b1 , w_9908 );
or ( w_9905 , \1981_b0 , \1982_b0 );
not ( \1982_b0 , w_9909 );
and ( w_9909 , w_9908 , \1982_b1 );
or ( \1989_b1 , \1984_b1 , w_9912 );
or ( \1989_b0 , \1984_b0 , w_9911 );
not ( w_9911 , w_9913 );
and ( w_9913 , w_9912 , w_9910 );
or ( w_9910 , \1987_b1 , w_9914 );
or ( w_9911 , \1987_b0 , \1988_b0 );
not ( \1988_b0 , w_9915 );
and ( w_9915 , w_9914 , \1988_b1 );
or ( \1995_b1 , \1990_b1 , w_9918 );
or ( \1995_b0 , \1990_b0 , w_9917 );
not ( w_9917 , w_9919 );
and ( w_9919 , w_9918 , w_9916 );
or ( w_9916 , \1993_b1 , w_9920 );
or ( w_9917 , \1993_b0 , \1994_b0 );
not ( \1994_b0 , w_9921 );
and ( w_9921 , w_9920 , \1994_b1 );
or ( \1999_b1 , \1996_b1 , w_9924 );
or ( \1999_b0 , \1996_b0 , w_9923 );
not ( w_9923 , w_9925 );
and ( w_9925 , w_9924 , w_9922 );
or ( w_9922 , \1997_b1 , w_9926 );
or ( w_9923 , \1997_b0 , \1998_b0 );
not ( \1998_b0 , w_9927 );
and ( w_9927 , w_9926 , \1998_b1 );
or ( \2003_b1 , \2000_b1 , w_9930 );
or ( \2003_b0 , \2000_b0 , w_9929 );
not ( w_9929 , w_9931 );
and ( w_9931 , w_9930 , w_9928 );
or ( w_9928 , \2001_b1 , w_9932 );
or ( w_9929 , \2001_b0 , \2002_b0 );
not ( \2002_b0 , w_9933 );
and ( w_9933 , w_9932 , \2002_b1 );
or ( \2013_b1 , \2008_b1 , w_9936 );
or ( \2013_b0 , \2008_b0 , w_9935 );
not ( w_9935 , w_9937 );
and ( w_9937 , w_9936 , w_9934 );
or ( w_9934 , \2011_b1 , w_9938 );
or ( w_9935 , \2011_b0 , \2012_b0 );
not ( \2012_b0 , w_9939 );
and ( w_9939 , w_9938 , \2012_b1 );
or ( \2017_b1 , \2014_b1 , w_9942 );
or ( \2017_b0 , \2014_b0 , w_9941 );
not ( w_9941 , w_9943 );
and ( w_9943 , w_9942 , w_9940 );
or ( w_9940 , \2015_b1 , w_9944 );
or ( w_9941 , \2015_b0 , \2016_b0 );
not ( \2016_b0 , w_9945 );
and ( w_9945 , w_9944 , \2016_b1 );
or ( \2021_b1 , \2018_b1 , w_9948 );
or ( \2021_b0 , \2018_b0 , w_9947 );
not ( w_9947 , w_9949 );
and ( w_9949 , w_9948 , w_9946 );
or ( w_9946 , \2019_b1 , w_9950 );
or ( w_9947 , \2019_b0 , \2020_b0 );
not ( \2020_b0 , w_9951 );
and ( w_9951 , w_9950 , \2020_b1 );
or ( \2054_b1 , \2051_b1 , w_9954 );
or ( \2054_b0 , \2051_b0 , w_9953 );
not ( w_9953 , w_9955 );
and ( w_9955 , w_9954 , w_9952 );
or ( w_9952 , \2052_b1 , w_9956 );
or ( w_9953 , \2052_b0 , \2053_b0 );
not ( \2053_b0 , w_9957 );
and ( w_9957 , w_9956 , \2053_b1 );
or ( \2058_b1 , \2055_b1 , w_9960 );
or ( \2058_b0 , \2055_b0 , w_9959 );
not ( w_9959 , w_9961 );
and ( w_9961 , w_9960 , w_9958 );
or ( w_9958 , \2056_b1 , w_9962 );
or ( w_9959 , \2056_b0 , \2057_b0 );
not ( \2057_b0 , w_9963 );
and ( w_9963 , w_9962 , \2057_b1 );
or ( \2062_b1 , \2059_b1 , w_9966 );
or ( \2062_b0 , \2059_b0 , w_9965 );
not ( w_9965 , w_9967 );
and ( w_9967 , w_9966 , w_9964 );
or ( w_9964 , \2060_b1 , w_9968 );
or ( w_9965 , \2060_b0 , \2061_b0 );
not ( \2061_b0 , w_9969 );
and ( w_9969 , w_9968 , \2061_b1 );
or ( \2067_b1 , \2064_b1 , w_9972 );
or ( \2067_b0 , \2064_b0 , w_9971 );
not ( w_9971 , w_9973 );
and ( w_9973 , w_9972 , w_9970 );
or ( w_9970 , \2065_b1 , w_9974 );
or ( w_9971 , \2065_b0 , \2066_b0 );
not ( \2066_b0 , w_9975 );
and ( w_9975 , w_9974 , \2066_b1 );
or ( \2100_b1 , \2095_b1 , w_9978 );
or ( \2100_b0 , \2095_b0 , w_9977 );
not ( w_9977 , w_9979 );
and ( w_9979 , w_9978 , w_9976 );
or ( w_9976 , \2098_b1 , w_9980 );
or ( w_9977 , \2098_b0 , \2099_b0 );
not ( \2099_b0 , w_9981 );
and ( w_9981 , w_9980 , \2099_b1 );
or ( \2105_b1 , \2102_b1 , w_9984 );
or ( \2105_b0 , \2102_b0 , w_9983 );
not ( w_9983 , w_9985 );
and ( w_9985 , w_9984 , w_9982 );
or ( w_9982 , \2103_b1 , w_9986 );
or ( w_9983 , \2103_b0 , \2104_b0 );
not ( \2104_b0 , w_9987 );
and ( w_9987 , w_9986 , \2104_b1 );
or ( \2109_b1 , \2106_b1 , w_9990 );
or ( \2109_b0 , \2106_b0 , w_9989 );
not ( w_9989 , w_9991 );
and ( w_9991 , w_9990 , w_9988 );
or ( w_9988 , \2107_b1 , w_9992 );
or ( w_9989 , \2107_b0 , \2108_b0 );
not ( \2108_b0 , w_9993 );
and ( w_9993 , w_9992 , \2108_b1 );
or ( \2113_b1 , \2110_b1 , w_9996 );
or ( \2113_b0 , \2110_b0 , w_9995 );
not ( w_9995 , w_9997 );
and ( w_9997 , w_9996 , w_9994 );
or ( w_9994 , \2111_b1 , w_9998 );
or ( w_9995 , \2111_b0 , \2112_b0 );
not ( \2112_b0 , w_9999 );
and ( w_9999 , w_9998 , \2112_b1 );
or ( \2117_b1 , \2114_b1 , w_10002 );
or ( \2117_b0 , \2114_b0 , w_10001 );
not ( w_10001 , w_10003 );
and ( w_10003 , w_10002 , w_10000 );
or ( w_10000 , \2115_b1 , w_10004 );
or ( w_10001 , \2115_b0 , \2116_b0 );
not ( \2116_b0 , w_10005 );
and ( w_10005 , w_10004 , \2116_b1 );
or ( \2138_b1 , \2135_b1 , w_10008 );
or ( \2138_b0 , \2135_b0 , w_10007 );
not ( w_10007 , w_10009 );
and ( w_10009 , w_10008 , w_10006 );
or ( w_10006 , \2136_b1 , w_10010 );
or ( w_10007 , \2136_b0 , \2137_b0 );
not ( \2137_b0 , w_10011 );
and ( w_10011 , w_10010 , \2137_b1 );
or ( \2142_b1 , \2139_b1 , w_10014 );
or ( \2142_b0 , \2139_b0 , w_10013 );
not ( w_10013 , w_10015 );
and ( w_10015 , w_10014 , w_10012 );
or ( w_10012 , \2140_b1 , w_10016 );
or ( w_10013 , \2140_b0 , \2141_b0 );
not ( \2141_b0 , w_10017 );
and ( w_10017 , w_10016 , \2141_b1 );
or ( \2189_b1 , \2186_b1 , w_10020 );
or ( \2189_b0 , \2186_b0 , w_10019 );
not ( w_10019 , w_10021 );
and ( w_10021 , w_10020 , w_10018 );
or ( w_10018 , \2187_b1 , w_10022 );
or ( w_10019 , \2187_b0 , \2188_b0 );
not ( \2188_b0 , w_10023 );
and ( w_10023 , w_10022 , \2188_b1 );
or ( \2193_b1 , \2190_b1 , w_10026 );
or ( \2193_b0 , \2190_b0 , w_10025 );
not ( w_10025 , w_10027 );
and ( w_10027 , w_10026 , w_10024 );
or ( w_10024 , \2191_b1 , w_10028 );
or ( w_10025 , \2191_b0 , \2192_b0 );
not ( \2192_b0 , w_10029 );
and ( w_10029 , w_10028 , \2192_b1 );
or ( \2198_b1 , \2195_b1 , w_10032 );
or ( \2198_b0 , \2195_b0 , w_10031 );
not ( w_10031 , w_10033 );
and ( w_10033 , w_10032 , w_10030 );
or ( w_10030 , \2196_b1 , w_10034 );
or ( w_10031 , \2196_b0 , \2197_b0 );
not ( \2197_b0 , w_10035 );
and ( w_10035 , w_10034 , \2197_b1 );
or ( \2202_b1 , \2199_b1 , w_10038 );
or ( \2202_b0 , \2199_b0 , w_10037 );
not ( w_10037 , w_10039 );
and ( w_10039 , w_10038 , w_10036 );
or ( w_10036 , \2200_b1 , w_10040 );
or ( w_10037 , \2200_b0 , \2201_b0 );
not ( \2201_b0 , w_10041 );
and ( w_10041 , w_10040 , \2201_b1 );
or ( \2207_b1 , \2204_b1 , w_10044 );
or ( \2207_b0 , \2204_b0 , w_10043 );
not ( w_10043 , w_10045 );
and ( w_10045 , w_10044 , w_10042 );
or ( w_10042 , \2205_b1 , w_10046 );
or ( w_10043 , \2205_b0 , \2206_b0 );
not ( \2206_b0 , w_10047 );
and ( w_10047 , w_10046 , \2206_b1 );
or ( \2211_b1 , \2208_b1 , w_10050 );
or ( \2211_b0 , \2208_b0 , w_10049 );
not ( w_10049 , w_10051 );
and ( w_10051 , w_10050 , w_10048 );
or ( w_10048 , \2209_b1 , w_10052 );
or ( w_10049 , \2209_b0 , \2210_b0 );
not ( \2210_b0 , w_10053 );
and ( w_10053 , w_10052 , \2210_b1 );
or ( \2264_b1 , \2259_b1 , w_10056 );
or ( \2264_b0 , \2259_b0 , w_10055 );
not ( w_10055 , w_10057 );
and ( w_10057 , w_10056 , w_10054 );
or ( w_10054 , \2262_b1 , w_10058 );
or ( w_10055 , \2262_b0 , \2263_b0 );
not ( \2263_b0 , w_10059 );
and ( w_10059 , w_10058 , \2263_b1 );
or ( \2272_b1 , \2267_b1 , w_10062 );
or ( \2272_b0 , \2267_b0 , w_10061 );
not ( w_10061 , w_10063 );
and ( w_10063 , w_10062 , w_10060 );
or ( w_10060 , \2270_b1 , w_10064 );
or ( w_10061 , \2270_b0 , \2271_b0 );
not ( \2271_b0 , w_10065 );
and ( w_10065 , w_10064 , \2271_b1 );
or ( \2280_b1 , \2275_b1 , w_10068 );
or ( \2280_b0 , \2275_b0 , w_10067 );
not ( w_10067 , w_10069 );
and ( w_10069 , w_10068 , w_10066 );
or ( w_10066 , \2278_b1 , w_10070 );
or ( w_10067 , \2278_b0 , \2279_b0 );
not ( \2279_b0 , w_10071 );
and ( w_10071 , w_10070 , \2279_b1 );
or ( \2288_b1 , \2283_b1 , w_10074 );
or ( \2288_b0 , \2283_b0 , w_10073 );
not ( w_10073 , w_10075 );
and ( w_10075 , w_10074 , w_10072 );
or ( w_10072 , \2286_b1 , w_10076 );
or ( w_10073 , \2286_b0 , \2287_b0 );
not ( \2287_b0 , w_10077 );
and ( w_10077 , w_10076 , \2287_b1 );
or ( \2302_b1 , \2299_b1 , w_10080 );
or ( \2302_b0 , \2299_b0 , w_10079 );
not ( w_10079 , w_10081 );
and ( w_10081 , w_10080 , w_10078 );
or ( w_10078 , \2300_b1 , w_10082 );
or ( w_10079 , \2300_b0 , \2301_b0 );
not ( \2301_b0 , w_10083 );
and ( w_10083 , w_10082 , \2301_b1 );
or ( \2318_b1 , \2311_b1 , w_10086 );
or ( \2318_b0 , \2311_b0 , w_10085 );
not ( w_10085 , w_10087 );
and ( w_10087 , w_10086 , w_10084 );
or ( w_10084 , \2316_b1 , w_10088 );
or ( w_10085 , \2316_b0 , \2317_b0 );
not ( \2317_b0 , w_10089 );
and ( w_10089 , w_10088 , \2317_b1 );
or ( \2326_b1 , \2319_b1 , w_10092 );
or ( \2326_b0 , \2319_b0 , w_10091 );
not ( w_10091 , w_10093 );
and ( w_10093 , w_10092 , w_10090 );
or ( w_10090 , \2324_b1 , w_10094 );
or ( w_10091 , \2324_b0 , \2325_b0 );
not ( \2325_b0 , w_10095 );
and ( w_10095 , w_10094 , \2325_b1 );
or ( \2342_b1 , \2335_b1 , w_10098 );
or ( \2342_b0 , \2335_b0 , w_10097 );
not ( w_10097 , w_10099 );
and ( w_10099 , w_10098 , w_10096 );
or ( w_10096 , \2340_b1 , w_10100 );
or ( w_10097 , \2340_b0 , \2341_b0 );
not ( \2341_b0 , w_10101 );
and ( w_10101 , w_10100 , \2341_b1 );
or ( \2358_b1 , \2351_b1 , w_10104 );
or ( \2358_b0 , \2351_b0 , w_10103 );
not ( w_10103 , w_10105 );
and ( w_10105 , w_10104 , w_10102 );
or ( w_10102 , \2356_b1 , w_10106 );
or ( w_10103 , \2356_b0 , \2357_b0 );
not ( \2357_b0 , w_10107 );
and ( w_10107 , w_10106 , \2357_b1 );
or ( \2364_b1 , \2359_b1 , w_10110 );
or ( \2364_b0 , \2359_b0 , w_10109 );
not ( w_10109 , w_10111 );
and ( w_10111 , w_10110 , w_10108 );
or ( w_10108 , \2362_b1 , w_10112 );
or ( w_10109 , \2362_b0 , \2363_b0 );
not ( \2363_b0 , w_10113 );
and ( w_10113 , w_10112 , \2363_b1 );
or ( \2370_b1 , \2365_b1 , w_10116 );
or ( \2370_b0 , \2365_b0 , w_10115 );
not ( w_10115 , w_10117 );
and ( w_10117 , w_10116 , w_10114 );
or ( w_10114 , \2368_b1 , w_10118 );
or ( w_10115 , \2368_b0 , \2369_b0 );
not ( \2369_b0 , w_10119 );
and ( w_10119 , w_10118 , \2369_b1 );
or ( \2380_b1 , \2375_b1 , w_10122 );
or ( \2380_b0 , \2375_b0 , w_10121 );
not ( w_10121 , w_10123 );
and ( w_10123 , w_10122 , w_10120 );
or ( w_10120 , \2378_b1 , w_10124 );
or ( w_10121 , \2378_b0 , \2379_b0 );
not ( \2379_b0 , w_10125 );
and ( w_10125 , w_10124 , \2379_b1 );
or ( \2388_b1 , \2383_b1 , w_10128 );
or ( \2388_b0 , \2383_b0 , w_10127 );
not ( w_10127 , w_10129 );
and ( w_10129 , w_10128 , w_10126 );
or ( w_10126 , \2386_b1 , w_10130 );
or ( w_10127 , \2386_b0 , \2387_b0 );
not ( \2387_b0 , w_10131 );
and ( w_10131 , w_10130 , \2387_b1 );
or ( \2394_b1 , \2389_b1 , w_10134 );
or ( \2394_b0 , \2389_b0 , w_10133 );
not ( w_10133 , w_10135 );
and ( w_10135 , w_10134 , w_10132 );
or ( w_10132 , \2392_b1 , w_10136 );
or ( w_10133 , \2392_b0 , \2393_b0 );
not ( \2393_b0 , w_10137 );
and ( w_10137 , w_10136 , \2393_b1 );
or ( \2402_b1 , \2397_b1 , w_10140 );
or ( \2402_b0 , \2397_b0 , w_10139 );
not ( w_10139 , w_10141 );
and ( w_10141 , w_10140 , w_10138 );
or ( w_10138 , \2400_b1 , w_10142 );
or ( w_10139 , \2400_b0 , \2401_b0 );
not ( \2401_b0 , w_10143 );
and ( w_10143 , w_10142 , \2401_b1 );
or ( \2424_b1 , \2417_b1 , w_10146 );
or ( \2424_b0 , \2417_b0 , w_10145 );
not ( w_10145 , w_10147 );
and ( w_10147 , w_10146 , w_10144 );
or ( w_10144 , \2422_b1 , w_10148 );
or ( w_10145 , \2422_b0 , \2423_b0 );
not ( \2423_b0 , w_10149 );
and ( w_10149 , w_10148 , \2423_b1 );
or ( \2441_b1 , \2434_b1 , w_10152 );
or ( \2441_b0 , \2434_b0 , w_10151 );
not ( w_10151 , w_10153 );
and ( w_10153 , w_10152 , w_10150 );
or ( w_10150 , \2439_b1 , w_10154 );
or ( w_10151 , \2439_b0 , \2440_b0 );
not ( \2440_b0 , w_10155 );
and ( w_10155 , w_10154 , \2440_b1 );
or ( \2457_b1 , \2450_b1 , w_10158 );
or ( \2457_b0 , \2450_b0 , w_10157 );
not ( w_10157 , w_10159 );
and ( w_10159 , w_10158 , w_10156 );
or ( w_10156 , \2455_b1 , w_10160 );
or ( w_10157 , \2455_b0 , \2456_b0 );
not ( \2456_b0 , w_10161 );
and ( w_10161 , w_10160 , \2456_b1 );
or ( \2472_b1 , \2466_b1 , w_10164 );
or ( \2472_b0 , \2466_b0 , w_10163 );
not ( w_10163 , w_10165 );
and ( w_10165 , w_10164 , w_10162 );
or ( w_10162 , \2470_b1 , w_10166 );
or ( w_10163 , \2470_b0 , \2471_b0 );
not ( \2471_b0 , w_10167 );
and ( w_10167 , w_10166 , \2471_b1 );
or ( \2478_b1 , \2473_b1 , w_10170 );
or ( \2478_b0 , \2473_b0 , w_10169 );
not ( w_10169 , w_10171 );
and ( w_10171 , w_10170 , w_10168 );
or ( w_10168 , \2476_b1 , w_10172 );
or ( w_10169 , \2476_b0 , \2477_b0 );
not ( \2477_b0 , w_10173 );
and ( w_10173 , w_10172 , \2477_b1 );
or ( \2484_b1 , \2479_b1 , w_10176 );
or ( \2484_b0 , \2479_b0 , w_10175 );
not ( w_10175 , w_10177 );
and ( w_10177 , w_10176 , w_10174 );
or ( w_10174 , \2482_b1 , w_10178 );
or ( w_10175 , \2482_b0 , \2483_b0 );
not ( \2483_b0 , w_10179 );
and ( w_10179 , w_10178 , \2483_b1 );
or ( \2494_b1 , \2489_b1 , w_10182 );
or ( \2494_b0 , \2489_b0 , w_10181 );
not ( w_10181 , w_10183 );
and ( w_10183 , w_10182 , w_10180 );
or ( w_10180 , \2492_b1 , w_10184 );
or ( w_10181 , \2492_b0 , \2493_b0 );
not ( \2493_b0 , w_10185 );
and ( w_10185 , w_10184 , \2493_b1 );
or ( \2502_b1 , \2497_b1 , w_10188 );
or ( \2502_b0 , \2497_b0 , w_10187 );
not ( w_10187 , w_10189 );
and ( w_10189 , w_10188 , w_10186 );
or ( w_10186 , \2500_b1 , w_10190 );
or ( w_10187 , \2500_b0 , \2501_b0 );
not ( \2501_b0 , w_10191 );
and ( w_10191 , w_10190 , \2501_b1 );
or ( \2508_b1 , \2503_b1 , w_10194 );
or ( \2508_b0 , \2503_b0 , w_10193 );
not ( w_10193 , w_10195 );
and ( w_10195 , w_10194 , w_10192 );
or ( w_10192 , \2506_b1 , w_10196 );
or ( w_10193 , \2506_b0 , \2507_b0 );
not ( \2507_b0 , w_10197 );
and ( w_10197 , w_10196 , \2507_b1 );
or ( \2516_b1 , \2511_b1 , w_10200 );
or ( \2516_b0 , \2511_b0 , w_10199 );
not ( w_10199 , w_10201 );
and ( w_10201 , w_10200 , w_10198 );
or ( w_10198 , \2514_b1 , w_10202 );
or ( w_10199 , \2514_b0 , \2515_b0 );
not ( \2515_b0 , w_10203 );
and ( w_10203 , w_10202 , \2515_b1 );
or ( \2532_b1 , \2529_b1 , w_10206 );
or ( \2532_b0 , \2529_b0 , w_10205 );
not ( w_10205 , w_10207 );
and ( w_10207 , w_10206 , w_10204 );
or ( w_10204 , \2530_b1 , w_10208 );
or ( w_10205 , \2530_b0 , \2531_b0 );
not ( \2531_b0 , w_10209 );
and ( w_10209 , w_10208 , \2531_b1 );
or ( \2548_b1 , \2541_b1 , w_10212 );
or ( \2548_b0 , \2541_b0 , w_10211 );
not ( w_10211 , w_10213 );
and ( w_10213 , w_10212 , w_10210 );
or ( w_10210 , \2546_b1 , w_10214 );
or ( w_10211 , \2546_b0 , \2547_b0 );
not ( \2547_b0 , w_10215 );
and ( w_10215 , w_10214 , \2547_b1 );
or ( \2565_b1 , \2558_b1 , w_10218 );
or ( \2565_b0 , \2558_b0 , w_10217 );
not ( w_10217 , w_10219 );
and ( w_10219 , w_10218 , w_10216 );
or ( w_10216 , \2563_b1 , w_10220 );
or ( w_10217 , \2563_b0 , \2564_b0 );
not ( \2564_b0 , w_10221 );
and ( w_10221 , w_10220 , \2564_b1 );
or ( \2568_b1 , \2549_b1 , w_10224 );
or ( \2568_b0 , \2549_b0 , w_10223 );
not ( w_10223 , w_10225 );
and ( w_10225 , w_10224 , w_10222 );
or ( w_10222 , \2566_b1 , w_10226 );
or ( w_10223 , \2566_b0 , \2567_b0 );
not ( \2567_b0 , w_10227 );
and ( w_10227 , w_10226 , \2567_b1 );
or ( \2581_b1 , \2574_b1 , w_10230 );
or ( \2581_b0 , \2574_b0 , w_10229 );
not ( w_10229 , w_10231 );
and ( w_10231 , w_10230 , w_10228 );
or ( w_10228 , \2579_b1 , w_10232 );
or ( w_10229 , \2579_b0 , \2580_b0 );
not ( \2580_b0 , w_10233 );
and ( w_10233 , w_10232 , \2580_b1 );
or ( \2587_b1 , \2582_b1 , w_10236 );
or ( \2587_b0 , \2582_b0 , w_10235 );
not ( w_10235 , w_10237 );
and ( w_10237 , w_10236 , w_10234 );
or ( w_10234 , \2585_b1 , w_10238 );
or ( w_10235 , \2585_b0 , \2586_b0 );
not ( \2586_b0 , w_10239 );
and ( w_10239 , w_10238 , \2586_b1 );
or ( \2603_b1 , \2596_b1 , w_10242 );
or ( \2603_b0 , \2596_b0 , w_10241 );
not ( w_10241 , w_10243 );
and ( w_10243 , w_10242 , w_10240 );
or ( w_10240 , \2601_b1 , w_10244 );
or ( w_10241 , \2601_b0 , \2602_b0 );
not ( \2602_b0 , w_10245 );
and ( w_10245 , w_10244 , \2602_b1 );
or ( \2611_b1 , \2606_b1 , w_10248 );
or ( \2611_b0 , \2606_b0 , w_10247 );
not ( w_10247 , w_10249 );
and ( w_10249 , w_10248 , w_10246 );
or ( w_10246 , \2609_b1 , w_10250 );
or ( w_10247 , \2609_b0 , \2610_b0 );
not ( \2610_b0 , w_10251 );
and ( w_10251 , w_10250 , \2610_b1 );
or ( \2619_b1 , \2614_b1 , w_10254 );
or ( \2619_b0 , \2614_b0 , w_10253 );
not ( w_10253 , w_10255 );
and ( w_10255 , w_10254 , w_10252 );
or ( w_10252 , \2617_b1 , w_10256 );
or ( w_10253 , \2617_b0 , \2618_b0 );
not ( \2618_b0 , w_10257 );
and ( w_10257 , w_10256 , \2618_b1 );
or ( \2625_b1 , \2620_b1 , w_10260 );
or ( \2625_b0 , \2620_b0 , w_10259 );
not ( w_10259 , w_10261 );
and ( w_10261 , w_10260 , w_10258 );
or ( w_10258 , \2623_b1 , w_10262 );
or ( w_10259 , \2623_b0 , \2624_b0 );
not ( \2624_b0 , w_10263 );
and ( w_10263 , w_10262 , \2624_b1 );
or ( \2633_b1 , \2628_b1 , w_10266 );
or ( \2633_b0 , \2628_b0 , w_10265 );
not ( w_10265 , w_10267 );
and ( w_10267 , w_10266 , w_10264 );
or ( w_10264 , \2631_b1 , w_10268 );
or ( w_10265 , \2631_b0 , \2632_b0 );
not ( \2632_b0 , w_10269 );
and ( w_10269 , w_10268 , \2632_b1 );
or ( \2653_b1 , \2646_b1 , w_10272 );
or ( \2653_b0 , \2646_b0 , w_10271 );
not ( w_10271 , w_10273 );
and ( w_10273 , w_10272 , w_10270 );
or ( w_10270 , \2651_b1 , w_10274 );
or ( w_10271 , \2651_b0 , \2652_b0 );
not ( \2652_b0 , w_10275 );
and ( w_10275 , w_10274 , \2652_b1 );
or ( \2669_b1 , \2662_b1 , w_10278 );
or ( \2669_b0 , \2662_b0 , w_10277 );
not ( w_10277 , w_10279 );
and ( w_10279 , w_10278 , w_10276 );
or ( w_10276 , \2667_b1 , w_10280 );
or ( w_10277 , \2667_b0 , \2668_b0 );
not ( \2668_b0 , w_10281 );
and ( w_10281 , w_10280 , \2668_b1 );
or ( \2681_b1 , \2670_b1 , w_10284 );
or ( \2681_b0 , \2670_b0 , w_10283 );
not ( w_10283 , w_10285 );
and ( w_10285 , w_10284 , w_10282 );
or ( w_10282 , \2679_b1 , w_10286 );
or ( w_10283 , \2679_b0 , \2680_b0 );
not ( \2680_b0 , w_10287 );
and ( w_10287 , w_10286 , \2680_b1 );
or ( \2689_b1 , \2684_b1 , w_10290 );
or ( \2689_b0 , \2684_b0 , w_10289 );
not ( w_10289 , w_10291 );
and ( w_10291 , w_10290 , w_10288 );
or ( w_10288 , \2687_b1 , w_10292 );
or ( w_10289 , \2687_b0 , \2688_b0 );
not ( \2688_b0 , w_10293 );
and ( w_10293 , w_10292 , \2688_b1 );
or ( \2705_b1 , \2698_b1 , w_10296 );
or ( \2705_b0 , \2698_b0 , w_10295 );
not ( w_10295 , w_10297 );
and ( w_10297 , w_10296 , w_10294 );
or ( w_10294 , \2703_b1 , w_10298 );
or ( w_10295 , \2703_b0 , \2704_b0 );
not ( \2704_b0 , w_10299 );
and ( w_10299 , w_10298 , \2704_b1 );
or ( \2713_b1 , \2708_b1 , w_10302 );
or ( \2713_b0 , \2708_b0 , w_10301 );
not ( w_10301 , w_10303 );
and ( w_10303 , w_10302 , w_10300 );
or ( w_10300 , \2711_b1 , w_10304 );
or ( w_10301 , \2711_b0 , \2712_b0 );
not ( \2712_b0 , w_10305 );
and ( w_10305 , w_10304 , \2712_b1 );
or ( \2726_b1 , \2723_b1 , w_10308 );
or ( \2726_b0 , \2723_b0 , w_10307 );
not ( w_10307 , w_10309 );
and ( w_10309 , w_10308 , w_10306 );
or ( w_10306 , \2724_b1 , w_10310 );
or ( w_10307 , \2724_b0 , \2725_b0 );
not ( \2725_b0 , w_10311 );
and ( w_10311 , w_10310 , \2725_b1 );
or ( \2734_b1 , \2727_b1 , w_10314 );
or ( \2734_b0 , \2727_b0 , w_10313 );
not ( w_10313 , w_10315 );
and ( w_10315 , w_10314 , w_10312 );
or ( w_10312 , \2732_b1 , w_10316 );
or ( w_10313 , \2732_b0 , \2733_b0 );
not ( \2733_b0 , w_10317 );
and ( w_10317 , w_10316 , \2733_b1 );
or ( \2742_b1 , \2737_b1 , w_10320 );
or ( \2742_b0 , \2737_b0 , w_10319 );
not ( w_10319 , w_10321 );
and ( w_10321 , w_10320 , w_10318 );
or ( w_10318 , \2740_b1 , w_10322 );
or ( w_10319 , \2740_b0 , \2741_b0 );
not ( \2741_b0 , w_10323 );
and ( w_10323 , w_10322 , \2741_b1 );
or ( \2748_b1 , \2743_b1 , w_10326 );
or ( \2748_b0 , \2743_b0 , w_10325 );
not ( w_10325 , w_10327 );
and ( w_10327 , w_10326 , w_10324 );
or ( w_10324 , \2746_b1 , w_10328 );
or ( w_10325 , \2746_b0 , \2747_b0 );
not ( \2747_b0 , w_10329 );
and ( w_10329 , w_10328 , \2747_b1 );
or ( \2754_b1 , \2749_b1 , w_10332 );
or ( \2754_b0 , \2749_b0 , w_10331 );
not ( w_10331 , w_10333 );
and ( w_10333 , w_10332 , w_10330 );
or ( w_10330 , \2752_b1 , w_10334 );
or ( w_10331 , \2752_b0 , \2753_b0 );
not ( \2753_b0 , w_10335 );
and ( w_10335 , w_10334 , \2753_b1 );
or ( \2762_b1 , \2757_b1 , w_10338 );
or ( \2762_b0 , \2757_b0 , w_10337 );
not ( w_10337 , w_10339 );
and ( w_10339 , w_10338 , w_10336 );
or ( w_10336 , \2760_b1 , w_10340 );
or ( w_10337 , \2760_b0 , \2761_b0 );
not ( \2761_b0 , w_10341 );
and ( w_10341 , w_10340 , \2761_b1 );
or ( \2782_b1 , \2775_b1 , w_10344 );
or ( \2782_b0 , \2775_b0 , w_10343 );
not ( w_10343 , w_10345 );
and ( w_10345 , w_10344 , w_10342 );
or ( w_10342 , \2780_b1 , w_10346 );
or ( w_10343 , \2780_b0 , \2781_b0 );
not ( \2781_b0 , w_10347 );
and ( w_10347 , w_10346 , \2781_b1 );
or ( \2798_b1 , \2791_b1 , w_10350 );
or ( \2798_b0 , \2791_b0 , w_10349 );
not ( w_10349 , w_10351 );
and ( w_10351 , w_10350 , w_10348 );
or ( w_10348 , \2796_b1 , w_10352 );
or ( w_10349 , \2796_b0 , \2797_b0 );
not ( \2797_b0 , w_10353 );
and ( w_10353 , w_10352 , \2797_b1 );
or ( \2804_b1 , \2799_b1 , w_10356 );
or ( \2804_b0 , \2799_b0 , w_10355 );
not ( w_10355 , w_10357 );
and ( w_10357 , w_10356 , w_10354 );
or ( w_10354 , \2802_b1 , w_10358 );
or ( w_10355 , \2802_b0 , \2803_b0 );
not ( \2803_b0 , w_10359 );
and ( w_10359 , w_10358 , \2803_b1 );
or ( \2824_b1 , \2817_b1 , w_10362 );
or ( \2824_b0 , \2817_b0 , w_10361 );
not ( w_10361 , w_10363 );
and ( w_10363 , w_10362 , w_10360 );
or ( w_10360 , \2822_b1 , w_10364 );
or ( w_10361 , \2822_b0 , \2823_b0 );
not ( \2823_b0 , w_10365 );
and ( w_10365 , w_10364 , \2823_b1 );
or ( \2832_b1 , \2827_b1 , w_10368 );
or ( \2832_b0 , \2827_b0 , w_10367 );
not ( w_10367 , w_10369 );
and ( w_10369 , w_10368 , w_10366 );
or ( w_10366 , \2830_b1 , w_10370 );
or ( w_10367 , \2830_b0 , \2831_b0 );
not ( \2831_b0 , w_10371 );
and ( w_10371 , w_10370 , \2831_b1 );
or ( \2838_b1 , \2833_b1 , w_10374 );
or ( \2838_b0 , \2833_b0 , w_10373 );
not ( w_10373 , w_10375 );
and ( w_10375 , w_10374 , w_10372 );
or ( w_10372 , \2836_b1 , w_10376 );
or ( w_10373 , \2836_b0 , \2837_b0 );
not ( \2837_b0 , w_10377 );
and ( w_10377 , w_10376 , \2837_b1 );
or ( \2846_b1 , \2841_b1 , w_10380 );
or ( \2846_b0 , \2841_b0 , w_10379 );
not ( w_10379 , w_10381 );
and ( w_10381 , w_10380 , w_10378 );
or ( w_10378 , \2844_b1 , w_10382 );
or ( w_10379 , \2844_b0 , \2845_b0 );
not ( \2845_b0 , w_10383 );
and ( w_10383 , w_10382 , \2845_b1 );
or ( \2854_b1 , \2849_b1 , w_10386 );
or ( \2854_b0 , \2849_b0 , w_10385 );
not ( w_10385 , w_10387 );
and ( w_10387 , w_10386 , w_10384 );
or ( w_10384 , \2852_b1 , w_10388 );
or ( w_10385 , \2852_b0 , \2853_b0 );
not ( \2853_b0 , w_10389 );
and ( w_10389 , w_10388 , \2853_b1 );
or ( \2874_b1 , \2867_b1 , w_10392 );
or ( \2874_b0 , \2867_b0 , w_10391 );
not ( w_10391 , w_10393 );
and ( w_10393 , w_10392 , w_10390 );
or ( w_10390 , \2872_b1 , w_10394 );
or ( w_10391 , \2872_b0 , \2873_b0 );
not ( \2873_b0 , w_10395 );
and ( w_10395 , w_10394 , \2873_b1 );
or ( \2890_b1 , \2883_b1 , w_10398 );
or ( \2890_b0 , \2883_b0 , w_10397 );
not ( w_10397 , w_10399 );
and ( w_10399 , w_10398 , w_10396 );
or ( w_10396 , \2888_b1 , w_10400 );
or ( w_10397 , \2888_b0 , \2889_b0 );
not ( \2889_b0 , w_10401 );
and ( w_10401 , w_10400 , \2889_b1 );
or ( \2896_b1 , \2891_b1 , w_10404 );
or ( \2896_b0 , \2891_b0 , w_10403 );
not ( w_10403 , w_10405 );
and ( w_10405 , w_10404 , w_10402 );
or ( w_10402 , \2894_b1 , w_10406 );
or ( w_10403 , \2894_b0 , \2895_b0 );
not ( \2895_b0 , w_10407 );
and ( w_10407 , w_10406 , \2895_b1 );
or ( \2904_b1 , \2899_b1 , w_10410 );
or ( \2904_b0 , \2899_b0 , w_10409 );
not ( w_10409 , w_10411 );
and ( w_10411 , w_10410 , w_10408 );
or ( w_10408 , \2902_b1 , w_10412 );
or ( w_10409 , \2902_b0 , \2903_b0 );
not ( \2903_b0 , w_10413 );
and ( w_10413 , w_10412 , \2903_b1 );
or ( \2912_b1 , \2907_b1 , w_10416 );
or ( \2912_b0 , \2907_b0 , w_10415 );
not ( w_10415 , w_10417 );
and ( w_10417 , w_10416 , w_10414 );
or ( w_10414 , \2910_b1 , w_10418 );
or ( w_10415 , \2910_b0 , \2911_b0 );
not ( \2911_b0 , w_10419 );
and ( w_10419 , w_10418 , \2911_b1 );
or ( \2920_b1 , \2915_b1 , w_10422 );
or ( \2920_b0 , \2915_b0 , w_10421 );
not ( w_10421 , w_10423 );
and ( w_10423 , w_10422 , w_10420 );
or ( w_10420 , \2918_b1 , w_10424 );
or ( w_10421 , \2918_b0 , \2919_b0 );
not ( \2919_b0 , w_10425 );
and ( w_10425 , w_10424 , \2919_b1 );
or ( \2935_b1 , \2928_b1 , w_10428 );
or ( \2935_b0 , \2928_b0 , w_10427 );
not ( w_10427 , w_10429 );
and ( w_10429 , w_10428 , w_10426 );
or ( w_10426 , \2933_b1 , w_10430 );
or ( w_10427 , \2933_b0 , \2934_b0 );
not ( \2934_b0 , w_10431 );
and ( w_10431 , w_10430 , \2934_b1 );
or ( \2943_b1 , \2938_b1 , w_10434 );
or ( \2943_b0 , \2938_b0 , w_10433 );
not ( w_10433 , w_10435 );
and ( w_10435 , w_10434 , w_10432 );
or ( w_10432 , \2941_b1 , w_10436 );
or ( w_10433 , \2941_b0 , \2942_b0 );
not ( \2942_b0 , w_10437 );
and ( w_10437 , w_10436 , \2942_b1 );
or ( \2955_b1 , \2952_b1 , w_10440 );
or ( \2955_b0 , \2952_b0 , w_10439 );
not ( w_10439 , w_10441 );
and ( w_10441 , w_10440 , w_10438 );
or ( w_10438 , \2953_b1 , w_10442 );
or ( w_10439 , \2953_b0 , \2954_b0 );
not ( \2954_b0 , w_10443 );
and ( w_10443 , w_10442 , \2954_b1 );
or ( \2971_b1 , \2964_b1 , w_10446 );
or ( \2971_b0 , \2964_b0 , w_10445 );
not ( w_10445 , w_10447 );
and ( w_10447 , w_10446 , w_10444 );
or ( w_10444 , \2969_b1 , w_10448 );
or ( w_10445 , \2969_b0 , \2970_b0 );
not ( \2970_b0 , w_10449 );
and ( w_10449 , w_10448 , \2970_b1 );
or ( \2979_b1 , \2972_b1 , w_10452 );
or ( \2979_b0 , \2972_b0 , w_10451 );
not ( w_10451 , w_10453 );
and ( w_10453 , w_10452 , w_10450 );
or ( w_10450 , \2977_b1 , w_10454 );
or ( w_10451 , \2977_b0 , \2978_b0 );
not ( \2978_b0 , w_10455 );
and ( w_10455 , w_10454 , \2978_b1 );
or ( \2987_b1 , \2982_b1 , w_10458 );
or ( \2987_b0 , \2982_b0 , w_10457 );
not ( w_10457 , w_10459 );
and ( w_10459 , w_10458 , w_10456 );
or ( w_10456 , \2985_b1 , w_10460 );
or ( w_10457 , \2985_b0 , \2986_b0 );
not ( \2986_b0 , w_10461 );
and ( w_10461 , w_10460 , \2986_b1 );
or ( \2993_b1 , \2988_b1 , w_10464 );
or ( \2993_b0 , \2988_b0 , w_10463 );
not ( w_10463 , w_10465 );
and ( w_10465 , w_10464 , w_10462 );
or ( w_10462 , \2991_b1 , w_10466 );
or ( w_10463 , \2991_b0 , \2992_b0 );
not ( \2992_b0 , w_10467 );
and ( w_10467 , w_10466 , \2992_b1 );
or ( \3001_b1 , \2996_b1 , w_10470 );
or ( \3001_b0 , \2996_b0 , w_10469 );
not ( w_10469 , w_10471 );
and ( w_10471 , w_10470 , w_10468 );
or ( w_10468 , \2999_b1 , w_10472 );
or ( w_10469 , \2999_b0 , \3000_b0 );
not ( \3000_b0 , w_10473 );
and ( w_10473 , w_10472 , \3000_b1 );
or ( \3023_b1 , \3016_b1 , w_10476 );
or ( \3023_b0 , \3016_b0 , w_10475 );
not ( w_10475 , w_10477 );
and ( w_10477 , w_10476 , w_10474 );
or ( w_10474 , \3021_b1 , w_10478 );
or ( w_10475 , \3021_b0 , \3022_b0 );
not ( \3022_b0 , w_10479 );
and ( w_10479 , w_10478 , \3022_b1 );
or ( \3031_b1 , \3026_b1 , w_10482 );
or ( \3031_b0 , \3026_b0 , w_10481 );
not ( w_10481 , w_10483 );
and ( w_10483 , w_10482 , w_10480 );
or ( w_10480 , \3029_b1 , w_10484 );
or ( w_10481 , \3029_b0 , \3030_b0 );
not ( \3030_b0 , w_10485 );
and ( w_10485 , w_10484 , \3030_b1 );
or ( \3049_b1 , \3044_b1 , w_10488 );
or ( \3049_b0 , \3044_b0 , w_10487 );
not ( w_10487 , w_10489 );
and ( w_10489 , w_10488 , w_10486 );
or ( w_10486 , \3047_b1 , w_10490 );
or ( w_10487 , \3047_b0 , \3048_b0 );
not ( \3048_b0 , w_10491 );
and ( w_10491 , w_10490 , \3048_b1 );
or ( \3057_b1 , \3052_b1 , w_10494 );
or ( \3057_b0 , \3052_b0 , w_10493 );
not ( w_10493 , w_10495 );
and ( w_10495 , w_10494 , w_10492 );
or ( w_10492 , \3055_b1 , w_10496 );
or ( w_10493 , \3055_b0 , \3056_b0 );
not ( \3056_b0 , w_10497 );
and ( w_10497 , w_10496 , \3056_b1 );
or ( \3063_b1 , \3058_b1 , w_10500 );
or ( \3063_b0 , \3058_b0 , w_10499 );
not ( w_10499 , w_10501 );
and ( w_10501 , w_10500 , w_10498 );
or ( w_10498 , \3061_b1 , w_10502 );
or ( w_10499 , \3061_b0 , \3062_b0 );
not ( \3062_b0 , w_10503 );
and ( w_10503 , w_10502 , \3062_b1 );
or ( \3071_b1 , \3066_b1 , w_10506 );
or ( \3071_b0 , \3066_b0 , w_10505 );
not ( w_10505 , w_10507 );
and ( w_10507 , w_10506 , w_10504 );
or ( w_10504 , \3069_b1 , w_10508 );
or ( w_10505 , \3069_b0 , \3070_b0 );
not ( \3070_b0 , w_10509 );
and ( w_10509 , w_10508 , \3070_b1 );
or ( \3091_b1 , \3084_b1 , w_10512 );
or ( \3091_b0 , \3084_b0 , w_10511 );
not ( w_10511 , w_10513 );
and ( w_10513 , w_10512 , w_10510 );
or ( w_10510 , \3089_b1 , w_10514 );
or ( w_10511 , \3089_b0 , \3090_b0 );
not ( \3090_b0 , w_10515 );
and ( w_10515 , w_10514 , \3090_b1 );
or ( \3107_b1 , \3100_b1 , w_10518 );
or ( \3107_b0 , \3100_b0 , w_10517 );
not ( w_10517 , w_10519 );
and ( w_10519 , w_10518 , w_10516 );
or ( w_10516 , \3105_b1 , w_10520 );
or ( w_10517 , \3105_b0 , \3106_b0 );
not ( \3106_b0 , w_10521 );
and ( w_10521 , w_10520 , \3106_b1 );
or ( \3121_b1 , \3114_b1 , w_10524 );
or ( \3121_b0 , \3114_b0 , w_10523 );
not ( w_10523 , w_10525 );
and ( w_10525 , w_10524 , w_10522 );
or ( w_10522 , \3119_b1 , w_10526 );
or ( w_10523 , \3119_b0 , \3120_b0 );
not ( \3120_b0 , w_10527 );
and ( w_10527 , w_10526 , \3120_b1 );
or ( \3124_b1 , \3108_b1 , w_10530 );
or ( \3124_b0 , \3108_b0 , w_10529 );
not ( w_10529 , w_10531 );
and ( w_10531 , w_10530 , w_10528 );
or ( w_10528 , \3122_b1 , w_10532 );
or ( w_10529 , \3122_b0 , \3123_b0 );
not ( \3123_b0 , w_10533 );
and ( w_10533 , w_10532 , \3123_b1 );
or ( \3140_b1 , \3133_b1 , w_10536 );
or ( \3140_b0 , \3133_b0 , w_10535 );
not ( w_10535 , w_10537 );
and ( w_10537 , w_10536 , w_10534 );
or ( w_10534 , \3138_b1 , w_10538 );
or ( w_10535 , \3138_b0 , \3139_b0 );
not ( \3139_b0 , w_10539 );
and ( w_10539 , w_10538 , \3139_b1 );
or ( \3156_b1 , \3149_b1 , w_10542 );
or ( \3156_b0 , \3149_b0 , w_10541 );
not ( w_10541 , w_10543 );
and ( w_10543 , w_10542 , w_10540 );
or ( w_10540 , \3154_b1 , w_10544 );
or ( w_10541 , \3154_b0 , \3155_b0 );
not ( \3155_b0 , w_10545 );
and ( w_10545 , w_10544 , \3155_b1 );
or ( \3169_b1 , \3166_b1 , w_10548 );
or ( \3169_b0 , \3166_b0 , w_10547 );
not ( w_10547 , w_10549 );
and ( w_10549 , w_10548 , w_10546 );
or ( w_10546 , \3167_b1 , w_10550 );
or ( w_10547 , \3167_b0 , \3168_b0 );
not ( \3168_b0 , w_10551 );
and ( w_10551 , w_10550 , \3168_b1 );
or ( \3172_b1 , \3157_b1 , w_10554 );
or ( \3172_b0 , \3157_b0 , w_10553 );
not ( w_10553 , w_10555 );
and ( w_10555 , w_10554 , w_10552 );
or ( w_10552 , \3170_b1 , w_10556 );
or ( w_10553 , \3170_b0 , \3171_b0 );
not ( \3171_b0 , w_10557 );
and ( w_10557 , w_10556 , \3171_b1 );
or ( \3180_b1 , \3175_b1 , w_10560 );
or ( \3180_b0 , \3175_b0 , w_10559 );
not ( w_10559 , w_10561 );
and ( w_10561 , w_10560 , w_10558 );
or ( w_10558 , \3178_b1 , w_10562 );
or ( w_10559 , \3178_b0 , \3179_b0 );
not ( \3179_b0 , w_10563 );
and ( w_10563 , w_10562 , \3179_b1 );
or ( \3186_b1 , \3181_b1 , w_10566 );
or ( \3186_b0 , \3181_b0 , w_10565 );
not ( w_10565 , w_10567 );
and ( w_10567 , w_10566 , w_10564 );
or ( w_10564 , \3184_b1 , w_10568 );
or ( w_10565 , \3184_b0 , \3185_b0 );
not ( \3185_b0 , w_10569 );
and ( w_10569 , w_10568 , \3185_b1 );
or ( \3194_b1 , \3189_b1 , w_10572 );
or ( \3194_b0 , \3189_b0 , w_10571 );
not ( w_10571 , w_10573 );
and ( w_10573 , w_10572 , w_10570 );
or ( w_10570 , \3192_b1 , w_10574 );
or ( w_10571 , \3192_b0 , \3193_b0 );
not ( \3193_b0 , w_10575 );
and ( w_10575 , w_10574 , \3193_b1 );
or ( \3208_b1 , \3203_b1 , w_10578 );
or ( \3208_b0 , \3203_b0 , w_10577 );
not ( w_10577 , w_10579 );
and ( w_10579 , w_10578 , w_10576 );
or ( w_10576 , \3206_b1 , w_10580 );
or ( w_10577 , \3206_b0 , \3207_b0 );
not ( \3207_b0 , w_10581 );
and ( w_10581 , w_10580 , \3207_b1 );
or ( \3216_b1 , \3211_b1 , w_10584 );
or ( \3216_b0 , \3211_b0 , w_10583 );
not ( w_10583 , w_10585 );
and ( w_10585 , w_10584 , w_10582 );
or ( w_10582 , \3214_b1 , w_10586 );
or ( w_10583 , \3214_b0 , \3215_b0 );
not ( \3215_b0 , w_10587 );
and ( w_10587 , w_10586 , \3215_b1 );
or ( \3224_b1 , \3219_b1 , w_10590 );
or ( \3224_b0 , \3219_b0 , w_10589 );
not ( w_10589 , w_10591 );
and ( w_10591 , w_10590 , w_10588 );
or ( w_10588 , \3222_b1 , w_10592 );
or ( w_10589 , \3222_b0 , \3223_b0 );
not ( \3223_b0 , w_10593 );
and ( w_10593 , w_10592 , \3223_b1 );
or ( \3244_b1 , \3237_b1 , w_10596 );
or ( \3244_b0 , \3237_b0 , w_10595 );
not ( w_10595 , w_10597 );
and ( w_10597 , w_10596 , w_10594 );
or ( w_10594 , \3242_b1 , w_10598 );
or ( w_10595 , \3242_b0 , \3243_b0 );
not ( \3243_b0 , w_10599 );
and ( w_10599 , w_10598 , \3243_b1 );
or ( \3252_b1 , \3247_b1 , w_10602 );
or ( \3252_b0 , \3247_b0 , w_10601 );
not ( w_10601 , w_10603 );
and ( w_10603 , w_10602 , w_10600 );
or ( w_10600 , \3250_b1 , w_10604 );
or ( w_10601 , \3250_b0 , \3251_b0 );
not ( \3251_b0 , w_10605 );
and ( w_10605 , w_10604 , \3251_b1 );
or ( \3268_b1 , \3261_b1 , w_10608 );
or ( \3268_b0 , \3261_b0 , w_10607 );
not ( w_10607 , w_10609 );
and ( w_10609 , w_10608 , w_10606 );
or ( w_10606 , \3266_b1 , w_10610 );
or ( w_10607 , \3266_b0 , \3267_b0 );
not ( \3267_b0 , w_10611 );
and ( w_10611 , w_10610 , \3267_b1 );
or ( \3282_b1 , \3277_b1 , w_10614 );
or ( \3282_b0 , \3277_b0 , w_10613 );
not ( w_10613 , w_10615 );
and ( w_10615 , w_10614 , w_10612 );
or ( w_10612 , \3280_b1 , w_10616 );
or ( w_10613 , \3280_b0 , \3281_b0 );
not ( \3281_b0 , w_10617 );
and ( w_10617 , w_10616 , \3281_b1 );
or ( \3288_b1 , \3283_b1 , w_10620 );
or ( \3288_b0 , \3283_b0 , w_10619 );
not ( w_10619 , w_10621 );
and ( w_10621 , w_10620 , w_10618 );
or ( w_10618 , \3286_b1 , w_10622 );
or ( w_10619 , \3286_b0 , \3287_b0 );
not ( \3287_b0 , w_10623 );
and ( w_10623 , w_10622 , \3287_b1 );
or ( \3296_b1 , \3291_b1 , w_10626 );
or ( \3296_b0 , \3291_b0 , w_10625 );
not ( w_10625 , w_10627 );
and ( w_10627 , w_10626 , w_10624 );
or ( w_10624 , \3294_b1 , w_10628 );
or ( w_10625 , \3294_b0 , \3295_b0 );
not ( \3295_b0 , w_10629 );
and ( w_10629 , w_10628 , \3295_b1 );
or ( \3311_b1 , \3308_b1 , w_10632 );
or ( \3311_b0 , \3308_b0 , w_10631 );
not ( w_10631 , w_10633 );
and ( w_10633 , w_10632 , w_10630 );
or ( w_10630 , \3309_b1 , w_10634 );
or ( w_10631 , \3309_b0 , \3310_b0 );
not ( \3310_b0 , w_10635 );
and ( w_10635 , w_10634 , \3310_b1 );
or ( \3319_b1 , \3312_b1 , w_10638 );
or ( \3319_b0 , \3312_b0 , w_10637 );
not ( w_10637 , w_10639 );
and ( w_10639 , w_10638 , w_10636 );
or ( w_10636 , \3317_b1 , w_10640 );
or ( w_10637 , \3317_b0 , \3318_b0 );
not ( \3318_b0 , w_10641 );
and ( w_10641 , w_10640 , \3318_b1 );
or ( \3335_b1 , \3328_b1 , w_10644 );
or ( \3335_b0 , \3328_b0 , w_10643 );
not ( w_10643 , w_10645 );
and ( w_10645 , w_10644 , w_10642 );
or ( w_10642 , \3333_b1 , w_10646 );
or ( w_10643 , \3333_b0 , \3334_b0 );
not ( \3334_b0 , w_10647 );
and ( w_10647 , w_10646 , \3334_b1 );
or ( \3343_b1 , \3338_b1 , w_10650 );
or ( \3343_b0 , \3338_b0 , w_10649 );
not ( w_10649 , w_10651 );
and ( w_10651 , w_10650 , w_10648 );
or ( w_10648 , \3341_b1 , w_10652 );
or ( w_10649 , \3341_b0 , \3342_b0 );
not ( \3342_b0 , w_10653 );
and ( w_10653 , w_10652 , \3342_b1 );
or ( \3349_b1 , \3344_b1 , w_10656 );
or ( \3349_b0 , \3344_b0 , w_10655 );
not ( w_10655 , w_10657 );
and ( w_10657 , w_10656 , w_10654 );
or ( w_10654 , \3347_b1 , w_10658 );
or ( w_10655 , \3347_b0 , \3348_b0 );
not ( \3348_b0 , w_10659 );
and ( w_10659 , w_10658 , \3348_b1 );
or ( \3357_b1 , \3352_b1 , w_10662 );
or ( \3357_b0 , \3352_b0 , w_10661 );
not ( w_10661 , w_10663 );
and ( w_10663 , w_10662 , w_10660 );
or ( w_10660 , \3355_b1 , w_10664 );
or ( w_10661 , \3355_b0 , \3356_b0 );
not ( \3356_b0 , w_10665 );
and ( w_10665 , w_10664 , \3356_b1 );
or ( \3383_b1 , \3376_b1 , w_10668 );
or ( \3383_b0 , \3376_b0 , w_10667 );
not ( w_10667 , w_10669 );
and ( w_10669 , w_10668 , w_10666 );
or ( w_10666 , \3381_b1 , w_10670 );
or ( w_10667 , \3381_b0 , \3382_b0 );
not ( \3382_b0 , w_10671 );
and ( w_10671 , w_10670 , \3382_b1 );
or ( \3399_b1 , \3392_b1 , w_10674 );
or ( \3399_b0 , \3392_b0 , w_10673 );
not ( w_10673 , w_10675 );
and ( w_10675 , w_10674 , w_10672 );
or ( w_10672 , \3397_b1 , w_10676 );
or ( w_10673 , \3397_b0 , \3398_b0 );
not ( \3398_b0 , w_10677 );
and ( w_10677 , w_10676 , \3398_b1 );
or ( \3415_b1 , \3408_b1 , w_10680 );
or ( \3415_b0 , \3408_b0 , w_10679 );
not ( w_10679 , w_10681 );
and ( w_10681 , w_10680 , w_10678 );
or ( w_10678 , \3413_b1 , w_10682 );
or ( w_10679 , \3413_b0 , \3414_b0 );
not ( \3414_b0 , w_10683 );
and ( w_10683 , w_10682 , \3414_b1 );
or ( \3421_b1 , \3416_b1 , w_10686 );
or ( \3421_b0 , \3416_b0 , w_10685 );
not ( w_10685 , w_10687 );
and ( w_10687 , w_10686 , w_10684 );
or ( w_10684 , \3419_b1 , w_10688 );
or ( w_10685 , \3419_b0 , \3420_b0 );
not ( \3420_b0 , w_10689 );
and ( w_10689 , w_10688 , \3420_b1 );
or ( \3427_b1 , \3422_b1 , w_10692 );
or ( \3427_b0 , \3422_b0 , w_10691 );
not ( w_10691 , w_10693 );
and ( w_10693 , w_10692 , w_10690 );
or ( w_10690 , \3425_b1 , w_10694 );
or ( w_10691 , \3425_b0 , \3426_b0 );
not ( \3426_b0 , w_10695 );
and ( w_10695 , w_10694 , \3426_b1 );
or ( \3435_b1 , \3430_b1 , w_10698 );
or ( \3435_b0 , \3430_b0 , w_10697 );
not ( w_10697 , w_10699 );
and ( w_10699 , w_10698 , w_10696 );
or ( w_10696 , \3433_b1 , w_10700 );
or ( w_10697 , \3433_b0 , \3434_b0 );
not ( \3434_b0 , w_10701 );
and ( w_10701 , w_10700 , \3434_b1 );
or ( \3452_b1 , \3449_b1 , w_10704 );
or ( \3452_b0 , \3449_b0 , w_10703 );
not ( w_10703 , w_10705 );
and ( w_10705 , w_10704 , w_10702 );
or ( w_10702 , \3450_b1 , w_10706 );
or ( w_10703 , \3450_b0 , \3451_b0 );
not ( \3451_b0 , w_10707 );
and ( w_10707 , w_10706 , \3451_b1 );
or ( \3469_b1 , \3462_b1 , w_10710 );
or ( \3469_b0 , \3462_b0 , w_10709 );
not ( w_10709 , w_10711 );
and ( w_10711 , w_10710 , w_10708 );
or ( w_10708 , \3467_b1 , w_10712 );
or ( w_10709 , \3467_b0 , \3468_b0 );
not ( \3468_b0 , w_10713 );
and ( w_10713 , w_10712 , \3468_b1 );
or ( \3472_b1 , \3453_b1 , w_10716 );
or ( \3472_b0 , \3453_b0 , w_10715 );
not ( w_10715 , w_10717 );
and ( w_10717 , w_10716 , w_10714 );
or ( w_10714 , \3470_b1 , w_10718 );
or ( w_10715 , \3470_b0 , \3471_b0 );
not ( \3471_b0 , w_10719 );
and ( w_10719 , w_10718 , \3471_b1 );
or ( \3480_b1 , \3475_b1 , w_10722 );
or ( \3480_b0 , \3475_b0 , w_10721 );
not ( w_10721 , w_10723 );
and ( w_10723 , w_10722 , w_10720 );
or ( w_10720 , \3478_b1 , w_10724 );
or ( w_10721 , \3478_b0 , \3479_b0 );
not ( \3479_b0 , w_10725 );
and ( w_10725 , w_10724 , \3479_b1 );
or ( \3488_b1 , \3483_b1 , w_10728 );
or ( \3488_b0 , \3483_b0 , w_10727 );
not ( w_10727 , w_10729 );
and ( w_10729 , w_10728 , w_10726 );
or ( w_10726 , \3486_b1 , w_10730 );
or ( w_10727 , \3486_b0 , \3487_b0 );
not ( \3487_b0 , w_10731 );
and ( w_10731 , w_10730 , \3487_b1 );
or ( \3508_b1 , \3501_b1 , w_10734 );
or ( \3508_b0 , \3501_b0 , w_10733 );
not ( w_10733 , w_10735 );
and ( w_10735 , w_10734 , w_10732 );
or ( w_10732 , \3506_b1 , w_10736 );
or ( w_10733 , \3506_b0 , \3507_b0 );
not ( \3507_b0 , w_10737 );
and ( w_10737 , w_10736 , \3507_b1 );
or ( \3524_b1 , \3517_b1 , w_10740 );
or ( \3524_b0 , \3517_b0 , w_10739 );
not ( w_10739 , w_10741 );
and ( w_10741 , w_10740 , w_10738 );
or ( w_10738 , \3522_b1 , w_10742 );
or ( w_10739 , \3522_b0 , \3523_b0 );
not ( \3523_b0 , w_10743 );
and ( w_10743 , w_10742 , \3523_b1 );
or ( \3532_b1 , \3527_b1 , w_10746 );
or ( \3532_b0 , \3527_b0 , w_10745 );
not ( w_10745 , w_10747 );
and ( w_10747 , w_10746 , w_10744 );
or ( w_10744 , \3530_b1 , w_10748 );
or ( w_10745 , \3530_b0 , \3531_b0 );
not ( \3531_b0 , w_10749 );
and ( w_10749 , w_10748 , \3531_b1 );
or ( \3540_b1 , \3535_b1 , w_10752 );
or ( \3540_b0 , \3535_b0 , w_10751 );
not ( w_10751 , w_10753 );
and ( w_10753 , w_10752 , w_10750 );
or ( w_10750 , \3538_b1 , w_10754 );
or ( w_10751 , \3538_b0 , \3539_b0 );
not ( \3539_b0 , w_10755 );
and ( w_10755 , w_10754 , \3539_b1 );
or ( \3557_b1 , \3550_b1 , w_10758 );
or ( \3557_b0 , \3550_b0 , w_10757 );
not ( w_10757 , w_10759 );
and ( w_10759 , w_10758 , w_10756 );
or ( w_10756 , \3555_b1 , w_10760 );
or ( w_10757 , \3555_b0 , \3556_b0 );
not ( \3556_b0 , w_10761 );
and ( w_10761 , w_10760 , \3556_b1 );
or ( \3565_b1 , \3560_b1 , w_10764 );
or ( \3565_b0 , \3560_b0 , w_10763 );
not ( w_10763 , w_10765 );
and ( w_10765 , w_10764 , w_10762 );
or ( w_10762 , \3563_b1 , w_10766 );
or ( w_10763 , \3563_b0 , \3564_b0 );
not ( \3564_b0 , w_10767 );
and ( w_10767 , w_10766 , \3564_b1 );
or ( \3573_b1 , \3568_b1 , w_10770 );
or ( \3573_b0 , \3568_b0 , w_10769 );
not ( w_10769 , w_10771 );
and ( w_10771 , w_10770 , w_10768 );
or ( w_10768 , \3571_b1 , w_10772 );
or ( w_10769 , \3571_b0 , \3572_b0 );
not ( \3572_b0 , w_10773 );
and ( w_10773 , w_10772 , \3572_b1 );
or ( \3589_b1 , \3586_b1 , w_10776 );
or ( \3589_b0 , \3586_b0 , w_10775 );
not ( w_10775 , w_10777 );
and ( w_10777 , w_10776 , w_10774 );
or ( w_10774 , \3587_b1 , w_10778 );
or ( w_10775 , \3587_b0 , \3588_b0 );
not ( \3588_b0 , w_10779 );
and ( w_10779 , w_10778 , \3588_b1 );
or ( \3605_b1 , \3598_b1 , w_10782 );
or ( \3605_b0 , \3598_b0 , w_10781 );
not ( w_10781 , w_10783 );
and ( w_10783 , w_10782 , w_10780 );
or ( w_10780 , \3603_b1 , w_10784 );
or ( w_10781 , \3603_b0 , \3604_b0 );
not ( \3604_b0 , w_10785 );
and ( w_10785 , w_10784 , \3604_b1 );
or ( \3611_b1 , \3606_b1 , w_10788 );
or ( \3611_b0 , \3606_b0 , w_10787 );
not ( w_10787 , w_10789 );
and ( w_10789 , w_10788 , w_10786 );
or ( w_10786 , \3609_b1 , w_10790 );
or ( w_10787 , \3609_b0 , \3610_b0 );
not ( \3610_b0 , w_10791 );
and ( w_10791 , w_10790 , \3610_b1 );
or ( \3619_b1 , \3614_b1 , w_10794 );
or ( \3619_b0 , \3614_b0 , w_10793 );
not ( w_10793 , w_10795 );
and ( w_10795 , w_10794 , w_10792 );
or ( w_10792 , \3617_b1 , w_10796 );
or ( w_10793 , \3617_b0 , \3618_b0 );
not ( \3618_b0 , w_10797 );
and ( w_10797 , w_10796 , \3618_b1 );
or ( \3639_b1 , \3632_b1 , w_10800 );
or ( \3639_b0 , \3632_b0 , w_10799 );
not ( w_10799 , w_10801 );
and ( w_10801 , w_10800 , w_10798 );
or ( w_10798 , \3637_b1 , w_10802 );
or ( w_10799 , \3637_b0 , \3638_b0 );
not ( \3638_b0 , w_10803 );
and ( w_10803 , w_10802 , \3638_b1 );
or ( \3653_b1 , \3648_b1 , w_10806 );
or ( \3653_b0 , \3648_b0 , w_10805 );
not ( w_10805 , w_10807 );
and ( w_10807 , w_10806 , w_10804 );
or ( w_10804 , \3651_b1 , w_10808 );
or ( w_10805 , \3651_b0 , \3652_b0 );
not ( \3652_b0 , w_10809 );
and ( w_10809 , w_10808 , \3652_b1 );
or ( \3661_b1 , \3656_b1 , w_10812 );
or ( \3661_b0 , \3656_b0 , w_10811 );
not ( w_10811 , w_10813 );
and ( w_10813 , w_10812 , w_10810 );
or ( w_10810 , \3659_b1 , w_10814 );
or ( w_10811 , \3659_b0 , \3660_b0 );
not ( \3660_b0 , w_10815 );
and ( w_10815 , w_10814 , \3660_b1 );
or ( \3676_b1 , \3673_b1 , w_10818 );
or ( \3676_b0 , \3673_b0 , w_10817 );
not ( w_10817 , w_10819 );
and ( w_10819 , w_10818 , w_10816 );
or ( w_10816 , \3674_b1 , w_10820 );
or ( w_10817 , \3674_b0 , \3675_b0 );
not ( \3675_b0 , w_10821 );
and ( w_10821 , w_10820 , \3675_b1 );
or ( \3684_b1 , \3677_b1 , w_10824 );
or ( \3684_b0 , \3677_b0 , w_10823 );
not ( w_10823 , w_10825 );
and ( w_10825 , w_10824 , w_10822 );
or ( w_10822 , \3682_b1 , w_10826 );
or ( w_10823 , \3682_b0 , \3683_b0 );
not ( \3683_b0 , w_10827 );
and ( w_10827 , w_10826 , \3683_b1 );
or ( \3692_b1 , \3687_b1 , w_10830 );
or ( \3692_b0 , \3687_b0 , w_10829 );
not ( w_10829 , w_10831 );
and ( w_10831 , w_10830 , w_10828 );
or ( w_10828 , \3690_b1 , w_10832 );
or ( w_10829 , \3690_b0 , \3691_b0 );
not ( \3691_b0 , w_10833 );
and ( w_10833 , w_10832 , \3691_b1 );
or ( \3718_b1 , \3711_b1 , w_10836 );
or ( \3718_b0 , \3711_b0 , w_10835 );
not ( w_10835 , w_10837 );
and ( w_10837 , w_10836 , w_10834 );
or ( w_10834 , \3716_b1 , w_10838 );
or ( w_10835 , \3716_b0 , \3717_b0 );
not ( \3717_b0 , w_10839 );
and ( w_10839 , w_10838 , \3717_b1 );
or ( \3726_b1 , \3721_b1 , w_10842 );
or ( \3726_b0 , \3721_b0 , w_10841 );
not ( w_10841 , w_10843 );
and ( w_10843 , w_10842 , w_10840 );
or ( w_10840 , \3724_b1 , w_10844 );
or ( w_10841 , \3724_b0 , \3725_b0 );
not ( \3725_b0 , w_10845 );
and ( w_10845 , w_10844 , \3725_b1 );
or ( \3746_b1 , \3739_b1 , w_10848 );
or ( \3746_b0 , \3739_b0 , w_10847 );
not ( w_10847 , w_10849 );
and ( w_10849 , w_10848 , w_10846 );
or ( w_10846 , \3744_b1 , w_10850 );
or ( w_10847 , \3744_b0 , \3745_b0 );
not ( \3745_b0 , w_10851 );
and ( w_10851 , w_10850 , \3745_b1 );
or ( \3754_b1 , \3749_b1 , w_10854 );
or ( \3754_b0 , \3749_b0 , w_10853 );
not ( w_10853 , w_10855 );
and ( w_10855 , w_10854 , w_10852 );
or ( w_10852 , \3752_b1 , w_10856 );
or ( w_10853 , \3752_b0 , \3753_b0 );
not ( \3753_b0 , w_10857 );
and ( w_10857 , w_10856 , \3753_b1 );
or ( \3769_b1 , \3766_b1 , w_10860 );
or ( \3769_b0 , \3766_b0 , w_10859 );
not ( w_10859 , w_10861 );
and ( w_10861 , w_10860 , w_10858 );
or ( w_10858 , \3767_b1 , w_10862 );
or ( w_10859 , \3767_b0 , \3768_b0 );
not ( \3768_b0 , w_10863 );
and ( w_10863 , w_10862 , \3768_b1 );
or ( \3775_b1 , \3770_b1 , w_10866 );
or ( \3775_b0 , \3770_b0 , w_10865 );
not ( w_10865 , w_10867 );
and ( w_10867 , w_10866 , w_10864 );
or ( w_10864 , \3773_b1 , w_10868 );
or ( w_10865 , \3773_b0 , \3774_b0 );
not ( \3774_b0 , w_10869 );
and ( w_10869 , w_10868 , \3774_b1 );
or ( \3799_b1 , \3794_b1 , w_10872 );
or ( \3799_b0 , \3794_b0 , w_10871 );
not ( w_10871 , w_10873 );
and ( w_10873 , w_10872 , w_10870 );
or ( w_10870 , \3797_b1 , w_10874 );
or ( w_10871 , \3797_b0 , \3798_b0 );
not ( \3798_b0 , w_10875 );
and ( w_10875 , w_10874 , \3798_b1 );
or ( \3816_b1 , \3809_b1 , w_10878 );
or ( \3816_b0 , \3809_b0 , w_10877 );
not ( w_10877 , w_10879 );
and ( w_10879 , w_10878 , w_10876 );
or ( w_10876 , \3814_b1 , w_10880 );
or ( w_10877 , \3814_b0 , \3815_b0 );
not ( \3815_b0 , w_10881 );
and ( w_10881 , w_10880 , \3815_b1 );
or ( \3830_b1 , \3827_b1 , w_10884 );
or ( \3830_b0 , \3827_b0 , w_10883 );
not ( w_10883 , w_10885 );
and ( w_10885 , w_10884 , w_10882 );
or ( w_10882 , \3828_b1 , w_10886 );
or ( w_10883 , \3828_b0 , \3829_b0 );
not ( \3829_b0 , w_10887 );
and ( w_10887 , w_10886 , \3829_b1 );
endmodule

