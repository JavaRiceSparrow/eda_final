// ...
module top(\a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,
		\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,
		\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,
		\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,\a[0]_b1 ,\a[0]_b0 ,\b[15]_b1 ,\b[15]_b0 ,\b[14]_b1 ,\b[14]_b0 ,
		\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,\b[10]_b0 ,\b[9]_b1 ,
		\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,\b[5]_b1 ,\b[5]_b0 ,
		\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,\b[1]_b0 ,\b[0]_b1 ,
		\b[0]_b0 ,\c[15]_b1 ,\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,
		\c[11]_b1 ,\c[11]_b0 ,\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,
		\c[7]_b0 ,\c[6]_b1 ,\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,
		\c[2]_b1 ,\c[2]_b0 ,\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,
		\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,
		\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,
		\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,
		\d[0]_b1 ,\d[0]_b0 ,\o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,
		\o[28]_b0 ,\o[27]_b1 ,\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,
		\o[23]_b1 ,\o[23]_b0 ,\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,
		\o[19]_b0 ,\o[18]_b1 ,\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,
		\o[14]_b1 ,\o[14]_b0 ,\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,
		\o[10]_b0 ,\o[9]_b1 ,\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,
		\o[5]_b1 ,\o[5]_b0 ,\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,
		\o[1]_b0 ,\o[0]_b1 ,\o[0]_b0 );
input \a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,
		\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,
		\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,
		\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,\a[0]_b1 ,\a[0]_b0 ,\b[15]_b1 ,\b[15]_b0 ,\b[14]_b1 ,\b[14]_b0 ,
		\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,\b[10]_b0 ,\b[9]_b1 ,
		\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,\b[5]_b1 ,\b[5]_b0 ,
		\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,\b[1]_b0 ,\b[0]_b1 ,
		\b[0]_b0 ,\c[15]_b1 ,\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,
		\c[11]_b1 ,\c[11]_b0 ,\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,
		\c[7]_b0 ,\c[6]_b1 ,\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,
		\c[2]_b1 ,\c[2]_b0 ,\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,
		\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,
		\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,
		\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,
		\d[0]_b1 ,\d[0]_b0 ;
output \o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,\o[28]_b0 ,\o[27]_b1 ,
		\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,\o[23]_b1 ,\o[23]_b0 ,
		\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,\o[19]_b0 ,\o[18]_b1 ,
		\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,\o[14]_b1 ,\o[14]_b0 ,
		\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,\o[10]_b0 ,\o[9]_b1 ,
		\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,\o[5]_b1 ,\o[5]_b0 ,
		\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,\o[1]_b0 ,\o[0]_b1 ,
		\o[0]_b0 ;

wire \97_n22[15]_b1 , \97_n22[15]_b0 , \98_n22[14]_b1 , \98_n22[14]_b0 , \99_n22[13]_b1 , \99_n22[13]_b0 , \100_n22[12]_b1 , \100_n22[12]_b0 , \101_n22[11]_b1 , \101_n22[11]_b0 , 
		\102_n22[10]_b1 , \102_n22[10]_b0 , \103_n22[9]_b1 , \103_n22[9]_b0 , \104_n22[8]_b1 , \104_n22[8]_b0 , \105_n22[7]_b1 , \105_n22[7]_b0 , \106_n22[6]_b1 , \106_n22[6]_b0 , 
		\107_n22[5]_b1 , \107_n22[5]_b0 , \108_n22[4]_b1 , \108_n22[4]_b0 , \109_n22[3]_b1 , \109_n22[3]_b0 , \110_n22[2]_b1 , \110_n22[2]_b0 , \111_n22[1]_b1 , \111_n22[1]_b0 , 
		\112_n22[0]_b1 , \112_n22[0]_b0 , \113_ZERO_b1 , \113_ZERO_b0 , \114_ZERO_b1 , \114_ZERO_b0 , \115_b1 , \115_b0 , \116_b1 , \116_b0 , 
		\117_b1 , \117_b0 , \118_b1 , \118_b0 , \119_b1 , \119_b0 , \120_b1 , \120_b0 , \121_b1 , \121_b0 , 
		\122_b1 , \122_b0 , \123_b1 , \123_b0 , \124_b1 , \124_b0 , \125_b1 , \125_b0 , \126_b1 , \126_b0 , 
		\127_b1 , \127_b0 , \128_b1 , \128_b0 , \129_b1 , \129_b0 , \130_b1 , \130_b0 , \131_b1 , \131_b0 , 
		\132_b1 , \132_b0 , \133_b1 , \133_b0 , \134_b1 , \134_b0 , \135_b1 , \135_b0 , \136_b1 , \136_b0 , 
		\137_b1 , \137_b0 , \138_b1 , \138_b0 , \139_b1 , \139_b0 , \140_b1 , \140_b0 , \141_b1 , \141_b0 , 
		\142_b1 , \142_b0 , \143_b1 , \143_b0 , \144_b1 , \144_b0 , \145_b1 , \145_b0 , \146_b1 , \146_b0 , 
		\147_b1 , \147_b0 , \148_b1 , \148_b0 , \149_b1 , \149_b0 , \150_b1 , \150_b0 , \151_b1 , \151_b0 , 
		\152_b1 , \152_b0 , \153_b1 , \153_b0 , \154_b1 , \154_b0 , \155_ONE_b1 , \155_ONE_b0 , \156_A[0]_b1 , \156_A[0]_b0 , 
		\157_B[0]_b1 , \157_B[0]_b0 , \158_b1 , \158_b0 , \159_Z[0]_b1 , \159_Z[0]_b0 , \160_b1 , \160_b0 , \161_A[1]_b1 , \161_A[1]_b0 , 
		\162_b1 , \162_b0 , \163_B[1]_b1 , \163_B[1]_b0 , \164_b1 , \164_b0 , \165_b1 , \165_b0 , \166_Z[1]_b1 , \166_Z[1]_b0 , 
		\167_A[2]_b1 , \167_A[2]_b0 , \168_b1 , \168_b0 , \169_b1 , \169_b0 , \170_b1 , \170_b0 , \171_b1 , \171_b0 , 
		\172_b1 , \172_b0 , \173_B[2]_b1 , \173_B[2]_b0 , \174_b1 , \174_b0 , \175_b1 , \175_b0 , \176_Z[2]_b1 , \176_Z[2]_b0 , 
		\177_A[3]_b1 , \177_A[3]_b0 , \178_b1 , \178_b0 , \179_b1 , \179_b0 , \180_b1 , \180_b0 , \181_b1 , \181_b0 , 
		\182_b1 , \182_b0 , \183_b1 , \183_b0 , \184_b1 , \184_b0 , \185_b1 , \185_b0 , \186_b1 , \186_b0 , 
		\187_b1 , \187_b0 , \188_b1 , \188_b0 , \189_B[3]_b1 , \189_B[3]_b0 , \190_b1 , \190_b0 , \191_b1 , \191_b0 , 
		\192_Z[3]_b1 , \192_Z[3]_b0 , \193_A[4]_b1 , \193_A[4]_b0 , \194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , 
		\197_b1 , \197_b0 , \198_b1 , \198_b0 , \199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , 
		\202_b1 , \202_b0 , \203_b1 , \203_b0 , \204_b1 , \204_b0 , \205_b1 , \205_b0 , \206_b1 , \206_b0 , 
		\207_b1 , \207_b0 , \208_b1 , \208_b0 , \209_b1 , \209_b0 , \210_b1 , \210_b0 , \211_B[4]_b1 , \211_B[4]_b0 , 
		\212_b1 , \212_b0 , \213_b1 , \213_b0 , \214_Z[4]_b1 , \214_Z[4]_b0 , \215_A[5]_b1 , \215_A[5]_b0 , \216_b1 , \216_b0 , 
		\217_b1 , \217_b0 , \218_b1 , \218_b0 , \219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , 
		\222_b1 , \222_b0 , \223_b1 , \223_b0 , \224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , 
		\227_b1 , \227_b0 , \228_b1 , \228_b0 , \229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , 
		\232_b1 , \232_b0 , \233_b1 , \233_b0 , \234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , 
		\237_b1 , \237_b0 , \238_b1 , \238_b0 , \239_B[5]_b1 , \239_B[5]_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , 
		\242_Z[5]_b1 , \242_Z[5]_b0 , \243_A[6]_b1 , \243_A[6]_b0 , \244_b1 , \244_b0 , \245_b1 , \245_b0 , \246_b1 , \246_b0 , 
		\247_b1 , \247_b0 , \248_b1 , \248_b0 , \249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , 
		\252_b1 , \252_b0 , \253_b1 , \253_b0 , \254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , 
		\257_b1 , \257_b0 , \258_b1 , \258_b0 , \259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , 
		\262_b1 , \262_b0 , \263_b1 , \263_b0 , \264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , 
		\267_b1 , \267_b0 , \268_b1 , \268_b0 , \269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , 
		\272_b1 , \272_b0 , \273_B[6]_b1 , \273_B[6]_b0 , \274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_Z[6]_b1 , \276_Z[6]_b0 , 
		\277_A[7]_b1 , \277_A[7]_b0 , \278_b1 , \278_b0 , \279_b1 , \279_b0 , \280_b1 , \280_b0 , \281_b1 , \281_b0 , 
		\282_b1 , \282_b0 , \283_b1 , \283_b0 , \284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , 
		\287_b1 , \287_b0 , \288_b1 , \288_b0 , \289_b1 , \289_b0 , \290_b1 , \290_b0 , \291_b1 , \291_b0 , 
		\292_b1 , \292_b0 , \293_b1 , \293_b0 , \294_b1 , \294_b0 , \295_b1 , \295_b0 , \296_b1 , \296_b0 , 
		\297_b1 , \297_b0 , \298_b1 , \298_b0 , \299_b1 , \299_b0 , \300_b1 , \300_b0 , \301_b1 , \301_b0 , 
		\302_b1 , \302_b0 , \303_b1 , \303_b0 , \304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , 
		\307_b1 , \307_b0 , \308_b1 , \308_b0 , \309_b1 , \309_b0 , \310_b1 , \310_b0 , \311_b1 , \311_b0 , 
		\312_b1 , \312_b0 , \313_B[7]_b1 , \313_B[7]_b0 , \314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_Z[7]_b1 , \316_Z[7]_b0 , 
		\317_A[8]_b1 , \317_A[8]_b0 , \318_b1 , \318_b0 , \319_b1 , \319_b0 , \320_b1 , \320_b0 , \321_b1 , \321_b0 , 
		\322_b1 , \322_b0 , \323_b1 , \323_b0 , \324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , 
		\327_b1 , \327_b0 , \328_b1 , \328_b0 , \329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_b1 , \331_b0 , 
		\332_b1 , \332_b0 , \333_b1 , \333_b0 , \334_b1 , \334_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , 
		\337_b1 , \337_b0 , \338_b1 , \338_b0 , \339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_b1 , \341_b0 , 
		\342_b1 , \342_b0 , \343_b1 , \343_b0 , \344_b1 , \344_b0 , \345_b1 , \345_b0 , \346_b1 , \346_b0 , 
		\347_b1 , \347_b0 , \348_b1 , \348_b0 , \349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , 
		\352_b1 , \352_b0 , \353_b1 , \353_b0 , \354_b1 , \354_b0 , \355_b1 , \355_b0 , \356_b1 , \356_b0 , 
		\357_b1 , \357_b0 , \358_b1 , \358_b0 , \359_B[8]_b1 , \359_B[8]_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , 
		\362_Z[8]_b1 , \362_Z[8]_b0 , \363_A[9]_b1 , \363_A[9]_b0 , \364_b1 , \364_b0 , \365_b1 , \365_b0 , \366_b1 , \366_b0 , 
		\367_b1 , \367_b0 , \368_b1 , \368_b0 , \369_b1 , \369_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , 
		\372_b1 , \372_b0 , \373_b1 , \373_b0 , \374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , 
		\377_b1 , \377_b0 , \378_b1 , \378_b0 , \379_b1 , \379_b0 , \380_b1 , \380_b0 , \381_b1 , \381_b0 , 
		\382_b1 , \382_b0 , \383_b1 , \383_b0 , \384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , 
		\387_b1 , \387_b0 , \388_b1 , \388_b0 , \389_b1 , \389_b0 , \390_b1 , \390_b0 , \391_b1 , \391_b0 , 
		\392_b1 , \392_b0 , \393_b1 , \393_b0 , \394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , 
		\397_b1 , \397_b0 , \398_b1 , \398_b0 , \399_b1 , \399_b0 , \400_b1 , \400_b0 , \401_b1 , \401_b0 , 
		\402_b1 , \402_b0 , \403_b1 , \403_b0 , \404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , 
		\407_b1 , \407_b0 , \408_b1 , \408_b0 , \409_b1 , \409_b0 , \410_b1 , \410_b0 , \411_B[9]_b1 , \411_B[9]_b0 , 
		\412_b1 , \412_b0 , \413_b1 , \413_b0 , \414_Z[9]_b1 , \414_Z[9]_b0 , \415_A[10]_b1 , \415_A[10]_b0 , \416_b1 , \416_b0 , 
		\417_b1 , \417_b0 , \418_b1 , \418_b0 , \419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , 
		\422_b1 , \422_b0 , \423_b1 , \423_b0 , \424_b1 , \424_b0 , \425_b1 , \425_b0 , \426_b1 , \426_b0 , 
		\427_b1 , \427_b0 , \428_b1 , \428_b0 , \429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , 
		\432_b1 , \432_b0 , \433_b1 , \433_b0 , \434_b1 , \434_b0 , \435_b1 , \435_b0 , \436_b1 , \436_b0 , 
		\437_b1 , \437_b0 , \438_b1 , \438_b0 , \439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , 
		\442_b1 , \442_b0 , \443_b1 , \443_b0 , \444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_b1 , \446_b0 , 
		\447_b1 , \447_b0 , \448_b1 , \448_b0 , \449_b1 , \449_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , 
		\452_b1 , \452_b0 , \453_b1 , \453_b0 , \454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_b1 , \456_b0 , 
		\457_b1 , \457_b0 , \458_b1 , \458_b0 , \459_b1 , \459_b0 , \460_b1 , \460_b0 , \461_b1 , \461_b0 , 
		\462_b1 , \462_b0 , \463_b1 , \463_b0 , \464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , 
		\467_b1 , \467_b0 , \468_b1 , \468_b0 , \469_B[10]_b1 , \469_B[10]_b0 , \470_b1 , \470_b0 , \471_b1 , \471_b0 , 
		\472_Z[10]_b1 , \472_Z[10]_b0 , \473_A[11]_b1 , \473_A[11]_b0 , \474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , 
		\477_b1 , \477_b0 , \478_b1 , \478_b0 , \479_b1 , \479_b0 , \480_b1 , \480_b0 , \481_b1 , \481_b0 , 
		\482_b1 , \482_b0 , \483_b1 , \483_b0 , \484_b1 , \484_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , 
		\487_b1 , \487_b0 , \488_b1 , \488_b0 , \489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , 
		\492_b1 , \492_b0 , \493_b1 , \493_b0 , \494_b1 , \494_b0 , \495_b1 , \495_b0 , \496_b1 , \496_b0 , 
		\497_b1 , \497_b0 , \498_b1 , \498_b0 , \499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , 
		\502_b1 , \502_b0 , \503_b1 , \503_b0 , \504_b1 , \504_b0 , \505_b1 , \505_b0 , \506_b1 , \506_b0 , 
		\507_b1 , \507_b0 , \508_b1 , \508_b0 , \509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , 
		\512_b1 , \512_b0 , \513_b1 , \513_b0 , \514_b1 , \514_b0 , \515_b1 , \515_b0 , \516_b1 , \516_b0 , 
		\517_b1 , \517_b0 , \518_b1 , \518_b0 , \519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , 
		\522_b1 , \522_b0 , \523_b1 , \523_b0 , \524_b1 , \524_b0 , \525_b1 , \525_b0 , \526_b1 , \526_b0 , 
		\527_b1 , \527_b0 , \528_b1 , \528_b0 , \529_b1 , \529_b0 , \530_b1 , \530_b0 , \531_b1 , \531_b0 , 
		\532_b1 , \532_b0 , \533_B[11]_b1 , \533_B[11]_b0 , \534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_Z[11]_b1 , \536_Z[11]_b0 , 
		\537_A[12]_b1 , \537_A[12]_b0 , \538_b1 , \538_b0 , \539_b1 , \539_b0 , \540_b1 , \540_b0 , \541_b1 , \541_b0 , 
		\542_b1 , \542_b0 , \543_b1 , \543_b0 , \544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , 
		\547_b1 , \547_b0 , \548_b1 , \548_b0 , \549_b1 , \549_b0 , \550_b1 , \550_b0 , \551_b1 , \551_b0 , 
		\552_b1 , \552_b0 , \553_b1 , \553_b0 , \554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , 
		\557_b1 , \557_b0 , \558_b1 , \558_b0 , \559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_b1 , \561_b0 , 
		\562_b1 , \562_b0 , \563_b1 , \563_b0 , \564_b1 , \564_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , 
		\567_b1 , \567_b0 , \568_b1 , \568_b0 , \569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_b1 , \571_b0 , 
		\572_b1 , \572_b0 , \573_b1 , \573_b0 , \574_b1 , \574_b0 , \575_b1 , \575_b0 , \576_b1 , \576_b0 , 
		\577_b1 , \577_b0 , \578_b1 , \578_b0 , \579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , 
		\582_b1 , \582_b0 , \583_b1 , \583_b0 , \584_b1 , \584_b0 , \585_b1 , \585_b0 , \586_b1 , \586_b0 , 
		\587_b1 , \587_b0 , \588_b1 , \588_b0 , \589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , 
		\592_b1 , \592_b0 , \593_b1 , \593_b0 , \594_b1 , \594_b0 , \595_b1 , \595_b0 , \596_b1 , \596_b0 , 
		\597_b1 , \597_b0 , \598_b1 , \598_b0 , \599_b1 , \599_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , 
		\602_b1 , \602_b0 , \603_B[12]_b1 , \603_B[12]_b0 , \604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_Z[12]_b1 , \606_Z[12]_b0 , 
		\607_A[13]_b1 , \607_A[13]_b0 , \608_b1 , \608_b0 , \609_b1 , \609_b0 , \610_b1 , \610_b0 , \611_b1 , \611_b0 , 
		\612_b1 , \612_b0 , \613_b1 , \613_b0 , \614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , 
		\617_b1 , \617_b0 , \618_b1 , \618_b0 , \619_b1 , \619_b0 , \620_b1 , \620_b0 , \621_b1 , \621_b0 , 
		\622_b1 , \622_b0 , \623_b1 , \623_b0 , \624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , 
		\627_b1 , \627_b0 , \628_b1 , \628_b0 , \629_b1 , \629_b0 , \630_b1 , \630_b0 , \631_b1 , \631_b0 , 
		\632_b1 , \632_b0 , \633_b1 , \633_b0 , \634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , 
		\637_b1 , \637_b0 , \638_b1 , \638_b0 , \639_b1 , \639_b0 , \640_b1 , \640_b0 , \641_b1 , \641_b0 , 
		\642_b1 , \642_b0 , \643_b1 , \643_b0 , \644_b1 , \644_b0 , \645_b1 , \645_b0 , \646_b1 , \646_b0 , 
		\647_b1 , \647_b0 , \648_b1 , \648_b0 , \649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , 
		\652_b1 , \652_b0 , \653_b1 , \653_b0 , \654_b1 , \654_b0 , \655_b1 , \655_b0 , \656_b1 , \656_b0 , 
		\657_b1 , \657_b0 , \658_b1 , \658_b0 , \659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , 
		\662_b1 , \662_b0 , \663_b1 , \663_b0 , \664_b1 , \664_b0 , \665_b1 , \665_b0 , \666_b1 , \666_b0 , 
		\667_b1 , \667_b0 , \668_b1 , \668_b0 , \669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , 
		\672_b1 , \672_b0 , \673_b1 , \673_b0 , \674_b1 , \674_b0 , \675_b1 , \675_b0 , \676_b1 , \676_b0 , 
		\677_b1 , \677_b0 , \678_b1 , \678_b0 , \679_B[13]_b1 , \679_B[13]_b0 , \680_b1 , \680_b0 , \681_b1 , \681_b0 , 
		\682_Z[13]_b1 , \682_Z[13]_b0 , \683_A[14]_b1 , \683_A[14]_b0 , \684_b1 , \684_b0 , \685_b1 , \685_b0 , \686_b1 , \686_b0 , 
		\687_b1 , \687_b0 , \688_b1 , \688_b0 , \689_b1 , \689_b0 , \690_b1 , \690_b0 , \691_b1 , \691_b0 , 
		\692_b1 , \692_b0 , \693_b1 , \693_b0 , \694_b1 , \694_b0 , \695_b1 , \695_b0 , \696_b1 , \696_b0 , 
		\697_b1 , \697_b0 , \698_b1 , \698_b0 , \699_b1 , \699_b0 , \700_b1 , \700_b0 , \701_b1 , \701_b0 , 
		\702_b1 , \702_b0 , \703_b1 , \703_b0 , \704_b1 , \704_b0 , \705_b1 , \705_b0 , \706_b1 , \706_b0 , 
		\707_b1 , \707_b0 , \708_b1 , \708_b0 , \709_b1 , \709_b0 , \710_b1 , \710_b0 , \711_b1 , \711_b0 , 
		\712_b1 , \712_b0 , \713_b1 , \713_b0 , \714_b1 , \714_b0 , \715_b1 , \715_b0 , \716_b1 , \716_b0 , 
		\717_b1 , \717_b0 , \718_b1 , \718_b0 , \719_b1 , \719_b0 , \720_b1 , \720_b0 , \721_b1 , \721_b0 , 
		\722_b1 , \722_b0 , \723_b1 , \723_b0 , \724_b1 , \724_b0 , \725_b1 , \725_b0 , \726_b1 , \726_b0 , 
		\727_b1 , \727_b0 , \728_b1 , \728_b0 , \729_b1 , \729_b0 , \730_b1 , \730_b0 , \731_b1 , \731_b0 , 
		\732_b1 , \732_b0 , \733_b1 , \733_b0 , \734_b1 , \734_b0 , \735_b1 , \735_b0 , \736_b1 , \736_b0 , 
		\737_b1 , \737_b0 , \738_b1 , \738_b0 , \739_b1 , \739_b0 , \740_b1 , \740_b0 , \741_b1 , \741_b0 , 
		\742_b1 , \742_b0 , \743_b1 , \743_b0 , \744_b1 , \744_b0 , \745_b1 , \745_b0 , \746_b1 , \746_b0 , 
		\747_b1 , \747_b0 , \748_b1 , \748_b0 , \749_b1 , \749_b0 , \750_b1 , \750_b0 , \751_b1 , \751_b0 , 
		\752_b1 , \752_b0 , \753_b1 , \753_b0 , \754_b1 , \754_b0 , \755_b1 , \755_b0 , \756_b1 , \756_b0 , 
		\757_b1 , \757_b0 , \758_b1 , \758_b0 , \759_b1 , \759_b0 , \760_b1 , \760_b0 , \761_B[14]_b1 , \761_B[14]_b0 , 
		\762_b1 , \762_b0 , \763_b1 , \763_b0 , \764_Z[14]_b1 , \764_Z[14]_b0 , \765_A[15]_b1 , \765_A[15]_b0 , \766_b1 , \766_b0 , 
		\767_b1 , \767_b0 , \768_b1 , \768_b0 , \769_b1 , \769_b0 , \770_b1 , \770_b0 , \771_b1 , \771_b0 , 
		\772_b1 , \772_b0 , \773_b1 , \773_b0 , \774_b1 , \774_b0 , \775_b1 , \775_b0 , \776_b1 , \776_b0 , 
		\777_b1 , \777_b0 , \778_b1 , \778_b0 , \779_b1 , \779_b0 , \780_b1 , \780_b0 , \781_b1 , \781_b0 , 
		\782_b1 , \782_b0 , \783_b1 , \783_b0 , \784_b1 , \784_b0 , \785_b1 , \785_b0 , \786_b1 , \786_b0 , 
		\787_b1 , \787_b0 , \788_b1 , \788_b0 , \789_b1 , \789_b0 , \790_b1 , \790_b0 , \791_b1 , \791_b0 , 
		\792_b1 , \792_b0 , \793_b1 , \793_b0 , \794_b1 , \794_b0 , \795_b1 , \795_b0 , \796_b1 , \796_b0 , 
		\797_b1 , \797_b0 , \798_b1 , \798_b0 , \799_b1 , \799_b0 , \800_b1 , \800_b0 , \801_b1 , \801_b0 , 
		\802_b1 , \802_b0 , \803_b1 , \803_b0 , \804_b1 , \804_b0 , \805_b1 , \805_b0 , \806_b1 , \806_b0 , 
		\807_b1 , \807_b0 , \808_b1 , \808_b0 , \809_b1 , \809_b0 , \810_b1 , \810_b0 , \811_b1 , \811_b0 , 
		\812_b1 , \812_b0 , \813_b1 , \813_b0 , \814_b1 , \814_b0 , \815_b1 , \815_b0 , \816_b1 , \816_b0 , 
		\817_b1 , \817_b0 , \818_b1 , \818_b0 , \819_b1 , \819_b0 , \820_b1 , \820_b0 , \821_b1 , \821_b0 , 
		\822_b1 , \822_b0 , \823_b1 , \823_b0 , \824_b1 , \824_b0 , \825_b1 , \825_b0 , \826_b1 , \826_b0 , 
		\827_b1 , \827_b0 , \828_b1 , \828_b0 , \829_b1 , \829_b0 , \830_b1 , \830_b0 , \831_b1 , \831_b0 , 
		\832_b1 , \832_b0 , \833_b1 , \833_b0 , \834_b1 , \834_b0 , \835_b1 , \835_b0 , \836_b1 , \836_b0 , 
		\837_b1 , \837_b0 , \838_b1 , \838_b0 , \839_b1 , \839_b0 , \840_b1 , \840_b0 , \841_b1 , \841_b0 , 
		\842_b1 , \842_b0 , \843_b1 , \843_b0 , \844_b1 , \844_b0 , \845_b1 , \845_b0 , \846_b1 , \846_b0 , 
		\847_b1 , \847_b0 , \848_b1 , \848_b0 , \849_B[15]_b1 , \849_B[15]_b0 , \850_b1 , \850_b0 , \851_b1 , \851_b0 , 
		\852_Z[15]_b1 , \852_Z[15]_b0 , \853_b1 , \853_b0 , \854_b1 , \854_b0 , \855_b1 , \855_b0 , \856_b1 , \856_b0 , 
		\857_b1 , \857_b0 , \858_b1 , \858_b0 , \859_b1 , \859_b0 , \860_b1 , \860_b0 , \861_b1 , \861_b0 , 
		\862_b1 , \862_b0 , \863_b1 , \863_b0 , \864_b1 , \864_b0 , \865_b1 , \865_b0 , \866_b1 , \866_b0 , 
		\867_b1 , \867_b0 , \868_b1 , \868_b0 , \869_b1 , \869_b0 , \870_b1 , \870_b0 , \871_b1 , \871_b0 , 
		\872_b1 , \872_b0 , \873_b1 , \873_b0 , \874_b1 , \874_b0 , \875_b1 , \875_b0 , \876_b1 , \876_b0 , 
		\877_b1 , \877_b0 , \878_b1 , \878_b0 , \879_b1 , \879_b0 , \880_b1 , \880_b0 , \881_b1 , \881_b0 , 
		\882_b1 , \882_b0 , \883_b1 , \883_b0 , \884_b1 , \884_b0 , \885_b1 , \885_b0 , \886_A[0]_b1 , \886_A[0]_b0 , 
		\887_B[0]_b1 , \887_B[0]_b0 , \888_b1 , \888_b0 , \889_Z[0]_b1 , \889_Z[0]_b0 , \890_b1 , \890_b0 , \891_A[0]_b1 , \891_A[0]_b0 , 
		\892_B[0]_b1 , \892_B[0]_b0 , \893_b1 , \893_b0 , \894_Z[0]_b1 , \894_Z[0]_b0 , \895_b1 , \895_b0 , \896_A[0]_b1 , \896_A[0]_b0 , 
		\897_B[0]_b1 , \897_B[0]_b0 , \898_b1 , \898_b0 , \899_SUM[0]_b1 , \899_SUM[0]_b0 , \900_b1 , \900_b0 , \901_A[0]_b1 , \901_A[0]_b0 , 
		\902_B[0]_b1 , \902_B[0]_b0 , \903_b1 , \903_b0 , \904_SUM[0]_b1 , \904_SUM[0]_b0 , \905_b1 , \905_b0 , \906_b1 , \906_b0 , 
		\907_b1 , \907_b0 , \908_b1 , \908_b0 , \909_b1 , \909_b0 , \910_b1 , \910_b0 , \911_b1 , \911_b0 , 
		\912_b1 , \912_b0 , \913_b1 , \913_b0 , \914_b1 , \914_b0 , \915_b1 , \915_b0 , \916_b1 , \916_b0 , 
		\917_b1 , \917_b0 , \918_b1 , \918_b0 , \919_b1 , \919_b0 , \920_A[1]_b1 , \920_A[1]_b0 , \921_b1 , \921_b0 , 
		\922_B[1]_b1 , \922_B[1]_b0 , \923_b1 , \923_b0 , \924_b1 , \924_b0 , \925_Z[1]_b1 , \925_Z[1]_b0 , \926_b1 , \926_b0 , 
		\927_A[1]_b1 , \927_A[1]_b0 , \928_b1 , \928_b0 , \929_B[1]_b1 , \929_B[1]_b0 , \930_b1 , \930_b0 , \931_b1 , \931_b0 , 
		\932_Z[1]_b1 , \932_Z[1]_b0 , \933_b1 , \933_b0 , \934_A[1]_b1 , \934_A[1]_b0 , \935_B[1]_b1 , \935_B[1]_b0 , \936_b1 , \936_b0 , 
		\937_b1 , \937_b0 , \938_b1 , \938_b0 , \939_SUM[1]_b1 , \939_SUM[1]_b0 , \940_b1 , \940_b0 , \941_A[1]_b1 , \941_A[1]_b0 , 
		\942_B[1]_b1 , \942_B[1]_b0 , \943_b1 , \943_b0 , \944_b1 , \944_b0 , \945_b1 , \945_b0 , \946_SUM[1]_b1 , \946_SUM[1]_b0 , 
		\947_b1 , \947_b0 , \948_b1 , \948_b0 , \949_b1 , \949_b0 , \950_b1 , \950_b0 , \951_b1 , \951_b0 , 
		\952_b1 , \952_b0 , \953_b1 , \953_b0 , \954_b1 , \954_b0 , \955_b1 , \955_b0 , \956_b1 , \956_b0 , 
		\957_b1 , \957_b0 , \958_b1 , \958_b0 , \959_b1 , \959_b0 , \960_b1 , \960_b0 , \961_b1 , \961_b0 , 
		\962_A[2]_b1 , \962_A[2]_b0 , \963_b1 , \963_b0 , \964_b1 , \964_b0 , \965_b1 , \965_b0 , \966_b1 , \966_b0 , 
		\967_b1 , \967_b0 , \968_B[2]_b1 , \968_B[2]_b0 , \969_b1 , \969_b0 , \970_b1 , \970_b0 , \971_Z[2]_b1 , \971_Z[2]_b0 , 
		\972_b1 , \972_b0 , \973_A[2]_b1 , \973_A[2]_b0 , \974_b1 , \974_b0 , \975_b1 , \975_b0 , \976_b1 , \976_b0 , 
		\977_b1 , \977_b0 , \978_b1 , \978_b0 , \979_B[2]_b1 , \979_B[2]_b0 , \980_b1 , \980_b0 , \981_b1 , \981_b0 , 
		\982_Z[2]_b1 , \982_Z[2]_b0 , \983_b1 , \983_b0 , \984_A[2]_b1 , \984_A[2]_b0 , \985_B[2]_b1 , \985_B[2]_b0 , \986_b1 , \986_b0 , 
		\987_b1 , \987_b0 , \988_b1 , \988_b0 , \989_b1 , \989_b0 , \990_b1 , \990_b0 , \991_b1 , \991_b0 , 
		\992_SUM[2]_b1 , \992_SUM[2]_b0 , \993_b1 , \993_b0 , \994_A[2]_b1 , \994_A[2]_b0 , \995_B[2]_b1 , \995_B[2]_b0 , \996_b1 , \996_b0 , 
		\997_b1 , \997_b0 , \998_b1 , \998_b0 , \999_b1 , \999_b0 , \1000_b1 , \1000_b0 , \1001_b1 , \1001_b0 , 
		\1002_SUM[2]_b1 , \1002_SUM[2]_b0 , \1003_b1 , \1003_b0 , \1004_b1 , \1004_b0 , \1005_b1 , \1005_b0 , \1006_b1 , \1006_b0 , 
		\1007_b1 , \1007_b0 , \1008_b1 , \1008_b0 , \1009_b1 , \1009_b0 , \1010_b1 , \1010_b0 , \1011_b1 , \1011_b0 , 
		\1012_b1 , \1012_b0 , \1013_b1 , \1013_b0 , \1014_b1 , \1014_b0 , \1015_b1 , \1015_b0 , \1016_b1 , \1016_b0 , 
		\1017_b1 , \1017_b0 , \1018_A[3]_b1 , \1018_A[3]_b0 , \1019_b1 , \1019_b0 , \1020_b1 , \1020_b0 , \1021_b1 , \1021_b0 , 
		\1022_b1 , \1022_b0 , \1023_b1 , \1023_b0 , \1024_b1 , \1024_b0 , \1025_b1 , \1025_b0 , \1026_b1 , \1026_b0 , 
		\1027_b1 , \1027_b0 , \1028_b1 , \1028_b0 , \1029_b1 , \1029_b0 , \1030_B[3]_b1 , \1030_B[3]_b0 , \1031_b1 , \1031_b0 , 
		\1032_b1 , \1032_b0 , \1033_Z[3]_b1 , \1033_Z[3]_b0 , \1034_b1 , \1034_b0 , \1035_A[3]_b1 , \1035_A[3]_b0 , \1036_b1 , \1036_b0 , 
		\1037_b1 , \1037_b0 , \1038_b1 , \1038_b0 , \1039_b1 , \1039_b0 , \1040_b1 , \1040_b0 , \1041_b1 , \1041_b0 , 
		\1042_b1 , \1042_b0 , \1043_b1 , \1043_b0 , \1044_b1 , \1044_b0 , \1045_b1 , \1045_b0 , \1046_b1 , \1046_b0 , 
		\1047_B[3]_b1 , \1047_B[3]_b0 , \1048_b1 , \1048_b0 , \1049_b1 , \1049_b0 , \1050_Z[3]_b1 , \1050_Z[3]_b0 , \1051_b1 , \1051_b0 , 
		\1052_A[3]_b1 , \1052_A[3]_b0 , \1053_B[3]_b1 , \1053_B[3]_b0 , \1054_b1 , \1054_b0 , \1055_b1 , \1055_b0 , \1056_b1 , \1056_b0 , 
		\1057_b1 , \1057_b0 , \1058_b1 , \1058_b0 , \1059_b1 , \1059_b0 , \1060_SUM[3]_b1 , \1060_SUM[3]_b0 , \1061_b1 , \1061_b0 , 
		\1062_A[3]_b1 , \1062_A[3]_b0 , \1063_B[3]_b1 , \1063_B[3]_b0 , \1064_b1 , \1064_b0 , \1065_b1 , \1065_b0 , \1066_b1 , \1066_b0 , 
		\1067_b1 , \1067_b0 , \1068_b1 , \1068_b0 , \1069_b1 , \1069_b0 , \1070_SUM[3]_b1 , \1070_SUM[3]_b0 , \1071_b1 , \1071_b0 , 
		\1072_b1 , \1072_b0 , \1073_b1 , \1073_b0 , \1074_b1 , \1074_b0 , \1075_b1 , \1075_b0 , \1076_b1 , \1076_b0 , 
		\1077_b1 , \1077_b0 , \1078_b1 , \1078_b0 , \1079_b1 , \1079_b0 , \1080_b1 , \1080_b0 , \1081_b1 , \1081_b0 , 
		\1082_b1 , \1082_b0 , \1083_b1 , \1083_b0 , \1084_b1 , \1084_b0 , \1085_b1 , \1085_b0 , \1086_A[4]_b1 , \1086_A[4]_b0 , 
		\1087_b1 , \1087_b0 , \1088_b1 , \1088_b0 , \1089_b1 , \1089_b0 , \1090_b1 , \1090_b0 , \1091_b1 , \1091_b0 , 
		\1092_b1 , \1092_b0 , \1093_b1 , \1093_b0 , \1094_b1 , \1094_b0 , \1095_b1 , \1095_b0 , \1096_b1 , \1096_b0 , 
		\1097_b1 , \1097_b0 , \1098_b1 , \1098_b0 , \1099_b1 , \1099_b0 , \1100_b1 , \1100_b0 , \1101_b1 , \1101_b0 , 
		\1102_b1 , \1102_b0 , \1103_b1 , \1103_b0 , \1104_B[4]_b1 , \1104_B[4]_b0 , \1105_b1 , \1105_b0 , \1106_b1 , \1106_b0 , 
		\1107_Z[4]_b1 , \1107_Z[4]_b0 , \1108_b1 , \1108_b0 , \1109_A[4]_b1 , \1109_A[4]_b0 , \1110_b1 , \1110_b0 , \1111_b1 , \1111_b0 , 
		\1112_b1 , \1112_b0 , \1113_b1 , \1113_b0 , \1114_b1 , \1114_b0 , \1115_b1 , \1115_b0 , \1116_b1 , \1116_b0 , 
		\1117_b1 , \1117_b0 , \1118_b1 , \1118_b0 , \1119_b1 , \1119_b0 , \1120_b1 , \1120_b0 , \1121_b1 , \1121_b0 , 
		\1122_b1 , \1122_b0 , \1123_b1 , \1123_b0 , \1124_b1 , \1124_b0 , \1125_b1 , \1125_b0 , \1126_b1 , \1126_b0 , 
		\1127_B[4]_b1 , \1127_B[4]_b0 , \1128_b1 , \1128_b0 , \1129_b1 , \1129_b0 , \1130_Z[4]_b1 , \1130_Z[4]_b0 , \1131_b1 , \1131_b0 , 
		\1132_A[4]_b1 , \1132_A[4]_b0 , \1133_B[4]_b1 , \1133_B[4]_b0 , \1134_b1 , \1134_b0 , \1135_b1 , \1135_b0 , \1136_b1 , \1136_b0 , 
		\1137_b1 , \1137_b0 , \1138_b1 , \1138_b0 , \1139_b1 , \1139_b0 , \1140_SUM[4]_b1 , \1140_SUM[4]_b0 , \1141_b1 , \1141_b0 , 
		\1142_A[4]_b1 , \1142_A[4]_b0 , \1143_B[4]_b1 , \1143_B[4]_b0 , \1144_b1 , \1144_b0 , \1145_b1 , \1145_b0 , \1146_b1 , \1146_b0 , 
		\1147_b1 , \1147_b0 , \1148_b1 , \1148_b0 , \1149_b1 , \1149_b0 , \1150_SUM[4]_b1 , \1150_SUM[4]_b0 , \1151_b1 , \1151_b0 , 
		\1152_b1 , \1152_b0 , \1153_b1 , \1153_b0 , \1154_b1 , \1154_b0 , \1155_b1 , \1155_b0 , \1156_b1 , \1156_b0 , 
		\1157_b1 , \1157_b0 , \1158_b1 , \1158_b0 , \1159_b1 , \1159_b0 , \1160_b1 , \1160_b0 , \1161_b1 , \1161_b0 , 
		\1162_b1 , \1162_b0 , \1163_b1 , \1163_b0 , \1164_b1 , \1164_b0 , \1165_b1 , \1165_b0 , \1166_A[5]_b1 , \1166_A[5]_b0 , 
		\1167_b1 , \1167_b0 , \1168_b1 , \1168_b0 , \1169_b1 , \1169_b0 , \1170_b1 , \1170_b0 , \1171_b1 , \1171_b0 , 
		\1172_b1 , \1172_b0 , \1173_b1 , \1173_b0 , \1174_b1 , \1174_b0 , \1175_b1 , \1175_b0 , \1176_b1 , \1176_b0 , 
		\1177_b1 , \1177_b0 , \1178_b1 , \1178_b0 , \1179_b1 , \1179_b0 , \1180_b1 , \1180_b0 , \1181_b1 , \1181_b0 , 
		\1182_b1 , \1182_b0 , \1183_b1 , \1183_b0 , \1184_b1 , \1184_b0 , \1185_b1 , \1185_b0 , \1186_b1 , \1186_b0 , 
		\1187_b1 , \1187_b0 , \1188_b1 , \1188_b0 , \1189_b1 , \1189_b0 , \1190_B[5]_b1 , \1190_B[5]_b0 , \1191_b1 , \1191_b0 , 
		\1192_b1 , \1192_b0 , \1193_Z[5]_b1 , \1193_Z[5]_b0 , \1194_b1 , \1194_b0 , \1195_A[5]_b1 , \1195_A[5]_b0 , \1196_b1 , \1196_b0 , 
		\1197_b1 , \1197_b0 , \1198_b1 , \1198_b0 , \1199_b1 , \1199_b0 , \1200_b1 , \1200_b0 , \1201_b1 , \1201_b0 , 
		\1202_b1 , \1202_b0 , \1203_b1 , \1203_b0 , \1204_b1 , \1204_b0 , \1205_b1 , \1205_b0 , \1206_b1 , \1206_b0 , 
		\1207_b1 , \1207_b0 , \1208_b1 , \1208_b0 , \1209_b1 , \1209_b0 , \1210_b1 , \1210_b0 , \1211_b1 , \1211_b0 , 
		\1212_b1 , \1212_b0 , \1213_b1 , \1213_b0 , \1214_b1 , \1214_b0 , \1215_b1 , \1215_b0 , \1216_b1 , \1216_b0 , 
		\1217_b1 , \1217_b0 , \1218_b1 , \1218_b0 , \1219_B[5]_b1 , \1219_B[5]_b0 , \1220_b1 , \1220_b0 , \1221_b1 , \1221_b0 , 
		\1222_Z[5]_b1 , \1222_Z[5]_b0 , \1223_b1 , \1223_b0 , \1224_A[5]_b1 , \1224_A[5]_b0 , \1225_B[5]_b1 , \1225_B[5]_b0 , \1226_b1 , \1226_b0 , 
		\1227_b1 , \1227_b0 , \1228_b1 , \1228_b0 , \1229_b1 , \1229_b0 , \1230_b1 , \1230_b0 , \1231_b1 , \1231_b0 , 
		\1232_SUM[5]_b1 , \1232_SUM[5]_b0 , \1233_b1 , \1233_b0 , \1234_A[5]_b1 , \1234_A[5]_b0 , \1235_B[5]_b1 , \1235_B[5]_b0 , \1236_b1 , \1236_b0 , 
		\1237_b1 , \1237_b0 , \1238_b1 , \1238_b0 , \1239_b1 , \1239_b0 , \1240_b1 , \1240_b0 , \1241_b1 , \1241_b0 , 
		\1242_SUM[5]_b1 , \1242_SUM[5]_b0 , \1243_b1 , \1243_b0 , \1244_b1 , \1244_b0 , \1245_b1 , \1245_b0 , \1246_b1 , \1246_b0 , 
		\1247_b1 , \1247_b0 , \1248_b1 , \1248_b0 , \1249_b1 , \1249_b0 , \1250_b1 , \1250_b0 , \1251_b1 , \1251_b0 , 
		\1252_b1 , \1252_b0 , \1253_b1 , \1253_b0 , \1254_b1 , \1254_b0 , \1255_b1 , \1255_b0 , \1256_b1 , \1256_b0 , 
		\1257_b1 , \1257_b0 , \1258_A[6]_b1 , \1258_A[6]_b0 , \1259_b1 , \1259_b0 , \1260_b1 , \1260_b0 , \1261_b1 , \1261_b0 , 
		\1262_b1 , \1262_b0 , \1263_b1 , \1263_b0 , \1264_b1 , \1264_b0 , \1265_b1 , \1265_b0 , \1266_b1 , \1266_b0 , 
		\1267_b1 , \1267_b0 , \1268_b1 , \1268_b0 , \1269_b1 , \1269_b0 , \1270_b1 , \1270_b0 , \1271_b1 , \1271_b0 , 
		\1272_b1 , \1272_b0 , \1273_b1 , \1273_b0 , \1274_b1 , \1274_b0 , \1275_b1 , \1275_b0 , \1276_b1 , \1276_b0 , 
		\1277_b1 , \1277_b0 , \1278_b1 , \1278_b0 , \1279_b1 , \1279_b0 , \1280_b1 , \1280_b0 , \1281_b1 , \1281_b0 , 
		\1282_b1 , \1282_b0 , \1283_b1 , \1283_b0 , \1284_b1 , \1284_b0 , \1285_b1 , \1285_b0 , \1286_b1 , \1286_b0 , 
		\1287_b1 , \1287_b0 , \1288_B[6]_b1 , \1288_B[6]_b0 , \1289_b1 , \1289_b0 , \1290_b1 , \1290_b0 , \1291_Z[6]_b1 , \1291_Z[6]_b0 , 
		\1292_b1 , \1292_b0 , \1293_A[6]_b1 , \1293_A[6]_b0 , \1294_b1 , \1294_b0 , \1295_b1 , \1295_b0 , \1296_b1 , \1296_b0 , 
		\1297_b1 , \1297_b0 , \1298_b1 , \1298_b0 , \1299_b1 , \1299_b0 , \1300_b1 , \1300_b0 , \1301_b1 , \1301_b0 , 
		\1302_b1 , \1302_b0 , \1303_b1 , \1303_b0 , \1304_b1 , \1304_b0 , \1305_b1 , \1305_b0 , \1306_b1 , \1306_b0 , 
		\1307_b1 , \1307_b0 , \1308_b1 , \1308_b0 , \1309_b1 , \1309_b0 , \1310_b1 , \1310_b0 , \1311_b1 , \1311_b0 , 
		\1312_b1 , \1312_b0 , \1313_b1 , \1313_b0 , \1314_b1 , \1314_b0 , \1315_b1 , \1315_b0 , \1316_b1 , \1316_b0 , 
		\1317_b1 , \1317_b0 , \1318_b1 , \1318_b0 , \1319_b1 , \1319_b0 , \1320_b1 , \1320_b0 , \1321_b1 , \1321_b0 , 
		\1322_b1 , \1322_b0 , \1323_B[6]_b1 , \1323_B[6]_b0 , \1324_b1 , \1324_b0 , \1325_b1 , \1325_b0 , \1326_Z[6]_b1 , \1326_Z[6]_b0 , 
		\1327_b1 , \1327_b0 , \1328_A[6]_b1 , \1328_A[6]_b0 , \1329_B[6]_b1 , \1329_B[6]_b0 , \1330_b1 , \1330_b0 , \1331_b1 , \1331_b0 , 
		\1332_b1 , \1332_b0 , \1333_b1 , \1333_b0 , \1334_b1 , \1334_b0 , \1335_b1 , \1335_b0 , \1336_SUM[6]_b1 , \1336_SUM[6]_b0 , 
		\1337_b1 , \1337_b0 , \1338_A[6]_b1 , \1338_A[6]_b0 , \1339_B[6]_b1 , \1339_B[6]_b0 , \1340_b1 , \1340_b0 , \1341_b1 , \1341_b0 , 
		\1342_b1 , \1342_b0 , \1343_b1 , \1343_b0 , \1344_b1 , \1344_b0 , \1345_b1 , \1345_b0 , \1346_SUM[6]_b1 , \1346_SUM[6]_b0 , 
		\1347_b1 , \1347_b0 , \1348_b1 , \1348_b0 , \1349_b1 , \1349_b0 , \1350_b1 , \1350_b0 , \1351_b1 , \1351_b0 , 
		\1352_b1 , \1352_b0 , \1353_b1 , \1353_b0 , \1354_b1 , \1354_b0 , \1355_b1 , \1355_b0 , \1356_b1 , \1356_b0 , 
		\1357_b1 , \1357_b0 , \1358_b1 , \1358_b0 , \1359_b1 , \1359_b0 , \1360_b1 , \1360_b0 , \1361_b1 , \1361_b0 , 
		\1362_A[7]_b1 , \1362_A[7]_b0 , \1363_b1 , \1363_b0 , \1364_b1 , \1364_b0 , \1365_b1 , \1365_b0 , \1366_b1 , \1366_b0 , 
		\1367_b1 , \1367_b0 , \1368_b1 , \1368_b0 , \1369_b1 , \1369_b0 , \1370_b1 , \1370_b0 , \1371_b1 , \1371_b0 , 
		\1372_b1 , \1372_b0 , \1373_b1 , \1373_b0 , \1374_b1 , \1374_b0 , \1375_b1 , \1375_b0 , \1376_b1 , \1376_b0 , 
		\1377_b1 , \1377_b0 , \1378_b1 , \1378_b0 , \1379_b1 , \1379_b0 , \1380_b1 , \1380_b0 , \1381_b1 , \1381_b0 , 
		\1382_b1 , \1382_b0 , \1383_b1 , \1383_b0 , \1384_b1 , \1384_b0 , \1385_b1 , \1385_b0 , \1386_b1 , \1386_b0 , 
		\1387_b1 , \1387_b0 , \1388_b1 , \1388_b0 , \1389_b1 , \1389_b0 , \1390_b1 , \1390_b0 , \1391_b1 , \1391_b0 , 
		\1392_b1 , \1392_b0 , \1393_b1 , \1393_b0 , \1394_b1 , \1394_b0 , \1395_b1 , \1395_b0 , \1396_b1 , \1396_b0 , 
		\1397_b1 , \1397_b0 , \1398_B[7]_b1 , \1398_B[7]_b0 , \1399_b1 , \1399_b0 , \1400_b1 , \1400_b0 , \1401_Z[7]_b1 , \1401_Z[7]_b0 , 
		\1402_b1 , \1402_b0 , \1403_A[7]_b1 , \1403_A[7]_b0 , \1404_b1 , \1404_b0 , \1405_b1 , \1405_b0 , \1406_b1 , \1406_b0 , 
		\1407_b1 , \1407_b0 , \1408_b1 , \1408_b0 , \1409_b1 , \1409_b0 , \1410_b1 , \1410_b0 , \1411_b1 , \1411_b0 , 
		\1412_b1 , \1412_b0 , \1413_b1 , \1413_b0 , \1414_b1 , \1414_b0 , \1415_b1 , \1415_b0 , \1416_b1 , \1416_b0 , 
		\1417_b1 , \1417_b0 , \1418_b1 , \1418_b0 , \1419_b1 , \1419_b0 , \1420_b1 , \1420_b0 , \1421_b1 , \1421_b0 , 
		\1422_b1 , \1422_b0 , \1423_b1 , \1423_b0 , \1424_b1 , \1424_b0 , \1425_b1 , \1425_b0 , \1426_b1 , \1426_b0 , 
		\1427_b1 , \1427_b0 , \1428_b1 , \1428_b0 , \1429_b1 , \1429_b0 , \1430_b1 , \1430_b0 , \1431_b1 , \1431_b0 , 
		\1432_b1 , \1432_b0 , \1433_b1 , \1433_b0 , \1434_b1 , \1434_b0 , \1435_b1 , \1435_b0 , \1436_b1 , \1436_b0 , 
		\1437_b1 , \1437_b0 , \1438_b1 , \1438_b0 , \1439_B[7]_b1 , \1439_B[7]_b0 , \1440_b1 , \1440_b0 , \1441_b1 , \1441_b0 , 
		\1442_Z[7]_b1 , \1442_Z[7]_b0 , \1443_b1 , \1443_b0 , \1444_A[7]_b1 , \1444_A[7]_b0 , \1445_B[7]_b1 , \1445_B[7]_b0 , \1446_b1 , \1446_b0 , 
		\1447_b1 , \1447_b0 , \1448_b1 , \1448_b0 , \1449_b1 , \1449_b0 , \1450_b1 , \1450_b0 , \1451_b1 , \1451_b0 , 
		\1452_SUM[7]_b1 , \1452_SUM[7]_b0 , \1453_b1 , \1453_b0 , \1454_A[7]_b1 , \1454_A[7]_b0 , \1455_B[7]_b1 , \1455_B[7]_b0 , \1456_b1 , \1456_b0 , 
		\1457_b1 , \1457_b0 , \1458_b1 , \1458_b0 , \1459_b1 , \1459_b0 , \1460_b1 , \1460_b0 , \1461_b1 , \1461_b0 , 
		\1462_SUM[7]_b1 , \1462_SUM[7]_b0 , \1463_b1 , \1463_b0 , \1464_b1 , \1464_b0 , \1465_b1 , \1465_b0 , \1466_b1 , \1466_b0 , 
		\1467_b1 , \1467_b0 , \1468_b1 , \1468_b0 , \1469_b1 , \1469_b0 , \1470_b1 , \1470_b0 , \1471_b1 , \1471_b0 , 
		\1472_b1 , \1472_b0 , \1473_b1 , \1473_b0 , \1474_b1 , \1474_b0 , \1475_b1 , \1475_b0 , \1476_b1 , \1476_b0 , 
		\1477_b1 , \1477_b0 , \1478_A[8]_b1 , \1478_A[8]_b0 , \1479_b1 , \1479_b0 , \1480_b1 , \1480_b0 , \1481_b1 , \1481_b0 , 
		\1482_b1 , \1482_b0 , \1483_b1 , \1483_b0 , \1484_b1 , \1484_b0 , \1485_b1 , \1485_b0 , \1486_b1 , \1486_b0 , 
		\1487_b1 , \1487_b0 , \1488_b1 , \1488_b0 , \1489_b1 , \1489_b0 , \1490_b1 , \1490_b0 , \1491_b1 , \1491_b0 , 
		\1492_b1 , \1492_b0 , \1493_b1 , \1493_b0 , \1494_b1 , \1494_b0 , \1495_b1 , \1495_b0 , \1496_b1 , \1496_b0 , 
		\1497_b1 , \1497_b0 , \1498_b1 , \1498_b0 , \1499_b1 , \1499_b0 , \1500_b1 , \1500_b0 , \1501_b1 , \1501_b0 , 
		\1502_b1 , \1502_b0 , \1503_b1 , \1503_b0 , \1504_b1 , \1504_b0 , \1505_b1 , \1505_b0 , \1506_b1 , \1506_b0 , 
		\1507_b1 , \1507_b0 , \1508_b1 , \1508_b0 , \1509_b1 , \1509_b0 , \1510_b1 , \1510_b0 , \1511_b1 , \1511_b0 , 
		\1512_b1 , \1512_b0 , \1513_b1 , \1513_b0 , \1514_b1 , \1514_b0 , \1515_b1 , \1515_b0 , \1516_b1 , \1516_b0 , 
		\1517_b1 , \1517_b0 , \1518_b1 , \1518_b0 , \1519_b1 , \1519_b0 , \1520_B[8]_b1 , \1520_B[8]_b0 , \1521_b1 , \1521_b0 , 
		\1522_b1 , \1522_b0 , \1523_Z[8]_b1 , \1523_Z[8]_b0 , \1524_b1 , \1524_b0 , \1525_A[8]_b1 , \1525_A[8]_b0 , \1526_b1 , \1526_b0 , 
		\1527_b1 , \1527_b0 , \1528_b1 , \1528_b0 , \1529_b1 , \1529_b0 , \1530_b1 , \1530_b0 , \1531_b1 , \1531_b0 , 
		\1532_b1 , \1532_b0 , \1533_b1 , \1533_b0 , \1534_b1 , \1534_b0 , \1535_b1 , \1535_b0 , \1536_b1 , \1536_b0 , 
		\1537_b1 , \1537_b0 , \1538_b1 , \1538_b0 , \1539_b1 , \1539_b0 , \1540_b1 , \1540_b0 , \1541_b1 , \1541_b0 , 
		\1542_b1 , \1542_b0 , \1543_b1 , \1543_b0 , \1544_b1 , \1544_b0 , \1545_b1 , \1545_b0 , \1546_b1 , \1546_b0 , 
		\1547_b1 , \1547_b0 , \1548_b1 , \1548_b0 , \1549_b1 , \1549_b0 , \1550_b1 , \1550_b0 , \1551_b1 , \1551_b0 , 
		\1552_b1 , \1552_b0 , \1553_b1 , \1553_b0 , \1554_b1 , \1554_b0 , \1555_b1 , \1555_b0 , \1556_b1 , \1556_b0 , 
		\1557_b1 , \1557_b0 , \1558_b1 , \1558_b0 , \1559_b1 , \1559_b0 , \1560_b1 , \1560_b0 , \1561_b1 , \1561_b0 , 
		\1562_b1 , \1562_b0 , \1563_b1 , \1563_b0 , \1564_b1 , \1564_b0 , \1565_b1 , \1565_b0 , \1566_b1 , \1566_b0 , 
		\1567_B[8]_b1 , \1567_B[8]_b0 , \1568_b1 , \1568_b0 , \1569_b1 , \1569_b0 , \1570_Z[8]_b1 , \1570_Z[8]_b0 , \1571_b1 , \1571_b0 , 
		\1572_A[8]_b1 , \1572_A[8]_b0 , \1573_B[8]_b1 , \1573_B[8]_b0 , \1574_b1 , \1574_b0 , \1575_b1 , \1575_b0 , \1576_b1 , \1576_b0 , 
		\1577_b1 , \1577_b0 , \1578_b1 , \1578_b0 , \1579_b1 , \1579_b0 , \1580_SUM[8]_b1 , \1580_SUM[8]_b0 , \1581_b1 , \1581_b0 , 
		\1582_A[8]_b1 , \1582_A[8]_b0 , \1583_B[8]_b1 , \1583_B[8]_b0 , \1584_b1 , \1584_b0 , \1585_b1 , \1585_b0 , \1586_b1 , \1586_b0 , 
		\1587_b1 , \1587_b0 , \1588_b1 , \1588_b0 , \1589_b1 , \1589_b0 , \1590_SUM[8]_b1 , \1590_SUM[8]_b0 , \1591_b1 , \1591_b0 , 
		\1592_b1 , \1592_b0 , \1593_b1 , \1593_b0 , \1594_b1 , \1594_b0 , \1595_b1 , \1595_b0 , \1596_b1 , \1596_b0 , 
		\1597_b1 , \1597_b0 , \1598_b1 , \1598_b0 , \1599_b1 , \1599_b0 , \1600_b1 , \1600_b0 , \1601_b1 , \1601_b0 , 
		\1602_b1 , \1602_b0 , \1603_b1 , \1603_b0 , \1604_b1 , \1604_b0 , \1605_b1 , \1605_b0 , \1606_A[9]_b1 , \1606_A[9]_b0 , 
		\1607_b1 , \1607_b0 , \1608_b1 , \1608_b0 , \1609_b1 , \1609_b0 , \1610_b1 , \1610_b0 , \1611_b1 , \1611_b0 , 
		\1612_b1 , \1612_b0 , \1613_b1 , \1613_b0 , \1614_b1 , \1614_b0 , \1615_b1 , \1615_b0 , \1616_b1 , \1616_b0 , 
		\1617_b1 , \1617_b0 , \1618_b1 , \1618_b0 , \1619_b1 , \1619_b0 , \1620_b1 , \1620_b0 , \1621_b1 , \1621_b0 , 
		\1622_b1 , \1622_b0 , \1623_b1 , \1623_b0 , \1624_b1 , \1624_b0 , \1625_b1 , \1625_b0 , \1626_b1 , \1626_b0 , 
		\1627_b1 , \1627_b0 , \1628_b1 , \1628_b0 , \1629_b1 , \1629_b0 , \1630_b1 , \1630_b0 , \1631_b1 , \1631_b0 , 
		\1632_b1 , \1632_b0 , \1633_b1 , \1633_b0 , \1634_b1 , \1634_b0 , \1635_b1 , \1635_b0 , \1636_b1 , \1636_b0 , 
		\1637_b1 , \1637_b0 , \1638_b1 , \1638_b0 , \1639_b1 , \1639_b0 , \1640_b1 , \1640_b0 , \1641_b1 , \1641_b0 , 
		\1642_b1 , \1642_b0 , \1643_b1 , \1643_b0 , \1644_b1 , \1644_b0 , \1645_b1 , \1645_b0 , \1646_b1 , \1646_b0 , 
		\1647_b1 , \1647_b0 , \1648_b1 , \1648_b0 , \1649_b1 , \1649_b0 , \1650_b1 , \1650_b0 , \1651_b1 , \1651_b0 , 
		\1652_b1 , \1652_b0 , \1653_b1 , \1653_b0 , \1654_B[9]_b1 , \1654_B[9]_b0 , \1655_b1 , \1655_b0 , \1656_b1 , \1656_b0 , 
		\1657_Z[9]_b1 , \1657_Z[9]_b0 , \1658_b1 , \1658_b0 , \1659_A[9]_b1 , \1659_A[9]_b0 , \1660_b1 , \1660_b0 , \1661_b1 , \1661_b0 , 
		\1662_b1 , \1662_b0 , \1663_b1 , \1663_b0 , \1664_b1 , \1664_b0 , \1665_b1 , \1665_b0 , \1666_b1 , \1666_b0 , 
		\1667_b1 , \1667_b0 , \1668_b1 , \1668_b0 , \1669_b1 , \1669_b0 , \1670_b1 , \1670_b0 , \1671_b1 , \1671_b0 , 
		\1672_b1 , \1672_b0 , \1673_b1 , \1673_b0 , \1674_b1 , \1674_b0 , \1675_b1 , \1675_b0 , \1676_b1 , \1676_b0 , 
		\1677_b1 , \1677_b0 , \1678_b1 , \1678_b0 , \1679_b1 , \1679_b0 , \1680_b1 , \1680_b0 , \1681_b1 , \1681_b0 , 
		\1682_b1 , \1682_b0 , \1683_b1 , \1683_b0 , \1684_b1 , \1684_b0 , \1685_b1 , \1685_b0 , \1686_b1 , \1686_b0 , 
		\1687_b1 , \1687_b0 , \1688_b1 , \1688_b0 , \1689_b1 , \1689_b0 , \1690_b1 , \1690_b0 , \1691_b1 , \1691_b0 , 
		\1692_b1 , \1692_b0 , \1693_b1 , \1693_b0 , \1694_b1 , \1694_b0 , \1695_b1 , \1695_b0 , \1696_b1 , \1696_b0 , 
		\1697_b1 , \1697_b0 , \1698_b1 , \1698_b0 , \1699_b1 , \1699_b0 , \1700_b1 , \1700_b0 , \1701_b1 , \1701_b0 , 
		\1702_b1 , \1702_b0 , \1703_b1 , \1703_b0 , \1704_b1 , \1704_b0 , \1705_b1 , \1705_b0 , \1706_b1 , \1706_b0 , 
		\1707_B[9]_b1 , \1707_B[9]_b0 , \1708_b1 , \1708_b0 , \1709_b1 , \1709_b0 , \1710_Z[9]_b1 , \1710_Z[9]_b0 , \1711_b1 , \1711_b0 , 
		\1712_A[9]_b1 , \1712_A[9]_b0 , \1713_B[9]_b1 , \1713_B[9]_b0 , \1714_b1 , \1714_b0 , \1715_b1 , \1715_b0 , \1716_b1 , \1716_b0 , 
		\1717_b1 , \1717_b0 , \1718_b1 , \1718_b0 , \1719_b1 , \1719_b0 , \1720_SUM[9]_b1 , \1720_SUM[9]_b0 , \1721_b1 , \1721_b0 , 
		\1722_A[9]_b1 , \1722_A[9]_b0 , \1723_B[9]_b1 , \1723_B[9]_b0 , \1724_b1 , \1724_b0 , \1725_b1 , \1725_b0 , \1726_b1 , \1726_b0 , 
		\1727_b1 , \1727_b0 , \1728_b1 , \1728_b0 , \1729_b1 , \1729_b0 , \1730_SUM[9]_b1 , \1730_SUM[9]_b0 , \1731_b1 , \1731_b0 , 
		\1732_b1 , \1732_b0 , \1733_b1 , \1733_b0 , \1734_b1 , \1734_b0 , \1735_b1 , \1735_b0 , \1736_b1 , \1736_b0 , 
		\1737_b1 , \1737_b0 , \1738_b1 , \1738_b0 , \1739_b1 , \1739_b0 , \1740_b1 , \1740_b0 , \1741_b1 , \1741_b0 , 
		\1742_b1 , \1742_b0 , \1743_b1 , \1743_b0 , \1744_b1 , \1744_b0 , \1745_b1 , \1745_b0 , \1746_A[10]_b1 , \1746_A[10]_b0 , 
		\1747_b1 , \1747_b0 , \1748_b1 , \1748_b0 , \1749_b1 , \1749_b0 , \1750_b1 , \1750_b0 , \1751_b1 , \1751_b0 , 
		\1752_b1 , \1752_b0 , \1753_b1 , \1753_b0 , \1754_b1 , \1754_b0 , \1755_b1 , \1755_b0 , \1756_b1 , \1756_b0 , 
		\1757_b1 , \1757_b0 , \1758_b1 , \1758_b0 , \1759_b1 , \1759_b0 , \1760_b1 , \1760_b0 , \1761_b1 , \1761_b0 , 
		\1762_b1 , \1762_b0 , \1763_b1 , \1763_b0 , \1764_b1 , \1764_b0 , \1765_b1 , \1765_b0 , \1766_b1 , \1766_b0 , 
		\1767_b1 , \1767_b0 , \1768_b1 , \1768_b0 , \1769_b1 , \1769_b0 , \1770_b1 , \1770_b0 , \1771_b1 , \1771_b0 , 
		\1772_b1 , \1772_b0 , \1773_b1 , \1773_b0 , \1774_b1 , \1774_b0 , \1775_b1 , \1775_b0 , \1776_b1 , \1776_b0 , 
		\1777_b1 , \1777_b0 , \1778_b1 , \1778_b0 , \1779_b1 , \1779_b0 , \1780_b1 , \1780_b0 , \1781_b1 , \1781_b0 , 
		\1782_b1 , \1782_b0 , \1783_b1 , \1783_b0 , \1784_b1 , \1784_b0 , \1785_b1 , \1785_b0 , \1786_b1 , \1786_b0 , 
		\1787_b1 , \1787_b0 , \1788_b1 , \1788_b0 , \1789_b1 , \1789_b0 , \1790_b1 , \1790_b0 , \1791_b1 , \1791_b0 , 
		\1792_b1 , \1792_b0 , \1793_b1 , \1793_b0 , \1794_b1 , \1794_b0 , \1795_b1 , \1795_b0 , \1796_b1 , \1796_b0 , 
		\1797_b1 , \1797_b0 , \1798_b1 , \1798_b0 , \1799_b1 , \1799_b0 , \1800_B[10]_b1 , \1800_B[10]_b0 , \1801_b1 , \1801_b0 , 
		\1802_b1 , \1802_b0 , \1803_Z[10]_b1 , \1803_Z[10]_b0 , \1804_b1 , \1804_b0 , \1805_A[10]_b1 , \1805_A[10]_b0 , \1806_b1 , \1806_b0 , 
		\1807_b1 , \1807_b0 , \1808_b1 , \1808_b0 , \1809_b1 , \1809_b0 , \1810_b1 , \1810_b0 , \1811_b1 , \1811_b0 , 
		\1812_b1 , \1812_b0 , \1813_b1 , \1813_b0 , \1814_b1 , \1814_b0 , \1815_b1 , \1815_b0 , \1816_b1 , \1816_b0 , 
		\1817_b1 , \1817_b0 , \1818_b1 , \1818_b0 , \1819_b1 , \1819_b0 , \1820_b1 , \1820_b0 , \1821_b1 , \1821_b0 , 
		\1822_b1 , \1822_b0 , \1823_b1 , \1823_b0 , \1824_b1 , \1824_b0 , \1825_b1 , \1825_b0 , \1826_b1 , \1826_b0 , 
		\1827_b1 , \1827_b0 , \1828_b1 , \1828_b0 , \1829_b1 , \1829_b0 , \1830_b1 , \1830_b0 , \1831_b1 , \1831_b0 , 
		\1832_b1 , \1832_b0 , \1833_b1 , \1833_b0 , \1834_b1 , \1834_b0 , \1835_b1 , \1835_b0 , \1836_b1 , \1836_b0 , 
		\1837_b1 , \1837_b0 , \1838_b1 , \1838_b0 , \1839_b1 , \1839_b0 , \1840_b1 , \1840_b0 , \1841_b1 , \1841_b0 , 
		\1842_b1 , \1842_b0 , \1843_b1 , \1843_b0 , \1844_b1 , \1844_b0 , \1845_b1 , \1845_b0 , \1846_b1 , \1846_b0 , 
		\1847_b1 , \1847_b0 , \1848_b1 , \1848_b0 , \1849_b1 , \1849_b0 , \1850_b1 , \1850_b0 , \1851_b1 , \1851_b0 , 
		\1852_b1 , \1852_b0 , \1853_b1 , \1853_b0 , \1854_b1 , \1854_b0 , \1855_b1 , \1855_b0 , \1856_b1 , \1856_b0 , 
		\1857_b1 , \1857_b0 , \1858_b1 , \1858_b0 , \1859_B[10]_b1 , \1859_B[10]_b0 , \1860_b1 , \1860_b0 , \1861_b1 , \1861_b0 , 
		\1862_Z[10]_b1 , \1862_Z[10]_b0 , \1863_b1 , \1863_b0 , \1864_A[10]_b1 , \1864_A[10]_b0 , \1865_B[10]_b1 , \1865_B[10]_b0 , \1866_b1 , \1866_b0 , 
		\1867_b1 , \1867_b0 , \1868_b1 , \1868_b0 , \1869_b1 , \1869_b0 , \1870_b1 , \1870_b0 , \1871_b1 , \1871_b0 , 
		\1872_SUM[10]_b1 , \1872_SUM[10]_b0 , \1873_b1 , \1873_b0 , \1874_A[10]_b1 , \1874_A[10]_b0 , \1875_B[10]_b1 , \1875_B[10]_b0 , \1876_b1 , \1876_b0 , 
		\1877_b1 , \1877_b0 , \1878_b1 , \1878_b0 , \1879_b1 , \1879_b0 , \1880_b1 , \1880_b0 , \1881_b1 , \1881_b0 , 
		\1882_SUM[10]_b1 , \1882_SUM[10]_b0 , \1883_b1 , \1883_b0 , \1884_b1 , \1884_b0 , \1885_b1 , \1885_b0 , \1886_b1 , \1886_b0 , 
		\1887_b1 , \1887_b0 , \1888_b1 , \1888_b0 , \1889_b1 , \1889_b0 , \1890_b1 , \1890_b0 , \1891_b1 , \1891_b0 , 
		\1892_b1 , \1892_b0 , \1893_b1 , \1893_b0 , \1894_b1 , \1894_b0 , \1895_b1 , \1895_b0 , \1896_b1 , \1896_b0 , 
		\1897_b1 , \1897_b0 , \1898_A[11]_b1 , \1898_A[11]_b0 , \1899_b1 , \1899_b0 , \1900_b1 , \1900_b0 , \1901_b1 , \1901_b0 , 
		\1902_b1 , \1902_b0 , \1903_b1 , \1903_b0 , \1904_b1 , \1904_b0 , \1905_b1 , \1905_b0 , \1906_b1 , \1906_b0 , 
		\1907_b1 , \1907_b0 , \1908_b1 , \1908_b0 , \1909_b1 , \1909_b0 , \1910_b1 , \1910_b0 , \1911_b1 , \1911_b0 , 
		\1912_b1 , \1912_b0 , \1913_b1 , \1913_b0 , \1914_b1 , \1914_b0 , \1915_b1 , \1915_b0 , \1916_b1 , \1916_b0 , 
		\1917_b1 , \1917_b0 , \1918_b1 , \1918_b0 , \1919_b1 , \1919_b0 , \1920_b1 , \1920_b0 , \1921_b1 , \1921_b0 , 
		\1922_b1 , \1922_b0 , \1923_b1 , \1923_b0 , \1924_b1 , \1924_b0 , \1925_b1 , \1925_b0 , \1926_b1 , \1926_b0 , 
		\1927_b1 , \1927_b0 , \1928_b1 , \1928_b0 , \1929_b1 , \1929_b0 , \1930_b1 , \1930_b0 , \1931_b1 , \1931_b0 , 
		\1932_b1 , \1932_b0 , \1933_b1 , \1933_b0 , \1934_b1 , \1934_b0 , \1935_b1 , \1935_b0 , \1936_b1 , \1936_b0 , 
		\1937_b1 , \1937_b0 , \1938_b1 , \1938_b0 , \1939_b1 , \1939_b0 , \1940_b1 , \1940_b0 , \1941_b1 , \1941_b0 , 
		\1942_b1 , \1942_b0 , \1943_b1 , \1943_b0 , \1944_b1 , \1944_b0 , \1945_b1 , \1945_b0 , \1946_b1 , \1946_b0 , 
		\1947_b1 , \1947_b0 , \1948_b1 , \1948_b0 , \1949_b1 , \1949_b0 , \1950_b1 , \1950_b0 , \1951_b1 , \1951_b0 , 
		\1952_b1 , \1952_b0 , \1953_b1 , \1953_b0 , \1954_b1 , \1954_b0 , \1955_b1 , \1955_b0 , \1956_b1 , \1956_b0 , 
		\1957_b1 , \1957_b0 , \1958_B[11]_b1 , \1958_B[11]_b0 , \1959_b1 , \1959_b0 , \1960_b1 , \1960_b0 , \1961_Z[11]_b1 , \1961_Z[11]_b0 , 
		\1962_b1 , \1962_b0 , \1963_A[11]_b1 , \1963_A[11]_b0 , \1964_b1 , \1964_b0 , \1965_b1 , \1965_b0 , \1966_b1 , \1966_b0 , 
		\1967_b1 , \1967_b0 , \1968_b1 , \1968_b0 , \1969_b1 , \1969_b0 , \1970_b1 , \1970_b0 , \1971_b1 , \1971_b0 , 
		\1972_b1 , \1972_b0 , \1973_b1 , \1973_b0 , \1974_b1 , \1974_b0 , \1975_b1 , \1975_b0 , \1976_b1 , \1976_b0 , 
		\1977_b1 , \1977_b0 , \1978_b1 , \1978_b0 , \1979_b1 , \1979_b0 , \1980_b1 , \1980_b0 , \1981_b1 , \1981_b0 , 
		\1982_b1 , \1982_b0 , \1983_b1 , \1983_b0 , \1984_b1 , \1984_b0 , \1985_b1 , \1985_b0 , \1986_b1 , \1986_b0 , 
		\1987_b1 , \1987_b0 , \1988_b1 , \1988_b0 , \1989_b1 , \1989_b0 , \1990_b1 , \1990_b0 , \1991_b1 , \1991_b0 , 
		\1992_b1 , \1992_b0 , \1993_b1 , \1993_b0 , \1994_b1 , \1994_b0 , \1995_b1 , \1995_b0 , \1996_b1 , \1996_b0 , 
		\1997_b1 , \1997_b0 , \1998_b1 , \1998_b0 , \1999_b1 , \1999_b0 , \2000_b1 , \2000_b0 , \2001_b1 , \2001_b0 , 
		\2002_b1 , \2002_b0 , \2003_b1 , \2003_b0 , \2004_b1 , \2004_b0 , \2005_b1 , \2005_b0 , \2006_b1 , \2006_b0 , 
		\2007_b1 , \2007_b0 , \2008_b1 , \2008_b0 , \2009_b1 , \2009_b0 , \2010_b1 , \2010_b0 , \2011_b1 , \2011_b0 , 
		\2012_b1 , \2012_b0 , \2013_b1 , \2013_b0 , \2014_b1 , \2014_b0 , \2015_b1 , \2015_b0 , \2016_b1 , \2016_b0 , 
		\2017_b1 , \2017_b0 , \2018_b1 , \2018_b0 , \2019_b1 , \2019_b0 , \2020_b1 , \2020_b0 , \2021_b1 , \2021_b0 , 
		\2022_b1 , \2022_b0 , \2023_B[11]_b1 , \2023_B[11]_b0 , \2024_b1 , \2024_b0 , \2025_b1 , \2025_b0 , \2026_Z[11]_b1 , \2026_Z[11]_b0 , 
		\2027_b1 , \2027_b0 , \2028_A[11]_b1 , \2028_A[11]_b0 , \2029_B[11]_b1 , \2029_B[11]_b0 , \2030_b1 , \2030_b0 , \2031_b1 , \2031_b0 , 
		\2032_b1 , \2032_b0 , \2033_b1 , \2033_b0 , \2034_b1 , \2034_b0 , \2035_b1 , \2035_b0 , \2036_SUM[11]_b1 , \2036_SUM[11]_b0 , 
		\2037_b1 , \2037_b0 , \2038_A[11]_b1 , \2038_A[11]_b0 , \2039_B[11]_b1 , \2039_B[11]_b0 , \2040_b1 , \2040_b0 , \2041_b1 , \2041_b0 , 
		\2042_b1 , \2042_b0 , \2043_b1 , \2043_b0 , \2044_b1 , \2044_b0 , \2045_b1 , \2045_b0 , \2046_SUM[11]_b1 , \2046_SUM[11]_b0 , 
		\2047_b1 , \2047_b0 , \2048_b1 , \2048_b0 , \2049_b1 , \2049_b0 , \2050_b1 , \2050_b0 , \2051_b1 , \2051_b0 , 
		\2052_b1 , \2052_b0 , \2053_b1 , \2053_b0 , \2054_b1 , \2054_b0 , \2055_b1 , \2055_b0 , \2056_b1 , \2056_b0 , 
		\2057_b1 , \2057_b0 , \2058_b1 , \2058_b0 , \2059_b1 , \2059_b0 , \2060_b1 , \2060_b0 , \2061_b1 , \2061_b0 , 
		\2062_A[12]_b1 , \2062_A[12]_b0 , \2063_b1 , \2063_b0 , \2064_b1 , \2064_b0 , \2065_b1 , \2065_b0 , \2066_b1 , \2066_b0 , 
		\2067_b1 , \2067_b0 , \2068_b1 , \2068_b0 , \2069_b1 , \2069_b0 , \2070_b1 , \2070_b0 , \2071_b1 , \2071_b0 , 
		\2072_b1 , \2072_b0 , \2073_b1 , \2073_b0 , \2074_b1 , \2074_b0 , \2075_b1 , \2075_b0 , \2076_b1 , \2076_b0 , 
		\2077_b1 , \2077_b0 , \2078_b1 , \2078_b0 , \2079_b1 , \2079_b0 , \2080_b1 , \2080_b0 , \2081_b1 , \2081_b0 , 
		\2082_b1 , \2082_b0 , \2083_b1 , \2083_b0 , \2084_b1 , \2084_b0 , \2085_b1 , \2085_b0 , \2086_b1 , \2086_b0 , 
		\2087_b1 , \2087_b0 , \2088_b1 , \2088_b0 , \2089_b1 , \2089_b0 , \2090_b1 , \2090_b0 , \2091_b1 , \2091_b0 , 
		\2092_b1 , \2092_b0 , \2093_b1 , \2093_b0 , \2094_b1 , \2094_b0 , \2095_b1 , \2095_b0 , \2096_b1 , \2096_b0 , 
		\2097_b1 , \2097_b0 , \2098_b1 , \2098_b0 , \2099_b1 , \2099_b0 , \2100_b1 , \2100_b0 , \2101_b1 , \2101_b0 , 
		\2102_b1 , \2102_b0 , \2103_b1 , \2103_b0 , \2104_b1 , \2104_b0 , \2105_b1 , \2105_b0 , \2106_b1 , \2106_b0 , 
		\2107_b1 , \2107_b0 , \2108_b1 , \2108_b0 , \2109_b1 , \2109_b0 , \2110_b1 , \2110_b0 , \2111_b1 , \2111_b0 , 
		\2112_b1 , \2112_b0 , \2113_b1 , \2113_b0 , \2114_b1 , \2114_b0 , \2115_b1 , \2115_b0 , \2116_b1 , \2116_b0 , 
		\2117_b1 , \2117_b0 , \2118_b1 , \2118_b0 , \2119_b1 , \2119_b0 , \2120_b1 , \2120_b0 , \2121_b1 , \2121_b0 , 
		\2122_b1 , \2122_b0 , \2123_b1 , \2123_b0 , \2124_b1 , \2124_b0 , \2125_b1 , \2125_b0 , \2126_b1 , \2126_b0 , 
		\2127_b1 , \2127_b0 , \2128_B[12]_b1 , \2128_B[12]_b0 , \2129_b1 , \2129_b0 , \2130_b1 , \2130_b0 , \2131_Z[12]_b1 , \2131_Z[12]_b0 , 
		\2132_b1 , \2132_b0 , \2133_A[12]_b1 , \2133_A[12]_b0 , \2134_b1 , \2134_b0 , \2135_b1 , \2135_b0 , \2136_b1 , \2136_b0 , 
		\2137_b1 , \2137_b0 , \2138_b1 , \2138_b0 , \2139_b1 , \2139_b0 , \2140_b1 , \2140_b0 , \2141_b1 , \2141_b0 , 
		\2142_b1 , \2142_b0 , \2143_b1 , \2143_b0 , \2144_b1 , \2144_b0 , \2145_b1 , \2145_b0 , \2146_b1 , \2146_b0 , 
		\2147_b1 , \2147_b0 , \2148_b1 , \2148_b0 , \2149_b1 , \2149_b0 , \2150_b1 , \2150_b0 , \2151_b1 , \2151_b0 , 
		\2152_b1 , \2152_b0 , \2153_b1 , \2153_b0 , \2154_b1 , \2154_b0 , \2155_b1 , \2155_b0 , \2156_b1 , \2156_b0 , 
		\2157_b1 , \2157_b0 , \2158_b1 , \2158_b0 , \2159_b1 , \2159_b0 , \2160_b1 , \2160_b0 , \2161_b1 , \2161_b0 , 
		\2162_b1 , \2162_b0 , \2163_b1 , \2163_b0 , \2164_b1 , \2164_b0 , \2165_b1 , \2165_b0 , \2166_b1 , \2166_b0 , 
		\2167_b1 , \2167_b0 , \2168_b1 , \2168_b0 , \2169_b1 , \2169_b0 , \2170_b1 , \2170_b0 , \2171_b1 , \2171_b0 , 
		\2172_b1 , \2172_b0 , \2173_b1 , \2173_b0 , \2174_b1 , \2174_b0 , \2175_b1 , \2175_b0 , \2176_b1 , \2176_b0 , 
		\2177_b1 , \2177_b0 , \2178_b1 , \2178_b0 , \2179_b1 , \2179_b0 , \2180_b1 , \2180_b0 , \2181_b1 , \2181_b0 , 
		\2182_b1 , \2182_b0 , \2183_b1 , \2183_b0 , \2184_b1 , \2184_b0 , \2185_b1 , \2185_b0 , \2186_b1 , \2186_b0 , 
		\2187_b1 , \2187_b0 , \2188_b1 , \2188_b0 , \2189_b1 , \2189_b0 , \2190_b1 , \2190_b0 , \2191_b1 , \2191_b0 , 
		\2192_b1 , \2192_b0 , \2193_b1 , \2193_b0 , \2194_b1 , \2194_b0 , \2195_b1 , \2195_b0 , \2196_b1 , \2196_b0 , 
		\2197_b1 , \2197_b0 , \2198_b1 , \2198_b0 , \2199_B[12]_b1 , \2199_B[12]_b0 , \2200_b1 , \2200_b0 , \2201_b1 , \2201_b0 , 
		\2202_Z[12]_b1 , \2202_Z[12]_b0 , \2203_b1 , \2203_b0 , \2204_A[12]_b1 , \2204_A[12]_b0 , \2205_B[12]_b1 , \2205_B[12]_b0 , \2206_b1 , \2206_b0 , 
		\2207_b1 , \2207_b0 , \2208_b1 , \2208_b0 , \2209_b1 , \2209_b0 , \2210_b1 , \2210_b0 , \2211_b1 , \2211_b0 , 
		\2212_SUM[12]_b1 , \2212_SUM[12]_b0 , \2213_b1 , \2213_b0 , \2214_A[12]_b1 , \2214_A[12]_b0 , \2215_B[12]_b1 , \2215_B[12]_b0 , \2216_b1 , \2216_b0 , 
		\2217_b1 , \2217_b0 , \2218_b1 , \2218_b0 , \2219_b1 , \2219_b0 , \2220_b1 , \2220_b0 , \2221_b1 , \2221_b0 , 
		\2222_SUM[12]_b1 , \2222_SUM[12]_b0 , \2223_b1 , \2223_b0 , \2224_b1 , \2224_b0 , \2225_b1 , \2225_b0 , \2226_b1 , \2226_b0 , 
		\2227_b1 , \2227_b0 , \2228_b1 , \2228_b0 , \2229_b1 , \2229_b0 , \2230_b1 , \2230_b0 , \2231_b1 , \2231_b0 , 
		\2232_b1 , \2232_b0 , \2233_b1 , \2233_b0 , \2234_b1 , \2234_b0 , \2235_b1 , \2235_b0 , \2236_b1 , \2236_b0 , 
		\2237_b1 , \2237_b0 , \2238_A[13]_b1 , \2238_A[13]_b0 , \2239_b1 , \2239_b0 , \2240_b1 , \2240_b0 , \2241_b1 , \2241_b0 , 
		\2242_b1 , \2242_b0 , \2243_b1 , \2243_b0 , \2244_b1 , \2244_b0 , \2245_b1 , \2245_b0 , \2246_b1 , \2246_b0 , 
		\2247_b1 , \2247_b0 , \2248_b1 , \2248_b0 , \2249_b1 , \2249_b0 , \2250_b1 , \2250_b0 , \2251_b1 , \2251_b0 , 
		\2252_b1 , \2252_b0 , \2253_b1 , \2253_b0 , \2254_b1 , \2254_b0 , \2255_b1 , \2255_b0 , \2256_b1 , \2256_b0 , 
		\2257_b1 , \2257_b0 , \2258_b1 , \2258_b0 , \2259_b1 , \2259_b0 , \2260_b1 , \2260_b0 , \2261_b1 , \2261_b0 , 
		\2262_b1 , \2262_b0 , \2263_b1 , \2263_b0 , \2264_b1 , \2264_b0 , \2265_b1 , \2265_b0 , \2266_b1 , \2266_b0 , 
		\2267_b1 , \2267_b0 , \2268_b1 , \2268_b0 , \2269_b1 , \2269_b0 , \2270_b1 , \2270_b0 , \2271_b1 , \2271_b0 , 
		\2272_b1 , \2272_b0 , \2273_b1 , \2273_b0 , \2274_b1 , \2274_b0 , \2275_b1 , \2275_b0 , \2276_b1 , \2276_b0 , 
		\2277_b1 , \2277_b0 , \2278_b1 , \2278_b0 , \2279_b1 , \2279_b0 , \2280_b1 , \2280_b0 , \2281_b1 , \2281_b0 , 
		\2282_b1 , \2282_b0 , \2283_b1 , \2283_b0 , \2284_b1 , \2284_b0 , \2285_b1 , \2285_b0 , \2286_b1 , \2286_b0 , 
		\2287_b1 , \2287_b0 , \2288_b1 , \2288_b0 , \2289_b1 , \2289_b0 , \2290_b1 , \2290_b0 , \2291_b1 , \2291_b0 , 
		\2292_b1 , \2292_b0 , \2293_b1 , \2293_b0 , \2294_b1 , \2294_b0 , \2295_b1 , \2295_b0 , \2296_b1 , \2296_b0 , 
		\2297_b1 , \2297_b0 , \2298_b1 , \2298_b0 , \2299_b1 , \2299_b0 , \2300_b1 , \2300_b0 , \2301_b1 , \2301_b0 , 
		\2302_b1 , \2302_b0 , \2303_b1 , \2303_b0 , \2304_b1 , \2304_b0 , \2305_b1 , \2305_b0 , \2306_b1 , \2306_b0 , 
		\2307_b1 , \2307_b0 , \2308_b1 , \2308_b0 , \2309_b1 , \2309_b0 , \2310_B[13]_b1 , \2310_B[13]_b0 , \2311_b1 , \2311_b0 , 
		\2312_b1 , \2312_b0 , \2313_Z[13]_b1 , \2313_Z[13]_b0 , \2314_b1 , \2314_b0 , \2315_A[13]_b1 , \2315_A[13]_b0 , \2316_b1 , \2316_b0 , 
		\2317_b1 , \2317_b0 , \2318_b1 , \2318_b0 , \2319_b1 , \2319_b0 , \2320_b1 , \2320_b0 , \2321_b1 , \2321_b0 , 
		\2322_b1 , \2322_b0 , \2323_b1 , \2323_b0 , \2324_b1 , \2324_b0 , \2325_b1 , \2325_b0 , \2326_b1 , \2326_b0 , 
		\2327_b1 , \2327_b0 , \2328_b1 , \2328_b0 , \2329_b1 , \2329_b0 , \2330_b1 , \2330_b0 , \2331_b1 , \2331_b0 , 
		\2332_b1 , \2332_b0 , \2333_b1 , \2333_b0 , \2334_b1 , \2334_b0 , \2335_b1 , \2335_b0 , \2336_b1 , \2336_b0 , 
		\2337_b1 , \2337_b0 , \2338_b1 , \2338_b0 , \2339_b1 , \2339_b0 , \2340_b1 , \2340_b0 , \2341_b1 , \2341_b0 , 
		\2342_b1 , \2342_b0 , \2343_b1 , \2343_b0 , \2344_b1 , \2344_b0 , \2345_b1 , \2345_b0 , \2346_b1 , \2346_b0 , 
		\2347_b1 , \2347_b0 , \2348_b1 , \2348_b0 , \2349_b1 , \2349_b0 , \2350_b1 , \2350_b0 , \2351_b1 , \2351_b0 , 
		\2352_b1 , \2352_b0 , \2353_b1 , \2353_b0 , \2354_b1 , \2354_b0 , \2355_b1 , \2355_b0 , \2356_b1 , \2356_b0 , 
		\2357_b1 , \2357_b0 , \2358_b1 , \2358_b0 , \2359_b1 , \2359_b0 , \2360_b1 , \2360_b0 , \2361_b1 , \2361_b0 , 
		\2362_b1 , \2362_b0 , \2363_b1 , \2363_b0 , \2364_b1 , \2364_b0 , \2365_b1 , \2365_b0 , \2366_b1 , \2366_b0 , 
		\2367_b1 , \2367_b0 , \2368_b1 , \2368_b0 , \2369_b1 , \2369_b0 , \2370_b1 , \2370_b0 , \2371_b1 , \2371_b0 , 
		\2372_b1 , \2372_b0 , \2373_b1 , \2373_b0 , \2374_b1 , \2374_b0 , \2375_b1 , \2375_b0 , \2376_b1 , \2376_b0 , 
		\2377_b1 , \2377_b0 , \2378_b1 , \2378_b0 , \2379_b1 , \2379_b0 , \2380_b1 , \2380_b0 , \2381_b1 , \2381_b0 , 
		\2382_b1 , \2382_b0 , \2383_b1 , \2383_b0 , \2384_b1 , \2384_b0 , \2385_b1 , \2385_b0 , \2386_b1 , \2386_b0 , 
		\2387_B[13]_b1 , \2387_B[13]_b0 , \2388_b1 , \2388_b0 , \2389_b1 , \2389_b0 , \2390_Z[13]_b1 , \2390_Z[13]_b0 , \2391_b1 , \2391_b0 , 
		\2392_A[13]_b1 , \2392_A[13]_b0 , \2393_B[13]_b1 , \2393_B[13]_b0 , \2394_b1 , \2394_b0 , \2395_b1 , \2395_b0 , \2396_b1 , \2396_b0 , 
		\2397_b1 , \2397_b0 , \2398_b1 , \2398_b0 , \2399_b1 , \2399_b0 , \2400_SUM[13]_b1 , \2400_SUM[13]_b0 , \2401_b1 , \2401_b0 , 
		\2402_A[13]_b1 , \2402_A[13]_b0 , \2403_B[13]_b1 , \2403_B[13]_b0 , \2404_b1 , \2404_b0 , \2405_b1 , \2405_b0 , \2406_b1 , \2406_b0 , 
		\2407_b1 , \2407_b0 , \2408_b1 , \2408_b0 , \2409_b1 , \2409_b0 , \2410_SUM[13]_b1 , \2410_SUM[13]_b0 , \2411_b1 , \2411_b0 , 
		\2412_b1 , \2412_b0 , \2413_b1 , \2413_b0 , \2414_b1 , \2414_b0 , \2415_b1 , \2415_b0 , \2416_b1 , \2416_b0 , 
		\2417_b1 , \2417_b0 , \2418_b1 , \2418_b0 , \2419_b1 , \2419_b0 , \2420_b1 , \2420_b0 , \2421_b1 , \2421_b0 , 
		\2422_b1 , \2422_b0 , \2423_b1 , \2423_b0 , \2424_b1 , \2424_b0 , \2425_b1 , \2425_b0 , \2426_A[14]_b1 , \2426_A[14]_b0 , 
		\2427_b1 , \2427_b0 , \2428_b1 , \2428_b0 , \2429_b1 , \2429_b0 , \2430_b1 , \2430_b0 , \2431_b1 , \2431_b0 , 
		\2432_b1 , \2432_b0 , \2433_b1 , \2433_b0 , \2434_b1 , \2434_b0 , \2435_b1 , \2435_b0 , \2436_b1 , \2436_b0 , 
		\2437_b1 , \2437_b0 , \2438_b1 , \2438_b0 , \2439_b1 , \2439_b0 , \2440_b1 , \2440_b0 , \2441_b1 , \2441_b0 , 
		\2442_b1 , \2442_b0 , \2443_b1 , \2443_b0 , \2444_b1 , \2444_b0 , \2445_b1 , \2445_b0 , \2446_b1 , \2446_b0 , 
		\2447_b1 , \2447_b0 , \2448_b1 , \2448_b0 , \2449_b1 , \2449_b0 , \2450_b1 , \2450_b0 , \2451_b1 , \2451_b0 , 
		\2452_b1 , \2452_b0 , \2453_b1 , \2453_b0 , \2454_b1 , \2454_b0 , \2455_b1 , \2455_b0 , \2456_b1 , \2456_b0 , 
		\2457_b1 , \2457_b0 , \2458_b1 , \2458_b0 , \2459_b1 , \2459_b0 , \2460_b1 , \2460_b0 , \2461_b1 , \2461_b0 , 
		\2462_b1 , \2462_b0 , \2463_b1 , \2463_b0 , \2464_b1 , \2464_b0 , \2465_b1 , \2465_b0 , \2466_b1 , \2466_b0 , 
		\2467_b1 , \2467_b0 , \2468_b1 , \2468_b0 , \2469_b1 , \2469_b0 , \2470_b1 , \2470_b0 , \2471_b1 , \2471_b0 , 
		\2472_b1 , \2472_b0 , \2473_b1 , \2473_b0 , \2474_b1 , \2474_b0 , \2475_b1 , \2475_b0 , \2476_b1 , \2476_b0 , 
		\2477_b1 , \2477_b0 , \2478_b1 , \2478_b0 , \2479_b1 , \2479_b0 , \2480_b1 , \2480_b0 , \2481_b1 , \2481_b0 , 
		\2482_b1 , \2482_b0 , \2483_b1 , \2483_b0 , \2484_b1 , \2484_b0 , \2485_b1 , \2485_b0 , \2486_b1 , \2486_b0 , 
		\2487_b1 , \2487_b0 , \2488_b1 , \2488_b0 , \2489_b1 , \2489_b0 , \2490_b1 , \2490_b0 , \2491_b1 , \2491_b0 , 
		\2492_b1 , \2492_b0 , \2493_b1 , \2493_b0 , \2494_b1 , \2494_b0 , \2495_b1 , \2495_b0 , \2496_b1 , \2496_b0 , 
		\2497_b1 , \2497_b0 , \2498_b1 , \2498_b0 , \2499_b1 , \2499_b0 , \2500_b1 , \2500_b0 , \2501_b1 , \2501_b0 , 
		\2502_b1 , \2502_b0 , \2503_b1 , \2503_b0 , \2504_B[14]_b1 , \2504_B[14]_b0 , \2505_b1 , \2505_b0 , \2506_b1 , \2506_b0 , 
		\2507_Z[14]_b1 , \2507_Z[14]_b0 , \2508_b1 , \2508_b0 , \2509_A[14]_b1 , \2509_A[14]_b0 , \2510_b1 , \2510_b0 , \2511_b1 , \2511_b0 , 
		\2512_b1 , \2512_b0 , \2513_b1 , \2513_b0 , \2514_b1 , \2514_b0 , \2515_b1 , \2515_b0 , \2516_b1 , \2516_b0 , 
		\2517_b1 , \2517_b0 , \2518_b1 , \2518_b0 , \2519_b1 , \2519_b0 , \2520_b1 , \2520_b0 , \2521_b1 , \2521_b0 , 
		\2522_b1 , \2522_b0 , \2523_b1 , \2523_b0 , \2524_b1 , \2524_b0 , \2525_b1 , \2525_b0 , \2526_b1 , \2526_b0 , 
		\2527_b1 , \2527_b0 , \2528_b1 , \2528_b0 , \2529_b1 , \2529_b0 , \2530_b1 , \2530_b0 , \2531_b1 , \2531_b0 , 
		\2532_b1 , \2532_b0 , \2533_b1 , \2533_b0 , \2534_b1 , \2534_b0 , \2535_b1 , \2535_b0 , \2536_b1 , \2536_b0 , 
		\2537_b1 , \2537_b0 , \2538_b1 , \2538_b0 , \2539_b1 , \2539_b0 , \2540_b1 , \2540_b0 , \2541_b1 , \2541_b0 , 
		\2542_b1 , \2542_b0 , \2543_b1 , \2543_b0 , \2544_b1 , \2544_b0 , \2545_b1 , \2545_b0 , \2546_b1 , \2546_b0 , 
		\2547_b1 , \2547_b0 , \2548_b1 , \2548_b0 , \2549_b1 , \2549_b0 , \2550_b1 , \2550_b0 , \2551_b1 , \2551_b0 , 
		\2552_b1 , \2552_b0 , \2553_b1 , \2553_b0 , \2554_b1 , \2554_b0 , \2555_b1 , \2555_b0 , \2556_b1 , \2556_b0 , 
		\2557_b1 , \2557_b0 , \2558_b1 , \2558_b0 , \2559_b1 , \2559_b0 , \2560_b1 , \2560_b0 , \2561_b1 , \2561_b0 , 
		\2562_b1 , \2562_b0 , \2563_b1 , \2563_b0 , \2564_b1 , \2564_b0 , \2565_b1 , \2565_b0 , \2566_b1 , \2566_b0 , 
		\2567_b1 , \2567_b0 , \2568_b1 , \2568_b0 , \2569_b1 , \2569_b0 , \2570_b1 , \2570_b0 , \2571_b1 , \2571_b0 , 
		\2572_b1 , \2572_b0 , \2573_b1 , \2573_b0 , \2574_b1 , \2574_b0 , \2575_b1 , \2575_b0 , \2576_b1 , \2576_b0 , 
		\2577_b1 , \2577_b0 , \2578_b1 , \2578_b0 , \2579_b1 , \2579_b0 , \2580_b1 , \2580_b0 , \2581_b1 , \2581_b0 , 
		\2582_b1 , \2582_b0 , \2583_b1 , \2583_b0 , \2584_b1 , \2584_b0 , \2585_b1 , \2585_b0 , \2586_b1 , \2586_b0 , 
		\2587_B[14]_b1 , \2587_B[14]_b0 , \2588_b1 , \2588_b0 , \2589_b1 , \2589_b0 , \2590_Z[14]_b1 , \2590_Z[14]_b0 , \2591_b1 , \2591_b0 , 
		\2592_A[14]_b1 , \2592_A[14]_b0 , \2593_B[14]_b1 , \2593_B[14]_b0 , \2594_b1 , \2594_b0 , \2595_b1 , \2595_b0 , \2596_b1 , \2596_b0 , 
		\2597_b1 , \2597_b0 , \2598_b1 , \2598_b0 , \2599_b1 , \2599_b0 , \2600_SUM[14]_b1 , \2600_SUM[14]_b0 , \2601_b1 , \2601_b0 , 
		\2602_A[14]_b1 , \2602_A[14]_b0 , \2603_B[14]_b1 , \2603_B[14]_b0 , \2604_b1 , \2604_b0 , \2605_b1 , \2605_b0 , \2606_b1 , \2606_b0 , 
		\2607_b1 , \2607_b0 , \2608_b1 , \2608_b0 , \2609_b1 , \2609_b0 , \2610_SUM[14]_b1 , \2610_SUM[14]_b0 , \2611_b1 , \2611_b0 , 
		\2612_b1 , \2612_b0 , \2613_b1 , \2613_b0 , \2614_b1 , \2614_b0 , \2615_b1 , \2615_b0 , \2616_b1 , \2616_b0 , 
		\2617_b1 , \2617_b0 , \2618_b1 , \2618_b0 , \2619_b1 , \2619_b0 , \2620_b1 , \2620_b0 , \2621_b1 , \2621_b0 , 
		\2622_b1 , \2622_b0 , \2623_b1 , \2623_b0 , \2624_b1 , \2624_b0 , \2625_b1 , \2625_b0 , \2626_A[15]_b1 , \2626_A[15]_b0 , 
		\2627_b1 , \2627_b0 , \2628_b1 , \2628_b0 , \2629_b1 , \2629_b0 , \2630_b1 , \2630_b0 , \2631_b1 , \2631_b0 , 
		\2632_b1 , \2632_b0 , \2633_b1 , \2633_b0 , \2634_b1 , \2634_b0 , \2635_b1 , \2635_b0 , \2636_b1 , \2636_b0 , 
		\2637_b1 , \2637_b0 , \2638_b1 , \2638_b0 , \2639_b1 , \2639_b0 , \2640_b1 , \2640_b0 , \2641_b1 , \2641_b0 , 
		\2642_b1 , \2642_b0 , \2643_b1 , \2643_b0 , \2644_b1 , \2644_b0 , \2645_b1 , \2645_b0 , \2646_b1 , \2646_b0 , 
		\2647_b1 , \2647_b0 , \2648_b1 , \2648_b0 , \2649_b1 , \2649_b0 , \2650_b1 , \2650_b0 , \2651_b1 , \2651_b0 , 
		\2652_b1 , \2652_b0 , \2653_b1 , \2653_b0 , \2654_b1 , \2654_b0 , \2655_b1 , \2655_b0 , \2656_b1 , \2656_b0 , 
		\2657_b1 , \2657_b0 , \2658_b1 , \2658_b0 , \2659_b1 , \2659_b0 , \2660_b1 , \2660_b0 , \2661_b1 , \2661_b0 , 
		\2662_b1 , \2662_b0 , \2663_b1 , \2663_b0 , \2664_b1 , \2664_b0 , \2665_b1 , \2665_b0 , \2666_b1 , \2666_b0 , 
		\2667_b1 , \2667_b0 , \2668_b1 , \2668_b0 , \2669_b1 , \2669_b0 , \2670_b1 , \2670_b0 , \2671_b1 , \2671_b0 , 
		\2672_b1 , \2672_b0 , \2673_b1 , \2673_b0 , \2674_b1 , \2674_b0 , \2675_b1 , \2675_b0 , \2676_b1 , \2676_b0 , 
		\2677_b1 , \2677_b0 , \2678_b1 , \2678_b0 , \2679_b1 , \2679_b0 , \2680_b1 , \2680_b0 , \2681_b1 , \2681_b0 , 
		\2682_b1 , \2682_b0 , \2683_b1 , \2683_b0 , \2684_b1 , \2684_b0 , \2685_b1 , \2685_b0 , \2686_b1 , \2686_b0 , 
		\2687_b1 , \2687_b0 , \2688_b1 , \2688_b0 , \2689_b1 , \2689_b0 , \2690_b1 , \2690_b0 , \2691_b1 , \2691_b0 , 
		\2692_b1 , \2692_b0 , \2693_b1 , \2693_b0 , \2694_b1 , \2694_b0 , \2695_b1 , \2695_b0 , \2696_b1 , \2696_b0 , 
		\2697_b1 , \2697_b0 , \2698_b1 , \2698_b0 , \2699_b1 , \2699_b0 , \2700_b1 , \2700_b0 , \2701_b1 , \2701_b0 , 
		\2702_b1 , \2702_b0 , \2703_b1 , \2703_b0 , \2704_b1 , \2704_b0 , \2705_b1 , \2705_b0 , \2706_b1 , \2706_b0 , 
		\2707_b1 , \2707_b0 , \2708_b1 , \2708_b0 , \2709_b1 , \2709_b0 , \2710_B[15]_b1 , \2710_B[15]_b0 , \2711_b1 , \2711_b0 , 
		\2712_b1 , \2712_b0 , \2713_Z[15]_b1 , \2713_Z[15]_b0 , \2714_b1 , \2714_b0 , \2715_A[15]_b1 , \2715_A[15]_b0 , \2716_b1 , \2716_b0 , 
		\2717_b1 , \2717_b0 , \2718_b1 , \2718_b0 , \2719_b1 , \2719_b0 , \2720_b1 , \2720_b0 , \2721_b1 , \2721_b0 , 
		\2722_b1 , \2722_b0 , \2723_b1 , \2723_b0 , \2724_b1 , \2724_b0 , \2725_b1 , \2725_b0 , \2726_b1 , \2726_b0 , 
		\2727_b1 , \2727_b0 , \2728_b1 , \2728_b0 , \2729_b1 , \2729_b0 , \2730_b1 , \2730_b0 , \2731_b1 , \2731_b0 , 
		\2732_b1 , \2732_b0 , \2733_b1 , \2733_b0 , \2734_b1 , \2734_b0 , \2735_b1 , \2735_b0 , \2736_b1 , \2736_b0 , 
		\2737_b1 , \2737_b0 , \2738_b1 , \2738_b0 , \2739_b1 , \2739_b0 , \2740_b1 , \2740_b0 , \2741_b1 , \2741_b0 , 
		\2742_b1 , \2742_b0 , \2743_b1 , \2743_b0 , \2744_b1 , \2744_b0 , \2745_b1 , \2745_b0 , \2746_b1 , \2746_b0 , 
		\2747_b1 , \2747_b0 , \2748_b1 , \2748_b0 , \2749_b1 , \2749_b0 , \2750_b1 , \2750_b0 , \2751_b1 , \2751_b0 , 
		\2752_b1 , \2752_b0 , \2753_b1 , \2753_b0 , \2754_b1 , \2754_b0 , \2755_b1 , \2755_b0 , \2756_b1 , \2756_b0 , 
		\2757_b1 , \2757_b0 , \2758_b1 , \2758_b0 , \2759_b1 , \2759_b0 , \2760_b1 , \2760_b0 , \2761_b1 , \2761_b0 , 
		\2762_b1 , \2762_b0 , \2763_b1 , \2763_b0 , \2764_b1 , \2764_b0 , \2765_b1 , \2765_b0 , \2766_b1 , \2766_b0 , 
		\2767_b1 , \2767_b0 , \2768_b1 , \2768_b0 , \2769_b1 , \2769_b0 , \2770_b1 , \2770_b0 , \2771_b1 , \2771_b0 , 
		\2772_b1 , \2772_b0 , \2773_b1 , \2773_b0 , \2774_b1 , \2774_b0 , \2775_b1 , \2775_b0 , \2776_b1 , \2776_b0 , 
		\2777_b1 , \2777_b0 , \2778_b1 , \2778_b0 , \2779_b1 , \2779_b0 , \2780_b1 , \2780_b0 , \2781_b1 , \2781_b0 , 
		\2782_b1 , \2782_b0 , \2783_b1 , \2783_b0 , \2784_b1 , \2784_b0 , \2785_b1 , \2785_b0 , \2786_b1 , \2786_b0 , 
		\2787_b1 , \2787_b0 , \2788_b1 , \2788_b0 , \2789_b1 , \2789_b0 , \2790_b1 , \2790_b0 , \2791_b1 , \2791_b0 , 
		\2792_b1 , \2792_b0 , \2793_b1 , \2793_b0 , \2794_b1 , \2794_b0 , \2795_b1 , \2795_b0 , \2796_b1 , \2796_b0 , 
		\2797_b1 , \2797_b0 , \2798_b1 , \2798_b0 , \2799_B[15]_b1 , \2799_B[15]_b0 , \2800_b1 , \2800_b0 , \2801_b1 , \2801_b0 , 
		\2802_Z[15]_b1 , \2802_Z[15]_b0 , \2803_b1 , \2803_b0 , \2804_A[15]_b1 , \2804_A[15]_b0 , \2805_B[15]_b1 , \2805_B[15]_b0 , \2806_b1 , \2806_b0 , 
		\2807_b1 , \2807_b0 , \2808_b1 , \2808_b0 , \2809_b1 , \2809_b0 , \2810_b1 , \2810_b0 , \2811_b1 , \2811_b0 , 
		\2812_SUM[15]_b1 , \2812_SUM[15]_b0 , \2813_b1 , \2813_b0 , \2814_A[15]_b1 , \2814_A[15]_b0 , \2815_B[15]_b1 , \2815_B[15]_b0 , \2816_b1 , \2816_b0 , 
		\2817_b1 , \2817_b0 , \2818_b1 , \2818_b0 , \2819_b1 , \2819_b0 , \2820_b1 , \2820_b0 , \2821_b1 , \2821_b0 , 
		\2822_SUM[15]_b1 , \2822_SUM[15]_b0 , \2823_b1 , \2823_b0 , \2824_b1 , \2824_b0 , \2825_b1 , \2825_b0 , \2826_b1 , \2826_b0 , 
		\2827_b1 , \2827_b0 , \2828_b1 , \2828_b0 , \2829_A[15]_b1 , \2829_A[15]_b0 , \2830_B[15]_b1 , \2830_B[15]_b0 , \2831_b1 , \2831_b0 , 
		\2832_A[14]_b1 , \2832_A[14]_b0 , \2833_B[14]_b1 , \2833_B[14]_b0 , \2834_b1 , \2834_b0 , \2835_A[13]_b1 , \2835_A[13]_b0 , \2836_B[13]_b1 , \2836_B[13]_b0 , 
		\2837_b1 , \2837_b0 , \2838_A[12]_b1 , \2838_A[12]_b0 , \2839_B[12]_b1 , \2839_B[12]_b0 , \2840_b1 , \2840_b0 , \2841_A[11]_b1 , \2841_A[11]_b0 , 
		\2842_B[11]_b1 , \2842_B[11]_b0 , \2843_b1 , \2843_b0 , \2844_A[10]_b1 , \2844_A[10]_b0 , \2845_B[10]_b1 , \2845_B[10]_b0 , \2846_b1 , \2846_b0 , 
		\2847_A[9]_b1 , \2847_A[9]_b0 , \2848_B[9]_b1 , \2848_B[9]_b0 , \2849_b1 , \2849_b0 , \2850_A[8]_b1 , \2850_A[8]_b0 , \2851_B[8]_b1 , \2851_B[8]_b0 , 
		\2852_b1 , \2852_b0 , \2853_A[7]_b1 , \2853_A[7]_b0 , \2854_B[7]_b1 , \2854_B[7]_b0 , \2855_b1 , \2855_b0 , \2856_A[6]_b1 , \2856_A[6]_b0 , 
		\2857_B[6]_b1 , \2857_B[6]_b0 , \2858_b1 , \2858_b0 , \2859_A[5]_b1 , \2859_A[5]_b0 , \2860_B[5]_b1 , \2860_B[5]_b0 , \2861_b1 , \2861_b0 , 
		\2862_A[4]_b1 , \2862_A[4]_b0 , \2863_B[4]_b1 , \2863_B[4]_b0 , \2864_b1 , \2864_b0 , \2865_A[3]_b1 , \2865_A[3]_b0 , \2866_B[3]_b1 , \2866_B[3]_b0 , 
		\2867_b1 , \2867_b0 , \2868_A[2]_b1 , \2868_A[2]_b0 , \2869_B[2]_b1 , \2869_B[2]_b0 , \2870_b1 , \2870_b0 , \2871_A[1]_b1 , \2871_A[1]_b0 , 
		\2872_B[1]_b1 , \2872_B[1]_b0 , \2873_b1 , \2873_b0 , \2874_A[0]_b1 , \2874_A[0]_b0 , \2875_B[0]_b1 , \2875_B[0]_b0 , \2876_b1 , \2876_b0 , 
		\2877_b1 , \2877_b0 , \2878_b1 , \2878_b0 , \2879_b1 , \2879_b0 , \2880_b1 , \2880_b0 , \2881_b1 , \2881_b0 , 
		\2882_b1 , \2882_b0 , \2883_b1 , \2883_b0 , \2884_b1 , \2884_b0 , \2885_b1 , \2885_b0 , \2886_b1 , \2886_b0 , 
		\2887_b1 , \2887_b0 , \2888_b1 , \2888_b0 , \2889_b1 , \2889_b0 , \2890_b1 , \2890_b0 , \2891_b1 , \2891_b0 , 
		\2892_b1 , \2892_b0 , \2893_b1 , \2893_b0 , \2894_b1 , \2894_b0 , \2895_b1 , \2895_b0 , \2896_b1 , \2896_b0 , 
		\2897_b1 , \2897_b0 , \2898_b1 , \2898_b0 , \2899_b1 , \2899_b0 , \2900_b1 , \2900_b0 , \2901_b1 , \2901_b0 , 
		\2902_b1 , \2902_b0 , \2903_b1 , \2903_b0 , \2904_b1 , \2904_b0 , \2905_b1 , \2905_b0 , \2906_b1 , \2906_b0 , 
		\2907_b1 , \2907_b0 , \2908_b1 , \2908_b0 , \2909_b1 , \2909_b0 , \2910_b1 , \2910_b0 , \2911_b1 , \2911_b0 , 
		\2912_b1 , \2912_b0 , \2913_b1 , \2913_b0 , \2914_b1 , \2914_b0 , \2915_b1 , \2915_b0 , \2916_b1 , \2916_b0 , 
		\2917_b1 , \2917_b0 , \2918_b1 , \2918_b0 , \2919_b1 , \2919_b0 , \2920_b1 , \2920_b0 , \2921_b1 , \2921_b0 , 
		\2922_SUM[16]_b1 , \2922_SUM[16]_b0 , \2923_A[16]_b1 , \2923_A[16]_b0 , \2924_b1 , \2924_b0 , \2925_b1 , \2925_b0 , \2926_SUM[15]_b1 , \2926_SUM[15]_b0 , 
		\2927_A[15]_b1 , \2927_A[15]_b0 , \2928_b1 , \2928_b0 , \2929_b1 , \2929_b0 , \2930_SUM[14]_b1 , \2930_SUM[14]_b0 , \2931_A[14]_b1 , \2931_A[14]_b0 , 
		\2932_b1 , \2932_b0 , \2933_b1 , \2933_b0 , \2934_SUM[13]_b1 , \2934_SUM[13]_b0 , \2935_A[13]_b1 , \2935_A[13]_b0 , \2936_b1 , \2936_b0 , 
		\2937_b1 , \2937_b0 , \2938_SUM[12]_b1 , \2938_SUM[12]_b0 , \2939_A[12]_b1 , \2939_A[12]_b0 , \2940_b1 , \2940_b0 , \2941_b1 , \2941_b0 , 
		\2942_SUM[11]_b1 , \2942_SUM[11]_b0 , \2943_A[11]_b1 , \2943_A[11]_b0 , \2944_b1 , \2944_b0 , \2945_b1 , \2945_b0 , \2946_SUM[10]_b1 , \2946_SUM[10]_b0 , 
		\2947_A[10]_b1 , \2947_A[10]_b0 , \2948_b1 , \2948_b0 , \2949_b1 , \2949_b0 , \2950_SUM[9]_b1 , \2950_SUM[9]_b0 , \2951_A[9]_b1 , \2951_A[9]_b0 , 
		\2952_b1 , \2952_b0 , \2953_b1 , \2953_b0 , \2954_SUM[8]_b1 , \2954_SUM[8]_b0 , \2955_A[8]_b1 , \2955_A[8]_b0 , \2956_b1 , \2956_b0 , 
		\2957_b1 , \2957_b0 , \2958_SUM[7]_b1 , \2958_SUM[7]_b0 , \2959_A[7]_b1 , \2959_A[7]_b0 , \2960_b1 , \2960_b0 , \2961_b1 , \2961_b0 , 
		\2962_SUM[6]_b1 , \2962_SUM[6]_b0 , \2963_A[6]_b1 , \2963_A[6]_b0 , \2964_b1 , \2964_b0 , \2965_b1 , \2965_b0 , \2966_SUM[5]_b1 , \2966_SUM[5]_b0 , 
		\2967_A[5]_b1 , \2967_A[5]_b0 , \2968_b1 , \2968_b0 , \2969_b1 , \2969_b0 , \2970_SUM[4]_b1 , \2970_SUM[4]_b0 , \2971_A[4]_b1 , \2971_A[4]_b0 , 
		\2972_b1 , \2972_b0 , \2973_b1 , \2973_b0 , \2974_SUM[3]_b1 , \2974_SUM[3]_b0 , \2975_A[3]_b1 , \2975_A[3]_b0 , \2976_b1 , \2976_b0 , 
		\2977_b1 , \2977_b0 , \2978_SUM[2]_b1 , \2978_SUM[2]_b0 , \2979_A[2]_b1 , \2979_A[2]_b0 , \2980_b1 , \2980_b0 , \2981_b1 , \2981_b0 , 
		\2982_SUM[1]_b1 , \2982_SUM[1]_b0 , \2983_A[1]_b1 , \2983_A[1]_b0 , \2984_b1 , \2984_b0 , \2985_SUM[0]_b1 , \2985_SUM[0]_b0 , \2986_A[0]_b1 , \2986_A[0]_b0 , 
		\2987_B[15]_b1 , \2987_B[15]_b0 , \2988_B[14]_b1 , \2988_B[14]_b0 , \2989_B[13]_b1 , \2989_B[13]_b0 , \2990_B[12]_b1 , \2990_B[12]_b0 , \2991_B[11]_b1 , \2991_B[11]_b0 , 
		\2992_B[10]_b1 , \2992_B[10]_b0 , \2993_B[9]_b1 , \2993_B[9]_b0 , \2994_B[8]_b1 , \2994_B[8]_b0 , \2995_B[7]_b1 , \2995_B[7]_b0 , \2996_B[6]_b1 , \2996_B[6]_b0 , 
		\2997_B[5]_b1 , \2997_B[5]_b0 , \2998_B[4]_b1 , \2998_B[4]_b0 , \2999_B[3]_b1 , \2999_B[3]_b0 , \3000_B[2]_b1 , \3000_B[2]_b0 , \3001_B[1]_b1 , \3001_B[1]_b0 , 
		\3002_B[0]_b1 , \3002_B[0]_b0 , \3003_b1 , \3003_b0 , \3004_b1 , \3004_b0 , \3005_b1 , \3005_b0 , \3006_b1 , \3006_b0 , 
		\3007_b1 , \3007_b0 , \3008_b1 , \3008_b0 , \3009_b1 , \3009_b0 , \3010_b1 , \3010_b0 , \3011_b1 , \3011_b0 , 
		\3012_b1 , \3012_b0 , \3013_b1 , \3013_b0 , \3014_b1 , \3014_b0 , \3015_b1 , \3015_b0 , \3016_b1 , \3016_b0 , 
		\3017_b1 , \3017_b0 , \3018_b1 , \3018_b0 , \3019_b1 , \3019_b0 , \3020_b1 , \3020_b0 , \3021_b1 , \3021_b0 , 
		\3022_b1 , \3022_b0 , \3023_b1 , \3023_b0 , \3024_b1 , \3024_b0 , \3025_b1 , \3025_b0 , \3026_b1 , \3026_b0 , 
		\3027_b1 , \3027_b0 , \3028_b1 , \3028_b0 , \3029_b1 , \3029_b0 , \3030_b1 , \3030_b0 , \3031_b1 , \3031_b0 , 
		\3032_b1 , \3032_b0 , \3033_b1 , \3033_b0 , \3034_b1 , \3034_b0 , \3035_b1 , \3035_b0 , \3036_b1 , \3036_b0 , 
		\3037_b1 , \3037_b0 , \3038_b1 , \3038_b0 , \3039_b1 , \3039_b0 , \3040_b1 , \3040_b0 , \3041_b1 , \3041_b0 , 
		\3042_b1 , \3042_b0 , \3043_b1 , \3043_b0 , \3044_b1 , \3044_b0 , \3045_b1 , \3045_b0 , \3046_b1 , \3046_b0 , 
		\3047_b1 , \3047_b0 , \3048_b1 , \3048_b0 , \3049_b1 , \3049_b0 , \3050_b1 , \3050_b0 , \3051_b1 , \3051_b0 , 
		\3052_b1 , \3052_b0 , \3053_b1 , \3053_b0 , \3054_b1 , \3054_b0 , \3055_b1 , \3055_b0 , \3056_b1 , \3056_b0 , 
		\3057_b1 , \3057_b0 , \3058_b1 , \3058_b0 , \3059_b1 , \3059_b0 , \3060_b1 , \3060_b0 , \3061_b1 , \3061_b0 , 
		\3062_b1 , \3062_b0 , \3063_b1 , \3063_b0 , \3064_b1 , \3064_b0 , \3065_b1 , \3065_b0 , \3066_b1 , \3066_b0 , 
		\3067_b1 , \3067_b0 , \3068_b1 , \3068_b0 , \3069_b1 , \3069_b0 , \3070_b1 , \3070_b0 , \3071_b1 , \3071_b0 , 
		\3072_b1 , \3072_b0 , \3073_b1 , \3073_b0 , \3074_b1 , \3074_b0 , \3075_b1 , \3075_b0 , \3076_b1 , \3076_b0 , 
		\3077_b1 , \3077_b0 , \3078_b1 , \3078_b0 , \3079_b1 , \3079_b0 , \3080_b1 , \3080_b0 , \3081_b1 , \3081_b0 , 
		\3082_b1 , \3082_b0 , \3083_b1 , \3083_b0 , \3084_b1 , \3084_b0 , \3085_b1 , \3085_b0 , \3086_b1 , \3086_b0 , 
		\3087_b1 , \3087_b0 , \3088_b1 , \3088_b0 , \3089_b1 , \3089_b0 , \3090_b1 , \3090_b0 , \3091_b1 , \3091_b0 , 
		\3092_b1 , \3092_b0 , \3093_b1 , \3093_b0 , \3094_b1 , \3094_b0 , \3095_b1 , \3095_b0 , \3096_b1 , \3096_b0 , 
		\3097_b1 , \3097_b0 , \3098_b1 , \3098_b0 , \3099_b1 , \3099_b0 , \3100_b1 , \3100_b0 , \3101_b1 , \3101_b0 , 
		\3102_b1 , \3102_b0 , \3103_b1 , \3103_b0 , \3104_b1 , \3104_b0 , \3105_b1 , \3105_b0 , \3106_b1 , \3106_b0 , 
		\3107_b1 , \3107_b0 , \3108_b1 , \3108_b0 , \3109_b1 , \3109_b0 , \3110_b1 , \3110_b0 , \3111_b1 , \3111_b0 , 
		\3112_b1 , \3112_b0 , \3113_b1 , \3113_b0 , \3114_b1 , \3114_b0 , \3115_b1 , \3115_b0 , \3116_b1 , \3116_b0 , 
		\3117_b1 , \3117_b0 , \3118_b1 , \3118_b0 , \3119_b1 , \3119_b0 , \3120_b1 , \3120_b0 , \3121_b1 , \3121_b0 , 
		\3122_b1 , \3122_b0 , \3123_b1 , \3123_b0 , \3124_b1 , \3124_b0 , \3125_b1 , \3125_b0 , \3126_b1 , \3126_b0 , 
		\3127_b1 , \3127_b0 , \3128_b1 , \3128_b0 , \3129_b1 , \3129_b0 , \3130_b1 , \3130_b0 , \3131_b1 , \3131_b0 , 
		\3132_b1 , \3132_b0 , \3133_b1 , \3133_b0 , \3134_b1 , \3134_b0 , \3135_b1 , \3135_b0 , \3136_b1 , \3136_b0 , 
		\3137_b1 , \3137_b0 , \3138_b1 , \3138_b0 , \3139_b1 , \3139_b0 , \3140_b1 , \3140_b0 , \3141_b1 , \3141_b0 , 
		\3142_b1 , \3142_b0 , \3143_b1 , \3143_b0 , \3144_b1 , \3144_b0 , \3145_b1 , \3145_b0 , \3146_b1 , \3146_b0 , 
		\3147_b1 , \3147_b0 , \3148_b1 , \3148_b0 , \3149_b1 , \3149_b0 , \3150_b1 , \3150_b0 , \3151_b1 , \3151_b0 , 
		\3152_b1 , \3152_b0 , \3153_b1 , \3153_b0 , \3154_b1 , \3154_b0 , \3155_b1 , \3155_b0 , \3156_b1 , \3156_b0 , 
		\3157_b1 , \3157_b0 , \3158_b1 , \3158_b0 , \3159_b1 , \3159_b0 , \3160_b1 , \3160_b0 , \3161_b1 , \3161_b0 , 
		\3162_b1 , \3162_b0 , \3163_b1 , \3163_b0 , \3164_b1 , \3164_b0 , \3165_b1 , \3165_b0 , \3166_b1 , \3166_b0 , 
		\3167_b1 , \3167_b0 , \3168_b1 , \3168_b0 , \3169_b1 , \3169_b0 , \3170_b1 , \3170_b0 , \3171_b1 , \3171_b0 , 
		\3172_b1 , \3172_b0 , \3173_b1 , \3173_b0 , \3174_b1 , \3174_b0 , \3175_b1 , \3175_b0 , \3176_b1 , \3176_b0 , 
		\3177_b1 , \3177_b0 , \3178_b1 , \3178_b0 , \3179_b1 , \3179_b0 , \3180_b1 , \3180_b0 , \3181_b1 , \3181_b0 , 
		\3182_b1 , \3182_b0 , \3183_b1 , \3183_b0 , \3184_b1 , \3184_b0 , \3185_b1 , \3185_b0 , \3186_b1 , \3186_b0 , 
		\3187_b1 , \3187_b0 , \3188_b1 , \3188_b0 , \3189_b1 , \3189_b0 , \3190_b1 , \3190_b0 , \3191_b1 , \3191_b0 , 
		\3192_b1 , \3192_b0 , \3193_b1 , \3193_b0 , \3194_b1 , \3194_b0 , \3195_b1 , \3195_b0 , \3196_b1 , \3196_b0 , 
		\3197_b1 , \3197_b0 , \3198_b1 , \3198_b0 , \3199_b1 , \3199_b0 , \3200_b1 , \3200_b0 , \3201_b1 , \3201_b0 , 
		\3202_b1 , \3202_b0 , \3203_b1 , \3203_b0 , \3204_b1 , \3204_b0 , \3205_b1 , \3205_b0 , \3206_b1 , \3206_b0 , 
		\3207_b1 , \3207_b0 , \3208_b1 , \3208_b0 , \3209_b1 , \3209_b0 , \3210_b1 , \3210_b0 , \3211_b1 , \3211_b0 , 
		\3212_b1 , \3212_b0 , \3213_b1 , \3213_b0 , \3214_b1 , \3214_b0 , \3215_b1 , \3215_b0 , \3216_b1 , \3216_b0 , 
		\3217_b1 , \3217_b0 , \3218_b1 , \3218_b0 , \3219_b1 , \3219_b0 , \3220_b1 , \3220_b0 , \3221_b1 , \3221_b0 , 
		\3222_b1 , \3222_b0 , \3223_b1 , \3223_b0 , \3224_b1 , \3224_b0 , \3225_b1 , \3225_b0 , \3226_b1 , \3226_b0 , 
		\3227_b1 , \3227_b0 , \3228_b1 , \3228_b0 , \3229_b1 , \3229_b0 , \3230_b1 , \3230_b0 , \3231_b1 , \3231_b0 , 
		\3232_b1 , \3232_b0 , \3233_b1 , \3233_b0 , \3234_b1 , \3234_b0 , \3235_b1 , \3235_b0 , \3236_b1 , \3236_b0 , 
		\3237_b1 , \3237_b0 , \3238_b1 , \3238_b0 , \3239_b1 , \3239_b0 , \3240_b1 , \3240_b0 , \3241_b1 , \3241_b0 , 
		\3242_b1 , \3242_b0 , \3243_b1 , \3243_b0 , \3244_b1 , \3244_b0 , \3245_b1 , \3245_b0 , \3246_b1 , \3246_b0 , 
		\3247_b1 , \3247_b0 , \3248_b1 , \3248_b0 , \3249_b1 , \3249_b0 , \3250_b1 , \3250_b0 , \3251_b1 , \3251_b0 , 
		\3252_b1 , \3252_b0 , \3253_b1 , \3253_b0 , \3254_b1 , \3254_b0 , \3255_b1 , \3255_b0 , \3256_b1 , \3256_b0 , 
		\3257_b1 , \3257_b0 , \3258_b1 , \3258_b0 , \3259_b1 , \3259_b0 , \3260_b1 , \3260_b0 , \3261_b1 , \3261_b0 , 
		\3262_b1 , \3262_b0 , \3263_b1 , \3263_b0 , \3264_b1 , \3264_b0 , \3265_b1 , \3265_b0 , \3266_b1 , \3266_b0 , 
		\3267_b1 , \3267_b0 , \3268_b1 , \3268_b0 , \3269_b1 , \3269_b0 , \3270_b1 , \3270_b0 , \3271_b1 , \3271_b0 , 
		\3272_b1 , \3272_b0 , \3273_b1 , \3273_b0 , \3274_b1 , \3274_b0 , \3275_b1 , \3275_b0 , \3276_b1 , \3276_b0 , 
		\3277_b1 , \3277_b0 , \3278_b1 , \3278_b0 , \3279_b1 , \3279_b0 , \3280_b1 , \3280_b0 , \3281_b1 , \3281_b0 , 
		\3282_b1 , \3282_b0 , \3283_b1 , \3283_b0 , \3284_b1 , \3284_b0 , \3285_b1 , \3285_b0 , \3286_b1 , \3286_b0 , 
		\3287_b1 , \3287_b0 , \3288_b1 , \3288_b0 , \3289_b1 , \3289_b0 , \3290_b1 , \3290_b0 , \3291_b1 , \3291_b0 , 
		\3292_b1 , \3292_b0 , \3293_b1 , \3293_b0 , \3294_b1 , \3294_b0 , \3295_b1 , \3295_b0 , \3296_b1 , \3296_b0 , 
		\3297_b1 , \3297_b0 , \3298_b1 , \3298_b0 , \3299_b1 , \3299_b0 , \3300_b1 , \3300_b0 , \3301_b1 , \3301_b0 , 
		\3302_b1 , \3302_b0 , \3303_b1 , \3303_b0 , \3304_b1 , \3304_b0 , \3305_b1 , \3305_b0 , \3306_b1 , \3306_b0 , 
		\3307_b1 , \3307_b0 , \3308_b1 , \3308_b0 , \3309_b1 , \3309_b0 , \3310_b1 , \3310_b0 , \3311_b1 , \3311_b0 , 
		\3312_b1 , \3312_b0 , \3313_b1 , \3313_b0 , \3314_b1 , \3314_b0 , \3315_b1 , \3315_b0 , \3316_b1 , \3316_b0 , 
		\3317_b1 , \3317_b0 , \3318_b1 , \3318_b0 , \3319_b1 , \3319_b0 , \3320_b1 , \3320_b0 , \3321_b1 , \3321_b0 , 
		\3322_b1 , \3322_b0 , \3323_b1 , \3323_b0 , \3324_b1 , \3324_b0 , \3325_b1 , \3325_b0 , \3326_b1 , \3326_b0 , 
		\3327_b1 , \3327_b0 , \3328_b1 , \3328_b0 , \3329_b1 , \3329_b0 , \3330_b1 , \3330_b0 , \3331_b1 , \3331_b0 , 
		\3332_b1 , \3332_b0 , \3333_b1 , \3333_b0 , \3334_b1 , \3334_b0 , \3335_b1 , \3335_b0 , \3336_b1 , \3336_b0 , 
		\3337_b1 , \3337_b0 , \3338_b1 , \3338_b0 , \3339_b1 , \3339_b0 , \3340_b1 , \3340_b0 , \3341_b1 , \3341_b0 , 
		\3342_b1 , \3342_b0 , \3343_b1 , \3343_b0 , \3344_b1 , \3344_b0 , \3345_b1 , \3345_b0 , \3346_b1 , \3346_b0 , 
		\3347_b1 , \3347_b0 , \3348_b1 , \3348_b0 , \3349_b1 , \3349_b0 , \3350_b1 , \3350_b0 , \3351_b1 , \3351_b0 , 
		\3352_b1 , \3352_b0 , \3353_b1 , \3353_b0 , \3354_b1 , \3354_b0 , \3355_b1 , \3355_b0 , \3356_b1 , \3356_b0 , 
		\3357_b1 , \3357_b0 , \3358_b1 , \3358_b0 , \3359_b1 , \3359_b0 , \3360_b1 , \3360_b0 , \3361_b1 , \3361_b0 , 
		\3362_b1 , \3362_b0 , \3363_b1 , \3363_b0 , \3364_b1 , \3364_b0 , \3365_b1 , \3365_b0 , \3366_b1 , \3366_b0 , 
		\3367_b1 , \3367_b0 , \3368_b1 , \3368_b0 , \3369_b1 , \3369_b0 , \3370_b1 , \3370_b0 , \3371_b1 , \3371_b0 , 
		\3372_b1 , \3372_b0 , \3373_b1 , \3373_b0 , \3374_b1 , \3374_b0 , \3375_b1 , \3375_b0 , \3376_b1 , \3376_b0 , 
		\3377_b1 , \3377_b0 , \3378_b1 , \3378_b0 , \3379_b1 , \3379_b0 , \3380_b1 , \3380_b0 , \3381_b1 , \3381_b0 , 
		\3382_b1 , \3382_b0 , \3383_b1 , \3383_b0 , \3384_b1 , \3384_b0 , \3385_b1 , \3385_b0 , \3386_b1 , \3386_b0 , 
		\3387_b1 , \3387_b0 , \3388_b1 , \3388_b0 , \3389_b1 , \3389_b0 , \3390_b1 , \3390_b0 , \3391_b1 , \3391_b0 , 
		\3392_b1 , \3392_b0 , \3393_b1 , \3393_b0 , \3394_b1 , \3394_b0 , \3395_b1 , \3395_b0 , \3396_b1 , \3396_b0 , 
		\3397_b1 , \3397_b0 , \3398_b1 , \3398_b0 , \3399_b1 , \3399_b0 , \3400_b1 , \3400_b0 , \3401_b1 , \3401_b0 , 
		\3402_b1 , \3402_b0 , \3403_b1 , \3403_b0 , \3404_b1 , \3404_b0 , \3405_b1 , \3405_b0 , \3406_b1 , \3406_b0 , 
		\3407_b1 , \3407_b0 , \3408_b1 , \3408_b0 , \3409_b1 , \3409_b0 , \3410_b1 , \3410_b0 , \3411_b1 , \3411_b0 , 
		\3412_b1 , \3412_b0 , \3413_b1 , \3413_b0 , \3414_b1 , \3414_b0 , \3415_b1 , \3415_b0 , \3416_b1 , \3416_b0 , 
		\3417_b1 , \3417_b0 , \3418_b1 , \3418_b0 , \3419_b1 , \3419_b0 , \3420_b1 , \3420_b0 , \3421_b1 , \3421_b0 , 
		\3422_b1 , \3422_b0 , \3423_b1 , \3423_b0 , \3424_b1 , \3424_b0 , \3425_b1 , \3425_b0 , \3426_b1 , \3426_b0 , 
		\3427_b1 , \3427_b0 , \3428_b1 , \3428_b0 , \3429_b1 , \3429_b0 , \3430_b1 , \3430_b0 , \3431_b1 , \3431_b0 , 
		\3432_b1 , \3432_b0 , \3433_b1 , \3433_b0 , \3434_b1 , \3434_b0 , \3435_b1 , \3435_b0 , \3436_b1 , \3436_b0 , 
		\3437_b1 , \3437_b0 , \3438_b1 , \3438_b0 , \3439_b1 , \3439_b0 , \3440_b1 , \3440_b0 , \3441_b1 , \3441_b0 , 
		\3442_b1 , \3442_b0 , \3443_b1 , \3443_b0 , \3444_b1 , \3444_b0 , \3445_b1 , \3445_b0 , \3446_b1 , \3446_b0 , 
		\3447_b1 , \3447_b0 , \3448_b1 , \3448_b0 , \3449_b1 , \3449_b0 , \3450_b1 , \3450_b0 , \3451_b1 , \3451_b0 , 
		\3452_b1 , \3452_b0 , \3453_b1 , \3453_b0 , \3454_b1 , \3454_b0 , \3455_b1 , \3455_b0 , \3456_b1 , \3456_b0 , 
		\3457_b1 , \3457_b0 , \3458_b1 , \3458_b0 , \3459_b1 , \3459_b0 , \3460_b1 , \3460_b0 , \3461_b1 , \3461_b0 , 
		\3462_b1 , \3462_b0 , \3463_b1 , \3463_b0 , \3464_b1 , \3464_b0 , \3465_b1 , \3465_b0 , \3466_b1 , \3466_b0 , 
		\3467_b1 , \3467_b0 , \3468_b1 , \3468_b0 , \3469_b1 , \3469_b0 , \3470_b1 , \3470_b0 , \3471_b1 , \3471_b0 , 
		\3472_b1 , \3472_b0 , \3473_b1 , \3473_b0 , \3474_b1 , \3474_b0 , \3475_b1 , \3475_b0 , \3476_b1 , \3476_b0 , 
		\3477_b1 , \3477_b0 , \3478_b1 , \3478_b0 , \3479_b1 , \3479_b0 , \3480_b1 , \3480_b0 , \3481_b1 , \3481_b0 , 
		\3482_b1 , \3482_b0 , \3483_b1 , \3483_b0 , \3484_b1 , \3484_b0 , \3485_b1 , \3485_b0 , \3486_b1 , \3486_b0 , 
		\3487_b1 , \3487_b0 , \3488_b1 , \3488_b0 , \3489_b1 , \3489_b0 , \3490_b1 , \3490_b0 , \3491_b1 , \3491_b0 , 
		\3492_b1 , \3492_b0 , \3493_b1 , \3493_b0 , \3494_b1 , \3494_b0 , \3495_b1 , \3495_b0 , \3496_b1 , \3496_b0 , 
		\3497_b1 , \3497_b0 , \3498_b1 , \3498_b0 , \3499_b1 , \3499_b0 , \3500_b1 , \3500_b0 , \3501_b1 , \3501_b0 , 
		\3502_b1 , \3502_b0 , \3503_b1 , \3503_b0 , \3504_b1 , \3504_b0 , \3505_b1 , \3505_b0 , \3506_b1 , \3506_b0 , 
		\3507_b1 , \3507_b0 , \3508_b1 , \3508_b0 , \3509_b1 , \3509_b0 , \3510_b1 , \3510_b0 , \3511_b1 , \3511_b0 , 
		\3512_b1 , \3512_b0 , \3513_b1 , \3513_b0 , \3514_b1 , \3514_b0 , \3515_b1 , \3515_b0 , \3516_b1 , \3516_b0 , 
		\3517_b1 , \3517_b0 , \3518_b1 , \3518_b0 , \3519_b1 , \3519_b0 , \3520_b1 , \3520_b0 , \3521_b1 , \3521_b0 , 
		\3522_b1 , \3522_b0 , \3523_b1 , \3523_b0 , \3524_b1 , \3524_b0 , \3525_b1 , \3525_b0 , \3526_b1 , \3526_b0 , 
		\3527_b1 , \3527_b0 , \3528_b1 , \3528_b0 , \3529_b1 , \3529_b0 , \3530_b1 , \3530_b0 , \3531_b1 , \3531_b0 , 
		\3532_b1 , \3532_b0 , \3533_b1 , \3533_b0 , \3534_b1 , \3534_b0 , \3535_b1 , \3535_b0 , \3536_b1 , \3536_b0 , 
		\3537_b1 , \3537_b0 , \3538_b1 , \3538_b0 , \3539_b1 , \3539_b0 , \3540_b1 , \3540_b0 , \3541_b1 , \3541_b0 , 
		\3542_b1 , \3542_b0 , \3543_b1 , \3543_b0 , \3544_b1 , \3544_b0 , \3545_b1 , \3545_b0 , \3546_b1 , \3546_b0 , 
		\3547_b1 , \3547_b0 , \3548_b1 , \3548_b0 , \3549_b1 , \3549_b0 , \3550_b1 , \3550_b0 , \3551_b1 , \3551_b0 , 
		\3552_b1 , \3552_b0 , \3553_b1 , \3553_b0 , \3554_b1 , \3554_b0 , \3555_b1 , \3555_b0 , \3556_b1 , \3556_b0 , 
		\3557_b1 , \3557_b0 , \3558_b1 , \3558_b0 , \3559_b1 , \3559_b0 , \3560_b1 , \3560_b0 , \3561_b1 , \3561_b0 , 
		\3562_b1 , \3562_b0 , \3563_b1 , \3563_b0 , \3564_b1 , \3564_b0 , \3565_b1 , \3565_b0 , \3566_b1 , \3566_b0 , 
		\3567_b1 , \3567_b0 , \3568_b1 , \3568_b0 , \3569_b1 , \3569_b0 , \3570_b1 , \3570_b0 , \3571_b1 , \3571_b0 , 
		\3572_b1 , \3572_b0 , \3573_b1 , \3573_b0 , \3574_b1 , \3574_b0 , \3575_b1 , \3575_b0 , \3576_b1 , \3576_b0 , 
		\3577_b1 , \3577_b0 , \3578_b1 , \3578_b0 , \3579_b1 , \3579_b0 , \3580_b1 , \3580_b0 , \3581_b1 , \3581_b0 , 
		\3582_b1 , \3582_b0 , \3583_b1 , \3583_b0 , \3584_b1 , \3584_b0 , \3585_b1 , \3585_b0 , \3586_b1 , \3586_b0 , 
		\3587_b1 , \3587_b0 , \3588_b1 , \3588_b0 , \3589_b1 , \3589_b0 , \3590_b1 , \3590_b0 , \3591_b1 , \3591_b0 , 
		\3592_b1 , \3592_b0 , \3593_b1 , \3593_b0 , \3594_b1 , \3594_b0 , \3595_b1 , \3595_b0 , \3596_b1 , \3596_b0 , 
		\3597_b1 , \3597_b0 , \3598_b1 , \3598_b0 , \3599_b1 , \3599_b0 , \3600_b1 , \3600_b0 , \3601_b1 , \3601_b0 , 
		\3602_b1 , \3602_b0 , \3603_b1 , \3603_b0 , \3604_b1 , \3604_b0 , \3605_b1 , \3605_b0 , \3606_b1 , \3606_b0 , 
		\3607_b1 , \3607_b0 , \3608_b1 , \3608_b0 , \3609_b1 , \3609_b0 , \3610_b1 , \3610_b0 , \3611_b1 , \3611_b0 , 
		\3612_b1 , \3612_b0 , \3613_b1 , \3613_b0 , \3614_b1 , \3614_b0 , \3615_b1 , \3615_b0 , \3616_b1 , \3616_b0 , 
		\3617_b1 , \3617_b0 , \3618_b1 , \3618_b0 , \3619_b1 , \3619_b0 , \3620_b1 , \3620_b0 , \3621_b1 , \3621_b0 , 
		\3622_b1 , \3622_b0 , \3623_b1 , \3623_b0 , \3624_b1 , \3624_b0 , \3625_b1 , \3625_b0 , \3626_b1 , \3626_b0 , 
		\3627_b1 , \3627_b0 , \3628_b1 , \3628_b0 , \3629_b1 , \3629_b0 , \3630_b1 , \3630_b0 , \3631_b1 , \3631_b0 , 
		\3632_b1 , \3632_b0 , \3633_b1 , \3633_b0 , \3634_b1 , \3634_b0 , \3635_b1 , \3635_b0 , \3636_b1 , \3636_b0 , 
		\3637_b1 , \3637_b0 , \3638_b1 , \3638_b0 , \3639_b1 , \3639_b0 , \3640_b1 , \3640_b0 , \3641_b1 , \3641_b0 , 
		\3642_b1 , \3642_b0 , \3643_b1 , \3643_b0 , \3644_b1 , \3644_b0 , \3645_b1 , \3645_b0 , \3646_b1 , \3646_b0 , 
		\3647_b1 , \3647_b0 , \3648_b1 , \3648_b0 , \3649_b1 , \3649_b0 , \3650_b1 , \3650_b0 , \3651_b1 , \3651_b0 , 
		\3652_b1 , \3652_b0 , \3653_b1 , \3653_b0 , \3654_b1 , \3654_b0 , \3655_b1 , \3655_b0 , \3656_b1 , \3656_b0 , 
		\3657_b1 , \3657_b0 , \3658_b1 , \3658_b0 , \3659_b1 , \3659_b0 , \3660_b1 , \3660_b0 , \3661_b1 , \3661_b0 , 
		\3662_b1 , \3662_b0 , \3663_b1 , \3663_b0 , \3664_b1 , \3664_b0 , \3665_b1 , \3665_b0 , \3666_b1 , \3666_b0 , 
		\3667_b1 , \3667_b0 , \3668_b1 , \3668_b0 , \3669_b1 , \3669_b0 , \3670_b1 , \3670_b0 , \3671_b1 , \3671_b0 , 
		\3672_b1 , \3672_b0 , \3673_b1 , \3673_b0 , \3674_b1 , \3674_b0 , \3675_b1 , \3675_b0 , \3676_b1 , \3676_b0 , 
		\3677_b1 , \3677_b0 , \3678_b1 , \3678_b0 , \3679_b1 , \3679_b0 , \3680_b1 , \3680_b0 , \3681_b1 , \3681_b0 , 
		\3682_b1 , \3682_b0 , \3683_b1 , \3683_b0 , \3684_b1 , \3684_b0 , \3685_b1 , \3685_b0 , \3686_b1 , \3686_b0 , 
		\3687_b1 , \3687_b0 , \3688_b1 , \3688_b0 , \3689_b1 , \3689_b0 , \3690_b1 , \3690_b0 , \3691_b1 , \3691_b0 , 
		\3692_b1 , \3692_b0 , \3693_b1 , \3693_b0 , \3694_b1 , \3694_b0 , \3695_b1 , \3695_b0 , \3696_b1 , \3696_b0 , 
		\3697_b1 , \3697_b0 , \3698_b1 , \3698_b0 , \3699_b1 , \3699_b0 , \3700_b1 , \3700_b0 , \3701_b1 , \3701_b0 , 
		\3702_b1 , \3702_b0 , \3703_b1 , \3703_b0 , \3704_b1 , \3704_b0 , \3705_b1 , \3705_b0 , \3706_b1 , \3706_b0 , 
		\3707_b1 , \3707_b0 , \3708_b1 , \3708_b0 , \3709_b1 , \3709_b0 , \3710_b1 , \3710_b0 , \3711_b1 , \3711_b0 , 
		\3712_b1 , \3712_b0 , \3713_b1 , \3713_b0 , \3714_b1 , \3714_b0 , \3715_b1 , \3715_b0 , \3716_b1 , \3716_b0 , 
		\3717_b1 , \3717_b0 , \3718_b1 , \3718_b0 , \3719_b1 , \3719_b0 , \3720_b1 , \3720_b0 , \3721_b1 , \3721_b0 , 
		\3722_b1 , \3722_b0 , \3723_b1 , \3723_b0 , \3724_b1 , \3724_b0 , \3725_b1 , \3725_b0 , \3726_b1 , \3726_b0 , 
		\3727_b1 , \3727_b0 , \3728_b1 , \3728_b0 , \3729_b1 , \3729_b0 , \3730_b1 , \3730_b0 , \3731_b1 , \3731_b0 , 
		\3732_b1 , \3732_b0 , \3733_b1 , \3733_b0 , \3734_b1 , \3734_b0 , \3735_b1 , \3735_b0 , \3736_b1 , \3736_b0 , 
		\3737_b1 , \3737_b0 , \3738_b1 , \3738_b0 , \3739_b1 , \3739_b0 , \3740_b1 , \3740_b0 , \3741_b1 , \3741_b0 , 
		\3742_b1 , \3742_b0 , \3743_b1 , \3743_b0 , \3744_b1 , \3744_b0 , \3745_b1 , \3745_b0 , \3746_b1 , \3746_b0 , 
		\3747_b1 , \3747_b0 , \3748_b1 , \3748_b0 , \3749_b1 , \3749_b0 , \3750_b1 , \3750_b0 , \3751_b1 , \3751_b0 , 
		\3752_b1 , \3752_b0 , \3753_b1 , \3753_b0 , \3754_b1 , \3754_b0 , \3755_b1 , \3755_b0 , \3756_b1 , \3756_b0 , 
		\3757_b1 , \3757_b0 , \3758_b1 , \3758_b0 , \3759_b1 , \3759_b0 , \3760_b1 , \3760_b0 , \3761_b1 , \3761_b0 , 
		\3762_b1 , \3762_b0 , \3763_b1 , \3763_b0 , \3764_b1 , \3764_b0 , \3765_b1 , \3765_b0 , \3766_b1 , \3766_b0 , 
		\3767_b1 , \3767_b0 , \3768_b1 , \3768_b0 , \3769_b1 , \3769_b0 , \3770_b1 , \3770_b0 , \3771_b1 , \3771_b0 , 
		\3772_b1 , \3772_b0 , \3773_b1 , \3773_b0 , \3774_b1 , \3774_b0 , \3775_b1 , \3775_b0 , \3776_b1 , \3776_b0 , 
		\3777_b1 , \3777_b0 , \3778_b1 , \3778_b0 , \3779_b1 , \3779_b0 , \3780_b1 , \3780_b0 , \3781_b1 , \3781_b0 , 
		\3782_b1 , \3782_b0 , \3783_b1 , \3783_b0 , \3784_b1 , \3784_b0 , \3785_b1 , \3785_b0 , \3786_b1 , \3786_b0 , 
		\3787_b1 , \3787_b0 , \3788_b1 , \3788_b0 , \3789_b1 , \3789_b0 , \3790_b1 , \3790_b0 , \3791_b1 , \3791_b0 , 
		\3792_b1 , \3792_b0 , \3793_b1 , \3793_b0 , \3794_b1 , \3794_b0 , \3795_b1 , \3795_b0 , \3796_b1 , \3796_b0 , 
		\3797_b1 , \3797_b0 , \3798_b1 , \3798_b0 , \3799_b1 , \3799_b0 , \3800_b1 , \3800_b0 , \3801_b1 , \3801_b0 , 
		\3802_b1 , \3802_b0 , \3803_b1 , \3803_b0 , \3804_b1 , \3804_b0 , \3805_b1 , \3805_b0 , \3806_b1 , \3806_b0 , 
		\3807_b1 , \3807_b0 , \3808_b1 , \3808_b0 , \3809_b1 , \3809_b0 , \3810_b1 , \3810_b0 , \3811_b1 , \3811_b0 , 
		\3812_b1 , \3812_b0 , \3813_b1 , \3813_b0 , \3814_b1 , \3814_b0 , \3815_b1 , \3815_b0 , \3816_b1 , \3816_b0 , 
		\3817_b1 , \3817_b0 , \3818_b1 , \3818_b0 , \3819_b1 , \3819_b0 , \3820_b1 , \3820_b0 , \3821_b1 , \3821_b0 , 
		\3822_b1 , \3822_b0 , \3823_b1 , \3823_b0 , \3824_b1 , \3824_b0 , \3825_b1 , \3825_b0 , \3826_b1 , \3826_b0 , 
		\3827_b1 , \3827_b0 , \3828_b1 , \3828_b0 , \3829_b1 , \3829_b0 , \3830_b1 , \3830_b0 , \3831_b1 , \3831_b0 , 
		\3832_b1 , \3832_b0 , \3833_b1 , \3833_b0 , \3834_b1 , \3834_b0 , \3835_b1 , \3835_b0 , \3836_b1 , \3836_b0 , 
		\3837_b1 , \3837_b0 , \3838_b1 , \3838_b0 , \3839_b1 , \3839_b0 , \3840_b1 , \3840_b0 , \3841_b1 , \3841_b0 , 
		\3842_b1 , \3842_b0 , \3843_b1 , \3843_b0 , \3844_b1 , \3844_b0 , \3845_b1 , \3845_b0 , \3846_b1 , \3846_b0 , 
		\3847_b1 , \3847_b0 , \3848_b1 , \3848_b0 , \3849_b1 , \3849_b0 , \3850_b1 , \3850_b0 , \3851_b1 , \3851_b0 , 
		\3852_b1 , \3852_b0 , \3853_b1 , \3853_b0 , \3854_b1 , \3854_b0 , \3855_b1 , \3855_b0 , \3856_b1 , \3856_b0 , 
		\3857_b1 , \3857_b0 , \3858_b1 , \3858_b0 , \3859_b1 , \3859_b0 , \3860_b1 , \3860_b0 , \3861_b1 , \3861_b0 , 
		\3862_b1 , \3862_b0 , \3863_b1 , \3863_b0 , \3864_b1 , \3864_b0 , \3865_b1 , \3865_b0 , \3866_b1 , \3866_b0 , 
		\3867_b1 , \3867_b0 , \3868_b1 , \3868_b0 , \3869_b1 , \3869_b0 , \3870_b1 , \3870_b0 , \3871_b1 , \3871_b0 , 
		\3872_b1 , \3872_b0 , \3873_b1 , \3873_b0 , \3874_b1 , \3874_b0 , \3875_b1 , \3875_b0 , \3876_b1 , \3876_b0 , 
		\3877_b1 , \3877_b0 , \3878_b1 , \3878_b0 , \3879_b1 , \3879_b0 , \3880_b1 , \3880_b0 , \3881_b1 , \3881_b0 , 
		\3882_b1 , \3882_b0 , \3883_b1 , \3883_b0 , \3884_b1 , \3884_b0 , \3885_b1 , \3885_b0 , \3886_b1 , \3886_b0 , 
		\3887_b1 , \3887_b0 , \3888_b1 , \3888_b0 , \3889_b1 , \3889_b0 , \3890_b1 , \3890_b0 , \3891_b1 , \3891_b0 , 
		\3892_b1 , \3892_b0 , \3893_b1 , \3893_b0 , \3894_b1 , \3894_b0 , \3895_b1 , \3895_b0 , \3896_b1 , \3896_b0 , 
		\3897_b1 , \3897_b0 , \3898_b1 , \3898_b0 , \3899_b1 , \3899_b0 , \3900_b1 , \3900_b0 , \3901_b1 , \3901_b0 , 
		\3902_b1 , \3902_b0 , \3903_b1 , \3903_b0 , \3904_b1 , \3904_b0 , \3905_b1 , \3905_b0 , \3906_b1 , \3906_b0 , 
		\3907_b1 , \3907_b0 , \3908_b1 , \3908_b0 , \3909_b1 , \3909_b0 , \3910_b1 , \3910_b0 , \3911_b1 , \3911_b0 , 
		\3912_b1 , \3912_b0 , \3913_b1 , \3913_b0 , \3914_b1 , \3914_b0 , \3915_b1 , \3915_b0 , \3916_b1 , \3916_b0 , 
		\3917_b1 , \3917_b0 , \3918_b1 , \3918_b0 , \3919_b1 , \3919_b0 , \3920_b1 , \3920_b0 , \3921_b1 , \3921_b0 , 
		\3922_b1 , \3922_b0 , \3923_b1 , \3923_b0 , \3924_b1 , \3924_b0 , \3925_b1 , \3925_b0 , \3926_b1 , \3926_b0 , 
		\3927_b1 , \3927_b0 , \3928_b1 , \3928_b0 , \3929_b1 , \3929_b0 , \3930_b1 , \3930_b0 , \3931_b1 , \3931_b0 , 
		\3932_b1 , \3932_b0 , \3933_b1 , \3933_b0 , \3934_b1 , \3934_b0 , \3935_b1 , \3935_b0 , \3936_b1 , \3936_b0 , 
		\3937_b1 , \3937_b0 , \3938_b1 , \3938_b0 , \3939_b1 , \3939_b0 , \3940_b1 , \3940_b0 , \3941_b1 , \3941_b0 , 
		\3942_b1 , \3942_b0 , \3943_b1 , \3943_b0 , \3944_b1 , \3944_b0 , \3945_b1 , \3945_b0 , \3946_b1 , \3946_b0 , 
		\3947_b1 , \3947_b0 , \3948_b1 , \3948_b0 , \3949_b1 , \3949_b0 , \3950_b1 , \3950_b0 , \3951_b1 , \3951_b0 , 
		\3952_b1 , \3952_b0 , \3953_b1 , \3953_b0 , \3954_b1 , \3954_b0 , \3955_b1 , \3955_b0 , \3956_b1 , \3956_b0 , 
		\3957_b1 , \3957_b0 , \3958_b1 , \3958_b0 , \3959_b1 , \3959_b0 , \3960_b1 , \3960_b0 , \3961_b1 , \3961_b0 , 
		\3962_b1 , \3962_b0 , \3963_b1 , \3963_b0 , \3964_b1 , \3964_b0 , \3965_b1 , \3965_b0 , \3966_b1 , \3966_b0 , 
		\3967_b1 , \3967_b0 , \3968_b1 , \3968_b0 , \3969_b1 , \3969_b0 , \3970_b1 , \3970_b0 , \3971_b1 , \3971_b0 , 
		\3972_b1 , \3972_b0 , \3973_b1 , \3973_b0 , \3974_b1 , \3974_b0 , \3975_b1 , \3975_b0 , \3976_b1 , \3976_b0 , 
		\3977_b1 , \3977_b0 , \3978_b1 , \3978_b0 , \3979_b1 , \3979_b0 , \3980_b1 , \3980_b0 , \3981_b1 , \3981_b0 , 
		\3982_b1 , \3982_b0 , \3983_b1 , \3983_b0 , \3984_b1 , \3984_b0 , \3985_b1 , \3985_b0 , \3986_b1 , \3986_b0 , 
		\3987_b1 , \3987_b0 , \3988_b1 , \3988_b0 , \3989_b1 , \3989_b0 , \3990_b1 , \3990_b0 , \3991_b1 , \3991_b0 , 
		\3992_b1 , \3992_b0 , \3993_b1 , \3993_b0 , \3994_b1 , \3994_b0 , \3995_b1 , \3995_b0 , \3996_b1 , \3996_b0 , 
		\3997_b1 , \3997_b0 , \3998_b1 , \3998_b0 , \3999_b1 , \3999_b0 , \4000_b1 , \4000_b0 , \4001_b1 , \4001_b0 , 
		\4002_b1 , \4002_b0 , \4003_b1 , \4003_b0 , \4004_b1 , \4004_b0 , \4005_b1 , \4005_b0 , \4006_b1 , \4006_b0 , 
		\4007_b1 , \4007_b0 , \4008_b1 , \4008_b0 , \4009_b1 , \4009_b0 , \4010_b1 , \4010_b0 , \4011_b1 , \4011_b0 , 
		\4012_b1 , \4012_b0 , \4013_b1 , \4013_b0 , \4014_b1 , \4014_b0 , \4015_b1 , \4015_b0 , \4016_b1 , \4016_b0 , 
		\4017_b1 , \4017_b0 , \4018_b1 , \4018_b0 , \4019_b1 , \4019_b0 , \4020_b1 , \4020_b0 , \4021_b1 , \4021_b0 , 
		\4022_b1 , \4022_b0 , \4023_b1 , \4023_b0 , \4024_b1 , \4024_b0 , \4025_b1 , \4025_b0 , \4026_b1 , \4026_b0 , 
		\4027_b1 , \4027_b0 , \4028_b1 , \4028_b0 , \4029_b1 , \4029_b0 , \4030_b1 , \4030_b0 , \4031_b1 , \4031_b0 , 
		\4032_b1 , \4032_b0 , \4033_b1 , \4033_b0 , \4034_b1 , \4034_b0 , \4035_b1 , \4035_b0 , \4036_b1 , \4036_b0 , 
		\4037_b1 , \4037_b0 , \4038_b1 , \4038_b0 , \4039_b1 , \4039_b0 , \4040_b1 , \4040_b0 , \4041_b1 , \4041_b0 , 
		\4042_b1 , \4042_b0 , \4043_b1 , \4043_b0 , \4044_b1 , \4044_b0 , \4045_b1 , \4045_b0 , \4046_b1 , \4046_b0 , 
		\4047_b1 , \4047_b0 , \4048_b1 , \4048_b0 , \4049_b1 , \4049_b0 , \4050_b1 , \4050_b0 , \4051_b1 , \4051_b0 , 
		\4052_b1 , \4052_b0 , \4053_b1 , \4053_b0 , \4054_b1 , \4054_b0 , \4055_b1 , \4055_b0 , \4056_b1 , \4056_b0 , 
		\4057_b1 , \4057_b0 , \4058_b1 , \4058_b0 , \4059_b1 , \4059_b0 , \4060_b1 , \4060_b0 , \4061_b1 , \4061_b0 , 
		\4062_b1 , \4062_b0 , \4063_b1 , \4063_b0 , \4064_b1 , \4064_b0 , \4065_b1 , \4065_b0 , \4066_b1 , \4066_b0 , 
		\4067_b1 , \4067_b0 , \4068_b1 , \4068_b0 , \4069_b1 , \4069_b0 , \4070_b1 , \4070_b0 , \4071_b1 , \4071_b0 , 
		\4072_b1 , \4072_b0 , \4073_b1 , \4073_b0 , \4074_b1 , \4074_b0 , \4075_b1 , \4075_b0 , \4076_b1 , \4076_b0 , 
		\4077_b1 , \4077_b0 , \4078_b1 , \4078_b0 , \4079_b1 , \4079_b0 , \4080_b1 , \4080_b0 , \4081_b1 , \4081_b0 , 
		\4082_b1 , \4082_b0 , \4083_b1 , \4083_b0 , \4084_b1 , \4084_b0 , \4085_b1 , \4085_b0 , \4086_b1 , \4086_b0 , 
		\4087_b1 , \4087_b0 , \4088_b1 , \4088_b0 , \4089_b1 , \4089_b0 , \4090_b1 , \4090_b0 , \4091_b1 , \4091_b0 , 
		\4092_b1 , \4092_b0 , \4093_b1 , \4093_b0 , \4094_b1 , \4094_b0 , \4095_b1 , \4095_b0 , \4096_b1 , \4096_b0 , 
		\4097_b1 , \4097_b0 , \4098_b1 , \4098_b0 , \4099_b1 , \4099_b0 , \4100_b1 , \4100_b0 , \4101_b1 , \4101_b0 , 
		\4102_b1 , \4102_b0 , \4103_b1 , \4103_b0 , \4104_b1 , \4104_b0 , \4105_b1 , \4105_b0 , \4106_b1 , \4106_b0 , 
		\4107_b1 , \4107_b0 , \4108_b1 , \4108_b0 , \4109_b1 , \4109_b0 , \4110_b1 , \4110_b0 , \4111_b1 , \4111_b0 , 
		\4112_b1 , \4112_b0 , \4113_b1 , \4113_b0 , \4114_b1 , \4114_b0 , \4115_b1 , \4115_b0 , \4116_b1 , \4116_b0 , 
		\4117_b1 , \4117_b0 , \4118_b1 , \4118_b0 , \4119_b1 , \4119_b0 , \4120_b1 , \4120_b0 , \4121_b1 , \4121_b0 , 
		\4122_b1 , \4122_b0 , \4123_b1 , \4123_b0 , \4124_b1 , \4124_b0 , \4125_b1 , \4125_b0 , \4126_b1 , \4126_b0 , 
		\4127_b1 , \4127_b0 , \4128_b1 , \4128_b0 , \4129_b1 , \4129_b0 , \4130_b1 , \4130_b0 , \4131_b1 , \4131_b0 , 
		\4132_b1 , \4132_b0 , \4133_b1 , \4133_b0 , \4134_b1 , \4134_b0 , \4135_b1 , \4135_b0 , \4136_b1 , \4136_b0 , 
		\4137_b1 , \4137_b0 , \4138_b1 , \4138_b0 , \4139_b1 , \4139_b0 , \4140_b1 , \4140_b0 , \4141_b1 , \4141_b0 , 
		\4142_b1 , \4142_b0 , \4143_b1 , \4143_b0 , \4144_b1 , \4144_b0 , \4145_b1 , \4145_b0 , \4146_b1 , \4146_b0 , 
		\4147_b1 , \4147_b0 , \4148_b1 , \4148_b0 , \4149_b1 , \4149_b0 , \4150_b1 , \4150_b0 , \4151_b1 , \4151_b0 , 
		\4152_b1 , \4152_b0 , \4153_b1 , \4153_b0 , \4154_b1 , \4154_b0 , \4155_b1 , \4155_b0 , \4156_b1 , \4156_b0 , 
		\4157_b1 , \4157_b0 , \4158_b1 , \4158_b0 , \4159_b1 , \4159_b0 , \4160_b1 , \4160_b0 , \4161_b1 , \4161_b0 , 
		\4162_b1 , \4162_b0 , \4163_b1 , \4163_b0 , \4164_b1 , \4164_b0 , \4165_b1 , \4165_b0 , \4166_b1 , \4166_b0 , 
		\4167_b1 , \4167_b0 , \4168_b1 , \4168_b0 , \4169_b1 , \4169_b0 , \4170_b1 , \4170_b0 , \4171_b1 , \4171_b0 , 
		\4172_b1 , \4172_b0 , \4173_b1 , \4173_b0 , \4174_b1 , \4174_b0 , \4175_b1 , \4175_b0 , \4176_b1 , \4176_b0 , 
		\4177_b1 , \4177_b0 , \4178_b1 , \4178_b0 , \4179_b1 , \4179_b0 , \4180_b1 , \4180_b0 , \4181_b1 , \4181_b0 , 
		\4182_b1 , \4182_b0 , \4183_b1 , \4183_b0 , \4184_b1 , \4184_b0 , \4185_b1 , \4185_b0 , \4186_b1 , \4186_b0 , 
		\4187_b1 , \4187_b0 , \4188_b1 , \4188_b0 , \4189_b1 , \4189_b0 , \4190_b1 , \4190_b0 , \4191_b1 , \4191_b0 , 
		\4192_b1 , \4192_b0 , \4193_b1 , \4193_b0 , \4194_b1 , \4194_b0 , \4195_b1 , \4195_b0 , \4196_b1 , \4196_b0 , 
		\4197_b1 , \4197_b0 , \4198_b1 , \4198_b0 , \4199_b1 , \4199_b0 , \4200_b1 , \4200_b0 , \4201_b1 , \4201_b0 , 
		\4202_b1 , \4202_b0 , \4203_b1 , \4203_b0 , \4204_b1 , \4204_b0 , \4205_b1 , \4205_b0 , \4206_b1 , \4206_b0 , 
		\4207_b1 , \4207_b0 , \4208_b1 , \4208_b0 , \4209_b1 , \4209_b0 , \4210_b1 , \4210_b0 , \4211_b1 , \4211_b0 , 
		\4212_b1 , \4212_b0 , \4213_b1 , \4213_b0 , \4214_b1 , \4214_b0 , \4215_b1 , \4215_b0 , \4216_b1 , \4216_b0 , 
		\4217_b1 , \4217_b0 , \4218_b1 , \4218_b0 , \4219_b1 , \4219_b0 , \4220_b1 , \4220_b0 , \4221_b1 , \4221_b0 , 
		\4222_b1 , \4222_b0 , \4223_b1 , \4223_b0 , \4224_b1 , \4224_b0 , \4225_b1 , \4225_b0 , \4226_b1 , \4226_b0 , 
		\4227_b1 , \4227_b0 , \4228_b1 , \4228_b0 , \4229_b1 , \4229_b0 , \4230_b1 , \4230_b0 , \4231_b1 , \4231_b0 , 
		\4232_b1 , \4232_b0 , \4233_b1 , \4233_b0 , \4234_b1 , \4234_b0 , \4235_b1 , \4235_b0 , \4236_b1 , \4236_b0 , 
		\4237_b1 , \4237_b0 , \4238_b1 , \4238_b0 , \4239_b1 , \4239_b0 , \4240_b1 , \4240_b0 , \4241_b1 , \4241_b0 , 
		\4242_b1 , \4242_b0 , \4243_b1 , \4243_b0 , \4244_b1 , \4244_b0 , \4245_b1 , \4245_b0 , \4246_b1 , \4246_b0 , 
		\4247_b1 , \4247_b0 , \4248_b1 , \4248_b0 , \4249_b1 , \4249_b0 , \4250_b1 , \4250_b0 , \4251_b1 , \4251_b0 , 
		\4252_b1 , \4252_b0 , \4253_b1 , \4253_b0 , \4254_b1 , \4254_b0 , \4255_b1 , \4255_b0 , \4256_b1 , \4256_b0 , 
		\4257_b1 , \4257_b0 , \4258_b1 , \4258_b0 , \4259_b1 , \4259_b0 , \4260_b1 , \4260_b0 , \4261_b1 , \4261_b0 , 
		\4262_b1 , \4262_b0 , \4263_b1 , \4263_b0 , \4264_b1 , \4264_b0 , \4265_b1 , \4265_b0 , \4266_b1 , \4266_b0 , 
		\4267_b1 , \4267_b0 , \4268_b1 , \4268_b0 , \4269_b1 , \4269_b0 , \4270_b1 , \4270_b0 , \4271_b1 , \4271_b0 , 
		\4272_b1 , \4272_b0 , \4273_b1 , \4273_b0 , \4274_b1 , \4274_b0 , \4275_b1 , \4275_b0 , \4276_b1 , \4276_b0 , 
		\4277_b1 , \4277_b0 , \4278_b1 , \4278_b0 , \4279_b1 , \4279_b0 , \4280_b1 , \4280_b0 , \4281_b1 , \4281_b0 , 
		\4282_b1 , \4282_b0 , \4283_b1 , \4283_b0 , \4284_b1 , \4284_b0 , \4285_b1 , \4285_b0 , \4286_b1 , \4286_b0 , 
		\4287_b1 , \4287_b0 , \4288_b1 , \4288_b0 , \4289_b1 , \4289_b0 , \4290_b1 , \4290_b0 , \4291_b1 , \4291_b0 , 
		\4292_b1 , \4292_b0 , \4293_b1 , \4293_b0 , \4294_b1 , \4294_b0 , \4295_b1 , \4295_b0 , \4296_b1 , \4296_b0 , 
		\4297_b1 , \4297_b0 , \4298_b1 , \4298_b0 , \4299_b1 , \4299_b0 , \4300_b1 , \4300_b0 , \4301_b1 , \4301_b0 , 
		\4302_b1 , \4302_b0 , \4303_b1 , \4303_b0 , \4304_b1 , \4304_b0 , \4305_b1 , \4305_b0 , \4306_b1 , \4306_b0 , 
		\4307_b1 , \4307_b0 , \4308_b1 , \4308_b0 , \4309_b1 , \4309_b0 , \4310_b1 , \4310_b0 , \4311_b1 , \4311_b0 , 
		\4312_b1 , \4312_b0 , \4313_b1 , \4313_b0 , \4314_b1 , \4314_b0 , \4315_b1 , \4315_b0 , \4316_b1 , \4316_b0 , 
		\4317_b1 , \4317_b0 , \4318_b1 , \4318_b0 , \4319_b1 , \4319_b0 , \4320_b1 , \4320_b0 , \4321_b1 , \4321_b0 , 
		\4322_b1 , \4322_b0 , \4323_b1 , \4323_b0 , \4324_b1 , \4324_b0 , \4325_b1 , \4325_b0 , \4326_b1 , \4326_b0 , 
		\4327_b1 , \4327_b0 , \4328_b1 , \4328_b0 , \4329_b1 , \4329_b0 , \4330_b1 , \4330_b0 , \4331_b1 , \4331_b0 , 
		\4332_b1 , \4332_b0 , \4333_b1 , \4333_b0 , \4334_b1 , \4334_b0 , \4335_b1 , \4335_b0 , \4336_b1 , \4336_b0 , 
		\4337_b1 , \4337_b0 , \4338_b1 , \4338_b0 , \4339_b1 , \4339_b0 , \4340_b1 , \4340_b0 , \4341_b1 , \4341_b0 , 
		\4342_b1 , \4342_b0 , \4343_b1 , \4343_b0 , \4344_b1 , \4344_b0 , \4345_b1 , \4345_b0 , \4346_b1 , \4346_b0 , 
		\4347_b1 , \4347_b0 , \4348_b1 , \4348_b0 , \4349_b1 , \4349_b0 , \4350_b1 , \4350_b0 , \4351_b1 , \4351_b0 , 
		\4352_b1 , \4352_b0 , \4353_b1 , \4353_b0 , \4354_b1 , \4354_b0 , \4355_b1 , \4355_b0 , \4356_b1 , \4356_b0 , 
		\4357_b1 , \4357_b0 , \4358_b1 , \4358_b0 , \4359_b1 , \4359_b0 , \4360_b1 , \4360_b0 , \4361_b1 , \4361_b0 , 
		\4362_b1 , \4362_b0 , \4363_b1 , \4363_b0 , \4364_b1 , \4364_b0 , \4365_b1 , \4365_b0 , \4366_b1 , \4366_b0 , 
		\4367_b1 , \4367_b0 , \4368_b1 , \4368_b0 , \4369_b1 , \4369_b0 , \4370_b1 , \4370_b0 , \4371_b1 , \4371_b0 , 
		\4372_b1 , \4372_b0 , \4373_b1 , \4373_b0 , \4374_b1 , \4374_b0 , \4375_b1 , \4375_b0 , \4376_b1 , \4376_b0 , 
		\4377_b1 , \4377_b0 , \4378_b1 , \4378_b0 , \4379_b1 , \4379_b0 , \4380_b1 , \4380_b0 , \4381_b1 , \4381_b0 , 
		\4382_b1 , \4382_b0 , \4383_b1 , \4383_b0 , \4384_b1 , \4384_b0 , \4385_b1 , \4385_b0 , \4386_b1 , \4386_b0 , 
		\4387_b1 , \4387_b0 , \4388_b1 , \4388_b0 , \4389_b1 , \4389_b0 , \4390_b1 , \4390_b0 , \4391_b1 , \4391_b0 , 
		\4392_b1 , \4392_b0 , \4393_b1 , \4393_b0 , \4394_b1 , \4394_b0 , \4395_b1 , \4395_b0 , \4396_b1 , \4396_b0 , 
		\4397_b1 , \4397_b0 , \4398_b1 , \4398_b0 , \4399_b1 , \4399_b0 , \4400_b1 , \4400_b0 , \4401_b1 , \4401_b0 , 
		\4402_b1 , \4402_b0 , \4403_b1 , \4403_b0 , \4404_b1 , \4404_b0 , \4405_b1 , \4405_b0 , \4406_b1 , \4406_b0 , 
		\4407_b1 , \4407_b0 , \4408_b1 , \4408_b0 , \4409_b1 , \4409_b0 , \4410_b1 , \4410_b0 , \4411_b1 , \4411_b0 , 
		\4412_b1 , \4412_b0 , \4413_b1 , \4413_b0 , \4414_b1 , \4414_b0 , \4415_b1 , \4415_b0 , \4416_b1 , \4416_b0 , 
		\4417_b1 , \4417_b0 , \4418_b1 , \4418_b0 , \4419_b1 , \4419_b0 , \4420_b1 , \4420_b0 , \4421_b1 , \4421_b0 , 
		\4422_b1 , \4422_b0 , \4423_b1 , \4423_b0 , \4424_b1 , \4424_b0 , \4425_b1 , \4425_b0 , \4426_b1 , \4426_b0 , 
		\4427_b1 , \4427_b0 , \4428_b1 , \4428_b0 , \4429_b1 , \4429_b0 , \4430_b1 , \4430_b0 , \4431_b1 , \4431_b0 , 
		\4432_b1 , \4432_b0 , \4433_b1 , \4433_b0 , \4434_b1 , \4434_b0 , \4435_b1 , \4435_b0 , \4436_b1 , \4436_b0 , 
		\4437_b1 , \4437_b0 , \4438_b1 , \4438_b0 , \4439_b1 , \4439_b0 , \4440_b1 , \4440_b0 , \4441_b1 , \4441_b0 , 
		\4442_b1 , \4442_b0 , \4443_b1 , \4443_b0 , \4444_b1 , \4444_b0 , \4445_b1 , \4445_b0 , \4446_b1 , \4446_b0 , 
		\4447_b1 , \4447_b0 , \4448_b1 , \4448_b0 , \4449_b1 , \4449_b0 , \4450_b1 , \4450_b0 , \4451_b1 , \4451_b0 , 
		\4452_b1 , \4452_b0 , \4453_b1 , \4453_b0 , \4454_b1 , \4454_b0 , \4455_b1 , \4455_b0 , \4456_b1 , \4456_b0 , 
		\4457_b1 , \4457_b0 , \4458_b1 , \4458_b0 , \4459_b1 , \4459_b0 , \4460_b1 , \4460_b0 , \4461_b1 , \4461_b0 , 
		\4462_b1 , \4462_b0 , \4463_b1 , \4463_b0 , \4464_b1 , \4464_b0 , \4465_b1 , \4465_b0 , \4466_b1 , \4466_b0 , 
		\4467_b1 , \4467_b0 , \4468_Z[31]_b1 , \4468_Z[31]_b0 , \4469_b1 , \4469_b0 , \4470_Z[30]_b1 , \4470_Z[30]_b0 , \4471_b1 , \4471_b0 , 
		\4472_Z[29]_b1 , \4472_Z[29]_b0 , \4473_b1 , \4473_b0 , \4474_Z[28]_b1 , \4474_Z[28]_b0 , \4475_b1 , \4475_b0 , \4476_Z[27]_b1 , \4476_Z[27]_b0 , 
		\4477_b1 , \4477_b0 , \4478_Z[26]_b1 , \4478_Z[26]_b0 , \4479_b1 , \4479_b0 , \4480_Z[25]_b1 , \4480_Z[25]_b0 , \4481_b1 , \4481_b0 , 
		\4482_Z[24]_b1 , \4482_Z[24]_b0 , \4483_b1 , \4483_b0 , \4484_Z[23]_b1 , \4484_Z[23]_b0 , \4485_b1 , \4485_b0 , \4486_Z[22]_b1 , \4486_Z[22]_b0 , 
		\4487_b1 , \4487_b0 , \4488_Z[21]_b1 , \4488_Z[21]_b0 , \4489_b1 , \4489_b0 , \4490_Z[20]_b1 , \4490_Z[20]_b0 , \4491_b1 , \4491_b0 , 
		\4492_Z[19]_b1 , \4492_Z[19]_b0 , \4493_b1 , \4493_b0 , \4494_Z[18]_b1 , \4494_Z[18]_b0 , \4495_b1 , \4495_b0 , \4496_Z[17]_b1 , \4496_Z[17]_b0 , 
		\4497_b1 , \4497_b0 , \4498_Z[16]_b1 , \4498_Z[16]_b0 , \4499_b1 , \4499_b0 , \4500_Z[15]_b1 , \4500_Z[15]_b0 , \4501_b1 , \4501_b0 , 
		\4502_Z[14]_b1 , \4502_Z[14]_b0 , \4503_b1 , \4503_b0 , \4504_Z[13]_b1 , \4504_Z[13]_b0 , \4505_b1 , \4505_b0 , \4506_Z[12]_b1 , \4506_Z[12]_b0 , 
		\4507_b1 , \4507_b0 , \4508_Z[11]_b1 , \4508_Z[11]_b0 , \4509_b1 , \4509_b0 , \4510_Z[10]_b1 , \4510_Z[10]_b0 , \4511_b1 , \4511_b0 , 
		\4512_Z[9]_b1 , \4512_Z[9]_b0 , \4513_b1 , \4513_b0 , \4514_Z[8]_b1 , \4514_Z[8]_b0 , \4515_b1 , \4515_b0 , \4516_Z[7]_b1 , \4516_Z[7]_b0 , 
		\4517_b1 , \4517_b0 , \4518_Z[6]_b1 , \4518_Z[6]_b0 , \4519_b1 , \4519_b0 , \4520_Z[5]_b1 , \4520_Z[5]_b0 , \4521_b1 , \4521_b0 , 
		\4522_Z[4]_b1 , \4522_Z[4]_b0 , \4523_b1 , \4523_b0 , \4524_Z[3]_b1 , \4524_Z[3]_b0 , \4525_b1 , \4525_b0 , \4526_Z[2]_b1 , \4526_Z[2]_b0 , 
		\4527_b1 , \4527_b0 , \4528_Z[1]_b1 , \4528_Z[1]_b0 , \4529_b1 , \4529_b0 , \4530_Z[0]_b1 , \4530_Z[0]_b0 , w_0 , w_1 , 
		w_2 , w_3 , w_4 , w_5 , w_6 , w_7 , w_8 , w_9 , w_10 , w_11 , 
		w_12 , w_13 , w_14 , w_15 , w_16 , w_17 , w_18 , w_19 , w_20 , w_21 , 
		w_22 , w_23 , w_24 , w_25 , w_26 , w_27 , w_28 , w_29 , w_30 , w_31 , 
		w_32 , w_33 , w_34 , w_35 , w_36 , w_37 , w_38 , w_39 , w_40 , w_41 , 
		w_42 , w_43 , w_44 , w_45 , w_46 , w_47 , w_48 , w_49 , w_50 , w_51 , 
		w_52 , w_53 , w_54 , w_55 , w_56 , w_57 , w_58 , w_59 , w_60 , w_61 , 
		w_62 , w_63 , w_64 , w_65 , w_66 , w_67 , w_68 , w_69 , w_70 , w_71 , 
		w_72 , w_73 , w_74 , w_75 , w_76 , w_77 , w_78 , w_79 , w_80 , w_81 , 
		w_82 , w_83 , w_84 , w_85 , w_86 , w_87 , w_88 , w_89 , w_90 , w_91 , 
		w_92 , w_93 , w_94 , w_95 , w_96 , w_97 , w_98 , w_99 , w_100 , w_101 , 
		w_102 , w_103 , w_104 , w_105 , w_106 , w_107 , w_108 , w_109 , w_110 , w_111 , 
		w_112 , w_113 , w_114 , w_115 , w_116 , w_117 , w_118 , w_119 , w_120 , w_121 , 
		w_122 , w_123 , w_124 , w_125 , w_126 , w_127 , w_128 , w_129 , w_130 , w_131 , 
		w_132 , w_133 , w_134 , w_135 , w_136 , w_137 , w_138 , w_139 , w_140 , w_141 , 
		w_142 , w_143 , w_144 , w_145 , w_146 , w_147 , w_148 , w_149 , w_150 , w_151 , 
		w_152 , w_153 , w_154 , w_155 , w_156 , w_157 , w_158 , w_159 , w_160 , w_161 , 
		w_162 , w_163 , w_164 , w_165 , w_166 , w_167 , w_168 , w_169 , w_170 , w_171 , 
		w_172 , w_173 , w_174 , w_175 , w_176 , w_177 , w_178 , w_179 , w_180 , w_181 , 
		w_182 , w_183 , w_184 , w_185 , w_186 , w_187 , w_188 , w_189 , w_190 , w_191 , 
		w_192 , w_193 , w_194 , w_195 , w_196 , w_197 , w_198 , w_199 , w_200 , w_201 , 
		w_202 , w_203 , w_204 , w_205 , w_206 , w_207 , w_208 , w_209 , w_210 , w_211 , 
		w_212 , w_213 , w_214 , w_215 , w_216 , w_217 , w_218 , w_219 , w_220 , w_221 , 
		w_222 , w_223 , w_224 , w_225 , w_226 , w_227 , w_228 , w_229 , w_230 , w_231 , 
		w_232 , w_233 , w_234 , w_235 , w_236 , w_237 , w_238 , w_239 , w_240 , w_241 , 
		w_242 , w_243 , w_244 , w_245 , w_246 , w_247 , w_248 , w_249 , w_250 , w_251 , 
		w_252 , w_253 , w_254 , w_255 , w_256 , w_257 , w_258 , w_259 , w_260 , w_261 , 
		w_262 , w_263 , w_264 , w_265 , w_266 , w_267 , w_268 , w_269 , w_270 , w_271 , 
		w_272 , w_273 , w_274 , w_275 , w_276 , w_277 , w_278 , w_279 , w_280 , w_281 , 
		w_282 , w_283 , w_284 , w_285 , w_286 , w_287 , w_288 , w_289 , w_290 , w_291 , 
		w_292 , w_293 , w_294 , w_295 , w_296 , w_297 , w_298 , w_299 , w_300 , w_301 , 
		w_302 , w_303 , w_304 , w_305 , w_306 , w_307 , w_308 , w_309 , w_310 , w_311 , 
		w_312 , w_313 , w_314 , w_315 , w_316 , w_317 , w_318 , w_319 , w_320 , w_321 , 
		w_322 , w_323 , w_324 , w_325 , w_326 , w_327 , w_328 , w_329 , w_330 , w_331 , 
		w_332 , w_333 , w_334 , w_335 , w_336 , w_337 , w_338 , w_339 , w_340 , w_341 , 
		w_342 , w_343 , w_344 , w_345 , w_346 , w_347 , w_348 , w_349 , w_350 , w_351 , 
		w_352 , w_353 , w_354 , w_355 , w_356 , w_357 , w_358 , w_359 , w_360 , w_361 , 
		w_362 , w_363 , w_364 , w_365 , w_366 , w_367 , w_368 , w_369 , w_370 , w_371 , 
		w_372 , w_373 , w_374 , w_375 , w_376 , w_377 , w_378 , w_379 , w_380 , w_381 , 
		w_382 , w_383 , w_384 , w_385 , w_386 , w_387 , w_388 , w_389 , w_390 , w_391 , 
		w_392 , w_393 , w_394 , w_395 , w_396 , w_397 , w_398 , w_399 , w_400 , w_401 , 
		w_402 , w_403 , w_404 , w_405 , w_406 , w_407 , w_408 , w_409 , w_410 , w_411 , 
		w_412 , w_413 , w_414 , w_415 , w_416 , w_417 , w_418 , w_419 , w_420 , w_421 , 
		w_422 , w_423 , w_424 , w_425 , w_426 , w_427 , w_428 , w_429 , w_430 , w_431 , 
		w_432 , w_433 , w_434 , w_435 , w_436 , w_437 , w_438 , w_439 , w_440 , w_441 , 
		w_442 , w_443 , w_444 , w_445 , w_446 , w_447 , w_448 , w_449 , w_450 , w_451 , 
		w_452 , w_453 , w_454 , w_455 , w_456 , w_457 , w_458 , w_459 , w_460 , w_461 , 
		w_462 , w_463 , w_464 , w_465 , w_466 , w_467 , w_468 , w_469 , w_470 , w_471 , 
		w_472 , w_473 , w_474 , w_475 , w_476 , w_477 , w_478 , w_479 , w_480 , w_481 , 
		w_482 , w_483 , w_484 , w_485 , w_486 , w_487 , w_488 , w_489 , w_490 , w_491 , 
		w_492 , w_493 , w_494 , w_495 , w_496 , w_497 , w_498 , w_499 , w_500 , w_501 , 
		w_502 , w_503 , w_504 , w_505 , w_506 , w_507 , w_508 , w_509 , w_510 , w_511 , 
		w_512 , w_513 , w_514 , w_515 , w_516 , w_517 , w_518 , w_519 , w_520 , w_521 , 
		w_522 , w_523 , w_524 , w_525 , w_526 , w_527 , w_528 , w_529 , w_530 , w_531 , 
		w_532 , w_533 , w_534 , w_535 , w_536 , w_537 , w_538 , w_539 , w_540 , w_541 , 
		w_542 , w_543 , w_544 , w_545 , w_546 , w_547 , w_548 , w_549 , w_550 , w_551 , 
		w_552 , w_553 , w_554 , w_555 , w_556 , w_557 , w_558 , w_559 , w_560 , w_561 , 
		w_562 , w_563 , w_564 , w_565 , w_566 , w_567 , w_568 , w_569 , w_570 , w_571 , 
		w_572 , w_573 , w_574 , w_575 , w_576 , w_577 , w_578 , w_579 , w_580 , w_581 , 
		w_582 , w_583 , w_584 , w_585 , w_586 , w_587 , w_588 , w_589 , w_590 , w_591 , 
		w_592 , w_593 , w_594 , w_595 , w_596 , w_597 , w_598 , w_599 , w_600 , w_601 , 
		w_602 , w_603 , w_604 , w_605 , w_606 , w_607 , w_608 , w_609 , w_610 , w_611 , 
		w_612 , w_613 , w_614 , w_615 , w_616 , w_617 , w_618 , w_619 , w_620 , w_621 , 
		w_622 , w_623 , w_624 , w_625 , w_626 , w_627 , w_628 , w_629 , w_630 , w_631 , 
		w_632 , w_633 , w_634 , w_635 , w_636 , w_637 , w_638 , w_639 , w_640 , w_641 , 
		w_642 , w_643 , w_644 , w_645 , w_646 , w_647 , w_648 , w_649 , w_650 , w_651 , 
		w_652 , w_653 , w_654 , w_655 , w_656 , w_657 , w_658 , w_659 , w_660 , w_661 , 
		w_662 , w_663 , w_664 , w_665 , w_666 , w_667 , w_668 , w_669 , w_670 , w_671 , 
		w_672 , w_673 , w_674 , w_675 , w_676 , w_677 , w_678 , w_679 , w_680 , w_681 , 
		w_682 , w_683 , w_684 , w_685 , w_686 , w_687 , w_688 , w_689 , w_690 , w_691 , 
		w_692 , w_693 , w_694 , w_695 , w_696 , w_697 , w_698 , w_699 , w_700 , w_701 , 
		w_702 , w_703 , w_704 , w_705 , w_706 , w_707 , w_708 , w_709 , w_710 , w_711 , 
		w_712 , w_713 , w_714 , w_715 , w_716 , w_717 , w_718 , w_719 , w_720 , w_721 , 
		w_722 , w_723 , w_724 , w_725 , w_726 , w_727 , w_728 , w_729 , w_730 , w_731 , 
		w_732 , w_733 , w_734 , w_735 , w_736 , w_737 , w_738 , w_739 , w_740 , w_741 , 
		w_742 , w_743 , w_744 , w_745 , w_746 , w_747 , w_748 , w_749 , w_750 , w_751 , 
		w_752 , w_753 , w_754 , w_755 , w_756 , w_757 , w_758 , w_759 , w_760 , w_761 , 
		w_762 , w_763 , w_764 , w_765 , w_766 , w_767 , w_768 , w_769 , w_770 , w_771 , 
		w_772 , w_773 , w_774 , w_775 , w_776 , w_777 , w_778 , w_779 , w_780 , w_781 , 
		w_782 , w_783 , w_784 , w_785 , w_786 , w_787 , w_788 , w_789 , w_790 , w_791 , 
		w_792 , w_793 , w_794 , w_795 , w_796 , w_797 , w_798 , w_799 , w_800 , w_801 , 
		w_802 , w_803 , w_804 , w_805 , w_806 , w_807 , w_808 , w_809 , w_810 , w_811 , 
		w_812 , w_813 , w_814 , w_815 , w_816 , w_817 , w_818 , w_819 , w_820 , w_821 , 
		w_822 , w_823 , w_824 , w_825 , w_826 , w_827 , w_828 , w_829 , w_830 , w_831 , 
		w_832 , w_833 , w_834 , w_835 , w_836 , w_837 , w_838 , w_839 , w_840 , w_841 , 
		w_842 , w_843 , w_844 , w_845 , w_846 , w_847 , w_848 , w_849 , w_850 , w_851 , 
		w_852 , w_853 , w_854 , w_855 , w_856 , w_857 , w_858 , w_859 , w_860 , w_861 , 
		w_862 , w_863 , w_864 , w_865 , w_866 , w_867 , w_868 , w_869 , w_870 , w_871 , 
		w_872 , w_873 , w_874 , w_875 , w_876 , w_877 , w_878 , w_879 , w_880 , w_881 , 
		w_882 , w_883 , w_884 , w_885 , w_886 , w_887 , w_888 , w_889 , w_890 , w_891 , 
		w_892 , w_893 , w_894 , w_895 , w_896 , w_897 , w_898 , w_899 , w_900 , w_901 , 
		w_902 , w_903 , w_904 , w_905 , w_906 , w_907 , w_908 , w_909 , w_910 , w_911 , 
		w_912 , w_913 , w_914 , w_915 , w_916 , w_917 , w_918 , w_919 , w_920 , w_921 , 
		w_922 , w_923 , w_924 , w_925 , w_926 , w_927 , w_928 , w_929 , w_930 , w_931 , 
		w_932 , w_933 , w_934 , w_935 , w_936 , w_937 , w_938 , w_939 , w_940 , w_941 , 
		w_942 , w_943 , w_944 , w_945 , w_946 , w_947 , w_948 , w_949 , w_950 , w_951 , 
		w_952 , w_953 , w_954 , w_955 , w_956 , w_957 , w_958 , w_959 , w_960 , w_961 , 
		w_962 , w_963 , w_964 , w_965 , w_966 , w_967 , w_968 , w_969 , w_970 , w_971 , 
		w_972 , w_973 , w_974 , w_975 , w_976 , w_977 , w_978 , w_979 , w_980 , w_981 , 
		w_982 , w_983 , w_984 , w_985 , w_986 , w_987 , w_988 , w_989 , w_990 , w_991 , 
		w_992 , w_993 , w_994 , w_995 , w_996 , w_997 , w_998 , w_999 , w_1000 , w_1001 , 
		w_1002 , w_1003 , w_1004 , w_1005 , w_1006 , w_1007 , w_1008 , w_1009 , w_1010 , w_1011 , 
		w_1012 , w_1013 , w_1014 , w_1015 , w_1016 , w_1017 , w_1018 , w_1019 , w_1020 , w_1021 , 
		w_1022 , w_1023 , w_1024 , w_1025 , w_1026 , w_1027 , w_1028 , w_1029 , w_1030 , w_1031 , 
		w_1032 , w_1033 , w_1034 , w_1035 , w_1036 , w_1037 , w_1038 , w_1039 , w_1040 , w_1041 , 
		w_1042 , w_1043 , w_1044 , w_1045 , w_1046 , w_1047 , w_1048 , w_1049 , w_1050 , w_1051 , 
		w_1052 , w_1053 , w_1054 , w_1055 , w_1056 , w_1057 , w_1058 , w_1059 , w_1060 , w_1061 , 
		w_1062 , w_1063 , w_1064 , w_1065 , w_1066 , w_1067 , w_1068 , w_1069 , w_1070 , w_1071 , 
		w_1072 , w_1073 , w_1074 , w_1075 , w_1076 , w_1077 , w_1078 , w_1079 , w_1080 , w_1081 , 
		w_1082 , w_1083 , w_1084 , w_1085 , w_1086 , w_1087 , w_1088 , w_1089 , w_1090 , w_1091 , 
		w_1092 , w_1093 , w_1094 , w_1095 , w_1096 , w_1097 , w_1098 , w_1099 , w_1100 , w_1101 , 
		w_1102 , w_1103 , w_1104 , w_1105 , w_1106 , w_1107 , w_1108 , w_1109 , w_1110 , w_1111 , 
		w_1112 , w_1113 , w_1114 , w_1115 , w_1116 , w_1117 , w_1118 , w_1119 , w_1120 , w_1121 , 
		w_1122 , w_1123 , w_1124 , w_1125 , w_1126 , w_1127 , w_1128 , w_1129 , w_1130 , w_1131 , 
		w_1132 , w_1133 , w_1134 , w_1135 , w_1136 , w_1137 , w_1138 , w_1139 , w_1140 , w_1141 , 
		w_1142 , w_1143 , w_1144 , w_1145 , w_1146 , w_1147 , w_1148 , w_1149 , w_1150 , w_1151 , 
		w_1152 , w_1153 , w_1154 , w_1155 , w_1156 , w_1157 , w_1158 , w_1159 , w_1160 , w_1161 , 
		w_1162 , w_1163 , w_1164 , w_1165 , w_1166 , w_1167 , w_1168 , w_1169 , w_1170 , w_1171 , 
		w_1172 , w_1173 , w_1174 , w_1175 , w_1176 , w_1177 , w_1178 , w_1179 , w_1180 , w_1181 , 
		w_1182 , w_1183 , w_1184 , w_1185 , w_1186 , w_1187 , w_1188 , w_1189 , w_1190 , w_1191 , 
		w_1192 , w_1193 , w_1194 , w_1195 , w_1196 , w_1197 , w_1198 , w_1199 , w_1200 , w_1201 , 
		w_1202 , w_1203 , w_1204 , w_1205 , w_1206 , w_1207 , w_1208 , w_1209 , w_1210 , w_1211 , 
		w_1212 , w_1213 , w_1214 , w_1215 , w_1216 , w_1217 , w_1218 , w_1219 , w_1220 , w_1221 , 
		w_1222 , w_1223 , w_1224 , w_1225 , w_1226 , w_1227 , w_1228 , w_1229 , w_1230 , w_1231 , 
		w_1232 , w_1233 , w_1234 , w_1235 , w_1236 , w_1237 , w_1238 , w_1239 , w_1240 , w_1241 , 
		w_1242 , w_1243 , w_1244 , w_1245 , w_1246 , w_1247 , w_1248 , w_1249 , w_1250 , w_1251 , 
		w_1252 , w_1253 , w_1254 , w_1255 , w_1256 , w_1257 , w_1258 , w_1259 , w_1260 , w_1261 , 
		w_1262 , w_1263 , w_1264 , w_1265 , w_1266 , w_1267 , w_1268 , w_1269 , w_1270 , w_1271 , 
		w_1272 , w_1273 , w_1274 , w_1275 , w_1276 , w_1277 , w_1278 , w_1279 , w_1280 , w_1281 , 
		w_1282 , w_1283 , w_1284 , w_1285 , w_1286 , w_1287 , w_1288 , w_1289 , w_1290 , w_1291 , 
		w_1292 , w_1293 , w_1294 , w_1295 , w_1296 , w_1297 , w_1298 , w_1299 , w_1300 , w_1301 , 
		w_1302 , w_1303 , w_1304 , w_1305 , w_1306 , w_1307 , w_1308 , w_1309 , w_1310 , w_1311 , 
		w_1312 , w_1313 , w_1314 , w_1315 , w_1316 , w_1317 , w_1318 , w_1319 , w_1320 , w_1321 , 
		w_1322 , w_1323 , w_1324 , w_1325 , w_1326 , w_1327 , w_1328 , w_1329 , w_1330 , w_1331 , 
		w_1332 , w_1333 , w_1334 , w_1335 , w_1336 , w_1337 , w_1338 , w_1339 , w_1340 , w_1341 , 
		w_1342 , w_1343 , w_1344 , w_1345 , w_1346 , w_1347 , w_1348 , w_1349 , w_1350 , w_1351 , 
		w_1352 , w_1353 , w_1354 , w_1355 , w_1356 , w_1357 , w_1358 , w_1359 , w_1360 , w_1361 , 
		w_1362 , w_1363 , w_1364 , w_1365 , w_1366 , w_1367 , w_1368 , w_1369 , w_1370 , w_1371 , 
		w_1372 , w_1373 , w_1374 , w_1375 , w_1376 , w_1377 , w_1378 , w_1379 , w_1380 , w_1381 , 
		w_1382 , w_1383 , w_1384 , w_1385 , w_1386 , w_1387 , w_1388 , w_1389 , w_1390 , w_1391 , 
		w_1392 , w_1393 , w_1394 , w_1395 , w_1396 , w_1397 , w_1398 , w_1399 , w_1400 , w_1401 , 
		w_1402 , w_1403 , w_1404 , w_1405 , w_1406 , w_1407 , w_1408 , w_1409 , w_1410 , w_1411 , 
		w_1412 , w_1413 , w_1414 , w_1415 , w_1416 , w_1417 , w_1418 , w_1419 , w_1420 , w_1421 , 
		w_1422 , w_1423 , w_1424 , w_1425 , w_1426 , w_1427 , w_1428 , w_1429 , w_1430 , w_1431 , 
		w_1432 , w_1433 , w_1434 , w_1435 , w_1436 , w_1437 , w_1438 , w_1439 , w_1440 , w_1441 , 
		w_1442 , w_1443 , w_1444 , w_1445 , w_1446 , w_1447 , w_1448 , w_1449 , w_1450 , w_1451 , 
		w_1452 , w_1453 , w_1454 , w_1455 , w_1456 , w_1457 , w_1458 , w_1459 , w_1460 , w_1461 , 
		w_1462 , w_1463 , w_1464 , w_1465 , w_1466 , w_1467 , w_1468 , w_1469 , w_1470 , w_1471 , 
		w_1472 , w_1473 , w_1474 , w_1475 , w_1476 , w_1477 , w_1478 , w_1479 , w_1480 , w_1481 , 
		w_1482 , w_1483 , w_1484 , w_1485 , w_1486 , w_1487 , w_1488 , w_1489 , w_1490 , w_1491 , 
		w_1492 , w_1493 , w_1494 , w_1495 , w_1496 , w_1497 , w_1498 , w_1499 , w_1500 , w_1501 , 
		w_1502 , w_1503 , w_1504 , w_1505 , w_1506 , w_1507 , w_1508 , w_1509 , w_1510 , w_1511 , 
		w_1512 , w_1513 , w_1514 , w_1515 , w_1516 , w_1517 , w_1518 , w_1519 , w_1520 , w_1521 , 
		w_1522 , w_1523 , w_1524 , w_1525 , w_1526 , w_1527 , w_1528 , w_1529 , w_1530 , w_1531 , 
		w_1532 , w_1533 , w_1534 , w_1535 , w_1536 , w_1537 , w_1538 , w_1539 , w_1540 , w_1541 , 
		w_1542 , w_1543 , w_1544 , w_1545 , w_1546 , w_1547 , w_1548 , w_1549 , w_1550 , w_1551 , 
		w_1552 , w_1553 , w_1554 , w_1555 , w_1556 , w_1557 , w_1558 , w_1559 , w_1560 , w_1561 , 
		w_1562 , w_1563 , w_1564 , w_1565 , w_1566 , w_1567 , w_1568 , w_1569 , w_1570 , w_1571 , 
		w_1572 , w_1573 , w_1574 , w_1575 , w_1576 , w_1577 , w_1578 , w_1579 , w_1580 , w_1581 , 
		w_1582 , w_1583 , w_1584 , w_1585 , w_1586 , w_1587 , w_1588 , w_1589 , w_1590 , w_1591 , 
		w_1592 , w_1593 , w_1594 , w_1595 , w_1596 , w_1597 , w_1598 , w_1599 , w_1600 , w_1601 , 
		w_1602 , w_1603 , w_1604 , w_1605 , w_1606 , w_1607 , w_1608 , w_1609 , w_1610 , w_1611 , 
		w_1612 , w_1613 , w_1614 , w_1615 , w_1616 , w_1617 , w_1618 , w_1619 , w_1620 , w_1621 , 
		w_1622 , w_1623 , w_1624 , w_1625 , w_1626 , w_1627 , w_1628 , w_1629 , w_1630 , w_1631 , 
		w_1632 , w_1633 , w_1634 , w_1635 , w_1636 , w_1637 , w_1638 , w_1639 , w_1640 , w_1641 , 
		w_1642 , w_1643 , w_1644 , w_1645 , w_1646 , w_1647 , w_1648 , w_1649 , w_1650 , w_1651 , 
		w_1652 , w_1653 , w_1654 , w_1655 , w_1656 , w_1657 , w_1658 , w_1659 , w_1660 , w_1661 , 
		w_1662 , w_1663 , w_1664 , w_1665 , w_1666 , w_1667 , w_1668 , w_1669 , w_1670 , w_1671 , 
		w_1672 , w_1673 , w_1674 , w_1675 , w_1676 , w_1677 , w_1678 , w_1679 , w_1680 , w_1681 , 
		w_1682 , w_1683 , w_1684 , w_1685 , w_1686 , w_1687 , w_1688 , w_1689 , w_1690 , w_1691 , 
		w_1692 , w_1693 , w_1694 , w_1695 , w_1696 , w_1697 , w_1698 , w_1699 , w_1700 , w_1701 , 
		w_1702 , w_1703 , w_1704 , w_1705 , w_1706 , w_1707 , w_1708 , w_1709 , w_1710 , w_1711 , 
		w_1712 , w_1713 , w_1714 , w_1715 , w_1716 , w_1717 , w_1718 , w_1719 , w_1720 , w_1721 , 
		w_1722 , w_1723 , w_1724 , w_1725 , w_1726 , w_1727 , w_1728 , w_1729 , w_1730 , w_1731 , 
		w_1732 , w_1733 , w_1734 , w_1735 , w_1736 , w_1737 , w_1738 , w_1739 , w_1740 , w_1741 , 
		w_1742 , w_1743 , w_1744 , w_1745 , w_1746 , w_1747 , w_1748 , w_1749 , w_1750 , w_1751 , 
		w_1752 , w_1753 , w_1754 , w_1755 , w_1756 , w_1757 , w_1758 , w_1759 , w_1760 , w_1761 , 
		w_1762 , w_1763 , w_1764 , w_1765 , w_1766 , w_1767 , w_1768 , w_1769 , w_1770 , w_1771 , 
		w_1772 , w_1773 , w_1774 , w_1775 , w_1776 , w_1777 , w_1778 , w_1779 , w_1780 , w_1781 , 
		w_1782 , w_1783 , w_1784 , w_1785 , w_1786 , w_1787 , w_1788 , w_1789 , w_1790 , w_1791 , 
		w_1792 , w_1793 , w_1794 , w_1795 , w_1796 , w_1797 , w_1798 , w_1799 , w_1800 , w_1801 , 
		w_1802 , w_1803 , w_1804 , w_1805 , w_1806 , w_1807 , w_1808 , w_1809 , w_1810 , w_1811 , 
		w_1812 , w_1813 , w_1814 , w_1815 , w_1816 , w_1817 , w_1818 , w_1819 , w_1820 , w_1821 , 
		w_1822 , w_1823 , w_1824 , w_1825 , w_1826 , w_1827 , w_1828 , w_1829 , w_1830 , w_1831 , 
		w_1832 , w_1833 , w_1834 , w_1835 , w_1836 , w_1837 , w_1838 , w_1839 , w_1840 , w_1841 , 
		w_1842 , w_1843 , w_1844 , w_1845 , w_1846 , w_1847 , w_1848 , w_1849 , w_1850 , w_1851 , 
		w_1852 , w_1853 , w_1854 , w_1855 , w_1856 , w_1857 , w_1858 , w_1859 , w_1860 , w_1861 , 
		w_1862 , w_1863 , w_1864 , w_1865 , w_1866 , w_1867 , w_1868 , w_1869 , w_1870 , w_1871 , 
		w_1872 , w_1873 , w_1874 , w_1875 , w_1876 , w_1877 , w_1878 , w_1879 , w_1880 , w_1881 , 
		w_1882 , w_1883 , w_1884 , w_1885 , w_1886 , w_1887 , w_1888 , w_1889 , w_1890 , w_1891 , 
		w_1892 , w_1893 , w_1894 , w_1895 , w_1896 , w_1897 , w_1898 , w_1899 , w_1900 , w_1901 , 
		w_1902 , w_1903 , w_1904 , w_1905 , w_1906 , w_1907 , w_1908 , w_1909 , w_1910 , w_1911 , 
		w_1912 , w_1913 , w_1914 , w_1915 , w_1916 , w_1917 , w_1918 , w_1919 , w_1920 , w_1921 , 
		w_1922 , w_1923 , w_1924 , w_1925 , w_1926 , w_1927 , w_1928 , w_1929 , w_1930 , w_1931 , 
		w_1932 , w_1933 , w_1934 , w_1935 , w_1936 , w_1937 , w_1938 , w_1939 , w_1940 , w_1941 , 
		w_1942 , w_1943 , w_1944 , w_1945 , w_1946 , w_1947 , w_1948 , w_1949 , w_1950 , w_1951 , 
		w_1952 , w_1953 , w_1954 , w_1955 , w_1956 , w_1957 , w_1958 , w_1959 , w_1960 , w_1961 , 
		w_1962 , w_1963 , w_1964 , w_1965 , w_1966 , w_1967 , w_1968 , w_1969 , w_1970 , w_1971 , 
		w_1972 , w_1973 , w_1974 , w_1975 , w_1976 , w_1977 , w_1978 , w_1979 , w_1980 , w_1981 , 
		w_1982 , w_1983 , w_1984 , w_1985 , w_1986 , w_1987 , w_1988 , w_1989 , w_1990 , w_1991 , 
		w_1992 , w_1993 , w_1994 , w_1995 , w_1996 , w_1997 , w_1998 , w_1999 , w_2000 , w_2001 , 
		w_2002 , w_2003 , w_2004 , w_2005 , w_2006 , w_2007 , w_2008 , w_2009 , w_2010 , w_2011 , 
		w_2012 , w_2013 , w_2014 , w_2015 , w_2016 , w_2017 , w_2018 , w_2019 , w_2020 , w_2021 , 
		w_2022 , w_2023 , w_2024 , w_2025 , w_2026 , w_2027 , w_2028 , w_2029 , w_2030 , w_2031 , 
		w_2032 , w_2033 , w_2034 , w_2035 , w_2036 , w_2037 , w_2038 , w_2039 , w_2040 , w_2041 , 
		w_2042 , w_2043 , w_2044 , w_2045 , w_2046 , w_2047 , w_2048 , w_2049 , w_2050 , w_2051 , 
		w_2052 , w_2053 , w_2054 , w_2055 , w_2056 , w_2057 , w_2058 , w_2059 , w_2060 , w_2061 , 
		w_2062 , w_2063 , w_2064 , w_2065 , w_2066 , w_2067 , w_2068 , w_2069 , w_2070 , w_2071 , 
		w_2072 , w_2073 , w_2074 , w_2075 , w_2076 , w_2077 , w_2078 , w_2079 , w_2080 , w_2081 , 
		w_2082 , w_2083 , w_2084 , w_2085 , w_2086 , w_2087 , w_2088 , w_2089 , w_2090 , w_2091 , 
		w_2092 , w_2093 , w_2094 , w_2095 , w_2096 , w_2097 , w_2098 , w_2099 , w_2100 , w_2101 , 
		w_2102 , w_2103 , w_2104 , w_2105 , w_2106 , w_2107 , w_2108 , w_2109 , w_2110 , w_2111 , 
		w_2112 , w_2113 , w_2114 , w_2115 , w_2116 , w_2117 , w_2118 , w_2119 , w_2120 , w_2121 , 
		w_2122 , w_2123 , w_2124 , w_2125 , w_2126 , w_2127 , w_2128 , w_2129 , w_2130 , w_2131 , 
		w_2132 , w_2133 , w_2134 , w_2135 , w_2136 , w_2137 , w_2138 , w_2139 , w_2140 , w_2141 , 
		w_2142 , w_2143 , w_2144 , w_2145 , w_2146 , w_2147 , w_2148 , w_2149 , w_2150 , w_2151 , 
		w_2152 , w_2153 , w_2154 , w_2155 , w_2156 , w_2157 , w_2158 , w_2159 , w_2160 , w_2161 , 
		w_2162 , w_2163 , w_2164 , w_2165 , w_2166 , w_2167 , w_2168 , w_2169 , w_2170 , w_2171 , 
		w_2172 , w_2173 , w_2174 , w_2175 , w_2176 , w_2177 , w_2178 , w_2179 , w_2180 , w_2181 , 
		w_2182 , w_2183 , w_2184 , w_2185 , w_2186 , w_2187 , w_2188 , w_2189 , w_2190 , w_2191 , 
		w_2192 , w_2193 , w_2194 , w_2195 , w_2196 , w_2197 , w_2198 , w_2199 , w_2200 , w_2201 , 
		w_2202 , w_2203 , w_2204 , w_2205 , w_2206 , w_2207 , w_2208 , w_2209 , w_2210 , w_2211 , 
		w_2212 , w_2213 , w_2214 , w_2215 , w_2216 , w_2217 , w_2218 , w_2219 , w_2220 , w_2221 , 
		w_2222 , w_2223 , w_2224 , w_2225 , w_2226 , w_2227 , w_2228 , w_2229 , w_2230 , w_2231 , 
		w_2232 , w_2233 , w_2234 , w_2235 , w_2236 , w_2237 , w_2238 , w_2239 , w_2240 , w_2241 , 
		w_2242 , w_2243 , w_2244 , w_2245 , w_2246 , w_2247 , w_2248 , w_2249 , w_2250 , w_2251 , 
		w_2252 , w_2253 , w_2254 , w_2255 , w_2256 , w_2257 , w_2258 , w_2259 , w_2260 , w_2261 , 
		w_2262 , w_2263 , w_2264 , w_2265 , w_2266 , w_2267 , w_2268 , w_2269 , w_2270 , w_2271 , 
		w_2272 , w_2273 , w_2274 , w_2275 , w_2276 , w_2277 , w_2278 , w_2279 , w_2280 , w_2281 , 
		w_2282 , w_2283 , w_2284 , w_2285 , w_2286 , w_2287 , w_2288 , w_2289 , w_2290 , w_2291 , 
		w_2292 , w_2293 , w_2294 , w_2295 , w_2296 , w_2297 , w_2298 , w_2299 , w_2300 , w_2301 , 
		w_2302 , w_2303 , w_2304 , w_2305 , w_2306 , w_2307 , w_2308 , w_2309 , w_2310 , w_2311 , 
		w_2312 , w_2313 , w_2314 , w_2315 , w_2316 , w_2317 , w_2318 , w_2319 , w_2320 , w_2321 , 
		w_2322 , w_2323 , w_2324 , w_2325 , w_2326 , w_2327 , w_2328 , w_2329 , w_2330 , w_2331 , 
		w_2332 , w_2333 , w_2334 , w_2335 , w_2336 , w_2337 , w_2338 , w_2339 , w_2340 , w_2341 , 
		w_2342 , w_2343 , w_2344 , w_2345 , w_2346 , w_2347 , w_2348 , w_2349 , w_2350 , w_2351 , 
		w_2352 , w_2353 , w_2354 , w_2355 , w_2356 , w_2357 , w_2358 , w_2359 , w_2360 , w_2361 , 
		w_2362 , w_2363 , w_2364 , w_2365 , w_2366 , w_2367 , w_2368 , w_2369 , w_2370 , w_2371 , 
		w_2372 , w_2373 , w_2374 , w_2375 , w_2376 , w_2377 , w_2378 , w_2379 , w_2380 , w_2381 , 
		w_2382 , w_2383 , w_2384 , w_2385 , w_2386 , w_2387 , w_2388 , w_2389 , w_2390 , w_2391 , 
		w_2392 , w_2393 , w_2394 , w_2395 , w_2396 , w_2397 , w_2398 , w_2399 , w_2400 , w_2401 , 
		w_2402 , w_2403 , w_2404 , w_2405 , w_2406 , w_2407 , w_2408 , w_2409 , w_2410 , w_2411 , 
		w_2412 , w_2413 , w_2414 , w_2415 , w_2416 , w_2417 , w_2418 , w_2419 , w_2420 , w_2421 , 
		w_2422 , w_2423 , w_2424 , w_2425 , w_2426 , w_2427 , w_2428 , w_2429 , w_2430 , w_2431 , 
		w_2432 , w_2433 , w_2434 , w_2435 , w_2436 , w_2437 , w_2438 , w_2439 , w_2440 , w_2441 , 
		w_2442 , w_2443 , w_2444 , w_2445 , w_2446 , w_2447 , w_2448 , w_2449 , w_2450 , w_2451 , 
		w_2452 , w_2453 , w_2454 , w_2455 , w_2456 , w_2457 , w_2458 , w_2459 , w_2460 , w_2461 , 
		w_2462 , w_2463 , w_2464 , w_2465 , w_2466 , w_2467 , w_2468 , w_2469 , w_2470 , w_2471 , 
		w_2472 , w_2473 , w_2474 , w_2475 , w_2476 , w_2477 , w_2478 , w_2479 , w_2480 , w_2481 , 
		w_2482 , w_2483 , w_2484 , w_2485 , w_2486 , w_2487 , w_2488 , w_2489 , w_2490 , w_2491 , 
		w_2492 , w_2493 , w_2494 , w_2495 , w_2496 , w_2497 , w_2498 , w_2499 , w_2500 , w_2501 , 
		w_2502 , w_2503 , w_2504 , w_2505 , w_2506 , w_2507 , w_2508 , w_2509 , w_2510 , w_2511 , 
		w_2512 , w_2513 , w_2514 , w_2515 , w_2516 , w_2517 , w_2518 , w_2519 , w_2520 , w_2521 , 
		w_2522 , w_2523 , w_2524 , w_2525 , w_2526 , w_2527 , w_2528 , w_2529 , w_2530 , w_2531 , 
		w_2532 , w_2533 , w_2534 , w_2535 , w_2536 , w_2537 , w_2538 , w_2539 , w_2540 , w_2541 , 
		w_2542 , w_2543 , w_2544 , w_2545 , w_2546 , w_2547 , w_2548 , w_2549 , w_2550 , w_2551 , 
		w_2552 , w_2553 , w_2554 , w_2555 , w_2556 , w_2557 , w_2558 , w_2559 , w_2560 , w_2561 , 
		w_2562 , w_2563 , w_2564 , w_2565 , w_2566 , w_2567 , w_2568 , w_2569 , w_2570 , w_2571 , 
		w_2572 , w_2573 , w_2574 , w_2575 , w_2576 , w_2577 , w_2578 , w_2579 , w_2580 , w_2581 , 
		w_2582 , w_2583 , w_2584 , w_2585 , w_2586 , w_2587 , w_2588 , w_2589 , w_2590 , w_2591 , 
		w_2592 , w_2593 , w_2594 , w_2595 , w_2596 , w_2597 , w_2598 , w_2599 , w_2600 , w_2601 , 
		w_2602 , w_2603 , w_2604 , w_2605 , w_2606 , w_2607 , w_2608 , w_2609 , w_2610 , w_2611 , 
		w_2612 , w_2613 , w_2614 , w_2615 , w_2616 , w_2617 , w_2618 , w_2619 , w_2620 , w_2621 , 
		w_2622 , w_2623 , w_2624 , w_2625 , w_2626 , w_2627 , w_2628 , w_2629 , w_2630 , w_2631 , 
		w_2632 , w_2633 , w_2634 , w_2635 , w_2636 , w_2637 , w_2638 , w_2639 , w_2640 , w_2641 , 
		w_2642 , w_2643 , w_2644 , w_2645 , w_2646 , w_2647 , w_2648 , w_2649 , w_2650 , w_2651 , 
		w_2652 , w_2653 , w_2654 , w_2655 , w_2656 , w_2657 , w_2658 , w_2659 , w_2660 , w_2661 , 
		w_2662 , w_2663 , w_2664 , w_2665 , w_2666 , w_2667 , w_2668 , w_2669 , w_2670 , w_2671 , 
		w_2672 , w_2673 , w_2674 , w_2675 , w_2676 , w_2677 , w_2678 , w_2679 , w_2680 , w_2681 , 
		w_2682 , w_2683 , w_2684 , w_2685 , w_2686 , w_2687 , w_2688 , w_2689 , w_2690 , w_2691 , 
		w_2692 , w_2693 , w_2694 , w_2695 , w_2696 , w_2697 , w_2698 , w_2699 , w_2700 , w_2701 , 
		w_2702 , w_2703 , w_2704 , w_2705 , w_2706 , w_2707 , w_2708 , w_2709 , w_2710 , w_2711 , 
		w_2712 , w_2713 , w_2714 , w_2715 , w_2716 , w_2717 , w_2718 , w_2719 , w_2720 , w_2721 , 
		w_2722 , w_2723 , w_2724 , w_2725 , w_2726 , w_2727 , w_2728 , w_2729 , w_2730 , w_2731 , 
		w_2732 , w_2733 , w_2734 , w_2735 , w_2736 , w_2737 , w_2738 , w_2739 , w_2740 , w_2741 , 
		w_2742 , w_2743 , w_2744 , w_2745 , w_2746 , w_2747 , w_2748 , w_2749 , w_2750 , w_2751 , 
		w_2752 , w_2753 , w_2754 , w_2755 , w_2756 , w_2757 , w_2758 , w_2759 , w_2760 , w_2761 , 
		w_2762 , w_2763 , w_2764 , w_2765 , w_2766 , w_2767 , w_2768 , w_2769 , w_2770 , w_2771 , 
		w_2772 , w_2773 , w_2774 , w_2775 , w_2776 , w_2777 , w_2778 , w_2779 , w_2780 , w_2781 , 
		w_2782 , w_2783 , w_2784 , w_2785 , w_2786 , w_2787 , w_2788 , w_2789 , w_2790 , w_2791 , 
		w_2792 , w_2793 , w_2794 , w_2795 , w_2796 , w_2797 , w_2798 , w_2799 , w_2800 , w_2801 , 
		w_2802 , w_2803 , w_2804 , w_2805 , w_2806 , w_2807 , w_2808 , w_2809 , w_2810 , w_2811 , 
		w_2812 , w_2813 , w_2814 , w_2815 , w_2816 , w_2817 , w_2818 , w_2819 , w_2820 , w_2821 , 
		w_2822 , w_2823 , w_2824 , w_2825 , w_2826 , w_2827 , w_2828 , w_2829 , w_2830 , w_2831 , 
		w_2832 , w_2833 , w_2834 , w_2835 , w_2836 , w_2837 , w_2838 , w_2839 , w_2840 , w_2841 , 
		w_2842 , w_2843 , w_2844 , w_2845 , w_2846 , w_2847 , w_2848 , w_2849 , w_2850 , w_2851 , 
		w_2852 , w_2853 , w_2854 , w_2855 , w_2856 , w_2857 , w_2858 , w_2859 , w_2860 , w_2861 , 
		w_2862 , w_2863 , w_2864 , w_2865 , w_2866 , w_2867 , w_2868 , w_2869 , w_2870 , w_2871 , 
		w_2872 , w_2873 , w_2874 , w_2875 , w_2876 , w_2877 , w_2878 , w_2879 , w_2880 , w_2881 , 
		w_2882 , w_2883 , w_2884 , w_2885 , w_2886 , w_2887 , w_2888 , w_2889 , w_2890 , w_2891 , 
		w_2892 , w_2893 , w_2894 , w_2895 , w_2896 , w_2897 , w_2898 , w_2899 , w_2900 , w_2901 , 
		w_2902 , w_2903 , w_2904 , w_2905 , w_2906 , w_2907 , w_2908 , w_2909 , w_2910 , w_2911 , 
		w_2912 , w_2913 , w_2914 , w_2915 , w_2916 , w_2917 , w_2918 , w_2919 , w_2920 , w_2921 , 
		w_2922 , w_2923 , w_2924 , w_2925 , w_2926 , w_2927 , w_2928 , w_2929 , w_2930 , w_2931 , 
		w_2932 , w_2933 , w_2934 , w_2935 , w_2936 , w_2937 , w_2938 , w_2939 , w_2940 , w_2941 , 
		w_2942 , w_2943 , w_2944 , w_2945 , w_2946 , w_2947 , w_2948 , w_2949 , w_2950 , w_2951 , 
		w_2952 , w_2953 , w_2954 , w_2955 , w_2956 , w_2957 , w_2958 , w_2959 , w_2960 , w_2961 , 
		w_2962 , w_2963 , w_2964 , w_2965 , w_2966 , w_2967 , w_2968 , w_2969 , w_2970 , w_2971 , 
		w_2972 , w_2973 , w_2974 , w_2975 , w_2976 , w_2977 , w_2978 , w_2979 , w_2980 , w_2981 , 
		w_2982 , w_2983 , w_2984 , w_2985 , w_2986 , w_2987 , w_2988 , w_2989 , w_2990 , w_2991 , 
		w_2992 , w_2993 , w_2994 , w_2995 , w_2996 , w_2997 , w_2998 , w_2999 , w_3000 , w_3001 , 
		w_3002 , w_3003 , w_3004 , w_3005 , w_3006 , w_3007 , w_3008 , w_3009 , w_3010 , w_3011 , 
		w_3012 , w_3013 , w_3014 , w_3015 , w_3016 , w_3017 , w_3018 , w_3019 , w_3020 , w_3021 , 
		w_3022 , w_3023 , w_3024 , w_3025 , w_3026 , w_3027 , w_3028 , w_3029 , w_3030 , w_3031 , 
		w_3032 , w_3033 , w_3034 , w_3035 , w_3036 , w_3037 , w_3038 , w_3039 , w_3040 , w_3041 , 
		w_3042 , w_3043 , w_3044 , w_3045 , w_3046 , w_3047 , w_3048 , w_3049 , w_3050 , w_3051 , 
		w_3052 , w_3053 , w_3054 , w_3055 , w_3056 , w_3057 , w_3058 , w_3059 , w_3060 , w_3061 , 
		w_3062 , w_3063 , w_3064 , w_3065 , w_3066 , w_3067 , w_3068 , w_3069 , w_3070 , w_3071 , 
		w_3072 , w_3073 , w_3074 , w_3075 , w_3076 , w_3077 , w_3078 , w_3079 , w_3080 , w_3081 , 
		w_3082 , w_3083 , w_3084 , w_3085 , w_3086 , w_3087 , w_3088 , w_3089 , w_3090 , w_3091 , 
		w_3092 , w_3093 , w_3094 , w_3095 , w_3096 , w_3097 , w_3098 , w_3099 , w_3100 , w_3101 , 
		w_3102 , w_3103 , w_3104 , w_3105 , w_3106 , w_3107 , w_3108 , w_3109 , w_3110 , w_3111 , 
		w_3112 , w_3113 , w_3114 , w_3115 , w_3116 , w_3117 , w_3118 , w_3119 , w_3120 , w_3121 , 
		w_3122 , w_3123 , w_3124 , w_3125 , w_3126 , w_3127 , w_3128 , w_3129 , w_3130 , w_3131 , 
		w_3132 , w_3133 , w_3134 , w_3135 , w_3136 , w_3137 , w_3138 , w_3139 , w_3140 , w_3141 , 
		w_3142 , w_3143 , w_3144 , w_3145 , w_3146 , w_3147 , w_3148 , w_3149 , w_3150 , w_3151 , 
		w_3152 , w_3153 , w_3154 , w_3155 , w_3156 , w_3157 , w_3158 , w_3159 , w_3160 , w_3161 , 
		w_3162 , w_3163 , w_3164 , w_3165 , w_3166 , w_3167 , w_3168 , w_3169 , w_3170 , w_3171 , 
		w_3172 , w_3173 , w_3174 , w_3175 , w_3176 , w_3177 , w_3178 , w_3179 , w_3180 , w_3181 , 
		w_3182 , w_3183 , w_3184 , w_3185 , w_3186 , w_3187 , w_3188 , w_3189 , w_3190 , w_3191 , 
		w_3192 , w_3193 , w_3194 , w_3195 , w_3196 , w_3197 , w_3198 , w_3199 , w_3200 , w_3201 , 
		w_3202 , w_3203 , w_3204 , w_3205 , w_3206 , w_3207 , w_3208 , w_3209 , w_3210 , w_3211 , 
		w_3212 , w_3213 , w_3214 , w_3215 , w_3216 , w_3217 , w_3218 , w_3219 , w_3220 , w_3221 , 
		w_3222 , w_3223 , w_3224 , w_3225 , w_3226 , w_3227 , w_3228 , w_3229 , w_3230 , w_3231 , 
		w_3232 , w_3233 , w_3234 , w_3235 , w_3236 , w_3237 , w_3238 , w_3239 , w_3240 , w_3241 , 
		w_3242 , w_3243 , w_3244 , w_3245 , w_3246 , w_3247 , w_3248 , w_3249 , w_3250 , w_3251 , 
		w_3252 , w_3253 , w_3254 , w_3255 , w_3256 , w_3257 , w_3258 , w_3259 , w_3260 , w_3261 , 
		w_3262 , w_3263 , w_3264 , w_3265 , w_3266 , w_3267 , w_3268 , w_3269 , w_3270 , w_3271 , 
		w_3272 , w_3273 , w_3274 , w_3275 , w_3276 , w_3277 , w_3278 , w_3279 , w_3280 , w_3281 , 
		w_3282 , w_3283 , w_3284 , w_3285 , w_3286 , w_3287 , w_3288 , w_3289 , w_3290 , w_3291 , 
		w_3292 , w_3293 , w_3294 , w_3295 , w_3296 , w_3297 , w_3298 , w_3299 , w_3300 , w_3301 , 
		w_3302 , w_3303 , w_3304 , w_3305 , w_3306 , w_3307 , w_3308 , w_3309 , w_3310 , w_3311 , 
		w_3312 , w_3313 , w_3314 , w_3315 , w_3316 , w_3317 , w_3318 , w_3319 , w_3320 , w_3321 , 
		w_3322 , w_3323 , w_3324 , w_3325 , w_3326 , w_3327 , w_3328 , w_3329 , w_3330 , w_3331 , 
		w_3332 , w_3333 , w_3334 , w_3335 , w_3336 , w_3337 , w_3338 , w_3339 , w_3340 , w_3341 , 
		w_3342 , w_3343 , w_3344 , w_3345 , w_3346 , w_3347 , w_3348 , w_3349 , w_3350 , w_3351 , 
		w_3352 , w_3353 , w_3354 , w_3355 , w_3356 , w_3357 , w_3358 , w_3359 , w_3360 , w_3361 , 
		w_3362 , w_3363 , w_3364 , w_3365 , w_3366 , w_3367 , w_3368 , w_3369 , w_3370 , w_3371 , 
		w_3372 , w_3373 , w_3374 , w_3375 , w_3376 , w_3377 , w_3378 , w_3379 , w_3380 , w_3381 , 
		w_3382 , w_3383 , w_3384 , w_3385 , w_3386 , w_3387 , w_3388 , w_3389 , w_3390 , w_3391 , 
		w_3392 , w_3393 , w_3394 , w_3395 , w_3396 , w_3397 , w_3398 , w_3399 , w_3400 , w_3401 , 
		w_3402 , w_3403 , w_3404 , w_3405 , w_3406 , w_3407 , w_3408 , w_3409 , w_3410 , w_3411 , 
		w_3412 , w_3413 , w_3414 , w_3415 , w_3416 , w_3417 , w_3418 , w_3419 , w_3420 , w_3421 , 
		w_3422 , w_3423 , w_3424 , w_3425 , w_3426 , w_3427 , w_3428 , w_3429 , w_3430 , w_3431 , 
		w_3432 , w_3433 , w_3434 , w_3435 , w_3436 , w_3437 , w_3438 , w_3439 , w_3440 , w_3441 , 
		w_3442 , w_3443 , w_3444 , w_3445 , w_3446 , w_3447 , w_3448 , w_3449 , w_3450 , w_3451 , 
		w_3452 , w_3453 , w_3454 , w_3455 , w_3456 , w_3457 , w_3458 , w_3459 , w_3460 , w_3461 , 
		w_3462 , w_3463 , w_3464 , w_3465 , w_3466 , w_3467 , w_3468 , w_3469 , w_3470 , w_3471 , 
		w_3472 , w_3473 , w_3474 , w_3475 , w_3476 , w_3477 , w_3478 , w_3479 , w_3480 , w_3481 , 
		w_3482 , w_3483 , w_3484 , w_3485 , w_3486 , w_3487 , w_3488 , w_3489 , w_3490 , w_3491 , 
		w_3492 , w_3493 , w_3494 , w_3495 , w_3496 , w_3497 , w_3498 , w_3499 , w_3500 , w_3501 , 
		w_3502 , w_3503 , w_3504 , w_3505 , w_3506 , w_3507 , w_3508 , w_3509 , w_3510 , w_3511 , 
		w_3512 , w_3513 , w_3514 , w_3515 , w_3516 , w_3517 , w_3518 , w_3519 , w_3520 , w_3521 , 
		w_3522 , w_3523 , w_3524 , w_3525 , w_3526 , w_3527 , w_3528 , w_3529 , w_3530 , w_3531 , 
		w_3532 , w_3533 , w_3534 , w_3535 , w_3536 , w_3537 , w_3538 , w_3539 , w_3540 , w_3541 , 
		w_3542 , w_3543 , w_3544 , w_3545 , w_3546 , w_3547 , w_3548 , w_3549 , w_3550 , w_3551 , 
		w_3552 , w_3553 , w_3554 , w_3555 , w_3556 , w_3557 , w_3558 , w_3559 , w_3560 , w_3561 , 
		w_3562 , w_3563 , w_3564 , w_3565 , w_3566 , w_3567 , w_3568 , w_3569 , w_3570 , w_3571 , 
		w_3572 , w_3573 , w_3574 , w_3575 , w_3576 , w_3577 , w_3578 , w_3579 , w_3580 , w_3581 , 
		w_3582 , w_3583 , w_3584 , w_3585 , w_3586 , w_3587 , w_3588 , w_3589 , w_3590 , w_3591 , 
		w_3592 , w_3593 , w_3594 , w_3595 , w_3596 , w_3597 , w_3598 , w_3599 , w_3600 , w_3601 , 
		w_3602 , w_3603 , w_3604 , w_3605 , w_3606 , w_3607 , w_3608 , w_3609 , w_3610 , w_3611 , 
		w_3612 , w_3613 , w_3614 , w_3615 , w_3616 , w_3617 , w_3618 , w_3619 , w_3620 , w_3621 , 
		w_3622 , w_3623 , w_3624 , w_3625 , w_3626 , w_3627 , w_3628 , w_3629 , w_3630 , w_3631 , 
		w_3632 , w_3633 , w_3634 , w_3635 , w_3636 , w_3637 , w_3638 , w_3639 , w_3640 , w_3641 , 
		w_3642 , w_3643 , w_3644 , w_3645 , w_3646 , w_3647 , w_3648 , w_3649 , w_3650 , w_3651 , 
		w_3652 , w_3653 , w_3654 , w_3655 , w_3656 , w_3657 , w_3658 , w_3659 , w_3660 , w_3661 , 
		w_3662 , w_3663 , w_3664 , w_3665 , w_3666 , w_3667 , w_3668 , w_3669 , w_3670 , w_3671 , 
		w_3672 , w_3673 , w_3674 , w_3675 , w_3676 , w_3677 , w_3678 , w_3679 , w_3680 , w_3681 , 
		w_3682 , w_3683 , w_3684 , w_3685 , w_3686 , w_3687 , w_3688 , w_3689 , w_3690 , w_3691 , 
		w_3692 , w_3693 , w_3694 , w_3695 , w_3696 , w_3697 , w_3698 , w_3699 , w_3700 , w_3701 , 
		w_3702 , w_3703 , w_3704 , w_3705 , w_3706 , w_3707 , w_3708 , w_3709 , w_3710 , w_3711 , 
		w_3712 , w_3713 , w_3714 , w_3715 , w_3716 , w_3717 , w_3718 , w_3719 , w_3720 , w_3721 , 
		w_3722 , w_3723 , w_3724 , w_3725 , w_3726 , w_3727 , w_3728 , w_3729 , w_3730 , w_3731 , 
		w_3732 , w_3733 , w_3734 , w_3735 , w_3736 , w_3737 , w_3738 , w_3739 , w_3740 , w_3741 , 
		w_3742 , w_3743 , w_3744 , w_3745 , w_3746 , w_3747 , w_3748 , w_3749 , w_3750 , w_3751 , 
		w_3752 , w_3753 , w_3754 , w_3755 , w_3756 , w_3757 , w_3758 , w_3759 , w_3760 , w_3761 , 
		w_3762 , w_3763 , w_3764 , w_3765 , w_3766 , w_3767 , w_3768 , w_3769 , w_3770 , w_3771 , 
		w_3772 , w_3773 , w_3774 , w_3775 , w_3776 , w_3777 , w_3778 , w_3779 , w_3780 , w_3781 , 
		w_3782 , w_3783 , w_3784 , w_3785 , w_3786 , w_3787 , w_3788 , w_3789 , w_3790 , w_3791 , 
		w_3792 , w_3793 , w_3794 , w_3795 , w_3796 , w_3797 , w_3798 , w_3799 , w_3800 , w_3801 , 
		w_3802 , w_3803 , w_3804 , w_3805 , w_3806 , w_3807 , w_3808 , w_3809 , w_3810 , w_3811 , 
		w_3812 , w_3813 , w_3814 , w_3815 , w_3816 , w_3817 , w_3818 , w_3819 , w_3820 , w_3821 , 
		w_3822 , w_3823 , w_3824 , w_3825 , w_3826 , w_3827 , w_3828 , w_3829 , w_3830 , w_3831 , 
		w_3832 , w_3833 , w_3834 , w_3835 , w_3836 , w_3837 , w_3838 , w_3839 , w_3840 , w_3841 , 
		w_3842 , w_3843 , w_3844 , w_3845 , w_3846 , w_3847 , w_3848 , w_3849 , w_3850 , w_3851 , 
		w_3852 , w_3853 , w_3854 , w_3855 , w_3856 , w_3857 , w_3858 , w_3859 , w_3860 , w_3861 , 
		w_3862 , w_3863 , w_3864 , w_3865 , w_3866 , w_3867 , w_3868 , w_3869 , w_3870 , w_3871 , 
		w_3872 , w_3873 , w_3874 , w_3875 , w_3876 , w_3877 , w_3878 , w_3879 , w_3880 , w_3881 , 
		w_3882 , w_3883 , w_3884 , w_3885 , w_3886 , w_3887 , w_3888 , w_3889 , w_3890 , w_3891 , 
		w_3892 , w_3893 , w_3894 , w_3895 , w_3896 , w_3897 , w_3898 , w_3899 , w_3900 , w_3901 , 
		w_3902 , w_3903 , w_3904 , w_3905 , w_3906 , w_3907 , w_3908 , w_3909 , w_3910 , w_3911 , 
		w_3912 , w_3913 , w_3914 , w_3915 , w_3916 , w_3917 , w_3918 , w_3919 , w_3920 , w_3921 , 
		w_3922 , w_3923 , w_3924 , w_3925 , w_3926 , w_3927 , w_3928 , w_3929 , w_3930 , w_3931 , 
		w_3932 , w_3933 , w_3934 , w_3935 , w_3936 , w_3937 , w_3938 , w_3939 , w_3940 , w_3941 , 
		w_3942 , w_3943 , w_3944 , w_3945 , w_3946 , w_3947 , w_3948 , w_3949 , w_3950 , w_3951 , 
		w_3952 , w_3953 , w_3954 , w_3955 , w_3956 , w_3957 , w_3958 , w_3959 , w_3960 , w_3961 , 
		w_3962 , w_3963 , w_3964 , w_3965 , w_3966 , w_3967 , w_3968 , w_3969 , w_3970 , w_3971 , 
		w_3972 , w_3973 , w_3974 , w_3975 , w_3976 , w_3977 , w_3978 , w_3979 , w_3980 , w_3981 , 
		w_3982 , w_3983 , w_3984 , w_3985 , w_3986 , w_3987 , w_3988 , w_3989 , w_3990 , w_3991 , 
		w_3992 , w_3993 , w_3994 , w_3995 , w_3996 , w_3997 , w_3998 , w_3999 , w_4000 , w_4001 , 
		w_4002 , w_4003 , w_4004 , w_4005 , w_4006 , w_4007 , w_4008 , w_4009 , w_4010 , w_4011 , 
		w_4012 , w_4013 , w_4014 , w_4015 , w_4016 , w_4017 , w_4018 , w_4019 , w_4020 , w_4021 , 
		w_4022 , w_4023 , w_4024 , w_4025 , w_4026 , w_4027 , w_4028 , w_4029 , w_4030 , w_4031 , 
		w_4032 , w_4033 , w_4034 , w_4035 , w_4036 , w_4037 , w_4038 , w_4039 , w_4040 , w_4041 , 
		w_4042 , w_4043 , w_4044 , w_4045 , w_4046 , w_4047 , w_4048 , w_4049 , w_4050 , w_4051 , 
		w_4052 , w_4053 , w_4054 , w_4055 , w_4056 , w_4057 , w_4058 , w_4059 , w_4060 , w_4061 , 
		w_4062 , w_4063 , w_4064 , w_4065 , w_4066 , w_4067 , w_4068 , w_4069 , w_4070 , w_4071 , 
		w_4072 , w_4073 , w_4074 , w_4075 , w_4076 , w_4077 , w_4078 , w_4079 , w_4080 , w_4081 , 
		w_4082 , w_4083 , w_4084 , w_4085 , w_4086 , w_4087 , w_4088 , w_4089 , w_4090 , w_4091 , 
		w_4092 , w_4093 , w_4094 , w_4095 , w_4096 , w_4097 , w_4098 , w_4099 , w_4100 , w_4101 , 
		w_4102 , w_4103 , w_4104 , w_4105 , w_4106 , w_4107 , w_4108 , w_4109 , w_4110 , w_4111 , 
		w_4112 , w_4113 , w_4114 , w_4115 , w_4116 , w_4117 , w_4118 , w_4119 , w_4120 , w_4121 , 
		w_4122 , w_4123 , w_4124 , w_4125 , w_4126 , w_4127 , w_4128 , w_4129 , w_4130 , w_4131 , 
		w_4132 , w_4133 , w_4134 , w_4135 , w_4136 , w_4137 , w_4138 , w_4139 , w_4140 , w_4141 , 
		w_4142 , w_4143 , w_4144 , w_4145 , w_4146 , w_4147 , w_4148 , w_4149 , w_4150 , w_4151 , 
		w_4152 , w_4153 , w_4154 , w_4155 , w_4156 , w_4157 , w_4158 , w_4159 , w_4160 , w_4161 , 
		w_4162 , w_4163 , w_4164 , w_4165 , w_4166 , w_4167 , w_4168 , w_4169 , w_4170 , w_4171 , 
		w_4172 , w_4173 , w_4174 , w_4175 , w_4176 , w_4177 , w_4178 , w_4179 , w_4180 , w_4181 , 
		w_4182 , w_4183 , w_4184 , w_4185 , w_4186 , w_4187 , w_4188 , w_4189 , w_4190 , w_4191 , 
		w_4192 , w_4193 , w_4194 , w_4195 , w_4196 , w_4197 , w_4198 , w_4199 , w_4200 , w_4201 , 
		w_4202 , w_4203 , w_4204 , w_4205 , w_4206 , w_4207 , w_4208 , w_4209 , w_4210 , w_4211 , 
		w_4212 , w_4213 , w_4214 , w_4215 , w_4216 , w_4217 , w_4218 , w_4219 , w_4220 , w_4221 , 
		w_4222 , w_4223 , w_4224 , w_4225 , w_4226 , w_4227 , w_4228 , w_4229 , w_4230 , w_4231 , 
		w_4232 , w_4233 , w_4234 , w_4235 , w_4236 , w_4237 , w_4238 , w_4239 , w_4240 , w_4241 , 
		w_4242 , w_4243 , w_4244 , w_4245 , w_4246 , w_4247 , w_4248 , w_4249 , w_4250 , w_4251 , 
		w_4252 , w_4253 , w_4254 , w_4255 , w_4256 , w_4257 , w_4258 , w_4259 , w_4260 , w_4261 , 
		w_4262 , w_4263 , w_4264 , w_4265 , w_4266 , w_4267 , w_4268 , w_4269 , w_4270 , w_4271 , 
		w_4272 , w_4273 , w_4274 , w_4275 , w_4276 , w_4277 , w_4278 , w_4279 , w_4280 , w_4281 , 
		w_4282 , w_4283 , w_4284 , w_4285 , w_4286 , w_4287 , w_4288 , w_4289 , w_4290 , w_4291 , 
		w_4292 , w_4293 , w_4294 , w_4295 , w_4296 , w_4297 , w_4298 , w_4299 , w_4300 , w_4301 , 
		w_4302 , w_4303 , w_4304 , w_4305 , w_4306 , w_4307 , w_4308 , w_4309 , w_4310 , w_4311 , 
		w_4312 , w_4313 , w_4314 , w_4315 , w_4316 , w_4317 , w_4318 , w_4319 , w_4320 , w_4321 , 
		w_4322 , w_4323 , w_4324 , w_4325 , w_4326 , w_4327 , w_4328 , w_4329 , w_4330 , w_4331 , 
		w_4332 , w_4333 , w_4334 , w_4335 , w_4336 , w_4337 , w_4338 , w_4339 , w_4340 , w_4341 , 
		w_4342 , w_4343 , w_4344 , w_4345 , w_4346 , w_4347 , w_4348 , w_4349 , w_4350 , w_4351 , 
		w_4352 , w_4353 , w_4354 , w_4355 , w_4356 , w_4357 , w_4358 , w_4359 , w_4360 , w_4361 , 
		w_4362 , w_4363 , w_4364 , w_4365 , w_4366 , w_4367 , w_4368 , w_4369 , w_4370 , w_4371 , 
		w_4372 , w_4373 , w_4374 , w_4375 , w_4376 , w_4377 , w_4378 , w_4379 , w_4380 , w_4381 , 
		w_4382 , w_4383 , w_4384 , w_4385 , w_4386 , w_4387 , w_4388 , w_4389 , w_4390 , w_4391 , 
		w_4392 , w_4393 , w_4394 , w_4395 , w_4396 , w_4397 , w_4398 , w_4399 , w_4400 , w_4401 , 
		w_4402 , w_4403 , w_4404 , w_4405 , w_4406 , w_4407 , w_4408 , w_4409 , w_4410 , w_4411 , 
		w_4412 , w_4413 , w_4414 , w_4415 , w_4416 , w_4417 , w_4418 , w_4419 , w_4420 , w_4421 , 
		w_4422 , w_4423 , w_4424 , w_4425 , w_4426 , w_4427 , w_4428 , w_4429 , w_4430 , w_4431 , 
		w_4432 , w_4433 , w_4434 , w_4435 , w_4436 , w_4437 , w_4438 , w_4439 , w_4440 , w_4441 , 
		w_4442 , w_4443 , w_4444 , w_4445 , w_4446 , w_4447 , w_4448 , w_4449 , w_4450 , w_4451 , 
		w_4452 , w_4453 , w_4454 , w_4455 , w_4456 , w_4457 , w_4458 , w_4459 , w_4460 , w_4461 , 
		w_4462 , w_4463 , w_4464 , w_4465 , w_4466 , w_4467 , w_4468 , w_4469 , w_4470 , w_4471 , 
		w_4472 , w_4473 , w_4474 , w_4475 , w_4476 , w_4477 , w_4478 , w_4479 , w_4480 , w_4481 , 
		w_4482 , w_4483 , w_4484 , w_4485 , w_4486 , w_4487 , w_4488 , w_4489 , w_4490 , w_4491 , 
		w_4492 , w_4493 , w_4494 , w_4495 , w_4496 , w_4497 , w_4498 , w_4499 , w_4500 , w_4501 , 
		w_4502 , w_4503 , w_4504 , w_4505 , w_4506 , w_4507 , w_4508 , w_4509 , w_4510 , w_4511 , 
		w_4512 , w_4513 , w_4514 , w_4515 , w_4516 , w_4517 , w_4518 , w_4519 , w_4520 , w_4521 , 
		w_4522 , w_4523 , w_4524 , w_4525 , w_4526 , w_4527 , w_4528 , w_4529 , w_4530 , w_4531 , 
		w_4532 , w_4533 , w_4534 , w_4535 , w_4536 , w_4537 , w_4538 , w_4539 , w_4540 , w_4541 , 
		w_4542 , w_4543 , w_4544 , w_4545 , w_4546 , w_4547 , w_4548 , w_4549 , w_4550 , w_4551 , 
		w_4552 , w_4553 , w_4554 , w_4555 , w_4556 , w_4557 , w_4558 , w_4559 , w_4560 , w_4561 , 
		w_4562 , w_4563 , w_4564 , w_4565 , w_4566 , w_4567 , w_4568 , w_4569 , w_4570 , w_4571 , 
		w_4572 , w_4573 , w_4574 , w_4575 , w_4576 , w_4577 , w_4578 , w_4579 , w_4580 , w_4581 , 
		w_4582 , w_4583 , w_4584 , w_4585 , w_4586 , w_4587 , w_4588 , w_4589 , w_4590 , w_4591 , 
		w_4592 , w_4593 , w_4594 , w_4595 , w_4596 , w_4597 , w_4598 , w_4599 , w_4600 , w_4601 , 
		w_4602 , w_4603 , w_4604 , w_4605 , w_4606 , w_4607 , w_4608 , w_4609 , w_4610 , w_4611 , 
		w_4612 , w_4613 , w_4614 , w_4615 , w_4616 , w_4617 , w_4618 , w_4619 , w_4620 , w_4621 , 
		w_4622 , w_4623 , w_4624 , w_4625 , w_4626 , w_4627 , w_4628 , w_4629 , w_4630 , w_4631 , 
		w_4632 , w_4633 , w_4634 , w_4635 , w_4636 , w_4637 , w_4638 , w_4639 , w_4640 , w_4641 , 
		w_4642 , w_4643 , w_4644 , w_4645 , w_4646 , w_4647 , w_4648 , w_4649 , w_4650 , w_4651 , 
		w_4652 , w_4653 , w_4654 , w_4655 , w_4656 , w_4657 , w_4658 , w_4659 , w_4660 , w_4661 , 
		w_4662 , w_4663 , w_4664 , w_4665 , w_4666 , w_4667 , w_4668 , w_4669 , w_4670 , w_4671 , 
		w_4672 , w_4673 , w_4674 , w_4675 , w_4676 , w_4677 , w_4678 , w_4679 , w_4680 , w_4681 , 
		w_4682 , w_4683 , w_4684 , w_4685 , w_4686 , w_4687 , w_4688 , w_4689 , w_4690 , w_4691 , 
		w_4692 , w_4693 , w_4694 , w_4695 , w_4696 , w_4697 , w_4698 , w_4699 , w_4700 , w_4701 , 
		w_4702 , w_4703 , w_4704 , w_4705 , w_4706 , w_4707 , w_4708 , w_4709 , w_4710 , w_4711 , 
		w_4712 , w_4713 , w_4714 , w_4715 , w_4716 , w_4717 , w_4718 , w_4719 , w_4720 , w_4721 , 
		w_4722 , w_4723 , w_4724 , w_4725 , w_4726 , w_4727 , w_4728 , w_4729 , w_4730 , w_4731 , 
		w_4732 , w_4733 , w_4734 , w_4735 , w_4736 , w_4737 , w_4738 , w_4739 , w_4740 , w_4741 , 
		w_4742 , w_4743 , w_4744 , w_4745 , w_4746 , w_4747 , w_4748 , w_4749 , w_4750 , w_4751 , 
		w_4752 , w_4753 , w_4754 , w_4755 , w_4756 , w_4757 , w_4758 , w_4759 , w_4760 , w_4761 , 
		w_4762 , w_4763 , w_4764 , w_4765 , w_4766 , w_4767 , w_4768 , w_4769 , w_4770 , w_4771 , 
		w_4772 , w_4773 , w_4774 , w_4775 , w_4776 , w_4777 , w_4778 , w_4779 , w_4780 , w_4781 , 
		w_4782 , w_4783 , w_4784 , w_4785 , w_4786 , w_4787 , w_4788 , w_4789 , w_4790 , w_4791 , 
		w_4792 , w_4793 , w_4794 , w_4795 , w_4796 , w_4797 , w_4798 , w_4799 , w_4800 , w_4801 , 
		w_4802 , w_4803 , w_4804 , w_4805 , w_4806 , w_4807 , w_4808 , w_4809 , w_4810 , w_4811 , 
		w_4812 , w_4813 , w_4814 , w_4815 , w_4816 , w_4817 , w_4818 , w_4819 , w_4820 , w_4821 , 
		w_4822 , w_4823 , w_4824 , w_4825 , w_4826 , w_4827 , w_4828 , w_4829 , w_4830 , w_4831 , 
		w_4832 , w_4833 , w_4834 , w_4835 , w_4836 , w_4837 , w_4838 , w_4839 , w_4840 , w_4841 , 
		w_4842 , w_4843 , w_4844 , w_4845 , w_4846 , w_4847 , w_4848 , w_4849 , w_4850 , w_4851 , 
		w_4852 , w_4853 , w_4854 , w_4855 , w_4856 , w_4857 , w_4858 , w_4859 , w_4860 , w_4861 , 
		w_4862 , w_4863 , w_4864 , w_4865 , w_4866 , w_4867 , w_4868 , w_4869 , w_4870 , w_4871 , 
		w_4872 , w_4873 , w_4874 , w_4875 , w_4876 , w_4877 , w_4878 , w_4879 , w_4880 , w_4881 , 
		w_4882 , w_4883 , w_4884 , w_4885 , w_4886 , w_4887 , w_4888 , w_4889 , w_4890 , w_4891 , 
		w_4892 , w_4893 , w_4894 , w_4895 , w_4896 , w_4897 , w_4898 , w_4899 , w_4900 , w_4901 , 
		w_4902 , w_4903 , w_4904 , w_4905 , w_4906 , w_4907 , w_4908 , w_4909 , w_4910 , w_4911 , 
		w_4912 , w_4913 , w_4914 , w_4915 , w_4916 , w_4917 , w_4918 , w_4919 , w_4920 , w_4921 , 
		w_4922 , w_4923 , w_4924 , w_4925 , w_4926 , w_4927 , w_4928 , w_4929 , w_4930 , w_4931 , 
		w_4932 , w_4933 , w_4934 , w_4935 , w_4936 , w_4937 , w_4938 , w_4939 , w_4940 , w_4941 , 
		w_4942 , w_4943 , w_4944 , w_4945 , w_4946 , w_4947 , w_4948 , w_4949 , w_4950 , w_4951 , 
		w_4952 , w_4953 , w_4954 , w_4955 , w_4956 , w_4957 , w_4958 , w_4959 , w_4960 , w_4961 , 
		w_4962 , w_4963 , w_4964 , w_4965 , w_4966 , w_4967 , w_4968 , w_4969 , w_4970 , w_4971 , 
		w_4972 , w_4973 , w_4974 , w_4975 , w_4976 , w_4977 , w_4978 , w_4979 , w_4980 , w_4981 , 
		w_4982 , w_4983 , w_4984 , w_4985 , w_4986 , w_4987 , w_4988 , w_4989 , w_4990 , w_4991 , 
		w_4992 , w_4993 , w_4994 , w_4995 , w_4996 , w_4997 , w_4998 , w_4999 , w_5000 , w_5001 , 
		w_5002 , w_5003 , w_5004 , w_5005 , w_5006 , w_5007 , w_5008 , w_5009 , w_5010 , w_5011 , 
		w_5012 , w_5013 , w_5014 , w_5015 , w_5016 , w_5017 , w_5018 , w_5019 , w_5020 , w_5021 , 
		w_5022 , w_5023 , w_5024 , w_5025 , w_5026 , w_5027 , w_5028 , w_5029 , w_5030 , w_5031 , 
		w_5032 , w_5033 , w_5034 , w_5035 , w_5036 , w_5037 , w_5038 , w_5039 , w_5040 , w_5041 , 
		w_5042 , w_5043 , w_5044 , w_5045 , w_5046 , w_5047 , w_5048 , w_5049 , w_5050 , w_5051 , 
		w_5052 , w_5053 , w_5054 , w_5055 , w_5056 , w_5057 , w_5058 , w_5059 , w_5060 , w_5061 , 
		w_5062 , w_5063 , w_5064 , w_5065 , w_5066 , w_5067 , w_5068 , w_5069 , w_5070 , w_5071 , 
		w_5072 , w_5073 , w_5074 , w_5075 , w_5076 , w_5077 , w_5078 , w_5079 , w_5080 , w_5081 , 
		w_5082 , w_5083 , w_5084 , w_5085 , w_5086 , w_5087 , w_5088 , w_5089 , w_5090 , w_5091 , 
		w_5092 , w_5093 , w_5094 , w_5095 , w_5096 , w_5097 , w_5098 , w_5099 , w_5100 , w_5101 , 
		w_5102 , w_5103 , w_5104 , w_5105 , w_5106 , w_5107 , w_5108 , w_5109 , w_5110 , w_5111 , 
		w_5112 , w_5113 , w_5114 , w_5115 , w_5116 , w_5117 , w_5118 , w_5119 , w_5120 , w_5121 , 
		w_5122 , w_5123 , w_5124 , w_5125 , w_5126 , w_5127 , w_5128 , w_5129 , w_5130 , w_5131 , 
		w_5132 , w_5133 , w_5134 , w_5135 , w_5136 , w_5137 , w_5138 , w_5139 , w_5140 , w_5141 , 
		w_5142 , w_5143 , w_5144 , w_5145 , w_5146 , w_5147 , w_5148 , w_5149 , w_5150 , w_5151 , 
		w_5152 , w_5153 , w_5154 , w_5155 , w_5156 , w_5157 , w_5158 , w_5159 , w_5160 , w_5161 , 
		w_5162 , w_5163 , w_5164 , w_5165 , w_5166 , w_5167 , w_5168 , w_5169 , w_5170 , w_5171 , 
		w_5172 , w_5173 , w_5174 , w_5175 , w_5176 , w_5177 , w_5178 , w_5179 , w_5180 , w_5181 , 
		w_5182 , w_5183 , w_5184 , w_5185 , w_5186 , w_5187 , w_5188 , w_5189 , w_5190 , w_5191 , 
		w_5192 , w_5193 , w_5194 , w_5195 , w_5196 , w_5197 , w_5198 , w_5199 , w_5200 , w_5201 , 
		w_5202 , w_5203 , w_5204 , w_5205 , w_5206 , w_5207 , w_5208 , w_5209 , w_5210 , w_5211 , 
		w_5212 , w_5213 , w_5214 , w_5215 , w_5216 , w_5217 , w_5218 , w_5219 , w_5220 , w_5221 , 
		w_5222 , w_5223 , w_5224 , w_5225 , w_5226 , w_5227 , w_5228 , w_5229 , w_5230 , w_5231 , 
		w_5232 , w_5233 , w_5234 , w_5235 , w_5236 , w_5237 , w_5238 , w_5239 , w_5240 , w_5241 , 
		w_5242 , w_5243 , w_5244 , w_5245 , w_5246 , w_5247 , w_5248 , w_5249 , w_5250 , w_5251 , 
		w_5252 , w_5253 , w_5254 , w_5255 , w_5256 , w_5257 , w_5258 , w_5259 , w_5260 , w_5261 , 
		w_5262 , w_5263 , w_5264 , w_5265 , w_5266 , w_5267 , w_5268 , w_5269 , w_5270 , w_5271 , 
		w_5272 , w_5273 , w_5274 , w_5275 , w_5276 , w_5277 , w_5278 , w_5279 , w_5280 , w_5281 , 
		w_5282 , w_5283 , w_5284 , w_5285 , w_5286 , w_5287 , w_5288 , w_5289 , w_5290 , w_5291 , 
		w_5292 , w_5293 , w_5294 , w_5295 , w_5296 , w_5297 , w_5298 , w_5299 , w_5300 , w_5301 , 
		w_5302 , w_5303 , w_5304 , w_5305 , w_5306 , w_5307 , w_5308 , w_5309 , w_5310 , w_5311 , 
		w_5312 , w_5313 , w_5314 , w_5315 , w_5316 , w_5317 , w_5318 , w_5319 , w_5320 , w_5321 , 
		w_5322 , w_5323 , w_5324 , w_5325 , w_5326 , w_5327 , w_5328 , w_5329 , w_5330 , w_5331 , 
		w_5332 , w_5333 , w_5334 , w_5335 , w_5336 , w_5337 , w_5338 , w_5339 , w_5340 , w_5341 , 
		w_5342 , w_5343 , w_5344 , w_5345 , w_5346 , w_5347 , w_5348 , w_5349 , w_5350 , w_5351 , 
		w_5352 , w_5353 , w_5354 , w_5355 , w_5356 , w_5357 , w_5358 , w_5359 , w_5360 , w_5361 , 
		w_5362 , w_5363 , w_5364 , w_5365 , w_5366 , w_5367 , w_5368 , w_5369 , w_5370 , w_5371 , 
		w_5372 , w_5373 , w_5374 , w_5375 , w_5376 , w_5377 , w_5378 , w_5379 , w_5380 , w_5381 , 
		w_5382 , w_5383 , w_5384 , w_5385 , w_5386 , w_5387 , w_5388 , w_5389 , w_5390 , w_5391 , 
		w_5392 , w_5393 , w_5394 , w_5395 , w_5396 , w_5397 , w_5398 , w_5399 , w_5400 , w_5401 , 
		w_5402 , w_5403 , w_5404 , w_5405 , w_5406 , w_5407 , w_5408 , w_5409 , w_5410 , w_5411 , 
		w_5412 , w_5413 , w_5414 , w_5415 , w_5416 , w_5417 , w_5418 , w_5419 , w_5420 , w_5421 , 
		w_5422 , w_5423 , w_5424 , w_5425 , w_5426 , w_5427 , w_5428 , w_5429 , w_5430 , w_5431 , 
		w_5432 , w_5433 , w_5434 , w_5435 , w_5436 , w_5437 , w_5438 , w_5439 , w_5440 , w_5441 , 
		w_5442 , w_5443 , w_5444 , w_5445 , w_5446 , w_5447 , w_5448 , w_5449 , w_5450 , w_5451 , 
		w_5452 , w_5453 , w_5454 , w_5455 , w_5456 , w_5457 , w_5458 , w_5459 , w_5460 , w_5461 , 
		w_5462 , w_5463 , w_5464 , w_5465 , w_5466 , w_5467 , w_5468 , w_5469 , w_5470 , w_5471 , 
		w_5472 , w_5473 , w_5474 , w_5475 , w_5476 , w_5477 , w_5478 , w_5479 , w_5480 , w_5481 , 
		w_5482 , w_5483 , w_5484 , w_5485 , w_5486 , w_5487 , w_5488 , w_5489 , w_5490 , w_5491 , 
		w_5492 , w_5493 , w_5494 , w_5495 , w_5496 , w_5497 , w_5498 , w_5499 , w_5500 , w_5501 , 
		w_5502 , w_5503 , w_5504 , w_5505 , w_5506 , w_5507 , w_5508 , w_5509 , w_5510 , w_5511 , 
		w_5512 , w_5513 , w_5514 , w_5515 , w_5516 , w_5517 , w_5518 , w_5519 , w_5520 , w_5521 , 
		w_5522 , w_5523 , w_5524 , w_5525 , w_5526 , w_5527 , w_5528 , w_5529 , w_5530 , w_5531 , 
		w_5532 , w_5533 , w_5534 , w_5535 , w_5536 , w_5537 , w_5538 , w_5539 , w_5540 , w_5541 , 
		w_5542 , w_5543 , w_5544 , w_5545 , w_5546 , w_5547 , w_5548 , w_5549 , w_5550 , w_5551 , 
		w_5552 , w_5553 , w_5554 , w_5555 , w_5556 , w_5557 , w_5558 , w_5559 , w_5560 , w_5561 , 
		w_5562 , w_5563 , w_5564 , w_5565 , w_5566 , w_5567 , w_5568 , w_5569 , w_5570 , w_5571 , 
		w_5572 , w_5573 , w_5574 , w_5575 , w_5576 , w_5577 , w_5578 , w_5579 , w_5580 , w_5581 , 
		w_5582 , w_5583 , w_5584 , w_5585 , w_5586 , w_5587 , w_5588 , w_5589 , w_5590 , w_5591 , 
		w_5592 , w_5593 , w_5594 , w_5595 , w_5596 , w_5597 , w_5598 , w_5599 , w_5600 , w_5601 , 
		w_5602 , w_5603 , w_5604 , w_5605 , w_5606 , w_5607 , w_5608 , w_5609 , w_5610 , w_5611 , 
		w_5612 , w_5613 , w_5614 , w_5615 , w_5616 , w_5617 , w_5618 , w_5619 , w_5620 , w_5621 , 
		w_5622 , w_5623 , w_5624 , w_5625 , w_5626 , w_5627 , w_5628 , w_5629 , w_5630 , w_5631 , 
		w_5632 , w_5633 , w_5634 , w_5635 , w_5636 , w_5637 , w_5638 , w_5639 , w_5640 , w_5641 , 
		w_5642 , w_5643 , w_5644 , w_5645 , w_5646 , w_5647 , w_5648 , w_5649 , w_5650 , w_5651 , 
		w_5652 , w_5653 , w_5654 , w_5655 , w_5656 , w_5657 , w_5658 , w_5659 , w_5660 , w_5661 , 
		w_5662 , w_5663 , w_5664 , w_5665 , w_5666 , w_5667 , w_5668 , w_5669 , w_5670 , w_5671 , 
		w_5672 , w_5673 , w_5674 , w_5675 , w_5676 , w_5677 , w_5678 , w_5679 , w_5680 , w_5681 , 
		w_5682 , w_5683 , w_5684 , w_5685 , w_5686 , w_5687 , w_5688 , w_5689 , w_5690 , w_5691 , 
		w_5692 , w_5693 , w_5694 , w_5695 , w_5696 , w_5697 , w_5698 , w_5699 , w_5700 , w_5701 , 
		w_5702 , w_5703 , w_5704 , w_5705 , w_5706 , w_5707 , w_5708 , w_5709 , w_5710 , w_5711 , 
		w_5712 , w_5713 , w_5714 , w_5715 , w_5716 , w_5717 , w_5718 , w_5719 , w_5720 , w_5721 , 
		w_5722 , w_5723 , w_5724 , w_5725 , w_5726 , w_5727 , w_5728 , w_5729 , w_5730 , w_5731 , 
		w_5732 , w_5733 , w_5734 , w_5735 , w_5736 , w_5737 , w_5738 , w_5739 , w_5740 , w_5741 , 
		w_5742 , w_5743 , w_5744 , w_5745 , w_5746 , w_5747 , w_5748 , w_5749 , w_5750 , w_5751 , 
		w_5752 , w_5753 , w_5754 , w_5755 , w_5756 , w_5757 , w_5758 , w_5759 , w_5760 , w_5761 , 
		w_5762 , w_5763 , w_5764 , w_5765 , w_5766 , w_5767 , w_5768 , w_5769 , w_5770 , w_5771 , 
		w_5772 , w_5773 , w_5774 , w_5775 , w_5776 , w_5777 , w_5778 , w_5779 , w_5780 , w_5781 , 
		w_5782 , w_5783 , w_5784 , w_5785 , w_5786 , w_5787 , w_5788 , w_5789 , w_5790 , w_5791 , 
		w_5792 , w_5793 , w_5794 , w_5795 , w_5796 , w_5797 , w_5798 , w_5799 , w_5800 , w_5801 , 
		w_5802 , w_5803 , w_5804 , w_5805 , w_5806 , w_5807 , w_5808 , w_5809 , w_5810 , w_5811 , 
		w_5812 , w_5813 , w_5814 , w_5815 , w_5816 , w_5817 , w_5818 , w_5819 , w_5820 , w_5821 , 
		w_5822 , w_5823 , w_5824 , w_5825 , w_5826 , w_5827 , w_5828 , w_5829 , w_5830 , w_5831 , 
		w_5832 , w_5833 , w_5834 , w_5835 , w_5836 , w_5837 , w_5838 , w_5839 , w_5840 , w_5841 , 
		w_5842 , w_5843 , w_5844 , w_5845 , w_5846 , w_5847 , w_5848 , w_5849 , w_5850 , w_5851 , 
		w_5852 , w_5853 , w_5854 , w_5855 , w_5856 , w_5857 , w_5858 , w_5859 , w_5860 , w_5861 , 
		w_5862 , w_5863 , w_5864 , w_5865 , w_5866 , w_5867 , w_5868 , w_5869 , w_5870 , w_5871 , 
		w_5872 , w_5873 , w_5874 , w_5875 , w_5876 , w_5877 , w_5878 , w_5879 , w_5880 , w_5881 , 
		w_5882 , w_5883 , w_5884 , w_5885 , w_5886 , w_5887 , w_5888 , w_5889 , w_5890 , w_5891 , 
		w_5892 , w_5893 , w_5894 , w_5895 , w_5896 , w_5897 , w_5898 , w_5899 , w_5900 , w_5901 , 
		w_5902 , w_5903 , w_5904 , w_5905 , w_5906 , w_5907 , w_5908 , w_5909 , w_5910 , w_5911 , 
		w_5912 , w_5913 , w_5914 , w_5915 , w_5916 , w_5917 , w_5918 , w_5919 , w_5920 , w_5921 , 
		w_5922 , w_5923 , w_5924 , w_5925 , w_5926 , w_5927 , w_5928 , w_5929 , w_5930 , w_5931 , 
		w_5932 , w_5933 , w_5934 , w_5935 , w_5936 , w_5937 , w_5938 , w_5939 , w_5940 , w_5941 , 
		w_5942 , w_5943 , w_5944 , w_5945 , w_5946 , w_5947 , w_5948 , w_5949 , w_5950 , w_5951 , 
		w_5952 , w_5953 , w_5954 , w_5955 , w_5956 , w_5957 , w_5958 , w_5959 , w_5960 , w_5961 , 
		w_5962 , w_5963 , w_5964 , w_5965 , w_5966 , w_5967 , w_5968 , w_5969 , w_5970 , w_5971 , 
		w_5972 , w_5973 , w_5974 , w_5975 , w_5976 , w_5977 , w_5978 , w_5979 , w_5980 , w_5981 , 
		w_5982 , w_5983 , w_5984 , w_5985 , w_5986 , w_5987 , w_5988 , w_5989 , w_5990 , w_5991 , 
		w_5992 , w_5993 , w_5994 , w_5995 , w_5996 , w_5997 , w_5998 , w_5999 , w_6000 , w_6001 , 
		w_6002 , w_6003 , w_6004 , w_6005 , w_6006 , w_6007 , w_6008 , w_6009 , w_6010 , w_6011 , 
		w_6012 , w_6013 , w_6014 , w_6015 , w_6016 , w_6017 , w_6018 , w_6019 , w_6020 , w_6021 , 
		w_6022 , w_6023 , w_6024 , w_6025 , w_6026 , w_6027 , w_6028 , w_6029 , w_6030 , w_6031 , 
		w_6032 , w_6033 , w_6034 , w_6035 , w_6036 , w_6037 , w_6038 , w_6039 , w_6040 , w_6041 , 
		w_6042 , w_6043 , w_6044 , w_6045 , w_6046 , w_6047 , w_6048 , w_6049 , w_6050 , w_6051 , 
		w_6052 , w_6053 , w_6054 , w_6055 , w_6056 , w_6057 , w_6058 , w_6059 , w_6060 , w_6061 , 
		w_6062 , w_6063 , w_6064 , w_6065 , w_6066 , w_6067 , w_6068 , w_6069 , w_6070 , w_6071 , 
		w_6072 , w_6073 , w_6074 , w_6075 , w_6076 , w_6077 , w_6078 , w_6079 , w_6080 , w_6081 , 
		w_6082 , w_6083 , w_6084 , w_6085 , w_6086 , w_6087 , w_6088 , w_6089 , w_6090 , w_6091 , 
		w_6092 , w_6093 , w_6094 , w_6095 , w_6096 , w_6097 , w_6098 , w_6099 , w_6100 , w_6101 , 
		w_6102 , w_6103 , w_6104 , w_6105 , w_6106 , w_6107 , w_6108 , w_6109 , w_6110 , w_6111 , 
		w_6112 , w_6113 , w_6114 , w_6115 , w_6116 , w_6117 , w_6118 , w_6119 , w_6120 , w_6121 , 
		w_6122 , w_6123 , w_6124 , w_6125 , w_6126 , w_6127 , w_6128 , w_6129 , w_6130 , w_6131 , 
		w_6132 , w_6133 , w_6134 , w_6135 , w_6136 , w_6137 , w_6138 , w_6139 , w_6140 , w_6141 , 
		w_6142 , w_6143 , w_6144 , w_6145 , w_6146 , w_6147 , w_6148 , w_6149 , w_6150 , w_6151 , 
		w_6152 , w_6153 , w_6154 , w_6155 , w_6156 , w_6157 , w_6158 , w_6159 , w_6160 , w_6161 , 
		w_6162 , w_6163 , w_6164 , w_6165 , w_6166 , w_6167 , w_6168 , w_6169 , w_6170 , w_6171 , 
		w_6172 , w_6173 , w_6174 , w_6175 , w_6176 , w_6177 , w_6178 , w_6179 , w_6180 , w_6181 , 
		w_6182 , w_6183 , w_6184 , w_6185 , w_6186 , w_6187 , w_6188 , w_6189 , w_6190 , w_6191 , 
		w_6192 , w_6193 , w_6194 , w_6195 , w_6196 , w_6197 , w_6198 , w_6199 , w_6200 , w_6201 , 
		w_6202 , w_6203 , w_6204 , w_6205 , w_6206 , w_6207 , w_6208 , w_6209 , w_6210 , w_6211 , 
		w_6212 , w_6213 , w_6214 , w_6215 , w_6216 , w_6217 , w_6218 , w_6219 , w_6220 , w_6221 , 
		w_6222 , w_6223 , w_6224 , w_6225 , w_6226 , w_6227 , w_6228 , w_6229 , w_6230 , w_6231 , 
		w_6232 , w_6233 , w_6234 , w_6235 , w_6236 , w_6237 , w_6238 , w_6239 , w_6240 , w_6241 , 
		w_6242 , w_6243 , w_6244 , w_6245 , w_6246 , w_6247 , w_6248 , w_6249 , w_6250 , w_6251 , 
		w_6252 , w_6253 , w_6254 , w_6255 , w_6256 , w_6257 , w_6258 , w_6259 , w_6260 , w_6261 , 
		w_6262 , w_6263 , w_6264 , w_6265 , w_6266 , w_6267 , w_6268 , w_6269 , w_6270 , w_6271 , 
		w_6272 , w_6273 , w_6274 , w_6275 , w_6276 , w_6277 , w_6278 , w_6279 , w_6280 , w_6281 , 
		w_6282 , w_6283 , w_6284 , w_6285 , w_6286 , w_6287 , w_6288 , w_6289 , w_6290 , w_6291 , 
		w_6292 , w_6293 , w_6294 , w_6295 , w_6296 , w_6297 , w_6298 , w_6299 , w_6300 , w_6301 , 
		w_6302 , w_6303 , w_6304 , w_6305 , w_6306 , w_6307 , w_6308 , w_6309 , w_6310 , w_6311 , 
		w_6312 , w_6313 , w_6314 , w_6315 , w_6316 , w_6317 , w_6318 , w_6319 , w_6320 , w_6321 , 
		w_6322 , w_6323 , w_6324 , w_6325 , w_6326 , w_6327 , w_6328 , w_6329 , w_6330 , w_6331 , 
		w_6332 , w_6333 , w_6334 , w_6335 , w_6336 , w_6337 , w_6338 , w_6339 , w_6340 , w_6341 , 
		w_6342 , w_6343 , w_6344 , w_6345 , w_6346 , w_6347 , w_6348 , w_6349 , w_6350 , w_6351 , 
		w_6352 , w_6353 , w_6354 , w_6355 , w_6356 , w_6357 , w_6358 , w_6359 , w_6360 , w_6361 , 
		w_6362 , w_6363 , w_6364 , w_6365 , w_6366 , w_6367 , w_6368 , w_6369 , w_6370 , w_6371 , 
		w_6372 , w_6373 , w_6374 , w_6375 , w_6376 , w_6377 , w_6378 , w_6379 , w_6380 , w_6381 , 
		w_6382 , w_6383 , w_6384 , w_6385 , w_6386 , w_6387 , w_6388 , w_6389 , w_6390 , w_6391 , 
		w_6392 , w_6393 , w_6394 , w_6395 , w_6396 , w_6397 , w_6398 , w_6399 , w_6400 , w_6401 , 
		w_6402 , w_6403 , w_6404 , w_6405 , w_6406 , w_6407 , w_6408 , w_6409 , w_6410 , w_6411 , 
		w_6412 , w_6413 , w_6414 , w_6415 , w_6416 , w_6417 , w_6418 , w_6419 , w_6420 , w_6421 , 
		w_6422 , w_6423 , w_6424 , w_6425 , w_6426 , w_6427 , w_6428 , w_6429 , w_6430 , w_6431 , 
		w_6432 , w_6433 , w_6434 , w_6435 , w_6436 , w_6437 , w_6438 , w_6439 , w_6440 , w_6441 , 
		w_6442 , w_6443 , w_6444 , w_6445 , w_6446 , w_6447 , w_6448 , w_6449 , w_6450 , w_6451 , 
		w_6452 , w_6453 , w_6454 , w_6455 , w_6456 , w_6457 , w_6458 , w_6459 , w_6460 , w_6461 , 
		w_6462 , w_6463 , w_6464 , w_6465 , w_6466 , w_6467 , w_6468 , w_6469 , w_6470 , w_6471 , 
		w_6472 , w_6473 , w_6474 , w_6475 , w_6476 , w_6477 , w_6478 , w_6479 , w_6480 , w_6481 , 
		w_6482 , w_6483 , w_6484 , w_6485 , w_6486 , w_6487 , w_6488 , w_6489 , w_6490 , w_6491 , 
		w_6492 , w_6493 , w_6494 , w_6495 , w_6496 , w_6497 , w_6498 , w_6499 , w_6500 , w_6501 , 
		w_6502 , w_6503 , w_6504 , w_6505 , w_6506 , w_6507 , w_6508 , w_6509 , w_6510 , w_6511 , 
		w_6512 , w_6513 , w_6514 , w_6515 , w_6516 , w_6517 , w_6518 , w_6519 , w_6520 , w_6521 , 
		w_6522 , w_6523 , w_6524 , w_6525 , w_6526 , w_6527 , w_6528 , w_6529 , w_6530 , w_6531 , 
		w_6532 , w_6533 , w_6534 , w_6535 , w_6536 , w_6537 , w_6538 , w_6539 , w_6540 , w_6541 , 
		w_6542 , w_6543 , w_6544 , w_6545 , w_6546 , w_6547 , w_6548 , w_6549 , w_6550 , w_6551 , 
		w_6552 , w_6553 , w_6554 , w_6555 , w_6556 , w_6557 , w_6558 , w_6559 , w_6560 , w_6561 , 
		w_6562 , w_6563 , w_6564 , w_6565 , w_6566 , w_6567 , w_6568 , w_6569 , w_6570 , w_6571 , 
		w_6572 , w_6573 , w_6574 , w_6575 , w_6576 , w_6577 , w_6578 , w_6579 , w_6580 , w_6581 , 
		w_6582 , w_6583 , w_6584 , w_6585 , w_6586 , w_6587 , w_6588 , w_6589 , w_6590 , w_6591 , 
		w_6592 , w_6593 , w_6594 , w_6595 , w_6596 , w_6597 , w_6598 , w_6599 , w_6600 , w_6601 , 
		w_6602 , w_6603 , w_6604 , w_6605 , w_6606 , w_6607 , w_6608 , w_6609 , w_6610 , w_6611 , 
		w_6612 , w_6613 , w_6614 , w_6615 , w_6616 , w_6617 , w_6618 , w_6619 , w_6620 , w_6621 , 
		w_6622 , w_6623 , w_6624 , w_6625 , w_6626 , w_6627 , w_6628 , w_6629 , w_6630 , w_6631 , 
		w_6632 , w_6633 , w_6634 , w_6635 , w_6636 , w_6637 , w_6638 , w_6639 , w_6640 , w_6641 , 
		w_6642 , w_6643 , w_6644 , w_6645 , w_6646 , w_6647 , w_6648 , w_6649 , w_6650 , w_6651 , 
		w_6652 , w_6653 , w_6654 , w_6655 , w_6656 , w_6657 , w_6658 , w_6659 , w_6660 , w_6661 , 
		w_6662 , w_6663 , w_6664 , w_6665 , w_6666 , w_6667 , w_6668 , w_6669 , w_6670 , w_6671 , 
		w_6672 , w_6673 , w_6674 , w_6675 , w_6676 , w_6677 , w_6678 , w_6679 , w_6680 , w_6681 , 
		w_6682 , w_6683 , w_6684 , w_6685 , w_6686 , w_6687 , w_6688 , w_6689 , w_6690 , w_6691 , 
		w_6692 , w_6693 , w_6694 , w_6695 , w_6696 , w_6697 , w_6698 , w_6699 , w_6700 , w_6701 , 
		w_6702 , w_6703 , w_6704 , w_6705 , w_6706 , w_6707 , w_6708 , w_6709 , w_6710 , w_6711 , 
		w_6712 , w_6713 , w_6714 , w_6715 , w_6716 , w_6717 , w_6718 , w_6719 , w_6720 , w_6721 , 
		w_6722 , w_6723 , w_6724 , w_6725 , w_6726 , w_6727 , w_6728 , w_6729 , w_6730 , w_6731 , 
		w_6732 , w_6733 , w_6734 , w_6735 , w_6736 , w_6737 , w_6738 , w_6739 , w_6740 , w_6741 , 
		w_6742 , w_6743 , w_6744 , w_6745 , w_6746 , w_6747 , w_6748 , w_6749 , w_6750 , w_6751 , 
		w_6752 , w_6753 , w_6754 , w_6755 , w_6756 , w_6757 , w_6758 , w_6759 , w_6760 , w_6761 , 
		w_6762 , w_6763 , w_6764 , w_6765 , w_6766 , w_6767 , w_6768 , w_6769 , w_6770 , w_6771 , 
		w_6772 , w_6773 , w_6774 , w_6775 , w_6776 , w_6777 , w_6778 , w_6779 , w_6780 , w_6781 , 
		w_6782 , w_6783 , w_6784 , w_6785 , w_6786 , w_6787 , w_6788 , w_6789 , w_6790 , w_6791 , 
		w_6792 , w_6793 , w_6794 , w_6795 , w_6796 , w_6797 , w_6798 , w_6799 , w_6800 , w_6801 , 
		w_6802 , w_6803 , w_6804 , w_6805 , w_6806 , w_6807 , w_6808 , w_6809 , w_6810 , w_6811 , 
		w_6812 , w_6813 , w_6814 , w_6815 , w_6816 , w_6817 , w_6818 , w_6819 , w_6820 , w_6821 , 
		w_6822 , w_6823 , w_6824 , w_6825 , w_6826 , w_6827 , w_6828 , w_6829 , w_6830 , w_6831 , 
		w_6832 , w_6833 , w_6834 , w_6835 , w_6836 , w_6837 , w_6838 , w_6839 , w_6840 , w_6841 , 
		w_6842 , w_6843 , w_6844 , w_6845 , w_6846 , w_6847 , w_6848 , w_6849 , w_6850 , w_6851 , 
		w_6852 , w_6853 , w_6854 , w_6855 , w_6856 , w_6857 , w_6858 , w_6859 , w_6860 , w_6861 , 
		w_6862 , w_6863 , w_6864 , w_6865 , w_6866 , w_6867 , w_6868 , w_6869 , w_6870 , w_6871 , 
		w_6872 , w_6873 , w_6874 , w_6875 , w_6876 , w_6877 , w_6878 , w_6879 , w_6880 , w_6881 , 
		w_6882 , w_6883 , w_6884 , w_6885 , w_6886 , w_6887 , w_6888 , w_6889 , w_6890 , w_6891 , 
		w_6892 , w_6893 , w_6894 , w_6895 , w_6896 , w_6897 , w_6898 , w_6899 , w_6900 , w_6901 , 
		w_6902 , w_6903 , w_6904 , w_6905 , w_6906 , w_6907 , w_6908 , w_6909 , w_6910 , w_6911 , 
		w_6912 , w_6913 , w_6914 , w_6915 , w_6916 , w_6917 , w_6918 , w_6919 , w_6920 , w_6921 , 
		w_6922 , w_6923 , w_6924 , w_6925 , w_6926 , w_6927 , w_6928 , w_6929 , w_6930 , w_6931 , 
		w_6932 , w_6933 , w_6934 , w_6935 , w_6936 , w_6937 , w_6938 , w_6939 , w_6940 , w_6941 , 
		w_6942 , w_6943 , w_6944 , w_6945 , w_6946 , w_6947 , w_6948 , w_6949 , w_6950 , w_6951 , 
		w_6952 , w_6953 , w_6954 , w_6955 , w_6956 , w_6957 , w_6958 , w_6959 , w_6960 , w_6961 , 
		w_6962 , w_6963 , w_6964 , w_6965 , w_6966 , w_6967 , w_6968 , w_6969 , w_6970 , w_6971 , 
		w_6972 , w_6973 , w_6974 , w_6975 , w_6976 , w_6977 , w_6978 , w_6979 , w_6980 , w_6981 , 
		w_6982 , w_6983 , w_6984 , w_6985 , w_6986 , w_6987 , w_6988 , w_6989 , w_6990 , w_6991 , 
		w_6992 , w_6993 , w_6994 , w_6995 , w_6996 , w_6997 , w_6998 , w_6999 , w_7000 , w_7001 , 
		w_7002 , w_7003 , w_7004 , w_7005 , w_7006 , w_7007 , w_7008 , w_7009 , w_7010 , w_7011 , 
		w_7012 , w_7013 , w_7014 , w_7015 , w_7016 , w_7017 , w_7018 , w_7019 , w_7020 , w_7021 , 
		w_7022 , w_7023 , w_7024 , w_7025 , w_7026 , w_7027 , w_7028 , w_7029 , w_7030 , w_7031 , 
		w_7032 , w_7033 , w_7034 , w_7035 , w_7036 , w_7037 , w_7038 , w_7039 , w_7040 , w_7041 , 
		w_7042 , w_7043 , w_7044 , w_7045 , w_7046 , w_7047 , w_7048 , w_7049 , w_7050 , w_7051 , 
		w_7052 , w_7053 , w_7054 , w_7055 , w_7056 , w_7057 , w_7058 , w_7059 , w_7060 , w_7061 , 
		w_7062 , w_7063 , w_7064 , w_7065 , w_7066 , w_7067 , w_7068 , w_7069 , w_7070 , w_7071 , 
		w_7072 , w_7073 , w_7074 , w_7075 , w_7076 , w_7077 , w_7078 , w_7079 , w_7080 , w_7081 , 
		w_7082 , w_7083 , w_7084 , w_7085 , w_7086 , w_7087 , w_7088 , w_7089 , w_7090 , w_7091 , 
		w_7092 , w_7093 , w_7094 , w_7095 , w_7096 , w_7097 , w_7098 , w_7099 , w_7100 , w_7101 , 
		w_7102 , w_7103 , w_7104 , w_7105 , w_7106 , w_7107 , w_7108 , w_7109 , w_7110 , w_7111 , 
		w_7112 , w_7113 , w_7114 , w_7115 , w_7116 , w_7117 , w_7118 , w_7119 , w_7120 , w_7121 , 
		w_7122 , w_7123 , w_7124 , w_7125 , w_7126 , w_7127 , w_7128 , w_7129 , w_7130 , w_7131 , 
		w_7132 , w_7133 , w_7134 , w_7135 , w_7136 , w_7137 , w_7138 , w_7139 , w_7140 , w_7141 , 
		w_7142 , w_7143 , w_7144 , w_7145 , w_7146 , w_7147 , w_7148 , w_7149 , w_7150 , w_7151 , 
		w_7152 , w_7153 , w_7154 , w_7155 , w_7156 , w_7157 , w_7158 , w_7159 , w_7160 , w_7161 , 
		w_7162 , w_7163 , w_7164 , w_7165 , w_7166 , w_7167 , w_7168 , w_7169 , w_7170 , w_7171 , 
		w_7172 , w_7173 , w_7174 , w_7175 , w_7176 , w_7177 , w_7178 , w_7179 , w_7180 , w_7181 , 
		w_7182 , w_7183 , w_7184 , w_7185 , w_7186 , w_7187 , w_7188 , w_7189 , w_7190 , w_7191 , 
		w_7192 , w_7193 , w_7194 , w_7195 , w_7196 , w_7197 , w_7198 , w_7199 , w_7200 , w_7201 , 
		w_7202 , w_7203 , w_7204 , w_7205 , w_7206 , w_7207 , w_7208 , w_7209 , w_7210 , w_7211 , 
		w_7212 , w_7213 , w_7214 , w_7215 , w_7216 , w_7217 , w_7218 , w_7219 , w_7220 , w_7221 , 
		w_7222 , w_7223 , w_7224 , w_7225 , w_7226 , w_7227 , w_7228 , w_7229 , w_7230 , w_7231 , 
		w_7232 , w_7233 , w_7234 , w_7235 , w_7236 , w_7237 , w_7238 , w_7239 , w_7240 , w_7241 , 
		w_7242 , w_7243 , w_7244 , w_7245 , w_7246 , w_7247 , w_7248 , w_7249 , w_7250 , w_7251 , 
		w_7252 , w_7253 , w_7254 , w_7255 , w_7256 , w_7257 , w_7258 , w_7259 , w_7260 , w_7261 , 
		w_7262 , w_7263 , w_7264 , w_7265 , w_7266 , w_7267 , w_7268 , w_7269 , w_7270 , w_7271 , 
		w_7272 , w_7273 , w_7274 , w_7275 , w_7276 , w_7277 , w_7278 , w_7279 , w_7280 , w_7281 , 
		w_7282 , w_7283 , w_7284 , w_7285 , w_7286 , w_7287 , w_7288 , w_7289 , w_7290 , w_7291 , 
		w_7292 , w_7293 , w_7294 , w_7295 , w_7296 , w_7297 , w_7298 , w_7299 , w_7300 , w_7301 , 
		w_7302 , w_7303 , w_7304 , w_7305 , w_7306 , w_7307 , w_7308 , w_7309 , w_7310 , w_7311 , 
		w_7312 , w_7313 , w_7314 , w_7315 , w_7316 , w_7317 , w_7318 , w_7319 , w_7320 , w_7321 , 
		w_7322 , w_7323 , w_7324 , w_7325 , w_7326 , w_7327 , w_7328 , w_7329 , w_7330 , w_7331 , 
		w_7332 , w_7333 , w_7334 , w_7335 , w_7336 , w_7337 , w_7338 , w_7339 , w_7340 , w_7341 , 
		w_7342 , w_7343 , w_7344 , w_7345 , w_7346 , w_7347 , w_7348 , w_7349 , w_7350 , w_7351 , 
		w_7352 , w_7353 , w_7354 , w_7355 , w_7356 , w_7357 , w_7358 , w_7359 , w_7360 , w_7361 , 
		w_7362 , w_7363 , w_7364 , w_7365 , w_7366 , w_7367 , w_7368 , w_7369 , w_7370 , w_7371 , 
		w_7372 , w_7373 , w_7374 , w_7375 , w_7376 , w_7377 , w_7378 , w_7379 , w_7380 , w_7381 , 
		w_7382 , w_7383 , w_7384 , w_7385 , w_7386 , w_7387 , w_7388 , w_7389 , w_7390 , w_7391 , 
		w_7392 , w_7393 , w_7394 , w_7395 , w_7396 , w_7397 , w_7398 , w_7399 , w_7400 , w_7401 , 
		w_7402 , w_7403 , w_7404 , w_7405 , w_7406 , w_7407 , w_7408 , w_7409 , w_7410 , w_7411 , 
		w_7412 , w_7413 , w_7414 , w_7415 , w_7416 , w_7417 , w_7418 , w_7419 , w_7420 , w_7421 , 
		w_7422 , w_7423 , w_7424 , w_7425 , w_7426 , w_7427 , w_7428 , w_7429 , w_7430 , w_7431 , 
		w_7432 , w_7433 , w_7434 , w_7435 , w_7436 , w_7437 , w_7438 , w_7439 , w_7440 , w_7441 , 
		w_7442 , w_7443 , w_7444 , w_7445 , w_7446 , w_7447 , w_7448 , w_7449 , w_7450 , w_7451 , 
		w_7452 , w_7453 , w_7454 , w_7455 , w_7456 , w_7457 , w_7458 , w_7459 , w_7460 , w_7461 , 
		w_7462 , w_7463 , w_7464 , w_7465 , w_7466 , w_7467 , w_7468 , w_7469 , w_7470 , w_7471 , 
		w_7472 , w_7473 , w_7474 , w_7475 , w_7476 , w_7477 , w_7478 , w_7479 , w_7480 , w_7481 , 
		w_7482 , w_7483 , w_7484 , w_7485 , w_7486 , w_7487 , w_7488 , w_7489 , w_7490 , w_7491 , 
		w_7492 , w_7493 , w_7494 , w_7495 , w_7496 , w_7497 , w_7498 , w_7499 , w_7500 , w_7501 , 
		w_7502 , w_7503 , w_7504 , w_7505 , w_7506 , w_7507 , w_7508 , w_7509 , w_7510 , w_7511 , 
		w_7512 , w_7513 , w_7514 , w_7515 , w_7516 , w_7517 , w_7518 , w_7519 , w_7520 , w_7521 , 
		w_7522 , w_7523 , w_7524 , w_7525 , w_7526 , w_7527 , w_7528 , w_7529 , w_7530 , w_7531 , 
		w_7532 , w_7533 , w_7534 , w_7535 , w_7536 , w_7537 , w_7538 , w_7539 , w_7540 , w_7541 , 
		w_7542 , w_7543 , w_7544 , w_7545 , w_7546 , w_7547 , w_7548 , w_7549 , w_7550 , w_7551 , 
		w_7552 , w_7553 , w_7554 , w_7555 , w_7556 , w_7557 , w_7558 , w_7559 , w_7560 , w_7561 , 
		w_7562 , w_7563 , w_7564 , w_7565 , w_7566 , w_7567 , w_7568 , w_7569 , w_7570 , w_7571 , 
		w_7572 , w_7573 , w_7574 , w_7575 , w_7576 , w_7577 , w_7578 , w_7579 , w_7580 , w_7581 , 
		w_7582 , w_7583 , w_7584 , w_7585 , w_7586 , w_7587 , w_7588 , w_7589 , w_7590 , w_7591 , 
		w_7592 , w_7593 , w_7594 , w_7595 , w_7596 , w_7597 , w_7598 , w_7599 , w_7600 , w_7601 , 
		w_7602 , w_7603 , w_7604 , w_7605 , w_7606 , w_7607 , w_7608 , w_7609 , w_7610 , w_7611 , 
		w_7612 , w_7613 , w_7614 , w_7615 , w_7616 , w_7617 , w_7618 , w_7619 , w_7620 , w_7621 , 
		w_7622 , w_7623 , w_7624 , w_7625 , w_7626 , w_7627 , w_7628 , w_7629 , w_7630 , w_7631 , 
		w_7632 , w_7633 , w_7634 , w_7635 , w_7636 , w_7637 , w_7638 , w_7639 , w_7640 , w_7641 , 
		w_7642 , w_7643 , w_7644 , w_7645 , w_7646 , w_7647 , w_7648 , w_7649 , w_7650 , w_7651 , 
		w_7652 , w_7653 , w_7654 , w_7655 , w_7656 , w_7657 , w_7658 , w_7659 , w_7660 , w_7661 , 
		w_7662 , w_7663 , w_7664 , w_7665 , w_7666 , w_7667 , w_7668 , w_7669 , w_7670 , w_7671 , 
		w_7672 , w_7673 , w_7674 , w_7675 , w_7676 , w_7677 , w_7678 , w_7679 , w_7680 , w_7681 , 
		w_7682 , w_7683 , w_7684 , w_7685 , w_7686 , w_7687 , w_7688 , w_7689 , w_7690 , w_7691 , 
		w_7692 , w_7693 , w_7694 , w_7695 , w_7696 , w_7697 , w_7698 , w_7699 , w_7700 , w_7701 , 
		w_7702 , w_7703 , w_7704 , w_7705 , w_7706 , w_7707 , w_7708 , w_7709 , w_7710 , w_7711 , 
		w_7712 , w_7713 , w_7714 , w_7715 , w_7716 , w_7717 , w_7718 , w_7719 , w_7720 , w_7721 , 
		w_7722 , w_7723 , w_7724 , w_7725 , w_7726 , w_7727 , w_7728 , w_7729 , w_7730 , w_7731 , 
		w_7732 , w_7733 , w_7734 , w_7735 , w_7736 , w_7737 , w_7738 , w_7739 , w_7740 , w_7741 , 
		w_7742 , w_7743 , w_7744 , w_7745 , w_7746 , w_7747 , w_7748 , w_7749 , w_7750 , w_7751 , 
		w_7752 , w_7753 , w_7754 , w_7755 , w_7756 , w_7757 , w_7758 , w_7759 , w_7760 , w_7761 , 
		w_7762 , w_7763 , w_7764 , w_7765 , w_7766 , w_7767 , w_7768 , w_7769 , w_7770 , w_7771 , 
		w_7772 , w_7773 , w_7774 , w_7775 , w_7776 , w_7777 , w_7778 , w_7779 , w_7780 , w_7781 , 
		w_7782 , w_7783 , w_7784 , w_7785 , w_7786 , w_7787 , w_7788 , w_7789 , w_7790 , w_7791 , 
		w_7792 , w_7793 , w_7794 , w_7795 , w_7796 , w_7797 , w_7798 , w_7799 , w_7800 , w_7801 , 
		w_7802 , w_7803 , w_7804 , w_7805 , w_7806 , w_7807 , w_7808 , w_7809 , w_7810 , w_7811 , 
		w_7812 , w_7813 , w_7814 , w_7815 , w_7816 , w_7817 , w_7818 , w_7819 , w_7820 , w_7821 , 
		w_7822 , w_7823 , w_7824 , w_7825 , w_7826 , w_7827 , w_7828 , w_7829 , w_7830 , w_7831 , 
		w_7832 , w_7833 , w_7834 , w_7835 , w_7836 , w_7837 , w_7838 , w_7839 , w_7840 , w_7841 , 
		w_7842 , w_7843 , w_7844 , w_7845 , w_7846 , w_7847 , w_7848 , w_7849 , w_7850 , w_7851 , 
		w_7852 , w_7853 , w_7854 , w_7855 , w_7856 , w_7857 , w_7858 , w_7859 , w_7860 , w_7861 , 
		w_7862 , w_7863 , w_7864 , w_7865 , w_7866 , w_7867 , w_7868 , w_7869 , w_7870 , w_7871 , 
		w_7872 , w_7873 , w_7874 , w_7875 , w_7876 , w_7877 , w_7878 , w_7879 , w_7880 , w_7881 , 
		w_7882 , w_7883 , w_7884 , w_7885 , w_7886 , w_7887 , w_7888 , w_7889 , w_7890 , w_7891 , 
		w_7892 , w_7893 , w_7894 , w_7895 , w_7896 , w_7897 , w_7898 , w_7899 , w_7900 , w_7901 , 
		w_7902 , w_7903 , w_7904 , w_7905 , w_7906 , w_7907 , w_7908 , w_7909 , w_7910 , w_7911 , 
		w_7912 , w_7913 , w_7914 , w_7915 , w_7916 , w_7917 , w_7918 , w_7919 , w_7920 , w_7921 , 
		w_7922 , w_7923 , w_7924 , w_7925 , w_7926 , w_7927 , w_7928 , w_7929 , w_7930 , w_7931 , 
		w_7932 , w_7933 , w_7934 , w_7935 , w_7936 , w_7937 , w_7938 , w_7939 , w_7940 , w_7941 , 
		w_7942 , w_7943 , w_7944 , w_7945 , w_7946 , w_7947 , w_7948 , w_7949 , w_7950 , w_7951 , 
		w_7952 , w_7953 , w_7954 , w_7955 , w_7956 , w_7957 , w_7958 , w_7959 , w_7960 , w_7961 , 
		w_7962 , w_7963 , w_7964 , w_7965 , w_7966 , w_7967 , w_7968 , w_7969 , w_7970 , w_7971 , 
		w_7972 , w_7973 , w_7974 , w_7975 , w_7976 , w_7977 , w_7978 , w_7979 , w_7980 , w_7981 , 
		w_7982 , w_7983 , w_7984 , w_7985 , w_7986 , w_7987 , w_7988 , w_7989 , w_7990 , w_7991 , 
		w_7992 , w_7993 , w_7994 , w_7995 , w_7996 , w_7997 , w_7998 , w_7999 , w_8000 , w_8001 , 
		w_8002 , w_8003 , w_8004 , w_8005 , w_8006 , w_8007 , w_8008 , w_8009 , w_8010 , w_8011 , 
		w_8012 , w_8013 , w_8014 , w_8015 , w_8016 , w_8017 , w_8018 , w_8019 , w_8020 , w_8021 , 
		w_8022 , w_8023 , w_8024 , w_8025 , w_8026 , w_8027 , w_8028 , w_8029 , w_8030 , w_8031 , 
		w_8032 , w_8033 , w_8034 , w_8035 , w_8036 , w_8037 , w_8038 , w_8039 , w_8040 , w_8041 , 
		w_8042 , w_8043 , w_8044 , w_8045 , w_8046 , w_8047 , w_8048 , w_8049 , w_8050 , w_8051 , 
		w_8052 , w_8053 , w_8054 , w_8055 , w_8056 , w_8057 , w_8058 , w_8059 , w_8060 , w_8061 , 
		w_8062 , w_8063 , w_8064 , w_8065 , w_8066 , w_8067 , w_8068 , w_8069 , w_8070 , w_8071 , 
		w_8072 , w_8073 , w_8074 , w_8075 , w_8076 , w_8077 , w_8078 , w_8079 , w_8080 , w_8081 , 
		w_8082 , w_8083 , w_8084 , w_8085 , w_8086 , w_8087 , w_8088 , w_8089 , w_8090 , w_8091 , 
		w_8092 , w_8093 , w_8094 , w_8095 , w_8096 , w_8097 , w_8098 , w_8099 , w_8100 , w_8101 , 
		w_8102 , w_8103 , w_8104 , w_8105 , w_8106 , w_8107 , w_8108 , w_8109 , w_8110 , w_8111 , 
		w_8112 , w_8113 , w_8114 , w_8115 , w_8116 , w_8117 , w_8118 , w_8119 , w_8120 , w_8121 , 
		w_8122 , w_8123 , w_8124 , w_8125 , w_8126 , w_8127 , w_8128 , w_8129 , w_8130 , w_8131 , 
		w_8132 , w_8133 , w_8134 , w_8135 , w_8136 , w_8137 , w_8138 , w_8139 , w_8140 , w_8141 , 
		w_8142 , w_8143 , w_8144 , w_8145 , w_8146 , w_8147 , w_8148 , w_8149 , w_8150 , w_8151 , 
		w_8152 , w_8153 , w_8154 , w_8155 , w_8156 , w_8157 , w_8158 , w_8159 , w_8160 , w_8161 , 
		w_8162 , w_8163 , w_8164 , w_8165 , w_8166 , w_8167 , w_8168 , w_8169 , w_8170 , w_8171 , 
		w_8172 , w_8173 , w_8174 , w_8175 , w_8176 , w_8177 , w_8178 , w_8179 , w_8180 , w_8181 , 
		w_8182 , w_8183 , w_8184 , w_8185 , w_8186 , w_8187 , w_8188 , w_8189 , w_8190 , w_8191 , 
		w_8192 , w_8193 , w_8194 , w_8195 , w_8196 , w_8197 , w_8198 , w_8199 , w_8200 , w_8201 , 
		w_8202 , w_8203 , w_8204 , w_8205 , w_8206 , w_8207 , w_8208 , w_8209 , w_8210 , w_8211 , 
		w_8212 , w_8213 , w_8214 , w_8215 , w_8216 , w_8217 , w_8218 , w_8219 , w_8220 , w_8221 , 
		w_8222 , w_8223 , w_8224 , w_8225 , w_8226 , w_8227 , w_8228 , w_8229 , w_8230 , w_8231 , 
		w_8232 , w_8233 , w_8234 , w_8235 , w_8236 , w_8237 , w_8238 , w_8239 , w_8240 , w_8241 , 
		w_8242 , w_8243 , w_8244 , w_8245 , w_8246 , w_8247 , w_8248 , w_8249 , w_8250 , w_8251 , 
		w_8252 , w_8253 , w_8254 , w_8255 , w_8256 , w_8257 , w_8258 , w_8259 , w_8260 , w_8261 , 
		w_8262 , w_8263 , w_8264 , w_8265 , w_8266 , w_8267 , w_8268 , w_8269 , w_8270 , w_8271 , 
		w_8272 , w_8273 , w_8274 , w_8275 , w_8276 , w_8277 , w_8278 , w_8279 , w_8280 , w_8281 , 
		w_8282 , w_8283 , w_8284 , w_8285 , w_8286 , w_8287 , w_8288 , w_8289 , w_8290 , w_8291 , 
		w_8292 , w_8293 , w_8294 , w_8295 , w_8296 , w_8297 , w_8298 , w_8299 , w_8300 , w_8301 , 
		w_8302 , w_8303 , w_8304 , w_8305 , w_8306 , w_8307 , w_8308 , w_8309 , w_8310 , w_8311 , 
		w_8312 , w_8313 , w_8314 , w_8315 , w_8316 , w_8317 , w_8318 , w_8319 , w_8320 , w_8321 , 
		w_8322 , w_8323 , w_8324 , w_8325 , w_8326 , w_8327 , w_8328 , w_8329 , w_8330 , w_8331 , 
		w_8332 , w_8333 , w_8334 , w_8335 , w_8336 , w_8337 , w_8338 , w_8339 , w_8340 , w_8341 , 
		w_8342 , w_8343 , w_8344 , w_8345 , w_8346 , w_8347 , w_8348 , w_8349 , w_8350 , w_8351 , 
		w_8352 , w_8353 , w_8354 , w_8355 , w_8356 , w_8357 , w_8358 , w_8359 , w_8360 , w_8361 , 
		w_8362 , w_8363 , w_8364 , w_8365 , w_8366 , w_8367 , w_8368 , w_8369 , w_8370 , w_8371 , 
		w_8372 , w_8373 , w_8374 , w_8375 , w_8376 , w_8377 , w_8378 , w_8379 , w_8380 , w_8381 , 
		w_8382 , w_8383 , w_8384 , w_8385 , w_8386 , w_8387 , w_8388 , w_8389 , w_8390 , w_8391 , 
		w_8392 , w_8393 , w_8394 , w_8395 , w_8396 , w_8397 , w_8398 , w_8399 , w_8400 , w_8401 , 
		w_8402 , w_8403 , w_8404 , w_8405 , w_8406 , w_8407 , w_8408 , w_8409 , w_8410 , w_8411 , 
		w_8412 , w_8413 , w_8414 , w_8415 , w_8416 , w_8417 , w_8418 , w_8419 , w_8420 , w_8421 , 
		w_8422 , w_8423 , w_8424 , w_8425 , w_8426 , w_8427 , w_8428 , w_8429 , w_8430 , w_8431 , 
		w_8432 , w_8433 , w_8434 , w_8435 , w_8436 , w_8437 , w_8438 , w_8439 , w_8440 , w_8441 , 
		w_8442 , w_8443 , w_8444 , w_8445 , w_8446 , w_8447 , w_8448 , w_8449 , w_8450 , w_8451 , 
		w_8452 , w_8453 , w_8454 , w_8455 , w_8456 , w_8457 , w_8458 , w_8459 , w_8460 , w_8461 , 
		w_8462 , w_8463 , w_8464 , w_8465 , w_8466 , w_8467 , w_8468 , w_8469 , w_8470 , w_8471 , 
		w_8472 , w_8473 , w_8474 , w_8475 , w_8476 , w_8477 , w_8478 , w_8479 , w_8480 , w_8481 , 
		w_8482 , w_8483 , w_8484 , w_8485 , w_8486 , w_8487 , w_8488 , w_8489 , w_8490 , w_8491 , 
		w_8492 , w_8493 , w_8494 , w_8495 , w_8496 , w_8497 , w_8498 , w_8499 , w_8500 , w_8501 , 
		w_8502 , w_8503 , w_8504 , w_8505 , w_8506 , w_8507 , w_8508 , w_8509 , w_8510 , w_8511 , 
		w_8512 , w_8513 , w_8514 , w_8515 , w_8516 , w_8517 , w_8518 , w_8519 , w_8520 , w_8521 , 
		w_8522 , w_8523 , w_8524 , w_8525 , w_8526 , w_8527 , w_8528 , w_8529 , w_8530 , w_8531 , 
		w_8532 , w_8533 , w_8534 , w_8535 , w_8536 , w_8537 , w_8538 , w_8539 , w_8540 , w_8541 , 
		w_8542 , w_8543 , w_8544 , w_8545 , w_8546 , w_8547 , w_8548 , w_8549 , w_8550 , w_8551 , 
		w_8552 , w_8553 , w_8554 , w_8555 , w_8556 , w_8557 , w_8558 , w_8559 , w_8560 , w_8561 , 
		w_8562 , w_8563 , w_8564 , w_8565 , w_8566 , w_8567 , w_8568 , w_8569 , w_8570 , w_8571 , 
		w_8572 , w_8573 , w_8574 , w_8575 , w_8576 , w_8577 , w_8578 , w_8579 , w_8580 , w_8581 , 
		w_8582 , w_8583 , w_8584 , w_8585 , w_8586 , w_8587 , w_8588 , w_8589 , w_8590 , w_8591 , 
		w_8592 , w_8593 , w_8594 , w_8595 , w_8596 , w_8597 , w_8598 , w_8599 , w_8600 , w_8601 , 
		w_8602 , w_8603 , w_8604 , w_8605 , w_8606 , w_8607 , w_8608 , w_8609 , w_8610 , w_8611 , 
		w_8612 , w_8613 , w_8614 , w_8615 , w_8616 , w_8617 , w_8618 , w_8619 , w_8620 , w_8621 , 
		w_8622 , w_8623 , w_8624 , w_8625 , w_8626 , w_8627 , w_8628 , w_8629 , w_8630 , w_8631 , 
		w_8632 , w_8633 , w_8634 , w_8635 , w_8636 , w_8637 , w_8638 , w_8639 , w_8640 , w_8641 , 
		w_8642 , w_8643 , w_8644 , w_8645 , w_8646 , w_8647 , w_8648 , w_8649 , w_8650 , w_8651 , 
		w_8652 , w_8653 , w_8654 , w_8655 , w_8656 , w_8657 , w_8658 , w_8659 , w_8660 , w_8661 , 
		w_8662 , w_8663 , w_8664 , w_8665 , w_8666 , w_8667 , w_8668 , w_8669 , w_8670 , w_8671 , 
		w_8672 , w_8673 , w_8674 , w_8675 , w_8676 , w_8677 , w_8678 , w_8679 , w_8680 , w_8681 , 
		w_8682 , w_8683 , w_8684 , w_8685 , w_8686 , w_8687 , w_8688 , w_8689 , w_8690 , w_8691 , 
		w_8692 , w_8693 , w_8694 , w_8695 , w_8696 , w_8697 , w_8698 , w_8699 , w_8700 , w_8701 , 
		w_8702 , w_8703 , w_8704 , w_8705 , w_8706 , w_8707 , w_8708 , w_8709 , w_8710 , w_8711 , 
		w_8712 , w_8713 , w_8714 , w_8715 , w_8716 , w_8717 , w_8718 , w_8719 , w_8720 , w_8721 , 
		w_8722 , w_8723 , w_8724 , w_8725 , w_8726 , w_8727 , w_8728 , w_8729 , w_8730 , w_8731 , 
		w_8732 , w_8733 , w_8734 , w_8735 , w_8736 , w_8737 , w_8738 , w_8739 , w_8740 , w_8741 , 
		w_8742 , w_8743 , w_8744 , w_8745 , w_8746 , w_8747 , w_8748 , w_8749 , w_8750 , w_8751 , 
		w_8752 , w_8753 , w_8754 , w_8755 , w_8756 , w_8757 , w_8758 , w_8759 , w_8760 , w_8761 , 
		w_8762 , w_8763 , w_8764 , w_8765 , w_8766 , w_8767 , w_8768 , w_8769 , w_8770 , w_8771 , 
		w_8772 , w_8773 , w_8774 , w_8775 , w_8776 , w_8777 , w_8778 , w_8779 , w_8780 , w_8781 , 
		w_8782 , w_8783 , w_8784 , w_8785 , w_8786 , w_8787 , w_8788 , w_8789 , w_8790 , w_8791 , 
		w_8792 , w_8793 , w_8794 , w_8795 , w_8796 , w_8797 , w_8798 , w_8799 , w_8800 , w_8801 , 
		w_8802 , w_8803 , w_8804 , w_8805 , w_8806 , w_8807 , w_8808 , w_8809 , w_8810 , w_8811 , 
		w_8812 , w_8813 , w_8814 , w_8815 , w_8816 , w_8817 , w_8818 , w_8819 , w_8820 , w_8821 , 
		w_8822 , w_8823 , w_8824 , w_8825 , w_8826 , w_8827 , w_8828 , w_8829 , w_8830 , w_8831 , 
		w_8832 , w_8833 , w_8834 , w_8835 , w_8836 , w_8837 , w_8838 , w_8839 , w_8840 , w_8841 , 
		w_8842 , w_8843 , w_8844 , w_8845 , w_8846 , w_8847 , w_8848 , w_8849 , w_8850 , w_8851 , 
		w_8852 , w_8853 , w_8854 , w_8855 , w_8856 , w_8857 , w_8858 , w_8859 , w_8860 , w_8861 , 
		w_8862 , w_8863 , w_8864 , w_8865 , w_8866 , w_8867 , w_8868 , w_8869 , w_8870 , w_8871 , 
		w_8872 , w_8873 , w_8874 , w_8875 , w_8876 , w_8877 , w_8878 , w_8879 , w_8880 , w_8881 , 
		w_8882 , w_8883 , w_8884 , w_8885 , w_8886 , w_8887 , w_8888 , w_8889 , w_8890 , w_8891 , 
		w_8892 , w_8893 , w_8894 , w_8895 , w_8896 , w_8897 , w_8898 , w_8899 , w_8900 , w_8901 , 
		w_8902 , w_8903 , w_8904 , w_8905 , w_8906 , w_8907 , w_8908 , w_8909 , w_8910 , w_8911 , 
		w_8912 , w_8913 , w_8914 , w_8915 , w_8916 , w_8917 , w_8918 , w_8919 , w_8920 , w_8921 , 
		w_8922 , w_8923 , w_8924 , w_8925 , w_8926 , w_8927 , w_8928 , w_8929 , w_8930 , w_8931 , 
		w_8932 , w_8933 , w_8934 , w_8935 , w_8936 , w_8937 , w_8938 , w_8939 , w_8940 , w_8941 , 
		w_8942 , w_8943 , w_8944 , w_8945 , w_8946 , w_8947 , w_8948 , w_8949 , w_8950 , w_8951 , 
		w_8952 , w_8953 , w_8954 , w_8955 , w_8956 , w_8957 , w_8958 , w_8959 , w_8960 , w_8961 , 
		w_8962 , w_8963 , w_8964 , w_8965 , w_8966 , w_8967 , w_8968 , w_8969 , w_8970 , w_8971 , 
		w_8972 , w_8973 , w_8974 , w_8975 , w_8976 , w_8977 , w_8978 , w_8979 , w_8980 , w_8981 , 
		w_8982 , w_8983 , w_8984 , w_8985 , w_8986 , w_8987 , w_8988 , w_8989 , w_8990 , w_8991 , 
		w_8992 , w_8993 , w_8994 , w_8995 , w_8996 , w_8997 , w_8998 , w_8999 , w_9000 , w_9001 , 
		w_9002 , w_9003 , w_9004 , w_9005 , w_9006 , w_9007 , w_9008 , w_9009 , w_9010 , w_9011 , 
		w_9012 , w_9013 , w_9014 , w_9015 , w_9016 , w_9017 , w_9018 , w_9019 , w_9020 , w_9021 , 
		w_9022 , w_9023 , w_9024 , w_9025 , w_9026 , w_9027 , w_9028 , w_9029 , w_9030 , w_9031 , 
		w_9032 , w_9033 , w_9034 , w_9035 , w_9036 , w_9037 , w_9038 , w_9039 , w_9040 , w_9041 , 
		w_9042 , w_9043 , w_9044 , w_9045 , w_9046 , w_9047 , w_9048 , w_9049 , w_9050 , w_9051 , 
		w_9052 , w_9053 , w_9054 , w_9055 , w_9056 , w_9057 , w_9058 , w_9059 , w_9060 , w_9061 , 
		w_9062 , w_9063 , w_9064 , w_9065 , w_9066 , w_9067 , w_9068 , w_9069 , w_9070 , w_9071 , 
		w_9072 , w_9073 , w_9074 , w_9075 , w_9076 , w_9077 , w_9078 , w_9079 , w_9080 , w_9081 , 
		w_9082 , w_9083 , w_9084 , w_9085 , w_9086 , w_9087 , w_9088 , w_9089 , w_9090 , w_9091 , 
		w_9092 , w_9093 , w_9094 , w_9095 , w_9096 , w_9097 , w_9098 , w_9099 , w_9100 , w_9101 , 
		w_9102 , w_9103 , w_9104 , w_9105 , w_9106 , w_9107 , w_9108 , w_9109 , w_9110 , w_9111 , 
		w_9112 , w_9113 , w_9114 , w_9115 , w_9116 , w_9117 , w_9118 , w_9119 , w_9120 , w_9121 , 
		w_9122 , w_9123 , w_9124 , w_9125 , w_9126 , w_9127 , w_9128 , w_9129 , w_9130 , w_9131 , 
		w_9132 , w_9133 , w_9134 , w_9135 , w_9136 , w_9137 , w_9138 , w_9139 , w_9140 , w_9141 , 
		w_9142 , w_9143 , w_9144 , w_9145 , w_9146 , w_9147 , w_9148 , w_9149 , w_9150 , w_9151 , 
		w_9152 , w_9153 , w_9154 , w_9155 , w_9156 , w_9157 , w_9158 , w_9159 , w_9160 , w_9161 , 
		w_9162 , w_9163 , w_9164 , w_9165 , w_9166 , w_9167 , w_9168 , w_9169 , w_9170 , w_9171 , 
		w_9172 , w_9173 , w_9174 , w_9175 , w_9176 , w_9177 , w_9178 , w_9179 , w_9180 , w_9181 , 
		w_9182 , w_9183 , w_9184 , w_9185 , w_9186 , w_9187 , w_9188 , w_9189 , w_9190 , w_9191 , 
		w_9192 , w_9193 , w_9194 , w_9195 , w_9196 , w_9197 , w_9198 , w_9199 , w_9200 , w_9201 , 
		w_9202 , w_9203 , w_9204 , w_9205 , w_9206 , w_9207 , w_9208 , w_9209 , w_9210 , w_9211 , 
		w_9212 , w_9213 , w_9214 , w_9215 , w_9216 , w_9217 , w_9218 , w_9219 , w_9220 , w_9221 , 
		w_9222 , w_9223 , w_9224 , w_9225 , w_9226 , w_9227 , w_9228 , w_9229 , w_9230 , w_9231 , 
		w_9232 , w_9233 , w_9234 , w_9235 , w_9236 , w_9237 , w_9238 , w_9239 , w_9240 , w_9241 , 
		w_9242 , w_9243 , w_9244 , w_9245 , w_9246 , w_9247 , w_9248 , w_9249 , w_9250 , w_9251 , 
		w_9252 , w_9253 , w_9254 , w_9255 , w_9256 , w_9257 , w_9258 , w_9259 , w_9260 , w_9261 , 
		w_9262 , w_9263 , w_9264 , w_9265 , w_9266 , w_9267 , w_9268 , w_9269 , w_9270 , w_9271 , 
		w_9272 , w_9273 , w_9274 , w_9275 , w_9276 , w_9277 , w_9278 , w_9279 , w_9280 , w_9281 , 
		w_9282 , w_9283 , w_9284 , w_9285 , w_9286 , w_9287 , w_9288 , w_9289 , w_9290 , w_9291 , 
		w_9292 , w_9293 , w_9294 , w_9295 , w_9296 , w_9297 , w_9298 , w_9299 , w_9300 , w_9301 , 
		w_9302 , w_9303 , w_9304 , w_9305 , w_9306 , w_9307 , w_9308 , w_9309 , w_9310 , w_9311 , 
		w_9312 , w_9313 , w_9314 , w_9315 , w_9316 , w_9317 , w_9318 , w_9319 , w_9320 , w_9321 , 
		w_9322 , w_9323 , w_9324 , w_9325 , w_9326 , w_9327 , w_9328 , w_9329 , w_9330 , w_9331 , 
		w_9332 , w_9333 , w_9334 , w_9335 , w_9336 , w_9337 , w_9338 , w_9339 , w_9340 , w_9341 , 
		w_9342 , w_9343 , w_9344 , w_9345 , w_9346 , w_9347 , w_9348 , w_9349 , w_9350 , w_9351 , 
		w_9352 , w_9353 , w_9354 , w_9355 , w_9356 , w_9357 , w_9358 , w_9359 , w_9360 , w_9361 , 
		w_9362 , w_9363 , w_9364 , w_9365 , w_9366 , w_9367 , w_9368 , w_9369 , w_9370 , w_9371 , 
		w_9372 , w_9373 , w_9374 , w_9375 , w_9376 , w_9377 , w_9378 , w_9379 , w_9380 , w_9381 , 
		w_9382 , w_9383 , w_9384 , w_9385 , w_9386 , w_9387 , w_9388 , w_9389 , w_9390 , w_9391 , 
		w_9392 , w_9393 , w_9394 , w_9395 , w_9396 , w_9397 , w_9398 , w_9399 , w_9400 , w_9401 , 
		w_9402 , w_9403 , w_9404 , w_9405 , w_9406 , w_9407 , w_9408 , w_9409 , w_9410 , w_9411 , 
		w_9412 , w_9413 , w_9414 , w_9415 , w_9416 , w_9417 , w_9418 , w_9419 , w_9420 , w_9421 , 
		w_9422 , w_9423 , w_9424 , w_9425 , w_9426 , w_9427 , w_9428 , w_9429 , w_9430 , w_9431 , 
		w_9432 , w_9433 , w_9434 , w_9435 , w_9436 , w_9437 , w_9438 , w_9439 , w_9440 , w_9441 , 
		w_9442 , w_9443 , w_9444 , w_9445 , w_9446 , w_9447 , w_9448 , w_9449 , w_9450 , w_9451 , 
		w_9452 , w_9453 , w_9454 , w_9455 , w_9456 , w_9457 , w_9458 , w_9459 , w_9460 , w_9461 , 
		w_9462 , w_9463 , w_9464 , w_9465 , w_9466 , w_9467 , w_9468 , w_9469 , w_9470 , w_9471 , 
		w_9472 , w_9473 , w_9474 , w_9475 , w_9476 , w_9477 , w_9478 , w_9479 , w_9480 , w_9481 , 
		w_9482 , w_9483 , w_9484 , w_9485 , w_9486 , w_9487 , w_9488 , w_9489 , w_9490 , w_9491 , 
		w_9492 , w_9493 , w_9494 , w_9495 , w_9496 , w_9497 , w_9498 , w_9499 , w_9500 , w_9501 , 
		w_9502 , w_9503 , w_9504 , w_9505 , w_9506 , w_9507 , w_9508 , w_9509 , w_9510 , w_9511 , 
		w_9512 , w_9513 , w_9514 , w_9515 , w_9516 , w_9517 , w_9518 , w_9519 , w_9520 , w_9521 , 
		w_9522 , w_9523 , w_9524 , w_9525 , w_9526 , w_9527 , w_9528 , w_9529 , w_9530 , w_9531 , 
		w_9532 , w_9533 , w_9534 , w_9535 , w_9536 , w_9537 , w_9538 , w_9539 , w_9540 , w_9541 , 
		w_9542 , w_9543 , w_9544 , w_9545 , w_9546 , w_9547 , w_9548 , w_9549 , w_9550 , w_9551 , 
		w_9552 , w_9553 , w_9554 , w_9555 , w_9556 , w_9557 , w_9558 , w_9559 , w_9560 , w_9561 , 
		w_9562 , w_9563 , w_9564 , w_9565 , w_9566 , w_9567 , w_9568 , w_9569 , w_9570 , w_9571 , 
		w_9572 , w_9573 , w_9574 , w_9575 , w_9576 , w_9577 , w_9578 , w_9579 , w_9580 , w_9581 , 
		w_9582 , w_9583 , w_9584 , w_9585 , w_9586 , w_9587 , w_9588 , w_9589 , w_9590 , w_9591 , 
		w_9592 , w_9593 , w_9594 , w_9595 , w_9596 , w_9597 , w_9598 , w_9599 , w_9600 , w_9601 , 
		w_9602 , w_9603 , w_9604 , w_9605 , w_9606 , w_9607 , w_9608 , w_9609 , w_9610 , w_9611 , 
		w_9612 , w_9613 , w_9614 , w_9615 , w_9616 , w_9617 , w_9618 , w_9619 , w_9620 , w_9621 , 
		w_9622 , w_9623 , w_9624 , w_9625 , w_9626 , w_9627 , w_9628 , w_9629 , w_9630 , w_9631 , 
		w_9632 , w_9633 , w_9634 , w_9635 , w_9636 , w_9637 , w_9638 , w_9639 , w_9640 , w_9641 , 
		w_9642 , w_9643 , w_9644 , w_9645 , w_9646 , w_9647 , w_9648 , w_9649 , w_9650 , w_9651 , 
		w_9652 , w_9653 , w_9654 , w_9655 , w_9656 , w_9657 , w_9658 , w_9659 , w_9660 , w_9661 , 
		w_9662 , w_9663 , w_9664 , w_9665 , w_9666 , w_9667 , w_9668 , w_9669 , w_9670 , w_9671 , 
		w_9672 , w_9673 , w_9674 , w_9675 , w_9676 , w_9677 , w_9678 , w_9679 , w_9680 , w_9681 ;
buf ( \o[31]_b1 , \4468_Z[31]_b1 );
buf ( \o[31]_b0 , \4468_Z[31]_b0 );
buf ( \o[30]_b1 , \4470_Z[30]_b1 );
buf ( \o[30]_b0 , \4470_Z[30]_b0 );
buf ( \o[29]_b1 , \4472_Z[29]_b1 );
buf ( \o[29]_b0 , \4472_Z[29]_b0 );
buf ( \o[28]_b1 , \4474_Z[28]_b1 );
buf ( \o[28]_b0 , \4474_Z[28]_b0 );
buf ( \o[27]_b1 , \4476_Z[27]_b1 );
buf ( \o[27]_b0 , \4476_Z[27]_b0 );
buf ( \o[26]_b1 , \4478_Z[26]_b1 );
buf ( \o[26]_b0 , \4478_Z[26]_b0 );
buf ( \o[25]_b1 , \4480_Z[25]_b1 );
buf ( \o[25]_b0 , \4480_Z[25]_b0 );
buf ( \o[24]_b1 , \4482_Z[24]_b1 );
buf ( \o[24]_b0 , \4482_Z[24]_b0 );
buf ( \o[23]_b1 , \4484_Z[23]_b1 );
buf ( \o[23]_b0 , \4484_Z[23]_b0 );
buf ( \o[22]_b1 , \4486_Z[22]_b1 );
buf ( \o[22]_b0 , \4486_Z[22]_b0 );
buf ( \o[21]_b1 , \4488_Z[21]_b1 );
buf ( \o[21]_b0 , \4488_Z[21]_b0 );
buf ( \o[20]_b1 , \4490_Z[20]_b1 );
buf ( \o[20]_b0 , \4490_Z[20]_b0 );
buf ( \o[19]_b1 , \4492_Z[19]_b1 );
buf ( \o[19]_b0 , \4492_Z[19]_b0 );
buf ( \o[18]_b1 , \4494_Z[18]_b1 );
buf ( \o[18]_b0 , \4494_Z[18]_b0 );
buf ( \o[17]_b1 , \4496_Z[17]_b1 );
buf ( \o[17]_b0 , \4496_Z[17]_b0 );
buf ( \o[16]_b1 , \4498_Z[16]_b1 );
buf ( \o[16]_b0 , \4498_Z[16]_b0 );
buf ( \o[15]_b1 , \4500_Z[15]_b1 );
buf ( \o[15]_b0 , \4500_Z[15]_b0 );
buf ( \o[14]_b1 , \4502_Z[14]_b1 );
buf ( \o[14]_b0 , \4502_Z[14]_b0 );
buf ( \o[13]_b1 , \4504_Z[13]_b1 );
buf ( \o[13]_b0 , \4504_Z[13]_b0 );
buf ( \o[12]_b1 , \4506_Z[12]_b1 );
buf ( \o[12]_b0 , \4506_Z[12]_b0 );
buf ( \o[11]_b1 , \4508_Z[11]_b1 );
buf ( \o[11]_b0 , \4508_Z[11]_b0 );
buf ( \o[10]_b1 , \4510_Z[10]_b1 );
buf ( \o[10]_b0 , \4510_Z[10]_b0 );
buf ( \o[9]_b1 , \4512_Z[9]_b1 );
buf ( \o[9]_b0 , \4512_Z[9]_b0 );
buf ( \o[8]_b1 , \4514_Z[8]_b1 );
buf ( \o[8]_b0 , \4514_Z[8]_b0 );
buf ( \o[7]_b1 , \4516_Z[7]_b1 );
buf ( \o[7]_b0 , \4516_Z[7]_b0 );
buf ( \o[6]_b1 , \4518_Z[6]_b1 );
buf ( \o[6]_b0 , \4518_Z[6]_b0 );
buf ( \o[5]_b1 , \4520_Z[5]_b1 );
buf ( \o[5]_b0 , \4520_Z[5]_b0 );
buf ( \o[4]_b1 , \4522_Z[4]_b1 );
buf ( \o[4]_b0 , \4522_Z[4]_b0 );
buf ( \o[3]_b1 , \4524_Z[3]_b1 );
buf ( \o[3]_b0 , \4524_Z[3]_b0 );
buf ( \o[2]_b1 , \4526_Z[2]_b1 );
buf ( \o[2]_b0 , \4526_Z[2]_b0 );
buf ( \o[1]_b1 , \4528_Z[1]_b1 );
buf ( \o[1]_b0 , \4528_Z[1]_b0 );
buf ( \o[0]_b1 , \4530_Z[0]_b1 );
buf ( \o[0]_b0 , \4530_Z[0]_b0 );
buf ( \156_A[0]_b1 , \a[0]_b1 );
buf ( \156_A[0]_b0 , \a[0]_b0 );
buf ( \157_B[0]_b1 , \b[0]_b1 );
buf ( \157_B[0]_b0 , \b[0]_b0 );
or ( \158_b1 , \156_A[0]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_0 );
and ( \158_b0 , \156_A[0]_b0 , w_1 );
and ( w_0 , w_1 , \157_B[0]_b0 );
buf ( \159_Z[0]_b1 , \158_b1 );
buf ( \159_Z[0]_b0 , \158_b0 );
buf ( \160_b1 , \159_Z[0]_b1 );
not ( \160_b1 , w_2 );
not ( \160_b0 , w_3 );
and ( w_2 , w_3 , \159_Z[0]_b0 );
buf ( \161_A[1]_b1 , \a[1]_b1 );
buf ( \161_A[1]_b0 , \a[1]_b0 );
or ( \162_b1 , \161_A[1]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_4 );
and ( \162_b0 , \161_A[1]_b0 , w_5 );
and ( w_4 , w_5 , \157_B[0]_b0 );
buf ( \163_B[1]_b1 , \b[1]_b1 );
buf ( \163_B[1]_b0 , \b[1]_b0 );
or ( \164_b1 , \156_A[0]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_6 );
and ( \164_b0 , \156_A[0]_b0 , w_7 );
and ( w_6 , w_7 , \163_B[1]_b0 );
or ( \165_b1 , \162_b1 , \164_b1 );
xor ( \165_b0 , \162_b0 , w_8 );
not ( w_8 , w_9 );
and ( w_9 , \164_b1 , \164_b0 );
buf ( \166_Z[1]_b1 , \165_b1 );
buf ( \166_Z[1]_b0 , \165_b0 );
buf ( \167_A[2]_b1 , \a[2]_b1 );
buf ( \167_A[2]_b0 , \a[2]_b0 );
or ( \168_b1 , \167_A[2]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_10 );
and ( \168_b0 , \167_A[2]_b0 , w_11 );
and ( w_10 , w_11 , \157_B[0]_b0 );
or ( \169_b1 , \161_A[1]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_12 );
and ( \169_b0 , \161_A[1]_b0 , w_13 );
and ( w_12 , w_13 , \163_B[1]_b0 );
or ( \170_b1 , \168_b1 , \169_b1 );
xor ( \170_b0 , \168_b0 , w_14 );
not ( w_14 , w_15 );
and ( w_15 , \169_b1 , \169_b0 );
or ( \171_b1 , \162_b1 , \164_b1 );
not ( \164_b1 , w_16 );
and ( \171_b0 , \162_b0 , w_17 );
and ( w_16 , w_17 , \164_b0 );
or ( \172_b1 , \170_b1 , \171_b1 );
xor ( \172_b0 , \170_b0 , w_18 );
not ( w_18 , w_19 );
and ( w_19 , \171_b1 , \171_b0 );
buf ( \173_B[2]_b1 , \b[2]_b1 );
buf ( \173_B[2]_b0 , \b[2]_b0 );
or ( \174_b1 , \156_A[0]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_20 );
and ( \174_b0 , \156_A[0]_b0 , w_21 );
and ( w_20 , w_21 , \173_B[2]_b0 );
or ( \175_b1 , \172_b1 , \174_b1 );
xor ( \175_b0 , \172_b0 , w_22 );
not ( w_22 , w_23 );
and ( w_23 , \174_b1 , \174_b0 );
buf ( \176_Z[2]_b1 , \175_b1 );
buf ( \176_Z[2]_b0 , \175_b0 );
buf ( \177_A[3]_b1 , \a[3]_b1 );
buf ( \177_A[3]_b0 , \a[3]_b0 );
or ( \178_b1 , \177_A[3]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_24 );
and ( \178_b0 , \177_A[3]_b0 , w_25 );
and ( w_24 , w_25 , \157_B[0]_b0 );
or ( \179_b1 , \167_A[2]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_26 );
and ( \179_b0 , \167_A[2]_b0 , w_27 );
and ( w_26 , w_27 , \163_B[1]_b0 );
or ( \180_b1 , \178_b1 , \179_b1 );
xor ( \180_b0 , \178_b0 , w_28 );
not ( w_28 , w_29 );
and ( w_29 , \179_b1 , \179_b0 );
or ( \181_b1 , \168_b1 , \169_b1 );
not ( \169_b1 , w_30 );
and ( \181_b0 , \168_b0 , w_31 );
and ( w_30 , w_31 , \169_b0 );
or ( \182_b1 , \170_b1 , \171_b1 );
not ( \171_b1 , w_32 );
and ( \182_b0 , \170_b0 , w_33 );
and ( w_32 , w_33 , \171_b0 );
or ( \183_b1 , \181_b1 , w_34 );
or ( \183_b0 , \181_b0 , \182_b0 );
not ( \182_b0 , w_35 );
and ( w_35 , w_34 , \182_b1 );
or ( \184_b1 , \180_b1 , \183_b1 );
xor ( \184_b0 , \180_b0 , w_36 );
not ( w_36 , w_37 );
and ( w_37 , \183_b1 , \183_b0 );
or ( \185_b1 , \161_A[1]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_38 );
and ( \185_b0 , \161_A[1]_b0 , w_39 );
and ( w_38 , w_39 , \173_B[2]_b0 );
or ( \186_b1 , \184_b1 , \185_b1 );
xor ( \186_b0 , \184_b0 , w_40 );
not ( w_40 , w_41 );
and ( w_41 , \185_b1 , \185_b0 );
or ( \187_b1 , \172_b1 , \174_b1 );
not ( \174_b1 , w_42 );
and ( \187_b0 , \172_b0 , w_43 );
and ( w_42 , w_43 , \174_b0 );
or ( \188_b1 , \186_b1 , \187_b1 );
xor ( \188_b0 , \186_b0 , w_44 );
not ( w_44 , w_45 );
and ( w_45 , \187_b1 , \187_b0 );
buf ( \189_B[3]_b1 , \b[3]_b1 );
buf ( \189_B[3]_b0 , \b[3]_b0 );
or ( \190_b1 , \156_A[0]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_46 );
and ( \190_b0 , \156_A[0]_b0 , w_47 );
and ( w_46 , w_47 , \189_B[3]_b0 );
or ( \191_b1 , \188_b1 , \190_b1 );
xor ( \191_b0 , \188_b0 , w_48 );
not ( w_48 , w_49 );
and ( w_49 , \190_b1 , \190_b0 );
buf ( \192_Z[3]_b1 , \191_b1 );
buf ( \192_Z[3]_b0 , \191_b0 );
buf ( \193_A[4]_b1 , \a[4]_b1 );
buf ( \193_A[4]_b0 , \a[4]_b0 );
or ( \194_b1 , \193_A[4]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_50 );
and ( \194_b0 , \193_A[4]_b0 , w_51 );
and ( w_50 , w_51 , \157_B[0]_b0 );
or ( \195_b1 , \177_A[3]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_52 );
and ( \195_b0 , \177_A[3]_b0 , w_53 );
and ( w_52 , w_53 , \163_B[1]_b0 );
or ( \196_b1 , \194_b1 , \195_b1 );
xor ( \196_b0 , \194_b0 , w_54 );
not ( w_54 , w_55 );
and ( w_55 , \195_b1 , \195_b0 );
or ( \197_b1 , \178_b1 , \179_b1 );
not ( \179_b1 , w_56 );
and ( \197_b0 , \178_b0 , w_57 );
and ( w_56 , w_57 , \179_b0 );
or ( \198_b1 , \180_b1 , \183_b1 );
not ( \183_b1 , w_58 );
and ( \198_b0 , \180_b0 , w_59 );
and ( w_58 , w_59 , \183_b0 );
or ( \199_b1 , \197_b1 , w_60 );
or ( \199_b0 , \197_b0 , \198_b0 );
not ( \198_b0 , w_61 );
and ( w_61 , w_60 , \198_b1 );
or ( \200_b1 , \196_b1 , \199_b1 );
xor ( \200_b0 , \196_b0 , w_62 );
not ( w_62 , w_63 );
and ( w_63 , \199_b1 , \199_b0 );
or ( \201_b1 , \167_A[2]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_64 );
and ( \201_b0 , \167_A[2]_b0 , w_65 );
and ( w_64 , w_65 , \173_B[2]_b0 );
or ( \202_b1 , \200_b1 , \201_b1 );
xor ( \202_b0 , \200_b0 , w_66 );
not ( w_66 , w_67 );
and ( w_67 , \201_b1 , \201_b0 );
or ( \203_b1 , \184_b1 , \185_b1 );
not ( \185_b1 , w_68 );
and ( \203_b0 , \184_b0 , w_69 );
and ( w_68 , w_69 , \185_b0 );
or ( \204_b1 , \186_b1 , \187_b1 );
not ( \187_b1 , w_70 );
and ( \204_b0 , \186_b0 , w_71 );
and ( w_70 , w_71 , \187_b0 );
or ( \205_b1 , \203_b1 , w_72 );
or ( \205_b0 , \203_b0 , \204_b0 );
not ( \204_b0 , w_73 );
and ( w_73 , w_72 , \204_b1 );
or ( \206_b1 , \202_b1 , \205_b1 );
xor ( \206_b0 , \202_b0 , w_74 );
not ( w_74 , w_75 );
and ( w_75 , \205_b1 , \205_b0 );
or ( \207_b1 , \161_A[1]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_76 );
and ( \207_b0 , \161_A[1]_b0 , w_77 );
and ( w_76 , w_77 , \189_B[3]_b0 );
or ( \208_b1 , \206_b1 , \207_b1 );
xor ( \208_b0 , \206_b0 , w_78 );
not ( w_78 , w_79 );
and ( w_79 , \207_b1 , \207_b0 );
or ( \209_b1 , \188_b1 , \190_b1 );
not ( \190_b1 , w_80 );
and ( \209_b0 , \188_b0 , w_81 );
and ( w_80 , w_81 , \190_b0 );
or ( \210_b1 , \208_b1 , \209_b1 );
xor ( \210_b0 , \208_b0 , w_82 );
not ( w_82 , w_83 );
and ( w_83 , \209_b1 , \209_b0 );
buf ( \211_B[4]_b1 , \b[4]_b1 );
buf ( \211_B[4]_b0 , \b[4]_b0 );
or ( \212_b1 , \156_A[0]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_84 );
and ( \212_b0 , \156_A[0]_b0 , w_85 );
and ( w_84 , w_85 , \211_B[4]_b0 );
or ( \213_b1 , \210_b1 , \212_b1 );
xor ( \213_b0 , \210_b0 , w_86 );
not ( w_86 , w_87 );
and ( w_87 , \212_b1 , \212_b0 );
buf ( \214_Z[4]_b1 , \213_b1 );
buf ( \214_Z[4]_b0 , \213_b0 );
buf ( \215_A[5]_b1 , \a[5]_b1 );
buf ( \215_A[5]_b0 , \a[5]_b0 );
or ( \216_b1 , \215_A[5]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_88 );
and ( \216_b0 , \215_A[5]_b0 , w_89 );
and ( w_88 , w_89 , \157_B[0]_b0 );
or ( \217_b1 , \193_A[4]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_90 );
and ( \217_b0 , \193_A[4]_b0 , w_91 );
and ( w_90 , w_91 , \163_B[1]_b0 );
or ( \218_b1 , \216_b1 , \217_b1 );
xor ( \218_b0 , \216_b0 , w_92 );
not ( w_92 , w_93 );
and ( w_93 , \217_b1 , \217_b0 );
or ( \219_b1 , \194_b1 , \195_b1 );
not ( \195_b1 , w_94 );
and ( \219_b0 , \194_b0 , w_95 );
and ( w_94 , w_95 , \195_b0 );
or ( \220_b1 , \196_b1 , \199_b1 );
not ( \199_b1 , w_96 );
and ( \220_b0 , \196_b0 , w_97 );
and ( w_96 , w_97 , \199_b0 );
or ( \221_b1 , \219_b1 , w_98 );
or ( \221_b0 , \219_b0 , \220_b0 );
not ( \220_b0 , w_99 );
and ( w_99 , w_98 , \220_b1 );
or ( \222_b1 , \218_b1 , \221_b1 );
xor ( \222_b0 , \218_b0 , w_100 );
not ( w_100 , w_101 );
and ( w_101 , \221_b1 , \221_b0 );
or ( \223_b1 , \177_A[3]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_102 );
and ( \223_b0 , \177_A[3]_b0 , w_103 );
and ( w_102 , w_103 , \173_B[2]_b0 );
or ( \224_b1 , \222_b1 , \223_b1 );
xor ( \224_b0 , \222_b0 , w_104 );
not ( w_104 , w_105 );
and ( w_105 , \223_b1 , \223_b0 );
or ( \225_b1 , \200_b1 , \201_b1 );
not ( \201_b1 , w_106 );
and ( \225_b0 , \200_b0 , w_107 );
and ( w_106 , w_107 , \201_b0 );
or ( \226_b1 , \202_b1 , \205_b1 );
not ( \205_b1 , w_108 );
and ( \226_b0 , \202_b0 , w_109 );
and ( w_108 , w_109 , \205_b0 );
or ( \227_b1 , \225_b1 , w_110 );
or ( \227_b0 , \225_b0 , \226_b0 );
not ( \226_b0 , w_111 );
and ( w_111 , w_110 , \226_b1 );
or ( \228_b1 , \224_b1 , \227_b1 );
xor ( \228_b0 , \224_b0 , w_112 );
not ( w_112 , w_113 );
and ( w_113 , \227_b1 , \227_b0 );
or ( \229_b1 , \167_A[2]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_114 );
and ( \229_b0 , \167_A[2]_b0 , w_115 );
and ( w_114 , w_115 , \189_B[3]_b0 );
or ( \230_b1 , \228_b1 , \229_b1 );
xor ( \230_b0 , \228_b0 , w_116 );
not ( w_116 , w_117 );
and ( w_117 , \229_b1 , \229_b0 );
or ( \231_b1 , \206_b1 , \207_b1 );
not ( \207_b1 , w_118 );
and ( \231_b0 , \206_b0 , w_119 );
and ( w_118 , w_119 , \207_b0 );
or ( \232_b1 , \208_b1 , \209_b1 );
not ( \209_b1 , w_120 );
and ( \232_b0 , \208_b0 , w_121 );
and ( w_120 , w_121 , \209_b0 );
or ( \233_b1 , \231_b1 , w_122 );
or ( \233_b0 , \231_b0 , \232_b0 );
not ( \232_b0 , w_123 );
and ( w_123 , w_122 , \232_b1 );
or ( \234_b1 , \230_b1 , \233_b1 );
xor ( \234_b0 , \230_b0 , w_124 );
not ( w_124 , w_125 );
and ( w_125 , \233_b1 , \233_b0 );
or ( \235_b1 , \161_A[1]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_126 );
and ( \235_b0 , \161_A[1]_b0 , w_127 );
and ( w_126 , w_127 , \211_B[4]_b0 );
or ( \236_b1 , \234_b1 , \235_b1 );
xor ( \236_b0 , \234_b0 , w_128 );
not ( w_128 , w_129 );
and ( w_129 , \235_b1 , \235_b0 );
or ( \237_b1 , \210_b1 , \212_b1 );
not ( \212_b1 , w_130 );
and ( \237_b0 , \210_b0 , w_131 );
and ( w_130 , w_131 , \212_b0 );
or ( \238_b1 , \236_b1 , \237_b1 );
xor ( \238_b0 , \236_b0 , w_132 );
not ( w_132 , w_133 );
and ( w_133 , \237_b1 , \237_b0 );
buf ( \239_B[5]_b1 , \b[5]_b1 );
buf ( \239_B[5]_b0 , \b[5]_b0 );
or ( \240_b1 , \156_A[0]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_134 );
and ( \240_b0 , \156_A[0]_b0 , w_135 );
and ( w_134 , w_135 , \239_B[5]_b0 );
or ( \241_b1 , \238_b1 , \240_b1 );
xor ( \241_b0 , \238_b0 , w_136 );
not ( w_136 , w_137 );
and ( w_137 , \240_b1 , \240_b0 );
buf ( \242_Z[5]_b1 , \241_b1 );
buf ( \242_Z[5]_b0 , \241_b0 );
buf ( \243_A[6]_b1 , \a[6]_b1 );
buf ( \243_A[6]_b0 , \a[6]_b0 );
or ( \244_b1 , \243_A[6]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_138 );
and ( \244_b0 , \243_A[6]_b0 , w_139 );
and ( w_138 , w_139 , \157_B[0]_b0 );
or ( \245_b1 , \215_A[5]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_140 );
and ( \245_b0 , \215_A[5]_b0 , w_141 );
and ( w_140 , w_141 , \163_B[1]_b0 );
or ( \246_b1 , \244_b1 , \245_b1 );
xor ( \246_b0 , \244_b0 , w_142 );
not ( w_142 , w_143 );
and ( w_143 , \245_b1 , \245_b0 );
or ( \247_b1 , \216_b1 , \217_b1 );
not ( \217_b1 , w_144 );
and ( \247_b0 , \216_b0 , w_145 );
and ( w_144 , w_145 , \217_b0 );
or ( \248_b1 , \218_b1 , \221_b1 );
not ( \221_b1 , w_146 );
and ( \248_b0 , \218_b0 , w_147 );
and ( w_146 , w_147 , \221_b0 );
or ( \249_b1 , \247_b1 , w_148 );
or ( \249_b0 , \247_b0 , \248_b0 );
not ( \248_b0 , w_149 );
and ( w_149 , w_148 , \248_b1 );
or ( \250_b1 , \246_b1 , \249_b1 );
xor ( \250_b0 , \246_b0 , w_150 );
not ( w_150 , w_151 );
and ( w_151 , \249_b1 , \249_b0 );
or ( \251_b1 , \193_A[4]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_152 );
and ( \251_b0 , \193_A[4]_b0 , w_153 );
and ( w_152 , w_153 , \173_B[2]_b0 );
or ( \252_b1 , \250_b1 , \251_b1 );
xor ( \252_b0 , \250_b0 , w_154 );
not ( w_154 , w_155 );
and ( w_155 , \251_b1 , \251_b0 );
or ( \253_b1 , \222_b1 , \223_b1 );
not ( \223_b1 , w_156 );
and ( \253_b0 , \222_b0 , w_157 );
and ( w_156 , w_157 , \223_b0 );
or ( \254_b1 , \224_b1 , \227_b1 );
not ( \227_b1 , w_158 );
and ( \254_b0 , \224_b0 , w_159 );
and ( w_158 , w_159 , \227_b0 );
or ( \255_b1 , \253_b1 , w_160 );
or ( \255_b0 , \253_b0 , \254_b0 );
not ( \254_b0 , w_161 );
and ( w_161 , w_160 , \254_b1 );
or ( \256_b1 , \252_b1 , \255_b1 );
xor ( \256_b0 , \252_b0 , w_162 );
not ( w_162 , w_163 );
and ( w_163 , \255_b1 , \255_b0 );
or ( \257_b1 , \177_A[3]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_164 );
and ( \257_b0 , \177_A[3]_b0 , w_165 );
and ( w_164 , w_165 , \189_B[3]_b0 );
or ( \258_b1 , \256_b1 , \257_b1 );
xor ( \258_b0 , \256_b0 , w_166 );
not ( w_166 , w_167 );
and ( w_167 , \257_b1 , \257_b0 );
or ( \259_b1 , \228_b1 , \229_b1 );
not ( \229_b1 , w_168 );
and ( \259_b0 , \228_b0 , w_169 );
and ( w_168 , w_169 , \229_b0 );
or ( \260_b1 , \230_b1 , \233_b1 );
not ( \233_b1 , w_170 );
and ( \260_b0 , \230_b0 , w_171 );
and ( w_170 , w_171 , \233_b0 );
or ( \261_b1 , \259_b1 , w_172 );
or ( \261_b0 , \259_b0 , \260_b0 );
not ( \260_b0 , w_173 );
and ( w_173 , w_172 , \260_b1 );
or ( \262_b1 , \258_b1 , \261_b1 );
xor ( \262_b0 , \258_b0 , w_174 );
not ( w_174 , w_175 );
and ( w_175 , \261_b1 , \261_b0 );
or ( \263_b1 , \167_A[2]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_176 );
and ( \263_b0 , \167_A[2]_b0 , w_177 );
and ( w_176 , w_177 , \211_B[4]_b0 );
or ( \264_b1 , \262_b1 , \263_b1 );
xor ( \264_b0 , \262_b0 , w_178 );
not ( w_178 , w_179 );
and ( w_179 , \263_b1 , \263_b0 );
or ( \265_b1 , \234_b1 , \235_b1 );
not ( \235_b1 , w_180 );
and ( \265_b0 , \234_b0 , w_181 );
and ( w_180 , w_181 , \235_b0 );
or ( \266_b1 , \236_b1 , \237_b1 );
not ( \237_b1 , w_182 );
and ( \266_b0 , \236_b0 , w_183 );
and ( w_182 , w_183 , \237_b0 );
or ( \267_b1 , \265_b1 , w_184 );
or ( \267_b0 , \265_b0 , \266_b0 );
not ( \266_b0 , w_185 );
and ( w_185 , w_184 , \266_b1 );
or ( \268_b1 , \264_b1 , \267_b1 );
xor ( \268_b0 , \264_b0 , w_186 );
not ( w_186 , w_187 );
and ( w_187 , \267_b1 , \267_b0 );
or ( \269_b1 , \161_A[1]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_188 );
and ( \269_b0 , \161_A[1]_b0 , w_189 );
and ( w_188 , w_189 , \239_B[5]_b0 );
or ( \270_b1 , \268_b1 , \269_b1 );
xor ( \270_b0 , \268_b0 , w_190 );
not ( w_190 , w_191 );
and ( w_191 , \269_b1 , \269_b0 );
or ( \271_b1 , \238_b1 , \240_b1 );
not ( \240_b1 , w_192 );
and ( \271_b0 , \238_b0 , w_193 );
and ( w_192 , w_193 , \240_b0 );
or ( \272_b1 , \270_b1 , \271_b1 );
xor ( \272_b0 , \270_b0 , w_194 );
not ( w_194 , w_195 );
and ( w_195 , \271_b1 , \271_b0 );
buf ( \273_B[6]_b1 , \b[6]_b1 );
buf ( \273_B[6]_b0 , \b[6]_b0 );
or ( \274_b1 , \156_A[0]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_196 );
and ( \274_b0 , \156_A[0]_b0 , w_197 );
and ( w_196 , w_197 , \273_B[6]_b0 );
or ( \275_b1 , \272_b1 , \274_b1 );
xor ( \275_b0 , \272_b0 , w_198 );
not ( w_198 , w_199 );
and ( w_199 , \274_b1 , \274_b0 );
buf ( \276_Z[6]_b1 , \275_b1 );
buf ( \276_Z[6]_b0 , \275_b0 );
buf ( \277_A[7]_b1 , \a[7]_b1 );
buf ( \277_A[7]_b0 , \a[7]_b0 );
or ( \278_b1 , \277_A[7]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_200 );
and ( \278_b0 , \277_A[7]_b0 , w_201 );
and ( w_200 , w_201 , \157_B[0]_b0 );
or ( \279_b1 , \243_A[6]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_202 );
and ( \279_b0 , \243_A[6]_b0 , w_203 );
and ( w_202 , w_203 , \163_B[1]_b0 );
or ( \280_b1 , \278_b1 , \279_b1 );
xor ( \280_b0 , \278_b0 , w_204 );
not ( w_204 , w_205 );
and ( w_205 , \279_b1 , \279_b0 );
or ( \281_b1 , \244_b1 , \245_b1 );
not ( \245_b1 , w_206 );
and ( \281_b0 , \244_b0 , w_207 );
and ( w_206 , w_207 , \245_b0 );
or ( \282_b1 , \246_b1 , \249_b1 );
not ( \249_b1 , w_208 );
and ( \282_b0 , \246_b0 , w_209 );
and ( w_208 , w_209 , \249_b0 );
or ( \283_b1 , \281_b1 , w_210 );
or ( \283_b0 , \281_b0 , \282_b0 );
not ( \282_b0 , w_211 );
and ( w_211 , w_210 , \282_b1 );
or ( \284_b1 , \280_b1 , \283_b1 );
xor ( \284_b0 , \280_b0 , w_212 );
not ( w_212 , w_213 );
and ( w_213 , \283_b1 , \283_b0 );
or ( \285_b1 , \215_A[5]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_214 );
and ( \285_b0 , \215_A[5]_b0 , w_215 );
and ( w_214 , w_215 , \173_B[2]_b0 );
or ( \286_b1 , \284_b1 , \285_b1 );
xor ( \286_b0 , \284_b0 , w_216 );
not ( w_216 , w_217 );
and ( w_217 , \285_b1 , \285_b0 );
or ( \287_b1 , \250_b1 , \251_b1 );
not ( \251_b1 , w_218 );
and ( \287_b0 , \250_b0 , w_219 );
and ( w_218 , w_219 , \251_b0 );
or ( \288_b1 , \252_b1 , \255_b1 );
not ( \255_b1 , w_220 );
and ( \288_b0 , \252_b0 , w_221 );
and ( w_220 , w_221 , \255_b0 );
or ( \289_b1 , \287_b1 , w_222 );
or ( \289_b0 , \287_b0 , \288_b0 );
not ( \288_b0 , w_223 );
and ( w_223 , w_222 , \288_b1 );
or ( \290_b1 , \286_b1 , \289_b1 );
xor ( \290_b0 , \286_b0 , w_224 );
not ( w_224 , w_225 );
and ( w_225 , \289_b1 , \289_b0 );
or ( \291_b1 , \193_A[4]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_226 );
and ( \291_b0 , \193_A[4]_b0 , w_227 );
and ( w_226 , w_227 , \189_B[3]_b0 );
or ( \292_b1 , \290_b1 , \291_b1 );
xor ( \292_b0 , \290_b0 , w_228 );
not ( w_228 , w_229 );
and ( w_229 , \291_b1 , \291_b0 );
or ( \293_b1 , \256_b1 , \257_b1 );
not ( \257_b1 , w_230 );
and ( \293_b0 , \256_b0 , w_231 );
and ( w_230 , w_231 , \257_b0 );
or ( \294_b1 , \258_b1 , \261_b1 );
not ( \261_b1 , w_232 );
and ( \294_b0 , \258_b0 , w_233 );
and ( w_232 , w_233 , \261_b0 );
or ( \295_b1 , \293_b1 , w_234 );
or ( \295_b0 , \293_b0 , \294_b0 );
not ( \294_b0 , w_235 );
and ( w_235 , w_234 , \294_b1 );
or ( \296_b1 , \292_b1 , \295_b1 );
xor ( \296_b0 , \292_b0 , w_236 );
not ( w_236 , w_237 );
and ( w_237 , \295_b1 , \295_b0 );
or ( \297_b1 , \177_A[3]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_238 );
and ( \297_b0 , \177_A[3]_b0 , w_239 );
and ( w_238 , w_239 , \211_B[4]_b0 );
or ( \298_b1 , \296_b1 , \297_b1 );
xor ( \298_b0 , \296_b0 , w_240 );
not ( w_240 , w_241 );
and ( w_241 , \297_b1 , \297_b0 );
or ( \299_b1 , \262_b1 , \263_b1 );
not ( \263_b1 , w_242 );
and ( \299_b0 , \262_b0 , w_243 );
and ( w_242 , w_243 , \263_b0 );
or ( \300_b1 , \264_b1 , \267_b1 );
not ( \267_b1 , w_244 );
and ( \300_b0 , \264_b0 , w_245 );
and ( w_244 , w_245 , \267_b0 );
or ( \301_b1 , \299_b1 , w_246 );
or ( \301_b0 , \299_b0 , \300_b0 );
not ( \300_b0 , w_247 );
and ( w_247 , w_246 , \300_b1 );
or ( \302_b1 , \298_b1 , \301_b1 );
xor ( \302_b0 , \298_b0 , w_248 );
not ( w_248 , w_249 );
and ( w_249 , \301_b1 , \301_b0 );
or ( \303_b1 , \167_A[2]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_250 );
and ( \303_b0 , \167_A[2]_b0 , w_251 );
and ( w_250 , w_251 , \239_B[5]_b0 );
or ( \304_b1 , \302_b1 , \303_b1 );
xor ( \304_b0 , \302_b0 , w_252 );
not ( w_252 , w_253 );
and ( w_253 , \303_b1 , \303_b0 );
or ( \305_b1 , \268_b1 , \269_b1 );
not ( \269_b1 , w_254 );
and ( \305_b0 , \268_b0 , w_255 );
and ( w_254 , w_255 , \269_b0 );
or ( \306_b1 , \270_b1 , \271_b1 );
not ( \271_b1 , w_256 );
and ( \306_b0 , \270_b0 , w_257 );
and ( w_256 , w_257 , \271_b0 );
or ( \307_b1 , \305_b1 , w_258 );
or ( \307_b0 , \305_b0 , \306_b0 );
not ( \306_b0 , w_259 );
and ( w_259 , w_258 , \306_b1 );
or ( \308_b1 , \304_b1 , \307_b1 );
xor ( \308_b0 , \304_b0 , w_260 );
not ( w_260 , w_261 );
and ( w_261 , \307_b1 , \307_b0 );
or ( \309_b1 , \161_A[1]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_262 );
and ( \309_b0 , \161_A[1]_b0 , w_263 );
and ( w_262 , w_263 , \273_B[6]_b0 );
or ( \310_b1 , \308_b1 , \309_b1 );
xor ( \310_b0 , \308_b0 , w_264 );
not ( w_264 , w_265 );
and ( w_265 , \309_b1 , \309_b0 );
or ( \311_b1 , \272_b1 , \274_b1 );
not ( \274_b1 , w_266 );
and ( \311_b0 , \272_b0 , w_267 );
and ( w_266 , w_267 , \274_b0 );
or ( \312_b1 , \310_b1 , \311_b1 );
xor ( \312_b0 , \310_b0 , w_268 );
not ( w_268 , w_269 );
and ( w_269 , \311_b1 , \311_b0 );
buf ( \313_B[7]_b1 , \b[7]_b1 );
buf ( \313_B[7]_b0 , \b[7]_b0 );
or ( \314_b1 , \156_A[0]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_270 );
and ( \314_b0 , \156_A[0]_b0 , w_271 );
and ( w_270 , w_271 , \313_B[7]_b0 );
or ( \315_b1 , \312_b1 , \314_b1 );
xor ( \315_b0 , \312_b0 , w_272 );
not ( w_272 , w_273 );
and ( w_273 , \314_b1 , \314_b0 );
buf ( \316_Z[7]_b1 , \315_b1 );
buf ( \316_Z[7]_b0 , \315_b0 );
buf ( \317_A[8]_b1 , \a[8]_b1 );
buf ( \317_A[8]_b0 , \a[8]_b0 );
or ( \318_b1 , \317_A[8]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_274 );
and ( \318_b0 , \317_A[8]_b0 , w_275 );
and ( w_274 , w_275 , \157_B[0]_b0 );
or ( \319_b1 , \277_A[7]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_276 );
and ( \319_b0 , \277_A[7]_b0 , w_277 );
and ( w_276 , w_277 , \163_B[1]_b0 );
or ( \320_b1 , \318_b1 , \319_b1 );
xor ( \320_b0 , \318_b0 , w_278 );
not ( w_278 , w_279 );
and ( w_279 , \319_b1 , \319_b0 );
or ( \321_b1 , \278_b1 , \279_b1 );
not ( \279_b1 , w_280 );
and ( \321_b0 , \278_b0 , w_281 );
and ( w_280 , w_281 , \279_b0 );
or ( \322_b1 , \280_b1 , \283_b1 );
not ( \283_b1 , w_282 );
and ( \322_b0 , \280_b0 , w_283 );
and ( w_282 , w_283 , \283_b0 );
or ( \323_b1 , \321_b1 , w_284 );
or ( \323_b0 , \321_b0 , \322_b0 );
not ( \322_b0 , w_285 );
and ( w_285 , w_284 , \322_b1 );
or ( \324_b1 , \320_b1 , \323_b1 );
xor ( \324_b0 , \320_b0 , w_286 );
not ( w_286 , w_287 );
and ( w_287 , \323_b1 , \323_b0 );
or ( \325_b1 , \243_A[6]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_288 );
and ( \325_b0 , \243_A[6]_b0 , w_289 );
and ( w_288 , w_289 , \173_B[2]_b0 );
or ( \326_b1 , \324_b1 , \325_b1 );
xor ( \326_b0 , \324_b0 , w_290 );
not ( w_290 , w_291 );
and ( w_291 , \325_b1 , \325_b0 );
or ( \327_b1 , \284_b1 , \285_b1 );
not ( \285_b1 , w_292 );
and ( \327_b0 , \284_b0 , w_293 );
and ( w_292 , w_293 , \285_b0 );
or ( \328_b1 , \286_b1 , \289_b1 );
not ( \289_b1 , w_294 );
and ( \328_b0 , \286_b0 , w_295 );
and ( w_294 , w_295 , \289_b0 );
or ( \329_b1 , \327_b1 , w_296 );
or ( \329_b0 , \327_b0 , \328_b0 );
not ( \328_b0 , w_297 );
and ( w_297 , w_296 , \328_b1 );
or ( \330_b1 , \326_b1 , \329_b1 );
xor ( \330_b0 , \326_b0 , w_298 );
not ( w_298 , w_299 );
and ( w_299 , \329_b1 , \329_b0 );
or ( \331_b1 , \215_A[5]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_300 );
and ( \331_b0 , \215_A[5]_b0 , w_301 );
and ( w_300 , w_301 , \189_B[3]_b0 );
or ( \332_b1 , \330_b1 , \331_b1 );
xor ( \332_b0 , \330_b0 , w_302 );
not ( w_302 , w_303 );
and ( w_303 , \331_b1 , \331_b0 );
or ( \333_b1 , \290_b1 , \291_b1 );
not ( \291_b1 , w_304 );
and ( \333_b0 , \290_b0 , w_305 );
and ( w_304 , w_305 , \291_b0 );
or ( \334_b1 , \292_b1 , \295_b1 );
not ( \295_b1 , w_306 );
and ( \334_b0 , \292_b0 , w_307 );
and ( w_306 , w_307 , \295_b0 );
or ( \335_b1 , \333_b1 , w_308 );
or ( \335_b0 , \333_b0 , \334_b0 );
not ( \334_b0 , w_309 );
and ( w_309 , w_308 , \334_b1 );
or ( \336_b1 , \332_b1 , \335_b1 );
xor ( \336_b0 , \332_b0 , w_310 );
not ( w_310 , w_311 );
and ( w_311 , \335_b1 , \335_b0 );
or ( \337_b1 , \193_A[4]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_312 );
and ( \337_b0 , \193_A[4]_b0 , w_313 );
and ( w_312 , w_313 , \211_B[4]_b0 );
or ( \338_b1 , \336_b1 , \337_b1 );
xor ( \338_b0 , \336_b0 , w_314 );
not ( w_314 , w_315 );
and ( w_315 , \337_b1 , \337_b0 );
or ( \339_b1 , \296_b1 , \297_b1 );
not ( \297_b1 , w_316 );
and ( \339_b0 , \296_b0 , w_317 );
and ( w_316 , w_317 , \297_b0 );
or ( \340_b1 , \298_b1 , \301_b1 );
not ( \301_b1 , w_318 );
and ( \340_b0 , \298_b0 , w_319 );
and ( w_318 , w_319 , \301_b0 );
or ( \341_b1 , \339_b1 , w_320 );
or ( \341_b0 , \339_b0 , \340_b0 );
not ( \340_b0 , w_321 );
and ( w_321 , w_320 , \340_b1 );
or ( \342_b1 , \338_b1 , \341_b1 );
xor ( \342_b0 , \338_b0 , w_322 );
not ( w_322 , w_323 );
and ( w_323 , \341_b1 , \341_b0 );
or ( \343_b1 , \177_A[3]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_324 );
and ( \343_b0 , \177_A[3]_b0 , w_325 );
and ( w_324 , w_325 , \239_B[5]_b0 );
or ( \344_b1 , \342_b1 , \343_b1 );
xor ( \344_b0 , \342_b0 , w_326 );
not ( w_326 , w_327 );
and ( w_327 , \343_b1 , \343_b0 );
or ( \345_b1 , \302_b1 , \303_b1 );
not ( \303_b1 , w_328 );
and ( \345_b0 , \302_b0 , w_329 );
and ( w_328 , w_329 , \303_b0 );
or ( \346_b1 , \304_b1 , \307_b1 );
not ( \307_b1 , w_330 );
and ( \346_b0 , \304_b0 , w_331 );
and ( w_330 , w_331 , \307_b0 );
or ( \347_b1 , \345_b1 , w_332 );
or ( \347_b0 , \345_b0 , \346_b0 );
not ( \346_b0 , w_333 );
and ( w_333 , w_332 , \346_b1 );
or ( \348_b1 , \344_b1 , \347_b1 );
xor ( \348_b0 , \344_b0 , w_334 );
not ( w_334 , w_335 );
and ( w_335 , \347_b1 , \347_b0 );
or ( \349_b1 , \167_A[2]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_336 );
and ( \349_b0 , \167_A[2]_b0 , w_337 );
and ( w_336 , w_337 , \273_B[6]_b0 );
or ( \350_b1 , \348_b1 , \349_b1 );
xor ( \350_b0 , \348_b0 , w_338 );
not ( w_338 , w_339 );
and ( w_339 , \349_b1 , \349_b0 );
or ( \351_b1 , \308_b1 , \309_b1 );
not ( \309_b1 , w_340 );
and ( \351_b0 , \308_b0 , w_341 );
and ( w_340 , w_341 , \309_b0 );
or ( \352_b1 , \310_b1 , \311_b1 );
not ( \311_b1 , w_342 );
and ( \352_b0 , \310_b0 , w_343 );
and ( w_342 , w_343 , \311_b0 );
or ( \353_b1 , \351_b1 , w_344 );
or ( \353_b0 , \351_b0 , \352_b0 );
not ( \352_b0 , w_345 );
and ( w_345 , w_344 , \352_b1 );
or ( \354_b1 , \350_b1 , \353_b1 );
xor ( \354_b0 , \350_b0 , w_346 );
not ( w_346 , w_347 );
and ( w_347 , \353_b1 , \353_b0 );
or ( \355_b1 , \161_A[1]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_348 );
and ( \355_b0 , \161_A[1]_b0 , w_349 );
and ( w_348 , w_349 , \313_B[7]_b0 );
or ( \356_b1 , \354_b1 , \355_b1 );
xor ( \356_b0 , \354_b0 , w_350 );
not ( w_350 , w_351 );
and ( w_351 , \355_b1 , \355_b0 );
or ( \357_b1 , \312_b1 , \314_b1 );
not ( \314_b1 , w_352 );
and ( \357_b0 , \312_b0 , w_353 );
and ( w_352 , w_353 , \314_b0 );
or ( \358_b1 , \356_b1 , \357_b1 );
xor ( \358_b0 , \356_b0 , w_354 );
not ( w_354 , w_355 );
and ( w_355 , \357_b1 , \357_b0 );
buf ( \359_B[8]_b1 , \b[8]_b1 );
buf ( \359_B[8]_b0 , \b[8]_b0 );
or ( \360_b1 , \156_A[0]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_356 );
and ( \360_b0 , \156_A[0]_b0 , w_357 );
and ( w_356 , w_357 , \359_B[8]_b0 );
or ( \361_b1 , \358_b1 , \360_b1 );
xor ( \361_b0 , \358_b0 , w_358 );
not ( w_358 , w_359 );
and ( w_359 , \360_b1 , \360_b0 );
buf ( \362_Z[8]_b1 , \361_b1 );
buf ( \362_Z[8]_b0 , \361_b0 );
buf ( \363_A[9]_b1 , \a[9]_b1 );
buf ( \363_A[9]_b0 , \a[9]_b0 );
or ( \364_b1 , \363_A[9]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_360 );
and ( \364_b0 , \363_A[9]_b0 , w_361 );
and ( w_360 , w_361 , \157_B[0]_b0 );
or ( \365_b1 , \317_A[8]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_362 );
and ( \365_b0 , \317_A[8]_b0 , w_363 );
and ( w_362 , w_363 , \163_B[1]_b0 );
or ( \366_b1 , \364_b1 , \365_b1 );
xor ( \366_b0 , \364_b0 , w_364 );
not ( w_364 , w_365 );
and ( w_365 , \365_b1 , \365_b0 );
or ( \367_b1 , \318_b1 , \319_b1 );
not ( \319_b1 , w_366 );
and ( \367_b0 , \318_b0 , w_367 );
and ( w_366 , w_367 , \319_b0 );
or ( \368_b1 , \320_b1 , \323_b1 );
not ( \323_b1 , w_368 );
and ( \368_b0 , \320_b0 , w_369 );
and ( w_368 , w_369 , \323_b0 );
or ( \369_b1 , \367_b1 , w_370 );
or ( \369_b0 , \367_b0 , \368_b0 );
not ( \368_b0 , w_371 );
and ( w_371 , w_370 , \368_b1 );
or ( \370_b1 , \366_b1 , \369_b1 );
xor ( \370_b0 , \366_b0 , w_372 );
not ( w_372 , w_373 );
and ( w_373 , \369_b1 , \369_b0 );
or ( \371_b1 , \277_A[7]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_374 );
and ( \371_b0 , \277_A[7]_b0 , w_375 );
and ( w_374 , w_375 , \173_B[2]_b0 );
or ( \372_b1 , \370_b1 , \371_b1 );
xor ( \372_b0 , \370_b0 , w_376 );
not ( w_376 , w_377 );
and ( w_377 , \371_b1 , \371_b0 );
or ( \373_b1 , \324_b1 , \325_b1 );
not ( \325_b1 , w_378 );
and ( \373_b0 , \324_b0 , w_379 );
and ( w_378 , w_379 , \325_b0 );
or ( \374_b1 , \326_b1 , \329_b1 );
not ( \329_b1 , w_380 );
and ( \374_b0 , \326_b0 , w_381 );
and ( w_380 , w_381 , \329_b0 );
or ( \375_b1 , \373_b1 , w_382 );
or ( \375_b0 , \373_b0 , \374_b0 );
not ( \374_b0 , w_383 );
and ( w_383 , w_382 , \374_b1 );
or ( \376_b1 , \372_b1 , \375_b1 );
xor ( \376_b0 , \372_b0 , w_384 );
not ( w_384 , w_385 );
and ( w_385 , \375_b1 , \375_b0 );
or ( \377_b1 , \243_A[6]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_386 );
and ( \377_b0 , \243_A[6]_b0 , w_387 );
and ( w_386 , w_387 , \189_B[3]_b0 );
or ( \378_b1 , \376_b1 , \377_b1 );
xor ( \378_b0 , \376_b0 , w_388 );
not ( w_388 , w_389 );
and ( w_389 , \377_b1 , \377_b0 );
or ( \379_b1 , \330_b1 , \331_b1 );
not ( \331_b1 , w_390 );
and ( \379_b0 , \330_b0 , w_391 );
and ( w_390 , w_391 , \331_b0 );
or ( \380_b1 , \332_b1 , \335_b1 );
not ( \335_b1 , w_392 );
and ( \380_b0 , \332_b0 , w_393 );
and ( w_392 , w_393 , \335_b0 );
or ( \381_b1 , \379_b1 , w_394 );
or ( \381_b0 , \379_b0 , \380_b0 );
not ( \380_b0 , w_395 );
and ( w_395 , w_394 , \380_b1 );
or ( \382_b1 , \378_b1 , \381_b1 );
xor ( \382_b0 , \378_b0 , w_396 );
not ( w_396 , w_397 );
and ( w_397 , \381_b1 , \381_b0 );
or ( \383_b1 , \215_A[5]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_398 );
and ( \383_b0 , \215_A[5]_b0 , w_399 );
and ( w_398 , w_399 , \211_B[4]_b0 );
or ( \384_b1 , \382_b1 , \383_b1 );
xor ( \384_b0 , \382_b0 , w_400 );
not ( w_400 , w_401 );
and ( w_401 , \383_b1 , \383_b0 );
or ( \385_b1 , \336_b1 , \337_b1 );
not ( \337_b1 , w_402 );
and ( \385_b0 , \336_b0 , w_403 );
and ( w_402 , w_403 , \337_b0 );
or ( \386_b1 , \338_b1 , \341_b1 );
not ( \341_b1 , w_404 );
and ( \386_b0 , \338_b0 , w_405 );
and ( w_404 , w_405 , \341_b0 );
or ( \387_b1 , \385_b1 , w_406 );
or ( \387_b0 , \385_b0 , \386_b0 );
not ( \386_b0 , w_407 );
and ( w_407 , w_406 , \386_b1 );
or ( \388_b1 , \384_b1 , \387_b1 );
xor ( \388_b0 , \384_b0 , w_408 );
not ( w_408 , w_409 );
and ( w_409 , \387_b1 , \387_b0 );
or ( \389_b1 , \193_A[4]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_410 );
and ( \389_b0 , \193_A[4]_b0 , w_411 );
and ( w_410 , w_411 , \239_B[5]_b0 );
or ( \390_b1 , \388_b1 , \389_b1 );
xor ( \390_b0 , \388_b0 , w_412 );
not ( w_412 , w_413 );
and ( w_413 , \389_b1 , \389_b0 );
or ( \391_b1 , \342_b1 , \343_b1 );
not ( \343_b1 , w_414 );
and ( \391_b0 , \342_b0 , w_415 );
and ( w_414 , w_415 , \343_b0 );
or ( \392_b1 , \344_b1 , \347_b1 );
not ( \347_b1 , w_416 );
and ( \392_b0 , \344_b0 , w_417 );
and ( w_416 , w_417 , \347_b0 );
or ( \393_b1 , \391_b1 , w_418 );
or ( \393_b0 , \391_b0 , \392_b0 );
not ( \392_b0 , w_419 );
and ( w_419 , w_418 , \392_b1 );
or ( \394_b1 , \390_b1 , \393_b1 );
xor ( \394_b0 , \390_b0 , w_420 );
not ( w_420 , w_421 );
and ( w_421 , \393_b1 , \393_b0 );
or ( \395_b1 , \177_A[3]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_422 );
and ( \395_b0 , \177_A[3]_b0 , w_423 );
and ( w_422 , w_423 , \273_B[6]_b0 );
or ( \396_b1 , \394_b1 , \395_b1 );
xor ( \396_b0 , \394_b0 , w_424 );
not ( w_424 , w_425 );
and ( w_425 , \395_b1 , \395_b0 );
or ( \397_b1 , \348_b1 , \349_b1 );
not ( \349_b1 , w_426 );
and ( \397_b0 , \348_b0 , w_427 );
and ( w_426 , w_427 , \349_b0 );
or ( \398_b1 , \350_b1 , \353_b1 );
not ( \353_b1 , w_428 );
and ( \398_b0 , \350_b0 , w_429 );
and ( w_428 , w_429 , \353_b0 );
or ( \399_b1 , \397_b1 , w_430 );
or ( \399_b0 , \397_b0 , \398_b0 );
not ( \398_b0 , w_431 );
and ( w_431 , w_430 , \398_b1 );
or ( \400_b1 , \396_b1 , \399_b1 );
xor ( \400_b0 , \396_b0 , w_432 );
not ( w_432 , w_433 );
and ( w_433 , \399_b1 , \399_b0 );
or ( \401_b1 , \167_A[2]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_434 );
and ( \401_b0 , \167_A[2]_b0 , w_435 );
and ( w_434 , w_435 , \313_B[7]_b0 );
or ( \402_b1 , \400_b1 , \401_b1 );
xor ( \402_b0 , \400_b0 , w_436 );
not ( w_436 , w_437 );
and ( w_437 , \401_b1 , \401_b0 );
or ( \403_b1 , \354_b1 , \355_b1 );
not ( \355_b1 , w_438 );
and ( \403_b0 , \354_b0 , w_439 );
and ( w_438 , w_439 , \355_b0 );
or ( \404_b1 , \356_b1 , \357_b1 );
not ( \357_b1 , w_440 );
and ( \404_b0 , \356_b0 , w_441 );
and ( w_440 , w_441 , \357_b0 );
or ( \405_b1 , \403_b1 , w_442 );
or ( \405_b0 , \403_b0 , \404_b0 );
not ( \404_b0 , w_443 );
and ( w_443 , w_442 , \404_b1 );
or ( \406_b1 , \402_b1 , \405_b1 );
xor ( \406_b0 , \402_b0 , w_444 );
not ( w_444 , w_445 );
and ( w_445 , \405_b1 , \405_b0 );
or ( \407_b1 , \161_A[1]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_446 );
and ( \407_b0 , \161_A[1]_b0 , w_447 );
and ( w_446 , w_447 , \359_B[8]_b0 );
or ( \408_b1 , \406_b1 , \407_b1 );
xor ( \408_b0 , \406_b0 , w_448 );
not ( w_448 , w_449 );
and ( w_449 , \407_b1 , \407_b0 );
or ( \409_b1 , \358_b1 , \360_b1 );
not ( \360_b1 , w_450 );
and ( \409_b0 , \358_b0 , w_451 );
and ( w_450 , w_451 , \360_b0 );
or ( \410_b1 , \408_b1 , \409_b1 );
xor ( \410_b0 , \408_b0 , w_452 );
not ( w_452 , w_453 );
and ( w_453 , \409_b1 , \409_b0 );
buf ( \411_B[9]_b1 , \b[9]_b1 );
buf ( \411_B[9]_b0 , \b[9]_b0 );
or ( \412_b1 , \156_A[0]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_454 );
and ( \412_b0 , \156_A[0]_b0 , w_455 );
and ( w_454 , w_455 , \411_B[9]_b0 );
or ( \413_b1 , \410_b1 , \412_b1 );
xor ( \413_b0 , \410_b0 , w_456 );
not ( w_456 , w_457 );
and ( w_457 , \412_b1 , \412_b0 );
buf ( \414_Z[9]_b1 , \413_b1 );
buf ( \414_Z[9]_b0 , \413_b0 );
buf ( \415_A[10]_b1 , \a[10]_b1 );
buf ( \415_A[10]_b0 , \a[10]_b0 );
or ( \416_b1 , \415_A[10]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_458 );
and ( \416_b0 , \415_A[10]_b0 , w_459 );
and ( w_458 , w_459 , \157_B[0]_b0 );
or ( \417_b1 , \363_A[9]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_460 );
and ( \417_b0 , \363_A[9]_b0 , w_461 );
and ( w_460 , w_461 , \163_B[1]_b0 );
or ( \418_b1 , \416_b1 , \417_b1 );
xor ( \418_b0 , \416_b0 , w_462 );
not ( w_462 , w_463 );
and ( w_463 , \417_b1 , \417_b0 );
or ( \419_b1 , \364_b1 , \365_b1 );
not ( \365_b1 , w_464 );
and ( \419_b0 , \364_b0 , w_465 );
and ( w_464 , w_465 , \365_b0 );
or ( \420_b1 , \366_b1 , \369_b1 );
not ( \369_b1 , w_466 );
and ( \420_b0 , \366_b0 , w_467 );
and ( w_466 , w_467 , \369_b0 );
or ( \421_b1 , \419_b1 , w_468 );
or ( \421_b0 , \419_b0 , \420_b0 );
not ( \420_b0 , w_469 );
and ( w_469 , w_468 , \420_b1 );
or ( \422_b1 , \418_b1 , \421_b1 );
xor ( \422_b0 , \418_b0 , w_470 );
not ( w_470 , w_471 );
and ( w_471 , \421_b1 , \421_b0 );
or ( \423_b1 , \317_A[8]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_472 );
and ( \423_b0 , \317_A[8]_b0 , w_473 );
and ( w_472 , w_473 , \173_B[2]_b0 );
or ( \424_b1 , \422_b1 , \423_b1 );
xor ( \424_b0 , \422_b0 , w_474 );
not ( w_474 , w_475 );
and ( w_475 , \423_b1 , \423_b0 );
or ( \425_b1 , \370_b1 , \371_b1 );
not ( \371_b1 , w_476 );
and ( \425_b0 , \370_b0 , w_477 );
and ( w_476 , w_477 , \371_b0 );
or ( \426_b1 , \372_b1 , \375_b1 );
not ( \375_b1 , w_478 );
and ( \426_b0 , \372_b0 , w_479 );
and ( w_478 , w_479 , \375_b0 );
or ( \427_b1 , \425_b1 , w_480 );
or ( \427_b0 , \425_b0 , \426_b0 );
not ( \426_b0 , w_481 );
and ( w_481 , w_480 , \426_b1 );
or ( \428_b1 , \424_b1 , \427_b1 );
xor ( \428_b0 , \424_b0 , w_482 );
not ( w_482 , w_483 );
and ( w_483 , \427_b1 , \427_b0 );
or ( \429_b1 , \277_A[7]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_484 );
and ( \429_b0 , \277_A[7]_b0 , w_485 );
and ( w_484 , w_485 , \189_B[3]_b0 );
or ( \430_b1 , \428_b1 , \429_b1 );
xor ( \430_b0 , \428_b0 , w_486 );
not ( w_486 , w_487 );
and ( w_487 , \429_b1 , \429_b0 );
or ( \431_b1 , \376_b1 , \377_b1 );
not ( \377_b1 , w_488 );
and ( \431_b0 , \376_b0 , w_489 );
and ( w_488 , w_489 , \377_b0 );
or ( \432_b1 , \378_b1 , \381_b1 );
not ( \381_b1 , w_490 );
and ( \432_b0 , \378_b0 , w_491 );
and ( w_490 , w_491 , \381_b0 );
or ( \433_b1 , \431_b1 , w_492 );
or ( \433_b0 , \431_b0 , \432_b0 );
not ( \432_b0 , w_493 );
and ( w_493 , w_492 , \432_b1 );
or ( \434_b1 , \430_b1 , \433_b1 );
xor ( \434_b0 , \430_b0 , w_494 );
not ( w_494 , w_495 );
and ( w_495 , \433_b1 , \433_b0 );
or ( \435_b1 , \243_A[6]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_496 );
and ( \435_b0 , \243_A[6]_b0 , w_497 );
and ( w_496 , w_497 , \211_B[4]_b0 );
or ( \436_b1 , \434_b1 , \435_b1 );
xor ( \436_b0 , \434_b0 , w_498 );
not ( w_498 , w_499 );
and ( w_499 , \435_b1 , \435_b0 );
or ( \437_b1 , \382_b1 , \383_b1 );
not ( \383_b1 , w_500 );
and ( \437_b0 , \382_b0 , w_501 );
and ( w_500 , w_501 , \383_b0 );
or ( \438_b1 , \384_b1 , \387_b1 );
not ( \387_b1 , w_502 );
and ( \438_b0 , \384_b0 , w_503 );
and ( w_502 , w_503 , \387_b0 );
or ( \439_b1 , \437_b1 , w_504 );
or ( \439_b0 , \437_b0 , \438_b0 );
not ( \438_b0 , w_505 );
and ( w_505 , w_504 , \438_b1 );
or ( \440_b1 , \436_b1 , \439_b1 );
xor ( \440_b0 , \436_b0 , w_506 );
not ( w_506 , w_507 );
and ( w_507 , \439_b1 , \439_b0 );
or ( \441_b1 , \215_A[5]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_508 );
and ( \441_b0 , \215_A[5]_b0 , w_509 );
and ( w_508 , w_509 , \239_B[5]_b0 );
or ( \442_b1 , \440_b1 , \441_b1 );
xor ( \442_b0 , \440_b0 , w_510 );
not ( w_510 , w_511 );
and ( w_511 , \441_b1 , \441_b0 );
or ( \443_b1 , \388_b1 , \389_b1 );
not ( \389_b1 , w_512 );
and ( \443_b0 , \388_b0 , w_513 );
and ( w_512 , w_513 , \389_b0 );
or ( \444_b1 , \390_b1 , \393_b1 );
not ( \393_b1 , w_514 );
and ( \444_b0 , \390_b0 , w_515 );
and ( w_514 , w_515 , \393_b0 );
or ( \445_b1 , \443_b1 , w_516 );
or ( \445_b0 , \443_b0 , \444_b0 );
not ( \444_b0 , w_517 );
and ( w_517 , w_516 , \444_b1 );
or ( \446_b1 , \442_b1 , \445_b1 );
xor ( \446_b0 , \442_b0 , w_518 );
not ( w_518 , w_519 );
and ( w_519 , \445_b1 , \445_b0 );
or ( \447_b1 , \193_A[4]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_520 );
and ( \447_b0 , \193_A[4]_b0 , w_521 );
and ( w_520 , w_521 , \273_B[6]_b0 );
or ( \448_b1 , \446_b1 , \447_b1 );
xor ( \448_b0 , \446_b0 , w_522 );
not ( w_522 , w_523 );
and ( w_523 , \447_b1 , \447_b0 );
or ( \449_b1 , \394_b1 , \395_b1 );
not ( \395_b1 , w_524 );
and ( \449_b0 , \394_b0 , w_525 );
and ( w_524 , w_525 , \395_b0 );
or ( \450_b1 , \396_b1 , \399_b1 );
not ( \399_b1 , w_526 );
and ( \450_b0 , \396_b0 , w_527 );
and ( w_526 , w_527 , \399_b0 );
or ( \451_b1 , \449_b1 , w_528 );
or ( \451_b0 , \449_b0 , \450_b0 );
not ( \450_b0 , w_529 );
and ( w_529 , w_528 , \450_b1 );
or ( \452_b1 , \448_b1 , \451_b1 );
xor ( \452_b0 , \448_b0 , w_530 );
not ( w_530 , w_531 );
and ( w_531 , \451_b1 , \451_b0 );
or ( \453_b1 , \177_A[3]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_532 );
and ( \453_b0 , \177_A[3]_b0 , w_533 );
and ( w_532 , w_533 , \313_B[7]_b0 );
or ( \454_b1 , \452_b1 , \453_b1 );
xor ( \454_b0 , \452_b0 , w_534 );
not ( w_534 , w_535 );
and ( w_535 , \453_b1 , \453_b0 );
or ( \455_b1 , \400_b1 , \401_b1 );
not ( \401_b1 , w_536 );
and ( \455_b0 , \400_b0 , w_537 );
and ( w_536 , w_537 , \401_b0 );
or ( \456_b1 , \402_b1 , \405_b1 );
not ( \405_b1 , w_538 );
and ( \456_b0 , \402_b0 , w_539 );
and ( w_538 , w_539 , \405_b0 );
or ( \457_b1 , \455_b1 , w_540 );
or ( \457_b0 , \455_b0 , \456_b0 );
not ( \456_b0 , w_541 );
and ( w_541 , w_540 , \456_b1 );
or ( \458_b1 , \454_b1 , \457_b1 );
xor ( \458_b0 , \454_b0 , w_542 );
not ( w_542 , w_543 );
and ( w_543 , \457_b1 , \457_b0 );
or ( \459_b1 , \167_A[2]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_544 );
and ( \459_b0 , \167_A[2]_b0 , w_545 );
and ( w_544 , w_545 , \359_B[8]_b0 );
or ( \460_b1 , \458_b1 , \459_b1 );
xor ( \460_b0 , \458_b0 , w_546 );
not ( w_546 , w_547 );
and ( w_547 , \459_b1 , \459_b0 );
or ( \461_b1 , \406_b1 , \407_b1 );
not ( \407_b1 , w_548 );
and ( \461_b0 , \406_b0 , w_549 );
and ( w_548 , w_549 , \407_b0 );
or ( \462_b1 , \408_b1 , \409_b1 );
not ( \409_b1 , w_550 );
and ( \462_b0 , \408_b0 , w_551 );
and ( w_550 , w_551 , \409_b0 );
or ( \463_b1 , \461_b1 , w_552 );
or ( \463_b0 , \461_b0 , \462_b0 );
not ( \462_b0 , w_553 );
and ( w_553 , w_552 , \462_b1 );
or ( \464_b1 , \460_b1 , \463_b1 );
xor ( \464_b0 , \460_b0 , w_554 );
not ( w_554 , w_555 );
and ( w_555 , \463_b1 , \463_b0 );
or ( \465_b1 , \161_A[1]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_556 );
and ( \465_b0 , \161_A[1]_b0 , w_557 );
and ( w_556 , w_557 , \411_B[9]_b0 );
or ( \466_b1 , \464_b1 , \465_b1 );
xor ( \466_b0 , \464_b0 , w_558 );
not ( w_558 , w_559 );
and ( w_559 , \465_b1 , \465_b0 );
or ( \467_b1 , \410_b1 , \412_b1 );
not ( \412_b1 , w_560 );
and ( \467_b0 , \410_b0 , w_561 );
and ( w_560 , w_561 , \412_b0 );
or ( \468_b1 , \466_b1 , \467_b1 );
xor ( \468_b0 , \466_b0 , w_562 );
not ( w_562 , w_563 );
and ( w_563 , \467_b1 , \467_b0 );
buf ( \469_B[10]_b1 , \b[10]_b1 );
buf ( \469_B[10]_b0 , \b[10]_b0 );
or ( \470_b1 , \156_A[0]_b1 , \469_B[10]_b1 );
not ( \469_B[10]_b1 , w_564 );
and ( \470_b0 , \156_A[0]_b0 , w_565 );
and ( w_564 , w_565 , \469_B[10]_b0 );
or ( \471_b1 , \468_b1 , \470_b1 );
xor ( \471_b0 , \468_b0 , w_566 );
not ( w_566 , w_567 );
and ( w_567 , \470_b1 , \470_b0 );
buf ( \472_Z[10]_b1 , \471_b1 );
buf ( \472_Z[10]_b0 , \471_b0 );
buf ( \473_A[11]_b1 , \a[11]_b1 );
buf ( \473_A[11]_b0 , \a[11]_b0 );
or ( \474_b1 , \473_A[11]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_568 );
and ( \474_b0 , \473_A[11]_b0 , w_569 );
and ( w_568 , w_569 , \157_B[0]_b0 );
or ( \475_b1 , \415_A[10]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_570 );
and ( \475_b0 , \415_A[10]_b0 , w_571 );
and ( w_570 , w_571 , \163_B[1]_b0 );
or ( \476_b1 , \474_b1 , \475_b1 );
xor ( \476_b0 , \474_b0 , w_572 );
not ( w_572 , w_573 );
and ( w_573 , \475_b1 , \475_b0 );
or ( \477_b1 , \416_b1 , \417_b1 );
not ( \417_b1 , w_574 );
and ( \477_b0 , \416_b0 , w_575 );
and ( w_574 , w_575 , \417_b0 );
or ( \478_b1 , \418_b1 , \421_b1 );
not ( \421_b1 , w_576 );
and ( \478_b0 , \418_b0 , w_577 );
and ( w_576 , w_577 , \421_b0 );
or ( \479_b1 , \477_b1 , w_578 );
or ( \479_b0 , \477_b0 , \478_b0 );
not ( \478_b0 , w_579 );
and ( w_579 , w_578 , \478_b1 );
or ( \480_b1 , \476_b1 , \479_b1 );
xor ( \480_b0 , \476_b0 , w_580 );
not ( w_580 , w_581 );
and ( w_581 , \479_b1 , \479_b0 );
or ( \481_b1 , \363_A[9]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_582 );
and ( \481_b0 , \363_A[9]_b0 , w_583 );
and ( w_582 , w_583 , \173_B[2]_b0 );
or ( \482_b1 , \480_b1 , \481_b1 );
xor ( \482_b0 , \480_b0 , w_584 );
not ( w_584 , w_585 );
and ( w_585 , \481_b1 , \481_b0 );
or ( \483_b1 , \422_b1 , \423_b1 );
not ( \423_b1 , w_586 );
and ( \483_b0 , \422_b0 , w_587 );
and ( w_586 , w_587 , \423_b0 );
or ( \484_b1 , \424_b1 , \427_b1 );
not ( \427_b1 , w_588 );
and ( \484_b0 , \424_b0 , w_589 );
and ( w_588 , w_589 , \427_b0 );
or ( \485_b1 , \483_b1 , w_590 );
or ( \485_b0 , \483_b0 , \484_b0 );
not ( \484_b0 , w_591 );
and ( w_591 , w_590 , \484_b1 );
or ( \486_b1 , \482_b1 , \485_b1 );
xor ( \486_b0 , \482_b0 , w_592 );
not ( w_592 , w_593 );
and ( w_593 , \485_b1 , \485_b0 );
or ( \487_b1 , \317_A[8]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_594 );
and ( \487_b0 , \317_A[8]_b0 , w_595 );
and ( w_594 , w_595 , \189_B[3]_b0 );
or ( \488_b1 , \486_b1 , \487_b1 );
xor ( \488_b0 , \486_b0 , w_596 );
not ( w_596 , w_597 );
and ( w_597 , \487_b1 , \487_b0 );
or ( \489_b1 , \428_b1 , \429_b1 );
not ( \429_b1 , w_598 );
and ( \489_b0 , \428_b0 , w_599 );
and ( w_598 , w_599 , \429_b0 );
or ( \490_b1 , \430_b1 , \433_b1 );
not ( \433_b1 , w_600 );
and ( \490_b0 , \430_b0 , w_601 );
and ( w_600 , w_601 , \433_b0 );
or ( \491_b1 , \489_b1 , w_602 );
or ( \491_b0 , \489_b0 , \490_b0 );
not ( \490_b0 , w_603 );
and ( w_603 , w_602 , \490_b1 );
or ( \492_b1 , \488_b1 , \491_b1 );
xor ( \492_b0 , \488_b0 , w_604 );
not ( w_604 , w_605 );
and ( w_605 , \491_b1 , \491_b0 );
or ( \493_b1 , \277_A[7]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_606 );
and ( \493_b0 , \277_A[7]_b0 , w_607 );
and ( w_606 , w_607 , \211_B[4]_b0 );
or ( \494_b1 , \492_b1 , \493_b1 );
xor ( \494_b0 , \492_b0 , w_608 );
not ( w_608 , w_609 );
and ( w_609 , \493_b1 , \493_b0 );
or ( \495_b1 , \434_b1 , \435_b1 );
not ( \435_b1 , w_610 );
and ( \495_b0 , \434_b0 , w_611 );
and ( w_610 , w_611 , \435_b0 );
or ( \496_b1 , \436_b1 , \439_b1 );
not ( \439_b1 , w_612 );
and ( \496_b0 , \436_b0 , w_613 );
and ( w_612 , w_613 , \439_b0 );
or ( \497_b1 , \495_b1 , w_614 );
or ( \497_b0 , \495_b0 , \496_b0 );
not ( \496_b0 , w_615 );
and ( w_615 , w_614 , \496_b1 );
or ( \498_b1 , \494_b1 , \497_b1 );
xor ( \498_b0 , \494_b0 , w_616 );
not ( w_616 , w_617 );
and ( w_617 , \497_b1 , \497_b0 );
or ( \499_b1 , \243_A[6]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_618 );
and ( \499_b0 , \243_A[6]_b0 , w_619 );
and ( w_618 , w_619 , \239_B[5]_b0 );
or ( \500_b1 , \498_b1 , \499_b1 );
xor ( \500_b0 , \498_b0 , w_620 );
not ( w_620 , w_621 );
and ( w_621 , \499_b1 , \499_b0 );
or ( \501_b1 , \440_b1 , \441_b1 );
not ( \441_b1 , w_622 );
and ( \501_b0 , \440_b0 , w_623 );
and ( w_622 , w_623 , \441_b0 );
or ( \502_b1 , \442_b1 , \445_b1 );
not ( \445_b1 , w_624 );
and ( \502_b0 , \442_b0 , w_625 );
and ( w_624 , w_625 , \445_b0 );
or ( \503_b1 , \501_b1 , w_626 );
or ( \503_b0 , \501_b0 , \502_b0 );
not ( \502_b0 , w_627 );
and ( w_627 , w_626 , \502_b1 );
or ( \504_b1 , \500_b1 , \503_b1 );
xor ( \504_b0 , \500_b0 , w_628 );
not ( w_628 , w_629 );
and ( w_629 , \503_b1 , \503_b0 );
or ( \505_b1 , \215_A[5]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_630 );
and ( \505_b0 , \215_A[5]_b0 , w_631 );
and ( w_630 , w_631 , \273_B[6]_b0 );
or ( \506_b1 , \504_b1 , \505_b1 );
xor ( \506_b0 , \504_b0 , w_632 );
not ( w_632 , w_633 );
and ( w_633 , \505_b1 , \505_b0 );
or ( \507_b1 , \446_b1 , \447_b1 );
not ( \447_b1 , w_634 );
and ( \507_b0 , \446_b0 , w_635 );
and ( w_634 , w_635 , \447_b0 );
or ( \508_b1 , \448_b1 , \451_b1 );
not ( \451_b1 , w_636 );
and ( \508_b0 , \448_b0 , w_637 );
and ( w_636 , w_637 , \451_b0 );
or ( \509_b1 , \507_b1 , w_638 );
or ( \509_b0 , \507_b0 , \508_b0 );
not ( \508_b0 , w_639 );
and ( w_639 , w_638 , \508_b1 );
or ( \510_b1 , \506_b1 , \509_b1 );
xor ( \510_b0 , \506_b0 , w_640 );
not ( w_640 , w_641 );
and ( w_641 , \509_b1 , \509_b0 );
or ( \511_b1 , \193_A[4]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_642 );
and ( \511_b0 , \193_A[4]_b0 , w_643 );
and ( w_642 , w_643 , \313_B[7]_b0 );
or ( \512_b1 , \510_b1 , \511_b1 );
xor ( \512_b0 , \510_b0 , w_644 );
not ( w_644 , w_645 );
and ( w_645 , \511_b1 , \511_b0 );
or ( \513_b1 , \452_b1 , \453_b1 );
not ( \453_b1 , w_646 );
and ( \513_b0 , \452_b0 , w_647 );
and ( w_646 , w_647 , \453_b0 );
or ( \514_b1 , \454_b1 , \457_b1 );
not ( \457_b1 , w_648 );
and ( \514_b0 , \454_b0 , w_649 );
and ( w_648 , w_649 , \457_b0 );
or ( \515_b1 , \513_b1 , w_650 );
or ( \515_b0 , \513_b0 , \514_b0 );
not ( \514_b0 , w_651 );
and ( w_651 , w_650 , \514_b1 );
or ( \516_b1 , \512_b1 , \515_b1 );
xor ( \516_b0 , \512_b0 , w_652 );
not ( w_652 , w_653 );
and ( w_653 , \515_b1 , \515_b0 );
or ( \517_b1 , \177_A[3]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_654 );
and ( \517_b0 , \177_A[3]_b0 , w_655 );
and ( w_654 , w_655 , \359_B[8]_b0 );
or ( \518_b1 , \516_b1 , \517_b1 );
xor ( \518_b0 , \516_b0 , w_656 );
not ( w_656 , w_657 );
and ( w_657 , \517_b1 , \517_b0 );
or ( \519_b1 , \458_b1 , \459_b1 );
not ( \459_b1 , w_658 );
and ( \519_b0 , \458_b0 , w_659 );
and ( w_658 , w_659 , \459_b0 );
or ( \520_b1 , \460_b1 , \463_b1 );
not ( \463_b1 , w_660 );
and ( \520_b0 , \460_b0 , w_661 );
and ( w_660 , w_661 , \463_b0 );
or ( \521_b1 , \519_b1 , w_662 );
or ( \521_b0 , \519_b0 , \520_b0 );
not ( \520_b0 , w_663 );
and ( w_663 , w_662 , \520_b1 );
or ( \522_b1 , \518_b1 , \521_b1 );
xor ( \522_b0 , \518_b0 , w_664 );
not ( w_664 , w_665 );
and ( w_665 , \521_b1 , \521_b0 );
or ( \523_b1 , \167_A[2]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_666 );
and ( \523_b0 , \167_A[2]_b0 , w_667 );
and ( w_666 , w_667 , \411_B[9]_b0 );
or ( \524_b1 , \522_b1 , \523_b1 );
xor ( \524_b0 , \522_b0 , w_668 );
not ( w_668 , w_669 );
and ( w_669 , \523_b1 , \523_b0 );
or ( \525_b1 , \464_b1 , \465_b1 );
not ( \465_b1 , w_670 );
and ( \525_b0 , \464_b0 , w_671 );
and ( w_670 , w_671 , \465_b0 );
or ( \526_b1 , \466_b1 , \467_b1 );
not ( \467_b1 , w_672 );
and ( \526_b0 , \466_b0 , w_673 );
and ( w_672 , w_673 , \467_b0 );
or ( \527_b1 , \525_b1 , w_674 );
or ( \527_b0 , \525_b0 , \526_b0 );
not ( \526_b0 , w_675 );
and ( w_675 , w_674 , \526_b1 );
or ( \528_b1 , \524_b1 , \527_b1 );
xor ( \528_b0 , \524_b0 , w_676 );
not ( w_676 , w_677 );
and ( w_677 , \527_b1 , \527_b0 );
or ( \529_b1 , \161_A[1]_b1 , \469_B[10]_b1 );
not ( \469_B[10]_b1 , w_678 );
and ( \529_b0 , \161_A[1]_b0 , w_679 );
and ( w_678 , w_679 , \469_B[10]_b0 );
or ( \530_b1 , \528_b1 , \529_b1 );
xor ( \530_b0 , \528_b0 , w_680 );
not ( w_680 , w_681 );
and ( w_681 , \529_b1 , \529_b0 );
or ( \531_b1 , \468_b1 , \470_b1 );
not ( \470_b1 , w_682 );
and ( \531_b0 , \468_b0 , w_683 );
and ( w_682 , w_683 , \470_b0 );
or ( \532_b1 , \530_b1 , \531_b1 );
xor ( \532_b0 , \530_b0 , w_684 );
not ( w_684 , w_685 );
and ( w_685 , \531_b1 , \531_b0 );
buf ( \533_B[11]_b1 , \b[11]_b1 );
buf ( \533_B[11]_b0 , \b[11]_b0 );
or ( \534_b1 , \156_A[0]_b1 , \533_B[11]_b1 );
not ( \533_B[11]_b1 , w_686 );
and ( \534_b0 , \156_A[0]_b0 , w_687 );
and ( w_686 , w_687 , \533_B[11]_b0 );
or ( \535_b1 , \532_b1 , \534_b1 );
xor ( \535_b0 , \532_b0 , w_688 );
not ( w_688 , w_689 );
and ( w_689 , \534_b1 , \534_b0 );
buf ( \536_Z[11]_b1 , \535_b1 );
buf ( \536_Z[11]_b0 , \535_b0 );
buf ( \537_A[12]_b1 , \a[12]_b1 );
buf ( \537_A[12]_b0 , \a[12]_b0 );
or ( \538_b1 , \537_A[12]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_690 );
and ( \538_b0 , \537_A[12]_b0 , w_691 );
and ( w_690 , w_691 , \157_B[0]_b0 );
or ( \539_b1 , \473_A[11]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_692 );
and ( \539_b0 , \473_A[11]_b0 , w_693 );
and ( w_692 , w_693 , \163_B[1]_b0 );
or ( \540_b1 , \538_b1 , \539_b1 );
xor ( \540_b0 , \538_b0 , w_694 );
not ( w_694 , w_695 );
and ( w_695 , \539_b1 , \539_b0 );
or ( \541_b1 , \474_b1 , \475_b1 );
not ( \475_b1 , w_696 );
and ( \541_b0 , \474_b0 , w_697 );
and ( w_696 , w_697 , \475_b0 );
or ( \542_b1 , \476_b1 , \479_b1 );
not ( \479_b1 , w_698 );
and ( \542_b0 , \476_b0 , w_699 );
and ( w_698 , w_699 , \479_b0 );
or ( \543_b1 , \541_b1 , w_700 );
or ( \543_b0 , \541_b0 , \542_b0 );
not ( \542_b0 , w_701 );
and ( w_701 , w_700 , \542_b1 );
or ( \544_b1 , \540_b1 , \543_b1 );
xor ( \544_b0 , \540_b0 , w_702 );
not ( w_702 , w_703 );
and ( w_703 , \543_b1 , \543_b0 );
or ( \545_b1 , \415_A[10]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_704 );
and ( \545_b0 , \415_A[10]_b0 , w_705 );
and ( w_704 , w_705 , \173_B[2]_b0 );
or ( \546_b1 , \544_b1 , \545_b1 );
xor ( \546_b0 , \544_b0 , w_706 );
not ( w_706 , w_707 );
and ( w_707 , \545_b1 , \545_b0 );
or ( \547_b1 , \480_b1 , \481_b1 );
not ( \481_b1 , w_708 );
and ( \547_b0 , \480_b0 , w_709 );
and ( w_708 , w_709 , \481_b0 );
or ( \548_b1 , \482_b1 , \485_b1 );
not ( \485_b1 , w_710 );
and ( \548_b0 , \482_b0 , w_711 );
and ( w_710 , w_711 , \485_b0 );
or ( \549_b1 , \547_b1 , w_712 );
or ( \549_b0 , \547_b0 , \548_b0 );
not ( \548_b0 , w_713 );
and ( w_713 , w_712 , \548_b1 );
or ( \550_b1 , \546_b1 , \549_b1 );
xor ( \550_b0 , \546_b0 , w_714 );
not ( w_714 , w_715 );
and ( w_715 , \549_b1 , \549_b0 );
or ( \551_b1 , \363_A[9]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_716 );
and ( \551_b0 , \363_A[9]_b0 , w_717 );
and ( w_716 , w_717 , \189_B[3]_b0 );
or ( \552_b1 , \550_b1 , \551_b1 );
xor ( \552_b0 , \550_b0 , w_718 );
not ( w_718 , w_719 );
and ( w_719 , \551_b1 , \551_b0 );
or ( \553_b1 , \486_b1 , \487_b1 );
not ( \487_b1 , w_720 );
and ( \553_b0 , \486_b0 , w_721 );
and ( w_720 , w_721 , \487_b0 );
or ( \554_b1 , \488_b1 , \491_b1 );
not ( \491_b1 , w_722 );
and ( \554_b0 , \488_b0 , w_723 );
and ( w_722 , w_723 , \491_b0 );
or ( \555_b1 , \553_b1 , w_724 );
or ( \555_b0 , \553_b0 , \554_b0 );
not ( \554_b0 , w_725 );
and ( w_725 , w_724 , \554_b1 );
or ( \556_b1 , \552_b1 , \555_b1 );
xor ( \556_b0 , \552_b0 , w_726 );
not ( w_726 , w_727 );
and ( w_727 , \555_b1 , \555_b0 );
or ( \557_b1 , \317_A[8]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_728 );
and ( \557_b0 , \317_A[8]_b0 , w_729 );
and ( w_728 , w_729 , \211_B[4]_b0 );
or ( \558_b1 , \556_b1 , \557_b1 );
xor ( \558_b0 , \556_b0 , w_730 );
not ( w_730 , w_731 );
and ( w_731 , \557_b1 , \557_b0 );
or ( \559_b1 , \492_b1 , \493_b1 );
not ( \493_b1 , w_732 );
and ( \559_b0 , \492_b0 , w_733 );
and ( w_732 , w_733 , \493_b0 );
or ( \560_b1 , \494_b1 , \497_b1 );
not ( \497_b1 , w_734 );
and ( \560_b0 , \494_b0 , w_735 );
and ( w_734 , w_735 , \497_b0 );
or ( \561_b1 , \559_b1 , w_736 );
or ( \561_b0 , \559_b0 , \560_b0 );
not ( \560_b0 , w_737 );
and ( w_737 , w_736 , \560_b1 );
or ( \562_b1 , \558_b1 , \561_b1 );
xor ( \562_b0 , \558_b0 , w_738 );
not ( w_738 , w_739 );
and ( w_739 , \561_b1 , \561_b0 );
or ( \563_b1 , \277_A[7]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_740 );
and ( \563_b0 , \277_A[7]_b0 , w_741 );
and ( w_740 , w_741 , \239_B[5]_b0 );
or ( \564_b1 , \562_b1 , \563_b1 );
xor ( \564_b0 , \562_b0 , w_742 );
not ( w_742 , w_743 );
and ( w_743 , \563_b1 , \563_b0 );
or ( \565_b1 , \498_b1 , \499_b1 );
not ( \499_b1 , w_744 );
and ( \565_b0 , \498_b0 , w_745 );
and ( w_744 , w_745 , \499_b0 );
or ( \566_b1 , \500_b1 , \503_b1 );
not ( \503_b1 , w_746 );
and ( \566_b0 , \500_b0 , w_747 );
and ( w_746 , w_747 , \503_b0 );
or ( \567_b1 , \565_b1 , w_748 );
or ( \567_b0 , \565_b0 , \566_b0 );
not ( \566_b0 , w_749 );
and ( w_749 , w_748 , \566_b1 );
or ( \568_b1 , \564_b1 , \567_b1 );
xor ( \568_b0 , \564_b0 , w_750 );
not ( w_750 , w_751 );
and ( w_751 , \567_b1 , \567_b0 );
or ( \569_b1 , \243_A[6]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_752 );
and ( \569_b0 , \243_A[6]_b0 , w_753 );
and ( w_752 , w_753 , \273_B[6]_b0 );
or ( \570_b1 , \568_b1 , \569_b1 );
xor ( \570_b0 , \568_b0 , w_754 );
not ( w_754 , w_755 );
and ( w_755 , \569_b1 , \569_b0 );
or ( \571_b1 , \504_b1 , \505_b1 );
not ( \505_b1 , w_756 );
and ( \571_b0 , \504_b0 , w_757 );
and ( w_756 , w_757 , \505_b0 );
or ( \572_b1 , \506_b1 , \509_b1 );
not ( \509_b1 , w_758 );
and ( \572_b0 , \506_b0 , w_759 );
and ( w_758 , w_759 , \509_b0 );
or ( \573_b1 , \571_b1 , w_760 );
or ( \573_b0 , \571_b0 , \572_b0 );
not ( \572_b0 , w_761 );
and ( w_761 , w_760 , \572_b1 );
or ( \574_b1 , \570_b1 , \573_b1 );
xor ( \574_b0 , \570_b0 , w_762 );
not ( w_762 , w_763 );
and ( w_763 , \573_b1 , \573_b0 );
or ( \575_b1 , \215_A[5]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_764 );
and ( \575_b0 , \215_A[5]_b0 , w_765 );
and ( w_764 , w_765 , \313_B[7]_b0 );
or ( \576_b1 , \574_b1 , \575_b1 );
xor ( \576_b0 , \574_b0 , w_766 );
not ( w_766 , w_767 );
and ( w_767 , \575_b1 , \575_b0 );
or ( \577_b1 , \510_b1 , \511_b1 );
not ( \511_b1 , w_768 );
and ( \577_b0 , \510_b0 , w_769 );
and ( w_768 , w_769 , \511_b0 );
or ( \578_b1 , \512_b1 , \515_b1 );
not ( \515_b1 , w_770 );
and ( \578_b0 , \512_b0 , w_771 );
and ( w_770 , w_771 , \515_b0 );
or ( \579_b1 , \577_b1 , w_772 );
or ( \579_b0 , \577_b0 , \578_b0 );
not ( \578_b0 , w_773 );
and ( w_773 , w_772 , \578_b1 );
or ( \580_b1 , \576_b1 , \579_b1 );
xor ( \580_b0 , \576_b0 , w_774 );
not ( w_774 , w_775 );
and ( w_775 , \579_b1 , \579_b0 );
or ( \581_b1 , \193_A[4]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_776 );
and ( \581_b0 , \193_A[4]_b0 , w_777 );
and ( w_776 , w_777 , \359_B[8]_b0 );
or ( \582_b1 , \580_b1 , \581_b1 );
xor ( \582_b0 , \580_b0 , w_778 );
not ( w_778 , w_779 );
and ( w_779 , \581_b1 , \581_b0 );
or ( \583_b1 , \516_b1 , \517_b1 );
not ( \517_b1 , w_780 );
and ( \583_b0 , \516_b0 , w_781 );
and ( w_780 , w_781 , \517_b0 );
or ( \584_b1 , \518_b1 , \521_b1 );
not ( \521_b1 , w_782 );
and ( \584_b0 , \518_b0 , w_783 );
and ( w_782 , w_783 , \521_b0 );
or ( \585_b1 , \583_b1 , w_784 );
or ( \585_b0 , \583_b0 , \584_b0 );
not ( \584_b0 , w_785 );
and ( w_785 , w_784 , \584_b1 );
or ( \586_b1 , \582_b1 , \585_b1 );
xor ( \586_b0 , \582_b0 , w_786 );
not ( w_786 , w_787 );
and ( w_787 , \585_b1 , \585_b0 );
or ( \587_b1 , \177_A[3]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_788 );
and ( \587_b0 , \177_A[3]_b0 , w_789 );
and ( w_788 , w_789 , \411_B[9]_b0 );
or ( \588_b1 , \586_b1 , \587_b1 );
xor ( \588_b0 , \586_b0 , w_790 );
not ( w_790 , w_791 );
and ( w_791 , \587_b1 , \587_b0 );
or ( \589_b1 , \522_b1 , \523_b1 );
not ( \523_b1 , w_792 );
and ( \589_b0 , \522_b0 , w_793 );
and ( w_792 , w_793 , \523_b0 );
or ( \590_b1 , \524_b1 , \527_b1 );
not ( \527_b1 , w_794 );
and ( \590_b0 , \524_b0 , w_795 );
and ( w_794 , w_795 , \527_b0 );
or ( \591_b1 , \589_b1 , w_796 );
or ( \591_b0 , \589_b0 , \590_b0 );
not ( \590_b0 , w_797 );
and ( w_797 , w_796 , \590_b1 );
or ( \592_b1 , \588_b1 , \591_b1 );
xor ( \592_b0 , \588_b0 , w_798 );
not ( w_798 , w_799 );
and ( w_799 , \591_b1 , \591_b0 );
or ( \593_b1 , \167_A[2]_b1 , \469_B[10]_b1 );
not ( \469_B[10]_b1 , w_800 );
and ( \593_b0 , \167_A[2]_b0 , w_801 );
and ( w_800 , w_801 , \469_B[10]_b0 );
or ( \594_b1 , \592_b1 , \593_b1 );
xor ( \594_b0 , \592_b0 , w_802 );
not ( w_802 , w_803 );
and ( w_803 , \593_b1 , \593_b0 );
or ( \595_b1 , \528_b1 , \529_b1 );
not ( \529_b1 , w_804 );
and ( \595_b0 , \528_b0 , w_805 );
and ( w_804 , w_805 , \529_b0 );
or ( \596_b1 , \530_b1 , \531_b1 );
not ( \531_b1 , w_806 );
and ( \596_b0 , \530_b0 , w_807 );
and ( w_806 , w_807 , \531_b0 );
or ( \597_b1 , \595_b1 , w_808 );
or ( \597_b0 , \595_b0 , \596_b0 );
not ( \596_b0 , w_809 );
and ( w_809 , w_808 , \596_b1 );
or ( \598_b1 , \594_b1 , \597_b1 );
xor ( \598_b0 , \594_b0 , w_810 );
not ( w_810 , w_811 );
and ( w_811 , \597_b1 , \597_b0 );
or ( \599_b1 , \161_A[1]_b1 , \533_B[11]_b1 );
not ( \533_B[11]_b1 , w_812 );
and ( \599_b0 , \161_A[1]_b0 , w_813 );
and ( w_812 , w_813 , \533_B[11]_b0 );
or ( \600_b1 , \598_b1 , \599_b1 );
xor ( \600_b0 , \598_b0 , w_814 );
not ( w_814 , w_815 );
and ( w_815 , \599_b1 , \599_b0 );
or ( \601_b1 , \532_b1 , \534_b1 );
not ( \534_b1 , w_816 );
and ( \601_b0 , \532_b0 , w_817 );
and ( w_816 , w_817 , \534_b0 );
or ( \602_b1 , \600_b1 , \601_b1 );
xor ( \602_b0 , \600_b0 , w_818 );
not ( w_818 , w_819 );
and ( w_819 , \601_b1 , \601_b0 );
buf ( \603_B[12]_b1 , \b[12]_b1 );
buf ( \603_B[12]_b0 , \b[12]_b0 );
or ( \604_b1 , \156_A[0]_b1 , \603_B[12]_b1 );
not ( \603_B[12]_b1 , w_820 );
and ( \604_b0 , \156_A[0]_b0 , w_821 );
and ( w_820 , w_821 , \603_B[12]_b0 );
or ( \605_b1 , \602_b1 , \604_b1 );
xor ( \605_b0 , \602_b0 , w_822 );
not ( w_822 , w_823 );
and ( w_823 , \604_b1 , \604_b0 );
buf ( \606_Z[12]_b1 , \605_b1 );
buf ( \606_Z[12]_b0 , \605_b0 );
buf ( \607_A[13]_b1 , \a[13]_b1 );
buf ( \607_A[13]_b0 , \a[13]_b0 );
or ( \608_b1 , \607_A[13]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_824 );
and ( \608_b0 , \607_A[13]_b0 , w_825 );
and ( w_824 , w_825 , \157_B[0]_b0 );
or ( \609_b1 , \537_A[12]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_826 );
and ( \609_b0 , \537_A[12]_b0 , w_827 );
and ( w_826 , w_827 , \163_B[1]_b0 );
or ( \610_b1 , \608_b1 , \609_b1 );
xor ( \610_b0 , \608_b0 , w_828 );
not ( w_828 , w_829 );
and ( w_829 , \609_b1 , \609_b0 );
or ( \611_b1 , \538_b1 , \539_b1 );
not ( \539_b1 , w_830 );
and ( \611_b0 , \538_b0 , w_831 );
and ( w_830 , w_831 , \539_b0 );
or ( \612_b1 , \540_b1 , \543_b1 );
not ( \543_b1 , w_832 );
and ( \612_b0 , \540_b0 , w_833 );
and ( w_832 , w_833 , \543_b0 );
or ( \613_b1 , \611_b1 , w_834 );
or ( \613_b0 , \611_b0 , \612_b0 );
not ( \612_b0 , w_835 );
and ( w_835 , w_834 , \612_b1 );
or ( \614_b1 , \610_b1 , \613_b1 );
xor ( \614_b0 , \610_b0 , w_836 );
not ( w_836 , w_837 );
and ( w_837 , \613_b1 , \613_b0 );
or ( \615_b1 , \473_A[11]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_838 );
and ( \615_b0 , \473_A[11]_b0 , w_839 );
and ( w_838 , w_839 , \173_B[2]_b0 );
or ( \616_b1 , \614_b1 , \615_b1 );
xor ( \616_b0 , \614_b0 , w_840 );
not ( w_840 , w_841 );
and ( w_841 , \615_b1 , \615_b0 );
or ( \617_b1 , \544_b1 , \545_b1 );
not ( \545_b1 , w_842 );
and ( \617_b0 , \544_b0 , w_843 );
and ( w_842 , w_843 , \545_b0 );
or ( \618_b1 , \546_b1 , \549_b1 );
not ( \549_b1 , w_844 );
and ( \618_b0 , \546_b0 , w_845 );
and ( w_844 , w_845 , \549_b0 );
or ( \619_b1 , \617_b1 , w_846 );
or ( \619_b0 , \617_b0 , \618_b0 );
not ( \618_b0 , w_847 );
and ( w_847 , w_846 , \618_b1 );
or ( \620_b1 , \616_b1 , \619_b1 );
xor ( \620_b0 , \616_b0 , w_848 );
not ( w_848 , w_849 );
and ( w_849 , \619_b1 , \619_b0 );
or ( \621_b1 , \415_A[10]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_850 );
and ( \621_b0 , \415_A[10]_b0 , w_851 );
and ( w_850 , w_851 , \189_B[3]_b0 );
or ( \622_b1 , \620_b1 , \621_b1 );
xor ( \622_b0 , \620_b0 , w_852 );
not ( w_852 , w_853 );
and ( w_853 , \621_b1 , \621_b0 );
or ( \623_b1 , \550_b1 , \551_b1 );
not ( \551_b1 , w_854 );
and ( \623_b0 , \550_b0 , w_855 );
and ( w_854 , w_855 , \551_b0 );
or ( \624_b1 , \552_b1 , \555_b1 );
not ( \555_b1 , w_856 );
and ( \624_b0 , \552_b0 , w_857 );
and ( w_856 , w_857 , \555_b0 );
or ( \625_b1 , \623_b1 , w_858 );
or ( \625_b0 , \623_b0 , \624_b0 );
not ( \624_b0 , w_859 );
and ( w_859 , w_858 , \624_b1 );
or ( \626_b1 , \622_b1 , \625_b1 );
xor ( \626_b0 , \622_b0 , w_860 );
not ( w_860 , w_861 );
and ( w_861 , \625_b1 , \625_b0 );
or ( \627_b1 , \363_A[9]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_862 );
and ( \627_b0 , \363_A[9]_b0 , w_863 );
and ( w_862 , w_863 , \211_B[4]_b0 );
or ( \628_b1 , \626_b1 , \627_b1 );
xor ( \628_b0 , \626_b0 , w_864 );
not ( w_864 , w_865 );
and ( w_865 , \627_b1 , \627_b0 );
or ( \629_b1 , \556_b1 , \557_b1 );
not ( \557_b1 , w_866 );
and ( \629_b0 , \556_b0 , w_867 );
and ( w_866 , w_867 , \557_b0 );
or ( \630_b1 , \558_b1 , \561_b1 );
not ( \561_b1 , w_868 );
and ( \630_b0 , \558_b0 , w_869 );
and ( w_868 , w_869 , \561_b0 );
or ( \631_b1 , \629_b1 , w_870 );
or ( \631_b0 , \629_b0 , \630_b0 );
not ( \630_b0 , w_871 );
and ( w_871 , w_870 , \630_b1 );
or ( \632_b1 , \628_b1 , \631_b1 );
xor ( \632_b0 , \628_b0 , w_872 );
not ( w_872 , w_873 );
and ( w_873 , \631_b1 , \631_b0 );
or ( \633_b1 , \317_A[8]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_874 );
and ( \633_b0 , \317_A[8]_b0 , w_875 );
and ( w_874 , w_875 , \239_B[5]_b0 );
or ( \634_b1 , \632_b1 , \633_b1 );
xor ( \634_b0 , \632_b0 , w_876 );
not ( w_876 , w_877 );
and ( w_877 , \633_b1 , \633_b0 );
or ( \635_b1 , \562_b1 , \563_b1 );
not ( \563_b1 , w_878 );
and ( \635_b0 , \562_b0 , w_879 );
and ( w_878 , w_879 , \563_b0 );
or ( \636_b1 , \564_b1 , \567_b1 );
not ( \567_b1 , w_880 );
and ( \636_b0 , \564_b0 , w_881 );
and ( w_880 , w_881 , \567_b0 );
or ( \637_b1 , \635_b1 , w_882 );
or ( \637_b0 , \635_b0 , \636_b0 );
not ( \636_b0 , w_883 );
and ( w_883 , w_882 , \636_b1 );
or ( \638_b1 , \634_b1 , \637_b1 );
xor ( \638_b0 , \634_b0 , w_884 );
not ( w_884 , w_885 );
and ( w_885 , \637_b1 , \637_b0 );
or ( \639_b1 , \277_A[7]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_886 );
and ( \639_b0 , \277_A[7]_b0 , w_887 );
and ( w_886 , w_887 , \273_B[6]_b0 );
or ( \640_b1 , \638_b1 , \639_b1 );
xor ( \640_b0 , \638_b0 , w_888 );
not ( w_888 , w_889 );
and ( w_889 , \639_b1 , \639_b0 );
or ( \641_b1 , \568_b1 , \569_b1 );
not ( \569_b1 , w_890 );
and ( \641_b0 , \568_b0 , w_891 );
and ( w_890 , w_891 , \569_b0 );
or ( \642_b1 , \570_b1 , \573_b1 );
not ( \573_b1 , w_892 );
and ( \642_b0 , \570_b0 , w_893 );
and ( w_892 , w_893 , \573_b0 );
or ( \643_b1 , \641_b1 , w_894 );
or ( \643_b0 , \641_b0 , \642_b0 );
not ( \642_b0 , w_895 );
and ( w_895 , w_894 , \642_b1 );
or ( \644_b1 , \640_b1 , \643_b1 );
xor ( \644_b0 , \640_b0 , w_896 );
not ( w_896 , w_897 );
and ( w_897 , \643_b1 , \643_b0 );
or ( \645_b1 , \243_A[6]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_898 );
and ( \645_b0 , \243_A[6]_b0 , w_899 );
and ( w_898 , w_899 , \313_B[7]_b0 );
or ( \646_b1 , \644_b1 , \645_b1 );
xor ( \646_b0 , \644_b0 , w_900 );
not ( w_900 , w_901 );
and ( w_901 , \645_b1 , \645_b0 );
or ( \647_b1 , \574_b1 , \575_b1 );
not ( \575_b1 , w_902 );
and ( \647_b0 , \574_b0 , w_903 );
and ( w_902 , w_903 , \575_b0 );
or ( \648_b1 , \576_b1 , \579_b1 );
not ( \579_b1 , w_904 );
and ( \648_b0 , \576_b0 , w_905 );
and ( w_904 , w_905 , \579_b0 );
or ( \649_b1 , \647_b1 , w_906 );
or ( \649_b0 , \647_b0 , \648_b0 );
not ( \648_b0 , w_907 );
and ( w_907 , w_906 , \648_b1 );
or ( \650_b1 , \646_b1 , \649_b1 );
xor ( \650_b0 , \646_b0 , w_908 );
not ( w_908 , w_909 );
and ( w_909 , \649_b1 , \649_b0 );
or ( \651_b1 , \215_A[5]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_910 );
and ( \651_b0 , \215_A[5]_b0 , w_911 );
and ( w_910 , w_911 , \359_B[8]_b0 );
or ( \652_b1 , \650_b1 , \651_b1 );
xor ( \652_b0 , \650_b0 , w_912 );
not ( w_912 , w_913 );
and ( w_913 , \651_b1 , \651_b0 );
or ( \653_b1 , \580_b1 , \581_b1 );
not ( \581_b1 , w_914 );
and ( \653_b0 , \580_b0 , w_915 );
and ( w_914 , w_915 , \581_b0 );
or ( \654_b1 , \582_b1 , \585_b1 );
not ( \585_b1 , w_916 );
and ( \654_b0 , \582_b0 , w_917 );
and ( w_916 , w_917 , \585_b0 );
or ( \655_b1 , \653_b1 , w_918 );
or ( \655_b0 , \653_b0 , \654_b0 );
not ( \654_b0 , w_919 );
and ( w_919 , w_918 , \654_b1 );
or ( \656_b1 , \652_b1 , \655_b1 );
xor ( \656_b0 , \652_b0 , w_920 );
not ( w_920 , w_921 );
and ( w_921 , \655_b1 , \655_b0 );
or ( \657_b1 , \193_A[4]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_922 );
and ( \657_b0 , \193_A[4]_b0 , w_923 );
and ( w_922 , w_923 , \411_B[9]_b0 );
or ( \658_b1 , \656_b1 , \657_b1 );
xor ( \658_b0 , \656_b0 , w_924 );
not ( w_924 , w_925 );
and ( w_925 , \657_b1 , \657_b0 );
or ( \659_b1 , \586_b1 , \587_b1 );
not ( \587_b1 , w_926 );
and ( \659_b0 , \586_b0 , w_927 );
and ( w_926 , w_927 , \587_b0 );
or ( \660_b1 , \588_b1 , \591_b1 );
not ( \591_b1 , w_928 );
and ( \660_b0 , \588_b0 , w_929 );
and ( w_928 , w_929 , \591_b0 );
or ( \661_b1 , \659_b1 , w_930 );
or ( \661_b0 , \659_b0 , \660_b0 );
not ( \660_b0 , w_931 );
and ( w_931 , w_930 , \660_b1 );
or ( \662_b1 , \658_b1 , \661_b1 );
xor ( \662_b0 , \658_b0 , w_932 );
not ( w_932 , w_933 );
and ( w_933 , \661_b1 , \661_b0 );
or ( \663_b1 , \177_A[3]_b1 , \469_B[10]_b1 );
not ( \469_B[10]_b1 , w_934 );
and ( \663_b0 , \177_A[3]_b0 , w_935 );
and ( w_934 , w_935 , \469_B[10]_b0 );
or ( \664_b1 , \662_b1 , \663_b1 );
xor ( \664_b0 , \662_b0 , w_936 );
not ( w_936 , w_937 );
and ( w_937 , \663_b1 , \663_b0 );
or ( \665_b1 , \592_b1 , \593_b1 );
not ( \593_b1 , w_938 );
and ( \665_b0 , \592_b0 , w_939 );
and ( w_938 , w_939 , \593_b0 );
or ( \666_b1 , \594_b1 , \597_b1 );
not ( \597_b1 , w_940 );
and ( \666_b0 , \594_b0 , w_941 );
and ( w_940 , w_941 , \597_b0 );
or ( \667_b1 , \665_b1 , w_942 );
or ( \667_b0 , \665_b0 , \666_b0 );
not ( \666_b0 , w_943 );
and ( w_943 , w_942 , \666_b1 );
or ( \668_b1 , \664_b1 , \667_b1 );
xor ( \668_b0 , \664_b0 , w_944 );
not ( w_944 , w_945 );
and ( w_945 , \667_b1 , \667_b0 );
or ( \669_b1 , \167_A[2]_b1 , \533_B[11]_b1 );
not ( \533_B[11]_b1 , w_946 );
and ( \669_b0 , \167_A[2]_b0 , w_947 );
and ( w_946 , w_947 , \533_B[11]_b0 );
or ( \670_b1 , \668_b1 , \669_b1 );
xor ( \670_b0 , \668_b0 , w_948 );
not ( w_948 , w_949 );
and ( w_949 , \669_b1 , \669_b0 );
or ( \671_b1 , \598_b1 , \599_b1 );
not ( \599_b1 , w_950 );
and ( \671_b0 , \598_b0 , w_951 );
and ( w_950 , w_951 , \599_b0 );
or ( \672_b1 , \600_b1 , \601_b1 );
not ( \601_b1 , w_952 );
and ( \672_b0 , \600_b0 , w_953 );
and ( w_952 , w_953 , \601_b0 );
or ( \673_b1 , \671_b1 , w_954 );
or ( \673_b0 , \671_b0 , \672_b0 );
not ( \672_b0 , w_955 );
and ( w_955 , w_954 , \672_b1 );
or ( \674_b1 , \670_b1 , \673_b1 );
xor ( \674_b0 , \670_b0 , w_956 );
not ( w_956 , w_957 );
and ( w_957 , \673_b1 , \673_b0 );
or ( \675_b1 , \161_A[1]_b1 , \603_B[12]_b1 );
not ( \603_B[12]_b1 , w_958 );
and ( \675_b0 , \161_A[1]_b0 , w_959 );
and ( w_958 , w_959 , \603_B[12]_b0 );
or ( \676_b1 , \674_b1 , \675_b1 );
xor ( \676_b0 , \674_b0 , w_960 );
not ( w_960 , w_961 );
and ( w_961 , \675_b1 , \675_b0 );
or ( \677_b1 , \602_b1 , \604_b1 );
not ( \604_b1 , w_962 );
and ( \677_b0 , \602_b0 , w_963 );
and ( w_962 , w_963 , \604_b0 );
or ( \678_b1 , \676_b1 , \677_b1 );
xor ( \678_b0 , \676_b0 , w_964 );
not ( w_964 , w_965 );
and ( w_965 , \677_b1 , \677_b0 );
buf ( \679_B[13]_b1 , \b[13]_b1 );
buf ( \679_B[13]_b0 , \b[13]_b0 );
or ( \680_b1 , \156_A[0]_b1 , \679_B[13]_b1 );
not ( \679_B[13]_b1 , w_966 );
and ( \680_b0 , \156_A[0]_b0 , w_967 );
and ( w_966 , w_967 , \679_B[13]_b0 );
or ( \681_b1 , \678_b1 , \680_b1 );
xor ( \681_b0 , \678_b0 , w_968 );
not ( w_968 , w_969 );
and ( w_969 , \680_b1 , \680_b0 );
buf ( \682_Z[13]_b1 , \681_b1 );
buf ( \682_Z[13]_b0 , \681_b0 );
buf ( \683_A[14]_b1 , \a[14]_b1 );
buf ( \683_A[14]_b0 , \a[14]_b0 );
or ( \684_b1 , \683_A[14]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_970 );
and ( \684_b0 , \683_A[14]_b0 , w_971 );
and ( w_970 , w_971 , \157_B[0]_b0 );
or ( \685_b1 , \607_A[13]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_972 );
and ( \685_b0 , \607_A[13]_b0 , w_973 );
and ( w_972 , w_973 , \163_B[1]_b0 );
or ( \686_b1 , \684_b1 , \685_b1 );
xor ( \686_b0 , \684_b0 , w_974 );
not ( w_974 , w_975 );
and ( w_975 , \685_b1 , \685_b0 );
or ( \687_b1 , \608_b1 , \609_b1 );
not ( \609_b1 , w_976 );
and ( \687_b0 , \608_b0 , w_977 );
and ( w_976 , w_977 , \609_b0 );
or ( \688_b1 , \610_b1 , \613_b1 );
not ( \613_b1 , w_978 );
and ( \688_b0 , \610_b0 , w_979 );
and ( w_978 , w_979 , \613_b0 );
or ( \689_b1 , \687_b1 , w_980 );
or ( \689_b0 , \687_b0 , \688_b0 );
not ( \688_b0 , w_981 );
and ( w_981 , w_980 , \688_b1 );
or ( \690_b1 , \686_b1 , \689_b1 );
xor ( \690_b0 , \686_b0 , w_982 );
not ( w_982 , w_983 );
and ( w_983 , \689_b1 , \689_b0 );
or ( \691_b1 , \537_A[12]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_984 );
and ( \691_b0 , \537_A[12]_b0 , w_985 );
and ( w_984 , w_985 , \173_B[2]_b0 );
or ( \692_b1 , \690_b1 , \691_b1 );
xor ( \692_b0 , \690_b0 , w_986 );
not ( w_986 , w_987 );
and ( w_987 , \691_b1 , \691_b0 );
or ( \693_b1 , \614_b1 , \615_b1 );
not ( \615_b1 , w_988 );
and ( \693_b0 , \614_b0 , w_989 );
and ( w_988 , w_989 , \615_b0 );
or ( \694_b1 , \616_b1 , \619_b1 );
not ( \619_b1 , w_990 );
and ( \694_b0 , \616_b0 , w_991 );
and ( w_990 , w_991 , \619_b0 );
or ( \695_b1 , \693_b1 , w_992 );
or ( \695_b0 , \693_b0 , \694_b0 );
not ( \694_b0 , w_993 );
and ( w_993 , w_992 , \694_b1 );
or ( \696_b1 , \692_b1 , \695_b1 );
xor ( \696_b0 , \692_b0 , w_994 );
not ( w_994 , w_995 );
and ( w_995 , \695_b1 , \695_b0 );
or ( \697_b1 , \473_A[11]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_996 );
and ( \697_b0 , \473_A[11]_b0 , w_997 );
and ( w_996 , w_997 , \189_B[3]_b0 );
or ( \698_b1 , \696_b1 , \697_b1 );
xor ( \698_b0 , \696_b0 , w_998 );
not ( w_998 , w_999 );
and ( w_999 , \697_b1 , \697_b0 );
or ( \699_b1 , \620_b1 , \621_b1 );
not ( \621_b1 , w_1000 );
and ( \699_b0 , \620_b0 , w_1001 );
and ( w_1000 , w_1001 , \621_b0 );
or ( \700_b1 , \622_b1 , \625_b1 );
not ( \625_b1 , w_1002 );
and ( \700_b0 , \622_b0 , w_1003 );
and ( w_1002 , w_1003 , \625_b0 );
or ( \701_b1 , \699_b1 , w_1004 );
or ( \701_b0 , \699_b0 , \700_b0 );
not ( \700_b0 , w_1005 );
and ( w_1005 , w_1004 , \700_b1 );
or ( \702_b1 , \698_b1 , \701_b1 );
xor ( \702_b0 , \698_b0 , w_1006 );
not ( w_1006 , w_1007 );
and ( w_1007 , \701_b1 , \701_b0 );
or ( \703_b1 , \415_A[10]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_1008 );
and ( \703_b0 , \415_A[10]_b0 , w_1009 );
and ( w_1008 , w_1009 , \211_B[4]_b0 );
or ( \704_b1 , \702_b1 , \703_b1 );
xor ( \704_b0 , \702_b0 , w_1010 );
not ( w_1010 , w_1011 );
and ( w_1011 , \703_b1 , \703_b0 );
or ( \705_b1 , \626_b1 , \627_b1 );
not ( \627_b1 , w_1012 );
and ( \705_b0 , \626_b0 , w_1013 );
and ( w_1012 , w_1013 , \627_b0 );
or ( \706_b1 , \628_b1 , \631_b1 );
not ( \631_b1 , w_1014 );
and ( \706_b0 , \628_b0 , w_1015 );
and ( w_1014 , w_1015 , \631_b0 );
or ( \707_b1 , \705_b1 , w_1016 );
or ( \707_b0 , \705_b0 , \706_b0 );
not ( \706_b0 , w_1017 );
and ( w_1017 , w_1016 , \706_b1 );
or ( \708_b1 , \704_b1 , \707_b1 );
xor ( \708_b0 , \704_b0 , w_1018 );
not ( w_1018 , w_1019 );
and ( w_1019 , \707_b1 , \707_b0 );
or ( \709_b1 , \363_A[9]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_1020 );
and ( \709_b0 , \363_A[9]_b0 , w_1021 );
and ( w_1020 , w_1021 , \239_B[5]_b0 );
or ( \710_b1 , \708_b1 , \709_b1 );
xor ( \710_b0 , \708_b0 , w_1022 );
not ( w_1022 , w_1023 );
and ( w_1023 , \709_b1 , \709_b0 );
or ( \711_b1 , \632_b1 , \633_b1 );
not ( \633_b1 , w_1024 );
and ( \711_b0 , \632_b0 , w_1025 );
and ( w_1024 , w_1025 , \633_b0 );
or ( \712_b1 , \634_b1 , \637_b1 );
not ( \637_b1 , w_1026 );
and ( \712_b0 , \634_b0 , w_1027 );
and ( w_1026 , w_1027 , \637_b0 );
or ( \713_b1 , \711_b1 , w_1028 );
or ( \713_b0 , \711_b0 , \712_b0 );
not ( \712_b0 , w_1029 );
and ( w_1029 , w_1028 , \712_b1 );
or ( \714_b1 , \710_b1 , \713_b1 );
xor ( \714_b0 , \710_b0 , w_1030 );
not ( w_1030 , w_1031 );
and ( w_1031 , \713_b1 , \713_b0 );
or ( \715_b1 , \317_A[8]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_1032 );
and ( \715_b0 , \317_A[8]_b0 , w_1033 );
and ( w_1032 , w_1033 , \273_B[6]_b0 );
or ( \716_b1 , \714_b1 , \715_b1 );
xor ( \716_b0 , \714_b0 , w_1034 );
not ( w_1034 , w_1035 );
and ( w_1035 , \715_b1 , \715_b0 );
or ( \717_b1 , \638_b1 , \639_b1 );
not ( \639_b1 , w_1036 );
and ( \717_b0 , \638_b0 , w_1037 );
and ( w_1036 , w_1037 , \639_b0 );
or ( \718_b1 , \640_b1 , \643_b1 );
not ( \643_b1 , w_1038 );
and ( \718_b0 , \640_b0 , w_1039 );
and ( w_1038 , w_1039 , \643_b0 );
or ( \719_b1 , \717_b1 , w_1040 );
or ( \719_b0 , \717_b0 , \718_b0 );
not ( \718_b0 , w_1041 );
and ( w_1041 , w_1040 , \718_b1 );
or ( \720_b1 , \716_b1 , \719_b1 );
xor ( \720_b0 , \716_b0 , w_1042 );
not ( w_1042 , w_1043 );
and ( w_1043 , \719_b1 , \719_b0 );
or ( \721_b1 , \277_A[7]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_1044 );
and ( \721_b0 , \277_A[7]_b0 , w_1045 );
and ( w_1044 , w_1045 , \313_B[7]_b0 );
or ( \722_b1 , \720_b1 , \721_b1 );
xor ( \722_b0 , \720_b0 , w_1046 );
not ( w_1046 , w_1047 );
and ( w_1047 , \721_b1 , \721_b0 );
or ( \723_b1 , \644_b1 , \645_b1 );
not ( \645_b1 , w_1048 );
and ( \723_b0 , \644_b0 , w_1049 );
and ( w_1048 , w_1049 , \645_b0 );
or ( \724_b1 , \646_b1 , \649_b1 );
not ( \649_b1 , w_1050 );
and ( \724_b0 , \646_b0 , w_1051 );
and ( w_1050 , w_1051 , \649_b0 );
or ( \725_b1 , \723_b1 , w_1052 );
or ( \725_b0 , \723_b0 , \724_b0 );
not ( \724_b0 , w_1053 );
and ( w_1053 , w_1052 , \724_b1 );
or ( \726_b1 , \722_b1 , \725_b1 );
xor ( \726_b0 , \722_b0 , w_1054 );
not ( w_1054 , w_1055 );
and ( w_1055 , \725_b1 , \725_b0 );
or ( \727_b1 , \243_A[6]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_1056 );
and ( \727_b0 , \243_A[6]_b0 , w_1057 );
and ( w_1056 , w_1057 , \359_B[8]_b0 );
or ( \728_b1 , \726_b1 , \727_b1 );
xor ( \728_b0 , \726_b0 , w_1058 );
not ( w_1058 , w_1059 );
and ( w_1059 , \727_b1 , \727_b0 );
or ( \729_b1 , \650_b1 , \651_b1 );
not ( \651_b1 , w_1060 );
and ( \729_b0 , \650_b0 , w_1061 );
and ( w_1060 , w_1061 , \651_b0 );
or ( \730_b1 , \652_b1 , \655_b1 );
not ( \655_b1 , w_1062 );
and ( \730_b0 , \652_b0 , w_1063 );
and ( w_1062 , w_1063 , \655_b0 );
or ( \731_b1 , \729_b1 , w_1064 );
or ( \731_b0 , \729_b0 , \730_b0 );
not ( \730_b0 , w_1065 );
and ( w_1065 , w_1064 , \730_b1 );
or ( \732_b1 , \728_b1 , \731_b1 );
xor ( \732_b0 , \728_b0 , w_1066 );
not ( w_1066 , w_1067 );
and ( w_1067 , \731_b1 , \731_b0 );
or ( \733_b1 , \215_A[5]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_1068 );
and ( \733_b0 , \215_A[5]_b0 , w_1069 );
and ( w_1068 , w_1069 , \411_B[9]_b0 );
or ( \734_b1 , \732_b1 , \733_b1 );
xor ( \734_b0 , \732_b0 , w_1070 );
not ( w_1070 , w_1071 );
and ( w_1071 , \733_b1 , \733_b0 );
or ( \735_b1 , \656_b1 , \657_b1 );
not ( \657_b1 , w_1072 );
and ( \735_b0 , \656_b0 , w_1073 );
and ( w_1072 , w_1073 , \657_b0 );
or ( \736_b1 , \658_b1 , \661_b1 );
not ( \661_b1 , w_1074 );
and ( \736_b0 , \658_b0 , w_1075 );
and ( w_1074 , w_1075 , \661_b0 );
or ( \737_b1 , \735_b1 , w_1076 );
or ( \737_b0 , \735_b0 , \736_b0 );
not ( \736_b0 , w_1077 );
and ( w_1077 , w_1076 , \736_b1 );
or ( \738_b1 , \734_b1 , \737_b1 );
xor ( \738_b0 , \734_b0 , w_1078 );
not ( w_1078 , w_1079 );
and ( w_1079 , \737_b1 , \737_b0 );
or ( \739_b1 , \193_A[4]_b1 , \469_B[10]_b1 );
not ( \469_B[10]_b1 , w_1080 );
and ( \739_b0 , \193_A[4]_b0 , w_1081 );
and ( w_1080 , w_1081 , \469_B[10]_b0 );
or ( \740_b1 , \738_b1 , \739_b1 );
xor ( \740_b0 , \738_b0 , w_1082 );
not ( w_1082 , w_1083 );
and ( w_1083 , \739_b1 , \739_b0 );
or ( \741_b1 , \662_b1 , \663_b1 );
not ( \663_b1 , w_1084 );
and ( \741_b0 , \662_b0 , w_1085 );
and ( w_1084 , w_1085 , \663_b0 );
or ( \742_b1 , \664_b1 , \667_b1 );
not ( \667_b1 , w_1086 );
and ( \742_b0 , \664_b0 , w_1087 );
and ( w_1086 , w_1087 , \667_b0 );
or ( \743_b1 , \741_b1 , w_1088 );
or ( \743_b0 , \741_b0 , \742_b0 );
not ( \742_b0 , w_1089 );
and ( w_1089 , w_1088 , \742_b1 );
or ( \744_b1 , \740_b1 , \743_b1 );
xor ( \744_b0 , \740_b0 , w_1090 );
not ( w_1090 , w_1091 );
and ( w_1091 , \743_b1 , \743_b0 );
or ( \745_b1 , \177_A[3]_b1 , \533_B[11]_b1 );
not ( \533_B[11]_b1 , w_1092 );
and ( \745_b0 , \177_A[3]_b0 , w_1093 );
and ( w_1092 , w_1093 , \533_B[11]_b0 );
or ( \746_b1 , \744_b1 , \745_b1 );
xor ( \746_b0 , \744_b0 , w_1094 );
not ( w_1094 , w_1095 );
and ( w_1095 , \745_b1 , \745_b0 );
or ( \747_b1 , \668_b1 , \669_b1 );
not ( \669_b1 , w_1096 );
and ( \747_b0 , \668_b0 , w_1097 );
and ( w_1096 , w_1097 , \669_b0 );
or ( \748_b1 , \670_b1 , \673_b1 );
not ( \673_b1 , w_1098 );
and ( \748_b0 , \670_b0 , w_1099 );
and ( w_1098 , w_1099 , \673_b0 );
or ( \749_b1 , \747_b1 , w_1100 );
or ( \749_b0 , \747_b0 , \748_b0 );
not ( \748_b0 , w_1101 );
and ( w_1101 , w_1100 , \748_b1 );
or ( \750_b1 , \746_b1 , \749_b1 );
xor ( \750_b0 , \746_b0 , w_1102 );
not ( w_1102 , w_1103 );
and ( w_1103 , \749_b1 , \749_b0 );
or ( \751_b1 , \167_A[2]_b1 , \603_B[12]_b1 );
not ( \603_B[12]_b1 , w_1104 );
and ( \751_b0 , \167_A[2]_b0 , w_1105 );
and ( w_1104 , w_1105 , \603_B[12]_b0 );
or ( \752_b1 , \750_b1 , \751_b1 );
xor ( \752_b0 , \750_b0 , w_1106 );
not ( w_1106 , w_1107 );
and ( w_1107 , \751_b1 , \751_b0 );
or ( \753_b1 , \674_b1 , \675_b1 );
not ( \675_b1 , w_1108 );
and ( \753_b0 , \674_b0 , w_1109 );
and ( w_1108 , w_1109 , \675_b0 );
or ( \754_b1 , \676_b1 , \677_b1 );
not ( \677_b1 , w_1110 );
and ( \754_b0 , \676_b0 , w_1111 );
and ( w_1110 , w_1111 , \677_b0 );
or ( \755_b1 , \753_b1 , w_1112 );
or ( \755_b0 , \753_b0 , \754_b0 );
not ( \754_b0 , w_1113 );
and ( w_1113 , w_1112 , \754_b1 );
or ( \756_b1 , \752_b1 , \755_b1 );
xor ( \756_b0 , \752_b0 , w_1114 );
not ( w_1114 , w_1115 );
and ( w_1115 , \755_b1 , \755_b0 );
or ( \757_b1 , \161_A[1]_b1 , \679_B[13]_b1 );
not ( \679_B[13]_b1 , w_1116 );
and ( \757_b0 , \161_A[1]_b0 , w_1117 );
and ( w_1116 , w_1117 , \679_B[13]_b0 );
or ( \758_b1 , \756_b1 , \757_b1 );
xor ( \758_b0 , \756_b0 , w_1118 );
not ( w_1118 , w_1119 );
and ( w_1119 , \757_b1 , \757_b0 );
or ( \759_b1 , \678_b1 , \680_b1 );
not ( \680_b1 , w_1120 );
and ( \759_b0 , \678_b0 , w_1121 );
and ( w_1120 , w_1121 , \680_b0 );
or ( \760_b1 , \758_b1 , \759_b1 );
xor ( \760_b0 , \758_b0 , w_1122 );
not ( w_1122 , w_1123 );
and ( w_1123 , \759_b1 , \759_b0 );
buf ( \761_B[14]_b1 , \b[14]_b1 );
buf ( \761_B[14]_b0 , \b[14]_b0 );
or ( \762_b1 , \156_A[0]_b1 , \761_B[14]_b1 );
not ( \761_B[14]_b1 , w_1124 );
and ( \762_b0 , \156_A[0]_b0 , w_1125 );
and ( w_1124 , w_1125 , \761_B[14]_b0 );
or ( \763_b1 , \760_b1 , \762_b1 );
xor ( \763_b0 , \760_b0 , w_1126 );
not ( w_1126 , w_1127 );
and ( w_1127 , \762_b1 , \762_b0 );
buf ( \764_Z[14]_b1 , \763_b1 );
buf ( \764_Z[14]_b0 , \763_b0 );
buf ( \765_A[15]_b1 , \a[15]_b1 );
buf ( \765_A[15]_b0 , \a[15]_b0 );
or ( \766_b1 , \765_A[15]_b1 , \157_B[0]_b1 );
not ( \157_B[0]_b1 , w_1128 );
and ( \766_b0 , \765_A[15]_b0 , w_1129 );
and ( w_1128 , w_1129 , \157_B[0]_b0 );
or ( \767_b1 , \683_A[14]_b1 , \163_B[1]_b1 );
not ( \163_B[1]_b1 , w_1130 );
and ( \767_b0 , \683_A[14]_b0 , w_1131 );
and ( w_1130 , w_1131 , \163_B[1]_b0 );
or ( \768_b1 , \766_b1 , \767_b1 );
xor ( \768_b0 , \766_b0 , w_1132 );
not ( w_1132 , w_1133 );
and ( w_1133 , \767_b1 , \767_b0 );
or ( \769_b1 , \684_b1 , \685_b1 );
not ( \685_b1 , w_1134 );
and ( \769_b0 , \684_b0 , w_1135 );
and ( w_1134 , w_1135 , \685_b0 );
or ( \770_b1 , \686_b1 , \689_b1 );
not ( \689_b1 , w_1136 );
and ( \770_b0 , \686_b0 , w_1137 );
and ( w_1136 , w_1137 , \689_b0 );
or ( \771_b1 , \769_b1 , w_1138 );
or ( \771_b0 , \769_b0 , \770_b0 );
not ( \770_b0 , w_1139 );
and ( w_1139 , w_1138 , \770_b1 );
or ( \772_b1 , \768_b1 , \771_b1 );
xor ( \772_b0 , \768_b0 , w_1140 );
not ( w_1140 , w_1141 );
and ( w_1141 , \771_b1 , \771_b0 );
or ( \773_b1 , \607_A[13]_b1 , \173_B[2]_b1 );
not ( \173_B[2]_b1 , w_1142 );
and ( \773_b0 , \607_A[13]_b0 , w_1143 );
and ( w_1142 , w_1143 , \173_B[2]_b0 );
or ( \774_b1 , \772_b1 , \773_b1 );
xor ( \774_b0 , \772_b0 , w_1144 );
not ( w_1144 , w_1145 );
and ( w_1145 , \773_b1 , \773_b0 );
or ( \775_b1 , \690_b1 , \691_b1 );
not ( \691_b1 , w_1146 );
and ( \775_b0 , \690_b0 , w_1147 );
and ( w_1146 , w_1147 , \691_b0 );
or ( \776_b1 , \692_b1 , \695_b1 );
not ( \695_b1 , w_1148 );
and ( \776_b0 , \692_b0 , w_1149 );
and ( w_1148 , w_1149 , \695_b0 );
or ( \777_b1 , \775_b1 , w_1150 );
or ( \777_b0 , \775_b0 , \776_b0 );
not ( \776_b0 , w_1151 );
and ( w_1151 , w_1150 , \776_b1 );
or ( \778_b1 , \774_b1 , \777_b1 );
xor ( \778_b0 , \774_b0 , w_1152 );
not ( w_1152 , w_1153 );
and ( w_1153 , \777_b1 , \777_b0 );
or ( \779_b1 , \537_A[12]_b1 , \189_B[3]_b1 );
not ( \189_B[3]_b1 , w_1154 );
and ( \779_b0 , \537_A[12]_b0 , w_1155 );
and ( w_1154 , w_1155 , \189_B[3]_b0 );
or ( \780_b1 , \778_b1 , \779_b1 );
xor ( \780_b0 , \778_b0 , w_1156 );
not ( w_1156 , w_1157 );
and ( w_1157 , \779_b1 , \779_b0 );
or ( \781_b1 , \696_b1 , \697_b1 );
not ( \697_b1 , w_1158 );
and ( \781_b0 , \696_b0 , w_1159 );
and ( w_1158 , w_1159 , \697_b0 );
or ( \782_b1 , \698_b1 , \701_b1 );
not ( \701_b1 , w_1160 );
and ( \782_b0 , \698_b0 , w_1161 );
and ( w_1160 , w_1161 , \701_b0 );
or ( \783_b1 , \781_b1 , w_1162 );
or ( \783_b0 , \781_b0 , \782_b0 );
not ( \782_b0 , w_1163 );
and ( w_1163 , w_1162 , \782_b1 );
or ( \784_b1 , \780_b1 , \783_b1 );
xor ( \784_b0 , \780_b0 , w_1164 );
not ( w_1164 , w_1165 );
and ( w_1165 , \783_b1 , \783_b0 );
or ( \785_b1 , \473_A[11]_b1 , \211_B[4]_b1 );
not ( \211_B[4]_b1 , w_1166 );
and ( \785_b0 , \473_A[11]_b0 , w_1167 );
and ( w_1166 , w_1167 , \211_B[4]_b0 );
or ( \786_b1 , \784_b1 , \785_b1 );
xor ( \786_b0 , \784_b0 , w_1168 );
not ( w_1168 , w_1169 );
and ( w_1169 , \785_b1 , \785_b0 );
or ( \787_b1 , \702_b1 , \703_b1 );
not ( \703_b1 , w_1170 );
and ( \787_b0 , \702_b0 , w_1171 );
and ( w_1170 , w_1171 , \703_b0 );
or ( \788_b1 , \704_b1 , \707_b1 );
not ( \707_b1 , w_1172 );
and ( \788_b0 , \704_b0 , w_1173 );
and ( w_1172 , w_1173 , \707_b0 );
or ( \789_b1 , \787_b1 , w_1174 );
or ( \789_b0 , \787_b0 , \788_b0 );
not ( \788_b0 , w_1175 );
and ( w_1175 , w_1174 , \788_b1 );
or ( \790_b1 , \786_b1 , \789_b1 );
xor ( \790_b0 , \786_b0 , w_1176 );
not ( w_1176 , w_1177 );
and ( w_1177 , \789_b1 , \789_b0 );
or ( \791_b1 , \415_A[10]_b1 , \239_B[5]_b1 );
not ( \239_B[5]_b1 , w_1178 );
and ( \791_b0 , \415_A[10]_b0 , w_1179 );
and ( w_1178 , w_1179 , \239_B[5]_b0 );
or ( \792_b1 , \790_b1 , \791_b1 );
xor ( \792_b0 , \790_b0 , w_1180 );
not ( w_1180 , w_1181 );
and ( w_1181 , \791_b1 , \791_b0 );
or ( \793_b1 , \708_b1 , \709_b1 );
not ( \709_b1 , w_1182 );
and ( \793_b0 , \708_b0 , w_1183 );
and ( w_1182 , w_1183 , \709_b0 );
or ( \794_b1 , \710_b1 , \713_b1 );
not ( \713_b1 , w_1184 );
and ( \794_b0 , \710_b0 , w_1185 );
and ( w_1184 , w_1185 , \713_b0 );
or ( \795_b1 , \793_b1 , w_1186 );
or ( \795_b0 , \793_b0 , \794_b0 );
not ( \794_b0 , w_1187 );
and ( w_1187 , w_1186 , \794_b1 );
or ( \796_b1 , \792_b1 , \795_b1 );
xor ( \796_b0 , \792_b0 , w_1188 );
not ( w_1188 , w_1189 );
and ( w_1189 , \795_b1 , \795_b0 );
or ( \797_b1 , \363_A[9]_b1 , \273_B[6]_b1 );
not ( \273_B[6]_b1 , w_1190 );
and ( \797_b0 , \363_A[9]_b0 , w_1191 );
and ( w_1190 , w_1191 , \273_B[6]_b0 );
or ( \798_b1 , \796_b1 , \797_b1 );
xor ( \798_b0 , \796_b0 , w_1192 );
not ( w_1192 , w_1193 );
and ( w_1193 , \797_b1 , \797_b0 );
or ( \799_b1 , \714_b1 , \715_b1 );
not ( \715_b1 , w_1194 );
and ( \799_b0 , \714_b0 , w_1195 );
and ( w_1194 , w_1195 , \715_b0 );
or ( \800_b1 , \716_b1 , \719_b1 );
not ( \719_b1 , w_1196 );
and ( \800_b0 , \716_b0 , w_1197 );
and ( w_1196 , w_1197 , \719_b0 );
or ( \801_b1 , \799_b1 , w_1198 );
or ( \801_b0 , \799_b0 , \800_b0 );
not ( \800_b0 , w_1199 );
and ( w_1199 , w_1198 , \800_b1 );
or ( \802_b1 , \798_b1 , \801_b1 );
xor ( \802_b0 , \798_b0 , w_1200 );
not ( w_1200 , w_1201 );
and ( w_1201 , \801_b1 , \801_b0 );
or ( \803_b1 , \317_A[8]_b1 , \313_B[7]_b1 );
not ( \313_B[7]_b1 , w_1202 );
and ( \803_b0 , \317_A[8]_b0 , w_1203 );
and ( w_1202 , w_1203 , \313_B[7]_b0 );
or ( \804_b1 , \802_b1 , \803_b1 );
xor ( \804_b0 , \802_b0 , w_1204 );
not ( w_1204 , w_1205 );
and ( w_1205 , \803_b1 , \803_b0 );
or ( \805_b1 , \720_b1 , \721_b1 );
not ( \721_b1 , w_1206 );
and ( \805_b0 , \720_b0 , w_1207 );
and ( w_1206 , w_1207 , \721_b0 );
or ( \806_b1 , \722_b1 , \725_b1 );
not ( \725_b1 , w_1208 );
and ( \806_b0 , \722_b0 , w_1209 );
and ( w_1208 , w_1209 , \725_b0 );
or ( \807_b1 , \805_b1 , w_1210 );
or ( \807_b0 , \805_b0 , \806_b0 );
not ( \806_b0 , w_1211 );
and ( w_1211 , w_1210 , \806_b1 );
or ( \808_b1 , \804_b1 , \807_b1 );
xor ( \808_b0 , \804_b0 , w_1212 );
not ( w_1212 , w_1213 );
and ( w_1213 , \807_b1 , \807_b0 );
or ( \809_b1 , \277_A[7]_b1 , \359_B[8]_b1 );
not ( \359_B[8]_b1 , w_1214 );
and ( \809_b0 , \277_A[7]_b0 , w_1215 );
and ( w_1214 , w_1215 , \359_B[8]_b0 );
or ( \810_b1 , \808_b1 , \809_b1 );
xor ( \810_b0 , \808_b0 , w_1216 );
not ( w_1216 , w_1217 );
and ( w_1217 , \809_b1 , \809_b0 );
or ( \811_b1 , \726_b1 , \727_b1 );
not ( \727_b1 , w_1218 );
and ( \811_b0 , \726_b0 , w_1219 );
and ( w_1218 , w_1219 , \727_b0 );
or ( \812_b1 , \728_b1 , \731_b1 );
not ( \731_b1 , w_1220 );
and ( \812_b0 , \728_b0 , w_1221 );
and ( w_1220 , w_1221 , \731_b0 );
or ( \813_b1 , \811_b1 , w_1222 );
or ( \813_b0 , \811_b0 , \812_b0 );
not ( \812_b0 , w_1223 );
and ( w_1223 , w_1222 , \812_b1 );
or ( \814_b1 , \810_b1 , \813_b1 );
xor ( \814_b0 , \810_b0 , w_1224 );
not ( w_1224 , w_1225 );
and ( w_1225 , \813_b1 , \813_b0 );
or ( \815_b1 , \243_A[6]_b1 , \411_B[9]_b1 );
not ( \411_B[9]_b1 , w_1226 );
and ( \815_b0 , \243_A[6]_b0 , w_1227 );
and ( w_1226 , w_1227 , \411_B[9]_b0 );
or ( \816_b1 , \814_b1 , \815_b1 );
xor ( \816_b0 , \814_b0 , w_1228 );
not ( w_1228 , w_1229 );
and ( w_1229 , \815_b1 , \815_b0 );
or ( \817_b1 , \732_b1 , \733_b1 );
not ( \733_b1 , w_1230 );
and ( \817_b0 , \732_b0 , w_1231 );
and ( w_1230 , w_1231 , \733_b0 );
or ( \818_b1 , \734_b1 , \737_b1 );
not ( \737_b1 , w_1232 );
and ( \818_b0 , \734_b0 , w_1233 );
and ( w_1232 , w_1233 , \737_b0 );
or ( \819_b1 , \817_b1 , w_1234 );
or ( \819_b0 , \817_b0 , \818_b0 );
not ( \818_b0 , w_1235 );
and ( w_1235 , w_1234 , \818_b1 );
or ( \820_b1 , \816_b1 , \819_b1 );
xor ( \820_b0 , \816_b0 , w_1236 );
not ( w_1236 , w_1237 );
and ( w_1237 , \819_b1 , \819_b0 );
or ( \821_b1 , \215_A[5]_b1 , \469_B[10]_b1 );
not ( \469_B[10]_b1 , w_1238 );
and ( \821_b0 , \215_A[5]_b0 , w_1239 );
and ( w_1238 , w_1239 , \469_B[10]_b0 );
or ( \822_b1 , \820_b1 , \821_b1 );
xor ( \822_b0 , \820_b0 , w_1240 );
not ( w_1240 , w_1241 );
and ( w_1241 , \821_b1 , \821_b0 );
or ( \823_b1 , \738_b1 , \739_b1 );
not ( \739_b1 , w_1242 );
and ( \823_b0 , \738_b0 , w_1243 );
and ( w_1242 , w_1243 , \739_b0 );
or ( \824_b1 , \740_b1 , \743_b1 );
not ( \743_b1 , w_1244 );
and ( \824_b0 , \740_b0 , w_1245 );
and ( w_1244 , w_1245 , \743_b0 );
or ( \825_b1 , \823_b1 , w_1246 );
or ( \825_b0 , \823_b0 , \824_b0 );
not ( \824_b0 , w_1247 );
and ( w_1247 , w_1246 , \824_b1 );
or ( \826_b1 , \822_b1 , \825_b1 );
xor ( \826_b0 , \822_b0 , w_1248 );
not ( w_1248 , w_1249 );
and ( w_1249 , \825_b1 , \825_b0 );
or ( \827_b1 , \193_A[4]_b1 , \533_B[11]_b1 );
not ( \533_B[11]_b1 , w_1250 );
and ( \827_b0 , \193_A[4]_b0 , w_1251 );
and ( w_1250 , w_1251 , \533_B[11]_b0 );
or ( \828_b1 , \826_b1 , \827_b1 );
xor ( \828_b0 , \826_b0 , w_1252 );
not ( w_1252 , w_1253 );
and ( w_1253 , \827_b1 , \827_b0 );
or ( \829_b1 , \744_b1 , \745_b1 );
not ( \745_b1 , w_1254 );
and ( \829_b0 , \744_b0 , w_1255 );
and ( w_1254 , w_1255 , \745_b0 );
or ( \830_b1 , \746_b1 , \749_b1 );
not ( \749_b1 , w_1256 );
and ( \830_b0 , \746_b0 , w_1257 );
and ( w_1256 , w_1257 , \749_b0 );
or ( \831_b1 , \829_b1 , w_1258 );
or ( \831_b0 , \829_b0 , \830_b0 );
not ( \830_b0 , w_1259 );
and ( w_1259 , w_1258 , \830_b1 );
or ( \832_b1 , \828_b1 , \831_b1 );
xor ( \832_b0 , \828_b0 , w_1260 );
not ( w_1260 , w_1261 );
and ( w_1261 , \831_b1 , \831_b0 );
or ( \833_b1 , \177_A[3]_b1 , \603_B[12]_b1 );
not ( \603_B[12]_b1 , w_1262 );
and ( \833_b0 , \177_A[3]_b0 , w_1263 );
and ( w_1262 , w_1263 , \603_B[12]_b0 );
or ( \834_b1 , \832_b1 , \833_b1 );
xor ( \834_b0 , \832_b0 , w_1264 );
not ( w_1264 , w_1265 );
and ( w_1265 , \833_b1 , \833_b0 );
or ( \835_b1 , \750_b1 , \751_b1 );
not ( \751_b1 , w_1266 );
and ( \835_b0 , \750_b0 , w_1267 );
and ( w_1266 , w_1267 , \751_b0 );
or ( \836_b1 , \752_b1 , \755_b1 );
not ( \755_b1 , w_1268 );
and ( \836_b0 , \752_b0 , w_1269 );
and ( w_1268 , w_1269 , \755_b0 );
or ( \837_b1 , \835_b1 , w_1270 );
or ( \837_b0 , \835_b0 , \836_b0 );
not ( \836_b0 , w_1271 );
and ( w_1271 , w_1270 , \836_b1 );
or ( \838_b1 , \834_b1 , \837_b1 );
xor ( \838_b0 , \834_b0 , w_1272 );
not ( w_1272 , w_1273 );
and ( w_1273 , \837_b1 , \837_b0 );
or ( \839_b1 , \167_A[2]_b1 , \679_B[13]_b1 );
not ( \679_B[13]_b1 , w_1274 );
and ( \839_b0 , \167_A[2]_b0 , w_1275 );
and ( w_1274 , w_1275 , \679_B[13]_b0 );
or ( \840_b1 , \838_b1 , \839_b1 );
xor ( \840_b0 , \838_b0 , w_1276 );
not ( w_1276 , w_1277 );
and ( w_1277 , \839_b1 , \839_b0 );
or ( \841_b1 , \756_b1 , \757_b1 );
not ( \757_b1 , w_1278 );
and ( \841_b0 , \756_b0 , w_1279 );
and ( w_1278 , w_1279 , \757_b0 );
or ( \842_b1 , \758_b1 , \759_b1 );
not ( \759_b1 , w_1280 );
and ( \842_b0 , \758_b0 , w_1281 );
and ( w_1280 , w_1281 , \759_b0 );
or ( \843_b1 , \841_b1 , w_1282 );
or ( \843_b0 , \841_b0 , \842_b0 );
not ( \842_b0 , w_1283 );
and ( w_1283 , w_1282 , \842_b1 );
or ( \844_b1 , \840_b1 , \843_b1 );
xor ( \844_b0 , \840_b0 , w_1284 );
not ( w_1284 , w_1285 );
and ( w_1285 , \843_b1 , \843_b0 );
or ( \845_b1 , \161_A[1]_b1 , \761_B[14]_b1 );
not ( \761_B[14]_b1 , w_1286 );
and ( \845_b0 , \161_A[1]_b0 , w_1287 );
and ( w_1286 , w_1287 , \761_B[14]_b0 );
or ( \846_b1 , \844_b1 , \845_b1 );
xor ( \846_b0 , \844_b0 , w_1288 );
not ( w_1288 , w_1289 );
and ( w_1289 , \845_b1 , \845_b0 );
or ( \847_b1 , \760_b1 , \762_b1 );
not ( \762_b1 , w_1290 );
and ( \847_b0 , \760_b0 , w_1291 );
and ( w_1290 , w_1291 , \762_b0 );
or ( \848_b1 , \846_b1 , \847_b1 );
xor ( \848_b0 , \846_b0 , w_1292 );
not ( w_1292 , w_1293 );
and ( w_1293 , \847_b1 , \847_b0 );
buf ( \849_B[15]_b1 , \b[15]_b1 );
buf ( \849_B[15]_b0 , \b[15]_b0 );
or ( \850_b1 , \156_A[0]_b1 , \849_B[15]_b1 );
not ( \849_B[15]_b1 , w_1294 );
and ( \850_b0 , \156_A[0]_b0 , w_1295 );
and ( w_1294 , w_1295 , \849_B[15]_b0 );
or ( \851_b1 , \848_b1 , \850_b1 );
xor ( \851_b0 , \848_b0 , w_1296 );
not ( w_1296 , w_1297 );
and ( w_1297 , \850_b1 , \850_b0 );
buf ( \852_Z[15]_b1 , \851_b1 );
buf ( \852_Z[15]_b0 , \851_b0 );
buf ( \854_b1 , \166_Z[1]_b1 );
not ( \854_b1 , w_1298 );
not ( \854_b0 , w_1299 );
and ( w_1298 , w_1299 , \166_Z[1]_b0 );
buf ( \856_b1 , \176_Z[2]_b1 );
not ( \856_b1 , w_1300 );
not ( \856_b0 , w_1301 );
and ( w_1300 , w_1301 , \176_Z[2]_b0 );
buf ( \858_b1 , \192_Z[3]_b1 );
not ( \858_b1 , w_1302 );
not ( \858_b0 , w_1303 );
and ( w_1302 , w_1303 , \192_Z[3]_b0 );
buf ( \860_b1 , \214_Z[4]_b1 );
not ( \860_b1 , w_1304 );
not ( \860_b0 , w_1305 );
and ( w_1304 , w_1305 , \214_Z[4]_b0 );
buf ( \862_b1 , \242_Z[5]_b1 );
not ( \862_b1 , w_1306 );
not ( \862_b0 , w_1307 );
and ( w_1306 , w_1307 , \242_Z[5]_b0 );
buf ( \864_b1 , \276_Z[6]_b1 );
not ( \864_b1 , w_1308 );
not ( \864_b0 , w_1309 );
and ( w_1308 , w_1309 , \276_Z[6]_b0 );
buf ( \866_b1 , \316_Z[7]_b1 );
not ( \866_b1 , w_1310 );
not ( \866_b0 , w_1311 );
and ( w_1310 , w_1311 , \316_Z[7]_b0 );
buf ( \868_b1 , \362_Z[8]_b1 );
not ( \868_b1 , w_1312 );
not ( \868_b0 , w_1313 );
and ( w_1312 , w_1313 , \362_Z[8]_b0 );
buf ( \870_b1 , \414_Z[9]_b1 );
not ( \870_b1 , w_1314 );
not ( \870_b0 , w_1315 );
and ( w_1314 , w_1315 , \414_Z[9]_b0 );
buf ( \872_b1 , \472_Z[10]_b1 );
not ( \872_b1 , w_1316 );
not ( \872_b0 , w_1317 );
and ( w_1316 , w_1317 , \472_Z[10]_b0 );
buf ( \874_b1 , \536_Z[11]_b1 );
not ( \874_b1 , w_1318 );
not ( \874_b0 , w_1319 );
and ( w_1318 , w_1319 , \536_Z[11]_b0 );
and ( \877_b1 , 1'b0_b1 , w_1320 );
xor ( w_1320 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1321 );
and ( \877_b0 , w_1321 , \876_b0 );
or ( \878_b1 , \a[0]_b1 , w_1322 );
or ( \878_b0 , \a[0]_b0 , \d[0]_b0 );
not ( \d[0]_b0 , w_1323 );
and ( w_1323 , w_1322 , \d[0]_b1 );
or ( \879_b1 , \878_b1 , \875_b1 );
not ( \875_b1 , w_1324 );
and ( \879_b0 , \878_b0 , w_1325 );
and ( w_1324 , w_1325 , \875_b0 );
or ( \880_b1 , \b[0]_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_1326 );
and ( \880_b0 , \b[0]_b0 , w_1327 );
and ( w_1326 , w_1327 , \c[0]_b0 );
or ( \881_b1 , \880_b1 , \873_b1 );
not ( \873_b1 , w_1328 );
and ( \881_b0 , \880_b0 , w_1329 );
and ( w_1328 , w_1329 , \873_b0 );
or ( \882_b1 , \a[0]_b1 , w_1330 );
or ( \882_b0 , \a[0]_b0 , \b[0]_b0 );
not ( \b[0]_b0 , w_1331 );
and ( w_1331 , w_1330 , \b[0]_b1 );
or ( \883_b1 , \882_b1 , \871_b1 );
not ( \871_b1 , w_1332 );
and ( \883_b0 , \882_b0 , w_1333 );
and ( w_1332 , w_1333 , \871_b0 );
or ( \884_b1 , \c[0]_b1 , \d[0]_b1 );
xor ( \884_b0 , \c[0]_b0 , w_1334 );
not ( w_1334 , w_1335 );
and ( w_1335 , \d[0]_b1 , \d[0]_b0 );
or ( \885_b1 , \884_b1 , \869_b1 );
not ( \869_b1 , w_1336 );
and ( \885_b0 , \884_b0 , w_1337 );
and ( w_1336 , w_1337 , \869_b0 );
buf ( \886_A[0]_b1 , \b[0]_b1 );
buf ( \886_A[0]_b0 , \b[0]_b0 );
buf ( \887_B[0]_b1 , \c[0]_b1 );
buf ( \887_B[0]_b0 , \c[0]_b0 );
or ( \888_b1 , \886_A[0]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1338 );
and ( \888_b0 , \886_A[0]_b0 , w_1339 );
and ( w_1338 , w_1339 , \887_B[0]_b0 );
buf ( \889_Z[0]_b1 , \888_b1 );
buf ( \889_Z[0]_b0 , \888_b0 );
or ( \890_b1 , \889_Z[0]_b1 , \867_b1 );
not ( \867_b1 , w_1340 );
and ( \890_b0 , \889_Z[0]_b0 , w_1341 );
and ( w_1340 , w_1341 , \867_b0 );
buf ( \891_A[0]_b1 , \a[0]_b1 );
buf ( \891_A[0]_b0 , \a[0]_b0 );
buf ( \892_B[0]_b1 , \d[0]_b1 );
buf ( \892_B[0]_b0 , \d[0]_b0 );
or ( \893_b1 , \891_A[0]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1342 );
and ( \893_b0 , \891_A[0]_b0 , w_1343 );
and ( w_1342 , w_1343 , \892_B[0]_b0 );
buf ( \894_Z[0]_b1 , \893_b1 );
buf ( \894_Z[0]_b0 , \893_b0 );
or ( \895_b1 , \894_Z[0]_b1 , \865_b1 );
not ( \865_b1 , w_1344 );
and ( \895_b0 , \894_Z[0]_b0 , w_1345 );
and ( w_1344 , w_1345 , \865_b0 );
buf ( \896_A[0]_b1 , \b[0]_b1 );
buf ( \896_A[0]_b0 , \b[0]_b0 );
buf ( \897_B[0]_b1 , \d[0]_b1 );
buf ( \897_B[0]_b0 , \d[0]_b0 );
or ( \898_b1 , \896_A[0]_b1 , \897_B[0]_b1 );
xor ( \898_b0 , \896_A[0]_b0 , w_1346 );
not ( w_1346 , w_1347 );
and ( w_1347 , \897_B[0]_b1 , \897_B[0]_b0 );
buf ( \899_SUM[0]_b1 , \898_b1 );
buf ( \899_SUM[0]_b0 , \898_b0 );
or ( \900_b1 , \899_SUM[0]_b1 , \863_b1 );
not ( \863_b1 , w_1348 );
and ( \900_b0 , \899_SUM[0]_b0 , w_1349 );
and ( w_1348 , w_1349 , \863_b0 );
buf ( \901_A[0]_b1 , \a[0]_b1 );
buf ( \901_A[0]_b0 , \a[0]_b0 );
buf ( \902_B[0]_b1 , \c[0]_b1 );
buf ( \902_B[0]_b0 , \c[0]_b0 );
or ( \903_b1 , \901_A[0]_b1 , \902_B[0]_b1 );
xor ( \903_b0 , \901_A[0]_b0 , w_1350 );
not ( w_1350 , w_1351 );
and ( w_1351 , \902_B[0]_b1 , \902_B[0]_b0 );
buf ( \904_SUM[0]_b1 , \903_b1 );
buf ( \904_SUM[0]_b0 , \903_b0 );
or ( \905_b1 , \904_SUM[0]_b1 , \861_b1 );
not ( \861_b1 , w_1352 );
and ( \905_b0 , \904_SUM[0]_b0 , w_1353 );
and ( w_1352 , w_1353 , \861_b0 );
or ( \906_b1 , \d[0]_b1 , \859_b1 );
not ( \859_b1 , w_1354 );
and ( \906_b0 , \d[0]_b0 , w_1355 );
and ( w_1354 , w_1355 , \859_b0 );
or ( \907_b1 , \c[0]_b1 , \857_b1 );
not ( \857_b1 , w_1356 );
and ( \907_b0 , \c[0]_b0 , w_1357 );
and ( w_1356 , w_1357 , \857_b0 );
or ( \908_b1 , \b[0]_b1 , \855_b1 );
not ( \855_b1 , w_1358 );
and ( \908_b0 , \b[0]_b0 , w_1359 );
and ( w_1358 , w_1359 , \855_b0 );
or ( \909_b1 , \a[0]_b1 , \853_b1 );
not ( \853_b1 , w_1360 );
and ( \909_b0 , \a[0]_b0 , w_1361 );
and ( w_1360 , w_1361 , \853_b0 );
and ( \911_b1 , 1'b0_b1 , w_1362 );
xor ( w_1362 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1363 );
and ( \911_b0 , w_1363 , \876_b0 );
or ( \912_b1 , \a[1]_b1 , w_1364 );
or ( \912_b0 , \a[1]_b0 , \d[1]_b0 );
not ( \d[1]_b0 , w_1365 );
and ( w_1365 , w_1364 , \d[1]_b1 );
or ( \913_b1 , \912_b1 , \875_b1 );
not ( \875_b1 , w_1366 );
and ( \913_b0 , \912_b0 , w_1367 );
and ( w_1366 , w_1367 , \875_b0 );
or ( \914_b1 , \b[1]_b1 , \c[1]_b1 );
not ( \c[1]_b1 , w_1368 );
and ( \914_b0 , \b[1]_b0 , w_1369 );
and ( w_1368 , w_1369 , \c[1]_b0 );
or ( \915_b1 , \914_b1 , \873_b1 );
not ( \873_b1 , w_1370 );
and ( \915_b0 , \914_b0 , w_1371 );
and ( w_1370 , w_1371 , \873_b0 );
or ( \916_b1 , \a[1]_b1 , w_1372 );
or ( \916_b0 , \a[1]_b0 , \b[1]_b0 );
not ( \b[1]_b0 , w_1373 );
and ( w_1373 , w_1372 , \b[1]_b1 );
or ( \917_b1 , \916_b1 , \871_b1 );
not ( \871_b1 , w_1374 );
and ( \917_b0 , \916_b0 , w_1375 );
and ( w_1374 , w_1375 , \871_b0 );
or ( \918_b1 , \c[1]_b1 , \d[1]_b1 );
xor ( \918_b0 , \c[1]_b0 , w_1376 );
not ( w_1376 , w_1377 );
and ( w_1377 , \d[1]_b1 , \d[1]_b0 );
or ( \919_b1 , \918_b1 , \869_b1 );
not ( \869_b1 , w_1378 );
and ( \919_b0 , \918_b0 , w_1379 );
and ( w_1378 , w_1379 , \869_b0 );
buf ( \920_A[1]_b1 , \b[1]_b1 );
buf ( \920_A[1]_b0 , \b[1]_b0 );
or ( \921_b1 , \920_A[1]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1380 );
and ( \921_b0 , \920_A[1]_b0 , w_1381 );
and ( w_1380 , w_1381 , \887_B[0]_b0 );
buf ( \922_B[1]_b1 , \c[1]_b1 );
buf ( \922_B[1]_b0 , \c[1]_b0 );
or ( \923_b1 , \886_A[0]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_1382 );
and ( \923_b0 , \886_A[0]_b0 , w_1383 );
and ( w_1382 , w_1383 , \922_B[1]_b0 );
or ( \924_b1 , \921_b1 , \923_b1 );
xor ( \924_b0 , \921_b0 , w_1384 );
not ( w_1384 , w_1385 );
and ( w_1385 , \923_b1 , \923_b0 );
buf ( \925_Z[1]_b1 , \924_b1 );
buf ( \925_Z[1]_b0 , \924_b0 );
or ( \926_b1 , \925_Z[1]_b1 , \867_b1 );
not ( \867_b1 , w_1386 );
and ( \926_b0 , \925_Z[1]_b0 , w_1387 );
and ( w_1386 , w_1387 , \867_b0 );
buf ( \927_A[1]_b1 , \a[1]_b1 );
buf ( \927_A[1]_b0 , \a[1]_b0 );
or ( \928_b1 , \927_A[1]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1388 );
and ( \928_b0 , \927_A[1]_b0 , w_1389 );
and ( w_1388 , w_1389 , \892_B[0]_b0 );
buf ( \929_B[1]_b1 , \d[1]_b1 );
buf ( \929_B[1]_b0 , \d[1]_b0 );
or ( \930_b1 , \891_A[0]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_1390 );
and ( \930_b0 , \891_A[0]_b0 , w_1391 );
and ( w_1390 , w_1391 , \929_B[1]_b0 );
or ( \931_b1 , \928_b1 , \930_b1 );
xor ( \931_b0 , \928_b0 , w_1392 );
not ( w_1392 , w_1393 );
and ( w_1393 , \930_b1 , \930_b0 );
buf ( \932_Z[1]_b1 , \931_b1 );
buf ( \932_Z[1]_b0 , \931_b0 );
or ( \933_b1 , \932_Z[1]_b1 , \865_b1 );
not ( \865_b1 , w_1394 );
and ( \933_b0 , \932_Z[1]_b0 , w_1395 );
and ( w_1394 , w_1395 , \865_b0 );
buf ( \934_A[1]_b1 , \b[1]_b1 );
buf ( \934_A[1]_b0 , \b[1]_b0 );
buf ( \935_B[1]_b1 , \d[1]_b1 );
buf ( \935_B[1]_b0 , \d[1]_b0 );
or ( \936_b1 , \934_A[1]_b1 , \935_B[1]_b1 );
xor ( \936_b0 , \934_A[1]_b0 , w_1396 );
not ( w_1396 , w_1397 );
and ( w_1397 , \935_B[1]_b1 , \935_B[1]_b0 );
or ( \937_b1 , \896_A[0]_b1 , \897_B[0]_b1 );
not ( \897_B[0]_b1 , w_1398 );
and ( \937_b0 , \896_A[0]_b0 , w_1399 );
and ( w_1398 , w_1399 , \897_B[0]_b0 );
or ( \938_b1 , \936_b1 , \937_b1 );
xor ( \938_b0 , \936_b0 , w_1400 );
not ( w_1400 , w_1401 );
and ( w_1401 , \937_b1 , \937_b0 );
buf ( \939_SUM[1]_b1 , \938_b1 );
buf ( \939_SUM[1]_b0 , \938_b0 );
or ( \940_b1 , \939_SUM[1]_b1 , \863_b1 );
not ( \863_b1 , w_1402 );
and ( \940_b0 , \939_SUM[1]_b0 , w_1403 );
and ( w_1402 , w_1403 , \863_b0 );
buf ( \941_A[1]_b1 , \a[1]_b1 );
buf ( \941_A[1]_b0 , \a[1]_b0 );
buf ( \942_B[1]_b1 , \c[1]_b1 );
buf ( \942_B[1]_b0 , \c[1]_b0 );
or ( \943_b1 , \941_A[1]_b1 , \942_B[1]_b1 );
xor ( \943_b0 , \941_A[1]_b0 , w_1404 );
not ( w_1404 , w_1405 );
and ( w_1405 , \942_B[1]_b1 , \942_B[1]_b0 );
or ( \944_b1 , \901_A[0]_b1 , \902_B[0]_b1 );
not ( \902_B[0]_b1 , w_1406 );
and ( \944_b0 , \901_A[0]_b0 , w_1407 );
and ( w_1406 , w_1407 , \902_B[0]_b0 );
or ( \945_b1 , \943_b1 , \944_b1 );
xor ( \945_b0 , \943_b0 , w_1408 );
not ( w_1408 , w_1409 );
and ( w_1409 , \944_b1 , \944_b0 );
buf ( \946_SUM[1]_b1 , \945_b1 );
buf ( \946_SUM[1]_b0 , \945_b0 );
or ( \947_b1 , \946_SUM[1]_b1 , \861_b1 );
not ( \861_b1 , w_1410 );
and ( \947_b0 , \946_SUM[1]_b0 , w_1411 );
and ( w_1410 , w_1411 , \861_b0 );
or ( \948_b1 , \d[1]_b1 , \859_b1 );
not ( \859_b1 , w_1412 );
and ( \948_b0 , \d[1]_b0 , w_1413 );
and ( w_1412 , w_1413 , \859_b0 );
or ( \949_b1 , \c[1]_b1 , \857_b1 );
not ( \857_b1 , w_1414 );
and ( \949_b0 , \c[1]_b0 , w_1415 );
and ( w_1414 , w_1415 , \857_b0 );
or ( \950_b1 , \b[1]_b1 , \855_b1 );
not ( \855_b1 , w_1416 );
and ( \950_b0 , \b[1]_b0 , w_1417 );
and ( w_1416 , w_1417 , \855_b0 );
or ( \951_b1 , \a[1]_b1 , \853_b1 );
not ( \853_b1 , w_1418 );
and ( \951_b0 , \a[1]_b0 , w_1419 );
and ( w_1418 , w_1419 , \853_b0 );
and ( \953_b1 , 1'b0_b1 , w_1420 );
xor ( w_1420 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1421 );
and ( \953_b0 , w_1421 , \876_b0 );
or ( \954_b1 , \a[2]_b1 , w_1422 );
or ( \954_b0 , \a[2]_b0 , \d[2]_b0 );
not ( \d[2]_b0 , w_1423 );
and ( w_1423 , w_1422 , \d[2]_b1 );
or ( \955_b1 , \954_b1 , \875_b1 );
not ( \875_b1 , w_1424 );
and ( \955_b0 , \954_b0 , w_1425 );
and ( w_1424 , w_1425 , \875_b0 );
or ( \956_b1 , \b[2]_b1 , \c[2]_b1 );
not ( \c[2]_b1 , w_1426 );
and ( \956_b0 , \b[2]_b0 , w_1427 );
and ( w_1426 , w_1427 , \c[2]_b0 );
or ( \957_b1 , \956_b1 , \873_b1 );
not ( \873_b1 , w_1428 );
and ( \957_b0 , \956_b0 , w_1429 );
and ( w_1428 , w_1429 , \873_b0 );
or ( \958_b1 , \a[2]_b1 , w_1430 );
or ( \958_b0 , \a[2]_b0 , \b[2]_b0 );
not ( \b[2]_b0 , w_1431 );
and ( w_1431 , w_1430 , \b[2]_b1 );
or ( \959_b1 , \958_b1 , \871_b1 );
not ( \871_b1 , w_1432 );
and ( \959_b0 , \958_b0 , w_1433 );
and ( w_1432 , w_1433 , \871_b0 );
or ( \960_b1 , \c[2]_b1 , \d[2]_b1 );
xor ( \960_b0 , \c[2]_b0 , w_1434 );
not ( w_1434 , w_1435 );
and ( w_1435 , \d[2]_b1 , \d[2]_b0 );
or ( \961_b1 , \960_b1 , \869_b1 );
not ( \869_b1 , w_1436 );
and ( \961_b0 , \960_b0 , w_1437 );
and ( w_1436 , w_1437 , \869_b0 );
buf ( \962_A[2]_b1 , \b[2]_b1 );
buf ( \962_A[2]_b0 , \b[2]_b0 );
or ( \963_b1 , \962_A[2]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1438 );
and ( \963_b0 , \962_A[2]_b0 , w_1439 );
and ( w_1438 , w_1439 , \887_B[0]_b0 );
or ( \964_b1 , \920_A[1]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_1440 );
and ( \964_b0 , \920_A[1]_b0 , w_1441 );
and ( w_1440 , w_1441 , \922_B[1]_b0 );
or ( \965_b1 , \963_b1 , \964_b1 );
xor ( \965_b0 , \963_b0 , w_1442 );
not ( w_1442 , w_1443 );
and ( w_1443 , \964_b1 , \964_b0 );
or ( \966_b1 , \921_b1 , \923_b1 );
not ( \923_b1 , w_1444 );
and ( \966_b0 , \921_b0 , w_1445 );
and ( w_1444 , w_1445 , \923_b0 );
or ( \967_b1 , \965_b1 , \966_b1 );
xor ( \967_b0 , \965_b0 , w_1446 );
not ( w_1446 , w_1447 );
and ( w_1447 , \966_b1 , \966_b0 );
buf ( \968_B[2]_b1 , \c[2]_b1 );
buf ( \968_B[2]_b0 , \c[2]_b0 );
or ( \969_b1 , \886_A[0]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_1448 );
and ( \969_b0 , \886_A[0]_b0 , w_1449 );
and ( w_1448 , w_1449 , \968_B[2]_b0 );
or ( \970_b1 , \967_b1 , \969_b1 );
xor ( \970_b0 , \967_b0 , w_1450 );
not ( w_1450 , w_1451 );
and ( w_1451 , \969_b1 , \969_b0 );
buf ( \971_Z[2]_b1 , \970_b1 );
buf ( \971_Z[2]_b0 , \970_b0 );
or ( \972_b1 , \971_Z[2]_b1 , \867_b1 );
not ( \867_b1 , w_1452 );
and ( \972_b0 , \971_Z[2]_b0 , w_1453 );
and ( w_1452 , w_1453 , \867_b0 );
buf ( \973_A[2]_b1 , \a[2]_b1 );
buf ( \973_A[2]_b0 , \a[2]_b0 );
or ( \974_b1 , \973_A[2]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1454 );
and ( \974_b0 , \973_A[2]_b0 , w_1455 );
and ( w_1454 , w_1455 , \892_B[0]_b0 );
or ( \975_b1 , \927_A[1]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_1456 );
and ( \975_b0 , \927_A[1]_b0 , w_1457 );
and ( w_1456 , w_1457 , \929_B[1]_b0 );
or ( \976_b1 , \974_b1 , \975_b1 );
xor ( \976_b0 , \974_b0 , w_1458 );
not ( w_1458 , w_1459 );
and ( w_1459 , \975_b1 , \975_b0 );
or ( \977_b1 , \928_b1 , \930_b1 );
not ( \930_b1 , w_1460 );
and ( \977_b0 , \928_b0 , w_1461 );
and ( w_1460 , w_1461 , \930_b0 );
or ( \978_b1 , \976_b1 , \977_b1 );
xor ( \978_b0 , \976_b0 , w_1462 );
not ( w_1462 , w_1463 );
and ( w_1463 , \977_b1 , \977_b0 );
buf ( \979_B[2]_b1 , \d[2]_b1 );
buf ( \979_B[2]_b0 , \d[2]_b0 );
or ( \980_b1 , \891_A[0]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_1464 );
and ( \980_b0 , \891_A[0]_b0 , w_1465 );
and ( w_1464 , w_1465 , \979_B[2]_b0 );
or ( \981_b1 , \978_b1 , \980_b1 );
xor ( \981_b0 , \978_b0 , w_1466 );
not ( w_1466 , w_1467 );
and ( w_1467 , \980_b1 , \980_b0 );
buf ( \982_Z[2]_b1 , \981_b1 );
buf ( \982_Z[2]_b0 , \981_b0 );
or ( \983_b1 , \982_Z[2]_b1 , \865_b1 );
not ( \865_b1 , w_1468 );
and ( \983_b0 , \982_Z[2]_b0 , w_1469 );
and ( w_1468 , w_1469 , \865_b0 );
buf ( \984_A[2]_b1 , \b[2]_b1 );
buf ( \984_A[2]_b0 , \b[2]_b0 );
buf ( \985_B[2]_b1 , \d[2]_b1 );
buf ( \985_B[2]_b0 , \d[2]_b0 );
or ( \986_b1 , \984_A[2]_b1 , \985_B[2]_b1 );
xor ( \986_b0 , \984_A[2]_b0 , w_1470 );
not ( w_1470 , w_1471 );
and ( w_1471 , \985_B[2]_b1 , \985_B[2]_b0 );
or ( \987_b1 , \934_A[1]_b1 , \935_B[1]_b1 );
not ( \935_B[1]_b1 , w_1472 );
and ( \987_b0 , \934_A[1]_b0 , w_1473 );
and ( w_1472 , w_1473 , \935_B[1]_b0 );
or ( \988_b1 , \935_B[1]_b1 , \937_b1 );
not ( \937_b1 , w_1474 );
and ( \988_b0 , \935_B[1]_b0 , w_1475 );
and ( w_1474 , w_1475 , \937_b0 );
or ( \989_b1 , \934_A[1]_b1 , \937_b1 );
not ( \937_b1 , w_1476 );
and ( \989_b0 , \934_A[1]_b0 , w_1477 );
and ( w_1476 , w_1477 , \937_b0 );
or ( \991_b1 , \986_b1 , \990_b1 );
xor ( \991_b0 , \986_b0 , w_1478 );
not ( w_1478 , w_1479 );
and ( w_1479 , \990_b1 , \990_b0 );
buf ( \992_SUM[2]_b1 , \991_b1 );
buf ( \992_SUM[2]_b0 , \991_b0 );
or ( \993_b1 , \992_SUM[2]_b1 , \863_b1 );
not ( \863_b1 , w_1480 );
and ( \993_b0 , \992_SUM[2]_b0 , w_1481 );
and ( w_1480 , w_1481 , \863_b0 );
buf ( \994_A[2]_b1 , \a[2]_b1 );
buf ( \994_A[2]_b0 , \a[2]_b0 );
buf ( \995_B[2]_b1 , \c[2]_b1 );
buf ( \995_B[2]_b0 , \c[2]_b0 );
or ( \996_b1 , \994_A[2]_b1 , \995_B[2]_b1 );
xor ( \996_b0 , \994_A[2]_b0 , w_1482 );
not ( w_1482 , w_1483 );
and ( w_1483 , \995_B[2]_b1 , \995_B[2]_b0 );
or ( \997_b1 , \941_A[1]_b1 , \942_B[1]_b1 );
not ( \942_B[1]_b1 , w_1484 );
and ( \997_b0 , \941_A[1]_b0 , w_1485 );
and ( w_1484 , w_1485 , \942_B[1]_b0 );
or ( \998_b1 , \942_B[1]_b1 , \944_b1 );
not ( \944_b1 , w_1486 );
and ( \998_b0 , \942_B[1]_b0 , w_1487 );
and ( w_1486 , w_1487 , \944_b0 );
or ( \999_b1 , \941_A[1]_b1 , \944_b1 );
not ( \944_b1 , w_1488 );
and ( \999_b0 , \941_A[1]_b0 , w_1489 );
and ( w_1488 , w_1489 , \944_b0 );
or ( \1001_b1 , \996_b1 , \1000_b1 );
xor ( \1001_b0 , \996_b0 , w_1490 );
not ( w_1490 , w_1491 );
and ( w_1491 , \1000_b1 , \1000_b0 );
buf ( \1002_SUM[2]_b1 , \1001_b1 );
buf ( \1002_SUM[2]_b0 , \1001_b0 );
or ( \1003_b1 , \1002_SUM[2]_b1 , \861_b1 );
not ( \861_b1 , w_1492 );
and ( \1003_b0 , \1002_SUM[2]_b0 , w_1493 );
and ( w_1492 , w_1493 , \861_b0 );
or ( \1004_b1 , \d[2]_b1 , \859_b1 );
not ( \859_b1 , w_1494 );
and ( \1004_b0 , \d[2]_b0 , w_1495 );
and ( w_1494 , w_1495 , \859_b0 );
or ( \1005_b1 , \c[2]_b1 , \857_b1 );
not ( \857_b1 , w_1496 );
and ( \1005_b0 , \c[2]_b0 , w_1497 );
and ( w_1496 , w_1497 , \857_b0 );
or ( \1006_b1 , \b[2]_b1 , \855_b1 );
not ( \855_b1 , w_1498 );
and ( \1006_b0 , \b[2]_b0 , w_1499 );
and ( w_1498 , w_1499 , \855_b0 );
or ( \1007_b1 , \a[2]_b1 , \853_b1 );
not ( \853_b1 , w_1500 );
and ( \1007_b0 , \a[2]_b0 , w_1501 );
and ( w_1500 , w_1501 , \853_b0 );
and ( \1009_b1 , 1'b0_b1 , w_1502 );
xor ( w_1502 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1503 );
and ( \1009_b0 , w_1503 , \876_b0 );
or ( \1010_b1 , \a[3]_b1 , w_1504 );
or ( \1010_b0 , \a[3]_b0 , \d[3]_b0 );
not ( \d[3]_b0 , w_1505 );
and ( w_1505 , w_1504 , \d[3]_b1 );
or ( \1011_b1 , \1010_b1 , \875_b1 );
not ( \875_b1 , w_1506 );
and ( \1011_b0 , \1010_b0 , w_1507 );
and ( w_1506 , w_1507 , \875_b0 );
or ( \1012_b1 , \b[3]_b1 , \c[3]_b1 );
not ( \c[3]_b1 , w_1508 );
and ( \1012_b0 , \b[3]_b0 , w_1509 );
and ( w_1508 , w_1509 , \c[3]_b0 );
or ( \1013_b1 , \1012_b1 , \873_b1 );
not ( \873_b1 , w_1510 );
and ( \1013_b0 , \1012_b0 , w_1511 );
and ( w_1510 , w_1511 , \873_b0 );
or ( \1014_b1 , \a[3]_b1 , w_1512 );
or ( \1014_b0 , \a[3]_b0 , \b[3]_b0 );
not ( \b[3]_b0 , w_1513 );
and ( w_1513 , w_1512 , \b[3]_b1 );
or ( \1015_b1 , \1014_b1 , \871_b1 );
not ( \871_b1 , w_1514 );
and ( \1015_b0 , \1014_b0 , w_1515 );
and ( w_1514 , w_1515 , \871_b0 );
or ( \1016_b1 , \c[3]_b1 , \d[3]_b1 );
xor ( \1016_b0 , \c[3]_b0 , w_1516 );
not ( w_1516 , w_1517 );
and ( w_1517 , \d[3]_b1 , \d[3]_b0 );
or ( \1017_b1 , \1016_b1 , \869_b1 );
not ( \869_b1 , w_1518 );
and ( \1017_b0 , \1016_b0 , w_1519 );
and ( w_1518 , w_1519 , \869_b0 );
buf ( \1018_A[3]_b1 , \b[3]_b1 );
buf ( \1018_A[3]_b0 , \b[3]_b0 );
or ( \1019_b1 , \1018_A[3]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1520 );
and ( \1019_b0 , \1018_A[3]_b0 , w_1521 );
and ( w_1520 , w_1521 , \887_B[0]_b0 );
or ( \1020_b1 , \962_A[2]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_1522 );
and ( \1020_b0 , \962_A[2]_b0 , w_1523 );
and ( w_1522 , w_1523 , \922_B[1]_b0 );
or ( \1021_b1 , \1019_b1 , \1020_b1 );
xor ( \1021_b0 , \1019_b0 , w_1524 );
not ( w_1524 , w_1525 );
and ( w_1525 , \1020_b1 , \1020_b0 );
or ( \1022_b1 , \963_b1 , \964_b1 );
not ( \964_b1 , w_1526 );
and ( \1022_b0 , \963_b0 , w_1527 );
and ( w_1526 , w_1527 , \964_b0 );
or ( \1023_b1 , \965_b1 , \966_b1 );
not ( \966_b1 , w_1528 );
and ( \1023_b0 , \965_b0 , w_1529 );
and ( w_1528 , w_1529 , \966_b0 );
or ( \1024_b1 , \1022_b1 , w_1530 );
or ( \1024_b0 , \1022_b0 , \1023_b0 );
not ( \1023_b0 , w_1531 );
and ( w_1531 , w_1530 , \1023_b1 );
or ( \1025_b1 , \1021_b1 , \1024_b1 );
xor ( \1025_b0 , \1021_b0 , w_1532 );
not ( w_1532 , w_1533 );
and ( w_1533 , \1024_b1 , \1024_b0 );
or ( \1026_b1 , \920_A[1]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_1534 );
and ( \1026_b0 , \920_A[1]_b0 , w_1535 );
and ( w_1534 , w_1535 , \968_B[2]_b0 );
or ( \1027_b1 , \1025_b1 , \1026_b1 );
xor ( \1027_b0 , \1025_b0 , w_1536 );
not ( w_1536 , w_1537 );
and ( w_1537 , \1026_b1 , \1026_b0 );
or ( \1028_b1 , \967_b1 , \969_b1 );
not ( \969_b1 , w_1538 );
and ( \1028_b0 , \967_b0 , w_1539 );
and ( w_1538 , w_1539 , \969_b0 );
or ( \1029_b1 , \1027_b1 , \1028_b1 );
xor ( \1029_b0 , \1027_b0 , w_1540 );
not ( w_1540 , w_1541 );
and ( w_1541 , \1028_b1 , \1028_b0 );
buf ( \1030_B[3]_b1 , \c[3]_b1 );
buf ( \1030_B[3]_b0 , \c[3]_b0 );
or ( \1031_b1 , \886_A[0]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_1542 );
and ( \1031_b0 , \886_A[0]_b0 , w_1543 );
and ( w_1542 , w_1543 , \1030_B[3]_b0 );
or ( \1032_b1 , \1029_b1 , \1031_b1 );
xor ( \1032_b0 , \1029_b0 , w_1544 );
not ( w_1544 , w_1545 );
and ( w_1545 , \1031_b1 , \1031_b0 );
buf ( \1033_Z[3]_b1 , \1032_b1 );
buf ( \1033_Z[3]_b0 , \1032_b0 );
or ( \1034_b1 , \1033_Z[3]_b1 , \867_b1 );
not ( \867_b1 , w_1546 );
and ( \1034_b0 , \1033_Z[3]_b0 , w_1547 );
and ( w_1546 , w_1547 , \867_b0 );
buf ( \1035_A[3]_b1 , \a[3]_b1 );
buf ( \1035_A[3]_b0 , \a[3]_b0 );
or ( \1036_b1 , \1035_A[3]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1548 );
and ( \1036_b0 , \1035_A[3]_b0 , w_1549 );
and ( w_1548 , w_1549 , \892_B[0]_b0 );
or ( \1037_b1 , \973_A[2]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_1550 );
and ( \1037_b0 , \973_A[2]_b0 , w_1551 );
and ( w_1550 , w_1551 , \929_B[1]_b0 );
or ( \1038_b1 , \1036_b1 , \1037_b1 );
xor ( \1038_b0 , \1036_b0 , w_1552 );
not ( w_1552 , w_1553 );
and ( w_1553 , \1037_b1 , \1037_b0 );
or ( \1039_b1 , \974_b1 , \975_b1 );
not ( \975_b1 , w_1554 );
and ( \1039_b0 , \974_b0 , w_1555 );
and ( w_1554 , w_1555 , \975_b0 );
or ( \1040_b1 , \976_b1 , \977_b1 );
not ( \977_b1 , w_1556 );
and ( \1040_b0 , \976_b0 , w_1557 );
and ( w_1556 , w_1557 , \977_b0 );
or ( \1041_b1 , \1039_b1 , w_1558 );
or ( \1041_b0 , \1039_b0 , \1040_b0 );
not ( \1040_b0 , w_1559 );
and ( w_1559 , w_1558 , \1040_b1 );
or ( \1042_b1 , \1038_b1 , \1041_b1 );
xor ( \1042_b0 , \1038_b0 , w_1560 );
not ( w_1560 , w_1561 );
and ( w_1561 , \1041_b1 , \1041_b0 );
or ( \1043_b1 , \927_A[1]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_1562 );
and ( \1043_b0 , \927_A[1]_b0 , w_1563 );
and ( w_1562 , w_1563 , \979_B[2]_b0 );
or ( \1044_b1 , \1042_b1 , \1043_b1 );
xor ( \1044_b0 , \1042_b0 , w_1564 );
not ( w_1564 , w_1565 );
and ( w_1565 , \1043_b1 , \1043_b0 );
or ( \1045_b1 , \978_b1 , \980_b1 );
not ( \980_b1 , w_1566 );
and ( \1045_b0 , \978_b0 , w_1567 );
and ( w_1566 , w_1567 , \980_b0 );
or ( \1046_b1 , \1044_b1 , \1045_b1 );
xor ( \1046_b0 , \1044_b0 , w_1568 );
not ( w_1568 , w_1569 );
and ( w_1569 , \1045_b1 , \1045_b0 );
buf ( \1047_B[3]_b1 , \d[3]_b1 );
buf ( \1047_B[3]_b0 , \d[3]_b0 );
or ( \1048_b1 , \891_A[0]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_1570 );
and ( \1048_b0 , \891_A[0]_b0 , w_1571 );
and ( w_1570 , w_1571 , \1047_B[3]_b0 );
or ( \1049_b1 , \1046_b1 , \1048_b1 );
xor ( \1049_b0 , \1046_b0 , w_1572 );
not ( w_1572 , w_1573 );
and ( w_1573 , \1048_b1 , \1048_b0 );
buf ( \1050_Z[3]_b1 , \1049_b1 );
buf ( \1050_Z[3]_b0 , \1049_b0 );
or ( \1051_b1 , \1050_Z[3]_b1 , \865_b1 );
not ( \865_b1 , w_1574 );
and ( \1051_b0 , \1050_Z[3]_b0 , w_1575 );
and ( w_1574 , w_1575 , \865_b0 );
buf ( \1052_A[3]_b1 , \b[3]_b1 );
buf ( \1052_A[3]_b0 , \b[3]_b0 );
buf ( \1053_B[3]_b1 , \d[3]_b1 );
buf ( \1053_B[3]_b0 , \d[3]_b0 );
or ( \1054_b1 , \1052_A[3]_b1 , \1053_B[3]_b1 );
xor ( \1054_b0 , \1052_A[3]_b0 , w_1576 );
not ( w_1576 , w_1577 );
and ( w_1577 , \1053_B[3]_b1 , \1053_B[3]_b0 );
or ( \1055_b1 , \984_A[2]_b1 , \985_B[2]_b1 );
not ( \985_B[2]_b1 , w_1578 );
and ( \1055_b0 , \984_A[2]_b0 , w_1579 );
and ( w_1578 , w_1579 , \985_B[2]_b0 );
or ( \1056_b1 , \985_B[2]_b1 , \990_b1 );
not ( \990_b1 , w_1580 );
and ( \1056_b0 , \985_B[2]_b0 , w_1581 );
and ( w_1580 , w_1581 , \990_b0 );
or ( \1057_b1 , \984_A[2]_b1 , \990_b1 );
not ( \990_b1 , w_1582 );
and ( \1057_b0 , \984_A[2]_b0 , w_1583 );
and ( w_1582 , w_1583 , \990_b0 );
or ( \1059_b1 , \1054_b1 , \1058_b1 );
xor ( \1059_b0 , \1054_b0 , w_1584 );
not ( w_1584 , w_1585 );
and ( w_1585 , \1058_b1 , \1058_b0 );
buf ( \1060_SUM[3]_b1 , \1059_b1 );
buf ( \1060_SUM[3]_b0 , \1059_b0 );
or ( \1061_b1 , \1060_SUM[3]_b1 , \863_b1 );
not ( \863_b1 , w_1586 );
and ( \1061_b0 , \1060_SUM[3]_b0 , w_1587 );
and ( w_1586 , w_1587 , \863_b0 );
buf ( \1062_A[3]_b1 , \a[3]_b1 );
buf ( \1062_A[3]_b0 , \a[3]_b0 );
buf ( \1063_B[3]_b1 , \c[3]_b1 );
buf ( \1063_B[3]_b0 , \c[3]_b0 );
or ( \1064_b1 , \1062_A[3]_b1 , \1063_B[3]_b1 );
xor ( \1064_b0 , \1062_A[3]_b0 , w_1588 );
not ( w_1588 , w_1589 );
and ( w_1589 , \1063_B[3]_b1 , \1063_B[3]_b0 );
or ( \1065_b1 , \994_A[2]_b1 , \995_B[2]_b1 );
not ( \995_B[2]_b1 , w_1590 );
and ( \1065_b0 , \994_A[2]_b0 , w_1591 );
and ( w_1590 , w_1591 , \995_B[2]_b0 );
or ( \1066_b1 , \995_B[2]_b1 , \1000_b1 );
not ( \1000_b1 , w_1592 );
and ( \1066_b0 , \995_B[2]_b0 , w_1593 );
and ( w_1592 , w_1593 , \1000_b0 );
or ( \1067_b1 , \994_A[2]_b1 , \1000_b1 );
not ( \1000_b1 , w_1594 );
and ( \1067_b0 , \994_A[2]_b0 , w_1595 );
and ( w_1594 , w_1595 , \1000_b0 );
or ( \1069_b1 , \1064_b1 , \1068_b1 );
xor ( \1069_b0 , \1064_b0 , w_1596 );
not ( w_1596 , w_1597 );
and ( w_1597 , \1068_b1 , \1068_b0 );
buf ( \1070_SUM[3]_b1 , \1069_b1 );
buf ( \1070_SUM[3]_b0 , \1069_b0 );
or ( \1071_b1 , \1070_SUM[3]_b1 , \861_b1 );
not ( \861_b1 , w_1598 );
and ( \1071_b0 , \1070_SUM[3]_b0 , w_1599 );
and ( w_1598 , w_1599 , \861_b0 );
or ( \1072_b1 , \d[3]_b1 , \859_b1 );
not ( \859_b1 , w_1600 );
and ( \1072_b0 , \d[3]_b0 , w_1601 );
and ( w_1600 , w_1601 , \859_b0 );
or ( \1073_b1 , \c[3]_b1 , \857_b1 );
not ( \857_b1 , w_1602 );
and ( \1073_b0 , \c[3]_b0 , w_1603 );
and ( w_1602 , w_1603 , \857_b0 );
or ( \1074_b1 , \b[3]_b1 , \855_b1 );
not ( \855_b1 , w_1604 );
and ( \1074_b0 , \b[3]_b0 , w_1605 );
and ( w_1604 , w_1605 , \855_b0 );
or ( \1075_b1 , \a[3]_b1 , \853_b1 );
not ( \853_b1 , w_1606 );
and ( \1075_b0 , \a[3]_b0 , w_1607 );
and ( w_1606 , w_1607 , \853_b0 );
and ( \1077_b1 , 1'b0_b1 , w_1608 );
xor ( w_1608 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1609 );
and ( \1077_b0 , w_1609 , \876_b0 );
or ( \1078_b1 , \a[4]_b1 , w_1610 );
or ( \1078_b0 , \a[4]_b0 , \d[4]_b0 );
not ( \d[4]_b0 , w_1611 );
and ( w_1611 , w_1610 , \d[4]_b1 );
or ( \1079_b1 , \1078_b1 , \875_b1 );
not ( \875_b1 , w_1612 );
and ( \1079_b0 , \1078_b0 , w_1613 );
and ( w_1612 , w_1613 , \875_b0 );
or ( \1080_b1 , \b[4]_b1 , \c[4]_b1 );
not ( \c[4]_b1 , w_1614 );
and ( \1080_b0 , \b[4]_b0 , w_1615 );
and ( w_1614 , w_1615 , \c[4]_b0 );
or ( \1081_b1 , \1080_b1 , \873_b1 );
not ( \873_b1 , w_1616 );
and ( \1081_b0 , \1080_b0 , w_1617 );
and ( w_1616 , w_1617 , \873_b0 );
or ( \1082_b1 , \a[4]_b1 , w_1618 );
or ( \1082_b0 , \a[4]_b0 , \b[4]_b0 );
not ( \b[4]_b0 , w_1619 );
and ( w_1619 , w_1618 , \b[4]_b1 );
or ( \1083_b1 , \1082_b1 , \871_b1 );
not ( \871_b1 , w_1620 );
and ( \1083_b0 , \1082_b0 , w_1621 );
and ( w_1620 , w_1621 , \871_b0 );
or ( \1084_b1 , \c[4]_b1 , \d[4]_b1 );
xor ( \1084_b0 , \c[4]_b0 , w_1622 );
not ( w_1622 , w_1623 );
and ( w_1623 , \d[4]_b1 , \d[4]_b0 );
or ( \1085_b1 , \1084_b1 , \869_b1 );
not ( \869_b1 , w_1624 );
and ( \1085_b0 , \1084_b0 , w_1625 );
and ( w_1624 , w_1625 , \869_b0 );
buf ( \1086_A[4]_b1 , \b[4]_b1 );
buf ( \1086_A[4]_b0 , \b[4]_b0 );
or ( \1087_b1 , \1086_A[4]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1626 );
and ( \1087_b0 , \1086_A[4]_b0 , w_1627 );
and ( w_1626 , w_1627 , \887_B[0]_b0 );
or ( \1088_b1 , \1018_A[3]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_1628 );
and ( \1088_b0 , \1018_A[3]_b0 , w_1629 );
and ( w_1628 , w_1629 , \922_B[1]_b0 );
or ( \1089_b1 , \1087_b1 , \1088_b1 );
xor ( \1089_b0 , \1087_b0 , w_1630 );
not ( w_1630 , w_1631 );
and ( w_1631 , \1088_b1 , \1088_b0 );
or ( \1090_b1 , \1019_b1 , \1020_b1 );
not ( \1020_b1 , w_1632 );
and ( \1090_b0 , \1019_b0 , w_1633 );
and ( w_1632 , w_1633 , \1020_b0 );
or ( \1091_b1 , \1021_b1 , \1024_b1 );
not ( \1024_b1 , w_1634 );
and ( \1091_b0 , \1021_b0 , w_1635 );
and ( w_1634 , w_1635 , \1024_b0 );
or ( \1092_b1 , \1090_b1 , w_1636 );
or ( \1092_b0 , \1090_b0 , \1091_b0 );
not ( \1091_b0 , w_1637 );
and ( w_1637 , w_1636 , \1091_b1 );
or ( \1093_b1 , \1089_b1 , \1092_b1 );
xor ( \1093_b0 , \1089_b0 , w_1638 );
not ( w_1638 , w_1639 );
and ( w_1639 , \1092_b1 , \1092_b0 );
or ( \1094_b1 , \962_A[2]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_1640 );
and ( \1094_b0 , \962_A[2]_b0 , w_1641 );
and ( w_1640 , w_1641 , \968_B[2]_b0 );
or ( \1095_b1 , \1093_b1 , \1094_b1 );
xor ( \1095_b0 , \1093_b0 , w_1642 );
not ( w_1642 , w_1643 );
and ( w_1643 , \1094_b1 , \1094_b0 );
or ( \1096_b1 , \1025_b1 , \1026_b1 );
not ( \1026_b1 , w_1644 );
and ( \1096_b0 , \1025_b0 , w_1645 );
and ( w_1644 , w_1645 , \1026_b0 );
or ( \1097_b1 , \1027_b1 , \1028_b1 );
not ( \1028_b1 , w_1646 );
and ( \1097_b0 , \1027_b0 , w_1647 );
and ( w_1646 , w_1647 , \1028_b0 );
or ( \1098_b1 , \1096_b1 , w_1648 );
or ( \1098_b0 , \1096_b0 , \1097_b0 );
not ( \1097_b0 , w_1649 );
and ( w_1649 , w_1648 , \1097_b1 );
or ( \1099_b1 , \1095_b1 , \1098_b1 );
xor ( \1099_b0 , \1095_b0 , w_1650 );
not ( w_1650 , w_1651 );
and ( w_1651 , \1098_b1 , \1098_b0 );
or ( \1100_b1 , \920_A[1]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_1652 );
and ( \1100_b0 , \920_A[1]_b0 , w_1653 );
and ( w_1652 , w_1653 , \1030_B[3]_b0 );
or ( \1101_b1 , \1099_b1 , \1100_b1 );
xor ( \1101_b0 , \1099_b0 , w_1654 );
not ( w_1654 , w_1655 );
and ( w_1655 , \1100_b1 , \1100_b0 );
or ( \1102_b1 , \1029_b1 , \1031_b1 );
not ( \1031_b1 , w_1656 );
and ( \1102_b0 , \1029_b0 , w_1657 );
and ( w_1656 , w_1657 , \1031_b0 );
or ( \1103_b1 , \1101_b1 , \1102_b1 );
xor ( \1103_b0 , \1101_b0 , w_1658 );
not ( w_1658 , w_1659 );
and ( w_1659 , \1102_b1 , \1102_b0 );
buf ( \1104_B[4]_b1 , \c[4]_b1 );
buf ( \1104_B[4]_b0 , \c[4]_b0 );
or ( \1105_b1 , \886_A[0]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_1660 );
and ( \1105_b0 , \886_A[0]_b0 , w_1661 );
and ( w_1660 , w_1661 , \1104_B[4]_b0 );
or ( \1106_b1 , \1103_b1 , \1105_b1 );
xor ( \1106_b0 , \1103_b0 , w_1662 );
not ( w_1662 , w_1663 );
and ( w_1663 , \1105_b1 , \1105_b0 );
buf ( \1107_Z[4]_b1 , \1106_b1 );
buf ( \1107_Z[4]_b0 , \1106_b0 );
or ( \1108_b1 , \1107_Z[4]_b1 , \867_b1 );
not ( \867_b1 , w_1664 );
and ( \1108_b0 , \1107_Z[4]_b0 , w_1665 );
and ( w_1664 , w_1665 , \867_b0 );
buf ( \1109_A[4]_b1 , \a[4]_b1 );
buf ( \1109_A[4]_b0 , \a[4]_b0 );
or ( \1110_b1 , \1109_A[4]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1666 );
and ( \1110_b0 , \1109_A[4]_b0 , w_1667 );
and ( w_1666 , w_1667 , \892_B[0]_b0 );
or ( \1111_b1 , \1035_A[3]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_1668 );
and ( \1111_b0 , \1035_A[3]_b0 , w_1669 );
and ( w_1668 , w_1669 , \929_B[1]_b0 );
or ( \1112_b1 , \1110_b1 , \1111_b1 );
xor ( \1112_b0 , \1110_b0 , w_1670 );
not ( w_1670 , w_1671 );
and ( w_1671 , \1111_b1 , \1111_b0 );
or ( \1113_b1 , \1036_b1 , \1037_b1 );
not ( \1037_b1 , w_1672 );
and ( \1113_b0 , \1036_b0 , w_1673 );
and ( w_1672 , w_1673 , \1037_b0 );
or ( \1114_b1 , \1038_b1 , \1041_b1 );
not ( \1041_b1 , w_1674 );
and ( \1114_b0 , \1038_b0 , w_1675 );
and ( w_1674 , w_1675 , \1041_b0 );
or ( \1115_b1 , \1113_b1 , w_1676 );
or ( \1115_b0 , \1113_b0 , \1114_b0 );
not ( \1114_b0 , w_1677 );
and ( w_1677 , w_1676 , \1114_b1 );
or ( \1116_b1 , \1112_b1 , \1115_b1 );
xor ( \1116_b0 , \1112_b0 , w_1678 );
not ( w_1678 , w_1679 );
and ( w_1679 , \1115_b1 , \1115_b0 );
or ( \1117_b1 , \973_A[2]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_1680 );
and ( \1117_b0 , \973_A[2]_b0 , w_1681 );
and ( w_1680 , w_1681 , \979_B[2]_b0 );
or ( \1118_b1 , \1116_b1 , \1117_b1 );
xor ( \1118_b0 , \1116_b0 , w_1682 );
not ( w_1682 , w_1683 );
and ( w_1683 , \1117_b1 , \1117_b0 );
or ( \1119_b1 , \1042_b1 , \1043_b1 );
not ( \1043_b1 , w_1684 );
and ( \1119_b0 , \1042_b0 , w_1685 );
and ( w_1684 , w_1685 , \1043_b0 );
or ( \1120_b1 , \1044_b1 , \1045_b1 );
not ( \1045_b1 , w_1686 );
and ( \1120_b0 , \1044_b0 , w_1687 );
and ( w_1686 , w_1687 , \1045_b0 );
or ( \1121_b1 , \1119_b1 , w_1688 );
or ( \1121_b0 , \1119_b0 , \1120_b0 );
not ( \1120_b0 , w_1689 );
and ( w_1689 , w_1688 , \1120_b1 );
or ( \1122_b1 , \1118_b1 , \1121_b1 );
xor ( \1122_b0 , \1118_b0 , w_1690 );
not ( w_1690 , w_1691 );
and ( w_1691 , \1121_b1 , \1121_b0 );
or ( \1123_b1 , \927_A[1]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_1692 );
and ( \1123_b0 , \927_A[1]_b0 , w_1693 );
and ( w_1692 , w_1693 , \1047_B[3]_b0 );
or ( \1124_b1 , \1122_b1 , \1123_b1 );
xor ( \1124_b0 , \1122_b0 , w_1694 );
not ( w_1694 , w_1695 );
and ( w_1695 , \1123_b1 , \1123_b0 );
or ( \1125_b1 , \1046_b1 , \1048_b1 );
not ( \1048_b1 , w_1696 );
and ( \1125_b0 , \1046_b0 , w_1697 );
and ( w_1696 , w_1697 , \1048_b0 );
or ( \1126_b1 , \1124_b1 , \1125_b1 );
xor ( \1126_b0 , \1124_b0 , w_1698 );
not ( w_1698 , w_1699 );
and ( w_1699 , \1125_b1 , \1125_b0 );
buf ( \1127_B[4]_b1 , \d[4]_b1 );
buf ( \1127_B[4]_b0 , \d[4]_b0 );
or ( \1128_b1 , \891_A[0]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_1700 );
and ( \1128_b0 , \891_A[0]_b0 , w_1701 );
and ( w_1700 , w_1701 , \1127_B[4]_b0 );
or ( \1129_b1 , \1126_b1 , \1128_b1 );
xor ( \1129_b0 , \1126_b0 , w_1702 );
not ( w_1702 , w_1703 );
and ( w_1703 , \1128_b1 , \1128_b0 );
buf ( \1130_Z[4]_b1 , \1129_b1 );
buf ( \1130_Z[4]_b0 , \1129_b0 );
or ( \1131_b1 , \1130_Z[4]_b1 , \865_b1 );
not ( \865_b1 , w_1704 );
and ( \1131_b0 , \1130_Z[4]_b0 , w_1705 );
and ( w_1704 , w_1705 , \865_b0 );
buf ( \1132_A[4]_b1 , \b[4]_b1 );
buf ( \1132_A[4]_b0 , \b[4]_b0 );
buf ( \1133_B[4]_b1 , \d[4]_b1 );
buf ( \1133_B[4]_b0 , \d[4]_b0 );
or ( \1134_b1 , \1132_A[4]_b1 , \1133_B[4]_b1 );
xor ( \1134_b0 , \1132_A[4]_b0 , w_1706 );
not ( w_1706 , w_1707 );
and ( w_1707 , \1133_B[4]_b1 , \1133_B[4]_b0 );
or ( \1135_b1 , \1052_A[3]_b1 , \1053_B[3]_b1 );
not ( \1053_B[3]_b1 , w_1708 );
and ( \1135_b0 , \1052_A[3]_b0 , w_1709 );
and ( w_1708 , w_1709 , \1053_B[3]_b0 );
or ( \1136_b1 , \1053_B[3]_b1 , \1058_b1 );
not ( \1058_b1 , w_1710 );
and ( \1136_b0 , \1053_B[3]_b0 , w_1711 );
and ( w_1710 , w_1711 , \1058_b0 );
or ( \1137_b1 , \1052_A[3]_b1 , \1058_b1 );
not ( \1058_b1 , w_1712 );
and ( \1137_b0 , \1052_A[3]_b0 , w_1713 );
and ( w_1712 , w_1713 , \1058_b0 );
or ( \1139_b1 , \1134_b1 , \1138_b1 );
xor ( \1139_b0 , \1134_b0 , w_1714 );
not ( w_1714 , w_1715 );
and ( w_1715 , \1138_b1 , \1138_b0 );
buf ( \1140_SUM[4]_b1 , \1139_b1 );
buf ( \1140_SUM[4]_b0 , \1139_b0 );
or ( \1141_b1 , \1140_SUM[4]_b1 , \863_b1 );
not ( \863_b1 , w_1716 );
and ( \1141_b0 , \1140_SUM[4]_b0 , w_1717 );
and ( w_1716 , w_1717 , \863_b0 );
buf ( \1142_A[4]_b1 , \a[4]_b1 );
buf ( \1142_A[4]_b0 , \a[4]_b0 );
buf ( \1143_B[4]_b1 , \c[4]_b1 );
buf ( \1143_B[4]_b0 , \c[4]_b0 );
or ( \1144_b1 , \1142_A[4]_b1 , \1143_B[4]_b1 );
xor ( \1144_b0 , \1142_A[4]_b0 , w_1718 );
not ( w_1718 , w_1719 );
and ( w_1719 , \1143_B[4]_b1 , \1143_B[4]_b0 );
or ( \1145_b1 , \1062_A[3]_b1 , \1063_B[3]_b1 );
not ( \1063_B[3]_b1 , w_1720 );
and ( \1145_b0 , \1062_A[3]_b0 , w_1721 );
and ( w_1720 , w_1721 , \1063_B[3]_b0 );
or ( \1146_b1 , \1063_B[3]_b1 , \1068_b1 );
not ( \1068_b1 , w_1722 );
and ( \1146_b0 , \1063_B[3]_b0 , w_1723 );
and ( w_1722 , w_1723 , \1068_b0 );
or ( \1147_b1 , \1062_A[3]_b1 , \1068_b1 );
not ( \1068_b1 , w_1724 );
and ( \1147_b0 , \1062_A[3]_b0 , w_1725 );
and ( w_1724 , w_1725 , \1068_b0 );
or ( \1149_b1 , \1144_b1 , \1148_b1 );
xor ( \1149_b0 , \1144_b0 , w_1726 );
not ( w_1726 , w_1727 );
and ( w_1727 , \1148_b1 , \1148_b0 );
buf ( \1150_SUM[4]_b1 , \1149_b1 );
buf ( \1150_SUM[4]_b0 , \1149_b0 );
or ( \1151_b1 , \1150_SUM[4]_b1 , \861_b1 );
not ( \861_b1 , w_1728 );
and ( \1151_b0 , \1150_SUM[4]_b0 , w_1729 );
and ( w_1728 , w_1729 , \861_b0 );
or ( \1152_b1 , \d[4]_b1 , \859_b1 );
not ( \859_b1 , w_1730 );
and ( \1152_b0 , \d[4]_b0 , w_1731 );
and ( w_1730 , w_1731 , \859_b0 );
or ( \1153_b1 , \c[4]_b1 , \857_b1 );
not ( \857_b1 , w_1732 );
and ( \1153_b0 , \c[4]_b0 , w_1733 );
and ( w_1732 , w_1733 , \857_b0 );
or ( \1154_b1 , \b[4]_b1 , \855_b1 );
not ( \855_b1 , w_1734 );
and ( \1154_b0 , \b[4]_b0 , w_1735 );
and ( w_1734 , w_1735 , \855_b0 );
or ( \1155_b1 , \a[4]_b1 , \853_b1 );
not ( \853_b1 , w_1736 );
and ( \1155_b0 , \a[4]_b0 , w_1737 );
and ( w_1736 , w_1737 , \853_b0 );
and ( \1157_b1 , 1'b0_b1 , w_1738 );
xor ( w_1738 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1739 );
and ( \1157_b0 , w_1739 , \876_b0 );
or ( \1158_b1 , \a[5]_b1 , w_1740 );
or ( \1158_b0 , \a[5]_b0 , \d[5]_b0 );
not ( \d[5]_b0 , w_1741 );
and ( w_1741 , w_1740 , \d[5]_b1 );
or ( \1159_b1 , \1158_b1 , \875_b1 );
not ( \875_b1 , w_1742 );
and ( \1159_b0 , \1158_b0 , w_1743 );
and ( w_1742 , w_1743 , \875_b0 );
or ( \1160_b1 , \b[5]_b1 , \c[5]_b1 );
not ( \c[5]_b1 , w_1744 );
and ( \1160_b0 , \b[5]_b0 , w_1745 );
and ( w_1744 , w_1745 , \c[5]_b0 );
or ( \1161_b1 , \1160_b1 , \873_b1 );
not ( \873_b1 , w_1746 );
and ( \1161_b0 , \1160_b0 , w_1747 );
and ( w_1746 , w_1747 , \873_b0 );
or ( \1162_b1 , \a[5]_b1 , w_1748 );
or ( \1162_b0 , \a[5]_b0 , \b[5]_b0 );
not ( \b[5]_b0 , w_1749 );
and ( w_1749 , w_1748 , \b[5]_b1 );
or ( \1163_b1 , \1162_b1 , \871_b1 );
not ( \871_b1 , w_1750 );
and ( \1163_b0 , \1162_b0 , w_1751 );
and ( w_1750 , w_1751 , \871_b0 );
or ( \1164_b1 , \c[5]_b1 , \d[5]_b1 );
xor ( \1164_b0 , \c[5]_b0 , w_1752 );
not ( w_1752 , w_1753 );
and ( w_1753 , \d[5]_b1 , \d[5]_b0 );
or ( \1165_b1 , \1164_b1 , \869_b1 );
not ( \869_b1 , w_1754 );
and ( \1165_b0 , \1164_b0 , w_1755 );
and ( w_1754 , w_1755 , \869_b0 );
buf ( \1166_A[5]_b1 , \b[5]_b1 );
buf ( \1166_A[5]_b0 , \b[5]_b0 );
or ( \1167_b1 , \1166_A[5]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1756 );
and ( \1167_b0 , \1166_A[5]_b0 , w_1757 );
and ( w_1756 , w_1757 , \887_B[0]_b0 );
or ( \1168_b1 , \1086_A[4]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_1758 );
and ( \1168_b0 , \1086_A[4]_b0 , w_1759 );
and ( w_1758 , w_1759 , \922_B[1]_b0 );
or ( \1169_b1 , \1167_b1 , \1168_b1 );
xor ( \1169_b0 , \1167_b0 , w_1760 );
not ( w_1760 , w_1761 );
and ( w_1761 , \1168_b1 , \1168_b0 );
or ( \1170_b1 , \1087_b1 , \1088_b1 );
not ( \1088_b1 , w_1762 );
and ( \1170_b0 , \1087_b0 , w_1763 );
and ( w_1762 , w_1763 , \1088_b0 );
or ( \1171_b1 , \1089_b1 , \1092_b1 );
not ( \1092_b1 , w_1764 );
and ( \1171_b0 , \1089_b0 , w_1765 );
and ( w_1764 , w_1765 , \1092_b0 );
or ( \1172_b1 , \1170_b1 , w_1766 );
or ( \1172_b0 , \1170_b0 , \1171_b0 );
not ( \1171_b0 , w_1767 );
and ( w_1767 , w_1766 , \1171_b1 );
or ( \1173_b1 , \1169_b1 , \1172_b1 );
xor ( \1173_b0 , \1169_b0 , w_1768 );
not ( w_1768 , w_1769 );
and ( w_1769 , \1172_b1 , \1172_b0 );
or ( \1174_b1 , \1018_A[3]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_1770 );
and ( \1174_b0 , \1018_A[3]_b0 , w_1771 );
and ( w_1770 , w_1771 , \968_B[2]_b0 );
or ( \1175_b1 , \1173_b1 , \1174_b1 );
xor ( \1175_b0 , \1173_b0 , w_1772 );
not ( w_1772 , w_1773 );
and ( w_1773 , \1174_b1 , \1174_b0 );
or ( \1176_b1 , \1093_b1 , \1094_b1 );
not ( \1094_b1 , w_1774 );
and ( \1176_b0 , \1093_b0 , w_1775 );
and ( w_1774 , w_1775 , \1094_b0 );
or ( \1177_b1 , \1095_b1 , \1098_b1 );
not ( \1098_b1 , w_1776 );
and ( \1177_b0 , \1095_b0 , w_1777 );
and ( w_1776 , w_1777 , \1098_b0 );
or ( \1178_b1 , \1176_b1 , w_1778 );
or ( \1178_b0 , \1176_b0 , \1177_b0 );
not ( \1177_b0 , w_1779 );
and ( w_1779 , w_1778 , \1177_b1 );
or ( \1179_b1 , \1175_b1 , \1178_b1 );
xor ( \1179_b0 , \1175_b0 , w_1780 );
not ( w_1780 , w_1781 );
and ( w_1781 , \1178_b1 , \1178_b0 );
or ( \1180_b1 , \962_A[2]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_1782 );
and ( \1180_b0 , \962_A[2]_b0 , w_1783 );
and ( w_1782 , w_1783 , \1030_B[3]_b0 );
or ( \1181_b1 , \1179_b1 , \1180_b1 );
xor ( \1181_b0 , \1179_b0 , w_1784 );
not ( w_1784 , w_1785 );
and ( w_1785 , \1180_b1 , \1180_b0 );
or ( \1182_b1 , \1099_b1 , \1100_b1 );
not ( \1100_b1 , w_1786 );
and ( \1182_b0 , \1099_b0 , w_1787 );
and ( w_1786 , w_1787 , \1100_b0 );
or ( \1183_b1 , \1101_b1 , \1102_b1 );
not ( \1102_b1 , w_1788 );
and ( \1183_b0 , \1101_b0 , w_1789 );
and ( w_1788 , w_1789 , \1102_b0 );
or ( \1184_b1 , \1182_b1 , w_1790 );
or ( \1184_b0 , \1182_b0 , \1183_b0 );
not ( \1183_b0 , w_1791 );
and ( w_1791 , w_1790 , \1183_b1 );
or ( \1185_b1 , \1181_b1 , \1184_b1 );
xor ( \1185_b0 , \1181_b0 , w_1792 );
not ( w_1792 , w_1793 );
and ( w_1793 , \1184_b1 , \1184_b0 );
or ( \1186_b1 , \920_A[1]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_1794 );
and ( \1186_b0 , \920_A[1]_b0 , w_1795 );
and ( w_1794 , w_1795 , \1104_B[4]_b0 );
or ( \1187_b1 , \1185_b1 , \1186_b1 );
xor ( \1187_b0 , \1185_b0 , w_1796 );
not ( w_1796 , w_1797 );
and ( w_1797 , \1186_b1 , \1186_b0 );
or ( \1188_b1 , \1103_b1 , \1105_b1 );
not ( \1105_b1 , w_1798 );
and ( \1188_b0 , \1103_b0 , w_1799 );
and ( w_1798 , w_1799 , \1105_b0 );
or ( \1189_b1 , \1187_b1 , \1188_b1 );
xor ( \1189_b0 , \1187_b0 , w_1800 );
not ( w_1800 , w_1801 );
and ( w_1801 , \1188_b1 , \1188_b0 );
buf ( \1190_B[5]_b1 , \c[5]_b1 );
buf ( \1190_B[5]_b0 , \c[5]_b0 );
or ( \1191_b1 , \886_A[0]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_1802 );
and ( \1191_b0 , \886_A[0]_b0 , w_1803 );
and ( w_1802 , w_1803 , \1190_B[5]_b0 );
or ( \1192_b1 , \1189_b1 , \1191_b1 );
xor ( \1192_b0 , \1189_b0 , w_1804 );
not ( w_1804 , w_1805 );
and ( w_1805 , \1191_b1 , \1191_b0 );
buf ( \1193_Z[5]_b1 , \1192_b1 );
buf ( \1193_Z[5]_b0 , \1192_b0 );
or ( \1194_b1 , \1193_Z[5]_b1 , \867_b1 );
not ( \867_b1 , w_1806 );
and ( \1194_b0 , \1193_Z[5]_b0 , w_1807 );
and ( w_1806 , w_1807 , \867_b0 );
buf ( \1195_A[5]_b1 , \a[5]_b1 );
buf ( \1195_A[5]_b0 , \a[5]_b0 );
or ( \1196_b1 , \1195_A[5]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1808 );
and ( \1196_b0 , \1195_A[5]_b0 , w_1809 );
and ( w_1808 , w_1809 , \892_B[0]_b0 );
or ( \1197_b1 , \1109_A[4]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_1810 );
and ( \1197_b0 , \1109_A[4]_b0 , w_1811 );
and ( w_1810 , w_1811 , \929_B[1]_b0 );
or ( \1198_b1 , \1196_b1 , \1197_b1 );
xor ( \1198_b0 , \1196_b0 , w_1812 );
not ( w_1812 , w_1813 );
and ( w_1813 , \1197_b1 , \1197_b0 );
or ( \1199_b1 , \1110_b1 , \1111_b1 );
not ( \1111_b1 , w_1814 );
and ( \1199_b0 , \1110_b0 , w_1815 );
and ( w_1814 , w_1815 , \1111_b0 );
or ( \1200_b1 , \1112_b1 , \1115_b1 );
not ( \1115_b1 , w_1816 );
and ( \1200_b0 , \1112_b0 , w_1817 );
and ( w_1816 , w_1817 , \1115_b0 );
or ( \1201_b1 , \1199_b1 , w_1818 );
or ( \1201_b0 , \1199_b0 , \1200_b0 );
not ( \1200_b0 , w_1819 );
and ( w_1819 , w_1818 , \1200_b1 );
or ( \1202_b1 , \1198_b1 , \1201_b1 );
xor ( \1202_b0 , \1198_b0 , w_1820 );
not ( w_1820 , w_1821 );
and ( w_1821 , \1201_b1 , \1201_b0 );
or ( \1203_b1 , \1035_A[3]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_1822 );
and ( \1203_b0 , \1035_A[3]_b0 , w_1823 );
and ( w_1822 , w_1823 , \979_B[2]_b0 );
or ( \1204_b1 , \1202_b1 , \1203_b1 );
xor ( \1204_b0 , \1202_b0 , w_1824 );
not ( w_1824 , w_1825 );
and ( w_1825 , \1203_b1 , \1203_b0 );
or ( \1205_b1 , \1116_b1 , \1117_b1 );
not ( \1117_b1 , w_1826 );
and ( \1205_b0 , \1116_b0 , w_1827 );
and ( w_1826 , w_1827 , \1117_b0 );
or ( \1206_b1 , \1118_b1 , \1121_b1 );
not ( \1121_b1 , w_1828 );
and ( \1206_b0 , \1118_b0 , w_1829 );
and ( w_1828 , w_1829 , \1121_b0 );
or ( \1207_b1 , \1205_b1 , w_1830 );
or ( \1207_b0 , \1205_b0 , \1206_b0 );
not ( \1206_b0 , w_1831 );
and ( w_1831 , w_1830 , \1206_b1 );
or ( \1208_b1 , \1204_b1 , \1207_b1 );
xor ( \1208_b0 , \1204_b0 , w_1832 );
not ( w_1832 , w_1833 );
and ( w_1833 , \1207_b1 , \1207_b0 );
or ( \1209_b1 , \973_A[2]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_1834 );
and ( \1209_b0 , \973_A[2]_b0 , w_1835 );
and ( w_1834 , w_1835 , \1047_B[3]_b0 );
or ( \1210_b1 , \1208_b1 , \1209_b1 );
xor ( \1210_b0 , \1208_b0 , w_1836 );
not ( w_1836 , w_1837 );
and ( w_1837 , \1209_b1 , \1209_b0 );
or ( \1211_b1 , \1122_b1 , \1123_b1 );
not ( \1123_b1 , w_1838 );
and ( \1211_b0 , \1122_b0 , w_1839 );
and ( w_1838 , w_1839 , \1123_b0 );
or ( \1212_b1 , \1124_b1 , \1125_b1 );
not ( \1125_b1 , w_1840 );
and ( \1212_b0 , \1124_b0 , w_1841 );
and ( w_1840 , w_1841 , \1125_b0 );
or ( \1213_b1 , \1211_b1 , w_1842 );
or ( \1213_b0 , \1211_b0 , \1212_b0 );
not ( \1212_b0 , w_1843 );
and ( w_1843 , w_1842 , \1212_b1 );
or ( \1214_b1 , \1210_b1 , \1213_b1 );
xor ( \1214_b0 , \1210_b0 , w_1844 );
not ( w_1844 , w_1845 );
and ( w_1845 , \1213_b1 , \1213_b0 );
or ( \1215_b1 , \927_A[1]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_1846 );
and ( \1215_b0 , \927_A[1]_b0 , w_1847 );
and ( w_1846 , w_1847 , \1127_B[4]_b0 );
or ( \1216_b1 , \1214_b1 , \1215_b1 );
xor ( \1216_b0 , \1214_b0 , w_1848 );
not ( w_1848 , w_1849 );
and ( w_1849 , \1215_b1 , \1215_b0 );
or ( \1217_b1 , \1126_b1 , \1128_b1 );
not ( \1128_b1 , w_1850 );
and ( \1217_b0 , \1126_b0 , w_1851 );
and ( w_1850 , w_1851 , \1128_b0 );
or ( \1218_b1 , \1216_b1 , \1217_b1 );
xor ( \1218_b0 , \1216_b0 , w_1852 );
not ( w_1852 , w_1853 );
and ( w_1853 , \1217_b1 , \1217_b0 );
buf ( \1219_B[5]_b1 , \d[5]_b1 );
buf ( \1219_B[5]_b0 , \d[5]_b0 );
or ( \1220_b1 , \891_A[0]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_1854 );
and ( \1220_b0 , \891_A[0]_b0 , w_1855 );
and ( w_1854 , w_1855 , \1219_B[5]_b0 );
or ( \1221_b1 , \1218_b1 , \1220_b1 );
xor ( \1221_b0 , \1218_b0 , w_1856 );
not ( w_1856 , w_1857 );
and ( w_1857 , \1220_b1 , \1220_b0 );
buf ( \1222_Z[5]_b1 , \1221_b1 );
buf ( \1222_Z[5]_b0 , \1221_b0 );
or ( \1223_b1 , \1222_Z[5]_b1 , \865_b1 );
not ( \865_b1 , w_1858 );
and ( \1223_b0 , \1222_Z[5]_b0 , w_1859 );
and ( w_1858 , w_1859 , \865_b0 );
buf ( \1224_A[5]_b1 , \b[5]_b1 );
buf ( \1224_A[5]_b0 , \b[5]_b0 );
buf ( \1225_B[5]_b1 , \d[5]_b1 );
buf ( \1225_B[5]_b0 , \d[5]_b0 );
or ( \1226_b1 , \1224_A[5]_b1 , \1225_B[5]_b1 );
xor ( \1226_b0 , \1224_A[5]_b0 , w_1860 );
not ( w_1860 , w_1861 );
and ( w_1861 , \1225_B[5]_b1 , \1225_B[5]_b0 );
or ( \1227_b1 , \1132_A[4]_b1 , \1133_B[4]_b1 );
not ( \1133_B[4]_b1 , w_1862 );
and ( \1227_b0 , \1132_A[4]_b0 , w_1863 );
and ( w_1862 , w_1863 , \1133_B[4]_b0 );
or ( \1228_b1 , \1133_B[4]_b1 , \1138_b1 );
not ( \1138_b1 , w_1864 );
and ( \1228_b0 , \1133_B[4]_b0 , w_1865 );
and ( w_1864 , w_1865 , \1138_b0 );
or ( \1229_b1 , \1132_A[4]_b1 , \1138_b1 );
not ( \1138_b1 , w_1866 );
and ( \1229_b0 , \1132_A[4]_b0 , w_1867 );
and ( w_1866 , w_1867 , \1138_b0 );
or ( \1231_b1 , \1226_b1 , \1230_b1 );
xor ( \1231_b0 , \1226_b0 , w_1868 );
not ( w_1868 , w_1869 );
and ( w_1869 , \1230_b1 , \1230_b0 );
buf ( \1232_SUM[5]_b1 , \1231_b1 );
buf ( \1232_SUM[5]_b0 , \1231_b0 );
or ( \1233_b1 , \1232_SUM[5]_b1 , \863_b1 );
not ( \863_b1 , w_1870 );
and ( \1233_b0 , \1232_SUM[5]_b0 , w_1871 );
and ( w_1870 , w_1871 , \863_b0 );
buf ( \1234_A[5]_b1 , \a[5]_b1 );
buf ( \1234_A[5]_b0 , \a[5]_b0 );
buf ( \1235_B[5]_b1 , \c[5]_b1 );
buf ( \1235_B[5]_b0 , \c[5]_b0 );
or ( \1236_b1 , \1234_A[5]_b1 , \1235_B[5]_b1 );
xor ( \1236_b0 , \1234_A[5]_b0 , w_1872 );
not ( w_1872 , w_1873 );
and ( w_1873 , \1235_B[5]_b1 , \1235_B[5]_b0 );
or ( \1237_b1 , \1142_A[4]_b1 , \1143_B[4]_b1 );
not ( \1143_B[4]_b1 , w_1874 );
and ( \1237_b0 , \1142_A[4]_b0 , w_1875 );
and ( w_1874 , w_1875 , \1143_B[4]_b0 );
or ( \1238_b1 , \1143_B[4]_b1 , \1148_b1 );
not ( \1148_b1 , w_1876 );
and ( \1238_b0 , \1143_B[4]_b0 , w_1877 );
and ( w_1876 , w_1877 , \1148_b0 );
or ( \1239_b1 , \1142_A[4]_b1 , \1148_b1 );
not ( \1148_b1 , w_1878 );
and ( \1239_b0 , \1142_A[4]_b0 , w_1879 );
and ( w_1878 , w_1879 , \1148_b0 );
or ( \1241_b1 , \1236_b1 , \1240_b1 );
xor ( \1241_b0 , \1236_b0 , w_1880 );
not ( w_1880 , w_1881 );
and ( w_1881 , \1240_b1 , \1240_b0 );
buf ( \1242_SUM[5]_b1 , \1241_b1 );
buf ( \1242_SUM[5]_b0 , \1241_b0 );
or ( \1243_b1 , \1242_SUM[5]_b1 , \861_b1 );
not ( \861_b1 , w_1882 );
and ( \1243_b0 , \1242_SUM[5]_b0 , w_1883 );
and ( w_1882 , w_1883 , \861_b0 );
or ( \1244_b1 , \d[5]_b1 , \859_b1 );
not ( \859_b1 , w_1884 );
and ( \1244_b0 , \d[5]_b0 , w_1885 );
and ( w_1884 , w_1885 , \859_b0 );
or ( \1245_b1 , \c[5]_b1 , \857_b1 );
not ( \857_b1 , w_1886 );
and ( \1245_b0 , \c[5]_b0 , w_1887 );
and ( w_1886 , w_1887 , \857_b0 );
or ( \1246_b1 , \b[5]_b1 , \855_b1 );
not ( \855_b1 , w_1888 );
and ( \1246_b0 , \b[5]_b0 , w_1889 );
and ( w_1888 , w_1889 , \855_b0 );
or ( \1247_b1 , \a[5]_b1 , \853_b1 );
not ( \853_b1 , w_1890 );
and ( \1247_b0 , \a[5]_b0 , w_1891 );
and ( w_1890 , w_1891 , \853_b0 );
and ( \1249_b1 , 1'b0_b1 , w_1892 );
xor ( w_1892 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_1893 );
and ( \1249_b0 , w_1893 , \876_b0 );
or ( \1250_b1 , \a[6]_b1 , w_1894 );
or ( \1250_b0 , \a[6]_b0 , \d[6]_b0 );
not ( \d[6]_b0 , w_1895 );
and ( w_1895 , w_1894 , \d[6]_b1 );
or ( \1251_b1 , \1250_b1 , \875_b1 );
not ( \875_b1 , w_1896 );
and ( \1251_b0 , \1250_b0 , w_1897 );
and ( w_1896 , w_1897 , \875_b0 );
or ( \1252_b1 , \b[6]_b1 , \c[6]_b1 );
not ( \c[6]_b1 , w_1898 );
and ( \1252_b0 , \b[6]_b0 , w_1899 );
and ( w_1898 , w_1899 , \c[6]_b0 );
or ( \1253_b1 , \1252_b1 , \873_b1 );
not ( \873_b1 , w_1900 );
and ( \1253_b0 , \1252_b0 , w_1901 );
and ( w_1900 , w_1901 , \873_b0 );
or ( \1254_b1 , \a[6]_b1 , w_1902 );
or ( \1254_b0 , \a[6]_b0 , \b[6]_b0 );
not ( \b[6]_b0 , w_1903 );
and ( w_1903 , w_1902 , \b[6]_b1 );
or ( \1255_b1 , \1254_b1 , \871_b1 );
not ( \871_b1 , w_1904 );
and ( \1255_b0 , \1254_b0 , w_1905 );
and ( w_1904 , w_1905 , \871_b0 );
or ( \1256_b1 , \c[6]_b1 , \d[6]_b1 );
xor ( \1256_b0 , \c[6]_b0 , w_1906 );
not ( w_1906 , w_1907 );
and ( w_1907 , \d[6]_b1 , \d[6]_b0 );
or ( \1257_b1 , \1256_b1 , \869_b1 );
not ( \869_b1 , w_1908 );
and ( \1257_b0 , \1256_b0 , w_1909 );
and ( w_1908 , w_1909 , \869_b0 );
buf ( \1258_A[6]_b1 , \b[6]_b1 );
buf ( \1258_A[6]_b0 , \b[6]_b0 );
or ( \1259_b1 , \1258_A[6]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_1910 );
and ( \1259_b0 , \1258_A[6]_b0 , w_1911 );
and ( w_1910 , w_1911 , \887_B[0]_b0 );
or ( \1260_b1 , \1166_A[5]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_1912 );
and ( \1260_b0 , \1166_A[5]_b0 , w_1913 );
and ( w_1912 , w_1913 , \922_B[1]_b0 );
or ( \1261_b1 , \1259_b1 , \1260_b1 );
xor ( \1261_b0 , \1259_b0 , w_1914 );
not ( w_1914 , w_1915 );
and ( w_1915 , \1260_b1 , \1260_b0 );
or ( \1262_b1 , \1167_b1 , \1168_b1 );
not ( \1168_b1 , w_1916 );
and ( \1262_b0 , \1167_b0 , w_1917 );
and ( w_1916 , w_1917 , \1168_b0 );
or ( \1263_b1 , \1169_b1 , \1172_b1 );
not ( \1172_b1 , w_1918 );
and ( \1263_b0 , \1169_b0 , w_1919 );
and ( w_1918 , w_1919 , \1172_b0 );
or ( \1264_b1 , \1262_b1 , w_1920 );
or ( \1264_b0 , \1262_b0 , \1263_b0 );
not ( \1263_b0 , w_1921 );
and ( w_1921 , w_1920 , \1263_b1 );
or ( \1265_b1 , \1261_b1 , \1264_b1 );
xor ( \1265_b0 , \1261_b0 , w_1922 );
not ( w_1922 , w_1923 );
and ( w_1923 , \1264_b1 , \1264_b0 );
or ( \1266_b1 , \1086_A[4]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_1924 );
and ( \1266_b0 , \1086_A[4]_b0 , w_1925 );
and ( w_1924 , w_1925 , \968_B[2]_b0 );
or ( \1267_b1 , \1265_b1 , \1266_b1 );
xor ( \1267_b0 , \1265_b0 , w_1926 );
not ( w_1926 , w_1927 );
and ( w_1927 , \1266_b1 , \1266_b0 );
or ( \1268_b1 , \1173_b1 , \1174_b1 );
not ( \1174_b1 , w_1928 );
and ( \1268_b0 , \1173_b0 , w_1929 );
and ( w_1928 , w_1929 , \1174_b0 );
or ( \1269_b1 , \1175_b1 , \1178_b1 );
not ( \1178_b1 , w_1930 );
and ( \1269_b0 , \1175_b0 , w_1931 );
and ( w_1930 , w_1931 , \1178_b0 );
or ( \1270_b1 , \1268_b1 , w_1932 );
or ( \1270_b0 , \1268_b0 , \1269_b0 );
not ( \1269_b0 , w_1933 );
and ( w_1933 , w_1932 , \1269_b1 );
or ( \1271_b1 , \1267_b1 , \1270_b1 );
xor ( \1271_b0 , \1267_b0 , w_1934 );
not ( w_1934 , w_1935 );
and ( w_1935 , \1270_b1 , \1270_b0 );
or ( \1272_b1 , \1018_A[3]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_1936 );
and ( \1272_b0 , \1018_A[3]_b0 , w_1937 );
and ( w_1936 , w_1937 , \1030_B[3]_b0 );
or ( \1273_b1 , \1271_b1 , \1272_b1 );
xor ( \1273_b0 , \1271_b0 , w_1938 );
not ( w_1938 , w_1939 );
and ( w_1939 , \1272_b1 , \1272_b0 );
or ( \1274_b1 , \1179_b1 , \1180_b1 );
not ( \1180_b1 , w_1940 );
and ( \1274_b0 , \1179_b0 , w_1941 );
and ( w_1940 , w_1941 , \1180_b0 );
or ( \1275_b1 , \1181_b1 , \1184_b1 );
not ( \1184_b1 , w_1942 );
and ( \1275_b0 , \1181_b0 , w_1943 );
and ( w_1942 , w_1943 , \1184_b0 );
or ( \1276_b1 , \1274_b1 , w_1944 );
or ( \1276_b0 , \1274_b0 , \1275_b0 );
not ( \1275_b0 , w_1945 );
and ( w_1945 , w_1944 , \1275_b1 );
or ( \1277_b1 , \1273_b1 , \1276_b1 );
xor ( \1277_b0 , \1273_b0 , w_1946 );
not ( w_1946 , w_1947 );
and ( w_1947 , \1276_b1 , \1276_b0 );
or ( \1278_b1 , \962_A[2]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_1948 );
and ( \1278_b0 , \962_A[2]_b0 , w_1949 );
and ( w_1948 , w_1949 , \1104_B[4]_b0 );
or ( \1279_b1 , \1277_b1 , \1278_b1 );
xor ( \1279_b0 , \1277_b0 , w_1950 );
not ( w_1950 , w_1951 );
and ( w_1951 , \1278_b1 , \1278_b0 );
or ( \1280_b1 , \1185_b1 , \1186_b1 );
not ( \1186_b1 , w_1952 );
and ( \1280_b0 , \1185_b0 , w_1953 );
and ( w_1952 , w_1953 , \1186_b0 );
or ( \1281_b1 , \1187_b1 , \1188_b1 );
not ( \1188_b1 , w_1954 );
and ( \1281_b0 , \1187_b0 , w_1955 );
and ( w_1954 , w_1955 , \1188_b0 );
or ( \1282_b1 , \1280_b1 , w_1956 );
or ( \1282_b0 , \1280_b0 , \1281_b0 );
not ( \1281_b0 , w_1957 );
and ( w_1957 , w_1956 , \1281_b1 );
or ( \1283_b1 , \1279_b1 , \1282_b1 );
xor ( \1283_b0 , \1279_b0 , w_1958 );
not ( w_1958 , w_1959 );
and ( w_1959 , \1282_b1 , \1282_b0 );
or ( \1284_b1 , \920_A[1]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_1960 );
and ( \1284_b0 , \920_A[1]_b0 , w_1961 );
and ( w_1960 , w_1961 , \1190_B[5]_b0 );
or ( \1285_b1 , \1283_b1 , \1284_b1 );
xor ( \1285_b0 , \1283_b0 , w_1962 );
not ( w_1962 , w_1963 );
and ( w_1963 , \1284_b1 , \1284_b0 );
or ( \1286_b1 , \1189_b1 , \1191_b1 );
not ( \1191_b1 , w_1964 );
and ( \1286_b0 , \1189_b0 , w_1965 );
and ( w_1964 , w_1965 , \1191_b0 );
or ( \1287_b1 , \1285_b1 , \1286_b1 );
xor ( \1287_b0 , \1285_b0 , w_1966 );
not ( w_1966 , w_1967 );
and ( w_1967 , \1286_b1 , \1286_b0 );
buf ( \1288_B[6]_b1 , \c[6]_b1 );
buf ( \1288_B[6]_b0 , \c[6]_b0 );
or ( \1289_b1 , \886_A[0]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_1968 );
and ( \1289_b0 , \886_A[0]_b0 , w_1969 );
and ( w_1968 , w_1969 , \1288_B[6]_b0 );
or ( \1290_b1 , \1287_b1 , \1289_b1 );
xor ( \1290_b0 , \1287_b0 , w_1970 );
not ( w_1970 , w_1971 );
and ( w_1971 , \1289_b1 , \1289_b0 );
buf ( \1291_Z[6]_b1 , \1290_b1 );
buf ( \1291_Z[6]_b0 , \1290_b0 );
or ( \1292_b1 , \1291_Z[6]_b1 , \867_b1 );
not ( \867_b1 , w_1972 );
and ( \1292_b0 , \1291_Z[6]_b0 , w_1973 );
and ( w_1972 , w_1973 , \867_b0 );
buf ( \1293_A[6]_b1 , \a[6]_b1 );
buf ( \1293_A[6]_b0 , \a[6]_b0 );
or ( \1294_b1 , \1293_A[6]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_1974 );
and ( \1294_b0 , \1293_A[6]_b0 , w_1975 );
and ( w_1974 , w_1975 , \892_B[0]_b0 );
or ( \1295_b1 , \1195_A[5]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_1976 );
and ( \1295_b0 , \1195_A[5]_b0 , w_1977 );
and ( w_1976 , w_1977 , \929_B[1]_b0 );
or ( \1296_b1 , \1294_b1 , \1295_b1 );
xor ( \1296_b0 , \1294_b0 , w_1978 );
not ( w_1978 , w_1979 );
and ( w_1979 , \1295_b1 , \1295_b0 );
or ( \1297_b1 , \1196_b1 , \1197_b1 );
not ( \1197_b1 , w_1980 );
and ( \1297_b0 , \1196_b0 , w_1981 );
and ( w_1980 , w_1981 , \1197_b0 );
or ( \1298_b1 , \1198_b1 , \1201_b1 );
not ( \1201_b1 , w_1982 );
and ( \1298_b0 , \1198_b0 , w_1983 );
and ( w_1982 , w_1983 , \1201_b0 );
or ( \1299_b1 , \1297_b1 , w_1984 );
or ( \1299_b0 , \1297_b0 , \1298_b0 );
not ( \1298_b0 , w_1985 );
and ( w_1985 , w_1984 , \1298_b1 );
or ( \1300_b1 , \1296_b1 , \1299_b1 );
xor ( \1300_b0 , \1296_b0 , w_1986 );
not ( w_1986 , w_1987 );
and ( w_1987 , \1299_b1 , \1299_b0 );
or ( \1301_b1 , \1109_A[4]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_1988 );
and ( \1301_b0 , \1109_A[4]_b0 , w_1989 );
and ( w_1988 , w_1989 , \979_B[2]_b0 );
or ( \1302_b1 , \1300_b1 , \1301_b1 );
xor ( \1302_b0 , \1300_b0 , w_1990 );
not ( w_1990 , w_1991 );
and ( w_1991 , \1301_b1 , \1301_b0 );
or ( \1303_b1 , \1202_b1 , \1203_b1 );
not ( \1203_b1 , w_1992 );
and ( \1303_b0 , \1202_b0 , w_1993 );
and ( w_1992 , w_1993 , \1203_b0 );
or ( \1304_b1 , \1204_b1 , \1207_b1 );
not ( \1207_b1 , w_1994 );
and ( \1304_b0 , \1204_b0 , w_1995 );
and ( w_1994 , w_1995 , \1207_b0 );
or ( \1305_b1 , \1303_b1 , w_1996 );
or ( \1305_b0 , \1303_b0 , \1304_b0 );
not ( \1304_b0 , w_1997 );
and ( w_1997 , w_1996 , \1304_b1 );
or ( \1306_b1 , \1302_b1 , \1305_b1 );
xor ( \1306_b0 , \1302_b0 , w_1998 );
not ( w_1998 , w_1999 );
and ( w_1999 , \1305_b1 , \1305_b0 );
or ( \1307_b1 , \1035_A[3]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_2000 );
and ( \1307_b0 , \1035_A[3]_b0 , w_2001 );
and ( w_2000 , w_2001 , \1047_B[3]_b0 );
or ( \1308_b1 , \1306_b1 , \1307_b1 );
xor ( \1308_b0 , \1306_b0 , w_2002 );
not ( w_2002 , w_2003 );
and ( w_2003 , \1307_b1 , \1307_b0 );
or ( \1309_b1 , \1208_b1 , \1209_b1 );
not ( \1209_b1 , w_2004 );
and ( \1309_b0 , \1208_b0 , w_2005 );
and ( w_2004 , w_2005 , \1209_b0 );
or ( \1310_b1 , \1210_b1 , \1213_b1 );
not ( \1213_b1 , w_2006 );
and ( \1310_b0 , \1210_b0 , w_2007 );
and ( w_2006 , w_2007 , \1213_b0 );
or ( \1311_b1 , \1309_b1 , w_2008 );
or ( \1311_b0 , \1309_b0 , \1310_b0 );
not ( \1310_b0 , w_2009 );
and ( w_2009 , w_2008 , \1310_b1 );
or ( \1312_b1 , \1308_b1 , \1311_b1 );
xor ( \1312_b0 , \1308_b0 , w_2010 );
not ( w_2010 , w_2011 );
and ( w_2011 , \1311_b1 , \1311_b0 );
or ( \1313_b1 , \973_A[2]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_2012 );
and ( \1313_b0 , \973_A[2]_b0 , w_2013 );
and ( w_2012 , w_2013 , \1127_B[4]_b0 );
or ( \1314_b1 , \1312_b1 , \1313_b1 );
xor ( \1314_b0 , \1312_b0 , w_2014 );
not ( w_2014 , w_2015 );
and ( w_2015 , \1313_b1 , \1313_b0 );
or ( \1315_b1 , \1214_b1 , \1215_b1 );
not ( \1215_b1 , w_2016 );
and ( \1315_b0 , \1214_b0 , w_2017 );
and ( w_2016 , w_2017 , \1215_b0 );
or ( \1316_b1 , \1216_b1 , \1217_b1 );
not ( \1217_b1 , w_2018 );
and ( \1316_b0 , \1216_b0 , w_2019 );
and ( w_2018 , w_2019 , \1217_b0 );
or ( \1317_b1 , \1315_b1 , w_2020 );
or ( \1317_b0 , \1315_b0 , \1316_b0 );
not ( \1316_b0 , w_2021 );
and ( w_2021 , w_2020 , \1316_b1 );
or ( \1318_b1 , \1314_b1 , \1317_b1 );
xor ( \1318_b0 , \1314_b0 , w_2022 );
not ( w_2022 , w_2023 );
and ( w_2023 , \1317_b1 , \1317_b0 );
or ( \1319_b1 , \927_A[1]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_2024 );
and ( \1319_b0 , \927_A[1]_b0 , w_2025 );
and ( w_2024 , w_2025 , \1219_B[5]_b0 );
or ( \1320_b1 , \1318_b1 , \1319_b1 );
xor ( \1320_b0 , \1318_b0 , w_2026 );
not ( w_2026 , w_2027 );
and ( w_2027 , \1319_b1 , \1319_b0 );
or ( \1321_b1 , \1218_b1 , \1220_b1 );
not ( \1220_b1 , w_2028 );
and ( \1321_b0 , \1218_b0 , w_2029 );
and ( w_2028 , w_2029 , \1220_b0 );
or ( \1322_b1 , \1320_b1 , \1321_b1 );
xor ( \1322_b0 , \1320_b0 , w_2030 );
not ( w_2030 , w_2031 );
and ( w_2031 , \1321_b1 , \1321_b0 );
buf ( \1323_B[6]_b1 , \d[6]_b1 );
buf ( \1323_B[6]_b0 , \d[6]_b0 );
or ( \1324_b1 , \891_A[0]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_2032 );
and ( \1324_b0 , \891_A[0]_b0 , w_2033 );
and ( w_2032 , w_2033 , \1323_B[6]_b0 );
or ( \1325_b1 , \1322_b1 , \1324_b1 );
xor ( \1325_b0 , \1322_b0 , w_2034 );
not ( w_2034 , w_2035 );
and ( w_2035 , \1324_b1 , \1324_b0 );
buf ( \1326_Z[6]_b1 , \1325_b1 );
buf ( \1326_Z[6]_b0 , \1325_b0 );
or ( \1327_b1 , \1326_Z[6]_b1 , \865_b1 );
not ( \865_b1 , w_2036 );
and ( \1327_b0 , \1326_Z[6]_b0 , w_2037 );
and ( w_2036 , w_2037 , \865_b0 );
buf ( \1328_A[6]_b1 , \b[6]_b1 );
buf ( \1328_A[6]_b0 , \b[6]_b0 );
buf ( \1329_B[6]_b1 , \d[6]_b1 );
buf ( \1329_B[6]_b0 , \d[6]_b0 );
or ( \1330_b1 , \1328_A[6]_b1 , \1329_B[6]_b1 );
xor ( \1330_b0 , \1328_A[6]_b0 , w_2038 );
not ( w_2038 , w_2039 );
and ( w_2039 , \1329_B[6]_b1 , \1329_B[6]_b0 );
or ( \1331_b1 , \1224_A[5]_b1 , \1225_B[5]_b1 );
not ( \1225_B[5]_b1 , w_2040 );
and ( \1331_b0 , \1224_A[5]_b0 , w_2041 );
and ( w_2040 , w_2041 , \1225_B[5]_b0 );
or ( \1332_b1 , \1225_B[5]_b1 , \1230_b1 );
not ( \1230_b1 , w_2042 );
and ( \1332_b0 , \1225_B[5]_b0 , w_2043 );
and ( w_2042 , w_2043 , \1230_b0 );
or ( \1333_b1 , \1224_A[5]_b1 , \1230_b1 );
not ( \1230_b1 , w_2044 );
and ( \1333_b0 , \1224_A[5]_b0 , w_2045 );
and ( w_2044 , w_2045 , \1230_b0 );
or ( \1335_b1 , \1330_b1 , \1334_b1 );
xor ( \1335_b0 , \1330_b0 , w_2046 );
not ( w_2046 , w_2047 );
and ( w_2047 , \1334_b1 , \1334_b0 );
buf ( \1336_SUM[6]_b1 , \1335_b1 );
buf ( \1336_SUM[6]_b0 , \1335_b0 );
or ( \1337_b1 , \1336_SUM[6]_b1 , \863_b1 );
not ( \863_b1 , w_2048 );
and ( \1337_b0 , \1336_SUM[6]_b0 , w_2049 );
and ( w_2048 , w_2049 , \863_b0 );
buf ( \1338_A[6]_b1 , \a[6]_b1 );
buf ( \1338_A[6]_b0 , \a[6]_b0 );
buf ( \1339_B[6]_b1 , \c[6]_b1 );
buf ( \1339_B[6]_b0 , \c[6]_b0 );
or ( \1340_b1 , \1338_A[6]_b1 , \1339_B[6]_b1 );
xor ( \1340_b0 , \1338_A[6]_b0 , w_2050 );
not ( w_2050 , w_2051 );
and ( w_2051 , \1339_B[6]_b1 , \1339_B[6]_b0 );
or ( \1341_b1 , \1234_A[5]_b1 , \1235_B[5]_b1 );
not ( \1235_B[5]_b1 , w_2052 );
and ( \1341_b0 , \1234_A[5]_b0 , w_2053 );
and ( w_2052 , w_2053 , \1235_B[5]_b0 );
or ( \1342_b1 , \1235_B[5]_b1 , \1240_b1 );
not ( \1240_b1 , w_2054 );
and ( \1342_b0 , \1235_B[5]_b0 , w_2055 );
and ( w_2054 , w_2055 , \1240_b0 );
or ( \1343_b1 , \1234_A[5]_b1 , \1240_b1 );
not ( \1240_b1 , w_2056 );
and ( \1343_b0 , \1234_A[5]_b0 , w_2057 );
and ( w_2056 , w_2057 , \1240_b0 );
or ( \1345_b1 , \1340_b1 , \1344_b1 );
xor ( \1345_b0 , \1340_b0 , w_2058 );
not ( w_2058 , w_2059 );
and ( w_2059 , \1344_b1 , \1344_b0 );
buf ( \1346_SUM[6]_b1 , \1345_b1 );
buf ( \1346_SUM[6]_b0 , \1345_b0 );
or ( \1347_b1 , \1346_SUM[6]_b1 , \861_b1 );
not ( \861_b1 , w_2060 );
and ( \1347_b0 , \1346_SUM[6]_b0 , w_2061 );
and ( w_2060 , w_2061 , \861_b0 );
or ( \1348_b1 , \d[6]_b1 , \859_b1 );
not ( \859_b1 , w_2062 );
and ( \1348_b0 , \d[6]_b0 , w_2063 );
and ( w_2062 , w_2063 , \859_b0 );
or ( \1349_b1 , \c[6]_b1 , \857_b1 );
not ( \857_b1 , w_2064 );
and ( \1349_b0 , \c[6]_b0 , w_2065 );
and ( w_2064 , w_2065 , \857_b0 );
or ( \1350_b1 , \b[6]_b1 , \855_b1 );
not ( \855_b1 , w_2066 );
and ( \1350_b0 , \b[6]_b0 , w_2067 );
and ( w_2066 , w_2067 , \855_b0 );
or ( \1351_b1 , \a[6]_b1 , \853_b1 );
not ( \853_b1 , w_2068 );
and ( \1351_b0 , \a[6]_b0 , w_2069 );
and ( w_2068 , w_2069 , \853_b0 );
and ( \1353_b1 , 1'b0_b1 , w_2070 );
xor ( w_2070 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_2071 );
and ( \1353_b0 , w_2071 , \876_b0 );
or ( \1354_b1 , \a[7]_b1 , w_2072 );
or ( \1354_b0 , \a[7]_b0 , \d[7]_b0 );
not ( \d[7]_b0 , w_2073 );
and ( w_2073 , w_2072 , \d[7]_b1 );
or ( \1355_b1 , \1354_b1 , \875_b1 );
not ( \875_b1 , w_2074 );
and ( \1355_b0 , \1354_b0 , w_2075 );
and ( w_2074 , w_2075 , \875_b0 );
or ( \1356_b1 , \b[7]_b1 , \c[7]_b1 );
not ( \c[7]_b1 , w_2076 );
and ( \1356_b0 , \b[7]_b0 , w_2077 );
and ( w_2076 , w_2077 , \c[7]_b0 );
or ( \1357_b1 , \1356_b1 , \873_b1 );
not ( \873_b1 , w_2078 );
and ( \1357_b0 , \1356_b0 , w_2079 );
and ( w_2078 , w_2079 , \873_b0 );
or ( \1358_b1 , \a[7]_b1 , w_2080 );
or ( \1358_b0 , \a[7]_b0 , \b[7]_b0 );
not ( \b[7]_b0 , w_2081 );
and ( w_2081 , w_2080 , \b[7]_b1 );
or ( \1359_b1 , \1358_b1 , \871_b1 );
not ( \871_b1 , w_2082 );
and ( \1359_b0 , \1358_b0 , w_2083 );
and ( w_2082 , w_2083 , \871_b0 );
or ( \1360_b1 , \c[7]_b1 , \d[7]_b1 );
xor ( \1360_b0 , \c[7]_b0 , w_2084 );
not ( w_2084 , w_2085 );
and ( w_2085 , \d[7]_b1 , \d[7]_b0 );
or ( \1361_b1 , \1360_b1 , \869_b1 );
not ( \869_b1 , w_2086 );
and ( \1361_b0 , \1360_b0 , w_2087 );
and ( w_2086 , w_2087 , \869_b0 );
buf ( \1362_A[7]_b1 , \b[7]_b1 );
buf ( \1362_A[7]_b0 , \b[7]_b0 );
or ( \1363_b1 , \1362_A[7]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_2088 );
and ( \1363_b0 , \1362_A[7]_b0 , w_2089 );
and ( w_2088 , w_2089 , \887_B[0]_b0 );
or ( \1364_b1 , \1258_A[6]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_2090 );
and ( \1364_b0 , \1258_A[6]_b0 , w_2091 );
and ( w_2090 , w_2091 , \922_B[1]_b0 );
or ( \1365_b1 , \1363_b1 , \1364_b1 );
xor ( \1365_b0 , \1363_b0 , w_2092 );
not ( w_2092 , w_2093 );
and ( w_2093 , \1364_b1 , \1364_b0 );
or ( \1366_b1 , \1259_b1 , \1260_b1 );
not ( \1260_b1 , w_2094 );
and ( \1366_b0 , \1259_b0 , w_2095 );
and ( w_2094 , w_2095 , \1260_b0 );
or ( \1367_b1 , \1261_b1 , \1264_b1 );
not ( \1264_b1 , w_2096 );
and ( \1367_b0 , \1261_b0 , w_2097 );
and ( w_2096 , w_2097 , \1264_b0 );
or ( \1368_b1 , \1366_b1 , w_2098 );
or ( \1368_b0 , \1366_b0 , \1367_b0 );
not ( \1367_b0 , w_2099 );
and ( w_2099 , w_2098 , \1367_b1 );
or ( \1369_b1 , \1365_b1 , \1368_b1 );
xor ( \1369_b0 , \1365_b0 , w_2100 );
not ( w_2100 , w_2101 );
and ( w_2101 , \1368_b1 , \1368_b0 );
or ( \1370_b1 , \1166_A[5]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_2102 );
and ( \1370_b0 , \1166_A[5]_b0 , w_2103 );
and ( w_2102 , w_2103 , \968_B[2]_b0 );
or ( \1371_b1 , \1369_b1 , \1370_b1 );
xor ( \1371_b0 , \1369_b0 , w_2104 );
not ( w_2104 , w_2105 );
and ( w_2105 , \1370_b1 , \1370_b0 );
or ( \1372_b1 , \1265_b1 , \1266_b1 );
not ( \1266_b1 , w_2106 );
and ( \1372_b0 , \1265_b0 , w_2107 );
and ( w_2106 , w_2107 , \1266_b0 );
or ( \1373_b1 , \1267_b1 , \1270_b1 );
not ( \1270_b1 , w_2108 );
and ( \1373_b0 , \1267_b0 , w_2109 );
and ( w_2108 , w_2109 , \1270_b0 );
or ( \1374_b1 , \1372_b1 , w_2110 );
or ( \1374_b0 , \1372_b0 , \1373_b0 );
not ( \1373_b0 , w_2111 );
and ( w_2111 , w_2110 , \1373_b1 );
or ( \1375_b1 , \1371_b1 , \1374_b1 );
xor ( \1375_b0 , \1371_b0 , w_2112 );
not ( w_2112 , w_2113 );
and ( w_2113 , \1374_b1 , \1374_b0 );
or ( \1376_b1 , \1086_A[4]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_2114 );
and ( \1376_b0 , \1086_A[4]_b0 , w_2115 );
and ( w_2114 , w_2115 , \1030_B[3]_b0 );
or ( \1377_b1 , \1375_b1 , \1376_b1 );
xor ( \1377_b0 , \1375_b0 , w_2116 );
not ( w_2116 , w_2117 );
and ( w_2117 , \1376_b1 , \1376_b0 );
or ( \1378_b1 , \1271_b1 , \1272_b1 );
not ( \1272_b1 , w_2118 );
and ( \1378_b0 , \1271_b0 , w_2119 );
and ( w_2118 , w_2119 , \1272_b0 );
or ( \1379_b1 , \1273_b1 , \1276_b1 );
not ( \1276_b1 , w_2120 );
and ( \1379_b0 , \1273_b0 , w_2121 );
and ( w_2120 , w_2121 , \1276_b0 );
or ( \1380_b1 , \1378_b1 , w_2122 );
or ( \1380_b0 , \1378_b0 , \1379_b0 );
not ( \1379_b0 , w_2123 );
and ( w_2123 , w_2122 , \1379_b1 );
or ( \1381_b1 , \1377_b1 , \1380_b1 );
xor ( \1381_b0 , \1377_b0 , w_2124 );
not ( w_2124 , w_2125 );
and ( w_2125 , \1380_b1 , \1380_b0 );
or ( \1382_b1 , \1018_A[3]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_2126 );
and ( \1382_b0 , \1018_A[3]_b0 , w_2127 );
and ( w_2126 , w_2127 , \1104_B[4]_b0 );
or ( \1383_b1 , \1381_b1 , \1382_b1 );
xor ( \1383_b0 , \1381_b0 , w_2128 );
not ( w_2128 , w_2129 );
and ( w_2129 , \1382_b1 , \1382_b0 );
or ( \1384_b1 , \1277_b1 , \1278_b1 );
not ( \1278_b1 , w_2130 );
and ( \1384_b0 , \1277_b0 , w_2131 );
and ( w_2130 , w_2131 , \1278_b0 );
or ( \1385_b1 , \1279_b1 , \1282_b1 );
not ( \1282_b1 , w_2132 );
and ( \1385_b0 , \1279_b0 , w_2133 );
and ( w_2132 , w_2133 , \1282_b0 );
or ( \1386_b1 , \1384_b1 , w_2134 );
or ( \1386_b0 , \1384_b0 , \1385_b0 );
not ( \1385_b0 , w_2135 );
and ( w_2135 , w_2134 , \1385_b1 );
or ( \1387_b1 , \1383_b1 , \1386_b1 );
xor ( \1387_b0 , \1383_b0 , w_2136 );
not ( w_2136 , w_2137 );
and ( w_2137 , \1386_b1 , \1386_b0 );
or ( \1388_b1 , \962_A[2]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_2138 );
and ( \1388_b0 , \962_A[2]_b0 , w_2139 );
and ( w_2138 , w_2139 , \1190_B[5]_b0 );
or ( \1389_b1 , \1387_b1 , \1388_b1 );
xor ( \1389_b0 , \1387_b0 , w_2140 );
not ( w_2140 , w_2141 );
and ( w_2141 , \1388_b1 , \1388_b0 );
or ( \1390_b1 , \1283_b1 , \1284_b1 );
not ( \1284_b1 , w_2142 );
and ( \1390_b0 , \1283_b0 , w_2143 );
and ( w_2142 , w_2143 , \1284_b0 );
or ( \1391_b1 , \1285_b1 , \1286_b1 );
not ( \1286_b1 , w_2144 );
and ( \1391_b0 , \1285_b0 , w_2145 );
and ( w_2144 , w_2145 , \1286_b0 );
or ( \1392_b1 , \1390_b1 , w_2146 );
or ( \1392_b0 , \1390_b0 , \1391_b0 );
not ( \1391_b0 , w_2147 );
and ( w_2147 , w_2146 , \1391_b1 );
or ( \1393_b1 , \1389_b1 , \1392_b1 );
xor ( \1393_b0 , \1389_b0 , w_2148 );
not ( w_2148 , w_2149 );
and ( w_2149 , \1392_b1 , \1392_b0 );
or ( \1394_b1 , \920_A[1]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_2150 );
and ( \1394_b0 , \920_A[1]_b0 , w_2151 );
and ( w_2150 , w_2151 , \1288_B[6]_b0 );
or ( \1395_b1 , \1393_b1 , \1394_b1 );
xor ( \1395_b0 , \1393_b0 , w_2152 );
not ( w_2152 , w_2153 );
and ( w_2153 , \1394_b1 , \1394_b0 );
or ( \1396_b1 , \1287_b1 , \1289_b1 );
not ( \1289_b1 , w_2154 );
and ( \1396_b0 , \1287_b0 , w_2155 );
and ( w_2154 , w_2155 , \1289_b0 );
or ( \1397_b1 , \1395_b1 , \1396_b1 );
xor ( \1397_b0 , \1395_b0 , w_2156 );
not ( w_2156 , w_2157 );
and ( w_2157 , \1396_b1 , \1396_b0 );
buf ( \1398_B[7]_b1 , \c[7]_b1 );
buf ( \1398_B[7]_b0 , \c[7]_b0 );
or ( \1399_b1 , \886_A[0]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_2158 );
and ( \1399_b0 , \886_A[0]_b0 , w_2159 );
and ( w_2158 , w_2159 , \1398_B[7]_b0 );
or ( \1400_b1 , \1397_b1 , \1399_b1 );
xor ( \1400_b0 , \1397_b0 , w_2160 );
not ( w_2160 , w_2161 );
and ( w_2161 , \1399_b1 , \1399_b0 );
buf ( \1401_Z[7]_b1 , \1400_b1 );
buf ( \1401_Z[7]_b0 , \1400_b0 );
or ( \1402_b1 , \1401_Z[7]_b1 , \867_b1 );
not ( \867_b1 , w_2162 );
and ( \1402_b0 , \1401_Z[7]_b0 , w_2163 );
and ( w_2162 , w_2163 , \867_b0 );
buf ( \1403_A[7]_b1 , \a[7]_b1 );
buf ( \1403_A[7]_b0 , \a[7]_b0 );
or ( \1404_b1 , \1403_A[7]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_2164 );
and ( \1404_b0 , \1403_A[7]_b0 , w_2165 );
and ( w_2164 , w_2165 , \892_B[0]_b0 );
or ( \1405_b1 , \1293_A[6]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_2166 );
and ( \1405_b0 , \1293_A[6]_b0 , w_2167 );
and ( w_2166 , w_2167 , \929_B[1]_b0 );
or ( \1406_b1 , \1404_b1 , \1405_b1 );
xor ( \1406_b0 , \1404_b0 , w_2168 );
not ( w_2168 , w_2169 );
and ( w_2169 , \1405_b1 , \1405_b0 );
or ( \1407_b1 , \1294_b1 , \1295_b1 );
not ( \1295_b1 , w_2170 );
and ( \1407_b0 , \1294_b0 , w_2171 );
and ( w_2170 , w_2171 , \1295_b0 );
or ( \1408_b1 , \1296_b1 , \1299_b1 );
not ( \1299_b1 , w_2172 );
and ( \1408_b0 , \1296_b0 , w_2173 );
and ( w_2172 , w_2173 , \1299_b0 );
or ( \1409_b1 , \1407_b1 , w_2174 );
or ( \1409_b0 , \1407_b0 , \1408_b0 );
not ( \1408_b0 , w_2175 );
and ( w_2175 , w_2174 , \1408_b1 );
or ( \1410_b1 , \1406_b1 , \1409_b1 );
xor ( \1410_b0 , \1406_b0 , w_2176 );
not ( w_2176 , w_2177 );
and ( w_2177 , \1409_b1 , \1409_b0 );
or ( \1411_b1 , \1195_A[5]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_2178 );
and ( \1411_b0 , \1195_A[5]_b0 , w_2179 );
and ( w_2178 , w_2179 , \979_B[2]_b0 );
or ( \1412_b1 , \1410_b1 , \1411_b1 );
xor ( \1412_b0 , \1410_b0 , w_2180 );
not ( w_2180 , w_2181 );
and ( w_2181 , \1411_b1 , \1411_b0 );
or ( \1413_b1 , \1300_b1 , \1301_b1 );
not ( \1301_b1 , w_2182 );
and ( \1413_b0 , \1300_b0 , w_2183 );
and ( w_2182 , w_2183 , \1301_b0 );
or ( \1414_b1 , \1302_b1 , \1305_b1 );
not ( \1305_b1 , w_2184 );
and ( \1414_b0 , \1302_b0 , w_2185 );
and ( w_2184 , w_2185 , \1305_b0 );
or ( \1415_b1 , \1413_b1 , w_2186 );
or ( \1415_b0 , \1413_b0 , \1414_b0 );
not ( \1414_b0 , w_2187 );
and ( w_2187 , w_2186 , \1414_b1 );
or ( \1416_b1 , \1412_b1 , \1415_b1 );
xor ( \1416_b0 , \1412_b0 , w_2188 );
not ( w_2188 , w_2189 );
and ( w_2189 , \1415_b1 , \1415_b0 );
or ( \1417_b1 , \1109_A[4]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_2190 );
and ( \1417_b0 , \1109_A[4]_b0 , w_2191 );
and ( w_2190 , w_2191 , \1047_B[3]_b0 );
or ( \1418_b1 , \1416_b1 , \1417_b1 );
xor ( \1418_b0 , \1416_b0 , w_2192 );
not ( w_2192 , w_2193 );
and ( w_2193 , \1417_b1 , \1417_b0 );
or ( \1419_b1 , \1306_b1 , \1307_b1 );
not ( \1307_b1 , w_2194 );
and ( \1419_b0 , \1306_b0 , w_2195 );
and ( w_2194 , w_2195 , \1307_b0 );
or ( \1420_b1 , \1308_b1 , \1311_b1 );
not ( \1311_b1 , w_2196 );
and ( \1420_b0 , \1308_b0 , w_2197 );
and ( w_2196 , w_2197 , \1311_b0 );
or ( \1421_b1 , \1419_b1 , w_2198 );
or ( \1421_b0 , \1419_b0 , \1420_b0 );
not ( \1420_b0 , w_2199 );
and ( w_2199 , w_2198 , \1420_b1 );
or ( \1422_b1 , \1418_b1 , \1421_b1 );
xor ( \1422_b0 , \1418_b0 , w_2200 );
not ( w_2200 , w_2201 );
and ( w_2201 , \1421_b1 , \1421_b0 );
or ( \1423_b1 , \1035_A[3]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_2202 );
and ( \1423_b0 , \1035_A[3]_b0 , w_2203 );
and ( w_2202 , w_2203 , \1127_B[4]_b0 );
or ( \1424_b1 , \1422_b1 , \1423_b1 );
xor ( \1424_b0 , \1422_b0 , w_2204 );
not ( w_2204 , w_2205 );
and ( w_2205 , \1423_b1 , \1423_b0 );
or ( \1425_b1 , \1312_b1 , \1313_b1 );
not ( \1313_b1 , w_2206 );
and ( \1425_b0 , \1312_b0 , w_2207 );
and ( w_2206 , w_2207 , \1313_b0 );
or ( \1426_b1 , \1314_b1 , \1317_b1 );
not ( \1317_b1 , w_2208 );
and ( \1426_b0 , \1314_b0 , w_2209 );
and ( w_2208 , w_2209 , \1317_b0 );
or ( \1427_b1 , \1425_b1 , w_2210 );
or ( \1427_b0 , \1425_b0 , \1426_b0 );
not ( \1426_b0 , w_2211 );
and ( w_2211 , w_2210 , \1426_b1 );
or ( \1428_b1 , \1424_b1 , \1427_b1 );
xor ( \1428_b0 , \1424_b0 , w_2212 );
not ( w_2212 , w_2213 );
and ( w_2213 , \1427_b1 , \1427_b0 );
or ( \1429_b1 , \973_A[2]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_2214 );
and ( \1429_b0 , \973_A[2]_b0 , w_2215 );
and ( w_2214 , w_2215 , \1219_B[5]_b0 );
or ( \1430_b1 , \1428_b1 , \1429_b1 );
xor ( \1430_b0 , \1428_b0 , w_2216 );
not ( w_2216 , w_2217 );
and ( w_2217 , \1429_b1 , \1429_b0 );
or ( \1431_b1 , \1318_b1 , \1319_b1 );
not ( \1319_b1 , w_2218 );
and ( \1431_b0 , \1318_b0 , w_2219 );
and ( w_2218 , w_2219 , \1319_b0 );
or ( \1432_b1 , \1320_b1 , \1321_b1 );
not ( \1321_b1 , w_2220 );
and ( \1432_b0 , \1320_b0 , w_2221 );
and ( w_2220 , w_2221 , \1321_b0 );
or ( \1433_b1 , \1431_b1 , w_2222 );
or ( \1433_b0 , \1431_b0 , \1432_b0 );
not ( \1432_b0 , w_2223 );
and ( w_2223 , w_2222 , \1432_b1 );
or ( \1434_b1 , \1430_b1 , \1433_b1 );
xor ( \1434_b0 , \1430_b0 , w_2224 );
not ( w_2224 , w_2225 );
and ( w_2225 , \1433_b1 , \1433_b0 );
or ( \1435_b1 , \927_A[1]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_2226 );
and ( \1435_b0 , \927_A[1]_b0 , w_2227 );
and ( w_2226 , w_2227 , \1323_B[6]_b0 );
or ( \1436_b1 , \1434_b1 , \1435_b1 );
xor ( \1436_b0 , \1434_b0 , w_2228 );
not ( w_2228 , w_2229 );
and ( w_2229 , \1435_b1 , \1435_b0 );
or ( \1437_b1 , \1322_b1 , \1324_b1 );
not ( \1324_b1 , w_2230 );
and ( \1437_b0 , \1322_b0 , w_2231 );
and ( w_2230 , w_2231 , \1324_b0 );
or ( \1438_b1 , \1436_b1 , \1437_b1 );
xor ( \1438_b0 , \1436_b0 , w_2232 );
not ( w_2232 , w_2233 );
and ( w_2233 , \1437_b1 , \1437_b0 );
buf ( \1439_B[7]_b1 , \d[7]_b1 );
buf ( \1439_B[7]_b0 , \d[7]_b0 );
or ( \1440_b1 , \891_A[0]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_2234 );
and ( \1440_b0 , \891_A[0]_b0 , w_2235 );
and ( w_2234 , w_2235 , \1439_B[7]_b0 );
or ( \1441_b1 , \1438_b1 , \1440_b1 );
xor ( \1441_b0 , \1438_b0 , w_2236 );
not ( w_2236 , w_2237 );
and ( w_2237 , \1440_b1 , \1440_b0 );
buf ( \1442_Z[7]_b1 , \1441_b1 );
buf ( \1442_Z[7]_b0 , \1441_b0 );
or ( \1443_b1 , \1442_Z[7]_b1 , \865_b1 );
not ( \865_b1 , w_2238 );
and ( \1443_b0 , \1442_Z[7]_b0 , w_2239 );
and ( w_2238 , w_2239 , \865_b0 );
buf ( \1444_A[7]_b1 , \b[7]_b1 );
buf ( \1444_A[7]_b0 , \b[7]_b0 );
buf ( \1445_B[7]_b1 , \d[7]_b1 );
buf ( \1445_B[7]_b0 , \d[7]_b0 );
or ( \1446_b1 , \1444_A[7]_b1 , \1445_B[7]_b1 );
xor ( \1446_b0 , \1444_A[7]_b0 , w_2240 );
not ( w_2240 , w_2241 );
and ( w_2241 , \1445_B[7]_b1 , \1445_B[7]_b0 );
or ( \1447_b1 , \1328_A[6]_b1 , \1329_B[6]_b1 );
not ( \1329_B[6]_b1 , w_2242 );
and ( \1447_b0 , \1328_A[6]_b0 , w_2243 );
and ( w_2242 , w_2243 , \1329_B[6]_b0 );
or ( \1448_b1 , \1329_B[6]_b1 , \1334_b1 );
not ( \1334_b1 , w_2244 );
and ( \1448_b0 , \1329_B[6]_b0 , w_2245 );
and ( w_2244 , w_2245 , \1334_b0 );
or ( \1449_b1 , \1328_A[6]_b1 , \1334_b1 );
not ( \1334_b1 , w_2246 );
and ( \1449_b0 , \1328_A[6]_b0 , w_2247 );
and ( w_2246 , w_2247 , \1334_b0 );
or ( \1451_b1 , \1446_b1 , \1450_b1 );
xor ( \1451_b0 , \1446_b0 , w_2248 );
not ( w_2248 , w_2249 );
and ( w_2249 , \1450_b1 , \1450_b0 );
buf ( \1452_SUM[7]_b1 , \1451_b1 );
buf ( \1452_SUM[7]_b0 , \1451_b0 );
or ( \1453_b1 , \1452_SUM[7]_b1 , \863_b1 );
not ( \863_b1 , w_2250 );
and ( \1453_b0 , \1452_SUM[7]_b0 , w_2251 );
and ( w_2250 , w_2251 , \863_b0 );
buf ( \1454_A[7]_b1 , \a[7]_b1 );
buf ( \1454_A[7]_b0 , \a[7]_b0 );
buf ( \1455_B[7]_b1 , \c[7]_b1 );
buf ( \1455_B[7]_b0 , \c[7]_b0 );
or ( \1456_b1 , \1454_A[7]_b1 , \1455_B[7]_b1 );
xor ( \1456_b0 , \1454_A[7]_b0 , w_2252 );
not ( w_2252 , w_2253 );
and ( w_2253 , \1455_B[7]_b1 , \1455_B[7]_b0 );
or ( \1457_b1 , \1338_A[6]_b1 , \1339_B[6]_b1 );
not ( \1339_B[6]_b1 , w_2254 );
and ( \1457_b0 , \1338_A[6]_b0 , w_2255 );
and ( w_2254 , w_2255 , \1339_B[6]_b0 );
or ( \1458_b1 , \1339_B[6]_b1 , \1344_b1 );
not ( \1344_b1 , w_2256 );
and ( \1458_b0 , \1339_B[6]_b0 , w_2257 );
and ( w_2256 , w_2257 , \1344_b0 );
or ( \1459_b1 , \1338_A[6]_b1 , \1344_b1 );
not ( \1344_b1 , w_2258 );
and ( \1459_b0 , \1338_A[6]_b0 , w_2259 );
and ( w_2258 , w_2259 , \1344_b0 );
or ( \1461_b1 , \1456_b1 , \1460_b1 );
xor ( \1461_b0 , \1456_b0 , w_2260 );
not ( w_2260 , w_2261 );
and ( w_2261 , \1460_b1 , \1460_b0 );
buf ( \1462_SUM[7]_b1 , \1461_b1 );
buf ( \1462_SUM[7]_b0 , \1461_b0 );
or ( \1463_b1 , \1462_SUM[7]_b1 , \861_b1 );
not ( \861_b1 , w_2262 );
and ( \1463_b0 , \1462_SUM[7]_b0 , w_2263 );
and ( w_2262 , w_2263 , \861_b0 );
or ( \1464_b1 , \d[7]_b1 , \859_b1 );
not ( \859_b1 , w_2264 );
and ( \1464_b0 , \d[7]_b0 , w_2265 );
and ( w_2264 , w_2265 , \859_b0 );
or ( \1465_b1 , \c[7]_b1 , \857_b1 );
not ( \857_b1 , w_2266 );
and ( \1465_b0 , \c[7]_b0 , w_2267 );
and ( w_2266 , w_2267 , \857_b0 );
or ( \1466_b1 , \b[7]_b1 , \855_b1 );
not ( \855_b1 , w_2268 );
and ( \1466_b0 , \b[7]_b0 , w_2269 );
and ( w_2268 , w_2269 , \855_b0 );
or ( \1467_b1 , \a[7]_b1 , \853_b1 );
not ( \853_b1 , w_2270 );
and ( \1467_b0 , \a[7]_b0 , w_2271 );
and ( w_2270 , w_2271 , \853_b0 );
and ( \1469_b1 , 1'b0_b1 , w_2272 );
xor ( w_2272 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_2273 );
and ( \1469_b0 , w_2273 , \876_b0 );
or ( \1470_b1 , \a[8]_b1 , w_2274 );
or ( \1470_b0 , \a[8]_b0 , \d[8]_b0 );
not ( \d[8]_b0 , w_2275 );
and ( w_2275 , w_2274 , \d[8]_b1 );
or ( \1471_b1 , \1470_b1 , \875_b1 );
not ( \875_b1 , w_2276 );
and ( \1471_b0 , \1470_b0 , w_2277 );
and ( w_2276 , w_2277 , \875_b0 );
or ( \1472_b1 , \b[8]_b1 , \c[8]_b1 );
not ( \c[8]_b1 , w_2278 );
and ( \1472_b0 , \b[8]_b0 , w_2279 );
and ( w_2278 , w_2279 , \c[8]_b0 );
or ( \1473_b1 , \1472_b1 , \873_b1 );
not ( \873_b1 , w_2280 );
and ( \1473_b0 , \1472_b0 , w_2281 );
and ( w_2280 , w_2281 , \873_b0 );
or ( \1474_b1 , \a[8]_b1 , w_2282 );
or ( \1474_b0 , \a[8]_b0 , \b[8]_b0 );
not ( \b[8]_b0 , w_2283 );
and ( w_2283 , w_2282 , \b[8]_b1 );
or ( \1475_b1 , \1474_b1 , \871_b1 );
not ( \871_b1 , w_2284 );
and ( \1475_b0 , \1474_b0 , w_2285 );
and ( w_2284 , w_2285 , \871_b0 );
or ( \1476_b1 , \c[8]_b1 , \d[8]_b1 );
xor ( \1476_b0 , \c[8]_b0 , w_2286 );
not ( w_2286 , w_2287 );
and ( w_2287 , \d[8]_b1 , \d[8]_b0 );
or ( \1477_b1 , \1476_b1 , \869_b1 );
not ( \869_b1 , w_2288 );
and ( \1477_b0 , \1476_b0 , w_2289 );
and ( w_2288 , w_2289 , \869_b0 );
buf ( \1478_A[8]_b1 , \b[8]_b1 );
buf ( \1478_A[8]_b0 , \b[8]_b0 );
or ( \1479_b1 , \1478_A[8]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_2290 );
and ( \1479_b0 , \1478_A[8]_b0 , w_2291 );
and ( w_2290 , w_2291 , \887_B[0]_b0 );
or ( \1480_b1 , \1362_A[7]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_2292 );
and ( \1480_b0 , \1362_A[7]_b0 , w_2293 );
and ( w_2292 , w_2293 , \922_B[1]_b0 );
or ( \1481_b1 , \1479_b1 , \1480_b1 );
xor ( \1481_b0 , \1479_b0 , w_2294 );
not ( w_2294 , w_2295 );
and ( w_2295 , \1480_b1 , \1480_b0 );
or ( \1482_b1 , \1363_b1 , \1364_b1 );
not ( \1364_b1 , w_2296 );
and ( \1482_b0 , \1363_b0 , w_2297 );
and ( w_2296 , w_2297 , \1364_b0 );
or ( \1483_b1 , \1365_b1 , \1368_b1 );
not ( \1368_b1 , w_2298 );
and ( \1483_b0 , \1365_b0 , w_2299 );
and ( w_2298 , w_2299 , \1368_b0 );
or ( \1484_b1 , \1482_b1 , w_2300 );
or ( \1484_b0 , \1482_b0 , \1483_b0 );
not ( \1483_b0 , w_2301 );
and ( w_2301 , w_2300 , \1483_b1 );
or ( \1485_b1 , \1481_b1 , \1484_b1 );
xor ( \1485_b0 , \1481_b0 , w_2302 );
not ( w_2302 , w_2303 );
and ( w_2303 , \1484_b1 , \1484_b0 );
or ( \1486_b1 , \1258_A[6]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_2304 );
and ( \1486_b0 , \1258_A[6]_b0 , w_2305 );
and ( w_2304 , w_2305 , \968_B[2]_b0 );
or ( \1487_b1 , \1485_b1 , \1486_b1 );
xor ( \1487_b0 , \1485_b0 , w_2306 );
not ( w_2306 , w_2307 );
and ( w_2307 , \1486_b1 , \1486_b0 );
or ( \1488_b1 , \1369_b1 , \1370_b1 );
not ( \1370_b1 , w_2308 );
and ( \1488_b0 , \1369_b0 , w_2309 );
and ( w_2308 , w_2309 , \1370_b0 );
or ( \1489_b1 , \1371_b1 , \1374_b1 );
not ( \1374_b1 , w_2310 );
and ( \1489_b0 , \1371_b0 , w_2311 );
and ( w_2310 , w_2311 , \1374_b0 );
or ( \1490_b1 , \1488_b1 , w_2312 );
or ( \1490_b0 , \1488_b0 , \1489_b0 );
not ( \1489_b0 , w_2313 );
and ( w_2313 , w_2312 , \1489_b1 );
or ( \1491_b1 , \1487_b1 , \1490_b1 );
xor ( \1491_b0 , \1487_b0 , w_2314 );
not ( w_2314 , w_2315 );
and ( w_2315 , \1490_b1 , \1490_b0 );
or ( \1492_b1 , \1166_A[5]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_2316 );
and ( \1492_b0 , \1166_A[5]_b0 , w_2317 );
and ( w_2316 , w_2317 , \1030_B[3]_b0 );
or ( \1493_b1 , \1491_b1 , \1492_b1 );
xor ( \1493_b0 , \1491_b0 , w_2318 );
not ( w_2318 , w_2319 );
and ( w_2319 , \1492_b1 , \1492_b0 );
or ( \1494_b1 , \1375_b1 , \1376_b1 );
not ( \1376_b1 , w_2320 );
and ( \1494_b0 , \1375_b0 , w_2321 );
and ( w_2320 , w_2321 , \1376_b0 );
or ( \1495_b1 , \1377_b1 , \1380_b1 );
not ( \1380_b1 , w_2322 );
and ( \1495_b0 , \1377_b0 , w_2323 );
and ( w_2322 , w_2323 , \1380_b0 );
or ( \1496_b1 , \1494_b1 , w_2324 );
or ( \1496_b0 , \1494_b0 , \1495_b0 );
not ( \1495_b0 , w_2325 );
and ( w_2325 , w_2324 , \1495_b1 );
or ( \1497_b1 , \1493_b1 , \1496_b1 );
xor ( \1497_b0 , \1493_b0 , w_2326 );
not ( w_2326 , w_2327 );
and ( w_2327 , \1496_b1 , \1496_b0 );
or ( \1498_b1 , \1086_A[4]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_2328 );
and ( \1498_b0 , \1086_A[4]_b0 , w_2329 );
and ( w_2328 , w_2329 , \1104_B[4]_b0 );
or ( \1499_b1 , \1497_b1 , \1498_b1 );
xor ( \1499_b0 , \1497_b0 , w_2330 );
not ( w_2330 , w_2331 );
and ( w_2331 , \1498_b1 , \1498_b0 );
or ( \1500_b1 , \1381_b1 , \1382_b1 );
not ( \1382_b1 , w_2332 );
and ( \1500_b0 , \1381_b0 , w_2333 );
and ( w_2332 , w_2333 , \1382_b0 );
or ( \1501_b1 , \1383_b1 , \1386_b1 );
not ( \1386_b1 , w_2334 );
and ( \1501_b0 , \1383_b0 , w_2335 );
and ( w_2334 , w_2335 , \1386_b0 );
or ( \1502_b1 , \1500_b1 , w_2336 );
or ( \1502_b0 , \1500_b0 , \1501_b0 );
not ( \1501_b0 , w_2337 );
and ( w_2337 , w_2336 , \1501_b1 );
or ( \1503_b1 , \1499_b1 , \1502_b1 );
xor ( \1503_b0 , \1499_b0 , w_2338 );
not ( w_2338 , w_2339 );
and ( w_2339 , \1502_b1 , \1502_b0 );
or ( \1504_b1 , \1018_A[3]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_2340 );
and ( \1504_b0 , \1018_A[3]_b0 , w_2341 );
and ( w_2340 , w_2341 , \1190_B[5]_b0 );
or ( \1505_b1 , \1503_b1 , \1504_b1 );
xor ( \1505_b0 , \1503_b0 , w_2342 );
not ( w_2342 , w_2343 );
and ( w_2343 , \1504_b1 , \1504_b0 );
or ( \1506_b1 , \1387_b1 , \1388_b1 );
not ( \1388_b1 , w_2344 );
and ( \1506_b0 , \1387_b0 , w_2345 );
and ( w_2344 , w_2345 , \1388_b0 );
or ( \1507_b1 , \1389_b1 , \1392_b1 );
not ( \1392_b1 , w_2346 );
and ( \1507_b0 , \1389_b0 , w_2347 );
and ( w_2346 , w_2347 , \1392_b0 );
or ( \1508_b1 , \1506_b1 , w_2348 );
or ( \1508_b0 , \1506_b0 , \1507_b0 );
not ( \1507_b0 , w_2349 );
and ( w_2349 , w_2348 , \1507_b1 );
or ( \1509_b1 , \1505_b1 , \1508_b1 );
xor ( \1509_b0 , \1505_b0 , w_2350 );
not ( w_2350 , w_2351 );
and ( w_2351 , \1508_b1 , \1508_b0 );
or ( \1510_b1 , \962_A[2]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_2352 );
and ( \1510_b0 , \962_A[2]_b0 , w_2353 );
and ( w_2352 , w_2353 , \1288_B[6]_b0 );
or ( \1511_b1 , \1509_b1 , \1510_b1 );
xor ( \1511_b0 , \1509_b0 , w_2354 );
not ( w_2354 , w_2355 );
and ( w_2355 , \1510_b1 , \1510_b0 );
or ( \1512_b1 , \1393_b1 , \1394_b1 );
not ( \1394_b1 , w_2356 );
and ( \1512_b0 , \1393_b0 , w_2357 );
and ( w_2356 , w_2357 , \1394_b0 );
or ( \1513_b1 , \1395_b1 , \1396_b1 );
not ( \1396_b1 , w_2358 );
and ( \1513_b0 , \1395_b0 , w_2359 );
and ( w_2358 , w_2359 , \1396_b0 );
or ( \1514_b1 , \1512_b1 , w_2360 );
or ( \1514_b0 , \1512_b0 , \1513_b0 );
not ( \1513_b0 , w_2361 );
and ( w_2361 , w_2360 , \1513_b1 );
or ( \1515_b1 , \1511_b1 , \1514_b1 );
xor ( \1515_b0 , \1511_b0 , w_2362 );
not ( w_2362 , w_2363 );
and ( w_2363 , \1514_b1 , \1514_b0 );
or ( \1516_b1 , \920_A[1]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_2364 );
and ( \1516_b0 , \920_A[1]_b0 , w_2365 );
and ( w_2364 , w_2365 , \1398_B[7]_b0 );
or ( \1517_b1 , \1515_b1 , \1516_b1 );
xor ( \1517_b0 , \1515_b0 , w_2366 );
not ( w_2366 , w_2367 );
and ( w_2367 , \1516_b1 , \1516_b0 );
or ( \1518_b1 , \1397_b1 , \1399_b1 );
not ( \1399_b1 , w_2368 );
and ( \1518_b0 , \1397_b0 , w_2369 );
and ( w_2368 , w_2369 , \1399_b0 );
or ( \1519_b1 , \1517_b1 , \1518_b1 );
xor ( \1519_b0 , \1517_b0 , w_2370 );
not ( w_2370 , w_2371 );
and ( w_2371 , \1518_b1 , \1518_b0 );
buf ( \1520_B[8]_b1 , \c[8]_b1 );
buf ( \1520_B[8]_b0 , \c[8]_b0 );
or ( \1521_b1 , \886_A[0]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_2372 );
and ( \1521_b0 , \886_A[0]_b0 , w_2373 );
and ( w_2372 , w_2373 , \1520_B[8]_b0 );
or ( \1522_b1 , \1519_b1 , \1521_b1 );
xor ( \1522_b0 , \1519_b0 , w_2374 );
not ( w_2374 , w_2375 );
and ( w_2375 , \1521_b1 , \1521_b0 );
buf ( \1523_Z[8]_b1 , \1522_b1 );
buf ( \1523_Z[8]_b0 , \1522_b0 );
or ( \1524_b1 , \1523_Z[8]_b1 , \867_b1 );
not ( \867_b1 , w_2376 );
and ( \1524_b0 , \1523_Z[8]_b0 , w_2377 );
and ( w_2376 , w_2377 , \867_b0 );
buf ( \1525_A[8]_b1 , \a[8]_b1 );
buf ( \1525_A[8]_b0 , \a[8]_b0 );
or ( \1526_b1 , \1525_A[8]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_2378 );
and ( \1526_b0 , \1525_A[8]_b0 , w_2379 );
and ( w_2378 , w_2379 , \892_B[0]_b0 );
or ( \1527_b1 , \1403_A[7]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_2380 );
and ( \1527_b0 , \1403_A[7]_b0 , w_2381 );
and ( w_2380 , w_2381 , \929_B[1]_b0 );
or ( \1528_b1 , \1526_b1 , \1527_b1 );
xor ( \1528_b0 , \1526_b0 , w_2382 );
not ( w_2382 , w_2383 );
and ( w_2383 , \1527_b1 , \1527_b0 );
or ( \1529_b1 , \1404_b1 , \1405_b1 );
not ( \1405_b1 , w_2384 );
and ( \1529_b0 , \1404_b0 , w_2385 );
and ( w_2384 , w_2385 , \1405_b0 );
or ( \1530_b1 , \1406_b1 , \1409_b1 );
not ( \1409_b1 , w_2386 );
and ( \1530_b0 , \1406_b0 , w_2387 );
and ( w_2386 , w_2387 , \1409_b0 );
or ( \1531_b1 , \1529_b1 , w_2388 );
or ( \1531_b0 , \1529_b0 , \1530_b0 );
not ( \1530_b0 , w_2389 );
and ( w_2389 , w_2388 , \1530_b1 );
or ( \1532_b1 , \1528_b1 , \1531_b1 );
xor ( \1532_b0 , \1528_b0 , w_2390 );
not ( w_2390 , w_2391 );
and ( w_2391 , \1531_b1 , \1531_b0 );
or ( \1533_b1 , \1293_A[6]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_2392 );
and ( \1533_b0 , \1293_A[6]_b0 , w_2393 );
and ( w_2392 , w_2393 , \979_B[2]_b0 );
or ( \1534_b1 , \1532_b1 , \1533_b1 );
xor ( \1534_b0 , \1532_b0 , w_2394 );
not ( w_2394 , w_2395 );
and ( w_2395 , \1533_b1 , \1533_b0 );
or ( \1535_b1 , \1410_b1 , \1411_b1 );
not ( \1411_b1 , w_2396 );
and ( \1535_b0 , \1410_b0 , w_2397 );
and ( w_2396 , w_2397 , \1411_b0 );
or ( \1536_b1 , \1412_b1 , \1415_b1 );
not ( \1415_b1 , w_2398 );
and ( \1536_b0 , \1412_b0 , w_2399 );
and ( w_2398 , w_2399 , \1415_b0 );
or ( \1537_b1 , \1535_b1 , w_2400 );
or ( \1537_b0 , \1535_b0 , \1536_b0 );
not ( \1536_b0 , w_2401 );
and ( w_2401 , w_2400 , \1536_b1 );
or ( \1538_b1 , \1534_b1 , \1537_b1 );
xor ( \1538_b0 , \1534_b0 , w_2402 );
not ( w_2402 , w_2403 );
and ( w_2403 , \1537_b1 , \1537_b0 );
or ( \1539_b1 , \1195_A[5]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_2404 );
and ( \1539_b0 , \1195_A[5]_b0 , w_2405 );
and ( w_2404 , w_2405 , \1047_B[3]_b0 );
or ( \1540_b1 , \1538_b1 , \1539_b1 );
xor ( \1540_b0 , \1538_b0 , w_2406 );
not ( w_2406 , w_2407 );
and ( w_2407 , \1539_b1 , \1539_b0 );
or ( \1541_b1 , \1416_b1 , \1417_b1 );
not ( \1417_b1 , w_2408 );
and ( \1541_b0 , \1416_b0 , w_2409 );
and ( w_2408 , w_2409 , \1417_b0 );
or ( \1542_b1 , \1418_b1 , \1421_b1 );
not ( \1421_b1 , w_2410 );
and ( \1542_b0 , \1418_b0 , w_2411 );
and ( w_2410 , w_2411 , \1421_b0 );
or ( \1543_b1 , \1541_b1 , w_2412 );
or ( \1543_b0 , \1541_b0 , \1542_b0 );
not ( \1542_b0 , w_2413 );
and ( w_2413 , w_2412 , \1542_b1 );
or ( \1544_b1 , \1540_b1 , \1543_b1 );
xor ( \1544_b0 , \1540_b0 , w_2414 );
not ( w_2414 , w_2415 );
and ( w_2415 , \1543_b1 , \1543_b0 );
or ( \1545_b1 , \1109_A[4]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_2416 );
and ( \1545_b0 , \1109_A[4]_b0 , w_2417 );
and ( w_2416 , w_2417 , \1127_B[4]_b0 );
or ( \1546_b1 , \1544_b1 , \1545_b1 );
xor ( \1546_b0 , \1544_b0 , w_2418 );
not ( w_2418 , w_2419 );
and ( w_2419 , \1545_b1 , \1545_b0 );
or ( \1547_b1 , \1422_b1 , \1423_b1 );
not ( \1423_b1 , w_2420 );
and ( \1547_b0 , \1422_b0 , w_2421 );
and ( w_2420 , w_2421 , \1423_b0 );
or ( \1548_b1 , \1424_b1 , \1427_b1 );
not ( \1427_b1 , w_2422 );
and ( \1548_b0 , \1424_b0 , w_2423 );
and ( w_2422 , w_2423 , \1427_b0 );
or ( \1549_b1 , \1547_b1 , w_2424 );
or ( \1549_b0 , \1547_b0 , \1548_b0 );
not ( \1548_b0 , w_2425 );
and ( w_2425 , w_2424 , \1548_b1 );
or ( \1550_b1 , \1546_b1 , \1549_b1 );
xor ( \1550_b0 , \1546_b0 , w_2426 );
not ( w_2426 , w_2427 );
and ( w_2427 , \1549_b1 , \1549_b0 );
or ( \1551_b1 , \1035_A[3]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_2428 );
and ( \1551_b0 , \1035_A[3]_b0 , w_2429 );
and ( w_2428 , w_2429 , \1219_B[5]_b0 );
or ( \1552_b1 , \1550_b1 , \1551_b1 );
xor ( \1552_b0 , \1550_b0 , w_2430 );
not ( w_2430 , w_2431 );
and ( w_2431 , \1551_b1 , \1551_b0 );
or ( \1553_b1 , \1428_b1 , \1429_b1 );
not ( \1429_b1 , w_2432 );
and ( \1553_b0 , \1428_b0 , w_2433 );
and ( w_2432 , w_2433 , \1429_b0 );
or ( \1554_b1 , \1430_b1 , \1433_b1 );
not ( \1433_b1 , w_2434 );
and ( \1554_b0 , \1430_b0 , w_2435 );
and ( w_2434 , w_2435 , \1433_b0 );
or ( \1555_b1 , \1553_b1 , w_2436 );
or ( \1555_b0 , \1553_b0 , \1554_b0 );
not ( \1554_b0 , w_2437 );
and ( w_2437 , w_2436 , \1554_b1 );
or ( \1556_b1 , \1552_b1 , \1555_b1 );
xor ( \1556_b0 , \1552_b0 , w_2438 );
not ( w_2438 , w_2439 );
and ( w_2439 , \1555_b1 , \1555_b0 );
or ( \1557_b1 , \973_A[2]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_2440 );
and ( \1557_b0 , \973_A[2]_b0 , w_2441 );
and ( w_2440 , w_2441 , \1323_B[6]_b0 );
or ( \1558_b1 , \1556_b1 , \1557_b1 );
xor ( \1558_b0 , \1556_b0 , w_2442 );
not ( w_2442 , w_2443 );
and ( w_2443 , \1557_b1 , \1557_b0 );
or ( \1559_b1 , \1434_b1 , \1435_b1 );
not ( \1435_b1 , w_2444 );
and ( \1559_b0 , \1434_b0 , w_2445 );
and ( w_2444 , w_2445 , \1435_b0 );
or ( \1560_b1 , \1436_b1 , \1437_b1 );
not ( \1437_b1 , w_2446 );
and ( \1560_b0 , \1436_b0 , w_2447 );
and ( w_2446 , w_2447 , \1437_b0 );
or ( \1561_b1 , \1559_b1 , w_2448 );
or ( \1561_b0 , \1559_b0 , \1560_b0 );
not ( \1560_b0 , w_2449 );
and ( w_2449 , w_2448 , \1560_b1 );
or ( \1562_b1 , \1558_b1 , \1561_b1 );
xor ( \1562_b0 , \1558_b0 , w_2450 );
not ( w_2450 , w_2451 );
and ( w_2451 , \1561_b1 , \1561_b0 );
or ( \1563_b1 , \927_A[1]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_2452 );
and ( \1563_b0 , \927_A[1]_b0 , w_2453 );
and ( w_2452 , w_2453 , \1439_B[7]_b0 );
or ( \1564_b1 , \1562_b1 , \1563_b1 );
xor ( \1564_b0 , \1562_b0 , w_2454 );
not ( w_2454 , w_2455 );
and ( w_2455 , \1563_b1 , \1563_b0 );
or ( \1565_b1 , \1438_b1 , \1440_b1 );
not ( \1440_b1 , w_2456 );
and ( \1565_b0 , \1438_b0 , w_2457 );
and ( w_2456 , w_2457 , \1440_b0 );
or ( \1566_b1 , \1564_b1 , \1565_b1 );
xor ( \1566_b0 , \1564_b0 , w_2458 );
not ( w_2458 , w_2459 );
and ( w_2459 , \1565_b1 , \1565_b0 );
buf ( \1567_B[8]_b1 , \d[8]_b1 );
buf ( \1567_B[8]_b0 , \d[8]_b0 );
or ( \1568_b1 , \891_A[0]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_2460 );
and ( \1568_b0 , \891_A[0]_b0 , w_2461 );
and ( w_2460 , w_2461 , \1567_B[8]_b0 );
or ( \1569_b1 , \1566_b1 , \1568_b1 );
xor ( \1569_b0 , \1566_b0 , w_2462 );
not ( w_2462 , w_2463 );
and ( w_2463 , \1568_b1 , \1568_b0 );
buf ( \1570_Z[8]_b1 , \1569_b1 );
buf ( \1570_Z[8]_b0 , \1569_b0 );
or ( \1571_b1 , \1570_Z[8]_b1 , \865_b1 );
not ( \865_b1 , w_2464 );
and ( \1571_b0 , \1570_Z[8]_b0 , w_2465 );
and ( w_2464 , w_2465 , \865_b0 );
buf ( \1572_A[8]_b1 , \b[8]_b1 );
buf ( \1572_A[8]_b0 , \b[8]_b0 );
buf ( \1573_B[8]_b1 , \d[8]_b1 );
buf ( \1573_B[8]_b0 , \d[8]_b0 );
or ( \1574_b1 , \1572_A[8]_b1 , \1573_B[8]_b1 );
xor ( \1574_b0 , \1572_A[8]_b0 , w_2466 );
not ( w_2466 , w_2467 );
and ( w_2467 , \1573_B[8]_b1 , \1573_B[8]_b0 );
or ( \1575_b1 , \1444_A[7]_b1 , \1445_B[7]_b1 );
not ( \1445_B[7]_b1 , w_2468 );
and ( \1575_b0 , \1444_A[7]_b0 , w_2469 );
and ( w_2468 , w_2469 , \1445_B[7]_b0 );
or ( \1576_b1 , \1445_B[7]_b1 , \1450_b1 );
not ( \1450_b1 , w_2470 );
and ( \1576_b0 , \1445_B[7]_b0 , w_2471 );
and ( w_2470 , w_2471 , \1450_b0 );
or ( \1577_b1 , \1444_A[7]_b1 , \1450_b1 );
not ( \1450_b1 , w_2472 );
and ( \1577_b0 , \1444_A[7]_b0 , w_2473 );
and ( w_2472 , w_2473 , \1450_b0 );
or ( \1579_b1 , \1574_b1 , \1578_b1 );
xor ( \1579_b0 , \1574_b0 , w_2474 );
not ( w_2474 , w_2475 );
and ( w_2475 , \1578_b1 , \1578_b0 );
buf ( \1580_SUM[8]_b1 , \1579_b1 );
buf ( \1580_SUM[8]_b0 , \1579_b0 );
or ( \1581_b1 , \1580_SUM[8]_b1 , \863_b1 );
not ( \863_b1 , w_2476 );
and ( \1581_b0 , \1580_SUM[8]_b0 , w_2477 );
and ( w_2476 , w_2477 , \863_b0 );
buf ( \1582_A[8]_b1 , \a[8]_b1 );
buf ( \1582_A[8]_b0 , \a[8]_b0 );
buf ( \1583_B[8]_b1 , \c[8]_b1 );
buf ( \1583_B[8]_b0 , \c[8]_b0 );
or ( \1584_b1 , \1582_A[8]_b1 , \1583_B[8]_b1 );
xor ( \1584_b0 , \1582_A[8]_b0 , w_2478 );
not ( w_2478 , w_2479 );
and ( w_2479 , \1583_B[8]_b1 , \1583_B[8]_b0 );
or ( \1585_b1 , \1454_A[7]_b1 , \1455_B[7]_b1 );
not ( \1455_B[7]_b1 , w_2480 );
and ( \1585_b0 , \1454_A[7]_b0 , w_2481 );
and ( w_2480 , w_2481 , \1455_B[7]_b0 );
or ( \1586_b1 , \1455_B[7]_b1 , \1460_b1 );
not ( \1460_b1 , w_2482 );
and ( \1586_b0 , \1455_B[7]_b0 , w_2483 );
and ( w_2482 , w_2483 , \1460_b0 );
or ( \1587_b1 , \1454_A[7]_b1 , \1460_b1 );
not ( \1460_b1 , w_2484 );
and ( \1587_b0 , \1454_A[7]_b0 , w_2485 );
and ( w_2484 , w_2485 , \1460_b0 );
or ( \1589_b1 , \1584_b1 , \1588_b1 );
xor ( \1589_b0 , \1584_b0 , w_2486 );
not ( w_2486 , w_2487 );
and ( w_2487 , \1588_b1 , \1588_b0 );
buf ( \1590_SUM[8]_b1 , \1589_b1 );
buf ( \1590_SUM[8]_b0 , \1589_b0 );
or ( \1591_b1 , \1590_SUM[8]_b1 , \861_b1 );
not ( \861_b1 , w_2488 );
and ( \1591_b0 , \1590_SUM[8]_b0 , w_2489 );
and ( w_2488 , w_2489 , \861_b0 );
or ( \1592_b1 , \d[8]_b1 , \859_b1 );
not ( \859_b1 , w_2490 );
and ( \1592_b0 , \d[8]_b0 , w_2491 );
and ( w_2490 , w_2491 , \859_b0 );
or ( \1593_b1 , \c[8]_b1 , \857_b1 );
not ( \857_b1 , w_2492 );
and ( \1593_b0 , \c[8]_b0 , w_2493 );
and ( w_2492 , w_2493 , \857_b0 );
or ( \1594_b1 , \b[8]_b1 , \855_b1 );
not ( \855_b1 , w_2494 );
and ( \1594_b0 , \b[8]_b0 , w_2495 );
and ( w_2494 , w_2495 , \855_b0 );
or ( \1595_b1 , \a[8]_b1 , \853_b1 );
not ( \853_b1 , w_2496 );
and ( \1595_b0 , \a[8]_b0 , w_2497 );
and ( w_2496 , w_2497 , \853_b0 );
and ( \1597_b1 , 1'b0_b1 , w_2498 );
xor ( w_2498 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_2499 );
and ( \1597_b0 , w_2499 , \876_b0 );
or ( \1598_b1 , \a[9]_b1 , w_2500 );
or ( \1598_b0 , \a[9]_b0 , \d[9]_b0 );
not ( \d[9]_b0 , w_2501 );
and ( w_2501 , w_2500 , \d[9]_b1 );
or ( \1599_b1 , \1598_b1 , \875_b1 );
not ( \875_b1 , w_2502 );
and ( \1599_b0 , \1598_b0 , w_2503 );
and ( w_2502 , w_2503 , \875_b0 );
or ( \1600_b1 , \b[9]_b1 , \c[9]_b1 );
not ( \c[9]_b1 , w_2504 );
and ( \1600_b0 , \b[9]_b0 , w_2505 );
and ( w_2504 , w_2505 , \c[9]_b0 );
or ( \1601_b1 , \1600_b1 , \873_b1 );
not ( \873_b1 , w_2506 );
and ( \1601_b0 , \1600_b0 , w_2507 );
and ( w_2506 , w_2507 , \873_b0 );
or ( \1602_b1 , \a[9]_b1 , w_2508 );
or ( \1602_b0 , \a[9]_b0 , \b[9]_b0 );
not ( \b[9]_b0 , w_2509 );
and ( w_2509 , w_2508 , \b[9]_b1 );
or ( \1603_b1 , \1602_b1 , \871_b1 );
not ( \871_b1 , w_2510 );
and ( \1603_b0 , \1602_b0 , w_2511 );
and ( w_2510 , w_2511 , \871_b0 );
or ( \1604_b1 , \c[9]_b1 , \d[9]_b1 );
xor ( \1604_b0 , \c[9]_b0 , w_2512 );
not ( w_2512 , w_2513 );
and ( w_2513 , \d[9]_b1 , \d[9]_b0 );
or ( \1605_b1 , \1604_b1 , \869_b1 );
not ( \869_b1 , w_2514 );
and ( \1605_b0 , \1604_b0 , w_2515 );
and ( w_2514 , w_2515 , \869_b0 );
buf ( \1606_A[9]_b1 , \b[9]_b1 );
buf ( \1606_A[9]_b0 , \b[9]_b0 );
or ( \1607_b1 , \1606_A[9]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_2516 );
and ( \1607_b0 , \1606_A[9]_b0 , w_2517 );
and ( w_2516 , w_2517 , \887_B[0]_b0 );
or ( \1608_b1 , \1478_A[8]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_2518 );
and ( \1608_b0 , \1478_A[8]_b0 , w_2519 );
and ( w_2518 , w_2519 , \922_B[1]_b0 );
or ( \1609_b1 , \1607_b1 , \1608_b1 );
xor ( \1609_b0 , \1607_b0 , w_2520 );
not ( w_2520 , w_2521 );
and ( w_2521 , \1608_b1 , \1608_b0 );
or ( \1610_b1 , \1479_b1 , \1480_b1 );
not ( \1480_b1 , w_2522 );
and ( \1610_b0 , \1479_b0 , w_2523 );
and ( w_2522 , w_2523 , \1480_b0 );
or ( \1611_b1 , \1481_b1 , \1484_b1 );
not ( \1484_b1 , w_2524 );
and ( \1611_b0 , \1481_b0 , w_2525 );
and ( w_2524 , w_2525 , \1484_b0 );
or ( \1612_b1 , \1610_b1 , w_2526 );
or ( \1612_b0 , \1610_b0 , \1611_b0 );
not ( \1611_b0 , w_2527 );
and ( w_2527 , w_2526 , \1611_b1 );
or ( \1613_b1 , \1609_b1 , \1612_b1 );
xor ( \1613_b0 , \1609_b0 , w_2528 );
not ( w_2528 , w_2529 );
and ( w_2529 , \1612_b1 , \1612_b0 );
or ( \1614_b1 , \1362_A[7]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_2530 );
and ( \1614_b0 , \1362_A[7]_b0 , w_2531 );
and ( w_2530 , w_2531 , \968_B[2]_b0 );
or ( \1615_b1 , \1613_b1 , \1614_b1 );
xor ( \1615_b0 , \1613_b0 , w_2532 );
not ( w_2532 , w_2533 );
and ( w_2533 , \1614_b1 , \1614_b0 );
or ( \1616_b1 , \1485_b1 , \1486_b1 );
not ( \1486_b1 , w_2534 );
and ( \1616_b0 , \1485_b0 , w_2535 );
and ( w_2534 , w_2535 , \1486_b0 );
or ( \1617_b1 , \1487_b1 , \1490_b1 );
not ( \1490_b1 , w_2536 );
and ( \1617_b0 , \1487_b0 , w_2537 );
and ( w_2536 , w_2537 , \1490_b0 );
or ( \1618_b1 , \1616_b1 , w_2538 );
or ( \1618_b0 , \1616_b0 , \1617_b0 );
not ( \1617_b0 , w_2539 );
and ( w_2539 , w_2538 , \1617_b1 );
or ( \1619_b1 , \1615_b1 , \1618_b1 );
xor ( \1619_b0 , \1615_b0 , w_2540 );
not ( w_2540 , w_2541 );
and ( w_2541 , \1618_b1 , \1618_b0 );
or ( \1620_b1 , \1258_A[6]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_2542 );
and ( \1620_b0 , \1258_A[6]_b0 , w_2543 );
and ( w_2542 , w_2543 , \1030_B[3]_b0 );
or ( \1621_b1 , \1619_b1 , \1620_b1 );
xor ( \1621_b0 , \1619_b0 , w_2544 );
not ( w_2544 , w_2545 );
and ( w_2545 , \1620_b1 , \1620_b0 );
or ( \1622_b1 , \1491_b1 , \1492_b1 );
not ( \1492_b1 , w_2546 );
and ( \1622_b0 , \1491_b0 , w_2547 );
and ( w_2546 , w_2547 , \1492_b0 );
or ( \1623_b1 , \1493_b1 , \1496_b1 );
not ( \1496_b1 , w_2548 );
and ( \1623_b0 , \1493_b0 , w_2549 );
and ( w_2548 , w_2549 , \1496_b0 );
or ( \1624_b1 , \1622_b1 , w_2550 );
or ( \1624_b0 , \1622_b0 , \1623_b0 );
not ( \1623_b0 , w_2551 );
and ( w_2551 , w_2550 , \1623_b1 );
or ( \1625_b1 , \1621_b1 , \1624_b1 );
xor ( \1625_b0 , \1621_b0 , w_2552 );
not ( w_2552 , w_2553 );
and ( w_2553 , \1624_b1 , \1624_b0 );
or ( \1626_b1 , \1166_A[5]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_2554 );
and ( \1626_b0 , \1166_A[5]_b0 , w_2555 );
and ( w_2554 , w_2555 , \1104_B[4]_b0 );
or ( \1627_b1 , \1625_b1 , \1626_b1 );
xor ( \1627_b0 , \1625_b0 , w_2556 );
not ( w_2556 , w_2557 );
and ( w_2557 , \1626_b1 , \1626_b0 );
or ( \1628_b1 , \1497_b1 , \1498_b1 );
not ( \1498_b1 , w_2558 );
and ( \1628_b0 , \1497_b0 , w_2559 );
and ( w_2558 , w_2559 , \1498_b0 );
or ( \1629_b1 , \1499_b1 , \1502_b1 );
not ( \1502_b1 , w_2560 );
and ( \1629_b0 , \1499_b0 , w_2561 );
and ( w_2560 , w_2561 , \1502_b0 );
or ( \1630_b1 , \1628_b1 , w_2562 );
or ( \1630_b0 , \1628_b0 , \1629_b0 );
not ( \1629_b0 , w_2563 );
and ( w_2563 , w_2562 , \1629_b1 );
or ( \1631_b1 , \1627_b1 , \1630_b1 );
xor ( \1631_b0 , \1627_b0 , w_2564 );
not ( w_2564 , w_2565 );
and ( w_2565 , \1630_b1 , \1630_b0 );
or ( \1632_b1 , \1086_A[4]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_2566 );
and ( \1632_b0 , \1086_A[4]_b0 , w_2567 );
and ( w_2566 , w_2567 , \1190_B[5]_b0 );
or ( \1633_b1 , \1631_b1 , \1632_b1 );
xor ( \1633_b0 , \1631_b0 , w_2568 );
not ( w_2568 , w_2569 );
and ( w_2569 , \1632_b1 , \1632_b0 );
or ( \1634_b1 , \1503_b1 , \1504_b1 );
not ( \1504_b1 , w_2570 );
and ( \1634_b0 , \1503_b0 , w_2571 );
and ( w_2570 , w_2571 , \1504_b0 );
or ( \1635_b1 , \1505_b1 , \1508_b1 );
not ( \1508_b1 , w_2572 );
and ( \1635_b0 , \1505_b0 , w_2573 );
and ( w_2572 , w_2573 , \1508_b0 );
or ( \1636_b1 , \1634_b1 , w_2574 );
or ( \1636_b0 , \1634_b0 , \1635_b0 );
not ( \1635_b0 , w_2575 );
and ( w_2575 , w_2574 , \1635_b1 );
or ( \1637_b1 , \1633_b1 , \1636_b1 );
xor ( \1637_b0 , \1633_b0 , w_2576 );
not ( w_2576 , w_2577 );
and ( w_2577 , \1636_b1 , \1636_b0 );
or ( \1638_b1 , \1018_A[3]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_2578 );
and ( \1638_b0 , \1018_A[3]_b0 , w_2579 );
and ( w_2578 , w_2579 , \1288_B[6]_b0 );
or ( \1639_b1 , \1637_b1 , \1638_b1 );
xor ( \1639_b0 , \1637_b0 , w_2580 );
not ( w_2580 , w_2581 );
and ( w_2581 , \1638_b1 , \1638_b0 );
or ( \1640_b1 , \1509_b1 , \1510_b1 );
not ( \1510_b1 , w_2582 );
and ( \1640_b0 , \1509_b0 , w_2583 );
and ( w_2582 , w_2583 , \1510_b0 );
or ( \1641_b1 , \1511_b1 , \1514_b1 );
not ( \1514_b1 , w_2584 );
and ( \1641_b0 , \1511_b0 , w_2585 );
and ( w_2584 , w_2585 , \1514_b0 );
or ( \1642_b1 , \1640_b1 , w_2586 );
or ( \1642_b0 , \1640_b0 , \1641_b0 );
not ( \1641_b0 , w_2587 );
and ( w_2587 , w_2586 , \1641_b1 );
or ( \1643_b1 , \1639_b1 , \1642_b1 );
xor ( \1643_b0 , \1639_b0 , w_2588 );
not ( w_2588 , w_2589 );
and ( w_2589 , \1642_b1 , \1642_b0 );
or ( \1644_b1 , \962_A[2]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_2590 );
and ( \1644_b0 , \962_A[2]_b0 , w_2591 );
and ( w_2590 , w_2591 , \1398_B[7]_b0 );
or ( \1645_b1 , \1643_b1 , \1644_b1 );
xor ( \1645_b0 , \1643_b0 , w_2592 );
not ( w_2592 , w_2593 );
and ( w_2593 , \1644_b1 , \1644_b0 );
or ( \1646_b1 , \1515_b1 , \1516_b1 );
not ( \1516_b1 , w_2594 );
and ( \1646_b0 , \1515_b0 , w_2595 );
and ( w_2594 , w_2595 , \1516_b0 );
or ( \1647_b1 , \1517_b1 , \1518_b1 );
not ( \1518_b1 , w_2596 );
and ( \1647_b0 , \1517_b0 , w_2597 );
and ( w_2596 , w_2597 , \1518_b0 );
or ( \1648_b1 , \1646_b1 , w_2598 );
or ( \1648_b0 , \1646_b0 , \1647_b0 );
not ( \1647_b0 , w_2599 );
and ( w_2599 , w_2598 , \1647_b1 );
or ( \1649_b1 , \1645_b1 , \1648_b1 );
xor ( \1649_b0 , \1645_b0 , w_2600 );
not ( w_2600 , w_2601 );
and ( w_2601 , \1648_b1 , \1648_b0 );
or ( \1650_b1 , \920_A[1]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_2602 );
and ( \1650_b0 , \920_A[1]_b0 , w_2603 );
and ( w_2602 , w_2603 , \1520_B[8]_b0 );
or ( \1651_b1 , \1649_b1 , \1650_b1 );
xor ( \1651_b0 , \1649_b0 , w_2604 );
not ( w_2604 , w_2605 );
and ( w_2605 , \1650_b1 , \1650_b0 );
or ( \1652_b1 , \1519_b1 , \1521_b1 );
not ( \1521_b1 , w_2606 );
and ( \1652_b0 , \1519_b0 , w_2607 );
and ( w_2606 , w_2607 , \1521_b0 );
or ( \1653_b1 , \1651_b1 , \1652_b1 );
xor ( \1653_b0 , \1651_b0 , w_2608 );
not ( w_2608 , w_2609 );
and ( w_2609 , \1652_b1 , \1652_b0 );
buf ( \1654_B[9]_b1 , \c[9]_b1 );
buf ( \1654_B[9]_b0 , \c[9]_b0 );
or ( \1655_b1 , \886_A[0]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_2610 );
and ( \1655_b0 , \886_A[0]_b0 , w_2611 );
and ( w_2610 , w_2611 , \1654_B[9]_b0 );
or ( \1656_b1 , \1653_b1 , \1655_b1 );
xor ( \1656_b0 , \1653_b0 , w_2612 );
not ( w_2612 , w_2613 );
and ( w_2613 , \1655_b1 , \1655_b0 );
buf ( \1657_Z[9]_b1 , \1656_b1 );
buf ( \1657_Z[9]_b0 , \1656_b0 );
or ( \1658_b1 , \1657_Z[9]_b1 , \867_b1 );
not ( \867_b1 , w_2614 );
and ( \1658_b0 , \1657_Z[9]_b0 , w_2615 );
and ( w_2614 , w_2615 , \867_b0 );
buf ( \1659_A[9]_b1 , \a[9]_b1 );
buf ( \1659_A[9]_b0 , \a[9]_b0 );
or ( \1660_b1 , \1659_A[9]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_2616 );
and ( \1660_b0 , \1659_A[9]_b0 , w_2617 );
and ( w_2616 , w_2617 , \892_B[0]_b0 );
or ( \1661_b1 , \1525_A[8]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_2618 );
and ( \1661_b0 , \1525_A[8]_b0 , w_2619 );
and ( w_2618 , w_2619 , \929_B[1]_b0 );
or ( \1662_b1 , \1660_b1 , \1661_b1 );
xor ( \1662_b0 , \1660_b0 , w_2620 );
not ( w_2620 , w_2621 );
and ( w_2621 , \1661_b1 , \1661_b0 );
or ( \1663_b1 , \1526_b1 , \1527_b1 );
not ( \1527_b1 , w_2622 );
and ( \1663_b0 , \1526_b0 , w_2623 );
and ( w_2622 , w_2623 , \1527_b0 );
or ( \1664_b1 , \1528_b1 , \1531_b1 );
not ( \1531_b1 , w_2624 );
and ( \1664_b0 , \1528_b0 , w_2625 );
and ( w_2624 , w_2625 , \1531_b0 );
or ( \1665_b1 , \1663_b1 , w_2626 );
or ( \1665_b0 , \1663_b0 , \1664_b0 );
not ( \1664_b0 , w_2627 );
and ( w_2627 , w_2626 , \1664_b1 );
or ( \1666_b1 , \1662_b1 , \1665_b1 );
xor ( \1666_b0 , \1662_b0 , w_2628 );
not ( w_2628 , w_2629 );
and ( w_2629 , \1665_b1 , \1665_b0 );
or ( \1667_b1 , \1403_A[7]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_2630 );
and ( \1667_b0 , \1403_A[7]_b0 , w_2631 );
and ( w_2630 , w_2631 , \979_B[2]_b0 );
or ( \1668_b1 , \1666_b1 , \1667_b1 );
xor ( \1668_b0 , \1666_b0 , w_2632 );
not ( w_2632 , w_2633 );
and ( w_2633 , \1667_b1 , \1667_b0 );
or ( \1669_b1 , \1532_b1 , \1533_b1 );
not ( \1533_b1 , w_2634 );
and ( \1669_b0 , \1532_b0 , w_2635 );
and ( w_2634 , w_2635 , \1533_b0 );
or ( \1670_b1 , \1534_b1 , \1537_b1 );
not ( \1537_b1 , w_2636 );
and ( \1670_b0 , \1534_b0 , w_2637 );
and ( w_2636 , w_2637 , \1537_b0 );
or ( \1671_b1 , \1669_b1 , w_2638 );
or ( \1671_b0 , \1669_b0 , \1670_b0 );
not ( \1670_b0 , w_2639 );
and ( w_2639 , w_2638 , \1670_b1 );
or ( \1672_b1 , \1668_b1 , \1671_b1 );
xor ( \1672_b0 , \1668_b0 , w_2640 );
not ( w_2640 , w_2641 );
and ( w_2641 , \1671_b1 , \1671_b0 );
or ( \1673_b1 , \1293_A[6]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_2642 );
and ( \1673_b0 , \1293_A[6]_b0 , w_2643 );
and ( w_2642 , w_2643 , \1047_B[3]_b0 );
or ( \1674_b1 , \1672_b1 , \1673_b1 );
xor ( \1674_b0 , \1672_b0 , w_2644 );
not ( w_2644 , w_2645 );
and ( w_2645 , \1673_b1 , \1673_b0 );
or ( \1675_b1 , \1538_b1 , \1539_b1 );
not ( \1539_b1 , w_2646 );
and ( \1675_b0 , \1538_b0 , w_2647 );
and ( w_2646 , w_2647 , \1539_b0 );
or ( \1676_b1 , \1540_b1 , \1543_b1 );
not ( \1543_b1 , w_2648 );
and ( \1676_b0 , \1540_b0 , w_2649 );
and ( w_2648 , w_2649 , \1543_b0 );
or ( \1677_b1 , \1675_b1 , w_2650 );
or ( \1677_b0 , \1675_b0 , \1676_b0 );
not ( \1676_b0 , w_2651 );
and ( w_2651 , w_2650 , \1676_b1 );
or ( \1678_b1 , \1674_b1 , \1677_b1 );
xor ( \1678_b0 , \1674_b0 , w_2652 );
not ( w_2652 , w_2653 );
and ( w_2653 , \1677_b1 , \1677_b0 );
or ( \1679_b1 , \1195_A[5]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_2654 );
and ( \1679_b0 , \1195_A[5]_b0 , w_2655 );
and ( w_2654 , w_2655 , \1127_B[4]_b0 );
or ( \1680_b1 , \1678_b1 , \1679_b1 );
xor ( \1680_b0 , \1678_b0 , w_2656 );
not ( w_2656 , w_2657 );
and ( w_2657 , \1679_b1 , \1679_b0 );
or ( \1681_b1 , \1544_b1 , \1545_b1 );
not ( \1545_b1 , w_2658 );
and ( \1681_b0 , \1544_b0 , w_2659 );
and ( w_2658 , w_2659 , \1545_b0 );
or ( \1682_b1 , \1546_b1 , \1549_b1 );
not ( \1549_b1 , w_2660 );
and ( \1682_b0 , \1546_b0 , w_2661 );
and ( w_2660 , w_2661 , \1549_b0 );
or ( \1683_b1 , \1681_b1 , w_2662 );
or ( \1683_b0 , \1681_b0 , \1682_b0 );
not ( \1682_b0 , w_2663 );
and ( w_2663 , w_2662 , \1682_b1 );
or ( \1684_b1 , \1680_b1 , \1683_b1 );
xor ( \1684_b0 , \1680_b0 , w_2664 );
not ( w_2664 , w_2665 );
and ( w_2665 , \1683_b1 , \1683_b0 );
or ( \1685_b1 , \1109_A[4]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_2666 );
and ( \1685_b0 , \1109_A[4]_b0 , w_2667 );
and ( w_2666 , w_2667 , \1219_B[5]_b0 );
or ( \1686_b1 , \1684_b1 , \1685_b1 );
xor ( \1686_b0 , \1684_b0 , w_2668 );
not ( w_2668 , w_2669 );
and ( w_2669 , \1685_b1 , \1685_b0 );
or ( \1687_b1 , \1550_b1 , \1551_b1 );
not ( \1551_b1 , w_2670 );
and ( \1687_b0 , \1550_b0 , w_2671 );
and ( w_2670 , w_2671 , \1551_b0 );
or ( \1688_b1 , \1552_b1 , \1555_b1 );
not ( \1555_b1 , w_2672 );
and ( \1688_b0 , \1552_b0 , w_2673 );
and ( w_2672 , w_2673 , \1555_b0 );
or ( \1689_b1 , \1687_b1 , w_2674 );
or ( \1689_b0 , \1687_b0 , \1688_b0 );
not ( \1688_b0 , w_2675 );
and ( w_2675 , w_2674 , \1688_b1 );
or ( \1690_b1 , \1686_b1 , \1689_b1 );
xor ( \1690_b0 , \1686_b0 , w_2676 );
not ( w_2676 , w_2677 );
and ( w_2677 , \1689_b1 , \1689_b0 );
or ( \1691_b1 , \1035_A[3]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_2678 );
and ( \1691_b0 , \1035_A[3]_b0 , w_2679 );
and ( w_2678 , w_2679 , \1323_B[6]_b0 );
or ( \1692_b1 , \1690_b1 , \1691_b1 );
xor ( \1692_b0 , \1690_b0 , w_2680 );
not ( w_2680 , w_2681 );
and ( w_2681 , \1691_b1 , \1691_b0 );
or ( \1693_b1 , \1556_b1 , \1557_b1 );
not ( \1557_b1 , w_2682 );
and ( \1693_b0 , \1556_b0 , w_2683 );
and ( w_2682 , w_2683 , \1557_b0 );
or ( \1694_b1 , \1558_b1 , \1561_b1 );
not ( \1561_b1 , w_2684 );
and ( \1694_b0 , \1558_b0 , w_2685 );
and ( w_2684 , w_2685 , \1561_b0 );
or ( \1695_b1 , \1693_b1 , w_2686 );
or ( \1695_b0 , \1693_b0 , \1694_b0 );
not ( \1694_b0 , w_2687 );
and ( w_2687 , w_2686 , \1694_b1 );
or ( \1696_b1 , \1692_b1 , \1695_b1 );
xor ( \1696_b0 , \1692_b0 , w_2688 );
not ( w_2688 , w_2689 );
and ( w_2689 , \1695_b1 , \1695_b0 );
or ( \1697_b1 , \973_A[2]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_2690 );
and ( \1697_b0 , \973_A[2]_b0 , w_2691 );
and ( w_2690 , w_2691 , \1439_B[7]_b0 );
or ( \1698_b1 , \1696_b1 , \1697_b1 );
xor ( \1698_b0 , \1696_b0 , w_2692 );
not ( w_2692 , w_2693 );
and ( w_2693 , \1697_b1 , \1697_b0 );
or ( \1699_b1 , \1562_b1 , \1563_b1 );
not ( \1563_b1 , w_2694 );
and ( \1699_b0 , \1562_b0 , w_2695 );
and ( w_2694 , w_2695 , \1563_b0 );
or ( \1700_b1 , \1564_b1 , \1565_b1 );
not ( \1565_b1 , w_2696 );
and ( \1700_b0 , \1564_b0 , w_2697 );
and ( w_2696 , w_2697 , \1565_b0 );
or ( \1701_b1 , \1699_b1 , w_2698 );
or ( \1701_b0 , \1699_b0 , \1700_b0 );
not ( \1700_b0 , w_2699 );
and ( w_2699 , w_2698 , \1700_b1 );
or ( \1702_b1 , \1698_b1 , \1701_b1 );
xor ( \1702_b0 , \1698_b0 , w_2700 );
not ( w_2700 , w_2701 );
and ( w_2701 , \1701_b1 , \1701_b0 );
or ( \1703_b1 , \927_A[1]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_2702 );
and ( \1703_b0 , \927_A[1]_b0 , w_2703 );
and ( w_2702 , w_2703 , \1567_B[8]_b0 );
or ( \1704_b1 , \1702_b1 , \1703_b1 );
xor ( \1704_b0 , \1702_b0 , w_2704 );
not ( w_2704 , w_2705 );
and ( w_2705 , \1703_b1 , \1703_b0 );
or ( \1705_b1 , \1566_b1 , \1568_b1 );
not ( \1568_b1 , w_2706 );
and ( \1705_b0 , \1566_b0 , w_2707 );
and ( w_2706 , w_2707 , \1568_b0 );
or ( \1706_b1 , \1704_b1 , \1705_b1 );
xor ( \1706_b0 , \1704_b0 , w_2708 );
not ( w_2708 , w_2709 );
and ( w_2709 , \1705_b1 , \1705_b0 );
buf ( \1707_B[9]_b1 , \d[9]_b1 );
buf ( \1707_B[9]_b0 , \d[9]_b0 );
or ( \1708_b1 , \891_A[0]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_2710 );
and ( \1708_b0 , \891_A[0]_b0 , w_2711 );
and ( w_2710 , w_2711 , \1707_B[9]_b0 );
or ( \1709_b1 , \1706_b1 , \1708_b1 );
xor ( \1709_b0 , \1706_b0 , w_2712 );
not ( w_2712 , w_2713 );
and ( w_2713 , \1708_b1 , \1708_b0 );
buf ( \1710_Z[9]_b1 , \1709_b1 );
buf ( \1710_Z[9]_b0 , \1709_b0 );
or ( \1711_b1 , \1710_Z[9]_b1 , \865_b1 );
not ( \865_b1 , w_2714 );
and ( \1711_b0 , \1710_Z[9]_b0 , w_2715 );
and ( w_2714 , w_2715 , \865_b0 );
buf ( \1712_A[9]_b1 , \b[9]_b1 );
buf ( \1712_A[9]_b0 , \b[9]_b0 );
buf ( \1713_B[9]_b1 , \d[9]_b1 );
buf ( \1713_B[9]_b0 , \d[9]_b0 );
or ( \1714_b1 , \1712_A[9]_b1 , \1713_B[9]_b1 );
xor ( \1714_b0 , \1712_A[9]_b0 , w_2716 );
not ( w_2716 , w_2717 );
and ( w_2717 , \1713_B[9]_b1 , \1713_B[9]_b0 );
or ( \1715_b1 , \1572_A[8]_b1 , \1573_B[8]_b1 );
not ( \1573_B[8]_b1 , w_2718 );
and ( \1715_b0 , \1572_A[8]_b0 , w_2719 );
and ( w_2718 , w_2719 , \1573_B[8]_b0 );
or ( \1716_b1 , \1573_B[8]_b1 , \1578_b1 );
not ( \1578_b1 , w_2720 );
and ( \1716_b0 , \1573_B[8]_b0 , w_2721 );
and ( w_2720 , w_2721 , \1578_b0 );
or ( \1717_b1 , \1572_A[8]_b1 , \1578_b1 );
not ( \1578_b1 , w_2722 );
and ( \1717_b0 , \1572_A[8]_b0 , w_2723 );
and ( w_2722 , w_2723 , \1578_b0 );
or ( \1719_b1 , \1714_b1 , \1718_b1 );
xor ( \1719_b0 , \1714_b0 , w_2724 );
not ( w_2724 , w_2725 );
and ( w_2725 , \1718_b1 , \1718_b0 );
buf ( \1720_SUM[9]_b1 , \1719_b1 );
buf ( \1720_SUM[9]_b0 , \1719_b0 );
or ( \1721_b1 , \1720_SUM[9]_b1 , \863_b1 );
not ( \863_b1 , w_2726 );
and ( \1721_b0 , \1720_SUM[9]_b0 , w_2727 );
and ( w_2726 , w_2727 , \863_b0 );
buf ( \1722_A[9]_b1 , \a[9]_b1 );
buf ( \1722_A[9]_b0 , \a[9]_b0 );
buf ( \1723_B[9]_b1 , \c[9]_b1 );
buf ( \1723_B[9]_b0 , \c[9]_b0 );
or ( \1724_b1 , \1722_A[9]_b1 , \1723_B[9]_b1 );
xor ( \1724_b0 , \1722_A[9]_b0 , w_2728 );
not ( w_2728 , w_2729 );
and ( w_2729 , \1723_B[9]_b1 , \1723_B[9]_b0 );
or ( \1725_b1 , \1582_A[8]_b1 , \1583_B[8]_b1 );
not ( \1583_B[8]_b1 , w_2730 );
and ( \1725_b0 , \1582_A[8]_b0 , w_2731 );
and ( w_2730 , w_2731 , \1583_B[8]_b0 );
or ( \1726_b1 , \1583_B[8]_b1 , \1588_b1 );
not ( \1588_b1 , w_2732 );
and ( \1726_b0 , \1583_B[8]_b0 , w_2733 );
and ( w_2732 , w_2733 , \1588_b0 );
or ( \1727_b1 , \1582_A[8]_b1 , \1588_b1 );
not ( \1588_b1 , w_2734 );
and ( \1727_b0 , \1582_A[8]_b0 , w_2735 );
and ( w_2734 , w_2735 , \1588_b0 );
or ( \1729_b1 , \1724_b1 , \1728_b1 );
xor ( \1729_b0 , \1724_b0 , w_2736 );
not ( w_2736 , w_2737 );
and ( w_2737 , \1728_b1 , \1728_b0 );
buf ( \1730_SUM[9]_b1 , \1729_b1 );
buf ( \1730_SUM[9]_b0 , \1729_b0 );
or ( \1731_b1 , \1730_SUM[9]_b1 , \861_b1 );
not ( \861_b1 , w_2738 );
and ( \1731_b0 , \1730_SUM[9]_b0 , w_2739 );
and ( w_2738 , w_2739 , \861_b0 );
or ( \1732_b1 , \d[9]_b1 , \859_b1 );
not ( \859_b1 , w_2740 );
and ( \1732_b0 , \d[9]_b0 , w_2741 );
and ( w_2740 , w_2741 , \859_b0 );
or ( \1733_b1 , \c[9]_b1 , \857_b1 );
not ( \857_b1 , w_2742 );
and ( \1733_b0 , \c[9]_b0 , w_2743 );
and ( w_2742 , w_2743 , \857_b0 );
or ( \1734_b1 , \b[9]_b1 , \855_b1 );
not ( \855_b1 , w_2744 );
and ( \1734_b0 , \b[9]_b0 , w_2745 );
and ( w_2744 , w_2745 , \855_b0 );
or ( \1735_b1 , \a[9]_b1 , \853_b1 );
not ( \853_b1 , w_2746 );
and ( \1735_b0 , \a[9]_b0 , w_2747 );
and ( w_2746 , w_2747 , \853_b0 );
and ( \1737_b1 , 1'b0_b1 , w_2748 );
xor ( w_2748 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_2749 );
and ( \1737_b0 , w_2749 , \876_b0 );
or ( \1738_b1 , \a[10]_b1 , w_2750 );
or ( \1738_b0 , \a[10]_b0 , \d[10]_b0 );
not ( \d[10]_b0 , w_2751 );
and ( w_2751 , w_2750 , \d[10]_b1 );
or ( \1739_b1 , \1738_b1 , \875_b1 );
not ( \875_b1 , w_2752 );
and ( \1739_b0 , \1738_b0 , w_2753 );
and ( w_2752 , w_2753 , \875_b0 );
or ( \1740_b1 , \b[10]_b1 , \c[10]_b1 );
not ( \c[10]_b1 , w_2754 );
and ( \1740_b0 , \b[10]_b0 , w_2755 );
and ( w_2754 , w_2755 , \c[10]_b0 );
or ( \1741_b1 , \1740_b1 , \873_b1 );
not ( \873_b1 , w_2756 );
and ( \1741_b0 , \1740_b0 , w_2757 );
and ( w_2756 , w_2757 , \873_b0 );
or ( \1742_b1 , \a[10]_b1 , w_2758 );
or ( \1742_b0 , \a[10]_b0 , \b[10]_b0 );
not ( \b[10]_b0 , w_2759 );
and ( w_2759 , w_2758 , \b[10]_b1 );
or ( \1743_b1 , \1742_b1 , \871_b1 );
not ( \871_b1 , w_2760 );
and ( \1743_b0 , \1742_b0 , w_2761 );
and ( w_2760 , w_2761 , \871_b0 );
or ( \1744_b1 , \c[10]_b1 , \d[10]_b1 );
xor ( \1744_b0 , \c[10]_b0 , w_2762 );
not ( w_2762 , w_2763 );
and ( w_2763 , \d[10]_b1 , \d[10]_b0 );
or ( \1745_b1 , \1744_b1 , \869_b1 );
not ( \869_b1 , w_2764 );
and ( \1745_b0 , \1744_b0 , w_2765 );
and ( w_2764 , w_2765 , \869_b0 );
buf ( \1746_A[10]_b1 , \b[10]_b1 );
buf ( \1746_A[10]_b0 , \b[10]_b0 );
or ( \1747_b1 , \1746_A[10]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_2766 );
and ( \1747_b0 , \1746_A[10]_b0 , w_2767 );
and ( w_2766 , w_2767 , \887_B[0]_b0 );
or ( \1748_b1 , \1606_A[9]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_2768 );
and ( \1748_b0 , \1606_A[9]_b0 , w_2769 );
and ( w_2768 , w_2769 , \922_B[1]_b0 );
or ( \1749_b1 , \1747_b1 , \1748_b1 );
xor ( \1749_b0 , \1747_b0 , w_2770 );
not ( w_2770 , w_2771 );
and ( w_2771 , \1748_b1 , \1748_b0 );
or ( \1750_b1 , \1607_b1 , \1608_b1 );
not ( \1608_b1 , w_2772 );
and ( \1750_b0 , \1607_b0 , w_2773 );
and ( w_2772 , w_2773 , \1608_b0 );
or ( \1751_b1 , \1609_b1 , \1612_b1 );
not ( \1612_b1 , w_2774 );
and ( \1751_b0 , \1609_b0 , w_2775 );
and ( w_2774 , w_2775 , \1612_b0 );
or ( \1752_b1 , \1750_b1 , w_2776 );
or ( \1752_b0 , \1750_b0 , \1751_b0 );
not ( \1751_b0 , w_2777 );
and ( w_2777 , w_2776 , \1751_b1 );
or ( \1753_b1 , \1749_b1 , \1752_b1 );
xor ( \1753_b0 , \1749_b0 , w_2778 );
not ( w_2778 , w_2779 );
and ( w_2779 , \1752_b1 , \1752_b0 );
or ( \1754_b1 , \1478_A[8]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_2780 );
and ( \1754_b0 , \1478_A[8]_b0 , w_2781 );
and ( w_2780 , w_2781 , \968_B[2]_b0 );
or ( \1755_b1 , \1753_b1 , \1754_b1 );
xor ( \1755_b0 , \1753_b0 , w_2782 );
not ( w_2782 , w_2783 );
and ( w_2783 , \1754_b1 , \1754_b0 );
or ( \1756_b1 , \1613_b1 , \1614_b1 );
not ( \1614_b1 , w_2784 );
and ( \1756_b0 , \1613_b0 , w_2785 );
and ( w_2784 , w_2785 , \1614_b0 );
or ( \1757_b1 , \1615_b1 , \1618_b1 );
not ( \1618_b1 , w_2786 );
and ( \1757_b0 , \1615_b0 , w_2787 );
and ( w_2786 , w_2787 , \1618_b0 );
or ( \1758_b1 , \1756_b1 , w_2788 );
or ( \1758_b0 , \1756_b0 , \1757_b0 );
not ( \1757_b0 , w_2789 );
and ( w_2789 , w_2788 , \1757_b1 );
or ( \1759_b1 , \1755_b1 , \1758_b1 );
xor ( \1759_b0 , \1755_b0 , w_2790 );
not ( w_2790 , w_2791 );
and ( w_2791 , \1758_b1 , \1758_b0 );
or ( \1760_b1 , \1362_A[7]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_2792 );
and ( \1760_b0 , \1362_A[7]_b0 , w_2793 );
and ( w_2792 , w_2793 , \1030_B[3]_b0 );
or ( \1761_b1 , \1759_b1 , \1760_b1 );
xor ( \1761_b0 , \1759_b0 , w_2794 );
not ( w_2794 , w_2795 );
and ( w_2795 , \1760_b1 , \1760_b0 );
or ( \1762_b1 , \1619_b1 , \1620_b1 );
not ( \1620_b1 , w_2796 );
and ( \1762_b0 , \1619_b0 , w_2797 );
and ( w_2796 , w_2797 , \1620_b0 );
or ( \1763_b1 , \1621_b1 , \1624_b1 );
not ( \1624_b1 , w_2798 );
and ( \1763_b0 , \1621_b0 , w_2799 );
and ( w_2798 , w_2799 , \1624_b0 );
or ( \1764_b1 , \1762_b1 , w_2800 );
or ( \1764_b0 , \1762_b0 , \1763_b0 );
not ( \1763_b0 , w_2801 );
and ( w_2801 , w_2800 , \1763_b1 );
or ( \1765_b1 , \1761_b1 , \1764_b1 );
xor ( \1765_b0 , \1761_b0 , w_2802 );
not ( w_2802 , w_2803 );
and ( w_2803 , \1764_b1 , \1764_b0 );
or ( \1766_b1 , \1258_A[6]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_2804 );
and ( \1766_b0 , \1258_A[6]_b0 , w_2805 );
and ( w_2804 , w_2805 , \1104_B[4]_b0 );
or ( \1767_b1 , \1765_b1 , \1766_b1 );
xor ( \1767_b0 , \1765_b0 , w_2806 );
not ( w_2806 , w_2807 );
and ( w_2807 , \1766_b1 , \1766_b0 );
or ( \1768_b1 , \1625_b1 , \1626_b1 );
not ( \1626_b1 , w_2808 );
and ( \1768_b0 , \1625_b0 , w_2809 );
and ( w_2808 , w_2809 , \1626_b0 );
or ( \1769_b1 , \1627_b1 , \1630_b1 );
not ( \1630_b1 , w_2810 );
and ( \1769_b0 , \1627_b0 , w_2811 );
and ( w_2810 , w_2811 , \1630_b0 );
or ( \1770_b1 , \1768_b1 , w_2812 );
or ( \1770_b0 , \1768_b0 , \1769_b0 );
not ( \1769_b0 , w_2813 );
and ( w_2813 , w_2812 , \1769_b1 );
or ( \1771_b1 , \1767_b1 , \1770_b1 );
xor ( \1771_b0 , \1767_b0 , w_2814 );
not ( w_2814 , w_2815 );
and ( w_2815 , \1770_b1 , \1770_b0 );
or ( \1772_b1 , \1166_A[5]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_2816 );
and ( \1772_b0 , \1166_A[5]_b0 , w_2817 );
and ( w_2816 , w_2817 , \1190_B[5]_b0 );
or ( \1773_b1 , \1771_b1 , \1772_b1 );
xor ( \1773_b0 , \1771_b0 , w_2818 );
not ( w_2818 , w_2819 );
and ( w_2819 , \1772_b1 , \1772_b0 );
or ( \1774_b1 , \1631_b1 , \1632_b1 );
not ( \1632_b1 , w_2820 );
and ( \1774_b0 , \1631_b0 , w_2821 );
and ( w_2820 , w_2821 , \1632_b0 );
or ( \1775_b1 , \1633_b1 , \1636_b1 );
not ( \1636_b1 , w_2822 );
and ( \1775_b0 , \1633_b0 , w_2823 );
and ( w_2822 , w_2823 , \1636_b0 );
or ( \1776_b1 , \1774_b1 , w_2824 );
or ( \1776_b0 , \1774_b0 , \1775_b0 );
not ( \1775_b0 , w_2825 );
and ( w_2825 , w_2824 , \1775_b1 );
or ( \1777_b1 , \1773_b1 , \1776_b1 );
xor ( \1777_b0 , \1773_b0 , w_2826 );
not ( w_2826 , w_2827 );
and ( w_2827 , \1776_b1 , \1776_b0 );
or ( \1778_b1 , \1086_A[4]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_2828 );
and ( \1778_b0 , \1086_A[4]_b0 , w_2829 );
and ( w_2828 , w_2829 , \1288_B[6]_b0 );
or ( \1779_b1 , \1777_b1 , \1778_b1 );
xor ( \1779_b0 , \1777_b0 , w_2830 );
not ( w_2830 , w_2831 );
and ( w_2831 , \1778_b1 , \1778_b0 );
or ( \1780_b1 , \1637_b1 , \1638_b1 );
not ( \1638_b1 , w_2832 );
and ( \1780_b0 , \1637_b0 , w_2833 );
and ( w_2832 , w_2833 , \1638_b0 );
or ( \1781_b1 , \1639_b1 , \1642_b1 );
not ( \1642_b1 , w_2834 );
and ( \1781_b0 , \1639_b0 , w_2835 );
and ( w_2834 , w_2835 , \1642_b0 );
or ( \1782_b1 , \1780_b1 , w_2836 );
or ( \1782_b0 , \1780_b0 , \1781_b0 );
not ( \1781_b0 , w_2837 );
and ( w_2837 , w_2836 , \1781_b1 );
or ( \1783_b1 , \1779_b1 , \1782_b1 );
xor ( \1783_b0 , \1779_b0 , w_2838 );
not ( w_2838 , w_2839 );
and ( w_2839 , \1782_b1 , \1782_b0 );
or ( \1784_b1 , \1018_A[3]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_2840 );
and ( \1784_b0 , \1018_A[3]_b0 , w_2841 );
and ( w_2840 , w_2841 , \1398_B[7]_b0 );
or ( \1785_b1 , \1783_b1 , \1784_b1 );
xor ( \1785_b0 , \1783_b0 , w_2842 );
not ( w_2842 , w_2843 );
and ( w_2843 , \1784_b1 , \1784_b0 );
or ( \1786_b1 , \1643_b1 , \1644_b1 );
not ( \1644_b1 , w_2844 );
and ( \1786_b0 , \1643_b0 , w_2845 );
and ( w_2844 , w_2845 , \1644_b0 );
or ( \1787_b1 , \1645_b1 , \1648_b1 );
not ( \1648_b1 , w_2846 );
and ( \1787_b0 , \1645_b0 , w_2847 );
and ( w_2846 , w_2847 , \1648_b0 );
or ( \1788_b1 , \1786_b1 , w_2848 );
or ( \1788_b0 , \1786_b0 , \1787_b0 );
not ( \1787_b0 , w_2849 );
and ( w_2849 , w_2848 , \1787_b1 );
or ( \1789_b1 , \1785_b1 , \1788_b1 );
xor ( \1789_b0 , \1785_b0 , w_2850 );
not ( w_2850 , w_2851 );
and ( w_2851 , \1788_b1 , \1788_b0 );
or ( \1790_b1 , \962_A[2]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_2852 );
and ( \1790_b0 , \962_A[2]_b0 , w_2853 );
and ( w_2852 , w_2853 , \1520_B[8]_b0 );
or ( \1791_b1 , \1789_b1 , \1790_b1 );
xor ( \1791_b0 , \1789_b0 , w_2854 );
not ( w_2854 , w_2855 );
and ( w_2855 , \1790_b1 , \1790_b0 );
or ( \1792_b1 , \1649_b1 , \1650_b1 );
not ( \1650_b1 , w_2856 );
and ( \1792_b0 , \1649_b0 , w_2857 );
and ( w_2856 , w_2857 , \1650_b0 );
or ( \1793_b1 , \1651_b1 , \1652_b1 );
not ( \1652_b1 , w_2858 );
and ( \1793_b0 , \1651_b0 , w_2859 );
and ( w_2858 , w_2859 , \1652_b0 );
or ( \1794_b1 , \1792_b1 , w_2860 );
or ( \1794_b0 , \1792_b0 , \1793_b0 );
not ( \1793_b0 , w_2861 );
and ( w_2861 , w_2860 , \1793_b1 );
or ( \1795_b1 , \1791_b1 , \1794_b1 );
xor ( \1795_b0 , \1791_b0 , w_2862 );
not ( w_2862 , w_2863 );
and ( w_2863 , \1794_b1 , \1794_b0 );
or ( \1796_b1 , \920_A[1]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_2864 );
and ( \1796_b0 , \920_A[1]_b0 , w_2865 );
and ( w_2864 , w_2865 , \1654_B[9]_b0 );
or ( \1797_b1 , \1795_b1 , \1796_b1 );
xor ( \1797_b0 , \1795_b0 , w_2866 );
not ( w_2866 , w_2867 );
and ( w_2867 , \1796_b1 , \1796_b0 );
or ( \1798_b1 , \1653_b1 , \1655_b1 );
not ( \1655_b1 , w_2868 );
and ( \1798_b0 , \1653_b0 , w_2869 );
and ( w_2868 , w_2869 , \1655_b0 );
or ( \1799_b1 , \1797_b1 , \1798_b1 );
xor ( \1799_b0 , \1797_b0 , w_2870 );
not ( w_2870 , w_2871 );
and ( w_2871 , \1798_b1 , \1798_b0 );
buf ( \1800_B[10]_b1 , \c[10]_b1 );
buf ( \1800_B[10]_b0 , \c[10]_b0 );
or ( \1801_b1 , \886_A[0]_b1 , \1800_B[10]_b1 );
not ( \1800_B[10]_b1 , w_2872 );
and ( \1801_b0 , \886_A[0]_b0 , w_2873 );
and ( w_2872 , w_2873 , \1800_B[10]_b0 );
or ( \1802_b1 , \1799_b1 , \1801_b1 );
xor ( \1802_b0 , \1799_b0 , w_2874 );
not ( w_2874 , w_2875 );
and ( w_2875 , \1801_b1 , \1801_b0 );
buf ( \1803_Z[10]_b1 , \1802_b1 );
buf ( \1803_Z[10]_b0 , \1802_b0 );
or ( \1804_b1 , \1803_Z[10]_b1 , \867_b1 );
not ( \867_b1 , w_2876 );
and ( \1804_b0 , \1803_Z[10]_b0 , w_2877 );
and ( w_2876 , w_2877 , \867_b0 );
buf ( \1805_A[10]_b1 , \a[10]_b1 );
buf ( \1805_A[10]_b0 , \a[10]_b0 );
or ( \1806_b1 , \1805_A[10]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_2878 );
and ( \1806_b0 , \1805_A[10]_b0 , w_2879 );
and ( w_2878 , w_2879 , \892_B[0]_b0 );
or ( \1807_b1 , \1659_A[9]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_2880 );
and ( \1807_b0 , \1659_A[9]_b0 , w_2881 );
and ( w_2880 , w_2881 , \929_B[1]_b0 );
or ( \1808_b1 , \1806_b1 , \1807_b1 );
xor ( \1808_b0 , \1806_b0 , w_2882 );
not ( w_2882 , w_2883 );
and ( w_2883 , \1807_b1 , \1807_b0 );
or ( \1809_b1 , \1660_b1 , \1661_b1 );
not ( \1661_b1 , w_2884 );
and ( \1809_b0 , \1660_b0 , w_2885 );
and ( w_2884 , w_2885 , \1661_b0 );
or ( \1810_b1 , \1662_b1 , \1665_b1 );
not ( \1665_b1 , w_2886 );
and ( \1810_b0 , \1662_b0 , w_2887 );
and ( w_2886 , w_2887 , \1665_b0 );
or ( \1811_b1 , \1809_b1 , w_2888 );
or ( \1811_b0 , \1809_b0 , \1810_b0 );
not ( \1810_b0 , w_2889 );
and ( w_2889 , w_2888 , \1810_b1 );
or ( \1812_b1 , \1808_b1 , \1811_b1 );
xor ( \1812_b0 , \1808_b0 , w_2890 );
not ( w_2890 , w_2891 );
and ( w_2891 , \1811_b1 , \1811_b0 );
or ( \1813_b1 , \1525_A[8]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_2892 );
and ( \1813_b0 , \1525_A[8]_b0 , w_2893 );
and ( w_2892 , w_2893 , \979_B[2]_b0 );
or ( \1814_b1 , \1812_b1 , \1813_b1 );
xor ( \1814_b0 , \1812_b0 , w_2894 );
not ( w_2894 , w_2895 );
and ( w_2895 , \1813_b1 , \1813_b0 );
or ( \1815_b1 , \1666_b1 , \1667_b1 );
not ( \1667_b1 , w_2896 );
and ( \1815_b0 , \1666_b0 , w_2897 );
and ( w_2896 , w_2897 , \1667_b0 );
or ( \1816_b1 , \1668_b1 , \1671_b1 );
not ( \1671_b1 , w_2898 );
and ( \1816_b0 , \1668_b0 , w_2899 );
and ( w_2898 , w_2899 , \1671_b0 );
or ( \1817_b1 , \1815_b1 , w_2900 );
or ( \1817_b0 , \1815_b0 , \1816_b0 );
not ( \1816_b0 , w_2901 );
and ( w_2901 , w_2900 , \1816_b1 );
or ( \1818_b1 , \1814_b1 , \1817_b1 );
xor ( \1818_b0 , \1814_b0 , w_2902 );
not ( w_2902 , w_2903 );
and ( w_2903 , \1817_b1 , \1817_b0 );
or ( \1819_b1 , \1403_A[7]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_2904 );
and ( \1819_b0 , \1403_A[7]_b0 , w_2905 );
and ( w_2904 , w_2905 , \1047_B[3]_b0 );
or ( \1820_b1 , \1818_b1 , \1819_b1 );
xor ( \1820_b0 , \1818_b0 , w_2906 );
not ( w_2906 , w_2907 );
and ( w_2907 , \1819_b1 , \1819_b0 );
or ( \1821_b1 , \1672_b1 , \1673_b1 );
not ( \1673_b1 , w_2908 );
and ( \1821_b0 , \1672_b0 , w_2909 );
and ( w_2908 , w_2909 , \1673_b0 );
or ( \1822_b1 , \1674_b1 , \1677_b1 );
not ( \1677_b1 , w_2910 );
and ( \1822_b0 , \1674_b0 , w_2911 );
and ( w_2910 , w_2911 , \1677_b0 );
or ( \1823_b1 , \1821_b1 , w_2912 );
or ( \1823_b0 , \1821_b0 , \1822_b0 );
not ( \1822_b0 , w_2913 );
and ( w_2913 , w_2912 , \1822_b1 );
or ( \1824_b1 , \1820_b1 , \1823_b1 );
xor ( \1824_b0 , \1820_b0 , w_2914 );
not ( w_2914 , w_2915 );
and ( w_2915 , \1823_b1 , \1823_b0 );
or ( \1825_b1 , \1293_A[6]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_2916 );
and ( \1825_b0 , \1293_A[6]_b0 , w_2917 );
and ( w_2916 , w_2917 , \1127_B[4]_b0 );
or ( \1826_b1 , \1824_b1 , \1825_b1 );
xor ( \1826_b0 , \1824_b0 , w_2918 );
not ( w_2918 , w_2919 );
and ( w_2919 , \1825_b1 , \1825_b0 );
or ( \1827_b1 , \1678_b1 , \1679_b1 );
not ( \1679_b1 , w_2920 );
and ( \1827_b0 , \1678_b0 , w_2921 );
and ( w_2920 , w_2921 , \1679_b0 );
or ( \1828_b1 , \1680_b1 , \1683_b1 );
not ( \1683_b1 , w_2922 );
and ( \1828_b0 , \1680_b0 , w_2923 );
and ( w_2922 , w_2923 , \1683_b0 );
or ( \1829_b1 , \1827_b1 , w_2924 );
or ( \1829_b0 , \1827_b0 , \1828_b0 );
not ( \1828_b0 , w_2925 );
and ( w_2925 , w_2924 , \1828_b1 );
or ( \1830_b1 , \1826_b1 , \1829_b1 );
xor ( \1830_b0 , \1826_b0 , w_2926 );
not ( w_2926 , w_2927 );
and ( w_2927 , \1829_b1 , \1829_b0 );
or ( \1831_b1 , \1195_A[5]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_2928 );
and ( \1831_b0 , \1195_A[5]_b0 , w_2929 );
and ( w_2928 , w_2929 , \1219_B[5]_b0 );
or ( \1832_b1 , \1830_b1 , \1831_b1 );
xor ( \1832_b0 , \1830_b0 , w_2930 );
not ( w_2930 , w_2931 );
and ( w_2931 , \1831_b1 , \1831_b0 );
or ( \1833_b1 , \1684_b1 , \1685_b1 );
not ( \1685_b1 , w_2932 );
and ( \1833_b0 , \1684_b0 , w_2933 );
and ( w_2932 , w_2933 , \1685_b0 );
or ( \1834_b1 , \1686_b1 , \1689_b1 );
not ( \1689_b1 , w_2934 );
and ( \1834_b0 , \1686_b0 , w_2935 );
and ( w_2934 , w_2935 , \1689_b0 );
or ( \1835_b1 , \1833_b1 , w_2936 );
or ( \1835_b0 , \1833_b0 , \1834_b0 );
not ( \1834_b0 , w_2937 );
and ( w_2937 , w_2936 , \1834_b1 );
or ( \1836_b1 , \1832_b1 , \1835_b1 );
xor ( \1836_b0 , \1832_b0 , w_2938 );
not ( w_2938 , w_2939 );
and ( w_2939 , \1835_b1 , \1835_b0 );
or ( \1837_b1 , \1109_A[4]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_2940 );
and ( \1837_b0 , \1109_A[4]_b0 , w_2941 );
and ( w_2940 , w_2941 , \1323_B[6]_b0 );
or ( \1838_b1 , \1836_b1 , \1837_b1 );
xor ( \1838_b0 , \1836_b0 , w_2942 );
not ( w_2942 , w_2943 );
and ( w_2943 , \1837_b1 , \1837_b0 );
or ( \1839_b1 , \1690_b1 , \1691_b1 );
not ( \1691_b1 , w_2944 );
and ( \1839_b0 , \1690_b0 , w_2945 );
and ( w_2944 , w_2945 , \1691_b0 );
or ( \1840_b1 , \1692_b1 , \1695_b1 );
not ( \1695_b1 , w_2946 );
and ( \1840_b0 , \1692_b0 , w_2947 );
and ( w_2946 , w_2947 , \1695_b0 );
or ( \1841_b1 , \1839_b1 , w_2948 );
or ( \1841_b0 , \1839_b0 , \1840_b0 );
not ( \1840_b0 , w_2949 );
and ( w_2949 , w_2948 , \1840_b1 );
or ( \1842_b1 , \1838_b1 , \1841_b1 );
xor ( \1842_b0 , \1838_b0 , w_2950 );
not ( w_2950 , w_2951 );
and ( w_2951 , \1841_b1 , \1841_b0 );
or ( \1843_b1 , \1035_A[3]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_2952 );
and ( \1843_b0 , \1035_A[3]_b0 , w_2953 );
and ( w_2952 , w_2953 , \1439_B[7]_b0 );
or ( \1844_b1 , \1842_b1 , \1843_b1 );
xor ( \1844_b0 , \1842_b0 , w_2954 );
not ( w_2954 , w_2955 );
and ( w_2955 , \1843_b1 , \1843_b0 );
or ( \1845_b1 , \1696_b1 , \1697_b1 );
not ( \1697_b1 , w_2956 );
and ( \1845_b0 , \1696_b0 , w_2957 );
and ( w_2956 , w_2957 , \1697_b0 );
or ( \1846_b1 , \1698_b1 , \1701_b1 );
not ( \1701_b1 , w_2958 );
and ( \1846_b0 , \1698_b0 , w_2959 );
and ( w_2958 , w_2959 , \1701_b0 );
or ( \1847_b1 , \1845_b1 , w_2960 );
or ( \1847_b0 , \1845_b0 , \1846_b0 );
not ( \1846_b0 , w_2961 );
and ( w_2961 , w_2960 , \1846_b1 );
or ( \1848_b1 , \1844_b1 , \1847_b1 );
xor ( \1848_b0 , \1844_b0 , w_2962 );
not ( w_2962 , w_2963 );
and ( w_2963 , \1847_b1 , \1847_b0 );
or ( \1849_b1 , \973_A[2]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_2964 );
and ( \1849_b0 , \973_A[2]_b0 , w_2965 );
and ( w_2964 , w_2965 , \1567_B[8]_b0 );
or ( \1850_b1 , \1848_b1 , \1849_b1 );
xor ( \1850_b0 , \1848_b0 , w_2966 );
not ( w_2966 , w_2967 );
and ( w_2967 , \1849_b1 , \1849_b0 );
or ( \1851_b1 , \1702_b1 , \1703_b1 );
not ( \1703_b1 , w_2968 );
and ( \1851_b0 , \1702_b0 , w_2969 );
and ( w_2968 , w_2969 , \1703_b0 );
or ( \1852_b1 , \1704_b1 , \1705_b1 );
not ( \1705_b1 , w_2970 );
and ( \1852_b0 , \1704_b0 , w_2971 );
and ( w_2970 , w_2971 , \1705_b0 );
or ( \1853_b1 , \1851_b1 , w_2972 );
or ( \1853_b0 , \1851_b0 , \1852_b0 );
not ( \1852_b0 , w_2973 );
and ( w_2973 , w_2972 , \1852_b1 );
or ( \1854_b1 , \1850_b1 , \1853_b1 );
xor ( \1854_b0 , \1850_b0 , w_2974 );
not ( w_2974 , w_2975 );
and ( w_2975 , \1853_b1 , \1853_b0 );
or ( \1855_b1 , \927_A[1]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_2976 );
and ( \1855_b0 , \927_A[1]_b0 , w_2977 );
and ( w_2976 , w_2977 , \1707_B[9]_b0 );
or ( \1856_b1 , \1854_b1 , \1855_b1 );
xor ( \1856_b0 , \1854_b0 , w_2978 );
not ( w_2978 , w_2979 );
and ( w_2979 , \1855_b1 , \1855_b0 );
or ( \1857_b1 , \1706_b1 , \1708_b1 );
not ( \1708_b1 , w_2980 );
and ( \1857_b0 , \1706_b0 , w_2981 );
and ( w_2980 , w_2981 , \1708_b0 );
or ( \1858_b1 , \1856_b1 , \1857_b1 );
xor ( \1858_b0 , \1856_b0 , w_2982 );
not ( w_2982 , w_2983 );
and ( w_2983 , \1857_b1 , \1857_b0 );
buf ( \1859_B[10]_b1 , \d[10]_b1 );
buf ( \1859_B[10]_b0 , \d[10]_b0 );
or ( \1860_b1 , \891_A[0]_b1 , \1859_B[10]_b1 );
not ( \1859_B[10]_b1 , w_2984 );
and ( \1860_b0 , \891_A[0]_b0 , w_2985 );
and ( w_2984 , w_2985 , \1859_B[10]_b0 );
or ( \1861_b1 , \1858_b1 , \1860_b1 );
xor ( \1861_b0 , \1858_b0 , w_2986 );
not ( w_2986 , w_2987 );
and ( w_2987 , \1860_b1 , \1860_b0 );
buf ( \1862_Z[10]_b1 , \1861_b1 );
buf ( \1862_Z[10]_b0 , \1861_b0 );
or ( \1863_b1 , \1862_Z[10]_b1 , \865_b1 );
not ( \865_b1 , w_2988 );
and ( \1863_b0 , \1862_Z[10]_b0 , w_2989 );
and ( w_2988 , w_2989 , \865_b0 );
buf ( \1864_A[10]_b1 , \b[10]_b1 );
buf ( \1864_A[10]_b0 , \b[10]_b0 );
buf ( \1865_B[10]_b1 , \d[10]_b1 );
buf ( \1865_B[10]_b0 , \d[10]_b0 );
or ( \1866_b1 , \1864_A[10]_b1 , \1865_B[10]_b1 );
xor ( \1866_b0 , \1864_A[10]_b0 , w_2990 );
not ( w_2990 , w_2991 );
and ( w_2991 , \1865_B[10]_b1 , \1865_B[10]_b0 );
or ( \1867_b1 , \1712_A[9]_b1 , \1713_B[9]_b1 );
not ( \1713_B[9]_b1 , w_2992 );
and ( \1867_b0 , \1712_A[9]_b0 , w_2993 );
and ( w_2992 , w_2993 , \1713_B[9]_b0 );
or ( \1868_b1 , \1713_B[9]_b1 , \1718_b1 );
not ( \1718_b1 , w_2994 );
and ( \1868_b0 , \1713_B[9]_b0 , w_2995 );
and ( w_2994 , w_2995 , \1718_b0 );
or ( \1869_b1 , \1712_A[9]_b1 , \1718_b1 );
not ( \1718_b1 , w_2996 );
and ( \1869_b0 , \1712_A[9]_b0 , w_2997 );
and ( w_2996 , w_2997 , \1718_b0 );
or ( \1871_b1 , \1866_b1 , \1870_b1 );
xor ( \1871_b0 , \1866_b0 , w_2998 );
not ( w_2998 , w_2999 );
and ( w_2999 , \1870_b1 , \1870_b0 );
buf ( \1872_SUM[10]_b1 , \1871_b1 );
buf ( \1872_SUM[10]_b0 , \1871_b0 );
or ( \1873_b1 , \1872_SUM[10]_b1 , \863_b1 );
not ( \863_b1 , w_3000 );
and ( \1873_b0 , \1872_SUM[10]_b0 , w_3001 );
and ( w_3000 , w_3001 , \863_b0 );
buf ( \1874_A[10]_b1 , \a[10]_b1 );
buf ( \1874_A[10]_b0 , \a[10]_b0 );
buf ( \1875_B[10]_b1 , \c[10]_b1 );
buf ( \1875_B[10]_b0 , \c[10]_b0 );
or ( \1876_b1 , \1874_A[10]_b1 , \1875_B[10]_b1 );
xor ( \1876_b0 , \1874_A[10]_b0 , w_3002 );
not ( w_3002 , w_3003 );
and ( w_3003 , \1875_B[10]_b1 , \1875_B[10]_b0 );
or ( \1877_b1 , \1722_A[9]_b1 , \1723_B[9]_b1 );
not ( \1723_B[9]_b1 , w_3004 );
and ( \1877_b0 , \1722_A[9]_b0 , w_3005 );
and ( w_3004 , w_3005 , \1723_B[9]_b0 );
or ( \1878_b1 , \1723_B[9]_b1 , \1728_b1 );
not ( \1728_b1 , w_3006 );
and ( \1878_b0 , \1723_B[9]_b0 , w_3007 );
and ( w_3006 , w_3007 , \1728_b0 );
or ( \1879_b1 , \1722_A[9]_b1 , \1728_b1 );
not ( \1728_b1 , w_3008 );
and ( \1879_b0 , \1722_A[9]_b0 , w_3009 );
and ( w_3008 , w_3009 , \1728_b0 );
or ( \1881_b1 , \1876_b1 , \1880_b1 );
xor ( \1881_b0 , \1876_b0 , w_3010 );
not ( w_3010 , w_3011 );
and ( w_3011 , \1880_b1 , \1880_b0 );
buf ( \1882_SUM[10]_b1 , \1881_b1 );
buf ( \1882_SUM[10]_b0 , \1881_b0 );
or ( \1883_b1 , \1882_SUM[10]_b1 , \861_b1 );
not ( \861_b1 , w_3012 );
and ( \1883_b0 , \1882_SUM[10]_b0 , w_3013 );
and ( w_3012 , w_3013 , \861_b0 );
or ( \1884_b1 , \d[10]_b1 , \859_b1 );
not ( \859_b1 , w_3014 );
and ( \1884_b0 , \d[10]_b0 , w_3015 );
and ( w_3014 , w_3015 , \859_b0 );
or ( \1885_b1 , \c[10]_b1 , \857_b1 );
not ( \857_b1 , w_3016 );
and ( \1885_b0 , \c[10]_b0 , w_3017 );
and ( w_3016 , w_3017 , \857_b0 );
or ( \1886_b1 , \b[10]_b1 , \855_b1 );
not ( \855_b1 , w_3018 );
and ( \1886_b0 , \b[10]_b0 , w_3019 );
and ( w_3018 , w_3019 , \855_b0 );
or ( \1887_b1 , \a[10]_b1 , \853_b1 );
not ( \853_b1 , w_3020 );
and ( \1887_b0 , \a[10]_b0 , w_3021 );
and ( w_3020 , w_3021 , \853_b0 );
and ( \1889_b1 , 1'b0_b1 , w_3022 );
xor ( w_3022 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_3023 );
and ( \1889_b0 , w_3023 , \876_b0 );
or ( \1890_b1 , \a[11]_b1 , w_3024 );
or ( \1890_b0 , \a[11]_b0 , \d[11]_b0 );
not ( \d[11]_b0 , w_3025 );
and ( w_3025 , w_3024 , \d[11]_b1 );
or ( \1891_b1 , \1890_b1 , \875_b1 );
not ( \875_b1 , w_3026 );
and ( \1891_b0 , \1890_b0 , w_3027 );
and ( w_3026 , w_3027 , \875_b0 );
or ( \1892_b1 , \b[11]_b1 , \c[11]_b1 );
not ( \c[11]_b1 , w_3028 );
and ( \1892_b0 , \b[11]_b0 , w_3029 );
and ( w_3028 , w_3029 , \c[11]_b0 );
or ( \1893_b1 , \1892_b1 , \873_b1 );
not ( \873_b1 , w_3030 );
and ( \1893_b0 , \1892_b0 , w_3031 );
and ( w_3030 , w_3031 , \873_b0 );
or ( \1894_b1 , \a[11]_b1 , w_3032 );
or ( \1894_b0 , \a[11]_b0 , \b[11]_b0 );
not ( \b[11]_b0 , w_3033 );
and ( w_3033 , w_3032 , \b[11]_b1 );
or ( \1895_b1 , \1894_b1 , \871_b1 );
not ( \871_b1 , w_3034 );
and ( \1895_b0 , \1894_b0 , w_3035 );
and ( w_3034 , w_3035 , \871_b0 );
or ( \1896_b1 , \c[11]_b1 , \d[11]_b1 );
xor ( \1896_b0 , \c[11]_b0 , w_3036 );
not ( w_3036 , w_3037 );
and ( w_3037 , \d[11]_b1 , \d[11]_b0 );
or ( \1897_b1 , \1896_b1 , \869_b1 );
not ( \869_b1 , w_3038 );
and ( \1897_b0 , \1896_b0 , w_3039 );
and ( w_3038 , w_3039 , \869_b0 );
buf ( \1898_A[11]_b1 , \b[11]_b1 );
buf ( \1898_A[11]_b0 , \b[11]_b0 );
or ( \1899_b1 , \1898_A[11]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_3040 );
and ( \1899_b0 , \1898_A[11]_b0 , w_3041 );
and ( w_3040 , w_3041 , \887_B[0]_b0 );
or ( \1900_b1 , \1746_A[10]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_3042 );
and ( \1900_b0 , \1746_A[10]_b0 , w_3043 );
and ( w_3042 , w_3043 , \922_B[1]_b0 );
or ( \1901_b1 , \1899_b1 , \1900_b1 );
xor ( \1901_b0 , \1899_b0 , w_3044 );
not ( w_3044 , w_3045 );
and ( w_3045 , \1900_b1 , \1900_b0 );
or ( \1902_b1 , \1747_b1 , \1748_b1 );
not ( \1748_b1 , w_3046 );
and ( \1902_b0 , \1747_b0 , w_3047 );
and ( w_3046 , w_3047 , \1748_b0 );
or ( \1903_b1 , \1749_b1 , \1752_b1 );
not ( \1752_b1 , w_3048 );
and ( \1903_b0 , \1749_b0 , w_3049 );
and ( w_3048 , w_3049 , \1752_b0 );
or ( \1904_b1 , \1902_b1 , w_3050 );
or ( \1904_b0 , \1902_b0 , \1903_b0 );
not ( \1903_b0 , w_3051 );
and ( w_3051 , w_3050 , \1903_b1 );
or ( \1905_b1 , \1901_b1 , \1904_b1 );
xor ( \1905_b0 , \1901_b0 , w_3052 );
not ( w_3052 , w_3053 );
and ( w_3053 , \1904_b1 , \1904_b0 );
or ( \1906_b1 , \1606_A[9]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_3054 );
and ( \1906_b0 , \1606_A[9]_b0 , w_3055 );
and ( w_3054 , w_3055 , \968_B[2]_b0 );
or ( \1907_b1 , \1905_b1 , \1906_b1 );
xor ( \1907_b0 , \1905_b0 , w_3056 );
not ( w_3056 , w_3057 );
and ( w_3057 , \1906_b1 , \1906_b0 );
or ( \1908_b1 , \1753_b1 , \1754_b1 );
not ( \1754_b1 , w_3058 );
and ( \1908_b0 , \1753_b0 , w_3059 );
and ( w_3058 , w_3059 , \1754_b0 );
or ( \1909_b1 , \1755_b1 , \1758_b1 );
not ( \1758_b1 , w_3060 );
and ( \1909_b0 , \1755_b0 , w_3061 );
and ( w_3060 , w_3061 , \1758_b0 );
or ( \1910_b1 , \1908_b1 , w_3062 );
or ( \1910_b0 , \1908_b0 , \1909_b0 );
not ( \1909_b0 , w_3063 );
and ( w_3063 , w_3062 , \1909_b1 );
or ( \1911_b1 , \1907_b1 , \1910_b1 );
xor ( \1911_b0 , \1907_b0 , w_3064 );
not ( w_3064 , w_3065 );
and ( w_3065 , \1910_b1 , \1910_b0 );
or ( \1912_b1 , \1478_A[8]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_3066 );
and ( \1912_b0 , \1478_A[8]_b0 , w_3067 );
and ( w_3066 , w_3067 , \1030_B[3]_b0 );
or ( \1913_b1 , \1911_b1 , \1912_b1 );
xor ( \1913_b0 , \1911_b0 , w_3068 );
not ( w_3068 , w_3069 );
and ( w_3069 , \1912_b1 , \1912_b0 );
or ( \1914_b1 , \1759_b1 , \1760_b1 );
not ( \1760_b1 , w_3070 );
and ( \1914_b0 , \1759_b0 , w_3071 );
and ( w_3070 , w_3071 , \1760_b0 );
or ( \1915_b1 , \1761_b1 , \1764_b1 );
not ( \1764_b1 , w_3072 );
and ( \1915_b0 , \1761_b0 , w_3073 );
and ( w_3072 , w_3073 , \1764_b0 );
or ( \1916_b1 , \1914_b1 , w_3074 );
or ( \1916_b0 , \1914_b0 , \1915_b0 );
not ( \1915_b0 , w_3075 );
and ( w_3075 , w_3074 , \1915_b1 );
or ( \1917_b1 , \1913_b1 , \1916_b1 );
xor ( \1917_b0 , \1913_b0 , w_3076 );
not ( w_3076 , w_3077 );
and ( w_3077 , \1916_b1 , \1916_b0 );
or ( \1918_b1 , \1362_A[7]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_3078 );
and ( \1918_b0 , \1362_A[7]_b0 , w_3079 );
and ( w_3078 , w_3079 , \1104_B[4]_b0 );
or ( \1919_b1 , \1917_b1 , \1918_b1 );
xor ( \1919_b0 , \1917_b0 , w_3080 );
not ( w_3080 , w_3081 );
and ( w_3081 , \1918_b1 , \1918_b0 );
or ( \1920_b1 , \1765_b1 , \1766_b1 );
not ( \1766_b1 , w_3082 );
and ( \1920_b0 , \1765_b0 , w_3083 );
and ( w_3082 , w_3083 , \1766_b0 );
or ( \1921_b1 , \1767_b1 , \1770_b1 );
not ( \1770_b1 , w_3084 );
and ( \1921_b0 , \1767_b0 , w_3085 );
and ( w_3084 , w_3085 , \1770_b0 );
or ( \1922_b1 , \1920_b1 , w_3086 );
or ( \1922_b0 , \1920_b0 , \1921_b0 );
not ( \1921_b0 , w_3087 );
and ( w_3087 , w_3086 , \1921_b1 );
or ( \1923_b1 , \1919_b1 , \1922_b1 );
xor ( \1923_b0 , \1919_b0 , w_3088 );
not ( w_3088 , w_3089 );
and ( w_3089 , \1922_b1 , \1922_b0 );
or ( \1924_b1 , \1258_A[6]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_3090 );
and ( \1924_b0 , \1258_A[6]_b0 , w_3091 );
and ( w_3090 , w_3091 , \1190_B[5]_b0 );
or ( \1925_b1 , \1923_b1 , \1924_b1 );
xor ( \1925_b0 , \1923_b0 , w_3092 );
not ( w_3092 , w_3093 );
and ( w_3093 , \1924_b1 , \1924_b0 );
or ( \1926_b1 , \1771_b1 , \1772_b1 );
not ( \1772_b1 , w_3094 );
and ( \1926_b0 , \1771_b0 , w_3095 );
and ( w_3094 , w_3095 , \1772_b0 );
or ( \1927_b1 , \1773_b1 , \1776_b1 );
not ( \1776_b1 , w_3096 );
and ( \1927_b0 , \1773_b0 , w_3097 );
and ( w_3096 , w_3097 , \1776_b0 );
or ( \1928_b1 , \1926_b1 , w_3098 );
or ( \1928_b0 , \1926_b0 , \1927_b0 );
not ( \1927_b0 , w_3099 );
and ( w_3099 , w_3098 , \1927_b1 );
or ( \1929_b1 , \1925_b1 , \1928_b1 );
xor ( \1929_b0 , \1925_b0 , w_3100 );
not ( w_3100 , w_3101 );
and ( w_3101 , \1928_b1 , \1928_b0 );
or ( \1930_b1 , \1166_A[5]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_3102 );
and ( \1930_b0 , \1166_A[5]_b0 , w_3103 );
and ( w_3102 , w_3103 , \1288_B[6]_b0 );
or ( \1931_b1 , \1929_b1 , \1930_b1 );
xor ( \1931_b0 , \1929_b0 , w_3104 );
not ( w_3104 , w_3105 );
and ( w_3105 , \1930_b1 , \1930_b0 );
or ( \1932_b1 , \1777_b1 , \1778_b1 );
not ( \1778_b1 , w_3106 );
and ( \1932_b0 , \1777_b0 , w_3107 );
and ( w_3106 , w_3107 , \1778_b0 );
or ( \1933_b1 , \1779_b1 , \1782_b1 );
not ( \1782_b1 , w_3108 );
and ( \1933_b0 , \1779_b0 , w_3109 );
and ( w_3108 , w_3109 , \1782_b0 );
or ( \1934_b1 , \1932_b1 , w_3110 );
or ( \1934_b0 , \1932_b0 , \1933_b0 );
not ( \1933_b0 , w_3111 );
and ( w_3111 , w_3110 , \1933_b1 );
or ( \1935_b1 , \1931_b1 , \1934_b1 );
xor ( \1935_b0 , \1931_b0 , w_3112 );
not ( w_3112 , w_3113 );
and ( w_3113 , \1934_b1 , \1934_b0 );
or ( \1936_b1 , \1086_A[4]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_3114 );
and ( \1936_b0 , \1086_A[4]_b0 , w_3115 );
and ( w_3114 , w_3115 , \1398_B[7]_b0 );
or ( \1937_b1 , \1935_b1 , \1936_b1 );
xor ( \1937_b0 , \1935_b0 , w_3116 );
not ( w_3116 , w_3117 );
and ( w_3117 , \1936_b1 , \1936_b0 );
or ( \1938_b1 , \1783_b1 , \1784_b1 );
not ( \1784_b1 , w_3118 );
and ( \1938_b0 , \1783_b0 , w_3119 );
and ( w_3118 , w_3119 , \1784_b0 );
or ( \1939_b1 , \1785_b1 , \1788_b1 );
not ( \1788_b1 , w_3120 );
and ( \1939_b0 , \1785_b0 , w_3121 );
and ( w_3120 , w_3121 , \1788_b0 );
or ( \1940_b1 , \1938_b1 , w_3122 );
or ( \1940_b0 , \1938_b0 , \1939_b0 );
not ( \1939_b0 , w_3123 );
and ( w_3123 , w_3122 , \1939_b1 );
or ( \1941_b1 , \1937_b1 , \1940_b1 );
xor ( \1941_b0 , \1937_b0 , w_3124 );
not ( w_3124 , w_3125 );
and ( w_3125 , \1940_b1 , \1940_b0 );
or ( \1942_b1 , \1018_A[3]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_3126 );
and ( \1942_b0 , \1018_A[3]_b0 , w_3127 );
and ( w_3126 , w_3127 , \1520_B[8]_b0 );
or ( \1943_b1 , \1941_b1 , \1942_b1 );
xor ( \1943_b0 , \1941_b0 , w_3128 );
not ( w_3128 , w_3129 );
and ( w_3129 , \1942_b1 , \1942_b0 );
or ( \1944_b1 , \1789_b1 , \1790_b1 );
not ( \1790_b1 , w_3130 );
and ( \1944_b0 , \1789_b0 , w_3131 );
and ( w_3130 , w_3131 , \1790_b0 );
or ( \1945_b1 , \1791_b1 , \1794_b1 );
not ( \1794_b1 , w_3132 );
and ( \1945_b0 , \1791_b0 , w_3133 );
and ( w_3132 , w_3133 , \1794_b0 );
or ( \1946_b1 , \1944_b1 , w_3134 );
or ( \1946_b0 , \1944_b0 , \1945_b0 );
not ( \1945_b0 , w_3135 );
and ( w_3135 , w_3134 , \1945_b1 );
or ( \1947_b1 , \1943_b1 , \1946_b1 );
xor ( \1947_b0 , \1943_b0 , w_3136 );
not ( w_3136 , w_3137 );
and ( w_3137 , \1946_b1 , \1946_b0 );
or ( \1948_b1 , \962_A[2]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_3138 );
and ( \1948_b0 , \962_A[2]_b0 , w_3139 );
and ( w_3138 , w_3139 , \1654_B[9]_b0 );
or ( \1949_b1 , \1947_b1 , \1948_b1 );
xor ( \1949_b0 , \1947_b0 , w_3140 );
not ( w_3140 , w_3141 );
and ( w_3141 , \1948_b1 , \1948_b0 );
or ( \1950_b1 , \1795_b1 , \1796_b1 );
not ( \1796_b1 , w_3142 );
and ( \1950_b0 , \1795_b0 , w_3143 );
and ( w_3142 , w_3143 , \1796_b0 );
or ( \1951_b1 , \1797_b1 , \1798_b1 );
not ( \1798_b1 , w_3144 );
and ( \1951_b0 , \1797_b0 , w_3145 );
and ( w_3144 , w_3145 , \1798_b0 );
or ( \1952_b1 , \1950_b1 , w_3146 );
or ( \1952_b0 , \1950_b0 , \1951_b0 );
not ( \1951_b0 , w_3147 );
and ( w_3147 , w_3146 , \1951_b1 );
or ( \1953_b1 , \1949_b1 , \1952_b1 );
xor ( \1953_b0 , \1949_b0 , w_3148 );
not ( w_3148 , w_3149 );
and ( w_3149 , \1952_b1 , \1952_b0 );
or ( \1954_b1 , \920_A[1]_b1 , \1800_B[10]_b1 );
not ( \1800_B[10]_b1 , w_3150 );
and ( \1954_b0 , \920_A[1]_b0 , w_3151 );
and ( w_3150 , w_3151 , \1800_B[10]_b0 );
or ( \1955_b1 , \1953_b1 , \1954_b1 );
xor ( \1955_b0 , \1953_b0 , w_3152 );
not ( w_3152 , w_3153 );
and ( w_3153 , \1954_b1 , \1954_b0 );
or ( \1956_b1 , \1799_b1 , \1801_b1 );
not ( \1801_b1 , w_3154 );
and ( \1956_b0 , \1799_b0 , w_3155 );
and ( w_3154 , w_3155 , \1801_b0 );
or ( \1957_b1 , \1955_b1 , \1956_b1 );
xor ( \1957_b0 , \1955_b0 , w_3156 );
not ( w_3156 , w_3157 );
and ( w_3157 , \1956_b1 , \1956_b0 );
buf ( \1958_B[11]_b1 , \c[11]_b1 );
buf ( \1958_B[11]_b0 , \c[11]_b0 );
or ( \1959_b1 , \886_A[0]_b1 , \1958_B[11]_b1 );
not ( \1958_B[11]_b1 , w_3158 );
and ( \1959_b0 , \886_A[0]_b0 , w_3159 );
and ( w_3158 , w_3159 , \1958_B[11]_b0 );
or ( \1960_b1 , \1957_b1 , \1959_b1 );
xor ( \1960_b0 , \1957_b0 , w_3160 );
not ( w_3160 , w_3161 );
and ( w_3161 , \1959_b1 , \1959_b0 );
buf ( \1961_Z[11]_b1 , \1960_b1 );
buf ( \1961_Z[11]_b0 , \1960_b0 );
or ( \1962_b1 , \1961_Z[11]_b1 , \867_b1 );
not ( \867_b1 , w_3162 );
and ( \1962_b0 , \1961_Z[11]_b0 , w_3163 );
and ( w_3162 , w_3163 , \867_b0 );
buf ( \1963_A[11]_b1 , \a[11]_b1 );
buf ( \1963_A[11]_b0 , \a[11]_b0 );
or ( \1964_b1 , \1963_A[11]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_3164 );
and ( \1964_b0 , \1963_A[11]_b0 , w_3165 );
and ( w_3164 , w_3165 , \892_B[0]_b0 );
or ( \1965_b1 , \1805_A[10]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_3166 );
and ( \1965_b0 , \1805_A[10]_b0 , w_3167 );
and ( w_3166 , w_3167 , \929_B[1]_b0 );
or ( \1966_b1 , \1964_b1 , \1965_b1 );
xor ( \1966_b0 , \1964_b0 , w_3168 );
not ( w_3168 , w_3169 );
and ( w_3169 , \1965_b1 , \1965_b0 );
or ( \1967_b1 , \1806_b1 , \1807_b1 );
not ( \1807_b1 , w_3170 );
and ( \1967_b0 , \1806_b0 , w_3171 );
and ( w_3170 , w_3171 , \1807_b0 );
or ( \1968_b1 , \1808_b1 , \1811_b1 );
not ( \1811_b1 , w_3172 );
and ( \1968_b0 , \1808_b0 , w_3173 );
and ( w_3172 , w_3173 , \1811_b0 );
or ( \1969_b1 , \1967_b1 , w_3174 );
or ( \1969_b0 , \1967_b0 , \1968_b0 );
not ( \1968_b0 , w_3175 );
and ( w_3175 , w_3174 , \1968_b1 );
or ( \1970_b1 , \1966_b1 , \1969_b1 );
xor ( \1970_b0 , \1966_b0 , w_3176 );
not ( w_3176 , w_3177 );
and ( w_3177 , \1969_b1 , \1969_b0 );
or ( \1971_b1 , \1659_A[9]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_3178 );
and ( \1971_b0 , \1659_A[9]_b0 , w_3179 );
and ( w_3178 , w_3179 , \979_B[2]_b0 );
or ( \1972_b1 , \1970_b1 , \1971_b1 );
xor ( \1972_b0 , \1970_b0 , w_3180 );
not ( w_3180 , w_3181 );
and ( w_3181 , \1971_b1 , \1971_b0 );
or ( \1973_b1 , \1812_b1 , \1813_b1 );
not ( \1813_b1 , w_3182 );
and ( \1973_b0 , \1812_b0 , w_3183 );
and ( w_3182 , w_3183 , \1813_b0 );
or ( \1974_b1 , \1814_b1 , \1817_b1 );
not ( \1817_b1 , w_3184 );
and ( \1974_b0 , \1814_b0 , w_3185 );
and ( w_3184 , w_3185 , \1817_b0 );
or ( \1975_b1 , \1973_b1 , w_3186 );
or ( \1975_b0 , \1973_b0 , \1974_b0 );
not ( \1974_b0 , w_3187 );
and ( w_3187 , w_3186 , \1974_b1 );
or ( \1976_b1 , \1972_b1 , \1975_b1 );
xor ( \1976_b0 , \1972_b0 , w_3188 );
not ( w_3188 , w_3189 );
and ( w_3189 , \1975_b1 , \1975_b0 );
or ( \1977_b1 , \1525_A[8]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_3190 );
and ( \1977_b0 , \1525_A[8]_b0 , w_3191 );
and ( w_3190 , w_3191 , \1047_B[3]_b0 );
or ( \1978_b1 , \1976_b1 , \1977_b1 );
xor ( \1978_b0 , \1976_b0 , w_3192 );
not ( w_3192 , w_3193 );
and ( w_3193 , \1977_b1 , \1977_b0 );
or ( \1979_b1 , \1818_b1 , \1819_b1 );
not ( \1819_b1 , w_3194 );
and ( \1979_b0 , \1818_b0 , w_3195 );
and ( w_3194 , w_3195 , \1819_b0 );
or ( \1980_b1 , \1820_b1 , \1823_b1 );
not ( \1823_b1 , w_3196 );
and ( \1980_b0 , \1820_b0 , w_3197 );
and ( w_3196 , w_3197 , \1823_b0 );
or ( \1981_b1 , \1979_b1 , w_3198 );
or ( \1981_b0 , \1979_b0 , \1980_b0 );
not ( \1980_b0 , w_3199 );
and ( w_3199 , w_3198 , \1980_b1 );
or ( \1982_b1 , \1978_b1 , \1981_b1 );
xor ( \1982_b0 , \1978_b0 , w_3200 );
not ( w_3200 , w_3201 );
and ( w_3201 , \1981_b1 , \1981_b0 );
or ( \1983_b1 , \1403_A[7]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_3202 );
and ( \1983_b0 , \1403_A[7]_b0 , w_3203 );
and ( w_3202 , w_3203 , \1127_B[4]_b0 );
or ( \1984_b1 , \1982_b1 , \1983_b1 );
xor ( \1984_b0 , \1982_b0 , w_3204 );
not ( w_3204 , w_3205 );
and ( w_3205 , \1983_b1 , \1983_b0 );
or ( \1985_b1 , \1824_b1 , \1825_b1 );
not ( \1825_b1 , w_3206 );
and ( \1985_b0 , \1824_b0 , w_3207 );
and ( w_3206 , w_3207 , \1825_b0 );
or ( \1986_b1 , \1826_b1 , \1829_b1 );
not ( \1829_b1 , w_3208 );
and ( \1986_b0 , \1826_b0 , w_3209 );
and ( w_3208 , w_3209 , \1829_b0 );
or ( \1987_b1 , \1985_b1 , w_3210 );
or ( \1987_b0 , \1985_b0 , \1986_b0 );
not ( \1986_b0 , w_3211 );
and ( w_3211 , w_3210 , \1986_b1 );
or ( \1988_b1 , \1984_b1 , \1987_b1 );
xor ( \1988_b0 , \1984_b0 , w_3212 );
not ( w_3212 , w_3213 );
and ( w_3213 , \1987_b1 , \1987_b0 );
or ( \1989_b1 , \1293_A[6]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_3214 );
and ( \1989_b0 , \1293_A[6]_b0 , w_3215 );
and ( w_3214 , w_3215 , \1219_B[5]_b0 );
or ( \1990_b1 , \1988_b1 , \1989_b1 );
xor ( \1990_b0 , \1988_b0 , w_3216 );
not ( w_3216 , w_3217 );
and ( w_3217 , \1989_b1 , \1989_b0 );
or ( \1991_b1 , \1830_b1 , \1831_b1 );
not ( \1831_b1 , w_3218 );
and ( \1991_b0 , \1830_b0 , w_3219 );
and ( w_3218 , w_3219 , \1831_b0 );
or ( \1992_b1 , \1832_b1 , \1835_b1 );
not ( \1835_b1 , w_3220 );
and ( \1992_b0 , \1832_b0 , w_3221 );
and ( w_3220 , w_3221 , \1835_b0 );
or ( \1993_b1 , \1991_b1 , w_3222 );
or ( \1993_b0 , \1991_b0 , \1992_b0 );
not ( \1992_b0 , w_3223 );
and ( w_3223 , w_3222 , \1992_b1 );
or ( \1994_b1 , \1990_b1 , \1993_b1 );
xor ( \1994_b0 , \1990_b0 , w_3224 );
not ( w_3224 , w_3225 );
and ( w_3225 , \1993_b1 , \1993_b0 );
or ( \1995_b1 , \1195_A[5]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_3226 );
and ( \1995_b0 , \1195_A[5]_b0 , w_3227 );
and ( w_3226 , w_3227 , \1323_B[6]_b0 );
or ( \1996_b1 , \1994_b1 , \1995_b1 );
xor ( \1996_b0 , \1994_b0 , w_3228 );
not ( w_3228 , w_3229 );
and ( w_3229 , \1995_b1 , \1995_b0 );
or ( \1997_b1 , \1836_b1 , \1837_b1 );
not ( \1837_b1 , w_3230 );
and ( \1997_b0 , \1836_b0 , w_3231 );
and ( w_3230 , w_3231 , \1837_b0 );
or ( \1998_b1 , \1838_b1 , \1841_b1 );
not ( \1841_b1 , w_3232 );
and ( \1998_b0 , \1838_b0 , w_3233 );
and ( w_3232 , w_3233 , \1841_b0 );
or ( \1999_b1 , \1997_b1 , w_3234 );
or ( \1999_b0 , \1997_b0 , \1998_b0 );
not ( \1998_b0 , w_3235 );
and ( w_3235 , w_3234 , \1998_b1 );
or ( \2000_b1 , \1996_b1 , \1999_b1 );
xor ( \2000_b0 , \1996_b0 , w_3236 );
not ( w_3236 , w_3237 );
and ( w_3237 , \1999_b1 , \1999_b0 );
or ( \2001_b1 , \1109_A[4]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_3238 );
and ( \2001_b0 , \1109_A[4]_b0 , w_3239 );
and ( w_3238 , w_3239 , \1439_B[7]_b0 );
or ( \2002_b1 , \2000_b1 , \2001_b1 );
xor ( \2002_b0 , \2000_b0 , w_3240 );
not ( w_3240 , w_3241 );
and ( w_3241 , \2001_b1 , \2001_b0 );
or ( \2003_b1 , \1842_b1 , \1843_b1 );
not ( \1843_b1 , w_3242 );
and ( \2003_b0 , \1842_b0 , w_3243 );
and ( w_3242 , w_3243 , \1843_b0 );
or ( \2004_b1 , \1844_b1 , \1847_b1 );
not ( \1847_b1 , w_3244 );
and ( \2004_b0 , \1844_b0 , w_3245 );
and ( w_3244 , w_3245 , \1847_b0 );
or ( \2005_b1 , \2003_b1 , w_3246 );
or ( \2005_b0 , \2003_b0 , \2004_b0 );
not ( \2004_b0 , w_3247 );
and ( w_3247 , w_3246 , \2004_b1 );
or ( \2006_b1 , \2002_b1 , \2005_b1 );
xor ( \2006_b0 , \2002_b0 , w_3248 );
not ( w_3248 , w_3249 );
and ( w_3249 , \2005_b1 , \2005_b0 );
or ( \2007_b1 , \1035_A[3]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_3250 );
and ( \2007_b0 , \1035_A[3]_b0 , w_3251 );
and ( w_3250 , w_3251 , \1567_B[8]_b0 );
or ( \2008_b1 , \2006_b1 , \2007_b1 );
xor ( \2008_b0 , \2006_b0 , w_3252 );
not ( w_3252 , w_3253 );
and ( w_3253 , \2007_b1 , \2007_b0 );
or ( \2009_b1 , \1848_b1 , \1849_b1 );
not ( \1849_b1 , w_3254 );
and ( \2009_b0 , \1848_b0 , w_3255 );
and ( w_3254 , w_3255 , \1849_b0 );
or ( \2010_b1 , \1850_b1 , \1853_b1 );
not ( \1853_b1 , w_3256 );
and ( \2010_b0 , \1850_b0 , w_3257 );
and ( w_3256 , w_3257 , \1853_b0 );
or ( \2011_b1 , \2009_b1 , w_3258 );
or ( \2011_b0 , \2009_b0 , \2010_b0 );
not ( \2010_b0 , w_3259 );
and ( w_3259 , w_3258 , \2010_b1 );
or ( \2012_b1 , \2008_b1 , \2011_b1 );
xor ( \2012_b0 , \2008_b0 , w_3260 );
not ( w_3260 , w_3261 );
and ( w_3261 , \2011_b1 , \2011_b0 );
or ( \2013_b1 , \973_A[2]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_3262 );
and ( \2013_b0 , \973_A[2]_b0 , w_3263 );
and ( w_3262 , w_3263 , \1707_B[9]_b0 );
or ( \2014_b1 , \2012_b1 , \2013_b1 );
xor ( \2014_b0 , \2012_b0 , w_3264 );
not ( w_3264 , w_3265 );
and ( w_3265 , \2013_b1 , \2013_b0 );
or ( \2015_b1 , \1854_b1 , \1855_b1 );
not ( \1855_b1 , w_3266 );
and ( \2015_b0 , \1854_b0 , w_3267 );
and ( w_3266 , w_3267 , \1855_b0 );
or ( \2016_b1 , \1856_b1 , \1857_b1 );
not ( \1857_b1 , w_3268 );
and ( \2016_b0 , \1856_b0 , w_3269 );
and ( w_3268 , w_3269 , \1857_b0 );
or ( \2017_b1 , \2015_b1 , w_3270 );
or ( \2017_b0 , \2015_b0 , \2016_b0 );
not ( \2016_b0 , w_3271 );
and ( w_3271 , w_3270 , \2016_b1 );
or ( \2018_b1 , \2014_b1 , \2017_b1 );
xor ( \2018_b0 , \2014_b0 , w_3272 );
not ( w_3272 , w_3273 );
and ( w_3273 , \2017_b1 , \2017_b0 );
or ( \2019_b1 , \927_A[1]_b1 , \1859_B[10]_b1 );
not ( \1859_B[10]_b1 , w_3274 );
and ( \2019_b0 , \927_A[1]_b0 , w_3275 );
and ( w_3274 , w_3275 , \1859_B[10]_b0 );
or ( \2020_b1 , \2018_b1 , \2019_b1 );
xor ( \2020_b0 , \2018_b0 , w_3276 );
not ( w_3276 , w_3277 );
and ( w_3277 , \2019_b1 , \2019_b0 );
or ( \2021_b1 , \1858_b1 , \1860_b1 );
not ( \1860_b1 , w_3278 );
and ( \2021_b0 , \1858_b0 , w_3279 );
and ( w_3278 , w_3279 , \1860_b0 );
or ( \2022_b1 , \2020_b1 , \2021_b1 );
xor ( \2022_b0 , \2020_b0 , w_3280 );
not ( w_3280 , w_3281 );
and ( w_3281 , \2021_b1 , \2021_b0 );
buf ( \2023_B[11]_b1 , \d[11]_b1 );
buf ( \2023_B[11]_b0 , \d[11]_b0 );
or ( \2024_b1 , \891_A[0]_b1 , \2023_B[11]_b1 );
not ( \2023_B[11]_b1 , w_3282 );
and ( \2024_b0 , \891_A[0]_b0 , w_3283 );
and ( w_3282 , w_3283 , \2023_B[11]_b0 );
or ( \2025_b1 , \2022_b1 , \2024_b1 );
xor ( \2025_b0 , \2022_b0 , w_3284 );
not ( w_3284 , w_3285 );
and ( w_3285 , \2024_b1 , \2024_b0 );
buf ( \2026_Z[11]_b1 , \2025_b1 );
buf ( \2026_Z[11]_b0 , \2025_b0 );
or ( \2027_b1 , \2026_Z[11]_b1 , \865_b1 );
not ( \865_b1 , w_3286 );
and ( \2027_b0 , \2026_Z[11]_b0 , w_3287 );
and ( w_3286 , w_3287 , \865_b0 );
buf ( \2028_A[11]_b1 , \b[11]_b1 );
buf ( \2028_A[11]_b0 , \b[11]_b0 );
buf ( \2029_B[11]_b1 , \d[11]_b1 );
buf ( \2029_B[11]_b0 , \d[11]_b0 );
or ( \2030_b1 , \2028_A[11]_b1 , \2029_B[11]_b1 );
xor ( \2030_b0 , \2028_A[11]_b0 , w_3288 );
not ( w_3288 , w_3289 );
and ( w_3289 , \2029_B[11]_b1 , \2029_B[11]_b0 );
or ( \2031_b1 , \1864_A[10]_b1 , \1865_B[10]_b1 );
not ( \1865_B[10]_b1 , w_3290 );
and ( \2031_b0 , \1864_A[10]_b0 , w_3291 );
and ( w_3290 , w_3291 , \1865_B[10]_b0 );
or ( \2032_b1 , \1865_B[10]_b1 , \1870_b1 );
not ( \1870_b1 , w_3292 );
and ( \2032_b0 , \1865_B[10]_b0 , w_3293 );
and ( w_3292 , w_3293 , \1870_b0 );
or ( \2033_b1 , \1864_A[10]_b1 , \1870_b1 );
not ( \1870_b1 , w_3294 );
and ( \2033_b0 , \1864_A[10]_b0 , w_3295 );
and ( w_3294 , w_3295 , \1870_b0 );
or ( \2035_b1 , \2030_b1 , \2034_b1 );
xor ( \2035_b0 , \2030_b0 , w_3296 );
not ( w_3296 , w_3297 );
and ( w_3297 , \2034_b1 , \2034_b0 );
buf ( \2036_SUM[11]_b1 , \2035_b1 );
buf ( \2036_SUM[11]_b0 , \2035_b0 );
or ( \2037_b1 , \2036_SUM[11]_b1 , \863_b1 );
not ( \863_b1 , w_3298 );
and ( \2037_b0 , \2036_SUM[11]_b0 , w_3299 );
and ( w_3298 , w_3299 , \863_b0 );
buf ( \2038_A[11]_b1 , \a[11]_b1 );
buf ( \2038_A[11]_b0 , \a[11]_b0 );
buf ( \2039_B[11]_b1 , \c[11]_b1 );
buf ( \2039_B[11]_b0 , \c[11]_b0 );
or ( \2040_b1 , \2038_A[11]_b1 , \2039_B[11]_b1 );
xor ( \2040_b0 , \2038_A[11]_b0 , w_3300 );
not ( w_3300 , w_3301 );
and ( w_3301 , \2039_B[11]_b1 , \2039_B[11]_b0 );
or ( \2041_b1 , \1874_A[10]_b1 , \1875_B[10]_b1 );
not ( \1875_B[10]_b1 , w_3302 );
and ( \2041_b0 , \1874_A[10]_b0 , w_3303 );
and ( w_3302 , w_3303 , \1875_B[10]_b0 );
or ( \2042_b1 , \1875_B[10]_b1 , \1880_b1 );
not ( \1880_b1 , w_3304 );
and ( \2042_b0 , \1875_B[10]_b0 , w_3305 );
and ( w_3304 , w_3305 , \1880_b0 );
or ( \2043_b1 , \1874_A[10]_b1 , \1880_b1 );
not ( \1880_b1 , w_3306 );
and ( \2043_b0 , \1874_A[10]_b0 , w_3307 );
and ( w_3306 , w_3307 , \1880_b0 );
or ( \2045_b1 , \2040_b1 , \2044_b1 );
xor ( \2045_b0 , \2040_b0 , w_3308 );
not ( w_3308 , w_3309 );
and ( w_3309 , \2044_b1 , \2044_b0 );
buf ( \2046_SUM[11]_b1 , \2045_b1 );
buf ( \2046_SUM[11]_b0 , \2045_b0 );
or ( \2047_b1 , \2046_SUM[11]_b1 , \861_b1 );
not ( \861_b1 , w_3310 );
and ( \2047_b0 , \2046_SUM[11]_b0 , w_3311 );
and ( w_3310 , w_3311 , \861_b0 );
or ( \2048_b1 , \d[11]_b1 , \859_b1 );
not ( \859_b1 , w_3312 );
and ( \2048_b0 , \d[11]_b0 , w_3313 );
and ( w_3312 , w_3313 , \859_b0 );
or ( \2049_b1 , \c[11]_b1 , \857_b1 );
not ( \857_b1 , w_3314 );
and ( \2049_b0 , \c[11]_b0 , w_3315 );
and ( w_3314 , w_3315 , \857_b0 );
or ( \2050_b1 , \b[11]_b1 , \855_b1 );
not ( \855_b1 , w_3316 );
and ( \2050_b0 , \b[11]_b0 , w_3317 );
and ( w_3316 , w_3317 , \855_b0 );
or ( \2051_b1 , \a[11]_b1 , \853_b1 );
not ( \853_b1 , w_3318 );
and ( \2051_b0 , \a[11]_b0 , w_3319 );
and ( w_3318 , w_3319 , \853_b0 );
and ( \2053_b1 , 1'b0_b1 , w_3320 );
xor ( w_3320 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_3321 );
and ( \2053_b0 , w_3321 , \876_b0 );
or ( \2054_b1 , \a[12]_b1 , w_3322 );
or ( \2054_b0 , \a[12]_b0 , \d[12]_b0 );
not ( \d[12]_b0 , w_3323 );
and ( w_3323 , w_3322 , \d[12]_b1 );
or ( \2055_b1 , \2054_b1 , \875_b1 );
not ( \875_b1 , w_3324 );
and ( \2055_b0 , \2054_b0 , w_3325 );
and ( w_3324 , w_3325 , \875_b0 );
or ( \2056_b1 , \b[12]_b1 , \c[12]_b1 );
not ( \c[12]_b1 , w_3326 );
and ( \2056_b0 , \b[12]_b0 , w_3327 );
and ( w_3326 , w_3327 , \c[12]_b0 );
or ( \2057_b1 , \2056_b1 , \873_b1 );
not ( \873_b1 , w_3328 );
and ( \2057_b0 , \2056_b0 , w_3329 );
and ( w_3328 , w_3329 , \873_b0 );
or ( \2058_b1 , \a[12]_b1 , w_3330 );
or ( \2058_b0 , \a[12]_b0 , \b[12]_b0 );
not ( \b[12]_b0 , w_3331 );
and ( w_3331 , w_3330 , \b[12]_b1 );
or ( \2059_b1 , \2058_b1 , \871_b1 );
not ( \871_b1 , w_3332 );
and ( \2059_b0 , \2058_b0 , w_3333 );
and ( w_3332 , w_3333 , \871_b0 );
or ( \2060_b1 , \c[12]_b1 , \d[12]_b1 );
xor ( \2060_b0 , \c[12]_b0 , w_3334 );
not ( w_3334 , w_3335 );
and ( w_3335 , \d[12]_b1 , \d[12]_b0 );
or ( \2061_b1 , \2060_b1 , \869_b1 );
not ( \869_b1 , w_3336 );
and ( \2061_b0 , \2060_b0 , w_3337 );
and ( w_3336 , w_3337 , \869_b0 );
buf ( \2062_A[12]_b1 , \b[12]_b1 );
buf ( \2062_A[12]_b0 , \b[12]_b0 );
or ( \2063_b1 , \2062_A[12]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_3338 );
and ( \2063_b0 , \2062_A[12]_b0 , w_3339 );
and ( w_3338 , w_3339 , \887_B[0]_b0 );
or ( \2064_b1 , \1898_A[11]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_3340 );
and ( \2064_b0 , \1898_A[11]_b0 , w_3341 );
and ( w_3340 , w_3341 , \922_B[1]_b0 );
or ( \2065_b1 , \2063_b1 , \2064_b1 );
xor ( \2065_b0 , \2063_b0 , w_3342 );
not ( w_3342 , w_3343 );
and ( w_3343 , \2064_b1 , \2064_b0 );
or ( \2066_b1 , \1899_b1 , \1900_b1 );
not ( \1900_b1 , w_3344 );
and ( \2066_b0 , \1899_b0 , w_3345 );
and ( w_3344 , w_3345 , \1900_b0 );
or ( \2067_b1 , \1901_b1 , \1904_b1 );
not ( \1904_b1 , w_3346 );
and ( \2067_b0 , \1901_b0 , w_3347 );
and ( w_3346 , w_3347 , \1904_b0 );
or ( \2068_b1 , \2066_b1 , w_3348 );
or ( \2068_b0 , \2066_b0 , \2067_b0 );
not ( \2067_b0 , w_3349 );
and ( w_3349 , w_3348 , \2067_b1 );
or ( \2069_b1 , \2065_b1 , \2068_b1 );
xor ( \2069_b0 , \2065_b0 , w_3350 );
not ( w_3350 , w_3351 );
and ( w_3351 , \2068_b1 , \2068_b0 );
or ( \2070_b1 , \1746_A[10]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_3352 );
and ( \2070_b0 , \1746_A[10]_b0 , w_3353 );
and ( w_3352 , w_3353 , \968_B[2]_b0 );
or ( \2071_b1 , \2069_b1 , \2070_b1 );
xor ( \2071_b0 , \2069_b0 , w_3354 );
not ( w_3354 , w_3355 );
and ( w_3355 , \2070_b1 , \2070_b0 );
or ( \2072_b1 , \1905_b1 , \1906_b1 );
not ( \1906_b1 , w_3356 );
and ( \2072_b0 , \1905_b0 , w_3357 );
and ( w_3356 , w_3357 , \1906_b0 );
or ( \2073_b1 , \1907_b1 , \1910_b1 );
not ( \1910_b1 , w_3358 );
and ( \2073_b0 , \1907_b0 , w_3359 );
and ( w_3358 , w_3359 , \1910_b0 );
or ( \2074_b1 , \2072_b1 , w_3360 );
or ( \2074_b0 , \2072_b0 , \2073_b0 );
not ( \2073_b0 , w_3361 );
and ( w_3361 , w_3360 , \2073_b1 );
or ( \2075_b1 , \2071_b1 , \2074_b1 );
xor ( \2075_b0 , \2071_b0 , w_3362 );
not ( w_3362 , w_3363 );
and ( w_3363 , \2074_b1 , \2074_b0 );
or ( \2076_b1 , \1606_A[9]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_3364 );
and ( \2076_b0 , \1606_A[9]_b0 , w_3365 );
and ( w_3364 , w_3365 , \1030_B[3]_b0 );
or ( \2077_b1 , \2075_b1 , \2076_b1 );
xor ( \2077_b0 , \2075_b0 , w_3366 );
not ( w_3366 , w_3367 );
and ( w_3367 , \2076_b1 , \2076_b0 );
or ( \2078_b1 , \1911_b1 , \1912_b1 );
not ( \1912_b1 , w_3368 );
and ( \2078_b0 , \1911_b0 , w_3369 );
and ( w_3368 , w_3369 , \1912_b0 );
or ( \2079_b1 , \1913_b1 , \1916_b1 );
not ( \1916_b1 , w_3370 );
and ( \2079_b0 , \1913_b0 , w_3371 );
and ( w_3370 , w_3371 , \1916_b0 );
or ( \2080_b1 , \2078_b1 , w_3372 );
or ( \2080_b0 , \2078_b0 , \2079_b0 );
not ( \2079_b0 , w_3373 );
and ( w_3373 , w_3372 , \2079_b1 );
or ( \2081_b1 , \2077_b1 , \2080_b1 );
xor ( \2081_b0 , \2077_b0 , w_3374 );
not ( w_3374 , w_3375 );
and ( w_3375 , \2080_b1 , \2080_b0 );
or ( \2082_b1 , \1478_A[8]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_3376 );
and ( \2082_b0 , \1478_A[8]_b0 , w_3377 );
and ( w_3376 , w_3377 , \1104_B[4]_b0 );
or ( \2083_b1 , \2081_b1 , \2082_b1 );
xor ( \2083_b0 , \2081_b0 , w_3378 );
not ( w_3378 , w_3379 );
and ( w_3379 , \2082_b1 , \2082_b0 );
or ( \2084_b1 , \1917_b1 , \1918_b1 );
not ( \1918_b1 , w_3380 );
and ( \2084_b0 , \1917_b0 , w_3381 );
and ( w_3380 , w_3381 , \1918_b0 );
or ( \2085_b1 , \1919_b1 , \1922_b1 );
not ( \1922_b1 , w_3382 );
and ( \2085_b0 , \1919_b0 , w_3383 );
and ( w_3382 , w_3383 , \1922_b0 );
or ( \2086_b1 , \2084_b1 , w_3384 );
or ( \2086_b0 , \2084_b0 , \2085_b0 );
not ( \2085_b0 , w_3385 );
and ( w_3385 , w_3384 , \2085_b1 );
or ( \2087_b1 , \2083_b1 , \2086_b1 );
xor ( \2087_b0 , \2083_b0 , w_3386 );
not ( w_3386 , w_3387 );
and ( w_3387 , \2086_b1 , \2086_b0 );
or ( \2088_b1 , \1362_A[7]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_3388 );
and ( \2088_b0 , \1362_A[7]_b0 , w_3389 );
and ( w_3388 , w_3389 , \1190_B[5]_b0 );
or ( \2089_b1 , \2087_b1 , \2088_b1 );
xor ( \2089_b0 , \2087_b0 , w_3390 );
not ( w_3390 , w_3391 );
and ( w_3391 , \2088_b1 , \2088_b0 );
or ( \2090_b1 , \1923_b1 , \1924_b1 );
not ( \1924_b1 , w_3392 );
and ( \2090_b0 , \1923_b0 , w_3393 );
and ( w_3392 , w_3393 , \1924_b0 );
or ( \2091_b1 , \1925_b1 , \1928_b1 );
not ( \1928_b1 , w_3394 );
and ( \2091_b0 , \1925_b0 , w_3395 );
and ( w_3394 , w_3395 , \1928_b0 );
or ( \2092_b1 , \2090_b1 , w_3396 );
or ( \2092_b0 , \2090_b0 , \2091_b0 );
not ( \2091_b0 , w_3397 );
and ( w_3397 , w_3396 , \2091_b1 );
or ( \2093_b1 , \2089_b1 , \2092_b1 );
xor ( \2093_b0 , \2089_b0 , w_3398 );
not ( w_3398 , w_3399 );
and ( w_3399 , \2092_b1 , \2092_b0 );
or ( \2094_b1 , \1258_A[6]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_3400 );
and ( \2094_b0 , \1258_A[6]_b0 , w_3401 );
and ( w_3400 , w_3401 , \1288_B[6]_b0 );
or ( \2095_b1 , \2093_b1 , \2094_b1 );
xor ( \2095_b0 , \2093_b0 , w_3402 );
not ( w_3402 , w_3403 );
and ( w_3403 , \2094_b1 , \2094_b0 );
or ( \2096_b1 , \1929_b1 , \1930_b1 );
not ( \1930_b1 , w_3404 );
and ( \2096_b0 , \1929_b0 , w_3405 );
and ( w_3404 , w_3405 , \1930_b0 );
or ( \2097_b1 , \1931_b1 , \1934_b1 );
not ( \1934_b1 , w_3406 );
and ( \2097_b0 , \1931_b0 , w_3407 );
and ( w_3406 , w_3407 , \1934_b0 );
or ( \2098_b1 , \2096_b1 , w_3408 );
or ( \2098_b0 , \2096_b0 , \2097_b0 );
not ( \2097_b0 , w_3409 );
and ( w_3409 , w_3408 , \2097_b1 );
or ( \2099_b1 , \2095_b1 , \2098_b1 );
xor ( \2099_b0 , \2095_b0 , w_3410 );
not ( w_3410 , w_3411 );
and ( w_3411 , \2098_b1 , \2098_b0 );
or ( \2100_b1 , \1166_A[5]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_3412 );
and ( \2100_b0 , \1166_A[5]_b0 , w_3413 );
and ( w_3412 , w_3413 , \1398_B[7]_b0 );
or ( \2101_b1 , \2099_b1 , \2100_b1 );
xor ( \2101_b0 , \2099_b0 , w_3414 );
not ( w_3414 , w_3415 );
and ( w_3415 , \2100_b1 , \2100_b0 );
or ( \2102_b1 , \1935_b1 , \1936_b1 );
not ( \1936_b1 , w_3416 );
and ( \2102_b0 , \1935_b0 , w_3417 );
and ( w_3416 , w_3417 , \1936_b0 );
or ( \2103_b1 , \1937_b1 , \1940_b1 );
not ( \1940_b1 , w_3418 );
and ( \2103_b0 , \1937_b0 , w_3419 );
and ( w_3418 , w_3419 , \1940_b0 );
or ( \2104_b1 , \2102_b1 , w_3420 );
or ( \2104_b0 , \2102_b0 , \2103_b0 );
not ( \2103_b0 , w_3421 );
and ( w_3421 , w_3420 , \2103_b1 );
or ( \2105_b1 , \2101_b1 , \2104_b1 );
xor ( \2105_b0 , \2101_b0 , w_3422 );
not ( w_3422 , w_3423 );
and ( w_3423 , \2104_b1 , \2104_b0 );
or ( \2106_b1 , \1086_A[4]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_3424 );
and ( \2106_b0 , \1086_A[4]_b0 , w_3425 );
and ( w_3424 , w_3425 , \1520_B[8]_b0 );
or ( \2107_b1 , \2105_b1 , \2106_b1 );
xor ( \2107_b0 , \2105_b0 , w_3426 );
not ( w_3426 , w_3427 );
and ( w_3427 , \2106_b1 , \2106_b0 );
or ( \2108_b1 , \1941_b1 , \1942_b1 );
not ( \1942_b1 , w_3428 );
and ( \2108_b0 , \1941_b0 , w_3429 );
and ( w_3428 , w_3429 , \1942_b0 );
or ( \2109_b1 , \1943_b1 , \1946_b1 );
not ( \1946_b1 , w_3430 );
and ( \2109_b0 , \1943_b0 , w_3431 );
and ( w_3430 , w_3431 , \1946_b0 );
or ( \2110_b1 , \2108_b1 , w_3432 );
or ( \2110_b0 , \2108_b0 , \2109_b0 );
not ( \2109_b0 , w_3433 );
and ( w_3433 , w_3432 , \2109_b1 );
or ( \2111_b1 , \2107_b1 , \2110_b1 );
xor ( \2111_b0 , \2107_b0 , w_3434 );
not ( w_3434 , w_3435 );
and ( w_3435 , \2110_b1 , \2110_b0 );
or ( \2112_b1 , \1018_A[3]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_3436 );
and ( \2112_b0 , \1018_A[3]_b0 , w_3437 );
and ( w_3436 , w_3437 , \1654_B[9]_b0 );
or ( \2113_b1 , \2111_b1 , \2112_b1 );
xor ( \2113_b0 , \2111_b0 , w_3438 );
not ( w_3438 , w_3439 );
and ( w_3439 , \2112_b1 , \2112_b0 );
or ( \2114_b1 , \1947_b1 , \1948_b1 );
not ( \1948_b1 , w_3440 );
and ( \2114_b0 , \1947_b0 , w_3441 );
and ( w_3440 , w_3441 , \1948_b0 );
or ( \2115_b1 , \1949_b1 , \1952_b1 );
not ( \1952_b1 , w_3442 );
and ( \2115_b0 , \1949_b0 , w_3443 );
and ( w_3442 , w_3443 , \1952_b0 );
or ( \2116_b1 , \2114_b1 , w_3444 );
or ( \2116_b0 , \2114_b0 , \2115_b0 );
not ( \2115_b0 , w_3445 );
and ( w_3445 , w_3444 , \2115_b1 );
or ( \2117_b1 , \2113_b1 , \2116_b1 );
xor ( \2117_b0 , \2113_b0 , w_3446 );
not ( w_3446 , w_3447 );
and ( w_3447 , \2116_b1 , \2116_b0 );
or ( \2118_b1 , \962_A[2]_b1 , \1800_B[10]_b1 );
not ( \1800_B[10]_b1 , w_3448 );
and ( \2118_b0 , \962_A[2]_b0 , w_3449 );
and ( w_3448 , w_3449 , \1800_B[10]_b0 );
or ( \2119_b1 , \2117_b1 , \2118_b1 );
xor ( \2119_b0 , \2117_b0 , w_3450 );
not ( w_3450 , w_3451 );
and ( w_3451 , \2118_b1 , \2118_b0 );
or ( \2120_b1 , \1953_b1 , \1954_b1 );
not ( \1954_b1 , w_3452 );
and ( \2120_b0 , \1953_b0 , w_3453 );
and ( w_3452 , w_3453 , \1954_b0 );
or ( \2121_b1 , \1955_b1 , \1956_b1 );
not ( \1956_b1 , w_3454 );
and ( \2121_b0 , \1955_b0 , w_3455 );
and ( w_3454 , w_3455 , \1956_b0 );
or ( \2122_b1 , \2120_b1 , w_3456 );
or ( \2122_b0 , \2120_b0 , \2121_b0 );
not ( \2121_b0 , w_3457 );
and ( w_3457 , w_3456 , \2121_b1 );
or ( \2123_b1 , \2119_b1 , \2122_b1 );
xor ( \2123_b0 , \2119_b0 , w_3458 );
not ( w_3458 , w_3459 );
and ( w_3459 , \2122_b1 , \2122_b0 );
or ( \2124_b1 , \920_A[1]_b1 , \1958_B[11]_b1 );
not ( \1958_B[11]_b1 , w_3460 );
and ( \2124_b0 , \920_A[1]_b0 , w_3461 );
and ( w_3460 , w_3461 , \1958_B[11]_b0 );
or ( \2125_b1 , \2123_b1 , \2124_b1 );
xor ( \2125_b0 , \2123_b0 , w_3462 );
not ( w_3462 , w_3463 );
and ( w_3463 , \2124_b1 , \2124_b0 );
or ( \2126_b1 , \1957_b1 , \1959_b1 );
not ( \1959_b1 , w_3464 );
and ( \2126_b0 , \1957_b0 , w_3465 );
and ( w_3464 , w_3465 , \1959_b0 );
or ( \2127_b1 , \2125_b1 , \2126_b1 );
xor ( \2127_b0 , \2125_b0 , w_3466 );
not ( w_3466 , w_3467 );
and ( w_3467 , \2126_b1 , \2126_b0 );
buf ( \2128_B[12]_b1 , \c[12]_b1 );
buf ( \2128_B[12]_b0 , \c[12]_b0 );
or ( \2129_b1 , \886_A[0]_b1 , \2128_B[12]_b1 );
not ( \2128_B[12]_b1 , w_3468 );
and ( \2129_b0 , \886_A[0]_b0 , w_3469 );
and ( w_3468 , w_3469 , \2128_B[12]_b0 );
or ( \2130_b1 , \2127_b1 , \2129_b1 );
xor ( \2130_b0 , \2127_b0 , w_3470 );
not ( w_3470 , w_3471 );
and ( w_3471 , \2129_b1 , \2129_b0 );
buf ( \2131_Z[12]_b1 , \2130_b1 );
buf ( \2131_Z[12]_b0 , \2130_b0 );
or ( \2132_b1 , \2131_Z[12]_b1 , \867_b1 );
not ( \867_b1 , w_3472 );
and ( \2132_b0 , \2131_Z[12]_b0 , w_3473 );
and ( w_3472 , w_3473 , \867_b0 );
buf ( \2133_A[12]_b1 , \a[12]_b1 );
buf ( \2133_A[12]_b0 , \a[12]_b0 );
or ( \2134_b1 , \2133_A[12]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_3474 );
and ( \2134_b0 , \2133_A[12]_b0 , w_3475 );
and ( w_3474 , w_3475 , \892_B[0]_b0 );
or ( \2135_b1 , \1963_A[11]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_3476 );
and ( \2135_b0 , \1963_A[11]_b0 , w_3477 );
and ( w_3476 , w_3477 , \929_B[1]_b0 );
or ( \2136_b1 , \2134_b1 , \2135_b1 );
xor ( \2136_b0 , \2134_b0 , w_3478 );
not ( w_3478 , w_3479 );
and ( w_3479 , \2135_b1 , \2135_b0 );
or ( \2137_b1 , \1964_b1 , \1965_b1 );
not ( \1965_b1 , w_3480 );
and ( \2137_b0 , \1964_b0 , w_3481 );
and ( w_3480 , w_3481 , \1965_b0 );
or ( \2138_b1 , \1966_b1 , \1969_b1 );
not ( \1969_b1 , w_3482 );
and ( \2138_b0 , \1966_b0 , w_3483 );
and ( w_3482 , w_3483 , \1969_b0 );
or ( \2139_b1 , \2137_b1 , w_3484 );
or ( \2139_b0 , \2137_b0 , \2138_b0 );
not ( \2138_b0 , w_3485 );
and ( w_3485 , w_3484 , \2138_b1 );
or ( \2140_b1 , \2136_b1 , \2139_b1 );
xor ( \2140_b0 , \2136_b0 , w_3486 );
not ( w_3486 , w_3487 );
and ( w_3487 , \2139_b1 , \2139_b0 );
or ( \2141_b1 , \1805_A[10]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_3488 );
and ( \2141_b0 , \1805_A[10]_b0 , w_3489 );
and ( w_3488 , w_3489 , \979_B[2]_b0 );
or ( \2142_b1 , \2140_b1 , \2141_b1 );
xor ( \2142_b0 , \2140_b0 , w_3490 );
not ( w_3490 , w_3491 );
and ( w_3491 , \2141_b1 , \2141_b0 );
or ( \2143_b1 , \1970_b1 , \1971_b1 );
not ( \1971_b1 , w_3492 );
and ( \2143_b0 , \1970_b0 , w_3493 );
and ( w_3492 , w_3493 , \1971_b0 );
or ( \2144_b1 , \1972_b1 , \1975_b1 );
not ( \1975_b1 , w_3494 );
and ( \2144_b0 , \1972_b0 , w_3495 );
and ( w_3494 , w_3495 , \1975_b0 );
or ( \2145_b1 , \2143_b1 , w_3496 );
or ( \2145_b0 , \2143_b0 , \2144_b0 );
not ( \2144_b0 , w_3497 );
and ( w_3497 , w_3496 , \2144_b1 );
or ( \2146_b1 , \2142_b1 , \2145_b1 );
xor ( \2146_b0 , \2142_b0 , w_3498 );
not ( w_3498 , w_3499 );
and ( w_3499 , \2145_b1 , \2145_b0 );
or ( \2147_b1 , \1659_A[9]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_3500 );
and ( \2147_b0 , \1659_A[9]_b0 , w_3501 );
and ( w_3500 , w_3501 , \1047_B[3]_b0 );
or ( \2148_b1 , \2146_b1 , \2147_b1 );
xor ( \2148_b0 , \2146_b0 , w_3502 );
not ( w_3502 , w_3503 );
and ( w_3503 , \2147_b1 , \2147_b0 );
or ( \2149_b1 , \1976_b1 , \1977_b1 );
not ( \1977_b1 , w_3504 );
and ( \2149_b0 , \1976_b0 , w_3505 );
and ( w_3504 , w_3505 , \1977_b0 );
or ( \2150_b1 , \1978_b1 , \1981_b1 );
not ( \1981_b1 , w_3506 );
and ( \2150_b0 , \1978_b0 , w_3507 );
and ( w_3506 , w_3507 , \1981_b0 );
or ( \2151_b1 , \2149_b1 , w_3508 );
or ( \2151_b0 , \2149_b0 , \2150_b0 );
not ( \2150_b0 , w_3509 );
and ( w_3509 , w_3508 , \2150_b1 );
or ( \2152_b1 , \2148_b1 , \2151_b1 );
xor ( \2152_b0 , \2148_b0 , w_3510 );
not ( w_3510 , w_3511 );
and ( w_3511 , \2151_b1 , \2151_b0 );
or ( \2153_b1 , \1525_A[8]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_3512 );
and ( \2153_b0 , \1525_A[8]_b0 , w_3513 );
and ( w_3512 , w_3513 , \1127_B[4]_b0 );
or ( \2154_b1 , \2152_b1 , \2153_b1 );
xor ( \2154_b0 , \2152_b0 , w_3514 );
not ( w_3514 , w_3515 );
and ( w_3515 , \2153_b1 , \2153_b0 );
or ( \2155_b1 , \1982_b1 , \1983_b1 );
not ( \1983_b1 , w_3516 );
and ( \2155_b0 , \1982_b0 , w_3517 );
and ( w_3516 , w_3517 , \1983_b0 );
or ( \2156_b1 , \1984_b1 , \1987_b1 );
not ( \1987_b1 , w_3518 );
and ( \2156_b0 , \1984_b0 , w_3519 );
and ( w_3518 , w_3519 , \1987_b0 );
or ( \2157_b1 , \2155_b1 , w_3520 );
or ( \2157_b0 , \2155_b0 , \2156_b0 );
not ( \2156_b0 , w_3521 );
and ( w_3521 , w_3520 , \2156_b1 );
or ( \2158_b1 , \2154_b1 , \2157_b1 );
xor ( \2158_b0 , \2154_b0 , w_3522 );
not ( w_3522 , w_3523 );
and ( w_3523 , \2157_b1 , \2157_b0 );
or ( \2159_b1 , \1403_A[7]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_3524 );
and ( \2159_b0 , \1403_A[7]_b0 , w_3525 );
and ( w_3524 , w_3525 , \1219_B[5]_b0 );
or ( \2160_b1 , \2158_b1 , \2159_b1 );
xor ( \2160_b0 , \2158_b0 , w_3526 );
not ( w_3526 , w_3527 );
and ( w_3527 , \2159_b1 , \2159_b0 );
or ( \2161_b1 , \1988_b1 , \1989_b1 );
not ( \1989_b1 , w_3528 );
and ( \2161_b0 , \1988_b0 , w_3529 );
and ( w_3528 , w_3529 , \1989_b0 );
or ( \2162_b1 , \1990_b1 , \1993_b1 );
not ( \1993_b1 , w_3530 );
and ( \2162_b0 , \1990_b0 , w_3531 );
and ( w_3530 , w_3531 , \1993_b0 );
or ( \2163_b1 , \2161_b1 , w_3532 );
or ( \2163_b0 , \2161_b0 , \2162_b0 );
not ( \2162_b0 , w_3533 );
and ( w_3533 , w_3532 , \2162_b1 );
or ( \2164_b1 , \2160_b1 , \2163_b1 );
xor ( \2164_b0 , \2160_b0 , w_3534 );
not ( w_3534 , w_3535 );
and ( w_3535 , \2163_b1 , \2163_b0 );
or ( \2165_b1 , \1293_A[6]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_3536 );
and ( \2165_b0 , \1293_A[6]_b0 , w_3537 );
and ( w_3536 , w_3537 , \1323_B[6]_b0 );
or ( \2166_b1 , \2164_b1 , \2165_b1 );
xor ( \2166_b0 , \2164_b0 , w_3538 );
not ( w_3538 , w_3539 );
and ( w_3539 , \2165_b1 , \2165_b0 );
or ( \2167_b1 , \1994_b1 , \1995_b1 );
not ( \1995_b1 , w_3540 );
and ( \2167_b0 , \1994_b0 , w_3541 );
and ( w_3540 , w_3541 , \1995_b0 );
or ( \2168_b1 , \1996_b1 , \1999_b1 );
not ( \1999_b1 , w_3542 );
and ( \2168_b0 , \1996_b0 , w_3543 );
and ( w_3542 , w_3543 , \1999_b0 );
or ( \2169_b1 , \2167_b1 , w_3544 );
or ( \2169_b0 , \2167_b0 , \2168_b0 );
not ( \2168_b0 , w_3545 );
and ( w_3545 , w_3544 , \2168_b1 );
or ( \2170_b1 , \2166_b1 , \2169_b1 );
xor ( \2170_b0 , \2166_b0 , w_3546 );
not ( w_3546 , w_3547 );
and ( w_3547 , \2169_b1 , \2169_b0 );
or ( \2171_b1 , \1195_A[5]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_3548 );
and ( \2171_b0 , \1195_A[5]_b0 , w_3549 );
and ( w_3548 , w_3549 , \1439_B[7]_b0 );
or ( \2172_b1 , \2170_b1 , \2171_b1 );
xor ( \2172_b0 , \2170_b0 , w_3550 );
not ( w_3550 , w_3551 );
and ( w_3551 , \2171_b1 , \2171_b0 );
or ( \2173_b1 , \2000_b1 , \2001_b1 );
not ( \2001_b1 , w_3552 );
and ( \2173_b0 , \2000_b0 , w_3553 );
and ( w_3552 , w_3553 , \2001_b0 );
or ( \2174_b1 , \2002_b1 , \2005_b1 );
not ( \2005_b1 , w_3554 );
and ( \2174_b0 , \2002_b0 , w_3555 );
and ( w_3554 , w_3555 , \2005_b0 );
or ( \2175_b1 , \2173_b1 , w_3556 );
or ( \2175_b0 , \2173_b0 , \2174_b0 );
not ( \2174_b0 , w_3557 );
and ( w_3557 , w_3556 , \2174_b1 );
or ( \2176_b1 , \2172_b1 , \2175_b1 );
xor ( \2176_b0 , \2172_b0 , w_3558 );
not ( w_3558 , w_3559 );
and ( w_3559 , \2175_b1 , \2175_b0 );
or ( \2177_b1 , \1109_A[4]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_3560 );
and ( \2177_b0 , \1109_A[4]_b0 , w_3561 );
and ( w_3560 , w_3561 , \1567_B[8]_b0 );
or ( \2178_b1 , \2176_b1 , \2177_b1 );
xor ( \2178_b0 , \2176_b0 , w_3562 );
not ( w_3562 , w_3563 );
and ( w_3563 , \2177_b1 , \2177_b0 );
or ( \2179_b1 , \2006_b1 , \2007_b1 );
not ( \2007_b1 , w_3564 );
and ( \2179_b0 , \2006_b0 , w_3565 );
and ( w_3564 , w_3565 , \2007_b0 );
or ( \2180_b1 , \2008_b1 , \2011_b1 );
not ( \2011_b1 , w_3566 );
and ( \2180_b0 , \2008_b0 , w_3567 );
and ( w_3566 , w_3567 , \2011_b0 );
or ( \2181_b1 , \2179_b1 , w_3568 );
or ( \2181_b0 , \2179_b0 , \2180_b0 );
not ( \2180_b0 , w_3569 );
and ( w_3569 , w_3568 , \2180_b1 );
or ( \2182_b1 , \2178_b1 , \2181_b1 );
xor ( \2182_b0 , \2178_b0 , w_3570 );
not ( w_3570 , w_3571 );
and ( w_3571 , \2181_b1 , \2181_b0 );
or ( \2183_b1 , \1035_A[3]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_3572 );
and ( \2183_b0 , \1035_A[3]_b0 , w_3573 );
and ( w_3572 , w_3573 , \1707_B[9]_b0 );
or ( \2184_b1 , \2182_b1 , \2183_b1 );
xor ( \2184_b0 , \2182_b0 , w_3574 );
not ( w_3574 , w_3575 );
and ( w_3575 , \2183_b1 , \2183_b0 );
or ( \2185_b1 , \2012_b1 , \2013_b1 );
not ( \2013_b1 , w_3576 );
and ( \2185_b0 , \2012_b0 , w_3577 );
and ( w_3576 , w_3577 , \2013_b0 );
or ( \2186_b1 , \2014_b1 , \2017_b1 );
not ( \2017_b1 , w_3578 );
and ( \2186_b0 , \2014_b0 , w_3579 );
and ( w_3578 , w_3579 , \2017_b0 );
or ( \2187_b1 , \2185_b1 , w_3580 );
or ( \2187_b0 , \2185_b0 , \2186_b0 );
not ( \2186_b0 , w_3581 );
and ( w_3581 , w_3580 , \2186_b1 );
or ( \2188_b1 , \2184_b1 , \2187_b1 );
xor ( \2188_b0 , \2184_b0 , w_3582 );
not ( w_3582 , w_3583 );
and ( w_3583 , \2187_b1 , \2187_b0 );
or ( \2189_b1 , \973_A[2]_b1 , \1859_B[10]_b1 );
not ( \1859_B[10]_b1 , w_3584 );
and ( \2189_b0 , \973_A[2]_b0 , w_3585 );
and ( w_3584 , w_3585 , \1859_B[10]_b0 );
or ( \2190_b1 , \2188_b1 , \2189_b1 );
xor ( \2190_b0 , \2188_b0 , w_3586 );
not ( w_3586 , w_3587 );
and ( w_3587 , \2189_b1 , \2189_b0 );
or ( \2191_b1 , \2018_b1 , \2019_b1 );
not ( \2019_b1 , w_3588 );
and ( \2191_b0 , \2018_b0 , w_3589 );
and ( w_3588 , w_3589 , \2019_b0 );
or ( \2192_b1 , \2020_b1 , \2021_b1 );
not ( \2021_b1 , w_3590 );
and ( \2192_b0 , \2020_b0 , w_3591 );
and ( w_3590 , w_3591 , \2021_b0 );
or ( \2193_b1 , \2191_b1 , w_3592 );
or ( \2193_b0 , \2191_b0 , \2192_b0 );
not ( \2192_b0 , w_3593 );
and ( w_3593 , w_3592 , \2192_b1 );
or ( \2194_b1 , \2190_b1 , \2193_b1 );
xor ( \2194_b0 , \2190_b0 , w_3594 );
not ( w_3594 , w_3595 );
and ( w_3595 , \2193_b1 , \2193_b0 );
or ( \2195_b1 , \927_A[1]_b1 , \2023_B[11]_b1 );
not ( \2023_B[11]_b1 , w_3596 );
and ( \2195_b0 , \927_A[1]_b0 , w_3597 );
and ( w_3596 , w_3597 , \2023_B[11]_b0 );
or ( \2196_b1 , \2194_b1 , \2195_b1 );
xor ( \2196_b0 , \2194_b0 , w_3598 );
not ( w_3598 , w_3599 );
and ( w_3599 , \2195_b1 , \2195_b0 );
or ( \2197_b1 , \2022_b1 , \2024_b1 );
not ( \2024_b1 , w_3600 );
and ( \2197_b0 , \2022_b0 , w_3601 );
and ( w_3600 , w_3601 , \2024_b0 );
or ( \2198_b1 , \2196_b1 , \2197_b1 );
xor ( \2198_b0 , \2196_b0 , w_3602 );
not ( w_3602 , w_3603 );
and ( w_3603 , \2197_b1 , \2197_b0 );
buf ( \2199_B[12]_b1 , \d[12]_b1 );
buf ( \2199_B[12]_b0 , \d[12]_b0 );
or ( \2200_b1 , \891_A[0]_b1 , \2199_B[12]_b1 );
not ( \2199_B[12]_b1 , w_3604 );
and ( \2200_b0 , \891_A[0]_b0 , w_3605 );
and ( w_3604 , w_3605 , \2199_B[12]_b0 );
or ( \2201_b1 , \2198_b1 , \2200_b1 );
xor ( \2201_b0 , \2198_b0 , w_3606 );
not ( w_3606 , w_3607 );
and ( w_3607 , \2200_b1 , \2200_b0 );
buf ( \2202_Z[12]_b1 , \2201_b1 );
buf ( \2202_Z[12]_b0 , \2201_b0 );
or ( \2203_b1 , \2202_Z[12]_b1 , \865_b1 );
not ( \865_b1 , w_3608 );
and ( \2203_b0 , \2202_Z[12]_b0 , w_3609 );
and ( w_3608 , w_3609 , \865_b0 );
buf ( \2204_A[12]_b1 , \b[12]_b1 );
buf ( \2204_A[12]_b0 , \b[12]_b0 );
buf ( \2205_B[12]_b1 , \d[12]_b1 );
buf ( \2205_B[12]_b0 , \d[12]_b0 );
or ( \2206_b1 , \2204_A[12]_b1 , \2205_B[12]_b1 );
xor ( \2206_b0 , \2204_A[12]_b0 , w_3610 );
not ( w_3610 , w_3611 );
and ( w_3611 , \2205_B[12]_b1 , \2205_B[12]_b0 );
or ( \2207_b1 , \2028_A[11]_b1 , \2029_B[11]_b1 );
not ( \2029_B[11]_b1 , w_3612 );
and ( \2207_b0 , \2028_A[11]_b0 , w_3613 );
and ( w_3612 , w_3613 , \2029_B[11]_b0 );
or ( \2208_b1 , \2029_B[11]_b1 , \2034_b1 );
not ( \2034_b1 , w_3614 );
and ( \2208_b0 , \2029_B[11]_b0 , w_3615 );
and ( w_3614 , w_3615 , \2034_b0 );
or ( \2209_b1 , \2028_A[11]_b1 , \2034_b1 );
not ( \2034_b1 , w_3616 );
and ( \2209_b0 , \2028_A[11]_b0 , w_3617 );
and ( w_3616 , w_3617 , \2034_b0 );
or ( \2211_b1 , \2206_b1 , \2210_b1 );
xor ( \2211_b0 , \2206_b0 , w_3618 );
not ( w_3618 , w_3619 );
and ( w_3619 , \2210_b1 , \2210_b0 );
buf ( \2212_SUM[12]_b1 , \2211_b1 );
buf ( \2212_SUM[12]_b0 , \2211_b0 );
or ( \2213_b1 , \2212_SUM[12]_b1 , \863_b1 );
not ( \863_b1 , w_3620 );
and ( \2213_b0 , \2212_SUM[12]_b0 , w_3621 );
and ( w_3620 , w_3621 , \863_b0 );
buf ( \2214_A[12]_b1 , \a[12]_b1 );
buf ( \2214_A[12]_b0 , \a[12]_b0 );
buf ( \2215_B[12]_b1 , \c[12]_b1 );
buf ( \2215_B[12]_b0 , \c[12]_b0 );
or ( \2216_b1 , \2214_A[12]_b1 , \2215_B[12]_b1 );
xor ( \2216_b0 , \2214_A[12]_b0 , w_3622 );
not ( w_3622 , w_3623 );
and ( w_3623 , \2215_B[12]_b1 , \2215_B[12]_b0 );
or ( \2217_b1 , \2038_A[11]_b1 , \2039_B[11]_b1 );
not ( \2039_B[11]_b1 , w_3624 );
and ( \2217_b0 , \2038_A[11]_b0 , w_3625 );
and ( w_3624 , w_3625 , \2039_B[11]_b0 );
or ( \2218_b1 , \2039_B[11]_b1 , \2044_b1 );
not ( \2044_b1 , w_3626 );
and ( \2218_b0 , \2039_B[11]_b0 , w_3627 );
and ( w_3626 , w_3627 , \2044_b0 );
or ( \2219_b1 , \2038_A[11]_b1 , \2044_b1 );
not ( \2044_b1 , w_3628 );
and ( \2219_b0 , \2038_A[11]_b0 , w_3629 );
and ( w_3628 , w_3629 , \2044_b0 );
or ( \2221_b1 , \2216_b1 , \2220_b1 );
xor ( \2221_b0 , \2216_b0 , w_3630 );
not ( w_3630 , w_3631 );
and ( w_3631 , \2220_b1 , \2220_b0 );
buf ( \2222_SUM[12]_b1 , \2221_b1 );
buf ( \2222_SUM[12]_b0 , \2221_b0 );
or ( \2223_b1 , \2222_SUM[12]_b1 , \861_b1 );
not ( \861_b1 , w_3632 );
and ( \2223_b0 , \2222_SUM[12]_b0 , w_3633 );
and ( w_3632 , w_3633 , \861_b0 );
or ( \2224_b1 , \d[12]_b1 , \859_b1 );
not ( \859_b1 , w_3634 );
and ( \2224_b0 , \d[12]_b0 , w_3635 );
and ( w_3634 , w_3635 , \859_b0 );
or ( \2225_b1 , \c[12]_b1 , \857_b1 );
not ( \857_b1 , w_3636 );
and ( \2225_b0 , \c[12]_b0 , w_3637 );
and ( w_3636 , w_3637 , \857_b0 );
or ( \2226_b1 , \b[12]_b1 , \855_b1 );
not ( \855_b1 , w_3638 );
and ( \2226_b0 , \b[12]_b0 , w_3639 );
and ( w_3638 , w_3639 , \855_b0 );
or ( \2227_b1 , \a[12]_b1 , \853_b1 );
not ( \853_b1 , w_3640 );
and ( \2227_b0 , \a[12]_b0 , w_3641 );
and ( w_3640 , w_3641 , \853_b0 );
and ( \2229_b1 , 1'b0_b1 , w_3642 );
xor ( w_3642 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_3643 );
and ( \2229_b0 , w_3643 , \876_b0 );
or ( \2230_b1 , \a[13]_b1 , w_3644 );
or ( \2230_b0 , \a[13]_b0 , \d[13]_b0 );
not ( \d[13]_b0 , w_3645 );
and ( w_3645 , w_3644 , \d[13]_b1 );
or ( \2231_b1 , \2230_b1 , \875_b1 );
not ( \875_b1 , w_3646 );
and ( \2231_b0 , \2230_b0 , w_3647 );
and ( w_3646 , w_3647 , \875_b0 );
or ( \2232_b1 , \b[13]_b1 , \c[13]_b1 );
not ( \c[13]_b1 , w_3648 );
and ( \2232_b0 , \b[13]_b0 , w_3649 );
and ( w_3648 , w_3649 , \c[13]_b0 );
or ( \2233_b1 , \2232_b1 , \873_b1 );
not ( \873_b1 , w_3650 );
and ( \2233_b0 , \2232_b0 , w_3651 );
and ( w_3650 , w_3651 , \873_b0 );
or ( \2234_b1 , \a[13]_b1 , w_3652 );
or ( \2234_b0 , \a[13]_b0 , \b[13]_b0 );
not ( \b[13]_b0 , w_3653 );
and ( w_3653 , w_3652 , \b[13]_b1 );
or ( \2235_b1 , \2234_b1 , \871_b1 );
not ( \871_b1 , w_3654 );
and ( \2235_b0 , \2234_b0 , w_3655 );
and ( w_3654 , w_3655 , \871_b0 );
or ( \2236_b1 , \c[13]_b1 , \d[13]_b1 );
xor ( \2236_b0 , \c[13]_b0 , w_3656 );
not ( w_3656 , w_3657 );
and ( w_3657 , \d[13]_b1 , \d[13]_b0 );
or ( \2237_b1 , \2236_b1 , \869_b1 );
not ( \869_b1 , w_3658 );
and ( \2237_b0 , \2236_b0 , w_3659 );
and ( w_3658 , w_3659 , \869_b0 );
buf ( \2238_A[13]_b1 , \b[13]_b1 );
buf ( \2238_A[13]_b0 , \b[13]_b0 );
or ( \2239_b1 , \2238_A[13]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_3660 );
and ( \2239_b0 , \2238_A[13]_b0 , w_3661 );
and ( w_3660 , w_3661 , \887_B[0]_b0 );
or ( \2240_b1 , \2062_A[12]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_3662 );
and ( \2240_b0 , \2062_A[12]_b0 , w_3663 );
and ( w_3662 , w_3663 , \922_B[1]_b0 );
or ( \2241_b1 , \2239_b1 , \2240_b1 );
xor ( \2241_b0 , \2239_b0 , w_3664 );
not ( w_3664 , w_3665 );
and ( w_3665 , \2240_b1 , \2240_b0 );
or ( \2242_b1 , \2063_b1 , \2064_b1 );
not ( \2064_b1 , w_3666 );
and ( \2242_b0 , \2063_b0 , w_3667 );
and ( w_3666 , w_3667 , \2064_b0 );
or ( \2243_b1 , \2065_b1 , \2068_b1 );
not ( \2068_b1 , w_3668 );
and ( \2243_b0 , \2065_b0 , w_3669 );
and ( w_3668 , w_3669 , \2068_b0 );
or ( \2244_b1 , \2242_b1 , w_3670 );
or ( \2244_b0 , \2242_b0 , \2243_b0 );
not ( \2243_b0 , w_3671 );
and ( w_3671 , w_3670 , \2243_b1 );
or ( \2245_b1 , \2241_b1 , \2244_b1 );
xor ( \2245_b0 , \2241_b0 , w_3672 );
not ( w_3672 , w_3673 );
and ( w_3673 , \2244_b1 , \2244_b0 );
or ( \2246_b1 , \1898_A[11]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_3674 );
and ( \2246_b0 , \1898_A[11]_b0 , w_3675 );
and ( w_3674 , w_3675 , \968_B[2]_b0 );
or ( \2247_b1 , \2245_b1 , \2246_b1 );
xor ( \2247_b0 , \2245_b0 , w_3676 );
not ( w_3676 , w_3677 );
and ( w_3677 , \2246_b1 , \2246_b0 );
or ( \2248_b1 , \2069_b1 , \2070_b1 );
not ( \2070_b1 , w_3678 );
and ( \2248_b0 , \2069_b0 , w_3679 );
and ( w_3678 , w_3679 , \2070_b0 );
or ( \2249_b1 , \2071_b1 , \2074_b1 );
not ( \2074_b1 , w_3680 );
and ( \2249_b0 , \2071_b0 , w_3681 );
and ( w_3680 , w_3681 , \2074_b0 );
or ( \2250_b1 , \2248_b1 , w_3682 );
or ( \2250_b0 , \2248_b0 , \2249_b0 );
not ( \2249_b0 , w_3683 );
and ( w_3683 , w_3682 , \2249_b1 );
or ( \2251_b1 , \2247_b1 , \2250_b1 );
xor ( \2251_b0 , \2247_b0 , w_3684 );
not ( w_3684 , w_3685 );
and ( w_3685 , \2250_b1 , \2250_b0 );
or ( \2252_b1 , \1746_A[10]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_3686 );
and ( \2252_b0 , \1746_A[10]_b0 , w_3687 );
and ( w_3686 , w_3687 , \1030_B[3]_b0 );
or ( \2253_b1 , \2251_b1 , \2252_b1 );
xor ( \2253_b0 , \2251_b0 , w_3688 );
not ( w_3688 , w_3689 );
and ( w_3689 , \2252_b1 , \2252_b0 );
or ( \2254_b1 , \2075_b1 , \2076_b1 );
not ( \2076_b1 , w_3690 );
and ( \2254_b0 , \2075_b0 , w_3691 );
and ( w_3690 , w_3691 , \2076_b0 );
or ( \2255_b1 , \2077_b1 , \2080_b1 );
not ( \2080_b1 , w_3692 );
and ( \2255_b0 , \2077_b0 , w_3693 );
and ( w_3692 , w_3693 , \2080_b0 );
or ( \2256_b1 , \2254_b1 , w_3694 );
or ( \2256_b0 , \2254_b0 , \2255_b0 );
not ( \2255_b0 , w_3695 );
and ( w_3695 , w_3694 , \2255_b1 );
or ( \2257_b1 , \2253_b1 , \2256_b1 );
xor ( \2257_b0 , \2253_b0 , w_3696 );
not ( w_3696 , w_3697 );
and ( w_3697 , \2256_b1 , \2256_b0 );
or ( \2258_b1 , \1606_A[9]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_3698 );
and ( \2258_b0 , \1606_A[9]_b0 , w_3699 );
and ( w_3698 , w_3699 , \1104_B[4]_b0 );
or ( \2259_b1 , \2257_b1 , \2258_b1 );
xor ( \2259_b0 , \2257_b0 , w_3700 );
not ( w_3700 , w_3701 );
and ( w_3701 , \2258_b1 , \2258_b0 );
or ( \2260_b1 , \2081_b1 , \2082_b1 );
not ( \2082_b1 , w_3702 );
and ( \2260_b0 , \2081_b0 , w_3703 );
and ( w_3702 , w_3703 , \2082_b0 );
or ( \2261_b1 , \2083_b1 , \2086_b1 );
not ( \2086_b1 , w_3704 );
and ( \2261_b0 , \2083_b0 , w_3705 );
and ( w_3704 , w_3705 , \2086_b0 );
or ( \2262_b1 , \2260_b1 , w_3706 );
or ( \2262_b0 , \2260_b0 , \2261_b0 );
not ( \2261_b0 , w_3707 );
and ( w_3707 , w_3706 , \2261_b1 );
or ( \2263_b1 , \2259_b1 , \2262_b1 );
xor ( \2263_b0 , \2259_b0 , w_3708 );
not ( w_3708 , w_3709 );
and ( w_3709 , \2262_b1 , \2262_b0 );
or ( \2264_b1 , \1478_A[8]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_3710 );
and ( \2264_b0 , \1478_A[8]_b0 , w_3711 );
and ( w_3710 , w_3711 , \1190_B[5]_b0 );
or ( \2265_b1 , \2263_b1 , \2264_b1 );
xor ( \2265_b0 , \2263_b0 , w_3712 );
not ( w_3712 , w_3713 );
and ( w_3713 , \2264_b1 , \2264_b0 );
or ( \2266_b1 , \2087_b1 , \2088_b1 );
not ( \2088_b1 , w_3714 );
and ( \2266_b0 , \2087_b0 , w_3715 );
and ( w_3714 , w_3715 , \2088_b0 );
or ( \2267_b1 , \2089_b1 , \2092_b1 );
not ( \2092_b1 , w_3716 );
and ( \2267_b0 , \2089_b0 , w_3717 );
and ( w_3716 , w_3717 , \2092_b0 );
or ( \2268_b1 , \2266_b1 , w_3718 );
or ( \2268_b0 , \2266_b0 , \2267_b0 );
not ( \2267_b0 , w_3719 );
and ( w_3719 , w_3718 , \2267_b1 );
or ( \2269_b1 , \2265_b1 , \2268_b1 );
xor ( \2269_b0 , \2265_b0 , w_3720 );
not ( w_3720 , w_3721 );
and ( w_3721 , \2268_b1 , \2268_b0 );
or ( \2270_b1 , \1362_A[7]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_3722 );
and ( \2270_b0 , \1362_A[7]_b0 , w_3723 );
and ( w_3722 , w_3723 , \1288_B[6]_b0 );
or ( \2271_b1 , \2269_b1 , \2270_b1 );
xor ( \2271_b0 , \2269_b0 , w_3724 );
not ( w_3724 , w_3725 );
and ( w_3725 , \2270_b1 , \2270_b0 );
or ( \2272_b1 , \2093_b1 , \2094_b1 );
not ( \2094_b1 , w_3726 );
and ( \2272_b0 , \2093_b0 , w_3727 );
and ( w_3726 , w_3727 , \2094_b0 );
or ( \2273_b1 , \2095_b1 , \2098_b1 );
not ( \2098_b1 , w_3728 );
and ( \2273_b0 , \2095_b0 , w_3729 );
and ( w_3728 , w_3729 , \2098_b0 );
or ( \2274_b1 , \2272_b1 , w_3730 );
or ( \2274_b0 , \2272_b0 , \2273_b0 );
not ( \2273_b0 , w_3731 );
and ( w_3731 , w_3730 , \2273_b1 );
or ( \2275_b1 , \2271_b1 , \2274_b1 );
xor ( \2275_b0 , \2271_b0 , w_3732 );
not ( w_3732 , w_3733 );
and ( w_3733 , \2274_b1 , \2274_b0 );
or ( \2276_b1 , \1258_A[6]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_3734 );
and ( \2276_b0 , \1258_A[6]_b0 , w_3735 );
and ( w_3734 , w_3735 , \1398_B[7]_b0 );
or ( \2277_b1 , \2275_b1 , \2276_b1 );
xor ( \2277_b0 , \2275_b0 , w_3736 );
not ( w_3736 , w_3737 );
and ( w_3737 , \2276_b1 , \2276_b0 );
or ( \2278_b1 , \2099_b1 , \2100_b1 );
not ( \2100_b1 , w_3738 );
and ( \2278_b0 , \2099_b0 , w_3739 );
and ( w_3738 , w_3739 , \2100_b0 );
or ( \2279_b1 , \2101_b1 , \2104_b1 );
not ( \2104_b1 , w_3740 );
and ( \2279_b0 , \2101_b0 , w_3741 );
and ( w_3740 , w_3741 , \2104_b0 );
or ( \2280_b1 , \2278_b1 , w_3742 );
or ( \2280_b0 , \2278_b0 , \2279_b0 );
not ( \2279_b0 , w_3743 );
and ( w_3743 , w_3742 , \2279_b1 );
or ( \2281_b1 , \2277_b1 , \2280_b1 );
xor ( \2281_b0 , \2277_b0 , w_3744 );
not ( w_3744 , w_3745 );
and ( w_3745 , \2280_b1 , \2280_b0 );
or ( \2282_b1 , \1166_A[5]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_3746 );
and ( \2282_b0 , \1166_A[5]_b0 , w_3747 );
and ( w_3746 , w_3747 , \1520_B[8]_b0 );
or ( \2283_b1 , \2281_b1 , \2282_b1 );
xor ( \2283_b0 , \2281_b0 , w_3748 );
not ( w_3748 , w_3749 );
and ( w_3749 , \2282_b1 , \2282_b0 );
or ( \2284_b1 , \2105_b1 , \2106_b1 );
not ( \2106_b1 , w_3750 );
and ( \2284_b0 , \2105_b0 , w_3751 );
and ( w_3750 , w_3751 , \2106_b0 );
or ( \2285_b1 , \2107_b1 , \2110_b1 );
not ( \2110_b1 , w_3752 );
and ( \2285_b0 , \2107_b0 , w_3753 );
and ( w_3752 , w_3753 , \2110_b0 );
or ( \2286_b1 , \2284_b1 , w_3754 );
or ( \2286_b0 , \2284_b0 , \2285_b0 );
not ( \2285_b0 , w_3755 );
and ( w_3755 , w_3754 , \2285_b1 );
or ( \2287_b1 , \2283_b1 , \2286_b1 );
xor ( \2287_b0 , \2283_b0 , w_3756 );
not ( w_3756 , w_3757 );
and ( w_3757 , \2286_b1 , \2286_b0 );
or ( \2288_b1 , \1086_A[4]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_3758 );
and ( \2288_b0 , \1086_A[4]_b0 , w_3759 );
and ( w_3758 , w_3759 , \1654_B[9]_b0 );
or ( \2289_b1 , \2287_b1 , \2288_b1 );
xor ( \2289_b0 , \2287_b0 , w_3760 );
not ( w_3760 , w_3761 );
and ( w_3761 , \2288_b1 , \2288_b0 );
or ( \2290_b1 , \2111_b1 , \2112_b1 );
not ( \2112_b1 , w_3762 );
and ( \2290_b0 , \2111_b0 , w_3763 );
and ( w_3762 , w_3763 , \2112_b0 );
or ( \2291_b1 , \2113_b1 , \2116_b1 );
not ( \2116_b1 , w_3764 );
and ( \2291_b0 , \2113_b0 , w_3765 );
and ( w_3764 , w_3765 , \2116_b0 );
or ( \2292_b1 , \2290_b1 , w_3766 );
or ( \2292_b0 , \2290_b0 , \2291_b0 );
not ( \2291_b0 , w_3767 );
and ( w_3767 , w_3766 , \2291_b1 );
or ( \2293_b1 , \2289_b1 , \2292_b1 );
xor ( \2293_b0 , \2289_b0 , w_3768 );
not ( w_3768 , w_3769 );
and ( w_3769 , \2292_b1 , \2292_b0 );
or ( \2294_b1 , \1018_A[3]_b1 , \1800_B[10]_b1 );
not ( \1800_B[10]_b1 , w_3770 );
and ( \2294_b0 , \1018_A[3]_b0 , w_3771 );
and ( w_3770 , w_3771 , \1800_B[10]_b0 );
or ( \2295_b1 , \2293_b1 , \2294_b1 );
xor ( \2295_b0 , \2293_b0 , w_3772 );
not ( w_3772 , w_3773 );
and ( w_3773 , \2294_b1 , \2294_b0 );
or ( \2296_b1 , \2117_b1 , \2118_b1 );
not ( \2118_b1 , w_3774 );
and ( \2296_b0 , \2117_b0 , w_3775 );
and ( w_3774 , w_3775 , \2118_b0 );
or ( \2297_b1 , \2119_b1 , \2122_b1 );
not ( \2122_b1 , w_3776 );
and ( \2297_b0 , \2119_b0 , w_3777 );
and ( w_3776 , w_3777 , \2122_b0 );
or ( \2298_b1 , \2296_b1 , w_3778 );
or ( \2298_b0 , \2296_b0 , \2297_b0 );
not ( \2297_b0 , w_3779 );
and ( w_3779 , w_3778 , \2297_b1 );
or ( \2299_b1 , \2295_b1 , \2298_b1 );
xor ( \2299_b0 , \2295_b0 , w_3780 );
not ( w_3780 , w_3781 );
and ( w_3781 , \2298_b1 , \2298_b0 );
or ( \2300_b1 , \962_A[2]_b1 , \1958_B[11]_b1 );
not ( \1958_B[11]_b1 , w_3782 );
and ( \2300_b0 , \962_A[2]_b0 , w_3783 );
and ( w_3782 , w_3783 , \1958_B[11]_b0 );
or ( \2301_b1 , \2299_b1 , \2300_b1 );
xor ( \2301_b0 , \2299_b0 , w_3784 );
not ( w_3784 , w_3785 );
and ( w_3785 , \2300_b1 , \2300_b0 );
or ( \2302_b1 , \2123_b1 , \2124_b1 );
not ( \2124_b1 , w_3786 );
and ( \2302_b0 , \2123_b0 , w_3787 );
and ( w_3786 , w_3787 , \2124_b0 );
or ( \2303_b1 , \2125_b1 , \2126_b1 );
not ( \2126_b1 , w_3788 );
and ( \2303_b0 , \2125_b0 , w_3789 );
and ( w_3788 , w_3789 , \2126_b0 );
or ( \2304_b1 , \2302_b1 , w_3790 );
or ( \2304_b0 , \2302_b0 , \2303_b0 );
not ( \2303_b0 , w_3791 );
and ( w_3791 , w_3790 , \2303_b1 );
or ( \2305_b1 , \2301_b1 , \2304_b1 );
xor ( \2305_b0 , \2301_b0 , w_3792 );
not ( w_3792 , w_3793 );
and ( w_3793 , \2304_b1 , \2304_b0 );
or ( \2306_b1 , \920_A[1]_b1 , \2128_B[12]_b1 );
not ( \2128_B[12]_b1 , w_3794 );
and ( \2306_b0 , \920_A[1]_b0 , w_3795 );
and ( w_3794 , w_3795 , \2128_B[12]_b0 );
or ( \2307_b1 , \2305_b1 , \2306_b1 );
xor ( \2307_b0 , \2305_b0 , w_3796 );
not ( w_3796 , w_3797 );
and ( w_3797 , \2306_b1 , \2306_b0 );
or ( \2308_b1 , \2127_b1 , \2129_b1 );
not ( \2129_b1 , w_3798 );
and ( \2308_b0 , \2127_b0 , w_3799 );
and ( w_3798 , w_3799 , \2129_b0 );
or ( \2309_b1 , \2307_b1 , \2308_b1 );
xor ( \2309_b0 , \2307_b0 , w_3800 );
not ( w_3800 , w_3801 );
and ( w_3801 , \2308_b1 , \2308_b0 );
buf ( \2310_B[13]_b1 , \c[13]_b1 );
buf ( \2310_B[13]_b0 , \c[13]_b0 );
or ( \2311_b1 , \886_A[0]_b1 , \2310_B[13]_b1 );
not ( \2310_B[13]_b1 , w_3802 );
and ( \2311_b0 , \886_A[0]_b0 , w_3803 );
and ( w_3802 , w_3803 , \2310_B[13]_b0 );
or ( \2312_b1 , \2309_b1 , \2311_b1 );
xor ( \2312_b0 , \2309_b0 , w_3804 );
not ( w_3804 , w_3805 );
and ( w_3805 , \2311_b1 , \2311_b0 );
buf ( \2313_Z[13]_b1 , \2312_b1 );
buf ( \2313_Z[13]_b0 , \2312_b0 );
or ( \2314_b1 , \2313_Z[13]_b1 , \867_b1 );
not ( \867_b1 , w_3806 );
and ( \2314_b0 , \2313_Z[13]_b0 , w_3807 );
and ( w_3806 , w_3807 , \867_b0 );
buf ( \2315_A[13]_b1 , \a[13]_b1 );
buf ( \2315_A[13]_b0 , \a[13]_b0 );
or ( \2316_b1 , \2315_A[13]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_3808 );
and ( \2316_b0 , \2315_A[13]_b0 , w_3809 );
and ( w_3808 , w_3809 , \892_B[0]_b0 );
or ( \2317_b1 , \2133_A[12]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_3810 );
and ( \2317_b0 , \2133_A[12]_b0 , w_3811 );
and ( w_3810 , w_3811 , \929_B[1]_b0 );
or ( \2318_b1 , \2316_b1 , \2317_b1 );
xor ( \2318_b0 , \2316_b0 , w_3812 );
not ( w_3812 , w_3813 );
and ( w_3813 , \2317_b1 , \2317_b0 );
or ( \2319_b1 , \2134_b1 , \2135_b1 );
not ( \2135_b1 , w_3814 );
and ( \2319_b0 , \2134_b0 , w_3815 );
and ( w_3814 , w_3815 , \2135_b0 );
or ( \2320_b1 , \2136_b1 , \2139_b1 );
not ( \2139_b1 , w_3816 );
and ( \2320_b0 , \2136_b0 , w_3817 );
and ( w_3816 , w_3817 , \2139_b0 );
or ( \2321_b1 , \2319_b1 , w_3818 );
or ( \2321_b0 , \2319_b0 , \2320_b0 );
not ( \2320_b0 , w_3819 );
and ( w_3819 , w_3818 , \2320_b1 );
or ( \2322_b1 , \2318_b1 , \2321_b1 );
xor ( \2322_b0 , \2318_b0 , w_3820 );
not ( w_3820 , w_3821 );
and ( w_3821 , \2321_b1 , \2321_b0 );
or ( \2323_b1 , \1963_A[11]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_3822 );
and ( \2323_b0 , \1963_A[11]_b0 , w_3823 );
and ( w_3822 , w_3823 , \979_B[2]_b0 );
or ( \2324_b1 , \2322_b1 , \2323_b1 );
xor ( \2324_b0 , \2322_b0 , w_3824 );
not ( w_3824 , w_3825 );
and ( w_3825 , \2323_b1 , \2323_b0 );
or ( \2325_b1 , \2140_b1 , \2141_b1 );
not ( \2141_b1 , w_3826 );
and ( \2325_b0 , \2140_b0 , w_3827 );
and ( w_3826 , w_3827 , \2141_b0 );
or ( \2326_b1 , \2142_b1 , \2145_b1 );
not ( \2145_b1 , w_3828 );
and ( \2326_b0 , \2142_b0 , w_3829 );
and ( w_3828 , w_3829 , \2145_b0 );
or ( \2327_b1 , \2325_b1 , w_3830 );
or ( \2327_b0 , \2325_b0 , \2326_b0 );
not ( \2326_b0 , w_3831 );
and ( w_3831 , w_3830 , \2326_b1 );
or ( \2328_b1 , \2324_b1 , \2327_b1 );
xor ( \2328_b0 , \2324_b0 , w_3832 );
not ( w_3832 , w_3833 );
and ( w_3833 , \2327_b1 , \2327_b0 );
or ( \2329_b1 , \1805_A[10]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_3834 );
and ( \2329_b0 , \1805_A[10]_b0 , w_3835 );
and ( w_3834 , w_3835 , \1047_B[3]_b0 );
or ( \2330_b1 , \2328_b1 , \2329_b1 );
xor ( \2330_b0 , \2328_b0 , w_3836 );
not ( w_3836 , w_3837 );
and ( w_3837 , \2329_b1 , \2329_b0 );
or ( \2331_b1 , \2146_b1 , \2147_b1 );
not ( \2147_b1 , w_3838 );
and ( \2331_b0 , \2146_b0 , w_3839 );
and ( w_3838 , w_3839 , \2147_b0 );
or ( \2332_b1 , \2148_b1 , \2151_b1 );
not ( \2151_b1 , w_3840 );
and ( \2332_b0 , \2148_b0 , w_3841 );
and ( w_3840 , w_3841 , \2151_b0 );
or ( \2333_b1 , \2331_b1 , w_3842 );
or ( \2333_b0 , \2331_b0 , \2332_b0 );
not ( \2332_b0 , w_3843 );
and ( w_3843 , w_3842 , \2332_b1 );
or ( \2334_b1 , \2330_b1 , \2333_b1 );
xor ( \2334_b0 , \2330_b0 , w_3844 );
not ( w_3844 , w_3845 );
and ( w_3845 , \2333_b1 , \2333_b0 );
or ( \2335_b1 , \1659_A[9]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_3846 );
and ( \2335_b0 , \1659_A[9]_b0 , w_3847 );
and ( w_3846 , w_3847 , \1127_B[4]_b0 );
or ( \2336_b1 , \2334_b1 , \2335_b1 );
xor ( \2336_b0 , \2334_b0 , w_3848 );
not ( w_3848 , w_3849 );
and ( w_3849 , \2335_b1 , \2335_b0 );
or ( \2337_b1 , \2152_b1 , \2153_b1 );
not ( \2153_b1 , w_3850 );
and ( \2337_b0 , \2152_b0 , w_3851 );
and ( w_3850 , w_3851 , \2153_b0 );
or ( \2338_b1 , \2154_b1 , \2157_b1 );
not ( \2157_b1 , w_3852 );
and ( \2338_b0 , \2154_b0 , w_3853 );
and ( w_3852 , w_3853 , \2157_b0 );
or ( \2339_b1 , \2337_b1 , w_3854 );
or ( \2339_b0 , \2337_b0 , \2338_b0 );
not ( \2338_b0 , w_3855 );
and ( w_3855 , w_3854 , \2338_b1 );
or ( \2340_b1 , \2336_b1 , \2339_b1 );
xor ( \2340_b0 , \2336_b0 , w_3856 );
not ( w_3856 , w_3857 );
and ( w_3857 , \2339_b1 , \2339_b0 );
or ( \2341_b1 , \1525_A[8]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_3858 );
and ( \2341_b0 , \1525_A[8]_b0 , w_3859 );
and ( w_3858 , w_3859 , \1219_B[5]_b0 );
or ( \2342_b1 , \2340_b1 , \2341_b1 );
xor ( \2342_b0 , \2340_b0 , w_3860 );
not ( w_3860 , w_3861 );
and ( w_3861 , \2341_b1 , \2341_b0 );
or ( \2343_b1 , \2158_b1 , \2159_b1 );
not ( \2159_b1 , w_3862 );
and ( \2343_b0 , \2158_b0 , w_3863 );
and ( w_3862 , w_3863 , \2159_b0 );
or ( \2344_b1 , \2160_b1 , \2163_b1 );
not ( \2163_b1 , w_3864 );
and ( \2344_b0 , \2160_b0 , w_3865 );
and ( w_3864 , w_3865 , \2163_b0 );
or ( \2345_b1 , \2343_b1 , w_3866 );
or ( \2345_b0 , \2343_b0 , \2344_b0 );
not ( \2344_b0 , w_3867 );
and ( w_3867 , w_3866 , \2344_b1 );
or ( \2346_b1 , \2342_b1 , \2345_b1 );
xor ( \2346_b0 , \2342_b0 , w_3868 );
not ( w_3868 , w_3869 );
and ( w_3869 , \2345_b1 , \2345_b0 );
or ( \2347_b1 , \1403_A[7]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_3870 );
and ( \2347_b0 , \1403_A[7]_b0 , w_3871 );
and ( w_3870 , w_3871 , \1323_B[6]_b0 );
or ( \2348_b1 , \2346_b1 , \2347_b1 );
xor ( \2348_b0 , \2346_b0 , w_3872 );
not ( w_3872 , w_3873 );
and ( w_3873 , \2347_b1 , \2347_b0 );
or ( \2349_b1 , \2164_b1 , \2165_b1 );
not ( \2165_b1 , w_3874 );
and ( \2349_b0 , \2164_b0 , w_3875 );
and ( w_3874 , w_3875 , \2165_b0 );
or ( \2350_b1 , \2166_b1 , \2169_b1 );
not ( \2169_b1 , w_3876 );
and ( \2350_b0 , \2166_b0 , w_3877 );
and ( w_3876 , w_3877 , \2169_b0 );
or ( \2351_b1 , \2349_b1 , w_3878 );
or ( \2351_b0 , \2349_b0 , \2350_b0 );
not ( \2350_b0 , w_3879 );
and ( w_3879 , w_3878 , \2350_b1 );
or ( \2352_b1 , \2348_b1 , \2351_b1 );
xor ( \2352_b0 , \2348_b0 , w_3880 );
not ( w_3880 , w_3881 );
and ( w_3881 , \2351_b1 , \2351_b0 );
or ( \2353_b1 , \1293_A[6]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_3882 );
and ( \2353_b0 , \1293_A[6]_b0 , w_3883 );
and ( w_3882 , w_3883 , \1439_B[7]_b0 );
or ( \2354_b1 , \2352_b1 , \2353_b1 );
xor ( \2354_b0 , \2352_b0 , w_3884 );
not ( w_3884 , w_3885 );
and ( w_3885 , \2353_b1 , \2353_b0 );
or ( \2355_b1 , \2170_b1 , \2171_b1 );
not ( \2171_b1 , w_3886 );
and ( \2355_b0 , \2170_b0 , w_3887 );
and ( w_3886 , w_3887 , \2171_b0 );
or ( \2356_b1 , \2172_b1 , \2175_b1 );
not ( \2175_b1 , w_3888 );
and ( \2356_b0 , \2172_b0 , w_3889 );
and ( w_3888 , w_3889 , \2175_b0 );
or ( \2357_b1 , \2355_b1 , w_3890 );
or ( \2357_b0 , \2355_b0 , \2356_b0 );
not ( \2356_b0 , w_3891 );
and ( w_3891 , w_3890 , \2356_b1 );
or ( \2358_b1 , \2354_b1 , \2357_b1 );
xor ( \2358_b0 , \2354_b0 , w_3892 );
not ( w_3892 , w_3893 );
and ( w_3893 , \2357_b1 , \2357_b0 );
or ( \2359_b1 , \1195_A[5]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_3894 );
and ( \2359_b0 , \1195_A[5]_b0 , w_3895 );
and ( w_3894 , w_3895 , \1567_B[8]_b0 );
or ( \2360_b1 , \2358_b1 , \2359_b1 );
xor ( \2360_b0 , \2358_b0 , w_3896 );
not ( w_3896 , w_3897 );
and ( w_3897 , \2359_b1 , \2359_b0 );
or ( \2361_b1 , \2176_b1 , \2177_b1 );
not ( \2177_b1 , w_3898 );
and ( \2361_b0 , \2176_b0 , w_3899 );
and ( w_3898 , w_3899 , \2177_b0 );
or ( \2362_b1 , \2178_b1 , \2181_b1 );
not ( \2181_b1 , w_3900 );
and ( \2362_b0 , \2178_b0 , w_3901 );
and ( w_3900 , w_3901 , \2181_b0 );
or ( \2363_b1 , \2361_b1 , w_3902 );
or ( \2363_b0 , \2361_b0 , \2362_b0 );
not ( \2362_b0 , w_3903 );
and ( w_3903 , w_3902 , \2362_b1 );
or ( \2364_b1 , \2360_b1 , \2363_b1 );
xor ( \2364_b0 , \2360_b0 , w_3904 );
not ( w_3904 , w_3905 );
and ( w_3905 , \2363_b1 , \2363_b0 );
or ( \2365_b1 , \1109_A[4]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_3906 );
and ( \2365_b0 , \1109_A[4]_b0 , w_3907 );
and ( w_3906 , w_3907 , \1707_B[9]_b0 );
or ( \2366_b1 , \2364_b1 , \2365_b1 );
xor ( \2366_b0 , \2364_b0 , w_3908 );
not ( w_3908 , w_3909 );
and ( w_3909 , \2365_b1 , \2365_b0 );
or ( \2367_b1 , \2182_b1 , \2183_b1 );
not ( \2183_b1 , w_3910 );
and ( \2367_b0 , \2182_b0 , w_3911 );
and ( w_3910 , w_3911 , \2183_b0 );
or ( \2368_b1 , \2184_b1 , \2187_b1 );
not ( \2187_b1 , w_3912 );
and ( \2368_b0 , \2184_b0 , w_3913 );
and ( w_3912 , w_3913 , \2187_b0 );
or ( \2369_b1 , \2367_b1 , w_3914 );
or ( \2369_b0 , \2367_b0 , \2368_b0 );
not ( \2368_b0 , w_3915 );
and ( w_3915 , w_3914 , \2368_b1 );
or ( \2370_b1 , \2366_b1 , \2369_b1 );
xor ( \2370_b0 , \2366_b0 , w_3916 );
not ( w_3916 , w_3917 );
and ( w_3917 , \2369_b1 , \2369_b0 );
or ( \2371_b1 , \1035_A[3]_b1 , \1859_B[10]_b1 );
not ( \1859_B[10]_b1 , w_3918 );
and ( \2371_b0 , \1035_A[3]_b0 , w_3919 );
and ( w_3918 , w_3919 , \1859_B[10]_b0 );
or ( \2372_b1 , \2370_b1 , \2371_b1 );
xor ( \2372_b0 , \2370_b0 , w_3920 );
not ( w_3920 , w_3921 );
and ( w_3921 , \2371_b1 , \2371_b0 );
or ( \2373_b1 , \2188_b1 , \2189_b1 );
not ( \2189_b1 , w_3922 );
and ( \2373_b0 , \2188_b0 , w_3923 );
and ( w_3922 , w_3923 , \2189_b0 );
or ( \2374_b1 , \2190_b1 , \2193_b1 );
not ( \2193_b1 , w_3924 );
and ( \2374_b0 , \2190_b0 , w_3925 );
and ( w_3924 , w_3925 , \2193_b0 );
or ( \2375_b1 , \2373_b1 , w_3926 );
or ( \2375_b0 , \2373_b0 , \2374_b0 );
not ( \2374_b0 , w_3927 );
and ( w_3927 , w_3926 , \2374_b1 );
or ( \2376_b1 , \2372_b1 , \2375_b1 );
xor ( \2376_b0 , \2372_b0 , w_3928 );
not ( w_3928 , w_3929 );
and ( w_3929 , \2375_b1 , \2375_b0 );
or ( \2377_b1 , \973_A[2]_b1 , \2023_B[11]_b1 );
not ( \2023_B[11]_b1 , w_3930 );
and ( \2377_b0 , \973_A[2]_b0 , w_3931 );
and ( w_3930 , w_3931 , \2023_B[11]_b0 );
or ( \2378_b1 , \2376_b1 , \2377_b1 );
xor ( \2378_b0 , \2376_b0 , w_3932 );
not ( w_3932 , w_3933 );
and ( w_3933 , \2377_b1 , \2377_b0 );
or ( \2379_b1 , \2194_b1 , \2195_b1 );
not ( \2195_b1 , w_3934 );
and ( \2379_b0 , \2194_b0 , w_3935 );
and ( w_3934 , w_3935 , \2195_b0 );
or ( \2380_b1 , \2196_b1 , \2197_b1 );
not ( \2197_b1 , w_3936 );
and ( \2380_b0 , \2196_b0 , w_3937 );
and ( w_3936 , w_3937 , \2197_b0 );
or ( \2381_b1 , \2379_b1 , w_3938 );
or ( \2381_b0 , \2379_b0 , \2380_b0 );
not ( \2380_b0 , w_3939 );
and ( w_3939 , w_3938 , \2380_b1 );
or ( \2382_b1 , \2378_b1 , \2381_b1 );
xor ( \2382_b0 , \2378_b0 , w_3940 );
not ( w_3940 , w_3941 );
and ( w_3941 , \2381_b1 , \2381_b0 );
or ( \2383_b1 , \927_A[1]_b1 , \2199_B[12]_b1 );
not ( \2199_B[12]_b1 , w_3942 );
and ( \2383_b0 , \927_A[1]_b0 , w_3943 );
and ( w_3942 , w_3943 , \2199_B[12]_b0 );
or ( \2384_b1 , \2382_b1 , \2383_b1 );
xor ( \2384_b0 , \2382_b0 , w_3944 );
not ( w_3944 , w_3945 );
and ( w_3945 , \2383_b1 , \2383_b0 );
or ( \2385_b1 , \2198_b1 , \2200_b1 );
not ( \2200_b1 , w_3946 );
and ( \2385_b0 , \2198_b0 , w_3947 );
and ( w_3946 , w_3947 , \2200_b0 );
or ( \2386_b1 , \2384_b1 , \2385_b1 );
xor ( \2386_b0 , \2384_b0 , w_3948 );
not ( w_3948 , w_3949 );
and ( w_3949 , \2385_b1 , \2385_b0 );
buf ( \2387_B[13]_b1 , \d[13]_b1 );
buf ( \2387_B[13]_b0 , \d[13]_b0 );
or ( \2388_b1 , \891_A[0]_b1 , \2387_B[13]_b1 );
not ( \2387_B[13]_b1 , w_3950 );
and ( \2388_b0 , \891_A[0]_b0 , w_3951 );
and ( w_3950 , w_3951 , \2387_B[13]_b0 );
or ( \2389_b1 , \2386_b1 , \2388_b1 );
xor ( \2389_b0 , \2386_b0 , w_3952 );
not ( w_3952 , w_3953 );
and ( w_3953 , \2388_b1 , \2388_b0 );
buf ( \2390_Z[13]_b1 , \2389_b1 );
buf ( \2390_Z[13]_b0 , \2389_b0 );
or ( \2391_b1 , \2390_Z[13]_b1 , \865_b1 );
not ( \865_b1 , w_3954 );
and ( \2391_b0 , \2390_Z[13]_b0 , w_3955 );
and ( w_3954 , w_3955 , \865_b0 );
buf ( \2392_A[13]_b1 , \b[13]_b1 );
buf ( \2392_A[13]_b0 , \b[13]_b0 );
buf ( \2393_B[13]_b1 , \d[13]_b1 );
buf ( \2393_B[13]_b0 , \d[13]_b0 );
or ( \2394_b1 , \2392_A[13]_b1 , \2393_B[13]_b1 );
xor ( \2394_b0 , \2392_A[13]_b0 , w_3956 );
not ( w_3956 , w_3957 );
and ( w_3957 , \2393_B[13]_b1 , \2393_B[13]_b0 );
or ( \2395_b1 , \2204_A[12]_b1 , \2205_B[12]_b1 );
not ( \2205_B[12]_b1 , w_3958 );
and ( \2395_b0 , \2204_A[12]_b0 , w_3959 );
and ( w_3958 , w_3959 , \2205_B[12]_b0 );
or ( \2396_b1 , \2205_B[12]_b1 , \2210_b1 );
not ( \2210_b1 , w_3960 );
and ( \2396_b0 , \2205_B[12]_b0 , w_3961 );
and ( w_3960 , w_3961 , \2210_b0 );
or ( \2397_b1 , \2204_A[12]_b1 , \2210_b1 );
not ( \2210_b1 , w_3962 );
and ( \2397_b0 , \2204_A[12]_b0 , w_3963 );
and ( w_3962 , w_3963 , \2210_b0 );
or ( \2399_b1 , \2394_b1 , \2398_b1 );
xor ( \2399_b0 , \2394_b0 , w_3964 );
not ( w_3964 , w_3965 );
and ( w_3965 , \2398_b1 , \2398_b0 );
buf ( \2400_SUM[13]_b1 , \2399_b1 );
buf ( \2400_SUM[13]_b0 , \2399_b0 );
or ( \2401_b1 , \2400_SUM[13]_b1 , \863_b1 );
not ( \863_b1 , w_3966 );
and ( \2401_b0 , \2400_SUM[13]_b0 , w_3967 );
and ( w_3966 , w_3967 , \863_b0 );
buf ( \2402_A[13]_b1 , \a[13]_b1 );
buf ( \2402_A[13]_b0 , \a[13]_b0 );
buf ( \2403_B[13]_b1 , \c[13]_b1 );
buf ( \2403_B[13]_b0 , \c[13]_b0 );
or ( \2404_b1 , \2402_A[13]_b1 , \2403_B[13]_b1 );
xor ( \2404_b0 , \2402_A[13]_b0 , w_3968 );
not ( w_3968 , w_3969 );
and ( w_3969 , \2403_B[13]_b1 , \2403_B[13]_b0 );
or ( \2405_b1 , \2214_A[12]_b1 , \2215_B[12]_b1 );
not ( \2215_B[12]_b1 , w_3970 );
and ( \2405_b0 , \2214_A[12]_b0 , w_3971 );
and ( w_3970 , w_3971 , \2215_B[12]_b0 );
or ( \2406_b1 , \2215_B[12]_b1 , \2220_b1 );
not ( \2220_b1 , w_3972 );
and ( \2406_b0 , \2215_B[12]_b0 , w_3973 );
and ( w_3972 , w_3973 , \2220_b0 );
or ( \2407_b1 , \2214_A[12]_b1 , \2220_b1 );
not ( \2220_b1 , w_3974 );
and ( \2407_b0 , \2214_A[12]_b0 , w_3975 );
and ( w_3974 , w_3975 , \2220_b0 );
or ( \2409_b1 , \2404_b1 , \2408_b1 );
xor ( \2409_b0 , \2404_b0 , w_3976 );
not ( w_3976 , w_3977 );
and ( w_3977 , \2408_b1 , \2408_b0 );
buf ( \2410_SUM[13]_b1 , \2409_b1 );
buf ( \2410_SUM[13]_b0 , \2409_b0 );
or ( \2411_b1 , \2410_SUM[13]_b1 , \861_b1 );
not ( \861_b1 , w_3978 );
and ( \2411_b0 , \2410_SUM[13]_b0 , w_3979 );
and ( w_3978 , w_3979 , \861_b0 );
or ( \2412_b1 , \d[13]_b1 , \859_b1 );
not ( \859_b1 , w_3980 );
and ( \2412_b0 , \d[13]_b0 , w_3981 );
and ( w_3980 , w_3981 , \859_b0 );
or ( \2413_b1 , \c[13]_b1 , \857_b1 );
not ( \857_b1 , w_3982 );
and ( \2413_b0 , \c[13]_b0 , w_3983 );
and ( w_3982 , w_3983 , \857_b0 );
or ( \2414_b1 , \b[13]_b1 , \855_b1 );
not ( \855_b1 , w_3984 );
and ( \2414_b0 , \b[13]_b0 , w_3985 );
and ( w_3984 , w_3985 , \855_b0 );
or ( \2415_b1 , \a[13]_b1 , \853_b1 );
not ( \853_b1 , w_3986 );
and ( \2415_b0 , \a[13]_b0 , w_3987 );
and ( w_3986 , w_3987 , \853_b0 );
and ( \2417_b1 , 1'b0_b1 , w_3988 );
xor ( w_3988 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_3989 );
and ( \2417_b0 , w_3989 , \876_b0 );
or ( \2418_b1 , \a[14]_b1 , w_3990 );
or ( \2418_b0 , \a[14]_b0 , \d[14]_b0 );
not ( \d[14]_b0 , w_3991 );
and ( w_3991 , w_3990 , \d[14]_b1 );
or ( \2419_b1 , \2418_b1 , \875_b1 );
not ( \875_b1 , w_3992 );
and ( \2419_b0 , \2418_b0 , w_3993 );
and ( w_3992 , w_3993 , \875_b0 );
or ( \2420_b1 , \b[14]_b1 , \c[14]_b1 );
not ( \c[14]_b1 , w_3994 );
and ( \2420_b0 , \b[14]_b0 , w_3995 );
and ( w_3994 , w_3995 , \c[14]_b0 );
or ( \2421_b1 , \2420_b1 , \873_b1 );
not ( \873_b1 , w_3996 );
and ( \2421_b0 , \2420_b0 , w_3997 );
and ( w_3996 , w_3997 , \873_b0 );
or ( \2422_b1 , \a[14]_b1 , w_3998 );
or ( \2422_b0 , \a[14]_b0 , \b[14]_b0 );
not ( \b[14]_b0 , w_3999 );
and ( w_3999 , w_3998 , \b[14]_b1 );
or ( \2423_b1 , \2422_b1 , \871_b1 );
not ( \871_b1 , w_4000 );
and ( \2423_b0 , \2422_b0 , w_4001 );
and ( w_4000 , w_4001 , \871_b0 );
or ( \2424_b1 , \c[14]_b1 , \d[14]_b1 );
xor ( \2424_b0 , \c[14]_b0 , w_4002 );
not ( w_4002 , w_4003 );
and ( w_4003 , \d[14]_b1 , \d[14]_b0 );
or ( \2425_b1 , \2424_b1 , \869_b1 );
not ( \869_b1 , w_4004 );
and ( \2425_b0 , \2424_b0 , w_4005 );
and ( w_4004 , w_4005 , \869_b0 );
buf ( \2426_A[14]_b1 , \b[14]_b1 );
buf ( \2426_A[14]_b0 , \b[14]_b0 );
or ( \2427_b1 , \2426_A[14]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_4006 );
and ( \2427_b0 , \2426_A[14]_b0 , w_4007 );
and ( w_4006 , w_4007 , \887_B[0]_b0 );
or ( \2428_b1 , \2238_A[13]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_4008 );
and ( \2428_b0 , \2238_A[13]_b0 , w_4009 );
and ( w_4008 , w_4009 , \922_B[1]_b0 );
or ( \2429_b1 , \2427_b1 , \2428_b1 );
xor ( \2429_b0 , \2427_b0 , w_4010 );
not ( w_4010 , w_4011 );
and ( w_4011 , \2428_b1 , \2428_b0 );
or ( \2430_b1 , \2239_b1 , \2240_b1 );
not ( \2240_b1 , w_4012 );
and ( \2430_b0 , \2239_b0 , w_4013 );
and ( w_4012 , w_4013 , \2240_b0 );
or ( \2431_b1 , \2241_b1 , \2244_b1 );
not ( \2244_b1 , w_4014 );
and ( \2431_b0 , \2241_b0 , w_4015 );
and ( w_4014 , w_4015 , \2244_b0 );
or ( \2432_b1 , \2430_b1 , w_4016 );
or ( \2432_b0 , \2430_b0 , \2431_b0 );
not ( \2431_b0 , w_4017 );
and ( w_4017 , w_4016 , \2431_b1 );
or ( \2433_b1 , \2429_b1 , \2432_b1 );
xor ( \2433_b0 , \2429_b0 , w_4018 );
not ( w_4018 , w_4019 );
and ( w_4019 , \2432_b1 , \2432_b0 );
or ( \2434_b1 , \2062_A[12]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_4020 );
and ( \2434_b0 , \2062_A[12]_b0 , w_4021 );
and ( w_4020 , w_4021 , \968_B[2]_b0 );
or ( \2435_b1 , \2433_b1 , \2434_b1 );
xor ( \2435_b0 , \2433_b0 , w_4022 );
not ( w_4022 , w_4023 );
and ( w_4023 , \2434_b1 , \2434_b0 );
or ( \2436_b1 , \2245_b1 , \2246_b1 );
not ( \2246_b1 , w_4024 );
and ( \2436_b0 , \2245_b0 , w_4025 );
and ( w_4024 , w_4025 , \2246_b0 );
or ( \2437_b1 , \2247_b1 , \2250_b1 );
not ( \2250_b1 , w_4026 );
and ( \2437_b0 , \2247_b0 , w_4027 );
and ( w_4026 , w_4027 , \2250_b0 );
or ( \2438_b1 , \2436_b1 , w_4028 );
or ( \2438_b0 , \2436_b0 , \2437_b0 );
not ( \2437_b0 , w_4029 );
and ( w_4029 , w_4028 , \2437_b1 );
or ( \2439_b1 , \2435_b1 , \2438_b1 );
xor ( \2439_b0 , \2435_b0 , w_4030 );
not ( w_4030 , w_4031 );
and ( w_4031 , \2438_b1 , \2438_b0 );
or ( \2440_b1 , \1898_A[11]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_4032 );
and ( \2440_b0 , \1898_A[11]_b0 , w_4033 );
and ( w_4032 , w_4033 , \1030_B[3]_b0 );
or ( \2441_b1 , \2439_b1 , \2440_b1 );
xor ( \2441_b0 , \2439_b0 , w_4034 );
not ( w_4034 , w_4035 );
and ( w_4035 , \2440_b1 , \2440_b0 );
or ( \2442_b1 , \2251_b1 , \2252_b1 );
not ( \2252_b1 , w_4036 );
and ( \2442_b0 , \2251_b0 , w_4037 );
and ( w_4036 , w_4037 , \2252_b0 );
or ( \2443_b1 , \2253_b1 , \2256_b1 );
not ( \2256_b1 , w_4038 );
and ( \2443_b0 , \2253_b0 , w_4039 );
and ( w_4038 , w_4039 , \2256_b0 );
or ( \2444_b1 , \2442_b1 , w_4040 );
or ( \2444_b0 , \2442_b0 , \2443_b0 );
not ( \2443_b0 , w_4041 );
and ( w_4041 , w_4040 , \2443_b1 );
or ( \2445_b1 , \2441_b1 , \2444_b1 );
xor ( \2445_b0 , \2441_b0 , w_4042 );
not ( w_4042 , w_4043 );
and ( w_4043 , \2444_b1 , \2444_b0 );
or ( \2446_b1 , \1746_A[10]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_4044 );
and ( \2446_b0 , \1746_A[10]_b0 , w_4045 );
and ( w_4044 , w_4045 , \1104_B[4]_b0 );
or ( \2447_b1 , \2445_b1 , \2446_b1 );
xor ( \2447_b0 , \2445_b0 , w_4046 );
not ( w_4046 , w_4047 );
and ( w_4047 , \2446_b1 , \2446_b0 );
or ( \2448_b1 , \2257_b1 , \2258_b1 );
not ( \2258_b1 , w_4048 );
and ( \2448_b0 , \2257_b0 , w_4049 );
and ( w_4048 , w_4049 , \2258_b0 );
or ( \2449_b1 , \2259_b1 , \2262_b1 );
not ( \2262_b1 , w_4050 );
and ( \2449_b0 , \2259_b0 , w_4051 );
and ( w_4050 , w_4051 , \2262_b0 );
or ( \2450_b1 , \2448_b1 , w_4052 );
or ( \2450_b0 , \2448_b0 , \2449_b0 );
not ( \2449_b0 , w_4053 );
and ( w_4053 , w_4052 , \2449_b1 );
or ( \2451_b1 , \2447_b1 , \2450_b1 );
xor ( \2451_b0 , \2447_b0 , w_4054 );
not ( w_4054 , w_4055 );
and ( w_4055 , \2450_b1 , \2450_b0 );
or ( \2452_b1 , \1606_A[9]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_4056 );
and ( \2452_b0 , \1606_A[9]_b0 , w_4057 );
and ( w_4056 , w_4057 , \1190_B[5]_b0 );
or ( \2453_b1 , \2451_b1 , \2452_b1 );
xor ( \2453_b0 , \2451_b0 , w_4058 );
not ( w_4058 , w_4059 );
and ( w_4059 , \2452_b1 , \2452_b0 );
or ( \2454_b1 , \2263_b1 , \2264_b1 );
not ( \2264_b1 , w_4060 );
and ( \2454_b0 , \2263_b0 , w_4061 );
and ( w_4060 , w_4061 , \2264_b0 );
or ( \2455_b1 , \2265_b1 , \2268_b1 );
not ( \2268_b1 , w_4062 );
and ( \2455_b0 , \2265_b0 , w_4063 );
and ( w_4062 , w_4063 , \2268_b0 );
or ( \2456_b1 , \2454_b1 , w_4064 );
or ( \2456_b0 , \2454_b0 , \2455_b0 );
not ( \2455_b0 , w_4065 );
and ( w_4065 , w_4064 , \2455_b1 );
or ( \2457_b1 , \2453_b1 , \2456_b1 );
xor ( \2457_b0 , \2453_b0 , w_4066 );
not ( w_4066 , w_4067 );
and ( w_4067 , \2456_b1 , \2456_b0 );
or ( \2458_b1 , \1478_A[8]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_4068 );
and ( \2458_b0 , \1478_A[8]_b0 , w_4069 );
and ( w_4068 , w_4069 , \1288_B[6]_b0 );
or ( \2459_b1 , \2457_b1 , \2458_b1 );
xor ( \2459_b0 , \2457_b0 , w_4070 );
not ( w_4070 , w_4071 );
and ( w_4071 , \2458_b1 , \2458_b0 );
or ( \2460_b1 , \2269_b1 , \2270_b1 );
not ( \2270_b1 , w_4072 );
and ( \2460_b0 , \2269_b0 , w_4073 );
and ( w_4072 , w_4073 , \2270_b0 );
or ( \2461_b1 , \2271_b1 , \2274_b1 );
not ( \2274_b1 , w_4074 );
and ( \2461_b0 , \2271_b0 , w_4075 );
and ( w_4074 , w_4075 , \2274_b0 );
or ( \2462_b1 , \2460_b1 , w_4076 );
or ( \2462_b0 , \2460_b0 , \2461_b0 );
not ( \2461_b0 , w_4077 );
and ( w_4077 , w_4076 , \2461_b1 );
or ( \2463_b1 , \2459_b1 , \2462_b1 );
xor ( \2463_b0 , \2459_b0 , w_4078 );
not ( w_4078 , w_4079 );
and ( w_4079 , \2462_b1 , \2462_b0 );
or ( \2464_b1 , \1362_A[7]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_4080 );
and ( \2464_b0 , \1362_A[7]_b0 , w_4081 );
and ( w_4080 , w_4081 , \1398_B[7]_b0 );
or ( \2465_b1 , \2463_b1 , \2464_b1 );
xor ( \2465_b0 , \2463_b0 , w_4082 );
not ( w_4082 , w_4083 );
and ( w_4083 , \2464_b1 , \2464_b0 );
or ( \2466_b1 , \2275_b1 , \2276_b1 );
not ( \2276_b1 , w_4084 );
and ( \2466_b0 , \2275_b0 , w_4085 );
and ( w_4084 , w_4085 , \2276_b0 );
or ( \2467_b1 , \2277_b1 , \2280_b1 );
not ( \2280_b1 , w_4086 );
and ( \2467_b0 , \2277_b0 , w_4087 );
and ( w_4086 , w_4087 , \2280_b0 );
or ( \2468_b1 , \2466_b1 , w_4088 );
or ( \2468_b0 , \2466_b0 , \2467_b0 );
not ( \2467_b0 , w_4089 );
and ( w_4089 , w_4088 , \2467_b1 );
or ( \2469_b1 , \2465_b1 , \2468_b1 );
xor ( \2469_b0 , \2465_b0 , w_4090 );
not ( w_4090 , w_4091 );
and ( w_4091 , \2468_b1 , \2468_b0 );
or ( \2470_b1 , \1258_A[6]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_4092 );
and ( \2470_b0 , \1258_A[6]_b0 , w_4093 );
and ( w_4092 , w_4093 , \1520_B[8]_b0 );
or ( \2471_b1 , \2469_b1 , \2470_b1 );
xor ( \2471_b0 , \2469_b0 , w_4094 );
not ( w_4094 , w_4095 );
and ( w_4095 , \2470_b1 , \2470_b0 );
or ( \2472_b1 , \2281_b1 , \2282_b1 );
not ( \2282_b1 , w_4096 );
and ( \2472_b0 , \2281_b0 , w_4097 );
and ( w_4096 , w_4097 , \2282_b0 );
or ( \2473_b1 , \2283_b1 , \2286_b1 );
not ( \2286_b1 , w_4098 );
and ( \2473_b0 , \2283_b0 , w_4099 );
and ( w_4098 , w_4099 , \2286_b0 );
or ( \2474_b1 , \2472_b1 , w_4100 );
or ( \2474_b0 , \2472_b0 , \2473_b0 );
not ( \2473_b0 , w_4101 );
and ( w_4101 , w_4100 , \2473_b1 );
or ( \2475_b1 , \2471_b1 , \2474_b1 );
xor ( \2475_b0 , \2471_b0 , w_4102 );
not ( w_4102 , w_4103 );
and ( w_4103 , \2474_b1 , \2474_b0 );
or ( \2476_b1 , \1166_A[5]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_4104 );
and ( \2476_b0 , \1166_A[5]_b0 , w_4105 );
and ( w_4104 , w_4105 , \1654_B[9]_b0 );
or ( \2477_b1 , \2475_b1 , \2476_b1 );
xor ( \2477_b0 , \2475_b0 , w_4106 );
not ( w_4106 , w_4107 );
and ( w_4107 , \2476_b1 , \2476_b0 );
or ( \2478_b1 , \2287_b1 , \2288_b1 );
not ( \2288_b1 , w_4108 );
and ( \2478_b0 , \2287_b0 , w_4109 );
and ( w_4108 , w_4109 , \2288_b0 );
or ( \2479_b1 , \2289_b1 , \2292_b1 );
not ( \2292_b1 , w_4110 );
and ( \2479_b0 , \2289_b0 , w_4111 );
and ( w_4110 , w_4111 , \2292_b0 );
or ( \2480_b1 , \2478_b1 , w_4112 );
or ( \2480_b0 , \2478_b0 , \2479_b0 );
not ( \2479_b0 , w_4113 );
and ( w_4113 , w_4112 , \2479_b1 );
or ( \2481_b1 , \2477_b1 , \2480_b1 );
xor ( \2481_b0 , \2477_b0 , w_4114 );
not ( w_4114 , w_4115 );
and ( w_4115 , \2480_b1 , \2480_b0 );
or ( \2482_b1 , \1086_A[4]_b1 , \1800_B[10]_b1 );
not ( \1800_B[10]_b1 , w_4116 );
and ( \2482_b0 , \1086_A[4]_b0 , w_4117 );
and ( w_4116 , w_4117 , \1800_B[10]_b0 );
or ( \2483_b1 , \2481_b1 , \2482_b1 );
xor ( \2483_b0 , \2481_b0 , w_4118 );
not ( w_4118 , w_4119 );
and ( w_4119 , \2482_b1 , \2482_b0 );
or ( \2484_b1 , \2293_b1 , \2294_b1 );
not ( \2294_b1 , w_4120 );
and ( \2484_b0 , \2293_b0 , w_4121 );
and ( w_4120 , w_4121 , \2294_b0 );
or ( \2485_b1 , \2295_b1 , \2298_b1 );
not ( \2298_b1 , w_4122 );
and ( \2485_b0 , \2295_b0 , w_4123 );
and ( w_4122 , w_4123 , \2298_b0 );
or ( \2486_b1 , \2484_b1 , w_4124 );
or ( \2486_b0 , \2484_b0 , \2485_b0 );
not ( \2485_b0 , w_4125 );
and ( w_4125 , w_4124 , \2485_b1 );
or ( \2487_b1 , \2483_b1 , \2486_b1 );
xor ( \2487_b0 , \2483_b0 , w_4126 );
not ( w_4126 , w_4127 );
and ( w_4127 , \2486_b1 , \2486_b0 );
or ( \2488_b1 , \1018_A[3]_b1 , \1958_B[11]_b1 );
not ( \1958_B[11]_b1 , w_4128 );
and ( \2488_b0 , \1018_A[3]_b0 , w_4129 );
and ( w_4128 , w_4129 , \1958_B[11]_b0 );
or ( \2489_b1 , \2487_b1 , \2488_b1 );
xor ( \2489_b0 , \2487_b0 , w_4130 );
not ( w_4130 , w_4131 );
and ( w_4131 , \2488_b1 , \2488_b0 );
or ( \2490_b1 , \2299_b1 , \2300_b1 );
not ( \2300_b1 , w_4132 );
and ( \2490_b0 , \2299_b0 , w_4133 );
and ( w_4132 , w_4133 , \2300_b0 );
or ( \2491_b1 , \2301_b1 , \2304_b1 );
not ( \2304_b1 , w_4134 );
and ( \2491_b0 , \2301_b0 , w_4135 );
and ( w_4134 , w_4135 , \2304_b0 );
or ( \2492_b1 , \2490_b1 , w_4136 );
or ( \2492_b0 , \2490_b0 , \2491_b0 );
not ( \2491_b0 , w_4137 );
and ( w_4137 , w_4136 , \2491_b1 );
or ( \2493_b1 , \2489_b1 , \2492_b1 );
xor ( \2493_b0 , \2489_b0 , w_4138 );
not ( w_4138 , w_4139 );
and ( w_4139 , \2492_b1 , \2492_b0 );
or ( \2494_b1 , \962_A[2]_b1 , \2128_B[12]_b1 );
not ( \2128_B[12]_b1 , w_4140 );
and ( \2494_b0 , \962_A[2]_b0 , w_4141 );
and ( w_4140 , w_4141 , \2128_B[12]_b0 );
or ( \2495_b1 , \2493_b1 , \2494_b1 );
xor ( \2495_b0 , \2493_b0 , w_4142 );
not ( w_4142 , w_4143 );
and ( w_4143 , \2494_b1 , \2494_b0 );
or ( \2496_b1 , \2305_b1 , \2306_b1 );
not ( \2306_b1 , w_4144 );
and ( \2496_b0 , \2305_b0 , w_4145 );
and ( w_4144 , w_4145 , \2306_b0 );
or ( \2497_b1 , \2307_b1 , \2308_b1 );
not ( \2308_b1 , w_4146 );
and ( \2497_b0 , \2307_b0 , w_4147 );
and ( w_4146 , w_4147 , \2308_b0 );
or ( \2498_b1 , \2496_b1 , w_4148 );
or ( \2498_b0 , \2496_b0 , \2497_b0 );
not ( \2497_b0 , w_4149 );
and ( w_4149 , w_4148 , \2497_b1 );
or ( \2499_b1 , \2495_b1 , \2498_b1 );
xor ( \2499_b0 , \2495_b0 , w_4150 );
not ( w_4150 , w_4151 );
and ( w_4151 , \2498_b1 , \2498_b0 );
or ( \2500_b1 , \920_A[1]_b1 , \2310_B[13]_b1 );
not ( \2310_B[13]_b1 , w_4152 );
and ( \2500_b0 , \920_A[1]_b0 , w_4153 );
and ( w_4152 , w_4153 , \2310_B[13]_b0 );
or ( \2501_b1 , \2499_b1 , \2500_b1 );
xor ( \2501_b0 , \2499_b0 , w_4154 );
not ( w_4154 , w_4155 );
and ( w_4155 , \2500_b1 , \2500_b0 );
or ( \2502_b1 , \2309_b1 , \2311_b1 );
not ( \2311_b1 , w_4156 );
and ( \2502_b0 , \2309_b0 , w_4157 );
and ( w_4156 , w_4157 , \2311_b0 );
or ( \2503_b1 , \2501_b1 , \2502_b1 );
xor ( \2503_b0 , \2501_b0 , w_4158 );
not ( w_4158 , w_4159 );
and ( w_4159 , \2502_b1 , \2502_b0 );
buf ( \2504_B[14]_b1 , \c[14]_b1 );
buf ( \2504_B[14]_b0 , \c[14]_b0 );
or ( \2505_b1 , \886_A[0]_b1 , \2504_B[14]_b1 );
not ( \2504_B[14]_b1 , w_4160 );
and ( \2505_b0 , \886_A[0]_b0 , w_4161 );
and ( w_4160 , w_4161 , \2504_B[14]_b0 );
or ( \2506_b1 , \2503_b1 , \2505_b1 );
xor ( \2506_b0 , \2503_b0 , w_4162 );
not ( w_4162 , w_4163 );
and ( w_4163 , \2505_b1 , \2505_b0 );
buf ( \2507_Z[14]_b1 , \2506_b1 );
buf ( \2507_Z[14]_b0 , \2506_b0 );
or ( \2508_b1 , \2507_Z[14]_b1 , \867_b1 );
not ( \867_b1 , w_4164 );
and ( \2508_b0 , \2507_Z[14]_b0 , w_4165 );
and ( w_4164 , w_4165 , \867_b0 );
buf ( \2509_A[14]_b1 , \a[14]_b1 );
buf ( \2509_A[14]_b0 , \a[14]_b0 );
or ( \2510_b1 , \2509_A[14]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_4166 );
and ( \2510_b0 , \2509_A[14]_b0 , w_4167 );
and ( w_4166 , w_4167 , \892_B[0]_b0 );
or ( \2511_b1 , \2315_A[13]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_4168 );
and ( \2511_b0 , \2315_A[13]_b0 , w_4169 );
and ( w_4168 , w_4169 , \929_B[1]_b0 );
or ( \2512_b1 , \2510_b1 , \2511_b1 );
xor ( \2512_b0 , \2510_b0 , w_4170 );
not ( w_4170 , w_4171 );
and ( w_4171 , \2511_b1 , \2511_b0 );
or ( \2513_b1 , \2316_b1 , \2317_b1 );
not ( \2317_b1 , w_4172 );
and ( \2513_b0 , \2316_b0 , w_4173 );
and ( w_4172 , w_4173 , \2317_b0 );
or ( \2514_b1 , \2318_b1 , \2321_b1 );
not ( \2321_b1 , w_4174 );
and ( \2514_b0 , \2318_b0 , w_4175 );
and ( w_4174 , w_4175 , \2321_b0 );
or ( \2515_b1 , \2513_b1 , w_4176 );
or ( \2515_b0 , \2513_b0 , \2514_b0 );
not ( \2514_b0 , w_4177 );
and ( w_4177 , w_4176 , \2514_b1 );
or ( \2516_b1 , \2512_b1 , \2515_b1 );
xor ( \2516_b0 , \2512_b0 , w_4178 );
not ( w_4178 , w_4179 );
and ( w_4179 , \2515_b1 , \2515_b0 );
or ( \2517_b1 , \2133_A[12]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_4180 );
and ( \2517_b0 , \2133_A[12]_b0 , w_4181 );
and ( w_4180 , w_4181 , \979_B[2]_b0 );
or ( \2518_b1 , \2516_b1 , \2517_b1 );
xor ( \2518_b0 , \2516_b0 , w_4182 );
not ( w_4182 , w_4183 );
and ( w_4183 , \2517_b1 , \2517_b0 );
or ( \2519_b1 , \2322_b1 , \2323_b1 );
not ( \2323_b1 , w_4184 );
and ( \2519_b0 , \2322_b0 , w_4185 );
and ( w_4184 , w_4185 , \2323_b0 );
or ( \2520_b1 , \2324_b1 , \2327_b1 );
not ( \2327_b1 , w_4186 );
and ( \2520_b0 , \2324_b0 , w_4187 );
and ( w_4186 , w_4187 , \2327_b0 );
or ( \2521_b1 , \2519_b1 , w_4188 );
or ( \2521_b0 , \2519_b0 , \2520_b0 );
not ( \2520_b0 , w_4189 );
and ( w_4189 , w_4188 , \2520_b1 );
or ( \2522_b1 , \2518_b1 , \2521_b1 );
xor ( \2522_b0 , \2518_b0 , w_4190 );
not ( w_4190 , w_4191 );
and ( w_4191 , \2521_b1 , \2521_b0 );
or ( \2523_b1 , \1963_A[11]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_4192 );
and ( \2523_b0 , \1963_A[11]_b0 , w_4193 );
and ( w_4192 , w_4193 , \1047_B[3]_b0 );
or ( \2524_b1 , \2522_b1 , \2523_b1 );
xor ( \2524_b0 , \2522_b0 , w_4194 );
not ( w_4194 , w_4195 );
and ( w_4195 , \2523_b1 , \2523_b0 );
or ( \2525_b1 , \2328_b1 , \2329_b1 );
not ( \2329_b1 , w_4196 );
and ( \2525_b0 , \2328_b0 , w_4197 );
and ( w_4196 , w_4197 , \2329_b0 );
or ( \2526_b1 , \2330_b1 , \2333_b1 );
not ( \2333_b1 , w_4198 );
and ( \2526_b0 , \2330_b0 , w_4199 );
and ( w_4198 , w_4199 , \2333_b0 );
or ( \2527_b1 , \2525_b1 , w_4200 );
or ( \2527_b0 , \2525_b0 , \2526_b0 );
not ( \2526_b0 , w_4201 );
and ( w_4201 , w_4200 , \2526_b1 );
or ( \2528_b1 , \2524_b1 , \2527_b1 );
xor ( \2528_b0 , \2524_b0 , w_4202 );
not ( w_4202 , w_4203 );
and ( w_4203 , \2527_b1 , \2527_b0 );
or ( \2529_b1 , \1805_A[10]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_4204 );
and ( \2529_b0 , \1805_A[10]_b0 , w_4205 );
and ( w_4204 , w_4205 , \1127_B[4]_b0 );
or ( \2530_b1 , \2528_b1 , \2529_b1 );
xor ( \2530_b0 , \2528_b0 , w_4206 );
not ( w_4206 , w_4207 );
and ( w_4207 , \2529_b1 , \2529_b0 );
or ( \2531_b1 , \2334_b1 , \2335_b1 );
not ( \2335_b1 , w_4208 );
and ( \2531_b0 , \2334_b0 , w_4209 );
and ( w_4208 , w_4209 , \2335_b0 );
or ( \2532_b1 , \2336_b1 , \2339_b1 );
not ( \2339_b1 , w_4210 );
and ( \2532_b0 , \2336_b0 , w_4211 );
and ( w_4210 , w_4211 , \2339_b0 );
or ( \2533_b1 , \2531_b1 , w_4212 );
or ( \2533_b0 , \2531_b0 , \2532_b0 );
not ( \2532_b0 , w_4213 );
and ( w_4213 , w_4212 , \2532_b1 );
or ( \2534_b1 , \2530_b1 , \2533_b1 );
xor ( \2534_b0 , \2530_b0 , w_4214 );
not ( w_4214 , w_4215 );
and ( w_4215 , \2533_b1 , \2533_b0 );
or ( \2535_b1 , \1659_A[9]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_4216 );
and ( \2535_b0 , \1659_A[9]_b0 , w_4217 );
and ( w_4216 , w_4217 , \1219_B[5]_b0 );
or ( \2536_b1 , \2534_b1 , \2535_b1 );
xor ( \2536_b0 , \2534_b0 , w_4218 );
not ( w_4218 , w_4219 );
and ( w_4219 , \2535_b1 , \2535_b0 );
or ( \2537_b1 , \2340_b1 , \2341_b1 );
not ( \2341_b1 , w_4220 );
and ( \2537_b0 , \2340_b0 , w_4221 );
and ( w_4220 , w_4221 , \2341_b0 );
or ( \2538_b1 , \2342_b1 , \2345_b1 );
not ( \2345_b1 , w_4222 );
and ( \2538_b0 , \2342_b0 , w_4223 );
and ( w_4222 , w_4223 , \2345_b0 );
or ( \2539_b1 , \2537_b1 , w_4224 );
or ( \2539_b0 , \2537_b0 , \2538_b0 );
not ( \2538_b0 , w_4225 );
and ( w_4225 , w_4224 , \2538_b1 );
or ( \2540_b1 , \2536_b1 , \2539_b1 );
xor ( \2540_b0 , \2536_b0 , w_4226 );
not ( w_4226 , w_4227 );
and ( w_4227 , \2539_b1 , \2539_b0 );
or ( \2541_b1 , \1525_A[8]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_4228 );
and ( \2541_b0 , \1525_A[8]_b0 , w_4229 );
and ( w_4228 , w_4229 , \1323_B[6]_b0 );
or ( \2542_b1 , \2540_b1 , \2541_b1 );
xor ( \2542_b0 , \2540_b0 , w_4230 );
not ( w_4230 , w_4231 );
and ( w_4231 , \2541_b1 , \2541_b0 );
or ( \2543_b1 , \2346_b1 , \2347_b1 );
not ( \2347_b1 , w_4232 );
and ( \2543_b0 , \2346_b0 , w_4233 );
and ( w_4232 , w_4233 , \2347_b0 );
or ( \2544_b1 , \2348_b1 , \2351_b1 );
not ( \2351_b1 , w_4234 );
and ( \2544_b0 , \2348_b0 , w_4235 );
and ( w_4234 , w_4235 , \2351_b0 );
or ( \2545_b1 , \2543_b1 , w_4236 );
or ( \2545_b0 , \2543_b0 , \2544_b0 );
not ( \2544_b0 , w_4237 );
and ( w_4237 , w_4236 , \2544_b1 );
or ( \2546_b1 , \2542_b1 , \2545_b1 );
xor ( \2546_b0 , \2542_b0 , w_4238 );
not ( w_4238 , w_4239 );
and ( w_4239 , \2545_b1 , \2545_b0 );
or ( \2547_b1 , \1403_A[7]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_4240 );
and ( \2547_b0 , \1403_A[7]_b0 , w_4241 );
and ( w_4240 , w_4241 , \1439_B[7]_b0 );
or ( \2548_b1 , \2546_b1 , \2547_b1 );
xor ( \2548_b0 , \2546_b0 , w_4242 );
not ( w_4242 , w_4243 );
and ( w_4243 , \2547_b1 , \2547_b0 );
or ( \2549_b1 , \2352_b1 , \2353_b1 );
not ( \2353_b1 , w_4244 );
and ( \2549_b0 , \2352_b0 , w_4245 );
and ( w_4244 , w_4245 , \2353_b0 );
or ( \2550_b1 , \2354_b1 , \2357_b1 );
not ( \2357_b1 , w_4246 );
and ( \2550_b0 , \2354_b0 , w_4247 );
and ( w_4246 , w_4247 , \2357_b0 );
or ( \2551_b1 , \2549_b1 , w_4248 );
or ( \2551_b0 , \2549_b0 , \2550_b0 );
not ( \2550_b0 , w_4249 );
and ( w_4249 , w_4248 , \2550_b1 );
or ( \2552_b1 , \2548_b1 , \2551_b1 );
xor ( \2552_b0 , \2548_b0 , w_4250 );
not ( w_4250 , w_4251 );
and ( w_4251 , \2551_b1 , \2551_b0 );
or ( \2553_b1 , \1293_A[6]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_4252 );
and ( \2553_b0 , \1293_A[6]_b0 , w_4253 );
and ( w_4252 , w_4253 , \1567_B[8]_b0 );
or ( \2554_b1 , \2552_b1 , \2553_b1 );
xor ( \2554_b0 , \2552_b0 , w_4254 );
not ( w_4254 , w_4255 );
and ( w_4255 , \2553_b1 , \2553_b0 );
or ( \2555_b1 , \2358_b1 , \2359_b1 );
not ( \2359_b1 , w_4256 );
and ( \2555_b0 , \2358_b0 , w_4257 );
and ( w_4256 , w_4257 , \2359_b0 );
or ( \2556_b1 , \2360_b1 , \2363_b1 );
not ( \2363_b1 , w_4258 );
and ( \2556_b0 , \2360_b0 , w_4259 );
and ( w_4258 , w_4259 , \2363_b0 );
or ( \2557_b1 , \2555_b1 , w_4260 );
or ( \2557_b0 , \2555_b0 , \2556_b0 );
not ( \2556_b0 , w_4261 );
and ( w_4261 , w_4260 , \2556_b1 );
or ( \2558_b1 , \2554_b1 , \2557_b1 );
xor ( \2558_b0 , \2554_b0 , w_4262 );
not ( w_4262 , w_4263 );
and ( w_4263 , \2557_b1 , \2557_b0 );
or ( \2559_b1 , \1195_A[5]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_4264 );
and ( \2559_b0 , \1195_A[5]_b0 , w_4265 );
and ( w_4264 , w_4265 , \1707_B[9]_b0 );
or ( \2560_b1 , \2558_b1 , \2559_b1 );
xor ( \2560_b0 , \2558_b0 , w_4266 );
not ( w_4266 , w_4267 );
and ( w_4267 , \2559_b1 , \2559_b0 );
or ( \2561_b1 , \2364_b1 , \2365_b1 );
not ( \2365_b1 , w_4268 );
and ( \2561_b0 , \2364_b0 , w_4269 );
and ( w_4268 , w_4269 , \2365_b0 );
or ( \2562_b1 , \2366_b1 , \2369_b1 );
not ( \2369_b1 , w_4270 );
and ( \2562_b0 , \2366_b0 , w_4271 );
and ( w_4270 , w_4271 , \2369_b0 );
or ( \2563_b1 , \2561_b1 , w_4272 );
or ( \2563_b0 , \2561_b0 , \2562_b0 );
not ( \2562_b0 , w_4273 );
and ( w_4273 , w_4272 , \2562_b1 );
or ( \2564_b1 , \2560_b1 , \2563_b1 );
xor ( \2564_b0 , \2560_b0 , w_4274 );
not ( w_4274 , w_4275 );
and ( w_4275 , \2563_b1 , \2563_b0 );
or ( \2565_b1 , \1109_A[4]_b1 , \1859_B[10]_b1 );
not ( \1859_B[10]_b1 , w_4276 );
and ( \2565_b0 , \1109_A[4]_b0 , w_4277 );
and ( w_4276 , w_4277 , \1859_B[10]_b0 );
or ( \2566_b1 , \2564_b1 , \2565_b1 );
xor ( \2566_b0 , \2564_b0 , w_4278 );
not ( w_4278 , w_4279 );
and ( w_4279 , \2565_b1 , \2565_b0 );
or ( \2567_b1 , \2370_b1 , \2371_b1 );
not ( \2371_b1 , w_4280 );
and ( \2567_b0 , \2370_b0 , w_4281 );
and ( w_4280 , w_4281 , \2371_b0 );
or ( \2568_b1 , \2372_b1 , \2375_b1 );
not ( \2375_b1 , w_4282 );
and ( \2568_b0 , \2372_b0 , w_4283 );
and ( w_4282 , w_4283 , \2375_b0 );
or ( \2569_b1 , \2567_b1 , w_4284 );
or ( \2569_b0 , \2567_b0 , \2568_b0 );
not ( \2568_b0 , w_4285 );
and ( w_4285 , w_4284 , \2568_b1 );
or ( \2570_b1 , \2566_b1 , \2569_b1 );
xor ( \2570_b0 , \2566_b0 , w_4286 );
not ( w_4286 , w_4287 );
and ( w_4287 , \2569_b1 , \2569_b0 );
or ( \2571_b1 , \1035_A[3]_b1 , \2023_B[11]_b1 );
not ( \2023_B[11]_b1 , w_4288 );
and ( \2571_b0 , \1035_A[3]_b0 , w_4289 );
and ( w_4288 , w_4289 , \2023_B[11]_b0 );
or ( \2572_b1 , \2570_b1 , \2571_b1 );
xor ( \2572_b0 , \2570_b0 , w_4290 );
not ( w_4290 , w_4291 );
and ( w_4291 , \2571_b1 , \2571_b0 );
or ( \2573_b1 , \2376_b1 , \2377_b1 );
not ( \2377_b1 , w_4292 );
and ( \2573_b0 , \2376_b0 , w_4293 );
and ( w_4292 , w_4293 , \2377_b0 );
or ( \2574_b1 , \2378_b1 , \2381_b1 );
not ( \2381_b1 , w_4294 );
and ( \2574_b0 , \2378_b0 , w_4295 );
and ( w_4294 , w_4295 , \2381_b0 );
or ( \2575_b1 , \2573_b1 , w_4296 );
or ( \2575_b0 , \2573_b0 , \2574_b0 );
not ( \2574_b0 , w_4297 );
and ( w_4297 , w_4296 , \2574_b1 );
or ( \2576_b1 , \2572_b1 , \2575_b1 );
xor ( \2576_b0 , \2572_b0 , w_4298 );
not ( w_4298 , w_4299 );
and ( w_4299 , \2575_b1 , \2575_b0 );
or ( \2577_b1 , \973_A[2]_b1 , \2199_B[12]_b1 );
not ( \2199_B[12]_b1 , w_4300 );
and ( \2577_b0 , \973_A[2]_b0 , w_4301 );
and ( w_4300 , w_4301 , \2199_B[12]_b0 );
or ( \2578_b1 , \2576_b1 , \2577_b1 );
xor ( \2578_b0 , \2576_b0 , w_4302 );
not ( w_4302 , w_4303 );
and ( w_4303 , \2577_b1 , \2577_b0 );
or ( \2579_b1 , \2382_b1 , \2383_b1 );
not ( \2383_b1 , w_4304 );
and ( \2579_b0 , \2382_b0 , w_4305 );
and ( w_4304 , w_4305 , \2383_b0 );
or ( \2580_b1 , \2384_b1 , \2385_b1 );
not ( \2385_b1 , w_4306 );
and ( \2580_b0 , \2384_b0 , w_4307 );
and ( w_4306 , w_4307 , \2385_b0 );
or ( \2581_b1 , \2579_b1 , w_4308 );
or ( \2581_b0 , \2579_b0 , \2580_b0 );
not ( \2580_b0 , w_4309 );
and ( w_4309 , w_4308 , \2580_b1 );
or ( \2582_b1 , \2578_b1 , \2581_b1 );
xor ( \2582_b0 , \2578_b0 , w_4310 );
not ( w_4310 , w_4311 );
and ( w_4311 , \2581_b1 , \2581_b0 );
or ( \2583_b1 , \927_A[1]_b1 , \2387_B[13]_b1 );
not ( \2387_B[13]_b1 , w_4312 );
and ( \2583_b0 , \927_A[1]_b0 , w_4313 );
and ( w_4312 , w_4313 , \2387_B[13]_b0 );
or ( \2584_b1 , \2582_b1 , \2583_b1 );
xor ( \2584_b0 , \2582_b0 , w_4314 );
not ( w_4314 , w_4315 );
and ( w_4315 , \2583_b1 , \2583_b0 );
or ( \2585_b1 , \2386_b1 , \2388_b1 );
not ( \2388_b1 , w_4316 );
and ( \2585_b0 , \2386_b0 , w_4317 );
and ( w_4316 , w_4317 , \2388_b0 );
or ( \2586_b1 , \2584_b1 , \2585_b1 );
xor ( \2586_b0 , \2584_b0 , w_4318 );
not ( w_4318 , w_4319 );
and ( w_4319 , \2585_b1 , \2585_b0 );
buf ( \2587_B[14]_b1 , \d[14]_b1 );
buf ( \2587_B[14]_b0 , \d[14]_b0 );
or ( \2588_b1 , \891_A[0]_b1 , \2587_B[14]_b1 );
not ( \2587_B[14]_b1 , w_4320 );
and ( \2588_b0 , \891_A[0]_b0 , w_4321 );
and ( w_4320 , w_4321 , \2587_B[14]_b0 );
or ( \2589_b1 , \2586_b1 , \2588_b1 );
xor ( \2589_b0 , \2586_b0 , w_4322 );
not ( w_4322 , w_4323 );
and ( w_4323 , \2588_b1 , \2588_b0 );
buf ( \2590_Z[14]_b1 , \2589_b1 );
buf ( \2590_Z[14]_b0 , \2589_b0 );
or ( \2591_b1 , \2590_Z[14]_b1 , \865_b1 );
not ( \865_b1 , w_4324 );
and ( \2591_b0 , \2590_Z[14]_b0 , w_4325 );
and ( w_4324 , w_4325 , \865_b0 );
buf ( \2592_A[14]_b1 , \b[14]_b1 );
buf ( \2592_A[14]_b0 , \b[14]_b0 );
buf ( \2593_B[14]_b1 , \d[14]_b1 );
buf ( \2593_B[14]_b0 , \d[14]_b0 );
or ( \2594_b1 , \2592_A[14]_b1 , \2593_B[14]_b1 );
xor ( \2594_b0 , \2592_A[14]_b0 , w_4326 );
not ( w_4326 , w_4327 );
and ( w_4327 , \2593_B[14]_b1 , \2593_B[14]_b0 );
or ( \2595_b1 , \2392_A[13]_b1 , \2393_B[13]_b1 );
not ( \2393_B[13]_b1 , w_4328 );
and ( \2595_b0 , \2392_A[13]_b0 , w_4329 );
and ( w_4328 , w_4329 , \2393_B[13]_b0 );
or ( \2596_b1 , \2393_B[13]_b1 , \2398_b1 );
not ( \2398_b1 , w_4330 );
and ( \2596_b0 , \2393_B[13]_b0 , w_4331 );
and ( w_4330 , w_4331 , \2398_b0 );
or ( \2597_b1 , \2392_A[13]_b1 , \2398_b1 );
not ( \2398_b1 , w_4332 );
and ( \2597_b0 , \2392_A[13]_b0 , w_4333 );
and ( w_4332 , w_4333 , \2398_b0 );
or ( \2599_b1 , \2594_b1 , \2598_b1 );
xor ( \2599_b0 , \2594_b0 , w_4334 );
not ( w_4334 , w_4335 );
and ( w_4335 , \2598_b1 , \2598_b0 );
buf ( \2600_SUM[14]_b1 , \2599_b1 );
buf ( \2600_SUM[14]_b0 , \2599_b0 );
or ( \2601_b1 , \2600_SUM[14]_b1 , \863_b1 );
not ( \863_b1 , w_4336 );
and ( \2601_b0 , \2600_SUM[14]_b0 , w_4337 );
and ( w_4336 , w_4337 , \863_b0 );
buf ( \2602_A[14]_b1 , \a[14]_b1 );
buf ( \2602_A[14]_b0 , \a[14]_b0 );
buf ( \2603_B[14]_b1 , \c[14]_b1 );
buf ( \2603_B[14]_b0 , \c[14]_b0 );
or ( \2604_b1 , \2602_A[14]_b1 , \2603_B[14]_b1 );
xor ( \2604_b0 , \2602_A[14]_b0 , w_4338 );
not ( w_4338 , w_4339 );
and ( w_4339 , \2603_B[14]_b1 , \2603_B[14]_b0 );
or ( \2605_b1 , \2402_A[13]_b1 , \2403_B[13]_b1 );
not ( \2403_B[13]_b1 , w_4340 );
and ( \2605_b0 , \2402_A[13]_b0 , w_4341 );
and ( w_4340 , w_4341 , \2403_B[13]_b0 );
or ( \2606_b1 , \2403_B[13]_b1 , \2408_b1 );
not ( \2408_b1 , w_4342 );
and ( \2606_b0 , \2403_B[13]_b0 , w_4343 );
and ( w_4342 , w_4343 , \2408_b0 );
or ( \2607_b1 , \2402_A[13]_b1 , \2408_b1 );
not ( \2408_b1 , w_4344 );
and ( \2607_b0 , \2402_A[13]_b0 , w_4345 );
and ( w_4344 , w_4345 , \2408_b0 );
or ( \2609_b1 , \2604_b1 , \2608_b1 );
xor ( \2609_b0 , \2604_b0 , w_4346 );
not ( w_4346 , w_4347 );
and ( w_4347 , \2608_b1 , \2608_b0 );
buf ( \2610_SUM[14]_b1 , \2609_b1 );
buf ( \2610_SUM[14]_b0 , \2609_b0 );
or ( \2611_b1 , \2610_SUM[14]_b1 , \861_b1 );
not ( \861_b1 , w_4348 );
and ( \2611_b0 , \2610_SUM[14]_b0 , w_4349 );
and ( w_4348 , w_4349 , \861_b0 );
or ( \2612_b1 , \d[14]_b1 , \859_b1 );
not ( \859_b1 , w_4350 );
and ( \2612_b0 , \d[14]_b0 , w_4351 );
and ( w_4350 , w_4351 , \859_b0 );
or ( \2613_b1 , \c[14]_b1 , \857_b1 );
not ( \857_b1 , w_4352 );
and ( \2613_b0 , \c[14]_b0 , w_4353 );
and ( w_4352 , w_4353 , \857_b0 );
or ( \2614_b1 , \b[14]_b1 , \855_b1 );
not ( \855_b1 , w_4354 );
and ( \2614_b0 , \b[14]_b0 , w_4355 );
and ( w_4354 , w_4355 , \855_b0 );
or ( \2615_b1 , \a[14]_b1 , \853_b1 );
not ( \853_b1 , w_4356 );
and ( \2615_b0 , \a[14]_b0 , w_4357 );
and ( w_4356 , w_4357 , \853_b0 );
and ( \2617_b1 , 1'b0_b1 , w_4358 );
xor ( w_4358 , 1'b0_b0 , \876_b1 );
not ( \876_b1 , w_4359 );
and ( \2617_b0 , w_4359 , \876_b0 );
or ( \2618_b1 , \a[15]_b1 , w_4360 );
or ( \2618_b0 , \a[15]_b0 , \d[15]_b0 );
not ( \d[15]_b0 , w_4361 );
and ( w_4361 , w_4360 , \d[15]_b1 );
or ( \2619_b1 , \2618_b1 , \875_b1 );
not ( \875_b1 , w_4362 );
and ( \2619_b0 , \2618_b0 , w_4363 );
and ( w_4362 , w_4363 , \875_b0 );
or ( \2620_b1 , \b[15]_b1 , \c[15]_b1 );
not ( \c[15]_b1 , w_4364 );
and ( \2620_b0 , \b[15]_b0 , w_4365 );
and ( w_4364 , w_4365 , \c[15]_b0 );
or ( \2621_b1 , \2620_b1 , \873_b1 );
not ( \873_b1 , w_4366 );
and ( \2621_b0 , \2620_b0 , w_4367 );
and ( w_4366 , w_4367 , \873_b0 );
or ( \2622_b1 , \a[15]_b1 , w_4368 );
or ( \2622_b0 , \a[15]_b0 , \b[15]_b0 );
not ( \b[15]_b0 , w_4369 );
and ( w_4369 , w_4368 , \b[15]_b1 );
or ( \2623_b1 , \2622_b1 , \871_b1 );
not ( \871_b1 , w_4370 );
and ( \2623_b0 , \2622_b0 , w_4371 );
and ( w_4370 , w_4371 , \871_b0 );
or ( \2624_b1 , \c[15]_b1 , \d[15]_b1 );
xor ( \2624_b0 , \c[15]_b0 , w_4372 );
not ( w_4372 , w_4373 );
and ( w_4373 , \d[15]_b1 , \d[15]_b0 );
or ( \2625_b1 , \2624_b1 , \869_b1 );
not ( \869_b1 , w_4374 );
and ( \2625_b0 , \2624_b0 , w_4375 );
and ( w_4374 , w_4375 , \869_b0 );
buf ( \2626_A[15]_b1 , \b[15]_b1 );
buf ( \2626_A[15]_b0 , \b[15]_b0 );
or ( \2627_b1 , \2626_A[15]_b1 , \887_B[0]_b1 );
not ( \887_B[0]_b1 , w_4376 );
and ( \2627_b0 , \2626_A[15]_b0 , w_4377 );
and ( w_4376 , w_4377 , \887_B[0]_b0 );
or ( \2628_b1 , \2426_A[14]_b1 , \922_B[1]_b1 );
not ( \922_B[1]_b1 , w_4378 );
and ( \2628_b0 , \2426_A[14]_b0 , w_4379 );
and ( w_4378 , w_4379 , \922_B[1]_b0 );
or ( \2629_b1 , \2627_b1 , \2628_b1 );
xor ( \2629_b0 , \2627_b0 , w_4380 );
not ( w_4380 , w_4381 );
and ( w_4381 , \2628_b1 , \2628_b0 );
or ( \2630_b1 , \2427_b1 , \2428_b1 );
not ( \2428_b1 , w_4382 );
and ( \2630_b0 , \2427_b0 , w_4383 );
and ( w_4382 , w_4383 , \2428_b0 );
or ( \2631_b1 , \2429_b1 , \2432_b1 );
not ( \2432_b1 , w_4384 );
and ( \2631_b0 , \2429_b0 , w_4385 );
and ( w_4384 , w_4385 , \2432_b0 );
or ( \2632_b1 , \2630_b1 , w_4386 );
or ( \2632_b0 , \2630_b0 , \2631_b0 );
not ( \2631_b0 , w_4387 );
and ( w_4387 , w_4386 , \2631_b1 );
or ( \2633_b1 , \2629_b1 , \2632_b1 );
xor ( \2633_b0 , \2629_b0 , w_4388 );
not ( w_4388 , w_4389 );
and ( w_4389 , \2632_b1 , \2632_b0 );
or ( \2634_b1 , \2238_A[13]_b1 , \968_B[2]_b1 );
not ( \968_B[2]_b1 , w_4390 );
and ( \2634_b0 , \2238_A[13]_b0 , w_4391 );
and ( w_4390 , w_4391 , \968_B[2]_b0 );
or ( \2635_b1 , \2633_b1 , \2634_b1 );
xor ( \2635_b0 , \2633_b0 , w_4392 );
not ( w_4392 , w_4393 );
and ( w_4393 , \2634_b1 , \2634_b0 );
or ( \2636_b1 , \2433_b1 , \2434_b1 );
not ( \2434_b1 , w_4394 );
and ( \2636_b0 , \2433_b0 , w_4395 );
and ( w_4394 , w_4395 , \2434_b0 );
or ( \2637_b1 , \2435_b1 , \2438_b1 );
not ( \2438_b1 , w_4396 );
and ( \2637_b0 , \2435_b0 , w_4397 );
and ( w_4396 , w_4397 , \2438_b0 );
or ( \2638_b1 , \2636_b1 , w_4398 );
or ( \2638_b0 , \2636_b0 , \2637_b0 );
not ( \2637_b0 , w_4399 );
and ( w_4399 , w_4398 , \2637_b1 );
or ( \2639_b1 , \2635_b1 , \2638_b1 );
xor ( \2639_b0 , \2635_b0 , w_4400 );
not ( w_4400 , w_4401 );
and ( w_4401 , \2638_b1 , \2638_b0 );
or ( \2640_b1 , \2062_A[12]_b1 , \1030_B[3]_b1 );
not ( \1030_B[3]_b1 , w_4402 );
and ( \2640_b0 , \2062_A[12]_b0 , w_4403 );
and ( w_4402 , w_4403 , \1030_B[3]_b0 );
or ( \2641_b1 , \2639_b1 , \2640_b1 );
xor ( \2641_b0 , \2639_b0 , w_4404 );
not ( w_4404 , w_4405 );
and ( w_4405 , \2640_b1 , \2640_b0 );
or ( \2642_b1 , \2439_b1 , \2440_b1 );
not ( \2440_b1 , w_4406 );
and ( \2642_b0 , \2439_b0 , w_4407 );
and ( w_4406 , w_4407 , \2440_b0 );
or ( \2643_b1 , \2441_b1 , \2444_b1 );
not ( \2444_b1 , w_4408 );
and ( \2643_b0 , \2441_b0 , w_4409 );
and ( w_4408 , w_4409 , \2444_b0 );
or ( \2644_b1 , \2642_b1 , w_4410 );
or ( \2644_b0 , \2642_b0 , \2643_b0 );
not ( \2643_b0 , w_4411 );
and ( w_4411 , w_4410 , \2643_b1 );
or ( \2645_b1 , \2641_b1 , \2644_b1 );
xor ( \2645_b0 , \2641_b0 , w_4412 );
not ( w_4412 , w_4413 );
and ( w_4413 , \2644_b1 , \2644_b0 );
or ( \2646_b1 , \1898_A[11]_b1 , \1104_B[4]_b1 );
not ( \1104_B[4]_b1 , w_4414 );
and ( \2646_b0 , \1898_A[11]_b0 , w_4415 );
and ( w_4414 , w_4415 , \1104_B[4]_b0 );
or ( \2647_b1 , \2645_b1 , \2646_b1 );
xor ( \2647_b0 , \2645_b0 , w_4416 );
not ( w_4416 , w_4417 );
and ( w_4417 , \2646_b1 , \2646_b0 );
or ( \2648_b1 , \2445_b1 , \2446_b1 );
not ( \2446_b1 , w_4418 );
and ( \2648_b0 , \2445_b0 , w_4419 );
and ( w_4418 , w_4419 , \2446_b0 );
or ( \2649_b1 , \2447_b1 , \2450_b1 );
not ( \2450_b1 , w_4420 );
and ( \2649_b0 , \2447_b0 , w_4421 );
and ( w_4420 , w_4421 , \2450_b0 );
or ( \2650_b1 , \2648_b1 , w_4422 );
or ( \2650_b0 , \2648_b0 , \2649_b0 );
not ( \2649_b0 , w_4423 );
and ( w_4423 , w_4422 , \2649_b1 );
or ( \2651_b1 , \2647_b1 , \2650_b1 );
xor ( \2651_b0 , \2647_b0 , w_4424 );
not ( w_4424 , w_4425 );
and ( w_4425 , \2650_b1 , \2650_b0 );
or ( \2652_b1 , \1746_A[10]_b1 , \1190_B[5]_b1 );
not ( \1190_B[5]_b1 , w_4426 );
and ( \2652_b0 , \1746_A[10]_b0 , w_4427 );
and ( w_4426 , w_4427 , \1190_B[5]_b0 );
or ( \2653_b1 , \2651_b1 , \2652_b1 );
xor ( \2653_b0 , \2651_b0 , w_4428 );
not ( w_4428 , w_4429 );
and ( w_4429 , \2652_b1 , \2652_b0 );
or ( \2654_b1 , \2451_b1 , \2452_b1 );
not ( \2452_b1 , w_4430 );
and ( \2654_b0 , \2451_b0 , w_4431 );
and ( w_4430 , w_4431 , \2452_b0 );
or ( \2655_b1 , \2453_b1 , \2456_b1 );
not ( \2456_b1 , w_4432 );
and ( \2655_b0 , \2453_b0 , w_4433 );
and ( w_4432 , w_4433 , \2456_b0 );
or ( \2656_b1 , \2654_b1 , w_4434 );
or ( \2656_b0 , \2654_b0 , \2655_b0 );
not ( \2655_b0 , w_4435 );
and ( w_4435 , w_4434 , \2655_b1 );
or ( \2657_b1 , \2653_b1 , \2656_b1 );
xor ( \2657_b0 , \2653_b0 , w_4436 );
not ( w_4436 , w_4437 );
and ( w_4437 , \2656_b1 , \2656_b0 );
or ( \2658_b1 , \1606_A[9]_b1 , \1288_B[6]_b1 );
not ( \1288_B[6]_b1 , w_4438 );
and ( \2658_b0 , \1606_A[9]_b0 , w_4439 );
and ( w_4438 , w_4439 , \1288_B[6]_b0 );
or ( \2659_b1 , \2657_b1 , \2658_b1 );
xor ( \2659_b0 , \2657_b0 , w_4440 );
not ( w_4440 , w_4441 );
and ( w_4441 , \2658_b1 , \2658_b0 );
or ( \2660_b1 , \2457_b1 , \2458_b1 );
not ( \2458_b1 , w_4442 );
and ( \2660_b0 , \2457_b0 , w_4443 );
and ( w_4442 , w_4443 , \2458_b0 );
or ( \2661_b1 , \2459_b1 , \2462_b1 );
not ( \2462_b1 , w_4444 );
and ( \2661_b0 , \2459_b0 , w_4445 );
and ( w_4444 , w_4445 , \2462_b0 );
or ( \2662_b1 , \2660_b1 , w_4446 );
or ( \2662_b0 , \2660_b0 , \2661_b0 );
not ( \2661_b0 , w_4447 );
and ( w_4447 , w_4446 , \2661_b1 );
or ( \2663_b1 , \2659_b1 , \2662_b1 );
xor ( \2663_b0 , \2659_b0 , w_4448 );
not ( w_4448 , w_4449 );
and ( w_4449 , \2662_b1 , \2662_b0 );
or ( \2664_b1 , \1478_A[8]_b1 , \1398_B[7]_b1 );
not ( \1398_B[7]_b1 , w_4450 );
and ( \2664_b0 , \1478_A[8]_b0 , w_4451 );
and ( w_4450 , w_4451 , \1398_B[7]_b0 );
or ( \2665_b1 , \2663_b1 , \2664_b1 );
xor ( \2665_b0 , \2663_b0 , w_4452 );
not ( w_4452 , w_4453 );
and ( w_4453 , \2664_b1 , \2664_b0 );
or ( \2666_b1 , \2463_b1 , \2464_b1 );
not ( \2464_b1 , w_4454 );
and ( \2666_b0 , \2463_b0 , w_4455 );
and ( w_4454 , w_4455 , \2464_b0 );
or ( \2667_b1 , \2465_b1 , \2468_b1 );
not ( \2468_b1 , w_4456 );
and ( \2667_b0 , \2465_b0 , w_4457 );
and ( w_4456 , w_4457 , \2468_b0 );
or ( \2668_b1 , \2666_b1 , w_4458 );
or ( \2668_b0 , \2666_b0 , \2667_b0 );
not ( \2667_b0 , w_4459 );
and ( w_4459 , w_4458 , \2667_b1 );
or ( \2669_b1 , \2665_b1 , \2668_b1 );
xor ( \2669_b0 , \2665_b0 , w_4460 );
not ( w_4460 , w_4461 );
and ( w_4461 , \2668_b1 , \2668_b0 );
or ( \2670_b1 , \1362_A[7]_b1 , \1520_B[8]_b1 );
not ( \1520_B[8]_b1 , w_4462 );
and ( \2670_b0 , \1362_A[7]_b0 , w_4463 );
and ( w_4462 , w_4463 , \1520_B[8]_b0 );
or ( \2671_b1 , \2669_b1 , \2670_b1 );
xor ( \2671_b0 , \2669_b0 , w_4464 );
not ( w_4464 , w_4465 );
and ( w_4465 , \2670_b1 , \2670_b0 );
or ( \2672_b1 , \2469_b1 , \2470_b1 );
not ( \2470_b1 , w_4466 );
and ( \2672_b0 , \2469_b0 , w_4467 );
and ( w_4466 , w_4467 , \2470_b0 );
or ( \2673_b1 , \2471_b1 , \2474_b1 );
not ( \2474_b1 , w_4468 );
and ( \2673_b0 , \2471_b0 , w_4469 );
and ( w_4468 , w_4469 , \2474_b0 );
or ( \2674_b1 , \2672_b1 , w_4470 );
or ( \2674_b0 , \2672_b0 , \2673_b0 );
not ( \2673_b0 , w_4471 );
and ( w_4471 , w_4470 , \2673_b1 );
or ( \2675_b1 , \2671_b1 , \2674_b1 );
xor ( \2675_b0 , \2671_b0 , w_4472 );
not ( w_4472 , w_4473 );
and ( w_4473 , \2674_b1 , \2674_b0 );
or ( \2676_b1 , \1258_A[6]_b1 , \1654_B[9]_b1 );
not ( \1654_B[9]_b1 , w_4474 );
and ( \2676_b0 , \1258_A[6]_b0 , w_4475 );
and ( w_4474 , w_4475 , \1654_B[9]_b0 );
or ( \2677_b1 , \2675_b1 , \2676_b1 );
xor ( \2677_b0 , \2675_b0 , w_4476 );
not ( w_4476 , w_4477 );
and ( w_4477 , \2676_b1 , \2676_b0 );
or ( \2678_b1 , \2475_b1 , \2476_b1 );
not ( \2476_b1 , w_4478 );
and ( \2678_b0 , \2475_b0 , w_4479 );
and ( w_4478 , w_4479 , \2476_b0 );
or ( \2679_b1 , \2477_b1 , \2480_b1 );
not ( \2480_b1 , w_4480 );
and ( \2679_b0 , \2477_b0 , w_4481 );
and ( w_4480 , w_4481 , \2480_b0 );
or ( \2680_b1 , \2678_b1 , w_4482 );
or ( \2680_b0 , \2678_b0 , \2679_b0 );
not ( \2679_b0 , w_4483 );
and ( w_4483 , w_4482 , \2679_b1 );
or ( \2681_b1 , \2677_b1 , \2680_b1 );
xor ( \2681_b0 , \2677_b0 , w_4484 );
not ( w_4484 , w_4485 );
and ( w_4485 , \2680_b1 , \2680_b0 );
or ( \2682_b1 , \1166_A[5]_b1 , \1800_B[10]_b1 );
not ( \1800_B[10]_b1 , w_4486 );
and ( \2682_b0 , \1166_A[5]_b0 , w_4487 );
and ( w_4486 , w_4487 , \1800_B[10]_b0 );
or ( \2683_b1 , \2681_b1 , \2682_b1 );
xor ( \2683_b0 , \2681_b0 , w_4488 );
not ( w_4488 , w_4489 );
and ( w_4489 , \2682_b1 , \2682_b0 );
or ( \2684_b1 , \2481_b1 , \2482_b1 );
not ( \2482_b1 , w_4490 );
and ( \2684_b0 , \2481_b0 , w_4491 );
and ( w_4490 , w_4491 , \2482_b0 );
or ( \2685_b1 , \2483_b1 , \2486_b1 );
not ( \2486_b1 , w_4492 );
and ( \2685_b0 , \2483_b0 , w_4493 );
and ( w_4492 , w_4493 , \2486_b0 );
or ( \2686_b1 , \2684_b1 , w_4494 );
or ( \2686_b0 , \2684_b0 , \2685_b0 );
not ( \2685_b0 , w_4495 );
and ( w_4495 , w_4494 , \2685_b1 );
or ( \2687_b1 , \2683_b1 , \2686_b1 );
xor ( \2687_b0 , \2683_b0 , w_4496 );
not ( w_4496 , w_4497 );
and ( w_4497 , \2686_b1 , \2686_b0 );
or ( \2688_b1 , \1086_A[4]_b1 , \1958_B[11]_b1 );
not ( \1958_B[11]_b1 , w_4498 );
and ( \2688_b0 , \1086_A[4]_b0 , w_4499 );
and ( w_4498 , w_4499 , \1958_B[11]_b0 );
or ( \2689_b1 , \2687_b1 , \2688_b1 );
xor ( \2689_b0 , \2687_b0 , w_4500 );
not ( w_4500 , w_4501 );
and ( w_4501 , \2688_b1 , \2688_b0 );
or ( \2690_b1 , \2487_b1 , \2488_b1 );
not ( \2488_b1 , w_4502 );
and ( \2690_b0 , \2487_b0 , w_4503 );
and ( w_4502 , w_4503 , \2488_b0 );
or ( \2691_b1 , \2489_b1 , \2492_b1 );
not ( \2492_b1 , w_4504 );
and ( \2691_b0 , \2489_b0 , w_4505 );
and ( w_4504 , w_4505 , \2492_b0 );
or ( \2692_b1 , \2690_b1 , w_4506 );
or ( \2692_b0 , \2690_b0 , \2691_b0 );
not ( \2691_b0 , w_4507 );
and ( w_4507 , w_4506 , \2691_b1 );
or ( \2693_b1 , \2689_b1 , \2692_b1 );
xor ( \2693_b0 , \2689_b0 , w_4508 );
not ( w_4508 , w_4509 );
and ( w_4509 , \2692_b1 , \2692_b0 );
or ( \2694_b1 , \1018_A[3]_b1 , \2128_B[12]_b1 );
not ( \2128_B[12]_b1 , w_4510 );
and ( \2694_b0 , \1018_A[3]_b0 , w_4511 );
and ( w_4510 , w_4511 , \2128_B[12]_b0 );
or ( \2695_b1 , \2693_b1 , \2694_b1 );
xor ( \2695_b0 , \2693_b0 , w_4512 );
not ( w_4512 , w_4513 );
and ( w_4513 , \2694_b1 , \2694_b0 );
or ( \2696_b1 , \2493_b1 , \2494_b1 );
not ( \2494_b1 , w_4514 );
and ( \2696_b0 , \2493_b0 , w_4515 );
and ( w_4514 , w_4515 , \2494_b0 );
or ( \2697_b1 , \2495_b1 , \2498_b1 );
not ( \2498_b1 , w_4516 );
and ( \2697_b0 , \2495_b0 , w_4517 );
and ( w_4516 , w_4517 , \2498_b0 );
or ( \2698_b1 , \2696_b1 , w_4518 );
or ( \2698_b0 , \2696_b0 , \2697_b0 );
not ( \2697_b0 , w_4519 );
and ( w_4519 , w_4518 , \2697_b1 );
or ( \2699_b1 , \2695_b1 , \2698_b1 );
xor ( \2699_b0 , \2695_b0 , w_4520 );
not ( w_4520 , w_4521 );
and ( w_4521 , \2698_b1 , \2698_b0 );
or ( \2700_b1 , \962_A[2]_b1 , \2310_B[13]_b1 );
not ( \2310_B[13]_b1 , w_4522 );
and ( \2700_b0 , \962_A[2]_b0 , w_4523 );
and ( w_4522 , w_4523 , \2310_B[13]_b0 );
or ( \2701_b1 , \2699_b1 , \2700_b1 );
xor ( \2701_b0 , \2699_b0 , w_4524 );
not ( w_4524 , w_4525 );
and ( w_4525 , \2700_b1 , \2700_b0 );
or ( \2702_b1 , \2499_b1 , \2500_b1 );
not ( \2500_b1 , w_4526 );
and ( \2702_b0 , \2499_b0 , w_4527 );
and ( w_4526 , w_4527 , \2500_b0 );
or ( \2703_b1 , \2501_b1 , \2502_b1 );
not ( \2502_b1 , w_4528 );
and ( \2703_b0 , \2501_b0 , w_4529 );
and ( w_4528 , w_4529 , \2502_b0 );
or ( \2704_b1 , \2702_b1 , w_4530 );
or ( \2704_b0 , \2702_b0 , \2703_b0 );
not ( \2703_b0 , w_4531 );
and ( w_4531 , w_4530 , \2703_b1 );
or ( \2705_b1 , \2701_b1 , \2704_b1 );
xor ( \2705_b0 , \2701_b0 , w_4532 );
not ( w_4532 , w_4533 );
and ( w_4533 , \2704_b1 , \2704_b0 );
or ( \2706_b1 , \920_A[1]_b1 , \2504_B[14]_b1 );
not ( \2504_B[14]_b1 , w_4534 );
and ( \2706_b0 , \920_A[1]_b0 , w_4535 );
and ( w_4534 , w_4535 , \2504_B[14]_b0 );
or ( \2707_b1 , \2705_b1 , \2706_b1 );
xor ( \2707_b0 , \2705_b0 , w_4536 );
not ( w_4536 , w_4537 );
and ( w_4537 , \2706_b1 , \2706_b0 );
or ( \2708_b1 , \2503_b1 , \2505_b1 );
not ( \2505_b1 , w_4538 );
and ( \2708_b0 , \2503_b0 , w_4539 );
and ( w_4538 , w_4539 , \2505_b0 );
or ( \2709_b1 , \2707_b1 , \2708_b1 );
xor ( \2709_b0 , \2707_b0 , w_4540 );
not ( w_4540 , w_4541 );
and ( w_4541 , \2708_b1 , \2708_b0 );
buf ( \2710_B[15]_b1 , \c[15]_b1 );
buf ( \2710_B[15]_b0 , \c[15]_b0 );
or ( \2711_b1 , \886_A[0]_b1 , \2710_B[15]_b1 );
not ( \2710_B[15]_b1 , w_4542 );
and ( \2711_b0 , \886_A[0]_b0 , w_4543 );
and ( w_4542 , w_4543 , \2710_B[15]_b0 );
or ( \2712_b1 , \2709_b1 , \2711_b1 );
xor ( \2712_b0 , \2709_b0 , w_4544 );
not ( w_4544 , w_4545 );
and ( w_4545 , \2711_b1 , \2711_b0 );
buf ( \2713_Z[15]_b1 , \2712_b1 );
buf ( \2713_Z[15]_b0 , \2712_b0 );
or ( \2714_b1 , \2713_Z[15]_b1 , \867_b1 );
not ( \867_b1 , w_4546 );
and ( \2714_b0 , \2713_Z[15]_b0 , w_4547 );
and ( w_4546 , w_4547 , \867_b0 );
buf ( \2715_A[15]_b1 , \a[15]_b1 );
buf ( \2715_A[15]_b0 , \a[15]_b0 );
or ( \2716_b1 , \2715_A[15]_b1 , \892_B[0]_b1 );
not ( \892_B[0]_b1 , w_4548 );
and ( \2716_b0 , \2715_A[15]_b0 , w_4549 );
and ( w_4548 , w_4549 , \892_B[0]_b0 );
or ( \2717_b1 , \2509_A[14]_b1 , \929_B[1]_b1 );
not ( \929_B[1]_b1 , w_4550 );
and ( \2717_b0 , \2509_A[14]_b0 , w_4551 );
and ( w_4550 , w_4551 , \929_B[1]_b0 );
or ( \2718_b1 , \2716_b1 , \2717_b1 );
xor ( \2718_b0 , \2716_b0 , w_4552 );
not ( w_4552 , w_4553 );
and ( w_4553 , \2717_b1 , \2717_b0 );
or ( \2719_b1 , \2510_b1 , \2511_b1 );
not ( \2511_b1 , w_4554 );
and ( \2719_b0 , \2510_b0 , w_4555 );
and ( w_4554 , w_4555 , \2511_b0 );
or ( \2720_b1 , \2512_b1 , \2515_b1 );
not ( \2515_b1 , w_4556 );
and ( \2720_b0 , \2512_b0 , w_4557 );
and ( w_4556 , w_4557 , \2515_b0 );
or ( \2721_b1 , \2719_b1 , w_4558 );
or ( \2721_b0 , \2719_b0 , \2720_b0 );
not ( \2720_b0 , w_4559 );
and ( w_4559 , w_4558 , \2720_b1 );
or ( \2722_b1 , \2718_b1 , \2721_b1 );
xor ( \2722_b0 , \2718_b0 , w_4560 );
not ( w_4560 , w_4561 );
and ( w_4561 , \2721_b1 , \2721_b0 );
or ( \2723_b1 , \2315_A[13]_b1 , \979_B[2]_b1 );
not ( \979_B[2]_b1 , w_4562 );
and ( \2723_b0 , \2315_A[13]_b0 , w_4563 );
and ( w_4562 , w_4563 , \979_B[2]_b0 );
or ( \2724_b1 , \2722_b1 , \2723_b1 );
xor ( \2724_b0 , \2722_b0 , w_4564 );
not ( w_4564 , w_4565 );
and ( w_4565 , \2723_b1 , \2723_b0 );
or ( \2725_b1 , \2516_b1 , \2517_b1 );
not ( \2517_b1 , w_4566 );
and ( \2725_b0 , \2516_b0 , w_4567 );
and ( w_4566 , w_4567 , \2517_b0 );
or ( \2726_b1 , \2518_b1 , \2521_b1 );
not ( \2521_b1 , w_4568 );
and ( \2726_b0 , \2518_b0 , w_4569 );
and ( w_4568 , w_4569 , \2521_b0 );
or ( \2727_b1 , \2725_b1 , w_4570 );
or ( \2727_b0 , \2725_b0 , \2726_b0 );
not ( \2726_b0 , w_4571 );
and ( w_4571 , w_4570 , \2726_b1 );
or ( \2728_b1 , \2724_b1 , \2727_b1 );
xor ( \2728_b0 , \2724_b0 , w_4572 );
not ( w_4572 , w_4573 );
and ( w_4573 , \2727_b1 , \2727_b0 );
or ( \2729_b1 , \2133_A[12]_b1 , \1047_B[3]_b1 );
not ( \1047_B[3]_b1 , w_4574 );
and ( \2729_b0 , \2133_A[12]_b0 , w_4575 );
and ( w_4574 , w_4575 , \1047_B[3]_b0 );
or ( \2730_b1 , \2728_b1 , \2729_b1 );
xor ( \2730_b0 , \2728_b0 , w_4576 );
not ( w_4576 , w_4577 );
and ( w_4577 , \2729_b1 , \2729_b0 );
or ( \2731_b1 , \2522_b1 , \2523_b1 );
not ( \2523_b1 , w_4578 );
and ( \2731_b0 , \2522_b0 , w_4579 );
and ( w_4578 , w_4579 , \2523_b0 );
or ( \2732_b1 , \2524_b1 , \2527_b1 );
not ( \2527_b1 , w_4580 );
and ( \2732_b0 , \2524_b0 , w_4581 );
and ( w_4580 , w_4581 , \2527_b0 );
or ( \2733_b1 , \2731_b1 , w_4582 );
or ( \2733_b0 , \2731_b0 , \2732_b0 );
not ( \2732_b0 , w_4583 );
and ( w_4583 , w_4582 , \2732_b1 );
or ( \2734_b1 , \2730_b1 , \2733_b1 );
xor ( \2734_b0 , \2730_b0 , w_4584 );
not ( w_4584 , w_4585 );
and ( w_4585 , \2733_b1 , \2733_b0 );
or ( \2735_b1 , \1963_A[11]_b1 , \1127_B[4]_b1 );
not ( \1127_B[4]_b1 , w_4586 );
and ( \2735_b0 , \1963_A[11]_b0 , w_4587 );
and ( w_4586 , w_4587 , \1127_B[4]_b0 );
or ( \2736_b1 , \2734_b1 , \2735_b1 );
xor ( \2736_b0 , \2734_b0 , w_4588 );
not ( w_4588 , w_4589 );
and ( w_4589 , \2735_b1 , \2735_b0 );
or ( \2737_b1 , \2528_b1 , \2529_b1 );
not ( \2529_b1 , w_4590 );
and ( \2737_b0 , \2528_b0 , w_4591 );
and ( w_4590 , w_4591 , \2529_b0 );
or ( \2738_b1 , \2530_b1 , \2533_b1 );
not ( \2533_b1 , w_4592 );
and ( \2738_b0 , \2530_b0 , w_4593 );
and ( w_4592 , w_4593 , \2533_b0 );
or ( \2739_b1 , \2737_b1 , w_4594 );
or ( \2739_b0 , \2737_b0 , \2738_b0 );
not ( \2738_b0 , w_4595 );
and ( w_4595 , w_4594 , \2738_b1 );
or ( \2740_b1 , \2736_b1 , \2739_b1 );
xor ( \2740_b0 , \2736_b0 , w_4596 );
not ( w_4596 , w_4597 );
and ( w_4597 , \2739_b1 , \2739_b0 );
or ( \2741_b1 , \1805_A[10]_b1 , \1219_B[5]_b1 );
not ( \1219_B[5]_b1 , w_4598 );
and ( \2741_b0 , \1805_A[10]_b0 , w_4599 );
and ( w_4598 , w_4599 , \1219_B[5]_b0 );
or ( \2742_b1 , \2740_b1 , \2741_b1 );
xor ( \2742_b0 , \2740_b0 , w_4600 );
not ( w_4600 , w_4601 );
and ( w_4601 , \2741_b1 , \2741_b0 );
or ( \2743_b1 , \2534_b1 , \2535_b1 );
not ( \2535_b1 , w_4602 );
and ( \2743_b0 , \2534_b0 , w_4603 );
and ( w_4602 , w_4603 , \2535_b0 );
or ( \2744_b1 , \2536_b1 , \2539_b1 );
not ( \2539_b1 , w_4604 );
and ( \2744_b0 , \2536_b0 , w_4605 );
and ( w_4604 , w_4605 , \2539_b0 );
or ( \2745_b1 , \2743_b1 , w_4606 );
or ( \2745_b0 , \2743_b0 , \2744_b0 );
not ( \2744_b0 , w_4607 );
and ( w_4607 , w_4606 , \2744_b1 );
or ( \2746_b1 , \2742_b1 , \2745_b1 );
xor ( \2746_b0 , \2742_b0 , w_4608 );
not ( w_4608 , w_4609 );
and ( w_4609 , \2745_b1 , \2745_b0 );
or ( \2747_b1 , \1659_A[9]_b1 , \1323_B[6]_b1 );
not ( \1323_B[6]_b1 , w_4610 );
and ( \2747_b0 , \1659_A[9]_b0 , w_4611 );
and ( w_4610 , w_4611 , \1323_B[6]_b0 );
or ( \2748_b1 , \2746_b1 , \2747_b1 );
xor ( \2748_b0 , \2746_b0 , w_4612 );
not ( w_4612 , w_4613 );
and ( w_4613 , \2747_b1 , \2747_b0 );
or ( \2749_b1 , \2540_b1 , \2541_b1 );
not ( \2541_b1 , w_4614 );
and ( \2749_b0 , \2540_b0 , w_4615 );
and ( w_4614 , w_4615 , \2541_b0 );
or ( \2750_b1 , \2542_b1 , \2545_b1 );
not ( \2545_b1 , w_4616 );
and ( \2750_b0 , \2542_b0 , w_4617 );
and ( w_4616 , w_4617 , \2545_b0 );
or ( \2751_b1 , \2749_b1 , w_4618 );
or ( \2751_b0 , \2749_b0 , \2750_b0 );
not ( \2750_b0 , w_4619 );
and ( w_4619 , w_4618 , \2750_b1 );
or ( \2752_b1 , \2748_b1 , \2751_b1 );
xor ( \2752_b0 , \2748_b0 , w_4620 );
not ( w_4620 , w_4621 );
and ( w_4621 , \2751_b1 , \2751_b0 );
or ( \2753_b1 , \1525_A[8]_b1 , \1439_B[7]_b1 );
not ( \1439_B[7]_b1 , w_4622 );
and ( \2753_b0 , \1525_A[8]_b0 , w_4623 );
and ( w_4622 , w_4623 , \1439_B[7]_b0 );
or ( \2754_b1 , \2752_b1 , \2753_b1 );
xor ( \2754_b0 , \2752_b0 , w_4624 );
not ( w_4624 , w_4625 );
and ( w_4625 , \2753_b1 , \2753_b0 );
or ( \2755_b1 , \2546_b1 , \2547_b1 );
not ( \2547_b1 , w_4626 );
and ( \2755_b0 , \2546_b0 , w_4627 );
and ( w_4626 , w_4627 , \2547_b0 );
or ( \2756_b1 , \2548_b1 , \2551_b1 );
not ( \2551_b1 , w_4628 );
and ( \2756_b0 , \2548_b0 , w_4629 );
and ( w_4628 , w_4629 , \2551_b0 );
or ( \2757_b1 , \2755_b1 , w_4630 );
or ( \2757_b0 , \2755_b0 , \2756_b0 );
not ( \2756_b0 , w_4631 );
and ( w_4631 , w_4630 , \2756_b1 );
or ( \2758_b1 , \2754_b1 , \2757_b1 );
xor ( \2758_b0 , \2754_b0 , w_4632 );
not ( w_4632 , w_4633 );
and ( w_4633 , \2757_b1 , \2757_b0 );
or ( \2759_b1 , \1403_A[7]_b1 , \1567_B[8]_b1 );
not ( \1567_B[8]_b1 , w_4634 );
and ( \2759_b0 , \1403_A[7]_b0 , w_4635 );
and ( w_4634 , w_4635 , \1567_B[8]_b0 );
or ( \2760_b1 , \2758_b1 , \2759_b1 );
xor ( \2760_b0 , \2758_b0 , w_4636 );
not ( w_4636 , w_4637 );
and ( w_4637 , \2759_b1 , \2759_b0 );
or ( \2761_b1 , \2552_b1 , \2553_b1 );
not ( \2553_b1 , w_4638 );
and ( \2761_b0 , \2552_b0 , w_4639 );
and ( w_4638 , w_4639 , \2553_b0 );
or ( \2762_b1 , \2554_b1 , \2557_b1 );
not ( \2557_b1 , w_4640 );
and ( \2762_b0 , \2554_b0 , w_4641 );
and ( w_4640 , w_4641 , \2557_b0 );
or ( \2763_b1 , \2761_b1 , w_4642 );
or ( \2763_b0 , \2761_b0 , \2762_b0 );
not ( \2762_b0 , w_4643 );
and ( w_4643 , w_4642 , \2762_b1 );
or ( \2764_b1 , \2760_b1 , \2763_b1 );
xor ( \2764_b0 , \2760_b0 , w_4644 );
not ( w_4644 , w_4645 );
and ( w_4645 , \2763_b1 , \2763_b0 );
or ( \2765_b1 , \1293_A[6]_b1 , \1707_B[9]_b1 );
not ( \1707_B[9]_b1 , w_4646 );
and ( \2765_b0 , \1293_A[6]_b0 , w_4647 );
and ( w_4646 , w_4647 , \1707_B[9]_b0 );
or ( \2766_b1 , \2764_b1 , \2765_b1 );
xor ( \2766_b0 , \2764_b0 , w_4648 );
not ( w_4648 , w_4649 );
and ( w_4649 , \2765_b1 , \2765_b0 );
or ( \2767_b1 , \2558_b1 , \2559_b1 );
not ( \2559_b1 , w_4650 );
and ( \2767_b0 , \2558_b0 , w_4651 );
and ( w_4650 , w_4651 , \2559_b0 );
or ( \2768_b1 , \2560_b1 , \2563_b1 );
not ( \2563_b1 , w_4652 );
and ( \2768_b0 , \2560_b0 , w_4653 );
and ( w_4652 , w_4653 , \2563_b0 );
or ( \2769_b1 , \2767_b1 , w_4654 );
or ( \2769_b0 , \2767_b0 , \2768_b0 );
not ( \2768_b0 , w_4655 );
and ( w_4655 , w_4654 , \2768_b1 );
or ( \2770_b1 , \2766_b1 , \2769_b1 );
xor ( \2770_b0 , \2766_b0 , w_4656 );
not ( w_4656 , w_4657 );
and ( w_4657 , \2769_b1 , \2769_b0 );
or ( \2771_b1 , \1195_A[5]_b1 , \1859_B[10]_b1 );
not ( \1859_B[10]_b1 , w_4658 );
and ( \2771_b0 , \1195_A[5]_b0 , w_4659 );
and ( w_4658 , w_4659 , \1859_B[10]_b0 );
or ( \2772_b1 , \2770_b1 , \2771_b1 );
xor ( \2772_b0 , \2770_b0 , w_4660 );
not ( w_4660 , w_4661 );
and ( w_4661 , \2771_b1 , \2771_b0 );
or ( \2773_b1 , \2564_b1 , \2565_b1 );
not ( \2565_b1 , w_4662 );
and ( \2773_b0 , \2564_b0 , w_4663 );
and ( w_4662 , w_4663 , \2565_b0 );
or ( \2774_b1 , \2566_b1 , \2569_b1 );
not ( \2569_b1 , w_4664 );
and ( \2774_b0 , \2566_b0 , w_4665 );
and ( w_4664 , w_4665 , \2569_b0 );
or ( \2775_b1 , \2773_b1 , w_4666 );
or ( \2775_b0 , \2773_b0 , \2774_b0 );
not ( \2774_b0 , w_4667 );
and ( w_4667 , w_4666 , \2774_b1 );
or ( \2776_b1 , \2772_b1 , \2775_b1 );
xor ( \2776_b0 , \2772_b0 , w_4668 );
not ( w_4668 , w_4669 );
and ( w_4669 , \2775_b1 , \2775_b0 );
or ( \2777_b1 , \1109_A[4]_b1 , \2023_B[11]_b1 );
not ( \2023_B[11]_b1 , w_4670 );
and ( \2777_b0 , \1109_A[4]_b0 , w_4671 );
and ( w_4670 , w_4671 , \2023_B[11]_b0 );
or ( \2778_b1 , \2776_b1 , \2777_b1 );
xor ( \2778_b0 , \2776_b0 , w_4672 );
not ( w_4672 , w_4673 );
and ( w_4673 , \2777_b1 , \2777_b0 );
or ( \2779_b1 , \2570_b1 , \2571_b1 );
not ( \2571_b1 , w_4674 );
and ( \2779_b0 , \2570_b0 , w_4675 );
and ( w_4674 , w_4675 , \2571_b0 );
or ( \2780_b1 , \2572_b1 , \2575_b1 );
not ( \2575_b1 , w_4676 );
and ( \2780_b0 , \2572_b0 , w_4677 );
and ( w_4676 , w_4677 , \2575_b0 );
or ( \2781_b1 , \2779_b1 , w_4678 );
or ( \2781_b0 , \2779_b0 , \2780_b0 );
not ( \2780_b0 , w_4679 );
and ( w_4679 , w_4678 , \2780_b1 );
or ( \2782_b1 , \2778_b1 , \2781_b1 );
xor ( \2782_b0 , \2778_b0 , w_4680 );
not ( w_4680 , w_4681 );
and ( w_4681 , \2781_b1 , \2781_b0 );
or ( \2783_b1 , \1035_A[3]_b1 , \2199_B[12]_b1 );
not ( \2199_B[12]_b1 , w_4682 );
and ( \2783_b0 , \1035_A[3]_b0 , w_4683 );
and ( w_4682 , w_4683 , \2199_B[12]_b0 );
or ( \2784_b1 , \2782_b1 , \2783_b1 );
xor ( \2784_b0 , \2782_b0 , w_4684 );
not ( w_4684 , w_4685 );
and ( w_4685 , \2783_b1 , \2783_b0 );
or ( \2785_b1 , \2576_b1 , \2577_b1 );
not ( \2577_b1 , w_4686 );
and ( \2785_b0 , \2576_b0 , w_4687 );
and ( w_4686 , w_4687 , \2577_b0 );
or ( \2786_b1 , \2578_b1 , \2581_b1 );
not ( \2581_b1 , w_4688 );
and ( \2786_b0 , \2578_b0 , w_4689 );
and ( w_4688 , w_4689 , \2581_b0 );
or ( \2787_b1 , \2785_b1 , w_4690 );
or ( \2787_b0 , \2785_b0 , \2786_b0 );
not ( \2786_b0 , w_4691 );
and ( w_4691 , w_4690 , \2786_b1 );
or ( \2788_b1 , \2784_b1 , \2787_b1 );
xor ( \2788_b0 , \2784_b0 , w_4692 );
not ( w_4692 , w_4693 );
and ( w_4693 , \2787_b1 , \2787_b0 );
or ( \2789_b1 , \973_A[2]_b1 , \2387_B[13]_b1 );
not ( \2387_B[13]_b1 , w_4694 );
and ( \2789_b0 , \973_A[2]_b0 , w_4695 );
and ( w_4694 , w_4695 , \2387_B[13]_b0 );
or ( \2790_b1 , \2788_b1 , \2789_b1 );
xor ( \2790_b0 , \2788_b0 , w_4696 );
not ( w_4696 , w_4697 );
and ( w_4697 , \2789_b1 , \2789_b0 );
or ( \2791_b1 , \2582_b1 , \2583_b1 );
not ( \2583_b1 , w_4698 );
and ( \2791_b0 , \2582_b0 , w_4699 );
and ( w_4698 , w_4699 , \2583_b0 );
or ( \2792_b1 , \2584_b1 , \2585_b1 );
not ( \2585_b1 , w_4700 );
and ( \2792_b0 , \2584_b0 , w_4701 );
and ( w_4700 , w_4701 , \2585_b0 );
or ( \2793_b1 , \2791_b1 , w_4702 );
or ( \2793_b0 , \2791_b0 , \2792_b0 );
not ( \2792_b0 , w_4703 );
and ( w_4703 , w_4702 , \2792_b1 );
or ( \2794_b1 , \2790_b1 , \2793_b1 );
xor ( \2794_b0 , \2790_b0 , w_4704 );
not ( w_4704 , w_4705 );
and ( w_4705 , \2793_b1 , \2793_b0 );
or ( \2795_b1 , \927_A[1]_b1 , \2587_B[14]_b1 );
not ( \2587_B[14]_b1 , w_4706 );
and ( \2795_b0 , \927_A[1]_b0 , w_4707 );
and ( w_4706 , w_4707 , \2587_B[14]_b0 );
or ( \2796_b1 , \2794_b1 , \2795_b1 );
xor ( \2796_b0 , \2794_b0 , w_4708 );
not ( w_4708 , w_4709 );
and ( w_4709 , \2795_b1 , \2795_b0 );
or ( \2797_b1 , \2586_b1 , \2588_b1 );
not ( \2588_b1 , w_4710 );
and ( \2797_b0 , \2586_b0 , w_4711 );
and ( w_4710 , w_4711 , \2588_b0 );
or ( \2798_b1 , \2796_b1 , \2797_b1 );
xor ( \2798_b0 , \2796_b0 , w_4712 );
not ( w_4712 , w_4713 );
and ( w_4713 , \2797_b1 , \2797_b0 );
buf ( \2799_B[15]_b1 , \d[15]_b1 );
buf ( \2799_B[15]_b0 , \d[15]_b0 );
or ( \2800_b1 , \891_A[0]_b1 , \2799_B[15]_b1 );
not ( \2799_B[15]_b1 , w_4714 );
and ( \2800_b0 , \891_A[0]_b0 , w_4715 );
and ( w_4714 , w_4715 , \2799_B[15]_b0 );
or ( \2801_b1 , \2798_b1 , \2800_b1 );
xor ( \2801_b0 , \2798_b0 , w_4716 );
not ( w_4716 , w_4717 );
and ( w_4717 , \2800_b1 , \2800_b0 );
buf ( \2802_Z[15]_b1 , \2801_b1 );
buf ( \2802_Z[15]_b0 , \2801_b0 );
or ( \2803_b1 , \2802_Z[15]_b1 , \865_b1 );
not ( \865_b1 , w_4718 );
and ( \2803_b0 , \2802_Z[15]_b0 , w_4719 );
and ( w_4718 , w_4719 , \865_b0 );
buf ( \2804_A[15]_b1 , \b[15]_b1 );
buf ( \2804_A[15]_b0 , \b[15]_b0 );
buf ( \2805_B[15]_b1 , \d[15]_b1 );
buf ( \2805_B[15]_b0 , \d[15]_b0 );
or ( \2806_b1 , \2804_A[15]_b1 , \2805_B[15]_b1 );
xor ( \2806_b0 , \2804_A[15]_b0 , w_4720 );
not ( w_4720 , w_4721 );
and ( w_4721 , \2805_B[15]_b1 , \2805_B[15]_b0 );
or ( \2807_b1 , \2592_A[14]_b1 , \2593_B[14]_b1 );
not ( \2593_B[14]_b1 , w_4722 );
and ( \2807_b0 , \2592_A[14]_b0 , w_4723 );
and ( w_4722 , w_4723 , \2593_B[14]_b0 );
or ( \2808_b1 , \2593_B[14]_b1 , \2598_b1 );
not ( \2598_b1 , w_4724 );
and ( \2808_b0 , \2593_B[14]_b0 , w_4725 );
and ( w_4724 , w_4725 , \2598_b0 );
or ( \2809_b1 , \2592_A[14]_b1 , \2598_b1 );
not ( \2598_b1 , w_4726 );
and ( \2809_b0 , \2592_A[14]_b0 , w_4727 );
and ( w_4726 , w_4727 , \2598_b0 );
or ( \2811_b1 , \2806_b1 , \2810_b1 );
xor ( \2811_b0 , \2806_b0 , w_4728 );
not ( w_4728 , w_4729 );
and ( w_4729 , \2810_b1 , \2810_b0 );
buf ( \2812_SUM[15]_b1 , \2811_b1 );
buf ( \2812_SUM[15]_b0 , \2811_b0 );
or ( \2813_b1 , \2812_SUM[15]_b1 , \863_b1 );
not ( \863_b1 , w_4730 );
and ( \2813_b0 , \2812_SUM[15]_b0 , w_4731 );
and ( w_4730 , w_4731 , \863_b0 );
buf ( \2814_A[15]_b1 , \a[15]_b1 );
buf ( \2814_A[15]_b0 , \a[15]_b0 );
buf ( \2815_B[15]_b1 , \c[15]_b1 );
buf ( \2815_B[15]_b0 , \c[15]_b0 );
or ( \2816_b1 , \2814_A[15]_b1 , \2815_B[15]_b1 );
xor ( \2816_b0 , \2814_A[15]_b0 , w_4732 );
not ( w_4732 , w_4733 );
and ( w_4733 , \2815_B[15]_b1 , \2815_B[15]_b0 );
or ( \2817_b1 , \2602_A[14]_b1 , \2603_B[14]_b1 );
not ( \2603_B[14]_b1 , w_4734 );
and ( \2817_b0 , \2602_A[14]_b0 , w_4735 );
and ( w_4734 , w_4735 , \2603_B[14]_b0 );
or ( \2818_b1 , \2603_B[14]_b1 , \2608_b1 );
not ( \2608_b1 , w_4736 );
and ( \2818_b0 , \2603_B[14]_b0 , w_4737 );
and ( w_4736 , w_4737 , \2608_b0 );
or ( \2819_b1 , \2602_A[14]_b1 , \2608_b1 );
not ( \2608_b1 , w_4738 );
and ( \2819_b0 , \2602_A[14]_b0 , w_4739 );
and ( w_4738 , w_4739 , \2608_b0 );
or ( \2821_b1 , \2816_b1 , \2820_b1 );
xor ( \2821_b0 , \2816_b0 , w_4740 );
not ( w_4740 , w_4741 );
and ( w_4741 , \2820_b1 , \2820_b0 );
buf ( \2822_SUM[15]_b1 , \2821_b1 );
buf ( \2822_SUM[15]_b0 , \2821_b0 );
or ( \2823_b1 , \2822_SUM[15]_b1 , \861_b1 );
not ( \861_b1 , w_4742 );
and ( \2823_b0 , \2822_SUM[15]_b0 , w_4743 );
and ( w_4742 , w_4743 , \861_b0 );
or ( \2824_b1 , \d[15]_b1 , \859_b1 );
not ( \859_b1 , w_4744 );
and ( \2824_b0 , \d[15]_b0 , w_4745 );
and ( w_4744 , w_4745 , \859_b0 );
or ( \2825_b1 , \c[15]_b1 , \857_b1 );
not ( \857_b1 , w_4746 );
and ( \2825_b0 , \c[15]_b0 , w_4747 );
and ( w_4746 , w_4747 , \857_b0 );
or ( \2826_b1 , \b[15]_b1 , \855_b1 );
not ( \855_b1 , w_4748 );
and ( \2826_b0 , \b[15]_b0 , w_4749 );
and ( w_4748 , w_4749 , \855_b0 );
or ( \2827_b1 , \a[15]_b1 , \853_b1 );
not ( \853_b1 , w_4750 );
and ( \2827_b0 , \a[15]_b0 , w_4751 );
and ( w_4750 , w_4751 , \853_b0 );
buf ( \2829_A[15]_b1 , \c[15]_b1 );
buf ( \2829_A[15]_b0 , \c[15]_b0 );
buf ( \2830_B[15]_b1 , \d[15]_b1 );
buf ( \2830_B[15]_b0 , \d[15]_b0 );
or ( \2831_b1 , \2829_A[15]_b1 , \2830_B[15]_b1 );
not ( \2830_B[15]_b1 , w_4752 );
and ( \2831_b0 , \2829_A[15]_b0 , w_4753 );
and ( w_4752 , w_4753 , \2830_B[15]_b0 );
buf ( \2832_A[14]_b1 , \c[14]_b1 );
buf ( \2832_A[14]_b0 , \c[14]_b0 );
buf ( \2833_B[14]_b1 , \d[14]_b1 );
buf ( \2833_B[14]_b0 , \d[14]_b0 );
or ( \2834_b1 , \2832_A[14]_b1 , \2833_B[14]_b1 );
not ( \2833_B[14]_b1 , w_4754 );
and ( \2834_b0 , \2832_A[14]_b0 , w_4755 );
and ( w_4754 , w_4755 , \2833_B[14]_b0 );
buf ( \2835_A[13]_b1 , \c[13]_b1 );
buf ( \2835_A[13]_b0 , \c[13]_b0 );
buf ( \2836_B[13]_b1 , \d[13]_b1 );
buf ( \2836_B[13]_b0 , \d[13]_b0 );
or ( \2837_b1 , \2835_A[13]_b1 , \2836_B[13]_b1 );
not ( \2836_B[13]_b1 , w_4756 );
and ( \2837_b0 , \2835_A[13]_b0 , w_4757 );
and ( w_4756 , w_4757 , \2836_B[13]_b0 );
buf ( \2838_A[12]_b1 , \c[12]_b1 );
buf ( \2838_A[12]_b0 , \c[12]_b0 );
buf ( \2839_B[12]_b1 , \d[12]_b1 );
buf ( \2839_B[12]_b0 , \d[12]_b0 );
or ( \2840_b1 , \2838_A[12]_b1 , \2839_B[12]_b1 );
not ( \2839_B[12]_b1 , w_4758 );
and ( \2840_b0 , \2838_A[12]_b0 , w_4759 );
and ( w_4758 , w_4759 , \2839_B[12]_b0 );
buf ( \2841_A[11]_b1 , \c[11]_b1 );
buf ( \2841_A[11]_b0 , \c[11]_b0 );
buf ( \2842_B[11]_b1 , \d[11]_b1 );
buf ( \2842_B[11]_b0 , \d[11]_b0 );
or ( \2843_b1 , \2841_A[11]_b1 , \2842_B[11]_b1 );
not ( \2842_B[11]_b1 , w_4760 );
and ( \2843_b0 , \2841_A[11]_b0 , w_4761 );
and ( w_4760 , w_4761 , \2842_B[11]_b0 );
buf ( \2844_A[10]_b1 , \c[10]_b1 );
buf ( \2844_A[10]_b0 , \c[10]_b0 );
buf ( \2845_B[10]_b1 , \d[10]_b1 );
buf ( \2845_B[10]_b0 , \d[10]_b0 );
or ( \2846_b1 , \2844_A[10]_b1 , \2845_B[10]_b1 );
not ( \2845_B[10]_b1 , w_4762 );
and ( \2846_b0 , \2844_A[10]_b0 , w_4763 );
and ( w_4762 , w_4763 , \2845_B[10]_b0 );
buf ( \2847_A[9]_b1 , \c[9]_b1 );
buf ( \2847_A[9]_b0 , \c[9]_b0 );
buf ( \2848_B[9]_b1 , \d[9]_b1 );
buf ( \2848_B[9]_b0 , \d[9]_b0 );
or ( \2849_b1 , \2847_A[9]_b1 , \2848_B[9]_b1 );
not ( \2848_B[9]_b1 , w_4764 );
and ( \2849_b0 , \2847_A[9]_b0 , w_4765 );
and ( w_4764 , w_4765 , \2848_B[9]_b0 );
buf ( \2850_A[8]_b1 , \c[8]_b1 );
buf ( \2850_A[8]_b0 , \c[8]_b0 );
buf ( \2851_B[8]_b1 , \d[8]_b1 );
buf ( \2851_B[8]_b0 , \d[8]_b0 );
or ( \2852_b1 , \2850_A[8]_b1 , \2851_B[8]_b1 );
not ( \2851_B[8]_b1 , w_4766 );
and ( \2852_b0 , \2850_A[8]_b0 , w_4767 );
and ( w_4766 , w_4767 , \2851_B[8]_b0 );
buf ( \2853_A[7]_b1 , \c[7]_b1 );
buf ( \2853_A[7]_b0 , \c[7]_b0 );
buf ( \2854_B[7]_b1 , \d[7]_b1 );
buf ( \2854_B[7]_b0 , \d[7]_b0 );
or ( \2855_b1 , \2853_A[7]_b1 , \2854_B[7]_b1 );
not ( \2854_B[7]_b1 , w_4768 );
and ( \2855_b0 , \2853_A[7]_b0 , w_4769 );
and ( w_4768 , w_4769 , \2854_B[7]_b0 );
buf ( \2856_A[6]_b1 , \c[6]_b1 );
buf ( \2856_A[6]_b0 , \c[6]_b0 );
buf ( \2857_B[6]_b1 , \d[6]_b1 );
buf ( \2857_B[6]_b0 , \d[6]_b0 );
or ( \2858_b1 , \2856_A[6]_b1 , \2857_B[6]_b1 );
not ( \2857_B[6]_b1 , w_4770 );
and ( \2858_b0 , \2856_A[6]_b0 , w_4771 );
and ( w_4770 , w_4771 , \2857_B[6]_b0 );
buf ( \2859_A[5]_b1 , \c[5]_b1 );
buf ( \2859_A[5]_b0 , \c[5]_b0 );
buf ( \2860_B[5]_b1 , \d[5]_b1 );
buf ( \2860_B[5]_b0 , \d[5]_b0 );
or ( \2861_b1 , \2859_A[5]_b1 , \2860_B[5]_b1 );
not ( \2860_B[5]_b1 , w_4772 );
and ( \2861_b0 , \2859_A[5]_b0 , w_4773 );
and ( w_4772 , w_4773 , \2860_B[5]_b0 );
buf ( \2862_A[4]_b1 , \c[4]_b1 );
buf ( \2862_A[4]_b0 , \c[4]_b0 );
buf ( \2863_B[4]_b1 , \d[4]_b1 );
buf ( \2863_B[4]_b0 , \d[4]_b0 );
or ( \2864_b1 , \2862_A[4]_b1 , \2863_B[4]_b1 );
not ( \2863_B[4]_b1 , w_4774 );
and ( \2864_b0 , \2862_A[4]_b0 , w_4775 );
and ( w_4774 , w_4775 , \2863_B[4]_b0 );
buf ( \2865_A[3]_b1 , \c[3]_b1 );
buf ( \2865_A[3]_b0 , \c[3]_b0 );
buf ( \2866_B[3]_b1 , \d[3]_b1 );
buf ( \2866_B[3]_b0 , \d[3]_b0 );
or ( \2867_b1 , \2865_A[3]_b1 , \2866_B[3]_b1 );
not ( \2866_B[3]_b1 , w_4776 );
and ( \2867_b0 , \2865_A[3]_b0 , w_4777 );
and ( w_4776 , w_4777 , \2866_B[3]_b0 );
buf ( \2868_A[2]_b1 , \c[2]_b1 );
buf ( \2868_A[2]_b0 , \c[2]_b0 );
buf ( \2869_B[2]_b1 , \d[2]_b1 );
buf ( \2869_B[2]_b0 , \d[2]_b0 );
or ( \2870_b1 , \2868_A[2]_b1 , \2869_B[2]_b1 );
not ( \2869_B[2]_b1 , w_4778 );
and ( \2870_b0 , \2868_A[2]_b0 , w_4779 );
and ( w_4778 , w_4779 , \2869_B[2]_b0 );
buf ( \2871_A[1]_b1 , \c[1]_b1 );
buf ( \2871_A[1]_b0 , \c[1]_b0 );
buf ( \2872_B[1]_b1 , \d[1]_b1 );
buf ( \2872_B[1]_b0 , \d[1]_b0 );
or ( \2873_b1 , \2871_A[1]_b1 , \2872_B[1]_b1 );
not ( \2872_B[1]_b1 , w_4780 );
and ( \2873_b0 , \2871_A[1]_b0 , w_4781 );
and ( w_4780 , w_4781 , \2872_B[1]_b0 );
buf ( \2874_A[0]_b1 , \c[0]_b1 );
buf ( \2874_A[0]_b0 , \c[0]_b0 );
buf ( \2875_B[0]_b1 , \d[0]_b1 );
buf ( \2875_B[0]_b0 , \d[0]_b0 );
or ( \2876_b1 , \2874_A[0]_b1 , \2875_B[0]_b1 );
not ( \2875_B[0]_b1 , w_4782 );
and ( \2876_b0 , \2874_A[0]_b0 , w_4783 );
and ( w_4782 , w_4783 , \2875_B[0]_b0 );
or ( \2877_b1 , \2872_B[1]_b1 , \2876_b1 );
not ( \2876_b1 , w_4784 );
and ( \2877_b0 , \2872_B[1]_b0 , w_4785 );
and ( w_4784 , w_4785 , \2876_b0 );
or ( \2878_b1 , \2871_A[1]_b1 , \2876_b1 );
not ( \2876_b1 , w_4786 );
and ( \2878_b0 , \2871_A[1]_b0 , w_4787 );
and ( w_4786 , w_4787 , \2876_b0 );
or ( \2880_b1 , \2869_B[2]_b1 , \2879_b1 );
not ( \2879_b1 , w_4788 );
and ( \2880_b0 , \2869_B[2]_b0 , w_4789 );
and ( w_4788 , w_4789 , \2879_b0 );
or ( \2881_b1 , \2868_A[2]_b1 , \2879_b1 );
not ( \2879_b1 , w_4790 );
and ( \2881_b0 , \2868_A[2]_b0 , w_4791 );
and ( w_4790 , w_4791 , \2879_b0 );
or ( \2883_b1 , \2866_B[3]_b1 , \2882_b1 );
not ( \2882_b1 , w_4792 );
and ( \2883_b0 , \2866_B[3]_b0 , w_4793 );
and ( w_4792 , w_4793 , \2882_b0 );
or ( \2884_b1 , \2865_A[3]_b1 , \2882_b1 );
not ( \2882_b1 , w_4794 );
and ( \2884_b0 , \2865_A[3]_b0 , w_4795 );
and ( w_4794 , w_4795 , \2882_b0 );
or ( \2886_b1 , \2863_B[4]_b1 , \2885_b1 );
not ( \2885_b1 , w_4796 );
and ( \2886_b0 , \2863_B[4]_b0 , w_4797 );
and ( w_4796 , w_4797 , \2885_b0 );
or ( \2887_b1 , \2862_A[4]_b1 , \2885_b1 );
not ( \2885_b1 , w_4798 );
and ( \2887_b0 , \2862_A[4]_b0 , w_4799 );
and ( w_4798 , w_4799 , \2885_b0 );
or ( \2889_b1 , \2860_B[5]_b1 , \2888_b1 );
not ( \2888_b1 , w_4800 );
and ( \2889_b0 , \2860_B[5]_b0 , w_4801 );
and ( w_4800 , w_4801 , \2888_b0 );
or ( \2890_b1 , \2859_A[5]_b1 , \2888_b1 );
not ( \2888_b1 , w_4802 );
and ( \2890_b0 , \2859_A[5]_b0 , w_4803 );
and ( w_4802 , w_4803 , \2888_b0 );
or ( \2892_b1 , \2857_B[6]_b1 , \2891_b1 );
not ( \2891_b1 , w_4804 );
and ( \2892_b0 , \2857_B[6]_b0 , w_4805 );
and ( w_4804 , w_4805 , \2891_b0 );
or ( \2893_b1 , \2856_A[6]_b1 , \2891_b1 );
not ( \2891_b1 , w_4806 );
and ( \2893_b0 , \2856_A[6]_b0 , w_4807 );
and ( w_4806 , w_4807 , \2891_b0 );
or ( \2895_b1 , \2854_B[7]_b1 , \2894_b1 );
not ( \2894_b1 , w_4808 );
and ( \2895_b0 , \2854_B[7]_b0 , w_4809 );
and ( w_4808 , w_4809 , \2894_b0 );
or ( \2896_b1 , \2853_A[7]_b1 , \2894_b1 );
not ( \2894_b1 , w_4810 );
and ( \2896_b0 , \2853_A[7]_b0 , w_4811 );
and ( w_4810 , w_4811 , \2894_b0 );
or ( \2898_b1 , \2851_B[8]_b1 , \2897_b1 );
not ( \2897_b1 , w_4812 );
and ( \2898_b0 , \2851_B[8]_b0 , w_4813 );
and ( w_4812 , w_4813 , \2897_b0 );
or ( \2899_b1 , \2850_A[8]_b1 , \2897_b1 );
not ( \2897_b1 , w_4814 );
and ( \2899_b0 , \2850_A[8]_b0 , w_4815 );
and ( w_4814 , w_4815 , \2897_b0 );
or ( \2901_b1 , \2848_B[9]_b1 , \2900_b1 );
not ( \2900_b1 , w_4816 );
and ( \2901_b0 , \2848_B[9]_b0 , w_4817 );
and ( w_4816 , w_4817 , \2900_b0 );
or ( \2902_b1 , \2847_A[9]_b1 , \2900_b1 );
not ( \2900_b1 , w_4818 );
and ( \2902_b0 , \2847_A[9]_b0 , w_4819 );
and ( w_4818 , w_4819 , \2900_b0 );
or ( \2904_b1 , \2845_B[10]_b1 , \2903_b1 );
not ( \2903_b1 , w_4820 );
and ( \2904_b0 , \2845_B[10]_b0 , w_4821 );
and ( w_4820 , w_4821 , \2903_b0 );
or ( \2905_b1 , \2844_A[10]_b1 , \2903_b1 );
not ( \2903_b1 , w_4822 );
and ( \2905_b0 , \2844_A[10]_b0 , w_4823 );
and ( w_4822 , w_4823 , \2903_b0 );
or ( \2907_b1 , \2842_B[11]_b1 , \2906_b1 );
not ( \2906_b1 , w_4824 );
and ( \2907_b0 , \2842_B[11]_b0 , w_4825 );
and ( w_4824 , w_4825 , \2906_b0 );
or ( \2908_b1 , \2841_A[11]_b1 , \2906_b1 );
not ( \2906_b1 , w_4826 );
and ( \2908_b0 , \2841_A[11]_b0 , w_4827 );
and ( w_4826 , w_4827 , \2906_b0 );
or ( \2910_b1 , \2839_B[12]_b1 , \2909_b1 );
not ( \2909_b1 , w_4828 );
and ( \2910_b0 , \2839_B[12]_b0 , w_4829 );
and ( w_4828 , w_4829 , \2909_b0 );
or ( \2911_b1 , \2838_A[12]_b1 , \2909_b1 );
not ( \2909_b1 , w_4830 );
and ( \2911_b0 , \2838_A[12]_b0 , w_4831 );
and ( w_4830 , w_4831 , \2909_b0 );
or ( \2913_b1 , \2836_B[13]_b1 , \2912_b1 );
not ( \2912_b1 , w_4832 );
and ( \2913_b0 , \2836_B[13]_b0 , w_4833 );
and ( w_4832 , w_4833 , \2912_b0 );
or ( \2914_b1 , \2835_A[13]_b1 , \2912_b1 );
not ( \2912_b1 , w_4834 );
and ( \2914_b0 , \2835_A[13]_b0 , w_4835 );
and ( w_4834 , w_4835 , \2912_b0 );
or ( \2916_b1 , \2833_B[14]_b1 , \2915_b1 );
not ( \2915_b1 , w_4836 );
and ( \2916_b0 , \2833_B[14]_b0 , w_4837 );
and ( w_4836 , w_4837 , \2915_b0 );
or ( \2917_b1 , \2832_A[14]_b1 , \2915_b1 );
not ( \2915_b1 , w_4838 );
and ( \2917_b0 , \2832_A[14]_b0 , w_4839 );
and ( w_4838 , w_4839 , \2915_b0 );
or ( \2919_b1 , \2830_B[15]_b1 , \2918_b1 );
not ( \2918_b1 , w_4840 );
and ( \2919_b0 , \2830_B[15]_b0 , w_4841 );
and ( w_4840 , w_4841 , \2918_b0 );
or ( \2920_b1 , \2829_A[15]_b1 , \2918_b1 );
not ( \2918_b1 , w_4842 );
and ( \2920_b0 , \2829_A[15]_b0 , w_4843 );
and ( w_4842 , w_4843 , \2918_b0 );
buf ( \2922_SUM[16]_b1 , \2921_b1 );
buf ( \2922_SUM[16]_b0 , \2921_b0 );
buf ( \2923_A[16]_b1 , \2922_SUM[16]_b1 );
buf ( \2923_A[16]_b0 , \2922_SUM[16]_b0 );
or ( \2924_b1 , \2829_A[15]_b1 , \2830_B[15]_b1 );
xor ( \2924_b0 , \2829_A[15]_b0 , w_4844 );
not ( w_4844 , w_4845 );
and ( w_4845 , \2830_B[15]_b1 , \2830_B[15]_b0 );
or ( \2925_b1 , \2924_b1 , \2918_b1 );
xor ( \2925_b0 , \2924_b0 , w_4846 );
not ( w_4846 , w_4847 );
and ( w_4847 , \2918_b1 , \2918_b0 );
buf ( \2926_SUM[15]_b1 , \2925_b1 );
buf ( \2926_SUM[15]_b0 , \2925_b0 );
buf ( \2927_A[15]_b1 , \2926_SUM[15]_b1 );
buf ( \2927_A[15]_b0 , \2926_SUM[15]_b0 );
or ( \2928_b1 , \2832_A[14]_b1 , \2833_B[14]_b1 );
xor ( \2928_b0 , \2832_A[14]_b0 , w_4848 );
not ( w_4848 , w_4849 );
and ( w_4849 , \2833_B[14]_b1 , \2833_B[14]_b0 );
or ( \2929_b1 , \2928_b1 , \2915_b1 );
xor ( \2929_b0 , \2928_b0 , w_4850 );
not ( w_4850 , w_4851 );
and ( w_4851 , \2915_b1 , \2915_b0 );
buf ( \2930_SUM[14]_b1 , \2929_b1 );
buf ( \2930_SUM[14]_b0 , \2929_b0 );
buf ( \2931_A[14]_b1 , \2930_SUM[14]_b1 );
buf ( \2931_A[14]_b0 , \2930_SUM[14]_b0 );
or ( \2932_b1 , \2835_A[13]_b1 , \2836_B[13]_b1 );
xor ( \2932_b0 , \2835_A[13]_b0 , w_4852 );
not ( w_4852 , w_4853 );
and ( w_4853 , \2836_B[13]_b1 , \2836_B[13]_b0 );
or ( \2933_b1 , \2932_b1 , \2912_b1 );
xor ( \2933_b0 , \2932_b0 , w_4854 );
not ( w_4854 , w_4855 );
and ( w_4855 , \2912_b1 , \2912_b0 );
buf ( \2934_SUM[13]_b1 , \2933_b1 );
buf ( \2934_SUM[13]_b0 , \2933_b0 );
buf ( \2935_A[13]_b1 , \2934_SUM[13]_b1 );
buf ( \2935_A[13]_b0 , \2934_SUM[13]_b0 );
or ( \2936_b1 , \2838_A[12]_b1 , \2839_B[12]_b1 );
xor ( \2936_b0 , \2838_A[12]_b0 , w_4856 );
not ( w_4856 , w_4857 );
and ( w_4857 , \2839_B[12]_b1 , \2839_B[12]_b0 );
or ( \2937_b1 , \2936_b1 , \2909_b1 );
xor ( \2937_b0 , \2936_b0 , w_4858 );
not ( w_4858 , w_4859 );
and ( w_4859 , \2909_b1 , \2909_b0 );
buf ( \2938_SUM[12]_b1 , \2937_b1 );
buf ( \2938_SUM[12]_b0 , \2937_b0 );
buf ( \2939_A[12]_b1 , \2938_SUM[12]_b1 );
buf ( \2939_A[12]_b0 , \2938_SUM[12]_b0 );
or ( \2940_b1 , \2841_A[11]_b1 , \2842_B[11]_b1 );
xor ( \2940_b0 , \2841_A[11]_b0 , w_4860 );
not ( w_4860 , w_4861 );
and ( w_4861 , \2842_B[11]_b1 , \2842_B[11]_b0 );
or ( \2941_b1 , \2940_b1 , \2906_b1 );
xor ( \2941_b0 , \2940_b0 , w_4862 );
not ( w_4862 , w_4863 );
and ( w_4863 , \2906_b1 , \2906_b0 );
buf ( \2942_SUM[11]_b1 , \2941_b1 );
buf ( \2942_SUM[11]_b0 , \2941_b0 );
buf ( \2943_A[11]_b1 , \2942_SUM[11]_b1 );
buf ( \2943_A[11]_b0 , \2942_SUM[11]_b0 );
or ( \2944_b1 , \2844_A[10]_b1 , \2845_B[10]_b1 );
xor ( \2944_b0 , \2844_A[10]_b0 , w_4864 );
not ( w_4864 , w_4865 );
and ( w_4865 , \2845_B[10]_b1 , \2845_B[10]_b0 );
or ( \2945_b1 , \2944_b1 , \2903_b1 );
xor ( \2945_b0 , \2944_b0 , w_4866 );
not ( w_4866 , w_4867 );
and ( w_4867 , \2903_b1 , \2903_b0 );
buf ( \2946_SUM[10]_b1 , \2945_b1 );
buf ( \2946_SUM[10]_b0 , \2945_b0 );
buf ( \2947_A[10]_b1 , \2946_SUM[10]_b1 );
buf ( \2947_A[10]_b0 , \2946_SUM[10]_b0 );
or ( \2948_b1 , \2847_A[9]_b1 , \2848_B[9]_b1 );
xor ( \2948_b0 , \2847_A[9]_b0 , w_4868 );
not ( w_4868 , w_4869 );
and ( w_4869 , \2848_B[9]_b1 , \2848_B[9]_b0 );
or ( \2949_b1 , \2948_b1 , \2900_b1 );
xor ( \2949_b0 , \2948_b0 , w_4870 );
not ( w_4870 , w_4871 );
and ( w_4871 , \2900_b1 , \2900_b0 );
buf ( \2950_SUM[9]_b1 , \2949_b1 );
buf ( \2950_SUM[9]_b0 , \2949_b0 );
buf ( \2951_A[9]_b1 , \2950_SUM[9]_b1 );
buf ( \2951_A[9]_b0 , \2950_SUM[9]_b0 );
or ( \2952_b1 , \2850_A[8]_b1 , \2851_B[8]_b1 );
xor ( \2952_b0 , \2850_A[8]_b0 , w_4872 );
not ( w_4872 , w_4873 );
and ( w_4873 , \2851_B[8]_b1 , \2851_B[8]_b0 );
or ( \2953_b1 , \2952_b1 , \2897_b1 );
xor ( \2953_b0 , \2952_b0 , w_4874 );
not ( w_4874 , w_4875 );
and ( w_4875 , \2897_b1 , \2897_b0 );
buf ( \2954_SUM[8]_b1 , \2953_b1 );
buf ( \2954_SUM[8]_b0 , \2953_b0 );
buf ( \2955_A[8]_b1 , \2954_SUM[8]_b1 );
buf ( \2955_A[8]_b0 , \2954_SUM[8]_b0 );
or ( \2956_b1 , \2853_A[7]_b1 , \2854_B[7]_b1 );
xor ( \2956_b0 , \2853_A[7]_b0 , w_4876 );
not ( w_4876 , w_4877 );
and ( w_4877 , \2854_B[7]_b1 , \2854_B[7]_b0 );
or ( \2957_b1 , \2956_b1 , \2894_b1 );
xor ( \2957_b0 , \2956_b0 , w_4878 );
not ( w_4878 , w_4879 );
and ( w_4879 , \2894_b1 , \2894_b0 );
buf ( \2958_SUM[7]_b1 , \2957_b1 );
buf ( \2958_SUM[7]_b0 , \2957_b0 );
buf ( \2959_A[7]_b1 , \2958_SUM[7]_b1 );
buf ( \2959_A[7]_b0 , \2958_SUM[7]_b0 );
or ( \2960_b1 , \2856_A[6]_b1 , \2857_B[6]_b1 );
xor ( \2960_b0 , \2856_A[6]_b0 , w_4880 );
not ( w_4880 , w_4881 );
and ( w_4881 , \2857_B[6]_b1 , \2857_B[6]_b0 );
or ( \2961_b1 , \2960_b1 , \2891_b1 );
xor ( \2961_b0 , \2960_b0 , w_4882 );
not ( w_4882 , w_4883 );
and ( w_4883 , \2891_b1 , \2891_b0 );
buf ( \2962_SUM[6]_b1 , \2961_b1 );
buf ( \2962_SUM[6]_b0 , \2961_b0 );
buf ( \2963_A[6]_b1 , \2962_SUM[6]_b1 );
buf ( \2963_A[6]_b0 , \2962_SUM[6]_b0 );
or ( \2964_b1 , \2859_A[5]_b1 , \2860_B[5]_b1 );
xor ( \2964_b0 , \2859_A[5]_b0 , w_4884 );
not ( w_4884 , w_4885 );
and ( w_4885 , \2860_B[5]_b1 , \2860_B[5]_b0 );
or ( \2965_b1 , \2964_b1 , \2888_b1 );
xor ( \2965_b0 , \2964_b0 , w_4886 );
not ( w_4886 , w_4887 );
and ( w_4887 , \2888_b1 , \2888_b0 );
buf ( \2966_SUM[5]_b1 , \2965_b1 );
buf ( \2966_SUM[5]_b0 , \2965_b0 );
buf ( \2967_A[5]_b1 , \2966_SUM[5]_b1 );
buf ( \2967_A[5]_b0 , \2966_SUM[5]_b0 );
or ( \2968_b1 , \2862_A[4]_b1 , \2863_B[4]_b1 );
xor ( \2968_b0 , \2862_A[4]_b0 , w_4888 );
not ( w_4888 , w_4889 );
and ( w_4889 , \2863_B[4]_b1 , \2863_B[4]_b0 );
or ( \2969_b1 , \2968_b1 , \2885_b1 );
xor ( \2969_b0 , \2968_b0 , w_4890 );
not ( w_4890 , w_4891 );
and ( w_4891 , \2885_b1 , \2885_b0 );
buf ( \2970_SUM[4]_b1 , \2969_b1 );
buf ( \2970_SUM[4]_b0 , \2969_b0 );
buf ( \2971_A[4]_b1 , \2970_SUM[4]_b1 );
buf ( \2971_A[4]_b0 , \2970_SUM[4]_b0 );
or ( \2972_b1 , \2865_A[3]_b1 , \2866_B[3]_b1 );
xor ( \2972_b0 , \2865_A[3]_b0 , w_4892 );
not ( w_4892 , w_4893 );
and ( w_4893 , \2866_B[3]_b1 , \2866_B[3]_b0 );
or ( \2973_b1 , \2972_b1 , \2882_b1 );
xor ( \2973_b0 , \2972_b0 , w_4894 );
not ( w_4894 , w_4895 );
and ( w_4895 , \2882_b1 , \2882_b0 );
buf ( \2974_SUM[3]_b1 , \2973_b1 );
buf ( \2974_SUM[3]_b0 , \2973_b0 );
buf ( \2975_A[3]_b1 , \2974_SUM[3]_b1 );
buf ( \2975_A[3]_b0 , \2974_SUM[3]_b0 );
or ( \2976_b1 , \2868_A[2]_b1 , \2869_B[2]_b1 );
xor ( \2976_b0 , \2868_A[2]_b0 , w_4896 );
not ( w_4896 , w_4897 );
and ( w_4897 , \2869_B[2]_b1 , \2869_B[2]_b0 );
or ( \2977_b1 , \2976_b1 , \2879_b1 );
xor ( \2977_b0 , \2976_b0 , w_4898 );
not ( w_4898 , w_4899 );
and ( w_4899 , \2879_b1 , \2879_b0 );
buf ( \2978_SUM[2]_b1 , \2977_b1 );
buf ( \2978_SUM[2]_b0 , \2977_b0 );
buf ( \2979_A[2]_b1 , \2978_SUM[2]_b1 );
buf ( \2979_A[2]_b0 , \2978_SUM[2]_b0 );
or ( \2980_b1 , \2871_A[1]_b1 , \2872_B[1]_b1 );
xor ( \2980_b0 , \2871_A[1]_b0 , w_4900 );
not ( w_4900 , w_4901 );
and ( w_4901 , \2872_B[1]_b1 , \2872_B[1]_b0 );
or ( \2981_b1 , \2980_b1 , \2876_b1 );
xor ( \2981_b0 , \2980_b0 , w_4902 );
not ( w_4902 , w_4903 );
and ( w_4903 , \2876_b1 , \2876_b0 );
buf ( \2982_SUM[1]_b1 , \2981_b1 );
buf ( \2982_SUM[1]_b0 , \2981_b0 );
buf ( \2983_A[1]_b1 , \2982_SUM[1]_b1 );
buf ( \2983_A[1]_b0 , \2982_SUM[1]_b0 );
or ( \2984_b1 , \2874_A[0]_b1 , \2875_B[0]_b1 );
xor ( \2984_b0 , \2874_A[0]_b0 , w_4904 );
not ( w_4904 , w_4905 );
and ( w_4905 , \2875_B[0]_b1 , \2875_B[0]_b0 );
buf ( \2985_SUM[0]_b1 , \2984_b1 );
buf ( \2985_SUM[0]_b0 , \2984_b0 );
buf ( \2986_A[0]_b1 , \2985_SUM[0]_b1 );
buf ( \2986_A[0]_b0 , \2985_SUM[0]_b0 );
buf ( \2987_B[15]_b1 , \2828_b1 );
buf ( \2987_B[15]_b0 , \2828_b0 );
buf ( \2988_B[14]_b1 , \2616_b1 );
buf ( \2988_B[14]_b0 , \2616_b0 );
buf ( \2989_B[13]_b1 , \2416_b1 );
buf ( \2989_B[13]_b0 , \2416_b0 );
buf ( \2990_B[12]_b1 , \2228_b1 );
buf ( \2990_B[12]_b0 , \2228_b0 );
buf ( \2991_B[11]_b1 , \2052_b1 );
buf ( \2991_B[11]_b0 , \2052_b0 );
buf ( \2992_B[10]_b1 , \1888_b1 );
buf ( \2992_B[10]_b0 , \1888_b0 );
buf ( \2993_B[9]_b1 , \1736_b1 );
buf ( \2993_B[9]_b0 , \1736_b0 );
buf ( \2994_B[8]_b1 , \1596_b1 );
buf ( \2994_B[8]_b0 , \1596_b0 );
buf ( \2995_B[7]_b1 , \1468_b1 );
buf ( \2995_B[7]_b0 , \1468_b0 );
buf ( \2996_B[6]_b1 , \1352_b1 );
buf ( \2996_B[6]_b0 , \1352_b0 );
buf ( \2997_B[5]_b1 , \1248_b1 );
buf ( \2997_B[5]_b0 , \1248_b0 );
buf ( \2998_B[4]_b1 , \1156_b1 );
buf ( \2998_B[4]_b0 , \1156_b0 );
buf ( \2999_B[3]_b1 , \1076_b1 );
buf ( \2999_B[3]_b0 , \1076_b0 );
buf ( \3000_B[2]_b1 , \1008_b1 );
buf ( \3000_B[2]_b0 , \1008_b0 );
buf ( \3001_B[1]_b1 , \952_b1 );
buf ( \3001_B[1]_b0 , \952_b0 );
buf ( \3002_B[0]_b1 , \910_b1 );
buf ( \3002_B[0]_b0 , \910_b0 );
or ( \3003_b1 , \2923_A[16]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4906 );
and ( \3003_b0 , \2923_A[16]_b0 , w_4907 );
and ( w_4906 , w_4907 , \3001_B[1]_b0 );
or ( \3004_b1 , \2923_A[16]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4908 );
and ( \3004_b0 , \2923_A[16]_b0 , w_4909 );
and ( w_4908 , w_4909 , \3002_B[0]_b0 );
or ( \3005_b1 , \2927_A[15]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4910 );
and ( \3005_b0 , \2927_A[15]_b0 , w_4911 );
and ( w_4910 , w_4911 , \3001_B[1]_b0 );
or ( \3006_b1 , \3004_b1 , \3005_b1 );
not ( \3005_b1 , w_4912 );
and ( \3006_b0 , \3004_b0 , w_4913 );
and ( w_4912 , w_4913 , \3005_b0 );
or ( \3007_b1 , \3004_b1 , \3005_b1 );
xor ( \3007_b0 , \3004_b0 , w_4914 );
not ( w_4914 , w_4915 );
and ( w_4915 , \3005_b1 , \3005_b0 );
or ( \3008_b1 , \2927_A[15]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4916 );
and ( \3008_b0 , \2927_A[15]_b0 , w_4917 );
and ( w_4916 , w_4917 , \3002_B[0]_b0 );
or ( \3009_b1 , \2931_A[14]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4918 );
and ( \3009_b0 , \2931_A[14]_b0 , w_4919 );
and ( w_4918 , w_4919 , \3001_B[1]_b0 );
or ( \3010_b1 , \3008_b1 , \3009_b1 );
not ( \3009_b1 , w_4920 );
and ( \3010_b0 , \3008_b0 , w_4921 );
and ( w_4920 , w_4921 , \3009_b0 );
or ( \3011_b1 , \3008_b1 , \3009_b1 );
xor ( \3011_b0 , \3008_b0 , w_4922 );
not ( w_4922 , w_4923 );
and ( w_4923 , \3009_b1 , \3009_b0 );
or ( \3012_b1 , \2931_A[14]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4924 );
and ( \3012_b0 , \2931_A[14]_b0 , w_4925 );
and ( w_4924 , w_4925 , \3002_B[0]_b0 );
or ( \3013_b1 , \2935_A[13]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4926 );
and ( \3013_b0 , \2935_A[13]_b0 , w_4927 );
and ( w_4926 , w_4927 , \3001_B[1]_b0 );
or ( \3014_b1 , \3012_b1 , \3013_b1 );
not ( \3013_b1 , w_4928 );
and ( \3014_b0 , \3012_b0 , w_4929 );
and ( w_4928 , w_4929 , \3013_b0 );
or ( \3015_b1 , \3012_b1 , \3013_b1 );
xor ( \3015_b0 , \3012_b0 , w_4930 );
not ( w_4930 , w_4931 );
and ( w_4931 , \3013_b1 , \3013_b0 );
or ( \3016_b1 , \2935_A[13]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4932 );
and ( \3016_b0 , \2935_A[13]_b0 , w_4933 );
and ( w_4932 , w_4933 , \3002_B[0]_b0 );
or ( \3017_b1 , \2939_A[12]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4934 );
and ( \3017_b0 , \2939_A[12]_b0 , w_4935 );
and ( w_4934 , w_4935 , \3001_B[1]_b0 );
or ( \3018_b1 , \3016_b1 , \3017_b1 );
not ( \3017_b1 , w_4936 );
and ( \3018_b0 , \3016_b0 , w_4937 );
and ( w_4936 , w_4937 , \3017_b0 );
or ( \3019_b1 , \3016_b1 , \3017_b1 );
xor ( \3019_b0 , \3016_b0 , w_4938 );
not ( w_4938 , w_4939 );
and ( w_4939 , \3017_b1 , \3017_b0 );
or ( \3020_b1 , \2939_A[12]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4940 );
and ( \3020_b0 , \2939_A[12]_b0 , w_4941 );
and ( w_4940 , w_4941 , \3002_B[0]_b0 );
or ( \3021_b1 , \2943_A[11]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4942 );
and ( \3021_b0 , \2943_A[11]_b0 , w_4943 );
and ( w_4942 , w_4943 , \3001_B[1]_b0 );
or ( \3022_b1 , \3020_b1 , \3021_b1 );
not ( \3021_b1 , w_4944 );
and ( \3022_b0 , \3020_b0 , w_4945 );
and ( w_4944 , w_4945 , \3021_b0 );
or ( \3023_b1 , \3020_b1 , \3021_b1 );
xor ( \3023_b0 , \3020_b0 , w_4946 );
not ( w_4946 , w_4947 );
and ( w_4947 , \3021_b1 , \3021_b0 );
or ( \3024_b1 , \2943_A[11]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4948 );
and ( \3024_b0 , \2943_A[11]_b0 , w_4949 );
and ( w_4948 , w_4949 , \3002_B[0]_b0 );
or ( \3025_b1 , \2947_A[10]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4950 );
and ( \3025_b0 , \2947_A[10]_b0 , w_4951 );
and ( w_4950 , w_4951 , \3001_B[1]_b0 );
or ( \3026_b1 , \3024_b1 , \3025_b1 );
not ( \3025_b1 , w_4952 );
and ( \3026_b0 , \3024_b0 , w_4953 );
and ( w_4952 , w_4953 , \3025_b0 );
or ( \3027_b1 , \3024_b1 , \3025_b1 );
xor ( \3027_b0 , \3024_b0 , w_4954 );
not ( w_4954 , w_4955 );
and ( w_4955 , \3025_b1 , \3025_b0 );
or ( \3028_b1 , \2947_A[10]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4956 );
and ( \3028_b0 , \2947_A[10]_b0 , w_4957 );
and ( w_4956 , w_4957 , \3002_B[0]_b0 );
or ( \3029_b1 , \2951_A[9]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4958 );
and ( \3029_b0 , \2951_A[9]_b0 , w_4959 );
and ( w_4958 , w_4959 , \3001_B[1]_b0 );
or ( \3030_b1 , \3028_b1 , \3029_b1 );
not ( \3029_b1 , w_4960 );
and ( \3030_b0 , \3028_b0 , w_4961 );
and ( w_4960 , w_4961 , \3029_b0 );
or ( \3031_b1 , \3028_b1 , \3029_b1 );
xor ( \3031_b0 , \3028_b0 , w_4962 );
not ( w_4962 , w_4963 );
and ( w_4963 , \3029_b1 , \3029_b0 );
or ( \3032_b1 , \2951_A[9]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4964 );
and ( \3032_b0 , \2951_A[9]_b0 , w_4965 );
and ( w_4964 , w_4965 , \3002_B[0]_b0 );
or ( \3033_b1 , \2955_A[8]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4966 );
and ( \3033_b0 , \2955_A[8]_b0 , w_4967 );
and ( w_4966 , w_4967 , \3001_B[1]_b0 );
or ( \3034_b1 , \3032_b1 , \3033_b1 );
not ( \3033_b1 , w_4968 );
and ( \3034_b0 , \3032_b0 , w_4969 );
and ( w_4968 , w_4969 , \3033_b0 );
or ( \3035_b1 , \3032_b1 , \3033_b1 );
xor ( \3035_b0 , \3032_b0 , w_4970 );
not ( w_4970 , w_4971 );
and ( w_4971 , \3033_b1 , \3033_b0 );
or ( \3036_b1 , \2955_A[8]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4972 );
and ( \3036_b0 , \2955_A[8]_b0 , w_4973 );
and ( w_4972 , w_4973 , \3002_B[0]_b0 );
or ( \3037_b1 , \2959_A[7]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4974 );
and ( \3037_b0 , \2959_A[7]_b0 , w_4975 );
and ( w_4974 , w_4975 , \3001_B[1]_b0 );
or ( \3038_b1 , \3036_b1 , \3037_b1 );
not ( \3037_b1 , w_4976 );
and ( \3038_b0 , \3036_b0 , w_4977 );
and ( w_4976 , w_4977 , \3037_b0 );
or ( \3039_b1 , \3036_b1 , \3037_b1 );
xor ( \3039_b0 , \3036_b0 , w_4978 );
not ( w_4978 , w_4979 );
and ( w_4979 , \3037_b1 , \3037_b0 );
or ( \3040_b1 , \2959_A[7]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4980 );
and ( \3040_b0 , \2959_A[7]_b0 , w_4981 );
and ( w_4980 , w_4981 , \3002_B[0]_b0 );
or ( \3041_b1 , \2963_A[6]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4982 );
and ( \3041_b0 , \2963_A[6]_b0 , w_4983 );
and ( w_4982 , w_4983 , \3001_B[1]_b0 );
or ( \3042_b1 , \3040_b1 , \3041_b1 );
not ( \3041_b1 , w_4984 );
and ( \3042_b0 , \3040_b0 , w_4985 );
and ( w_4984 , w_4985 , \3041_b0 );
or ( \3043_b1 , \3040_b1 , \3041_b1 );
xor ( \3043_b0 , \3040_b0 , w_4986 );
not ( w_4986 , w_4987 );
and ( w_4987 , \3041_b1 , \3041_b0 );
or ( \3044_b1 , \2963_A[6]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4988 );
and ( \3044_b0 , \2963_A[6]_b0 , w_4989 );
and ( w_4988 , w_4989 , \3002_B[0]_b0 );
or ( \3045_b1 , \2967_A[5]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4990 );
and ( \3045_b0 , \2967_A[5]_b0 , w_4991 );
and ( w_4990 , w_4991 , \3001_B[1]_b0 );
or ( \3046_b1 , \3044_b1 , \3045_b1 );
not ( \3045_b1 , w_4992 );
and ( \3046_b0 , \3044_b0 , w_4993 );
and ( w_4992 , w_4993 , \3045_b0 );
or ( \3047_b1 , \3044_b1 , \3045_b1 );
xor ( \3047_b0 , \3044_b0 , w_4994 );
not ( w_4994 , w_4995 );
and ( w_4995 , \3045_b1 , \3045_b0 );
or ( \3048_b1 , \2967_A[5]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_4996 );
and ( \3048_b0 , \2967_A[5]_b0 , w_4997 );
and ( w_4996 , w_4997 , \3002_B[0]_b0 );
or ( \3049_b1 , \2971_A[4]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_4998 );
and ( \3049_b0 , \2971_A[4]_b0 , w_4999 );
and ( w_4998 , w_4999 , \3001_B[1]_b0 );
or ( \3050_b1 , \3048_b1 , \3049_b1 );
not ( \3049_b1 , w_5000 );
and ( \3050_b0 , \3048_b0 , w_5001 );
and ( w_5000 , w_5001 , \3049_b0 );
or ( \3051_b1 , \3048_b1 , \3049_b1 );
xor ( \3051_b0 , \3048_b0 , w_5002 );
not ( w_5002 , w_5003 );
and ( w_5003 , \3049_b1 , \3049_b0 );
or ( \3052_b1 , \2971_A[4]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_5004 );
and ( \3052_b0 , \2971_A[4]_b0 , w_5005 );
and ( w_5004 , w_5005 , \3002_B[0]_b0 );
or ( \3053_b1 , \2975_A[3]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_5006 );
and ( \3053_b0 , \2975_A[3]_b0 , w_5007 );
and ( w_5006 , w_5007 , \3001_B[1]_b0 );
or ( \3054_b1 , \3052_b1 , \3053_b1 );
not ( \3053_b1 , w_5008 );
and ( \3054_b0 , \3052_b0 , w_5009 );
and ( w_5008 , w_5009 , \3053_b0 );
or ( \3055_b1 , \3052_b1 , \3053_b1 );
xor ( \3055_b0 , \3052_b0 , w_5010 );
not ( w_5010 , w_5011 );
and ( w_5011 , \3053_b1 , \3053_b0 );
or ( \3056_b1 , \2975_A[3]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_5012 );
and ( \3056_b0 , \2975_A[3]_b0 , w_5013 );
and ( w_5012 , w_5013 , \3002_B[0]_b0 );
or ( \3057_b1 , \2979_A[2]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_5014 );
and ( \3057_b0 , \2979_A[2]_b0 , w_5015 );
and ( w_5014 , w_5015 , \3001_B[1]_b0 );
or ( \3058_b1 , \3056_b1 , \3057_b1 );
not ( \3057_b1 , w_5016 );
and ( \3058_b0 , \3056_b0 , w_5017 );
and ( w_5016 , w_5017 , \3057_b0 );
or ( \3059_b1 , \3056_b1 , \3057_b1 );
xor ( \3059_b0 , \3056_b0 , w_5018 );
not ( w_5018 , w_5019 );
and ( w_5019 , \3057_b1 , \3057_b0 );
or ( \3060_b1 , \2979_A[2]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_5020 );
and ( \3060_b0 , \2979_A[2]_b0 , w_5021 );
and ( w_5020 , w_5021 , \3002_B[0]_b0 );
or ( \3061_b1 , \2983_A[1]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_5022 );
and ( \3061_b0 , \2983_A[1]_b0 , w_5023 );
and ( w_5022 , w_5023 , \3001_B[1]_b0 );
or ( \3062_b1 , \3060_b1 , \3061_b1 );
not ( \3061_b1 , w_5024 );
and ( \3062_b0 , \3060_b0 , w_5025 );
and ( w_5024 , w_5025 , \3061_b0 );
or ( \3063_b1 , \3060_b1 , \3061_b1 );
xor ( \3063_b0 , \3060_b0 , w_5026 );
not ( w_5026 , w_5027 );
and ( w_5027 , \3061_b1 , \3061_b0 );
or ( \3064_b1 , \2983_A[1]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_5028 );
and ( \3064_b0 , \2983_A[1]_b0 , w_5029 );
and ( w_5028 , w_5029 , \3002_B[0]_b0 );
or ( \3065_b1 , \2986_A[0]_b1 , \3001_B[1]_b1 );
not ( \3001_B[1]_b1 , w_5030 );
and ( \3065_b0 , \2986_A[0]_b0 , w_5031 );
and ( w_5030 , w_5031 , \3001_B[1]_b0 );
or ( \3066_b1 , \3064_b1 , \3065_b1 );
not ( \3065_b1 , w_5032 );
and ( \3066_b0 , \3064_b0 , w_5033 );
and ( w_5032 , w_5033 , \3065_b0 );
or ( \3067_b1 , \3063_b1 , \3066_b1 );
not ( \3066_b1 , w_5034 );
and ( \3067_b0 , \3063_b0 , w_5035 );
and ( w_5034 , w_5035 , \3066_b0 );
or ( \3068_b1 , \3062_b1 , w_5036 );
or ( \3068_b0 , \3062_b0 , \3067_b0 );
not ( \3067_b0 , w_5037 );
and ( w_5037 , w_5036 , \3067_b1 );
or ( \3069_b1 , \3059_b1 , \3068_b1 );
not ( \3068_b1 , w_5038 );
and ( \3069_b0 , \3059_b0 , w_5039 );
and ( w_5038 , w_5039 , \3068_b0 );
or ( \3070_b1 , \3058_b1 , w_5040 );
or ( \3070_b0 , \3058_b0 , \3069_b0 );
not ( \3069_b0 , w_5041 );
and ( w_5041 , w_5040 , \3069_b1 );
or ( \3071_b1 , \3055_b1 , \3070_b1 );
not ( \3070_b1 , w_5042 );
and ( \3071_b0 , \3055_b0 , w_5043 );
and ( w_5042 , w_5043 , \3070_b0 );
or ( \3072_b1 , \3054_b1 , w_5044 );
or ( \3072_b0 , \3054_b0 , \3071_b0 );
not ( \3071_b0 , w_5045 );
and ( w_5045 , w_5044 , \3071_b1 );
or ( \3073_b1 , \3051_b1 , \3072_b1 );
not ( \3072_b1 , w_5046 );
and ( \3073_b0 , \3051_b0 , w_5047 );
and ( w_5046 , w_5047 , \3072_b0 );
or ( \3074_b1 , \3050_b1 , w_5048 );
or ( \3074_b0 , \3050_b0 , \3073_b0 );
not ( \3073_b0 , w_5049 );
and ( w_5049 , w_5048 , \3073_b1 );
or ( \3075_b1 , \3047_b1 , \3074_b1 );
not ( \3074_b1 , w_5050 );
and ( \3075_b0 , \3047_b0 , w_5051 );
and ( w_5050 , w_5051 , \3074_b0 );
or ( \3076_b1 , \3046_b1 , w_5052 );
or ( \3076_b0 , \3046_b0 , \3075_b0 );
not ( \3075_b0 , w_5053 );
and ( w_5053 , w_5052 , \3075_b1 );
or ( \3077_b1 , \3043_b1 , \3076_b1 );
not ( \3076_b1 , w_5054 );
and ( \3077_b0 , \3043_b0 , w_5055 );
and ( w_5054 , w_5055 , \3076_b0 );
or ( \3078_b1 , \3042_b1 , w_5056 );
or ( \3078_b0 , \3042_b0 , \3077_b0 );
not ( \3077_b0 , w_5057 );
and ( w_5057 , w_5056 , \3077_b1 );
or ( \3079_b1 , \3039_b1 , \3078_b1 );
not ( \3078_b1 , w_5058 );
and ( \3079_b0 , \3039_b0 , w_5059 );
and ( w_5058 , w_5059 , \3078_b0 );
or ( \3080_b1 , \3038_b1 , w_5060 );
or ( \3080_b0 , \3038_b0 , \3079_b0 );
not ( \3079_b0 , w_5061 );
and ( w_5061 , w_5060 , \3079_b1 );
or ( \3081_b1 , \3035_b1 , \3080_b1 );
not ( \3080_b1 , w_5062 );
and ( \3081_b0 , \3035_b0 , w_5063 );
and ( w_5062 , w_5063 , \3080_b0 );
or ( \3082_b1 , \3034_b1 , w_5064 );
or ( \3082_b0 , \3034_b0 , \3081_b0 );
not ( \3081_b0 , w_5065 );
and ( w_5065 , w_5064 , \3081_b1 );
or ( \3083_b1 , \3031_b1 , \3082_b1 );
not ( \3082_b1 , w_5066 );
and ( \3083_b0 , \3031_b0 , w_5067 );
and ( w_5066 , w_5067 , \3082_b0 );
or ( \3084_b1 , \3030_b1 , w_5068 );
or ( \3084_b0 , \3030_b0 , \3083_b0 );
not ( \3083_b0 , w_5069 );
and ( w_5069 , w_5068 , \3083_b1 );
or ( \3085_b1 , \3027_b1 , \3084_b1 );
not ( \3084_b1 , w_5070 );
and ( \3085_b0 , \3027_b0 , w_5071 );
and ( w_5070 , w_5071 , \3084_b0 );
or ( \3086_b1 , \3026_b1 , w_5072 );
or ( \3086_b0 , \3026_b0 , \3085_b0 );
not ( \3085_b0 , w_5073 );
and ( w_5073 , w_5072 , \3085_b1 );
or ( \3087_b1 , \3023_b1 , \3086_b1 );
not ( \3086_b1 , w_5074 );
and ( \3087_b0 , \3023_b0 , w_5075 );
and ( w_5074 , w_5075 , \3086_b0 );
or ( \3088_b1 , \3022_b1 , w_5076 );
or ( \3088_b0 , \3022_b0 , \3087_b0 );
not ( \3087_b0 , w_5077 );
and ( w_5077 , w_5076 , \3087_b1 );
or ( \3089_b1 , \3019_b1 , \3088_b1 );
not ( \3088_b1 , w_5078 );
and ( \3089_b0 , \3019_b0 , w_5079 );
and ( w_5078 , w_5079 , \3088_b0 );
or ( \3090_b1 , \3018_b1 , w_5080 );
or ( \3090_b0 , \3018_b0 , \3089_b0 );
not ( \3089_b0 , w_5081 );
and ( w_5081 , w_5080 , \3089_b1 );
or ( \3091_b1 , \3015_b1 , \3090_b1 );
not ( \3090_b1 , w_5082 );
and ( \3091_b0 , \3015_b0 , w_5083 );
and ( w_5082 , w_5083 , \3090_b0 );
or ( \3092_b1 , \3014_b1 , w_5084 );
or ( \3092_b0 , \3014_b0 , \3091_b0 );
not ( \3091_b0 , w_5085 );
and ( w_5085 , w_5084 , \3091_b1 );
or ( \3093_b1 , \3011_b1 , \3092_b1 );
not ( \3092_b1 , w_5086 );
and ( \3093_b0 , \3011_b0 , w_5087 );
and ( w_5086 , w_5087 , \3092_b0 );
or ( \3094_b1 , \3010_b1 , w_5088 );
or ( \3094_b0 , \3010_b0 , \3093_b0 );
not ( \3093_b0 , w_5089 );
and ( w_5089 , w_5088 , \3093_b1 );
or ( \3095_b1 , \3007_b1 , \3094_b1 );
not ( \3094_b1 , w_5090 );
and ( \3095_b0 , \3007_b0 , w_5091 );
and ( w_5090 , w_5091 , \3094_b0 );
or ( \3096_b1 , \3006_b1 , w_5092 );
or ( \3096_b0 , \3006_b0 , \3095_b0 );
not ( \3095_b0 , w_5093 );
and ( w_5093 , w_5092 , \3095_b1 );
or ( \3097_b1 , \3003_b1 , \3096_b1 );
not ( \3096_b1 , w_5094 );
and ( \3097_b0 , \3003_b0 , w_5095 );
and ( w_5094 , w_5095 , \3096_b0 );
or ( \3098_b1 , \2923_A[16]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5096 );
and ( \3098_b0 , \2923_A[16]_b0 , w_5097 );
and ( w_5096 , w_5097 , \3000_B[2]_b0 );
or ( \3099_b1 , \3097_b1 , \3098_b1 );
not ( \3098_b1 , w_5098 );
and ( \3099_b0 , \3097_b0 , w_5099 );
and ( w_5098 , w_5099 , \3098_b0 );
or ( \3100_b1 , \3097_b1 , \3098_b1 );
xor ( \3100_b0 , \3097_b0 , w_5100 );
not ( w_5100 , w_5101 );
and ( w_5101 , \3098_b1 , \3098_b0 );
or ( \3101_b1 , \3003_b1 , \3096_b1 );
xor ( \3101_b0 , \3003_b0 , w_5102 );
not ( w_5102 , w_5103 );
and ( w_5103 , \3096_b1 , \3096_b0 );
or ( \3102_b1 , \2927_A[15]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5104 );
and ( \3102_b0 , \2927_A[15]_b0 , w_5105 );
and ( w_5104 , w_5105 , \3000_B[2]_b0 );
or ( \3103_b1 , \3101_b1 , \3102_b1 );
not ( \3102_b1 , w_5106 );
and ( \3103_b0 , \3101_b0 , w_5107 );
and ( w_5106 , w_5107 , \3102_b0 );
or ( \3104_b1 , \3101_b1 , \3102_b1 );
xor ( \3104_b0 , \3101_b0 , w_5108 );
not ( w_5108 , w_5109 );
and ( w_5109 , \3102_b1 , \3102_b0 );
or ( \3105_b1 , \3007_b1 , \3094_b1 );
xor ( \3105_b0 , \3007_b0 , w_5110 );
not ( w_5110 , w_5111 );
and ( w_5111 , \3094_b1 , \3094_b0 );
or ( \3106_b1 , \2931_A[14]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5112 );
and ( \3106_b0 , \2931_A[14]_b0 , w_5113 );
and ( w_5112 , w_5113 , \3000_B[2]_b0 );
or ( \3107_b1 , \3105_b1 , \3106_b1 );
not ( \3106_b1 , w_5114 );
and ( \3107_b0 , \3105_b0 , w_5115 );
and ( w_5114 , w_5115 , \3106_b0 );
or ( \3108_b1 , \3105_b1 , \3106_b1 );
xor ( \3108_b0 , \3105_b0 , w_5116 );
not ( w_5116 , w_5117 );
and ( w_5117 , \3106_b1 , \3106_b0 );
or ( \3109_b1 , \3011_b1 , \3092_b1 );
xor ( \3109_b0 , \3011_b0 , w_5118 );
not ( w_5118 , w_5119 );
and ( w_5119 , \3092_b1 , \3092_b0 );
or ( \3110_b1 , \2935_A[13]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5120 );
and ( \3110_b0 , \2935_A[13]_b0 , w_5121 );
and ( w_5120 , w_5121 , \3000_B[2]_b0 );
or ( \3111_b1 , \3109_b1 , \3110_b1 );
not ( \3110_b1 , w_5122 );
and ( \3111_b0 , \3109_b0 , w_5123 );
and ( w_5122 , w_5123 , \3110_b0 );
or ( \3112_b1 , \3109_b1 , \3110_b1 );
xor ( \3112_b0 , \3109_b0 , w_5124 );
not ( w_5124 , w_5125 );
and ( w_5125 , \3110_b1 , \3110_b0 );
or ( \3113_b1 , \3015_b1 , \3090_b1 );
xor ( \3113_b0 , \3015_b0 , w_5126 );
not ( w_5126 , w_5127 );
and ( w_5127 , \3090_b1 , \3090_b0 );
or ( \3114_b1 , \2939_A[12]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5128 );
and ( \3114_b0 , \2939_A[12]_b0 , w_5129 );
and ( w_5128 , w_5129 , \3000_B[2]_b0 );
or ( \3115_b1 , \3113_b1 , \3114_b1 );
not ( \3114_b1 , w_5130 );
and ( \3115_b0 , \3113_b0 , w_5131 );
and ( w_5130 , w_5131 , \3114_b0 );
or ( \3116_b1 , \3113_b1 , \3114_b1 );
xor ( \3116_b0 , \3113_b0 , w_5132 );
not ( w_5132 , w_5133 );
and ( w_5133 , \3114_b1 , \3114_b0 );
or ( \3117_b1 , \3019_b1 , \3088_b1 );
xor ( \3117_b0 , \3019_b0 , w_5134 );
not ( w_5134 , w_5135 );
and ( w_5135 , \3088_b1 , \3088_b0 );
or ( \3118_b1 , \2943_A[11]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5136 );
and ( \3118_b0 , \2943_A[11]_b0 , w_5137 );
and ( w_5136 , w_5137 , \3000_B[2]_b0 );
or ( \3119_b1 , \3117_b1 , \3118_b1 );
not ( \3118_b1 , w_5138 );
and ( \3119_b0 , \3117_b0 , w_5139 );
and ( w_5138 , w_5139 , \3118_b0 );
or ( \3120_b1 , \3117_b1 , \3118_b1 );
xor ( \3120_b0 , \3117_b0 , w_5140 );
not ( w_5140 , w_5141 );
and ( w_5141 , \3118_b1 , \3118_b0 );
or ( \3121_b1 , \3023_b1 , \3086_b1 );
xor ( \3121_b0 , \3023_b0 , w_5142 );
not ( w_5142 , w_5143 );
and ( w_5143 , \3086_b1 , \3086_b0 );
or ( \3122_b1 , \2947_A[10]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5144 );
and ( \3122_b0 , \2947_A[10]_b0 , w_5145 );
and ( w_5144 , w_5145 , \3000_B[2]_b0 );
or ( \3123_b1 , \3121_b1 , \3122_b1 );
not ( \3122_b1 , w_5146 );
and ( \3123_b0 , \3121_b0 , w_5147 );
and ( w_5146 , w_5147 , \3122_b0 );
or ( \3124_b1 , \3121_b1 , \3122_b1 );
xor ( \3124_b0 , \3121_b0 , w_5148 );
not ( w_5148 , w_5149 );
and ( w_5149 , \3122_b1 , \3122_b0 );
or ( \3125_b1 , \3027_b1 , \3084_b1 );
xor ( \3125_b0 , \3027_b0 , w_5150 );
not ( w_5150 , w_5151 );
and ( w_5151 , \3084_b1 , \3084_b0 );
or ( \3126_b1 , \2951_A[9]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5152 );
and ( \3126_b0 , \2951_A[9]_b0 , w_5153 );
and ( w_5152 , w_5153 , \3000_B[2]_b0 );
or ( \3127_b1 , \3125_b1 , \3126_b1 );
not ( \3126_b1 , w_5154 );
and ( \3127_b0 , \3125_b0 , w_5155 );
and ( w_5154 , w_5155 , \3126_b0 );
or ( \3128_b1 , \3125_b1 , \3126_b1 );
xor ( \3128_b0 , \3125_b0 , w_5156 );
not ( w_5156 , w_5157 );
and ( w_5157 , \3126_b1 , \3126_b0 );
or ( \3129_b1 , \3031_b1 , \3082_b1 );
xor ( \3129_b0 , \3031_b0 , w_5158 );
not ( w_5158 , w_5159 );
and ( w_5159 , \3082_b1 , \3082_b0 );
or ( \3130_b1 , \2955_A[8]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5160 );
and ( \3130_b0 , \2955_A[8]_b0 , w_5161 );
and ( w_5160 , w_5161 , \3000_B[2]_b0 );
or ( \3131_b1 , \3129_b1 , \3130_b1 );
not ( \3130_b1 , w_5162 );
and ( \3131_b0 , \3129_b0 , w_5163 );
and ( w_5162 , w_5163 , \3130_b0 );
or ( \3132_b1 , \3129_b1 , \3130_b1 );
xor ( \3132_b0 , \3129_b0 , w_5164 );
not ( w_5164 , w_5165 );
and ( w_5165 , \3130_b1 , \3130_b0 );
or ( \3133_b1 , \3035_b1 , \3080_b1 );
xor ( \3133_b0 , \3035_b0 , w_5166 );
not ( w_5166 , w_5167 );
and ( w_5167 , \3080_b1 , \3080_b0 );
or ( \3134_b1 , \2959_A[7]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5168 );
and ( \3134_b0 , \2959_A[7]_b0 , w_5169 );
and ( w_5168 , w_5169 , \3000_B[2]_b0 );
or ( \3135_b1 , \3133_b1 , \3134_b1 );
not ( \3134_b1 , w_5170 );
and ( \3135_b0 , \3133_b0 , w_5171 );
and ( w_5170 , w_5171 , \3134_b0 );
or ( \3136_b1 , \3133_b1 , \3134_b1 );
xor ( \3136_b0 , \3133_b0 , w_5172 );
not ( w_5172 , w_5173 );
and ( w_5173 , \3134_b1 , \3134_b0 );
or ( \3137_b1 , \3039_b1 , \3078_b1 );
xor ( \3137_b0 , \3039_b0 , w_5174 );
not ( w_5174 , w_5175 );
and ( w_5175 , \3078_b1 , \3078_b0 );
or ( \3138_b1 , \2963_A[6]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5176 );
and ( \3138_b0 , \2963_A[6]_b0 , w_5177 );
and ( w_5176 , w_5177 , \3000_B[2]_b0 );
or ( \3139_b1 , \3137_b1 , \3138_b1 );
not ( \3138_b1 , w_5178 );
and ( \3139_b0 , \3137_b0 , w_5179 );
and ( w_5178 , w_5179 , \3138_b0 );
or ( \3140_b1 , \3137_b1 , \3138_b1 );
xor ( \3140_b0 , \3137_b0 , w_5180 );
not ( w_5180 , w_5181 );
and ( w_5181 , \3138_b1 , \3138_b0 );
or ( \3141_b1 , \3043_b1 , \3076_b1 );
xor ( \3141_b0 , \3043_b0 , w_5182 );
not ( w_5182 , w_5183 );
and ( w_5183 , \3076_b1 , \3076_b0 );
or ( \3142_b1 , \2967_A[5]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5184 );
and ( \3142_b0 , \2967_A[5]_b0 , w_5185 );
and ( w_5184 , w_5185 , \3000_B[2]_b0 );
or ( \3143_b1 , \3141_b1 , \3142_b1 );
not ( \3142_b1 , w_5186 );
and ( \3143_b0 , \3141_b0 , w_5187 );
and ( w_5186 , w_5187 , \3142_b0 );
or ( \3144_b1 , \3141_b1 , \3142_b1 );
xor ( \3144_b0 , \3141_b0 , w_5188 );
not ( w_5188 , w_5189 );
and ( w_5189 , \3142_b1 , \3142_b0 );
or ( \3145_b1 , \3047_b1 , \3074_b1 );
xor ( \3145_b0 , \3047_b0 , w_5190 );
not ( w_5190 , w_5191 );
and ( w_5191 , \3074_b1 , \3074_b0 );
or ( \3146_b1 , \2971_A[4]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5192 );
and ( \3146_b0 , \2971_A[4]_b0 , w_5193 );
and ( w_5192 , w_5193 , \3000_B[2]_b0 );
or ( \3147_b1 , \3145_b1 , \3146_b1 );
not ( \3146_b1 , w_5194 );
and ( \3147_b0 , \3145_b0 , w_5195 );
and ( w_5194 , w_5195 , \3146_b0 );
or ( \3148_b1 , \3145_b1 , \3146_b1 );
xor ( \3148_b0 , \3145_b0 , w_5196 );
not ( w_5196 , w_5197 );
and ( w_5197 , \3146_b1 , \3146_b0 );
or ( \3149_b1 , \3051_b1 , \3072_b1 );
xor ( \3149_b0 , \3051_b0 , w_5198 );
not ( w_5198 , w_5199 );
and ( w_5199 , \3072_b1 , \3072_b0 );
or ( \3150_b1 , \2975_A[3]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5200 );
and ( \3150_b0 , \2975_A[3]_b0 , w_5201 );
and ( w_5200 , w_5201 , \3000_B[2]_b0 );
or ( \3151_b1 , \3149_b1 , \3150_b1 );
not ( \3150_b1 , w_5202 );
and ( \3151_b0 , \3149_b0 , w_5203 );
and ( w_5202 , w_5203 , \3150_b0 );
or ( \3152_b1 , \3149_b1 , \3150_b1 );
xor ( \3152_b0 , \3149_b0 , w_5204 );
not ( w_5204 , w_5205 );
and ( w_5205 , \3150_b1 , \3150_b0 );
or ( \3153_b1 , \3055_b1 , \3070_b1 );
xor ( \3153_b0 , \3055_b0 , w_5206 );
not ( w_5206 , w_5207 );
and ( w_5207 , \3070_b1 , \3070_b0 );
or ( \3154_b1 , \2979_A[2]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5208 );
and ( \3154_b0 , \2979_A[2]_b0 , w_5209 );
and ( w_5208 , w_5209 , \3000_B[2]_b0 );
or ( \3155_b1 , \3153_b1 , \3154_b1 );
not ( \3154_b1 , w_5210 );
and ( \3155_b0 , \3153_b0 , w_5211 );
and ( w_5210 , w_5211 , \3154_b0 );
or ( \3156_b1 , \3153_b1 , \3154_b1 );
xor ( \3156_b0 , \3153_b0 , w_5212 );
not ( w_5212 , w_5213 );
and ( w_5213 , \3154_b1 , \3154_b0 );
or ( \3157_b1 , \3059_b1 , \3068_b1 );
xor ( \3157_b0 , \3059_b0 , w_5214 );
not ( w_5214 , w_5215 );
and ( w_5215 , \3068_b1 , \3068_b0 );
or ( \3158_b1 , \2983_A[1]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5216 );
and ( \3158_b0 , \2983_A[1]_b0 , w_5217 );
and ( w_5216 , w_5217 , \3000_B[2]_b0 );
or ( \3159_b1 , \3157_b1 , \3158_b1 );
not ( \3158_b1 , w_5218 );
and ( \3159_b0 , \3157_b0 , w_5219 );
and ( w_5218 , w_5219 , \3158_b0 );
or ( \3160_b1 , \3157_b1 , \3158_b1 );
xor ( \3160_b0 , \3157_b0 , w_5220 );
not ( w_5220 , w_5221 );
and ( w_5221 , \3158_b1 , \3158_b0 );
or ( \3161_b1 , \3063_b1 , \3066_b1 );
xor ( \3161_b0 , \3063_b0 , w_5222 );
not ( w_5222 , w_5223 );
and ( w_5223 , \3066_b1 , \3066_b0 );
or ( \3162_b1 , \2986_A[0]_b1 , \3000_B[2]_b1 );
not ( \3000_B[2]_b1 , w_5224 );
and ( \3162_b0 , \2986_A[0]_b0 , w_5225 );
and ( w_5224 , w_5225 , \3000_B[2]_b0 );
or ( \3163_b1 , \3161_b1 , \3162_b1 );
not ( \3162_b1 , w_5226 );
and ( \3163_b0 , \3161_b0 , w_5227 );
and ( w_5226 , w_5227 , \3162_b0 );
or ( \3164_b1 , \3160_b1 , \3163_b1 );
not ( \3163_b1 , w_5228 );
and ( \3164_b0 , \3160_b0 , w_5229 );
and ( w_5228 , w_5229 , \3163_b0 );
or ( \3165_b1 , \3159_b1 , w_5230 );
or ( \3165_b0 , \3159_b0 , \3164_b0 );
not ( \3164_b0 , w_5231 );
and ( w_5231 , w_5230 , \3164_b1 );
or ( \3166_b1 , \3156_b1 , \3165_b1 );
not ( \3165_b1 , w_5232 );
and ( \3166_b0 , \3156_b0 , w_5233 );
and ( w_5232 , w_5233 , \3165_b0 );
or ( \3167_b1 , \3155_b1 , w_5234 );
or ( \3167_b0 , \3155_b0 , \3166_b0 );
not ( \3166_b0 , w_5235 );
and ( w_5235 , w_5234 , \3166_b1 );
or ( \3168_b1 , \3152_b1 , \3167_b1 );
not ( \3167_b1 , w_5236 );
and ( \3168_b0 , \3152_b0 , w_5237 );
and ( w_5236 , w_5237 , \3167_b0 );
or ( \3169_b1 , \3151_b1 , w_5238 );
or ( \3169_b0 , \3151_b0 , \3168_b0 );
not ( \3168_b0 , w_5239 );
and ( w_5239 , w_5238 , \3168_b1 );
or ( \3170_b1 , \3148_b1 , \3169_b1 );
not ( \3169_b1 , w_5240 );
and ( \3170_b0 , \3148_b0 , w_5241 );
and ( w_5240 , w_5241 , \3169_b0 );
or ( \3171_b1 , \3147_b1 , w_5242 );
or ( \3171_b0 , \3147_b0 , \3170_b0 );
not ( \3170_b0 , w_5243 );
and ( w_5243 , w_5242 , \3170_b1 );
or ( \3172_b1 , \3144_b1 , \3171_b1 );
not ( \3171_b1 , w_5244 );
and ( \3172_b0 , \3144_b0 , w_5245 );
and ( w_5244 , w_5245 , \3171_b0 );
or ( \3173_b1 , \3143_b1 , w_5246 );
or ( \3173_b0 , \3143_b0 , \3172_b0 );
not ( \3172_b0 , w_5247 );
and ( w_5247 , w_5246 , \3172_b1 );
or ( \3174_b1 , \3140_b1 , \3173_b1 );
not ( \3173_b1 , w_5248 );
and ( \3174_b0 , \3140_b0 , w_5249 );
and ( w_5248 , w_5249 , \3173_b0 );
or ( \3175_b1 , \3139_b1 , w_5250 );
or ( \3175_b0 , \3139_b0 , \3174_b0 );
not ( \3174_b0 , w_5251 );
and ( w_5251 , w_5250 , \3174_b1 );
or ( \3176_b1 , \3136_b1 , \3175_b1 );
not ( \3175_b1 , w_5252 );
and ( \3176_b0 , \3136_b0 , w_5253 );
and ( w_5252 , w_5253 , \3175_b0 );
or ( \3177_b1 , \3135_b1 , w_5254 );
or ( \3177_b0 , \3135_b0 , \3176_b0 );
not ( \3176_b0 , w_5255 );
and ( w_5255 , w_5254 , \3176_b1 );
or ( \3178_b1 , \3132_b1 , \3177_b1 );
not ( \3177_b1 , w_5256 );
and ( \3178_b0 , \3132_b0 , w_5257 );
and ( w_5256 , w_5257 , \3177_b0 );
or ( \3179_b1 , \3131_b1 , w_5258 );
or ( \3179_b0 , \3131_b0 , \3178_b0 );
not ( \3178_b0 , w_5259 );
and ( w_5259 , w_5258 , \3178_b1 );
or ( \3180_b1 , \3128_b1 , \3179_b1 );
not ( \3179_b1 , w_5260 );
and ( \3180_b0 , \3128_b0 , w_5261 );
and ( w_5260 , w_5261 , \3179_b0 );
or ( \3181_b1 , \3127_b1 , w_5262 );
or ( \3181_b0 , \3127_b0 , \3180_b0 );
not ( \3180_b0 , w_5263 );
and ( w_5263 , w_5262 , \3180_b1 );
or ( \3182_b1 , \3124_b1 , \3181_b1 );
not ( \3181_b1 , w_5264 );
and ( \3182_b0 , \3124_b0 , w_5265 );
and ( w_5264 , w_5265 , \3181_b0 );
or ( \3183_b1 , \3123_b1 , w_5266 );
or ( \3183_b0 , \3123_b0 , \3182_b0 );
not ( \3182_b0 , w_5267 );
and ( w_5267 , w_5266 , \3182_b1 );
or ( \3184_b1 , \3120_b1 , \3183_b1 );
not ( \3183_b1 , w_5268 );
and ( \3184_b0 , \3120_b0 , w_5269 );
and ( w_5268 , w_5269 , \3183_b0 );
or ( \3185_b1 , \3119_b1 , w_5270 );
or ( \3185_b0 , \3119_b0 , \3184_b0 );
not ( \3184_b0 , w_5271 );
and ( w_5271 , w_5270 , \3184_b1 );
or ( \3186_b1 , \3116_b1 , \3185_b1 );
not ( \3185_b1 , w_5272 );
and ( \3186_b0 , \3116_b0 , w_5273 );
and ( w_5272 , w_5273 , \3185_b0 );
or ( \3187_b1 , \3115_b1 , w_5274 );
or ( \3187_b0 , \3115_b0 , \3186_b0 );
not ( \3186_b0 , w_5275 );
and ( w_5275 , w_5274 , \3186_b1 );
or ( \3188_b1 , \3112_b1 , \3187_b1 );
not ( \3187_b1 , w_5276 );
and ( \3188_b0 , \3112_b0 , w_5277 );
and ( w_5276 , w_5277 , \3187_b0 );
or ( \3189_b1 , \3111_b1 , w_5278 );
or ( \3189_b0 , \3111_b0 , \3188_b0 );
not ( \3188_b0 , w_5279 );
and ( w_5279 , w_5278 , \3188_b1 );
or ( \3190_b1 , \3108_b1 , \3189_b1 );
not ( \3189_b1 , w_5280 );
and ( \3190_b0 , \3108_b0 , w_5281 );
and ( w_5280 , w_5281 , \3189_b0 );
or ( \3191_b1 , \3107_b1 , w_5282 );
or ( \3191_b0 , \3107_b0 , \3190_b0 );
not ( \3190_b0 , w_5283 );
and ( w_5283 , w_5282 , \3190_b1 );
or ( \3192_b1 , \3104_b1 , \3191_b1 );
not ( \3191_b1 , w_5284 );
and ( \3192_b0 , \3104_b0 , w_5285 );
and ( w_5284 , w_5285 , \3191_b0 );
or ( \3193_b1 , \3103_b1 , w_5286 );
or ( \3193_b0 , \3103_b0 , \3192_b0 );
not ( \3192_b0 , w_5287 );
and ( w_5287 , w_5286 , \3192_b1 );
or ( \3194_b1 , \3100_b1 , \3193_b1 );
not ( \3193_b1 , w_5288 );
and ( \3194_b0 , \3100_b0 , w_5289 );
and ( w_5288 , w_5289 , \3193_b0 );
or ( \3195_b1 , \3099_b1 , w_5290 );
or ( \3195_b0 , \3099_b0 , \3194_b0 );
not ( \3194_b0 , w_5291 );
and ( w_5291 , w_5290 , \3194_b1 );
or ( \3196_b1 , \2923_A[16]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5292 );
and ( \3196_b0 , \2923_A[16]_b0 , w_5293 );
and ( w_5292 , w_5293 , \2999_B[3]_b0 );
or ( \3197_b1 , \3195_b1 , \3196_b1 );
not ( \3196_b1 , w_5294 );
and ( \3197_b0 , \3195_b0 , w_5295 );
and ( w_5294 , w_5295 , \3196_b0 );
or ( \3198_b1 , \3195_b1 , \3196_b1 );
xor ( \3198_b0 , \3195_b0 , w_5296 );
not ( w_5296 , w_5297 );
and ( w_5297 , \3196_b1 , \3196_b0 );
or ( \3199_b1 , \3100_b1 , \3193_b1 );
xor ( \3199_b0 , \3100_b0 , w_5298 );
not ( w_5298 , w_5299 );
and ( w_5299 , \3193_b1 , \3193_b0 );
or ( \3200_b1 , \2927_A[15]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5300 );
and ( \3200_b0 , \2927_A[15]_b0 , w_5301 );
and ( w_5300 , w_5301 , \2999_B[3]_b0 );
or ( \3201_b1 , \3199_b1 , \3200_b1 );
not ( \3200_b1 , w_5302 );
and ( \3201_b0 , \3199_b0 , w_5303 );
and ( w_5302 , w_5303 , \3200_b0 );
or ( \3202_b1 , \3199_b1 , \3200_b1 );
xor ( \3202_b0 , \3199_b0 , w_5304 );
not ( w_5304 , w_5305 );
and ( w_5305 , \3200_b1 , \3200_b0 );
or ( \3203_b1 , \3104_b1 , \3191_b1 );
xor ( \3203_b0 , \3104_b0 , w_5306 );
not ( w_5306 , w_5307 );
and ( w_5307 , \3191_b1 , \3191_b0 );
or ( \3204_b1 , \2931_A[14]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5308 );
and ( \3204_b0 , \2931_A[14]_b0 , w_5309 );
and ( w_5308 , w_5309 , \2999_B[3]_b0 );
or ( \3205_b1 , \3203_b1 , \3204_b1 );
not ( \3204_b1 , w_5310 );
and ( \3205_b0 , \3203_b0 , w_5311 );
and ( w_5310 , w_5311 , \3204_b0 );
or ( \3206_b1 , \3203_b1 , \3204_b1 );
xor ( \3206_b0 , \3203_b0 , w_5312 );
not ( w_5312 , w_5313 );
and ( w_5313 , \3204_b1 , \3204_b0 );
or ( \3207_b1 , \3108_b1 , \3189_b1 );
xor ( \3207_b0 , \3108_b0 , w_5314 );
not ( w_5314 , w_5315 );
and ( w_5315 , \3189_b1 , \3189_b0 );
or ( \3208_b1 , \2935_A[13]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5316 );
and ( \3208_b0 , \2935_A[13]_b0 , w_5317 );
and ( w_5316 , w_5317 , \2999_B[3]_b0 );
or ( \3209_b1 , \3207_b1 , \3208_b1 );
not ( \3208_b1 , w_5318 );
and ( \3209_b0 , \3207_b0 , w_5319 );
and ( w_5318 , w_5319 , \3208_b0 );
or ( \3210_b1 , \3207_b1 , \3208_b1 );
xor ( \3210_b0 , \3207_b0 , w_5320 );
not ( w_5320 , w_5321 );
and ( w_5321 , \3208_b1 , \3208_b0 );
or ( \3211_b1 , \3112_b1 , \3187_b1 );
xor ( \3211_b0 , \3112_b0 , w_5322 );
not ( w_5322 , w_5323 );
and ( w_5323 , \3187_b1 , \3187_b0 );
or ( \3212_b1 , \2939_A[12]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5324 );
and ( \3212_b0 , \2939_A[12]_b0 , w_5325 );
and ( w_5324 , w_5325 , \2999_B[3]_b0 );
or ( \3213_b1 , \3211_b1 , \3212_b1 );
not ( \3212_b1 , w_5326 );
and ( \3213_b0 , \3211_b0 , w_5327 );
and ( w_5326 , w_5327 , \3212_b0 );
or ( \3214_b1 , \3211_b1 , \3212_b1 );
xor ( \3214_b0 , \3211_b0 , w_5328 );
not ( w_5328 , w_5329 );
and ( w_5329 , \3212_b1 , \3212_b0 );
or ( \3215_b1 , \3116_b1 , \3185_b1 );
xor ( \3215_b0 , \3116_b0 , w_5330 );
not ( w_5330 , w_5331 );
and ( w_5331 , \3185_b1 , \3185_b0 );
or ( \3216_b1 , \2943_A[11]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5332 );
and ( \3216_b0 , \2943_A[11]_b0 , w_5333 );
and ( w_5332 , w_5333 , \2999_B[3]_b0 );
or ( \3217_b1 , \3215_b1 , \3216_b1 );
not ( \3216_b1 , w_5334 );
and ( \3217_b0 , \3215_b0 , w_5335 );
and ( w_5334 , w_5335 , \3216_b0 );
or ( \3218_b1 , \3215_b1 , \3216_b1 );
xor ( \3218_b0 , \3215_b0 , w_5336 );
not ( w_5336 , w_5337 );
and ( w_5337 , \3216_b1 , \3216_b0 );
or ( \3219_b1 , \3120_b1 , \3183_b1 );
xor ( \3219_b0 , \3120_b0 , w_5338 );
not ( w_5338 , w_5339 );
and ( w_5339 , \3183_b1 , \3183_b0 );
or ( \3220_b1 , \2947_A[10]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5340 );
and ( \3220_b0 , \2947_A[10]_b0 , w_5341 );
and ( w_5340 , w_5341 , \2999_B[3]_b0 );
or ( \3221_b1 , \3219_b1 , \3220_b1 );
not ( \3220_b1 , w_5342 );
and ( \3221_b0 , \3219_b0 , w_5343 );
and ( w_5342 , w_5343 , \3220_b0 );
or ( \3222_b1 , \3219_b1 , \3220_b1 );
xor ( \3222_b0 , \3219_b0 , w_5344 );
not ( w_5344 , w_5345 );
and ( w_5345 , \3220_b1 , \3220_b0 );
or ( \3223_b1 , \3124_b1 , \3181_b1 );
xor ( \3223_b0 , \3124_b0 , w_5346 );
not ( w_5346 , w_5347 );
and ( w_5347 , \3181_b1 , \3181_b0 );
or ( \3224_b1 , \2951_A[9]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5348 );
and ( \3224_b0 , \2951_A[9]_b0 , w_5349 );
and ( w_5348 , w_5349 , \2999_B[3]_b0 );
or ( \3225_b1 , \3223_b1 , \3224_b1 );
not ( \3224_b1 , w_5350 );
and ( \3225_b0 , \3223_b0 , w_5351 );
and ( w_5350 , w_5351 , \3224_b0 );
or ( \3226_b1 , \3223_b1 , \3224_b1 );
xor ( \3226_b0 , \3223_b0 , w_5352 );
not ( w_5352 , w_5353 );
and ( w_5353 , \3224_b1 , \3224_b0 );
or ( \3227_b1 , \3128_b1 , \3179_b1 );
xor ( \3227_b0 , \3128_b0 , w_5354 );
not ( w_5354 , w_5355 );
and ( w_5355 , \3179_b1 , \3179_b0 );
or ( \3228_b1 , \2955_A[8]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5356 );
and ( \3228_b0 , \2955_A[8]_b0 , w_5357 );
and ( w_5356 , w_5357 , \2999_B[3]_b0 );
or ( \3229_b1 , \3227_b1 , \3228_b1 );
not ( \3228_b1 , w_5358 );
and ( \3229_b0 , \3227_b0 , w_5359 );
and ( w_5358 , w_5359 , \3228_b0 );
or ( \3230_b1 , \3227_b1 , \3228_b1 );
xor ( \3230_b0 , \3227_b0 , w_5360 );
not ( w_5360 , w_5361 );
and ( w_5361 , \3228_b1 , \3228_b0 );
or ( \3231_b1 , \3132_b1 , \3177_b1 );
xor ( \3231_b0 , \3132_b0 , w_5362 );
not ( w_5362 , w_5363 );
and ( w_5363 , \3177_b1 , \3177_b0 );
or ( \3232_b1 , \2959_A[7]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5364 );
and ( \3232_b0 , \2959_A[7]_b0 , w_5365 );
and ( w_5364 , w_5365 , \2999_B[3]_b0 );
or ( \3233_b1 , \3231_b1 , \3232_b1 );
not ( \3232_b1 , w_5366 );
and ( \3233_b0 , \3231_b0 , w_5367 );
and ( w_5366 , w_5367 , \3232_b0 );
or ( \3234_b1 , \3231_b1 , \3232_b1 );
xor ( \3234_b0 , \3231_b0 , w_5368 );
not ( w_5368 , w_5369 );
and ( w_5369 , \3232_b1 , \3232_b0 );
or ( \3235_b1 , \3136_b1 , \3175_b1 );
xor ( \3235_b0 , \3136_b0 , w_5370 );
not ( w_5370 , w_5371 );
and ( w_5371 , \3175_b1 , \3175_b0 );
or ( \3236_b1 , \2963_A[6]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5372 );
and ( \3236_b0 , \2963_A[6]_b0 , w_5373 );
and ( w_5372 , w_5373 , \2999_B[3]_b0 );
or ( \3237_b1 , \3235_b1 , \3236_b1 );
not ( \3236_b1 , w_5374 );
and ( \3237_b0 , \3235_b0 , w_5375 );
and ( w_5374 , w_5375 , \3236_b0 );
or ( \3238_b1 , \3235_b1 , \3236_b1 );
xor ( \3238_b0 , \3235_b0 , w_5376 );
not ( w_5376 , w_5377 );
and ( w_5377 , \3236_b1 , \3236_b0 );
or ( \3239_b1 , \3140_b1 , \3173_b1 );
xor ( \3239_b0 , \3140_b0 , w_5378 );
not ( w_5378 , w_5379 );
and ( w_5379 , \3173_b1 , \3173_b0 );
or ( \3240_b1 , \2967_A[5]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5380 );
and ( \3240_b0 , \2967_A[5]_b0 , w_5381 );
and ( w_5380 , w_5381 , \2999_B[3]_b0 );
or ( \3241_b1 , \3239_b1 , \3240_b1 );
not ( \3240_b1 , w_5382 );
and ( \3241_b0 , \3239_b0 , w_5383 );
and ( w_5382 , w_5383 , \3240_b0 );
or ( \3242_b1 , \3239_b1 , \3240_b1 );
xor ( \3242_b0 , \3239_b0 , w_5384 );
not ( w_5384 , w_5385 );
and ( w_5385 , \3240_b1 , \3240_b0 );
or ( \3243_b1 , \3144_b1 , \3171_b1 );
xor ( \3243_b0 , \3144_b0 , w_5386 );
not ( w_5386 , w_5387 );
and ( w_5387 , \3171_b1 , \3171_b0 );
or ( \3244_b1 , \2971_A[4]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5388 );
and ( \3244_b0 , \2971_A[4]_b0 , w_5389 );
and ( w_5388 , w_5389 , \2999_B[3]_b0 );
or ( \3245_b1 , \3243_b1 , \3244_b1 );
not ( \3244_b1 , w_5390 );
and ( \3245_b0 , \3243_b0 , w_5391 );
and ( w_5390 , w_5391 , \3244_b0 );
or ( \3246_b1 , \3243_b1 , \3244_b1 );
xor ( \3246_b0 , \3243_b0 , w_5392 );
not ( w_5392 , w_5393 );
and ( w_5393 , \3244_b1 , \3244_b0 );
or ( \3247_b1 , \3148_b1 , \3169_b1 );
xor ( \3247_b0 , \3148_b0 , w_5394 );
not ( w_5394 , w_5395 );
and ( w_5395 , \3169_b1 , \3169_b0 );
or ( \3248_b1 , \2975_A[3]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5396 );
and ( \3248_b0 , \2975_A[3]_b0 , w_5397 );
and ( w_5396 , w_5397 , \2999_B[3]_b0 );
or ( \3249_b1 , \3247_b1 , \3248_b1 );
not ( \3248_b1 , w_5398 );
and ( \3249_b0 , \3247_b0 , w_5399 );
and ( w_5398 , w_5399 , \3248_b0 );
or ( \3250_b1 , \3247_b1 , \3248_b1 );
xor ( \3250_b0 , \3247_b0 , w_5400 );
not ( w_5400 , w_5401 );
and ( w_5401 , \3248_b1 , \3248_b0 );
or ( \3251_b1 , \3152_b1 , \3167_b1 );
xor ( \3251_b0 , \3152_b0 , w_5402 );
not ( w_5402 , w_5403 );
and ( w_5403 , \3167_b1 , \3167_b0 );
or ( \3252_b1 , \2979_A[2]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5404 );
and ( \3252_b0 , \2979_A[2]_b0 , w_5405 );
and ( w_5404 , w_5405 , \2999_B[3]_b0 );
or ( \3253_b1 , \3251_b1 , \3252_b1 );
not ( \3252_b1 , w_5406 );
and ( \3253_b0 , \3251_b0 , w_5407 );
and ( w_5406 , w_5407 , \3252_b0 );
or ( \3254_b1 , \3251_b1 , \3252_b1 );
xor ( \3254_b0 , \3251_b0 , w_5408 );
not ( w_5408 , w_5409 );
and ( w_5409 , \3252_b1 , \3252_b0 );
or ( \3255_b1 , \3156_b1 , \3165_b1 );
xor ( \3255_b0 , \3156_b0 , w_5410 );
not ( w_5410 , w_5411 );
and ( w_5411 , \3165_b1 , \3165_b0 );
or ( \3256_b1 , \2983_A[1]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5412 );
and ( \3256_b0 , \2983_A[1]_b0 , w_5413 );
and ( w_5412 , w_5413 , \2999_B[3]_b0 );
or ( \3257_b1 , \3255_b1 , \3256_b1 );
not ( \3256_b1 , w_5414 );
and ( \3257_b0 , \3255_b0 , w_5415 );
and ( w_5414 , w_5415 , \3256_b0 );
or ( \3258_b1 , \3255_b1 , \3256_b1 );
xor ( \3258_b0 , \3255_b0 , w_5416 );
not ( w_5416 , w_5417 );
and ( w_5417 , \3256_b1 , \3256_b0 );
or ( \3259_b1 , \3160_b1 , \3163_b1 );
xor ( \3259_b0 , \3160_b0 , w_5418 );
not ( w_5418 , w_5419 );
and ( w_5419 , \3163_b1 , \3163_b0 );
or ( \3260_b1 , \2986_A[0]_b1 , \2999_B[3]_b1 );
not ( \2999_B[3]_b1 , w_5420 );
and ( \3260_b0 , \2986_A[0]_b0 , w_5421 );
and ( w_5420 , w_5421 , \2999_B[3]_b0 );
or ( \3261_b1 , \3259_b1 , \3260_b1 );
not ( \3260_b1 , w_5422 );
and ( \3261_b0 , \3259_b0 , w_5423 );
and ( w_5422 , w_5423 , \3260_b0 );
or ( \3262_b1 , \3258_b1 , \3261_b1 );
not ( \3261_b1 , w_5424 );
and ( \3262_b0 , \3258_b0 , w_5425 );
and ( w_5424 , w_5425 , \3261_b0 );
or ( \3263_b1 , \3257_b1 , w_5426 );
or ( \3263_b0 , \3257_b0 , \3262_b0 );
not ( \3262_b0 , w_5427 );
and ( w_5427 , w_5426 , \3262_b1 );
or ( \3264_b1 , \3254_b1 , \3263_b1 );
not ( \3263_b1 , w_5428 );
and ( \3264_b0 , \3254_b0 , w_5429 );
and ( w_5428 , w_5429 , \3263_b0 );
or ( \3265_b1 , \3253_b1 , w_5430 );
or ( \3265_b0 , \3253_b0 , \3264_b0 );
not ( \3264_b0 , w_5431 );
and ( w_5431 , w_5430 , \3264_b1 );
or ( \3266_b1 , \3250_b1 , \3265_b1 );
not ( \3265_b1 , w_5432 );
and ( \3266_b0 , \3250_b0 , w_5433 );
and ( w_5432 , w_5433 , \3265_b0 );
or ( \3267_b1 , \3249_b1 , w_5434 );
or ( \3267_b0 , \3249_b0 , \3266_b0 );
not ( \3266_b0 , w_5435 );
and ( w_5435 , w_5434 , \3266_b1 );
or ( \3268_b1 , \3246_b1 , \3267_b1 );
not ( \3267_b1 , w_5436 );
and ( \3268_b0 , \3246_b0 , w_5437 );
and ( w_5436 , w_5437 , \3267_b0 );
or ( \3269_b1 , \3245_b1 , w_5438 );
or ( \3269_b0 , \3245_b0 , \3268_b0 );
not ( \3268_b0 , w_5439 );
and ( w_5439 , w_5438 , \3268_b1 );
or ( \3270_b1 , \3242_b1 , \3269_b1 );
not ( \3269_b1 , w_5440 );
and ( \3270_b0 , \3242_b0 , w_5441 );
and ( w_5440 , w_5441 , \3269_b0 );
or ( \3271_b1 , \3241_b1 , w_5442 );
or ( \3271_b0 , \3241_b0 , \3270_b0 );
not ( \3270_b0 , w_5443 );
and ( w_5443 , w_5442 , \3270_b1 );
or ( \3272_b1 , \3238_b1 , \3271_b1 );
not ( \3271_b1 , w_5444 );
and ( \3272_b0 , \3238_b0 , w_5445 );
and ( w_5444 , w_5445 , \3271_b0 );
or ( \3273_b1 , \3237_b1 , w_5446 );
or ( \3273_b0 , \3237_b0 , \3272_b0 );
not ( \3272_b0 , w_5447 );
and ( w_5447 , w_5446 , \3272_b1 );
or ( \3274_b1 , \3234_b1 , \3273_b1 );
not ( \3273_b1 , w_5448 );
and ( \3274_b0 , \3234_b0 , w_5449 );
and ( w_5448 , w_5449 , \3273_b0 );
or ( \3275_b1 , \3233_b1 , w_5450 );
or ( \3275_b0 , \3233_b0 , \3274_b0 );
not ( \3274_b0 , w_5451 );
and ( w_5451 , w_5450 , \3274_b1 );
or ( \3276_b1 , \3230_b1 , \3275_b1 );
not ( \3275_b1 , w_5452 );
and ( \3276_b0 , \3230_b0 , w_5453 );
and ( w_5452 , w_5453 , \3275_b0 );
or ( \3277_b1 , \3229_b1 , w_5454 );
or ( \3277_b0 , \3229_b0 , \3276_b0 );
not ( \3276_b0 , w_5455 );
and ( w_5455 , w_5454 , \3276_b1 );
or ( \3278_b1 , \3226_b1 , \3277_b1 );
not ( \3277_b1 , w_5456 );
and ( \3278_b0 , \3226_b0 , w_5457 );
and ( w_5456 , w_5457 , \3277_b0 );
or ( \3279_b1 , \3225_b1 , w_5458 );
or ( \3279_b0 , \3225_b0 , \3278_b0 );
not ( \3278_b0 , w_5459 );
and ( w_5459 , w_5458 , \3278_b1 );
or ( \3280_b1 , \3222_b1 , \3279_b1 );
not ( \3279_b1 , w_5460 );
and ( \3280_b0 , \3222_b0 , w_5461 );
and ( w_5460 , w_5461 , \3279_b0 );
or ( \3281_b1 , \3221_b1 , w_5462 );
or ( \3281_b0 , \3221_b0 , \3280_b0 );
not ( \3280_b0 , w_5463 );
and ( w_5463 , w_5462 , \3280_b1 );
or ( \3282_b1 , \3218_b1 , \3281_b1 );
not ( \3281_b1 , w_5464 );
and ( \3282_b0 , \3218_b0 , w_5465 );
and ( w_5464 , w_5465 , \3281_b0 );
or ( \3283_b1 , \3217_b1 , w_5466 );
or ( \3283_b0 , \3217_b0 , \3282_b0 );
not ( \3282_b0 , w_5467 );
and ( w_5467 , w_5466 , \3282_b1 );
or ( \3284_b1 , \3214_b1 , \3283_b1 );
not ( \3283_b1 , w_5468 );
and ( \3284_b0 , \3214_b0 , w_5469 );
and ( w_5468 , w_5469 , \3283_b0 );
or ( \3285_b1 , \3213_b1 , w_5470 );
or ( \3285_b0 , \3213_b0 , \3284_b0 );
not ( \3284_b0 , w_5471 );
and ( w_5471 , w_5470 , \3284_b1 );
or ( \3286_b1 , \3210_b1 , \3285_b1 );
not ( \3285_b1 , w_5472 );
and ( \3286_b0 , \3210_b0 , w_5473 );
and ( w_5472 , w_5473 , \3285_b0 );
or ( \3287_b1 , \3209_b1 , w_5474 );
or ( \3287_b0 , \3209_b0 , \3286_b0 );
not ( \3286_b0 , w_5475 );
and ( w_5475 , w_5474 , \3286_b1 );
or ( \3288_b1 , \3206_b1 , \3287_b1 );
not ( \3287_b1 , w_5476 );
and ( \3288_b0 , \3206_b0 , w_5477 );
and ( w_5476 , w_5477 , \3287_b0 );
or ( \3289_b1 , \3205_b1 , w_5478 );
or ( \3289_b0 , \3205_b0 , \3288_b0 );
not ( \3288_b0 , w_5479 );
and ( w_5479 , w_5478 , \3288_b1 );
or ( \3290_b1 , \3202_b1 , \3289_b1 );
not ( \3289_b1 , w_5480 );
and ( \3290_b0 , \3202_b0 , w_5481 );
and ( w_5480 , w_5481 , \3289_b0 );
or ( \3291_b1 , \3201_b1 , w_5482 );
or ( \3291_b0 , \3201_b0 , \3290_b0 );
not ( \3290_b0 , w_5483 );
and ( w_5483 , w_5482 , \3290_b1 );
or ( \3292_b1 , \3198_b1 , \3291_b1 );
not ( \3291_b1 , w_5484 );
and ( \3292_b0 , \3198_b0 , w_5485 );
and ( w_5484 , w_5485 , \3291_b0 );
or ( \3293_b1 , \3197_b1 , w_5486 );
or ( \3293_b0 , \3197_b0 , \3292_b0 );
not ( \3292_b0 , w_5487 );
and ( w_5487 , w_5486 , \3292_b1 );
or ( \3294_b1 , \2923_A[16]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5488 );
and ( \3294_b0 , \2923_A[16]_b0 , w_5489 );
and ( w_5488 , w_5489 , \2998_B[4]_b0 );
or ( \3295_b1 , \3293_b1 , \3294_b1 );
not ( \3294_b1 , w_5490 );
and ( \3295_b0 , \3293_b0 , w_5491 );
and ( w_5490 , w_5491 , \3294_b0 );
or ( \3296_b1 , \3293_b1 , \3294_b1 );
xor ( \3296_b0 , \3293_b0 , w_5492 );
not ( w_5492 , w_5493 );
and ( w_5493 , \3294_b1 , \3294_b0 );
or ( \3297_b1 , \3198_b1 , \3291_b1 );
xor ( \3297_b0 , \3198_b0 , w_5494 );
not ( w_5494 , w_5495 );
and ( w_5495 , \3291_b1 , \3291_b0 );
or ( \3298_b1 , \2927_A[15]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5496 );
and ( \3298_b0 , \2927_A[15]_b0 , w_5497 );
and ( w_5496 , w_5497 , \2998_B[4]_b0 );
or ( \3299_b1 , \3297_b1 , \3298_b1 );
not ( \3298_b1 , w_5498 );
and ( \3299_b0 , \3297_b0 , w_5499 );
and ( w_5498 , w_5499 , \3298_b0 );
or ( \3300_b1 , \3297_b1 , \3298_b1 );
xor ( \3300_b0 , \3297_b0 , w_5500 );
not ( w_5500 , w_5501 );
and ( w_5501 , \3298_b1 , \3298_b0 );
or ( \3301_b1 , \3202_b1 , \3289_b1 );
xor ( \3301_b0 , \3202_b0 , w_5502 );
not ( w_5502 , w_5503 );
and ( w_5503 , \3289_b1 , \3289_b0 );
or ( \3302_b1 , \2931_A[14]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5504 );
and ( \3302_b0 , \2931_A[14]_b0 , w_5505 );
and ( w_5504 , w_5505 , \2998_B[4]_b0 );
or ( \3303_b1 , \3301_b1 , \3302_b1 );
not ( \3302_b1 , w_5506 );
and ( \3303_b0 , \3301_b0 , w_5507 );
and ( w_5506 , w_5507 , \3302_b0 );
or ( \3304_b1 , \3301_b1 , \3302_b1 );
xor ( \3304_b0 , \3301_b0 , w_5508 );
not ( w_5508 , w_5509 );
and ( w_5509 , \3302_b1 , \3302_b0 );
or ( \3305_b1 , \3206_b1 , \3287_b1 );
xor ( \3305_b0 , \3206_b0 , w_5510 );
not ( w_5510 , w_5511 );
and ( w_5511 , \3287_b1 , \3287_b0 );
or ( \3306_b1 , \2935_A[13]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5512 );
and ( \3306_b0 , \2935_A[13]_b0 , w_5513 );
and ( w_5512 , w_5513 , \2998_B[4]_b0 );
or ( \3307_b1 , \3305_b1 , \3306_b1 );
not ( \3306_b1 , w_5514 );
and ( \3307_b0 , \3305_b0 , w_5515 );
and ( w_5514 , w_5515 , \3306_b0 );
or ( \3308_b1 , \3305_b1 , \3306_b1 );
xor ( \3308_b0 , \3305_b0 , w_5516 );
not ( w_5516 , w_5517 );
and ( w_5517 , \3306_b1 , \3306_b0 );
or ( \3309_b1 , \3210_b1 , \3285_b1 );
xor ( \3309_b0 , \3210_b0 , w_5518 );
not ( w_5518 , w_5519 );
and ( w_5519 , \3285_b1 , \3285_b0 );
or ( \3310_b1 , \2939_A[12]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5520 );
and ( \3310_b0 , \2939_A[12]_b0 , w_5521 );
and ( w_5520 , w_5521 , \2998_B[4]_b0 );
or ( \3311_b1 , \3309_b1 , \3310_b1 );
not ( \3310_b1 , w_5522 );
and ( \3311_b0 , \3309_b0 , w_5523 );
and ( w_5522 , w_5523 , \3310_b0 );
or ( \3312_b1 , \3309_b1 , \3310_b1 );
xor ( \3312_b0 , \3309_b0 , w_5524 );
not ( w_5524 , w_5525 );
and ( w_5525 , \3310_b1 , \3310_b0 );
or ( \3313_b1 , \3214_b1 , \3283_b1 );
xor ( \3313_b0 , \3214_b0 , w_5526 );
not ( w_5526 , w_5527 );
and ( w_5527 , \3283_b1 , \3283_b0 );
or ( \3314_b1 , \2943_A[11]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5528 );
and ( \3314_b0 , \2943_A[11]_b0 , w_5529 );
and ( w_5528 , w_5529 , \2998_B[4]_b0 );
or ( \3315_b1 , \3313_b1 , \3314_b1 );
not ( \3314_b1 , w_5530 );
and ( \3315_b0 , \3313_b0 , w_5531 );
and ( w_5530 , w_5531 , \3314_b0 );
or ( \3316_b1 , \3313_b1 , \3314_b1 );
xor ( \3316_b0 , \3313_b0 , w_5532 );
not ( w_5532 , w_5533 );
and ( w_5533 , \3314_b1 , \3314_b0 );
or ( \3317_b1 , \3218_b1 , \3281_b1 );
xor ( \3317_b0 , \3218_b0 , w_5534 );
not ( w_5534 , w_5535 );
and ( w_5535 , \3281_b1 , \3281_b0 );
or ( \3318_b1 , \2947_A[10]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5536 );
and ( \3318_b0 , \2947_A[10]_b0 , w_5537 );
and ( w_5536 , w_5537 , \2998_B[4]_b0 );
or ( \3319_b1 , \3317_b1 , \3318_b1 );
not ( \3318_b1 , w_5538 );
and ( \3319_b0 , \3317_b0 , w_5539 );
and ( w_5538 , w_5539 , \3318_b0 );
or ( \3320_b1 , \3317_b1 , \3318_b1 );
xor ( \3320_b0 , \3317_b0 , w_5540 );
not ( w_5540 , w_5541 );
and ( w_5541 , \3318_b1 , \3318_b0 );
or ( \3321_b1 , \3222_b1 , \3279_b1 );
xor ( \3321_b0 , \3222_b0 , w_5542 );
not ( w_5542 , w_5543 );
and ( w_5543 , \3279_b1 , \3279_b0 );
or ( \3322_b1 , \2951_A[9]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5544 );
and ( \3322_b0 , \2951_A[9]_b0 , w_5545 );
and ( w_5544 , w_5545 , \2998_B[4]_b0 );
or ( \3323_b1 , \3321_b1 , \3322_b1 );
not ( \3322_b1 , w_5546 );
and ( \3323_b0 , \3321_b0 , w_5547 );
and ( w_5546 , w_5547 , \3322_b0 );
or ( \3324_b1 , \3321_b1 , \3322_b1 );
xor ( \3324_b0 , \3321_b0 , w_5548 );
not ( w_5548 , w_5549 );
and ( w_5549 , \3322_b1 , \3322_b0 );
or ( \3325_b1 , \3226_b1 , \3277_b1 );
xor ( \3325_b0 , \3226_b0 , w_5550 );
not ( w_5550 , w_5551 );
and ( w_5551 , \3277_b1 , \3277_b0 );
or ( \3326_b1 , \2955_A[8]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5552 );
and ( \3326_b0 , \2955_A[8]_b0 , w_5553 );
and ( w_5552 , w_5553 , \2998_B[4]_b0 );
or ( \3327_b1 , \3325_b1 , \3326_b1 );
not ( \3326_b1 , w_5554 );
and ( \3327_b0 , \3325_b0 , w_5555 );
and ( w_5554 , w_5555 , \3326_b0 );
or ( \3328_b1 , \3325_b1 , \3326_b1 );
xor ( \3328_b0 , \3325_b0 , w_5556 );
not ( w_5556 , w_5557 );
and ( w_5557 , \3326_b1 , \3326_b0 );
or ( \3329_b1 , \3230_b1 , \3275_b1 );
xor ( \3329_b0 , \3230_b0 , w_5558 );
not ( w_5558 , w_5559 );
and ( w_5559 , \3275_b1 , \3275_b0 );
or ( \3330_b1 , \2959_A[7]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5560 );
and ( \3330_b0 , \2959_A[7]_b0 , w_5561 );
and ( w_5560 , w_5561 , \2998_B[4]_b0 );
or ( \3331_b1 , \3329_b1 , \3330_b1 );
not ( \3330_b1 , w_5562 );
and ( \3331_b0 , \3329_b0 , w_5563 );
and ( w_5562 , w_5563 , \3330_b0 );
or ( \3332_b1 , \3329_b1 , \3330_b1 );
xor ( \3332_b0 , \3329_b0 , w_5564 );
not ( w_5564 , w_5565 );
and ( w_5565 , \3330_b1 , \3330_b0 );
or ( \3333_b1 , \3234_b1 , \3273_b1 );
xor ( \3333_b0 , \3234_b0 , w_5566 );
not ( w_5566 , w_5567 );
and ( w_5567 , \3273_b1 , \3273_b0 );
or ( \3334_b1 , \2963_A[6]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5568 );
and ( \3334_b0 , \2963_A[6]_b0 , w_5569 );
and ( w_5568 , w_5569 , \2998_B[4]_b0 );
or ( \3335_b1 , \3333_b1 , \3334_b1 );
not ( \3334_b1 , w_5570 );
and ( \3335_b0 , \3333_b0 , w_5571 );
and ( w_5570 , w_5571 , \3334_b0 );
or ( \3336_b1 , \3333_b1 , \3334_b1 );
xor ( \3336_b0 , \3333_b0 , w_5572 );
not ( w_5572 , w_5573 );
and ( w_5573 , \3334_b1 , \3334_b0 );
or ( \3337_b1 , \3238_b1 , \3271_b1 );
xor ( \3337_b0 , \3238_b0 , w_5574 );
not ( w_5574 , w_5575 );
and ( w_5575 , \3271_b1 , \3271_b0 );
or ( \3338_b1 , \2967_A[5]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5576 );
and ( \3338_b0 , \2967_A[5]_b0 , w_5577 );
and ( w_5576 , w_5577 , \2998_B[4]_b0 );
or ( \3339_b1 , \3337_b1 , \3338_b1 );
not ( \3338_b1 , w_5578 );
and ( \3339_b0 , \3337_b0 , w_5579 );
and ( w_5578 , w_5579 , \3338_b0 );
or ( \3340_b1 , \3337_b1 , \3338_b1 );
xor ( \3340_b0 , \3337_b0 , w_5580 );
not ( w_5580 , w_5581 );
and ( w_5581 , \3338_b1 , \3338_b0 );
or ( \3341_b1 , \3242_b1 , \3269_b1 );
xor ( \3341_b0 , \3242_b0 , w_5582 );
not ( w_5582 , w_5583 );
and ( w_5583 , \3269_b1 , \3269_b0 );
or ( \3342_b1 , \2971_A[4]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5584 );
and ( \3342_b0 , \2971_A[4]_b0 , w_5585 );
and ( w_5584 , w_5585 , \2998_B[4]_b0 );
or ( \3343_b1 , \3341_b1 , \3342_b1 );
not ( \3342_b1 , w_5586 );
and ( \3343_b0 , \3341_b0 , w_5587 );
and ( w_5586 , w_5587 , \3342_b0 );
or ( \3344_b1 , \3341_b1 , \3342_b1 );
xor ( \3344_b0 , \3341_b0 , w_5588 );
not ( w_5588 , w_5589 );
and ( w_5589 , \3342_b1 , \3342_b0 );
or ( \3345_b1 , \3246_b1 , \3267_b1 );
xor ( \3345_b0 , \3246_b0 , w_5590 );
not ( w_5590 , w_5591 );
and ( w_5591 , \3267_b1 , \3267_b0 );
or ( \3346_b1 , \2975_A[3]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5592 );
and ( \3346_b0 , \2975_A[3]_b0 , w_5593 );
and ( w_5592 , w_5593 , \2998_B[4]_b0 );
or ( \3347_b1 , \3345_b1 , \3346_b1 );
not ( \3346_b1 , w_5594 );
and ( \3347_b0 , \3345_b0 , w_5595 );
and ( w_5594 , w_5595 , \3346_b0 );
or ( \3348_b1 , \3345_b1 , \3346_b1 );
xor ( \3348_b0 , \3345_b0 , w_5596 );
not ( w_5596 , w_5597 );
and ( w_5597 , \3346_b1 , \3346_b0 );
or ( \3349_b1 , \3250_b1 , \3265_b1 );
xor ( \3349_b0 , \3250_b0 , w_5598 );
not ( w_5598 , w_5599 );
and ( w_5599 , \3265_b1 , \3265_b0 );
or ( \3350_b1 , \2979_A[2]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5600 );
and ( \3350_b0 , \2979_A[2]_b0 , w_5601 );
and ( w_5600 , w_5601 , \2998_B[4]_b0 );
or ( \3351_b1 , \3349_b1 , \3350_b1 );
not ( \3350_b1 , w_5602 );
and ( \3351_b0 , \3349_b0 , w_5603 );
and ( w_5602 , w_5603 , \3350_b0 );
or ( \3352_b1 , \3349_b1 , \3350_b1 );
xor ( \3352_b0 , \3349_b0 , w_5604 );
not ( w_5604 , w_5605 );
and ( w_5605 , \3350_b1 , \3350_b0 );
or ( \3353_b1 , \3254_b1 , \3263_b1 );
xor ( \3353_b0 , \3254_b0 , w_5606 );
not ( w_5606 , w_5607 );
and ( w_5607 , \3263_b1 , \3263_b0 );
or ( \3354_b1 , \2983_A[1]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5608 );
and ( \3354_b0 , \2983_A[1]_b0 , w_5609 );
and ( w_5608 , w_5609 , \2998_B[4]_b0 );
or ( \3355_b1 , \3353_b1 , \3354_b1 );
not ( \3354_b1 , w_5610 );
and ( \3355_b0 , \3353_b0 , w_5611 );
and ( w_5610 , w_5611 , \3354_b0 );
or ( \3356_b1 , \3353_b1 , \3354_b1 );
xor ( \3356_b0 , \3353_b0 , w_5612 );
not ( w_5612 , w_5613 );
and ( w_5613 , \3354_b1 , \3354_b0 );
or ( \3357_b1 , \3258_b1 , \3261_b1 );
xor ( \3357_b0 , \3258_b0 , w_5614 );
not ( w_5614 , w_5615 );
and ( w_5615 , \3261_b1 , \3261_b0 );
or ( \3358_b1 , \2986_A[0]_b1 , \2998_B[4]_b1 );
not ( \2998_B[4]_b1 , w_5616 );
and ( \3358_b0 , \2986_A[0]_b0 , w_5617 );
and ( w_5616 , w_5617 , \2998_B[4]_b0 );
or ( \3359_b1 , \3357_b1 , \3358_b1 );
not ( \3358_b1 , w_5618 );
and ( \3359_b0 , \3357_b0 , w_5619 );
and ( w_5618 , w_5619 , \3358_b0 );
or ( \3360_b1 , \3356_b1 , \3359_b1 );
not ( \3359_b1 , w_5620 );
and ( \3360_b0 , \3356_b0 , w_5621 );
and ( w_5620 , w_5621 , \3359_b0 );
or ( \3361_b1 , \3355_b1 , w_5622 );
or ( \3361_b0 , \3355_b0 , \3360_b0 );
not ( \3360_b0 , w_5623 );
and ( w_5623 , w_5622 , \3360_b1 );
or ( \3362_b1 , \3352_b1 , \3361_b1 );
not ( \3361_b1 , w_5624 );
and ( \3362_b0 , \3352_b0 , w_5625 );
and ( w_5624 , w_5625 , \3361_b0 );
or ( \3363_b1 , \3351_b1 , w_5626 );
or ( \3363_b0 , \3351_b0 , \3362_b0 );
not ( \3362_b0 , w_5627 );
and ( w_5627 , w_5626 , \3362_b1 );
or ( \3364_b1 , \3348_b1 , \3363_b1 );
not ( \3363_b1 , w_5628 );
and ( \3364_b0 , \3348_b0 , w_5629 );
and ( w_5628 , w_5629 , \3363_b0 );
or ( \3365_b1 , \3347_b1 , w_5630 );
or ( \3365_b0 , \3347_b0 , \3364_b0 );
not ( \3364_b0 , w_5631 );
and ( w_5631 , w_5630 , \3364_b1 );
or ( \3366_b1 , \3344_b1 , \3365_b1 );
not ( \3365_b1 , w_5632 );
and ( \3366_b0 , \3344_b0 , w_5633 );
and ( w_5632 , w_5633 , \3365_b0 );
or ( \3367_b1 , \3343_b1 , w_5634 );
or ( \3367_b0 , \3343_b0 , \3366_b0 );
not ( \3366_b0 , w_5635 );
and ( w_5635 , w_5634 , \3366_b1 );
or ( \3368_b1 , \3340_b1 , \3367_b1 );
not ( \3367_b1 , w_5636 );
and ( \3368_b0 , \3340_b0 , w_5637 );
and ( w_5636 , w_5637 , \3367_b0 );
or ( \3369_b1 , \3339_b1 , w_5638 );
or ( \3369_b0 , \3339_b0 , \3368_b0 );
not ( \3368_b0 , w_5639 );
and ( w_5639 , w_5638 , \3368_b1 );
or ( \3370_b1 , \3336_b1 , \3369_b1 );
not ( \3369_b1 , w_5640 );
and ( \3370_b0 , \3336_b0 , w_5641 );
and ( w_5640 , w_5641 , \3369_b0 );
or ( \3371_b1 , \3335_b1 , w_5642 );
or ( \3371_b0 , \3335_b0 , \3370_b0 );
not ( \3370_b0 , w_5643 );
and ( w_5643 , w_5642 , \3370_b1 );
or ( \3372_b1 , \3332_b1 , \3371_b1 );
not ( \3371_b1 , w_5644 );
and ( \3372_b0 , \3332_b0 , w_5645 );
and ( w_5644 , w_5645 , \3371_b0 );
or ( \3373_b1 , \3331_b1 , w_5646 );
or ( \3373_b0 , \3331_b0 , \3372_b0 );
not ( \3372_b0 , w_5647 );
and ( w_5647 , w_5646 , \3372_b1 );
or ( \3374_b1 , \3328_b1 , \3373_b1 );
not ( \3373_b1 , w_5648 );
and ( \3374_b0 , \3328_b0 , w_5649 );
and ( w_5648 , w_5649 , \3373_b0 );
or ( \3375_b1 , \3327_b1 , w_5650 );
or ( \3375_b0 , \3327_b0 , \3374_b0 );
not ( \3374_b0 , w_5651 );
and ( w_5651 , w_5650 , \3374_b1 );
or ( \3376_b1 , \3324_b1 , \3375_b1 );
not ( \3375_b1 , w_5652 );
and ( \3376_b0 , \3324_b0 , w_5653 );
and ( w_5652 , w_5653 , \3375_b0 );
or ( \3377_b1 , \3323_b1 , w_5654 );
or ( \3377_b0 , \3323_b0 , \3376_b0 );
not ( \3376_b0 , w_5655 );
and ( w_5655 , w_5654 , \3376_b1 );
or ( \3378_b1 , \3320_b1 , \3377_b1 );
not ( \3377_b1 , w_5656 );
and ( \3378_b0 , \3320_b0 , w_5657 );
and ( w_5656 , w_5657 , \3377_b0 );
or ( \3379_b1 , \3319_b1 , w_5658 );
or ( \3379_b0 , \3319_b0 , \3378_b0 );
not ( \3378_b0 , w_5659 );
and ( w_5659 , w_5658 , \3378_b1 );
or ( \3380_b1 , \3316_b1 , \3379_b1 );
not ( \3379_b1 , w_5660 );
and ( \3380_b0 , \3316_b0 , w_5661 );
and ( w_5660 , w_5661 , \3379_b0 );
or ( \3381_b1 , \3315_b1 , w_5662 );
or ( \3381_b0 , \3315_b0 , \3380_b0 );
not ( \3380_b0 , w_5663 );
and ( w_5663 , w_5662 , \3380_b1 );
or ( \3382_b1 , \3312_b1 , \3381_b1 );
not ( \3381_b1 , w_5664 );
and ( \3382_b0 , \3312_b0 , w_5665 );
and ( w_5664 , w_5665 , \3381_b0 );
or ( \3383_b1 , \3311_b1 , w_5666 );
or ( \3383_b0 , \3311_b0 , \3382_b0 );
not ( \3382_b0 , w_5667 );
and ( w_5667 , w_5666 , \3382_b1 );
or ( \3384_b1 , \3308_b1 , \3383_b1 );
not ( \3383_b1 , w_5668 );
and ( \3384_b0 , \3308_b0 , w_5669 );
and ( w_5668 , w_5669 , \3383_b0 );
or ( \3385_b1 , \3307_b1 , w_5670 );
or ( \3385_b0 , \3307_b0 , \3384_b0 );
not ( \3384_b0 , w_5671 );
and ( w_5671 , w_5670 , \3384_b1 );
or ( \3386_b1 , \3304_b1 , \3385_b1 );
not ( \3385_b1 , w_5672 );
and ( \3386_b0 , \3304_b0 , w_5673 );
and ( w_5672 , w_5673 , \3385_b0 );
or ( \3387_b1 , \3303_b1 , w_5674 );
or ( \3387_b0 , \3303_b0 , \3386_b0 );
not ( \3386_b0 , w_5675 );
and ( w_5675 , w_5674 , \3386_b1 );
or ( \3388_b1 , \3300_b1 , \3387_b1 );
not ( \3387_b1 , w_5676 );
and ( \3388_b0 , \3300_b0 , w_5677 );
and ( w_5676 , w_5677 , \3387_b0 );
or ( \3389_b1 , \3299_b1 , w_5678 );
or ( \3389_b0 , \3299_b0 , \3388_b0 );
not ( \3388_b0 , w_5679 );
and ( w_5679 , w_5678 , \3388_b1 );
or ( \3390_b1 , \3296_b1 , \3389_b1 );
not ( \3389_b1 , w_5680 );
and ( \3390_b0 , \3296_b0 , w_5681 );
and ( w_5680 , w_5681 , \3389_b0 );
or ( \3391_b1 , \3295_b1 , w_5682 );
or ( \3391_b0 , \3295_b0 , \3390_b0 );
not ( \3390_b0 , w_5683 );
and ( w_5683 , w_5682 , \3390_b1 );
or ( \3392_b1 , \2923_A[16]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5684 );
and ( \3392_b0 , \2923_A[16]_b0 , w_5685 );
and ( w_5684 , w_5685 , \2997_B[5]_b0 );
or ( \3393_b1 , \3391_b1 , \3392_b1 );
not ( \3392_b1 , w_5686 );
and ( \3393_b0 , \3391_b0 , w_5687 );
and ( w_5686 , w_5687 , \3392_b0 );
or ( \3394_b1 , \3391_b1 , \3392_b1 );
xor ( \3394_b0 , \3391_b0 , w_5688 );
not ( w_5688 , w_5689 );
and ( w_5689 , \3392_b1 , \3392_b0 );
or ( \3395_b1 , \3296_b1 , \3389_b1 );
xor ( \3395_b0 , \3296_b0 , w_5690 );
not ( w_5690 , w_5691 );
and ( w_5691 , \3389_b1 , \3389_b0 );
or ( \3396_b1 , \2927_A[15]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5692 );
and ( \3396_b0 , \2927_A[15]_b0 , w_5693 );
and ( w_5692 , w_5693 , \2997_B[5]_b0 );
or ( \3397_b1 , \3395_b1 , \3396_b1 );
not ( \3396_b1 , w_5694 );
and ( \3397_b0 , \3395_b0 , w_5695 );
and ( w_5694 , w_5695 , \3396_b0 );
or ( \3398_b1 , \3395_b1 , \3396_b1 );
xor ( \3398_b0 , \3395_b0 , w_5696 );
not ( w_5696 , w_5697 );
and ( w_5697 , \3396_b1 , \3396_b0 );
or ( \3399_b1 , \3300_b1 , \3387_b1 );
xor ( \3399_b0 , \3300_b0 , w_5698 );
not ( w_5698 , w_5699 );
and ( w_5699 , \3387_b1 , \3387_b0 );
or ( \3400_b1 , \2931_A[14]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5700 );
and ( \3400_b0 , \2931_A[14]_b0 , w_5701 );
and ( w_5700 , w_5701 , \2997_B[5]_b0 );
or ( \3401_b1 , \3399_b1 , \3400_b1 );
not ( \3400_b1 , w_5702 );
and ( \3401_b0 , \3399_b0 , w_5703 );
and ( w_5702 , w_5703 , \3400_b0 );
or ( \3402_b1 , \3399_b1 , \3400_b1 );
xor ( \3402_b0 , \3399_b0 , w_5704 );
not ( w_5704 , w_5705 );
and ( w_5705 , \3400_b1 , \3400_b0 );
or ( \3403_b1 , \3304_b1 , \3385_b1 );
xor ( \3403_b0 , \3304_b0 , w_5706 );
not ( w_5706 , w_5707 );
and ( w_5707 , \3385_b1 , \3385_b0 );
or ( \3404_b1 , \2935_A[13]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5708 );
and ( \3404_b0 , \2935_A[13]_b0 , w_5709 );
and ( w_5708 , w_5709 , \2997_B[5]_b0 );
or ( \3405_b1 , \3403_b1 , \3404_b1 );
not ( \3404_b1 , w_5710 );
and ( \3405_b0 , \3403_b0 , w_5711 );
and ( w_5710 , w_5711 , \3404_b0 );
or ( \3406_b1 , \3403_b1 , \3404_b1 );
xor ( \3406_b0 , \3403_b0 , w_5712 );
not ( w_5712 , w_5713 );
and ( w_5713 , \3404_b1 , \3404_b0 );
or ( \3407_b1 , \3308_b1 , \3383_b1 );
xor ( \3407_b0 , \3308_b0 , w_5714 );
not ( w_5714 , w_5715 );
and ( w_5715 , \3383_b1 , \3383_b0 );
or ( \3408_b1 , \2939_A[12]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5716 );
and ( \3408_b0 , \2939_A[12]_b0 , w_5717 );
and ( w_5716 , w_5717 , \2997_B[5]_b0 );
or ( \3409_b1 , \3407_b1 , \3408_b1 );
not ( \3408_b1 , w_5718 );
and ( \3409_b0 , \3407_b0 , w_5719 );
and ( w_5718 , w_5719 , \3408_b0 );
or ( \3410_b1 , \3407_b1 , \3408_b1 );
xor ( \3410_b0 , \3407_b0 , w_5720 );
not ( w_5720 , w_5721 );
and ( w_5721 , \3408_b1 , \3408_b0 );
or ( \3411_b1 , \3312_b1 , \3381_b1 );
xor ( \3411_b0 , \3312_b0 , w_5722 );
not ( w_5722 , w_5723 );
and ( w_5723 , \3381_b1 , \3381_b0 );
or ( \3412_b1 , \2943_A[11]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5724 );
and ( \3412_b0 , \2943_A[11]_b0 , w_5725 );
and ( w_5724 , w_5725 , \2997_B[5]_b0 );
or ( \3413_b1 , \3411_b1 , \3412_b1 );
not ( \3412_b1 , w_5726 );
and ( \3413_b0 , \3411_b0 , w_5727 );
and ( w_5726 , w_5727 , \3412_b0 );
or ( \3414_b1 , \3411_b1 , \3412_b1 );
xor ( \3414_b0 , \3411_b0 , w_5728 );
not ( w_5728 , w_5729 );
and ( w_5729 , \3412_b1 , \3412_b0 );
or ( \3415_b1 , \3316_b1 , \3379_b1 );
xor ( \3415_b0 , \3316_b0 , w_5730 );
not ( w_5730 , w_5731 );
and ( w_5731 , \3379_b1 , \3379_b0 );
or ( \3416_b1 , \2947_A[10]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5732 );
and ( \3416_b0 , \2947_A[10]_b0 , w_5733 );
and ( w_5732 , w_5733 , \2997_B[5]_b0 );
or ( \3417_b1 , \3415_b1 , \3416_b1 );
not ( \3416_b1 , w_5734 );
and ( \3417_b0 , \3415_b0 , w_5735 );
and ( w_5734 , w_5735 , \3416_b0 );
or ( \3418_b1 , \3415_b1 , \3416_b1 );
xor ( \3418_b0 , \3415_b0 , w_5736 );
not ( w_5736 , w_5737 );
and ( w_5737 , \3416_b1 , \3416_b0 );
or ( \3419_b1 , \3320_b1 , \3377_b1 );
xor ( \3419_b0 , \3320_b0 , w_5738 );
not ( w_5738 , w_5739 );
and ( w_5739 , \3377_b1 , \3377_b0 );
or ( \3420_b1 , \2951_A[9]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5740 );
and ( \3420_b0 , \2951_A[9]_b0 , w_5741 );
and ( w_5740 , w_5741 , \2997_B[5]_b0 );
or ( \3421_b1 , \3419_b1 , \3420_b1 );
not ( \3420_b1 , w_5742 );
and ( \3421_b0 , \3419_b0 , w_5743 );
and ( w_5742 , w_5743 , \3420_b0 );
or ( \3422_b1 , \3419_b1 , \3420_b1 );
xor ( \3422_b0 , \3419_b0 , w_5744 );
not ( w_5744 , w_5745 );
and ( w_5745 , \3420_b1 , \3420_b0 );
or ( \3423_b1 , \3324_b1 , \3375_b1 );
xor ( \3423_b0 , \3324_b0 , w_5746 );
not ( w_5746 , w_5747 );
and ( w_5747 , \3375_b1 , \3375_b0 );
or ( \3424_b1 , \2955_A[8]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5748 );
and ( \3424_b0 , \2955_A[8]_b0 , w_5749 );
and ( w_5748 , w_5749 , \2997_B[5]_b0 );
or ( \3425_b1 , \3423_b1 , \3424_b1 );
not ( \3424_b1 , w_5750 );
and ( \3425_b0 , \3423_b0 , w_5751 );
and ( w_5750 , w_5751 , \3424_b0 );
or ( \3426_b1 , \3423_b1 , \3424_b1 );
xor ( \3426_b0 , \3423_b0 , w_5752 );
not ( w_5752 , w_5753 );
and ( w_5753 , \3424_b1 , \3424_b0 );
or ( \3427_b1 , \3328_b1 , \3373_b1 );
xor ( \3427_b0 , \3328_b0 , w_5754 );
not ( w_5754 , w_5755 );
and ( w_5755 , \3373_b1 , \3373_b0 );
or ( \3428_b1 , \2959_A[7]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5756 );
and ( \3428_b0 , \2959_A[7]_b0 , w_5757 );
and ( w_5756 , w_5757 , \2997_B[5]_b0 );
or ( \3429_b1 , \3427_b1 , \3428_b1 );
not ( \3428_b1 , w_5758 );
and ( \3429_b0 , \3427_b0 , w_5759 );
and ( w_5758 , w_5759 , \3428_b0 );
or ( \3430_b1 , \3427_b1 , \3428_b1 );
xor ( \3430_b0 , \3427_b0 , w_5760 );
not ( w_5760 , w_5761 );
and ( w_5761 , \3428_b1 , \3428_b0 );
or ( \3431_b1 , \3332_b1 , \3371_b1 );
xor ( \3431_b0 , \3332_b0 , w_5762 );
not ( w_5762 , w_5763 );
and ( w_5763 , \3371_b1 , \3371_b0 );
or ( \3432_b1 , \2963_A[6]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5764 );
and ( \3432_b0 , \2963_A[6]_b0 , w_5765 );
and ( w_5764 , w_5765 , \2997_B[5]_b0 );
or ( \3433_b1 , \3431_b1 , \3432_b1 );
not ( \3432_b1 , w_5766 );
and ( \3433_b0 , \3431_b0 , w_5767 );
and ( w_5766 , w_5767 , \3432_b0 );
or ( \3434_b1 , \3431_b1 , \3432_b1 );
xor ( \3434_b0 , \3431_b0 , w_5768 );
not ( w_5768 , w_5769 );
and ( w_5769 , \3432_b1 , \3432_b0 );
or ( \3435_b1 , \3336_b1 , \3369_b1 );
xor ( \3435_b0 , \3336_b0 , w_5770 );
not ( w_5770 , w_5771 );
and ( w_5771 , \3369_b1 , \3369_b0 );
or ( \3436_b1 , \2967_A[5]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5772 );
and ( \3436_b0 , \2967_A[5]_b0 , w_5773 );
and ( w_5772 , w_5773 , \2997_B[5]_b0 );
or ( \3437_b1 , \3435_b1 , \3436_b1 );
not ( \3436_b1 , w_5774 );
and ( \3437_b0 , \3435_b0 , w_5775 );
and ( w_5774 , w_5775 , \3436_b0 );
or ( \3438_b1 , \3435_b1 , \3436_b1 );
xor ( \3438_b0 , \3435_b0 , w_5776 );
not ( w_5776 , w_5777 );
and ( w_5777 , \3436_b1 , \3436_b0 );
or ( \3439_b1 , \3340_b1 , \3367_b1 );
xor ( \3439_b0 , \3340_b0 , w_5778 );
not ( w_5778 , w_5779 );
and ( w_5779 , \3367_b1 , \3367_b0 );
or ( \3440_b1 , \2971_A[4]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5780 );
and ( \3440_b0 , \2971_A[4]_b0 , w_5781 );
and ( w_5780 , w_5781 , \2997_B[5]_b0 );
or ( \3441_b1 , \3439_b1 , \3440_b1 );
not ( \3440_b1 , w_5782 );
and ( \3441_b0 , \3439_b0 , w_5783 );
and ( w_5782 , w_5783 , \3440_b0 );
or ( \3442_b1 , \3439_b1 , \3440_b1 );
xor ( \3442_b0 , \3439_b0 , w_5784 );
not ( w_5784 , w_5785 );
and ( w_5785 , \3440_b1 , \3440_b0 );
or ( \3443_b1 , \3344_b1 , \3365_b1 );
xor ( \3443_b0 , \3344_b0 , w_5786 );
not ( w_5786 , w_5787 );
and ( w_5787 , \3365_b1 , \3365_b0 );
or ( \3444_b1 , \2975_A[3]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5788 );
and ( \3444_b0 , \2975_A[3]_b0 , w_5789 );
and ( w_5788 , w_5789 , \2997_B[5]_b0 );
or ( \3445_b1 , \3443_b1 , \3444_b1 );
not ( \3444_b1 , w_5790 );
and ( \3445_b0 , \3443_b0 , w_5791 );
and ( w_5790 , w_5791 , \3444_b0 );
or ( \3446_b1 , \3443_b1 , \3444_b1 );
xor ( \3446_b0 , \3443_b0 , w_5792 );
not ( w_5792 , w_5793 );
and ( w_5793 , \3444_b1 , \3444_b0 );
or ( \3447_b1 , \3348_b1 , \3363_b1 );
xor ( \3447_b0 , \3348_b0 , w_5794 );
not ( w_5794 , w_5795 );
and ( w_5795 , \3363_b1 , \3363_b0 );
or ( \3448_b1 , \2979_A[2]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5796 );
and ( \3448_b0 , \2979_A[2]_b0 , w_5797 );
and ( w_5796 , w_5797 , \2997_B[5]_b0 );
or ( \3449_b1 , \3447_b1 , \3448_b1 );
not ( \3448_b1 , w_5798 );
and ( \3449_b0 , \3447_b0 , w_5799 );
and ( w_5798 , w_5799 , \3448_b0 );
or ( \3450_b1 , \3447_b1 , \3448_b1 );
xor ( \3450_b0 , \3447_b0 , w_5800 );
not ( w_5800 , w_5801 );
and ( w_5801 , \3448_b1 , \3448_b0 );
or ( \3451_b1 , \3352_b1 , \3361_b1 );
xor ( \3451_b0 , \3352_b0 , w_5802 );
not ( w_5802 , w_5803 );
and ( w_5803 , \3361_b1 , \3361_b0 );
or ( \3452_b1 , \2983_A[1]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5804 );
and ( \3452_b0 , \2983_A[1]_b0 , w_5805 );
and ( w_5804 , w_5805 , \2997_B[5]_b0 );
or ( \3453_b1 , \3451_b1 , \3452_b1 );
not ( \3452_b1 , w_5806 );
and ( \3453_b0 , \3451_b0 , w_5807 );
and ( w_5806 , w_5807 , \3452_b0 );
or ( \3454_b1 , \3451_b1 , \3452_b1 );
xor ( \3454_b0 , \3451_b0 , w_5808 );
not ( w_5808 , w_5809 );
and ( w_5809 , \3452_b1 , \3452_b0 );
or ( \3455_b1 , \3356_b1 , \3359_b1 );
xor ( \3455_b0 , \3356_b0 , w_5810 );
not ( w_5810 , w_5811 );
and ( w_5811 , \3359_b1 , \3359_b0 );
or ( \3456_b1 , \2986_A[0]_b1 , \2997_B[5]_b1 );
not ( \2997_B[5]_b1 , w_5812 );
and ( \3456_b0 , \2986_A[0]_b0 , w_5813 );
and ( w_5812 , w_5813 , \2997_B[5]_b0 );
or ( \3457_b1 , \3455_b1 , \3456_b1 );
not ( \3456_b1 , w_5814 );
and ( \3457_b0 , \3455_b0 , w_5815 );
and ( w_5814 , w_5815 , \3456_b0 );
or ( \3458_b1 , \3454_b1 , \3457_b1 );
not ( \3457_b1 , w_5816 );
and ( \3458_b0 , \3454_b0 , w_5817 );
and ( w_5816 , w_5817 , \3457_b0 );
or ( \3459_b1 , \3453_b1 , w_5818 );
or ( \3459_b0 , \3453_b0 , \3458_b0 );
not ( \3458_b0 , w_5819 );
and ( w_5819 , w_5818 , \3458_b1 );
or ( \3460_b1 , \3450_b1 , \3459_b1 );
not ( \3459_b1 , w_5820 );
and ( \3460_b0 , \3450_b0 , w_5821 );
and ( w_5820 , w_5821 , \3459_b0 );
or ( \3461_b1 , \3449_b1 , w_5822 );
or ( \3461_b0 , \3449_b0 , \3460_b0 );
not ( \3460_b0 , w_5823 );
and ( w_5823 , w_5822 , \3460_b1 );
or ( \3462_b1 , \3446_b1 , \3461_b1 );
not ( \3461_b1 , w_5824 );
and ( \3462_b0 , \3446_b0 , w_5825 );
and ( w_5824 , w_5825 , \3461_b0 );
or ( \3463_b1 , \3445_b1 , w_5826 );
or ( \3463_b0 , \3445_b0 , \3462_b0 );
not ( \3462_b0 , w_5827 );
and ( w_5827 , w_5826 , \3462_b1 );
or ( \3464_b1 , \3442_b1 , \3463_b1 );
not ( \3463_b1 , w_5828 );
and ( \3464_b0 , \3442_b0 , w_5829 );
and ( w_5828 , w_5829 , \3463_b0 );
or ( \3465_b1 , \3441_b1 , w_5830 );
or ( \3465_b0 , \3441_b0 , \3464_b0 );
not ( \3464_b0 , w_5831 );
and ( w_5831 , w_5830 , \3464_b1 );
or ( \3466_b1 , \3438_b1 , \3465_b1 );
not ( \3465_b1 , w_5832 );
and ( \3466_b0 , \3438_b0 , w_5833 );
and ( w_5832 , w_5833 , \3465_b0 );
or ( \3467_b1 , \3437_b1 , w_5834 );
or ( \3467_b0 , \3437_b0 , \3466_b0 );
not ( \3466_b0 , w_5835 );
and ( w_5835 , w_5834 , \3466_b1 );
or ( \3468_b1 , \3434_b1 , \3467_b1 );
not ( \3467_b1 , w_5836 );
and ( \3468_b0 , \3434_b0 , w_5837 );
and ( w_5836 , w_5837 , \3467_b0 );
or ( \3469_b1 , \3433_b1 , w_5838 );
or ( \3469_b0 , \3433_b0 , \3468_b0 );
not ( \3468_b0 , w_5839 );
and ( w_5839 , w_5838 , \3468_b1 );
or ( \3470_b1 , \3430_b1 , \3469_b1 );
not ( \3469_b1 , w_5840 );
and ( \3470_b0 , \3430_b0 , w_5841 );
and ( w_5840 , w_5841 , \3469_b0 );
or ( \3471_b1 , \3429_b1 , w_5842 );
or ( \3471_b0 , \3429_b0 , \3470_b0 );
not ( \3470_b0 , w_5843 );
and ( w_5843 , w_5842 , \3470_b1 );
or ( \3472_b1 , \3426_b1 , \3471_b1 );
not ( \3471_b1 , w_5844 );
and ( \3472_b0 , \3426_b0 , w_5845 );
and ( w_5844 , w_5845 , \3471_b0 );
or ( \3473_b1 , \3425_b1 , w_5846 );
or ( \3473_b0 , \3425_b0 , \3472_b0 );
not ( \3472_b0 , w_5847 );
and ( w_5847 , w_5846 , \3472_b1 );
or ( \3474_b1 , \3422_b1 , \3473_b1 );
not ( \3473_b1 , w_5848 );
and ( \3474_b0 , \3422_b0 , w_5849 );
and ( w_5848 , w_5849 , \3473_b0 );
or ( \3475_b1 , \3421_b1 , w_5850 );
or ( \3475_b0 , \3421_b0 , \3474_b0 );
not ( \3474_b0 , w_5851 );
and ( w_5851 , w_5850 , \3474_b1 );
or ( \3476_b1 , \3418_b1 , \3475_b1 );
not ( \3475_b1 , w_5852 );
and ( \3476_b0 , \3418_b0 , w_5853 );
and ( w_5852 , w_5853 , \3475_b0 );
or ( \3477_b1 , \3417_b1 , w_5854 );
or ( \3477_b0 , \3417_b0 , \3476_b0 );
not ( \3476_b0 , w_5855 );
and ( w_5855 , w_5854 , \3476_b1 );
or ( \3478_b1 , \3414_b1 , \3477_b1 );
not ( \3477_b1 , w_5856 );
and ( \3478_b0 , \3414_b0 , w_5857 );
and ( w_5856 , w_5857 , \3477_b0 );
or ( \3479_b1 , \3413_b1 , w_5858 );
or ( \3479_b0 , \3413_b0 , \3478_b0 );
not ( \3478_b0 , w_5859 );
and ( w_5859 , w_5858 , \3478_b1 );
or ( \3480_b1 , \3410_b1 , \3479_b1 );
not ( \3479_b1 , w_5860 );
and ( \3480_b0 , \3410_b0 , w_5861 );
and ( w_5860 , w_5861 , \3479_b0 );
or ( \3481_b1 , \3409_b1 , w_5862 );
or ( \3481_b0 , \3409_b0 , \3480_b0 );
not ( \3480_b0 , w_5863 );
and ( w_5863 , w_5862 , \3480_b1 );
or ( \3482_b1 , \3406_b1 , \3481_b1 );
not ( \3481_b1 , w_5864 );
and ( \3482_b0 , \3406_b0 , w_5865 );
and ( w_5864 , w_5865 , \3481_b0 );
or ( \3483_b1 , \3405_b1 , w_5866 );
or ( \3483_b0 , \3405_b0 , \3482_b0 );
not ( \3482_b0 , w_5867 );
and ( w_5867 , w_5866 , \3482_b1 );
or ( \3484_b1 , \3402_b1 , \3483_b1 );
not ( \3483_b1 , w_5868 );
and ( \3484_b0 , \3402_b0 , w_5869 );
and ( w_5868 , w_5869 , \3483_b0 );
or ( \3485_b1 , \3401_b1 , w_5870 );
or ( \3485_b0 , \3401_b0 , \3484_b0 );
not ( \3484_b0 , w_5871 );
and ( w_5871 , w_5870 , \3484_b1 );
or ( \3486_b1 , \3398_b1 , \3485_b1 );
not ( \3485_b1 , w_5872 );
and ( \3486_b0 , \3398_b0 , w_5873 );
and ( w_5872 , w_5873 , \3485_b0 );
or ( \3487_b1 , \3397_b1 , w_5874 );
or ( \3487_b0 , \3397_b0 , \3486_b0 );
not ( \3486_b0 , w_5875 );
and ( w_5875 , w_5874 , \3486_b1 );
or ( \3488_b1 , \3394_b1 , \3487_b1 );
not ( \3487_b1 , w_5876 );
and ( \3488_b0 , \3394_b0 , w_5877 );
and ( w_5876 , w_5877 , \3487_b0 );
or ( \3489_b1 , \3393_b1 , w_5878 );
or ( \3489_b0 , \3393_b0 , \3488_b0 );
not ( \3488_b0 , w_5879 );
and ( w_5879 , w_5878 , \3488_b1 );
or ( \3490_b1 , \2923_A[16]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5880 );
and ( \3490_b0 , \2923_A[16]_b0 , w_5881 );
and ( w_5880 , w_5881 , \2996_B[6]_b0 );
or ( \3491_b1 , \3489_b1 , \3490_b1 );
not ( \3490_b1 , w_5882 );
and ( \3491_b0 , \3489_b0 , w_5883 );
and ( w_5882 , w_5883 , \3490_b0 );
or ( \3492_b1 , \3489_b1 , \3490_b1 );
xor ( \3492_b0 , \3489_b0 , w_5884 );
not ( w_5884 , w_5885 );
and ( w_5885 , \3490_b1 , \3490_b0 );
or ( \3493_b1 , \3394_b1 , \3487_b1 );
xor ( \3493_b0 , \3394_b0 , w_5886 );
not ( w_5886 , w_5887 );
and ( w_5887 , \3487_b1 , \3487_b0 );
or ( \3494_b1 , \2927_A[15]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5888 );
and ( \3494_b0 , \2927_A[15]_b0 , w_5889 );
and ( w_5888 , w_5889 , \2996_B[6]_b0 );
or ( \3495_b1 , \3493_b1 , \3494_b1 );
not ( \3494_b1 , w_5890 );
and ( \3495_b0 , \3493_b0 , w_5891 );
and ( w_5890 , w_5891 , \3494_b0 );
or ( \3496_b1 , \3493_b1 , \3494_b1 );
xor ( \3496_b0 , \3493_b0 , w_5892 );
not ( w_5892 , w_5893 );
and ( w_5893 , \3494_b1 , \3494_b0 );
or ( \3497_b1 , \3398_b1 , \3485_b1 );
xor ( \3497_b0 , \3398_b0 , w_5894 );
not ( w_5894 , w_5895 );
and ( w_5895 , \3485_b1 , \3485_b0 );
or ( \3498_b1 , \2931_A[14]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5896 );
and ( \3498_b0 , \2931_A[14]_b0 , w_5897 );
and ( w_5896 , w_5897 , \2996_B[6]_b0 );
or ( \3499_b1 , \3497_b1 , \3498_b1 );
not ( \3498_b1 , w_5898 );
and ( \3499_b0 , \3497_b0 , w_5899 );
and ( w_5898 , w_5899 , \3498_b0 );
or ( \3500_b1 , \3497_b1 , \3498_b1 );
xor ( \3500_b0 , \3497_b0 , w_5900 );
not ( w_5900 , w_5901 );
and ( w_5901 , \3498_b1 , \3498_b0 );
or ( \3501_b1 , \3402_b1 , \3483_b1 );
xor ( \3501_b0 , \3402_b0 , w_5902 );
not ( w_5902 , w_5903 );
and ( w_5903 , \3483_b1 , \3483_b0 );
or ( \3502_b1 , \2935_A[13]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5904 );
and ( \3502_b0 , \2935_A[13]_b0 , w_5905 );
and ( w_5904 , w_5905 , \2996_B[6]_b0 );
or ( \3503_b1 , \3501_b1 , \3502_b1 );
not ( \3502_b1 , w_5906 );
and ( \3503_b0 , \3501_b0 , w_5907 );
and ( w_5906 , w_5907 , \3502_b0 );
or ( \3504_b1 , \3501_b1 , \3502_b1 );
xor ( \3504_b0 , \3501_b0 , w_5908 );
not ( w_5908 , w_5909 );
and ( w_5909 , \3502_b1 , \3502_b0 );
or ( \3505_b1 , \3406_b1 , \3481_b1 );
xor ( \3505_b0 , \3406_b0 , w_5910 );
not ( w_5910 , w_5911 );
and ( w_5911 , \3481_b1 , \3481_b0 );
or ( \3506_b1 , \2939_A[12]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5912 );
and ( \3506_b0 , \2939_A[12]_b0 , w_5913 );
and ( w_5912 , w_5913 , \2996_B[6]_b0 );
or ( \3507_b1 , \3505_b1 , \3506_b1 );
not ( \3506_b1 , w_5914 );
and ( \3507_b0 , \3505_b0 , w_5915 );
and ( w_5914 , w_5915 , \3506_b0 );
or ( \3508_b1 , \3505_b1 , \3506_b1 );
xor ( \3508_b0 , \3505_b0 , w_5916 );
not ( w_5916 , w_5917 );
and ( w_5917 , \3506_b1 , \3506_b0 );
or ( \3509_b1 , \3410_b1 , \3479_b1 );
xor ( \3509_b0 , \3410_b0 , w_5918 );
not ( w_5918 , w_5919 );
and ( w_5919 , \3479_b1 , \3479_b0 );
or ( \3510_b1 , \2943_A[11]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5920 );
and ( \3510_b0 , \2943_A[11]_b0 , w_5921 );
and ( w_5920 , w_5921 , \2996_B[6]_b0 );
or ( \3511_b1 , \3509_b1 , \3510_b1 );
not ( \3510_b1 , w_5922 );
and ( \3511_b0 , \3509_b0 , w_5923 );
and ( w_5922 , w_5923 , \3510_b0 );
or ( \3512_b1 , \3509_b1 , \3510_b1 );
xor ( \3512_b0 , \3509_b0 , w_5924 );
not ( w_5924 , w_5925 );
and ( w_5925 , \3510_b1 , \3510_b0 );
or ( \3513_b1 , \3414_b1 , \3477_b1 );
xor ( \3513_b0 , \3414_b0 , w_5926 );
not ( w_5926 , w_5927 );
and ( w_5927 , \3477_b1 , \3477_b0 );
or ( \3514_b1 , \2947_A[10]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5928 );
and ( \3514_b0 , \2947_A[10]_b0 , w_5929 );
and ( w_5928 , w_5929 , \2996_B[6]_b0 );
or ( \3515_b1 , \3513_b1 , \3514_b1 );
not ( \3514_b1 , w_5930 );
and ( \3515_b0 , \3513_b0 , w_5931 );
and ( w_5930 , w_5931 , \3514_b0 );
or ( \3516_b1 , \3513_b1 , \3514_b1 );
xor ( \3516_b0 , \3513_b0 , w_5932 );
not ( w_5932 , w_5933 );
and ( w_5933 , \3514_b1 , \3514_b0 );
or ( \3517_b1 , \3418_b1 , \3475_b1 );
xor ( \3517_b0 , \3418_b0 , w_5934 );
not ( w_5934 , w_5935 );
and ( w_5935 , \3475_b1 , \3475_b0 );
or ( \3518_b1 , \2951_A[9]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5936 );
and ( \3518_b0 , \2951_A[9]_b0 , w_5937 );
and ( w_5936 , w_5937 , \2996_B[6]_b0 );
or ( \3519_b1 , \3517_b1 , \3518_b1 );
not ( \3518_b1 , w_5938 );
and ( \3519_b0 , \3517_b0 , w_5939 );
and ( w_5938 , w_5939 , \3518_b0 );
or ( \3520_b1 , \3517_b1 , \3518_b1 );
xor ( \3520_b0 , \3517_b0 , w_5940 );
not ( w_5940 , w_5941 );
and ( w_5941 , \3518_b1 , \3518_b0 );
or ( \3521_b1 , \3422_b1 , \3473_b1 );
xor ( \3521_b0 , \3422_b0 , w_5942 );
not ( w_5942 , w_5943 );
and ( w_5943 , \3473_b1 , \3473_b0 );
or ( \3522_b1 , \2955_A[8]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5944 );
and ( \3522_b0 , \2955_A[8]_b0 , w_5945 );
and ( w_5944 , w_5945 , \2996_B[6]_b0 );
or ( \3523_b1 , \3521_b1 , \3522_b1 );
not ( \3522_b1 , w_5946 );
and ( \3523_b0 , \3521_b0 , w_5947 );
and ( w_5946 , w_5947 , \3522_b0 );
or ( \3524_b1 , \3521_b1 , \3522_b1 );
xor ( \3524_b0 , \3521_b0 , w_5948 );
not ( w_5948 , w_5949 );
and ( w_5949 , \3522_b1 , \3522_b0 );
or ( \3525_b1 , \3426_b1 , \3471_b1 );
xor ( \3525_b0 , \3426_b0 , w_5950 );
not ( w_5950 , w_5951 );
and ( w_5951 , \3471_b1 , \3471_b0 );
or ( \3526_b1 , \2959_A[7]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5952 );
and ( \3526_b0 , \2959_A[7]_b0 , w_5953 );
and ( w_5952 , w_5953 , \2996_B[6]_b0 );
or ( \3527_b1 , \3525_b1 , \3526_b1 );
not ( \3526_b1 , w_5954 );
and ( \3527_b0 , \3525_b0 , w_5955 );
and ( w_5954 , w_5955 , \3526_b0 );
or ( \3528_b1 , \3525_b1 , \3526_b1 );
xor ( \3528_b0 , \3525_b0 , w_5956 );
not ( w_5956 , w_5957 );
and ( w_5957 , \3526_b1 , \3526_b0 );
or ( \3529_b1 , \3430_b1 , \3469_b1 );
xor ( \3529_b0 , \3430_b0 , w_5958 );
not ( w_5958 , w_5959 );
and ( w_5959 , \3469_b1 , \3469_b0 );
or ( \3530_b1 , \2963_A[6]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5960 );
and ( \3530_b0 , \2963_A[6]_b0 , w_5961 );
and ( w_5960 , w_5961 , \2996_B[6]_b0 );
or ( \3531_b1 , \3529_b1 , \3530_b1 );
not ( \3530_b1 , w_5962 );
and ( \3531_b0 , \3529_b0 , w_5963 );
and ( w_5962 , w_5963 , \3530_b0 );
or ( \3532_b1 , \3529_b1 , \3530_b1 );
xor ( \3532_b0 , \3529_b0 , w_5964 );
not ( w_5964 , w_5965 );
and ( w_5965 , \3530_b1 , \3530_b0 );
or ( \3533_b1 , \3434_b1 , \3467_b1 );
xor ( \3533_b0 , \3434_b0 , w_5966 );
not ( w_5966 , w_5967 );
and ( w_5967 , \3467_b1 , \3467_b0 );
or ( \3534_b1 , \2967_A[5]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5968 );
and ( \3534_b0 , \2967_A[5]_b0 , w_5969 );
and ( w_5968 , w_5969 , \2996_B[6]_b0 );
or ( \3535_b1 , \3533_b1 , \3534_b1 );
not ( \3534_b1 , w_5970 );
and ( \3535_b0 , \3533_b0 , w_5971 );
and ( w_5970 , w_5971 , \3534_b0 );
or ( \3536_b1 , \3533_b1 , \3534_b1 );
xor ( \3536_b0 , \3533_b0 , w_5972 );
not ( w_5972 , w_5973 );
and ( w_5973 , \3534_b1 , \3534_b0 );
or ( \3537_b1 , \3438_b1 , \3465_b1 );
xor ( \3537_b0 , \3438_b0 , w_5974 );
not ( w_5974 , w_5975 );
and ( w_5975 , \3465_b1 , \3465_b0 );
or ( \3538_b1 , \2971_A[4]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5976 );
and ( \3538_b0 , \2971_A[4]_b0 , w_5977 );
and ( w_5976 , w_5977 , \2996_B[6]_b0 );
or ( \3539_b1 , \3537_b1 , \3538_b1 );
not ( \3538_b1 , w_5978 );
and ( \3539_b0 , \3537_b0 , w_5979 );
and ( w_5978 , w_5979 , \3538_b0 );
or ( \3540_b1 , \3537_b1 , \3538_b1 );
xor ( \3540_b0 , \3537_b0 , w_5980 );
not ( w_5980 , w_5981 );
and ( w_5981 , \3538_b1 , \3538_b0 );
or ( \3541_b1 , \3442_b1 , \3463_b1 );
xor ( \3541_b0 , \3442_b0 , w_5982 );
not ( w_5982 , w_5983 );
and ( w_5983 , \3463_b1 , \3463_b0 );
or ( \3542_b1 , \2975_A[3]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5984 );
and ( \3542_b0 , \2975_A[3]_b0 , w_5985 );
and ( w_5984 , w_5985 , \2996_B[6]_b0 );
or ( \3543_b1 , \3541_b1 , \3542_b1 );
not ( \3542_b1 , w_5986 );
and ( \3543_b0 , \3541_b0 , w_5987 );
and ( w_5986 , w_5987 , \3542_b0 );
or ( \3544_b1 , \3541_b1 , \3542_b1 );
xor ( \3544_b0 , \3541_b0 , w_5988 );
not ( w_5988 , w_5989 );
and ( w_5989 , \3542_b1 , \3542_b0 );
or ( \3545_b1 , \3446_b1 , \3461_b1 );
xor ( \3545_b0 , \3446_b0 , w_5990 );
not ( w_5990 , w_5991 );
and ( w_5991 , \3461_b1 , \3461_b0 );
or ( \3546_b1 , \2979_A[2]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_5992 );
and ( \3546_b0 , \2979_A[2]_b0 , w_5993 );
and ( w_5992 , w_5993 , \2996_B[6]_b0 );
or ( \3547_b1 , \3545_b1 , \3546_b1 );
not ( \3546_b1 , w_5994 );
and ( \3547_b0 , \3545_b0 , w_5995 );
and ( w_5994 , w_5995 , \3546_b0 );
or ( \3548_b1 , \3545_b1 , \3546_b1 );
xor ( \3548_b0 , \3545_b0 , w_5996 );
not ( w_5996 , w_5997 );
and ( w_5997 , \3546_b1 , \3546_b0 );
or ( \3549_b1 , \3450_b1 , \3459_b1 );
xor ( \3549_b0 , \3450_b0 , w_5998 );
not ( w_5998 , w_5999 );
and ( w_5999 , \3459_b1 , \3459_b0 );
or ( \3550_b1 , \2983_A[1]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_6000 );
and ( \3550_b0 , \2983_A[1]_b0 , w_6001 );
and ( w_6000 , w_6001 , \2996_B[6]_b0 );
or ( \3551_b1 , \3549_b1 , \3550_b1 );
not ( \3550_b1 , w_6002 );
and ( \3551_b0 , \3549_b0 , w_6003 );
and ( w_6002 , w_6003 , \3550_b0 );
or ( \3552_b1 , \3549_b1 , \3550_b1 );
xor ( \3552_b0 , \3549_b0 , w_6004 );
not ( w_6004 , w_6005 );
and ( w_6005 , \3550_b1 , \3550_b0 );
or ( \3553_b1 , \3454_b1 , \3457_b1 );
xor ( \3553_b0 , \3454_b0 , w_6006 );
not ( w_6006 , w_6007 );
and ( w_6007 , \3457_b1 , \3457_b0 );
or ( \3554_b1 , \2986_A[0]_b1 , \2996_B[6]_b1 );
not ( \2996_B[6]_b1 , w_6008 );
and ( \3554_b0 , \2986_A[0]_b0 , w_6009 );
and ( w_6008 , w_6009 , \2996_B[6]_b0 );
or ( \3555_b1 , \3553_b1 , \3554_b1 );
not ( \3554_b1 , w_6010 );
and ( \3555_b0 , \3553_b0 , w_6011 );
and ( w_6010 , w_6011 , \3554_b0 );
or ( \3556_b1 , \3552_b1 , \3555_b1 );
not ( \3555_b1 , w_6012 );
and ( \3556_b0 , \3552_b0 , w_6013 );
and ( w_6012 , w_6013 , \3555_b0 );
or ( \3557_b1 , \3551_b1 , w_6014 );
or ( \3557_b0 , \3551_b0 , \3556_b0 );
not ( \3556_b0 , w_6015 );
and ( w_6015 , w_6014 , \3556_b1 );
or ( \3558_b1 , \3548_b1 , \3557_b1 );
not ( \3557_b1 , w_6016 );
and ( \3558_b0 , \3548_b0 , w_6017 );
and ( w_6016 , w_6017 , \3557_b0 );
or ( \3559_b1 , \3547_b1 , w_6018 );
or ( \3559_b0 , \3547_b0 , \3558_b0 );
not ( \3558_b0 , w_6019 );
and ( w_6019 , w_6018 , \3558_b1 );
or ( \3560_b1 , \3544_b1 , \3559_b1 );
not ( \3559_b1 , w_6020 );
and ( \3560_b0 , \3544_b0 , w_6021 );
and ( w_6020 , w_6021 , \3559_b0 );
or ( \3561_b1 , \3543_b1 , w_6022 );
or ( \3561_b0 , \3543_b0 , \3560_b0 );
not ( \3560_b0 , w_6023 );
and ( w_6023 , w_6022 , \3560_b1 );
or ( \3562_b1 , \3540_b1 , \3561_b1 );
not ( \3561_b1 , w_6024 );
and ( \3562_b0 , \3540_b0 , w_6025 );
and ( w_6024 , w_6025 , \3561_b0 );
or ( \3563_b1 , \3539_b1 , w_6026 );
or ( \3563_b0 , \3539_b0 , \3562_b0 );
not ( \3562_b0 , w_6027 );
and ( w_6027 , w_6026 , \3562_b1 );
or ( \3564_b1 , \3536_b1 , \3563_b1 );
not ( \3563_b1 , w_6028 );
and ( \3564_b0 , \3536_b0 , w_6029 );
and ( w_6028 , w_6029 , \3563_b0 );
or ( \3565_b1 , \3535_b1 , w_6030 );
or ( \3565_b0 , \3535_b0 , \3564_b0 );
not ( \3564_b0 , w_6031 );
and ( w_6031 , w_6030 , \3564_b1 );
or ( \3566_b1 , \3532_b1 , \3565_b1 );
not ( \3565_b1 , w_6032 );
and ( \3566_b0 , \3532_b0 , w_6033 );
and ( w_6032 , w_6033 , \3565_b0 );
or ( \3567_b1 , \3531_b1 , w_6034 );
or ( \3567_b0 , \3531_b0 , \3566_b0 );
not ( \3566_b0 , w_6035 );
and ( w_6035 , w_6034 , \3566_b1 );
or ( \3568_b1 , \3528_b1 , \3567_b1 );
not ( \3567_b1 , w_6036 );
and ( \3568_b0 , \3528_b0 , w_6037 );
and ( w_6036 , w_6037 , \3567_b0 );
or ( \3569_b1 , \3527_b1 , w_6038 );
or ( \3569_b0 , \3527_b0 , \3568_b0 );
not ( \3568_b0 , w_6039 );
and ( w_6039 , w_6038 , \3568_b1 );
or ( \3570_b1 , \3524_b1 , \3569_b1 );
not ( \3569_b1 , w_6040 );
and ( \3570_b0 , \3524_b0 , w_6041 );
and ( w_6040 , w_6041 , \3569_b0 );
or ( \3571_b1 , \3523_b1 , w_6042 );
or ( \3571_b0 , \3523_b0 , \3570_b0 );
not ( \3570_b0 , w_6043 );
and ( w_6043 , w_6042 , \3570_b1 );
or ( \3572_b1 , \3520_b1 , \3571_b1 );
not ( \3571_b1 , w_6044 );
and ( \3572_b0 , \3520_b0 , w_6045 );
and ( w_6044 , w_6045 , \3571_b0 );
or ( \3573_b1 , \3519_b1 , w_6046 );
or ( \3573_b0 , \3519_b0 , \3572_b0 );
not ( \3572_b0 , w_6047 );
and ( w_6047 , w_6046 , \3572_b1 );
or ( \3574_b1 , \3516_b1 , \3573_b1 );
not ( \3573_b1 , w_6048 );
and ( \3574_b0 , \3516_b0 , w_6049 );
and ( w_6048 , w_6049 , \3573_b0 );
or ( \3575_b1 , \3515_b1 , w_6050 );
or ( \3575_b0 , \3515_b0 , \3574_b0 );
not ( \3574_b0 , w_6051 );
and ( w_6051 , w_6050 , \3574_b1 );
or ( \3576_b1 , \3512_b1 , \3575_b1 );
not ( \3575_b1 , w_6052 );
and ( \3576_b0 , \3512_b0 , w_6053 );
and ( w_6052 , w_6053 , \3575_b0 );
or ( \3577_b1 , \3511_b1 , w_6054 );
or ( \3577_b0 , \3511_b0 , \3576_b0 );
not ( \3576_b0 , w_6055 );
and ( w_6055 , w_6054 , \3576_b1 );
or ( \3578_b1 , \3508_b1 , \3577_b1 );
not ( \3577_b1 , w_6056 );
and ( \3578_b0 , \3508_b0 , w_6057 );
and ( w_6056 , w_6057 , \3577_b0 );
or ( \3579_b1 , \3507_b1 , w_6058 );
or ( \3579_b0 , \3507_b0 , \3578_b0 );
not ( \3578_b0 , w_6059 );
and ( w_6059 , w_6058 , \3578_b1 );
or ( \3580_b1 , \3504_b1 , \3579_b1 );
not ( \3579_b1 , w_6060 );
and ( \3580_b0 , \3504_b0 , w_6061 );
and ( w_6060 , w_6061 , \3579_b0 );
or ( \3581_b1 , \3503_b1 , w_6062 );
or ( \3581_b0 , \3503_b0 , \3580_b0 );
not ( \3580_b0 , w_6063 );
and ( w_6063 , w_6062 , \3580_b1 );
or ( \3582_b1 , \3500_b1 , \3581_b1 );
not ( \3581_b1 , w_6064 );
and ( \3582_b0 , \3500_b0 , w_6065 );
and ( w_6064 , w_6065 , \3581_b0 );
or ( \3583_b1 , \3499_b1 , w_6066 );
or ( \3583_b0 , \3499_b0 , \3582_b0 );
not ( \3582_b0 , w_6067 );
and ( w_6067 , w_6066 , \3582_b1 );
or ( \3584_b1 , \3496_b1 , \3583_b1 );
not ( \3583_b1 , w_6068 );
and ( \3584_b0 , \3496_b0 , w_6069 );
and ( w_6068 , w_6069 , \3583_b0 );
or ( \3585_b1 , \3495_b1 , w_6070 );
or ( \3585_b0 , \3495_b0 , \3584_b0 );
not ( \3584_b0 , w_6071 );
and ( w_6071 , w_6070 , \3584_b1 );
or ( \3586_b1 , \3492_b1 , \3585_b1 );
not ( \3585_b1 , w_6072 );
and ( \3586_b0 , \3492_b0 , w_6073 );
and ( w_6072 , w_6073 , \3585_b0 );
or ( \3587_b1 , \3491_b1 , w_6074 );
or ( \3587_b0 , \3491_b0 , \3586_b0 );
not ( \3586_b0 , w_6075 );
and ( w_6075 , w_6074 , \3586_b1 );
or ( \3588_b1 , \2923_A[16]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6076 );
and ( \3588_b0 , \2923_A[16]_b0 , w_6077 );
and ( w_6076 , w_6077 , \2995_B[7]_b0 );
or ( \3589_b1 , \3587_b1 , \3588_b1 );
not ( \3588_b1 , w_6078 );
and ( \3589_b0 , \3587_b0 , w_6079 );
and ( w_6078 , w_6079 , \3588_b0 );
or ( \3590_b1 , \3587_b1 , \3588_b1 );
xor ( \3590_b0 , \3587_b0 , w_6080 );
not ( w_6080 , w_6081 );
and ( w_6081 , \3588_b1 , \3588_b0 );
or ( \3591_b1 , \3492_b1 , \3585_b1 );
xor ( \3591_b0 , \3492_b0 , w_6082 );
not ( w_6082 , w_6083 );
and ( w_6083 , \3585_b1 , \3585_b0 );
or ( \3592_b1 , \2927_A[15]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6084 );
and ( \3592_b0 , \2927_A[15]_b0 , w_6085 );
and ( w_6084 , w_6085 , \2995_B[7]_b0 );
or ( \3593_b1 , \3591_b1 , \3592_b1 );
not ( \3592_b1 , w_6086 );
and ( \3593_b0 , \3591_b0 , w_6087 );
and ( w_6086 , w_6087 , \3592_b0 );
or ( \3594_b1 , \3591_b1 , \3592_b1 );
xor ( \3594_b0 , \3591_b0 , w_6088 );
not ( w_6088 , w_6089 );
and ( w_6089 , \3592_b1 , \3592_b0 );
or ( \3595_b1 , \3496_b1 , \3583_b1 );
xor ( \3595_b0 , \3496_b0 , w_6090 );
not ( w_6090 , w_6091 );
and ( w_6091 , \3583_b1 , \3583_b0 );
or ( \3596_b1 , \2931_A[14]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6092 );
and ( \3596_b0 , \2931_A[14]_b0 , w_6093 );
and ( w_6092 , w_6093 , \2995_B[7]_b0 );
or ( \3597_b1 , \3595_b1 , \3596_b1 );
not ( \3596_b1 , w_6094 );
and ( \3597_b0 , \3595_b0 , w_6095 );
and ( w_6094 , w_6095 , \3596_b0 );
or ( \3598_b1 , \3595_b1 , \3596_b1 );
xor ( \3598_b0 , \3595_b0 , w_6096 );
not ( w_6096 , w_6097 );
and ( w_6097 , \3596_b1 , \3596_b0 );
or ( \3599_b1 , \3500_b1 , \3581_b1 );
xor ( \3599_b0 , \3500_b0 , w_6098 );
not ( w_6098 , w_6099 );
and ( w_6099 , \3581_b1 , \3581_b0 );
or ( \3600_b1 , \2935_A[13]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6100 );
and ( \3600_b0 , \2935_A[13]_b0 , w_6101 );
and ( w_6100 , w_6101 , \2995_B[7]_b0 );
or ( \3601_b1 , \3599_b1 , \3600_b1 );
not ( \3600_b1 , w_6102 );
and ( \3601_b0 , \3599_b0 , w_6103 );
and ( w_6102 , w_6103 , \3600_b0 );
or ( \3602_b1 , \3599_b1 , \3600_b1 );
xor ( \3602_b0 , \3599_b0 , w_6104 );
not ( w_6104 , w_6105 );
and ( w_6105 , \3600_b1 , \3600_b0 );
or ( \3603_b1 , \3504_b1 , \3579_b1 );
xor ( \3603_b0 , \3504_b0 , w_6106 );
not ( w_6106 , w_6107 );
and ( w_6107 , \3579_b1 , \3579_b0 );
or ( \3604_b1 , \2939_A[12]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6108 );
and ( \3604_b0 , \2939_A[12]_b0 , w_6109 );
and ( w_6108 , w_6109 , \2995_B[7]_b0 );
or ( \3605_b1 , \3603_b1 , \3604_b1 );
not ( \3604_b1 , w_6110 );
and ( \3605_b0 , \3603_b0 , w_6111 );
and ( w_6110 , w_6111 , \3604_b0 );
or ( \3606_b1 , \3603_b1 , \3604_b1 );
xor ( \3606_b0 , \3603_b0 , w_6112 );
not ( w_6112 , w_6113 );
and ( w_6113 , \3604_b1 , \3604_b0 );
or ( \3607_b1 , \3508_b1 , \3577_b1 );
xor ( \3607_b0 , \3508_b0 , w_6114 );
not ( w_6114 , w_6115 );
and ( w_6115 , \3577_b1 , \3577_b0 );
or ( \3608_b1 , \2943_A[11]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6116 );
and ( \3608_b0 , \2943_A[11]_b0 , w_6117 );
and ( w_6116 , w_6117 , \2995_B[7]_b0 );
or ( \3609_b1 , \3607_b1 , \3608_b1 );
not ( \3608_b1 , w_6118 );
and ( \3609_b0 , \3607_b0 , w_6119 );
and ( w_6118 , w_6119 , \3608_b0 );
or ( \3610_b1 , \3607_b1 , \3608_b1 );
xor ( \3610_b0 , \3607_b0 , w_6120 );
not ( w_6120 , w_6121 );
and ( w_6121 , \3608_b1 , \3608_b0 );
or ( \3611_b1 , \3512_b1 , \3575_b1 );
xor ( \3611_b0 , \3512_b0 , w_6122 );
not ( w_6122 , w_6123 );
and ( w_6123 , \3575_b1 , \3575_b0 );
or ( \3612_b1 , \2947_A[10]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6124 );
and ( \3612_b0 , \2947_A[10]_b0 , w_6125 );
and ( w_6124 , w_6125 , \2995_B[7]_b0 );
or ( \3613_b1 , \3611_b1 , \3612_b1 );
not ( \3612_b1 , w_6126 );
and ( \3613_b0 , \3611_b0 , w_6127 );
and ( w_6126 , w_6127 , \3612_b0 );
or ( \3614_b1 , \3611_b1 , \3612_b1 );
xor ( \3614_b0 , \3611_b0 , w_6128 );
not ( w_6128 , w_6129 );
and ( w_6129 , \3612_b1 , \3612_b0 );
or ( \3615_b1 , \3516_b1 , \3573_b1 );
xor ( \3615_b0 , \3516_b0 , w_6130 );
not ( w_6130 , w_6131 );
and ( w_6131 , \3573_b1 , \3573_b0 );
or ( \3616_b1 , \2951_A[9]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6132 );
and ( \3616_b0 , \2951_A[9]_b0 , w_6133 );
and ( w_6132 , w_6133 , \2995_B[7]_b0 );
or ( \3617_b1 , \3615_b1 , \3616_b1 );
not ( \3616_b1 , w_6134 );
and ( \3617_b0 , \3615_b0 , w_6135 );
and ( w_6134 , w_6135 , \3616_b0 );
or ( \3618_b1 , \3615_b1 , \3616_b1 );
xor ( \3618_b0 , \3615_b0 , w_6136 );
not ( w_6136 , w_6137 );
and ( w_6137 , \3616_b1 , \3616_b0 );
or ( \3619_b1 , \3520_b1 , \3571_b1 );
xor ( \3619_b0 , \3520_b0 , w_6138 );
not ( w_6138 , w_6139 );
and ( w_6139 , \3571_b1 , \3571_b0 );
or ( \3620_b1 , \2955_A[8]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6140 );
and ( \3620_b0 , \2955_A[8]_b0 , w_6141 );
and ( w_6140 , w_6141 , \2995_B[7]_b0 );
or ( \3621_b1 , \3619_b1 , \3620_b1 );
not ( \3620_b1 , w_6142 );
and ( \3621_b0 , \3619_b0 , w_6143 );
and ( w_6142 , w_6143 , \3620_b0 );
or ( \3622_b1 , \3619_b1 , \3620_b1 );
xor ( \3622_b0 , \3619_b0 , w_6144 );
not ( w_6144 , w_6145 );
and ( w_6145 , \3620_b1 , \3620_b0 );
or ( \3623_b1 , \3524_b1 , \3569_b1 );
xor ( \3623_b0 , \3524_b0 , w_6146 );
not ( w_6146 , w_6147 );
and ( w_6147 , \3569_b1 , \3569_b0 );
or ( \3624_b1 , \2959_A[7]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6148 );
and ( \3624_b0 , \2959_A[7]_b0 , w_6149 );
and ( w_6148 , w_6149 , \2995_B[7]_b0 );
or ( \3625_b1 , \3623_b1 , \3624_b1 );
not ( \3624_b1 , w_6150 );
and ( \3625_b0 , \3623_b0 , w_6151 );
and ( w_6150 , w_6151 , \3624_b0 );
or ( \3626_b1 , \3623_b1 , \3624_b1 );
xor ( \3626_b0 , \3623_b0 , w_6152 );
not ( w_6152 , w_6153 );
and ( w_6153 , \3624_b1 , \3624_b0 );
or ( \3627_b1 , \3528_b1 , \3567_b1 );
xor ( \3627_b0 , \3528_b0 , w_6154 );
not ( w_6154 , w_6155 );
and ( w_6155 , \3567_b1 , \3567_b0 );
or ( \3628_b1 , \2963_A[6]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6156 );
and ( \3628_b0 , \2963_A[6]_b0 , w_6157 );
and ( w_6156 , w_6157 , \2995_B[7]_b0 );
or ( \3629_b1 , \3627_b1 , \3628_b1 );
not ( \3628_b1 , w_6158 );
and ( \3629_b0 , \3627_b0 , w_6159 );
and ( w_6158 , w_6159 , \3628_b0 );
or ( \3630_b1 , \3627_b1 , \3628_b1 );
xor ( \3630_b0 , \3627_b0 , w_6160 );
not ( w_6160 , w_6161 );
and ( w_6161 , \3628_b1 , \3628_b0 );
or ( \3631_b1 , \3532_b1 , \3565_b1 );
xor ( \3631_b0 , \3532_b0 , w_6162 );
not ( w_6162 , w_6163 );
and ( w_6163 , \3565_b1 , \3565_b0 );
or ( \3632_b1 , \2967_A[5]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6164 );
and ( \3632_b0 , \2967_A[5]_b0 , w_6165 );
and ( w_6164 , w_6165 , \2995_B[7]_b0 );
or ( \3633_b1 , \3631_b1 , \3632_b1 );
not ( \3632_b1 , w_6166 );
and ( \3633_b0 , \3631_b0 , w_6167 );
and ( w_6166 , w_6167 , \3632_b0 );
or ( \3634_b1 , \3631_b1 , \3632_b1 );
xor ( \3634_b0 , \3631_b0 , w_6168 );
not ( w_6168 , w_6169 );
and ( w_6169 , \3632_b1 , \3632_b0 );
or ( \3635_b1 , \3536_b1 , \3563_b1 );
xor ( \3635_b0 , \3536_b0 , w_6170 );
not ( w_6170 , w_6171 );
and ( w_6171 , \3563_b1 , \3563_b0 );
or ( \3636_b1 , \2971_A[4]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6172 );
and ( \3636_b0 , \2971_A[4]_b0 , w_6173 );
and ( w_6172 , w_6173 , \2995_B[7]_b0 );
or ( \3637_b1 , \3635_b1 , \3636_b1 );
not ( \3636_b1 , w_6174 );
and ( \3637_b0 , \3635_b0 , w_6175 );
and ( w_6174 , w_6175 , \3636_b0 );
or ( \3638_b1 , \3635_b1 , \3636_b1 );
xor ( \3638_b0 , \3635_b0 , w_6176 );
not ( w_6176 , w_6177 );
and ( w_6177 , \3636_b1 , \3636_b0 );
or ( \3639_b1 , \3540_b1 , \3561_b1 );
xor ( \3639_b0 , \3540_b0 , w_6178 );
not ( w_6178 , w_6179 );
and ( w_6179 , \3561_b1 , \3561_b0 );
or ( \3640_b1 , \2975_A[3]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6180 );
and ( \3640_b0 , \2975_A[3]_b0 , w_6181 );
and ( w_6180 , w_6181 , \2995_B[7]_b0 );
or ( \3641_b1 , \3639_b1 , \3640_b1 );
not ( \3640_b1 , w_6182 );
and ( \3641_b0 , \3639_b0 , w_6183 );
and ( w_6182 , w_6183 , \3640_b0 );
or ( \3642_b1 , \3639_b1 , \3640_b1 );
xor ( \3642_b0 , \3639_b0 , w_6184 );
not ( w_6184 , w_6185 );
and ( w_6185 , \3640_b1 , \3640_b0 );
or ( \3643_b1 , \3544_b1 , \3559_b1 );
xor ( \3643_b0 , \3544_b0 , w_6186 );
not ( w_6186 , w_6187 );
and ( w_6187 , \3559_b1 , \3559_b0 );
or ( \3644_b1 , \2979_A[2]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6188 );
and ( \3644_b0 , \2979_A[2]_b0 , w_6189 );
and ( w_6188 , w_6189 , \2995_B[7]_b0 );
or ( \3645_b1 , \3643_b1 , \3644_b1 );
not ( \3644_b1 , w_6190 );
and ( \3645_b0 , \3643_b0 , w_6191 );
and ( w_6190 , w_6191 , \3644_b0 );
or ( \3646_b1 , \3643_b1 , \3644_b1 );
xor ( \3646_b0 , \3643_b0 , w_6192 );
not ( w_6192 , w_6193 );
and ( w_6193 , \3644_b1 , \3644_b0 );
or ( \3647_b1 , \3548_b1 , \3557_b1 );
xor ( \3647_b0 , \3548_b0 , w_6194 );
not ( w_6194 , w_6195 );
and ( w_6195 , \3557_b1 , \3557_b0 );
or ( \3648_b1 , \2983_A[1]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6196 );
and ( \3648_b0 , \2983_A[1]_b0 , w_6197 );
and ( w_6196 , w_6197 , \2995_B[7]_b0 );
or ( \3649_b1 , \3647_b1 , \3648_b1 );
not ( \3648_b1 , w_6198 );
and ( \3649_b0 , \3647_b0 , w_6199 );
and ( w_6198 , w_6199 , \3648_b0 );
or ( \3650_b1 , \3647_b1 , \3648_b1 );
xor ( \3650_b0 , \3647_b0 , w_6200 );
not ( w_6200 , w_6201 );
and ( w_6201 , \3648_b1 , \3648_b0 );
or ( \3651_b1 , \3552_b1 , \3555_b1 );
xor ( \3651_b0 , \3552_b0 , w_6202 );
not ( w_6202 , w_6203 );
and ( w_6203 , \3555_b1 , \3555_b0 );
or ( \3652_b1 , \2986_A[0]_b1 , \2995_B[7]_b1 );
not ( \2995_B[7]_b1 , w_6204 );
and ( \3652_b0 , \2986_A[0]_b0 , w_6205 );
and ( w_6204 , w_6205 , \2995_B[7]_b0 );
or ( \3653_b1 , \3651_b1 , \3652_b1 );
not ( \3652_b1 , w_6206 );
and ( \3653_b0 , \3651_b0 , w_6207 );
and ( w_6206 , w_6207 , \3652_b0 );
or ( \3654_b1 , \3650_b1 , \3653_b1 );
not ( \3653_b1 , w_6208 );
and ( \3654_b0 , \3650_b0 , w_6209 );
and ( w_6208 , w_6209 , \3653_b0 );
or ( \3655_b1 , \3649_b1 , w_6210 );
or ( \3655_b0 , \3649_b0 , \3654_b0 );
not ( \3654_b0 , w_6211 );
and ( w_6211 , w_6210 , \3654_b1 );
or ( \3656_b1 , \3646_b1 , \3655_b1 );
not ( \3655_b1 , w_6212 );
and ( \3656_b0 , \3646_b0 , w_6213 );
and ( w_6212 , w_6213 , \3655_b0 );
or ( \3657_b1 , \3645_b1 , w_6214 );
or ( \3657_b0 , \3645_b0 , \3656_b0 );
not ( \3656_b0 , w_6215 );
and ( w_6215 , w_6214 , \3656_b1 );
or ( \3658_b1 , \3642_b1 , \3657_b1 );
not ( \3657_b1 , w_6216 );
and ( \3658_b0 , \3642_b0 , w_6217 );
and ( w_6216 , w_6217 , \3657_b0 );
or ( \3659_b1 , \3641_b1 , w_6218 );
or ( \3659_b0 , \3641_b0 , \3658_b0 );
not ( \3658_b0 , w_6219 );
and ( w_6219 , w_6218 , \3658_b1 );
or ( \3660_b1 , \3638_b1 , \3659_b1 );
not ( \3659_b1 , w_6220 );
and ( \3660_b0 , \3638_b0 , w_6221 );
and ( w_6220 , w_6221 , \3659_b0 );
or ( \3661_b1 , \3637_b1 , w_6222 );
or ( \3661_b0 , \3637_b0 , \3660_b0 );
not ( \3660_b0 , w_6223 );
and ( w_6223 , w_6222 , \3660_b1 );
or ( \3662_b1 , \3634_b1 , \3661_b1 );
not ( \3661_b1 , w_6224 );
and ( \3662_b0 , \3634_b0 , w_6225 );
and ( w_6224 , w_6225 , \3661_b0 );
or ( \3663_b1 , \3633_b1 , w_6226 );
or ( \3663_b0 , \3633_b0 , \3662_b0 );
not ( \3662_b0 , w_6227 );
and ( w_6227 , w_6226 , \3662_b1 );
or ( \3664_b1 , \3630_b1 , \3663_b1 );
not ( \3663_b1 , w_6228 );
and ( \3664_b0 , \3630_b0 , w_6229 );
and ( w_6228 , w_6229 , \3663_b0 );
or ( \3665_b1 , \3629_b1 , w_6230 );
or ( \3665_b0 , \3629_b0 , \3664_b0 );
not ( \3664_b0 , w_6231 );
and ( w_6231 , w_6230 , \3664_b1 );
or ( \3666_b1 , \3626_b1 , \3665_b1 );
not ( \3665_b1 , w_6232 );
and ( \3666_b0 , \3626_b0 , w_6233 );
and ( w_6232 , w_6233 , \3665_b0 );
or ( \3667_b1 , \3625_b1 , w_6234 );
or ( \3667_b0 , \3625_b0 , \3666_b0 );
not ( \3666_b0 , w_6235 );
and ( w_6235 , w_6234 , \3666_b1 );
or ( \3668_b1 , \3622_b1 , \3667_b1 );
not ( \3667_b1 , w_6236 );
and ( \3668_b0 , \3622_b0 , w_6237 );
and ( w_6236 , w_6237 , \3667_b0 );
or ( \3669_b1 , \3621_b1 , w_6238 );
or ( \3669_b0 , \3621_b0 , \3668_b0 );
not ( \3668_b0 , w_6239 );
and ( w_6239 , w_6238 , \3668_b1 );
or ( \3670_b1 , \3618_b1 , \3669_b1 );
not ( \3669_b1 , w_6240 );
and ( \3670_b0 , \3618_b0 , w_6241 );
and ( w_6240 , w_6241 , \3669_b0 );
or ( \3671_b1 , \3617_b1 , w_6242 );
or ( \3671_b0 , \3617_b0 , \3670_b0 );
not ( \3670_b0 , w_6243 );
and ( w_6243 , w_6242 , \3670_b1 );
or ( \3672_b1 , \3614_b1 , \3671_b1 );
not ( \3671_b1 , w_6244 );
and ( \3672_b0 , \3614_b0 , w_6245 );
and ( w_6244 , w_6245 , \3671_b0 );
or ( \3673_b1 , \3613_b1 , w_6246 );
or ( \3673_b0 , \3613_b0 , \3672_b0 );
not ( \3672_b0 , w_6247 );
and ( w_6247 , w_6246 , \3672_b1 );
or ( \3674_b1 , \3610_b1 , \3673_b1 );
not ( \3673_b1 , w_6248 );
and ( \3674_b0 , \3610_b0 , w_6249 );
and ( w_6248 , w_6249 , \3673_b0 );
or ( \3675_b1 , \3609_b1 , w_6250 );
or ( \3675_b0 , \3609_b0 , \3674_b0 );
not ( \3674_b0 , w_6251 );
and ( w_6251 , w_6250 , \3674_b1 );
or ( \3676_b1 , \3606_b1 , \3675_b1 );
not ( \3675_b1 , w_6252 );
and ( \3676_b0 , \3606_b0 , w_6253 );
and ( w_6252 , w_6253 , \3675_b0 );
or ( \3677_b1 , \3605_b1 , w_6254 );
or ( \3677_b0 , \3605_b0 , \3676_b0 );
not ( \3676_b0 , w_6255 );
and ( w_6255 , w_6254 , \3676_b1 );
or ( \3678_b1 , \3602_b1 , \3677_b1 );
not ( \3677_b1 , w_6256 );
and ( \3678_b0 , \3602_b0 , w_6257 );
and ( w_6256 , w_6257 , \3677_b0 );
or ( \3679_b1 , \3601_b1 , w_6258 );
or ( \3679_b0 , \3601_b0 , \3678_b0 );
not ( \3678_b0 , w_6259 );
and ( w_6259 , w_6258 , \3678_b1 );
or ( \3680_b1 , \3598_b1 , \3679_b1 );
not ( \3679_b1 , w_6260 );
and ( \3680_b0 , \3598_b0 , w_6261 );
and ( w_6260 , w_6261 , \3679_b0 );
or ( \3681_b1 , \3597_b1 , w_6262 );
or ( \3681_b0 , \3597_b0 , \3680_b0 );
not ( \3680_b0 , w_6263 );
and ( w_6263 , w_6262 , \3680_b1 );
or ( \3682_b1 , \3594_b1 , \3681_b1 );
not ( \3681_b1 , w_6264 );
and ( \3682_b0 , \3594_b0 , w_6265 );
and ( w_6264 , w_6265 , \3681_b0 );
or ( \3683_b1 , \3593_b1 , w_6266 );
or ( \3683_b0 , \3593_b0 , \3682_b0 );
not ( \3682_b0 , w_6267 );
and ( w_6267 , w_6266 , \3682_b1 );
or ( \3684_b1 , \3590_b1 , \3683_b1 );
not ( \3683_b1 , w_6268 );
and ( \3684_b0 , \3590_b0 , w_6269 );
and ( w_6268 , w_6269 , \3683_b0 );
or ( \3685_b1 , \3589_b1 , w_6270 );
or ( \3685_b0 , \3589_b0 , \3684_b0 );
not ( \3684_b0 , w_6271 );
and ( w_6271 , w_6270 , \3684_b1 );
or ( \3686_b1 , \2923_A[16]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6272 );
and ( \3686_b0 , \2923_A[16]_b0 , w_6273 );
and ( w_6272 , w_6273 , \2994_B[8]_b0 );
or ( \3687_b1 , \3685_b1 , \3686_b1 );
not ( \3686_b1 , w_6274 );
and ( \3687_b0 , \3685_b0 , w_6275 );
and ( w_6274 , w_6275 , \3686_b0 );
or ( \3688_b1 , \3685_b1 , \3686_b1 );
xor ( \3688_b0 , \3685_b0 , w_6276 );
not ( w_6276 , w_6277 );
and ( w_6277 , \3686_b1 , \3686_b0 );
or ( \3689_b1 , \3590_b1 , \3683_b1 );
xor ( \3689_b0 , \3590_b0 , w_6278 );
not ( w_6278 , w_6279 );
and ( w_6279 , \3683_b1 , \3683_b0 );
or ( \3690_b1 , \2927_A[15]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6280 );
and ( \3690_b0 , \2927_A[15]_b0 , w_6281 );
and ( w_6280 , w_6281 , \2994_B[8]_b0 );
or ( \3691_b1 , \3689_b1 , \3690_b1 );
not ( \3690_b1 , w_6282 );
and ( \3691_b0 , \3689_b0 , w_6283 );
and ( w_6282 , w_6283 , \3690_b0 );
or ( \3692_b1 , \3689_b1 , \3690_b1 );
xor ( \3692_b0 , \3689_b0 , w_6284 );
not ( w_6284 , w_6285 );
and ( w_6285 , \3690_b1 , \3690_b0 );
or ( \3693_b1 , \3594_b1 , \3681_b1 );
xor ( \3693_b0 , \3594_b0 , w_6286 );
not ( w_6286 , w_6287 );
and ( w_6287 , \3681_b1 , \3681_b0 );
or ( \3694_b1 , \2931_A[14]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6288 );
and ( \3694_b0 , \2931_A[14]_b0 , w_6289 );
and ( w_6288 , w_6289 , \2994_B[8]_b0 );
or ( \3695_b1 , \3693_b1 , \3694_b1 );
not ( \3694_b1 , w_6290 );
and ( \3695_b0 , \3693_b0 , w_6291 );
and ( w_6290 , w_6291 , \3694_b0 );
or ( \3696_b1 , \3693_b1 , \3694_b1 );
xor ( \3696_b0 , \3693_b0 , w_6292 );
not ( w_6292 , w_6293 );
and ( w_6293 , \3694_b1 , \3694_b0 );
or ( \3697_b1 , \3598_b1 , \3679_b1 );
xor ( \3697_b0 , \3598_b0 , w_6294 );
not ( w_6294 , w_6295 );
and ( w_6295 , \3679_b1 , \3679_b0 );
or ( \3698_b1 , \2935_A[13]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6296 );
and ( \3698_b0 , \2935_A[13]_b0 , w_6297 );
and ( w_6296 , w_6297 , \2994_B[8]_b0 );
or ( \3699_b1 , \3697_b1 , \3698_b1 );
not ( \3698_b1 , w_6298 );
and ( \3699_b0 , \3697_b0 , w_6299 );
and ( w_6298 , w_6299 , \3698_b0 );
or ( \3700_b1 , \3697_b1 , \3698_b1 );
xor ( \3700_b0 , \3697_b0 , w_6300 );
not ( w_6300 , w_6301 );
and ( w_6301 , \3698_b1 , \3698_b0 );
or ( \3701_b1 , \3602_b1 , \3677_b1 );
xor ( \3701_b0 , \3602_b0 , w_6302 );
not ( w_6302 , w_6303 );
and ( w_6303 , \3677_b1 , \3677_b0 );
or ( \3702_b1 , \2939_A[12]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6304 );
and ( \3702_b0 , \2939_A[12]_b0 , w_6305 );
and ( w_6304 , w_6305 , \2994_B[8]_b0 );
or ( \3703_b1 , \3701_b1 , \3702_b1 );
not ( \3702_b1 , w_6306 );
and ( \3703_b0 , \3701_b0 , w_6307 );
and ( w_6306 , w_6307 , \3702_b0 );
or ( \3704_b1 , \3701_b1 , \3702_b1 );
xor ( \3704_b0 , \3701_b0 , w_6308 );
not ( w_6308 , w_6309 );
and ( w_6309 , \3702_b1 , \3702_b0 );
or ( \3705_b1 , \3606_b1 , \3675_b1 );
xor ( \3705_b0 , \3606_b0 , w_6310 );
not ( w_6310 , w_6311 );
and ( w_6311 , \3675_b1 , \3675_b0 );
or ( \3706_b1 , \2943_A[11]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6312 );
and ( \3706_b0 , \2943_A[11]_b0 , w_6313 );
and ( w_6312 , w_6313 , \2994_B[8]_b0 );
or ( \3707_b1 , \3705_b1 , \3706_b1 );
not ( \3706_b1 , w_6314 );
and ( \3707_b0 , \3705_b0 , w_6315 );
and ( w_6314 , w_6315 , \3706_b0 );
or ( \3708_b1 , \3705_b1 , \3706_b1 );
xor ( \3708_b0 , \3705_b0 , w_6316 );
not ( w_6316 , w_6317 );
and ( w_6317 , \3706_b1 , \3706_b0 );
or ( \3709_b1 , \3610_b1 , \3673_b1 );
xor ( \3709_b0 , \3610_b0 , w_6318 );
not ( w_6318 , w_6319 );
and ( w_6319 , \3673_b1 , \3673_b0 );
or ( \3710_b1 , \2947_A[10]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6320 );
and ( \3710_b0 , \2947_A[10]_b0 , w_6321 );
and ( w_6320 , w_6321 , \2994_B[8]_b0 );
or ( \3711_b1 , \3709_b1 , \3710_b1 );
not ( \3710_b1 , w_6322 );
and ( \3711_b0 , \3709_b0 , w_6323 );
and ( w_6322 , w_6323 , \3710_b0 );
or ( \3712_b1 , \3709_b1 , \3710_b1 );
xor ( \3712_b0 , \3709_b0 , w_6324 );
not ( w_6324 , w_6325 );
and ( w_6325 , \3710_b1 , \3710_b0 );
or ( \3713_b1 , \3614_b1 , \3671_b1 );
xor ( \3713_b0 , \3614_b0 , w_6326 );
not ( w_6326 , w_6327 );
and ( w_6327 , \3671_b1 , \3671_b0 );
or ( \3714_b1 , \2951_A[9]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6328 );
and ( \3714_b0 , \2951_A[9]_b0 , w_6329 );
and ( w_6328 , w_6329 , \2994_B[8]_b0 );
or ( \3715_b1 , \3713_b1 , \3714_b1 );
not ( \3714_b1 , w_6330 );
and ( \3715_b0 , \3713_b0 , w_6331 );
and ( w_6330 , w_6331 , \3714_b0 );
or ( \3716_b1 , \3713_b1 , \3714_b1 );
xor ( \3716_b0 , \3713_b0 , w_6332 );
not ( w_6332 , w_6333 );
and ( w_6333 , \3714_b1 , \3714_b0 );
or ( \3717_b1 , \3618_b1 , \3669_b1 );
xor ( \3717_b0 , \3618_b0 , w_6334 );
not ( w_6334 , w_6335 );
and ( w_6335 , \3669_b1 , \3669_b0 );
or ( \3718_b1 , \2955_A[8]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6336 );
and ( \3718_b0 , \2955_A[8]_b0 , w_6337 );
and ( w_6336 , w_6337 , \2994_B[8]_b0 );
or ( \3719_b1 , \3717_b1 , \3718_b1 );
not ( \3718_b1 , w_6338 );
and ( \3719_b0 , \3717_b0 , w_6339 );
and ( w_6338 , w_6339 , \3718_b0 );
or ( \3720_b1 , \3717_b1 , \3718_b1 );
xor ( \3720_b0 , \3717_b0 , w_6340 );
not ( w_6340 , w_6341 );
and ( w_6341 , \3718_b1 , \3718_b0 );
or ( \3721_b1 , \3622_b1 , \3667_b1 );
xor ( \3721_b0 , \3622_b0 , w_6342 );
not ( w_6342 , w_6343 );
and ( w_6343 , \3667_b1 , \3667_b0 );
or ( \3722_b1 , \2959_A[7]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6344 );
and ( \3722_b0 , \2959_A[7]_b0 , w_6345 );
and ( w_6344 , w_6345 , \2994_B[8]_b0 );
or ( \3723_b1 , \3721_b1 , \3722_b1 );
not ( \3722_b1 , w_6346 );
and ( \3723_b0 , \3721_b0 , w_6347 );
and ( w_6346 , w_6347 , \3722_b0 );
or ( \3724_b1 , \3721_b1 , \3722_b1 );
xor ( \3724_b0 , \3721_b0 , w_6348 );
not ( w_6348 , w_6349 );
and ( w_6349 , \3722_b1 , \3722_b0 );
or ( \3725_b1 , \3626_b1 , \3665_b1 );
xor ( \3725_b0 , \3626_b0 , w_6350 );
not ( w_6350 , w_6351 );
and ( w_6351 , \3665_b1 , \3665_b0 );
or ( \3726_b1 , \2963_A[6]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6352 );
and ( \3726_b0 , \2963_A[6]_b0 , w_6353 );
and ( w_6352 , w_6353 , \2994_B[8]_b0 );
or ( \3727_b1 , \3725_b1 , \3726_b1 );
not ( \3726_b1 , w_6354 );
and ( \3727_b0 , \3725_b0 , w_6355 );
and ( w_6354 , w_6355 , \3726_b0 );
or ( \3728_b1 , \3725_b1 , \3726_b1 );
xor ( \3728_b0 , \3725_b0 , w_6356 );
not ( w_6356 , w_6357 );
and ( w_6357 , \3726_b1 , \3726_b0 );
or ( \3729_b1 , \3630_b1 , \3663_b1 );
xor ( \3729_b0 , \3630_b0 , w_6358 );
not ( w_6358 , w_6359 );
and ( w_6359 , \3663_b1 , \3663_b0 );
or ( \3730_b1 , \2967_A[5]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6360 );
and ( \3730_b0 , \2967_A[5]_b0 , w_6361 );
and ( w_6360 , w_6361 , \2994_B[8]_b0 );
or ( \3731_b1 , \3729_b1 , \3730_b1 );
not ( \3730_b1 , w_6362 );
and ( \3731_b0 , \3729_b0 , w_6363 );
and ( w_6362 , w_6363 , \3730_b0 );
or ( \3732_b1 , \3729_b1 , \3730_b1 );
xor ( \3732_b0 , \3729_b0 , w_6364 );
not ( w_6364 , w_6365 );
and ( w_6365 , \3730_b1 , \3730_b0 );
or ( \3733_b1 , \3634_b1 , \3661_b1 );
xor ( \3733_b0 , \3634_b0 , w_6366 );
not ( w_6366 , w_6367 );
and ( w_6367 , \3661_b1 , \3661_b0 );
or ( \3734_b1 , \2971_A[4]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6368 );
and ( \3734_b0 , \2971_A[4]_b0 , w_6369 );
and ( w_6368 , w_6369 , \2994_B[8]_b0 );
or ( \3735_b1 , \3733_b1 , \3734_b1 );
not ( \3734_b1 , w_6370 );
and ( \3735_b0 , \3733_b0 , w_6371 );
and ( w_6370 , w_6371 , \3734_b0 );
or ( \3736_b1 , \3733_b1 , \3734_b1 );
xor ( \3736_b0 , \3733_b0 , w_6372 );
not ( w_6372 , w_6373 );
and ( w_6373 , \3734_b1 , \3734_b0 );
or ( \3737_b1 , \3638_b1 , \3659_b1 );
xor ( \3737_b0 , \3638_b0 , w_6374 );
not ( w_6374 , w_6375 );
and ( w_6375 , \3659_b1 , \3659_b0 );
or ( \3738_b1 , \2975_A[3]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6376 );
and ( \3738_b0 , \2975_A[3]_b0 , w_6377 );
and ( w_6376 , w_6377 , \2994_B[8]_b0 );
or ( \3739_b1 , \3737_b1 , \3738_b1 );
not ( \3738_b1 , w_6378 );
and ( \3739_b0 , \3737_b0 , w_6379 );
and ( w_6378 , w_6379 , \3738_b0 );
or ( \3740_b1 , \3737_b1 , \3738_b1 );
xor ( \3740_b0 , \3737_b0 , w_6380 );
not ( w_6380 , w_6381 );
and ( w_6381 , \3738_b1 , \3738_b0 );
or ( \3741_b1 , \3642_b1 , \3657_b1 );
xor ( \3741_b0 , \3642_b0 , w_6382 );
not ( w_6382 , w_6383 );
and ( w_6383 , \3657_b1 , \3657_b0 );
or ( \3742_b1 , \2979_A[2]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6384 );
and ( \3742_b0 , \2979_A[2]_b0 , w_6385 );
and ( w_6384 , w_6385 , \2994_B[8]_b0 );
or ( \3743_b1 , \3741_b1 , \3742_b1 );
not ( \3742_b1 , w_6386 );
and ( \3743_b0 , \3741_b0 , w_6387 );
and ( w_6386 , w_6387 , \3742_b0 );
or ( \3744_b1 , \3741_b1 , \3742_b1 );
xor ( \3744_b0 , \3741_b0 , w_6388 );
not ( w_6388 , w_6389 );
and ( w_6389 , \3742_b1 , \3742_b0 );
or ( \3745_b1 , \3646_b1 , \3655_b1 );
xor ( \3745_b0 , \3646_b0 , w_6390 );
not ( w_6390 , w_6391 );
and ( w_6391 , \3655_b1 , \3655_b0 );
or ( \3746_b1 , \2983_A[1]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6392 );
and ( \3746_b0 , \2983_A[1]_b0 , w_6393 );
and ( w_6392 , w_6393 , \2994_B[8]_b0 );
or ( \3747_b1 , \3745_b1 , \3746_b1 );
not ( \3746_b1 , w_6394 );
and ( \3747_b0 , \3745_b0 , w_6395 );
and ( w_6394 , w_6395 , \3746_b0 );
or ( \3748_b1 , \3745_b1 , \3746_b1 );
xor ( \3748_b0 , \3745_b0 , w_6396 );
not ( w_6396 , w_6397 );
and ( w_6397 , \3746_b1 , \3746_b0 );
or ( \3749_b1 , \3650_b1 , \3653_b1 );
xor ( \3749_b0 , \3650_b0 , w_6398 );
not ( w_6398 , w_6399 );
and ( w_6399 , \3653_b1 , \3653_b0 );
or ( \3750_b1 , \2986_A[0]_b1 , \2994_B[8]_b1 );
not ( \2994_B[8]_b1 , w_6400 );
and ( \3750_b0 , \2986_A[0]_b0 , w_6401 );
and ( w_6400 , w_6401 , \2994_B[8]_b0 );
or ( \3751_b1 , \3749_b1 , \3750_b1 );
not ( \3750_b1 , w_6402 );
and ( \3751_b0 , \3749_b0 , w_6403 );
and ( w_6402 , w_6403 , \3750_b0 );
or ( \3752_b1 , \3748_b1 , \3751_b1 );
not ( \3751_b1 , w_6404 );
and ( \3752_b0 , \3748_b0 , w_6405 );
and ( w_6404 , w_6405 , \3751_b0 );
or ( \3753_b1 , \3747_b1 , w_6406 );
or ( \3753_b0 , \3747_b0 , \3752_b0 );
not ( \3752_b0 , w_6407 );
and ( w_6407 , w_6406 , \3752_b1 );
or ( \3754_b1 , \3744_b1 , \3753_b1 );
not ( \3753_b1 , w_6408 );
and ( \3754_b0 , \3744_b0 , w_6409 );
and ( w_6408 , w_6409 , \3753_b0 );
or ( \3755_b1 , \3743_b1 , w_6410 );
or ( \3755_b0 , \3743_b0 , \3754_b0 );
not ( \3754_b0 , w_6411 );
and ( w_6411 , w_6410 , \3754_b1 );
or ( \3756_b1 , \3740_b1 , \3755_b1 );
not ( \3755_b1 , w_6412 );
and ( \3756_b0 , \3740_b0 , w_6413 );
and ( w_6412 , w_6413 , \3755_b0 );
or ( \3757_b1 , \3739_b1 , w_6414 );
or ( \3757_b0 , \3739_b0 , \3756_b0 );
not ( \3756_b0 , w_6415 );
and ( w_6415 , w_6414 , \3756_b1 );
or ( \3758_b1 , \3736_b1 , \3757_b1 );
not ( \3757_b1 , w_6416 );
and ( \3758_b0 , \3736_b0 , w_6417 );
and ( w_6416 , w_6417 , \3757_b0 );
or ( \3759_b1 , \3735_b1 , w_6418 );
or ( \3759_b0 , \3735_b0 , \3758_b0 );
not ( \3758_b0 , w_6419 );
and ( w_6419 , w_6418 , \3758_b1 );
or ( \3760_b1 , \3732_b1 , \3759_b1 );
not ( \3759_b1 , w_6420 );
and ( \3760_b0 , \3732_b0 , w_6421 );
and ( w_6420 , w_6421 , \3759_b0 );
or ( \3761_b1 , \3731_b1 , w_6422 );
or ( \3761_b0 , \3731_b0 , \3760_b0 );
not ( \3760_b0 , w_6423 );
and ( w_6423 , w_6422 , \3760_b1 );
or ( \3762_b1 , \3728_b1 , \3761_b1 );
not ( \3761_b1 , w_6424 );
and ( \3762_b0 , \3728_b0 , w_6425 );
and ( w_6424 , w_6425 , \3761_b0 );
or ( \3763_b1 , \3727_b1 , w_6426 );
or ( \3763_b0 , \3727_b0 , \3762_b0 );
not ( \3762_b0 , w_6427 );
and ( w_6427 , w_6426 , \3762_b1 );
or ( \3764_b1 , \3724_b1 , \3763_b1 );
not ( \3763_b1 , w_6428 );
and ( \3764_b0 , \3724_b0 , w_6429 );
and ( w_6428 , w_6429 , \3763_b0 );
or ( \3765_b1 , \3723_b1 , w_6430 );
or ( \3765_b0 , \3723_b0 , \3764_b0 );
not ( \3764_b0 , w_6431 );
and ( w_6431 , w_6430 , \3764_b1 );
or ( \3766_b1 , \3720_b1 , \3765_b1 );
not ( \3765_b1 , w_6432 );
and ( \3766_b0 , \3720_b0 , w_6433 );
and ( w_6432 , w_6433 , \3765_b0 );
or ( \3767_b1 , \3719_b1 , w_6434 );
or ( \3767_b0 , \3719_b0 , \3766_b0 );
not ( \3766_b0 , w_6435 );
and ( w_6435 , w_6434 , \3766_b1 );
or ( \3768_b1 , \3716_b1 , \3767_b1 );
not ( \3767_b1 , w_6436 );
and ( \3768_b0 , \3716_b0 , w_6437 );
and ( w_6436 , w_6437 , \3767_b0 );
or ( \3769_b1 , \3715_b1 , w_6438 );
or ( \3769_b0 , \3715_b0 , \3768_b0 );
not ( \3768_b0 , w_6439 );
and ( w_6439 , w_6438 , \3768_b1 );
or ( \3770_b1 , \3712_b1 , \3769_b1 );
not ( \3769_b1 , w_6440 );
and ( \3770_b0 , \3712_b0 , w_6441 );
and ( w_6440 , w_6441 , \3769_b0 );
or ( \3771_b1 , \3711_b1 , w_6442 );
or ( \3771_b0 , \3711_b0 , \3770_b0 );
not ( \3770_b0 , w_6443 );
and ( w_6443 , w_6442 , \3770_b1 );
or ( \3772_b1 , \3708_b1 , \3771_b1 );
not ( \3771_b1 , w_6444 );
and ( \3772_b0 , \3708_b0 , w_6445 );
and ( w_6444 , w_6445 , \3771_b0 );
or ( \3773_b1 , \3707_b1 , w_6446 );
or ( \3773_b0 , \3707_b0 , \3772_b0 );
not ( \3772_b0 , w_6447 );
and ( w_6447 , w_6446 , \3772_b1 );
or ( \3774_b1 , \3704_b1 , \3773_b1 );
not ( \3773_b1 , w_6448 );
and ( \3774_b0 , \3704_b0 , w_6449 );
and ( w_6448 , w_6449 , \3773_b0 );
or ( \3775_b1 , \3703_b1 , w_6450 );
or ( \3775_b0 , \3703_b0 , \3774_b0 );
not ( \3774_b0 , w_6451 );
and ( w_6451 , w_6450 , \3774_b1 );
or ( \3776_b1 , \3700_b1 , \3775_b1 );
not ( \3775_b1 , w_6452 );
and ( \3776_b0 , \3700_b0 , w_6453 );
and ( w_6452 , w_6453 , \3775_b0 );
or ( \3777_b1 , \3699_b1 , w_6454 );
or ( \3777_b0 , \3699_b0 , \3776_b0 );
not ( \3776_b0 , w_6455 );
and ( w_6455 , w_6454 , \3776_b1 );
or ( \3778_b1 , \3696_b1 , \3777_b1 );
not ( \3777_b1 , w_6456 );
and ( \3778_b0 , \3696_b0 , w_6457 );
and ( w_6456 , w_6457 , \3777_b0 );
or ( \3779_b1 , \3695_b1 , w_6458 );
or ( \3779_b0 , \3695_b0 , \3778_b0 );
not ( \3778_b0 , w_6459 );
and ( w_6459 , w_6458 , \3778_b1 );
or ( \3780_b1 , \3692_b1 , \3779_b1 );
not ( \3779_b1 , w_6460 );
and ( \3780_b0 , \3692_b0 , w_6461 );
and ( w_6460 , w_6461 , \3779_b0 );
or ( \3781_b1 , \3691_b1 , w_6462 );
or ( \3781_b0 , \3691_b0 , \3780_b0 );
not ( \3780_b0 , w_6463 );
and ( w_6463 , w_6462 , \3780_b1 );
or ( \3782_b1 , \3688_b1 , \3781_b1 );
not ( \3781_b1 , w_6464 );
and ( \3782_b0 , \3688_b0 , w_6465 );
and ( w_6464 , w_6465 , \3781_b0 );
or ( \3783_b1 , \3687_b1 , w_6466 );
or ( \3783_b0 , \3687_b0 , \3782_b0 );
not ( \3782_b0 , w_6467 );
and ( w_6467 , w_6466 , \3782_b1 );
or ( \3784_b1 , \2923_A[16]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6468 );
and ( \3784_b0 , \2923_A[16]_b0 , w_6469 );
and ( w_6468 , w_6469 , \2993_B[9]_b0 );
or ( \3785_b1 , \3783_b1 , \3784_b1 );
not ( \3784_b1 , w_6470 );
and ( \3785_b0 , \3783_b0 , w_6471 );
and ( w_6470 , w_6471 , \3784_b0 );
or ( \3786_b1 , \3783_b1 , \3784_b1 );
xor ( \3786_b0 , \3783_b0 , w_6472 );
not ( w_6472 , w_6473 );
and ( w_6473 , \3784_b1 , \3784_b0 );
or ( \3787_b1 , \3688_b1 , \3781_b1 );
xor ( \3787_b0 , \3688_b0 , w_6474 );
not ( w_6474 , w_6475 );
and ( w_6475 , \3781_b1 , \3781_b0 );
or ( \3788_b1 , \2927_A[15]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6476 );
and ( \3788_b0 , \2927_A[15]_b0 , w_6477 );
and ( w_6476 , w_6477 , \2993_B[9]_b0 );
or ( \3789_b1 , \3787_b1 , \3788_b1 );
not ( \3788_b1 , w_6478 );
and ( \3789_b0 , \3787_b0 , w_6479 );
and ( w_6478 , w_6479 , \3788_b0 );
or ( \3790_b1 , \3787_b1 , \3788_b1 );
xor ( \3790_b0 , \3787_b0 , w_6480 );
not ( w_6480 , w_6481 );
and ( w_6481 , \3788_b1 , \3788_b0 );
or ( \3791_b1 , \3692_b1 , \3779_b1 );
xor ( \3791_b0 , \3692_b0 , w_6482 );
not ( w_6482 , w_6483 );
and ( w_6483 , \3779_b1 , \3779_b0 );
or ( \3792_b1 , \2931_A[14]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6484 );
and ( \3792_b0 , \2931_A[14]_b0 , w_6485 );
and ( w_6484 , w_6485 , \2993_B[9]_b0 );
or ( \3793_b1 , \3791_b1 , \3792_b1 );
not ( \3792_b1 , w_6486 );
and ( \3793_b0 , \3791_b0 , w_6487 );
and ( w_6486 , w_6487 , \3792_b0 );
or ( \3794_b1 , \3791_b1 , \3792_b1 );
xor ( \3794_b0 , \3791_b0 , w_6488 );
not ( w_6488 , w_6489 );
and ( w_6489 , \3792_b1 , \3792_b0 );
or ( \3795_b1 , \3696_b1 , \3777_b1 );
xor ( \3795_b0 , \3696_b0 , w_6490 );
not ( w_6490 , w_6491 );
and ( w_6491 , \3777_b1 , \3777_b0 );
or ( \3796_b1 , \2935_A[13]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6492 );
and ( \3796_b0 , \2935_A[13]_b0 , w_6493 );
and ( w_6492 , w_6493 , \2993_B[9]_b0 );
or ( \3797_b1 , \3795_b1 , \3796_b1 );
not ( \3796_b1 , w_6494 );
and ( \3797_b0 , \3795_b0 , w_6495 );
and ( w_6494 , w_6495 , \3796_b0 );
or ( \3798_b1 , \3795_b1 , \3796_b1 );
xor ( \3798_b0 , \3795_b0 , w_6496 );
not ( w_6496 , w_6497 );
and ( w_6497 , \3796_b1 , \3796_b0 );
or ( \3799_b1 , \3700_b1 , \3775_b1 );
xor ( \3799_b0 , \3700_b0 , w_6498 );
not ( w_6498 , w_6499 );
and ( w_6499 , \3775_b1 , \3775_b0 );
or ( \3800_b1 , \2939_A[12]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6500 );
and ( \3800_b0 , \2939_A[12]_b0 , w_6501 );
and ( w_6500 , w_6501 , \2993_B[9]_b0 );
or ( \3801_b1 , \3799_b1 , \3800_b1 );
not ( \3800_b1 , w_6502 );
and ( \3801_b0 , \3799_b0 , w_6503 );
and ( w_6502 , w_6503 , \3800_b0 );
or ( \3802_b1 , \3799_b1 , \3800_b1 );
xor ( \3802_b0 , \3799_b0 , w_6504 );
not ( w_6504 , w_6505 );
and ( w_6505 , \3800_b1 , \3800_b0 );
or ( \3803_b1 , \3704_b1 , \3773_b1 );
xor ( \3803_b0 , \3704_b0 , w_6506 );
not ( w_6506 , w_6507 );
and ( w_6507 , \3773_b1 , \3773_b0 );
or ( \3804_b1 , \2943_A[11]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6508 );
and ( \3804_b0 , \2943_A[11]_b0 , w_6509 );
and ( w_6508 , w_6509 , \2993_B[9]_b0 );
or ( \3805_b1 , \3803_b1 , \3804_b1 );
not ( \3804_b1 , w_6510 );
and ( \3805_b0 , \3803_b0 , w_6511 );
and ( w_6510 , w_6511 , \3804_b0 );
or ( \3806_b1 , \3803_b1 , \3804_b1 );
xor ( \3806_b0 , \3803_b0 , w_6512 );
not ( w_6512 , w_6513 );
and ( w_6513 , \3804_b1 , \3804_b0 );
or ( \3807_b1 , \3708_b1 , \3771_b1 );
xor ( \3807_b0 , \3708_b0 , w_6514 );
not ( w_6514 , w_6515 );
and ( w_6515 , \3771_b1 , \3771_b0 );
or ( \3808_b1 , \2947_A[10]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6516 );
and ( \3808_b0 , \2947_A[10]_b0 , w_6517 );
and ( w_6516 , w_6517 , \2993_B[9]_b0 );
or ( \3809_b1 , \3807_b1 , \3808_b1 );
not ( \3808_b1 , w_6518 );
and ( \3809_b0 , \3807_b0 , w_6519 );
and ( w_6518 , w_6519 , \3808_b0 );
or ( \3810_b1 , \3807_b1 , \3808_b1 );
xor ( \3810_b0 , \3807_b0 , w_6520 );
not ( w_6520 , w_6521 );
and ( w_6521 , \3808_b1 , \3808_b0 );
or ( \3811_b1 , \3712_b1 , \3769_b1 );
xor ( \3811_b0 , \3712_b0 , w_6522 );
not ( w_6522 , w_6523 );
and ( w_6523 , \3769_b1 , \3769_b0 );
or ( \3812_b1 , \2951_A[9]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6524 );
and ( \3812_b0 , \2951_A[9]_b0 , w_6525 );
and ( w_6524 , w_6525 , \2993_B[9]_b0 );
or ( \3813_b1 , \3811_b1 , \3812_b1 );
not ( \3812_b1 , w_6526 );
and ( \3813_b0 , \3811_b0 , w_6527 );
and ( w_6526 , w_6527 , \3812_b0 );
or ( \3814_b1 , \3811_b1 , \3812_b1 );
xor ( \3814_b0 , \3811_b0 , w_6528 );
not ( w_6528 , w_6529 );
and ( w_6529 , \3812_b1 , \3812_b0 );
or ( \3815_b1 , \3716_b1 , \3767_b1 );
xor ( \3815_b0 , \3716_b0 , w_6530 );
not ( w_6530 , w_6531 );
and ( w_6531 , \3767_b1 , \3767_b0 );
or ( \3816_b1 , \2955_A[8]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6532 );
and ( \3816_b0 , \2955_A[8]_b0 , w_6533 );
and ( w_6532 , w_6533 , \2993_B[9]_b0 );
or ( \3817_b1 , \3815_b1 , \3816_b1 );
not ( \3816_b1 , w_6534 );
and ( \3817_b0 , \3815_b0 , w_6535 );
and ( w_6534 , w_6535 , \3816_b0 );
or ( \3818_b1 , \3815_b1 , \3816_b1 );
xor ( \3818_b0 , \3815_b0 , w_6536 );
not ( w_6536 , w_6537 );
and ( w_6537 , \3816_b1 , \3816_b0 );
or ( \3819_b1 , \3720_b1 , \3765_b1 );
xor ( \3819_b0 , \3720_b0 , w_6538 );
not ( w_6538 , w_6539 );
and ( w_6539 , \3765_b1 , \3765_b0 );
or ( \3820_b1 , \2959_A[7]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6540 );
and ( \3820_b0 , \2959_A[7]_b0 , w_6541 );
and ( w_6540 , w_6541 , \2993_B[9]_b0 );
or ( \3821_b1 , \3819_b1 , \3820_b1 );
not ( \3820_b1 , w_6542 );
and ( \3821_b0 , \3819_b0 , w_6543 );
and ( w_6542 , w_6543 , \3820_b0 );
or ( \3822_b1 , \3819_b1 , \3820_b1 );
xor ( \3822_b0 , \3819_b0 , w_6544 );
not ( w_6544 , w_6545 );
and ( w_6545 , \3820_b1 , \3820_b0 );
or ( \3823_b1 , \3724_b1 , \3763_b1 );
xor ( \3823_b0 , \3724_b0 , w_6546 );
not ( w_6546 , w_6547 );
and ( w_6547 , \3763_b1 , \3763_b0 );
or ( \3824_b1 , \2963_A[6]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6548 );
and ( \3824_b0 , \2963_A[6]_b0 , w_6549 );
and ( w_6548 , w_6549 , \2993_B[9]_b0 );
or ( \3825_b1 , \3823_b1 , \3824_b1 );
not ( \3824_b1 , w_6550 );
and ( \3825_b0 , \3823_b0 , w_6551 );
and ( w_6550 , w_6551 , \3824_b0 );
or ( \3826_b1 , \3823_b1 , \3824_b1 );
xor ( \3826_b0 , \3823_b0 , w_6552 );
not ( w_6552 , w_6553 );
and ( w_6553 , \3824_b1 , \3824_b0 );
or ( \3827_b1 , \3728_b1 , \3761_b1 );
xor ( \3827_b0 , \3728_b0 , w_6554 );
not ( w_6554 , w_6555 );
and ( w_6555 , \3761_b1 , \3761_b0 );
or ( \3828_b1 , \2967_A[5]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6556 );
and ( \3828_b0 , \2967_A[5]_b0 , w_6557 );
and ( w_6556 , w_6557 , \2993_B[9]_b0 );
or ( \3829_b1 , \3827_b1 , \3828_b1 );
not ( \3828_b1 , w_6558 );
and ( \3829_b0 , \3827_b0 , w_6559 );
and ( w_6558 , w_6559 , \3828_b0 );
or ( \3830_b1 , \3827_b1 , \3828_b1 );
xor ( \3830_b0 , \3827_b0 , w_6560 );
not ( w_6560 , w_6561 );
and ( w_6561 , \3828_b1 , \3828_b0 );
or ( \3831_b1 , \3732_b1 , \3759_b1 );
xor ( \3831_b0 , \3732_b0 , w_6562 );
not ( w_6562 , w_6563 );
and ( w_6563 , \3759_b1 , \3759_b0 );
or ( \3832_b1 , \2971_A[4]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6564 );
and ( \3832_b0 , \2971_A[4]_b0 , w_6565 );
and ( w_6564 , w_6565 , \2993_B[9]_b0 );
or ( \3833_b1 , \3831_b1 , \3832_b1 );
not ( \3832_b1 , w_6566 );
and ( \3833_b0 , \3831_b0 , w_6567 );
and ( w_6566 , w_6567 , \3832_b0 );
or ( \3834_b1 , \3831_b1 , \3832_b1 );
xor ( \3834_b0 , \3831_b0 , w_6568 );
not ( w_6568 , w_6569 );
and ( w_6569 , \3832_b1 , \3832_b0 );
or ( \3835_b1 , \3736_b1 , \3757_b1 );
xor ( \3835_b0 , \3736_b0 , w_6570 );
not ( w_6570 , w_6571 );
and ( w_6571 , \3757_b1 , \3757_b0 );
or ( \3836_b1 , \2975_A[3]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6572 );
and ( \3836_b0 , \2975_A[3]_b0 , w_6573 );
and ( w_6572 , w_6573 , \2993_B[9]_b0 );
or ( \3837_b1 , \3835_b1 , \3836_b1 );
not ( \3836_b1 , w_6574 );
and ( \3837_b0 , \3835_b0 , w_6575 );
and ( w_6574 , w_6575 , \3836_b0 );
or ( \3838_b1 , \3835_b1 , \3836_b1 );
xor ( \3838_b0 , \3835_b0 , w_6576 );
not ( w_6576 , w_6577 );
and ( w_6577 , \3836_b1 , \3836_b0 );
or ( \3839_b1 , \3740_b1 , \3755_b1 );
xor ( \3839_b0 , \3740_b0 , w_6578 );
not ( w_6578 , w_6579 );
and ( w_6579 , \3755_b1 , \3755_b0 );
or ( \3840_b1 , \2979_A[2]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6580 );
and ( \3840_b0 , \2979_A[2]_b0 , w_6581 );
and ( w_6580 , w_6581 , \2993_B[9]_b0 );
or ( \3841_b1 , \3839_b1 , \3840_b1 );
not ( \3840_b1 , w_6582 );
and ( \3841_b0 , \3839_b0 , w_6583 );
and ( w_6582 , w_6583 , \3840_b0 );
or ( \3842_b1 , \3839_b1 , \3840_b1 );
xor ( \3842_b0 , \3839_b0 , w_6584 );
not ( w_6584 , w_6585 );
and ( w_6585 , \3840_b1 , \3840_b0 );
or ( \3843_b1 , \3744_b1 , \3753_b1 );
xor ( \3843_b0 , \3744_b0 , w_6586 );
not ( w_6586 , w_6587 );
and ( w_6587 , \3753_b1 , \3753_b0 );
or ( \3844_b1 , \2983_A[1]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6588 );
and ( \3844_b0 , \2983_A[1]_b0 , w_6589 );
and ( w_6588 , w_6589 , \2993_B[9]_b0 );
or ( \3845_b1 , \3843_b1 , \3844_b1 );
not ( \3844_b1 , w_6590 );
and ( \3845_b0 , \3843_b0 , w_6591 );
and ( w_6590 , w_6591 , \3844_b0 );
or ( \3846_b1 , \3843_b1 , \3844_b1 );
xor ( \3846_b0 , \3843_b0 , w_6592 );
not ( w_6592 , w_6593 );
and ( w_6593 , \3844_b1 , \3844_b0 );
or ( \3847_b1 , \3748_b1 , \3751_b1 );
xor ( \3847_b0 , \3748_b0 , w_6594 );
not ( w_6594 , w_6595 );
and ( w_6595 , \3751_b1 , \3751_b0 );
or ( \3848_b1 , \2986_A[0]_b1 , \2993_B[9]_b1 );
not ( \2993_B[9]_b1 , w_6596 );
and ( \3848_b0 , \2986_A[0]_b0 , w_6597 );
and ( w_6596 , w_6597 , \2993_B[9]_b0 );
or ( \3849_b1 , \3847_b1 , \3848_b1 );
not ( \3848_b1 , w_6598 );
and ( \3849_b0 , \3847_b0 , w_6599 );
and ( w_6598 , w_6599 , \3848_b0 );
or ( \3850_b1 , \3846_b1 , \3849_b1 );
not ( \3849_b1 , w_6600 );
and ( \3850_b0 , \3846_b0 , w_6601 );
and ( w_6600 , w_6601 , \3849_b0 );
or ( \3851_b1 , \3845_b1 , w_6602 );
or ( \3851_b0 , \3845_b0 , \3850_b0 );
not ( \3850_b0 , w_6603 );
and ( w_6603 , w_6602 , \3850_b1 );
or ( \3852_b1 , \3842_b1 , \3851_b1 );
not ( \3851_b1 , w_6604 );
and ( \3852_b0 , \3842_b0 , w_6605 );
and ( w_6604 , w_6605 , \3851_b0 );
or ( \3853_b1 , \3841_b1 , w_6606 );
or ( \3853_b0 , \3841_b0 , \3852_b0 );
not ( \3852_b0 , w_6607 );
and ( w_6607 , w_6606 , \3852_b1 );
or ( \3854_b1 , \3838_b1 , \3853_b1 );
not ( \3853_b1 , w_6608 );
and ( \3854_b0 , \3838_b0 , w_6609 );
and ( w_6608 , w_6609 , \3853_b0 );
or ( \3855_b1 , \3837_b1 , w_6610 );
or ( \3855_b0 , \3837_b0 , \3854_b0 );
not ( \3854_b0 , w_6611 );
and ( w_6611 , w_6610 , \3854_b1 );
or ( \3856_b1 , \3834_b1 , \3855_b1 );
not ( \3855_b1 , w_6612 );
and ( \3856_b0 , \3834_b0 , w_6613 );
and ( w_6612 , w_6613 , \3855_b0 );
or ( \3857_b1 , \3833_b1 , w_6614 );
or ( \3857_b0 , \3833_b0 , \3856_b0 );
not ( \3856_b0 , w_6615 );
and ( w_6615 , w_6614 , \3856_b1 );
or ( \3858_b1 , \3830_b1 , \3857_b1 );
not ( \3857_b1 , w_6616 );
and ( \3858_b0 , \3830_b0 , w_6617 );
and ( w_6616 , w_6617 , \3857_b0 );
or ( \3859_b1 , \3829_b1 , w_6618 );
or ( \3859_b0 , \3829_b0 , \3858_b0 );
not ( \3858_b0 , w_6619 );
and ( w_6619 , w_6618 , \3858_b1 );
or ( \3860_b1 , \3826_b1 , \3859_b1 );
not ( \3859_b1 , w_6620 );
and ( \3860_b0 , \3826_b0 , w_6621 );
and ( w_6620 , w_6621 , \3859_b0 );
or ( \3861_b1 , \3825_b1 , w_6622 );
or ( \3861_b0 , \3825_b0 , \3860_b0 );
not ( \3860_b0 , w_6623 );
and ( w_6623 , w_6622 , \3860_b1 );
or ( \3862_b1 , \3822_b1 , \3861_b1 );
not ( \3861_b1 , w_6624 );
and ( \3862_b0 , \3822_b0 , w_6625 );
and ( w_6624 , w_6625 , \3861_b0 );
or ( \3863_b1 , \3821_b1 , w_6626 );
or ( \3863_b0 , \3821_b0 , \3862_b0 );
not ( \3862_b0 , w_6627 );
and ( w_6627 , w_6626 , \3862_b1 );
or ( \3864_b1 , \3818_b1 , \3863_b1 );
not ( \3863_b1 , w_6628 );
and ( \3864_b0 , \3818_b0 , w_6629 );
and ( w_6628 , w_6629 , \3863_b0 );
or ( \3865_b1 , \3817_b1 , w_6630 );
or ( \3865_b0 , \3817_b0 , \3864_b0 );
not ( \3864_b0 , w_6631 );
and ( w_6631 , w_6630 , \3864_b1 );
or ( \3866_b1 , \3814_b1 , \3865_b1 );
not ( \3865_b1 , w_6632 );
and ( \3866_b0 , \3814_b0 , w_6633 );
and ( w_6632 , w_6633 , \3865_b0 );
or ( \3867_b1 , \3813_b1 , w_6634 );
or ( \3867_b0 , \3813_b0 , \3866_b0 );
not ( \3866_b0 , w_6635 );
and ( w_6635 , w_6634 , \3866_b1 );
or ( \3868_b1 , \3810_b1 , \3867_b1 );
not ( \3867_b1 , w_6636 );
and ( \3868_b0 , \3810_b0 , w_6637 );
and ( w_6636 , w_6637 , \3867_b0 );
or ( \3869_b1 , \3809_b1 , w_6638 );
or ( \3869_b0 , \3809_b0 , \3868_b0 );
not ( \3868_b0 , w_6639 );
and ( w_6639 , w_6638 , \3868_b1 );
or ( \3870_b1 , \3806_b1 , \3869_b1 );
not ( \3869_b1 , w_6640 );
and ( \3870_b0 , \3806_b0 , w_6641 );
and ( w_6640 , w_6641 , \3869_b0 );
or ( \3871_b1 , \3805_b1 , w_6642 );
or ( \3871_b0 , \3805_b0 , \3870_b0 );
not ( \3870_b0 , w_6643 );
and ( w_6643 , w_6642 , \3870_b1 );
or ( \3872_b1 , \3802_b1 , \3871_b1 );
not ( \3871_b1 , w_6644 );
and ( \3872_b0 , \3802_b0 , w_6645 );
and ( w_6644 , w_6645 , \3871_b0 );
or ( \3873_b1 , \3801_b1 , w_6646 );
or ( \3873_b0 , \3801_b0 , \3872_b0 );
not ( \3872_b0 , w_6647 );
and ( w_6647 , w_6646 , \3872_b1 );
or ( \3874_b1 , \3798_b1 , \3873_b1 );
not ( \3873_b1 , w_6648 );
and ( \3874_b0 , \3798_b0 , w_6649 );
and ( w_6648 , w_6649 , \3873_b0 );
or ( \3875_b1 , \3797_b1 , w_6650 );
or ( \3875_b0 , \3797_b0 , \3874_b0 );
not ( \3874_b0 , w_6651 );
and ( w_6651 , w_6650 , \3874_b1 );
or ( \3876_b1 , \3794_b1 , \3875_b1 );
not ( \3875_b1 , w_6652 );
and ( \3876_b0 , \3794_b0 , w_6653 );
and ( w_6652 , w_6653 , \3875_b0 );
or ( \3877_b1 , \3793_b1 , w_6654 );
or ( \3877_b0 , \3793_b0 , \3876_b0 );
not ( \3876_b0 , w_6655 );
and ( w_6655 , w_6654 , \3876_b1 );
or ( \3878_b1 , \3790_b1 , \3877_b1 );
not ( \3877_b1 , w_6656 );
and ( \3878_b0 , \3790_b0 , w_6657 );
and ( w_6656 , w_6657 , \3877_b0 );
or ( \3879_b1 , \3789_b1 , w_6658 );
or ( \3879_b0 , \3789_b0 , \3878_b0 );
not ( \3878_b0 , w_6659 );
and ( w_6659 , w_6658 , \3878_b1 );
or ( \3880_b1 , \3786_b1 , \3879_b1 );
not ( \3879_b1 , w_6660 );
and ( \3880_b0 , \3786_b0 , w_6661 );
and ( w_6660 , w_6661 , \3879_b0 );
or ( \3881_b1 , \3785_b1 , w_6662 );
or ( \3881_b0 , \3785_b0 , \3880_b0 );
not ( \3880_b0 , w_6663 );
and ( w_6663 , w_6662 , \3880_b1 );
or ( \3882_b1 , \2923_A[16]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6664 );
and ( \3882_b0 , \2923_A[16]_b0 , w_6665 );
and ( w_6664 , w_6665 , \2992_B[10]_b0 );
or ( \3883_b1 , \3881_b1 , \3882_b1 );
not ( \3882_b1 , w_6666 );
and ( \3883_b0 , \3881_b0 , w_6667 );
and ( w_6666 , w_6667 , \3882_b0 );
or ( \3884_b1 , \3881_b1 , \3882_b1 );
xor ( \3884_b0 , \3881_b0 , w_6668 );
not ( w_6668 , w_6669 );
and ( w_6669 , \3882_b1 , \3882_b0 );
or ( \3885_b1 , \3786_b1 , \3879_b1 );
xor ( \3885_b0 , \3786_b0 , w_6670 );
not ( w_6670 , w_6671 );
and ( w_6671 , \3879_b1 , \3879_b0 );
or ( \3886_b1 , \2927_A[15]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6672 );
and ( \3886_b0 , \2927_A[15]_b0 , w_6673 );
and ( w_6672 , w_6673 , \2992_B[10]_b0 );
or ( \3887_b1 , \3885_b1 , \3886_b1 );
not ( \3886_b1 , w_6674 );
and ( \3887_b0 , \3885_b0 , w_6675 );
and ( w_6674 , w_6675 , \3886_b0 );
or ( \3888_b1 , \3885_b1 , \3886_b1 );
xor ( \3888_b0 , \3885_b0 , w_6676 );
not ( w_6676 , w_6677 );
and ( w_6677 , \3886_b1 , \3886_b0 );
or ( \3889_b1 , \3790_b1 , \3877_b1 );
xor ( \3889_b0 , \3790_b0 , w_6678 );
not ( w_6678 , w_6679 );
and ( w_6679 , \3877_b1 , \3877_b0 );
or ( \3890_b1 , \2931_A[14]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6680 );
and ( \3890_b0 , \2931_A[14]_b0 , w_6681 );
and ( w_6680 , w_6681 , \2992_B[10]_b0 );
or ( \3891_b1 , \3889_b1 , \3890_b1 );
not ( \3890_b1 , w_6682 );
and ( \3891_b0 , \3889_b0 , w_6683 );
and ( w_6682 , w_6683 , \3890_b0 );
or ( \3892_b1 , \3889_b1 , \3890_b1 );
xor ( \3892_b0 , \3889_b0 , w_6684 );
not ( w_6684 , w_6685 );
and ( w_6685 , \3890_b1 , \3890_b0 );
or ( \3893_b1 , \3794_b1 , \3875_b1 );
xor ( \3893_b0 , \3794_b0 , w_6686 );
not ( w_6686 , w_6687 );
and ( w_6687 , \3875_b1 , \3875_b0 );
or ( \3894_b1 , \2935_A[13]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6688 );
and ( \3894_b0 , \2935_A[13]_b0 , w_6689 );
and ( w_6688 , w_6689 , \2992_B[10]_b0 );
or ( \3895_b1 , \3893_b1 , \3894_b1 );
not ( \3894_b1 , w_6690 );
and ( \3895_b0 , \3893_b0 , w_6691 );
and ( w_6690 , w_6691 , \3894_b0 );
or ( \3896_b1 , \3893_b1 , \3894_b1 );
xor ( \3896_b0 , \3893_b0 , w_6692 );
not ( w_6692 , w_6693 );
and ( w_6693 , \3894_b1 , \3894_b0 );
or ( \3897_b1 , \3798_b1 , \3873_b1 );
xor ( \3897_b0 , \3798_b0 , w_6694 );
not ( w_6694 , w_6695 );
and ( w_6695 , \3873_b1 , \3873_b0 );
or ( \3898_b1 , \2939_A[12]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6696 );
and ( \3898_b0 , \2939_A[12]_b0 , w_6697 );
and ( w_6696 , w_6697 , \2992_B[10]_b0 );
or ( \3899_b1 , \3897_b1 , \3898_b1 );
not ( \3898_b1 , w_6698 );
and ( \3899_b0 , \3897_b0 , w_6699 );
and ( w_6698 , w_6699 , \3898_b0 );
or ( \3900_b1 , \3897_b1 , \3898_b1 );
xor ( \3900_b0 , \3897_b0 , w_6700 );
not ( w_6700 , w_6701 );
and ( w_6701 , \3898_b1 , \3898_b0 );
or ( \3901_b1 , \3802_b1 , \3871_b1 );
xor ( \3901_b0 , \3802_b0 , w_6702 );
not ( w_6702 , w_6703 );
and ( w_6703 , \3871_b1 , \3871_b0 );
or ( \3902_b1 , \2943_A[11]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6704 );
and ( \3902_b0 , \2943_A[11]_b0 , w_6705 );
and ( w_6704 , w_6705 , \2992_B[10]_b0 );
or ( \3903_b1 , \3901_b1 , \3902_b1 );
not ( \3902_b1 , w_6706 );
and ( \3903_b0 , \3901_b0 , w_6707 );
and ( w_6706 , w_6707 , \3902_b0 );
or ( \3904_b1 , \3901_b1 , \3902_b1 );
xor ( \3904_b0 , \3901_b0 , w_6708 );
not ( w_6708 , w_6709 );
and ( w_6709 , \3902_b1 , \3902_b0 );
or ( \3905_b1 , \3806_b1 , \3869_b1 );
xor ( \3905_b0 , \3806_b0 , w_6710 );
not ( w_6710 , w_6711 );
and ( w_6711 , \3869_b1 , \3869_b0 );
or ( \3906_b1 , \2947_A[10]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6712 );
and ( \3906_b0 , \2947_A[10]_b0 , w_6713 );
and ( w_6712 , w_6713 , \2992_B[10]_b0 );
or ( \3907_b1 , \3905_b1 , \3906_b1 );
not ( \3906_b1 , w_6714 );
and ( \3907_b0 , \3905_b0 , w_6715 );
and ( w_6714 , w_6715 , \3906_b0 );
or ( \3908_b1 , \3905_b1 , \3906_b1 );
xor ( \3908_b0 , \3905_b0 , w_6716 );
not ( w_6716 , w_6717 );
and ( w_6717 , \3906_b1 , \3906_b0 );
or ( \3909_b1 , \3810_b1 , \3867_b1 );
xor ( \3909_b0 , \3810_b0 , w_6718 );
not ( w_6718 , w_6719 );
and ( w_6719 , \3867_b1 , \3867_b0 );
or ( \3910_b1 , \2951_A[9]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6720 );
and ( \3910_b0 , \2951_A[9]_b0 , w_6721 );
and ( w_6720 , w_6721 , \2992_B[10]_b0 );
or ( \3911_b1 , \3909_b1 , \3910_b1 );
not ( \3910_b1 , w_6722 );
and ( \3911_b0 , \3909_b0 , w_6723 );
and ( w_6722 , w_6723 , \3910_b0 );
or ( \3912_b1 , \3909_b1 , \3910_b1 );
xor ( \3912_b0 , \3909_b0 , w_6724 );
not ( w_6724 , w_6725 );
and ( w_6725 , \3910_b1 , \3910_b0 );
or ( \3913_b1 , \3814_b1 , \3865_b1 );
xor ( \3913_b0 , \3814_b0 , w_6726 );
not ( w_6726 , w_6727 );
and ( w_6727 , \3865_b1 , \3865_b0 );
or ( \3914_b1 , \2955_A[8]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6728 );
and ( \3914_b0 , \2955_A[8]_b0 , w_6729 );
and ( w_6728 , w_6729 , \2992_B[10]_b0 );
or ( \3915_b1 , \3913_b1 , \3914_b1 );
not ( \3914_b1 , w_6730 );
and ( \3915_b0 , \3913_b0 , w_6731 );
and ( w_6730 , w_6731 , \3914_b0 );
or ( \3916_b1 , \3913_b1 , \3914_b1 );
xor ( \3916_b0 , \3913_b0 , w_6732 );
not ( w_6732 , w_6733 );
and ( w_6733 , \3914_b1 , \3914_b0 );
or ( \3917_b1 , \3818_b1 , \3863_b1 );
xor ( \3917_b0 , \3818_b0 , w_6734 );
not ( w_6734 , w_6735 );
and ( w_6735 , \3863_b1 , \3863_b0 );
or ( \3918_b1 , \2959_A[7]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6736 );
and ( \3918_b0 , \2959_A[7]_b0 , w_6737 );
and ( w_6736 , w_6737 , \2992_B[10]_b0 );
or ( \3919_b1 , \3917_b1 , \3918_b1 );
not ( \3918_b1 , w_6738 );
and ( \3919_b0 , \3917_b0 , w_6739 );
and ( w_6738 , w_6739 , \3918_b0 );
or ( \3920_b1 , \3917_b1 , \3918_b1 );
xor ( \3920_b0 , \3917_b0 , w_6740 );
not ( w_6740 , w_6741 );
and ( w_6741 , \3918_b1 , \3918_b0 );
or ( \3921_b1 , \3822_b1 , \3861_b1 );
xor ( \3921_b0 , \3822_b0 , w_6742 );
not ( w_6742 , w_6743 );
and ( w_6743 , \3861_b1 , \3861_b0 );
or ( \3922_b1 , \2963_A[6]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6744 );
and ( \3922_b0 , \2963_A[6]_b0 , w_6745 );
and ( w_6744 , w_6745 , \2992_B[10]_b0 );
or ( \3923_b1 , \3921_b1 , \3922_b1 );
not ( \3922_b1 , w_6746 );
and ( \3923_b0 , \3921_b0 , w_6747 );
and ( w_6746 , w_6747 , \3922_b0 );
or ( \3924_b1 , \3921_b1 , \3922_b1 );
xor ( \3924_b0 , \3921_b0 , w_6748 );
not ( w_6748 , w_6749 );
and ( w_6749 , \3922_b1 , \3922_b0 );
or ( \3925_b1 , \3826_b1 , \3859_b1 );
xor ( \3925_b0 , \3826_b0 , w_6750 );
not ( w_6750 , w_6751 );
and ( w_6751 , \3859_b1 , \3859_b0 );
or ( \3926_b1 , \2967_A[5]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6752 );
and ( \3926_b0 , \2967_A[5]_b0 , w_6753 );
and ( w_6752 , w_6753 , \2992_B[10]_b0 );
or ( \3927_b1 , \3925_b1 , \3926_b1 );
not ( \3926_b1 , w_6754 );
and ( \3927_b0 , \3925_b0 , w_6755 );
and ( w_6754 , w_6755 , \3926_b0 );
or ( \3928_b1 , \3925_b1 , \3926_b1 );
xor ( \3928_b0 , \3925_b0 , w_6756 );
not ( w_6756 , w_6757 );
and ( w_6757 , \3926_b1 , \3926_b0 );
or ( \3929_b1 , \3830_b1 , \3857_b1 );
xor ( \3929_b0 , \3830_b0 , w_6758 );
not ( w_6758 , w_6759 );
and ( w_6759 , \3857_b1 , \3857_b0 );
or ( \3930_b1 , \2971_A[4]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6760 );
and ( \3930_b0 , \2971_A[4]_b0 , w_6761 );
and ( w_6760 , w_6761 , \2992_B[10]_b0 );
or ( \3931_b1 , \3929_b1 , \3930_b1 );
not ( \3930_b1 , w_6762 );
and ( \3931_b0 , \3929_b0 , w_6763 );
and ( w_6762 , w_6763 , \3930_b0 );
or ( \3932_b1 , \3929_b1 , \3930_b1 );
xor ( \3932_b0 , \3929_b0 , w_6764 );
not ( w_6764 , w_6765 );
and ( w_6765 , \3930_b1 , \3930_b0 );
or ( \3933_b1 , \3834_b1 , \3855_b1 );
xor ( \3933_b0 , \3834_b0 , w_6766 );
not ( w_6766 , w_6767 );
and ( w_6767 , \3855_b1 , \3855_b0 );
or ( \3934_b1 , \2975_A[3]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6768 );
and ( \3934_b0 , \2975_A[3]_b0 , w_6769 );
and ( w_6768 , w_6769 , \2992_B[10]_b0 );
or ( \3935_b1 , \3933_b1 , \3934_b1 );
not ( \3934_b1 , w_6770 );
and ( \3935_b0 , \3933_b0 , w_6771 );
and ( w_6770 , w_6771 , \3934_b0 );
or ( \3936_b1 , \3933_b1 , \3934_b1 );
xor ( \3936_b0 , \3933_b0 , w_6772 );
not ( w_6772 , w_6773 );
and ( w_6773 , \3934_b1 , \3934_b0 );
or ( \3937_b1 , \3838_b1 , \3853_b1 );
xor ( \3937_b0 , \3838_b0 , w_6774 );
not ( w_6774 , w_6775 );
and ( w_6775 , \3853_b1 , \3853_b0 );
or ( \3938_b1 , \2979_A[2]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6776 );
and ( \3938_b0 , \2979_A[2]_b0 , w_6777 );
and ( w_6776 , w_6777 , \2992_B[10]_b0 );
or ( \3939_b1 , \3937_b1 , \3938_b1 );
not ( \3938_b1 , w_6778 );
and ( \3939_b0 , \3937_b0 , w_6779 );
and ( w_6778 , w_6779 , \3938_b0 );
or ( \3940_b1 , \3937_b1 , \3938_b1 );
xor ( \3940_b0 , \3937_b0 , w_6780 );
not ( w_6780 , w_6781 );
and ( w_6781 , \3938_b1 , \3938_b0 );
or ( \3941_b1 , \3842_b1 , \3851_b1 );
xor ( \3941_b0 , \3842_b0 , w_6782 );
not ( w_6782 , w_6783 );
and ( w_6783 , \3851_b1 , \3851_b0 );
or ( \3942_b1 , \2983_A[1]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6784 );
and ( \3942_b0 , \2983_A[1]_b0 , w_6785 );
and ( w_6784 , w_6785 , \2992_B[10]_b0 );
or ( \3943_b1 , \3941_b1 , \3942_b1 );
not ( \3942_b1 , w_6786 );
and ( \3943_b0 , \3941_b0 , w_6787 );
and ( w_6786 , w_6787 , \3942_b0 );
or ( \3944_b1 , \3941_b1 , \3942_b1 );
xor ( \3944_b0 , \3941_b0 , w_6788 );
not ( w_6788 , w_6789 );
and ( w_6789 , \3942_b1 , \3942_b0 );
or ( \3945_b1 , \3846_b1 , \3849_b1 );
xor ( \3945_b0 , \3846_b0 , w_6790 );
not ( w_6790 , w_6791 );
and ( w_6791 , \3849_b1 , \3849_b0 );
or ( \3946_b1 , \2986_A[0]_b1 , \2992_B[10]_b1 );
not ( \2992_B[10]_b1 , w_6792 );
and ( \3946_b0 , \2986_A[0]_b0 , w_6793 );
and ( w_6792 , w_6793 , \2992_B[10]_b0 );
or ( \3947_b1 , \3945_b1 , \3946_b1 );
not ( \3946_b1 , w_6794 );
and ( \3947_b0 , \3945_b0 , w_6795 );
and ( w_6794 , w_6795 , \3946_b0 );
or ( \3948_b1 , \3944_b1 , \3947_b1 );
not ( \3947_b1 , w_6796 );
and ( \3948_b0 , \3944_b0 , w_6797 );
and ( w_6796 , w_6797 , \3947_b0 );
or ( \3949_b1 , \3943_b1 , w_6798 );
or ( \3949_b0 , \3943_b0 , \3948_b0 );
not ( \3948_b0 , w_6799 );
and ( w_6799 , w_6798 , \3948_b1 );
or ( \3950_b1 , \3940_b1 , \3949_b1 );
not ( \3949_b1 , w_6800 );
and ( \3950_b0 , \3940_b0 , w_6801 );
and ( w_6800 , w_6801 , \3949_b0 );
or ( \3951_b1 , \3939_b1 , w_6802 );
or ( \3951_b0 , \3939_b0 , \3950_b0 );
not ( \3950_b0 , w_6803 );
and ( w_6803 , w_6802 , \3950_b1 );
or ( \3952_b1 , \3936_b1 , \3951_b1 );
not ( \3951_b1 , w_6804 );
and ( \3952_b0 , \3936_b0 , w_6805 );
and ( w_6804 , w_6805 , \3951_b0 );
or ( \3953_b1 , \3935_b1 , w_6806 );
or ( \3953_b0 , \3935_b0 , \3952_b0 );
not ( \3952_b0 , w_6807 );
and ( w_6807 , w_6806 , \3952_b1 );
or ( \3954_b1 , \3932_b1 , \3953_b1 );
not ( \3953_b1 , w_6808 );
and ( \3954_b0 , \3932_b0 , w_6809 );
and ( w_6808 , w_6809 , \3953_b0 );
or ( \3955_b1 , \3931_b1 , w_6810 );
or ( \3955_b0 , \3931_b0 , \3954_b0 );
not ( \3954_b0 , w_6811 );
and ( w_6811 , w_6810 , \3954_b1 );
or ( \3956_b1 , \3928_b1 , \3955_b1 );
not ( \3955_b1 , w_6812 );
and ( \3956_b0 , \3928_b0 , w_6813 );
and ( w_6812 , w_6813 , \3955_b0 );
or ( \3957_b1 , \3927_b1 , w_6814 );
or ( \3957_b0 , \3927_b0 , \3956_b0 );
not ( \3956_b0 , w_6815 );
and ( w_6815 , w_6814 , \3956_b1 );
or ( \3958_b1 , \3924_b1 , \3957_b1 );
not ( \3957_b1 , w_6816 );
and ( \3958_b0 , \3924_b0 , w_6817 );
and ( w_6816 , w_6817 , \3957_b0 );
or ( \3959_b1 , \3923_b1 , w_6818 );
or ( \3959_b0 , \3923_b0 , \3958_b0 );
not ( \3958_b0 , w_6819 );
and ( w_6819 , w_6818 , \3958_b1 );
or ( \3960_b1 , \3920_b1 , \3959_b1 );
not ( \3959_b1 , w_6820 );
and ( \3960_b0 , \3920_b0 , w_6821 );
and ( w_6820 , w_6821 , \3959_b0 );
or ( \3961_b1 , \3919_b1 , w_6822 );
or ( \3961_b0 , \3919_b0 , \3960_b0 );
not ( \3960_b0 , w_6823 );
and ( w_6823 , w_6822 , \3960_b1 );
or ( \3962_b1 , \3916_b1 , \3961_b1 );
not ( \3961_b1 , w_6824 );
and ( \3962_b0 , \3916_b0 , w_6825 );
and ( w_6824 , w_6825 , \3961_b0 );
or ( \3963_b1 , \3915_b1 , w_6826 );
or ( \3963_b0 , \3915_b0 , \3962_b0 );
not ( \3962_b0 , w_6827 );
and ( w_6827 , w_6826 , \3962_b1 );
or ( \3964_b1 , \3912_b1 , \3963_b1 );
not ( \3963_b1 , w_6828 );
and ( \3964_b0 , \3912_b0 , w_6829 );
and ( w_6828 , w_6829 , \3963_b0 );
or ( \3965_b1 , \3911_b1 , w_6830 );
or ( \3965_b0 , \3911_b0 , \3964_b0 );
not ( \3964_b0 , w_6831 );
and ( w_6831 , w_6830 , \3964_b1 );
or ( \3966_b1 , \3908_b1 , \3965_b1 );
not ( \3965_b1 , w_6832 );
and ( \3966_b0 , \3908_b0 , w_6833 );
and ( w_6832 , w_6833 , \3965_b0 );
or ( \3967_b1 , \3907_b1 , w_6834 );
or ( \3967_b0 , \3907_b0 , \3966_b0 );
not ( \3966_b0 , w_6835 );
and ( w_6835 , w_6834 , \3966_b1 );
or ( \3968_b1 , \3904_b1 , \3967_b1 );
not ( \3967_b1 , w_6836 );
and ( \3968_b0 , \3904_b0 , w_6837 );
and ( w_6836 , w_6837 , \3967_b0 );
or ( \3969_b1 , \3903_b1 , w_6838 );
or ( \3969_b0 , \3903_b0 , \3968_b0 );
not ( \3968_b0 , w_6839 );
and ( w_6839 , w_6838 , \3968_b1 );
or ( \3970_b1 , \3900_b1 , \3969_b1 );
not ( \3969_b1 , w_6840 );
and ( \3970_b0 , \3900_b0 , w_6841 );
and ( w_6840 , w_6841 , \3969_b0 );
or ( \3971_b1 , \3899_b1 , w_6842 );
or ( \3971_b0 , \3899_b0 , \3970_b0 );
not ( \3970_b0 , w_6843 );
and ( w_6843 , w_6842 , \3970_b1 );
or ( \3972_b1 , \3896_b1 , \3971_b1 );
not ( \3971_b1 , w_6844 );
and ( \3972_b0 , \3896_b0 , w_6845 );
and ( w_6844 , w_6845 , \3971_b0 );
or ( \3973_b1 , \3895_b1 , w_6846 );
or ( \3973_b0 , \3895_b0 , \3972_b0 );
not ( \3972_b0 , w_6847 );
and ( w_6847 , w_6846 , \3972_b1 );
or ( \3974_b1 , \3892_b1 , \3973_b1 );
not ( \3973_b1 , w_6848 );
and ( \3974_b0 , \3892_b0 , w_6849 );
and ( w_6848 , w_6849 , \3973_b0 );
or ( \3975_b1 , \3891_b1 , w_6850 );
or ( \3975_b0 , \3891_b0 , \3974_b0 );
not ( \3974_b0 , w_6851 );
and ( w_6851 , w_6850 , \3974_b1 );
or ( \3976_b1 , \3888_b1 , \3975_b1 );
not ( \3975_b1 , w_6852 );
and ( \3976_b0 , \3888_b0 , w_6853 );
and ( w_6852 , w_6853 , \3975_b0 );
or ( \3977_b1 , \3887_b1 , w_6854 );
or ( \3977_b0 , \3887_b0 , \3976_b0 );
not ( \3976_b0 , w_6855 );
and ( w_6855 , w_6854 , \3976_b1 );
or ( \3978_b1 , \3884_b1 , \3977_b1 );
not ( \3977_b1 , w_6856 );
and ( \3978_b0 , \3884_b0 , w_6857 );
and ( w_6856 , w_6857 , \3977_b0 );
or ( \3979_b1 , \3883_b1 , w_6858 );
or ( \3979_b0 , \3883_b0 , \3978_b0 );
not ( \3978_b0 , w_6859 );
and ( w_6859 , w_6858 , \3978_b1 );
or ( \3980_b1 , \2923_A[16]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6860 );
and ( \3980_b0 , \2923_A[16]_b0 , w_6861 );
and ( w_6860 , w_6861 , \2991_B[11]_b0 );
or ( \3981_b1 , \3979_b1 , \3980_b1 );
not ( \3980_b1 , w_6862 );
and ( \3981_b0 , \3979_b0 , w_6863 );
and ( w_6862 , w_6863 , \3980_b0 );
or ( \3982_b1 , \3979_b1 , \3980_b1 );
xor ( \3982_b0 , \3979_b0 , w_6864 );
not ( w_6864 , w_6865 );
and ( w_6865 , \3980_b1 , \3980_b0 );
or ( \3983_b1 , \3884_b1 , \3977_b1 );
xor ( \3983_b0 , \3884_b0 , w_6866 );
not ( w_6866 , w_6867 );
and ( w_6867 , \3977_b1 , \3977_b0 );
or ( \3984_b1 , \2927_A[15]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6868 );
and ( \3984_b0 , \2927_A[15]_b0 , w_6869 );
and ( w_6868 , w_6869 , \2991_B[11]_b0 );
or ( \3985_b1 , \3983_b1 , \3984_b1 );
not ( \3984_b1 , w_6870 );
and ( \3985_b0 , \3983_b0 , w_6871 );
and ( w_6870 , w_6871 , \3984_b0 );
or ( \3986_b1 , \3983_b1 , \3984_b1 );
xor ( \3986_b0 , \3983_b0 , w_6872 );
not ( w_6872 , w_6873 );
and ( w_6873 , \3984_b1 , \3984_b0 );
or ( \3987_b1 , \3888_b1 , \3975_b1 );
xor ( \3987_b0 , \3888_b0 , w_6874 );
not ( w_6874 , w_6875 );
and ( w_6875 , \3975_b1 , \3975_b0 );
or ( \3988_b1 , \2931_A[14]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6876 );
and ( \3988_b0 , \2931_A[14]_b0 , w_6877 );
and ( w_6876 , w_6877 , \2991_B[11]_b0 );
or ( \3989_b1 , \3987_b1 , \3988_b1 );
not ( \3988_b1 , w_6878 );
and ( \3989_b0 , \3987_b0 , w_6879 );
and ( w_6878 , w_6879 , \3988_b0 );
or ( \3990_b1 , \3987_b1 , \3988_b1 );
xor ( \3990_b0 , \3987_b0 , w_6880 );
not ( w_6880 , w_6881 );
and ( w_6881 , \3988_b1 , \3988_b0 );
or ( \3991_b1 , \3892_b1 , \3973_b1 );
xor ( \3991_b0 , \3892_b0 , w_6882 );
not ( w_6882 , w_6883 );
and ( w_6883 , \3973_b1 , \3973_b0 );
or ( \3992_b1 , \2935_A[13]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6884 );
and ( \3992_b0 , \2935_A[13]_b0 , w_6885 );
and ( w_6884 , w_6885 , \2991_B[11]_b0 );
or ( \3993_b1 , \3991_b1 , \3992_b1 );
not ( \3992_b1 , w_6886 );
and ( \3993_b0 , \3991_b0 , w_6887 );
and ( w_6886 , w_6887 , \3992_b0 );
or ( \3994_b1 , \3991_b1 , \3992_b1 );
xor ( \3994_b0 , \3991_b0 , w_6888 );
not ( w_6888 , w_6889 );
and ( w_6889 , \3992_b1 , \3992_b0 );
or ( \3995_b1 , \3896_b1 , \3971_b1 );
xor ( \3995_b0 , \3896_b0 , w_6890 );
not ( w_6890 , w_6891 );
and ( w_6891 , \3971_b1 , \3971_b0 );
or ( \3996_b1 , \2939_A[12]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6892 );
and ( \3996_b0 , \2939_A[12]_b0 , w_6893 );
and ( w_6892 , w_6893 , \2991_B[11]_b0 );
or ( \3997_b1 , \3995_b1 , \3996_b1 );
not ( \3996_b1 , w_6894 );
and ( \3997_b0 , \3995_b0 , w_6895 );
and ( w_6894 , w_6895 , \3996_b0 );
or ( \3998_b1 , \3995_b1 , \3996_b1 );
xor ( \3998_b0 , \3995_b0 , w_6896 );
not ( w_6896 , w_6897 );
and ( w_6897 , \3996_b1 , \3996_b0 );
or ( \3999_b1 , \3900_b1 , \3969_b1 );
xor ( \3999_b0 , \3900_b0 , w_6898 );
not ( w_6898 , w_6899 );
and ( w_6899 , \3969_b1 , \3969_b0 );
or ( \4000_b1 , \2943_A[11]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6900 );
and ( \4000_b0 , \2943_A[11]_b0 , w_6901 );
and ( w_6900 , w_6901 , \2991_B[11]_b0 );
or ( \4001_b1 , \3999_b1 , \4000_b1 );
not ( \4000_b1 , w_6902 );
and ( \4001_b0 , \3999_b0 , w_6903 );
and ( w_6902 , w_6903 , \4000_b0 );
or ( \4002_b1 , \3999_b1 , \4000_b1 );
xor ( \4002_b0 , \3999_b0 , w_6904 );
not ( w_6904 , w_6905 );
and ( w_6905 , \4000_b1 , \4000_b0 );
or ( \4003_b1 , \3904_b1 , \3967_b1 );
xor ( \4003_b0 , \3904_b0 , w_6906 );
not ( w_6906 , w_6907 );
and ( w_6907 , \3967_b1 , \3967_b0 );
or ( \4004_b1 , \2947_A[10]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6908 );
and ( \4004_b0 , \2947_A[10]_b0 , w_6909 );
and ( w_6908 , w_6909 , \2991_B[11]_b0 );
or ( \4005_b1 , \4003_b1 , \4004_b1 );
not ( \4004_b1 , w_6910 );
and ( \4005_b0 , \4003_b0 , w_6911 );
and ( w_6910 , w_6911 , \4004_b0 );
or ( \4006_b1 , \4003_b1 , \4004_b1 );
xor ( \4006_b0 , \4003_b0 , w_6912 );
not ( w_6912 , w_6913 );
and ( w_6913 , \4004_b1 , \4004_b0 );
or ( \4007_b1 , \3908_b1 , \3965_b1 );
xor ( \4007_b0 , \3908_b0 , w_6914 );
not ( w_6914 , w_6915 );
and ( w_6915 , \3965_b1 , \3965_b0 );
or ( \4008_b1 , \2951_A[9]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6916 );
and ( \4008_b0 , \2951_A[9]_b0 , w_6917 );
and ( w_6916 , w_6917 , \2991_B[11]_b0 );
or ( \4009_b1 , \4007_b1 , \4008_b1 );
not ( \4008_b1 , w_6918 );
and ( \4009_b0 , \4007_b0 , w_6919 );
and ( w_6918 , w_6919 , \4008_b0 );
or ( \4010_b1 , \4007_b1 , \4008_b1 );
xor ( \4010_b0 , \4007_b0 , w_6920 );
not ( w_6920 , w_6921 );
and ( w_6921 , \4008_b1 , \4008_b0 );
or ( \4011_b1 , \3912_b1 , \3963_b1 );
xor ( \4011_b0 , \3912_b0 , w_6922 );
not ( w_6922 , w_6923 );
and ( w_6923 , \3963_b1 , \3963_b0 );
or ( \4012_b1 , \2955_A[8]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6924 );
and ( \4012_b0 , \2955_A[8]_b0 , w_6925 );
and ( w_6924 , w_6925 , \2991_B[11]_b0 );
or ( \4013_b1 , \4011_b1 , \4012_b1 );
not ( \4012_b1 , w_6926 );
and ( \4013_b0 , \4011_b0 , w_6927 );
and ( w_6926 , w_6927 , \4012_b0 );
or ( \4014_b1 , \4011_b1 , \4012_b1 );
xor ( \4014_b0 , \4011_b0 , w_6928 );
not ( w_6928 , w_6929 );
and ( w_6929 , \4012_b1 , \4012_b0 );
or ( \4015_b1 , \3916_b1 , \3961_b1 );
xor ( \4015_b0 , \3916_b0 , w_6930 );
not ( w_6930 , w_6931 );
and ( w_6931 , \3961_b1 , \3961_b0 );
or ( \4016_b1 , \2959_A[7]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6932 );
and ( \4016_b0 , \2959_A[7]_b0 , w_6933 );
and ( w_6932 , w_6933 , \2991_B[11]_b0 );
or ( \4017_b1 , \4015_b1 , \4016_b1 );
not ( \4016_b1 , w_6934 );
and ( \4017_b0 , \4015_b0 , w_6935 );
and ( w_6934 , w_6935 , \4016_b0 );
or ( \4018_b1 , \4015_b1 , \4016_b1 );
xor ( \4018_b0 , \4015_b0 , w_6936 );
not ( w_6936 , w_6937 );
and ( w_6937 , \4016_b1 , \4016_b0 );
or ( \4019_b1 , \3920_b1 , \3959_b1 );
xor ( \4019_b0 , \3920_b0 , w_6938 );
not ( w_6938 , w_6939 );
and ( w_6939 , \3959_b1 , \3959_b0 );
or ( \4020_b1 , \2963_A[6]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6940 );
and ( \4020_b0 , \2963_A[6]_b0 , w_6941 );
and ( w_6940 , w_6941 , \2991_B[11]_b0 );
or ( \4021_b1 , \4019_b1 , \4020_b1 );
not ( \4020_b1 , w_6942 );
and ( \4021_b0 , \4019_b0 , w_6943 );
and ( w_6942 , w_6943 , \4020_b0 );
or ( \4022_b1 , \4019_b1 , \4020_b1 );
xor ( \4022_b0 , \4019_b0 , w_6944 );
not ( w_6944 , w_6945 );
and ( w_6945 , \4020_b1 , \4020_b0 );
or ( \4023_b1 , \3924_b1 , \3957_b1 );
xor ( \4023_b0 , \3924_b0 , w_6946 );
not ( w_6946 , w_6947 );
and ( w_6947 , \3957_b1 , \3957_b0 );
or ( \4024_b1 , \2967_A[5]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6948 );
and ( \4024_b0 , \2967_A[5]_b0 , w_6949 );
and ( w_6948 , w_6949 , \2991_B[11]_b0 );
or ( \4025_b1 , \4023_b1 , \4024_b1 );
not ( \4024_b1 , w_6950 );
and ( \4025_b0 , \4023_b0 , w_6951 );
and ( w_6950 , w_6951 , \4024_b0 );
or ( \4026_b1 , \4023_b1 , \4024_b1 );
xor ( \4026_b0 , \4023_b0 , w_6952 );
not ( w_6952 , w_6953 );
and ( w_6953 , \4024_b1 , \4024_b0 );
or ( \4027_b1 , \3928_b1 , \3955_b1 );
xor ( \4027_b0 , \3928_b0 , w_6954 );
not ( w_6954 , w_6955 );
and ( w_6955 , \3955_b1 , \3955_b0 );
or ( \4028_b1 , \2971_A[4]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6956 );
and ( \4028_b0 , \2971_A[4]_b0 , w_6957 );
and ( w_6956 , w_6957 , \2991_B[11]_b0 );
or ( \4029_b1 , \4027_b1 , \4028_b1 );
not ( \4028_b1 , w_6958 );
and ( \4029_b0 , \4027_b0 , w_6959 );
and ( w_6958 , w_6959 , \4028_b0 );
or ( \4030_b1 , \4027_b1 , \4028_b1 );
xor ( \4030_b0 , \4027_b0 , w_6960 );
not ( w_6960 , w_6961 );
and ( w_6961 , \4028_b1 , \4028_b0 );
or ( \4031_b1 , \3932_b1 , \3953_b1 );
xor ( \4031_b0 , \3932_b0 , w_6962 );
not ( w_6962 , w_6963 );
and ( w_6963 , \3953_b1 , \3953_b0 );
or ( \4032_b1 , \2975_A[3]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6964 );
and ( \4032_b0 , \2975_A[3]_b0 , w_6965 );
and ( w_6964 , w_6965 , \2991_B[11]_b0 );
or ( \4033_b1 , \4031_b1 , \4032_b1 );
not ( \4032_b1 , w_6966 );
and ( \4033_b0 , \4031_b0 , w_6967 );
and ( w_6966 , w_6967 , \4032_b0 );
or ( \4034_b1 , \4031_b1 , \4032_b1 );
xor ( \4034_b0 , \4031_b0 , w_6968 );
not ( w_6968 , w_6969 );
and ( w_6969 , \4032_b1 , \4032_b0 );
or ( \4035_b1 , \3936_b1 , \3951_b1 );
xor ( \4035_b0 , \3936_b0 , w_6970 );
not ( w_6970 , w_6971 );
and ( w_6971 , \3951_b1 , \3951_b0 );
or ( \4036_b1 , \2979_A[2]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6972 );
and ( \4036_b0 , \2979_A[2]_b0 , w_6973 );
and ( w_6972 , w_6973 , \2991_B[11]_b0 );
or ( \4037_b1 , \4035_b1 , \4036_b1 );
not ( \4036_b1 , w_6974 );
and ( \4037_b0 , \4035_b0 , w_6975 );
and ( w_6974 , w_6975 , \4036_b0 );
or ( \4038_b1 , \4035_b1 , \4036_b1 );
xor ( \4038_b0 , \4035_b0 , w_6976 );
not ( w_6976 , w_6977 );
and ( w_6977 , \4036_b1 , \4036_b0 );
or ( \4039_b1 , \3940_b1 , \3949_b1 );
xor ( \4039_b0 , \3940_b0 , w_6978 );
not ( w_6978 , w_6979 );
and ( w_6979 , \3949_b1 , \3949_b0 );
or ( \4040_b1 , \2983_A[1]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6980 );
and ( \4040_b0 , \2983_A[1]_b0 , w_6981 );
and ( w_6980 , w_6981 , \2991_B[11]_b0 );
or ( \4041_b1 , \4039_b1 , \4040_b1 );
not ( \4040_b1 , w_6982 );
and ( \4041_b0 , \4039_b0 , w_6983 );
and ( w_6982 , w_6983 , \4040_b0 );
or ( \4042_b1 , \4039_b1 , \4040_b1 );
xor ( \4042_b0 , \4039_b0 , w_6984 );
not ( w_6984 , w_6985 );
and ( w_6985 , \4040_b1 , \4040_b0 );
or ( \4043_b1 , \3944_b1 , \3947_b1 );
xor ( \4043_b0 , \3944_b0 , w_6986 );
not ( w_6986 , w_6987 );
and ( w_6987 , \3947_b1 , \3947_b0 );
or ( \4044_b1 , \2986_A[0]_b1 , \2991_B[11]_b1 );
not ( \2991_B[11]_b1 , w_6988 );
and ( \4044_b0 , \2986_A[0]_b0 , w_6989 );
and ( w_6988 , w_6989 , \2991_B[11]_b0 );
or ( \4045_b1 , \4043_b1 , \4044_b1 );
not ( \4044_b1 , w_6990 );
and ( \4045_b0 , \4043_b0 , w_6991 );
and ( w_6990 , w_6991 , \4044_b0 );
or ( \4046_b1 , \4042_b1 , \4045_b1 );
not ( \4045_b1 , w_6992 );
and ( \4046_b0 , \4042_b0 , w_6993 );
and ( w_6992 , w_6993 , \4045_b0 );
or ( \4047_b1 , \4041_b1 , w_6994 );
or ( \4047_b0 , \4041_b0 , \4046_b0 );
not ( \4046_b0 , w_6995 );
and ( w_6995 , w_6994 , \4046_b1 );
or ( \4048_b1 , \4038_b1 , \4047_b1 );
not ( \4047_b1 , w_6996 );
and ( \4048_b0 , \4038_b0 , w_6997 );
and ( w_6996 , w_6997 , \4047_b0 );
or ( \4049_b1 , \4037_b1 , w_6998 );
or ( \4049_b0 , \4037_b0 , \4048_b0 );
not ( \4048_b0 , w_6999 );
and ( w_6999 , w_6998 , \4048_b1 );
or ( \4050_b1 , \4034_b1 , \4049_b1 );
not ( \4049_b1 , w_7000 );
and ( \4050_b0 , \4034_b0 , w_7001 );
and ( w_7000 , w_7001 , \4049_b0 );
or ( \4051_b1 , \4033_b1 , w_7002 );
or ( \4051_b0 , \4033_b0 , \4050_b0 );
not ( \4050_b0 , w_7003 );
and ( w_7003 , w_7002 , \4050_b1 );
or ( \4052_b1 , \4030_b1 , \4051_b1 );
not ( \4051_b1 , w_7004 );
and ( \4052_b0 , \4030_b0 , w_7005 );
and ( w_7004 , w_7005 , \4051_b0 );
or ( \4053_b1 , \4029_b1 , w_7006 );
or ( \4053_b0 , \4029_b0 , \4052_b0 );
not ( \4052_b0 , w_7007 );
and ( w_7007 , w_7006 , \4052_b1 );
or ( \4054_b1 , \4026_b1 , \4053_b1 );
not ( \4053_b1 , w_7008 );
and ( \4054_b0 , \4026_b0 , w_7009 );
and ( w_7008 , w_7009 , \4053_b0 );
or ( \4055_b1 , \4025_b1 , w_7010 );
or ( \4055_b0 , \4025_b0 , \4054_b0 );
not ( \4054_b0 , w_7011 );
and ( w_7011 , w_7010 , \4054_b1 );
or ( \4056_b1 , \4022_b1 , \4055_b1 );
not ( \4055_b1 , w_7012 );
and ( \4056_b0 , \4022_b0 , w_7013 );
and ( w_7012 , w_7013 , \4055_b0 );
or ( \4057_b1 , \4021_b1 , w_7014 );
or ( \4057_b0 , \4021_b0 , \4056_b0 );
not ( \4056_b0 , w_7015 );
and ( w_7015 , w_7014 , \4056_b1 );
or ( \4058_b1 , \4018_b1 , \4057_b1 );
not ( \4057_b1 , w_7016 );
and ( \4058_b0 , \4018_b0 , w_7017 );
and ( w_7016 , w_7017 , \4057_b0 );
or ( \4059_b1 , \4017_b1 , w_7018 );
or ( \4059_b0 , \4017_b0 , \4058_b0 );
not ( \4058_b0 , w_7019 );
and ( w_7019 , w_7018 , \4058_b1 );
or ( \4060_b1 , \4014_b1 , \4059_b1 );
not ( \4059_b1 , w_7020 );
and ( \4060_b0 , \4014_b0 , w_7021 );
and ( w_7020 , w_7021 , \4059_b0 );
or ( \4061_b1 , \4013_b1 , w_7022 );
or ( \4061_b0 , \4013_b0 , \4060_b0 );
not ( \4060_b0 , w_7023 );
and ( w_7023 , w_7022 , \4060_b1 );
or ( \4062_b1 , \4010_b1 , \4061_b1 );
not ( \4061_b1 , w_7024 );
and ( \4062_b0 , \4010_b0 , w_7025 );
and ( w_7024 , w_7025 , \4061_b0 );
or ( \4063_b1 , \4009_b1 , w_7026 );
or ( \4063_b0 , \4009_b0 , \4062_b0 );
not ( \4062_b0 , w_7027 );
and ( w_7027 , w_7026 , \4062_b1 );
or ( \4064_b1 , \4006_b1 , \4063_b1 );
not ( \4063_b1 , w_7028 );
and ( \4064_b0 , \4006_b0 , w_7029 );
and ( w_7028 , w_7029 , \4063_b0 );
or ( \4065_b1 , \4005_b1 , w_7030 );
or ( \4065_b0 , \4005_b0 , \4064_b0 );
not ( \4064_b0 , w_7031 );
and ( w_7031 , w_7030 , \4064_b1 );
or ( \4066_b1 , \4002_b1 , \4065_b1 );
not ( \4065_b1 , w_7032 );
and ( \4066_b0 , \4002_b0 , w_7033 );
and ( w_7032 , w_7033 , \4065_b0 );
or ( \4067_b1 , \4001_b1 , w_7034 );
or ( \4067_b0 , \4001_b0 , \4066_b0 );
not ( \4066_b0 , w_7035 );
and ( w_7035 , w_7034 , \4066_b1 );
or ( \4068_b1 , \3998_b1 , \4067_b1 );
not ( \4067_b1 , w_7036 );
and ( \4068_b0 , \3998_b0 , w_7037 );
and ( w_7036 , w_7037 , \4067_b0 );
or ( \4069_b1 , \3997_b1 , w_7038 );
or ( \4069_b0 , \3997_b0 , \4068_b0 );
not ( \4068_b0 , w_7039 );
and ( w_7039 , w_7038 , \4068_b1 );
or ( \4070_b1 , \3994_b1 , \4069_b1 );
not ( \4069_b1 , w_7040 );
and ( \4070_b0 , \3994_b0 , w_7041 );
and ( w_7040 , w_7041 , \4069_b0 );
or ( \4071_b1 , \3993_b1 , w_7042 );
or ( \4071_b0 , \3993_b0 , \4070_b0 );
not ( \4070_b0 , w_7043 );
and ( w_7043 , w_7042 , \4070_b1 );
or ( \4072_b1 , \3990_b1 , \4071_b1 );
not ( \4071_b1 , w_7044 );
and ( \4072_b0 , \3990_b0 , w_7045 );
and ( w_7044 , w_7045 , \4071_b0 );
or ( \4073_b1 , \3989_b1 , w_7046 );
or ( \4073_b0 , \3989_b0 , \4072_b0 );
not ( \4072_b0 , w_7047 );
and ( w_7047 , w_7046 , \4072_b1 );
or ( \4074_b1 , \3986_b1 , \4073_b1 );
not ( \4073_b1 , w_7048 );
and ( \4074_b0 , \3986_b0 , w_7049 );
and ( w_7048 , w_7049 , \4073_b0 );
or ( \4075_b1 , \3985_b1 , w_7050 );
or ( \4075_b0 , \3985_b0 , \4074_b0 );
not ( \4074_b0 , w_7051 );
and ( w_7051 , w_7050 , \4074_b1 );
or ( \4076_b1 , \3982_b1 , \4075_b1 );
not ( \4075_b1 , w_7052 );
and ( \4076_b0 , \3982_b0 , w_7053 );
and ( w_7052 , w_7053 , \4075_b0 );
or ( \4077_b1 , \3981_b1 , w_7054 );
or ( \4077_b0 , \3981_b0 , \4076_b0 );
not ( \4076_b0 , w_7055 );
and ( w_7055 , w_7054 , \4076_b1 );
or ( \4078_b1 , \2923_A[16]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7056 );
and ( \4078_b0 , \2923_A[16]_b0 , w_7057 );
and ( w_7056 , w_7057 , \2990_B[12]_b0 );
or ( \4079_b1 , \4077_b1 , \4078_b1 );
not ( \4078_b1 , w_7058 );
and ( \4079_b0 , \4077_b0 , w_7059 );
and ( w_7058 , w_7059 , \4078_b0 );
or ( \4080_b1 , \4077_b1 , \4078_b1 );
xor ( \4080_b0 , \4077_b0 , w_7060 );
not ( w_7060 , w_7061 );
and ( w_7061 , \4078_b1 , \4078_b0 );
or ( \4081_b1 , \3982_b1 , \4075_b1 );
xor ( \4081_b0 , \3982_b0 , w_7062 );
not ( w_7062 , w_7063 );
and ( w_7063 , \4075_b1 , \4075_b0 );
or ( \4082_b1 , \2927_A[15]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7064 );
and ( \4082_b0 , \2927_A[15]_b0 , w_7065 );
and ( w_7064 , w_7065 , \2990_B[12]_b0 );
or ( \4083_b1 , \4081_b1 , \4082_b1 );
not ( \4082_b1 , w_7066 );
and ( \4083_b0 , \4081_b0 , w_7067 );
and ( w_7066 , w_7067 , \4082_b0 );
or ( \4084_b1 , \4081_b1 , \4082_b1 );
xor ( \4084_b0 , \4081_b0 , w_7068 );
not ( w_7068 , w_7069 );
and ( w_7069 , \4082_b1 , \4082_b0 );
or ( \4085_b1 , \3986_b1 , \4073_b1 );
xor ( \4085_b0 , \3986_b0 , w_7070 );
not ( w_7070 , w_7071 );
and ( w_7071 , \4073_b1 , \4073_b0 );
or ( \4086_b1 , \2931_A[14]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7072 );
and ( \4086_b0 , \2931_A[14]_b0 , w_7073 );
and ( w_7072 , w_7073 , \2990_B[12]_b0 );
or ( \4087_b1 , \4085_b1 , \4086_b1 );
not ( \4086_b1 , w_7074 );
and ( \4087_b0 , \4085_b0 , w_7075 );
and ( w_7074 , w_7075 , \4086_b0 );
or ( \4088_b1 , \4085_b1 , \4086_b1 );
xor ( \4088_b0 , \4085_b0 , w_7076 );
not ( w_7076 , w_7077 );
and ( w_7077 , \4086_b1 , \4086_b0 );
or ( \4089_b1 , \3990_b1 , \4071_b1 );
xor ( \4089_b0 , \3990_b0 , w_7078 );
not ( w_7078 , w_7079 );
and ( w_7079 , \4071_b1 , \4071_b0 );
or ( \4090_b1 , \2935_A[13]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7080 );
and ( \4090_b0 , \2935_A[13]_b0 , w_7081 );
and ( w_7080 , w_7081 , \2990_B[12]_b0 );
or ( \4091_b1 , \4089_b1 , \4090_b1 );
not ( \4090_b1 , w_7082 );
and ( \4091_b0 , \4089_b0 , w_7083 );
and ( w_7082 , w_7083 , \4090_b0 );
or ( \4092_b1 , \4089_b1 , \4090_b1 );
xor ( \4092_b0 , \4089_b0 , w_7084 );
not ( w_7084 , w_7085 );
and ( w_7085 , \4090_b1 , \4090_b0 );
or ( \4093_b1 , \3994_b1 , \4069_b1 );
xor ( \4093_b0 , \3994_b0 , w_7086 );
not ( w_7086 , w_7087 );
and ( w_7087 , \4069_b1 , \4069_b0 );
or ( \4094_b1 , \2939_A[12]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7088 );
and ( \4094_b0 , \2939_A[12]_b0 , w_7089 );
and ( w_7088 , w_7089 , \2990_B[12]_b0 );
or ( \4095_b1 , \4093_b1 , \4094_b1 );
not ( \4094_b1 , w_7090 );
and ( \4095_b0 , \4093_b0 , w_7091 );
and ( w_7090 , w_7091 , \4094_b0 );
or ( \4096_b1 , \4093_b1 , \4094_b1 );
xor ( \4096_b0 , \4093_b0 , w_7092 );
not ( w_7092 , w_7093 );
and ( w_7093 , \4094_b1 , \4094_b0 );
or ( \4097_b1 , \3998_b1 , \4067_b1 );
xor ( \4097_b0 , \3998_b0 , w_7094 );
not ( w_7094 , w_7095 );
and ( w_7095 , \4067_b1 , \4067_b0 );
or ( \4098_b1 , \2943_A[11]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7096 );
and ( \4098_b0 , \2943_A[11]_b0 , w_7097 );
and ( w_7096 , w_7097 , \2990_B[12]_b0 );
or ( \4099_b1 , \4097_b1 , \4098_b1 );
not ( \4098_b1 , w_7098 );
and ( \4099_b0 , \4097_b0 , w_7099 );
and ( w_7098 , w_7099 , \4098_b0 );
or ( \4100_b1 , \4097_b1 , \4098_b1 );
xor ( \4100_b0 , \4097_b0 , w_7100 );
not ( w_7100 , w_7101 );
and ( w_7101 , \4098_b1 , \4098_b0 );
or ( \4101_b1 , \4002_b1 , \4065_b1 );
xor ( \4101_b0 , \4002_b0 , w_7102 );
not ( w_7102 , w_7103 );
and ( w_7103 , \4065_b1 , \4065_b0 );
or ( \4102_b1 , \2947_A[10]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7104 );
and ( \4102_b0 , \2947_A[10]_b0 , w_7105 );
and ( w_7104 , w_7105 , \2990_B[12]_b0 );
or ( \4103_b1 , \4101_b1 , \4102_b1 );
not ( \4102_b1 , w_7106 );
and ( \4103_b0 , \4101_b0 , w_7107 );
and ( w_7106 , w_7107 , \4102_b0 );
or ( \4104_b1 , \4101_b1 , \4102_b1 );
xor ( \4104_b0 , \4101_b0 , w_7108 );
not ( w_7108 , w_7109 );
and ( w_7109 , \4102_b1 , \4102_b0 );
or ( \4105_b1 , \4006_b1 , \4063_b1 );
xor ( \4105_b0 , \4006_b0 , w_7110 );
not ( w_7110 , w_7111 );
and ( w_7111 , \4063_b1 , \4063_b0 );
or ( \4106_b1 , \2951_A[9]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7112 );
and ( \4106_b0 , \2951_A[9]_b0 , w_7113 );
and ( w_7112 , w_7113 , \2990_B[12]_b0 );
or ( \4107_b1 , \4105_b1 , \4106_b1 );
not ( \4106_b1 , w_7114 );
and ( \4107_b0 , \4105_b0 , w_7115 );
and ( w_7114 , w_7115 , \4106_b0 );
or ( \4108_b1 , \4105_b1 , \4106_b1 );
xor ( \4108_b0 , \4105_b0 , w_7116 );
not ( w_7116 , w_7117 );
and ( w_7117 , \4106_b1 , \4106_b0 );
or ( \4109_b1 , \4010_b1 , \4061_b1 );
xor ( \4109_b0 , \4010_b0 , w_7118 );
not ( w_7118 , w_7119 );
and ( w_7119 , \4061_b1 , \4061_b0 );
or ( \4110_b1 , \2955_A[8]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7120 );
and ( \4110_b0 , \2955_A[8]_b0 , w_7121 );
and ( w_7120 , w_7121 , \2990_B[12]_b0 );
or ( \4111_b1 , \4109_b1 , \4110_b1 );
not ( \4110_b1 , w_7122 );
and ( \4111_b0 , \4109_b0 , w_7123 );
and ( w_7122 , w_7123 , \4110_b0 );
or ( \4112_b1 , \4109_b1 , \4110_b1 );
xor ( \4112_b0 , \4109_b0 , w_7124 );
not ( w_7124 , w_7125 );
and ( w_7125 , \4110_b1 , \4110_b0 );
or ( \4113_b1 , \4014_b1 , \4059_b1 );
xor ( \4113_b0 , \4014_b0 , w_7126 );
not ( w_7126 , w_7127 );
and ( w_7127 , \4059_b1 , \4059_b0 );
or ( \4114_b1 , \2959_A[7]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7128 );
and ( \4114_b0 , \2959_A[7]_b0 , w_7129 );
and ( w_7128 , w_7129 , \2990_B[12]_b0 );
or ( \4115_b1 , \4113_b1 , \4114_b1 );
not ( \4114_b1 , w_7130 );
and ( \4115_b0 , \4113_b0 , w_7131 );
and ( w_7130 , w_7131 , \4114_b0 );
or ( \4116_b1 , \4113_b1 , \4114_b1 );
xor ( \4116_b0 , \4113_b0 , w_7132 );
not ( w_7132 , w_7133 );
and ( w_7133 , \4114_b1 , \4114_b0 );
or ( \4117_b1 , \4018_b1 , \4057_b1 );
xor ( \4117_b0 , \4018_b0 , w_7134 );
not ( w_7134 , w_7135 );
and ( w_7135 , \4057_b1 , \4057_b0 );
or ( \4118_b1 , \2963_A[6]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7136 );
and ( \4118_b0 , \2963_A[6]_b0 , w_7137 );
and ( w_7136 , w_7137 , \2990_B[12]_b0 );
or ( \4119_b1 , \4117_b1 , \4118_b1 );
not ( \4118_b1 , w_7138 );
and ( \4119_b0 , \4117_b0 , w_7139 );
and ( w_7138 , w_7139 , \4118_b0 );
or ( \4120_b1 , \4117_b1 , \4118_b1 );
xor ( \4120_b0 , \4117_b0 , w_7140 );
not ( w_7140 , w_7141 );
and ( w_7141 , \4118_b1 , \4118_b0 );
or ( \4121_b1 , \4022_b1 , \4055_b1 );
xor ( \4121_b0 , \4022_b0 , w_7142 );
not ( w_7142 , w_7143 );
and ( w_7143 , \4055_b1 , \4055_b0 );
or ( \4122_b1 , \2967_A[5]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7144 );
and ( \4122_b0 , \2967_A[5]_b0 , w_7145 );
and ( w_7144 , w_7145 , \2990_B[12]_b0 );
or ( \4123_b1 , \4121_b1 , \4122_b1 );
not ( \4122_b1 , w_7146 );
and ( \4123_b0 , \4121_b0 , w_7147 );
and ( w_7146 , w_7147 , \4122_b0 );
or ( \4124_b1 , \4121_b1 , \4122_b1 );
xor ( \4124_b0 , \4121_b0 , w_7148 );
not ( w_7148 , w_7149 );
and ( w_7149 , \4122_b1 , \4122_b0 );
or ( \4125_b1 , \4026_b1 , \4053_b1 );
xor ( \4125_b0 , \4026_b0 , w_7150 );
not ( w_7150 , w_7151 );
and ( w_7151 , \4053_b1 , \4053_b0 );
or ( \4126_b1 , \2971_A[4]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7152 );
and ( \4126_b0 , \2971_A[4]_b0 , w_7153 );
and ( w_7152 , w_7153 , \2990_B[12]_b0 );
or ( \4127_b1 , \4125_b1 , \4126_b1 );
not ( \4126_b1 , w_7154 );
and ( \4127_b0 , \4125_b0 , w_7155 );
and ( w_7154 , w_7155 , \4126_b0 );
or ( \4128_b1 , \4125_b1 , \4126_b1 );
xor ( \4128_b0 , \4125_b0 , w_7156 );
not ( w_7156 , w_7157 );
and ( w_7157 , \4126_b1 , \4126_b0 );
or ( \4129_b1 , \4030_b1 , \4051_b1 );
xor ( \4129_b0 , \4030_b0 , w_7158 );
not ( w_7158 , w_7159 );
and ( w_7159 , \4051_b1 , \4051_b0 );
or ( \4130_b1 , \2975_A[3]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7160 );
and ( \4130_b0 , \2975_A[3]_b0 , w_7161 );
and ( w_7160 , w_7161 , \2990_B[12]_b0 );
or ( \4131_b1 , \4129_b1 , \4130_b1 );
not ( \4130_b1 , w_7162 );
and ( \4131_b0 , \4129_b0 , w_7163 );
and ( w_7162 , w_7163 , \4130_b0 );
or ( \4132_b1 , \4129_b1 , \4130_b1 );
xor ( \4132_b0 , \4129_b0 , w_7164 );
not ( w_7164 , w_7165 );
and ( w_7165 , \4130_b1 , \4130_b0 );
or ( \4133_b1 , \4034_b1 , \4049_b1 );
xor ( \4133_b0 , \4034_b0 , w_7166 );
not ( w_7166 , w_7167 );
and ( w_7167 , \4049_b1 , \4049_b0 );
or ( \4134_b1 , \2979_A[2]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7168 );
and ( \4134_b0 , \2979_A[2]_b0 , w_7169 );
and ( w_7168 , w_7169 , \2990_B[12]_b0 );
or ( \4135_b1 , \4133_b1 , \4134_b1 );
not ( \4134_b1 , w_7170 );
and ( \4135_b0 , \4133_b0 , w_7171 );
and ( w_7170 , w_7171 , \4134_b0 );
or ( \4136_b1 , \4133_b1 , \4134_b1 );
xor ( \4136_b0 , \4133_b0 , w_7172 );
not ( w_7172 , w_7173 );
and ( w_7173 , \4134_b1 , \4134_b0 );
or ( \4137_b1 , \4038_b1 , \4047_b1 );
xor ( \4137_b0 , \4038_b0 , w_7174 );
not ( w_7174 , w_7175 );
and ( w_7175 , \4047_b1 , \4047_b0 );
or ( \4138_b1 , \2983_A[1]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7176 );
and ( \4138_b0 , \2983_A[1]_b0 , w_7177 );
and ( w_7176 , w_7177 , \2990_B[12]_b0 );
or ( \4139_b1 , \4137_b1 , \4138_b1 );
not ( \4138_b1 , w_7178 );
and ( \4139_b0 , \4137_b0 , w_7179 );
and ( w_7178 , w_7179 , \4138_b0 );
or ( \4140_b1 , \4137_b1 , \4138_b1 );
xor ( \4140_b0 , \4137_b0 , w_7180 );
not ( w_7180 , w_7181 );
and ( w_7181 , \4138_b1 , \4138_b0 );
or ( \4141_b1 , \4042_b1 , \4045_b1 );
xor ( \4141_b0 , \4042_b0 , w_7182 );
not ( w_7182 , w_7183 );
and ( w_7183 , \4045_b1 , \4045_b0 );
or ( \4142_b1 , \2986_A[0]_b1 , \2990_B[12]_b1 );
not ( \2990_B[12]_b1 , w_7184 );
and ( \4142_b0 , \2986_A[0]_b0 , w_7185 );
and ( w_7184 , w_7185 , \2990_B[12]_b0 );
or ( \4143_b1 , \4141_b1 , \4142_b1 );
not ( \4142_b1 , w_7186 );
and ( \4143_b0 , \4141_b0 , w_7187 );
and ( w_7186 , w_7187 , \4142_b0 );
or ( \4144_b1 , \4140_b1 , \4143_b1 );
not ( \4143_b1 , w_7188 );
and ( \4144_b0 , \4140_b0 , w_7189 );
and ( w_7188 , w_7189 , \4143_b0 );
or ( \4145_b1 , \4139_b1 , w_7190 );
or ( \4145_b0 , \4139_b0 , \4144_b0 );
not ( \4144_b0 , w_7191 );
and ( w_7191 , w_7190 , \4144_b1 );
or ( \4146_b1 , \4136_b1 , \4145_b1 );
not ( \4145_b1 , w_7192 );
and ( \4146_b0 , \4136_b0 , w_7193 );
and ( w_7192 , w_7193 , \4145_b0 );
or ( \4147_b1 , \4135_b1 , w_7194 );
or ( \4147_b0 , \4135_b0 , \4146_b0 );
not ( \4146_b0 , w_7195 );
and ( w_7195 , w_7194 , \4146_b1 );
or ( \4148_b1 , \4132_b1 , \4147_b1 );
not ( \4147_b1 , w_7196 );
and ( \4148_b0 , \4132_b0 , w_7197 );
and ( w_7196 , w_7197 , \4147_b0 );
or ( \4149_b1 , \4131_b1 , w_7198 );
or ( \4149_b0 , \4131_b0 , \4148_b0 );
not ( \4148_b0 , w_7199 );
and ( w_7199 , w_7198 , \4148_b1 );
or ( \4150_b1 , \4128_b1 , \4149_b1 );
not ( \4149_b1 , w_7200 );
and ( \4150_b0 , \4128_b0 , w_7201 );
and ( w_7200 , w_7201 , \4149_b0 );
or ( \4151_b1 , \4127_b1 , w_7202 );
or ( \4151_b0 , \4127_b0 , \4150_b0 );
not ( \4150_b0 , w_7203 );
and ( w_7203 , w_7202 , \4150_b1 );
or ( \4152_b1 , \4124_b1 , \4151_b1 );
not ( \4151_b1 , w_7204 );
and ( \4152_b0 , \4124_b0 , w_7205 );
and ( w_7204 , w_7205 , \4151_b0 );
or ( \4153_b1 , \4123_b1 , w_7206 );
or ( \4153_b0 , \4123_b0 , \4152_b0 );
not ( \4152_b0 , w_7207 );
and ( w_7207 , w_7206 , \4152_b1 );
or ( \4154_b1 , \4120_b1 , \4153_b1 );
not ( \4153_b1 , w_7208 );
and ( \4154_b0 , \4120_b0 , w_7209 );
and ( w_7208 , w_7209 , \4153_b0 );
or ( \4155_b1 , \4119_b1 , w_7210 );
or ( \4155_b0 , \4119_b0 , \4154_b0 );
not ( \4154_b0 , w_7211 );
and ( w_7211 , w_7210 , \4154_b1 );
or ( \4156_b1 , \4116_b1 , \4155_b1 );
not ( \4155_b1 , w_7212 );
and ( \4156_b0 , \4116_b0 , w_7213 );
and ( w_7212 , w_7213 , \4155_b0 );
or ( \4157_b1 , \4115_b1 , w_7214 );
or ( \4157_b0 , \4115_b0 , \4156_b0 );
not ( \4156_b0 , w_7215 );
and ( w_7215 , w_7214 , \4156_b1 );
or ( \4158_b1 , \4112_b1 , \4157_b1 );
not ( \4157_b1 , w_7216 );
and ( \4158_b0 , \4112_b0 , w_7217 );
and ( w_7216 , w_7217 , \4157_b0 );
or ( \4159_b1 , \4111_b1 , w_7218 );
or ( \4159_b0 , \4111_b0 , \4158_b0 );
not ( \4158_b0 , w_7219 );
and ( w_7219 , w_7218 , \4158_b1 );
or ( \4160_b1 , \4108_b1 , \4159_b1 );
not ( \4159_b1 , w_7220 );
and ( \4160_b0 , \4108_b0 , w_7221 );
and ( w_7220 , w_7221 , \4159_b0 );
or ( \4161_b1 , \4107_b1 , w_7222 );
or ( \4161_b0 , \4107_b0 , \4160_b0 );
not ( \4160_b0 , w_7223 );
and ( w_7223 , w_7222 , \4160_b1 );
or ( \4162_b1 , \4104_b1 , \4161_b1 );
not ( \4161_b1 , w_7224 );
and ( \4162_b0 , \4104_b0 , w_7225 );
and ( w_7224 , w_7225 , \4161_b0 );
or ( \4163_b1 , \4103_b1 , w_7226 );
or ( \4163_b0 , \4103_b0 , \4162_b0 );
not ( \4162_b0 , w_7227 );
and ( w_7227 , w_7226 , \4162_b1 );
or ( \4164_b1 , \4100_b1 , \4163_b1 );
not ( \4163_b1 , w_7228 );
and ( \4164_b0 , \4100_b0 , w_7229 );
and ( w_7228 , w_7229 , \4163_b0 );
or ( \4165_b1 , \4099_b1 , w_7230 );
or ( \4165_b0 , \4099_b0 , \4164_b0 );
not ( \4164_b0 , w_7231 );
and ( w_7231 , w_7230 , \4164_b1 );
or ( \4166_b1 , \4096_b1 , \4165_b1 );
not ( \4165_b1 , w_7232 );
and ( \4166_b0 , \4096_b0 , w_7233 );
and ( w_7232 , w_7233 , \4165_b0 );
or ( \4167_b1 , \4095_b1 , w_7234 );
or ( \4167_b0 , \4095_b0 , \4166_b0 );
not ( \4166_b0 , w_7235 );
and ( w_7235 , w_7234 , \4166_b1 );
or ( \4168_b1 , \4092_b1 , \4167_b1 );
not ( \4167_b1 , w_7236 );
and ( \4168_b0 , \4092_b0 , w_7237 );
and ( w_7236 , w_7237 , \4167_b0 );
or ( \4169_b1 , \4091_b1 , w_7238 );
or ( \4169_b0 , \4091_b0 , \4168_b0 );
not ( \4168_b0 , w_7239 );
and ( w_7239 , w_7238 , \4168_b1 );
or ( \4170_b1 , \4088_b1 , \4169_b1 );
not ( \4169_b1 , w_7240 );
and ( \4170_b0 , \4088_b0 , w_7241 );
and ( w_7240 , w_7241 , \4169_b0 );
or ( \4171_b1 , \4087_b1 , w_7242 );
or ( \4171_b0 , \4087_b0 , \4170_b0 );
not ( \4170_b0 , w_7243 );
and ( w_7243 , w_7242 , \4170_b1 );
or ( \4172_b1 , \4084_b1 , \4171_b1 );
not ( \4171_b1 , w_7244 );
and ( \4172_b0 , \4084_b0 , w_7245 );
and ( w_7244 , w_7245 , \4171_b0 );
or ( \4173_b1 , \4083_b1 , w_7246 );
or ( \4173_b0 , \4083_b0 , \4172_b0 );
not ( \4172_b0 , w_7247 );
and ( w_7247 , w_7246 , \4172_b1 );
or ( \4174_b1 , \4080_b1 , \4173_b1 );
not ( \4173_b1 , w_7248 );
and ( \4174_b0 , \4080_b0 , w_7249 );
and ( w_7248 , w_7249 , \4173_b0 );
or ( \4175_b1 , \4079_b1 , w_7250 );
or ( \4175_b0 , \4079_b0 , \4174_b0 );
not ( \4174_b0 , w_7251 );
and ( w_7251 , w_7250 , \4174_b1 );
or ( \4176_b1 , \2923_A[16]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7252 );
and ( \4176_b0 , \2923_A[16]_b0 , w_7253 );
and ( w_7252 , w_7253 , \2989_B[13]_b0 );
or ( \4177_b1 , \4175_b1 , \4176_b1 );
not ( \4176_b1 , w_7254 );
and ( \4177_b0 , \4175_b0 , w_7255 );
and ( w_7254 , w_7255 , \4176_b0 );
or ( \4178_b1 , \4175_b1 , \4176_b1 );
xor ( \4178_b0 , \4175_b0 , w_7256 );
not ( w_7256 , w_7257 );
and ( w_7257 , \4176_b1 , \4176_b0 );
or ( \4179_b1 , \4080_b1 , \4173_b1 );
xor ( \4179_b0 , \4080_b0 , w_7258 );
not ( w_7258 , w_7259 );
and ( w_7259 , \4173_b1 , \4173_b0 );
or ( \4180_b1 , \2927_A[15]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7260 );
and ( \4180_b0 , \2927_A[15]_b0 , w_7261 );
and ( w_7260 , w_7261 , \2989_B[13]_b0 );
or ( \4181_b1 , \4179_b1 , \4180_b1 );
not ( \4180_b1 , w_7262 );
and ( \4181_b0 , \4179_b0 , w_7263 );
and ( w_7262 , w_7263 , \4180_b0 );
or ( \4182_b1 , \4179_b1 , \4180_b1 );
xor ( \4182_b0 , \4179_b0 , w_7264 );
not ( w_7264 , w_7265 );
and ( w_7265 , \4180_b1 , \4180_b0 );
or ( \4183_b1 , \4084_b1 , \4171_b1 );
xor ( \4183_b0 , \4084_b0 , w_7266 );
not ( w_7266 , w_7267 );
and ( w_7267 , \4171_b1 , \4171_b0 );
or ( \4184_b1 , \2931_A[14]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7268 );
and ( \4184_b0 , \2931_A[14]_b0 , w_7269 );
and ( w_7268 , w_7269 , \2989_B[13]_b0 );
or ( \4185_b1 , \4183_b1 , \4184_b1 );
not ( \4184_b1 , w_7270 );
and ( \4185_b0 , \4183_b0 , w_7271 );
and ( w_7270 , w_7271 , \4184_b0 );
or ( \4186_b1 , \4183_b1 , \4184_b1 );
xor ( \4186_b0 , \4183_b0 , w_7272 );
not ( w_7272 , w_7273 );
and ( w_7273 , \4184_b1 , \4184_b0 );
or ( \4187_b1 , \4088_b1 , \4169_b1 );
xor ( \4187_b0 , \4088_b0 , w_7274 );
not ( w_7274 , w_7275 );
and ( w_7275 , \4169_b1 , \4169_b0 );
or ( \4188_b1 , \2935_A[13]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7276 );
and ( \4188_b0 , \2935_A[13]_b0 , w_7277 );
and ( w_7276 , w_7277 , \2989_B[13]_b0 );
or ( \4189_b1 , \4187_b1 , \4188_b1 );
not ( \4188_b1 , w_7278 );
and ( \4189_b0 , \4187_b0 , w_7279 );
and ( w_7278 , w_7279 , \4188_b0 );
or ( \4190_b1 , \4187_b1 , \4188_b1 );
xor ( \4190_b0 , \4187_b0 , w_7280 );
not ( w_7280 , w_7281 );
and ( w_7281 , \4188_b1 , \4188_b0 );
or ( \4191_b1 , \4092_b1 , \4167_b1 );
xor ( \4191_b0 , \4092_b0 , w_7282 );
not ( w_7282 , w_7283 );
and ( w_7283 , \4167_b1 , \4167_b0 );
or ( \4192_b1 , \2939_A[12]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7284 );
and ( \4192_b0 , \2939_A[12]_b0 , w_7285 );
and ( w_7284 , w_7285 , \2989_B[13]_b0 );
or ( \4193_b1 , \4191_b1 , \4192_b1 );
not ( \4192_b1 , w_7286 );
and ( \4193_b0 , \4191_b0 , w_7287 );
and ( w_7286 , w_7287 , \4192_b0 );
or ( \4194_b1 , \4191_b1 , \4192_b1 );
xor ( \4194_b0 , \4191_b0 , w_7288 );
not ( w_7288 , w_7289 );
and ( w_7289 , \4192_b1 , \4192_b0 );
or ( \4195_b1 , \4096_b1 , \4165_b1 );
xor ( \4195_b0 , \4096_b0 , w_7290 );
not ( w_7290 , w_7291 );
and ( w_7291 , \4165_b1 , \4165_b0 );
or ( \4196_b1 , \2943_A[11]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7292 );
and ( \4196_b0 , \2943_A[11]_b0 , w_7293 );
and ( w_7292 , w_7293 , \2989_B[13]_b0 );
or ( \4197_b1 , \4195_b1 , \4196_b1 );
not ( \4196_b1 , w_7294 );
and ( \4197_b0 , \4195_b0 , w_7295 );
and ( w_7294 , w_7295 , \4196_b0 );
or ( \4198_b1 , \4195_b1 , \4196_b1 );
xor ( \4198_b0 , \4195_b0 , w_7296 );
not ( w_7296 , w_7297 );
and ( w_7297 , \4196_b1 , \4196_b0 );
or ( \4199_b1 , \4100_b1 , \4163_b1 );
xor ( \4199_b0 , \4100_b0 , w_7298 );
not ( w_7298 , w_7299 );
and ( w_7299 , \4163_b1 , \4163_b0 );
or ( \4200_b1 , \2947_A[10]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7300 );
and ( \4200_b0 , \2947_A[10]_b0 , w_7301 );
and ( w_7300 , w_7301 , \2989_B[13]_b0 );
or ( \4201_b1 , \4199_b1 , \4200_b1 );
not ( \4200_b1 , w_7302 );
and ( \4201_b0 , \4199_b0 , w_7303 );
and ( w_7302 , w_7303 , \4200_b0 );
or ( \4202_b1 , \4199_b1 , \4200_b1 );
xor ( \4202_b0 , \4199_b0 , w_7304 );
not ( w_7304 , w_7305 );
and ( w_7305 , \4200_b1 , \4200_b0 );
or ( \4203_b1 , \4104_b1 , \4161_b1 );
xor ( \4203_b0 , \4104_b0 , w_7306 );
not ( w_7306 , w_7307 );
and ( w_7307 , \4161_b1 , \4161_b0 );
or ( \4204_b1 , \2951_A[9]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7308 );
and ( \4204_b0 , \2951_A[9]_b0 , w_7309 );
and ( w_7308 , w_7309 , \2989_B[13]_b0 );
or ( \4205_b1 , \4203_b1 , \4204_b1 );
not ( \4204_b1 , w_7310 );
and ( \4205_b0 , \4203_b0 , w_7311 );
and ( w_7310 , w_7311 , \4204_b0 );
or ( \4206_b1 , \4203_b1 , \4204_b1 );
xor ( \4206_b0 , \4203_b0 , w_7312 );
not ( w_7312 , w_7313 );
and ( w_7313 , \4204_b1 , \4204_b0 );
or ( \4207_b1 , \4108_b1 , \4159_b1 );
xor ( \4207_b0 , \4108_b0 , w_7314 );
not ( w_7314 , w_7315 );
and ( w_7315 , \4159_b1 , \4159_b0 );
or ( \4208_b1 , \2955_A[8]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7316 );
and ( \4208_b0 , \2955_A[8]_b0 , w_7317 );
and ( w_7316 , w_7317 , \2989_B[13]_b0 );
or ( \4209_b1 , \4207_b1 , \4208_b1 );
not ( \4208_b1 , w_7318 );
and ( \4209_b0 , \4207_b0 , w_7319 );
and ( w_7318 , w_7319 , \4208_b0 );
or ( \4210_b1 , \4207_b1 , \4208_b1 );
xor ( \4210_b0 , \4207_b0 , w_7320 );
not ( w_7320 , w_7321 );
and ( w_7321 , \4208_b1 , \4208_b0 );
or ( \4211_b1 , \4112_b1 , \4157_b1 );
xor ( \4211_b0 , \4112_b0 , w_7322 );
not ( w_7322 , w_7323 );
and ( w_7323 , \4157_b1 , \4157_b0 );
or ( \4212_b1 , \2959_A[7]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7324 );
and ( \4212_b0 , \2959_A[7]_b0 , w_7325 );
and ( w_7324 , w_7325 , \2989_B[13]_b0 );
or ( \4213_b1 , \4211_b1 , \4212_b1 );
not ( \4212_b1 , w_7326 );
and ( \4213_b0 , \4211_b0 , w_7327 );
and ( w_7326 , w_7327 , \4212_b0 );
or ( \4214_b1 , \4211_b1 , \4212_b1 );
xor ( \4214_b0 , \4211_b0 , w_7328 );
not ( w_7328 , w_7329 );
and ( w_7329 , \4212_b1 , \4212_b0 );
or ( \4215_b1 , \4116_b1 , \4155_b1 );
xor ( \4215_b0 , \4116_b0 , w_7330 );
not ( w_7330 , w_7331 );
and ( w_7331 , \4155_b1 , \4155_b0 );
or ( \4216_b1 , \2963_A[6]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7332 );
and ( \4216_b0 , \2963_A[6]_b0 , w_7333 );
and ( w_7332 , w_7333 , \2989_B[13]_b0 );
or ( \4217_b1 , \4215_b1 , \4216_b1 );
not ( \4216_b1 , w_7334 );
and ( \4217_b0 , \4215_b0 , w_7335 );
and ( w_7334 , w_7335 , \4216_b0 );
or ( \4218_b1 , \4215_b1 , \4216_b1 );
xor ( \4218_b0 , \4215_b0 , w_7336 );
not ( w_7336 , w_7337 );
and ( w_7337 , \4216_b1 , \4216_b0 );
or ( \4219_b1 , \4120_b1 , \4153_b1 );
xor ( \4219_b0 , \4120_b0 , w_7338 );
not ( w_7338 , w_7339 );
and ( w_7339 , \4153_b1 , \4153_b0 );
or ( \4220_b1 , \2967_A[5]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7340 );
and ( \4220_b0 , \2967_A[5]_b0 , w_7341 );
and ( w_7340 , w_7341 , \2989_B[13]_b0 );
or ( \4221_b1 , \4219_b1 , \4220_b1 );
not ( \4220_b1 , w_7342 );
and ( \4221_b0 , \4219_b0 , w_7343 );
and ( w_7342 , w_7343 , \4220_b0 );
or ( \4222_b1 , \4219_b1 , \4220_b1 );
xor ( \4222_b0 , \4219_b0 , w_7344 );
not ( w_7344 , w_7345 );
and ( w_7345 , \4220_b1 , \4220_b0 );
or ( \4223_b1 , \4124_b1 , \4151_b1 );
xor ( \4223_b0 , \4124_b0 , w_7346 );
not ( w_7346 , w_7347 );
and ( w_7347 , \4151_b1 , \4151_b0 );
or ( \4224_b1 , \2971_A[4]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7348 );
and ( \4224_b0 , \2971_A[4]_b0 , w_7349 );
and ( w_7348 , w_7349 , \2989_B[13]_b0 );
or ( \4225_b1 , \4223_b1 , \4224_b1 );
not ( \4224_b1 , w_7350 );
and ( \4225_b0 , \4223_b0 , w_7351 );
and ( w_7350 , w_7351 , \4224_b0 );
or ( \4226_b1 , \4223_b1 , \4224_b1 );
xor ( \4226_b0 , \4223_b0 , w_7352 );
not ( w_7352 , w_7353 );
and ( w_7353 , \4224_b1 , \4224_b0 );
or ( \4227_b1 , \4128_b1 , \4149_b1 );
xor ( \4227_b0 , \4128_b0 , w_7354 );
not ( w_7354 , w_7355 );
and ( w_7355 , \4149_b1 , \4149_b0 );
or ( \4228_b1 , \2975_A[3]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7356 );
and ( \4228_b0 , \2975_A[3]_b0 , w_7357 );
and ( w_7356 , w_7357 , \2989_B[13]_b0 );
or ( \4229_b1 , \4227_b1 , \4228_b1 );
not ( \4228_b1 , w_7358 );
and ( \4229_b0 , \4227_b0 , w_7359 );
and ( w_7358 , w_7359 , \4228_b0 );
or ( \4230_b1 , \4227_b1 , \4228_b1 );
xor ( \4230_b0 , \4227_b0 , w_7360 );
not ( w_7360 , w_7361 );
and ( w_7361 , \4228_b1 , \4228_b0 );
or ( \4231_b1 , \4132_b1 , \4147_b1 );
xor ( \4231_b0 , \4132_b0 , w_7362 );
not ( w_7362 , w_7363 );
and ( w_7363 , \4147_b1 , \4147_b0 );
or ( \4232_b1 , \2979_A[2]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7364 );
and ( \4232_b0 , \2979_A[2]_b0 , w_7365 );
and ( w_7364 , w_7365 , \2989_B[13]_b0 );
or ( \4233_b1 , \4231_b1 , \4232_b1 );
not ( \4232_b1 , w_7366 );
and ( \4233_b0 , \4231_b0 , w_7367 );
and ( w_7366 , w_7367 , \4232_b0 );
or ( \4234_b1 , \4231_b1 , \4232_b1 );
xor ( \4234_b0 , \4231_b0 , w_7368 );
not ( w_7368 , w_7369 );
and ( w_7369 , \4232_b1 , \4232_b0 );
or ( \4235_b1 , \4136_b1 , \4145_b1 );
xor ( \4235_b0 , \4136_b0 , w_7370 );
not ( w_7370 , w_7371 );
and ( w_7371 , \4145_b1 , \4145_b0 );
or ( \4236_b1 , \2983_A[1]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7372 );
and ( \4236_b0 , \2983_A[1]_b0 , w_7373 );
and ( w_7372 , w_7373 , \2989_B[13]_b0 );
or ( \4237_b1 , \4235_b1 , \4236_b1 );
not ( \4236_b1 , w_7374 );
and ( \4237_b0 , \4235_b0 , w_7375 );
and ( w_7374 , w_7375 , \4236_b0 );
or ( \4238_b1 , \4235_b1 , \4236_b1 );
xor ( \4238_b0 , \4235_b0 , w_7376 );
not ( w_7376 , w_7377 );
and ( w_7377 , \4236_b1 , \4236_b0 );
or ( \4239_b1 , \4140_b1 , \4143_b1 );
xor ( \4239_b0 , \4140_b0 , w_7378 );
not ( w_7378 , w_7379 );
and ( w_7379 , \4143_b1 , \4143_b0 );
or ( \4240_b1 , \2986_A[0]_b1 , \2989_B[13]_b1 );
not ( \2989_B[13]_b1 , w_7380 );
and ( \4240_b0 , \2986_A[0]_b0 , w_7381 );
and ( w_7380 , w_7381 , \2989_B[13]_b0 );
or ( \4241_b1 , \4239_b1 , \4240_b1 );
not ( \4240_b1 , w_7382 );
and ( \4241_b0 , \4239_b0 , w_7383 );
and ( w_7382 , w_7383 , \4240_b0 );
or ( \4242_b1 , \4238_b1 , \4241_b1 );
not ( \4241_b1 , w_7384 );
and ( \4242_b0 , \4238_b0 , w_7385 );
and ( w_7384 , w_7385 , \4241_b0 );
or ( \4243_b1 , \4237_b1 , w_7386 );
or ( \4243_b0 , \4237_b0 , \4242_b0 );
not ( \4242_b0 , w_7387 );
and ( w_7387 , w_7386 , \4242_b1 );
or ( \4244_b1 , \4234_b1 , \4243_b1 );
not ( \4243_b1 , w_7388 );
and ( \4244_b0 , \4234_b0 , w_7389 );
and ( w_7388 , w_7389 , \4243_b0 );
or ( \4245_b1 , \4233_b1 , w_7390 );
or ( \4245_b0 , \4233_b0 , \4244_b0 );
not ( \4244_b0 , w_7391 );
and ( w_7391 , w_7390 , \4244_b1 );
or ( \4246_b1 , \4230_b1 , \4245_b1 );
not ( \4245_b1 , w_7392 );
and ( \4246_b0 , \4230_b0 , w_7393 );
and ( w_7392 , w_7393 , \4245_b0 );
or ( \4247_b1 , \4229_b1 , w_7394 );
or ( \4247_b0 , \4229_b0 , \4246_b0 );
not ( \4246_b0 , w_7395 );
and ( w_7395 , w_7394 , \4246_b1 );
or ( \4248_b1 , \4226_b1 , \4247_b1 );
not ( \4247_b1 , w_7396 );
and ( \4248_b0 , \4226_b0 , w_7397 );
and ( w_7396 , w_7397 , \4247_b0 );
or ( \4249_b1 , \4225_b1 , w_7398 );
or ( \4249_b0 , \4225_b0 , \4248_b0 );
not ( \4248_b0 , w_7399 );
and ( w_7399 , w_7398 , \4248_b1 );
or ( \4250_b1 , \4222_b1 , \4249_b1 );
not ( \4249_b1 , w_7400 );
and ( \4250_b0 , \4222_b0 , w_7401 );
and ( w_7400 , w_7401 , \4249_b0 );
or ( \4251_b1 , \4221_b1 , w_7402 );
or ( \4251_b0 , \4221_b0 , \4250_b0 );
not ( \4250_b0 , w_7403 );
and ( w_7403 , w_7402 , \4250_b1 );
or ( \4252_b1 , \4218_b1 , \4251_b1 );
not ( \4251_b1 , w_7404 );
and ( \4252_b0 , \4218_b0 , w_7405 );
and ( w_7404 , w_7405 , \4251_b0 );
or ( \4253_b1 , \4217_b1 , w_7406 );
or ( \4253_b0 , \4217_b0 , \4252_b0 );
not ( \4252_b0 , w_7407 );
and ( w_7407 , w_7406 , \4252_b1 );
or ( \4254_b1 , \4214_b1 , \4253_b1 );
not ( \4253_b1 , w_7408 );
and ( \4254_b0 , \4214_b0 , w_7409 );
and ( w_7408 , w_7409 , \4253_b0 );
or ( \4255_b1 , \4213_b1 , w_7410 );
or ( \4255_b0 , \4213_b0 , \4254_b0 );
not ( \4254_b0 , w_7411 );
and ( w_7411 , w_7410 , \4254_b1 );
or ( \4256_b1 , \4210_b1 , \4255_b1 );
not ( \4255_b1 , w_7412 );
and ( \4256_b0 , \4210_b0 , w_7413 );
and ( w_7412 , w_7413 , \4255_b0 );
or ( \4257_b1 , \4209_b1 , w_7414 );
or ( \4257_b0 , \4209_b0 , \4256_b0 );
not ( \4256_b0 , w_7415 );
and ( w_7415 , w_7414 , \4256_b1 );
or ( \4258_b1 , \4206_b1 , \4257_b1 );
not ( \4257_b1 , w_7416 );
and ( \4258_b0 , \4206_b0 , w_7417 );
and ( w_7416 , w_7417 , \4257_b0 );
or ( \4259_b1 , \4205_b1 , w_7418 );
or ( \4259_b0 , \4205_b0 , \4258_b0 );
not ( \4258_b0 , w_7419 );
and ( w_7419 , w_7418 , \4258_b1 );
or ( \4260_b1 , \4202_b1 , \4259_b1 );
not ( \4259_b1 , w_7420 );
and ( \4260_b0 , \4202_b0 , w_7421 );
and ( w_7420 , w_7421 , \4259_b0 );
or ( \4261_b1 , \4201_b1 , w_7422 );
or ( \4261_b0 , \4201_b0 , \4260_b0 );
not ( \4260_b0 , w_7423 );
and ( w_7423 , w_7422 , \4260_b1 );
or ( \4262_b1 , \4198_b1 , \4261_b1 );
not ( \4261_b1 , w_7424 );
and ( \4262_b0 , \4198_b0 , w_7425 );
and ( w_7424 , w_7425 , \4261_b0 );
or ( \4263_b1 , \4197_b1 , w_7426 );
or ( \4263_b0 , \4197_b0 , \4262_b0 );
not ( \4262_b0 , w_7427 );
and ( w_7427 , w_7426 , \4262_b1 );
or ( \4264_b1 , \4194_b1 , \4263_b1 );
not ( \4263_b1 , w_7428 );
and ( \4264_b0 , \4194_b0 , w_7429 );
and ( w_7428 , w_7429 , \4263_b0 );
or ( \4265_b1 , \4193_b1 , w_7430 );
or ( \4265_b0 , \4193_b0 , \4264_b0 );
not ( \4264_b0 , w_7431 );
and ( w_7431 , w_7430 , \4264_b1 );
or ( \4266_b1 , \4190_b1 , \4265_b1 );
not ( \4265_b1 , w_7432 );
and ( \4266_b0 , \4190_b0 , w_7433 );
and ( w_7432 , w_7433 , \4265_b0 );
or ( \4267_b1 , \4189_b1 , w_7434 );
or ( \4267_b0 , \4189_b0 , \4266_b0 );
not ( \4266_b0 , w_7435 );
and ( w_7435 , w_7434 , \4266_b1 );
or ( \4268_b1 , \4186_b1 , \4267_b1 );
not ( \4267_b1 , w_7436 );
and ( \4268_b0 , \4186_b0 , w_7437 );
and ( w_7436 , w_7437 , \4267_b0 );
or ( \4269_b1 , \4185_b1 , w_7438 );
or ( \4269_b0 , \4185_b0 , \4268_b0 );
not ( \4268_b0 , w_7439 );
and ( w_7439 , w_7438 , \4268_b1 );
or ( \4270_b1 , \4182_b1 , \4269_b1 );
not ( \4269_b1 , w_7440 );
and ( \4270_b0 , \4182_b0 , w_7441 );
and ( w_7440 , w_7441 , \4269_b0 );
or ( \4271_b1 , \4181_b1 , w_7442 );
or ( \4271_b0 , \4181_b0 , \4270_b0 );
not ( \4270_b0 , w_7443 );
and ( w_7443 , w_7442 , \4270_b1 );
or ( \4272_b1 , \4178_b1 , \4271_b1 );
not ( \4271_b1 , w_7444 );
and ( \4272_b0 , \4178_b0 , w_7445 );
and ( w_7444 , w_7445 , \4271_b0 );
or ( \4273_b1 , \4177_b1 , w_7446 );
or ( \4273_b0 , \4177_b0 , \4272_b0 );
not ( \4272_b0 , w_7447 );
and ( w_7447 , w_7446 , \4272_b1 );
or ( \4274_b1 , \2923_A[16]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7448 );
and ( \4274_b0 , \2923_A[16]_b0 , w_7449 );
and ( w_7448 , w_7449 , \2988_B[14]_b0 );
or ( \4275_b1 , \4273_b1 , \4274_b1 );
not ( \4274_b1 , w_7450 );
and ( \4275_b0 , \4273_b0 , w_7451 );
and ( w_7450 , w_7451 , \4274_b0 );
or ( \4276_b1 , \4273_b1 , \4274_b1 );
xor ( \4276_b0 , \4273_b0 , w_7452 );
not ( w_7452 , w_7453 );
and ( w_7453 , \4274_b1 , \4274_b0 );
or ( \4277_b1 , \4178_b1 , \4271_b1 );
xor ( \4277_b0 , \4178_b0 , w_7454 );
not ( w_7454 , w_7455 );
and ( w_7455 , \4271_b1 , \4271_b0 );
or ( \4278_b1 , \2927_A[15]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7456 );
and ( \4278_b0 , \2927_A[15]_b0 , w_7457 );
and ( w_7456 , w_7457 , \2988_B[14]_b0 );
or ( \4279_b1 , \4277_b1 , \4278_b1 );
not ( \4278_b1 , w_7458 );
and ( \4279_b0 , \4277_b0 , w_7459 );
and ( w_7458 , w_7459 , \4278_b0 );
or ( \4280_b1 , \4277_b1 , \4278_b1 );
xor ( \4280_b0 , \4277_b0 , w_7460 );
not ( w_7460 , w_7461 );
and ( w_7461 , \4278_b1 , \4278_b0 );
or ( \4281_b1 , \4182_b1 , \4269_b1 );
xor ( \4281_b0 , \4182_b0 , w_7462 );
not ( w_7462 , w_7463 );
and ( w_7463 , \4269_b1 , \4269_b0 );
or ( \4282_b1 , \2931_A[14]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7464 );
and ( \4282_b0 , \2931_A[14]_b0 , w_7465 );
and ( w_7464 , w_7465 , \2988_B[14]_b0 );
or ( \4283_b1 , \4281_b1 , \4282_b1 );
not ( \4282_b1 , w_7466 );
and ( \4283_b0 , \4281_b0 , w_7467 );
and ( w_7466 , w_7467 , \4282_b0 );
or ( \4284_b1 , \4281_b1 , \4282_b1 );
xor ( \4284_b0 , \4281_b0 , w_7468 );
not ( w_7468 , w_7469 );
and ( w_7469 , \4282_b1 , \4282_b0 );
or ( \4285_b1 , \4186_b1 , \4267_b1 );
xor ( \4285_b0 , \4186_b0 , w_7470 );
not ( w_7470 , w_7471 );
and ( w_7471 , \4267_b1 , \4267_b0 );
or ( \4286_b1 , \2935_A[13]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7472 );
and ( \4286_b0 , \2935_A[13]_b0 , w_7473 );
and ( w_7472 , w_7473 , \2988_B[14]_b0 );
or ( \4287_b1 , \4285_b1 , \4286_b1 );
not ( \4286_b1 , w_7474 );
and ( \4287_b0 , \4285_b0 , w_7475 );
and ( w_7474 , w_7475 , \4286_b0 );
or ( \4288_b1 , \4285_b1 , \4286_b1 );
xor ( \4288_b0 , \4285_b0 , w_7476 );
not ( w_7476 , w_7477 );
and ( w_7477 , \4286_b1 , \4286_b0 );
or ( \4289_b1 , \4190_b1 , \4265_b1 );
xor ( \4289_b0 , \4190_b0 , w_7478 );
not ( w_7478 , w_7479 );
and ( w_7479 , \4265_b1 , \4265_b0 );
or ( \4290_b1 , \2939_A[12]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7480 );
and ( \4290_b0 , \2939_A[12]_b0 , w_7481 );
and ( w_7480 , w_7481 , \2988_B[14]_b0 );
or ( \4291_b1 , \4289_b1 , \4290_b1 );
not ( \4290_b1 , w_7482 );
and ( \4291_b0 , \4289_b0 , w_7483 );
and ( w_7482 , w_7483 , \4290_b0 );
or ( \4292_b1 , \4289_b1 , \4290_b1 );
xor ( \4292_b0 , \4289_b0 , w_7484 );
not ( w_7484 , w_7485 );
and ( w_7485 , \4290_b1 , \4290_b0 );
or ( \4293_b1 , \4194_b1 , \4263_b1 );
xor ( \4293_b0 , \4194_b0 , w_7486 );
not ( w_7486 , w_7487 );
and ( w_7487 , \4263_b1 , \4263_b0 );
or ( \4294_b1 , \2943_A[11]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7488 );
and ( \4294_b0 , \2943_A[11]_b0 , w_7489 );
and ( w_7488 , w_7489 , \2988_B[14]_b0 );
or ( \4295_b1 , \4293_b1 , \4294_b1 );
not ( \4294_b1 , w_7490 );
and ( \4295_b0 , \4293_b0 , w_7491 );
and ( w_7490 , w_7491 , \4294_b0 );
or ( \4296_b1 , \4293_b1 , \4294_b1 );
xor ( \4296_b0 , \4293_b0 , w_7492 );
not ( w_7492 , w_7493 );
and ( w_7493 , \4294_b1 , \4294_b0 );
or ( \4297_b1 , \4198_b1 , \4261_b1 );
xor ( \4297_b0 , \4198_b0 , w_7494 );
not ( w_7494 , w_7495 );
and ( w_7495 , \4261_b1 , \4261_b0 );
or ( \4298_b1 , \2947_A[10]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7496 );
and ( \4298_b0 , \2947_A[10]_b0 , w_7497 );
and ( w_7496 , w_7497 , \2988_B[14]_b0 );
or ( \4299_b1 , \4297_b1 , \4298_b1 );
not ( \4298_b1 , w_7498 );
and ( \4299_b0 , \4297_b0 , w_7499 );
and ( w_7498 , w_7499 , \4298_b0 );
or ( \4300_b1 , \4297_b1 , \4298_b1 );
xor ( \4300_b0 , \4297_b0 , w_7500 );
not ( w_7500 , w_7501 );
and ( w_7501 , \4298_b1 , \4298_b0 );
or ( \4301_b1 , \4202_b1 , \4259_b1 );
xor ( \4301_b0 , \4202_b0 , w_7502 );
not ( w_7502 , w_7503 );
and ( w_7503 , \4259_b1 , \4259_b0 );
or ( \4302_b1 , \2951_A[9]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7504 );
and ( \4302_b0 , \2951_A[9]_b0 , w_7505 );
and ( w_7504 , w_7505 , \2988_B[14]_b0 );
or ( \4303_b1 , \4301_b1 , \4302_b1 );
not ( \4302_b1 , w_7506 );
and ( \4303_b0 , \4301_b0 , w_7507 );
and ( w_7506 , w_7507 , \4302_b0 );
or ( \4304_b1 , \4301_b1 , \4302_b1 );
xor ( \4304_b0 , \4301_b0 , w_7508 );
not ( w_7508 , w_7509 );
and ( w_7509 , \4302_b1 , \4302_b0 );
or ( \4305_b1 , \4206_b1 , \4257_b1 );
xor ( \4305_b0 , \4206_b0 , w_7510 );
not ( w_7510 , w_7511 );
and ( w_7511 , \4257_b1 , \4257_b0 );
or ( \4306_b1 , \2955_A[8]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7512 );
and ( \4306_b0 , \2955_A[8]_b0 , w_7513 );
and ( w_7512 , w_7513 , \2988_B[14]_b0 );
or ( \4307_b1 , \4305_b1 , \4306_b1 );
not ( \4306_b1 , w_7514 );
and ( \4307_b0 , \4305_b0 , w_7515 );
and ( w_7514 , w_7515 , \4306_b0 );
or ( \4308_b1 , \4305_b1 , \4306_b1 );
xor ( \4308_b0 , \4305_b0 , w_7516 );
not ( w_7516 , w_7517 );
and ( w_7517 , \4306_b1 , \4306_b0 );
or ( \4309_b1 , \4210_b1 , \4255_b1 );
xor ( \4309_b0 , \4210_b0 , w_7518 );
not ( w_7518 , w_7519 );
and ( w_7519 , \4255_b1 , \4255_b0 );
or ( \4310_b1 , \2959_A[7]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7520 );
and ( \4310_b0 , \2959_A[7]_b0 , w_7521 );
and ( w_7520 , w_7521 , \2988_B[14]_b0 );
or ( \4311_b1 , \4309_b1 , \4310_b1 );
not ( \4310_b1 , w_7522 );
and ( \4311_b0 , \4309_b0 , w_7523 );
and ( w_7522 , w_7523 , \4310_b0 );
or ( \4312_b1 , \4309_b1 , \4310_b1 );
xor ( \4312_b0 , \4309_b0 , w_7524 );
not ( w_7524 , w_7525 );
and ( w_7525 , \4310_b1 , \4310_b0 );
or ( \4313_b1 , \4214_b1 , \4253_b1 );
xor ( \4313_b0 , \4214_b0 , w_7526 );
not ( w_7526 , w_7527 );
and ( w_7527 , \4253_b1 , \4253_b0 );
or ( \4314_b1 , \2963_A[6]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7528 );
and ( \4314_b0 , \2963_A[6]_b0 , w_7529 );
and ( w_7528 , w_7529 , \2988_B[14]_b0 );
or ( \4315_b1 , \4313_b1 , \4314_b1 );
not ( \4314_b1 , w_7530 );
and ( \4315_b0 , \4313_b0 , w_7531 );
and ( w_7530 , w_7531 , \4314_b0 );
or ( \4316_b1 , \4313_b1 , \4314_b1 );
xor ( \4316_b0 , \4313_b0 , w_7532 );
not ( w_7532 , w_7533 );
and ( w_7533 , \4314_b1 , \4314_b0 );
or ( \4317_b1 , \4218_b1 , \4251_b1 );
xor ( \4317_b0 , \4218_b0 , w_7534 );
not ( w_7534 , w_7535 );
and ( w_7535 , \4251_b1 , \4251_b0 );
or ( \4318_b1 , \2967_A[5]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7536 );
and ( \4318_b0 , \2967_A[5]_b0 , w_7537 );
and ( w_7536 , w_7537 , \2988_B[14]_b0 );
or ( \4319_b1 , \4317_b1 , \4318_b1 );
not ( \4318_b1 , w_7538 );
and ( \4319_b0 , \4317_b0 , w_7539 );
and ( w_7538 , w_7539 , \4318_b0 );
or ( \4320_b1 , \4317_b1 , \4318_b1 );
xor ( \4320_b0 , \4317_b0 , w_7540 );
not ( w_7540 , w_7541 );
and ( w_7541 , \4318_b1 , \4318_b0 );
or ( \4321_b1 , \4222_b1 , \4249_b1 );
xor ( \4321_b0 , \4222_b0 , w_7542 );
not ( w_7542 , w_7543 );
and ( w_7543 , \4249_b1 , \4249_b0 );
or ( \4322_b1 , \2971_A[4]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7544 );
and ( \4322_b0 , \2971_A[4]_b0 , w_7545 );
and ( w_7544 , w_7545 , \2988_B[14]_b0 );
or ( \4323_b1 , \4321_b1 , \4322_b1 );
not ( \4322_b1 , w_7546 );
and ( \4323_b0 , \4321_b0 , w_7547 );
and ( w_7546 , w_7547 , \4322_b0 );
or ( \4324_b1 , \4321_b1 , \4322_b1 );
xor ( \4324_b0 , \4321_b0 , w_7548 );
not ( w_7548 , w_7549 );
and ( w_7549 , \4322_b1 , \4322_b0 );
or ( \4325_b1 , \4226_b1 , \4247_b1 );
xor ( \4325_b0 , \4226_b0 , w_7550 );
not ( w_7550 , w_7551 );
and ( w_7551 , \4247_b1 , \4247_b0 );
or ( \4326_b1 , \2975_A[3]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7552 );
and ( \4326_b0 , \2975_A[3]_b0 , w_7553 );
and ( w_7552 , w_7553 , \2988_B[14]_b0 );
or ( \4327_b1 , \4325_b1 , \4326_b1 );
not ( \4326_b1 , w_7554 );
and ( \4327_b0 , \4325_b0 , w_7555 );
and ( w_7554 , w_7555 , \4326_b0 );
or ( \4328_b1 , \4325_b1 , \4326_b1 );
xor ( \4328_b0 , \4325_b0 , w_7556 );
not ( w_7556 , w_7557 );
and ( w_7557 , \4326_b1 , \4326_b0 );
or ( \4329_b1 , \4230_b1 , \4245_b1 );
xor ( \4329_b0 , \4230_b0 , w_7558 );
not ( w_7558 , w_7559 );
and ( w_7559 , \4245_b1 , \4245_b0 );
or ( \4330_b1 , \2979_A[2]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7560 );
and ( \4330_b0 , \2979_A[2]_b0 , w_7561 );
and ( w_7560 , w_7561 , \2988_B[14]_b0 );
or ( \4331_b1 , \4329_b1 , \4330_b1 );
not ( \4330_b1 , w_7562 );
and ( \4331_b0 , \4329_b0 , w_7563 );
and ( w_7562 , w_7563 , \4330_b0 );
or ( \4332_b1 , \4329_b1 , \4330_b1 );
xor ( \4332_b0 , \4329_b0 , w_7564 );
not ( w_7564 , w_7565 );
and ( w_7565 , \4330_b1 , \4330_b0 );
or ( \4333_b1 , \4234_b1 , \4243_b1 );
xor ( \4333_b0 , \4234_b0 , w_7566 );
not ( w_7566 , w_7567 );
and ( w_7567 , \4243_b1 , \4243_b0 );
or ( \4334_b1 , \2983_A[1]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7568 );
and ( \4334_b0 , \2983_A[1]_b0 , w_7569 );
and ( w_7568 , w_7569 , \2988_B[14]_b0 );
or ( \4335_b1 , \4333_b1 , \4334_b1 );
not ( \4334_b1 , w_7570 );
and ( \4335_b0 , \4333_b0 , w_7571 );
and ( w_7570 , w_7571 , \4334_b0 );
or ( \4336_b1 , \4333_b1 , \4334_b1 );
xor ( \4336_b0 , \4333_b0 , w_7572 );
not ( w_7572 , w_7573 );
and ( w_7573 , \4334_b1 , \4334_b0 );
or ( \4337_b1 , \4238_b1 , \4241_b1 );
xor ( \4337_b0 , \4238_b0 , w_7574 );
not ( w_7574 , w_7575 );
and ( w_7575 , \4241_b1 , \4241_b0 );
or ( \4338_b1 , \2986_A[0]_b1 , \2988_B[14]_b1 );
not ( \2988_B[14]_b1 , w_7576 );
and ( \4338_b0 , \2986_A[0]_b0 , w_7577 );
and ( w_7576 , w_7577 , \2988_B[14]_b0 );
or ( \4339_b1 , \4337_b1 , \4338_b1 );
not ( \4338_b1 , w_7578 );
and ( \4339_b0 , \4337_b0 , w_7579 );
and ( w_7578 , w_7579 , \4338_b0 );
or ( \4340_b1 , \4336_b1 , \4339_b1 );
not ( \4339_b1 , w_7580 );
and ( \4340_b0 , \4336_b0 , w_7581 );
and ( w_7580 , w_7581 , \4339_b0 );
or ( \4341_b1 , \4335_b1 , w_7582 );
or ( \4341_b0 , \4335_b0 , \4340_b0 );
not ( \4340_b0 , w_7583 );
and ( w_7583 , w_7582 , \4340_b1 );
or ( \4342_b1 , \4332_b1 , \4341_b1 );
not ( \4341_b1 , w_7584 );
and ( \4342_b0 , \4332_b0 , w_7585 );
and ( w_7584 , w_7585 , \4341_b0 );
or ( \4343_b1 , \4331_b1 , w_7586 );
or ( \4343_b0 , \4331_b0 , \4342_b0 );
not ( \4342_b0 , w_7587 );
and ( w_7587 , w_7586 , \4342_b1 );
or ( \4344_b1 , \4328_b1 , \4343_b1 );
not ( \4343_b1 , w_7588 );
and ( \4344_b0 , \4328_b0 , w_7589 );
and ( w_7588 , w_7589 , \4343_b0 );
or ( \4345_b1 , \4327_b1 , w_7590 );
or ( \4345_b0 , \4327_b0 , \4344_b0 );
not ( \4344_b0 , w_7591 );
and ( w_7591 , w_7590 , \4344_b1 );
or ( \4346_b1 , \4324_b1 , \4345_b1 );
not ( \4345_b1 , w_7592 );
and ( \4346_b0 , \4324_b0 , w_7593 );
and ( w_7592 , w_7593 , \4345_b0 );
or ( \4347_b1 , \4323_b1 , w_7594 );
or ( \4347_b0 , \4323_b0 , \4346_b0 );
not ( \4346_b0 , w_7595 );
and ( w_7595 , w_7594 , \4346_b1 );
or ( \4348_b1 , \4320_b1 , \4347_b1 );
not ( \4347_b1 , w_7596 );
and ( \4348_b0 , \4320_b0 , w_7597 );
and ( w_7596 , w_7597 , \4347_b0 );
or ( \4349_b1 , \4319_b1 , w_7598 );
or ( \4349_b0 , \4319_b0 , \4348_b0 );
not ( \4348_b0 , w_7599 );
and ( w_7599 , w_7598 , \4348_b1 );
or ( \4350_b1 , \4316_b1 , \4349_b1 );
not ( \4349_b1 , w_7600 );
and ( \4350_b0 , \4316_b0 , w_7601 );
and ( w_7600 , w_7601 , \4349_b0 );
or ( \4351_b1 , \4315_b1 , w_7602 );
or ( \4351_b0 , \4315_b0 , \4350_b0 );
not ( \4350_b0 , w_7603 );
and ( w_7603 , w_7602 , \4350_b1 );
or ( \4352_b1 , \4312_b1 , \4351_b1 );
not ( \4351_b1 , w_7604 );
and ( \4352_b0 , \4312_b0 , w_7605 );
and ( w_7604 , w_7605 , \4351_b0 );
or ( \4353_b1 , \4311_b1 , w_7606 );
or ( \4353_b0 , \4311_b0 , \4352_b0 );
not ( \4352_b0 , w_7607 );
and ( w_7607 , w_7606 , \4352_b1 );
or ( \4354_b1 , \4308_b1 , \4353_b1 );
not ( \4353_b1 , w_7608 );
and ( \4354_b0 , \4308_b0 , w_7609 );
and ( w_7608 , w_7609 , \4353_b0 );
or ( \4355_b1 , \4307_b1 , w_7610 );
or ( \4355_b0 , \4307_b0 , \4354_b0 );
not ( \4354_b0 , w_7611 );
and ( w_7611 , w_7610 , \4354_b1 );
or ( \4356_b1 , \4304_b1 , \4355_b1 );
not ( \4355_b1 , w_7612 );
and ( \4356_b0 , \4304_b0 , w_7613 );
and ( w_7612 , w_7613 , \4355_b0 );
or ( \4357_b1 , \4303_b1 , w_7614 );
or ( \4357_b0 , \4303_b0 , \4356_b0 );
not ( \4356_b0 , w_7615 );
and ( w_7615 , w_7614 , \4356_b1 );
or ( \4358_b1 , \4300_b1 , \4357_b1 );
not ( \4357_b1 , w_7616 );
and ( \4358_b0 , \4300_b0 , w_7617 );
and ( w_7616 , w_7617 , \4357_b0 );
or ( \4359_b1 , \4299_b1 , w_7618 );
or ( \4359_b0 , \4299_b0 , \4358_b0 );
not ( \4358_b0 , w_7619 );
and ( w_7619 , w_7618 , \4358_b1 );
or ( \4360_b1 , \4296_b1 , \4359_b1 );
not ( \4359_b1 , w_7620 );
and ( \4360_b0 , \4296_b0 , w_7621 );
and ( w_7620 , w_7621 , \4359_b0 );
or ( \4361_b1 , \4295_b1 , w_7622 );
or ( \4361_b0 , \4295_b0 , \4360_b0 );
not ( \4360_b0 , w_7623 );
and ( w_7623 , w_7622 , \4360_b1 );
or ( \4362_b1 , \4292_b1 , \4361_b1 );
not ( \4361_b1 , w_7624 );
and ( \4362_b0 , \4292_b0 , w_7625 );
and ( w_7624 , w_7625 , \4361_b0 );
or ( \4363_b1 , \4291_b1 , w_7626 );
or ( \4363_b0 , \4291_b0 , \4362_b0 );
not ( \4362_b0 , w_7627 );
and ( w_7627 , w_7626 , \4362_b1 );
or ( \4364_b1 , \4288_b1 , \4363_b1 );
not ( \4363_b1 , w_7628 );
and ( \4364_b0 , \4288_b0 , w_7629 );
and ( w_7628 , w_7629 , \4363_b0 );
or ( \4365_b1 , \4287_b1 , w_7630 );
or ( \4365_b0 , \4287_b0 , \4364_b0 );
not ( \4364_b0 , w_7631 );
and ( w_7631 , w_7630 , \4364_b1 );
or ( \4366_b1 , \4284_b1 , \4365_b1 );
not ( \4365_b1 , w_7632 );
and ( \4366_b0 , \4284_b0 , w_7633 );
and ( w_7632 , w_7633 , \4365_b0 );
or ( \4367_b1 , \4283_b1 , w_7634 );
or ( \4367_b0 , \4283_b0 , \4366_b0 );
not ( \4366_b0 , w_7635 );
and ( w_7635 , w_7634 , \4366_b1 );
or ( \4368_b1 , \4280_b1 , \4367_b1 );
not ( \4367_b1 , w_7636 );
and ( \4368_b0 , \4280_b0 , w_7637 );
and ( w_7636 , w_7637 , \4367_b0 );
or ( \4369_b1 , \4279_b1 , w_7638 );
or ( \4369_b0 , \4279_b0 , \4368_b0 );
not ( \4368_b0 , w_7639 );
and ( w_7639 , w_7638 , \4368_b1 );
or ( \4370_b1 , \4276_b1 , \4369_b1 );
not ( \4369_b1 , w_7640 );
and ( \4370_b0 , \4276_b0 , w_7641 );
and ( w_7640 , w_7641 , \4369_b0 );
or ( \4371_b1 , \4275_b1 , w_7642 );
or ( \4371_b0 , \4275_b0 , \4370_b0 );
not ( \4370_b0 , w_7643 );
and ( w_7643 , w_7642 , \4370_b1 );
or ( \4372_b1 , \2923_A[16]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7644 );
and ( \4372_b0 , \2923_A[16]_b0 , w_7645 );
and ( w_7644 , w_7645 , \2987_B[15]_b0 );
or ( \4373_b1 , \4371_b1 , \4372_b1 );
xor ( \4373_b0 , \4371_b0 , w_7646 );
not ( w_7646 , w_7647 );
and ( w_7647 , \4372_b1 , \4372_b0 );
or ( \4374_b1 , \4276_b1 , \4369_b1 );
xor ( \4374_b0 , \4276_b0 , w_7648 );
not ( w_7648 , w_7649 );
and ( w_7649 , \4369_b1 , \4369_b0 );
or ( \4375_b1 , \2927_A[15]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7650 );
and ( \4375_b0 , \2927_A[15]_b0 , w_7651 );
and ( w_7650 , w_7651 , \2987_B[15]_b0 );
or ( \4376_b1 , \4374_b1 , \4375_b1 );
not ( \4375_b1 , w_7652 );
and ( \4376_b0 , \4374_b0 , w_7653 );
and ( w_7652 , w_7653 , \4375_b0 );
or ( \4377_b1 , \4374_b1 , \4375_b1 );
xor ( \4377_b0 , \4374_b0 , w_7654 );
not ( w_7654 , w_7655 );
and ( w_7655 , \4375_b1 , \4375_b0 );
or ( \4378_b1 , \4280_b1 , \4367_b1 );
xor ( \4378_b0 , \4280_b0 , w_7656 );
not ( w_7656 , w_7657 );
and ( w_7657 , \4367_b1 , \4367_b0 );
or ( \4379_b1 , \2931_A[14]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7658 );
and ( \4379_b0 , \2931_A[14]_b0 , w_7659 );
and ( w_7658 , w_7659 , \2987_B[15]_b0 );
or ( \4380_b1 , \4378_b1 , \4379_b1 );
not ( \4379_b1 , w_7660 );
and ( \4380_b0 , \4378_b0 , w_7661 );
and ( w_7660 , w_7661 , \4379_b0 );
or ( \4381_b1 , \4378_b1 , \4379_b1 );
xor ( \4381_b0 , \4378_b0 , w_7662 );
not ( w_7662 , w_7663 );
and ( w_7663 , \4379_b1 , \4379_b0 );
or ( \4382_b1 , \4284_b1 , \4365_b1 );
xor ( \4382_b0 , \4284_b0 , w_7664 );
not ( w_7664 , w_7665 );
and ( w_7665 , \4365_b1 , \4365_b0 );
or ( \4383_b1 , \2935_A[13]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7666 );
and ( \4383_b0 , \2935_A[13]_b0 , w_7667 );
and ( w_7666 , w_7667 , \2987_B[15]_b0 );
or ( \4384_b1 , \4382_b1 , \4383_b1 );
not ( \4383_b1 , w_7668 );
and ( \4384_b0 , \4382_b0 , w_7669 );
and ( w_7668 , w_7669 , \4383_b0 );
or ( \4385_b1 , \4382_b1 , \4383_b1 );
xor ( \4385_b0 , \4382_b0 , w_7670 );
not ( w_7670 , w_7671 );
and ( w_7671 , \4383_b1 , \4383_b0 );
or ( \4386_b1 , \4288_b1 , \4363_b1 );
xor ( \4386_b0 , \4288_b0 , w_7672 );
not ( w_7672 , w_7673 );
and ( w_7673 , \4363_b1 , \4363_b0 );
or ( \4387_b1 , \2939_A[12]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7674 );
and ( \4387_b0 , \2939_A[12]_b0 , w_7675 );
and ( w_7674 , w_7675 , \2987_B[15]_b0 );
or ( \4388_b1 , \4386_b1 , \4387_b1 );
not ( \4387_b1 , w_7676 );
and ( \4388_b0 , \4386_b0 , w_7677 );
and ( w_7676 , w_7677 , \4387_b0 );
or ( \4389_b1 , \4386_b1 , \4387_b1 );
xor ( \4389_b0 , \4386_b0 , w_7678 );
not ( w_7678 , w_7679 );
and ( w_7679 , \4387_b1 , \4387_b0 );
or ( \4390_b1 , \4292_b1 , \4361_b1 );
xor ( \4390_b0 , \4292_b0 , w_7680 );
not ( w_7680 , w_7681 );
and ( w_7681 , \4361_b1 , \4361_b0 );
or ( \4391_b1 , \2943_A[11]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7682 );
and ( \4391_b0 , \2943_A[11]_b0 , w_7683 );
and ( w_7682 , w_7683 , \2987_B[15]_b0 );
or ( \4392_b1 , \4390_b1 , \4391_b1 );
not ( \4391_b1 , w_7684 );
and ( \4392_b0 , \4390_b0 , w_7685 );
and ( w_7684 , w_7685 , \4391_b0 );
or ( \4393_b1 , \4390_b1 , \4391_b1 );
xor ( \4393_b0 , \4390_b0 , w_7686 );
not ( w_7686 , w_7687 );
and ( w_7687 , \4391_b1 , \4391_b0 );
or ( \4394_b1 , \4296_b1 , \4359_b1 );
xor ( \4394_b0 , \4296_b0 , w_7688 );
not ( w_7688 , w_7689 );
and ( w_7689 , \4359_b1 , \4359_b0 );
or ( \4395_b1 , \2947_A[10]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7690 );
and ( \4395_b0 , \2947_A[10]_b0 , w_7691 );
and ( w_7690 , w_7691 , \2987_B[15]_b0 );
or ( \4396_b1 , \4394_b1 , \4395_b1 );
not ( \4395_b1 , w_7692 );
and ( \4396_b0 , \4394_b0 , w_7693 );
and ( w_7692 , w_7693 , \4395_b0 );
or ( \4397_b1 , \4394_b1 , \4395_b1 );
xor ( \4397_b0 , \4394_b0 , w_7694 );
not ( w_7694 , w_7695 );
and ( w_7695 , \4395_b1 , \4395_b0 );
or ( \4398_b1 , \4300_b1 , \4357_b1 );
xor ( \4398_b0 , \4300_b0 , w_7696 );
not ( w_7696 , w_7697 );
and ( w_7697 , \4357_b1 , \4357_b0 );
or ( \4399_b1 , \2951_A[9]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7698 );
and ( \4399_b0 , \2951_A[9]_b0 , w_7699 );
and ( w_7698 , w_7699 , \2987_B[15]_b0 );
or ( \4400_b1 , \4398_b1 , \4399_b1 );
not ( \4399_b1 , w_7700 );
and ( \4400_b0 , \4398_b0 , w_7701 );
and ( w_7700 , w_7701 , \4399_b0 );
or ( \4401_b1 , \4398_b1 , \4399_b1 );
xor ( \4401_b0 , \4398_b0 , w_7702 );
not ( w_7702 , w_7703 );
and ( w_7703 , \4399_b1 , \4399_b0 );
or ( \4402_b1 , \4304_b1 , \4355_b1 );
xor ( \4402_b0 , \4304_b0 , w_7704 );
not ( w_7704 , w_7705 );
and ( w_7705 , \4355_b1 , \4355_b0 );
or ( \4403_b1 , \2955_A[8]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7706 );
and ( \4403_b0 , \2955_A[8]_b0 , w_7707 );
and ( w_7706 , w_7707 , \2987_B[15]_b0 );
or ( \4404_b1 , \4402_b1 , \4403_b1 );
not ( \4403_b1 , w_7708 );
and ( \4404_b0 , \4402_b0 , w_7709 );
and ( w_7708 , w_7709 , \4403_b0 );
or ( \4405_b1 , \4402_b1 , \4403_b1 );
xor ( \4405_b0 , \4402_b0 , w_7710 );
not ( w_7710 , w_7711 );
and ( w_7711 , \4403_b1 , \4403_b0 );
or ( \4406_b1 , \4308_b1 , \4353_b1 );
xor ( \4406_b0 , \4308_b0 , w_7712 );
not ( w_7712 , w_7713 );
and ( w_7713 , \4353_b1 , \4353_b0 );
or ( \4407_b1 , \2959_A[7]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7714 );
and ( \4407_b0 , \2959_A[7]_b0 , w_7715 );
and ( w_7714 , w_7715 , \2987_B[15]_b0 );
or ( \4408_b1 , \4406_b1 , \4407_b1 );
not ( \4407_b1 , w_7716 );
and ( \4408_b0 , \4406_b0 , w_7717 );
and ( w_7716 , w_7717 , \4407_b0 );
or ( \4409_b1 , \4406_b1 , \4407_b1 );
xor ( \4409_b0 , \4406_b0 , w_7718 );
not ( w_7718 , w_7719 );
and ( w_7719 , \4407_b1 , \4407_b0 );
or ( \4410_b1 , \4312_b1 , \4351_b1 );
xor ( \4410_b0 , \4312_b0 , w_7720 );
not ( w_7720 , w_7721 );
and ( w_7721 , \4351_b1 , \4351_b0 );
or ( \4411_b1 , \2963_A[6]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7722 );
and ( \4411_b0 , \2963_A[6]_b0 , w_7723 );
and ( w_7722 , w_7723 , \2987_B[15]_b0 );
or ( \4412_b1 , \4410_b1 , \4411_b1 );
not ( \4411_b1 , w_7724 );
and ( \4412_b0 , \4410_b0 , w_7725 );
and ( w_7724 , w_7725 , \4411_b0 );
or ( \4413_b1 , \4410_b1 , \4411_b1 );
xor ( \4413_b0 , \4410_b0 , w_7726 );
not ( w_7726 , w_7727 );
and ( w_7727 , \4411_b1 , \4411_b0 );
or ( \4414_b1 , \4316_b1 , \4349_b1 );
xor ( \4414_b0 , \4316_b0 , w_7728 );
not ( w_7728 , w_7729 );
and ( w_7729 , \4349_b1 , \4349_b0 );
or ( \4415_b1 , \2967_A[5]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7730 );
and ( \4415_b0 , \2967_A[5]_b0 , w_7731 );
and ( w_7730 , w_7731 , \2987_B[15]_b0 );
or ( \4416_b1 , \4414_b1 , \4415_b1 );
not ( \4415_b1 , w_7732 );
and ( \4416_b0 , \4414_b0 , w_7733 );
and ( w_7732 , w_7733 , \4415_b0 );
or ( \4417_b1 , \4414_b1 , \4415_b1 );
xor ( \4417_b0 , \4414_b0 , w_7734 );
not ( w_7734 , w_7735 );
and ( w_7735 , \4415_b1 , \4415_b0 );
or ( \4418_b1 , \4320_b1 , \4347_b1 );
xor ( \4418_b0 , \4320_b0 , w_7736 );
not ( w_7736 , w_7737 );
and ( w_7737 , \4347_b1 , \4347_b0 );
or ( \4419_b1 , \2971_A[4]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7738 );
and ( \4419_b0 , \2971_A[4]_b0 , w_7739 );
and ( w_7738 , w_7739 , \2987_B[15]_b0 );
or ( \4420_b1 , \4418_b1 , \4419_b1 );
not ( \4419_b1 , w_7740 );
and ( \4420_b0 , \4418_b0 , w_7741 );
and ( w_7740 , w_7741 , \4419_b0 );
or ( \4421_b1 , \4418_b1 , \4419_b1 );
xor ( \4421_b0 , \4418_b0 , w_7742 );
not ( w_7742 , w_7743 );
and ( w_7743 , \4419_b1 , \4419_b0 );
or ( \4422_b1 , \4324_b1 , \4345_b1 );
xor ( \4422_b0 , \4324_b0 , w_7744 );
not ( w_7744 , w_7745 );
and ( w_7745 , \4345_b1 , \4345_b0 );
or ( \4423_b1 , \2975_A[3]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7746 );
and ( \4423_b0 , \2975_A[3]_b0 , w_7747 );
and ( w_7746 , w_7747 , \2987_B[15]_b0 );
or ( \4424_b1 , \4422_b1 , \4423_b1 );
not ( \4423_b1 , w_7748 );
and ( \4424_b0 , \4422_b0 , w_7749 );
and ( w_7748 , w_7749 , \4423_b0 );
or ( \4425_b1 , \4422_b1 , \4423_b1 );
xor ( \4425_b0 , \4422_b0 , w_7750 );
not ( w_7750 , w_7751 );
and ( w_7751 , \4423_b1 , \4423_b0 );
or ( \4426_b1 , \4328_b1 , \4343_b1 );
xor ( \4426_b0 , \4328_b0 , w_7752 );
not ( w_7752 , w_7753 );
and ( w_7753 , \4343_b1 , \4343_b0 );
or ( \4427_b1 , \2979_A[2]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7754 );
and ( \4427_b0 , \2979_A[2]_b0 , w_7755 );
and ( w_7754 , w_7755 , \2987_B[15]_b0 );
or ( \4428_b1 , \4426_b1 , \4427_b1 );
not ( \4427_b1 , w_7756 );
and ( \4428_b0 , \4426_b0 , w_7757 );
and ( w_7756 , w_7757 , \4427_b0 );
or ( \4429_b1 , \4426_b1 , \4427_b1 );
xor ( \4429_b0 , \4426_b0 , w_7758 );
not ( w_7758 , w_7759 );
and ( w_7759 , \4427_b1 , \4427_b0 );
or ( \4430_b1 , \4332_b1 , \4341_b1 );
xor ( \4430_b0 , \4332_b0 , w_7760 );
not ( w_7760 , w_7761 );
and ( w_7761 , \4341_b1 , \4341_b0 );
or ( \4431_b1 , \2983_A[1]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7762 );
and ( \4431_b0 , \2983_A[1]_b0 , w_7763 );
and ( w_7762 , w_7763 , \2987_B[15]_b0 );
or ( \4432_b1 , \4430_b1 , \4431_b1 );
not ( \4431_b1 , w_7764 );
and ( \4432_b0 , \4430_b0 , w_7765 );
and ( w_7764 , w_7765 , \4431_b0 );
or ( \4433_b1 , \4430_b1 , \4431_b1 );
xor ( \4433_b0 , \4430_b0 , w_7766 );
not ( w_7766 , w_7767 );
and ( w_7767 , \4431_b1 , \4431_b0 );
or ( \4434_b1 , \4336_b1 , \4339_b1 );
xor ( \4434_b0 , \4336_b0 , w_7768 );
not ( w_7768 , w_7769 );
and ( w_7769 , \4339_b1 , \4339_b0 );
or ( \4435_b1 , \2986_A[0]_b1 , \2987_B[15]_b1 );
not ( \2987_B[15]_b1 , w_7770 );
and ( \4435_b0 , \2986_A[0]_b0 , w_7771 );
and ( w_7770 , w_7771 , \2987_B[15]_b0 );
or ( \4436_b1 , \4434_b1 , \4435_b1 );
not ( \4435_b1 , w_7772 );
and ( \4436_b0 , \4434_b0 , w_7773 );
and ( w_7772 , w_7773 , \4435_b0 );
or ( \4437_b1 , \4433_b1 , \4436_b1 );
not ( \4436_b1 , w_7774 );
and ( \4437_b0 , \4433_b0 , w_7775 );
and ( w_7774 , w_7775 , \4436_b0 );
or ( \4438_b1 , \4432_b1 , w_7776 );
or ( \4438_b0 , \4432_b0 , \4437_b0 );
not ( \4437_b0 , w_7777 );
and ( w_7777 , w_7776 , \4437_b1 );
or ( \4439_b1 , \4429_b1 , \4438_b1 );
not ( \4438_b1 , w_7778 );
and ( \4439_b0 , \4429_b0 , w_7779 );
and ( w_7778 , w_7779 , \4438_b0 );
or ( \4440_b1 , \4428_b1 , w_7780 );
or ( \4440_b0 , \4428_b0 , \4439_b0 );
not ( \4439_b0 , w_7781 );
and ( w_7781 , w_7780 , \4439_b1 );
or ( \4441_b1 , \4425_b1 , \4440_b1 );
not ( \4440_b1 , w_7782 );
and ( \4441_b0 , \4425_b0 , w_7783 );
and ( w_7782 , w_7783 , \4440_b0 );
or ( \4442_b1 , \4424_b1 , w_7784 );
or ( \4442_b0 , \4424_b0 , \4441_b0 );
not ( \4441_b0 , w_7785 );
and ( w_7785 , w_7784 , \4441_b1 );
or ( \4443_b1 , \4421_b1 , \4442_b1 );
not ( \4442_b1 , w_7786 );
and ( \4443_b0 , \4421_b0 , w_7787 );
and ( w_7786 , w_7787 , \4442_b0 );
or ( \4444_b1 , \4420_b1 , w_7788 );
or ( \4444_b0 , \4420_b0 , \4443_b0 );
not ( \4443_b0 , w_7789 );
and ( w_7789 , w_7788 , \4443_b1 );
or ( \4445_b1 , \4417_b1 , \4444_b1 );
not ( \4444_b1 , w_7790 );
and ( \4445_b0 , \4417_b0 , w_7791 );
and ( w_7790 , w_7791 , \4444_b0 );
or ( \4446_b1 , \4416_b1 , w_7792 );
or ( \4446_b0 , \4416_b0 , \4445_b0 );
not ( \4445_b0 , w_7793 );
and ( w_7793 , w_7792 , \4445_b1 );
or ( \4447_b1 , \4413_b1 , \4446_b1 );
not ( \4446_b1 , w_7794 );
and ( \4447_b0 , \4413_b0 , w_7795 );
and ( w_7794 , w_7795 , \4446_b0 );
or ( \4448_b1 , \4412_b1 , w_7796 );
or ( \4448_b0 , \4412_b0 , \4447_b0 );
not ( \4447_b0 , w_7797 );
and ( w_7797 , w_7796 , \4447_b1 );
or ( \4449_b1 , \4409_b1 , \4448_b1 );
not ( \4448_b1 , w_7798 );
and ( \4449_b0 , \4409_b0 , w_7799 );
and ( w_7798 , w_7799 , \4448_b0 );
or ( \4450_b1 , \4408_b1 , w_7800 );
or ( \4450_b0 , \4408_b0 , \4449_b0 );
not ( \4449_b0 , w_7801 );
and ( w_7801 , w_7800 , \4449_b1 );
or ( \4451_b1 , \4405_b1 , \4450_b1 );
not ( \4450_b1 , w_7802 );
and ( \4451_b0 , \4405_b0 , w_7803 );
and ( w_7802 , w_7803 , \4450_b0 );
or ( \4452_b1 , \4404_b1 , w_7804 );
or ( \4452_b0 , \4404_b0 , \4451_b0 );
not ( \4451_b0 , w_7805 );
and ( w_7805 , w_7804 , \4451_b1 );
or ( \4453_b1 , \4401_b1 , \4452_b1 );
not ( \4452_b1 , w_7806 );
and ( \4453_b0 , \4401_b0 , w_7807 );
and ( w_7806 , w_7807 , \4452_b0 );
or ( \4454_b1 , \4400_b1 , w_7808 );
or ( \4454_b0 , \4400_b0 , \4453_b0 );
not ( \4453_b0 , w_7809 );
and ( w_7809 , w_7808 , \4453_b1 );
or ( \4455_b1 , \4397_b1 , \4454_b1 );
not ( \4454_b1 , w_7810 );
and ( \4455_b0 , \4397_b0 , w_7811 );
and ( w_7810 , w_7811 , \4454_b0 );
or ( \4456_b1 , \4396_b1 , w_7812 );
or ( \4456_b0 , \4396_b0 , \4455_b0 );
not ( \4455_b0 , w_7813 );
and ( w_7813 , w_7812 , \4455_b1 );
or ( \4457_b1 , \4393_b1 , \4456_b1 );
not ( \4456_b1 , w_7814 );
and ( \4457_b0 , \4393_b0 , w_7815 );
and ( w_7814 , w_7815 , \4456_b0 );
or ( \4458_b1 , \4392_b1 , w_7816 );
or ( \4458_b0 , \4392_b0 , \4457_b0 );
not ( \4457_b0 , w_7817 );
and ( w_7817 , w_7816 , \4457_b1 );
or ( \4459_b1 , \4389_b1 , \4458_b1 );
not ( \4458_b1 , w_7818 );
and ( \4459_b0 , \4389_b0 , w_7819 );
and ( w_7818 , w_7819 , \4458_b0 );
or ( \4460_b1 , \4388_b1 , w_7820 );
or ( \4460_b0 , \4388_b0 , \4459_b0 );
not ( \4459_b0 , w_7821 );
and ( w_7821 , w_7820 , \4459_b1 );
or ( \4461_b1 , \4385_b1 , \4460_b1 );
not ( \4460_b1 , w_7822 );
and ( \4461_b0 , \4385_b0 , w_7823 );
and ( w_7822 , w_7823 , \4460_b0 );
or ( \4462_b1 , \4384_b1 , w_7824 );
or ( \4462_b0 , \4384_b0 , \4461_b0 );
not ( \4461_b0 , w_7825 );
and ( w_7825 , w_7824 , \4461_b1 );
or ( \4463_b1 , \4381_b1 , \4462_b1 );
not ( \4462_b1 , w_7826 );
and ( \4463_b0 , \4381_b0 , w_7827 );
and ( w_7826 , w_7827 , \4462_b0 );
or ( \4464_b1 , \4380_b1 , w_7828 );
or ( \4464_b0 , \4380_b0 , \4463_b0 );
not ( \4463_b0 , w_7829 );
and ( w_7829 , w_7828 , \4463_b1 );
or ( \4465_b1 , \4377_b1 , \4464_b1 );
not ( \4464_b1 , w_7830 );
and ( \4465_b0 , \4377_b0 , w_7831 );
and ( w_7830 , w_7831 , \4464_b0 );
or ( \4466_b1 , \4376_b1 , w_7832 );
or ( \4466_b0 , \4376_b0 , \4465_b0 );
not ( \4465_b0 , w_7833 );
and ( w_7833 , w_7832 , \4465_b1 );
or ( \4467_b1 , \4373_b1 , \4466_b1 );
xor ( \4467_b0 , \4373_b0 , w_7834 );
not ( w_7834 , w_7835 );
and ( w_7835 , \4466_b1 , \4466_b0 );
buf ( \4468_Z[31]_b1 , \4467_b1 );
buf ( \4468_Z[31]_b0 , \4467_b0 );
or ( \4469_b1 , \4377_b1 , \4464_b1 );
xor ( \4469_b0 , \4377_b0 , w_7836 );
not ( w_7836 , w_7837 );
and ( w_7837 , \4464_b1 , \4464_b0 );
buf ( \4470_Z[30]_b1 , \4469_b1 );
buf ( \4470_Z[30]_b0 , \4469_b0 );
or ( \4471_b1 , \4381_b1 , \4462_b1 );
xor ( \4471_b0 , \4381_b0 , w_7838 );
not ( w_7838 , w_7839 );
and ( w_7839 , \4462_b1 , \4462_b0 );
buf ( \4472_Z[29]_b1 , \4471_b1 );
buf ( \4472_Z[29]_b0 , \4471_b0 );
or ( \4473_b1 , \4385_b1 , \4460_b1 );
xor ( \4473_b0 , \4385_b0 , w_7840 );
not ( w_7840 , w_7841 );
and ( w_7841 , \4460_b1 , \4460_b0 );
buf ( \4474_Z[28]_b1 , \4473_b1 );
buf ( \4474_Z[28]_b0 , \4473_b0 );
or ( \4475_b1 , \4389_b1 , \4458_b1 );
xor ( \4475_b0 , \4389_b0 , w_7842 );
not ( w_7842 , w_7843 );
and ( w_7843 , \4458_b1 , \4458_b0 );
buf ( \4476_Z[27]_b1 , \4475_b1 );
buf ( \4476_Z[27]_b0 , \4475_b0 );
or ( \4477_b1 , \4393_b1 , \4456_b1 );
xor ( \4477_b0 , \4393_b0 , w_7844 );
not ( w_7844 , w_7845 );
and ( w_7845 , \4456_b1 , \4456_b0 );
buf ( \4478_Z[26]_b1 , \4477_b1 );
buf ( \4478_Z[26]_b0 , \4477_b0 );
or ( \4479_b1 , \4397_b1 , \4454_b1 );
xor ( \4479_b0 , \4397_b0 , w_7846 );
not ( w_7846 , w_7847 );
and ( w_7847 , \4454_b1 , \4454_b0 );
buf ( \4480_Z[25]_b1 , \4479_b1 );
buf ( \4480_Z[25]_b0 , \4479_b0 );
or ( \4481_b1 , \4401_b1 , \4452_b1 );
xor ( \4481_b0 , \4401_b0 , w_7848 );
not ( w_7848 , w_7849 );
and ( w_7849 , \4452_b1 , \4452_b0 );
buf ( \4482_Z[24]_b1 , \4481_b1 );
buf ( \4482_Z[24]_b0 , \4481_b0 );
or ( \4483_b1 , \4405_b1 , \4450_b1 );
xor ( \4483_b0 , \4405_b0 , w_7850 );
not ( w_7850 , w_7851 );
and ( w_7851 , \4450_b1 , \4450_b0 );
buf ( \4484_Z[23]_b1 , \4483_b1 );
buf ( \4484_Z[23]_b0 , \4483_b0 );
or ( \4485_b1 , \4409_b1 , \4448_b1 );
xor ( \4485_b0 , \4409_b0 , w_7852 );
not ( w_7852 , w_7853 );
and ( w_7853 , \4448_b1 , \4448_b0 );
buf ( \4486_Z[22]_b1 , \4485_b1 );
buf ( \4486_Z[22]_b0 , \4485_b0 );
or ( \4487_b1 , \4413_b1 , \4446_b1 );
xor ( \4487_b0 , \4413_b0 , w_7854 );
not ( w_7854 , w_7855 );
and ( w_7855 , \4446_b1 , \4446_b0 );
buf ( \4488_Z[21]_b1 , \4487_b1 );
buf ( \4488_Z[21]_b0 , \4487_b0 );
or ( \4489_b1 , \4417_b1 , \4444_b1 );
xor ( \4489_b0 , \4417_b0 , w_7856 );
not ( w_7856 , w_7857 );
and ( w_7857 , \4444_b1 , \4444_b0 );
buf ( \4490_Z[20]_b1 , \4489_b1 );
buf ( \4490_Z[20]_b0 , \4489_b0 );
or ( \4491_b1 , \4421_b1 , \4442_b1 );
xor ( \4491_b0 , \4421_b0 , w_7858 );
not ( w_7858 , w_7859 );
and ( w_7859 , \4442_b1 , \4442_b0 );
buf ( \4492_Z[19]_b1 , \4491_b1 );
buf ( \4492_Z[19]_b0 , \4491_b0 );
or ( \4493_b1 , \4425_b1 , \4440_b1 );
xor ( \4493_b0 , \4425_b0 , w_7860 );
not ( w_7860 , w_7861 );
and ( w_7861 , \4440_b1 , \4440_b0 );
buf ( \4494_Z[18]_b1 , \4493_b1 );
buf ( \4494_Z[18]_b0 , \4493_b0 );
or ( \4495_b1 , \4429_b1 , \4438_b1 );
xor ( \4495_b0 , \4429_b0 , w_7862 );
not ( w_7862 , w_7863 );
and ( w_7863 , \4438_b1 , \4438_b0 );
buf ( \4496_Z[17]_b1 , \4495_b1 );
buf ( \4496_Z[17]_b0 , \4495_b0 );
or ( \4497_b1 , \4433_b1 , \4436_b1 );
xor ( \4497_b0 , \4433_b0 , w_7864 );
not ( w_7864 , w_7865 );
and ( w_7865 , \4436_b1 , \4436_b0 );
buf ( \4498_Z[16]_b1 , \4497_b1 );
buf ( \4498_Z[16]_b0 , \4497_b0 );
or ( \4499_b1 , \4434_b1 , \4435_b1 );
xor ( \4499_b0 , \4434_b0 , w_7866 );
not ( w_7866 , w_7867 );
and ( w_7867 , \4435_b1 , \4435_b0 );
buf ( \4500_Z[15]_b1 , \4499_b1 );
buf ( \4500_Z[15]_b0 , \4499_b0 );
or ( \4501_b1 , \4337_b1 , \4338_b1 );
xor ( \4501_b0 , \4337_b0 , w_7868 );
not ( w_7868 , w_7869 );
and ( w_7869 , \4338_b1 , \4338_b0 );
buf ( \4502_Z[14]_b1 , \4501_b1 );
buf ( \4502_Z[14]_b0 , \4501_b0 );
or ( \4503_b1 , \4239_b1 , \4240_b1 );
xor ( \4503_b0 , \4239_b0 , w_7870 );
not ( w_7870 , w_7871 );
and ( w_7871 , \4240_b1 , \4240_b0 );
buf ( \4504_Z[13]_b1 , \4503_b1 );
buf ( \4504_Z[13]_b0 , \4503_b0 );
or ( \4505_b1 , \4141_b1 , \4142_b1 );
xor ( \4505_b0 , \4141_b0 , w_7872 );
not ( w_7872 , w_7873 );
and ( w_7873 , \4142_b1 , \4142_b0 );
buf ( \4506_Z[12]_b1 , \4505_b1 );
buf ( \4506_Z[12]_b0 , \4505_b0 );
or ( \4507_b1 , \4043_b1 , \4044_b1 );
xor ( \4507_b0 , \4043_b0 , w_7874 );
not ( w_7874 , w_7875 );
and ( w_7875 , \4044_b1 , \4044_b0 );
buf ( \4508_Z[11]_b1 , \4507_b1 );
buf ( \4508_Z[11]_b0 , \4507_b0 );
or ( \4509_b1 , \3945_b1 , \3946_b1 );
xor ( \4509_b0 , \3945_b0 , w_7876 );
not ( w_7876 , w_7877 );
and ( w_7877 , \3946_b1 , \3946_b0 );
buf ( \4510_Z[10]_b1 , \4509_b1 );
buf ( \4510_Z[10]_b0 , \4509_b0 );
or ( \4511_b1 , \3847_b1 , \3848_b1 );
xor ( \4511_b0 , \3847_b0 , w_7878 );
not ( w_7878 , w_7879 );
and ( w_7879 , \3848_b1 , \3848_b0 );
buf ( \4512_Z[9]_b1 , \4511_b1 );
buf ( \4512_Z[9]_b0 , \4511_b0 );
or ( \4513_b1 , \3749_b1 , \3750_b1 );
xor ( \4513_b0 , \3749_b0 , w_7880 );
not ( w_7880 , w_7881 );
and ( w_7881 , \3750_b1 , \3750_b0 );
buf ( \4514_Z[8]_b1 , \4513_b1 );
buf ( \4514_Z[8]_b0 , \4513_b0 );
or ( \4515_b1 , \3651_b1 , \3652_b1 );
xor ( \4515_b0 , \3651_b0 , w_7882 );
not ( w_7882 , w_7883 );
and ( w_7883 , \3652_b1 , \3652_b0 );
buf ( \4516_Z[7]_b1 , \4515_b1 );
buf ( \4516_Z[7]_b0 , \4515_b0 );
or ( \4517_b1 , \3553_b1 , \3554_b1 );
xor ( \4517_b0 , \3553_b0 , w_7884 );
not ( w_7884 , w_7885 );
and ( w_7885 , \3554_b1 , \3554_b0 );
buf ( \4518_Z[6]_b1 , \4517_b1 );
buf ( \4518_Z[6]_b0 , \4517_b0 );
or ( \4519_b1 , \3455_b1 , \3456_b1 );
xor ( \4519_b0 , \3455_b0 , w_7886 );
not ( w_7886 , w_7887 );
and ( w_7887 , \3456_b1 , \3456_b0 );
buf ( \4520_Z[5]_b1 , \4519_b1 );
buf ( \4520_Z[5]_b0 , \4519_b0 );
or ( \4521_b1 , \3357_b1 , \3358_b1 );
xor ( \4521_b0 , \3357_b0 , w_7888 );
not ( w_7888 , w_7889 );
and ( w_7889 , \3358_b1 , \3358_b0 );
buf ( \4522_Z[4]_b1 , \4521_b1 );
buf ( \4522_Z[4]_b0 , \4521_b0 );
or ( \4523_b1 , \3259_b1 , \3260_b1 );
xor ( \4523_b0 , \3259_b0 , w_7890 );
not ( w_7890 , w_7891 );
and ( w_7891 , \3260_b1 , \3260_b0 );
buf ( \4524_Z[3]_b1 , \4523_b1 );
buf ( \4524_Z[3]_b0 , \4523_b0 );
or ( \4525_b1 , \3161_b1 , \3162_b1 );
xor ( \4525_b0 , \3161_b0 , w_7892 );
not ( w_7892 , w_7893 );
and ( w_7893 , \3162_b1 , \3162_b0 );
buf ( \4526_Z[2]_b1 , \4525_b1 );
buf ( \4526_Z[2]_b0 , \4525_b0 );
or ( \4527_b1 , \3064_b1 , \3065_b1 );
xor ( \4527_b0 , \3064_b0 , w_7894 );
not ( w_7894 , w_7895 );
and ( w_7895 , \3065_b1 , \3065_b0 );
buf ( \4528_Z[1]_b1 , \4527_b1 );
buf ( \4528_Z[1]_b0 , \4527_b0 );
or ( \4529_b1 , \2986_A[0]_b1 , \3002_B[0]_b1 );
not ( \3002_B[0]_b1 , w_7896 );
and ( \4529_b0 , \2986_A[0]_b0 , w_7897 );
and ( w_7896 , w_7897 , \3002_B[0]_b0 );
buf ( \4530_Z[0]_b1 , \4529_b1 );
buf ( \4530_Z[0]_b0 , \4529_b0 );
or ( \853_b1 , \160_b1 , w_7928 );
or ( \853_b0 , \160_b0 , w_7899 );
not ( w_7899 , w_7929 );
and ( w_7929 , w_7928 , w_7898 );
or ( w_7898 , \166_Z[1]_b1 , w_7930 );
or ( w_7899 , \166_Z[1]_b0 , w_7901 );
not ( w_7901 , w_7931 );
and ( w_7931 , w_7930 , w_7900 );
or ( w_7900 , \176_Z[2]_b1 , w_7932 );
or ( w_7901 , \176_Z[2]_b0 , w_7903 );
not ( w_7903 , w_7933 );
and ( w_7933 , w_7932 , w_7902 );
or ( w_7902 , \192_Z[3]_b1 , w_7934 );
or ( w_7903 , \192_Z[3]_b0 , w_7905 );
not ( w_7905 , w_7935 );
and ( w_7935 , w_7934 , w_7904 );
or ( w_7904 , \214_Z[4]_b1 , w_7936 );
or ( w_7905 , \214_Z[4]_b0 , w_7907 );
not ( w_7907 , w_7937 );
and ( w_7937 , w_7936 , w_7906 );
or ( w_7906 , \242_Z[5]_b1 , w_7938 );
or ( w_7907 , \242_Z[5]_b0 , w_7909 );
not ( w_7909 , w_7939 );
and ( w_7939 , w_7938 , w_7908 );
or ( w_7908 , \276_Z[6]_b1 , w_7940 );
or ( w_7909 , \276_Z[6]_b0 , w_7911 );
not ( w_7911 , w_7941 );
and ( w_7941 , w_7940 , w_7910 );
or ( w_7910 , \316_Z[7]_b1 , w_7942 );
or ( w_7911 , \316_Z[7]_b0 , w_7913 );
not ( w_7913 , w_7943 );
and ( w_7943 , w_7942 , w_7912 );
or ( w_7912 , \362_Z[8]_b1 , w_7944 );
or ( w_7913 , \362_Z[8]_b0 , w_7915 );
not ( w_7915 , w_7945 );
and ( w_7945 , w_7944 , w_7914 );
or ( w_7914 , \414_Z[9]_b1 , w_7946 );
or ( w_7915 , \414_Z[9]_b0 , w_7917 );
not ( w_7917 , w_7947 );
and ( w_7947 , w_7946 , w_7916 );
or ( w_7916 , \472_Z[10]_b1 , w_7948 );
or ( w_7917 , \472_Z[10]_b0 , w_7919 );
not ( w_7919 , w_7949 );
and ( w_7949 , w_7948 , w_7918 );
or ( w_7918 , \536_Z[11]_b1 , w_7950 );
or ( w_7919 , \536_Z[11]_b0 , w_7921 );
not ( w_7921 , w_7951 );
and ( w_7951 , w_7950 , w_7920 );
or ( w_7920 , \606_Z[12]_b1 , w_7952 );
or ( w_7921 , \606_Z[12]_b0 , w_7923 );
not ( w_7923 , w_7953 );
and ( w_7953 , w_7952 , w_7922 );
or ( w_7922 , \682_Z[13]_b1 , w_7954 );
or ( w_7923 , \682_Z[13]_b0 , w_7925 );
not ( w_7925 , w_7955 );
and ( w_7955 , w_7954 , w_7924 );
or ( w_7924 , \764_Z[14]_b1 , w_7956 );
or ( w_7925 , \764_Z[14]_b0 , w_7927 );
not ( w_7927 , w_7957 );
and ( w_7957 , w_7956 , w_7926 );
buf ( w_7926 , \852_Z[15]_b1 );
not ( w_7926 , w_7958 );
not ( w_7927 , w_7959 );
and ( w_7958 , w_7959 , \852_Z[15]_b0 );
or ( \855_b1 , \159_Z[0]_b1 , w_7990 );
or ( \855_b0 , \159_Z[0]_b0 , w_7961 );
not ( w_7961 , w_7991 );
and ( w_7991 , w_7990 , w_7960 );
or ( w_7960 , \854_b1 , w_7992 );
or ( w_7961 , \854_b0 , w_7963 );
not ( w_7963 , w_7993 );
and ( w_7993 , w_7992 , w_7962 );
or ( w_7962 , \176_Z[2]_b1 , w_7994 );
or ( w_7963 , \176_Z[2]_b0 , w_7965 );
not ( w_7965 , w_7995 );
and ( w_7995 , w_7994 , w_7964 );
or ( w_7964 , \192_Z[3]_b1 , w_7996 );
or ( w_7965 , \192_Z[3]_b0 , w_7967 );
not ( w_7967 , w_7997 );
and ( w_7997 , w_7996 , w_7966 );
or ( w_7966 , \214_Z[4]_b1 , w_7998 );
or ( w_7967 , \214_Z[4]_b0 , w_7969 );
not ( w_7969 , w_7999 );
and ( w_7999 , w_7998 , w_7968 );
or ( w_7968 , \242_Z[5]_b1 , w_8000 );
or ( w_7969 , \242_Z[5]_b0 , w_7971 );
not ( w_7971 , w_8001 );
and ( w_8001 , w_8000 , w_7970 );
or ( w_7970 , \276_Z[6]_b1 , w_8002 );
or ( w_7971 , \276_Z[6]_b0 , w_7973 );
not ( w_7973 , w_8003 );
and ( w_8003 , w_8002 , w_7972 );
or ( w_7972 , \316_Z[7]_b1 , w_8004 );
or ( w_7973 , \316_Z[7]_b0 , w_7975 );
not ( w_7975 , w_8005 );
and ( w_8005 , w_8004 , w_7974 );
or ( w_7974 , \362_Z[8]_b1 , w_8006 );
or ( w_7975 , \362_Z[8]_b0 , w_7977 );
not ( w_7977 , w_8007 );
and ( w_8007 , w_8006 , w_7976 );
or ( w_7976 , \414_Z[9]_b1 , w_8008 );
or ( w_7977 , \414_Z[9]_b0 , w_7979 );
not ( w_7979 , w_8009 );
and ( w_8009 , w_8008 , w_7978 );
or ( w_7978 , \472_Z[10]_b1 , w_8010 );
or ( w_7979 , \472_Z[10]_b0 , w_7981 );
not ( w_7981 , w_8011 );
and ( w_8011 , w_8010 , w_7980 );
or ( w_7980 , \536_Z[11]_b1 , w_8012 );
or ( w_7981 , \536_Z[11]_b0 , w_7983 );
not ( w_7983 , w_8013 );
and ( w_8013 , w_8012 , w_7982 );
or ( w_7982 , \606_Z[12]_b1 , w_8014 );
or ( w_7983 , \606_Z[12]_b0 , w_7985 );
not ( w_7985 , w_8015 );
and ( w_8015 , w_8014 , w_7984 );
or ( w_7984 , \682_Z[13]_b1 , w_8016 );
or ( w_7985 , \682_Z[13]_b0 , w_7987 );
not ( w_7987 , w_8017 );
and ( w_8017 , w_8016 , w_7986 );
or ( w_7986 , \764_Z[14]_b1 , w_8018 );
or ( w_7987 , \764_Z[14]_b0 , w_7989 );
not ( w_7989 , w_8019 );
and ( w_8019 , w_8018 , w_7988 );
buf ( w_7988 , \852_Z[15]_b1 );
not ( w_7988 , w_8020 );
not ( w_7989 , w_8021 );
and ( w_8020 , w_8021 , \852_Z[15]_b0 );
or ( \857_b1 , \159_Z[0]_b1 , w_8052 );
or ( \857_b0 , \159_Z[0]_b0 , w_8023 );
not ( w_8023 , w_8053 );
and ( w_8053 , w_8052 , w_8022 );
or ( w_8022 , \166_Z[1]_b1 , w_8054 );
or ( w_8023 , \166_Z[1]_b0 , w_8025 );
not ( w_8025 , w_8055 );
and ( w_8055 , w_8054 , w_8024 );
or ( w_8024 , \856_b1 , w_8056 );
or ( w_8025 , \856_b0 , w_8027 );
not ( w_8027 , w_8057 );
and ( w_8057 , w_8056 , w_8026 );
or ( w_8026 , \192_Z[3]_b1 , w_8058 );
or ( w_8027 , \192_Z[3]_b0 , w_8029 );
not ( w_8029 , w_8059 );
and ( w_8059 , w_8058 , w_8028 );
or ( w_8028 , \214_Z[4]_b1 , w_8060 );
or ( w_8029 , \214_Z[4]_b0 , w_8031 );
not ( w_8031 , w_8061 );
and ( w_8061 , w_8060 , w_8030 );
or ( w_8030 , \242_Z[5]_b1 , w_8062 );
or ( w_8031 , \242_Z[5]_b0 , w_8033 );
not ( w_8033 , w_8063 );
and ( w_8063 , w_8062 , w_8032 );
or ( w_8032 , \276_Z[6]_b1 , w_8064 );
or ( w_8033 , \276_Z[6]_b0 , w_8035 );
not ( w_8035 , w_8065 );
and ( w_8065 , w_8064 , w_8034 );
or ( w_8034 , \316_Z[7]_b1 , w_8066 );
or ( w_8035 , \316_Z[7]_b0 , w_8037 );
not ( w_8037 , w_8067 );
and ( w_8067 , w_8066 , w_8036 );
or ( w_8036 , \362_Z[8]_b1 , w_8068 );
or ( w_8037 , \362_Z[8]_b0 , w_8039 );
not ( w_8039 , w_8069 );
and ( w_8069 , w_8068 , w_8038 );
or ( w_8038 , \414_Z[9]_b1 , w_8070 );
or ( w_8039 , \414_Z[9]_b0 , w_8041 );
not ( w_8041 , w_8071 );
and ( w_8071 , w_8070 , w_8040 );
or ( w_8040 , \472_Z[10]_b1 , w_8072 );
or ( w_8041 , \472_Z[10]_b0 , w_8043 );
not ( w_8043 , w_8073 );
and ( w_8073 , w_8072 , w_8042 );
or ( w_8042 , \536_Z[11]_b1 , w_8074 );
or ( w_8043 , \536_Z[11]_b0 , w_8045 );
not ( w_8045 , w_8075 );
and ( w_8075 , w_8074 , w_8044 );
or ( w_8044 , \606_Z[12]_b1 , w_8076 );
or ( w_8045 , \606_Z[12]_b0 , w_8047 );
not ( w_8047 , w_8077 );
and ( w_8077 , w_8076 , w_8046 );
or ( w_8046 , \682_Z[13]_b1 , w_8078 );
or ( w_8047 , \682_Z[13]_b0 , w_8049 );
not ( w_8049 , w_8079 );
and ( w_8079 , w_8078 , w_8048 );
or ( w_8048 , \764_Z[14]_b1 , w_8080 );
or ( w_8049 , \764_Z[14]_b0 , w_8051 );
not ( w_8051 , w_8081 );
and ( w_8081 , w_8080 , w_8050 );
buf ( w_8050 , \852_Z[15]_b1 );
not ( w_8050 , w_8082 );
not ( w_8051 , w_8083 );
and ( w_8082 , w_8083 , \852_Z[15]_b0 );
or ( \859_b1 , \159_Z[0]_b1 , w_8114 );
or ( \859_b0 , \159_Z[0]_b0 , w_8085 );
not ( w_8085 , w_8115 );
and ( w_8115 , w_8114 , w_8084 );
or ( w_8084 , \166_Z[1]_b1 , w_8116 );
or ( w_8085 , \166_Z[1]_b0 , w_8087 );
not ( w_8087 , w_8117 );
and ( w_8117 , w_8116 , w_8086 );
or ( w_8086 , \176_Z[2]_b1 , w_8118 );
or ( w_8087 , \176_Z[2]_b0 , w_8089 );
not ( w_8089 , w_8119 );
and ( w_8119 , w_8118 , w_8088 );
or ( w_8088 , \858_b1 , w_8120 );
or ( w_8089 , \858_b0 , w_8091 );
not ( w_8091 , w_8121 );
and ( w_8121 , w_8120 , w_8090 );
or ( w_8090 , \214_Z[4]_b1 , w_8122 );
or ( w_8091 , \214_Z[4]_b0 , w_8093 );
not ( w_8093 , w_8123 );
and ( w_8123 , w_8122 , w_8092 );
or ( w_8092 , \242_Z[5]_b1 , w_8124 );
or ( w_8093 , \242_Z[5]_b0 , w_8095 );
not ( w_8095 , w_8125 );
and ( w_8125 , w_8124 , w_8094 );
or ( w_8094 , \276_Z[6]_b1 , w_8126 );
or ( w_8095 , \276_Z[6]_b0 , w_8097 );
not ( w_8097 , w_8127 );
and ( w_8127 , w_8126 , w_8096 );
or ( w_8096 , \316_Z[7]_b1 , w_8128 );
or ( w_8097 , \316_Z[7]_b0 , w_8099 );
not ( w_8099 , w_8129 );
and ( w_8129 , w_8128 , w_8098 );
or ( w_8098 , \362_Z[8]_b1 , w_8130 );
or ( w_8099 , \362_Z[8]_b0 , w_8101 );
not ( w_8101 , w_8131 );
and ( w_8131 , w_8130 , w_8100 );
or ( w_8100 , \414_Z[9]_b1 , w_8132 );
or ( w_8101 , \414_Z[9]_b0 , w_8103 );
not ( w_8103 , w_8133 );
and ( w_8133 , w_8132 , w_8102 );
or ( w_8102 , \472_Z[10]_b1 , w_8134 );
or ( w_8103 , \472_Z[10]_b0 , w_8105 );
not ( w_8105 , w_8135 );
and ( w_8135 , w_8134 , w_8104 );
or ( w_8104 , \536_Z[11]_b1 , w_8136 );
or ( w_8105 , \536_Z[11]_b0 , w_8107 );
not ( w_8107 , w_8137 );
and ( w_8137 , w_8136 , w_8106 );
or ( w_8106 , \606_Z[12]_b1 , w_8138 );
or ( w_8107 , \606_Z[12]_b0 , w_8109 );
not ( w_8109 , w_8139 );
and ( w_8139 , w_8138 , w_8108 );
or ( w_8108 , \682_Z[13]_b1 , w_8140 );
or ( w_8109 , \682_Z[13]_b0 , w_8111 );
not ( w_8111 , w_8141 );
and ( w_8141 , w_8140 , w_8110 );
or ( w_8110 , \764_Z[14]_b1 , w_8142 );
or ( w_8111 , \764_Z[14]_b0 , w_8113 );
not ( w_8113 , w_8143 );
and ( w_8143 , w_8142 , w_8112 );
buf ( w_8112 , \852_Z[15]_b1 );
not ( w_8112 , w_8144 );
not ( w_8113 , w_8145 );
and ( w_8144 , w_8145 , \852_Z[15]_b0 );
or ( \861_b1 , \159_Z[0]_b1 , w_8176 );
or ( \861_b0 , \159_Z[0]_b0 , w_8147 );
not ( w_8147 , w_8177 );
and ( w_8177 , w_8176 , w_8146 );
or ( w_8146 , \166_Z[1]_b1 , w_8178 );
or ( w_8147 , \166_Z[1]_b0 , w_8149 );
not ( w_8149 , w_8179 );
and ( w_8179 , w_8178 , w_8148 );
or ( w_8148 , \176_Z[2]_b1 , w_8180 );
or ( w_8149 , \176_Z[2]_b0 , w_8151 );
not ( w_8151 , w_8181 );
and ( w_8181 , w_8180 , w_8150 );
or ( w_8150 , \192_Z[3]_b1 , w_8182 );
or ( w_8151 , \192_Z[3]_b0 , w_8153 );
not ( w_8153 , w_8183 );
and ( w_8183 , w_8182 , w_8152 );
or ( w_8152 , \860_b1 , w_8184 );
or ( w_8153 , \860_b0 , w_8155 );
not ( w_8155 , w_8185 );
and ( w_8185 , w_8184 , w_8154 );
or ( w_8154 , \242_Z[5]_b1 , w_8186 );
or ( w_8155 , \242_Z[5]_b0 , w_8157 );
not ( w_8157 , w_8187 );
and ( w_8187 , w_8186 , w_8156 );
or ( w_8156 , \276_Z[6]_b1 , w_8188 );
or ( w_8157 , \276_Z[6]_b0 , w_8159 );
not ( w_8159 , w_8189 );
and ( w_8189 , w_8188 , w_8158 );
or ( w_8158 , \316_Z[7]_b1 , w_8190 );
or ( w_8159 , \316_Z[7]_b0 , w_8161 );
not ( w_8161 , w_8191 );
and ( w_8191 , w_8190 , w_8160 );
or ( w_8160 , \362_Z[8]_b1 , w_8192 );
or ( w_8161 , \362_Z[8]_b0 , w_8163 );
not ( w_8163 , w_8193 );
and ( w_8193 , w_8192 , w_8162 );
or ( w_8162 , \414_Z[9]_b1 , w_8194 );
or ( w_8163 , \414_Z[9]_b0 , w_8165 );
not ( w_8165 , w_8195 );
and ( w_8195 , w_8194 , w_8164 );
or ( w_8164 , \472_Z[10]_b1 , w_8196 );
or ( w_8165 , \472_Z[10]_b0 , w_8167 );
not ( w_8167 , w_8197 );
and ( w_8197 , w_8196 , w_8166 );
or ( w_8166 , \536_Z[11]_b1 , w_8198 );
or ( w_8167 , \536_Z[11]_b0 , w_8169 );
not ( w_8169 , w_8199 );
and ( w_8199 , w_8198 , w_8168 );
or ( w_8168 , \606_Z[12]_b1 , w_8200 );
or ( w_8169 , \606_Z[12]_b0 , w_8171 );
not ( w_8171 , w_8201 );
and ( w_8201 , w_8200 , w_8170 );
or ( w_8170 , \682_Z[13]_b1 , w_8202 );
or ( w_8171 , \682_Z[13]_b0 , w_8173 );
not ( w_8173 , w_8203 );
and ( w_8203 , w_8202 , w_8172 );
or ( w_8172 , \764_Z[14]_b1 , w_8204 );
or ( w_8173 , \764_Z[14]_b0 , w_8175 );
not ( w_8175 , w_8205 );
and ( w_8205 , w_8204 , w_8174 );
buf ( w_8174 , \852_Z[15]_b1 );
not ( w_8174 , w_8206 );
not ( w_8175 , w_8207 );
and ( w_8206 , w_8207 , \852_Z[15]_b0 );
or ( \863_b1 , \159_Z[0]_b1 , w_8238 );
or ( \863_b0 , \159_Z[0]_b0 , w_8209 );
not ( w_8209 , w_8239 );
and ( w_8239 , w_8238 , w_8208 );
or ( w_8208 , \166_Z[1]_b1 , w_8240 );
or ( w_8209 , \166_Z[1]_b0 , w_8211 );
not ( w_8211 , w_8241 );
and ( w_8241 , w_8240 , w_8210 );
or ( w_8210 , \176_Z[2]_b1 , w_8242 );
or ( w_8211 , \176_Z[2]_b0 , w_8213 );
not ( w_8213 , w_8243 );
and ( w_8243 , w_8242 , w_8212 );
or ( w_8212 , \192_Z[3]_b1 , w_8244 );
or ( w_8213 , \192_Z[3]_b0 , w_8215 );
not ( w_8215 , w_8245 );
and ( w_8245 , w_8244 , w_8214 );
or ( w_8214 , \214_Z[4]_b1 , w_8246 );
or ( w_8215 , \214_Z[4]_b0 , w_8217 );
not ( w_8217 , w_8247 );
and ( w_8247 , w_8246 , w_8216 );
or ( w_8216 , \862_b1 , w_8248 );
or ( w_8217 , \862_b0 , w_8219 );
not ( w_8219 , w_8249 );
and ( w_8249 , w_8248 , w_8218 );
or ( w_8218 , \276_Z[6]_b1 , w_8250 );
or ( w_8219 , \276_Z[6]_b0 , w_8221 );
not ( w_8221 , w_8251 );
and ( w_8251 , w_8250 , w_8220 );
or ( w_8220 , \316_Z[7]_b1 , w_8252 );
or ( w_8221 , \316_Z[7]_b0 , w_8223 );
not ( w_8223 , w_8253 );
and ( w_8253 , w_8252 , w_8222 );
or ( w_8222 , \362_Z[8]_b1 , w_8254 );
or ( w_8223 , \362_Z[8]_b0 , w_8225 );
not ( w_8225 , w_8255 );
and ( w_8255 , w_8254 , w_8224 );
or ( w_8224 , \414_Z[9]_b1 , w_8256 );
or ( w_8225 , \414_Z[9]_b0 , w_8227 );
not ( w_8227 , w_8257 );
and ( w_8257 , w_8256 , w_8226 );
or ( w_8226 , \472_Z[10]_b1 , w_8258 );
or ( w_8227 , \472_Z[10]_b0 , w_8229 );
not ( w_8229 , w_8259 );
and ( w_8259 , w_8258 , w_8228 );
or ( w_8228 , \536_Z[11]_b1 , w_8260 );
or ( w_8229 , \536_Z[11]_b0 , w_8231 );
not ( w_8231 , w_8261 );
and ( w_8261 , w_8260 , w_8230 );
or ( w_8230 , \606_Z[12]_b1 , w_8262 );
or ( w_8231 , \606_Z[12]_b0 , w_8233 );
not ( w_8233 , w_8263 );
and ( w_8263 , w_8262 , w_8232 );
or ( w_8232 , \682_Z[13]_b1 , w_8264 );
or ( w_8233 , \682_Z[13]_b0 , w_8235 );
not ( w_8235 , w_8265 );
and ( w_8265 , w_8264 , w_8234 );
or ( w_8234 , \764_Z[14]_b1 , w_8266 );
or ( w_8235 , \764_Z[14]_b0 , w_8237 );
not ( w_8237 , w_8267 );
and ( w_8267 , w_8266 , w_8236 );
buf ( w_8236 , \852_Z[15]_b1 );
not ( w_8236 , w_8268 );
not ( w_8237 , w_8269 );
and ( w_8268 , w_8269 , \852_Z[15]_b0 );
or ( \865_b1 , \159_Z[0]_b1 , w_8300 );
or ( \865_b0 , \159_Z[0]_b0 , w_8271 );
not ( w_8271 , w_8301 );
and ( w_8301 , w_8300 , w_8270 );
or ( w_8270 , \166_Z[1]_b1 , w_8302 );
or ( w_8271 , \166_Z[1]_b0 , w_8273 );
not ( w_8273 , w_8303 );
and ( w_8303 , w_8302 , w_8272 );
or ( w_8272 , \176_Z[2]_b1 , w_8304 );
or ( w_8273 , \176_Z[2]_b0 , w_8275 );
not ( w_8275 , w_8305 );
and ( w_8305 , w_8304 , w_8274 );
or ( w_8274 , \192_Z[3]_b1 , w_8306 );
or ( w_8275 , \192_Z[3]_b0 , w_8277 );
not ( w_8277 , w_8307 );
and ( w_8307 , w_8306 , w_8276 );
or ( w_8276 , \214_Z[4]_b1 , w_8308 );
or ( w_8277 , \214_Z[4]_b0 , w_8279 );
not ( w_8279 , w_8309 );
and ( w_8309 , w_8308 , w_8278 );
or ( w_8278 , \242_Z[5]_b1 , w_8310 );
or ( w_8279 , \242_Z[5]_b0 , w_8281 );
not ( w_8281 , w_8311 );
and ( w_8311 , w_8310 , w_8280 );
or ( w_8280 , \864_b1 , w_8312 );
or ( w_8281 , \864_b0 , w_8283 );
not ( w_8283 , w_8313 );
and ( w_8313 , w_8312 , w_8282 );
or ( w_8282 , \316_Z[7]_b1 , w_8314 );
or ( w_8283 , \316_Z[7]_b0 , w_8285 );
not ( w_8285 , w_8315 );
and ( w_8315 , w_8314 , w_8284 );
or ( w_8284 , \362_Z[8]_b1 , w_8316 );
or ( w_8285 , \362_Z[8]_b0 , w_8287 );
not ( w_8287 , w_8317 );
and ( w_8317 , w_8316 , w_8286 );
or ( w_8286 , \414_Z[9]_b1 , w_8318 );
or ( w_8287 , \414_Z[9]_b0 , w_8289 );
not ( w_8289 , w_8319 );
and ( w_8319 , w_8318 , w_8288 );
or ( w_8288 , \472_Z[10]_b1 , w_8320 );
or ( w_8289 , \472_Z[10]_b0 , w_8291 );
not ( w_8291 , w_8321 );
and ( w_8321 , w_8320 , w_8290 );
or ( w_8290 , \536_Z[11]_b1 , w_8322 );
or ( w_8291 , \536_Z[11]_b0 , w_8293 );
not ( w_8293 , w_8323 );
and ( w_8323 , w_8322 , w_8292 );
or ( w_8292 , \606_Z[12]_b1 , w_8324 );
or ( w_8293 , \606_Z[12]_b0 , w_8295 );
not ( w_8295 , w_8325 );
and ( w_8325 , w_8324 , w_8294 );
or ( w_8294 , \682_Z[13]_b1 , w_8326 );
or ( w_8295 , \682_Z[13]_b0 , w_8297 );
not ( w_8297 , w_8327 );
and ( w_8327 , w_8326 , w_8296 );
or ( w_8296 , \764_Z[14]_b1 , w_8328 );
or ( w_8297 , \764_Z[14]_b0 , w_8299 );
not ( w_8299 , w_8329 );
and ( w_8329 , w_8328 , w_8298 );
buf ( w_8298 , \852_Z[15]_b1 );
not ( w_8298 , w_8330 );
not ( w_8299 , w_8331 );
and ( w_8330 , w_8331 , \852_Z[15]_b0 );
or ( \867_b1 , \159_Z[0]_b1 , w_8362 );
or ( \867_b0 , \159_Z[0]_b0 , w_8333 );
not ( w_8333 , w_8363 );
and ( w_8363 , w_8362 , w_8332 );
or ( w_8332 , \166_Z[1]_b1 , w_8364 );
or ( w_8333 , \166_Z[1]_b0 , w_8335 );
not ( w_8335 , w_8365 );
and ( w_8365 , w_8364 , w_8334 );
or ( w_8334 , \176_Z[2]_b1 , w_8366 );
or ( w_8335 , \176_Z[2]_b0 , w_8337 );
not ( w_8337 , w_8367 );
and ( w_8367 , w_8366 , w_8336 );
or ( w_8336 , \192_Z[3]_b1 , w_8368 );
or ( w_8337 , \192_Z[3]_b0 , w_8339 );
not ( w_8339 , w_8369 );
and ( w_8369 , w_8368 , w_8338 );
or ( w_8338 , \214_Z[4]_b1 , w_8370 );
or ( w_8339 , \214_Z[4]_b0 , w_8341 );
not ( w_8341 , w_8371 );
and ( w_8371 , w_8370 , w_8340 );
or ( w_8340 , \242_Z[5]_b1 , w_8372 );
or ( w_8341 , \242_Z[5]_b0 , w_8343 );
not ( w_8343 , w_8373 );
and ( w_8373 , w_8372 , w_8342 );
or ( w_8342 , \276_Z[6]_b1 , w_8374 );
or ( w_8343 , \276_Z[6]_b0 , w_8345 );
not ( w_8345 , w_8375 );
and ( w_8375 , w_8374 , w_8344 );
or ( w_8344 , \866_b1 , w_8376 );
or ( w_8345 , \866_b0 , w_8347 );
not ( w_8347 , w_8377 );
and ( w_8377 , w_8376 , w_8346 );
or ( w_8346 , \362_Z[8]_b1 , w_8378 );
or ( w_8347 , \362_Z[8]_b0 , w_8349 );
not ( w_8349 , w_8379 );
and ( w_8379 , w_8378 , w_8348 );
or ( w_8348 , \414_Z[9]_b1 , w_8380 );
or ( w_8349 , \414_Z[9]_b0 , w_8351 );
not ( w_8351 , w_8381 );
and ( w_8381 , w_8380 , w_8350 );
or ( w_8350 , \472_Z[10]_b1 , w_8382 );
or ( w_8351 , \472_Z[10]_b0 , w_8353 );
not ( w_8353 , w_8383 );
and ( w_8383 , w_8382 , w_8352 );
or ( w_8352 , \536_Z[11]_b1 , w_8384 );
or ( w_8353 , \536_Z[11]_b0 , w_8355 );
not ( w_8355 , w_8385 );
and ( w_8385 , w_8384 , w_8354 );
or ( w_8354 , \606_Z[12]_b1 , w_8386 );
or ( w_8355 , \606_Z[12]_b0 , w_8357 );
not ( w_8357 , w_8387 );
and ( w_8387 , w_8386 , w_8356 );
or ( w_8356 , \682_Z[13]_b1 , w_8388 );
or ( w_8357 , \682_Z[13]_b0 , w_8359 );
not ( w_8359 , w_8389 );
and ( w_8389 , w_8388 , w_8358 );
or ( w_8358 , \764_Z[14]_b1 , w_8390 );
or ( w_8359 , \764_Z[14]_b0 , w_8361 );
not ( w_8361 , w_8391 );
and ( w_8391 , w_8390 , w_8360 );
buf ( w_8360 , \852_Z[15]_b1 );
not ( w_8360 , w_8392 );
not ( w_8361 , w_8393 );
and ( w_8392 , w_8393 , \852_Z[15]_b0 );
or ( \869_b1 , \159_Z[0]_b1 , w_8424 );
or ( \869_b0 , \159_Z[0]_b0 , w_8395 );
not ( w_8395 , w_8425 );
and ( w_8425 , w_8424 , w_8394 );
or ( w_8394 , \166_Z[1]_b1 , w_8426 );
or ( w_8395 , \166_Z[1]_b0 , w_8397 );
not ( w_8397 , w_8427 );
and ( w_8427 , w_8426 , w_8396 );
or ( w_8396 , \176_Z[2]_b1 , w_8428 );
or ( w_8397 , \176_Z[2]_b0 , w_8399 );
not ( w_8399 , w_8429 );
and ( w_8429 , w_8428 , w_8398 );
or ( w_8398 , \192_Z[3]_b1 , w_8430 );
or ( w_8399 , \192_Z[3]_b0 , w_8401 );
not ( w_8401 , w_8431 );
and ( w_8431 , w_8430 , w_8400 );
or ( w_8400 , \214_Z[4]_b1 , w_8432 );
or ( w_8401 , \214_Z[4]_b0 , w_8403 );
not ( w_8403 , w_8433 );
and ( w_8433 , w_8432 , w_8402 );
or ( w_8402 , \242_Z[5]_b1 , w_8434 );
or ( w_8403 , \242_Z[5]_b0 , w_8405 );
not ( w_8405 , w_8435 );
and ( w_8435 , w_8434 , w_8404 );
or ( w_8404 , \276_Z[6]_b1 , w_8436 );
or ( w_8405 , \276_Z[6]_b0 , w_8407 );
not ( w_8407 , w_8437 );
and ( w_8437 , w_8436 , w_8406 );
or ( w_8406 , \316_Z[7]_b1 , w_8438 );
or ( w_8407 , \316_Z[7]_b0 , w_8409 );
not ( w_8409 , w_8439 );
and ( w_8439 , w_8438 , w_8408 );
or ( w_8408 , \868_b1 , w_8440 );
or ( w_8409 , \868_b0 , w_8411 );
not ( w_8411 , w_8441 );
and ( w_8441 , w_8440 , w_8410 );
or ( w_8410 , \414_Z[9]_b1 , w_8442 );
or ( w_8411 , \414_Z[9]_b0 , w_8413 );
not ( w_8413 , w_8443 );
and ( w_8443 , w_8442 , w_8412 );
or ( w_8412 , \472_Z[10]_b1 , w_8444 );
or ( w_8413 , \472_Z[10]_b0 , w_8415 );
not ( w_8415 , w_8445 );
and ( w_8445 , w_8444 , w_8414 );
or ( w_8414 , \536_Z[11]_b1 , w_8446 );
or ( w_8415 , \536_Z[11]_b0 , w_8417 );
not ( w_8417 , w_8447 );
and ( w_8447 , w_8446 , w_8416 );
or ( w_8416 , \606_Z[12]_b1 , w_8448 );
or ( w_8417 , \606_Z[12]_b0 , w_8419 );
not ( w_8419 , w_8449 );
and ( w_8449 , w_8448 , w_8418 );
or ( w_8418 , \682_Z[13]_b1 , w_8450 );
or ( w_8419 , \682_Z[13]_b0 , w_8421 );
not ( w_8421 , w_8451 );
and ( w_8451 , w_8450 , w_8420 );
or ( w_8420 , \764_Z[14]_b1 , w_8452 );
or ( w_8421 , \764_Z[14]_b0 , w_8423 );
not ( w_8423 , w_8453 );
and ( w_8453 , w_8452 , w_8422 );
buf ( w_8422 , \852_Z[15]_b1 );
not ( w_8422 , w_8454 );
not ( w_8423 , w_8455 );
and ( w_8454 , w_8455 , \852_Z[15]_b0 );
or ( \871_b1 , \159_Z[0]_b1 , w_8486 );
or ( \871_b0 , \159_Z[0]_b0 , w_8457 );
not ( w_8457 , w_8487 );
and ( w_8487 , w_8486 , w_8456 );
or ( w_8456 , \166_Z[1]_b1 , w_8488 );
or ( w_8457 , \166_Z[1]_b0 , w_8459 );
not ( w_8459 , w_8489 );
and ( w_8489 , w_8488 , w_8458 );
or ( w_8458 , \176_Z[2]_b1 , w_8490 );
or ( w_8459 , \176_Z[2]_b0 , w_8461 );
not ( w_8461 , w_8491 );
and ( w_8491 , w_8490 , w_8460 );
or ( w_8460 , \192_Z[3]_b1 , w_8492 );
or ( w_8461 , \192_Z[3]_b0 , w_8463 );
not ( w_8463 , w_8493 );
and ( w_8493 , w_8492 , w_8462 );
or ( w_8462 , \214_Z[4]_b1 , w_8494 );
or ( w_8463 , \214_Z[4]_b0 , w_8465 );
not ( w_8465 , w_8495 );
and ( w_8495 , w_8494 , w_8464 );
or ( w_8464 , \242_Z[5]_b1 , w_8496 );
or ( w_8465 , \242_Z[5]_b0 , w_8467 );
not ( w_8467 , w_8497 );
and ( w_8497 , w_8496 , w_8466 );
or ( w_8466 , \276_Z[6]_b1 , w_8498 );
or ( w_8467 , \276_Z[6]_b0 , w_8469 );
not ( w_8469 , w_8499 );
and ( w_8499 , w_8498 , w_8468 );
or ( w_8468 , \316_Z[7]_b1 , w_8500 );
or ( w_8469 , \316_Z[7]_b0 , w_8471 );
not ( w_8471 , w_8501 );
and ( w_8501 , w_8500 , w_8470 );
or ( w_8470 , \362_Z[8]_b1 , w_8502 );
or ( w_8471 , \362_Z[8]_b0 , w_8473 );
not ( w_8473 , w_8503 );
and ( w_8503 , w_8502 , w_8472 );
or ( w_8472 , \870_b1 , w_8504 );
or ( w_8473 , \870_b0 , w_8475 );
not ( w_8475 , w_8505 );
and ( w_8505 , w_8504 , w_8474 );
or ( w_8474 , \472_Z[10]_b1 , w_8506 );
or ( w_8475 , \472_Z[10]_b0 , w_8477 );
not ( w_8477 , w_8507 );
and ( w_8507 , w_8506 , w_8476 );
or ( w_8476 , \536_Z[11]_b1 , w_8508 );
or ( w_8477 , \536_Z[11]_b0 , w_8479 );
not ( w_8479 , w_8509 );
and ( w_8509 , w_8508 , w_8478 );
or ( w_8478 , \606_Z[12]_b1 , w_8510 );
or ( w_8479 , \606_Z[12]_b0 , w_8481 );
not ( w_8481 , w_8511 );
and ( w_8511 , w_8510 , w_8480 );
or ( w_8480 , \682_Z[13]_b1 , w_8512 );
or ( w_8481 , \682_Z[13]_b0 , w_8483 );
not ( w_8483 , w_8513 );
and ( w_8513 , w_8512 , w_8482 );
or ( w_8482 , \764_Z[14]_b1 , w_8514 );
or ( w_8483 , \764_Z[14]_b0 , w_8485 );
not ( w_8485 , w_8515 );
and ( w_8515 , w_8514 , w_8484 );
buf ( w_8484 , \852_Z[15]_b1 );
not ( w_8484 , w_8516 );
not ( w_8485 , w_8517 );
and ( w_8516 , w_8517 , \852_Z[15]_b0 );
or ( \873_b1 , \159_Z[0]_b1 , w_8548 );
or ( \873_b0 , \159_Z[0]_b0 , w_8519 );
not ( w_8519 , w_8549 );
and ( w_8549 , w_8548 , w_8518 );
or ( w_8518 , \166_Z[1]_b1 , w_8550 );
or ( w_8519 , \166_Z[1]_b0 , w_8521 );
not ( w_8521 , w_8551 );
and ( w_8551 , w_8550 , w_8520 );
or ( w_8520 , \176_Z[2]_b1 , w_8552 );
or ( w_8521 , \176_Z[2]_b0 , w_8523 );
not ( w_8523 , w_8553 );
and ( w_8553 , w_8552 , w_8522 );
or ( w_8522 , \192_Z[3]_b1 , w_8554 );
or ( w_8523 , \192_Z[3]_b0 , w_8525 );
not ( w_8525 , w_8555 );
and ( w_8555 , w_8554 , w_8524 );
or ( w_8524 , \214_Z[4]_b1 , w_8556 );
or ( w_8525 , \214_Z[4]_b0 , w_8527 );
not ( w_8527 , w_8557 );
and ( w_8557 , w_8556 , w_8526 );
or ( w_8526 , \242_Z[5]_b1 , w_8558 );
or ( w_8527 , \242_Z[5]_b0 , w_8529 );
not ( w_8529 , w_8559 );
and ( w_8559 , w_8558 , w_8528 );
or ( w_8528 , \276_Z[6]_b1 , w_8560 );
or ( w_8529 , \276_Z[6]_b0 , w_8531 );
not ( w_8531 , w_8561 );
and ( w_8561 , w_8560 , w_8530 );
or ( w_8530 , \316_Z[7]_b1 , w_8562 );
or ( w_8531 , \316_Z[7]_b0 , w_8533 );
not ( w_8533 , w_8563 );
and ( w_8563 , w_8562 , w_8532 );
or ( w_8532 , \362_Z[8]_b1 , w_8564 );
or ( w_8533 , \362_Z[8]_b0 , w_8535 );
not ( w_8535 , w_8565 );
and ( w_8565 , w_8564 , w_8534 );
or ( w_8534 , \414_Z[9]_b1 , w_8566 );
or ( w_8535 , \414_Z[9]_b0 , w_8537 );
not ( w_8537 , w_8567 );
and ( w_8567 , w_8566 , w_8536 );
or ( w_8536 , \872_b1 , w_8568 );
or ( w_8537 , \872_b0 , w_8539 );
not ( w_8539 , w_8569 );
and ( w_8569 , w_8568 , w_8538 );
or ( w_8538 , \536_Z[11]_b1 , w_8570 );
or ( w_8539 , \536_Z[11]_b0 , w_8541 );
not ( w_8541 , w_8571 );
and ( w_8571 , w_8570 , w_8540 );
or ( w_8540 , \606_Z[12]_b1 , w_8572 );
or ( w_8541 , \606_Z[12]_b0 , w_8543 );
not ( w_8543 , w_8573 );
and ( w_8573 , w_8572 , w_8542 );
or ( w_8542 , \682_Z[13]_b1 , w_8574 );
or ( w_8543 , \682_Z[13]_b0 , w_8545 );
not ( w_8545 , w_8575 );
and ( w_8575 , w_8574 , w_8544 );
or ( w_8544 , \764_Z[14]_b1 , w_8576 );
or ( w_8545 , \764_Z[14]_b0 , w_8547 );
not ( w_8547 , w_8577 );
and ( w_8577 , w_8576 , w_8546 );
buf ( w_8546 , \852_Z[15]_b1 );
not ( w_8546 , w_8578 );
not ( w_8547 , w_8579 );
and ( w_8578 , w_8579 , \852_Z[15]_b0 );
or ( \875_b1 , \159_Z[0]_b1 , w_8610 );
or ( \875_b0 , \159_Z[0]_b0 , w_8581 );
not ( w_8581 , w_8611 );
and ( w_8611 , w_8610 , w_8580 );
or ( w_8580 , \166_Z[1]_b1 , w_8612 );
or ( w_8581 , \166_Z[1]_b0 , w_8583 );
not ( w_8583 , w_8613 );
and ( w_8613 , w_8612 , w_8582 );
or ( w_8582 , \176_Z[2]_b1 , w_8614 );
or ( w_8583 , \176_Z[2]_b0 , w_8585 );
not ( w_8585 , w_8615 );
and ( w_8615 , w_8614 , w_8584 );
or ( w_8584 , \192_Z[3]_b1 , w_8616 );
or ( w_8585 , \192_Z[3]_b0 , w_8587 );
not ( w_8587 , w_8617 );
and ( w_8617 , w_8616 , w_8586 );
or ( w_8586 , \214_Z[4]_b1 , w_8618 );
or ( w_8587 , \214_Z[4]_b0 , w_8589 );
not ( w_8589 , w_8619 );
and ( w_8619 , w_8618 , w_8588 );
or ( w_8588 , \242_Z[5]_b1 , w_8620 );
or ( w_8589 , \242_Z[5]_b0 , w_8591 );
not ( w_8591 , w_8621 );
and ( w_8621 , w_8620 , w_8590 );
or ( w_8590 , \276_Z[6]_b1 , w_8622 );
or ( w_8591 , \276_Z[6]_b0 , w_8593 );
not ( w_8593 , w_8623 );
and ( w_8623 , w_8622 , w_8592 );
or ( w_8592 , \316_Z[7]_b1 , w_8624 );
or ( w_8593 , \316_Z[7]_b0 , w_8595 );
not ( w_8595 , w_8625 );
and ( w_8625 , w_8624 , w_8594 );
or ( w_8594 , \362_Z[8]_b1 , w_8626 );
or ( w_8595 , \362_Z[8]_b0 , w_8597 );
not ( w_8597 , w_8627 );
and ( w_8627 , w_8626 , w_8596 );
or ( w_8596 , \414_Z[9]_b1 , w_8628 );
or ( w_8597 , \414_Z[9]_b0 , w_8599 );
not ( w_8599 , w_8629 );
and ( w_8629 , w_8628 , w_8598 );
or ( w_8598 , \472_Z[10]_b1 , w_8630 );
or ( w_8599 , \472_Z[10]_b0 , w_8601 );
not ( w_8601 , w_8631 );
and ( w_8631 , w_8630 , w_8600 );
or ( w_8600 , \874_b1 , w_8632 );
or ( w_8601 , \874_b0 , w_8603 );
not ( w_8603 , w_8633 );
and ( w_8633 , w_8632 , w_8602 );
or ( w_8602 , \606_Z[12]_b1 , w_8634 );
or ( w_8603 , \606_Z[12]_b0 , w_8605 );
not ( w_8605 , w_8635 );
and ( w_8635 , w_8634 , w_8604 );
or ( w_8604 , \682_Z[13]_b1 , w_8636 );
or ( w_8605 , \682_Z[13]_b0 , w_8607 );
not ( w_8607 , w_8637 );
and ( w_8637 , w_8636 , w_8606 );
or ( w_8606 , \764_Z[14]_b1 , w_8638 );
or ( w_8607 , \764_Z[14]_b0 , w_8609 );
not ( w_8609 , w_8639 );
and ( w_8639 , w_8638 , w_8608 );
buf ( w_8608 , \852_Z[15]_b1 );
not ( w_8608 , w_8640 );
not ( w_8609 , w_8641 );
and ( w_8640 , w_8641 , \852_Z[15]_b0 );
or ( \876_b1 , \853_b1 , w_8664 );
or ( \876_b0 , \853_b0 , w_8643 );
not ( w_8643 , w_8665 );
and ( w_8665 , w_8664 , w_8642 );
or ( w_8642 , \855_b1 , w_8666 );
or ( w_8643 , \855_b0 , w_8645 );
not ( w_8645 , w_8667 );
and ( w_8667 , w_8666 , w_8644 );
or ( w_8644 , \857_b1 , w_8668 );
or ( w_8645 , \857_b0 , w_8647 );
not ( w_8647 , w_8669 );
and ( w_8669 , w_8668 , w_8646 );
or ( w_8646 , \859_b1 , w_8670 );
or ( w_8647 , \859_b0 , w_8649 );
not ( w_8649 , w_8671 );
and ( w_8671 , w_8670 , w_8648 );
or ( w_8648 , \861_b1 , w_8672 );
or ( w_8649 , \861_b0 , w_8651 );
not ( w_8651 , w_8673 );
and ( w_8673 , w_8672 , w_8650 );
or ( w_8650 , \863_b1 , w_8674 );
or ( w_8651 , \863_b0 , w_8653 );
not ( w_8653 , w_8675 );
and ( w_8675 , w_8674 , w_8652 );
or ( w_8652 , \865_b1 , w_8676 );
or ( w_8653 , \865_b0 , w_8655 );
not ( w_8655 , w_8677 );
and ( w_8677 , w_8676 , w_8654 );
or ( w_8654 , \867_b1 , w_8678 );
or ( w_8655 , \867_b0 , w_8657 );
not ( w_8657 , w_8679 );
and ( w_8679 , w_8678 , w_8656 );
or ( w_8656 , \869_b1 , w_8680 );
or ( w_8657 , \869_b0 , w_8659 );
not ( w_8659 , w_8681 );
and ( w_8681 , w_8680 , w_8658 );
or ( w_8658 , \871_b1 , w_8682 );
or ( w_8659 , \871_b0 , w_8661 );
not ( w_8661 , w_8683 );
and ( w_8683 , w_8682 , w_8660 );
or ( w_8660 , \873_b1 , w_8684 );
or ( w_8661 , \873_b0 , w_8663 );
not ( w_8663 , w_8685 );
and ( w_8685 , w_8684 , w_8662 );
buf ( w_8662 , \875_b1 );
not ( w_8662 , w_8686 );
not ( w_8663 , w_8687 );
and ( w_8686 , w_8687 , \875_b0 );
or ( \910_b1 , \877_b1 , w_8710 );
or ( \910_b0 , \877_b0 , w_8689 );
not ( w_8689 , w_8711 );
and ( w_8711 , w_8710 , w_8688 );
or ( w_8688 , \879_b1 , w_8712 );
or ( w_8689 , \879_b0 , w_8691 );
not ( w_8691 , w_8713 );
and ( w_8713 , w_8712 , w_8690 );
or ( w_8690 , \881_b1 , w_8714 );
or ( w_8691 , \881_b0 , w_8693 );
not ( w_8693 , w_8715 );
and ( w_8715 , w_8714 , w_8692 );
or ( w_8692 , \883_b1 , w_8716 );
or ( w_8693 , \883_b0 , w_8695 );
not ( w_8695 , w_8717 );
and ( w_8717 , w_8716 , w_8694 );
or ( w_8694 , \885_b1 , w_8718 );
or ( w_8695 , \885_b0 , w_8697 );
not ( w_8697 , w_8719 );
and ( w_8719 , w_8718 , w_8696 );
or ( w_8696 , \890_b1 , w_8720 );
or ( w_8697 , \890_b0 , w_8699 );
not ( w_8699 , w_8721 );
and ( w_8721 , w_8720 , w_8698 );
or ( w_8698 , \895_b1 , w_8722 );
or ( w_8699 , \895_b0 , w_8701 );
not ( w_8701 , w_8723 );
and ( w_8723 , w_8722 , w_8700 );
or ( w_8700 , \900_b1 , w_8724 );
or ( w_8701 , \900_b0 , w_8703 );
not ( w_8703 , w_8725 );
and ( w_8725 , w_8724 , w_8702 );
or ( w_8702 , \905_b1 , w_8726 );
or ( w_8703 , \905_b0 , w_8705 );
not ( w_8705 , w_8727 );
and ( w_8727 , w_8726 , w_8704 );
or ( w_8704 , \906_b1 , w_8728 );
or ( w_8705 , \906_b0 , w_8707 );
not ( w_8707 , w_8729 );
and ( w_8729 , w_8728 , w_8706 );
or ( w_8706 , \907_b1 , w_8730 );
or ( w_8707 , \907_b0 , w_8709 );
not ( w_8709 , w_8731 );
and ( w_8731 , w_8730 , w_8708 );
or ( w_8708 , \908_b1 , w_8732 );
or ( w_8709 , \908_b0 , \909_b0 );
not ( \909_b0 , w_8733 );
and ( w_8733 , w_8732 , \909_b1 );
or ( \952_b1 , \911_b1 , w_8756 );
or ( \952_b0 , \911_b0 , w_8735 );
not ( w_8735 , w_8757 );
and ( w_8757 , w_8756 , w_8734 );
or ( w_8734 , \913_b1 , w_8758 );
or ( w_8735 , \913_b0 , w_8737 );
not ( w_8737 , w_8759 );
and ( w_8759 , w_8758 , w_8736 );
or ( w_8736 , \915_b1 , w_8760 );
or ( w_8737 , \915_b0 , w_8739 );
not ( w_8739 , w_8761 );
and ( w_8761 , w_8760 , w_8738 );
or ( w_8738 , \917_b1 , w_8762 );
or ( w_8739 , \917_b0 , w_8741 );
not ( w_8741 , w_8763 );
and ( w_8763 , w_8762 , w_8740 );
or ( w_8740 , \919_b1 , w_8764 );
or ( w_8741 , \919_b0 , w_8743 );
not ( w_8743 , w_8765 );
and ( w_8765 , w_8764 , w_8742 );
or ( w_8742 , \926_b1 , w_8766 );
or ( w_8743 , \926_b0 , w_8745 );
not ( w_8745 , w_8767 );
and ( w_8767 , w_8766 , w_8744 );
or ( w_8744 , \933_b1 , w_8768 );
or ( w_8745 , \933_b0 , w_8747 );
not ( w_8747 , w_8769 );
and ( w_8769 , w_8768 , w_8746 );
or ( w_8746 , \940_b1 , w_8770 );
or ( w_8747 , \940_b0 , w_8749 );
not ( w_8749 , w_8771 );
and ( w_8771 , w_8770 , w_8748 );
or ( w_8748 , \947_b1 , w_8772 );
or ( w_8749 , \947_b0 , w_8751 );
not ( w_8751 , w_8773 );
and ( w_8773 , w_8772 , w_8750 );
or ( w_8750 , \948_b1 , w_8774 );
or ( w_8751 , \948_b0 , w_8753 );
not ( w_8753 , w_8775 );
and ( w_8775 , w_8774 , w_8752 );
or ( w_8752 , \949_b1 , w_8776 );
or ( w_8753 , \949_b0 , w_8755 );
not ( w_8755 , w_8777 );
and ( w_8777 , w_8776 , w_8754 );
or ( w_8754 , \950_b1 , w_8778 );
or ( w_8755 , \950_b0 , \951_b0 );
not ( \951_b0 , w_8779 );
and ( w_8779 , w_8778 , \951_b1 );
or ( \990_b1 , \987_b1 , w_8782 );
or ( \990_b0 , \987_b0 , w_8781 );
not ( w_8781 , w_8783 );
and ( w_8783 , w_8782 , w_8780 );
or ( w_8780 , \988_b1 , w_8784 );
or ( w_8781 , \988_b0 , \989_b0 );
not ( \989_b0 , w_8785 );
and ( w_8785 , w_8784 , \989_b1 );
or ( \1000_b1 , \997_b1 , w_8788 );
or ( \1000_b0 , \997_b0 , w_8787 );
not ( w_8787 , w_8789 );
and ( w_8789 , w_8788 , w_8786 );
or ( w_8786 , \998_b1 , w_8790 );
or ( w_8787 , \998_b0 , \999_b0 );
not ( \999_b0 , w_8791 );
and ( w_8791 , w_8790 , \999_b1 );
or ( \1008_b1 , \953_b1 , w_8814 );
or ( \1008_b0 , \953_b0 , w_8793 );
not ( w_8793 , w_8815 );
and ( w_8815 , w_8814 , w_8792 );
or ( w_8792 , \955_b1 , w_8816 );
or ( w_8793 , \955_b0 , w_8795 );
not ( w_8795 , w_8817 );
and ( w_8817 , w_8816 , w_8794 );
or ( w_8794 , \957_b1 , w_8818 );
or ( w_8795 , \957_b0 , w_8797 );
not ( w_8797 , w_8819 );
and ( w_8819 , w_8818 , w_8796 );
or ( w_8796 , \959_b1 , w_8820 );
or ( w_8797 , \959_b0 , w_8799 );
not ( w_8799 , w_8821 );
and ( w_8821 , w_8820 , w_8798 );
or ( w_8798 , \961_b1 , w_8822 );
or ( w_8799 , \961_b0 , w_8801 );
not ( w_8801 , w_8823 );
and ( w_8823 , w_8822 , w_8800 );
or ( w_8800 , \972_b1 , w_8824 );
or ( w_8801 , \972_b0 , w_8803 );
not ( w_8803 , w_8825 );
and ( w_8825 , w_8824 , w_8802 );
or ( w_8802 , \983_b1 , w_8826 );
or ( w_8803 , \983_b0 , w_8805 );
not ( w_8805 , w_8827 );
and ( w_8827 , w_8826 , w_8804 );
or ( w_8804 , \993_b1 , w_8828 );
or ( w_8805 , \993_b0 , w_8807 );
not ( w_8807 , w_8829 );
and ( w_8829 , w_8828 , w_8806 );
or ( w_8806 , \1003_b1 , w_8830 );
or ( w_8807 , \1003_b0 , w_8809 );
not ( w_8809 , w_8831 );
and ( w_8831 , w_8830 , w_8808 );
or ( w_8808 , \1004_b1 , w_8832 );
or ( w_8809 , \1004_b0 , w_8811 );
not ( w_8811 , w_8833 );
and ( w_8833 , w_8832 , w_8810 );
or ( w_8810 , \1005_b1 , w_8834 );
or ( w_8811 , \1005_b0 , w_8813 );
not ( w_8813 , w_8835 );
and ( w_8835 , w_8834 , w_8812 );
or ( w_8812 , \1006_b1 , w_8836 );
or ( w_8813 , \1006_b0 , \1007_b0 );
not ( \1007_b0 , w_8837 );
and ( w_8837 , w_8836 , \1007_b1 );
or ( \1058_b1 , \1055_b1 , w_8840 );
or ( \1058_b0 , \1055_b0 , w_8839 );
not ( w_8839 , w_8841 );
and ( w_8841 , w_8840 , w_8838 );
or ( w_8838 , \1056_b1 , w_8842 );
or ( w_8839 , \1056_b0 , \1057_b0 );
not ( \1057_b0 , w_8843 );
and ( w_8843 , w_8842 , \1057_b1 );
or ( \1068_b1 , \1065_b1 , w_8846 );
or ( \1068_b0 , \1065_b0 , w_8845 );
not ( w_8845 , w_8847 );
and ( w_8847 , w_8846 , w_8844 );
or ( w_8844 , \1066_b1 , w_8848 );
or ( w_8845 , \1066_b0 , \1067_b0 );
not ( \1067_b0 , w_8849 );
and ( w_8849 , w_8848 , \1067_b1 );
or ( \1076_b1 , \1009_b1 , w_8872 );
or ( \1076_b0 , \1009_b0 , w_8851 );
not ( w_8851 , w_8873 );
and ( w_8873 , w_8872 , w_8850 );
or ( w_8850 , \1011_b1 , w_8874 );
or ( w_8851 , \1011_b0 , w_8853 );
not ( w_8853 , w_8875 );
and ( w_8875 , w_8874 , w_8852 );
or ( w_8852 , \1013_b1 , w_8876 );
or ( w_8853 , \1013_b0 , w_8855 );
not ( w_8855 , w_8877 );
and ( w_8877 , w_8876 , w_8854 );
or ( w_8854 , \1015_b1 , w_8878 );
or ( w_8855 , \1015_b0 , w_8857 );
not ( w_8857 , w_8879 );
and ( w_8879 , w_8878 , w_8856 );
or ( w_8856 , \1017_b1 , w_8880 );
or ( w_8857 , \1017_b0 , w_8859 );
not ( w_8859 , w_8881 );
and ( w_8881 , w_8880 , w_8858 );
or ( w_8858 , \1034_b1 , w_8882 );
or ( w_8859 , \1034_b0 , w_8861 );
not ( w_8861 , w_8883 );
and ( w_8883 , w_8882 , w_8860 );
or ( w_8860 , \1051_b1 , w_8884 );
or ( w_8861 , \1051_b0 , w_8863 );
not ( w_8863 , w_8885 );
and ( w_8885 , w_8884 , w_8862 );
or ( w_8862 , \1061_b1 , w_8886 );
or ( w_8863 , \1061_b0 , w_8865 );
not ( w_8865 , w_8887 );
and ( w_8887 , w_8886 , w_8864 );
or ( w_8864 , \1071_b1 , w_8888 );
or ( w_8865 , \1071_b0 , w_8867 );
not ( w_8867 , w_8889 );
and ( w_8889 , w_8888 , w_8866 );
or ( w_8866 , \1072_b1 , w_8890 );
or ( w_8867 , \1072_b0 , w_8869 );
not ( w_8869 , w_8891 );
and ( w_8891 , w_8890 , w_8868 );
or ( w_8868 , \1073_b1 , w_8892 );
or ( w_8869 , \1073_b0 , w_8871 );
not ( w_8871 , w_8893 );
and ( w_8893 , w_8892 , w_8870 );
or ( w_8870 , \1074_b1 , w_8894 );
or ( w_8871 , \1074_b0 , \1075_b0 );
not ( \1075_b0 , w_8895 );
and ( w_8895 , w_8894 , \1075_b1 );
or ( \1138_b1 , \1135_b1 , w_8898 );
or ( \1138_b0 , \1135_b0 , w_8897 );
not ( w_8897 , w_8899 );
and ( w_8899 , w_8898 , w_8896 );
or ( w_8896 , \1136_b1 , w_8900 );
or ( w_8897 , \1136_b0 , \1137_b0 );
not ( \1137_b0 , w_8901 );
and ( w_8901 , w_8900 , \1137_b1 );
or ( \1148_b1 , \1145_b1 , w_8904 );
or ( \1148_b0 , \1145_b0 , w_8903 );
not ( w_8903 , w_8905 );
and ( w_8905 , w_8904 , w_8902 );
or ( w_8902 , \1146_b1 , w_8906 );
or ( w_8903 , \1146_b0 , \1147_b0 );
not ( \1147_b0 , w_8907 );
and ( w_8907 , w_8906 , \1147_b1 );
or ( \1156_b1 , \1077_b1 , w_8930 );
or ( \1156_b0 , \1077_b0 , w_8909 );
not ( w_8909 , w_8931 );
and ( w_8931 , w_8930 , w_8908 );
or ( w_8908 , \1079_b1 , w_8932 );
or ( w_8909 , \1079_b0 , w_8911 );
not ( w_8911 , w_8933 );
and ( w_8933 , w_8932 , w_8910 );
or ( w_8910 , \1081_b1 , w_8934 );
or ( w_8911 , \1081_b0 , w_8913 );
not ( w_8913 , w_8935 );
and ( w_8935 , w_8934 , w_8912 );
or ( w_8912 , \1083_b1 , w_8936 );
or ( w_8913 , \1083_b0 , w_8915 );
not ( w_8915 , w_8937 );
and ( w_8937 , w_8936 , w_8914 );
or ( w_8914 , \1085_b1 , w_8938 );
or ( w_8915 , \1085_b0 , w_8917 );
not ( w_8917 , w_8939 );
and ( w_8939 , w_8938 , w_8916 );
or ( w_8916 , \1108_b1 , w_8940 );
or ( w_8917 , \1108_b0 , w_8919 );
not ( w_8919 , w_8941 );
and ( w_8941 , w_8940 , w_8918 );
or ( w_8918 , \1131_b1 , w_8942 );
or ( w_8919 , \1131_b0 , w_8921 );
not ( w_8921 , w_8943 );
and ( w_8943 , w_8942 , w_8920 );
or ( w_8920 , \1141_b1 , w_8944 );
or ( w_8921 , \1141_b0 , w_8923 );
not ( w_8923 , w_8945 );
and ( w_8945 , w_8944 , w_8922 );
or ( w_8922 , \1151_b1 , w_8946 );
or ( w_8923 , \1151_b0 , w_8925 );
not ( w_8925 , w_8947 );
and ( w_8947 , w_8946 , w_8924 );
or ( w_8924 , \1152_b1 , w_8948 );
or ( w_8925 , \1152_b0 , w_8927 );
not ( w_8927 , w_8949 );
and ( w_8949 , w_8948 , w_8926 );
or ( w_8926 , \1153_b1 , w_8950 );
or ( w_8927 , \1153_b0 , w_8929 );
not ( w_8929 , w_8951 );
and ( w_8951 , w_8950 , w_8928 );
or ( w_8928 , \1154_b1 , w_8952 );
or ( w_8929 , \1154_b0 , \1155_b0 );
not ( \1155_b0 , w_8953 );
and ( w_8953 , w_8952 , \1155_b1 );
or ( \1230_b1 , \1227_b1 , w_8956 );
or ( \1230_b0 , \1227_b0 , w_8955 );
not ( w_8955 , w_8957 );
and ( w_8957 , w_8956 , w_8954 );
or ( w_8954 , \1228_b1 , w_8958 );
or ( w_8955 , \1228_b0 , \1229_b0 );
not ( \1229_b0 , w_8959 );
and ( w_8959 , w_8958 , \1229_b1 );
or ( \1240_b1 , \1237_b1 , w_8962 );
or ( \1240_b0 , \1237_b0 , w_8961 );
not ( w_8961 , w_8963 );
and ( w_8963 , w_8962 , w_8960 );
or ( w_8960 , \1238_b1 , w_8964 );
or ( w_8961 , \1238_b0 , \1239_b0 );
not ( \1239_b0 , w_8965 );
and ( w_8965 , w_8964 , \1239_b1 );
or ( \1248_b1 , \1157_b1 , w_8988 );
or ( \1248_b0 , \1157_b0 , w_8967 );
not ( w_8967 , w_8989 );
and ( w_8989 , w_8988 , w_8966 );
or ( w_8966 , \1159_b1 , w_8990 );
or ( w_8967 , \1159_b0 , w_8969 );
not ( w_8969 , w_8991 );
and ( w_8991 , w_8990 , w_8968 );
or ( w_8968 , \1161_b1 , w_8992 );
or ( w_8969 , \1161_b0 , w_8971 );
not ( w_8971 , w_8993 );
and ( w_8993 , w_8992 , w_8970 );
or ( w_8970 , \1163_b1 , w_8994 );
or ( w_8971 , \1163_b0 , w_8973 );
not ( w_8973 , w_8995 );
and ( w_8995 , w_8994 , w_8972 );
or ( w_8972 , \1165_b1 , w_8996 );
or ( w_8973 , \1165_b0 , w_8975 );
not ( w_8975 , w_8997 );
and ( w_8997 , w_8996 , w_8974 );
or ( w_8974 , \1194_b1 , w_8998 );
or ( w_8975 , \1194_b0 , w_8977 );
not ( w_8977 , w_8999 );
and ( w_8999 , w_8998 , w_8976 );
or ( w_8976 , \1223_b1 , w_9000 );
or ( w_8977 , \1223_b0 , w_8979 );
not ( w_8979 , w_9001 );
and ( w_9001 , w_9000 , w_8978 );
or ( w_8978 , \1233_b1 , w_9002 );
or ( w_8979 , \1233_b0 , w_8981 );
not ( w_8981 , w_9003 );
and ( w_9003 , w_9002 , w_8980 );
or ( w_8980 , \1243_b1 , w_9004 );
or ( w_8981 , \1243_b0 , w_8983 );
not ( w_8983 , w_9005 );
and ( w_9005 , w_9004 , w_8982 );
or ( w_8982 , \1244_b1 , w_9006 );
or ( w_8983 , \1244_b0 , w_8985 );
not ( w_8985 , w_9007 );
and ( w_9007 , w_9006 , w_8984 );
or ( w_8984 , \1245_b1 , w_9008 );
or ( w_8985 , \1245_b0 , w_8987 );
not ( w_8987 , w_9009 );
and ( w_9009 , w_9008 , w_8986 );
or ( w_8986 , \1246_b1 , w_9010 );
or ( w_8987 , \1246_b0 , \1247_b0 );
not ( \1247_b0 , w_9011 );
and ( w_9011 , w_9010 , \1247_b1 );
or ( \1334_b1 , \1331_b1 , w_9014 );
or ( \1334_b0 , \1331_b0 , w_9013 );
not ( w_9013 , w_9015 );
and ( w_9015 , w_9014 , w_9012 );
or ( w_9012 , \1332_b1 , w_9016 );
or ( w_9013 , \1332_b0 , \1333_b0 );
not ( \1333_b0 , w_9017 );
and ( w_9017 , w_9016 , \1333_b1 );
or ( \1344_b1 , \1341_b1 , w_9020 );
or ( \1344_b0 , \1341_b0 , w_9019 );
not ( w_9019 , w_9021 );
and ( w_9021 , w_9020 , w_9018 );
or ( w_9018 , \1342_b1 , w_9022 );
or ( w_9019 , \1342_b0 , \1343_b0 );
not ( \1343_b0 , w_9023 );
and ( w_9023 , w_9022 , \1343_b1 );
or ( \1352_b1 , \1249_b1 , w_9046 );
or ( \1352_b0 , \1249_b0 , w_9025 );
not ( w_9025 , w_9047 );
and ( w_9047 , w_9046 , w_9024 );
or ( w_9024 , \1251_b1 , w_9048 );
or ( w_9025 , \1251_b0 , w_9027 );
not ( w_9027 , w_9049 );
and ( w_9049 , w_9048 , w_9026 );
or ( w_9026 , \1253_b1 , w_9050 );
or ( w_9027 , \1253_b0 , w_9029 );
not ( w_9029 , w_9051 );
and ( w_9051 , w_9050 , w_9028 );
or ( w_9028 , \1255_b1 , w_9052 );
or ( w_9029 , \1255_b0 , w_9031 );
not ( w_9031 , w_9053 );
and ( w_9053 , w_9052 , w_9030 );
or ( w_9030 , \1257_b1 , w_9054 );
or ( w_9031 , \1257_b0 , w_9033 );
not ( w_9033 , w_9055 );
and ( w_9055 , w_9054 , w_9032 );
or ( w_9032 , \1292_b1 , w_9056 );
or ( w_9033 , \1292_b0 , w_9035 );
not ( w_9035 , w_9057 );
and ( w_9057 , w_9056 , w_9034 );
or ( w_9034 , \1327_b1 , w_9058 );
or ( w_9035 , \1327_b0 , w_9037 );
not ( w_9037 , w_9059 );
and ( w_9059 , w_9058 , w_9036 );
or ( w_9036 , \1337_b1 , w_9060 );
or ( w_9037 , \1337_b0 , w_9039 );
not ( w_9039 , w_9061 );
and ( w_9061 , w_9060 , w_9038 );
or ( w_9038 , \1347_b1 , w_9062 );
or ( w_9039 , \1347_b0 , w_9041 );
not ( w_9041 , w_9063 );
and ( w_9063 , w_9062 , w_9040 );
or ( w_9040 , \1348_b1 , w_9064 );
or ( w_9041 , \1348_b0 , w_9043 );
not ( w_9043 , w_9065 );
and ( w_9065 , w_9064 , w_9042 );
or ( w_9042 , \1349_b1 , w_9066 );
or ( w_9043 , \1349_b0 , w_9045 );
not ( w_9045 , w_9067 );
and ( w_9067 , w_9066 , w_9044 );
or ( w_9044 , \1350_b1 , w_9068 );
or ( w_9045 , \1350_b0 , \1351_b0 );
not ( \1351_b0 , w_9069 );
and ( w_9069 , w_9068 , \1351_b1 );
or ( \1450_b1 , \1447_b1 , w_9072 );
or ( \1450_b0 , \1447_b0 , w_9071 );
not ( w_9071 , w_9073 );
and ( w_9073 , w_9072 , w_9070 );
or ( w_9070 , \1448_b1 , w_9074 );
or ( w_9071 , \1448_b0 , \1449_b0 );
not ( \1449_b0 , w_9075 );
and ( w_9075 , w_9074 , \1449_b1 );
or ( \1460_b1 , \1457_b1 , w_9078 );
or ( \1460_b0 , \1457_b0 , w_9077 );
not ( w_9077 , w_9079 );
and ( w_9079 , w_9078 , w_9076 );
or ( w_9076 , \1458_b1 , w_9080 );
or ( w_9077 , \1458_b0 , \1459_b0 );
not ( \1459_b0 , w_9081 );
and ( w_9081 , w_9080 , \1459_b1 );
or ( \1468_b1 , \1353_b1 , w_9104 );
or ( \1468_b0 , \1353_b0 , w_9083 );
not ( w_9083 , w_9105 );
and ( w_9105 , w_9104 , w_9082 );
or ( w_9082 , \1355_b1 , w_9106 );
or ( w_9083 , \1355_b0 , w_9085 );
not ( w_9085 , w_9107 );
and ( w_9107 , w_9106 , w_9084 );
or ( w_9084 , \1357_b1 , w_9108 );
or ( w_9085 , \1357_b0 , w_9087 );
not ( w_9087 , w_9109 );
and ( w_9109 , w_9108 , w_9086 );
or ( w_9086 , \1359_b1 , w_9110 );
or ( w_9087 , \1359_b0 , w_9089 );
not ( w_9089 , w_9111 );
and ( w_9111 , w_9110 , w_9088 );
or ( w_9088 , \1361_b1 , w_9112 );
or ( w_9089 , \1361_b0 , w_9091 );
not ( w_9091 , w_9113 );
and ( w_9113 , w_9112 , w_9090 );
or ( w_9090 , \1402_b1 , w_9114 );
or ( w_9091 , \1402_b0 , w_9093 );
not ( w_9093 , w_9115 );
and ( w_9115 , w_9114 , w_9092 );
or ( w_9092 , \1443_b1 , w_9116 );
or ( w_9093 , \1443_b0 , w_9095 );
not ( w_9095 , w_9117 );
and ( w_9117 , w_9116 , w_9094 );
or ( w_9094 , \1453_b1 , w_9118 );
or ( w_9095 , \1453_b0 , w_9097 );
not ( w_9097 , w_9119 );
and ( w_9119 , w_9118 , w_9096 );
or ( w_9096 , \1463_b1 , w_9120 );
or ( w_9097 , \1463_b0 , w_9099 );
not ( w_9099 , w_9121 );
and ( w_9121 , w_9120 , w_9098 );
or ( w_9098 , \1464_b1 , w_9122 );
or ( w_9099 , \1464_b0 , w_9101 );
not ( w_9101 , w_9123 );
and ( w_9123 , w_9122 , w_9100 );
or ( w_9100 , \1465_b1 , w_9124 );
or ( w_9101 , \1465_b0 , w_9103 );
not ( w_9103 , w_9125 );
and ( w_9125 , w_9124 , w_9102 );
or ( w_9102 , \1466_b1 , w_9126 );
or ( w_9103 , \1466_b0 , \1467_b0 );
not ( \1467_b0 , w_9127 );
and ( w_9127 , w_9126 , \1467_b1 );
or ( \1578_b1 , \1575_b1 , w_9130 );
or ( \1578_b0 , \1575_b0 , w_9129 );
not ( w_9129 , w_9131 );
and ( w_9131 , w_9130 , w_9128 );
or ( w_9128 , \1576_b1 , w_9132 );
or ( w_9129 , \1576_b0 , \1577_b0 );
not ( \1577_b0 , w_9133 );
and ( w_9133 , w_9132 , \1577_b1 );
or ( \1588_b1 , \1585_b1 , w_9136 );
or ( \1588_b0 , \1585_b0 , w_9135 );
not ( w_9135 , w_9137 );
and ( w_9137 , w_9136 , w_9134 );
or ( w_9134 , \1586_b1 , w_9138 );
or ( w_9135 , \1586_b0 , \1587_b0 );
not ( \1587_b0 , w_9139 );
and ( w_9139 , w_9138 , \1587_b1 );
or ( \1596_b1 , \1469_b1 , w_9162 );
or ( \1596_b0 , \1469_b0 , w_9141 );
not ( w_9141 , w_9163 );
and ( w_9163 , w_9162 , w_9140 );
or ( w_9140 , \1471_b1 , w_9164 );
or ( w_9141 , \1471_b0 , w_9143 );
not ( w_9143 , w_9165 );
and ( w_9165 , w_9164 , w_9142 );
or ( w_9142 , \1473_b1 , w_9166 );
or ( w_9143 , \1473_b0 , w_9145 );
not ( w_9145 , w_9167 );
and ( w_9167 , w_9166 , w_9144 );
or ( w_9144 , \1475_b1 , w_9168 );
or ( w_9145 , \1475_b0 , w_9147 );
not ( w_9147 , w_9169 );
and ( w_9169 , w_9168 , w_9146 );
or ( w_9146 , \1477_b1 , w_9170 );
or ( w_9147 , \1477_b0 , w_9149 );
not ( w_9149 , w_9171 );
and ( w_9171 , w_9170 , w_9148 );
or ( w_9148 , \1524_b1 , w_9172 );
or ( w_9149 , \1524_b0 , w_9151 );
not ( w_9151 , w_9173 );
and ( w_9173 , w_9172 , w_9150 );
or ( w_9150 , \1571_b1 , w_9174 );
or ( w_9151 , \1571_b0 , w_9153 );
not ( w_9153 , w_9175 );
and ( w_9175 , w_9174 , w_9152 );
or ( w_9152 , \1581_b1 , w_9176 );
or ( w_9153 , \1581_b0 , w_9155 );
not ( w_9155 , w_9177 );
and ( w_9177 , w_9176 , w_9154 );
or ( w_9154 , \1591_b1 , w_9178 );
or ( w_9155 , \1591_b0 , w_9157 );
not ( w_9157 , w_9179 );
and ( w_9179 , w_9178 , w_9156 );
or ( w_9156 , \1592_b1 , w_9180 );
or ( w_9157 , \1592_b0 , w_9159 );
not ( w_9159 , w_9181 );
and ( w_9181 , w_9180 , w_9158 );
or ( w_9158 , \1593_b1 , w_9182 );
or ( w_9159 , \1593_b0 , w_9161 );
not ( w_9161 , w_9183 );
and ( w_9183 , w_9182 , w_9160 );
or ( w_9160 , \1594_b1 , w_9184 );
or ( w_9161 , \1594_b0 , \1595_b0 );
not ( \1595_b0 , w_9185 );
and ( w_9185 , w_9184 , \1595_b1 );
or ( \1718_b1 , \1715_b1 , w_9188 );
or ( \1718_b0 , \1715_b0 , w_9187 );
not ( w_9187 , w_9189 );
and ( w_9189 , w_9188 , w_9186 );
or ( w_9186 , \1716_b1 , w_9190 );
or ( w_9187 , \1716_b0 , \1717_b0 );
not ( \1717_b0 , w_9191 );
and ( w_9191 , w_9190 , \1717_b1 );
or ( \1728_b1 , \1725_b1 , w_9194 );
or ( \1728_b0 , \1725_b0 , w_9193 );
not ( w_9193 , w_9195 );
and ( w_9195 , w_9194 , w_9192 );
or ( w_9192 , \1726_b1 , w_9196 );
or ( w_9193 , \1726_b0 , \1727_b0 );
not ( \1727_b0 , w_9197 );
and ( w_9197 , w_9196 , \1727_b1 );
or ( \1736_b1 , \1597_b1 , w_9220 );
or ( \1736_b0 , \1597_b0 , w_9199 );
not ( w_9199 , w_9221 );
and ( w_9221 , w_9220 , w_9198 );
or ( w_9198 , \1599_b1 , w_9222 );
or ( w_9199 , \1599_b0 , w_9201 );
not ( w_9201 , w_9223 );
and ( w_9223 , w_9222 , w_9200 );
or ( w_9200 , \1601_b1 , w_9224 );
or ( w_9201 , \1601_b0 , w_9203 );
not ( w_9203 , w_9225 );
and ( w_9225 , w_9224 , w_9202 );
or ( w_9202 , \1603_b1 , w_9226 );
or ( w_9203 , \1603_b0 , w_9205 );
not ( w_9205 , w_9227 );
and ( w_9227 , w_9226 , w_9204 );
or ( w_9204 , \1605_b1 , w_9228 );
or ( w_9205 , \1605_b0 , w_9207 );
not ( w_9207 , w_9229 );
and ( w_9229 , w_9228 , w_9206 );
or ( w_9206 , \1658_b1 , w_9230 );
or ( w_9207 , \1658_b0 , w_9209 );
not ( w_9209 , w_9231 );
and ( w_9231 , w_9230 , w_9208 );
or ( w_9208 , \1711_b1 , w_9232 );
or ( w_9209 , \1711_b0 , w_9211 );
not ( w_9211 , w_9233 );
and ( w_9233 , w_9232 , w_9210 );
or ( w_9210 , \1721_b1 , w_9234 );
or ( w_9211 , \1721_b0 , w_9213 );
not ( w_9213 , w_9235 );
and ( w_9235 , w_9234 , w_9212 );
or ( w_9212 , \1731_b1 , w_9236 );
or ( w_9213 , \1731_b0 , w_9215 );
not ( w_9215 , w_9237 );
and ( w_9237 , w_9236 , w_9214 );
or ( w_9214 , \1732_b1 , w_9238 );
or ( w_9215 , \1732_b0 , w_9217 );
not ( w_9217 , w_9239 );
and ( w_9239 , w_9238 , w_9216 );
or ( w_9216 , \1733_b1 , w_9240 );
or ( w_9217 , \1733_b0 , w_9219 );
not ( w_9219 , w_9241 );
and ( w_9241 , w_9240 , w_9218 );
or ( w_9218 , \1734_b1 , w_9242 );
or ( w_9219 , \1734_b0 , \1735_b0 );
not ( \1735_b0 , w_9243 );
and ( w_9243 , w_9242 , \1735_b1 );
or ( \1870_b1 , \1867_b1 , w_9246 );
or ( \1870_b0 , \1867_b0 , w_9245 );
not ( w_9245 , w_9247 );
and ( w_9247 , w_9246 , w_9244 );
or ( w_9244 , \1868_b1 , w_9248 );
or ( w_9245 , \1868_b0 , \1869_b0 );
not ( \1869_b0 , w_9249 );
and ( w_9249 , w_9248 , \1869_b1 );
or ( \1880_b1 , \1877_b1 , w_9252 );
or ( \1880_b0 , \1877_b0 , w_9251 );
not ( w_9251 , w_9253 );
and ( w_9253 , w_9252 , w_9250 );
or ( w_9250 , \1878_b1 , w_9254 );
or ( w_9251 , \1878_b0 , \1879_b0 );
not ( \1879_b0 , w_9255 );
and ( w_9255 , w_9254 , \1879_b1 );
or ( \1888_b1 , \1737_b1 , w_9278 );
or ( \1888_b0 , \1737_b0 , w_9257 );
not ( w_9257 , w_9279 );
and ( w_9279 , w_9278 , w_9256 );
or ( w_9256 , \1739_b1 , w_9280 );
or ( w_9257 , \1739_b0 , w_9259 );
not ( w_9259 , w_9281 );
and ( w_9281 , w_9280 , w_9258 );
or ( w_9258 , \1741_b1 , w_9282 );
or ( w_9259 , \1741_b0 , w_9261 );
not ( w_9261 , w_9283 );
and ( w_9283 , w_9282 , w_9260 );
or ( w_9260 , \1743_b1 , w_9284 );
or ( w_9261 , \1743_b0 , w_9263 );
not ( w_9263 , w_9285 );
and ( w_9285 , w_9284 , w_9262 );
or ( w_9262 , \1745_b1 , w_9286 );
or ( w_9263 , \1745_b0 , w_9265 );
not ( w_9265 , w_9287 );
and ( w_9287 , w_9286 , w_9264 );
or ( w_9264 , \1804_b1 , w_9288 );
or ( w_9265 , \1804_b0 , w_9267 );
not ( w_9267 , w_9289 );
and ( w_9289 , w_9288 , w_9266 );
or ( w_9266 , \1863_b1 , w_9290 );
or ( w_9267 , \1863_b0 , w_9269 );
not ( w_9269 , w_9291 );
and ( w_9291 , w_9290 , w_9268 );
or ( w_9268 , \1873_b1 , w_9292 );
or ( w_9269 , \1873_b0 , w_9271 );
not ( w_9271 , w_9293 );
and ( w_9293 , w_9292 , w_9270 );
or ( w_9270 , \1883_b1 , w_9294 );
or ( w_9271 , \1883_b0 , w_9273 );
not ( w_9273 , w_9295 );
and ( w_9295 , w_9294 , w_9272 );
or ( w_9272 , \1884_b1 , w_9296 );
or ( w_9273 , \1884_b0 , w_9275 );
not ( w_9275 , w_9297 );
and ( w_9297 , w_9296 , w_9274 );
or ( w_9274 , \1885_b1 , w_9298 );
or ( w_9275 , \1885_b0 , w_9277 );
not ( w_9277 , w_9299 );
and ( w_9299 , w_9298 , w_9276 );
or ( w_9276 , \1886_b1 , w_9300 );
or ( w_9277 , \1886_b0 , \1887_b0 );
not ( \1887_b0 , w_9301 );
and ( w_9301 , w_9300 , \1887_b1 );
or ( \2034_b1 , \2031_b1 , w_9304 );
or ( \2034_b0 , \2031_b0 , w_9303 );
not ( w_9303 , w_9305 );
and ( w_9305 , w_9304 , w_9302 );
or ( w_9302 , \2032_b1 , w_9306 );
or ( w_9303 , \2032_b0 , \2033_b0 );
not ( \2033_b0 , w_9307 );
and ( w_9307 , w_9306 , \2033_b1 );
or ( \2044_b1 , \2041_b1 , w_9310 );
or ( \2044_b0 , \2041_b0 , w_9309 );
not ( w_9309 , w_9311 );
and ( w_9311 , w_9310 , w_9308 );
or ( w_9308 , \2042_b1 , w_9312 );
or ( w_9309 , \2042_b0 , \2043_b0 );
not ( \2043_b0 , w_9313 );
and ( w_9313 , w_9312 , \2043_b1 );
or ( \2052_b1 , \1889_b1 , w_9336 );
or ( \2052_b0 , \1889_b0 , w_9315 );
not ( w_9315 , w_9337 );
and ( w_9337 , w_9336 , w_9314 );
or ( w_9314 , \1891_b1 , w_9338 );
or ( w_9315 , \1891_b0 , w_9317 );
not ( w_9317 , w_9339 );
and ( w_9339 , w_9338 , w_9316 );
or ( w_9316 , \1893_b1 , w_9340 );
or ( w_9317 , \1893_b0 , w_9319 );
not ( w_9319 , w_9341 );
and ( w_9341 , w_9340 , w_9318 );
or ( w_9318 , \1895_b1 , w_9342 );
or ( w_9319 , \1895_b0 , w_9321 );
not ( w_9321 , w_9343 );
and ( w_9343 , w_9342 , w_9320 );
or ( w_9320 , \1897_b1 , w_9344 );
or ( w_9321 , \1897_b0 , w_9323 );
not ( w_9323 , w_9345 );
and ( w_9345 , w_9344 , w_9322 );
or ( w_9322 , \1962_b1 , w_9346 );
or ( w_9323 , \1962_b0 , w_9325 );
not ( w_9325 , w_9347 );
and ( w_9347 , w_9346 , w_9324 );
or ( w_9324 , \2027_b1 , w_9348 );
or ( w_9325 , \2027_b0 , w_9327 );
not ( w_9327 , w_9349 );
and ( w_9349 , w_9348 , w_9326 );
or ( w_9326 , \2037_b1 , w_9350 );
or ( w_9327 , \2037_b0 , w_9329 );
not ( w_9329 , w_9351 );
and ( w_9351 , w_9350 , w_9328 );
or ( w_9328 , \2047_b1 , w_9352 );
or ( w_9329 , \2047_b0 , w_9331 );
not ( w_9331 , w_9353 );
and ( w_9353 , w_9352 , w_9330 );
or ( w_9330 , \2048_b1 , w_9354 );
or ( w_9331 , \2048_b0 , w_9333 );
not ( w_9333 , w_9355 );
and ( w_9355 , w_9354 , w_9332 );
or ( w_9332 , \2049_b1 , w_9356 );
or ( w_9333 , \2049_b0 , w_9335 );
not ( w_9335 , w_9357 );
and ( w_9357 , w_9356 , w_9334 );
or ( w_9334 , \2050_b1 , w_9358 );
or ( w_9335 , \2050_b0 , \2051_b0 );
not ( \2051_b0 , w_9359 );
and ( w_9359 , w_9358 , \2051_b1 );
or ( \2210_b1 , \2207_b1 , w_9362 );
or ( \2210_b0 , \2207_b0 , w_9361 );
not ( w_9361 , w_9363 );
and ( w_9363 , w_9362 , w_9360 );
or ( w_9360 , \2208_b1 , w_9364 );
or ( w_9361 , \2208_b0 , \2209_b0 );
not ( \2209_b0 , w_9365 );
and ( w_9365 , w_9364 , \2209_b1 );
or ( \2220_b1 , \2217_b1 , w_9368 );
or ( \2220_b0 , \2217_b0 , w_9367 );
not ( w_9367 , w_9369 );
and ( w_9369 , w_9368 , w_9366 );
or ( w_9366 , \2218_b1 , w_9370 );
or ( w_9367 , \2218_b0 , \2219_b0 );
not ( \2219_b0 , w_9371 );
and ( w_9371 , w_9370 , \2219_b1 );
or ( \2228_b1 , \2053_b1 , w_9394 );
or ( \2228_b0 , \2053_b0 , w_9373 );
not ( w_9373 , w_9395 );
and ( w_9395 , w_9394 , w_9372 );
or ( w_9372 , \2055_b1 , w_9396 );
or ( w_9373 , \2055_b0 , w_9375 );
not ( w_9375 , w_9397 );
and ( w_9397 , w_9396 , w_9374 );
or ( w_9374 , \2057_b1 , w_9398 );
or ( w_9375 , \2057_b0 , w_9377 );
not ( w_9377 , w_9399 );
and ( w_9399 , w_9398 , w_9376 );
or ( w_9376 , \2059_b1 , w_9400 );
or ( w_9377 , \2059_b0 , w_9379 );
not ( w_9379 , w_9401 );
and ( w_9401 , w_9400 , w_9378 );
or ( w_9378 , \2061_b1 , w_9402 );
or ( w_9379 , \2061_b0 , w_9381 );
not ( w_9381 , w_9403 );
and ( w_9403 , w_9402 , w_9380 );
or ( w_9380 , \2132_b1 , w_9404 );
or ( w_9381 , \2132_b0 , w_9383 );
not ( w_9383 , w_9405 );
and ( w_9405 , w_9404 , w_9382 );
or ( w_9382 , \2203_b1 , w_9406 );
or ( w_9383 , \2203_b0 , w_9385 );
not ( w_9385 , w_9407 );
and ( w_9407 , w_9406 , w_9384 );
or ( w_9384 , \2213_b1 , w_9408 );
or ( w_9385 , \2213_b0 , w_9387 );
not ( w_9387 , w_9409 );
and ( w_9409 , w_9408 , w_9386 );
or ( w_9386 , \2223_b1 , w_9410 );
or ( w_9387 , \2223_b0 , w_9389 );
not ( w_9389 , w_9411 );
and ( w_9411 , w_9410 , w_9388 );
or ( w_9388 , \2224_b1 , w_9412 );
or ( w_9389 , \2224_b0 , w_9391 );
not ( w_9391 , w_9413 );
and ( w_9413 , w_9412 , w_9390 );
or ( w_9390 , \2225_b1 , w_9414 );
or ( w_9391 , \2225_b0 , w_9393 );
not ( w_9393 , w_9415 );
and ( w_9415 , w_9414 , w_9392 );
or ( w_9392 , \2226_b1 , w_9416 );
or ( w_9393 , \2226_b0 , \2227_b0 );
not ( \2227_b0 , w_9417 );
and ( w_9417 , w_9416 , \2227_b1 );
or ( \2398_b1 , \2395_b1 , w_9420 );
or ( \2398_b0 , \2395_b0 , w_9419 );
not ( w_9419 , w_9421 );
and ( w_9421 , w_9420 , w_9418 );
or ( w_9418 , \2396_b1 , w_9422 );
or ( w_9419 , \2396_b0 , \2397_b0 );
not ( \2397_b0 , w_9423 );
and ( w_9423 , w_9422 , \2397_b1 );
or ( \2408_b1 , \2405_b1 , w_9426 );
or ( \2408_b0 , \2405_b0 , w_9425 );
not ( w_9425 , w_9427 );
and ( w_9427 , w_9426 , w_9424 );
or ( w_9424 , \2406_b1 , w_9428 );
or ( w_9425 , \2406_b0 , \2407_b0 );
not ( \2407_b0 , w_9429 );
and ( w_9429 , w_9428 , \2407_b1 );
or ( \2416_b1 , \2229_b1 , w_9452 );
or ( \2416_b0 , \2229_b0 , w_9431 );
not ( w_9431 , w_9453 );
and ( w_9453 , w_9452 , w_9430 );
or ( w_9430 , \2231_b1 , w_9454 );
or ( w_9431 , \2231_b0 , w_9433 );
not ( w_9433 , w_9455 );
and ( w_9455 , w_9454 , w_9432 );
or ( w_9432 , \2233_b1 , w_9456 );
or ( w_9433 , \2233_b0 , w_9435 );
not ( w_9435 , w_9457 );
and ( w_9457 , w_9456 , w_9434 );
or ( w_9434 , \2235_b1 , w_9458 );
or ( w_9435 , \2235_b0 , w_9437 );
not ( w_9437 , w_9459 );
and ( w_9459 , w_9458 , w_9436 );
or ( w_9436 , \2237_b1 , w_9460 );
or ( w_9437 , \2237_b0 , w_9439 );
not ( w_9439 , w_9461 );
and ( w_9461 , w_9460 , w_9438 );
or ( w_9438 , \2314_b1 , w_9462 );
or ( w_9439 , \2314_b0 , w_9441 );
not ( w_9441 , w_9463 );
and ( w_9463 , w_9462 , w_9440 );
or ( w_9440 , \2391_b1 , w_9464 );
or ( w_9441 , \2391_b0 , w_9443 );
not ( w_9443 , w_9465 );
and ( w_9465 , w_9464 , w_9442 );
or ( w_9442 , \2401_b1 , w_9466 );
or ( w_9443 , \2401_b0 , w_9445 );
not ( w_9445 , w_9467 );
and ( w_9467 , w_9466 , w_9444 );
or ( w_9444 , \2411_b1 , w_9468 );
or ( w_9445 , \2411_b0 , w_9447 );
not ( w_9447 , w_9469 );
and ( w_9469 , w_9468 , w_9446 );
or ( w_9446 , \2412_b1 , w_9470 );
or ( w_9447 , \2412_b0 , w_9449 );
not ( w_9449 , w_9471 );
and ( w_9471 , w_9470 , w_9448 );
or ( w_9448 , \2413_b1 , w_9472 );
or ( w_9449 , \2413_b0 , w_9451 );
not ( w_9451 , w_9473 );
and ( w_9473 , w_9472 , w_9450 );
or ( w_9450 , \2414_b1 , w_9474 );
or ( w_9451 , \2414_b0 , \2415_b0 );
not ( \2415_b0 , w_9475 );
and ( w_9475 , w_9474 , \2415_b1 );
or ( \2598_b1 , \2595_b1 , w_9478 );
or ( \2598_b0 , \2595_b0 , w_9477 );
not ( w_9477 , w_9479 );
and ( w_9479 , w_9478 , w_9476 );
or ( w_9476 , \2596_b1 , w_9480 );
or ( w_9477 , \2596_b0 , \2597_b0 );
not ( \2597_b0 , w_9481 );
and ( w_9481 , w_9480 , \2597_b1 );
or ( \2608_b1 , \2605_b1 , w_9484 );
or ( \2608_b0 , \2605_b0 , w_9483 );
not ( w_9483 , w_9485 );
and ( w_9485 , w_9484 , w_9482 );
or ( w_9482 , \2606_b1 , w_9486 );
or ( w_9483 , \2606_b0 , \2607_b0 );
not ( \2607_b0 , w_9487 );
and ( w_9487 , w_9486 , \2607_b1 );
or ( \2616_b1 , \2417_b1 , w_9510 );
or ( \2616_b0 , \2417_b0 , w_9489 );
not ( w_9489 , w_9511 );
and ( w_9511 , w_9510 , w_9488 );
or ( w_9488 , \2419_b1 , w_9512 );
or ( w_9489 , \2419_b0 , w_9491 );
not ( w_9491 , w_9513 );
and ( w_9513 , w_9512 , w_9490 );
or ( w_9490 , \2421_b1 , w_9514 );
or ( w_9491 , \2421_b0 , w_9493 );
not ( w_9493 , w_9515 );
and ( w_9515 , w_9514 , w_9492 );
or ( w_9492 , \2423_b1 , w_9516 );
or ( w_9493 , \2423_b0 , w_9495 );
not ( w_9495 , w_9517 );
and ( w_9517 , w_9516 , w_9494 );
or ( w_9494 , \2425_b1 , w_9518 );
or ( w_9495 , \2425_b0 , w_9497 );
not ( w_9497 , w_9519 );
and ( w_9519 , w_9518 , w_9496 );
or ( w_9496 , \2508_b1 , w_9520 );
or ( w_9497 , \2508_b0 , w_9499 );
not ( w_9499 , w_9521 );
and ( w_9521 , w_9520 , w_9498 );
or ( w_9498 , \2591_b1 , w_9522 );
or ( w_9499 , \2591_b0 , w_9501 );
not ( w_9501 , w_9523 );
and ( w_9523 , w_9522 , w_9500 );
or ( w_9500 , \2601_b1 , w_9524 );
or ( w_9501 , \2601_b0 , w_9503 );
not ( w_9503 , w_9525 );
and ( w_9525 , w_9524 , w_9502 );
or ( w_9502 , \2611_b1 , w_9526 );
or ( w_9503 , \2611_b0 , w_9505 );
not ( w_9505 , w_9527 );
and ( w_9527 , w_9526 , w_9504 );
or ( w_9504 , \2612_b1 , w_9528 );
or ( w_9505 , \2612_b0 , w_9507 );
not ( w_9507 , w_9529 );
and ( w_9529 , w_9528 , w_9506 );
or ( w_9506 , \2613_b1 , w_9530 );
or ( w_9507 , \2613_b0 , w_9509 );
not ( w_9509 , w_9531 );
and ( w_9531 , w_9530 , w_9508 );
or ( w_9508 , \2614_b1 , w_9532 );
or ( w_9509 , \2614_b0 , \2615_b0 );
not ( \2615_b0 , w_9533 );
and ( w_9533 , w_9532 , \2615_b1 );
or ( \2810_b1 , \2807_b1 , w_9536 );
or ( \2810_b0 , \2807_b0 , w_9535 );
not ( w_9535 , w_9537 );
and ( w_9537 , w_9536 , w_9534 );
or ( w_9534 , \2808_b1 , w_9538 );
or ( w_9535 , \2808_b0 , \2809_b0 );
not ( \2809_b0 , w_9539 );
and ( w_9539 , w_9538 , \2809_b1 );
or ( \2820_b1 , \2817_b1 , w_9542 );
or ( \2820_b0 , \2817_b0 , w_9541 );
not ( w_9541 , w_9543 );
and ( w_9543 , w_9542 , w_9540 );
or ( w_9540 , \2818_b1 , w_9544 );
or ( w_9541 , \2818_b0 , \2819_b0 );
not ( \2819_b0 , w_9545 );
and ( w_9545 , w_9544 , \2819_b1 );
or ( \2828_b1 , \2617_b1 , w_9568 );
or ( \2828_b0 , \2617_b0 , w_9547 );
not ( w_9547 , w_9569 );
and ( w_9569 , w_9568 , w_9546 );
or ( w_9546 , \2619_b1 , w_9570 );
or ( w_9547 , \2619_b0 , w_9549 );
not ( w_9549 , w_9571 );
and ( w_9571 , w_9570 , w_9548 );
or ( w_9548 , \2621_b1 , w_9572 );
or ( w_9549 , \2621_b0 , w_9551 );
not ( w_9551 , w_9573 );
and ( w_9573 , w_9572 , w_9550 );
or ( w_9550 , \2623_b1 , w_9574 );
or ( w_9551 , \2623_b0 , w_9553 );
not ( w_9553 , w_9575 );
and ( w_9575 , w_9574 , w_9552 );
or ( w_9552 , \2625_b1 , w_9576 );
or ( w_9553 , \2625_b0 , w_9555 );
not ( w_9555 , w_9577 );
and ( w_9577 , w_9576 , w_9554 );
or ( w_9554 , \2714_b1 , w_9578 );
or ( w_9555 , \2714_b0 , w_9557 );
not ( w_9557 , w_9579 );
and ( w_9579 , w_9578 , w_9556 );
or ( w_9556 , \2803_b1 , w_9580 );
or ( w_9557 , \2803_b0 , w_9559 );
not ( w_9559 , w_9581 );
and ( w_9581 , w_9580 , w_9558 );
or ( w_9558 , \2813_b1 , w_9582 );
or ( w_9559 , \2813_b0 , w_9561 );
not ( w_9561 , w_9583 );
and ( w_9583 , w_9582 , w_9560 );
or ( w_9560 , \2823_b1 , w_9584 );
or ( w_9561 , \2823_b0 , w_9563 );
not ( w_9563 , w_9585 );
and ( w_9585 , w_9584 , w_9562 );
or ( w_9562 , \2824_b1 , w_9586 );
or ( w_9563 , \2824_b0 , w_9565 );
not ( w_9565 , w_9587 );
and ( w_9587 , w_9586 , w_9564 );
or ( w_9564 , \2825_b1 , w_9588 );
or ( w_9565 , \2825_b0 , w_9567 );
not ( w_9567 , w_9589 );
and ( w_9589 , w_9588 , w_9566 );
or ( w_9566 , \2826_b1 , w_9590 );
or ( w_9567 , \2826_b0 , \2827_b0 );
not ( \2827_b0 , w_9591 );
and ( w_9591 , w_9590 , \2827_b1 );
or ( \2879_b1 , \2873_b1 , w_9594 );
or ( \2879_b0 , \2873_b0 , w_9593 );
not ( w_9593 , w_9595 );
and ( w_9595 , w_9594 , w_9592 );
or ( w_9592 , \2877_b1 , w_9596 );
or ( w_9593 , \2877_b0 , \2878_b0 );
not ( \2878_b0 , w_9597 );
and ( w_9597 , w_9596 , \2878_b1 );
or ( \2882_b1 , \2870_b1 , w_9600 );
or ( \2882_b0 , \2870_b0 , w_9599 );
not ( w_9599 , w_9601 );
and ( w_9601 , w_9600 , w_9598 );
or ( w_9598 , \2880_b1 , w_9602 );
or ( w_9599 , \2880_b0 , \2881_b0 );
not ( \2881_b0 , w_9603 );
and ( w_9603 , w_9602 , \2881_b1 );
or ( \2885_b1 , \2867_b1 , w_9606 );
or ( \2885_b0 , \2867_b0 , w_9605 );
not ( w_9605 , w_9607 );
and ( w_9607 , w_9606 , w_9604 );
or ( w_9604 , \2883_b1 , w_9608 );
or ( w_9605 , \2883_b0 , \2884_b0 );
not ( \2884_b0 , w_9609 );
and ( w_9609 , w_9608 , \2884_b1 );
or ( \2888_b1 , \2864_b1 , w_9612 );
or ( \2888_b0 , \2864_b0 , w_9611 );
not ( w_9611 , w_9613 );
and ( w_9613 , w_9612 , w_9610 );
or ( w_9610 , \2886_b1 , w_9614 );
or ( w_9611 , \2886_b0 , \2887_b0 );
not ( \2887_b0 , w_9615 );
and ( w_9615 , w_9614 , \2887_b1 );
or ( \2891_b1 , \2861_b1 , w_9618 );
or ( \2891_b0 , \2861_b0 , w_9617 );
not ( w_9617 , w_9619 );
and ( w_9619 , w_9618 , w_9616 );
or ( w_9616 , \2889_b1 , w_9620 );
or ( w_9617 , \2889_b0 , \2890_b0 );
not ( \2890_b0 , w_9621 );
and ( w_9621 , w_9620 , \2890_b1 );
or ( \2894_b1 , \2858_b1 , w_9624 );
or ( \2894_b0 , \2858_b0 , w_9623 );
not ( w_9623 , w_9625 );
and ( w_9625 , w_9624 , w_9622 );
or ( w_9622 , \2892_b1 , w_9626 );
or ( w_9623 , \2892_b0 , \2893_b0 );
not ( \2893_b0 , w_9627 );
and ( w_9627 , w_9626 , \2893_b1 );
or ( \2897_b1 , \2855_b1 , w_9630 );
or ( \2897_b0 , \2855_b0 , w_9629 );
not ( w_9629 , w_9631 );
and ( w_9631 , w_9630 , w_9628 );
or ( w_9628 , \2895_b1 , w_9632 );
or ( w_9629 , \2895_b0 , \2896_b0 );
not ( \2896_b0 , w_9633 );
and ( w_9633 , w_9632 , \2896_b1 );
or ( \2900_b1 , \2852_b1 , w_9636 );
or ( \2900_b0 , \2852_b0 , w_9635 );
not ( w_9635 , w_9637 );
and ( w_9637 , w_9636 , w_9634 );
or ( w_9634 , \2898_b1 , w_9638 );
or ( w_9635 , \2898_b0 , \2899_b0 );
not ( \2899_b0 , w_9639 );
and ( w_9639 , w_9638 , \2899_b1 );
or ( \2903_b1 , \2849_b1 , w_9642 );
or ( \2903_b0 , \2849_b0 , w_9641 );
not ( w_9641 , w_9643 );
and ( w_9643 , w_9642 , w_9640 );
or ( w_9640 , \2901_b1 , w_9644 );
or ( w_9641 , \2901_b0 , \2902_b0 );
not ( \2902_b0 , w_9645 );
and ( w_9645 , w_9644 , \2902_b1 );
or ( \2906_b1 , \2846_b1 , w_9648 );
or ( \2906_b0 , \2846_b0 , w_9647 );
not ( w_9647 , w_9649 );
and ( w_9649 , w_9648 , w_9646 );
or ( w_9646 , \2904_b1 , w_9650 );
or ( w_9647 , \2904_b0 , \2905_b0 );
not ( \2905_b0 , w_9651 );
and ( w_9651 , w_9650 , \2905_b1 );
or ( \2909_b1 , \2843_b1 , w_9654 );
or ( \2909_b0 , \2843_b0 , w_9653 );
not ( w_9653 , w_9655 );
and ( w_9655 , w_9654 , w_9652 );
or ( w_9652 , \2907_b1 , w_9656 );
or ( w_9653 , \2907_b0 , \2908_b0 );
not ( \2908_b0 , w_9657 );
and ( w_9657 , w_9656 , \2908_b1 );
or ( \2912_b1 , \2840_b1 , w_9660 );
or ( \2912_b0 , \2840_b0 , w_9659 );
not ( w_9659 , w_9661 );
and ( w_9661 , w_9660 , w_9658 );
or ( w_9658 , \2910_b1 , w_9662 );
or ( w_9659 , \2910_b0 , \2911_b0 );
not ( \2911_b0 , w_9663 );
and ( w_9663 , w_9662 , \2911_b1 );
or ( \2915_b1 , \2837_b1 , w_9666 );
or ( \2915_b0 , \2837_b0 , w_9665 );
not ( w_9665 , w_9667 );
and ( w_9667 , w_9666 , w_9664 );
or ( w_9664 , \2913_b1 , w_9668 );
or ( w_9665 , \2913_b0 , \2914_b0 );
not ( \2914_b0 , w_9669 );
and ( w_9669 , w_9668 , \2914_b1 );
or ( \2918_b1 , \2834_b1 , w_9672 );
or ( \2918_b0 , \2834_b0 , w_9671 );
not ( w_9671 , w_9673 );
and ( w_9673 , w_9672 , w_9670 );
or ( w_9670 , \2916_b1 , w_9674 );
or ( w_9671 , \2916_b0 , \2917_b0 );
not ( \2917_b0 , w_9675 );
and ( w_9675 , w_9674 , \2917_b1 );
or ( \2921_b1 , \2831_b1 , w_9678 );
or ( \2921_b0 , \2831_b0 , w_9677 );
not ( w_9677 , w_9679 );
and ( w_9679 , w_9678 , w_9676 );
or ( w_9676 , \2919_b1 , w_9680 );
or ( w_9677 , \2919_b0 , \2920_b0 );
not ( \2920_b0 , w_9681 );
and ( w_9681 , w_9680 , \2920_b1 );
endmodule

