// ...
module top(\a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,
		\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,
		\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,
		\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,\a[0]_b1 ,\a[0]_b0 ,\b[15]_b1 ,\b[15]_b0 ,\b[14]_b1 ,\b[14]_b0 ,
		\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,\b[10]_b0 ,\b[9]_b1 ,
		\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,\b[5]_b1 ,\b[5]_b0 ,
		\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,\b[1]_b0 ,\b[0]_b1 ,
		\b[0]_b0 ,\c[15]_b1 ,\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,
		\c[11]_b1 ,\c[11]_b0 ,\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,
		\c[7]_b0 ,\c[6]_b1 ,\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,
		\c[2]_b1 ,\c[2]_b0 ,\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,
		\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,
		\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,
		\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,
		\d[0]_b1 ,\d[0]_b0 ,\o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,
		\o[28]_b0 ,\o[27]_b1 ,\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,
		\o[23]_b1 ,\o[23]_b0 ,\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,
		\o[19]_b0 ,\o[18]_b1 ,\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,
		\o[14]_b1 ,\o[14]_b0 ,\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,
		\o[10]_b0 ,\o[9]_b1 ,\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,
		\o[5]_b1 ,\o[5]_b0 ,\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,
		\o[1]_b0 ,\o[0]_b1 ,\o[0]_b0 );
input \a[15]_b1 ,\a[15]_b0 ,\a[14]_b1 ,\a[14]_b0 ,\a[13]_b1 ,\a[13]_b0 ,\a[12]_b1 ,\a[12]_b0 ,\a[11]_b1 ,
		\a[11]_b0 ,\a[10]_b1 ,\a[10]_b0 ,\a[9]_b1 ,\a[9]_b0 ,\a[8]_b1 ,\a[8]_b0 ,\a[7]_b1 ,\a[7]_b0 ,
		\a[6]_b1 ,\a[6]_b0 ,\a[5]_b1 ,\a[5]_b0 ,\a[4]_b1 ,\a[4]_b0 ,\a[3]_b1 ,\a[3]_b0 ,\a[2]_b1 ,
		\a[2]_b0 ,\a[1]_b1 ,\a[1]_b0 ,\a[0]_b1 ,\a[0]_b0 ,\b[15]_b1 ,\b[15]_b0 ,\b[14]_b1 ,\b[14]_b0 ,
		\b[13]_b1 ,\b[13]_b0 ,\b[12]_b1 ,\b[12]_b0 ,\b[11]_b1 ,\b[11]_b0 ,\b[10]_b1 ,\b[10]_b0 ,\b[9]_b1 ,
		\b[9]_b0 ,\b[8]_b1 ,\b[8]_b0 ,\b[7]_b1 ,\b[7]_b0 ,\b[6]_b1 ,\b[6]_b0 ,\b[5]_b1 ,\b[5]_b0 ,
		\b[4]_b1 ,\b[4]_b0 ,\b[3]_b1 ,\b[3]_b0 ,\b[2]_b1 ,\b[2]_b0 ,\b[1]_b1 ,\b[1]_b0 ,\b[0]_b1 ,
		\b[0]_b0 ,\c[15]_b1 ,\c[15]_b0 ,\c[14]_b1 ,\c[14]_b0 ,\c[13]_b1 ,\c[13]_b0 ,\c[12]_b1 ,\c[12]_b0 ,
		\c[11]_b1 ,\c[11]_b0 ,\c[10]_b1 ,\c[10]_b0 ,\c[9]_b1 ,\c[9]_b0 ,\c[8]_b1 ,\c[8]_b0 ,\c[7]_b1 ,
		\c[7]_b0 ,\c[6]_b1 ,\c[6]_b0 ,\c[5]_b1 ,\c[5]_b0 ,\c[4]_b1 ,\c[4]_b0 ,\c[3]_b1 ,\c[3]_b0 ,
		\c[2]_b1 ,\c[2]_b0 ,\c[1]_b1 ,\c[1]_b0 ,\c[0]_b1 ,\c[0]_b0 ,\d[15]_b1 ,\d[15]_b0 ,\d[14]_b1 ,
		\d[14]_b0 ,\d[13]_b1 ,\d[13]_b0 ,\d[12]_b1 ,\d[12]_b0 ,\d[11]_b1 ,\d[11]_b0 ,\d[10]_b1 ,\d[10]_b0 ,
		\d[9]_b1 ,\d[9]_b0 ,\d[8]_b1 ,\d[8]_b0 ,\d[7]_b1 ,\d[7]_b0 ,\d[6]_b1 ,\d[6]_b0 ,\d[5]_b1 ,
		\d[5]_b0 ,\d[4]_b1 ,\d[4]_b0 ,\d[3]_b1 ,\d[3]_b0 ,\d[2]_b1 ,\d[2]_b0 ,\d[1]_b1 ,\d[1]_b0 ,
		\d[0]_b1 ,\d[0]_b0 ;
output \o[31]_b1 ,\o[31]_b0 ,\o[30]_b1 ,\o[30]_b0 ,\o[29]_b1 ,\o[29]_b0 ,\o[28]_b1 ,\o[28]_b0 ,\o[27]_b1 ,
		\o[27]_b0 ,\o[26]_b1 ,\o[26]_b0 ,\o[25]_b1 ,\o[25]_b0 ,\o[24]_b1 ,\o[24]_b0 ,\o[23]_b1 ,\o[23]_b0 ,
		\o[22]_b1 ,\o[22]_b0 ,\o[21]_b1 ,\o[21]_b0 ,\o[20]_b1 ,\o[20]_b0 ,\o[19]_b1 ,\o[19]_b0 ,\o[18]_b1 ,
		\o[18]_b0 ,\o[17]_b1 ,\o[17]_b0 ,\o[16]_b1 ,\o[16]_b0 ,\o[15]_b1 ,\o[15]_b0 ,\o[14]_b1 ,\o[14]_b0 ,
		\o[13]_b1 ,\o[13]_b0 ,\o[12]_b1 ,\o[12]_b0 ,\o[11]_b1 ,\o[11]_b0 ,\o[10]_b1 ,\o[10]_b0 ,\o[9]_b1 ,
		\o[9]_b0 ,\o[8]_b1 ,\o[8]_b0 ,\o[7]_b1 ,\o[7]_b0 ,\o[6]_b1 ,\o[6]_b0 ,\o[5]_b1 ,\o[5]_b0 ,
		\o[4]_b1 ,\o[4]_b0 ,\o[3]_b1 ,\o[3]_b0 ,\o[2]_b1 ,\o[2]_b0 ,\o[1]_b1 ,\o[1]_b0 ,\o[0]_b1 ,
		\o[0]_b0 ;

wire \97_ZERO_b1 , \97_ZERO_b0 , \98_ONE_b1 , \98_ONE_b0 , \99_b1 , \99_b0 , \100_b1 , \100_b0 , \101_b1 , \101_b0 , 
		\102_b1 , \102_b0 , \103_b1 , \103_b0 , \104_b1 , \104_b0 , \105_b1 , \105_b0 , \106_b1 , \106_b0 , 
		\107_b1 , \107_b0 , \108_b1 , \108_b0 , \109_b1 , \109_b0 , \110_b1 , \110_b0 , \111_b1 , \111_b0 , 
		\112_b1 , \112_b0 , \113_b1 , \113_b0 , \114_b1 , \114_b0 , \115_b1 , \115_b0 , \116_b1 , \116_b0 , 
		\117_b1 , \117_b0 , \118_b1 , \118_b0 , \119_b1 , \119_b0 , \120_b1 , \120_b0 , \121_b1 , \121_b0 , 
		\122_b1 , \122_b0 , \123_b1 , \123_b0 , \124_b1 , \124_b0 , \125_b1 , \125_b0 , \126_b1 , \126_b0 , 
		\127_b1 , \127_b0 , \128_b1 , \128_b0 , \129_b1 , \129_b0 , \130_b1 , \130_b0 , \131_b1 , \131_b0 , 
		\132_b1 , \132_b0 , \133_b1 , \133_b0 , \134_b1 , \134_b0 , \135_b1 , \135_b0 , \136_b1 , \136_b0 , 
		\137_b1 , \137_b0 , \138_b1 , \138_b0 , \139_b1 , \139_b0 , \140_b1 , \140_b0 , \141_b1 , \141_b0 , 
		\142_b1 , \142_b0 , \143_b1 , \143_b0 , \144_b1 , \144_b0 , \145_b1 , \145_b0 , \146_b1 , \146_b0 , 
		\147_b1 , \147_b0 , \148_b1 , \148_b0 , \149_b1 , \149_b0 , \150_b1 , \150_b0 , \151_b1 , \151_b0 , 
		\152_b1 , \152_b0 , \153_b1 , \153_b0 , \154_b1 , \154_b0 , \155_b1 , \155_b0 , \156_b1 , \156_b0 , 
		\157_b1 , \157_b0 , \158_b1 , \158_b0 , \159_b1 , \159_b0 , \160_b1 , \160_b0 , \161_b1 , \161_b0 , 
		\162_b1 , \162_b0 , \163_b1 , \163_b0 , \164_b1 , \164_b0 , \165_b1 , \165_b0 , \166_b1 , \166_b0 , 
		\167_b1 , \167_b0 , \168_b1 , \168_b0 , \169_b1 , \169_b0 , \170_b1 , \170_b0 , \171_b1 , \171_b0 , 
		\172_b1 , \172_b0 , \173_b1 , \173_b0 , \174_b1 , \174_b0 , \175_b1 , \175_b0 , \176_b1 , \176_b0 , 
		\177_b1 , \177_b0 , \178_b1 , \178_b0 , \179_b1 , \179_b0 , \180_b1 , \180_b0 , \181_b1 , \181_b0 , 
		\182_b1 , \182_b0 , \183_b1 , \183_b0 , \184_b1 , \184_b0 , \185_b1 , \185_b0 , \186_b1 , \186_b0 , 
		\187_b1 , \187_b0 , \188_b1 , \188_b0 , \189_b1 , \189_b0 , \190_b1 , \190_b0 , \191_b1 , \191_b0 , 
		\192_b1 , \192_b0 , \193_b1 , \193_b0 , \194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , 
		\197_b1 , \197_b0 , \198_b1 , \198_b0 , \199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , 
		\202_b1 , \202_b0 , \203_b1 , \203_b0 , \204_b1 , \204_b0 , \205_b1 , \205_b0 , \206_b1 , \206_b0 , 
		\207_b1 , \207_b0 , \208_b1 , \208_b0 , \209_b1 , \209_b0 , \210_b1 , \210_b0 , \211_b1 , \211_b0 , 
		\212_b1 , \212_b0 , \213_b1 , \213_b0 , \214_b1 , \214_b0 , \215_b1 , \215_b0 , \216_b1 , \216_b0 , 
		\217_b1 , \217_b0 , \218_b1 , \218_b0 , \219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , 
		\222_b1 , \222_b0 , \223_b1 , \223_b0 , \224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , 
		\227_b1 , \227_b0 , \228_b1 , \228_b0 , \229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , 
		\232_b1 , \232_b0 , \233_b1 , \233_b0 , \234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , 
		\237_b1 , \237_b0 , \238_b1 , \238_b0 , \239_b1 , \239_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , 
		\242_b1 , \242_b0 , \243_b1 , \243_b0 , \244_b1 , \244_b0 , \245_b1 , \245_b0 , \246_b1 , \246_b0 , 
		\247_b1 , \247_b0 , \248_b1 , \248_b0 , \249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , 
		\252_b1 , \252_b0 , \253_b1 , \253_b0 , \254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , 
		\257_b1 , \257_b0 , \258_b1 , \258_b0 , \259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , 
		\262_b1 , \262_b0 , \263_b1 , \263_b0 , \264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , 
		\267_b1 , \267_b0 , \268_b1 , \268_b0 , \269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , 
		\272_b1 , \272_b0 , \273_b1 , \273_b0 , \274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_b1 , \276_b0 , 
		\277_b1 , \277_b0 , \278_b1 , \278_b0 , \279_b1 , \279_b0 , \280_b1 , \280_b0 , \281_b1 , \281_b0 , 
		\282_b1 , \282_b0 , \283_b1 , \283_b0 , \284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , 
		\287_b1 , \287_b0 , \288_b1 , \288_b0 , \289_b1 , \289_b0 , \290_b1 , \290_b0 , \291_b1 , \291_b0 , 
		\292_b1 , \292_b0 , \293_b1 , \293_b0 , \294_b1 , \294_b0 , \295_b1 , \295_b0 , \296_b1 , \296_b0 , 
		\297_b1 , \297_b0 , \298_b1 , \298_b0 , \299_b1 , \299_b0 , \300_b1 , \300_b0 , \301_b1 , \301_b0 , 
		\302_b1 , \302_b0 , \303_b1 , \303_b0 , \304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , 
		\307_b1 , \307_b0 , \308_b1 , \308_b0 , \309_b1 , \309_b0 , \310_b1 , \310_b0 , \311_b1 , \311_b0 , 
		\312_b1 , \312_b0 , \313_b1 , \313_b0 , \314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_b1 , \316_b0 , 
		\317_b1 , \317_b0 , \318_b1 , \318_b0 , \319_b1 , \319_b0 , \320_b1 , \320_b0 , \321_b1 , \321_b0 , 
		\322_b1 , \322_b0 , \323_b1 , \323_b0 , \324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , 
		\327_b1 , \327_b0 , \328_b1 , \328_b0 , \329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_b1 , \331_b0 , 
		\332_b1 , \332_b0 , \333_b1 , \333_b0 , \334_b1 , \334_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , 
		\337_b1 , \337_b0 , \338_b1 , \338_b0 , \339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_b1 , \341_b0 , 
		\342_b1 , \342_b0 , \343_b1 , \343_b0 , \344_b1 , \344_b0 , \345_b1 , \345_b0 , \346_b1 , \346_b0 , 
		\347_b1 , \347_b0 , \348_b1 , \348_b0 , \349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , 
		\352_b1 , \352_b0 , \353_b1 , \353_b0 , \354_b1 , \354_b0 , \355_b1 , \355_b0 , \356_b1 , \356_b0 , 
		\357_b1 , \357_b0 , \358_b1 , \358_b0 , \359_b1 , \359_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , 
		\362_b1 , \362_b0 , \363_b1 , \363_b0 , \364_b1 , \364_b0 , \365_b1 , \365_b0 , \366_b1 , \366_b0 , 
		\367_b1 , \367_b0 , \368_b1 , \368_b0 , \369_b1 , \369_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , 
		\372_b1 , \372_b0 , \373_b1 , \373_b0 , \374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , 
		\377_b1 , \377_b0 , \378_b1 , \378_b0 , \379_b1 , \379_b0 , \380_b1 , \380_b0 , \381_b1 , \381_b0 , 
		\382_b1 , \382_b0 , \383_b1 , \383_b0 , \384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , 
		\387_b1 , \387_b0 , \388_b1 , \388_b0 , \389_b1 , \389_b0 , \390_b1 , \390_b0 , \391_b1 , \391_b0 , 
		\392_b1 , \392_b0 , \393_b1 , \393_b0 , \394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , 
		\397_b1 , \397_b0 , \398_b1 , \398_b0 , \399_b1 , \399_b0 , \400_b1 , \400_b0 , \401_b1 , \401_b0 , 
		\402_b1 , \402_b0 , \403_b1 , \403_b0 , \404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , 
		\407_b1 , \407_b0 , \408_b1 , \408_b0 , \409_b1 , \409_b0 , \410_b1 , \410_b0 , \411_b1 , \411_b0 , 
		\412_b1 , \412_b0 , \413_b1 , \413_b0 , \414_b1 , \414_b0 , \415_b1 , \415_b0 , \416_b1 , \416_b0 , 
		\417_b1 , \417_b0 , \418_b1 , \418_b0 , \419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , 
		\422_b1 , \422_b0 , \423_b1 , \423_b0 , \424_b1 , \424_b0 , \425_b1 , \425_b0 , \426_b1 , \426_b0 , 
		\427_b1 , \427_b0 , \428_b1 , \428_b0 , \429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , 
		\432_b1 , \432_b0 , \433_b1 , \433_b0 , \434_b1 , \434_b0 , \435_b1 , \435_b0 , \436_b1 , \436_b0 , 
		\437_b1 , \437_b0 , \438_b1 , \438_b0 , \439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , 
		\442_b1 , \442_b0 , \443_b1 , \443_b0 , \444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_b1 , \446_b0 , 
		\447_b1 , \447_b0 , \448_b1 , \448_b0 , \449_b1 , \449_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , 
		\452_b1 , \452_b0 , \453_b1 , \453_b0 , \454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_b1 , \456_b0 , 
		\457_b1 , \457_b0 , \458_b1 , \458_b0 , \459_b1 , \459_b0 , \460_b1 , \460_b0 , \461_b1 , \461_b0 , 
		\462_b1 , \462_b0 , \463_b1 , \463_b0 , \464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , 
		\467_b1 , \467_b0 , \468_b1 , \468_b0 , \469_b1 , \469_b0 , \470_b1 , \470_b0 , \471_b1 , \471_b0 , 
		\472_b1 , \472_b0 , \473_b1 , \473_b0 , \474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , 
		\477_b1 , \477_b0 , \478_b1 , \478_b0 , \479_b1 , \479_b0 , \480_b1 , \480_b0 , \481_b1 , \481_b0 , 
		\482_b1 , \482_b0 , \483_b1 , \483_b0 , \484_b1 , \484_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , 
		\487_b1 , \487_b0 , \488_b1 , \488_b0 , \489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , 
		\492_b1 , \492_b0 , \493_b1 , \493_b0 , \494_b1 , \494_b0 , \495_b1 , \495_b0 , \496_b1 , \496_b0 , 
		\497_b1 , \497_b0 , \498_b1 , \498_b0 , \499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , 
		\502_b1 , \502_b0 , \503_b1 , \503_b0 , \504_b1 , \504_b0 , \505_b1 , \505_b0 , \506_b1 , \506_b0 , 
		\507_b1 , \507_b0 , \508_b1 , \508_b0 , \509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , 
		\512_b1 , \512_b0 , \513_b1 , \513_b0 , \514_b1 , \514_b0 , \515_b1 , \515_b0 , \516_b1 , \516_b0 , 
		\517_b1 , \517_b0 , \518_b1 , \518_b0 , \519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , 
		\522_b1 , \522_b0 , \523_b1 , \523_b0 , \524_b1 , \524_b0 , \525_b1 , \525_b0 , \526_b1 , \526_b0 , 
		\527_b1 , \527_b0 , \528_b1 , \528_b0 , \529_b1 , \529_b0 , \530_b1 , \530_b0 , \531_b1 , \531_b0 , 
		\532_b1 , \532_b0 , \533_b1 , \533_b0 , \534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_b1 , \536_b0 , 
		\537_b1 , \537_b0 , \538_b1 , \538_b0 , \539_b1 , \539_b0 , \540_b1 , \540_b0 , \541_b1 , \541_b0 , 
		\542_b1 , \542_b0 , \543_b1 , \543_b0 , \544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , 
		\547_b1 , \547_b0 , \548_b1 , \548_b0 , \549_b1 , \549_b0 , \550_b1 , \550_b0 , \551_b1 , \551_b0 , 
		\552_b1 , \552_b0 , \553_b1 , \553_b0 , \554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , 
		\557_b1 , \557_b0 , \558_b1 , \558_b0 , \559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_b1 , \561_b0 , 
		\562_b1 , \562_b0 , \563_b1 , \563_b0 , \564_b1 , \564_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , 
		\567_b1 , \567_b0 , \568_b1 , \568_b0 , \569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_b1 , \571_b0 , 
		\572_b1 , \572_b0 , \573_b1 , \573_b0 , \574_b1 , \574_b0 , \575_b1 , \575_b0 , \576_b1 , \576_b0 , 
		\577_b1 , \577_b0 , \578_b1 , \578_b0 , \579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , 
		\582_b1 , \582_b0 , \583_b1 , \583_b0 , \584_b1 , \584_b0 , \585_b1 , \585_b0 , \586_b1 , \586_b0 , 
		\587_b1 , \587_b0 , \588_b1 , \588_b0 , \589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , 
		\592_b1 , \592_b0 , \593_b1 , \593_b0 , \594_b1 , \594_b0 , \595_b1 , \595_b0 , \596_b1 , \596_b0 , 
		\597_b1 , \597_b0 , \598_b1 , \598_b0 , \599_b1 , \599_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , 
		\602_b1 , \602_b0 , \603_b1 , \603_b0 , \604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_b1 , \606_b0 , 
		\607_b1 , \607_b0 , \608_b1 , \608_b0 , \609_b1 , \609_b0 , \610_b1 , \610_b0 , \611_b1 , \611_b0 , 
		\612_b1 , \612_b0 , \613_b1 , \613_b0 , \614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , 
		\617_b1 , \617_b0 , \618_b1 , \618_b0 , \619_b1 , \619_b0 , \620_b1 , \620_b0 , \621_b1 , \621_b0 , 
		\622_b1 , \622_b0 , \623_b1 , \623_b0 , \624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , 
		\627_b1 , \627_b0 , \628_b1 , \628_b0 , \629_b1 , \629_b0 , \630_b1 , \630_b0 , \631_b1 , \631_b0 , 
		\632_b1 , \632_b0 , \633_b1 , \633_b0 , \634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , 
		\637_b1 , \637_b0 , \638_b1 , \638_b0 , \639_b1 , \639_b0 , \640_b1 , \640_b0 , \641_b1 , \641_b0 , 
		\642_b1 , \642_b0 , \643_b1 , \643_b0 , \644_b1 , \644_b0 , \645_b1 , \645_b0 , \646_b1 , \646_b0 , 
		\647_b1 , \647_b0 , \648_b1 , \648_b0 , \649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , 
		\652_b1 , \652_b0 , \653_b1 , \653_b0 , \654_b1 , \654_b0 , \655_b1 , \655_b0 , \656_b1 , \656_b0 , 
		\657_b1 , \657_b0 , \658_b1 , \658_b0 , \659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , 
		\662_b1 , \662_b0 , \663_b1 , \663_b0 , \664_b1 , \664_b0 , \665_b1 , \665_b0 , \666_b1 , \666_b0 , 
		\667_b1 , \667_b0 , \668_b1 , \668_b0 , \669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , 
		\672_b1 , \672_b0 , \673_b1 , \673_b0 , \674_b1 , \674_b0 , \675_b1 , \675_b0 , \676_b1 , \676_b0 , 
		\677_b1 , \677_b0 , \678_b1 , \678_b0 , \679_b1 , \679_b0 , \680_b1 , \680_b0 , \681_b1 , \681_b0 , 
		\682_b1 , \682_b0 , \683_b1 , \683_b0 , \684_b1 , \684_b0 , \685_b1 , \685_b0 , \686_b1 , \686_b0 , 
		\687_b1 , \687_b0 , \688_b1 , \688_b0 , \689_b1 , \689_b0 , \690_b1 , \690_b0 , \691_b1 , \691_b0 , 
		\692_b1 , \692_b0 , \693_b1 , \693_b0 , \694_b1 , \694_b0 , \695_b1 , \695_b0 , \696_b1 , \696_b0 , 
		\697_b1 , \697_b0 , \698_b1 , \698_b0 , \699_b1 , \699_b0 , \700_b1 , \700_b0 , \701_b1 , \701_b0 , 
		\702_b1 , \702_b0 , \703_b1 , \703_b0 , \704_b1 , \704_b0 , \705_b1 , \705_b0 , \706_b1 , \706_b0 , 
		\707_b1 , \707_b0 , \708_b1 , \708_b0 , \709_b1 , \709_b0 , \710_b1 , \710_b0 , \711_b1 , \711_b0 , 
		\712_b1 , \712_b0 , \713_b1 , \713_b0 , \714_b1 , \714_b0 , \715_b1 , \715_b0 , \716_b1 , \716_b0 , 
		\717_b1 , \717_b0 , \718_b1 , \718_b0 , \719_b1 , \719_b0 , \720_b1 , \720_b0 , \721_b1 , \721_b0 , 
		\722_b1 , \722_b0 , \723_b1 , \723_b0 , \724_b1 , \724_b0 , \725_b1 , \725_b0 , \726_b1 , \726_b0 , 
		\727_b1 , \727_b0 , \728_b1 , \728_b0 , \729_b1 , \729_b0 , \730_b1 , \730_b0 , \731_b1 , \731_b0 , 
		\732_b1 , \732_b0 , \733_b1 , \733_b0 , \734_b1 , \734_b0 , \735_b1 , \735_b0 , \736_b1 , \736_b0 , 
		\737_b1 , \737_b0 , \738_b1 , \738_b0 , \739_b1 , \739_b0 , \740_b1 , \740_b0 , \741_b1 , \741_b0 , 
		\742_b1 , \742_b0 , \743_b1 , \743_b0 , \744_b1 , \744_b0 , \745_b1 , \745_b0 , \746_b1 , \746_b0 , 
		\747_b1 , \747_b0 , \748_b1 , \748_b0 , \749_b1 , \749_b0 , \750_b1 , \750_b0 , \751_b1 , \751_b0 , 
		\752_b1 , \752_b0 , \753_b1 , \753_b0 , \754_b1 , \754_b0 , \755_b1 , \755_b0 , \756_b1 , \756_b0 , 
		\757_b1 , \757_b0 , \758_b1 , \758_b0 , \759_b1 , \759_b0 , \760_b1 , \760_b0 , \761_b1 , \761_b0 , 
		\762_b1 , \762_b0 , \763_b1 , \763_b0 , \764_b1 , \764_b0 , \765_b1 , \765_b0 , \766_b1 , \766_b0 , 
		\767_b1 , \767_b0 , \768_b1 , \768_b0 , \769_b1 , \769_b0 , \770_b1 , \770_b0 , \771_b1 , \771_b0 , 
		\772_b1 , \772_b0 , \773_b1 , \773_b0 , \774_b1 , \774_b0 , \775_b1 , \775_b0 , \776_b1 , \776_b0 , 
		\777_b1 , \777_b0 , \778_b1 , \778_b0 , \779_b1 , \779_b0 , \780_b1 , \780_b0 , \781_b1 , \781_b0 , 
		\782_b1 , \782_b0 , \783_b1 , \783_b0 , \784_b1 , \784_b0 , \785_b1 , \785_b0 , \786_b1 , \786_b0 , 
		\787_b1 , \787_b0 , \788_b1 , \788_b0 , \789_b1 , \789_b0 , \790_b1 , \790_b0 , \791_b1 , \791_b0 , 
		\792_b1 , \792_b0 , \793_b1 , \793_b0 , \794_b1 , \794_b0 , \795_b1 , \795_b0 , \796_b1 , \796_b0 , 
		\797_b1 , \797_b0 , \798_b1 , \798_b0 , \799_b1 , \799_b0 , \800_b1 , \800_b0 , \801_b1 , \801_b0 , 
		\802_b1 , \802_b0 , \803_b1 , \803_b0 , \804_b1 , \804_b0 , \805_b1 , \805_b0 , \806_b1 , \806_b0 , 
		\807_b1 , \807_b0 , \808_b1 , \808_b0 , \809_b1 , \809_b0 , \810_b1 , \810_b0 , \811_b1 , \811_b0 , 
		\812_b1 , \812_b0 , \813_b1 , \813_b0 , \814_b1 , \814_b0 , \815_b1 , \815_b0 , \816_b1 , \816_b0 , 
		\817_b1 , \817_b0 , \818_b1 , \818_b0 , \819_b1 , \819_b0 , \820_b1 , \820_b0 , \821_b1 , \821_b0 , 
		\822_b1 , \822_b0 , \823_b1 , \823_b0 , \824_b1 , \824_b0 , \825_b1 , \825_b0 , \826_b1 , \826_b0 , 
		\827_b1 , \827_b0 , \828_b1 , \828_b0 , \829_b1 , \829_b0 , \830_b1 , \830_b0 , \831_b1 , \831_b0 , 
		\832_b1 , \832_b0 , \833_b1 , \833_b0 , \834_b1 , \834_b0 , \835_b1 , \835_b0 , \836_b1 , \836_b0 , 
		\837_b1 , \837_b0 , \838_b1 , \838_b0 , \839_b1 , \839_b0 , \840_b1 , \840_b0 , \841_b1 , \841_b0 , 
		\842_b1 , \842_b0 , \843_b1 , \843_b0 , \844_b1 , \844_b0 , \845_b1 , \845_b0 , \846_b1 , \846_b0 , 
		\847_b1 , \847_b0 , \848_b1 , \848_b0 , \849_b1 , \849_b0 , \850_b1 , \850_b0 , \851_b1 , \851_b0 , 
		\852_b1 , \852_b0 , \853_b1 , \853_b0 , \854_b1 , \854_b0 , \855_b1 , \855_b0 , \856_b1 , \856_b0 , 
		\857_b1 , \857_b0 , \858_b1 , \858_b0 , \859_b1 , \859_b0 , \860_b1 , \860_b0 , \861_b1 , \861_b0 , 
		\862_b1 , \862_b0 , \863_b1 , \863_b0 , \864_b1 , \864_b0 , \865_b1 , \865_b0 , \866_b1 , \866_b0 , 
		\867_b1 , \867_b0 , \868_b1 , \868_b0 , \869_b1 , \869_b0 , \870_b1 , \870_b0 , \871_b1 , \871_b0 , 
		\872_b1 , \872_b0 , \873_b1 , \873_b0 , \874_b1 , \874_b0 , \875_b1 , \875_b0 , \876_b1 , \876_b0 , 
		\877_b1 , \877_b0 , \878_b1 , \878_b0 , \879_b1 , \879_b0 , \880_b1 , \880_b0 , \881_b1 , \881_b0 , 
		\882_b1 , \882_b0 , \883_b1 , \883_b0 , \884_b1 , \884_b0 , \885_b1 , \885_b0 , \886_b1 , \886_b0 , 
		\887_b1 , \887_b0 , \888_b1 , \888_b0 , \889_b1 , \889_b0 , \890_b1 , \890_b0 , \891_b1 , \891_b0 , 
		\892_b1 , \892_b0 , \893_b1 , \893_b0 , \894_b1 , \894_b0 , \895_b1 , \895_b0 , \896_b1 , \896_b0 , 
		\897_b1 , \897_b0 , \898_b1 , \898_b0 , \899_b1 , \899_b0 , \900_b1 , \900_b0 , \901_b1 , \901_b0 , 
		\902_b1 , \902_b0 , \903_b1 , \903_b0 , \904_b1 , \904_b0 , \905_b1 , \905_b0 , \906_b1 , \906_b0 , 
		\907_b1 , \907_b0 , \908_b1 , \908_b0 , \909_b1 , \909_b0 , \910_b1 , \910_b0 , \911_b1 , \911_b0 , 
		\912_b1 , \912_b0 , \913_b1 , \913_b0 , \914_b1 , \914_b0 , \915_b1 , \915_b0 , \916_b1 , \916_b0 , 
		\917_b1 , \917_b0 , \918_b1 , \918_b0 , \919_b1 , \919_b0 , \920_b1 , \920_b0 , \921_b1 , \921_b0 , 
		\922_b1 , \922_b0 , \923_b1 , \923_b0 , \924_b1 , \924_b0 , \925_b1 , \925_b0 , \926_b1 , \926_b0 , 
		\927_b1 , \927_b0 , \928_b1 , \928_b0 , \929_b1 , \929_b0 , \930_b1 , \930_b0 , \931_b1 , \931_b0 , 
		\932_b1 , \932_b0 , \933_b1 , \933_b0 , \934_b1 , \934_b0 , \935_b1 , \935_b0 , \936_b1 , \936_b0 , 
		\937_b1 , \937_b0 , \938_b1 , \938_b0 , \939_b1 , \939_b0 , \940_b1 , \940_b0 , \941_b1 , \941_b0 , 
		\942_b1 , \942_b0 , \943_b1 , \943_b0 , \944_b1 , \944_b0 , \945_b1 , \945_b0 , \946_b1 , \946_b0 , 
		\947_b1 , \947_b0 , \948_b1 , \948_b0 , \949_b1 , \949_b0 , \950_b1 , \950_b0 , \951_b1 , \951_b0 , 
		\952_b1 , \952_b0 , \953_b1 , \953_b0 , \954_b1 , \954_b0 , \955_b1 , \955_b0 , \956_b1 , \956_b0 , 
		\957_b1 , \957_b0 , \958_b1 , \958_b0 , \959_b1 , \959_b0 , \960_b1 , \960_b0 , \961_b1 , \961_b0 , 
		\962_b1 , \962_b0 , \963_b1 , \963_b0 , \964_b1 , \964_b0 , \965_b1 , \965_b0 , \966_b1 , \966_b0 , 
		\967_b1 , \967_b0 , \968_b1 , \968_b0 , \969_b1 , \969_b0 , \970_b1 , \970_b0 , \971_b1 , \971_b0 , 
		\972_b1 , \972_b0 , \973_b1 , \973_b0 , \974_b1 , \974_b0 , \975_b1 , \975_b0 , \976_b1 , \976_b0 , 
		\977_b1 , \977_b0 , \978_b1 , \978_b0 , \979_b1 , \979_b0 , \980_b1 , \980_b0 , \981_b1 , \981_b0 , 
		\982_b1 , \982_b0 , \983_b1 , \983_b0 , \984_b1 , \984_b0 , \985_b1 , \985_b0 , \986_b1 , \986_b0 , 
		\987_b1 , \987_b0 , \988_b1 , \988_b0 , \989_b1 , \989_b0 , \990_b1 , \990_b0 , \991_b1 , \991_b0 , 
		\992_b1 , \992_b0 , \993_b1 , \993_b0 , \994_b1 , \994_b0 , \995_b1 , \995_b0 , \996_b1 , \996_b0 , 
		\997_b1 , \997_b0 , \998_b1 , \998_b0 , \999_b1 , \999_b0 , \1000_b1 , \1000_b0 , \1001_b1 , \1001_b0 , 
		\1002_b1 , \1002_b0 , \1003_b1 , \1003_b0 , \1004_b1 , \1004_b0 , \1005_b1 , \1005_b0 , \1006_b1 , \1006_b0 , 
		\1007_b1 , \1007_b0 , \1008_b1 , \1008_b0 , \1009_b1 , \1009_b0 , \1010_b1 , \1010_b0 , \1011_b1 , \1011_b0 , 
		\1012_b1 , \1012_b0 , \1013_b1 , \1013_b0 , \1014_b1 , \1014_b0 , \1015_b1 , \1015_b0 , \1016_b1 , \1016_b0 , 
		\1017_b1 , \1017_b0 , \1018_b1 , \1018_b0 , \1019_b1 , \1019_b0 , \1020_b1 , \1020_b0 , \1021_b1 , \1021_b0 , 
		\1022_b1 , \1022_b0 , \1023_b1 , \1023_b0 , \1024_b1 , \1024_b0 , \1025_b1 , \1025_b0 , \1026_b1 , \1026_b0 , 
		\1027_b1 , \1027_b0 , \1028_b1 , \1028_b0 , \1029_b1 , \1029_b0 , \1030_b1 , \1030_b0 , \1031_b1 , \1031_b0 , 
		\1032_b1 , \1032_b0 , \1033_b1 , \1033_b0 , \1034_b1 , \1034_b0 , \1035_b1 , \1035_b0 , \1036_b1 , \1036_b0 , 
		\1037_b1 , \1037_b0 , \1038_b1 , \1038_b0 , \1039_b1 , \1039_b0 , \1040_b1 , \1040_b0 , \1041_b1 , \1041_b0 , 
		\1042_b1 , \1042_b0 , \1043_b1 , \1043_b0 , \1044_b1 , \1044_b0 , \1045_b1 , \1045_b0 , \1046_b1 , \1046_b0 , 
		\1047_b1 , \1047_b0 , \1048_b1 , \1048_b0 , \1049_b1 , \1049_b0 , \1050_b1 , \1050_b0 , \1051_b1 , \1051_b0 , 
		\1052_b1 , \1052_b0 , \1053_b1 , \1053_b0 , \1054_b1 , \1054_b0 , \1055_b1 , \1055_b0 , \1056_b1 , \1056_b0 , 
		\1057_b1 , \1057_b0 , \1058_b1 , \1058_b0 , \1059_b1 , \1059_b0 , \1060_b1 , \1060_b0 , \1061_b1 , \1061_b0 , 
		\1062_b1 , \1062_b0 , \1063_b1 , \1063_b0 , \1064_b1 , \1064_b0 , \1065_b1 , \1065_b0 , \1066_b1 , \1066_b0 , 
		\1067_b1 , \1067_b0 , \1068_b1 , \1068_b0 , \1069_b1 , \1069_b0 , \1070_b1 , \1070_b0 , \1071_b1 , \1071_b0 , 
		\1072_b1 , \1072_b0 , \1073_b1 , \1073_b0 , \1074_b1 , \1074_b0 , \1075_b1 , \1075_b0 , \1076_b1 , \1076_b0 , 
		\1077_b1 , \1077_b0 , \1078_b1 , \1078_b0 , \1079_b1 , \1079_b0 , \1080_b1 , \1080_b0 , \1081_b1 , \1081_b0 , 
		\1082_b1 , \1082_b0 , \1083_b1 , \1083_b0 , \1084_b1 , \1084_b0 , \1085_b1 , \1085_b0 , \1086_b1 , \1086_b0 , 
		\1087_b1 , \1087_b0 , \1088_b1 , \1088_b0 , \1089_b1 , \1089_b0 , \1090_b1 , \1090_b0 , \1091_b1 , \1091_b0 , 
		\1092_b1 , \1092_b0 , \1093_b1 , \1093_b0 , \1094_b1 , \1094_b0 , \1095_b1 , \1095_b0 , \1096_b1 , \1096_b0 , 
		\1097_b1 , \1097_b0 , \1098_b1 , \1098_b0 , \1099_b1 , \1099_b0 , \1100_b1 , \1100_b0 , \1101_b1 , \1101_b0 , 
		\1102_b1 , \1102_b0 , \1103_b1 , \1103_b0 , \1104_b1 , \1104_b0 , \1105_b1 , \1105_b0 , \1106_b1 , \1106_b0 , 
		\1107_b1 , \1107_b0 , \1108_b1 , \1108_b0 , \1109_b1 , \1109_b0 , \1110_b1 , \1110_b0 , \1111_b1 , \1111_b0 , 
		\1112_b1 , \1112_b0 , \1113_b1 , \1113_b0 , \1114_b1 , \1114_b0 , \1115_b1 , \1115_b0 , \1116_b1 , \1116_b0 , 
		\1117_b1 , \1117_b0 , \1118_b1 , \1118_b0 , \1119_b1 , \1119_b0 , \1120_b1 , \1120_b0 , \1121_b1 , \1121_b0 , 
		\1122_b1 , \1122_b0 , \1123_b1 , \1123_b0 , \1124_b1 , \1124_b0 , \1125_b1 , \1125_b0 , \1126_b1 , \1126_b0 , 
		\1127_b1 , \1127_b0 , \1128_b1 , \1128_b0 , \1129_b1 , \1129_b0 , \1130_b1 , \1130_b0 , \1131_b1 , \1131_b0 , 
		\1132_b1 , \1132_b0 , \1133_b1 , \1133_b0 , \1134_b1 , \1134_b0 , \1135_b1 , \1135_b0 , \1136_b1 , \1136_b0 , 
		\1137_b1 , \1137_b0 , \1138_b1 , \1138_b0 , \1139_b1 , \1139_b0 , \1140_b1 , \1140_b0 , \1141_b1 , \1141_b0 , 
		\1142_b1 , \1142_b0 , \1143_b1 , \1143_b0 , \1144_b1 , \1144_b0 , \1145_b1 , \1145_b0 , \1146_b1 , \1146_b0 , 
		\1147_b1 , \1147_b0 , \1148_b1 , \1148_b0 , \1149_b1 , \1149_b0 , \1150_b1 , \1150_b0 , \1151_b1 , \1151_b0 , 
		\1152_b1 , \1152_b0 , \1153_b1 , \1153_b0 , \1154_b1 , \1154_b0 , \1155_b1 , \1155_b0 , \1156_b1 , \1156_b0 , 
		\1157_b1 , \1157_b0 , \1158_b1 , \1158_b0 , \1159_b1 , \1159_b0 , \1160_b1 , \1160_b0 , \1161_b1 , \1161_b0 , 
		\1162_b1 , \1162_b0 , \1163_b1 , \1163_b0 , \1164_b1 , \1164_b0 , \1165_b1 , \1165_b0 , \1166_b1 , \1166_b0 , 
		\1167_b1 , \1167_b0 , \1168_b1 , \1168_b0 , \1169_b1 , \1169_b0 , \1170_b1 , \1170_b0 , \1171_b1 , \1171_b0 , 
		\1172_b1 , \1172_b0 , \1173_b1 , \1173_b0 , \1174_b1 , \1174_b0 , \1175_b1 , \1175_b0 , \1176_b1 , \1176_b0 , 
		\1177_b1 , \1177_b0 , \1178_b1 , \1178_b0 , \1179_b1 , \1179_b0 , \1180_b1 , \1180_b0 , \1181_b1 , \1181_b0 , 
		\1182_b1 , \1182_b0 , \1183_b1 , \1183_b0 , \1184_b1 , \1184_b0 , \1185_b1 , \1185_b0 , \1186_b1 , \1186_b0 , 
		\1187_b1 , \1187_b0 , \1188_b1 , \1188_b0 , \1189_b1 , \1189_b0 , \1190_b1 , \1190_b0 , \1191_b1 , \1191_b0 , 
		\1192_b1 , \1192_b0 , \1193_b1 , \1193_b0 , \1194_b1 , \1194_b0 , \1195_b1 , \1195_b0 , \1196_b1 , \1196_b0 , 
		\1197_b1 , \1197_b0 , \1198_b1 , \1198_b0 , \1199_b1 , \1199_b0 , \1200_b1 , \1200_b0 , \1201_b1 , \1201_b0 , 
		\1202_b1 , \1202_b0 , \1203_b1 , \1203_b0 , \1204_b1 , \1204_b0 , \1205_b1 , \1205_b0 , \1206_b1 , \1206_b0 , 
		\1207_b1 , \1207_b0 , \1208_b1 , \1208_b0 , \1209_b1 , \1209_b0 , \1210_b1 , \1210_b0 , \1211_b1 , \1211_b0 , 
		\1212_b1 , \1212_b0 , \1213_b1 , \1213_b0 , \1214_b1 , \1214_b0 , \1215_b1 , \1215_b0 , \1216_b1 , \1216_b0 , 
		\1217_b1 , \1217_b0 , \1218_b1 , \1218_b0 , \1219_b1 , \1219_b0 , \1220_b1 , \1220_b0 , \1221_b1 , \1221_b0 , 
		\1222_b1 , \1222_b0 , \1223_b1 , \1223_b0 , \1224_b1 , \1224_b0 , \1225_b1 , \1225_b0 , \1226_b1 , \1226_b0 , 
		\1227_b1 , \1227_b0 , \1228_b1 , \1228_b0 , \1229_b1 , \1229_b0 , \1230_b1 , \1230_b0 , \1231_b1 , \1231_b0 , 
		\1232_b1 , \1232_b0 , \1233_b1 , \1233_b0 , \1234_b1 , \1234_b0 , \1235_b1 , \1235_b0 , \1236_b1 , \1236_b0 , 
		\1237_b1 , \1237_b0 , \1238_b1 , \1238_b0 , \1239_b1 , \1239_b0 , \1240_b1 , \1240_b0 , \1241_b1 , \1241_b0 , 
		\1242_b1 , \1242_b0 , \1243_b1 , \1243_b0 , \1244_b1 , \1244_b0 , \1245_b1 , \1245_b0 , \1246_b1 , \1246_b0 , 
		\1247_b1 , \1247_b0 , \1248_b1 , \1248_b0 , \1249_b1 , \1249_b0 , \1250_b1 , \1250_b0 , \1251_b1 , \1251_b0 , 
		\1252_b1 , \1252_b0 , \1253_b1 , \1253_b0 , \1254_b1 , \1254_b0 , \1255_b1 , \1255_b0 , \1256_b1 , \1256_b0 , 
		\1257_b1 , \1257_b0 , \1258_b1 , \1258_b0 , \1259_b1 , \1259_b0 , \1260_b1 , \1260_b0 , \1261_b1 , \1261_b0 , 
		\1262_b1 , \1262_b0 , \1263_b1 , \1263_b0 , \1264_b1 , \1264_b0 , \1265_b1 , \1265_b0 , \1266_b1 , \1266_b0 , 
		\1267_b1 , \1267_b0 , \1268_b1 , \1268_b0 , \1269_b1 , \1269_b0 , \1270_b1 , \1270_b0 , \1271_b1 , \1271_b0 , 
		\1272_b1 , \1272_b0 , \1273_b1 , \1273_b0 , \1274_b1 , \1274_b0 , \1275_b1 , \1275_b0 , \1276_b1 , \1276_b0 , 
		\1277_b1 , \1277_b0 , \1278_b1 , \1278_b0 , \1279_b1 , \1279_b0 , \1280_b1 , \1280_b0 , \1281_b1 , \1281_b0 , 
		\1282_b1 , \1282_b0 , \1283_b1 , \1283_b0 , \1284_b1 , \1284_b0 , \1285_b1 , \1285_b0 , \1286_b1 , \1286_b0 , 
		\1287_b1 , \1287_b0 , \1288_b1 , \1288_b0 , \1289_b1 , \1289_b0 , \1290_b1 , \1290_b0 , \1291_b1 , \1291_b0 , 
		\1292_b1 , \1292_b0 , \1293_b1 , \1293_b0 , \1294_b1 , \1294_b0 , \1295_b1 , \1295_b0 , \1296_b1 , \1296_b0 , 
		\1297_b1 , \1297_b0 , \1298_b1 , \1298_b0 , \1299_b1 , \1299_b0 , \1300_b1 , \1300_b0 , \1301_b1 , \1301_b0 , 
		\1302_b1 , \1302_b0 , \1303_b1 , \1303_b0 , \1304_b1 , \1304_b0 , \1305_b1 , \1305_b0 , \1306_b1 , \1306_b0 , 
		\1307_b1 , \1307_b0 , \1308_b1 , \1308_b0 , \1309_b1 , \1309_b0 , \1310_b1 , \1310_b0 , \1311_b1 , \1311_b0 , 
		\1312_b1 , \1312_b0 , \1313_b1 , \1313_b0 , \1314_b1 , \1314_b0 , \1315_b1 , \1315_b0 , \1316_b1 , \1316_b0 , 
		\1317_b1 , \1317_b0 , \1318_b1 , \1318_b0 , \1319_b1 , \1319_b0 , \1320_b1 , \1320_b0 , \1321_b1 , \1321_b0 , 
		\1322_b1 , \1322_b0 , \1323_b1 , \1323_b0 , \1324_b1 , \1324_b0 , \1325_b1 , \1325_b0 , \1326_b1 , \1326_b0 , 
		\1327_b1 , \1327_b0 , \1328_b1 , \1328_b0 , \1329_b1 , \1329_b0 , \1330_b1 , \1330_b0 , \1331_b1 , \1331_b0 , 
		\1332_b1 , \1332_b0 , \1333_b1 , \1333_b0 , \1334_b1 , \1334_b0 , \1335_b1 , \1335_b0 , \1336_b1 , \1336_b0 , 
		\1337_b1 , \1337_b0 , \1338_b1 , \1338_b0 , \1339_b1 , \1339_b0 , \1340_b1 , \1340_b0 , \1341_b1 , \1341_b0 , 
		\1342_b1 , \1342_b0 , \1343_b1 , \1343_b0 , \1344_b1 , \1344_b0 , \1345_b1 , \1345_b0 , \1346_b1 , \1346_b0 , 
		\1347_b1 , \1347_b0 , \1348_b1 , \1348_b0 , \1349_b1 , \1349_b0 , \1350_b1 , \1350_b0 , \1351_b1 , \1351_b0 , 
		\1352_b1 , \1352_b0 , \1353_b1 , \1353_b0 , \1354_b1 , \1354_b0 , \1355_b1 , \1355_b0 , \1356_b1 , \1356_b0 , 
		\1357_b1 , \1357_b0 , \1358_b1 , \1358_b0 , \1359_b1 , \1359_b0 , \1360_b1 , \1360_b0 , \1361_b1 , \1361_b0 , 
		\1362_b1 , \1362_b0 , \1363_b1 , \1363_b0 , \1364_b1 , \1364_b0 , \1365_b1 , \1365_b0 , \1366_b1 , \1366_b0 , 
		\1367_b1 , \1367_b0 , \1368_b1 , \1368_b0 , \1369_b1 , \1369_b0 , \1370_b1 , \1370_b0 , \1371_b1 , \1371_b0 , 
		\1372_b1 , \1372_b0 , \1373_b1 , \1373_b0 , \1374_b1 , \1374_b0 , \1375_b1 , \1375_b0 , \1376_b1 , \1376_b0 , 
		\1377_b1 , \1377_b0 , \1378_b1 , \1378_b0 , \1379_b1 , \1379_b0 , \1380_b1 , \1380_b0 , \1381_b1 , \1381_b0 , 
		\1382_b1 , \1382_b0 , \1383_b1 , \1383_b0 , \1384_b1 , \1384_b0 , \1385_b1 , \1385_b0 , \1386_b1 , \1386_b0 , 
		\1387_b1 , \1387_b0 , \1388_b1 , \1388_b0 , \1389_b1 , \1389_b0 , \1390_b1 , \1390_b0 , \1391_b1 , \1391_b0 , 
		\1392_b1 , \1392_b0 , \1393_b1 , \1393_b0 , \1394_b1 , \1394_b0 , \1395_b1 , \1395_b0 , \1396_b1 , \1396_b0 , 
		\1397_b1 , \1397_b0 , \1398_b1 , \1398_b0 , \1399_b1 , \1399_b0 , \1400_b1 , \1400_b0 , \1401_b1 , \1401_b0 , 
		\1402_b1 , \1402_b0 , \1403_b1 , \1403_b0 , \1404_b1 , \1404_b0 , \1405_b1 , \1405_b0 , \1406_b1 , \1406_b0 , 
		\1407_b1 , \1407_b0 , \1408_b1 , \1408_b0 , \1409_b1 , \1409_b0 , \1410_b1 , \1410_b0 , \1411_b1 , \1411_b0 , 
		\1412_b1 , \1412_b0 , \1413_b1 , \1413_b0 , \1414_b1 , \1414_b0 , \1415_b1 , \1415_b0 , \1416_b1 , \1416_b0 , 
		\1417_b1 , \1417_b0 , \1418_b1 , \1418_b0 , \1419_b1 , \1419_b0 , \1420_b1 , \1420_b0 , \1421_b1 , \1421_b0 , 
		\1422_b1 , \1422_b0 , \1423_b1 , \1423_b0 , \1424_b1 , \1424_b0 , \1425_b1 , \1425_b0 , \1426_b1 , \1426_b0 , 
		\1427_b1 , \1427_b0 , \1428_b1 , \1428_b0 , \1429_b1 , \1429_b0 , \1430_b1 , \1430_b0 , \1431_b1 , \1431_b0 , 
		\1432_b1 , \1432_b0 , \1433_b1 , \1433_b0 , \1434_b1 , \1434_b0 , \1435_b1 , \1435_b0 , \1436_b1 , \1436_b0 , 
		\1437_b1 , \1437_b0 , \1438_b1 , \1438_b0 , \1439_b1 , \1439_b0 , \1440_b1 , \1440_b0 , \1441_b1 , \1441_b0 , 
		\1442_b1 , \1442_b0 , \1443_b1 , \1443_b0 , \1444_b1 , \1444_b0 , \1445_b1 , \1445_b0 , \1446_b1 , \1446_b0 , 
		\1447_b1 , \1447_b0 , \1448_b1 , \1448_b0 , \1449_b1 , \1449_b0 , \1450_b1 , \1450_b0 , \1451_b1 , \1451_b0 , 
		\1452_b1 , \1452_b0 , \1453_b1 , \1453_b0 , \1454_b1 , \1454_b0 , \1455_b1 , \1455_b0 , \1456_b1 , \1456_b0 , 
		\1457_b1 , \1457_b0 , \1458_b1 , \1458_b0 , \1459_b1 , \1459_b0 , \1460_b1 , \1460_b0 , \1461_b1 , \1461_b0 , 
		\1462_b1 , \1462_b0 , \1463_b1 , \1463_b0 , \1464_b1 , \1464_b0 , \1465_b1 , \1465_b0 , \1466_b1 , \1466_b0 , 
		\1467_b1 , \1467_b0 , \1468_b1 , \1468_b0 , \1469_b1 , \1469_b0 , \1470_b1 , \1470_b0 , \1471_b1 , \1471_b0 , 
		\1472_b1 , \1472_b0 , \1473_b1 , \1473_b0 , \1474_b1 , \1474_b0 , \1475_b1 , \1475_b0 , \1476_b1 , \1476_b0 , 
		\1477_b1 , \1477_b0 , \1478_b1 , \1478_b0 , \1479_b1 , \1479_b0 , \1480_b1 , \1480_b0 , \1481_b1 , \1481_b0 , 
		\1482_b1 , \1482_b0 , \1483_b1 , \1483_b0 , \1484_b1 , \1484_b0 , \1485_b1 , \1485_b0 , \1486_b1 , \1486_b0 , 
		\1487_b1 , \1487_b0 , \1488_b1 , \1488_b0 , \1489_b1 , \1489_b0 , \1490_b1 , \1490_b0 , \1491_b1 , \1491_b0 , 
		\1492_b1 , \1492_b0 , \1493_b1 , \1493_b0 , \1494_b1 , \1494_b0 , \1495_b1 , \1495_b0 , \1496_b1 , \1496_b0 , 
		\1497_b1 , \1497_b0 , \1498_b1 , \1498_b0 , \1499_b1 , \1499_b0 , \1500_b1 , \1500_b0 , \1501_b1 , \1501_b0 , 
		\1502_b1 , \1502_b0 , \1503_b1 , \1503_b0 , \1504_b1 , \1504_b0 , \1505_b1 , \1505_b0 , \1506_b1 , \1506_b0 , 
		\1507_b1 , \1507_b0 , \1508_b1 , \1508_b0 , \1509_b1 , \1509_b0 , \1510_b1 , \1510_b0 , \1511_b1 , \1511_b0 , 
		\1512_b1 , \1512_b0 , \1513_b1 , \1513_b0 , \1514_b1 , \1514_b0 , \1515_b1 , \1515_b0 , \1516_b1 , \1516_b0 , 
		\1517_b1 , \1517_b0 , \1518_b1 , \1518_b0 , \1519_b1 , \1519_b0 , \1520_b1 , \1520_b0 , \1521_b1 , \1521_b0 , 
		\1522_b1 , \1522_b0 , \1523_b1 , \1523_b0 , \1524_b1 , \1524_b0 , \1525_b1 , \1525_b0 , \1526_b1 , \1526_b0 , 
		\1527_b1 , \1527_b0 , \1528_b1 , \1528_b0 , \1529_b1 , \1529_b0 , \1530_b1 , \1530_b0 , \1531_b1 , \1531_b0 , 
		\1532_b1 , \1532_b0 , \1533_b1 , \1533_b0 , \1534_b1 , \1534_b0 , \1535_b1 , \1535_b0 , \1536_b1 , \1536_b0 , 
		\1537_b1 , \1537_b0 , \1538_b1 , \1538_b0 , \1539_b1 , \1539_b0 , \1540_b1 , \1540_b0 , \1541_b1 , \1541_b0 , 
		\1542_b1 , \1542_b0 , \1543_b1 , \1543_b0 , \1544_b1 , \1544_b0 , \1545_b1 , \1545_b0 , \1546_b1 , \1546_b0 , 
		\1547_b1 , \1547_b0 , \1548_b1 , \1548_b0 , \1549_b1 , \1549_b0 , \1550_b1 , \1550_b0 , \1551_b1 , \1551_b0 , 
		\1552_b1 , \1552_b0 , \1553_b1 , \1553_b0 , \1554_b1 , \1554_b0 , \1555_b1 , \1555_b0 , \1556_b1 , \1556_b0 , 
		\1557_b1 , \1557_b0 , \1558_b1 , \1558_b0 , \1559_b1 , \1559_b0 , \1560_b1 , \1560_b0 , \1561_b1 , \1561_b0 , 
		\1562_b1 , \1562_b0 , \1563_b1 , \1563_b0 , \1564_b1 , \1564_b0 , \1565_b1 , \1565_b0 , \1566_b1 , \1566_b0 , 
		\1567_b1 , \1567_b0 , \1568_b1 , \1568_b0 , \1569_b1 , \1569_b0 , \1570_b1 , \1570_b0 , \1571_b1 , \1571_b0 , 
		\1572_b1 , \1572_b0 , \1573_b1 , \1573_b0 , \1574_b1 , \1574_b0 , \1575_b1 , \1575_b0 , \1576_b1 , \1576_b0 , 
		\1577_b1 , \1577_b0 , \1578_b1 , \1578_b0 , \1579_b1 , \1579_b0 , \1580_b1 , \1580_b0 , \1581_b1 , \1581_b0 , 
		\1582_b1 , \1582_b0 , \1583_b1 , \1583_b0 , \1584_b1 , \1584_b0 , \1585_b1 , \1585_b0 , \1586_b1 , \1586_b0 , 
		\1587_b1 , \1587_b0 , \1588_b1 , \1588_b0 , \1589_b1 , \1589_b0 , \1590_b1 , \1590_b0 , \1591_b1 , \1591_b0 , 
		\1592_b1 , \1592_b0 , \1593_b1 , \1593_b0 , \1594_b1 , \1594_b0 , \1595_b1 , \1595_b0 , \1596_b1 , \1596_b0 , 
		\1597_b1 , \1597_b0 , \1598_b1 , \1598_b0 , \1599_b1 , \1599_b0 , \1600_b1 , \1600_b0 , \1601_b1 , \1601_b0 , 
		\1602_b1 , \1602_b0 , \1603_b1 , \1603_b0 , \1604_b1 , \1604_b0 , \1605_b1 , \1605_b0 , \1606_b1 , \1606_b0 , 
		\1607_b1 , \1607_b0 , \1608_b1 , \1608_b0 , \1609_b1 , \1609_b0 , \1610_b1 , \1610_b0 , \1611_b1 , \1611_b0 , 
		\1612_b1 , \1612_b0 , \1613_b1 , \1613_b0 , \1614_b1 , \1614_b0 , \1615_b1 , \1615_b0 , \1616_b1 , \1616_b0 , 
		\1617_b1 , \1617_b0 , \1618_b1 , \1618_b0 , \1619_b1 , \1619_b0 , \1620_b1 , \1620_b0 , \1621_b1 , \1621_b0 , 
		\1622_b1 , \1622_b0 , \1623_b1 , \1623_b0 , \1624_b1 , \1624_b0 , \1625_b1 , \1625_b0 , \1626_b1 , \1626_b0 , 
		\1627_b1 , \1627_b0 , \1628_b1 , \1628_b0 , \1629_b1 , \1629_b0 , \1630_b1 , \1630_b0 , \1631_b1 , \1631_b0 , 
		\1632_b1 , \1632_b0 , \1633_b1 , \1633_b0 , \1634_b1 , \1634_b0 , \1635_b1 , \1635_b0 , \1636_b1 , \1636_b0 , 
		\1637_b1 , \1637_b0 , \1638_b1 , \1638_b0 , \1639_b1 , \1639_b0 , \1640_b1 , \1640_b0 , \1641_b1 , \1641_b0 , 
		\1642_b1 , \1642_b0 , \1643_b1 , \1643_b0 , \1644_b1 , \1644_b0 , \1645_b1 , \1645_b0 , \1646_b1 , \1646_b0 , 
		\1647_b1 , \1647_b0 , \1648_b1 , \1648_b0 , \1649_b1 , \1649_b0 , \1650_b1 , \1650_b0 , \1651_b1 , \1651_b0 , 
		\1652_b1 , \1652_b0 , \1653_b1 , \1653_b0 , \1654_b1 , \1654_b0 , \1655_b1 , \1655_b0 , \1656_b1 , \1656_b0 , 
		\1657_b1 , \1657_b0 , \1658_b1 , \1658_b0 , \1659_b1 , \1659_b0 , \1660_b1 , \1660_b0 , \1661_b1 , \1661_b0 , 
		\1662_b1 , \1662_b0 , \1663_b1 , \1663_b0 , \1664_b1 , \1664_b0 , \1665_b1 , \1665_b0 , \1666_b1 , \1666_b0 , 
		\1667_b1 , \1667_b0 , \1668_b1 , \1668_b0 , \1669_b1 , \1669_b0 , \1670_b1 , \1670_b0 , \1671_b1 , \1671_b0 , 
		\1672_b1 , \1672_b0 , \1673_b1 , \1673_b0 , \1674_b1 , \1674_b0 , \1675_b1 , \1675_b0 , \1676_b1 , \1676_b0 , 
		\1677_b1 , \1677_b0 , \1678_b1 , \1678_b0 , \1679_b1 , \1679_b0 , \1680_b1 , \1680_b0 , \1681_b1 , \1681_b0 , 
		\1682_b1 , \1682_b0 , \1683_b1 , \1683_b0 , \1684_b1 , \1684_b0 , \1685_b1 , \1685_b0 , \1686_b1 , \1686_b0 , 
		\1687_b1 , \1687_b0 , \1688_b1 , \1688_b0 , \1689_b1 , \1689_b0 , \1690_b1 , \1690_b0 , \1691_b1 , \1691_b0 , 
		\1692_b1 , \1692_b0 , \1693_b1 , \1693_b0 , \1694_b1 , \1694_b0 , \1695_b1 , \1695_b0 , \1696_b1 , \1696_b0 , 
		\1697_b1 , \1697_b0 , \1698_b1 , \1698_b0 , \1699_b1 , \1699_b0 , \1700_b1 , \1700_b0 , \1701_b1 , \1701_b0 , 
		\1702_b1 , \1702_b0 , \1703_b1 , \1703_b0 , \1704_b1 , \1704_b0 , \1705_b1 , \1705_b0 , \1706_b1 , \1706_b0 , 
		\1707_b1 , \1707_b0 , \1708_b1 , \1708_b0 , \1709_b1 , \1709_b0 , \1710_b1 , \1710_b0 , \1711_b1 , \1711_b0 , 
		\1712_b1 , \1712_b0 , \1713_b1 , \1713_b0 , \1714_b1 , \1714_b0 , \1715_b1 , \1715_b0 , \1716_b1 , \1716_b0 , 
		\1717_b1 , \1717_b0 , \1718_b1 , \1718_b0 , \1719_b1 , \1719_b0 , \1720_b1 , \1720_b0 , \1721_b1 , \1721_b0 , 
		\1722_b1 , \1722_b0 , \1723_b1 , \1723_b0 , \1724_b1 , \1724_b0 , \1725_b1 , \1725_b0 , \1726_b1 , \1726_b0 , 
		\1727_b1 , \1727_b0 , \1728_b1 , \1728_b0 , \1729_b1 , \1729_b0 , \1730_b1 , \1730_b0 , \1731_b1 , \1731_b0 , 
		\1732_b1 , \1732_b0 , \1733_b1 , \1733_b0 , \1734_b1 , \1734_b0 , \1735_b1 , \1735_b0 , \1736_b1 , \1736_b0 , 
		\1737_b1 , \1737_b0 , \1738_b1 , \1738_b0 , \1739_b1 , \1739_b0 , \1740_b1 , \1740_b0 , \1741_b1 , \1741_b0 , 
		\1742_b1 , \1742_b0 , \1743_b1 , \1743_b0 , \1744_b1 , \1744_b0 , \1745_b1 , \1745_b0 , \1746_b1 , \1746_b0 , 
		\1747_b1 , \1747_b0 , \1748_b1 , \1748_b0 , \1749_b1 , \1749_b0 , \1750_b1 , \1750_b0 , \1751_b1 , \1751_b0 , 
		\1752_b1 , \1752_b0 , \1753_b1 , \1753_b0 , \1754_b1 , \1754_b0 , \1755_b1 , \1755_b0 , \1756_b1 , \1756_b0 , 
		\1757_b1 , \1757_b0 , \1758_b1 , \1758_b0 , \1759_b1 , \1759_b0 , \1760_b1 , \1760_b0 , \1761_b1 , \1761_b0 , 
		\1762_b1 , \1762_b0 , \1763_b1 , \1763_b0 , \1764_b1 , \1764_b0 , \1765_b1 , \1765_b0 , \1766_b1 , \1766_b0 , 
		\1767_b1 , \1767_b0 , \1768_b1 , \1768_b0 , \1769_b1 , \1769_b0 , \1770_b1 , \1770_b0 , \1771_b1 , \1771_b0 , 
		\1772_b1 , \1772_b0 , \1773_b1 , \1773_b0 , \1774_b1 , \1774_b0 , \1775_b1 , \1775_b0 , \1776_b1 , \1776_b0 , 
		\1777_b1 , \1777_b0 , \1778_b1 , \1778_b0 , \1779_b1 , \1779_b0 , \1780_b1 , \1780_b0 , \1781_b1 , \1781_b0 , 
		\1782_b1 , \1782_b0 , \1783_b1 , \1783_b0 , \1784_b1 , \1784_b0 , \1785_b1 , \1785_b0 , \1786_b1 , \1786_b0 , 
		\1787_b1 , \1787_b0 , \1788_b1 , \1788_b0 , \1789_b1 , \1789_b0 , \1790_b1 , \1790_b0 , \1791_b1 , \1791_b0 , 
		\1792_b1 , \1792_b0 , \1793_b1 , \1793_b0 , \1794_b1 , \1794_b0 , \1795_b1 , \1795_b0 , \1796_b1 , \1796_b0 , 
		\1797_b1 , \1797_b0 , \1798_b1 , \1798_b0 , \1799_b1 , \1799_b0 , \1800_b1 , \1800_b0 , \1801_b1 , \1801_b0 , 
		\1802_b1 , \1802_b0 , \1803_b1 , \1803_b0 , \1804_b1 , \1804_b0 , \1805_b1 , \1805_b0 , \1806_b1 , \1806_b0 , 
		\1807_b1 , \1807_b0 , \1808_b1 , \1808_b0 , \1809_b1 , \1809_b0 , \1810_b1 , \1810_b0 , \1811_b1 , \1811_b0 , 
		\1812_b1 , \1812_b0 , \1813_b1 , \1813_b0 , \1814_b1 , \1814_b0 , \1815_b1 , \1815_b0 , \1816_b1 , \1816_b0 , 
		\1817_b1 , \1817_b0 , \1818_b1 , \1818_b0 , \1819_b1 , \1819_b0 , \1820_b1 , \1820_b0 , \1821_b1 , \1821_b0 , 
		\1822_b1 , \1822_b0 , \1823_b1 , \1823_b0 , \1824_b1 , \1824_b0 , \1825_b1 , \1825_b0 , \1826_b1 , \1826_b0 , 
		\1827_b1 , \1827_b0 , \1828_b1 , \1828_b0 , \1829_b1 , \1829_b0 , \1830_b1 , \1830_b0 , \1831_b1 , \1831_b0 , 
		\1832_b1 , \1832_b0 , \1833_b1 , \1833_b0 , \1834_b1 , \1834_b0 , \1835_b1 , \1835_b0 , \1836_b1 , \1836_b0 , 
		\1837_b1 , \1837_b0 , \1838_b1 , \1838_b0 , \1839_b1 , \1839_b0 , \1840_b1 , \1840_b0 , \1841_b1 , \1841_b0 , 
		\1842_b1 , \1842_b0 , \1843_b1 , \1843_b0 , \1844_b1 , \1844_b0 , \1845_b1 , \1845_b0 , \1846_b1 , \1846_b0 , 
		\1847_b1 , \1847_b0 , \1848_b1 , \1848_b0 , \1849_b1 , \1849_b0 , \1850_b1 , \1850_b0 , \1851_b1 , \1851_b0 , 
		\1852_b1 , \1852_b0 , \1853_b1 , \1853_b0 , \1854_b1 , \1854_b0 , \1855_b1 , \1855_b0 , \1856_b1 , \1856_b0 , 
		\1857_b1 , \1857_b0 , \1858_b1 , \1858_b0 , \1859_b1 , \1859_b0 , \1860_b1 , \1860_b0 , \1861_b1 , \1861_b0 , 
		\1862_b1 , \1862_b0 , \1863_b1 , \1863_b0 , \1864_b1 , \1864_b0 , \1865_b1 , \1865_b0 , \1866_b1 , \1866_b0 , 
		\1867_b1 , \1867_b0 , \1868_b1 , \1868_b0 , \1869_b1 , \1869_b0 , \1870_b1 , \1870_b0 , \1871_b1 , \1871_b0 , 
		\1872_b1 , \1872_b0 , \1873_b1 , \1873_b0 , \1874_b1 , \1874_b0 , \1875_b1 , \1875_b0 , \1876_b1 , \1876_b0 , 
		\1877_b1 , \1877_b0 , \1878_b1 , \1878_b0 , \1879_b1 , \1879_b0 , \1880_b1 , \1880_b0 , \1881_b1 , \1881_b0 , 
		\1882_b1 , \1882_b0 , \1883_b1 , \1883_b0 , \1884_b1 , \1884_b0 , \1885_b1 , \1885_b0 , \1886_b1 , \1886_b0 , 
		\1887_b1 , \1887_b0 , \1888_b1 , \1888_b0 , \1889_b1 , \1889_b0 , \1890_b1 , \1890_b0 , \1891_b1 , \1891_b0 , 
		\1892_b1 , \1892_b0 , \1893_b1 , \1893_b0 , \1894_b1 , \1894_b0 , \1895_b1 , \1895_b0 , \1896_b1 , \1896_b0 , 
		\1897_b1 , \1897_b0 , \1898_b1 , \1898_b0 , \1899_b1 , \1899_b0 , \1900_b1 , \1900_b0 , \1901_b1 , \1901_b0 , 
		\1902_b1 , \1902_b0 , \1903_b1 , \1903_b0 , \1904_b1 , \1904_b0 , \1905_b1 , \1905_b0 , \1906_b1 , \1906_b0 , 
		\1907_b1 , \1907_b0 , \1908_b1 , \1908_b0 , \1909_b1 , \1909_b0 , \1910_b1 , \1910_b0 , \1911_b1 , \1911_b0 , 
		\1912_b1 , \1912_b0 , \1913_b1 , \1913_b0 , \1914_b1 , \1914_b0 , \1915_b1 , \1915_b0 , \1916_b1 , \1916_b0 , 
		\1917_b1 , \1917_b0 , \1918_b1 , \1918_b0 , \1919_b1 , \1919_b0 , \1920_b1 , \1920_b0 , \1921_b1 , \1921_b0 , 
		\1922_b1 , \1922_b0 , \1923_b1 , \1923_b0 , \1924_b1 , \1924_b0 , \1925_b1 , \1925_b0 , \1926_b1 , \1926_b0 , 
		\1927_b1 , \1927_b0 , \1928_b1 , \1928_b0 , \1929_b1 , \1929_b0 , \1930_b1 , \1930_b0 , \1931_b1 , \1931_b0 , 
		\1932_b1 , \1932_b0 , \1933_b1 , \1933_b0 , \1934_b1 , \1934_b0 , \1935_b1 , \1935_b0 , \1936_b1 , \1936_b0 , 
		\1937_b1 , \1937_b0 , \1938_b1 , \1938_b0 , \1939_b1 , \1939_b0 , \1940_b1 , \1940_b0 , \1941_b1 , \1941_b0 , 
		\1942_b1 , \1942_b0 , \1943_b1 , \1943_b0 , \1944_b1 , \1944_b0 , \1945_b1 , \1945_b0 , \1946_b1 , \1946_b0 , 
		\1947_b1 , \1947_b0 , \1948_b1 , \1948_b0 , \1949_b1 , \1949_b0 , \1950_b1 , \1950_b0 , \1951_b1 , \1951_b0 , 
		\1952_b1 , \1952_b0 , \1953_b1 , \1953_b0 , \1954_b1 , \1954_b0 , \1955_b1 , \1955_b0 , \1956_b1 , \1956_b0 , 
		\1957_b1 , \1957_b0 , \1958_b1 , \1958_b0 , \1959_b1 , \1959_b0 , \1960_b1 , \1960_b0 , \1961_b1 , \1961_b0 , 
		\1962_b1 , \1962_b0 , \1963_b1 , \1963_b0 , \1964_b1 , \1964_b0 , \1965_b1 , \1965_b0 , \1966_b1 , \1966_b0 , 
		\1967_b1 , \1967_b0 , \1968_b1 , \1968_b0 , \1969_b1 , \1969_b0 , \1970_b1 , \1970_b0 , \1971_b1 , \1971_b0 , 
		\1972_b1 , \1972_b0 , \1973_b1 , \1973_b0 , \1974_b1 , \1974_b0 , \1975_b1 , \1975_b0 , \1976_b1 , \1976_b0 , 
		\1977_b1 , \1977_b0 , \1978_b1 , \1978_b0 , \1979_b1 , \1979_b0 , \1980_b1 , \1980_b0 , \1981_b1 , \1981_b0 , 
		\1982_b1 , \1982_b0 , \1983_b1 , \1983_b0 , \1984_b1 , \1984_b0 , \1985_b1 , \1985_b0 , \1986_b1 , \1986_b0 , 
		\1987_b1 , \1987_b0 , \1988_b1 , \1988_b0 , \1989_b1 , \1989_b0 , \1990_b1 , \1990_b0 , \1991_b1 , \1991_b0 , 
		\1992_b1 , \1992_b0 , \1993_b1 , \1993_b0 , \1994_b1 , \1994_b0 , \1995_b1 , \1995_b0 , \1996_b1 , \1996_b0 , 
		\1997_b1 , \1997_b0 , \1998_b1 , \1998_b0 , \1999_b1 , \1999_b0 , \2000_b1 , \2000_b0 , \2001_b1 , \2001_b0 , 
		\2002_b1 , \2002_b0 , \2003_b1 , \2003_b0 , \2004_b1 , \2004_b0 , \2005_b1 , \2005_b0 , \2006_b1 , \2006_b0 , 
		\2007_b1 , \2007_b0 , \2008_b1 , \2008_b0 , \2009_b1 , \2009_b0 , \2010_b1 , \2010_b0 , \2011_b1 , \2011_b0 , 
		\2012_b1 , \2012_b0 , \2013_b1 , \2013_b0 , \2014_b1 , \2014_b0 , \2015_b1 , \2015_b0 , \2016_b1 , \2016_b0 , 
		\2017_b1 , \2017_b0 , \2018_b1 , \2018_b0 , \2019_b1 , \2019_b0 , \2020_b1 , \2020_b0 , \2021_b1 , \2021_b0 , 
		\2022_b1 , \2022_b0 , \2023_b1 , \2023_b0 , \2024_b1 , \2024_b0 , \2025_b1 , \2025_b0 , \2026_b1 , \2026_b0 , 
		\2027_b1 , \2027_b0 , \2028_b1 , \2028_b0 , \2029_b1 , \2029_b0 , \2030_b1 , \2030_b0 , \2031_b1 , \2031_b0 , 
		\2032_b1 , \2032_b0 , \2033_b1 , \2033_b0 , \2034_b1 , \2034_b0 , \2035_b1 , \2035_b0 , \2036_b1 , \2036_b0 , 
		\2037_b1 , \2037_b0 , \2038_b1 , \2038_b0 , \2039_b1 , \2039_b0 , \2040_b1 , \2040_b0 , \2041_b1 , \2041_b0 , 
		\2042_b1 , \2042_b0 , \2043_b1 , \2043_b0 , \2044_b1 , \2044_b0 , \2045_b1 , \2045_b0 , \2046_b1 , \2046_b0 , 
		\2047_b1 , \2047_b0 , \2048_b1 , \2048_b0 , \2049_b1 , \2049_b0 , \2050_b1 , \2050_b0 , \2051_b1 , \2051_b0 , 
		\2052_b1 , \2052_b0 , \2053_b1 , \2053_b0 , \2054_b1 , \2054_b0 , \2055_b1 , \2055_b0 , \2056_b1 , \2056_b0 , 
		\2057_b1 , \2057_b0 , \2058_b1 , \2058_b0 , \2059_b1 , \2059_b0 , \2060_b1 , \2060_b0 , \2061_b1 , \2061_b0 , 
		\2062_b1 , \2062_b0 , \2063_b1 , \2063_b0 , \2064_b1 , \2064_b0 , \2065_b1 , \2065_b0 , \2066_b1 , \2066_b0 , 
		\2067_b1 , \2067_b0 , \2068_b1 , \2068_b0 , \2069_b1 , \2069_b0 , \2070_b1 , \2070_b0 , \2071_b1 , \2071_b0 , 
		\2072_b1 , \2072_b0 , \2073_b1 , \2073_b0 , \2074_b1 , \2074_b0 , \2075_b1 , \2075_b0 , \2076_b1 , \2076_b0 , 
		\2077_b1 , \2077_b0 , \2078_b1 , \2078_b0 , \2079_b1 , \2079_b0 , \2080_b1 , \2080_b0 , \2081_b1 , \2081_b0 , 
		\2082_b1 , \2082_b0 , \2083_b1 , \2083_b0 , \2084_b1 , \2084_b0 , \2085_b1 , \2085_b0 , \2086_b1 , \2086_b0 , 
		\2087_b1 , \2087_b0 , \2088_b1 , \2088_b0 , \2089_b1 , \2089_b0 , \2090_b1 , \2090_b0 , \2091_b1 , \2091_b0 , 
		\2092_b1 , \2092_b0 , \2093_b1 , \2093_b0 , \2094_b1 , \2094_b0 , \2095_b1 , \2095_b0 , \2096_b1 , \2096_b0 , 
		\2097_b1 , \2097_b0 , \2098_b1 , \2098_b0 , \2099_b1 , \2099_b0 , \2100_b1 , \2100_b0 , \2101_b1 , \2101_b0 , 
		\2102_b1 , \2102_b0 , \2103_b1 , \2103_b0 , \2104_b1 , \2104_b0 , \2105_b1 , \2105_b0 , \2106_b1 , \2106_b0 , 
		\2107_b1 , \2107_b0 , \2108_b1 , \2108_b0 , \2109_b1 , \2109_b0 , \2110_b1 , \2110_b0 , \2111_b1 , \2111_b0 , 
		\2112_b1 , \2112_b0 , \2113_b1 , \2113_b0 , \2114_b1 , \2114_b0 , \2115_b1 , \2115_b0 , \2116_b1 , \2116_b0 , 
		\2117_b1 , \2117_b0 , \2118_b1 , \2118_b0 , \2119_b1 , \2119_b0 , \2120_b1 , \2120_b0 , \2121_b1 , \2121_b0 , 
		\2122_b1 , \2122_b0 , \2123_b1 , \2123_b0 , \2124_b1 , \2124_b0 , \2125_b1 , \2125_b0 , \2126_b1 , \2126_b0 , 
		\2127_b1 , \2127_b0 , \2128_b1 , \2128_b0 , \2129_b1 , \2129_b0 , \2130_b1 , \2130_b0 , \2131_b1 , \2131_b0 , 
		\2132_b1 , \2132_b0 , \2133_b1 , \2133_b0 , \2134_b1 , \2134_b0 , \2135_b1 , \2135_b0 , \2136_b1 , \2136_b0 , 
		\2137_b1 , \2137_b0 , \2138_b1 , \2138_b0 , \2139_b1 , \2139_b0 , \2140_b1 , \2140_b0 , \2141_b1 , \2141_b0 , 
		\2142_b1 , \2142_b0 , \2143_b1 , \2143_b0 , \2144_b1 , \2144_b0 , \2145_b1 , \2145_b0 , \2146_b1 , \2146_b0 , 
		\2147_b1 , \2147_b0 , \2148_b1 , \2148_b0 , \2149_b1 , \2149_b0 , \2150_b1 , \2150_b0 , \2151_b1 , \2151_b0 , 
		\2152_b1 , \2152_b0 , \2153_b1 , \2153_b0 , \2154_b1 , \2154_b0 , \2155_b1 , \2155_b0 , \2156_b1 , \2156_b0 , 
		\2157_b1 , \2157_b0 , \2158_b1 , \2158_b0 , \2159_b1 , \2159_b0 , \2160_b1 , \2160_b0 , \2161_b1 , \2161_b0 , 
		\2162_b1 , \2162_b0 , \2163_b1 , \2163_b0 , \2164_b1 , \2164_b0 , \2165_b1 , \2165_b0 , \2166_b1 , \2166_b0 , 
		\2167_b1 , \2167_b0 , \2168_b1 , \2168_b0 , \2169_b1 , \2169_b0 , \2170_b1 , \2170_b0 , \2171_b1 , \2171_b0 , 
		\2172_b1 , \2172_b0 , \2173_b1 , \2173_b0 , \2174_b1 , \2174_b0 , \2175_b1 , \2175_b0 , \2176_b1 , \2176_b0 , 
		\2177_b1 , \2177_b0 , \2178_b1 , \2178_b0 , \2179_b1 , \2179_b0 , \2180_b1 , \2180_b0 , \2181_b1 , \2181_b0 , 
		\2182_b1 , \2182_b0 , \2183_b1 , \2183_b0 , \2184_b1 , \2184_b0 , \2185_b1 , \2185_b0 , \2186_b1 , \2186_b0 , 
		\2187_b1 , \2187_b0 , \2188_b1 , \2188_b0 , \2189_b1 , \2189_b0 , \2190_b1 , \2190_b0 , \2191_b1 , \2191_b0 , 
		\2192_b1 , \2192_b0 , \2193_b1 , \2193_b0 , \2194_b1 , \2194_b0 , \2195_b1 , \2195_b0 , \2196_b1 , \2196_b0 , 
		\2197_b1 , \2197_b0 , \2198_b1 , \2198_b0 , \2199_b1 , \2199_b0 , \2200_b1 , \2200_b0 , \2201_b1 , \2201_b0 , 
		\2202_b1 , \2202_b0 , \2203_b1 , \2203_b0 , \2204_b1 , \2204_b0 , \2205_b1 , \2205_b0 , \2206_b1 , \2206_b0 , 
		\2207_b1 , \2207_b0 , \2208_b1 , \2208_b0 , \2209_b1 , \2209_b0 , \2210_b1 , \2210_b0 , \2211_b1 , \2211_b0 , 
		\2212_b1 , \2212_b0 , \2213_b1 , \2213_b0 , \2214_b1 , \2214_b0 , \2215_b1 , \2215_b0 , \2216_b1 , \2216_b0 , 
		\2217_b1 , \2217_b0 , \2218_b1 , \2218_b0 , \2219_b1 , \2219_b0 , \2220_b1 , \2220_b0 , \2221_b1 , \2221_b0 , 
		\2222_b1 , \2222_b0 , \2223_b1 , \2223_b0 , \2224_b1 , \2224_b0 , \2225_b1 , \2225_b0 , \2226_b1 , \2226_b0 , 
		\2227_b1 , \2227_b0 , \2228_b1 , \2228_b0 , \2229_b1 , \2229_b0 , \2230_b1 , \2230_b0 , \2231_b1 , \2231_b0 , 
		\2232_b1 , \2232_b0 , \2233_b1 , \2233_b0 , \2234_b1 , \2234_b0 , \2235_b1 , \2235_b0 , \2236_b1 , \2236_b0 , 
		\2237_b1 , \2237_b0 , \2238_b1 , \2238_b0 , \2239_b1 , \2239_b0 , \2240_b1 , \2240_b0 , \2241_b1 , \2241_b0 , 
		\2242_b1 , \2242_b0 , \2243_b1 , \2243_b0 , \2244_b1 , \2244_b0 , \2245_b1 , \2245_b0 , \2246_b1 , \2246_b0 , 
		\2247_b1 , \2247_b0 , \2248_b1 , \2248_b0 , \2249_b1 , \2249_b0 , \2250_b1 , \2250_b0 , \2251_b1 , \2251_b0 , 
		\2252_b1 , \2252_b0 , \2253_b1 , \2253_b0 , \2254_b1 , \2254_b0 , \2255_b1 , \2255_b0 , \2256_b1 , \2256_b0 , 
		\2257_b1 , \2257_b0 , \2258_b1 , \2258_b0 , \2259_b1 , \2259_b0 , \2260_b1 , \2260_b0 , \2261_b1 , \2261_b0 , 
		\2262_b1 , \2262_b0 , \2263_b1 , \2263_b0 , \2264_b1 , \2264_b0 , \2265_b1 , \2265_b0 , \2266_b1 , \2266_b0 , 
		\2267_b1 , \2267_b0 , \2268_b1 , \2268_b0 , \2269_b1 , \2269_b0 , \2270_b1 , \2270_b0 , \2271_b1 , \2271_b0 , 
		\2272_b1 , \2272_b0 , \2273_b1 , \2273_b0 , \2274_b1 , \2274_b0 , \2275_b1 , \2275_b0 , \2276_b1 , \2276_b0 , 
		\2277_b1 , \2277_b0 , \2278_b1 , \2278_b0 , \2279_b1 , \2279_b0 , \2280_b1 , \2280_b0 , \2281_b1 , \2281_b0 , 
		\2282_b1 , \2282_b0 , \2283_b1 , \2283_b0 , \2284_b1 , \2284_b0 , \2285_b1 , \2285_b0 , \2286_b1 , \2286_b0 , 
		\2287_b1 , \2287_b0 , \2288_b1 , \2288_b0 , \2289_b1 , \2289_b0 , \2290_b1 , \2290_b0 , \2291_b1 , \2291_b0 , 
		\2292_b1 , \2292_b0 , \2293_b1 , \2293_b0 , \2294_b1 , \2294_b0 , \2295_b1 , \2295_b0 , \2296_b1 , \2296_b0 , 
		\2297_b1 , \2297_b0 , \2298_b1 , \2298_b0 , \2299_b1 , \2299_b0 , \2300_b1 , \2300_b0 , \2301_b1 , \2301_b0 , 
		\2302_b1 , \2302_b0 , \2303_b1 , \2303_b0 , \2304_b1 , \2304_b0 , \2305_b1 , \2305_b0 , \2306_b1 , \2306_b0 , 
		\2307_b1 , \2307_b0 , \2308_b1 , \2308_b0 , \2309_b1 , \2309_b0 , \2310_b1 , \2310_b0 , \2311_b1 , \2311_b0 , 
		\2312_b1 , \2312_b0 , \2313_b1 , \2313_b0 , \2314_b1 , \2314_b0 , \2315_b1 , \2315_b0 , \2316_b1 , \2316_b0 , 
		\2317_b1 , \2317_b0 , \2318_b1 , \2318_b0 , \2319_b1 , \2319_b0 , \2320_b1 , \2320_b0 , \2321_b1 , \2321_b0 , 
		\2322_b1 , \2322_b0 , \2323_b1 , \2323_b0 , \2324_b1 , \2324_b0 , \2325_b1 , \2325_b0 , \2326_b1 , \2326_b0 , 
		\2327_b1 , \2327_b0 , \2328_b1 , \2328_b0 , \2329_b1 , \2329_b0 , \2330_b1 , \2330_b0 , \2331_b1 , \2331_b0 , 
		\2332_b1 , \2332_b0 , \2333_b1 , \2333_b0 , \2334_b1 , \2334_b0 , \2335_b1 , \2335_b0 , \2336_b1 , \2336_b0 , 
		\2337_b1 , \2337_b0 , \2338_b1 , \2338_b0 , \2339_b1 , \2339_b0 , \2340_b1 , \2340_b0 , \2341_b1 , \2341_b0 , 
		\2342_b1 , \2342_b0 , \2343_b1 , \2343_b0 , \2344_b1 , \2344_b0 , \2345_b1 , \2345_b0 , \2346_b1 , \2346_b0 , 
		\2347_b1 , \2347_b0 , \2348_b1 , \2348_b0 , \2349_b1 , \2349_b0 , \2350_b1 , \2350_b0 , \2351_b1 , \2351_b0 , 
		\2352_b1 , \2352_b0 , \2353_b1 , \2353_b0 , \2354_b1 , \2354_b0 , \2355_b1 , \2355_b0 , \2356_b1 , \2356_b0 , 
		\2357_b1 , \2357_b0 , \2358_b1 , \2358_b0 , \2359_b1 , \2359_b0 , \2360_b1 , \2360_b0 , \2361_b1 , \2361_b0 , 
		\2362_b1 , \2362_b0 , \2363_b1 , \2363_b0 , \2364_b1 , \2364_b0 , \2365_b1 , \2365_b0 , \2366_b1 , \2366_b0 , 
		\2367_b1 , \2367_b0 , \2368_b1 , \2368_b0 , \2369_b1 , \2369_b0 , \2370_b1 , \2370_b0 , \2371_b1 , \2371_b0 , 
		\2372_b1 , \2372_b0 , \2373_b1 , \2373_b0 , \2374_b1 , \2374_b0 , \2375_b1 , \2375_b0 , \2376_b1 , \2376_b0 , 
		\2377_b1 , \2377_b0 , \2378_b1 , \2378_b0 , \2379_b1 , \2379_b0 , \2380_b1 , \2380_b0 , \2381_b1 , \2381_b0 , 
		\2382_b1 , \2382_b0 , \2383_b1 , \2383_b0 , \2384_b1 , \2384_b0 , \2385_b1 , \2385_b0 , \2386_b1 , \2386_b0 , 
		\2387_b1 , \2387_b0 , \2388_b1 , \2388_b0 , \2389_b1 , \2389_b0 , \2390_b1 , \2390_b0 , \2391_b1 , \2391_b0 , 
		\2392_b1 , \2392_b0 , \2393_b1 , \2393_b0 , \2394_b1 , \2394_b0 , \2395_b1 , \2395_b0 , \2396_b1 , \2396_b0 , 
		\2397_b1 , \2397_b0 , \2398_b1 , \2398_b0 , \2399_b1 , \2399_b0 , \2400_b1 , \2400_b0 , \2401_b1 , \2401_b0 , 
		\2402_b1 , \2402_b0 , \2403_b1 , \2403_b0 , \2404_b1 , \2404_b0 , \2405_b1 , \2405_b0 , \2406_b1 , \2406_b0 , 
		\2407_b1 , \2407_b0 , \2408_b1 , \2408_b0 , \2409_b1 , \2409_b0 , \2410_b1 , \2410_b0 , \2411_b1 , \2411_b0 , 
		\2412_b1 , \2412_b0 , \2413_b1 , \2413_b0 , \2414_b1 , \2414_b0 , \2415_b1 , \2415_b0 , \2416_b1 , \2416_b0 , 
		\2417_b1 , \2417_b0 , \2418_b1 , \2418_b0 , \2419_b1 , \2419_b0 , \2420_b1 , \2420_b0 , \2421_b1 , \2421_b0 , 
		\2422_b1 , \2422_b0 , \2423_b1 , \2423_b0 , \2424_b1 , \2424_b0 , \2425_b1 , \2425_b0 , \2426_b1 , \2426_b0 , 
		\2427_b1 , \2427_b0 , \2428_b1 , \2428_b0 , \2429_b1 , \2429_b0 , \2430_b1 , \2430_b0 , \2431_b1 , \2431_b0 , 
		\2432_b1 , \2432_b0 , \2433_b1 , \2433_b0 , \2434_b1 , \2434_b0 , \2435_b1 , \2435_b0 , \2436_b1 , \2436_b0 , 
		\2437_b1 , \2437_b0 , \2438_b1 , \2438_b0 , \2439_b1 , \2439_b0 , \2440_b1 , \2440_b0 , \2441_b1 , \2441_b0 , 
		\2442_b1 , \2442_b0 , \2443_b1 , \2443_b0 , \2444_b1 , \2444_b0 , \2445_b1 , \2445_b0 , \2446_b1 , \2446_b0 , 
		\2447_b1 , \2447_b0 , \2448_b1 , \2448_b0 , \2449_b1 , \2449_b0 , \2450_b1 , \2450_b0 , \2451_b1 , \2451_b0 , 
		\2452_b1 , \2452_b0 , \2453_b1 , \2453_b0 , \2454_b1 , \2454_b0 , \2455_b1 , \2455_b0 , \2456_b1 , \2456_b0 , 
		\2457_b1 , \2457_b0 , \2458_b1 , \2458_b0 , \2459_b1 , \2459_b0 , \2460_b1 , \2460_b0 , \2461_b1 , \2461_b0 , 
		\2462_b1 , \2462_b0 , \2463_b1 , \2463_b0 , \2464_b1 , \2464_b0 , \2465_b1 , \2465_b0 , \2466_b1 , \2466_b0 , 
		\2467_b1 , \2467_b0 , \2468_b1 , \2468_b0 , \2469_b1 , \2469_b0 , \2470_b1 , \2470_b0 , \2471_b1 , \2471_b0 , 
		\2472_b1 , \2472_b0 , \2473_b1 , \2473_b0 , \2474_b1 , \2474_b0 , \2475_b1 , \2475_b0 , \2476_b1 , \2476_b0 , 
		\2477_b1 , \2477_b0 , \2478_b1 , \2478_b0 , \2479_b1 , \2479_b0 , \2480_b1 , \2480_b0 , \2481_b1 , \2481_b0 , 
		\2482_b1 , \2482_b0 , \2483_b1 , \2483_b0 , \2484_b1 , \2484_b0 , \2485_b1 , \2485_b0 , \2486_b1 , \2486_b0 , 
		\2487_b1 , \2487_b0 , \2488_b1 , \2488_b0 , \2489_b1 , \2489_b0 , \2490_b1 , \2490_b0 , \2491_b1 , \2491_b0 , 
		\2492_b1 , \2492_b0 , \2493_b1 , \2493_b0 , \2494_b1 , \2494_b0 , \2495_b1 , \2495_b0 , \2496_b1 , \2496_b0 , 
		\2497_b1 , \2497_b0 , \2498_b1 , \2498_b0 , \2499_b1 , \2499_b0 , \2500_b1 , \2500_b0 , \2501_b1 , \2501_b0 , 
		\2502_b1 , \2502_b0 , \2503_b1 , \2503_b0 , \2504_b1 , \2504_b0 , \2505_b1 , \2505_b0 , \2506_b1 , \2506_b0 , 
		\2507_b1 , \2507_b0 , \2508_b1 , \2508_b0 , \2509_b1 , \2509_b0 , \2510_b1 , \2510_b0 , \2511_b1 , \2511_b0 , 
		\2512_b1 , \2512_b0 , \2513_b1 , \2513_b0 , \2514_b1 , \2514_b0 , \2515_b1 , \2515_b0 , \2516_b1 , \2516_b0 , 
		\2517_b1 , \2517_b0 , \2518_b1 , \2518_b0 , \2519_b1 , \2519_b0 , \2520_b1 , \2520_b0 , \2521_b1 , \2521_b0 , 
		\2522_b1 , \2522_b0 , \2523_b1 , \2523_b0 , \2524_b1 , \2524_b0 , \2525_b1 , \2525_b0 , \2526_b1 , \2526_b0 , 
		\2527_b1 , \2527_b0 , \2528_b1 , \2528_b0 , \2529_b1 , \2529_b0 , \2530_b1 , \2530_b0 , \2531_b1 , \2531_b0 , 
		\2532_b1 , \2532_b0 , \2533_b1 , \2533_b0 , \2534_b1 , \2534_b0 , \2535_b1 , \2535_b0 , \2536_b1 , \2536_b0 , 
		\2537_b1 , \2537_b0 , \2538_b1 , \2538_b0 , \2539_b1 , \2539_b0 , \2540_b1 , \2540_b0 , \2541_b1 , \2541_b0 , 
		\2542_b1 , \2542_b0 , \2543_b1 , \2543_b0 , \2544_b1 , \2544_b0 , \2545_b1 , \2545_b0 , \2546_b1 , \2546_b0 , 
		\2547_b1 , \2547_b0 , \2548_b1 , \2548_b0 , \2549_b1 , \2549_b0 , \2550_b1 , \2550_b0 , \2551_b1 , \2551_b0 , 
		\2552_b1 , \2552_b0 , \2553_b1 , \2553_b0 , \2554_b1 , \2554_b0 , \2555_b1 , \2555_b0 , \2556_b1 , \2556_b0 , 
		\2557_b1 , \2557_b0 , \2558_b1 , \2558_b0 , \2559_b1 , \2559_b0 , \2560_b1 , \2560_b0 , \2561_b1 , \2561_b0 , 
		\2562_b1 , \2562_b0 , \2563_b1 , \2563_b0 , \2564_b1 , \2564_b0 , \2565_b1 , \2565_b0 , \2566_b1 , \2566_b0 , 
		\2567_b1 , \2567_b0 , \2568_b1 , \2568_b0 , \2569_b1 , \2569_b0 , \2570_b1 , \2570_b0 , \2571_b1 , \2571_b0 , 
		\2572_b1 , \2572_b0 , \2573_b1 , \2573_b0 , \2574_b1 , \2574_b0 , \2575_b1 , \2575_b0 , \2576_b1 , \2576_b0 , 
		\2577_b1 , \2577_b0 , \2578_b1 , \2578_b0 , \2579_b1 , \2579_b0 , \2580_b1 , \2580_b0 , \2581_b1 , \2581_b0 , 
		\2582_b1 , \2582_b0 , \2583_b1 , \2583_b0 , \2584_b1 , \2584_b0 , \2585_b1 , \2585_b0 , \2586_b1 , \2586_b0 , 
		\2587_b1 , \2587_b0 , \2588_b1 , \2588_b0 , \2589_b1 , \2589_b0 , \2590_b1 , \2590_b0 , \2591_b1 , \2591_b0 , 
		\2592_b1 , \2592_b0 , \2593_b1 , \2593_b0 , \2594_b1 , \2594_b0 , \2595_b1 , \2595_b0 , \2596_b1 , \2596_b0 , 
		\2597_b1 , \2597_b0 , \2598_b1 , \2598_b0 , \2599_b1 , \2599_b0 , \2600_b1 , \2600_b0 , \2601_b1 , \2601_b0 , 
		\2602_b1 , \2602_b0 , \2603_b1 , \2603_b0 , \2604_b1 , \2604_b0 , \2605_b1 , \2605_b0 , \2606_b1 , \2606_b0 , 
		\2607_b1 , \2607_b0 , \2608_b1 , \2608_b0 , \2609_b1 , \2609_b0 , \2610_b1 , \2610_b0 , \2611_b1 , \2611_b0 , 
		\2612_b1 , \2612_b0 , \2613_b1 , \2613_b0 , \2614_b1 , \2614_b0 , \2615_b1 , \2615_b0 , \2616_b1 , \2616_b0 , 
		\2617_b1 , \2617_b0 , \2618_b1 , \2618_b0 , \2619_b1 , \2619_b0 , \2620_b1 , \2620_b0 , \2621_b1 , \2621_b0 , 
		\2622_b1 , \2622_b0 , \2623_b1 , \2623_b0 , \2624_b1 , \2624_b0 , \2625_b1 , \2625_b0 , \2626_b1 , \2626_b0 , 
		\2627_b1 , \2627_b0 , \2628_b1 , \2628_b0 , \2629_b1 , \2629_b0 , \2630_b1 , \2630_b0 , \2631_b1 , \2631_b0 , 
		\2632_b1 , \2632_b0 , \2633_b1 , \2633_b0 , \2634_b1 , \2634_b0 , \2635_b1 , \2635_b0 , \2636_b1 , \2636_b0 , 
		\2637_b1 , \2637_b0 , \2638_b1 , \2638_b0 , \2639_b1 , \2639_b0 , \2640_b1 , \2640_b0 , \2641_b1 , \2641_b0 , 
		\2642_b1 , \2642_b0 , \2643_b1 , \2643_b0 , \2644_b1 , \2644_b0 , \2645_b1 , \2645_b0 , \2646_b1 , \2646_b0 , 
		\2647_b1 , \2647_b0 , \2648_b1 , \2648_b0 , \2649_b1 , \2649_b0 , \2650_b1 , \2650_b0 , \2651_b1 , \2651_b0 , 
		\2652_b1 , \2652_b0 , \2653_b1 , \2653_b0 , \2654_b1 , \2654_b0 , \2655_b1 , \2655_b0 , \2656_b1 , \2656_b0 , 
		\2657_b1 , \2657_b0 , \2658_b1 , \2658_b0 , \2659_b1 , \2659_b0 , \2660_b1 , \2660_b0 , \2661_b1 , \2661_b0 , 
		\2662_b1 , \2662_b0 , \2663_b1 , \2663_b0 , \2664_b1 , \2664_b0 , \2665_b1 , \2665_b0 , \2666_b1 , \2666_b0 , 
		\2667_b1 , \2667_b0 , \2668_b1 , \2668_b0 , \2669_b1 , \2669_b0 , \2670_b1 , \2670_b0 , \2671_b1 , \2671_b0 , 
		\2672_b1 , \2672_b0 , \2673_b1 , \2673_b0 , \2674_b1 , \2674_b0 , \2675_b1 , \2675_b0 , \2676_b1 , \2676_b0 , 
		\2677_b1 , \2677_b0 , \2678_b1 , \2678_b0 , \2679_b1 , \2679_b0 , \2680_b1 , \2680_b0 , \2681_b1 , \2681_b0 , 
		\2682_b1 , \2682_b0 , \2683_b1 , \2683_b0 , \2684_b1 , \2684_b0 , \2685_b1 , \2685_b0 , \2686_b1 , \2686_b0 , 
		\2687_b1 , \2687_b0 , \2688_b1 , \2688_b0 , \2689_b1 , \2689_b0 , \2690_b1 , \2690_b0 , \2691_b1 , \2691_b0 , 
		\2692_b1 , \2692_b0 , \2693_b1 , \2693_b0 , \2694_b1 , \2694_b0 , \2695_b1 , \2695_b0 , \2696_b1 , \2696_b0 , 
		\2697_b1 , \2697_b0 , \2698_b1 , \2698_b0 , \2699_b1 , \2699_b0 , \2700_b1 , \2700_b0 , \2701_b1 , \2701_b0 , 
		\2702_b1 , \2702_b0 , \2703_b1 , \2703_b0 , \2704_b1 , \2704_b0 , \2705_b1 , \2705_b0 , \2706_b1 , \2706_b0 , 
		\2707_b1 , \2707_b0 , \2708_b1 , \2708_b0 , \2709_b1 , \2709_b0 , \2710_b1 , \2710_b0 , \2711_b1 , \2711_b0 , 
		\2712_b1 , \2712_b0 , \2713_b1 , \2713_b0 , \2714_b1 , \2714_b0 , \2715_b1 , \2715_b0 , \2716_b1 , \2716_b0 , 
		\2717_b1 , \2717_b0 , \2718_b1 , \2718_b0 , \2719_b1 , \2719_b0 , \2720_b1 , \2720_b0 , \2721_b1 , \2721_b0 , 
		\2722_b1 , \2722_b0 , \2723_b1 , \2723_b0 , \2724_b1 , \2724_b0 , \2725_b1 , \2725_b0 , \2726_b1 , \2726_b0 , 
		\2727_b1 , \2727_b0 , \2728_b1 , \2728_b0 , \2729_b1 , \2729_b0 , \2730_b1 , \2730_b0 , \2731_b1 , \2731_b0 , 
		\2732_b1 , \2732_b0 , \2733_b1 , \2733_b0 , \2734_b1 , \2734_b0 , \2735_b1 , \2735_b0 , \2736_b1 , \2736_b0 , 
		\2737_b1 , \2737_b0 , \2738_b1 , \2738_b0 , \2739_b1 , \2739_b0 , \2740_b1 , \2740_b0 , \2741_b1 , \2741_b0 , 
		\2742_b1 , \2742_b0 , \2743_b1 , \2743_b0 , \2744_b1 , \2744_b0 , \2745_b1 , \2745_b0 , \2746_b1 , \2746_b0 , 
		\2747_b1 , \2747_b0 , \2748_b1 , \2748_b0 , \2749_b1 , \2749_b0 , \2750_b1 , \2750_b0 , \2751_b1 , \2751_b0 , 
		\2752_b1 , \2752_b0 , \2753_b1 , \2753_b0 , \2754_b1 , \2754_b0 , \2755_b1 , \2755_b0 , \2756_b1 , \2756_b0 , 
		\2757_b1 , \2757_b0 , \2758_b1 , \2758_b0 , \2759_b1 , \2759_b0 , \2760_b1 , \2760_b0 , \2761_b1 , \2761_b0 , 
		\2762_b1 , \2762_b0 , \2763_b1 , \2763_b0 , \2764_b1 , \2764_b0 , \2765_b1 , \2765_b0 , \2766_b1 , \2766_b0 , 
		\2767_b1 , \2767_b0 , \2768_b1 , \2768_b0 , \2769_b1 , \2769_b0 , \2770_b1 , \2770_b0 , \2771_b1 , \2771_b0 , 
		\2772_b1 , \2772_b0 , \2773_b1 , \2773_b0 , \2774_b1 , \2774_b0 , \2775_b1 , \2775_b0 , \2776_b1 , \2776_b0 , 
		\2777_b1 , \2777_b0 , \2778_b1 , \2778_b0 , \2779_b1 , \2779_b0 , \2780_b1 , \2780_b0 , \2781_b1 , \2781_b0 , 
		\2782_b1 , \2782_b0 , \2783_b1 , \2783_b0 , \2784_b1 , \2784_b0 , \2785_b1 , \2785_b0 , \2786_b1 , \2786_b0 , 
		\2787_b1 , \2787_b0 , \2788_b1 , \2788_b0 , \2789_b1 , \2789_b0 , \2790_b1 , \2790_b0 , \2791_b1 , \2791_b0 , 
		\2792_b1 , \2792_b0 , \2793_b1 , \2793_b0 , \2794_b1 , \2794_b0 , \2795_b1 , \2795_b0 , \2796_b1 , \2796_b0 , 
		\2797_b1 , \2797_b0 , \2798_b1 , \2798_b0 , \2799_b1 , \2799_b0 , \2800_b1 , \2800_b0 , \2801_b1 , \2801_b0 , 
		\2802_b1 , \2802_b0 , \2803_b1 , \2803_b0 , \2804_b1 , \2804_b0 , \2805_b1 , \2805_b0 , \2806_b1 , \2806_b0 , 
		\2807_b1 , \2807_b0 , \2808_b1 , \2808_b0 , \2809_b1 , \2809_b0 , \2810_b1 , \2810_b0 , \2811_b1 , \2811_b0 , 
		\2812_b1 , \2812_b0 , \2813_b1 , \2813_b0 , \2814_b1 , \2814_b0 , \2815_b1 , \2815_b0 , \2816_b1 , \2816_b0 , 
		\2817_b1 , \2817_b0 , \2818_b1 , \2818_b0 , \2819_b1 , \2819_b0 , \2820_b1 , \2820_b0 , \2821_b1 , \2821_b0 , 
		\2822_b1 , \2822_b0 , \2823_b1 , \2823_b0 , \2824_b1 , \2824_b0 , \2825_b1 , \2825_b0 , \2826_b1 , \2826_b0 , 
		\2827_b1 , \2827_b0 , \2828_b1 , \2828_b0 , \2829_b1 , \2829_b0 , \2830_b1 , \2830_b0 , \2831_b1 , \2831_b0 , 
		\2832_b1 , \2832_b0 , \2833_b1 , \2833_b0 , \2834_b1 , \2834_b0 , \2835_b1 , \2835_b0 , \2836_b1 , \2836_b0 , 
		\2837_b1 , \2837_b0 , \2838_b1 , \2838_b0 , \2839_b1 , \2839_b0 , \2840_b1 , \2840_b0 , \2841_b1 , \2841_b0 , 
		\2842_b1 , \2842_b0 , \2843_b1 , \2843_b0 , \2844_b1 , \2844_b0 , \2845_b1 , \2845_b0 , \2846_b1 , \2846_b0 , 
		\2847_b1 , \2847_b0 , \2848_b1 , \2848_b0 , \2849_b1 , \2849_b0 , \2850_b1 , \2850_b0 , \2851_b1 , \2851_b0 , 
		\2852_b1 , \2852_b0 , \2853_b1 , \2853_b0 , \2854_b1 , \2854_b0 , \2855_b1 , \2855_b0 , \2856_b1 , \2856_b0 , 
		\2857_b1 , \2857_b0 , \2858_b1 , \2858_b0 , \2859_b1 , \2859_b0 , \2860_b1 , \2860_b0 , \2861_b1 , \2861_b0 , 
		\2862_b1 , \2862_b0 , \2863_b1 , \2863_b0 , \2864_b1 , \2864_b0 , \2865_b1 , \2865_b0 , \2866_b1 , \2866_b0 , 
		\2867_b1 , \2867_b0 , \2868_b1 , \2868_b0 , \2869_b1 , \2869_b0 , \2870_b1 , \2870_b0 , \2871_b1 , \2871_b0 , 
		\2872_b1 , \2872_b0 , \2873_b1 , \2873_b0 , \2874_b1 , \2874_b0 , \2875_b1 , \2875_b0 , \2876_b1 , \2876_b0 , 
		\2877_b1 , \2877_b0 , \2878_b1 , \2878_b0 , \2879_b1 , \2879_b0 , \2880_b1 , \2880_b0 , \2881_b1 , \2881_b0 , 
		\2882_b1 , \2882_b0 , \2883_b1 , \2883_b0 , \2884_b1 , \2884_b0 , \2885_b1 , \2885_b0 , \2886_b1 , \2886_b0 , 
		\2887_b1 , \2887_b0 , \2888_b1 , \2888_b0 , \2889_b1 , \2889_b0 , \2890_b1 , \2890_b0 , \2891_b1 , \2891_b0 , 
		\2892_b1 , \2892_b0 , \2893_b1 , \2893_b0 , \2894_b1 , \2894_b0 , \2895_b1 , \2895_b0 , \2896_b1 , \2896_b0 , 
		\2897_b1 , \2897_b0 , \2898_b1 , \2898_b0 , \2899_b1 , \2899_b0 , \2900_b1 , \2900_b0 , \2901_b1 , \2901_b0 , 
		\2902_b1 , \2902_b0 , \2903_b1 , \2903_b0 , \2904_b1 , \2904_b0 , \2905_b1 , \2905_b0 , \2906_b1 , \2906_b0 , 
		\2907_b1 , \2907_b0 , \2908_b1 , \2908_b0 , \2909_b1 , \2909_b0 , \2910_b1 , \2910_b0 , \2911_b1 , \2911_b0 , 
		\2912_b1 , \2912_b0 , \2913_b1 , \2913_b0 , \2914_b1 , \2914_b0 , \2915_b1 , \2915_b0 , \2916_b1 , \2916_b0 , 
		\2917_b1 , \2917_b0 , \2918_b1 , \2918_b0 , \2919_b1 , \2919_b0 , \2920_b1 , \2920_b0 , \2921_b1 , \2921_b0 , 
		\2922_b1 , \2922_b0 , \2923_b1 , \2923_b0 , \2924_b1 , \2924_b0 , \2925_b1 , \2925_b0 , \2926_b1 , \2926_b0 , 
		\2927_b1 , \2927_b0 , \2928_b1 , \2928_b0 , \2929_b1 , \2929_b0 , \2930_b1 , \2930_b0 , \2931_b1 , \2931_b0 , 
		\2932_b1 , \2932_b0 , \2933_b1 , \2933_b0 , \2934_b1 , \2934_b0 , \2935_b1 , \2935_b0 , \2936_b1 , \2936_b0 , 
		\2937_b1 , \2937_b0 , \2938_b1 , \2938_b0 , \2939_b1 , \2939_b0 , \2940_b1 , \2940_b0 , \2941_b1 , \2941_b0 , 
		\2942_b1 , \2942_b0 , \2943_b1 , \2943_b0 , \2944_b1 , \2944_b0 , \2945_b1 , \2945_b0 , \2946_b1 , \2946_b0 , 
		\2947_b1 , \2947_b0 , \2948_b1 , \2948_b0 , \2949_b1 , \2949_b0 , \2950_b1 , \2950_b0 , \2951_b1 , \2951_b0 , 
		\2952_b1 , \2952_b0 , \2953_b1 , \2953_b0 , \2954_b1 , \2954_b0 , \2955_b1 , \2955_b0 , \2956_b1 , \2956_b0 , 
		\2957_b1 , \2957_b0 , \2958_b1 , \2958_b0 , \2959_b1 , \2959_b0 , \2960_b1 , \2960_b0 , \2961_b1 , \2961_b0 , 
		\2962_b1 , \2962_b0 , \2963_b1 , \2963_b0 , \2964_b1 , \2964_b0 , \2965_b1 , \2965_b0 , \2966_b1 , \2966_b0 , 
		\2967_b1 , \2967_b0 , \2968_b1 , \2968_b0 , \2969_b1 , \2969_b0 , \2970_b1 , \2970_b0 , \2971_b1 , \2971_b0 , 
		\2972_b1 , \2972_b0 , \2973_b1 , \2973_b0 , \2974_b1 , \2974_b0 , \2975_b1 , \2975_b0 , \2976_b1 , \2976_b0 , 
		\2977_b1 , \2977_b0 , \2978_b1 , \2978_b0 , \2979_b1 , \2979_b0 , \2980_b1 , \2980_b0 , \2981_b1 , \2981_b0 , 
		\2982_b1 , \2982_b0 , \2983_b1 , \2983_b0 , \2984_b1 , \2984_b0 , \2985_b1 , \2985_b0 , \2986_b1 , \2986_b0 , 
		\2987_b1 , \2987_b0 , \2988_b1 , \2988_b0 , \2989_b1 , \2989_b0 , \2990_b1 , \2990_b0 , \2991_b1 , \2991_b0 , 
		\2992_b1 , \2992_b0 , \2993_b1 , \2993_b0 , \2994_b1 , \2994_b0 , \2995_b1 , \2995_b0 , \2996_b1 , \2996_b0 , 
		\2997_b1 , \2997_b0 , \2998_b1 , \2998_b0 , \2999_b1 , \2999_b0 , \3000_b1 , \3000_b0 , \3001_b1 , \3001_b0 , 
		\3002_b1 , \3002_b0 , \3003_b1 , \3003_b0 , \3004_b1 , \3004_b0 , \3005_b1 , \3005_b0 , \3006_b1 , \3006_b0 , 
		\3007_b1 , \3007_b0 , \3008_b1 , \3008_b0 , \3009_b1 , \3009_b0 , \3010_b1 , \3010_b0 , \3011_b1 , \3011_b0 , 
		\3012_b1 , \3012_b0 , \3013_b1 , \3013_b0 , \3014_b1 , \3014_b0 , \3015_b1 , \3015_b0 , \3016_b1 , \3016_b0 , 
		\3017_b1 , \3017_b0 , \3018_b1 , \3018_b0 , \3019_b1 , \3019_b0 , \3020_b1 , \3020_b0 , \3021_b1 , \3021_b0 , 
		\3022_b1 , \3022_b0 , \3023_b1 , \3023_b0 , \3024_b1 , \3024_b0 , \3025_b1 , \3025_b0 , \3026_b1 , \3026_b0 , 
		\3027_b1 , \3027_b0 , \3028_b1 , \3028_b0 , \3029_b1 , \3029_b0 , \3030_b1 , \3030_b0 , \3031_b1 , \3031_b0 , 
		\3032_b1 , \3032_b0 , \3033_b1 , \3033_b0 , \3034_b1 , \3034_b0 , \3035_b1 , \3035_b0 , \3036_b1 , \3036_b0 , 
		\3037_b1 , \3037_b0 , \3038_b1 , \3038_b0 , \3039_b1 , \3039_b0 , \3040_b1 , \3040_b0 , \3041_b1 , \3041_b0 , 
		\3042_b1 , \3042_b0 , \3043_b1 , \3043_b0 , \3044_b1 , \3044_b0 , \3045_b1 , \3045_b0 , \3046_b1 , \3046_b0 , 
		\3047_b1 , \3047_b0 , \3048_b1 , \3048_b0 , \3049_b1 , \3049_b0 , \3050_b1 , \3050_b0 , \3051_b1 , \3051_b0 , 
		\3052_b1 , \3052_b0 , \3053_b1 , \3053_b0 , \3054_b1 , \3054_b0 , \3055_b1 , \3055_b0 , \3056_b1 , \3056_b0 , 
		\3057_b1 , \3057_b0 , \3058_b1 , \3058_b0 , \3059_b1 , \3059_b0 , \3060_b1 , \3060_b0 , \3061_b1 , \3061_b0 , 
		\3062_b1 , \3062_b0 , \3063_b1 , \3063_b0 , \3064_b1 , \3064_b0 , \3065_b1 , \3065_b0 , \3066_b1 , \3066_b0 , 
		\3067_b1 , \3067_b0 , \3068_b1 , \3068_b0 , \3069_b1 , \3069_b0 , \3070_b1 , \3070_b0 , \3071_b1 , \3071_b0 , 
		\3072_b1 , \3072_b0 , \3073_b1 , \3073_b0 , \3074_b1 , \3074_b0 , \3075_b1 , \3075_b0 , \3076_b1 , \3076_b0 , 
		\3077_b1 , \3077_b0 , \3078_b1 , \3078_b0 , \3079_b1 , \3079_b0 , \3080_b1 , \3080_b0 , \3081_b1 , \3081_b0 , 
		\3082_b1 , \3082_b0 , \3083_b1 , \3083_b0 , \3084_b1 , \3084_b0 , \3085_b1 , \3085_b0 , \3086_b1 , \3086_b0 , 
		\3087_b1 , \3087_b0 , \3088_b1 , \3088_b0 , \3089_b1 , \3089_b0 , \3090_b1 , \3090_b0 , \3091_b1 , \3091_b0 , 
		\3092_b1 , \3092_b0 , \3093_b1 , \3093_b0 , \3094_b1 , \3094_b0 , \3095_b1 , \3095_b0 , \3096_b1 , \3096_b0 , 
		\3097_b1 , \3097_b0 , \3098_b1 , \3098_b0 , \3099_b1 , \3099_b0 , \3100_b1 , \3100_b0 , \3101_b1 , \3101_b0 , 
		\3102_b1 , \3102_b0 , \3103_b1 , \3103_b0 , \3104_b1 , \3104_b0 , \3105_b1 , \3105_b0 , \3106_b1 , \3106_b0 , 
		\3107_b1 , \3107_b0 , \3108_b1 , \3108_b0 , \3109_b1 , \3109_b0 , \3110_b1 , \3110_b0 , \3111_b1 , \3111_b0 , 
		\3112_b1 , \3112_b0 , \3113_b1 , \3113_b0 , \3114_b1 , \3114_b0 , \3115_b1 , \3115_b0 , \3116_b1 , \3116_b0 , 
		\3117_b1 , \3117_b0 , \3118_b1 , \3118_b0 , \3119_b1 , \3119_b0 , \3120_b1 , \3120_b0 , \3121_b1 , \3121_b0 , 
		\3122_b1 , \3122_b0 , \3123_b1 , \3123_b0 , \3124_b1 , \3124_b0 , \3125_b1 , \3125_b0 , \3126_b1 , \3126_b0 , 
		\3127_b1 , \3127_b0 , \3128_b1 , \3128_b0 , \3129_b1 , \3129_b0 , \3130_b1 , \3130_b0 , \3131_b1 , \3131_b0 , 
		\3132_b1 , \3132_b0 , \3133_b1 , \3133_b0 , \3134_b1 , \3134_b0 , \3135_b1 , \3135_b0 , \3136_b1 , \3136_b0 , 
		\3137_b1 , \3137_b0 , \3138_b1 , \3138_b0 , \3139_b1 , \3139_b0 , \3140_b1 , \3140_b0 , \3141_b1 , \3141_b0 , 
		\3142_b1 , \3142_b0 , \3143_b1 , \3143_b0 , \3144_b1 , \3144_b0 , \3145_b1 , \3145_b0 , \3146_b1 , \3146_b0 , 
		\3147_b1 , \3147_b0 , \3148_b1 , \3148_b0 , \3149_b1 , \3149_b0 , \3150_b1 , \3150_b0 , \3151_b1 , \3151_b0 , 
		\3152_b1 , \3152_b0 , \3153_b1 , \3153_b0 , \3154_b1 , \3154_b0 , \3155_b1 , \3155_b0 , \3156_b1 , \3156_b0 , 
		\3157_b1 , \3157_b0 , \3158_b1 , \3158_b0 , \3159_b1 , \3159_b0 , \3160_b1 , \3160_b0 , \3161_b1 , \3161_b0 , 
		\3162_b1 , \3162_b0 , \3163_b1 , \3163_b0 , \3164_b1 , \3164_b0 , \3165_b1 , \3165_b0 , \3166_b1 , \3166_b0 , 
		\3167_b1 , \3167_b0 , \3168_b1 , \3168_b0 , \3169_b1 , \3169_b0 , \3170_b1 , \3170_b0 , \3171_b1 , \3171_b0 , 
		\3172_b1 , \3172_b0 , \3173_b1 , \3173_b0 , \3174_b1 , \3174_b0 , \3175_b1 , \3175_b0 , \3176_b1 , \3176_b0 , 
		\3177_b1 , \3177_b0 , \3178_b1 , \3178_b0 , \3179_b1 , \3179_b0 , \3180_b1 , \3180_b0 , \3181_b1 , \3181_b0 , 
		\3182_b1 , \3182_b0 , \3183_b1 , \3183_b0 , \3184_b1 , \3184_b0 , \3185_b1 , \3185_b0 , \3186_b1 , \3186_b0 , 
		\3187_b1 , \3187_b0 , \3188_b1 , \3188_b0 , \3189_b1 , \3189_b0 , \3190_b1 , \3190_b0 , \3191_b1 , \3191_b0 , 
		\3192_b1 , \3192_b0 , \3193_b1 , \3193_b0 , \3194_b1 , \3194_b0 , \3195_b1 , \3195_b0 , \3196_b1 , \3196_b0 , 
		\3197_b1 , \3197_b0 , \3198_b1 , \3198_b0 , \3199_b1 , \3199_b0 , \3200_b1 , \3200_b0 , \3201_b1 , \3201_b0 , 
		\3202_b1 , \3202_b0 , \3203_b1 , \3203_b0 , \3204_b1 , \3204_b0 , \3205_b1 , \3205_b0 , \3206_b1 , \3206_b0 , 
		\3207_b1 , \3207_b0 , \3208_b1 , \3208_b0 , \3209_b1 , \3209_b0 , \3210_b1 , \3210_b0 , \3211_b1 , \3211_b0 , 
		\3212_b1 , \3212_b0 , \3213_b1 , \3213_b0 , \3214_b1 , \3214_b0 , \3215_b1 , \3215_b0 , \3216_b1 , \3216_b0 , 
		\3217_b1 , \3217_b0 , \3218_b1 , \3218_b0 , \3219_b1 , \3219_b0 , \3220_b1 , \3220_b0 , \3221_b1 , \3221_b0 , 
		\3222_b1 , \3222_b0 , \3223_b1 , \3223_b0 , \3224_b1 , \3224_b0 , \3225_b1 , \3225_b0 , \3226_b1 , \3226_b0 , 
		\3227_b1 , \3227_b0 , \3228_b1 , \3228_b0 , \3229_b1 , \3229_b0 , \3230_b1 , \3230_b0 , \3231_b1 , \3231_b0 , 
		\3232_b1 , \3232_b0 , \3233_b1 , \3233_b0 , \3234_b1 , \3234_b0 , \3235_b1 , \3235_b0 , \3236_b1 , \3236_b0 , 
		\3237_b1 , \3237_b0 , \3238_b1 , \3238_b0 , \3239_b1 , \3239_b0 , \3240_b1 , \3240_b0 , \3241_b1 , \3241_b0 , 
		\3242_b1 , \3242_b0 , \3243_b1 , \3243_b0 , \3244_b1 , \3244_b0 , \3245_b1 , \3245_b0 , \3246_b1 , \3246_b0 , 
		\3247_b1 , \3247_b0 , \3248_b1 , \3248_b0 , \3249_b1 , \3249_b0 , \3250_b1 , \3250_b0 , \3251_b1 , \3251_b0 , 
		\3252_b1 , \3252_b0 , \3253_b1 , \3253_b0 , \3254_b1 , \3254_b0 , \3255_b1 , \3255_b0 , \3256_b1 , \3256_b0 , 
		\3257_b1 , \3257_b0 , \3258_b1 , \3258_b0 , \3259_b1 , \3259_b0 , \3260_b1 , \3260_b0 , \3261_b1 , \3261_b0 , 
		\3262_b1 , \3262_b0 , \3263_b1 , \3263_b0 , \3264_b1 , \3264_b0 , \3265_b1 , \3265_b0 , \3266_b1 , \3266_b0 , 
		\3267_b1 , \3267_b0 , \3268_b1 , \3268_b0 , \3269_b1 , \3269_b0 , \3270_b1 , \3270_b0 , \3271_b1 , \3271_b0 , 
		\3272_b1 , \3272_b0 , \3273_b1 , \3273_b0 , \3274_b1 , \3274_b0 , \3275_b1 , \3275_b0 , \3276_b1 , \3276_b0 , 
		\3277_b1 , \3277_b0 , \3278_b1 , \3278_b0 , \3279_b1 , \3279_b0 , \3280_b1 , \3280_b0 , \3281_b1 , \3281_b0 , 
		\3282_b1 , \3282_b0 , \3283_b1 , \3283_b0 , \3284_b1 , \3284_b0 , \3285_b1 , \3285_b0 , \3286_b1 , \3286_b0 , 
		\3287_b1 , \3287_b0 , \3288_b1 , \3288_b0 , \3289_b1 , \3289_b0 , \3290_b1 , \3290_b0 , \3291_b1 , \3291_b0 , 
		\3292_b1 , \3292_b0 , \3293_b1 , \3293_b0 , \3294_b1 , \3294_b0 , \3295_b1 , \3295_b0 , \3296_b1 , \3296_b0 , 
		\3297_b1 , \3297_b0 , \3298_b1 , \3298_b0 , \3299_b1 , \3299_b0 , \3300_b1 , \3300_b0 , \3301_b1 , \3301_b0 , 
		\3302_b1 , \3302_b0 , \3303_b1 , \3303_b0 , \3304_b1 , \3304_b0 , \3305_b1 , \3305_b0 , \3306_b1 , \3306_b0 , 
		\3307_b1 , \3307_b0 , \3308_b1 , \3308_b0 , \3309_b1 , \3309_b0 , \3310_b1 , \3310_b0 , \3311_b1 , \3311_b0 , 
		\3312_b1 , \3312_b0 , \3313_b1 , \3313_b0 , \3314_b1 , \3314_b0 , \3315_b1 , \3315_b0 , \3316_b1 , \3316_b0 , 
		\3317_b1 , \3317_b0 , \3318_b1 , \3318_b0 , \3319_b1 , \3319_b0 , \3320_b1 , \3320_b0 , \3321_b1 , \3321_b0 , 
		\3322_b1 , \3322_b0 , \3323_b1 , \3323_b0 , \3324_b1 , \3324_b0 , \3325_b1 , \3325_b0 , \3326_b1 , \3326_b0 , 
		\3327_b1 , \3327_b0 , \3328_b1 , \3328_b0 , \3329_b1 , \3329_b0 , \3330_b1 , \3330_b0 , \3331_b1 , \3331_b0 , 
		\3332_b1 , \3332_b0 , \3333_b1 , \3333_b0 , \3334_b1 , \3334_b0 , \3335_b1 , \3335_b0 , \3336_b1 , \3336_b0 , 
		\3337_b1 , \3337_b0 , \3338_b1 , \3338_b0 , \3339_b1 , \3339_b0 , \3340_b1 , \3340_b0 , \3341_b1 , \3341_b0 , 
		\3342_b1 , \3342_b0 , \3343_b1 , \3343_b0 , \3344_b1 , \3344_b0 , \3345_b1 , \3345_b0 , \3346_b1 , \3346_b0 , 
		\3347_b1 , \3347_b0 , \3348_b1 , \3348_b0 , \3349_b1 , \3349_b0 , \3350_b1 , \3350_b0 , \3351_b1 , \3351_b0 , 
		\3352_b1 , \3352_b0 , \3353_b1 , \3353_b0 , \3354_b1 , \3354_b0 , \3355_b1 , \3355_b0 , \3356_b1 , \3356_b0 , 
		\3357_b1 , \3357_b0 , \3358_b1 , \3358_b0 , \3359_b1 , \3359_b0 , \3360_b1 , \3360_b0 , \3361_b1 , \3361_b0 , 
		\3362_b1 , \3362_b0 , \3363_b1 , \3363_b0 , \3364_b1 , \3364_b0 , \3365_b1 , \3365_b0 , \3366_b1 , \3366_b0 , 
		\3367_b1 , \3367_b0 , \3368_b1 , \3368_b0 , \3369_b1 , \3369_b0 , \3370_b1 , \3370_b0 , \3371_b1 , \3371_b0 , 
		\3372_b1 , \3372_b0 , \3373_b1 , \3373_b0 , \3374_b1 , \3374_b0 , \3375_b1 , \3375_b0 , \3376_b1 , \3376_b0 , 
		\3377_b1 , \3377_b0 , \3378_b1 , \3378_b0 , \3379_b1 , \3379_b0 , \3380_b1 , \3380_b0 , \3381_b1 , \3381_b0 , 
		\3382_b1 , \3382_b0 , \3383_b1 , \3383_b0 , \3384_b1 , \3384_b0 , \3385_b1 , \3385_b0 , \3386_b1 , \3386_b0 , 
		\3387_b1 , \3387_b0 , \3388_b1 , \3388_b0 , \3389_b1 , \3389_b0 , \3390_b1 , \3390_b0 , \3391_b1 , \3391_b0 , 
		\3392_b1 , \3392_b0 , \3393_b1 , \3393_b0 , \3394_b1 , \3394_b0 , \3395_b1 , \3395_b0 , \3396_b1 , \3396_b0 , 
		\3397_b1 , \3397_b0 , \3398_b1 , \3398_b0 , \3399_b1 , \3399_b0 , \3400_b1 , \3400_b0 , \3401_b1 , \3401_b0 , 
		\3402_b1 , \3402_b0 , \3403_b1 , \3403_b0 , \3404_b1 , \3404_b0 , \3405_b1 , \3405_b0 , \3406_b1 , \3406_b0 , 
		\3407_b1 , \3407_b0 , \3408_b1 , \3408_b0 , \3409_b1 , \3409_b0 , \3410_b1 , \3410_b0 , \3411_b1 , \3411_b0 , 
		\3412_b1 , \3412_b0 , \3413_b1 , \3413_b0 , \3414_b1 , \3414_b0 , \3415_b1 , \3415_b0 , \3416_b1 , \3416_b0 , 
		\3417_b1 , \3417_b0 , \3418_b1 , \3418_b0 , \3419_b1 , \3419_b0 , \3420_b1 , \3420_b0 , \3421_b1 , \3421_b0 , 
		\3422_b1 , \3422_b0 , \3423_b1 , \3423_b0 , \3424_b1 , \3424_b0 , \3425_b1 , \3425_b0 , \3426_b1 , \3426_b0 , 
		\3427_b1 , \3427_b0 , \3428_b1 , \3428_b0 , \3429_b1 , \3429_b0 , \3430_b1 , \3430_b0 , \3431_b1 , \3431_b0 , 
		\3432_b1 , \3432_b0 , \3433_b1 , \3433_b0 , \3434_b1 , \3434_b0 , \3435_b1 , \3435_b0 , \3436_b1 , \3436_b0 , 
		\3437_b1 , \3437_b0 , \3438_b1 , \3438_b0 , \3439_b1 , \3439_b0 , \3440_b1 , \3440_b0 , \3441_b1 , \3441_b0 , 
		\3442_b1 , \3442_b0 , \3443_b1 , \3443_b0 , \3444_b1 , \3444_b0 , \3445_b1 , \3445_b0 , \3446_b1 , \3446_b0 , 
		\3447_b1 , \3447_b0 , \3448_b1 , \3448_b0 , \3449_b1 , \3449_b0 , \3450_b1 , \3450_b0 , \3451_b1 , \3451_b0 , 
		\3452_b1 , \3452_b0 , \3453_b1 , \3453_b0 , \3454_b1 , \3454_b0 , \3455_b1 , \3455_b0 , \3456_b1 , \3456_b0 , 
		\3457_b1 , \3457_b0 , \3458_b1 , \3458_b0 , \3459_b1 , \3459_b0 , \3460_b1 , \3460_b0 , \3461_b1 , \3461_b0 , 
		\3462_b1 , \3462_b0 , \3463_b1 , \3463_b0 , \3464_b1 , \3464_b0 , \3465_b1 , \3465_b0 , \3466_b1 , \3466_b0 , 
		\3467_b1 , \3467_b0 , \3468_b1 , \3468_b0 , \3469_b1 , \3469_b0 , \3470_b1 , \3470_b0 , \3471_b1 , \3471_b0 , 
		\3472_b1 , \3472_b0 , \3473_b1 , \3473_b0 , \3474_b1 , \3474_b0 , \3475_b1 , \3475_b0 , \3476_b1 , \3476_b0 , 
		\3477_b1 , \3477_b0 , \3478_b1 , \3478_b0 , \3479_b1 , \3479_b0 , \3480_b1 , \3480_b0 , \3481_b1 , \3481_b0 , 
		\3482_b1 , \3482_b0 , \3483_b1 , \3483_b0 , \3484_b1 , \3484_b0 , \3485_b1 , \3485_b0 , \3486_b1 , \3486_b0 , 
		\3487_b1 , \3487_b0 , \3488_b1 , \3488_b0 , \3489_b1 , \3489_b0 , \3490_b1 , \3490_b0 , \3491_b1 , \3491_b0 , 
		\3492_b1 , \3492_b0 , \3493_b1 , \3493_b0 , \3494_b1 , \3494_b0 , \3495_b1 , \3495_b0 , \3496_b1 , \3496_b0 , 
		\3497_b1 , \3497_b0 , \3498_b1 , \3498_b0 , \3499_b1 , \3499_b0 , \3500_b1 , \3500_b0 , \3501_b1 , \3501_b0 , 
		\3502_b1 , \3502_b0 , \3503_b1 , \3503_b0 , \3504_b1 , \3504_b0 , \3505_b1 , \3505_b0 , \3506_b1 , \3506_b0 , 
		\3507_b1 , \3507_b0 , \3508_b1 , \3508_b0 , \3509_b1 , \3509_b0 , \3510_b1 , \3510_b0 , \3511_b1 , \3511_b0 , 
		\3512_b1 , \3512_b0 , \3513_b1 , \3513_b0 , \3514_b1 , \3514_b0 , \3515_b1 , \3515_b0 , \3516_b1 , \3516_b0 , 
		\3517_b1 , \3517_b0 , \3518_b1 , \3518_b0 , \3519_b1 , \3519_b0 , \3520_b1 , \3520_b0 , \3521_b1 , \3521_b0 , 
		\3522_b1 , \3522_b0 , \3523_b1 , \3523_b0 , \3524_b1 , \3524_b0 , \3525_b1 , \3525_b0 , \3526_b1 , \3526_b0 , 
		\3527_b1 , \3527_b0 , \3528_b1 , \3528_b0 , \3529_b1 , \3529_b0 , \3530_b1 , \3530_b0 , \3531_b1 , \3531_b0 , 
		\3532_b1 , \3532_b0 , \3533_b1 , \3533_b0 , \3534_b1 , \3534_b0 , \3535_b1 , \3535_b0 , \3536_b1 , \3536_b0 , 
		\3537_b1 , \3537_b0 , \3538_b1 , \3538_b0 , \3539_b1 , \3539_b0 , \3540_b1 , \3540_b0 , \3541_b1 , \3541_b0 , 
		\3542_b1 , \3542_b0 , \3543_b1 , \3543_b0 , \3544_b1 , \3544_b0 , \3545_b1 , \3545_b0 , \3546_b1 , \3546_b0 , 
		\3547_b1 , \3547_b0 , \3548_b1 , \3548_b0 , \3549_b1 , \3549_b0 , \3550_b1 , \3550_b0 , \3551_b1 , \3551_b0 , 
		\3552_b1 , \3552_b0 , \3553_b1 , \3553_b0 , \3554_b1 , \3554_b0 , \3555_b1 , \3555_b0 , \3556_b1 , \3556_b0 , 
		\3557_b1 , \3557_b0 , \3558_b1 , \3558_b0 , \3559_b1 , \3559_b0 , \3560_b1 , \3560_b0 , \3561_b1 , \3561_b0 , 
		\3562_b1 , \3562_b0 , \3563_b1 , \3563_b0 , \3564_b1 , \3564_b0 , \3565_b1 , \3565_b0 , \3566_b1 , \3566_b0 , 
		\3567_b1 , \3567_b0 , \3568_b1 , \3568_b0 , \3569_b1 , \3569_b0 , \3570_b1 , \3570_b0 , \3571_b1 , \3571_b0 , 
		\3572_b1 , \3572_b0 , \3573_b1 , \3573_b0 , \3574_b1 , \3574_b0 , \3575_b1 , \3575_b0 , \3576_b1 , \3576_b0 , 
		\3577_b1 , \3577_b0 , \3578_b1 , \3578_b0 , \3579_b1 , \3579_b0 , \3580_b1 , \3580_b0 , \3581_b1 , \3581_b0 , 
		\3582_b1 , \3582_b0 , \3583_b1 , \3583_b0 , \3584_b1 , \3584_b0 , \3585_b1 , \3585_b0 , \3586_b1 , \3586_b0 , 
		\3587_b1 , \3587_b0 , \3588_b1 , \3588_b0 , \3589_b1 , \3589_b0 , \3590_b1 , \3590_b0 , \3591_b1 , \3591_b0 , 
		\3592_b1 , \3592_b0 , \3593_b1 , \3593_b0 , \3594_b1 , \3594_b0 , \3595_b1 , \3595_b0 , \3596_b1 , \3596_b0 , 
		\3597_b1 , \3597_b0 , \3598_b1 , \3598_b0 , \3599_b1 , \3599_b0 , \3600_b1 , \3600_b0 , \3601_b1 , \3601_b0 , 
		\3602_b1 , \3602_b0 , \3603_b1 , \3603_b0 , \3604_b1 , \3604_b0 , \3605_b1 , \3605_b0 , \3606_b1 , \3606_b0 , 
		\3607_b1 , \3607_b0 , \3608_b1 , \3608_b0 , \3609_b1 , \3609_b0 , \3610_b1 , \3610_b0 , \3611_b1 , \3611_b0 , 
		\3612_b1 , \3612_b0 , \3613_b1 , \3613_b0 , \3614_b1 , \3614_b0 , \3615_b1 , \3615_b0 , \3616_b1 , \3616_b0 , 
		\3617_b1 , \3617_b0 , \3618_b1 , \3618_b0 , \3619_b1 , \3619_b0 , \3620_b1 , \3620_b0 , \3621_b1 , \3621_b0 , 
		\3622_b1 , \3622_b0 , \3623_b1 , \3623_b0 , \3624_b1 , \3624_b0 , \3625_b1 , \3625_b0 , \3626_b1 , \3626_b0 , 
		\3627_b1 , \3627_b0 , \3628_b1 , \3628_b0 , \3629_b1 , \3629_b0 , \3630_b1 , \3630_b0 , \3631_b1 , \3631_b0 , 
		\3632_b1 , \3632_b0 , \3633_b1 , \3633_b0 , \3634_b1 , \3634_b0 , \3635_b1 , \3635_b0 , \3636_b1 , \3636_b0 , 
		\3637_b1 , \3637_b0 , \3638_b1 , \3638_b0 , \3639_b1 , \3639_b0 , \3640_b1 , \3640_b0 , \3641_b1 , \3641_b0 , 
		\3642_b1 , \3642_b0 , \3643_b1 , \3643_b0 , \3644_b1 , \3644_b0 , \3645_b1 , \3645_b0 , \3646_b1 , \3646_b0 , 
		\3647_b1 , \3647_b0 , \3648_b1 , \3648_b0 , \3649_b1 , \3649_b0 , \3650_b1 , \3650_b0 , \3651_b1 , \3651_b0 , 
		\3652_b1 , \3652_b0 , \3653_b1 , \3653_b0 , \3654_b1 , \3654_b0 , \3655_b1 , \3655_b0 , \3656_b1 , \3656_b0 , 
		\3657_b1 , \3657_b0 , \3658_b1 , \3658_b0 , \3659_b1 , \3659_b0 , \3660_b1 , \3660_b0 , \3661_b1 , \3661_b0 , 
		\3662_b1 , \3662_b0 , \3663_b1 , \3663_b0 , \3664_b1 , \3664_b0 , \3665_b1 , \3665_b0 , \3666_b1 , \3666_b0 , 
		\3667_b1 , \3667_b0 , \3668_b1 , \3668_b0 , \3669_b1 , \3669_b0 , \3670_b1 , \3670_b0 , \3671_b1 , \3671_b0 , 
		\3672_b1 , \3672_b0 , \3673_b1 , \3673_b0 , \3674_b1 , \3674_b0 , \3675_b1 , \3675_b0 , \3676_b1 , \3676_b0 , 
		\3677_b1 , \3677_b0 , \3678_b1 , \3678_b0 , \3679_b1 , \3679_b0 , \3680_b1 , \3680_b0 , \3681_b1 , \3681_b0 , 
		\3682_b1 , \3682_b0 , \3683_b1 , \3683_b0 , \3684_b1 , \3684_b0 , \3685_b1 , \3685_b0 , \3686_b1 , \3686_b0 , 
		\3687_b1 , \3687_b0 , \3688_b1 , \3688_b0 , \3689_b1 , \3689_b0 , \3690_b1 , \3690_b0 , \3691_b1 , \3691_b0 , 
		\3692_b1 , \3692_b0 , \3693_b1 , \3693_b0 , \3694_b1 , \3694_b0 , \3695_b1 , \3695_b0 , \3696_b1 , \3696_b0 , 
		\3697_b1 , \3697_b0 , \3698_b1 , \3698_b0 , \3699_b1 , \3699_b0 , \3700_b1 , \3700_b0 , \3701_b1 , \3701_b0 , 
		\3702_b1 , \3702_b0 , \3703_b1 , \3703_b0 , \3704_b1 , \3704_b0 , \3705_b1 , \3705_b0 , \3706_b1 , \3706_b0 , 
		\3707_b1 , \3707_b0 , \3708_b1 , \3708_b0 , \3709_b1 , \3709_b0 , \3710_b1 , \3710_b0 , \3711_b1 , \3711_b0 , 
		\3712_b1 , \3712_b0 , \3713_b1 , \3713_b0 , \3714_b1 , \3714_b0 , \3715_b1 , \3715_b0 , \3716_b1 , \3716_b0 , 
		\3717_b1 , \3717_b0 , \3718_b1 , \3718_b0 , \3719_b1 , \3719_b0 , \3720_b1 , \3720_b0 , \3721_b1 , \3721_b0 , 
		\3722_b1 , \3722_b0 , \3723_b1 , \3723_b0 , \3724_b1 , \3724_b0 , \3725_b1 , \3725_b0 , \3726_b1 , \3726_b0 , 
		\3727_b1 , \3727_b0 , \3728_b1 , \3728_b0 , \3729_b1 , \3729_b0 , \3730_b1 , \3730_b0 , \3731_b1 , \3731_b0 , 
		\3732_b1 , \3732_b0 , \3733_b1 , \3733_b0 , \3734_b1 , \3734_b0 , \3735_b1 , \3735_b0 , \3736_b1 , \3736_b0 , 
		\3737_b1 , \3737_b0 , \3738_b1 , \3738_b0 , \3739_b1 , \3739_b0 , \3740_b1 , \3740_b0 , \3741_b1 , \3741_b0 , 
		\3742_b1 , \3742_b0 , \3743_b1 , \3743_b0 , \3744_b1 , \3744_b0 , \3745_b1 , \3745_b0 , \3746_b1 , \3746_b0 , 
		\3747_b1 , \3747_b0 , \3748_b1 , \3748_b0 , \3749_b1 , \3749_b0 , \3750_b1 , \3750_b0 , \3751_b1 , \3751_b0 , 
		\3752_b1 , \3752_b0 , \3753_b1 , \3753_b0 , \3754_b1 , \3754_b0 , \3755_b1 , \3755_b0 , \3756_b1 , \3756_b0 , 
		\3757_b1 , \3757_b0 , \3758_b1 , \3758_b0 , \3759_b1 , \3759_b0 , \3760_b1 , \3760_b0 , \3761_b1 , \3761_b0 , 
		\3762_b1 , \3762_b0 , \3763_b1 , \3763_b0 , \3764_b1 , \3764_b0 , \3765_b1 , \3765_b0 , \3766_b1 , \3766_b0 , 
		\3767_b1 , \3767_b0 , \3768_b1 , \3768_b0 , \3769_b1 , \3769_b0 , \3770_b1 , \3770_b0 , \3771_b1 , \3771_b0 , 
		\3772_b1 , \3772_b0 , \3773_b1 , \3773_b0 , \3774_b1 , \3774_b0 , \3775_b1 , \3775_b0 , \3776_b1 , \3776_b0 , 
		\3777_b1 , \3777_b0 , \3778_b1 , \3778_b0 , \3779_b1 , \3779_b0 , \3780_b1 , \3780_b0 , \3781_b1 , \3781_b0 , 
		\3782_b1 , \3782_b0 , \3783_b1 , \3783_b0 , \3784_b1 , \3784_b0 , \3785_b1 , \3785_b0 , \3786_b1 , \3786_b0 , 
		\3787_b1 , \3787_b0 , \3788_b1 , \3788_b0 , \3789_b1 , \3789_b0 , \3790_b1 , \3790_b0 , \3791_b1 , \3791_b0 , 
		\3792_b1 , \3792_b0 , \3793_b1 , \3793_b0 , \3794_b1 , \3794_b0 , \3795_b1 , \3795_b0 , \3796_b1 , \3796_b0 , 
		\3797_b1 , \3797_b0 , \3798_b1 , \3798_b0 , \3799_b1 , \3799_b0 , \3800_b1 , \3800_b0 , \3801_b1 , \3801_b0 , 
		\3802_b1 , \3802_b0 , \3803_b1 , \3803_b0 , \3804_b1 , \3804_b0 , \3805_b1 , \3805_b0 , \3806_b1 , \3806_b0 , 
		\3807_b1 , \3807_b0 , \3808_b1 , \3808_b0 , \3809_b1 , \3809_b0 , \3810_b1 , \3810_b0 , \3811_b1 , \3811_b0 , 
		\3812_b1 , \3812_b0 , \3813_b1 , \3813_b0 , \3814_b1 , \3814_b0 , \3815_b1 , \3815_b0 , \3816_b1 , \3816_b0 , 
		\3817_b1 , \3817_b0 , \3818_b1 , \3818_b0 , \3819_b1 , \3819_b0 , \3820_b1 , \3820_b0 , \3821_b1 , \3821_b0 , 
		\3822_b1 , \3822_b0 , \3823_b1 , \3823_b0 , \3824_b1 , \3824_b0 , \3825_b1 , \3825_b0 , \3826_b1 , \3826_b0 , 
		\3827_b1 , \3827_b0 , \3828_b1 , \3828_b0 , \3829_b1 , \3829_b0 , \3830_b1 , \3830_b0 , \3831_b1 , \3831_b0 , 
		\3832_b1 , \3832_b0 , \3833_b1 , \3833_b0 , \3834_b1 , \3834_b0 , \3835_b1 , \3835_b0 , \3836_b1 , \3836_b0 , 
		\3837_b1 , \3837_b0 , \3838_b1 , \3838_b0 , \3839_b1 , \3839_b0 , \3840_b1 , \3840_b0 , \3841_b1 , \3841_b0 , 
		\3842_b1 , \3842_b0 , \3843_b1 , \3843_b0 , \3844_b1 , \3844_b0 , \3845_b1 , \3845_b0 , \3846_b1 , \3846_b0 , 
		\3847_b1 , \3847_b0 , \3848_b1 , \3848_b0 , \3849_b1 , \3849_b0 , \3850_b1 , \3850_b0 , \3851_b1 , \3851_b0 , 
		\3852_b1 , \3852_b0 , \3853_b1 , \3853_b0 , \3854_b1 , \3854_b0 , \3855_b1 , \3855_b0 , \3856_b1 , \3856_b0 , 
		\3857_b1 , \3857_b0 , \3858_b1 , \3858_b0 , \3859_b1 , \3859_b0 , \3860_b1 , \3860_b0 , \3861_b1 , \3861_b0 , 
		\3862_b1 , \3862_b0 , \3863_b1 , \3863_b0 , \3864_b1 , \3864_b0 , \3865_b1 , \3865_b0 , \3866_b1 , \3866_b0 , 
		\3867_b1 , \3867_b0 , \3868_b1 , \3868_b0 , \3869_b1 , \3869_b0 , \3870_b1 , \3870_b0 , \3871_b1 , \3871_b0 , 
		\3872_b1 , \3872_b0 , \3873_b1 , \3873_b0 , \3874_b1 , \3874_b0 , \3875_b1 , \3875_b0 , \3876_b1 , \3876_b0 , 
		\3877_b1 , \3877_b0 , \3878_b1 , \3878_b0 , \3879_b1 , \3879_b0 , \3880_b1 , \3880_b0 , \3881_b1 , \3881_b0 , 
		\3882_b1 , \3882_b0 , \3883_b1 , \3883_b0 , \3884_b1 , \3884_b0 , \3885_b1 , \3885_b0 , \3886_b1 , \3886_b0 , 
		\3887_b1 , \3887_b0 , \3888_b1 , \3888_b0 , \3889_b1 , \3889_b0 , \3890_b1 , \3890_b0 , \3891_b1 , \3891_b0 , 
		\3892_b1 , \3892_b0 , \3893_b1 , \3893_b0 , \3894_b1 , \3894_b0 , \3895_b1 , \3895_b0 , \3896_b1 , \3896_b0 , 
		\3897_b1 , \3897_b0 , \3898_b1 , \3898_b0 , \3899_b1 , \3899_b0 , \3900_b1 , \3900_b0 , \3901_b1 , \3901_b0 , 
		\3902_b1 , \3902_b0 , \3903_b1 , \3903_b0 , \3904_b1 , \3904_b0 , \3905_b1 , \3905_b0 , \3906_b1 , \3906_b0 , 
		\3907_b1 , \3907_b0 , \3908_b1 , \3908_b0 , \3909_b1 , \3909_b0 , \3910_b1 , \3910_b0 , \3911_b1 , \3911_b0 , 
		\3912_b1 , \3912_b0 , \3913_b1 , \3913_b0 , \3914_b1 , \3914_b0 , \3915_b1 , \3915_b0 , \3916_b1 , \3916_b0 , 
		\3917_b1 , \3917_b0 , \3918_b1 , \3918_b0 , \3919_b1 , \3919_b0 , \3920_b1 , \3920_b0 , \3921_b1 , \3921_b0 , 
		\3922_b1 , \3922_b0 , \3923_b1 , \3923_b0 , \3924_b1 , \3924_b0 , \3925_b1 , \3925_b0 , \3926_b1 , \3926_b0 , 
		\3927_b1 , \3927_b0 , \3928_b1 , \3928_b0 , \3929_b1 , \3929_b0 , \3930_b1 , \3930_b0 , \3931_b1 , \3931_b0 , 
		\3932_b1 , \3932_b0 , \3933_b1 , \3933_b0 , \3934_b1 , \3934_b0 , \3935_b1 , \3935_b0 , \3936_b1 , \3936_b0 , 
		\3937_b1 , \3937_b0 , \3938_b1 , \3938_b0 , \3939_b1 , \3939_b0 , \3940_b1 , \3940_b0 , \3941_b1 , \3941_b0 , 
		\3942_b1 , \3942_b0 , \3943_b1 , \3943_b0 , \3944_b1 , \3944_b0 , \3945_b1 , \3945_b0 , \3946_b1 , \3946_b0 , 
		\3947_b1 , \3947_b0 , \3948_b1 , \3948_b0 , \3949_b1 , \3949_b0 , \3950_b1 , \3950_b0 , \3951_b1 , \3951_b0 , 
		\3952_b1 , \3952_b0 , \3953_b1 , \3953_b0 , \3954_b1 , \3954_b0 , \3955_b1 , \3955_b0 , \3956_b1 , \3956_b0 , 
		\3957_b1 , \3957_b0 , \3958_b1 , \3958_b0 , \3959_b1 , \3959_b0 , \3960_b1 , \3960_b0 , \3961_b1 , \3961_b0 , 
		\3962_b1 , \3962_b0 , \3963_b1 , \3963_b0 , \3964_b1 , \3964_b0 , \3965_b1 , \3965_b0 , \3966_b1 , \3966_b0 , 
		\3967_b1 , \3967_b0 , \3968_b1 , \3968_b0 , \3969_b1 , \3969_b0 , \3970_b1 , \3970_b0 , \3971_b1 , \3971_b0 , 
		\3972_b1 , \3972_b0 , \3973_b1 , \3973_b0 , \3974_b1 , \3974_b0 , \3975_b1 , \3975_b0 , \3976_b1 , \3976_b0 , 
		\3977_b1 , \3977_b0 , \3978_b1 , \3978_b0 , \3979_b1 , \3979_b0 , \3980_b1 , \3980_b0 , \3981_b1 , \3981_b0 , 
		\3982_b1 , \3982_b0 , \3983_b1 , \3983_b0 , \3984_b1 , \3984_b0 , \3985_b1 , \3985_b0 , \3986_b1 , \3986_b0 , 
		\3987_b1 , \3987_b0 , \3988_b1 , \3988_b0 , \3989_b1 , \3989_b0 , \3990_b1 , \3990_b0 , \3991_b1 , \3991_b0 , 
		\3992_b1 , \3992_b0 , \3993_b1 , \3993_b0 , \3994_b1 , \3994_b0 , \3995_b1 , \3995_b0 , \3996_b1 , \3996_b0 , 
		\3997_b1 , \3997_b0 , \3998_b1 , \3998_b0 , \3999_b1 , \3999_b0 , \4000_b1 , \4000_b0 , \4001_b1 , \4001_b0 , 
		\4002_b1 , \4002_b0 , \4003_b1 , \4003_b0 , \4004_b1 , \4004_b0 , \4005_b1 , \4005_b0 , \4006_b1 , \4006_b0 , 
		\4007_b1 , \4007_b0 , \4008_b1 , \4008_b0 , \4009_b1 , \4009_b0 , \4010_b1 , \4010_b0 , \4011_b1 , \4011_b0 , 
		\4012_b1 , \4012_b0 , \4013_b1 , \4013_b0 , \4014_b1 , \4014_b0 , \4015_b1 , \4015_b0 , \4016_b1 , \4016_b0 , 
		\4017_b1 , \4017_b0 , \4018_b1 , \4018_b0 , \4019_b1 , \4019_b0 , \4020_b1 , \4020_b0 , \4021_b1 , \4021_b0 , 
		\4022_b1 , \4022_b0 , \4023_b1 , \4023_b0 , \4024_b1 , \4024_b0 , \4025_b1 , \4025_b0 , \4026_b1 , \4026_b0 , 
		\4027_b1 , \4027_b0 , \4028_b1 , \4028_b0 , \4029_b1 , \4029_b0 , \4030_b1 , \4030_b0 , \4031_b1 , \4031_b0 , 
		\4032_b1 , \4032_b0 , \4033_b1 , \4033_b0 , \4034_b1 , \4034_b0 , \4035_b1 , \4035_b0 , \4036_b1 , \4036_b0 , 
		\4037_b1 , \4037_b0 , \4038_b1 , \4038_b0 , \4039_b1 , \4039_b0 , \4040_b1 , \4040_b0 , \4041_b1 , \4041_b0 , 
		\4042_b1 , \4042_b0 , \4043_b1 , \4043_b0 , \4044_b1 , \4044_b0 , \4045_b1 , \4045_b0 , \4046_b1 , \4046_b0 , 
		\4047_b1 , \4047_b0 , \4048_b1 , \4048_b0 , \4049_b1 , \4049_b0 , \4050_b1 , \4050_b0 , \4051_b1 , \4051_b0 , 
		\4052_b1 , \4052_b0 , \4053_b1 , \4053_b0 , \4054_b1 , \4054_b0 , \4055_b1 , \4055_b0 , \4056_b1 , \4056_b0 , 
		\4057_b1 , \4057_b0 , \4058_b1 , \4058_b0 , \4059_b1 , \4059_b0 , \4060_b1 , \4060_b0 , \4061_b1 , \4061_b0 , 
		\4062_b1 , \4062_b0 , \4063_b1 , \4063_b0 , \4064_b1 , \4064_b0 , \4065_b1 , \4065_b0 , \4066_b1 , \4066_b0 , 
		\4067_b1 , \4067_b0 , \4068_b1 , \4068_b0 , \4069_b1 , \4069_b0 , \4070_b1 , \4070_b0 , \4071_b1 , \4071_b0 , 
		\4072_b1 , \4072_b0 , \4073_b1 , \4073_b0 , \4074_b1 , \4074_b0 , \4075_b1 , \4075_b0 , \4076_b1 , \4076_b0 , 
		\4077_b1 , \4077_b0 , \4078_b1 , \4078_b0 , \4079_b1 , \4079_b0 , \4080_b1 , \4080_b0 , \4081_b1 , \4081_b0 , 
		\4082_b1 , \4082_b0 , \4083_b1 , \4083_b0 , \4084_b1 , \4084_b0 , \4085_b1 , \4085_b0 , \4086_b1 , \4086_b0 , 
		\4087_b1 , \4087_b0 , \4088_b1 , \4088_b0 , \4089_b1 , \4089_b0 , \4090_b1 , \4090_b0 , \4091_b1 , \4091_b0 , 
		\4092_b1 , \4092_b0 , \4093_b1 , \4093_b0 , \4094_b1 , \4094_b0 , \4095_b1 , \4095_b0 , \4096_b1 , \4096_b0 , 
		\4097_b1 , \4097_b0 , \4098_b1 , \4098_b0 , \4099_b1 , \4099_b0 , \4100_b1 , \4100_b0 , \4101_b1 , \4101_b0 , 
		\4102_b1 , \4102_b0 , \4103_b1 , \4103_b0 , \4104_b1 , \4104_b0 , \4105_b1 , \4105_b0 , \4106_b1 , \4106_b0 , 
		\4107_b1 , \4107_b0 , \4108_b1 , \4108_b0 , \4109_b1 , \4109_b0 , \4110_b1 , \4110_b0 , \4111_b1 , \4111_b0 , 
		\4112_b1 , \4112_b0 , \4113_b1 , \4113_b0 , \4114_b1 , \4114_b0 , \4115_b1 , \4115_b0 , \4116_b1 , \4116_b0 , 
		\4117_b1 , \4117_b0 , \4118_b1 , \4118_b0 , \4119_b1 , \4119_b0 , \4120_b1 , \4120_b0 , \4121_b1 , \4121_b0 , 
		\4122_b1 , \4122_b0 , \4123_b1 , \4123_b0 , \4124_b1 , \4124_b0 , \4125_b1 , \4125_b0 , \4126_b1 , \4126_b0 , 
		\4127_b1 , \4127_b0 , \4128_b1 , \4128_b0 , \4129_b1 , \4129_b0 , \4130_b1 , \4130_b0 , \4131_b1 , \4131_b0 , 
		\4132_b1 , \4132_b0 , \4133_b1 , \4133_b0 , \4134_b1 , \4134_b0 , \4135_b1 , \4135_b0 , \4136_b1 , \4136_b0 , 
		\4137_b1 , \4137_b0 , \4138_b1 , \4138_b0 , \4139_b1 , \4139_b0 , \4140_b1 , \4140_b0 , \4141_b1 , \4141_b0 , 
		\4142_b1 , \4142_b0 , \4143_b1 , \4143_b0 , \4144_b1 , \4144_b0 , \4145_b1 , \4145_b0 , \4146_b1 , \4146_b0 , 
		\4147_b1 , \4147_b0 , \4148_b1 , \4148_b0 , \4149_b1 , \4149_b0 , \4150_b1 , \4150_b0 , \4151_b1 , \4151_b0 , 
		\4152_b1 , \4152_b0 , \4153_b1 , \4153_b0 , \4154_b1 , \4154_b0 , \4155_b1 , \4155_b0 , \4156_b1 , \4156_b0 , 
		\4157_b1 , \4157_b0 , \4158_b1 , \4158_b0 , \4159_b1 , \4159_b0 , \4160_b1 , \4160_b0 , \4161_b1 , \4161_b0 , 
		\4162_b1 , \4162_b0 , \4163_b1 , \4163_b0 , \4164_b1 , \4164_b0 , \4165_b1 , \4165_b0 , \4166_b1 , \4166_b0 , 
		\4167_b1 , \4167_b0 , \4168_b1 , \4168_b0 , \4169_b1 , \4169_b0 , \4170_b1 , \4170_b0 , \4171_b1 , \4171_b0 , 
		\4172_b1 , \4172_b0 , \4173_b1 , \4173_b0 , \4174_b1 , \4174_b0 , \4175_b1 , \4175_b0 , \4176_b1 , \4176_b0 , 
		\4177_b1 , \4177_b0 , \4178_b1 , \4178_b0 , \4179_b1 , \4179_b0 , \4180_b1 , \4180_b0 , \4181_b1 , \4181_b0 , 
		\4182_b1 , \4182_b0 , \4183_b1 , \4183_b0 , \4184_b1 , \4184_b0 , \4185_b1 , \4185_b0 , \4186_b1 , \4186_b0 , 
		\4187_b1 , \4187_b0 , \4188_b1 , \4188_b0 , \4189_b1 , \4189_b0 , \4190_b1 , \4190_b0 , \4191_b1 , \4191_b0 , 
		\4192_b1 , \4192_b0 , \4193_b1 , \4193_b0 , \4194_b1 , \4194_b0 , \4195_b1 , \4195_b0 , \4196_b1 , \4196_b0 , 
		\4197_b1 , \4197_b0 , \4198_b1 , \4198_b0 , \4199_b1 , \4199_b0 , \4200_b1 , \4200_b0 , \4201_b1 , \4201_b0 , 
		\4202_b1 , \4202_b0 , \4203_b1 , \4203_b0 , \4204_b1 , \4204_b0 , \4205_b1 , \4205_b0 , \4206_b1 , \4206_b0 , 
		\4207_b1 , \4207_b0 , \4208_b1 , \4208_b0 , \4209_b1 , \4209_b0 , \4210_b1 , \4210_b0 , \4211_b1 , \4211_b0 , 
		\4212_b1 , \4212_b0 , \4213_b1 , \4213_b0 , \4214_b1 , \4214_b0 , \4215_b1 , \4215_b0 , \4216_b1 , \4216_b0 , 
		\4217_b1 , \4217_b0 , \4218_b1 , \4218_b0 , \4219_b1 , \4219_b0 , \4220_b1 , \4220_b0 , \4221_b1 , \4221_b0 , 
		\4222_b1 , \4222_b0 , \4223_b1 , \4223_b0 , \4224_b1 , \4224_b0 , \4225_b1 , \4225_b0 , \4226_b1 , \4226_b0 , 
		\4227_b1 , \4227_b0 , \4228_b1 , \4228_b0 , \4229_b1 , \4229_b0 , \4230_b1 , \4230_b0 , \4231_b1 , \4231_b0 , 
		\4232_b1 , \4232_b0 , \4233_b1 , \4233_b0 , \4234_b1 , \4234_b0 , \4235_b1 , \4235_b0 , \4236_b1 , \4236_b0 , 
		\4237_b1 , \4237_b0 , \4238_b1 , \4238_b0 , \4239_b1 , \4239_b0 , \4240_b1 , \4240_b0 , \4241_b1 , \4241_b0 , 
		\4242_b1 , \4242_b0 , \4243_b1 , \4243_b0 , \4244_b1 , \4244_b0 , \4245_b1 , \4245_b0 , \4246_b1 , \4246_b0 , 
		\4247_b1 , \4247_b0 , \4248_b1 , \4248_b0 , \4249_b1 , \4249_b0 , \4250_b1 , \4250_b0 , \4251_b1 , \4251_b0 , 
		\4252_b1 , \4252_b0 , \4253_b1 , \4253_b0 , \4254_b1 , \4254_b0 , \4255_b1 , \4255_b0 , \4256_b1 , \4256_b0 , 
		\4257_b1 , \4257_b0 , \4258_b1 , \4258_b0 , \4259_b1 , \4259_b0 , \4260_b1 , \4260_b0 , \4261_b1 , \4261_b0 , 
		\4262_b1 , \4262_b0 , \4263_b1 , \4263_b0 , \4264_b1 , \4264_b0 , \4265_b1 , \4265_b0 , \4266_b1 , \4266_b0 , 
		\4267_b1 , \4267_b0 , \4268_b1 , \4268_b0 , \4269_b1 , \4269_b0 , \4270_b1 , \4270_b0 , \4271_b1 , \4271_b0 , 
		\4272_b1 , \4272_b0 , \4273_b1 , \4273_b0 , \4274_b1 , \4274_b0 , \4275_b1 , \4275_b0 , \4276_b1 , \4276_b0 , 
		\4277_b1 , \4277_b0 , \4278_b1 , \4278_b0 , \4279_b1 , \4279_b0 , \4280_b1 , \4280_b0 , \4281_b1 , \4281_b0 , 
		\4282_b1 , \4282_b0 , \4283_b1 , \4283_b0 , \4284_b1 , \4284_b0 , \4285_b1 , \4285_b0 , \4286_b1 , \4286_b0 , 
		\4287_b1 , \4287_b0 , \4288_b1 , \4288_b0 , \4289_b1 , \4289_b0 , \4290_b1 , \4290_b0 , \4291_b1 , \4291_b0 , 
		\4292_b1 , \4292_b0 , \4293_b1 , \4293_b0 , \4294_b1 , \4294_b0 , \4295_b1 , \4295_b0 , \4296_b1 , \4296_b0 , 
		\4297_b1 , \4297_b0 , \4298_b1 , \4298_b0 , \4299_b1 , \4299_b0 , \4300_b1 , \4300_b0 , \4301_b1 , \4301_b0 , 
		\4302_b1 , \4302_b0 , \4303_b1 , \4303_b0 , \4304_b1 , \4304_b0 , \4305_b1 , \4305_b0 , \4306_b1 , \4306_b0 , 
		\4307_b1 , \4307_b0 , \4308_b1 , \4308_b0 , \4309_b1 , \4309_b0 , \4310_b1 , \4310_b0 , \4311_b1 , \4311_b0 , 
		\4312_b1 , \4312_b0 , \4313_b1 , \4313_b0 , \4314_b1 , \4314_b0 , \4315_b1 , \4315_b0 , \4316_b1 , \4316_b0 , 
		\4317_b1 , \4317_b0 , \4318_b1 , \4318_b0 , \4319_b1 , \4319_b0 , \4320_b1 , \4320_b0 , \4321_b1 , \4321_b0 , 
		\4322_b1 , \4322_b0 , \4323_b1 , \4323_b0 , \4324_b1 , \4324_b0 , \4325_b1 , \4325_b0 , \4326_b1 , \4326_b0 , 
		\4327_b1 , \4327_b0 , \4328_b1 , \4328_b0 , \4329_b1 , \4329_b0 , \4330_b1 , \4330_b0 , \4331_b1 , \4331_b0 , 
		\4332_b1 , \4332_b0 , \4333_b1 , \4333_b0 , \4334_b1 , \4334_b0 , \4335_b1 , \4335_b0 , \4336_b1 , \4336_b0 , 
		\4337_b1 , \4337_b0 , \4338_b1 , \4338_b0 , \4339_b1 , \4339_b0 , \4340_b1 , \4340_b0 , \4341_b1 , \4341_b0 , 
		\4342_b1 , \4342_b0 , \4343_b1 , \4343_b0 , \4344_b1 , \4344_b0 , \4345_b1 , \4345_b0 , \4346_b1 , \4346_b0 , 
		\4347_b1 , \4347_b0 , \4348_b1 , \4348_b0 , \4349_b1 , \4349_b0 , \4350_b1 , \4350_b0 , \4351_b1 , \4351_b0 , 
		\4352_b1 , \4352_b0 , \4353_b1 , \4353_b0 , \4354_b1 , \4354_b0 , \4355_b1 , \4355_b0 , \4356_b1 , \4356_b0 , 
		\4357_b1 , \4357_b0 , \4358_b1 , \4358_b0 , \4359_b1 , \4359_b0 , \4360_b1 , \4360_b0 , \4361_b1 , \4361_b0 , 
		\4362_b1 , \4362_b0 , \4363_b1 , \4363_b0 , \4364_b1 , \4364_b0 , \4365_b1 , \4365_b0 , \4366_b1 , \4366_b0 , 
		\4367_b1 , \4367_b0 , \4368_b1 , \4368_b0 , \4369_b1 , \4369_b0 , \4370_b1 , \4370_b0 , \4371_b1 , \4371_b0 , 
		\4372_b1 , \4372_b0 , \4373_b1 , \4373_b0 , \4374_b1 , \4374_b0 , \4375_b1 , \4375_b0 , \4376_b1 , \4376_b0 , 
		\4377_b1 , \4377_b0 , \4378_b1 , \4378_b0 , \4379_b1 , \4379_b0 , \4380_b1 , \4380_b0 , \4381_b1 , \4381_b0 , 
		\4382_b1 , \4382_b0 , \4383_b1 , \4383_b0 , \4384_b1 , \4384_b0 , \4385_b1 , \4385_b0 , \4386_b1 , \4386_b0 , 
		\4387_b1 , \4387_b0 , \4388_b1 , \4388_b0 , \4389_b1 , \4389_b0 , \4390_b1 , \4390_b0 , \4391_b1 , \4391_b0 , 
		\4392_b1 , \4392_b0 , \4393_b1 , \4393_b0 , \4394_b1 , \4394_b0 , \4395_b1 , \4395_b0 , \4396_b1 , \4396_b0 , 
		\4397_b1 , \4397_b0 , \4398_b1 , \4398_b0 , \4399_b1 , \4399_b0 , \4400_b1 , \4400_b0 , \4401_b1 , \4401_b0 , 
		\4402_b1 , \4402_b0 , \4403_b1 , \4403_b0 , \4404_b1 , \4404_b0 , \4405_b1 , \4405_b0 , \4406_b1 , \4406_b0 , 
		\4407_b1 , \4407_b0 , \4408_b1 , \4408_b0 , \4409_b1 , \4409_b0 , \4410_b1 , \4410_b0 , \4411_b1 , \4411_b0 , 
		\4412_b1 , \4412_b0 , \4413_b1 , \4413_b0 , \4414_b1 , \4414_b0 , \4415_b1 , \4415_b0 , \4416_b1 , \4416_b0 , 
		\4417_b1 , \4417_b0 , \4418_b1 , \4418_b0 , \4419_b1 , \4419_b0 , \4420_b1 , \4420_b0 , \4421_b1 , \4421_b0 , 
		\4422_b1 , \4422_b0 , \4423_b1 , \4423_b0 , \4424_b1 , \4424_b0 , \4425_b1 , \4425_b0 , \4426_b1 , \4426_b0 , 
		\4427_b1 , \4427_b0 , \4428_b1 , \4428_b0 , \4429_b1 , \4429_b0 , \4430_b1 , \4430_b0 , \4431_b1 , \4431_b0 , 
		\4432_b1 , \4432_b0 , \4433_b1 , \4433_b0 , \4434_b1 , \4434_b0 , \4435_b1 , \4435_b0 , \4436_b1 , \4436_b0 , 
		\4437_b1 , \4437_b0 , \4438_b1 , \4438_b0 , \4439_b1 , \4439_b0 , \4440_b1 , \4440_b0 , \4441_b1 , \4441_b0 , 
		\4442_b1 , \4442_b0 , \4443_b1 , \4443_b0 , \4444_b1 , \4444_b0 , \4445_b1 , \4445_b0 , \4446_b1 , \4446_b0 , 
		\4447_b1 , \4447_b0 , \4448_b1 , \4448_b0 , \4449_b1 , \4449_b0 , \4450_b1 , \4450_b0 , \4451_b1 , \4451_b0 , 
		\4452_b1 , \4452_b0 , \4453_b1 , \4453_b0 , \4454_b1 , \4454_b0 , \4455_b1 , \4455_b0 , \4456_b1 , \4456_b0 , 
		\4457_b1 , \4457_b0 , \4458_b1 , \4458_b0 , \4459_b1 , \4459_b0 , \4460_b1 , \4460_b0 , \4461_b1 , \4461_b0 , 
		\4462_b1 , \4462_b0 , \4463_b1 , \4463_b0 , \4464_b1 , \4464_b0 , \4465_b1 , \4465_b0 , \4466_b1 , \4466_b0 , 
		\4467_b1 , \4467_b0 , \4468_b1 , \4468_b0 , \4469_b1 , \4469_b0 , \4470_b1 , \4470_b0 , \4471_b1 , \4471_b0 , 
		\4472_b1 , \4472_b0 , \4473_b1 , \4473_b0 , \4474_b1 , \4474_b0 , \4475_b1 , \4475_b0 , \4476_b1 , \4476_b0 , 
		\4477_b1 , \4477_b0 , \4478_b1 , \4478_b0 , \4479_b1 , \4479_b0 , \4480_b1 , \4480_b0 , \4481_b1 , \4481_b0 , 
		\4482_b1 , \4482_b0 , \4483_b1 , \4483_b0 , \4484_b1 , \4484_b0 , \4485_b1 , \4485_b0 , \4486_b1 , \4486_b0 , 
		\4487_b1 , \4487_b0 , \4488_b1 , \4488_b0 , \4489_b1 , \4489_b0 , \4490_b1 , \4490_b0 , \4491_b1 , \4491_b0 , 
		\4492_b1 , \4492_b0 , \4493_b1 , \4493_b0 , \4494_b1 , \4494_b0 , \4495_b1 , \4495_b0 , \4496_b1 , \4496_b0 , 
		\4497_b1 , \4497_b0 , \4498_b1 , \4498_b0 , \4499_b1 , \4499_b0 , \4500_b1 , \4500_b0 , \4501_b1 , \4501_b0 , 
		\4502_b1 , \4502_b0 , \4503_b1 , \4503_b0 , \4504_b1 , \4504_b0 , \4505_b1 , \4505_b0 , \4506_b1 , \4506_b0 , 
		\4507_b1 , \4507_b0 , \4508_b1 , \4508_b0 , \4509_b1 , \4509_b0 , \4510_b1 , \4510_b0 , \4511_b1 , \4511_b0 , 
		\4512_b1 , \4512_b0 , \4513_b1 , \4513_b0 , \4514_b1 , \4514_b0 , \4515_b1 , \4515_b0 , \4516_b1 , \4516_b0 , 
		\4517_b1 , \4517_b0 , \4518_b1 , \4518_b0 , \4519_b1 , \4519_b0 , \4520_b1 , \4520_b0 , \4521_b1 , \4521_b0 , 
		\4522_b1 , \4522_b0 , \4523_b1 , \4523_b0 , \4524_b1 , \4524_b0 , \4525_b1 , \4525_b0 , \4526_b1 , \4526_b0 , 
		\4527_b1 , \4527_b0 , \4528_b1 , \4528_b0 , \4529_b1 , \4529_b0 , \4530_b1 , \4530_b0 , \4531_b1 , \4531_b0 , 
		\4532_b1 , \4532_b0 , \4533_b1 , \4533_b0 , \4534_b1 , \4534_b0 , \4535_b1 , \4535_b0 , \4536_b1 , \4536_b0 , 
		\4537_b1 , \4537_b0 , \4538_b1 , \4538_b0 , \4539_b1 , \4539_b0 , \4540_b1 , \4540_b0 , \4541_b1 , \4541_b0 , 
		\4542_b1 , \4542_b0 , \4543_b1 , \4543_b0 , \4544_b1 , \4544_b0 , \4545_b1 , \4545_b0 , \4546_b1 , \4546_b0 , 
		\4547_b1 , \4547_b0 , \4548_b1 , \4548_b0 , \4549_b1 , \4549_b0 , \4550_b1 , \4550_b0 , \4551_b1 , \4551_b0 , 
		\4552_b1 , \4552_b0 , \4553_b1 , \4553_b0 , \4554_b1 , \4554_b0 , \4555_b1 , \4555_b0 , \4556_b1 , \4556_b0 , 
		\4557_b1 , \4557_b0 , \4558_b1 , \4558_b0 , \4559_b1 , \4559_b0 , \4560_b1 , \4560_b0 , \4561_b1 , \4561_b0 , 
		\4562_b1 , \4562_b0 , \4563_b1 , \4563_b0 , \4564_b1 , \4564_b0 , \4565_b1 , \4565_b0 , \4566_b1 , \4566_b0 , 
		\4567_b1 , \4567_b0 , \4568_b1 , \4568_b0 , \4569_b1 , \4569_b0 , \4570_b1 , \4570_b0 , \4571_b1 , \4571_b0 , 
		\4572_b1 , \4572_b0 , \4573_b1 , \4573_b0 , \4574_b1 , \4574_b0 , \4575_b1 , \4575_b0 , \4576_b1 , \4576_b0 , 
		\4577_b1 , \4577_b0 , \4578_b1 , \4578_b0 , \4579_b1 , \4579_b0 , \4580_b1 , \4580_b0 , \4581_b1 , \4581_b0 , 
		\4582_b1 , \4582_b0 , \4583_b1 , \4583_b0 , \4584_b1 , \4584_b0 , \4585_b1 , \4585_b0 , \4586_b1 , \4586_b0 , 
		\4587_b1 , \4587_b0 , \4588_b1 , \4588_b0 , \4589_b1 , \4589_b0 , \4590_b1 , \4590_b0 , \4591_b1 , \4591_b0 , 
		\4592_b1 , \4592_b0 , \4593_b1 , \4593_b0 , \4594_b1 , \4594_b0 , \4595_b1 , \4595_b0 , \4596_b1 , \4596_b0 , 
		\4597_b1 , \4597_b0 , \4598_b1 , \4598_b0 , \4599_b1 , \4599_b0 , \4600_b1 , \4600_b0 , \4601_b1 , \4601_b0 , 
		\4602_b1 , \4602_b0 , \4603_b1 , \4603_b0 , \4604_b1 , \4604_b0 , \4605_b1 , \4605_b0 , \4606_b1 , \4606_b0 , 
		\4607_b1 , \4607_b0 , \4608_b1 , \4608_b0 , \4609_b1 , \4609_b0 , \4610_b1 , \4610_b0 , \4611_b1 , \4611_b0 , 
		\4612_b1 , \4612_b0 , \4613_b1 , \4613_b0 , \4614_b1 , \4614_b0 , \4615_b1 , \4615_b0 , \4616_b1 , \4616_b0 , 
		\4617_b1 , \4617_b0 , \4618_b1 , \4618_b0 , \4619_b1 , \4619_b0 , \4620_b1 , \4620_b0 , \4621_b1 , \4621_b0 , 
		\4622_b1 , \4622_b0 , \4623_b1 , \4623_b0 , \4624_b1 , \4624_b0 , \4625_b1 , \4625_b0 , \4626_b1 , \4626_b0 , 
		\4627_b1 , \4627_b0 , \4628_b1 , \4628_b0 , \4629_b1 , \4629_b0 , \4630_b1 , \4630_b0 , \4631_b1 , \4631_b0 , 
		\4632_b1 , \4632_b0 , \4633_b1 , \4633_b0 , \4634_b1 , \4634_b0 , \4635_b1 , \4635_b0 , \4636_b1 , \4636_b0 , 
		\4637_b1 , \4637_b0 , \4638_b1 , \4638_b0 , \4639_b1 , \4639_b0 , \4640_b1 , \4640_b0 , \4641_b1 , \4641_b0 , 
		\4642_b1 , \4642_b0 , \4643_b1 , \4643_b0 , \4644_b1 , \4644_b0 , \4645_b1 , \4645_b0 , \4646_b1 , \4646_b0 , 
		\4647_b1 , \4647_b0 , \4648_b1 , \4648_b0 , \4649_b1 , \4649_b0 , \4650_b1 , \4650_b0 , \4651_b1 , \4651_b0 , 
		\4652_b1 , \4652_b0 , \4653_b1 , \4653_b0 , \4654_b1 , \4654_b0 , \4655_b1 , \4655_b0 , \4656_b1 , \4656_b0 , 
		\4657_b1 , \4657_b0 , \4658_b1 , \4658_b0 , \4659_b1 , \4659_b0 , \4660_b1 , \4660_b0 , \4661_b1 , \4661_b0 , 
		\4662_b1 , \4662_b0 , \4663_b1 , \4663_b0 , \4664_b1 , \4664_b0 , \4665_b1 , \4665_b0 , \4666_b1 , \4666_b0 , 
		\4667_b1 , \4667_b0 , \4668_b1 , \4668_b0 , \4669_b1 , \4669_b0 , \4670_b1 , \4670_b0 , \4671_b1 , \4671_b0 , 
		\4672_b1 , \4672_b0 , \4673_b1 , \4673_b0 , \4674_b1 , \4674_b0 , \4675_b1 , \4675_b0 , \4676_b1 , \4676_b0 , 
		\4677_b1 , \4677_b0 , \4678_b1 , \4678_b0 , \4679_b1 , \4679_b0 , \4680_b1 , \4680_b0 , \4681_b1 , \4681_b0 , 
		\4682_b1 , \4682_b0 , \4683_b1 , \4683_b0 , \4684_b1 , \4684_b0 , \4685_b1 , \4685_b0 , \4686_b1 , \4686_b0 , 
		\4687_b1 , \4687_b0 , \4688_b1 , \4688_b0 , \4689_b1 , \4689_b0 , \4690_b1 , \4690_b0 , \4691_b1 , \4691_b0 , 
		\4692_b1 , \4692_b0 , \4693_b1 , \4693_b0 , \4694_b1 , \4694_b0 , \4695_b1 , \4695_b0 , \4696_b1 , \4696_b0 , 
		\4697_b1 , \4697_b0 , \4698_b1 , \4698_b0 , \4699_b1 , \4699_b0 , \4700_b1 , \4700_b0 , \4701_b1 , \4701_b0 , 
		\4702_b1 , \4702_b0 , \4703_b1 , \4703_b0 , \4704_b1 , \4704_b0 , \4705_b1 , \4705_b0 , \4706_b1 , \4706_b0 , 
		\4707_b1 , \4707_b0 , \4708_b1 , \4708_b0 , \4709_b1 , \4709_b0 , \4710_b1 , \4710_b0 , \4711_b1 , \4711_b0 , 
		\4712_b1 , \4712_b0 , \4713_b1 , \4713_b0 , \4714_b1 , \4714_b0 , \4715_b1 , \4715_b0 , \4716_b1 , \4716_b0 , 
		\4717_b1 , \4717_b0 , \4718_b1 , \4718_b0 , \4719_b1 , \4719_b0 , \4720_b1 , \4720_b0 , \4721_b1 , \4721_b0 , 
		\4722_b1 , \4722_b0 , \4723_b1 , \4723_b0 , \4724_b1 , \4724_b0 , \4725_b1 , \4725_b0 , \4726_b1 , \4726_b0 , 
		\4727_b1 , \4727_b0 , \4728_b1 , \4728_b0 , \4729_b1 , \4729_b0 , \4730_b1 , \4730_b0 , \4731_b1 , \4731_b0 , 
		\4732_b1 , \4732_b0 , \4733_b1 , \4733_b0 , \4734_b1 , \4734_b0 , \4735_b1 , \4735_b0 , \4736_b1 , \4736_b0 , 
		\4737_b1 , \4737_b0 , \4738_b1 , \4738_b0 , \4739_b1 , \4739_b0 , \4740_b1 , \4740_b0 , \4741_b1 , \4741_b0 , 
		\4742_b1 , \4742_b0 , \4743_b1 , \4743_b0 , \4744_b1 , \4744_b0 , \4745_b1 , \4745_b0 , \4746_b1 , \4746_b0 , 
		\4747_b1 , \4747_b0 , \4748_b1 , \4748_b0 , \4749_b1 , \4749_b0 , \4750_b1 , \4750_b0 , \4751_b1 , \4751_b0 , 
		\4752_b1 , \4752_b0 , \4753_b1 , \4753_b0 , \4754_b1 , \4754_b0 , \4755_b1 , \4755_b0 , \4756_b1 , \4756_b0 , 
		\4757_b1 , \4757_b0 , \4758_b1 , \4758_b0 , \4759_b1 , \4759_b0 , \4760_b1 , \4760_b0 , \4761_b1 , \4761_b0 , 
		\4762_b1 , \4762_b0 , \4763_b1 , \4763_b0 , \4764_b1 , \4764_b0 , \4765_b1 , \4765_b0 , \4766_b1 , \4766_b0 , 
		\4767_b1 , \4767_b0 , \4768_b1 , \4768_b0 , \4769_b1 , \4769_b0 , \4770_b1 , \4770_b0 , \4771_b1 , \4771_b0 , 
		\4772_b1 , \4772_b0 , \4773_b1 , \4773_b0 , \4774_b1 , \4774_b0 , \4775_b1 , \4775_b0 , \4776_b1 , \4776_b0 , 
		\4777_b1 , \4777_b0 , \4778_b1 , \4778_b0 , \4779_b1 , \4779_b0 , \4780_b1 , \4780_b0 , \4781_b1 , \4781_b0 , 
		\4782_b1 , \4782_b0 , \4783_b1 , \4783_b0 , \4784_b1 , \4784_b0 , \4785_b1 , \4785_b0 , \4786_b1 , \4786_b0 , 
		\4787_b1 , \4787_b0 , \4788_b1 , \4788_b0 , \4789_b1 , \4789_b0 , \4790_b1 , \4790_b0 , \4791_b1 , \4791_b0 , 
		\4792_b1 , \4792_b0 , \4793_b1 , \4793_b0 , \4794_b1 , \4794_b0 , \4795_b1 , \4795_b0 , \4796_b1 , \4796_b0 , 
		\4797_b1 , \4797_b0 , \4798_b1 , \4798_b0 , \4799_b1 , \4799_b0 , \4800_b1 , \4800_b0 , \4801_b1 , \4801_b0 , 
		\4802_b1 , \4802_b0 , \4803_b1 , \4803_b0 , \4804_b1 , \4804_b0 , \4805_b1 , \4805_b0 , \4806_b1 , \4806_b0 , 
		\4807_b1 , \4807_b0 , \4808_b1 , \4808_b0 , \4809_b1 , \4809_b0 , \4810_b1 , \4810_b0 , \4811_b1 , \4811_b0 , 
		\4812_b1 , \4812_b0 , \4813_b1 , \4813_b0 , \4814_b1 , \4814_b0 , \4815_b1 , \4815_b0 , \4816_b1 , \4816_b0 , 
		\4817_b1 , \4817_b0 , \4818_b1 , \4818_b0 , \4819_b1 , \4819_b0 , \4820_b1 , \4820_b0 , \4821_b1 , \4821_b0 , 
		\4822_b1 , \4822_b0 , \4823_b1 , \4823_b0 , \4824_b1 , \4824_b0 , \4825_b1 , \4825_b0 , \4826_b1 , \4826_b0 , 
		\4827_b1 , \4827_b0 , \4828_b1 , \4828_b0 , \4829_b1 , \4829_b0 , \4830_b1 , \4830_b0 , \4831_b1 , \4831_b0 , 
		\4832_b1 , \4832_b0 , \4833_b1 , \4833_b0 , \4834_b1 , \4834_b0 , \4835_b1 , \4835_b0 , \4836_b1 , \4836_b0 , 
		\4837_b1 , \4837_b0 , \4838_b1 , \4838_b0 , \4839_b1 , \4839_b0 , \4840_b1 , \4840_b0 , \4841_b1 , \4841_b0 , 
		\4842_b1 , \4842_b0 , \4843_b1 , \4843_b0 , \4844_b1 , \4844_b0 , \4845_b1 , \4845_b0 , \4846_b1 , \4846_b0 , 
		\4847_b1 , \4847_b0 , \4848_b1 , \4848_b0 , \4849_b1 , \4849_b0 , \4850_b1 , \4850_b0 , \4851_b1 , \4851_b0 , 
		\4852_b1 , \4852_b0 , \4853_b1 , \4853_b0 , \4854_b1 , \4854_b0 , \4855_b1 , \4855_b0 , \4856_b1 , \4856_b0 , 
		\4857_b1 , \4857_b0 , \4858_b1 , \4858_b0 , \4859_b1 , \4859_b0 , \4860_b1 , \4860_b0 , \4861_b1 , \4861_b0 , 
		\4862_b1 , \4862_b0 , \4863_b1 , \4863_b0 , \4864_b1 , \4864_b0 , \4865_b1 , \4865_b0 , \4866_b1 , \4866_b0 , 
		\4867_b1 , \4867_b0 , \4868_b1 , \4868_b0 , \4869_b1 , \4869_b0 , \4870_b1 , \4870_b0 , \4871_b1 , \4871_b0 , 
		\4872_b1 , \4872_b0 , \4873_b1 , \4873_b0 , \4874_b1 , \4874_b0 , \4875_b1 , \4875_b0 , \4876_b1 , \4876_b0 , 
		\4877_b1 , \4877_b0 , \4878_b1 , \4878_b0 , \4879_b1 , \4879_b0 , \4880_b1 , \4880_b0 , \4881_b1 , \4881_b0 , 
		\4882_b1 , \4882_b0 , \4883_b1 , \4883_b0 , \4884_b1 , \4884_b0 , \4885_b1 , \4885_b0 , \4886_b1 , \4886_b0 , 
		\4887_b1 , \4887_b0 , \4888_b1 , \4888_b0 , \4889_b1 , \4889_b0 , \4890_b1 , \4890_b0 , \4891_b1 , \4891_b0 , 
		\4892_b1 , \4892_b0 , \4893_b1 , \4893_b0 , \4894_b1 , \4894_b0 , \4895_b1 , \4895_b0 , \4896_b1 , \4896_b0 , 
		\4897_b1 , \4897_b0 , \4898_b1 , \4898_b0 , \4899_b1 , \4899_b0 , \4900_b1 , \4900_b0 , \4901_b1 , \4901_b0 , 
		\4902_b1 , \4902_b0 , \4903_b1 , \4903_b0 , \4904_b1 , \4904_b0 , \4905_b1 , \4905_b0 , \4906_b1 , \4906_b0 , 
		\4907_b1 , \4907_b0 , \4908_b1 , \4908_b0 , \4909_b1 , \4909_b0 , \4910_b1 , \4910_b0 , \4911_b1 , \4911_b0 , 
		\4912_b1 , \4912_b0 , \4913_b1 , \4913_b0 , \4914_b1 , \4914_b0 , \4915_b1 , \4915_b0 , \4916_b1 , \4916_b0 , 
		\4917_b1 , \4917_b0 , \4918_b1 , \4918_b0 , \4919_b1 , \4919_b0 , \4920_b1 , \4920_b0 , \4921_b1 , \4921_b0 , 
		\4922_b1 , \4922_b0 , \4923_b1 , \4923_b0 , \4924_b1 , \4924_b0 , \4925_b1 , \4925_b0 , \4926_b1 , \4926_b0 , 
		\4927_b1 , \4927_b0 , \4928_b1 , \4928_b0 , \4929_b1 , \4929_b0 , \4930_b1 , \4930_b0 , \4931_b1 , \4931_b0 , 
		\4932_b1 , \4932_b0 , \4933_b1 , \4933_b0 , \4934_b1 , \4934_b0 , \4935_b1 , \4935_b0 , \4936_b1 , \4936_b0 , 
		\4937_b1 , \4937_b0 , \4938_b1 , \4938_b0 , \4939_b1 , \4939_b0 , \4940_b1 , \4940_b0 , \4941_b1 , \4941_b0 , 
		\4942_b1 , \4942_b0 , \4943_b1 , \4943_b0 , \4944_b1 , \4944_b0 , \4945_b1 , \4945_b0 , \4946_b1 , \4946_b0 , 
		\4947_b1 , \4947_b0 , \4948_b1 , \4948_b0 , \4949_b1 , \4949_b0 , \4950_b1 , \4950_b0 , \4951_b1 , \4951_b0 , 
		\4952_b1 , \4952_b0 , \4953_b1 , \4953_b0 , \4954_b1 , \4954_b0 , \4955_b1 , \4955_b0 , \4956_b1 , \4956_b0 , 
		\4957_b1 , \4957_b0 , \4958_b1 , \4958_b0 , \4959_b1 , \4959_b0 , \4960_b1 , \4960_b0 , \4961_b1 , \4961_b0 , 
		\4962_b1 , \4962_b0 , \4963_b1 , \4963_b0 , \4964_b1 , \4964_b0 , \4965_b1 , \4965_b0 , \4966_b1 , \4966_b0 , 
		\4967_b1 , \4967_b0 , \4968_b1 , \4968_b0 , \4969_b1 , \4969_b0 , \4970_b1 , \4970_b0 , \4971_b1 , \4971_b0 , 
		\4972_b1 , \4972_b0 , \4973_b1 , \4973_b0 , \4974_b1 , \4974_b0 , \4975_b1 , \4975_b0 , \4976_b1 , \4976_b0 , 
		\4977_b1 , \4977_b0 , \4978_b1 , \4978_b0 , \4979_b1 , \4979_b0 , \4980_b1 , \4980_b0 , \4981_b1 , \4981_b0 , 
		\4982_b1 , \4982_b0 , \4983_b1 , \4983_b0 , \4984_b1 , \4984_b0 , \4985_b1 , \4985_b0 , \4986_b1 , \4986_b0 , 
		\4987_b1 , \4987_b0 , \4988_b1 , \4988_b0 , \4989_b1 , \4989_b0 , \4990_b1 , \4990_b0 , \4991_b1 , \4991_b0 , 
		\4992_b1 , \4992_b0 , \4993_b1 , \4993_b0 , \4994_b1 , \4994_b0 , \4995_b1 , \4995_b0 , \4996_b1 , \4996_b0 , 
		\4997_b1 , \4997_b0 , \4998_b1 , \4998_b0 , \4999_b1 , \4999_b0 , \5000_b1 , \5000_b0 , \5001_b1 , \5001_b0 , 
		\5002_b1 , \5002_b0 , \5003_b1 , \5003_b0 , \5004_b1 , \5004_b0 , \5005_b1 , \5005_b0 , \5006_b1 , \5006_b0 , 
		\5007_b1 , \5007_b0 , \5008_b1 , \5008_b0 , \5009_b1 , \5009_b0 , \5010_b1 , \5010_b0 , \5011_b1 , \5011_b0 , 
		\5012_b1 , \5012_b0 , \5013_b1 , \5013_b0 , \5014_b1 , \5014_b0 , \5015_b1 , \5015_b0 , \5016_b1 , \5016_b0 , 
		\5017_b1 , \5017_b0 , \5018_b1 , \5018_b0 , \5019_b1 , \5019_b0 , \5020_b1 , \5020_b0 , \5021_b1 , \5021_b0 , 
		\5022_b1 , \5022_b0 , \5023_b1 , \5023_b0 , \5024_b1 , \5024_b0 , \5025_b1 , \5025_b0 , \5026_b1 , \5026_b0 , 
		\5027_b1 , \5027_b0 , \5028_b1 , \5028_b0 , \5029_b1 , \5029_b0 , \5030_b1 , \5030_b0 , \5031_b1 , \5031_b0 , 
		\5032_b1 , \5032_b0 , \5033_b1 , \5033_b0 , \5034_b1 , \5034_b0 , \5035_b1 , \5035_b0 , \5036_b1 , \5036_b0 , 
		\5037_b1 , \5037_b0 , \5038_b1 , \5038_b0 , \5039_b1 , \5039_b0 , \5040_b1 , \5040_b0 , \5041_b1 , \5041_b0 , 
		\5042_b1 , \5042_b0 , \5043_b1 , \5043_b0 , \5044_b1 , \5044_b0 , \5045_b1 , \5045_b0 , \5046_b1 , \5046_b0 , 
		\5047_b1 , \5047_b0 , \5048_b1 , \5048_b0 , \5049_b1 , \5049_b0 , \5050_b1 , \5050_b0 , \5051_b1 , \5051_b0 , 
		\5052_b1 , \5052_b0 , \5053_b1 , \5053_b0 , \5054_b1 , \5054_b0 , \5055_b1 , \5055_b0 , \5056_b1 , \5056_b0 , 
		\5057_b1 , \5057_b0 , \5058_b1 , \5058_b0 , \5059_b1 , \5059_b0 , \5060_b1 , \5060_b0 , \5061_b1 , \5061_b0 , 
		\5062_b1 , \5062_b0 , \5063_b1 , \5063_b0 , \5064_b1 , \5064_b0 , \5065_b1 , \5065_b0 , \5066_b1 , \5066_b0 , 
		\5067_b1 , \5067_b0 , \5068_b1 , \5068_b0 , \5069_b1 , \5069_b0 , \5070_b1 , \5070_b0 , \5071_b1 , \5071_b0 , 
		\5072_b1 , \5072_b0 , \5073_b1 , \5073_b0 , \5074_b1 , \5074_b0 , \5075_b1 , \5075_b0 , \5076_b1 , \5076_b0 , 
		\5077_b1 , \5077_b0 , \5078_b1 , \5078_b0 , \5079_b1 , \5079_b0 , \5080_b1 , \5080_b0 , \5081_b1 , \5081_b0 , 
		\5082_b1 , \5082_b0 , \5083_b1 , \5083_b0 , \5084_b1 , \5084_b0 , \5085_b1 , \5085_b0 , \5086_b1 , \5086_b0 , 
		\5087_b1 , \5087_b0 , \5088_b1 , \5088_b0 , \5089_b1 , \5089_b0 , \5090_b1 , \5090_b0 , \5091_b1 , \5091_b0 , 
		\5092_b1 , \5092_b0 , \5093_b1 , \5093_b0 , \5094_b1 , \5094_b0 , \5095_b1 , \5095_b0 , \5096_b1 , \5096_b0 , 
		\5097_b1 , \5097_b0 , \5098_b1 , \5098_b0 , \5099_b1 , \5099_b0 , \5100_b1 , \5100_b0 , \5101_b1 , \5101_b0 , 
		\5102_b1 , \5102_b0 , \5103_b1 , \5103_b0 , \5104_b1 , \5104_b0 , \5105_b1 , \5105_b0 , \5106_b1 , \5106_b0 , 
		\5107_b1 , \5107_b0 , \5108_b1 , \5108_b0 , \5109_b1 , \5109_b0 , \5110_b1 , \5110_b0 , \5111_b1 , \5111_b0 , 
		\5112_b1 , \5112_b0 , \5113_b1 , \5113_b0 , \5114_b1 , \5114_b0 , \5115_b1 , \5115_b0 , \5116_b1 , \5116_b0 , 
		\5117_b1 , \5117_b0 , \5118_b1 , \5118_b0 , \5119_b1 , \5119_b0 , \5120_b1 , \5120_b0 , \5121_b1 , \5121_b0 , 
		\5122_b1 , \5122_b0 , \5123_b1 , \5123_b0 , \5124_b1 , \5124_b0 , \5125_b1 , \5125_b0 , \5126_b1 , \5126_b0 , 
		\5127_b1 , \5127_b0 , \5128_b1 , \5128_b0 , \5129_b1 , \5129_b0 , \5130_b1 , \5130_b0 , \5131_b1 , \5131_b0 , 
		\5132_b1 , \5132_b0 , \5133_b1 , \5133_b0 , \5134_b1 , \5134_b0 , \5135_b1 , \5135_b0 , \5136_b1 , \5136_b0 , 
		\5137_b1 , \5137_b0 , \5138_b1 , \5138_b0 , \5139_b1 , \5139_b0 , \5140_b1 , \5140_b0 , \5141_b1 , \5141_b0 , 
		\5142_b1 , \5142_b0 , \5143_b1 , \5143_b0 , \5144_b1 , \5144_b0 , \5145_b1 , \5145_b0 , \5146_b1 , \5146_b0 , 
		\5147_b1 , \5147_b0 , \5148_b1 , \5148_b0 , \5149_b1 , \5149_b0 , \5150_b1 , \5150_b0 , \5151_b1 , \5151_b0 , 
		\5152_b1 , \5152_b0 , \5153_b1 , \5153_b0 , \5154_b1 , \5154_b0 , \5155_b1 , \5155_b0 , \5156_b1 , \5156_b0 , 
		\5157_b1 , \5157_b0 , \5158_b1 , \5158_b0 , \5159_b1 , \5159_b0 , \5160_b1 , \5160_b0 , \5161_b1 , \5161_b0 , 
		\5162_b1 , \5162_b0 , \5163_b1 , \5163_b0 , \5164_b1 , \5164_b0 , \5165_b1 , \5165_b0 , \5166_b1 , \5166_b0 , 
		\5167_b1 , \5167_b0 , \5168_b1 , \5168_b0 , \5169_b1 , \5169_b0 , \5170_b1 , \5170_b0 , \5171_b1 , \5171_b0 , 
		\5172_b1 , \5172_b0 , \5173_b1 , \5173_b0 , \5174_b1 , \5174_b0 , \5175_b1 , \5175_b0 , \5176_b1 , \5176_b0 , 
		\5177_b1 , \5177_b0 , \5178_b1 , \5178_b0 , \5179_b1 , \5179_b0 , \5180_b1 , \5180_b0 , \5181_b1 , \5181_b0 , 
		\5182_b1 , \5182_b0 , \5183_b1 , \5183_b0 , \5184_b1 , \5184_b0 , \5185_b1 , \5185_b0 , \5186_b1 , \5186_b0 , 
		\5187_b1 , \5187_b0 , \5188_b1 , \5188_b0 , \5189_b1 , \5189_b0 , \5190_b1 , \5190_b0 , \5191_b1 , \5191_b0 , 
		\5192_b1 , \5192_b0 , \5193_b1 , \5193_b0 , \5194_b1 , \5194_b0 , \5195_b1 , \5195_b0 , \5196_b1 , \5196_b0 , 
		\5197_b1 , \5197_b0 , \5198_b1 , \5198_b0 , \5199_b1 , \5199_b0 , \5200_b1 , \5200_b0 , \5201_b1 , \5201_b0 , 
		\5202_b1 , \5202_b0 , \5203_b1 , \5203_b0 , \5204_b1 , \5204_b0 , \5205_b1 , \5205_b0 , \5206_b1 , \5206_b0 , 
		\5207_b1 , \5207_b0 , \5208_b1 , \5208_b0 , \5209_b1 , \5209_b0 , \5210_b1 , \5210_b0 , \5211_b1 , \5211_b0 , 
		\5212_b1 , \5212_b0 , \5213_b1 , \5213_b0 , \5214_b1 , \5214_b0 , \5215_b1 , \5215_b0 , \5216_b1 , \5216_b0 , 
		\5217_b1 , \5217_b0 , \5218_b1 , \5218_b0 , \5219_b1 , \5219_b0 , \5220_b1 , \5220_b0 , \5221_b1 , \5221_b0 , 
		\5222_b1 , \5222_b0 , \5223_b1 , \5223_b0 , \5224_b1 , \5224_b0 , \5225_b1 , \5225_b0 , \5226_b1 , \5226_b0 , 
		\5227_b1 , \5227_b0 , \5228_b1 , \5228_b0 , \5229_b1 , \5229_b0 , \5230_b1 , \5230_b0 , \5231_b1 , \5231_b0 , 
		\5232_b1 , \5232_b0 , \5233_b1 , \5233_b0 , \5234_b1 , \5234_b0 , \5235_b1 , \5235_b0 , \5236_b1 , \5236_b0 , 
		\5237_b1 , \5237_b0 , \5238_b1 , \5238_b0 , \5239_b1 , \5239_b0 , \5240_b1 , \5240_b0 , \5241_b1 , \5241_b0 , 
		\5242_b1 , \5242_b0 , \5243_b1 , \5243_b0 , \5244_b1 , \5244_b0 , \5245_b1 , \5245_b0 , \5246_b1 , \5246_b0 , 
		\5247_b1 , \5247_b0 , \5248_b1 , \5248_b0 , \5249_b1 , \5249_b0 , \5250_b1 , \5250_b0 , \5251_b1 , \5251_b0 , 
		\5252_b1 , \5252_b0 , \5253_b1 , \5253_b0 , \5254_b1 , \5254_b0 , \5255_b1 , \5255_b0 , \5256_b1 , \5256_b0 , 
		\5257_b1 , \5257_b0 , \5258_b1 , \5258_b0 , \5259_b1 , \5259_b0 , \5260_b1 , \5260_b0 , \5261_b1 , \5261_b0 , 
		\5262_b1 , \5262_b0 , \5263_b1 , \5263_b0 , \5264_b1 , \5264_b0 , \5265_b1 , \5265_b0 , \5266_b1 , \5266_b0 , 
		\5267_b1 , \5267_b0 , \5268_b1 , \5268_b0 , \5269_b1 , \5269_b0 , \5270_b1 , \5270_b0 , \5271_b1 , \5271_b0 , 
		\5272_b1 , \5272_b0 , \5273_b1 , \5273_b0 , \5274_b1 , \5274_b0 , \5275_b1 , \5275_b0 , \5276_b1 , \5276_b0 , 
		\5277_b1 , \5277_b0 , \5278_b1 , \5278_b0 , \5279_b1 , \5279_b0 , \5280_b1 , \5280_b0 , \5281_b1 , \5281_b0 , 
		\5282_b1 , \5282_b0 , \5283_b1 , \5283_b0 , \5284_b1 , \5284_b0 , \5285_b1 , \5285_b0 , \5286_b1 , \5286_b0 , 
		\5287_b1 , \5287_b0 , \5288_b1 , \5288_b0 , \5289_b1 , \5289_b0 , \5290_b1 , \5290_b0 , \5291_b1 , \5291_b0 , 
		\5292_b1 , \5292_b0 , \5293_b1 , \5293_b0 , \5294_b1 , \5294_b0 , \5295_b1 , \5295_b0 , \5296_b1 , \5296_b0 , 
		\5297_b1 , \5297_b0 , \5298_b1 , \5298_b0 , \5299_b1 , \5299_b0 , \5300_b1 , \5300_b0 , \5301_b1 , \5301_b0 , 
		\5302_b1 , \5302_b0 , \5303_b1 , \5303_b0 , \5304_b1 , \5304_b0 , \5305_b1 , \5305_b0 , \5306_b1 , \5306_b0 , 
		\5307_b1 , \5307_b0 , \5308_b1 , \5308_b0 , \5309_b1 , \5309_b0 , \5310_b1 , \5310_b0 , \5311_b1 , \5311_b0 , 
		\5312_b1 , \5312_b0 , \5313_b1 , \5313_b0 , \5314_b1 , \5314_b0 , \5315_b1 , \5315_b0 , \5316_b1 , \5316_b0 , 
		\5317_b1 , \5317_b0 , \5318_b1 , \5318_b0 , \5319_b1 , \5319_b0 , \5320_b1 , \5320_b0 , \5321_b1 , \5321_b0 , 
		\5322_b1 , \5322_b0 , \5323_b1 , \5323_b0 , \5324_b1 , \5324_b0 , \5325_b1 , \5325_b0 , \5326_b1 , \5326_b0 , 
		\5327_b1 , \5327_b0 , \5328_b1 , \5328_b0 , \5329_b1 , \5329_b0 , \5330_b1 , \5330_b0 , \5331_b1 , \5331_b0 , 
		\5332_b1 , \5332_b0 , \5333_b1 , \5333_b0 , \5334_b1 , \5334_b0 , \5335_b1 , \5335_b0 , \5336_b1 , \5336_b0 , 
		\5337_b1 , \5337_b0 , \5338_b1 , \5338_b0 , \5339_b1 , \5339_b0 , \5340_b1 , \5340_b0 , \5341_b1 , \5341_b0 , 
		\5342_b1 , \5342_b0 , \5343_b1 , \5343_b0 , \5344_b1 , \5344_b0 , \5345_b1 , \5345_b0 , \5346_b1 , \5346_b0 , 
		\5347_b1 , \5347_b0 , \5348_b1 , \5348_b0 , \5349_b1 , \5349_b0 , \5350_b1 , \5350_b0 , \5351_b1 , \5351_b0 , 
		\5352_b1 , \5352_b0 , \5353_b1 , \5353_b0 , \5354_b1 , \5354_b0 , \5355_b1 , \5355_b0 , \5356_b1 , \5356_b0 , 
		\5357_b1 , \5357_b0 , \5358_b1 , \5358_b0 , \5359_b1 , \5359_b0 , \5360_b1 , \5360_b0 , \5361_b1 , \5361_b0 , 
		\5362_b1 , \5362_b0 , \5363_b1 , \5363_b0 , \5364_b1 , \5364_b0 , \5365_b1 , \5365_b0 , \5366_b1 , \5366_b0 , 
		\5367_b1 , \5367_b0 , \5368_b1 , \5368_b0 , \5369_b1 , \5369_b0 , \5370_b1 , \5370_b0 , \5371_b1 , \5371_b0 , 
		\5372_b1 , \5372_b0 , \5373_b1 , \5373_b0 , \5374_b1 , \5374_b0 , \5375_b1 , \5375_b0 , \5376_b1 , \5376_b0 , 
		\5377_b1 , \5377_b0 , \5378_b1 , \5378_b0 , \5379_b1 , \5379_b0 , \5380_b1 , \5380_b0 , \5381_b1 , \5381_b0 , 
		\5382_b1 , \5382_b0 , \5383_b1 , \5383_b0 , \5384_b1 , \5384_b0 , \5385_b1 , \5385_b0 , \5386_b1 , \5386_b0 , 
		\5387_b1 , \5387_b0 , \5388_b1 , \5388_b0 , \5389_b1 , \5389_b0 , \5390_b1 , \5390_b0 , \5391_b1 , \5391_b0 , 
		\5392_b1 , \5392_b0 , \5393_b1 , \5393_b0 , \5394_b1 , \5394_b0 , \5395_b1 , \5395_b0 , \5396_b1 , \5396_b0 , 
		\5397_b1 , \5397_b0 , \5398_b1 , \5398_b0 , \5399_b1 , \5399_b0 , \5400_b1 , \5400_b0 , \5401_b1 , \5401_b0 , 
		\5402_b1 , \5402_b0 , \5403_b1 , \5403_b0 , \5404_b1 , \5404_b0 , \5405_b1 , \5405_b0 , \5406_b1 , \5406_b0 , 
		\5407_b1 , \5407_b0 , \5408_b1 , \5408_b0 , \5409_b1 , \5409_b0 , \5410_b1 , \5410_b0 , \5411_b1 , \5411_b0 , 
		\5412_b1 , \5412_b0 , \5413_b1 , \5413_b0 , \5414_b1 , \5414_b0 , \5415_b1 , \5415_b0 , \5416_b1 , \5416_b0 , 
		\5417_b1 , \5417_b0 , \5418_b1 , \5418_b0 , \5419_b1 , \5419_b0 , \5420_b1 , \5420_b0 , \5421_b1 , \5421_b0 , 
		\5422_b1 , \5422_b0 , \5423_b1 , \5423_b0 , \5424_b1 , \5424_b0 , \5425_b1 , \5425_b0 , \5426_b1 , \5426_b0 , 
		\5427_b1 , \5427_b0 , \5428_b1 , \5428_b0 , \5429_b1 , \5429_b0 , \5430_b1 , \5430_b0 , \5431_b1 , \5431_b0 , 
		\5432_b1 , \5432_b0 , \5433_b1 , \5433_b0 , \5434_b1 , \5434_b0 , \5435_b1 , \5435_b0 , \5436_b1 , \5436_b0 , 
		\5437_b1 , \5437_b0 , \5438_b1 , \5438_b0 , \5439_b1 , \5439_b0 , \5440_b1 , \5440_b0 , \5441_b1 , \5441_b0 , 
		\5442_b1 , \5442_b0 , \5443_b1 , \5443_b0 , \5444_b1 , \5444_b0 , \5445_b1 , \5445_b0 , \5446_b1 , \5446_b0 , 
		\5447_b1 , \5447_b0 , \5448_b1 , \5448_b0 , \5449_b1 , \5449_b0 , \5450_b1 , \5450_b0 , \5451_b1 , \5451_b0 , 
		\5452_b1 , \5452_b0 , \5453_b1 , \5453_b0 , \5454_b1 , \5454_b0 , \5455_b1 , \5455_b0 , \5456_b1 , \5456_b0 , 
		\5457_b1 , \5457_b0 , \5458_b1 , \5458_b0 , \5459_b1 , \5459_b0 , \5460_b1 , \5460_b0 , \5461_b1 , \5461_b0 , 
		\5462_b1 , \5462_b0 , \5463_b1 , \5463_b0 , \5464_b1 , \5464_b0 , \5465_b1 , \5465_b0 , \5466_b1 , \5466_b0 , 
		\5467_b1 , \5467_b0 , \5468_b1 , \5468_b0 , \5469_b1 , \5469_b0 , \5470_b1 , \5470_b0 , \5471_b1 , \5471_b0 , 
		\5472_b1 , \5472_b0 , \5473_b1 , \5473_b0 , \5474_b1 , \5474_b0 , \5475_b1 , \5475_b0 , \5476_b1 , \5476_b0 , 
		\5477_b1 , \5477_b0 , \5478_b1 , \5478_b0 , \5479_b1 , \5479_b0 , \5480_b1 , \5480_b0 , \5481_b1 , \5481_b0 , 
		\5482_b1 , \5482_b0 , \5483_b1 , \5483_b0 , \5484_b1 , \5484_b0 , \5485_b1 , \5485_b0 , \5486_b1 , \5486_b0 , 
		\5487_b1 , \5487_b0 , \5488_b1 , \5488_b0 , \5489_b1 , \5489_b0 , \5490_b1 , \5490_b0 , \5491_b1 , \5491_b0 , 
		\5492_b1 , \5492_b0 , \5493_b1 , \5493_b0 , \5494_b1 , \5494_b0 , \5495_b1 , \5495_b0 , \5496_b1 , \5496_b0 , 
		\5497_b1 , \5497_b0 , \5498_b1 , \5498_b0 , \5499_b1 , \5499_b0 , \5500_b1 , \5500_b0 , \5501_b1 , \5501_b0 , 
		\5502_b1 , \5502_b0 , \5503_b1 , \5503_b0 , \5504_b1 , \5504_b0 , \5505_b1 , \5505_b0 , \5506_b1 , \5506_b0 , 
		\5507_b1 , \5507_b0 , \5508_b1 , \5508_b0 , \5509_b1 , \5509_b0 , \5510_b1 , \5510_b0 , \5511_b1 , \5511_b0 , 
		\5512_b1 , \5512_b0 , \5513_b1 , \5513_b0 , \5514_b1 , \5514_b0 , \5515_b1 , \5515_b0 , \5516_b1 , \5516_b0 , 
		\5517_b1 , \5517_b0 , \5518_b1 , \5518_b0 , \5519_b1 , \5519_b0 , \5520_b1 , \5520_b0 , \5521_b1 , \5521_b0 , 
		\5522_b1 , \5522_b0 , \5523_b1 , \5523_b0 , \5524_b1 , \5524_b0 , \5525_b1 , \5525_b0 , \5526_b1 , \5526_b0 , 
		\5527_b1 , \5527_b0 , \5528_b1 , \5528_b0 , \5529_b1 , \5529_b0 , \5530_b1 , \5530_b0 , \5531_b1 , \5531_b0 , 
		\5532_b1 , \5532_b0 , \5533_b1 , \5533_b0 , \5534_b1 , \5534_b0 , \5535_b1 , \5535_b0 , \5536_b1 , \5536_b0 , 
		\5537_b1 , \5537_b0 , \5538_b1 , \5538_b0 , \5539_b1 , \5539_b0 , \5540_b1 , \5540_b0 , \5541_b1 , \5541_b0 , 
		\5542_b1 , \5542_b0 , \5543_b1 , \5543_b0 , \5544_b1 , \5544_b0 , \5545_b1 , \5545_b0 , \5546_b1 , \5546_b0 , 
		\5547_b1 , \5547_b0 , \5548_b1 , \5548_b0 , \5549_b1 , \5549_b0 , \5550_b1 , \5550_b0 , \5551_b1 , \5551_b0 , 
		\5552_b1 , \5552_b0 , \5553_b1 , \5553_b0 , \5554_b1 , \5554_b0 , \5555_b1 , \5555_b0 , \5556_b1 , \5556_b0 , 
		\5557_b1 , \5557_b0 , \5558_b1 , \5558_b0 , \5559_b1 , \5559_b0 , \5560_b1 , \5560_b0 , \5561_b1 , \5561_b0 , 
		\5562_b1 , \5562_b0 , \5563_b1 , \5563_b0 , \5564_b1 , \5564_b0 , \5565_b1 , \5565_b0 , \5566_b1 , \5566_b0 , 
		\5567_b1 , \5567_b0 , \5568_b1 , \5568_b0 , \5569_b1 , \5569_b0 , \5570_b1 , \5570_b0 , \5571_b1 , \5571_b0 , 
		\5572_b1 , \5572_b0 , \5573_b1 , \5573_b0 , \5574_b1 , \5574_b0 , \5575_b1 , \5575_b0 , \5576_b1 , \5576_b0 , 
		\5577_b1 , \5577_b0 , \5578_b1 , \5578_b0 , \5579_b1 , \5579_b0 , \5580_b1 , \5580_b0 , \5581_b1 , \5581_b0 , 
		\5582_b1 , \5582_b0 , \5583_b1 , \5583_b0 , \5584_b1 , \5584_b0 , \5585_b1 , \5585_b0 , \5586_b1 , \5586_b0 , 
		\5587_b1 , \5587_b0 , \5588_b1 , \5588_b0 , \5589_b1 , \5589_b0 , \5590_b1 , \5590_b0 , \5591_b1 , \5591_b0 , 
		\5592_b1 , \5592_b0 , \5593_b1 , \5593_b0 , \5594_b1 , \5594_b0 , \5595_b1 , \5595_b0 , \5596_b1 , \5596_b0 , 
		\5597_b1 , \5597_b0 , \5598_b1 , \5598_b0 , \5599_b1 , \5599_b0 , \5600_b1 , \5600_b0 , \5601_b1 , \5601_b0 , 
		\5602_b1 , \5602_b0 , \5603_b1 , \5603_b0 , \5604_b1 , \5604_b0 , \5605_b1 , \5605_b0 , \5606_b1 , \5606_b0 , 
		\5607_b1 , \5607_b0 , \5608_b1 , \5608_b0 , \5609_b1 , \5609_b0 , \5610_b1 , \5610_b0 , \5611_b1 , \5611_b0 , 
		\5612_b1 , \5612_b0 , \5613_b1 , \5613_b0 , \5614_b1 , \5614_b0 , \5615_b1 , \5615_b0 , \5616_b1 , \5616_b0 , 
		\5617_b1 , \5617_b0 , \5618_b1 , \5618_b0 , \5619_b1 , \5619_b0 , \5620_b1 , \5620_b0 , \5621_b1 , \5621_b0 , 
		\5622_b1 , \5622_b0 , \5623_b1 , \5623_b0 , \5624_b1 , \5624_b0 , \5625_b1 , \5625_b0 , \5626_b1 , \5626_b0 , 
		\5627_b1 , \5627_b0 , \5628_b1 , \5628_b0 , \5629_b1 , \5629_b0 , \5630_b1 , \5630_b0 , \5631_b1 , \5631_b0 , 
		\5632_b1 , \5632_b0 , \5633_b1 , \5633_b0 , \5634_b1 , \5634_b0 , \5635_b1 , \5635_b0 , \5636_b1 , \5636_b0 , 
		\5637_b1 , \5637_b0 , \5638_b1 , \5638_b0 , \5639_b1 , \5639_b0 , \5640_b1 , \5640_b0 , \5641_b1 , \5641_b0 , 
		\5642_b1 , \5642_b0 , \5643_b1 , \5643_b0 , \5644_b1 , \5644_b0 , \5645_b1 , \5645_b0 , \5646_b1 , \5646_b0 , 
		\5647_b1 , \5647_b0 , \5648_b1 , \5648_b0 , \5649_b1 , \5649_b0 , \5650_b1 , \5650_b0 , \5651_b1 , \5651_b0 , 
		\5652_b1 , \5652_b0 , \5653_b1 , \5653_b0 , \5654_b1 , \5654_b0 , \5655_b1 , \5655_b0 , \5656_b1 , \5656_b0 , 
		\5657_b1 , \5657_b0 , \5658_b1 , \5658_b0 , \5659_b1 , \5659_b0 , \5660_b1 , \5660_b0 , \5661_b1 , \5661_b0 , 
		\5662_b1 , \5662_b0 , \5663_b1 , \5663_b0 , \5664_b1 , \5664_b0 , \5665_b1 , \5665_b0 , \5666_b1 , \5666_b0 , 
		\5667_b1 , \5667_b0 , \5668_b1 , \5668_b0 , \5669_b1 , \5669_b0 , \5670_b1 , \5670_b0 , \5671_b1 , \5671_b0 , 
		\5672_b1 , \5672_b0 , \5673_b1 , \5673_b0 , \5674_b1 , \5674_b0 , \5675_b1 , \5675_b0 , \5676_b1 , \5676_b0 , 
		\5677_b1 , \5677_b0 , \5678_b1 , \5678_b0 , \5679_b1 , \5679_b0 , \5680_b1 , \5680_b0 , \5681_b1 , \5681_b0 , 
		\5682_b1 , \5682_b0 , \5683_b1 , \5683_b0 , \5684_b1 , \5684_b0 , \5685_b1 , \5685_b0 , \5686_b1 , \5686_b0 , 
		\5687_b1 , \5687_b0 , \5688_b1 , \5688_b0 , \5689_b1 , \5689_b0 , \5690_b1 , \5690_b0 , \5691_b1 , \5691_b0 , 
		\5692_b1 , \5692_b0 , \5693_b1 , \5693_b0 , \5694_b1 , \5694_b0 , \5695_b1 , \5695_b0 , \5696_b1 , \5696_b0 , 
		\5697_b1 , \5697_b0 , \5698_b1 , \5698_b0 , \5699_b1 , \5699_b0 , \5700_b1 , \5700_b0 , \5701_b1 , \5701_b0 , 
		\5702_b1 , \5702_b0 , \5703_b1 , \5703_b0 , \5704_b1 , \5704_b0 , \5705_b1 , \5705_b0 , \5706_b1 , \5706_b0 , 
		\5707_b1 , \5707_b0 , \5708_b1 , \5708_b0 , \5709_b1 , \5709_b0 , \5710_b1 , \5710_b0 , \5711_b1 , \5711_b0 , 
		\5712_b1 , \5712_b0 , \5713_b1 , \5713_b0 , \5714_b1 , \5714_b0 , \5715_b1 , \5715_b0 , \5716_b1 , \5716_b0 , 
		\5717_b1 , \5717_b0 , \5718_b1 , \5718_b0 , \5719_b1 , \5719_b0 , \5720_b1 , \5720_b0 , \5721_b1 , \5721_b0 , 
		\5722_b1 , \5722_b0 , \5723_b1 , \5723_b0 , \5724_b1 , \5724_b0 , \5725_b1 , \5725_b0 , \5726_b1 , \5726_b0 , 
		\5727_b1 , \5727_b0 , \5728_b1 , \5728_b0 , \5729_b1 , \5729_b0 , \5730_b1 , \5730_b0 , \5731_b1 , \5731_b0 , 
		\5732_b1 , \5732_b0 , \5733_b1 , \5733_b0 , \5734_b1 , \5734_b0 , \5735_b1 , \5735_b0 , \5736_b1 , \5736_b0 , 
		\5737_b1 , \5737_b0 , \5738_b1 , \5738_b0 , \5739_b1 , \5739_b0 , \5740_b1 , \5740_b0 , \5741_b1 , \5741_b0 , 
		\5742_b1 , \5742_b0 , \5743_b1 , \5743_b0 , \5744_b1 , \5744_b0 , \5745_b1 , \5745_b0 , \5746_b1 , \5746_b0 , 
		\5747_b1 , \5747_b0 , \5748_b1 , \5748_b0 , \5749_b1 , \5749_b0 , \5750_b1 , \5750_b0 , \5751_b1 , \5751_b0 , 
		\5752_b1 , \5752_b0 , \5753_b1 , \5753_b0 , \5754_b1 , \5754_b0 , \5755_b1 , \5755_b0 , \5756_b1 , \5756_b0 , 
		\5757_b1 , \5757_b0 , \5758_b1 , \5758_b0 , \5759_b1 , \5759_b0 , \5760_b1 , \5760_b0 , \5761_b1 , \5761_b0 , 
		\5762_b1 , \5762_b0 , \5763_b1 , \5763_b0 , \5764_b1 , \5764_b0 , \5765_b1 , \5765_b0 , \5766_b1 , \5766_b0 , 
		\5767_b1 , \5767_b0 , \5768_b1 , \5768_b0 , \5769_b1 , \5769_b0 , \5770_b1 , \5770_b0 , \5771_b1 , \5771_b0 , 
		\5772_b1 , \5772_b0 , \5773_b1 , \5773_b0 , \5774_b1 , \5774_b0 , \5775_b1 , \5775_b0 , \5776_b1 , \5776_b0 , 
		\5777_b1 , \5777_b0 , \5778_b1 , \5778_b0 , \5779_b1 , \5779_b0 , \5780_b1 , \5780_b0 , \5781_b1 , \5781_b0 , 
		\5782_b1 , \5782_b0 , \5783_b1 , \5783_b0 , \5784_b1 , \5784_b0 , \5785_b1 , \5785_b0 , \5786_b1 , \5786_b0 , 
		\5787_b1 , \5787_b0 , \5788_b1 , \5788_b0 , \5789_b1 , \5789_b0 , \5790_b1 , \5790_b0 , \5791_b1 , \5791_b0 , 
		\5792_b1 , \5792_b0 , \5793_b1 , \5793_b0 , \5794_b1 , \5794_b0 , \5795_b1 , \5795_b0 , \5796_b1 , \5796_b0 , 
		\5797_b1 , \5797_b0 , \5798_b1 , \5798_b0 , \5799_b1 , \5799_b0 , \5800_b1 , \5800_b0 , \5801_b1 , \5801_b0 , 
		\5802_b1 , \5802_b0 , \5803_b1 , \5803_b0 , \5804_b1 , \5804_b0 , \5805_b1 , \5805_b0 , \5806_b1 , \5806_b0 , 
		\5807_b1 , \5807_b0 , \5808_b1 , \5808_b0 , \5809_b1 , \5809_b0 , \5810_b1 , \5810_b0 , \5811_b1 , \5811_b0 , 
		\5812_b1 , \5812_b0 , \5813_b1 , \5813_b0 , \5814_b1 , \5814_b0 , \5815_b1 , \5815_b0 , \5816_b1 , \5816_b0 , 
		\5817_b1 , \5817_b0 , \5818_b1 , \5818_b0 , \5819_b1 , \5819_b0 , \5820_b1 , \5820_b0 , \5821_b1 , \5821_b0 , 
		\5822_b1 , \5822_b0 , \5823_b1 , \5823_b0 , \5824_b1 , \5824_b0 , \5825_b1 , \5825_b0 , \5826_b1 , \5826_b0 , 
		\5827_b1 , \5827_b0 , \5828_b1 , \5828_b0 , \5829_b1 , \5829_b0 , \5830_b1 , \5830_b0 , \5831_b1 , \5831_b0 , 
		\5832_b1 , \5832_b0 , \5833_b1 , \5833_b0 , \5834_b1 , \5834_b0 , \5835_b1 , \5835_b0 , \5836_b1 , \5836_b0 , 
		\5837_b1 , \5837_b0 , \5838_b1 , \5838_b0 , \5839_b1 , \5839_b0 , \5840_b1 , \5840_b0 , \5841_b1 , \5841_b0 , 
		\5842_b1 , \5842_b0 , \5843_b1 , \5843_b0 , \5844_b1 , \5844_b0 , \5845_b1 , \5845_b0 , \5846_b1 , \5846_b0 , 
		\5847_b1 , \5847_b0 , \5848_b1 , \5848_b0 , \5849_b1 , \5849_b0 , \5850_b1 , \5850_b0 , \5851_b1 , \5851_b0 , 
		\5852_b1 , \5852_b0 , \5853_b1 , \5853_b0 , \5854_b1 , \5854_b0 , \5855_b1 , \5855_b0 , \5856_b1 , \5856_b0 , 
		\5857_b1 , \5857_b0 , \5858_b1 , \5858_b0 , \5859_b1 , \5859_b0 , \5860_b1 , \5860_b0 , \5861_b1 , \5861_b0 , 
		\5862_b1 , \5862_b0 , \5863_b1 , \5863_b0 , \5864_b1 , \5864_b0 , \5865_b1 , \5865_b0 , \5866_b1 , \5866_b0 , 
		\5867_b1 , \5867_b0 , \5868_b1 , \5868_b0 , \5869_b1 , \5869_b0 , \5870_b1 , \5870_b0 , \5871_b1 , \5871_b0 , 
		\5872_b1 , \5872_b0 , \5873_b1 , \5873_b0 , \5874_b1 , \5874_b0 , \5875_b1 , \5875_b0 , \5876_b1 , \5876_b0 , 
		\5877_b1 , \5877_b0 , \5878_b1 , \5878_b0 , \5879_b1 , \5879_b0 , \5880_b1 , \5880_b0 , \5881_b1 , \5881_b0 , 
		\5882_b1 , \5882_b0 , \5883_b1 , \5883_b0 , \5884_b1 , \5884_b0 , \5885_b1 , \5885_b0 , \5886_b1 , \5886_b0 , 
		\5887_b1 , \5887_b0 , \5888_b1 , \5888_b0 , \5889_b1 , \5889_b0 , \5890_b1 , \5890_b0 , \5891_b1 , \5891_b0 , 
		\5892_b1 , \5892_b0 , \5893_b1 , \5893_b0 , \5894_b1 , \5894_b0 , \5895_b1 , \5895_b0 , \5896_b1 , \5896_b0 , 
		\5897_b1 , \5897_b0 , \5898_b1 , \5898_b0 , \5899_b1 , \5899_b0 , \5900_b1 , \5900_b0 , \5901_b1 , \5901_b0 , 
		\5902_b1 , \5902_b0 , \5903_b1 , \5903_b0 , \5904_b1 , \5904_b0 , \5905_b1 , \5905_b0 , \5906_b1 , \5906_b0 , 
		\5907_b1 , \5907_b0 , \5908_b1 , \5908_b0 , \5909_b1 , \5909_b0 , \5910_b1 , \5910_b0 , \5911_b1 , \5911_b0 , 
		\5912_b1 , \5912_b0 , \5913_b1 , \5913_b0 , \5914_b1 , \5914_b0 , \5915_b1 , \5915_b0 , \5916_b1 , \5916_b0 , 
		\5917_b1 , \5917_b0 , \5918_b1 , \5918_b0 , \5919_b1 , \5919_b0 , \5920_b1 , \5920_b0 , \5921_b1 , \5921_b0 , 
		\5922_b1 , \5922_b0 , \5923_b1 , \5923_b0 , \5924_b1 , \5924_b0 , \5925_b1 , \5925_b0 , \5926_b1 , \5926_b0 , 
		\5927_b1 , \5927_b0 , \5928_b1 , \5928_b0 , \5929_b1 , \5929_b0 , \5930_b1 , \5930_b0 , \5931_b1 , \5931_b0 , 
		\5932_b1 , \5932_b0 , \5933_b1 , \5933_b0 , \5934_b1 , \5934_b0 , \5935_b1 , \5935_b0 , \5936_b1 , \5936_b0 , 
		\5937_b1 , \5937_b0 , \5938_b1 , \5938_b0 , \5939_b1 , \5939_b0 , \5940_b1 , \5940_b0 , \5941_b1 , \5941_b0 , 
		\5942_b1 , \5942_b0 , \5943_b1 , \5943_b0 , \5944_b1 , \5944_b0 , \5945_b1 , \5945_b0 , \5946_b1 , \5946_b0 , 
		\5947_b1 , \5947_b0 , \5948_b1 , \5948_b0 , \5949_b1 , \5949_b0 , \5950_b1 , \5950_b0 , \5951_b1 , \5951_b0 , 
		\5952_b1 , \5952_b0 , \5953_b1 , \5953_b0 , \5954_b1 , \5954_b0 , \5955_b1 , \5955_b0 , \5956_b1 , \5956_b0 , 
		\5957_b1 , \5957_b0 , \5958_b1 , \5958_b0 , \5959_b1 , \5959_b0 , \5960_b1 , \5960_b0 , \5961_b1 , \5961_b0 , 
		\5962_b1 , \5962_b0 , \5963_b1 , \5963_b0 , \5964_b1 , \5964_b0 , \5965_b1 , \5965_b0 , \5966_b1 , \5966_b0 , 
		\5967_b1 , \5967_b0 , \5968_b1 , \5968_b0 , \5969_b1 , \5969_b0 , \5970_b1 , \5970_b0 , \5971_b1 , \5971_b0 , 
		\5972_b1 , \5972_b0 , \5973_b1 , \5973_b0 , \5974_b1 , \5974_b0 , \5975_b1 , \5975_b0 , \5976_b1 , \5976_b0 , 
		\5977_b1 , \5977_b0 , \5978_b1 , \5978_b0 , \5979_b1 , \5979_b0 , \5980_b1 , \5980_b0 , \5981_b1 , \5981_b0 , 
		\5982_b1 , \5982_b0 , \5983_b1 , \5983_b0 , \5984_b1 , \5984_b0 , \5985_b1 , \5985_b0 , \5986_b1 , \5986_b0 , 
		\5987_b1 , \5987_b0 , \5988_b1 , \5988_b0 , \5989_b1 , \5989_b0 , \5990_b1 , \5990_b0 , \5991_b1 , \5991_b0 , 
		\5992_b1 , \5992_b0 , \5993_b1 , \5993_b0 , \5994_b1 , \5994_b0 , \5995_b1 , \5995_b0 , \5996_b1 , \5996_b0 , 
		\5997_b1 , \5997_b0 , \5998_b1 , \5998_b0 , \5999_b1 , \5999_b0 , \6000_b1 , \6000_b0 , \6001_b1 , \6001_b0 , 
		\6002_b1 , \6002_b0 , \6003_b1 , \6003_b0 , \6004_b1 , \6004_b0 , \6005_b1 , \6005_b0 , \6006_b1 , \6006_b0 , 
		\6007_b1 , \6007_b0 , \6008_b1 , \6008_b0 , \6009_b1 , \6009_b0 , \6010_b1 , \6010_b0 , \6011_b1 , \6011_b0 , 
		\6012_b1 , \6012_b0 , \6013_b1 , \6013_b0 , \6014_b1 , \6014_b0 , \6015_b1 , \6015_b0 , \6016_b1 , \6016_b0 , 
		\6017_b1 , \6017_b0 , \6018_b1 , \6018_b0 , \6019_b1 , \6019_b0 , \6020_b1 , \6020_b0 , \6021_b1 , \6021_b0 , 
		\6022_b1 , \6022_b0 , \6023_b1 , \6023_b0 , \6024_b1 , \6024_b0 , \6025_b1 , \6025_b0 , \6026_b1 , \6026_b0 , 
		\6027_b1 , \6027_b0 , \6028_b1 , \6028_b0 , \6029_b1 , \6029_b0 , \6030_b1 , \6030_b0 , \6031_b1 , \6031_b0 , 
		\6032_b1 , \6032_b0 , \6033_b1 , \6033_b0 , \6034_b1 , \6034_b0 , \6035_b1 , \6035_b0 , \6036_b1 , \6036_b0 , 
		\6037_b1 , \6037_b0 , \6038_b1 , \6038_b0 , \6039_b1 , \6039_b0 , \6040_b1 , \6040_b0 , \6041_b1 , \6041_b0 , 
		\6042_b1 , \6042_b0 , \6043_b1 , \6043_b0 , \6044_b1 , \6044_b0 , \6045_b1 , \6045_b0 , \6046_b1 , \6046_b0 , 
		\6047_b1 , \6047_b0 , \6048_b1 , \6048_b0 , \6049_b1 , \6049_b0 , \6050_b1 , \6050_b0 , \6051_b1 , \6051_b0 , 
		\6052_b1 , \6052_b0 , \6053_b1 , \6053_b0 , \6054_b1 , \6054_b0 , \6055_b1 , \6055_b0 , \6056_b1 , \6056_b0 , 
		\6057_b1 , \6057_b0 , \6058_b1 , \6058_b0 , \6059_b1 , \6059_b0 , \6060_b1 , \6060_b0 , \6061_b1 , \6061_b0 , 
		\6062_b1 , \6062_b0 , \6063_b1 , \6063_b0 , \6064_b1 , \6064_b0 , \6065_b1 , \6065_b0 , \6066_b1 , \6066_b0 , 
		\6067_b1 , \6067_b0 , \6068_b1 , \6068_b0 , \6069_b1 , \6069_b0 , \6070_b1 , \6070_b0 , \6071_b1 , \6071_b0 , 
		\6072_b1 , \6072_b0 , \6073_b1 , \6073_b0 , \6074_b1 , \6074_b0 , \6075_b1 , \6075_b0 , \6076_b1 , \6076_b0 , 
		\6077_b1 , \6077_b0 , \6078_b1 , \6078_b0 , \6079_b1 , \6079_b0 , \6080_b1 , \6080_b0 , \6081_b1 , \6081_b0 , 
		\6082_b1 , \6082_b0 , \6083_b1 , \6083_b0 , \6084_b1 , \6084_b0 , \6085_b1 , \6085_b0 , \6086_b1 , \6086_b0 , 
		\6087_b1 , \6087_b0 , \6088_b1 , \6088_b0 , \6089_b1 , \6089_b0 , \6090_b1 , \6090_b0 , \6091_b1 , \6091_b0 , 
		\6092_b1 , \6092_b0 , \6093_b1 , \6093_b0 , \6094_b1 , \6094_b0 , \6095_b1 , \6095_b0 , \6096_b1 , \6096_b0 , 
		\6097_b1 , \6097_b0 , \6098_b1 , \6098_b0 , \6099_b1 , \6099_b0 , \6100_b1 , \6100_b0 , \6101_b1 , \6101_b0 , 
		\6102_b1 , \6102_b0 , \6103_b1 , \6103_b0 , \6104_b1 , \6104_b0 , \6105_b1 , \6105_b0 , \6106_b1 , \6106_b0 , 
		\6107_b1 , \6107_b0 , \6108_b1 , \6108_b0 , \6109_b1 , \6109_b0 , \6110_b1 , \6110_b0 , \6111_b1 , \6111_b0 , 
		\6112_b1 , \6112_b0 , \6113_b1 , \6113_b0 , \6114_b1 , \6114_b0 , \6115_b1 , \6115_b0 , \6116_b1 , \6116_b0 , 
		\6117_b1 , \6117_b0 , \6118_b1 , \6118_b0 , \6119_b1 , \6119_b0 , \6120_b1 , \6120_b0 , \6121_b1 , \6121_b0 , 
		\6122_b1 , \6122_b0 , \6123_b1 , \6123_b0 , \6124_b1 , \6124_b0 , \6125_b1 , \6125_b0 , \6126_b1 , \6126_b0 , 
		\6127_b1 , \6127_b0 , \6128_b1 , \6128_b0 , \6129_b1 , \6129_b0 , \6130_b1 , \6130_b0 , \6131_b1 , \6131_b0 , 
		\6132_b1 , \6132_b0 , \6133_b1 , \6133_b0 , \6134_b1 , \6134_b0 , \6135_b1 , \6135_b0 , \6136_b1 , \6136_b0 , 
		\6137_b1 , \6137_b0 , \6138_b1 , \6138_b0 , \6139_b1 , \6139_b0 , \6140_b1 , \6140_b0 , \6141_b1 , \6141_b0 , 
		\6142_b1 , \6142_b0 , \6143_b1 , \6143_b0 , \6144_b1 , \6144_b0 , \6145_b1 , \6145_b0 , \6146_b1 , \6146_b0 , 
		\6147_b1 , \6147_b0 , \6148_b1 , \6148_b0 , \6149_b1 , \6149_b0 , \6150_b1 , \6150_b0 , \6151_b1 , \6151_b0 , 
		\6152_b1 , \6152_b0 , \6153_b1 , \6153_b0 , \6154_b1 , \6154_b0 , \6155_b1 , \6155_b0 , \6156_b1 , \6156_b0 , 
		\6157_b1 , \6157_b0 , \6158_b1 , \6158_b0 , \6159_b1 , \6159_b0 , \6160_b1 , \6160_b0 , \6161_b1 , \6161_b0 , 
		\6162_b1 , \6162_b0 , \6163_b1 , \6163_b0 , \6164_b1 , \6164_b0 , \6165_b1 , \6165_b0 , \6166_b1 , \6166_b0 , 
		\6167_b1 , \6167_b0 , \6168_b1 , \6168_b0 , \6169_b1 , \6169_b0 , \6170_b1 , \6170_b0 , \6171_b1 , \6171_b0 , 
		\6172_b1 , \6172_b0 , \6173_b1 , \6173_b0 , \6174_b1 , \6174_b0 , \6175_b1 , \6175_b0 , \6176_b1 , \6176_b0 , 
		\6177_b1 , \6177_b0 , \6178_b1 , \6178_b0 , \6179_b1 , \6179_b0 , \6180_b1 , \6180_b0 , \6181_b1 , \6181_b0 , 
		\6182_b1 , \6182_b0 , \6183_b1 , \6183_b0 , \6184_b1 , \6184_b0 , \6185_b1 , \6185_b0 , \6186_b1 , \6186_b0 , 
		\6187_b1 , \6187_b0 , \6188_b1 , \6188_b0 , \6189_b1 , \6189_b0 , \6190_b1 , \6190_b0 , \6191_b1 , \6191_b0 , 
		\6192_b1 , \6192_b0 , \6193_b1 , \6193_b0 , \6194_b1 , \6194_b0 , \6195_b1 , \6195_b0 , \6196_b1 , \6196_b0 , 
		\6197_b1 , \6197_b0 , \6198_b1 , \6198_b0 , \6199_b1 , \6199_b0 , \6200_b1 , \6200_b0 , \6201_b1 , \6201_b0 , 
		\6202_b1 , \6202_b0 , \6203_b1 , \6203_b0 , \6204_b1 , \6204_b0 , \6205_b1 , \6205_b0 , \6206_b1 , \6206_b0 , 
		\6207_b1 , \6207_b0 , \6208_b1 , \6208_b0 , \6209_b1 , \6209_b0 , \6210_b1 , \6210_b0 , \6211_b1 , \6211_b0 , 
		\6212_b1 , \6212_b0 , \6213_b1 , \6213_b0 , \6214_b1 , \6214_b0 , \6215_b1 , \6215_b0 , \6216_b1 , \6216_b0 , 
		\6217_b1 , \6217_b0 , \6218_b1 , \6218_b0 , \6219_b1 , \6219_b0 , \6220_b1 , \6220_b0 , \6221_b1 , \6221_b0 , 
		\6222_b1 , \6222_b0 , \6223_b1 , \6223_b0 , \6224_b1 , \6224_b0 , \6225_b1 , \6225_b0 , \6226_b1 , \6226_b0 , 
		\6227_b1 , \6227_b0 , \6228_b1 , \6228_b0 , \6229_b1 , \6229_b0 , \6230_b1 , \6230_b0 , \6231_b1 , \6231_b0 , 
		\6232_b1 , \6232_b0 , \6233_b1 , \6233_b0 , \6234_b1 , \6234_b0 , \6235_b1 , \6235_b0 , \6236_b1 , \6236_b0 , 
		\6237_b1 , \6237_b0 , \6238_b1 , \6238_b0 , \6239_b1 , \6239_b0 , \6240_b1 , \6240_b0 , \6241_b1 , \6241_b0 , 
		\6242_b1 , \6242_b0 , \6243_b1 , \6243_b0 , \6244_b1 , \6244_b0 , \6245_b1 , \6245_b0 , \6246_b1 , \6246_b0 , 
		\6247_b1 , \6247_b0 , \6248_b1 , \6248_b0 , \6249_b1 , \6249_b0 , \6250_b1 , \6250_b0 , \6251_b1 , \6251_b0 , 
		\6252_b1 , \6252_b0 , \6253_b1 , \6253_b0 , \6254_b1 , \6254_b0 , \6255_b1 , \6255_b0 , \6256_b1 , \6256_b0 , 
		\6257_b1 , \6257_b0 , \6258_b1 , \6258_b0 , \6259_b1 , \6259_b0 , \6260_b1 , \6260_b0 , \6261_b1 , \6261_b0 , 
		\6262_b1 , \6262_b0 , \6263_b1 , \6263_b0 , \6264_b1 , \6264_b0 , \6265_b1 , \6265_b0 , \6266_b1 , \6266_b0 , 
		\6267_b1 , \6267_b0 , \6268_b1 , \6268_b0 , \6269_b1 , \6269_b0 , \6270_b1 , \6270_b0 , \6271_b1 , \6271_b0 , 
		\6272_b1 , \6272_b0 , \6273_b1 , \6273_b0 , \6274_b1 , \6274_b0 , \6275_b1 , \6275_b0 , \6276_b1 , \6276_b0 , 
		\6277_b1 , \6277_b0 , \6278_b1 , \6278_b0 , \6279_b1 , \6279_b0 , \6280_b1 , \6280_b0 , \6281_b1 , \6281_b0 , 
		\6282_b1 , \6282_b0 , \6283_b1 , \6283_b0 , \6284_b1 , \6284_b0 , \6285_b1 , \6285_b0 , \6286_b1 , \6286_b0 , 
		\6287_b1 , \6287_b0 , \6288_b1 , \6288_b0 , \6289_b1 , \6289_b0 , \6290_b1 , \6290_b0 , \6291_b1 , \6291_b0 , 
		\6292_b1 , \6292_b0 , \6293_b1 , \6293_b0 , \6294_b1 , \6294_b0 , \6295_b1 , \6295_b0 , \6296_b1 , \6296_b0 , 
		\6297_b1 , \6297_b0 , \6298_b1 , \6298_b0 , \6299_b1 , \6299_b0 , \6300_b1 , \6300_b0 , \6301_b1 , \6301_b0 , 
		\6302_b1 , \6302_b0 , \6303_b1 , \6303_b0 , \6304_b1 , \6304_b0 , \6305_b1 , \6305_b0 , \6306_b1 , \6306_b0 , 
		\6307_b1 , \6307_b0 , \6308_b1 , \6308_b0 , \6309_b1 , \6309_b0 , \6310_b1 , \6310_b0 , \6311_b1 , \6311_b0 , 
		\6312_b1 , \6312_b0 , \6313_b1 , \6313_b0 , \6314_b1 , \6314_b0 , \6315_b1 , \6315_b0 , \6316_b1 , \6316_b0 , 
		\6317_b1 , \6317_b0 , \6318_b1 , \6318_b0 , \6319_b1 , \6319_b0 , \6320_b1 , \6320_b0 , \6321_b1 , \6321_b0 , 
		\6322_b1 , \6322_b0 , \6323_b1 , \6323_b0 , \6324_b1 , \6324_b0 , \6325_b1 , \6325_b0 , \6326_b1 , \6326_b0 , 
		\6327_b1 , \6327_b0 , \6328_b1 , \6328_b0 , \6329_b1 , \6329_b0 , \6330_b1 , \6330_b0 , \6331_b1 , \6331_b0 , 
		\6332_b1 , \6332_b0 , \6333_b1 , \6333_b0 , \6334_b1 , \6334_b0 , \6335_b1 , \6335_b0 , \6336_b1 , \6336_b0 , 
		\6337_b1 , \6337_b0 , \6338_b1 , \6338_b0 , \6339_b1 , \6339_b0 , \6340_b1 , \6340_b0 , \6341_b1 , \6341_b0 , 
		\6342_b1 , \6342_b0 , \6343_b1 , \6343_b0 , \6344_b1 , \6344_b0 , \6345_b1 , \6345_b0 , \6346_b1 , \6346_b0 , 
		\6347_b1 , \6347_b0 , \6348_b1 , \6348_b0 , \6349_b1 , \6349_b0 , \6350_b1 , \6350_b0 , \6351_b1 , \6351_b0 , 
		\6352_b1 , \6352_b0 , \6353_b1 , \6353_b0 , \6354_b1 , \6354_b0 , \6355_b1 , \6355_b0 , \6356_b1 , \6356_b0 , 
		\6357_b1 , \6357_b0 , \6358_b1 , \6358_b0 , \6359_b1 , \6359_b0 , \6360_b1 , \6360_b0 , \6361_b1 , \6361_b0 , 
		\6362_b1 , \6362_b0 , \6363_b1 , \6363_b0 , \6364_b1 , \6364_b0 , \6365_b1 , \6365_b0 , \6366_b1 , \6366_b0 , 
		\6367_b1 , \6367_b0 , \6368_b1 , \6368_b0 , \6369_b1 , \6369_b0 , \6370_b1 , \6370_b0 , \6371_b1 , \6371_b0 , 
		\6372_b1 , \6372_b0 , \6373_b1 , \6373_b0 , \6374_b1 , \6374_b0 , \6375_b1 , \6375_b0 , \6376_b1 , \6376_b0 , 
		\6377_b1 , \6377_b0 , \6378_b1 , \6378_b0 , \6379_b1 , \6379_b0 , \6380_b1 , \6380_b0 , \6381_b1 , \6381_b0 , 
		\6382_b1 , \6382_b0 , \6383_b1 , \6383_b0 , \6384_b1 , \6384_b0 , \6385_b1 , \6385_b0 , \6386_b1 , \6386_b0 , 
		\6387_b1 , \6387_b0 , \6388_b1 , \6388_b0 , \6389_b1 , \6389_b0 , \6390_b1 , \6390_b0 , \6391_b1 , \6391_b0 , 
		\6392_b1 , \6392_b0 , \6393_b1 , \6393_b0 , \6394_b1 , \6394_b0 , \6395_b1 , \6395_b0 , \6396_b1 , \6396_b0 , 
		\6397_b1 , \6397_b0 , \6398_b1 , \6398_b0 , \6399_b1 , \6399_b0 , \6400_b1 , \6400_b0 , \6401_b1 , \6401_b0 , 
		\6402_b1 , \6402_b0 , \6403_b1 , \6403_b0 , \6404_b1 , \6404_b0 , \6405_b1 , \6405_b0 , \6406_b1 , \6406_b0 , 
		\6407_b1 , \6407_b0 , \6408_b1 , \6408_b0 , \6409_b1 , \6409_b0 , \6410_b1 , \6410_b0 , \6411_b1 , \6411_b0 , 
		\6412_b1 , \6412_b0 , \6413_b1 , \6413_b0 , \6414_b1 , \6414_b0 , \6415_b1 , \6415_b0 , \6416_b1 , \6416_b0 , 
		\6417_b1 , \6417_b0 , \6418_b1 , \6418_b0 , \6419_b1 , \6419_b0 , \6420_b1 , \6420_b0 , \6421_b1 , \6421_b0 , 
		\6422_b1 , \6422_b0 , \6423_b1 , \6423_b0 , \6424_b1 , \6424_b0 , \6425_b1 , \6425_b0 , \6426_b1 , \6426_b0 , 
		\6427_b1 , \6427_b0 , \6428_b1 , \6428_b0 , \6429_b1 , \6429_b0 , \6430_b1 , \6430_b0 , \6431_b1 , \6431_b0 , 
		\6432_b1 , \6432_b0 , \6433_b1 , \6433_b0 , \6434_b1 , \6434_b0 , \6435_b1 , \6435_b0 , \6436_b1 , \6436_b0 , 
		\6437_b1 , \6437_b0 , \6438_b1 , \6438_b0 , \6439_b1 , \6439_b0 , \6440_b1 , \6440_b0 , \6441_b1 , \6441_b0 , 
		\6442_b1 , \6442_b0 , \6443_b1 , \6443_b0 , \6444_b1 , \6444_b0 , \6445_b1 , \6445_b0 , \6446_b1 , \6446_b0 , 
		\6447_b1 , \6447_b0 , \6448_b1 , \6448_b0 , \6449_b1 , \6449_b0 , \6450_b1 , \6450_b0 , \6451_b1 , \6451_b0 , 
		\6452_b1 , \6452_b0 , \6453_b1 , \6453_b0 , \6454_b1 , \6454_b0 , \6455_b1 , \6455_b0 , \6456_b1 , \6456_b0 , 
		\6457_b1 , \6457_b0 , \6458_b1 , \6458_b0 , \6459_b1 , \6459_b0 , \6460_b1 , \6460_b0 , \6461_b1 , \6461_b0 , 
		\6462_b1 , \6462_b0 , \6463_b1 , \6463_b0 , \6464_b1 , \6464_b0 , \6465_b1 , \6465_b0 , \6466_b1 , \6466_b0 , 
		\6467_b1 , \6467_b0 , \6468_b1 , \6468_b0 , \6469_b1 , \6469_b0 , \6470_b1 , \6470_b0 , \6471_b1 , \6471_b0 , 
		\6472_b1 , \6472_b0 , \6473_b1 , \6473_b0 , \6474_b1 , \6474_b0 , \6475_b1 , \6475_b0 , \6476_b1 , \6476_b0 , 
		\6477_b1 , \6477_b0 , \6478_b1 , \6478_b0 , \6479_b1 , \6479_b0 , \6480_b1 , \6480_b0 , \6481_b1 , \6481_b0 , 
		\6482_b1 , \6482_b0 , \6483_b1 , \6483_b0 , \6484_b1 , \6484_b0 , \6485_b1 , \6485_b0 , \6486_b1 , \6486_b0 , 
		\6487_b1 , \6487_b0 , \6488_b1 , \6488_b0 , \6489_b1 , \6489_b0 , \6490_b1 , \6490_b0 , \6491_b1 , \6491_b0 , 
		\6492_b1 , \6492_b0 , \6493_b1 , \6493_b0 , \6494_b1 , \6494_b0 , \6495_b1 , \6495_b0 , \6496_b1 , \6496_b0 , 
		\6497_b1 , \6497_b0 , \6498_b1 , \6498_b0 , \6499_b1 , \6499_b0 , \6500_b1 , \6500_b0 , \6501_b1 , \6501_b0 , 
		\6502_b1 , \6502_b0 , \6503_b1 , \6503_b0 , \6504_b1 , \6504_b0 , \6505_b1 , \6505_b0 , \6506_b1 , \6506_b0 , 
		\6507_b1 , \6507_b0 , \6508_b1 , \6508_b0 , \6509_b1 , \6509_b0 , \6510_b1 , \6510_b0 , \6511_b1 , \6511_b0 , 
		\6512_b1 , \6512_b0 , \6513_b1 , \6513_b0 , \6514_b1 , \6514_b0 , \6515_b1 , \6515_b0 , \6516_b1 , \6516_b0 , 
		\6517_b1 , \6517_b0 , \6518_b1 , \6518_b0 , \6519_b1 , \6519_b0 , \6520_b1 , \6520_b0 , \6521_b1 , \6521_b0 , 
		\6522_b1 , \6522_b0 , \6523_b1 , \6523_b0 , \6524_b1 , \6524_b0 , \6525_b1 , \6525_b0 , \6526_b1 , \6526_b0 , 
		\6527_b1 , \6527_b0 , \6528_b1 , \6528_b0 , \6529_b1 , \6529_b0 , \6530_b1 , \6530_b0 , \6531_b1 , \6531_b0 , 
		\6532_b1 , \6532_b0 , \6533_b1 , \6533_b0 , \6534_b1 , \6534_b0 , \6535_b1 , \6535_b0 , \6536_b1 , \6536_b0 , 
		\6537_b1 , \6537_b0 , \6538_b1 , \6538_b0 , \6539_b1 , \6539_b0 , \6540_b1 , \6540_b0 , \6541_b1 , \6541_b0 , 
		\6542_b1 , \6542_b0 , \6543_b1 , \6543_b0 , \6544_b1 , \6544_b0 , \6545_b1 , \6545_b0 , \6546_b1 , \6546_b0 , 
		\6547_b1 , \6547_b0 , \6548_b1 , \6548_b0 , \6549_b1 , \6549_b0 , \6550_b1 , \6550_b0 , \6551_b1 , \6551_b0 , 
		\6552_b1 , \6552_b0 , \6553_b1 , \6553_b0 , \6554_b1 , \6554_b0 , \6555_b1 , \6555_b0 , \6556_b1 , \6556_b0 , 
		\6557_b1 , \6557_b0 , \6558_b1 , \6558_b0 , \6559_b1 , \6559_b0 , \6560_b1 , \6560_b0 , \6561_b1 , \6561_b0 , 
		\6562_b1 , \6562_b0 , \6563_b1 , \6563_b0 , \6564_b1 , \6564_b0 , \6565_b1 , \6565_b0 , \6566_b1 , \6566_b0 , 
		\6567_b1 , \6567_b0 , \6568_b1 , \6568_b0 , \6569_b1 , \6569_b0 , \6570_b1 , \6570_b0 , \6571_b1 , \6571_b0 , 
		\6572_b1 , \6572_b0 , \6573_b1 , \6573_b0 , \6574_b1 , \6574_b0 , \6575_b1 , \6575_b0 , \6576_b1 , \6576_b0 , 
		\6577_b1 , \6577_b0 , \6578_b1 , \6578_b0 , \6579_b1 , \6579_b0 , \6580_b1 , \6580_b0 , \6581_b1 , \6581_b0 , 
		\6582_b1 , \6582_b0 , \6583_b1 , \6583_b0 , \6584_b1 , \6584_b0 , \6585_b1 , \6585_b0 , \6586_b1 , \6586_b0 , 
		\6587_b1 , \6587_b0 , \6588_b1 , \6588_b0 , \6589_b1 , \6589_b0 , \6590_b1 , \6590_b0 , \6591_b1 , \6591_b0 , 
		\6592_b1 , \6592_b0 , \6593_b1 , \6593_b0 , \6594_b1 , \6594_b0 , \6595_b1 , \6595_b0 , \6596_b1 , \6596_b0 , 
		\6597_b1 , \6597_b0 , \6598_b1 , \6598_b0 , \6599_b1 , \6599_b0 , \6600_b1 , \6600_b0 , \6601_b1 , \6601_b0 , 
		\6602_b1 , \6602_b0 , \6603_b1 , \6603_b0 , \6604_b1 , \6604_b0 , \6605_b1 , \6605_b0 , \6606_b1 , \6606_b0 , 
		\6607_b1 , \6607_b0 , \6608_b1 , \6608_b0 , \6609_b1 , \6609_b0 , \6610_b1 , \6610_b0 , \6611_b1 , \6611_b0 , 
		\6612_b1 , \6612_b0 , \6613_b1 , \6613_b0 , \6614_b1 , \6614_b0 , \6615_b1 , \6615_b0 , \6616_b1 , \6616_b0 , 
		\6617_b1 , \6617_b0 , \6618_b1 , \6618_b0 , \6619_b1 , \6619_b0 , \6620_b1 , \6620_b0 , \6621_b1 , \6621_b0 , 
		\6622_b1 , \6622_b0 , \6623_b1 , \6623_b0 , \6624_b1 , \6624_b0 , \6625_b1 , \6625_b0 , \6626_b1 , \6626_b0 , 
		\6627_b1 , \6627_b0 , \6628_b1 , \6628_b0 , \6629_b1 , \6629_b0 , \6630_b1 , \6630_b0 , \6631_b1 , \6631_b0 , 
		\6632_b1 , \6632_b0 , \6633_b1 , \6633_b0 , \6634_b1 , \6634_b0 , \6635_b1 , \6635_b0 , \6636_b1 , \6636_b0 , 
		\6637_b1 , \6637_b0 , \6638_b1 , \6638_b0 , \6639_b1 , \6639_b0 , \6640_b1 , \6640_b0 , \6641_b1 , \6641_b0 , 
		\6642_b1 , \6642_b0 , \6643_b1 , \6643_b0 , \6644_b1 , \6644_b0 , \6645_b1 , \6645_b0 , \6646_b1 , \6646_b0 , 
		\6647_b1 , \6647_b0 , \6648_b1 , \6648_b0 , \6649_b1 , \6649_b0 , \6650_b1 , \6650_b0 , \6651_b1 , \6651_b0 , 
		\6652_b1 , \6652_b0 , \6653_b1 , \6653_b0 , \6654_b1 , \6654_b0 , \6655_b1 , \6655_b0 , \6656_b1 , \6656_b0 , 
		\6657_b1 , \6657_b0 , \6658_b1 , \6658_b0 , \6659_b1 , \6659_b0 , \6660_b1 , \6660_b0 , \6661_b1 , \6661_b0 , 
		\6662_b1 , \6662_b0 , \6663_b1 , \6663_b0 , \6664_b1 , \6664_b0 , \6665_b1 , \6665_b0 , \6666_b1 , \6666_b0 , 
		\6667_b1 , \6667_b0 , \6668_b1 , \6668_b0 , \6669_b1 , \6669_b0 , \6670_b1 , \6670_b0 , \6671_b1 , \6671_b0 , 
		\6672_b1 , \6672_b0 , \6673_b1 , \6673_b0 , \6674_b1 , \6674_b0 , \6675_b1 , \6675_b0 , \6676_b1 , \6676_b0 , 
		\6677_b1 , \6677_b0 , \6678_b1 , \6678_b0 , \6679_b1 , \6679_b0 , \6680_b1 , \6680_b0 , \6681_b1 , \6681_b0 , 
		\6682_b1 , \6682_b0 , \6683_b1 , \6683_b0 , \6684_b1 , \6684_b0 , \6685_b1 , \6685_b0 , \6686_b1 , \6686_b0 , 
		\6687_b1 , \6687_b0 , \6688_b1 , \6688_b0 , \6689_b1 , \6689_b0 , \6690_b1 , \6690_b0 , \6691_b1 , \6691_b0 , 
		\6692_b1 , \6692_b0 , \6693_b1 , \6693_b0 , \6694_b1 , \6694_b0 , \6695_b1 , \6695_b0 , \6696_b1 , \6696_b0 , 
		\6697_b1 , \6697_b0 , \6698_b1 , \6698_b0 , \6699_b1 , \6699_b0 , \6700_b1 , \6700_b0 , \6701_b1 , \6701_b0 , 
		\6702_b1 , \6702_b0 , \6703_b1 , \6703_b0 , \6704_b1 , \6704_b0 , \6705_b1 , \6705_b0 , \6706_b1 , \6706_b0 , 
		\6707_b1 , \6707_b0 , \6708_b1 , \6708_b0 , \6709_b1 , \6709_b0 , \6710_b1 , \6710_b0 , \6711_b1 , \6711_b0 , 
		\6712_b1 , \6712_b0 , \6713_b1 , \6713_b0 , \6714_b1 , \6714_b0 , \6715_b1 , \6715_b0 , \6716_b1 , \6716_b0 , 
		\6717_b1 , \6717_b0 , \6718_b1 , \6718_b0 , \6719_b1 , \6719_b0 , \6720_b1 , \6720_b0 , \6721_b1 , \6721_b0 , 
		\6722_b1 , \6722_b0 , \6723_b1 , \6723_b0 , \6724_b1 , \6724_b0 , \6725_b1 , \6725_b0 , \6726_b1 , \6726_b0 , 
		\6727_b1 , \6727_b0 , \6728_b1 , \6728_b0 , \6729_b1 , \6729_b0 , \6730_b1 , \6730_b0 , \6731_b1 , \6731_b0 , 
		\6732_b1 , \6732_b0 , \6733_b1 , \6733_b0 , \6734_b1 , \6734_b0 , \6735_b1 , \6735_b0 , \6736_b1 , \6736_b0 , 
		\6737_b1 , \6737_b0 , \6738_b1 , \6738_b0 , \6739_b1 , \6739_b0 , \6740_b1 , \6740_b0 , \6741_b1 , \6741_b0 , 
		\6742_b1 , \6742_b0 , \6743_b1 , \6743_b0 , \6744_b1 , \6744_b0 , \6745_b1 , \6745_b0 , \6746_b1 , \6746_b0 , 
		\6747_b1 , \6747_b0 , \6748_b1 , \6748_b0 , \6749_b1 , \6749_b0 , \6750_b1 , \6750_b0 , \6751_b1 , \6751_b0 , 
		\6752_b1 , \6752_b0 , \6753_b1 , \6753_b0 , \6754_b1 , \6754_b0 , \6755_b1 , \6755_b0 , \6756_b1 , \6756_b0 , 
		\6757_b1 , \6757_b0 , \6758_b1 , \6758_b0 , \6759_b1 , \6759_b0 , \6760_b1 , \6760_b0 , \6761_b1 , \6761_b0 , 
		\6762_b1 , \6762_b0 , \6763_b1 , \6763_b0 , \6764_b1 , \6764_b0 , \6765_b1 , \6765_b0 , \6766_b1 , \6766_b0 , 
		\6767_b1 , \6767_b0 , \6768_b1 , \6768_b0 , \6769_b1 , \6769_b0 , \6770_b1 , \6770_b0 , \6771_b1 , \6771_b0 , 
		\6772_b1 , \6772_b0 , \6773_b1 , \6773_b0 , \6774_b1 , \6774_b0 , \6775_b1 , \6775_b0 , \6776_b1 , \6776_b0 , 
		\6777_b1 , \6777_b0 , \6778_b1 , \6778_b0 , \6779_b1 , \6779_b0 , \6780_b1 , \6780_b0 , \6781_b1 , \6781_b0 , 
		\6782_b1 , \6782_b0 , \6783_b1 , \6783_b0 , \6784_b1 , \6784_b0 , \6785_b1 , \6785_b0 , \6786_b1 , \6786_b0 , 
		\6787_b1 , \6787_b0 , \6788_b1 , \6788_b0 , \6789_b1 , \6789_b0 , \6790_b1 , \6790_b0 , \6791_b1 , \6791_b0 , 
		\6792_b1 , \6792_b0 , \6793_b1 , \6793_b0 , \6794_b1 , \6794_b0 , \6795_b1 , \6795_b0 , \6796_b1 , \6796_b0 , 
		\6797_b1 , \6797_b0 , \6798_b1 , \6798_b0 , \6799_b1 , \6799_b0 , \6800_b1 , \6800_b0 , \6801_b1 , \6801_b0 , 
		\6802_b1 , \6802_b0 , \6803_b1 , \6803_b0 , \6804_b1 , \6804_b0 , \6805_b1 , \6805_b0 , \6806_b1 , \6806_b0 , 
		\6807_b1 , \6807_b0 , \6808_b1 , \6808_b0 , \6809_b1 , \6809_b0 , \6810_b1 , \6810_b0 , \6811_b1 , \6811_b0 , 
		\6812_b1 , \6812_b0 , \6813_b1 , \6813_b0 , \6814_b1 , \6814_b0 , \6815_b1 , \6815_b0 , \6816_b1 , \6816_b0 , 
		\6817_b1 , \6817_b0 , \6818_b1 , \6818_b0 , \6819_b1 , \6819_b0 , \6820_b1 , \6820_b0 , \6821_b1 , \6821_b0 , 
		\6822_b1 , \6822_b0 , \6823_b1 , \6823_b0 , \6824_b1 , \6824_b0 , \6825_b1 , \6825_b0 , \6826_b1 , \6826_b0 , 
		\6827_b1 , \6827_b0 , \6828_b1 , \6828_b0 , \6829_b1 , \6829_b0 , \6830_b1 , \6830_b0 , \6831_b1 , \6831_b0 , 
		\6832_b1 , \6832_b0 , \6833_b1 , \6833_b0 , \6834_b1 , \6834_b0 , \6835_b1 , \6835_b0 , \6836_b1 , \6836_b0 , 
		\6837_b1 , \6837_b0 , \6838_b1 , \6838_b0 , \6839_b1 , \6839_b0 , \6840_b1 , \6840_b0 , \6841_b1 , \6841_b0 , 
		\6842_b1 , \6842_b0 , \6843_b1 , \6843_b0 , \6844_b1 , \6844_b0 , \6845_b1 , \6845_b0 , \6846_b1 , \6846_b0 , 
		\6847_b1 , \6847_b0 , \6848_b1 , \6848_b0 , \6849_b1 , \6849_b0 , \6850_b1 , \6850_b0 , \6851_b1 , \6851_b0 , 
		\6852_b1 , \6852_b0 , \6853_b1 , \6853_b0 , \6854_b1 , \6854_b0 , \6855_b1 , \6855_b0 , \6856_b1 , \6856_b0 , 
		\6857_b1 , \6857_b0 , \6858_b1 , \6858_b0 , \6859_b1 , \6859_b0 , \6860_b1 , \6860_b0 , \6861_b1 , \6861_b0 , 
		\6862_b1 , \6862_b0 , \6863_b1 , \6863_b0 , \6864_b1 , \6864_b0 , \6865_b1 , \6865_b0 , \6866_b1 , \6866_b0 , 
		\6867_b1 , \6867_b0 , \6868_b1 , \6868_b0 , \6869_b1 , \6869_b0 , \6870_b1 , \6870_b0 , \6871_b1 , \6871_b0 , 
		\6872_b1 , \6872_b0 , \6873_b1 , \6873_b0 , \6874_b1 , \6874_b0 , \6875_b1 , \6875_b0 , \6876_b1 , \6876_b0 , 
		\6877_b1 , \6877_b0 , \6878_b1 , \6878_b0 , \6879_b1 , \6879_b0 , \6880_b1 , \6880_b0 , \6881_b1 , \6881_b0 , 
		\6882_b1 , \6882_b0 , \6883_b1 , \6883_b0 , \6884_b1 , \6884_b0 , \6885_b1 , \6885_b0 , \6886_b1 , \6886_b0 , 
		\6887_b1 , \6887_b0 , \6888_b1 , \6888_b0 , \6889_b1 , \6889_b0 , \6890_b1 , \6890_b0 , \6891_b1 , \6891_b0 , 
		\6892_b1 , \6892_b0 , \6893_b1 , \6893_b0 , \6894_b1 , \6894_b0 , \6895_b1 , \6895_b0 , \6896_b1 , \6896_b0 , 
		\6897_b1 , \6897_b0 , \6898_b1 , \6898_b0 , \6899_b1 , \6899_b0 , \6900_b1 , \6900_b0 , \6901_b1 , \6901_b0 , 
		\6902_b1 , \6902_b0 , \6903_b1 , \6903_b0 , \6904_b1 , \6904_b0 , \6905_b1 , \6905_b0 , \6906_b1 , \6906_b0 , 
		\6907_b1 , \6907_b0 , \6908_b1 , \6908_b0 , \6909_b1 , \6909_b0 , \6910_b1 , \6910_b0 , \6911_b1 , \6911_b0 , 
		\6912_b1 , \6912_b0 , \6913_b1 , \6913_b0 , \6914_b1 , \6914_b0 , \6915_b1 , \6915_b0 , \6916_b1 , \6916_b0 , 
		\6917_b1 , \6917_b0 , \6918_b1 , \6918_b0 , \6919_b1 , \6919_b0 , \6920_b1 , \6920_b0 , \6921_b1 , \6921_b0 , 
		\6922_b1 , \6922_b0 , \6923_b1 , \6923_b0 , \6924_b1 , \6924_b0 , \6925_b1 , \6925_b0 , \6926_b1 , \6926_b0 , 
		\6927_b1 , \6927_b0 , \6928_b1 , \6928_b0 , \6929_b1 , \6929_b0 , \6930_b1 , \6930_b0 , \6931_b1 , \6931_b0 , 
		\6932_b1 , \6932_b0 , \6933_b1 , \6933_b0 , \6934_b1 , \6934_b0 , \6935_b1 , \6935_b0 , \6936_b1 , \6936_b0 , 
		\6937_b1 , \6937_b0 , \6938_b1 , \6938_b0 , \6939_b1 , \6939_b0 , \6940_b1 , \6940_b0 , \6941_b1 , \6941_b0 , 
		\6942_b1 , \6942_b0 , \6943_b1 , \6943_b0 , \6944_b1 , \6944_b0 , \6945_b1 , \6945_b0 , \6946_b1 , \6946_b0 , 
		\6947_b1 , \6947_b0 , \6948_b1 , \6948_b0 , \6949_b1 , \6949_b0 , \6950_b1 , \6950_b0 , \6951_b1 , \6951_b0 , 
		\6952_b1 , \6952_b0 , \6953_b1 , \6953_b0 , \6954_b1 , \6954_b0 , \6955_b1 , \6955_b0 , \6956_b1 , \6956_b0 , 
		\6957_b1 , \6957_b0 , \6958_b1 , \6958_b0 , \6959_b1 , \6959_b0 , \6960_b1 , \6960_b0 , \6961_b1 , \6961_b0 , 
		\6962_b1 , \6962_b0 , \6963_b1 , \6963_b0 , \6964_b1 , \6964_b0 , \6965_b1 , \6965_b0 , \6966_b1 , \6966_b0 , 
		\6967_b1 , \6967_b0 , \6968_b1 , \6968_b0 , \6969_b1 , \6969_b0 , \6970_b1 , \6970_b0 , \6971_b1 , \6971_b0 , 
		\6972_b1 , \6972_b0 , \6973_b1 , \6973_b0 , \6974_b1 , \6974_b0 , \6975_b1 , \6975_b0 , \6976_b1 , \6976_b0 , 
		\6977_b1 , \6977_b0 , \6978_b1 , \6978_b0 , \6979_b1 , \6979_b0 , \6980_b1 , \6980_b0 , \6981_b1 , \6981_b0 , 
		\6982_b1 , \6982_b0 , \6983_b1 , \6983_b0 , \6984_b1 , \6984_b0 , \6985_b1 , \6985_b0 , \6986_b1 , \6986_b0 , 
		\6987_b1 , \6987_b0 , \6988_b1 , \6988_b0 , \6989_b1 , \6989_b0 , \6990_b1 , \6990_b0 , \6991_b1 , \6991_b0 , 
		\6992_b1 , \6992_b0 , \6993_b1 , \6993_b0 , \6994_b1 , \6994_b0 , \6995_b1 , \6995_b0 , \6996_b1 , \6996_b0 , 
		\6997_b1 , \6997_b0 , \6998_b1 , \6998_b0 , \6999_b1 , \6999_b0 , \7000_b1 , \7000_b0 , \7001_b1 , \7001_b0 , 
		\7002_b1 , \7002_b0 , \7003_b1 , \7003_b0 , \7004_b1 , \7004_b0 , \7005_b1 , \7005_b0 , \7006_b1 , \7006_b0 , 
		\7007_b1 , \7007_b0 , \7008_b1 , \7008_b0 , \7009_b1 , \7009_b0 , \7010_b1 , \7010_b0 , \7011_b1 , \7011_b0 , 
		\7012_b1 , \7012_b0 , \7013_b1 , \7013_b0 , \7014_b1 , \7014_b0 , \7015_b1 , \7015_b0 , \7016_b1 , \7016_b0 , 
		\7017_b1 , \7017_b0 , \7018_b1 , \7018_b0 , \7019_b1 , \7019_b0 , \7020_b1 , \7020_b0 , \7021_b1 , \7021_b0 , 
		\7022_b1 , \7022_b0 , \7023_b1 , \7023_b0 , \7024_b1 , \7024_b0 , \7025_b1 , \7025_b0 , \7026_b1 , \7026_b0 , 
		\7027_b1 , \7027_b0 , \7028_b1 , \7028_b0 , \7029_b1 , \7029_b0 , \7030_b1 , \7030_b0 , \7031_b1 , \7031_b0 , 
		\7032_b1 , \7032_b0 , \7033_b1 , \7033_b0 , \7034_b1 , \7034_b0 , \7035_b1 , \7035_b0 , \7036_b1 , \7036_b0 , 
		\7037_b1 , \7037_b0 , \7038_b1 , \7038_b0 , \7039_b1 , \7039_b0 , \7040_b1 , \7040_b0 , \7041_b1 , \7041_b0 , 
		\7042_b1 , \7042_b0 , \7043_b1 , \7043_b0 , \7044_b1 , \7044_b0 , \7045_b1 , \7045_b0 , \7046_b1 , \7046_b0 , 
		\7047_b1 , \7047_b0 , \7048_b1 , \7048_b0 , \7049_b1 , \7049_b0 , \7050_b1 , \7050_b0 , \7051_b1 , \7051_b0 , 
		\7052_b1 , \7052_b0 , \7053_b1 , \7053_b0 , \7054_b1 , \7054_b0 , \7055_b1 , \7055_b0 , \7056_b1 , \7056_b0 , 
		\7057_b1 , \7057_b0 , \7058_b1 , \7058_b0 , \7059_b1 , \7059_b0 , \7060_b1 , \7060_b0 , \7061_b1 , \7061_b0 , 
		\7062_b1 , \7062_b0 , \7063_b1 , \7063_b0 , \7064_b1 , \7064_b0 , \7065_b1 , \7065_b0 , \7066_b1 , \7066_b0 , 
		\7067_b1 , \7067_b0 , \7068_b1 , \7068_b0 , \7069_b1 , \7069_b0 , \7070_b1 , \7070_b0 , \7071_b1 , \7071_b0 , 
		\7072_b1 , \7072_b0 , \7073_b1 , \7073_b0 , \7074_b1 , \7074_b0 , \7075_b1 , \7075_b0 , \7076_b1 , \7076_b0 , 
		\7077_b1 , \7077_b0 , \7078_b1 , \7078_b0 , \7079_b1 , \7079_b0 , \7080_b1 , \7080_b0 , \7081_b1 , \7081_b0 , 
		\7082_b1 , \7082_b0 , \7083_b1 , \7083_b0 , \7084_b1 , \7084_b0 , \7085_b1 , \7085_b0 , \7086_b1 , \7086_b0 , 
		\7087_b1 , \7087_b0 , \7088_b1 , \7088_b0 , \7089_b1 , \7089_b0 , \7090_b1 , \7090_b0 , \7091_b1 , \7091_b0 , 
		\7092_b1 , \7092_b0 , \7093_b1 , \7093_b0 , \7094_b1 , \7094_b0 , \7095_b1 , \7095_b0 , \7096_b1 , \7096_b0 , 
		\7097_b1 , \7097_b0 , \7098_b1 , \7098_b0 , \7099_b1 , \7099_b0 , \7100_b1 , \7100_b0 , \7101_b1 , \7101_b0 , 
		\7102_b1 , \7102_b0 , \7103_b1 , \7103_b0 , \7104_b1 , \7104_b0 , \7105_b1 , \7105_b0 , \7106_b1 , \7106_b0 , 
		\7107_b1 , \7107_b0 , \7108_b1 , \7108_b0 , \7109_b1 , \7109_b0 , \7110_b1 , \7110_b0 , \7111_b1 , \7111_b0 , 
		\7112_b1 , \7112_b0 , \7113_b1 , \7113_b0 , \7114_b1 , \7114_b0 , \7115_b1 , \7115_b0 , \7116_b1 , \7116_b0 , 
		\7117_b1 , \7117_b0 , \7118_b1 , \7118_b0 , \7119_b1 , \7119_b0 , \7120_b1 , \7120_b0 , \7121_b1 , \7121_b0 , 
		\7122_b1 , \7122_b0 , \7123_b1 , \7123_b0 , \7124_b1 , \7124_b0 , \7125_b1 , \7125_b0 , \7126_b1 , \7126_b0 , 
		\7127_b1 , \7127_b0 , \7128_b1 , \7128_b0 , \7129_b1 , \7129_b0 , \7130_b1 , \7130_b0 , \7131_b1 , \7131_b0 , 
		\7132_b1 , \7132_b0 , \7133_b1 , \7133_b0 , \7134_b1 , \7134_b0 , \7135_b1 , \7135_b0 , \7136_b1 , \7136_b0 , 
		\7137_b1 , \7137_b0 , \7138_b1 , \7138_b0 , \7139_b1 , \7139_b0 , \7140_b1 , \7140_b0 , \7141_b1 , \7141_b0 , 
		\7142_b1 , \7142_b0 , \7143_b1 , \7143_b0 , \7144_b1 , \7144_b0 , \7145_b1 , \7145_b0 , \7146_b1 , \7146_b0 , 
		\7147_b1 , \7147_b0 , \7148_b1 , \7148_b0 , \7149_b1 , \7149_b0 , \7150_b1 , \7150_b0 , \7151_b1 , \7151_b0 , 
		\7152_b1 , \7152_b0 , \7153_b1 , \7153_b0 , \7154_b1 , \7154_b0 , \7155_b1 , \7155_b0 , \7156_b1 , \7156_b0 , 
		\7157_b1 , \7157_b0 , \7158_b1 , \7158_b0 , \7159_b1 , \7159_b0 , \7160_b1 , \7160_b0 , \7161_b1 , \7161_b0 , 
		\7162_b1 , \7162_b0 , \7163_b1 , \7163_b0 , \7164_b1 , \7164_b0 , \7165_b1 , \7165_b0 , \7166_b1 , \7166_b0 , 
		\7167_b1 , \7167_b0 , \7168_b1 , \7168_b0 , \7169_b1 , \7169_b0 , \7170_b1 , \7170_b0 , \7171_b1 , \7171_b0 , 
		\7172_b1 , \7172_b0 , \7173_b1 , \7173_b0 , \7174_b1 , \7174_b0 , \7175_b1 , \7175_b0 , \7176_b1 , \7176_b0 , 
		\7177_b1 , \7177_b0 , \7178_b1 , \7178_b0 , \7179_b1 , \7179_b0 , \7180_b1 , \7180_b0 , \7181_b1 , \7181_b0 , 
		\7182_b1 , \7182_b0 , \7183_b1 , \7183_b0 , \7184_b1 , \7184_b0 , \7185_b1 , \7185_b0 , \7186_b1 , \7186_b0 , 
		\7187_b1 , \7187_b0 , \7188_b1 , \7188_b0 , \7189_b1 , \7189_b0 , \7190_b1 , \7190_b0 , \7191_b1 , \7191_b0 , 
		\7192_b1 , \7192_b0 , \7193_b1 , \7193_b0 , \7194_b1 , \7194_b0 , \7195_b1 , \7195_b0 , \7196_b1 , \7196_b0 , 
		\7197_b1 , \7197_b0 , \7198_b1 , \7198_b0 , \7199_b1 , \7199_b0 , \7200_b1 , \7200_b0 , \7201_b1 , \7201_b0 , 
		\7202_b1 , \7202_b0 , \7203_b1 , \7203_b0 , \7204_b1 , \7204_b0 , \7205_b1 , \7205_b0 , \7206_b1 , \7206_b0 , 
		\7207_b1 , \7207_b0 , \7208_b1 , \7208_b0 , \7209_b1 , \7209_b0 , \7210_b1 , \7210_b0 , \7211_b1 , \7211_b0 , 
		\7212_b1 , \7212_b0 , \7213_b1 , \7213_b0 , \7214_b1 , \7214_b0 , \7215_b1 , \7215_b0 , \7216_b1 , \7216_b0 , 
		w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , w_6 , w_7 , w_8 , w_9 , 
		w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , w_16 , w_17 , w_18 , w_19 , 
		w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , w_26 , w_27 , w_28 , w_29 , 
		w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , w_36 , w_37 , w_38 , w_39 , 
		w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , w_46 , w_47 , w_48 , w_49 , 
		w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , w_56 , w_57 , w_58 , w_59 , 
		w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , w_66 , w_67 , w_68 , w_69 , 
		w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , w_76 , w_77 , w_78 , w_79 , 
		w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , w_86 , w_87 , w_88 , w_89 , 
		w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , w_96 , w_97 , w_98 , w_99 , 
		w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , w_106 , w_107 , w_108 , w_109 , 
		w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , w_116 , w_117 , w_118 , w_119 , 
		w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , w_126 , w_127 , w_128 , w_129 , 
		w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , w_136 , w_137 , w_138 , w_139 , 
		w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , w_146 , w_147 , w_148 , w_149 , 
		w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , w_156 , w_157 , w_158 , w_159 , 
		w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , w_166 , w_167 , w_168 , w_169 , 
		w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , w_176 , w_177 , w_178 , w_179 , 
		w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , w_186 , w_187 , w_188 , w_189 , 
		w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , w_196 , w_197 , w_198 , w_199 , 
		w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , w_206 , w_207 , w_208 , w_209 , 
		w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , w_216 , w_217 , w_218 , w_219 , 
		w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , w_226 , w_227 , w_228 , w_229 , 
		w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , w_236 , w_237 , w_238 , w_239 , 
		w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , w_246 , w_247 , w_248 , w_249 , 
		w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , w_256 , w_257 , w_258 , w_259 , 
		w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , w_266 , w_267 , w_268 , w_269 , 
		w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , w_276 , w_277 , w_278 , w_279 , 
		w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , w_286 , w_287 , w_288 , w_289 , 
		w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , w_296 , w_297 , w_298 , w_299 , 
		w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , w_306 , w_307 , w_308 , w_309 , 
		w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , w_316 , w_317 , w_318 , w_319 , 
		w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , w_326 , w_327 , w_328 , w_329 , 
		w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , w_336 , w_337 , w_338 , w_339 , 
		w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , w_346 , w_347 , w_348 , w_349 , 
		w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , w_356 , w_357 , w_358 , w_359 , 
		w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , w_366 , w_367 , w_368 , w_369 , 
		w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , w_376 , w_377 , w_378 , w_379 , 
		w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , w_386 , w_387 , w_388 , w_389 , 
		w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , w_396 , w_397 , w_398 , w_399 , 
		w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , w_406 , w_407 , w_408 , w_409 , 
		w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , w_416 , w_417 , w_418 , w_419 , 
		w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , w_426 , w_427 , w_428 , w_429 , 
		w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , w_436 , w_437 , w_438 , w_439 , 
		w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , w_446 , w_447 , w_448 , w_449 , 
		w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , w_456 , w_457 , w_458 , w_459 , 
		w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , w_466 , w_467 , w_468 , w_469 , 
		w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , w_476 , w_477 , w_478 , w_479 , 
		w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , w_486 , w_487 , w_488 , w_489 , 
		w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , w_496 , w_497 , w_498 , w_499 , 
		w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , w_506 , w_507 , w_508 , w_509 , 
		w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , w_516 , w_517 , w_518 , w_519 , 
		w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , w_526 , w_527 , w_528 , w_529 , 
		w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , w_536 , w_537 , w_538 , w_539 , 
		w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , w_546 , w_547 , w_548 , w_549 , 
		w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , w_556 , w_557 , w_558 , w_559 , 
		w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , w_566 , w_567 , w_568 , w_569 , 
		w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , w_576 , w_577 , w_578 , w_579 , 
		w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , w_586 , w_587 , w_588 , w_589 , 
		w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , w_596 , w_597 , w_598 , w_599 , 
		w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , w_606 , w_607 , w_608 , w_609 , 
		w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , w_616 , w_617 , w_618 , w_619 , 
		w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , w_626 , w_627 , w_628 , w_629 , 
		w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , w_636 , w_637 , w_638 , w_639 , 
		w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , w_646 , w_647 , w_648 , w_649 , 
		w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , w_656 , w_657 , w_658 , w_659 , 
		w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , w_666 , w_667 , w_668 , w_669 , 
		w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , w_676 , w_677 , w_678 , w_679 , 
		w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , w_686 , w_687 , w_688 , w_689 , 
		w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , w_696 , w_697 , w_698 , w_699 , 
		w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , w_706 , w_707 , w_708 , w_709 , 
		w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , w_716 , w_717 , w_718 , w_719 , 
		w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , w_726 , w_727 , w_728 , w_729 , 
		w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , w_736 , w_737 , w_738 , w_739 , 
		w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , w_746 , w_747 , w_748 , w_749 , 
		w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , w_756 , w_757 , w_758 , w_759 , 
		w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , w_766 , w_767 , w_768 , w_769 , 
		w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , w_776 , w_777 , w_778 , w_779 , 
		w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , w_786 , w_787 , w_788 , w_789 , 
		w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , w_796 , w_797 , w_798 , w_799 , 
		w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , w_806 , w_807 , w_808 , w_809 , 
		w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , w_816 , w_817 , w_818 , w_819 , 
		w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , w_826 , w_827 , w_828 , w_829 , 
		w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , w_836 , w_837 , w_838 , w_839 , 
		w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , w_846 , w_847 , w_848 , w_849 , 
		w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , w_856 , w_857 , w_858 , w_859 , 
		w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , w_866 , w_867 , w_868 , w_869 , 
		w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , w_876 , w_877 , w_878 , w_879 , 
		w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , w_886 , w_887 , w_888 , w_889 , 
		w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , w_896 , w_897 , w_898 , w_899 , 
		w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , w_906 , w_907 , w_908 , w_909 , 
		w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , w_916 , w_917 , w_918 , w_919 , 
		w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , w_926 , w_927 , w_928 , w_929 , 
		w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , w_936 , w_937 , w_938 , w_939 , 
		w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , w_946 , w_947 , w_948 , w_949 , 
		w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , w_956 , w_957 , w_958 , w_959 , 
		w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , w_966 , w_967 , w_968 , w_969 , 
		w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , w_976 , w_977 , w_978 , w_979 , 
		w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , w_986 , w_987 , w_988 , w_989 , 
		w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , w_996 , w_997 , w_998 , w_999 , 
		w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , w_1006 , w_1007 , w_1008 , w_1009 , 
		w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , w_1016 , w_1017 , w_1018 , w_1019 , 
		w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , w_1026 , w_1027 , w_1028 , w_1029 , 
		w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , w_1036 , w_1037 , w_1038 , w_1039 , 
		w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , w_1046 , w_1047 , w_1048 , w_1049 , 
		w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , w_1056 , w_1057 , w_1058 , w_1059 , 
		w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , w_1066 , w_1067 , w_1068 , w_1069 , 
		w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , w_1076 , w_1077 , w_1078 , w_1079 , 
		w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , w_1086 , w_1087 , w_1088 , w_1089 , 
		w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , w_1096 , w_1097 , w_1098 , w_1099 , 
		w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , w_1106 , w_1107 , w_1108 , w_1109 , 
		w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , w_1116 , w_1117 , w_1118 , w_1119 , 
		w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , w_1126 , w_1127 , w_1128 , w_1129 , 
		w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , w_1136 , w_1137 , w_1138 , w_1139 , 
		w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , w_1146 , w_1147 , w_1148 , w_1149 , 
		w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , w_1156 , w_1157 , w_1158 , w_1159 , 
		w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , w_1166 , w_1167 , w_1168 , w_1169 , 
		w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , w_1176 , w_1177 , w_1178 , w_1179 , 
		w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , w_1186 , w_1187 , w_1188 , w_1189 , 
		w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , w_1196 , w_1197 , w_1198 , w_1199 , 
		w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , w_1206 , w_1207 , w_1208 , w_1209 , 
		w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , w_1216 , w_1217 , w_1218 , w_1219 , 
		w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , w_1226 , w_1227 , w_1228 , w_1229 , 
		w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , w_1236 , w_1237 , w_1238 , w_1239 , 
		w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , w_1246 , w_1247 , w_1248 , w_1249 , 
		w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , w_1256 , w_1257 , w_1258 , w_1259 , 
		w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , w_1266 , w_1267 , w_1268 , w_1269 , 
		w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , w_1276 , w_1277 , w_1278 , w_1279 , 
		w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , w_1286 , w_1287 , w_1288 , w_1289 , 
		w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , w_1296 , w_1297 , w_1298 , w_1299 , 
		w_1300 , w_1301 , w_1302 , w_1303 , w_1304 , w_1305 , w_1306 , w_1307 , w_1308 , w_1309 , 
		w_1310 , w_1311 , w_1312 , w_1313 , w_1314 , w_1315 , w_1316 , w_1317 , w_1318 , w_1319 , 
		w_1320 , w_1321 , w_1322 , w_1323 , w_1324 , w_1325 , w_1326 , w_1327 , w_1328 , w_1329 , 
		w_1330 , w_1331 , w_1332 , w_1333 , w_1334 , w_1335 , w_1336 , w_1337 , w_1338 , w_1339 , 
		w_1340 , w_1341 , w_1342 , w_1343 , w_1344 , w_1345 , w_1346 , w_1347 , w_1348 , w_1349 , 
		w_1350 , w_1351 , w_1352 , w_1353 , w_1354 , w_1355 , w_1356 , w_1357 , w_1358 , w_1359 , 
		w_1360 , w_1361 , w_1362 , w_1363 , w_1364 , w_1365 , w_1366 , w_1367 , w_1368 , w_1369 , 
		w_1370 , w_1371 , w_1372 , w_1373 , w_1374 , w_1375 , w_1376 , w_1377 , w_1378 , w_1379 , 
		w_1380 , w_1381 , w_1382 , w_1383 , w_1384 , w_1385 , w_1386 , w_1387 , w_1388 , w_1389 , 
		w_1390 , w_1391 , w_1392 , w_1393 , w_1394 , w_1395 , w_1396 , w_1397 , w_1398 , w_1399 , 
		w_1400 , w_1401 , w_1402 , w_1403 , w_1404 , w_1405 , w_1406 , w_1407 , w_1408 , w_1409 , 
		w_1410 , w_1411 , w_1412 , w_1413 , w_1414 , w_1415 , w_1416 , w_1417 , w_1418 , w_1419 , 
		w_1420 , w_1421 , w_1422 , w_1423 , w_1424 , w_1425 , w_1426 , w_1427 , w_1428 , w_1429 , 
		w_1430 , w_1431 , w_1432 , w_1433 , w_1434 , w_1435 , w_1436 , w_1437 , w_1438 , w_1439 , 
		w_1440 , w_1441 , w_1442 , w_1443 , w_1444 , w_1445 , w_1446 , w_1447 , w_1448 , w_1449 , 
		w_1450 , w_1451 , w_1452 , w_1453 , w_1454 , w_1455 , w_1456 , w_1457 , w_1458 , w_1459 , 
		w_1460 , w_1461 , w_1462 , w_1463 , w_1464 , w_1465 , w_1466 , w_1467 , w_1468 , w_1469 , 
		w_1470 , w_1471 , w_1472 , w_1473 , w_1474 , w_1475 , w_1476 , w_1477 , w_1478 , w_1479 , 
		w_1480 , w_1481 , w_1482 , w_1483 , w_1484 , w_1485 , w_1486 , w_1487 , w_1488 , w_1489 , 
		w_1490 , w_1491 , w_1492 , w_1493 , w_1494 , w_1495 , w_1496 , w_1497 , w_1498 , w_1499 , 
		w_1500 , w_1501 , w_1502 , w_1503 , w_1504 , w_1505 , w_1506 , w_1507 , w_1508 , w_1509 , 
		w_1510 , w_1511 , w_1512 , w_1513 , w_1514 , w_1515 , w_1516 , w_1517 , w_1518 , w_1519 , 
		w_1520 , w_1521 , w_1522 , w_1523 , w_1524 , w_1525 , w_1526 , w_1527 , w_1528 , w_1529 , 
		w_1530 , w_1531 , w_1532 , w_1533 , w_1534 , w_1535 , w_1536 , w_1537 , w_1538 , w_1539 , 
		w_1540 , w_1541 , w_1542 , w_1543 , w_1544 , w_1545 , w_1546 , w_1547 , w_1548 , w_1549 , 
		w_1550 , w_1551 , w_1552 , w_1553 , w_1554 , w_1555 , w_1556 , w_1557 , w_1558 , w_1559 , 
		w_1560 , w_1561 , w_1562 , w_1563 , w_1564 , w_1565 , w_1566 , w_1567 , w_1568 , w_1569 , 
		w_1570 , w_1571 , w_1572 , w_1573 , w_1574 , w_1575 , w_1576 , w_1577 , w_1578 , w_1579 , 
		w_1580 , w_1581 , w_1582 , w_1583 , w_1584 , w_1585 , w_1586 , w_1587 , w_1588 , w_1589 , 
		w_1590 , w_1591 , w_1592 , w_1593 , w_1594 , w_1595 , w_1596 , w_1597 , w_1598 , w_1599 , 
		w_1600 , w_1601 , w_1602 , w_1603 , w_1604 , w_1605 , w_1606 , w_1607 , w_1608 , w_1609 , 
		w_1610 , w_1611 , w_1612 , w_1613 , w_1614 , w_1615 , w_1616 , w_1617 , w_1618 , w_1619 , 
		w_1620 , w_1621 , w_1622 , w_1623 , w_1624 , w_1625 , w_1626 , w_1627 , w_1628 , w_1629 , 
		w_1630 , w_1631 , w_1632 , w_1633 , w_1634 , w_1635 , w_1636 , w_1637 , w_1638 , w_1639 , 
		w_1640 , w_1641 , w_1642 , w_1643 , w_1644 , w_1645 , w_1646 , w_1647 , w_1648 , w_1649 , 
		w_1650 , w_1651 , w_1652 , w_1653 , w_1654 , w_1655 , w_1656 , w_1657 , w_1658 , w_1659 , 
		w_1660 , w_1661 , w_1662 , w_1663 , w_1664 , w_1665 , w_1666 , w_1667 , w_1668 , w_1669 , 
		w_1670 , w_1671 , w_1672 , w_1673 , w_1674 , w_1675 , w_1676 , w_1677 , w_1678 , w_1679 , 
		w_1680 , w_1681 , w_1682 , w_1683 , w_1684 , w_1685 , w_1686 , w_1687 , w_1688 , w_1689 , 
		w_1690 , w_1691 , w_1692 , w_1693 , w_1694 , w_1695 , w_1696 , w_1697 , w_1698 , w_1699 , 
		w_1700 , w_1701 , w_1702 , w_1703 , w_1704 , w_1705 , w_1706 , w_1707 , w_1708 , w_1709 , 
		w_1710 , w_1711 , w_1712 , w_1713 , w_1714 , w_1715 , w_1716 , w_1717 , w_1718 , w_1719 , 
		w_1720 , w_1721 , w_1722 , w_1723 , w_1724 , w_1725 , w_1726 , w_1727 , w_1728 , w_1729 , 
		w_1730 , w_1731 , w_1732 , w_1733 , w_1734 , w_1735 , w_1736 , w_1737 , w_1738 , w_1739 , 
		w_1740 , w_1741 , w_1742 , w_1743 , w_1744 , w_1745 , w_1746 , w_1747 , w_1748 , w_1749 , 
		w_1750 , w_1751 , w_1752 , w_1753 , w_1754 , w_1755 , w_1756 , w_1757 , w_1758 , w_1759 , 
		w_1760 , w_1761 , w_1762 , w_1763 , w_1764 , w_1765 , w_1766 , w_1767 , w_1768 , w_1769 , 
		w_1770 , w_1771 , w_1772 , w_1773 , w_1774 , w_1775 , w_1776 , w_1777 , w_1778 , w_1779 , 
		w_1780 , w_1781 , w_1782 , w_1783 , w_1784 , w_1785 , w_1786 , w_1787 , w_1788 , w_1789 , 
		w_1790 , w_1791 , w_1792 , w_1793 , w_1794 , w_1795 , w_1796 , w_1797 , w_1798 , w_1799 , 
		w_1800 , w_1801 , w_1802 , w_1803 , w_1804 , w_1805 , w_1806 , w_1807 , w_1808 , w_1809 , 
		w_1810 , w_1811 , w_1812 , w_1813 , w_1814 , w_1815 , w_1816 , w_1817 , w_1818 , w_1819 , 
		w_1820 , w_1821 , w_1822 , w_1823 , w_1824 , w_1825 , w_1826 , w_1827 , w_1828 , w_1829 , 
		w_1830 , w_1831 , w_1832 , w_1833 , w_1834 , w_1835 , w_1836 , w_1837 , w_1838 , w_1839 , 
		w_1840 , w_1841 , w_1842 , w_1843 , w_1844 , w_1845 , w_1846 , w_1847 , w_1848 , w_1849 , 
		w_1850 , w_1851 , w_1852 , w_1853 , w_1854 , w_1855 , w_1856 , w_1857 , w_1858 , w_1859 , 
		w_1860 , w_1861 , w_1862 , w_1863 , w_1864 , w_1865 , w_1866 , w_1867 , w_1868 , w_1869 , 
		w_1870 , w_1871 , w_1872 , w_1873 , w_1874 , w_1875 , w_1876 , w_1877 , w_1878 , w_1879 , 
		w_1880 , w_1881 , w_1882 , w_1883 , w_1884 , w_1885 , w_1886 , w_1887 , w_1888 , w_1889 , 
		w_1890 , w_1891 , w_1892 , w_1893 , w_1894 , w_1895 , w_1896 , w_1897 , w_1898 , w_1899 , 
		w_1900 , w_1901 , w_1902 , w_1903 , w_1904 , w_1905 , w_1906 , w_1907 , w_1908 , w_1909 , 
		w_1910 , w_1911 , w_1912 , w_1913 , w_1914 , w_1915 , w_1916 , w_1917 , w_1918 , w_1919 , 
		w_1920 , w_1921 , w_1922 , w_1923 , w_1924 , w_1925 , w_1926 , w_1927 , w_1928 , w_1929 , 
		w_1930 , w_1931 , w_1932 , w_1933 , w_1934 , w_1935 , w_1936 , w_1937 , w_1938 , w_1939 , 
		w_1940 , w_1941 , w_1942 , w_1943 , w_1944 , w_1945 , w_1946 , w_1947 , w_1948 , w_1949 , 
		w_1950 , w_1951 , w_1952 , w_1953 , w_1954 , w_1955 , w_1956 , w_1957 , w_1958 , w_1959 , 
		w_1960 , w_1961 , w_1962 , w_1963 , w_1964 , w_1965 , w_1966 , w_1967 , w_1968 , w_1969 , 
		w_1970 , w_1971 , w_1972 , w_1973 , w_1974 , w_1975 , w_1976 , w_1977 , w_1978 , w_1979 , 
		w_1980 , w_1981 , w_1982 , w_1983 , w_1984 , w_1985 , w_1986 , w_1987 , w_1988 , w_1989 , 
		w_1990 , w_1991 , w_1992 , w_1993 , w_1994 , w_1995 , w_1996 , w_1997 , w_1998 , w_1999 , 
		w_2000 , w_2001 , w_2002 , w_2003 , w_2004 , w_2005 , w_2006 , w_2007 , w_2008 , w_2009 , 
		w_2010 , w_2011 , w_2012 , w_2013 , w_2014 , w_2015 , w_2016 , w_2017 , w_2018 , w_2019 , 
		w_2020 , w_2021 , w_2022 , w_2023 , w_2024 , w_2025 , w_2026 , w_2027 , w_2028 , w_2029 , 
		w_2030 , w_2031 , w_2032 , w_2033 , w_2034 , w_2035 , w_2036 , w_2037 , w_2038 , w_2039 , 
		w_2040 , w_2041 , w_2042 , w_2043 , w_2044 , w_2045 , w_2046 , w_2047 , w_2048 , w_2049 , 
		w_2050 , w_2051 , w_2052 , w_2053 , w_2054 , w_2055 , w_2056 , w_2057 , w_2058 , w_2059 , 
		w_2060 , w_2061 , w_2062 , w_2063 , w_2064 , w_2065 , w_2066 , w_2067 , w_2068 , w_2069 , 
		w_2070 , w_2071 , w_2072 , w_2073 , w_2074 , w_2075 , w_2076 , w_2077 , w_2078 , w_2079 , 
		w_2080 , w_2081 , w_2082 , w_2083 , w_2084 , w_2085 , w_2086 , w_2087 , w_2088 , w_2089 , 
		w_2090 , w_2091 , w_2092 , w_2093 , w_2094 , w_2095 , w_2096 , w_2097 , w_2098 , w_2099 , 
		w_2100 , w_2101 , w_2102 , w_2103 , w_2104 , w_2105 , w_2106 , w_2107 , w_2108 , w_2109 , 
		w_2110 , w_2111 , w_2112 , w_2113 , w_2114 , w_2115 , w_2116 , w_2117 , w_2118 , w_2119 , 
		w_2120 , w_2121 , w_2122 , w_2123 , w_2124 , w_2125 , w_2126 , w_2127 , w_2128 , w_2129 , 
		w_2130 , w_2131 , w_2132 , w_2133 , w_2134 , w_2135 , w_2136 , w_2137 , w_2138 , w_2139 , 
		w_2140 , w_2141 , w_2142 , w_2143 , w_2144 , w_2145 , w_2146 , w_2147 , w_2148 , w_2149 , 
		w_2150 , w_2151 , w_2152 , w_2153 , w_2154 , w_2155 , w_2156 , w_2157 , w_2158 , w_2159 , 
		w_2160 , w_2161 , w_2162 , w_2163 , w_2164 , w_2165 , w_2166 , w_2167 , w_2168 , w_2169 , 
		w_2170 , w_2171 , w_2172 , w_2173 , w_2174 , w_2175 , w_2176 , w_2177 , w_2178 , w_2179 , 
		w_2180 , w_2181 , w_2182 , w_2183 , w_2184 , w_2185 , w_2186 , w_2187 , w_2188 , w_2189 , 
		w_2190 , w_2191 , w_2192 , w_2193 , w_2194 , w_2195 , w_2196 , w_2197 , w_2198 , w_2199 , 
		w_2200 , w_2201 , w_2202 , w_2203 , w_2204 , w_2205 , w_2206 , w_2207 , w_2208 , w_2209 , 
		w_2210 , w_2211 , w_2212 , w_2213 , w_2214 , w_2215 , w_2216 , w_2217 , w_2218 , w_2219 , 
		w_2220 , w_2221 , w_2222 , w_2223 , w_2224 , w_2225 , w_2226 , w_2227 , w_2228 , w_2229 , 
		w_2230 , w_2231 , w_2232 , w_2233 , w_2234 , w_2235 , w_2236 , w_2237 , w_2238 , w_2239 , 
		w_2240 , w_2241 , w_2242 , w_2243 , w_2244 , w_2245 , w_2246 , w_2247 , w_2248 , w_2249 , 
		w_2250 , w_2251 , w_2252 , w_2253 , w_2254 , w_2255 , w_2256 , w_2257 , w_2258 , w_2259 , 
		w_2260 , w_2261 , w_2262 , w_2263 , w_2264 , w_2265 , w_2266 , w_2267 , w_2268 , w_2269 , 
		w_2270 , w_2271 , w_2272 , w_2273 , w_2274 , w_2275 , w_2276 , w_2277 , w_2278 , w_2279 , 
		w_2280 , w_2281 , w_2282 , w_2283 , w_2284 , w_2285 , w_2286 , w_2287 , w_2288 , w_2289 , 
		w_2290 , w_2291 , w_2292 , w_2293 , w_2294 , w_2295 , w_2296 , w_2297 , w_2298 , w_2299 , 
		w_2300 , w_2301 , w_2302 , w_2303 , w_2304 , w_2305 , w_2306 , w_2307 , w_2308 , w_2309 , 
		w_2310 , w_2311 , w_2312 , w_2313 , w_2314 , w_2315 , w_2316 , w_2317 , w_2318 , w_2319 , 
		w_2320 , w_2321 , w_2322 , w_2323 , w_2324 , w_2325 , w_2326 , w_2327 , w_2328 , w_2329 , 
		w_2330 , w_2331 , w_2332 , w_2333 , w_2334 , w_2335 , w_2336 , w_2337 , w_2338 , w_2339 , 
		w_2340 , w_2341 , w_2342 , w_2343 , w_2344 , w_2345 , w_2346 , w_2347 , w_2348 , w_2349 , 
		w_2350 , w_2351 , w_2352 , w_2353 , w_2354 , w_2355 , w_2356 , w_2357 , w_2358 , w_2359 , 
		w_2360 , w_2361 , w_2362 , w_2363 , w_2364 , w_2365 , w_2366 , w_2367 , w_2368 , w_2369 , 
		w_2370 , w_2371 , w_2372 , w_2373 , w_2374 , w_2375 , w_2376 , w_2377 , w_2378 , w_2379 , 
		w_2380 , w_2381 , w_2382 , w_2383 , w_2384 , w_2385 , w_2386 , w_2387 , w_2388 , w_2389 , 
		w_2390 , w_2391 , w_2392 , w_2393 , w_2394 , w_2395 , w_2396 , w_2397 , w_2398 , w_2399 , 
		w_2400 , w_2401 , w_2402 , w_2403 , w_2404 , w_2405 , w_2406 , w_2407 , w_2408 , w_2409 , 
		w_2410 , w_2411 , w_2412 , w_2413 , w_2414 , w_2415 , w_2416 , w_2417 , w_2418 , w_2419 , 
		w_2420 , w_2421 , w_2422 , w_2423 , w_2424 , w_2425 , w_2426 , w_2427 , w_2428 , w_2429 , 
		w_2430 , w_2431 , w_2432 , w_2433 , w_2434 , w_2435 , w_2436 , w_2437 , w_2438 , w_2439 , 
		w_2440 , w_2441 , w_2442 , w_2443 , w_2444 , w_2445 , w_2446 , w_2447 , w_2448 , w_2449 , 
		w_2450 , w_2451 , w_2452 , w_2453 , w_2454 , w_2455 , w_2456 , w_2457 , w_2458 , w_2459 , 
		w_2460 , w_2461 , w_2462 , w_2463 , w_2464 , w_2465 , w_2466 , w_2467 , w_2468 , w_2469 , 
		w_2470 , w_2471 , w_2472 , w_2473 , w_2474 , w_2475 , w_2476 , w_2477 , w_2478 , w_2479 , 
		w_2480 , w_2481 , w_2482 , w_2483 , w_2484 , w_2485 , w_2486 , w_2487 , w_2488 , w_2489 , 
		w_2490 , w_2491 , w_2492 , w_2493 , w_2494 , w_2495 , w_2496 , w_2497 , w_2498 , w_2499 , 
		w_2500 , w_2501 , w_2502 , w_2503 , w_2504 , w_2505 , w_2506 , w_2507 , w_2508 , w_2509 , 
		w_2510 , w_2511 , w_2512 , w_2513 , w_2514 , w_2515 , w_2516 , w_2517 , w_2518 , w_2519 , 
		w_2520 , w_2521 , w_2522 , w_2523 , w_2524 , w_2525 , w_2526 , w_2527 , w_2528 , w_2529 , 
		w_2530 , w_2531 , w_2532 , w_2533 , w_2534 , w_2535 , w_2536 , w_2537 , w_2538 , w_2539 , 
		w_2540 , w_2541 , w_2542 , w_2543 , w_2544 , w_2545 , w_2546 , w_2547 , w_2548 , w_2549 , 
		w_2550 , w_2551 , w_2552 , w_2553 , w_2554 , w_2555 , w_2556 , w_2557 , w_2558 , w_2559 , 
		w_2560 , w_2561 , w_2562 , w_2563 , w_2564 , w_2565 , w_2566 , w_2567 , w_2568 , w_2569 , 
		w_2570 , w_2571 , w_2572 , w_2573 , w_2574 , w_2575 , w_2576 , w_2577 , w_2578 , w_2579 , 
		w_2580 , w_2581 , w_2582 , w_2583 , w_2584 , w_2585 , w_2586 , w_2587 , w_2588 , w_2589 , 
		w_2590 , w_2591 , w_2592 , w_2593 , w_2594 , w_2595 , w_2596 , w_2597 , w_2598 , w_2599 , 
		w_2600 , w_2601 , w_2602 , w_2603 , w_2604 , w_2605 , w_2606 , w_2607 , w_2608 , w_2609 , 
		w_2610 , w_2611 , w_2612 , w_2613 , w_2614 , w_2615 , w_2616 , w_2617 , w_2618 , w_2619 , 
		w_2620 , w_2621 , w_2622 , w_2623 , w_2624 , w_2625 , w_2626 , w_2627 , w_2628 , w_2629 , 
		w_2630 , w_2631 , w_2632 , w_2633 , w_2634 , w_2635 , w_2636 , w_2637 , w_2638 , w_2639 , 
		w_2640 , w_2641 , w_2642 , w_2643 , w_2644 , w_2645 , w_2646 , w_2647 , w_2648 , w_2649 , 
		w_2650 , w_2651 , w_2652 , w_2653 , w_2654 , w_2655 , w_2656 , w_2657 , w_2658 , w_2659 , 
		w_2660 , w_2661 , w_2662 , w_2663 , w_2664 , w_2665 , w_2666 , w_2667 , w_2668 , w_2669 , 
		w_2670 , w_2671 , w_2672 , w_2673 , w_2674 , w_2675 , w_2676 , w_2677 , w_2678 , w_2679 , 
		w_2680 , w_2681 , w_2682 , w_2683 , w_2684 , w_2685 , w_2686 , w_2687 , w_2688 , w_2689 , 
		w_2690 , w_2691 , w_2692 , w_2693 , w_2694 , w_2695 , w_2696 , w_2697 , w_2698 , w_2699 , 
		w_2700 , w_2701 , w_2702 , w_2703 , w_2704 , w_2705 , w_2706 , w_2707 , w_2708 , w_2709 , 
		w_2710 , w_2711 , w_2712 , w_2713 , w_2714 , w_2715 , w_2716 , w_2717 , w_2718 , w_2719 , 
		w_2720 , w_2721 , w_2722 , w_2723 , w_2724 , w_2725 , w_2726 , w_2727 , w_2728 , w_2729 , 
		w_2730 , w_2731 , w_2732 , w_2733 , w_2734 , w_2735 , w_2736 , w_2737 , w_2738 , w_2739 , 
		w_2740 , w_2741 , w_2742 , w_2743 , w_2744 , w_2745 , w_2746 , w_2747 , w_2748 , w_2749 , 
		w_2750 , w_2751 , w_2752 , w_2753 , w_2754 , w_2755 , w_2756 , w_2757 , w_2758 , w_2759 , 
		w_2760 , w_2761 , w_2762 , w_2763 , w_2764 , w_2765 , w_2766 , w_2767 , w_2768 , w_2769 , 
		w_2770 , w_2771 , w_2772 , w_2773 , w_2774 , w_2775 , w_2776 , w_2777 , w_2778 , w_2779 , 
		w_2780 , w_2781 , w_2782 , w_2783 , w_2784 , w_2785 , w_2786 , w_2787 , w_2788 , w_2789 , 
		w_2790 , w_2791 , w_2792 , w_2793 , w_2794 , w_2795 , w_2796 , w_2797 , w_2798 , w_2799 , 
		w_2800 , w_2801 , w_2802 , w_2803 , w_2804 , w_2805 , w_2806 , w_2807 , w_2808 , w_2809 , 
		w_2810 , w_2811 , w_2812 , w_2813 , w_2814 , w_2815 , w_2816 , w_2817 , w_2818 , w_2819 , 
		w_2820 , w_2821 , w_2822 , w_2823 , w_2824 , w_2825 , w_2826 , w_2827 , w_2828 , w_2829 , 
		w_2830 , w_2831 , w_2832 , w_2833 , w_2834 , w_2835 , w_2836 , w_2837 , w_2838 , w_2839 , 
		w_2840 , w_2841 , w_2842 , w_2843 , w_2844 , w_2845 , w_2846 , w_2847 , w_2848 , w_2849 , 
		w_2850 , w_2851 , w_2852 , w_2853 , w_2854 , w_2855 , w_2856 , w_2857 , w_2858 , w_2859 , 
		w_2860 , w_2861 , w_2862 , w_2863 , w_2864 , w_2865 , w_2866 , w_2867 , w_2868 , w_2869 , 
		w_2870 , w_2871 , w_2872 , w_2873 , w_2874 , w_2875 , w_2876 , w_2877 , w_2878 , w_2879 , 
		w_2880 , w_2881 , w_2882 , w_2883 , w_2884 , w_2885 , w_2886 , w_2887 , w_2888 , w_2889 , 
		w_2890 , w_2891 , w_2892 , w_2893 , w_2894 , w_2895 , w_2896 , w_2897 , w_2898 , w_2899 , 
		w_2900 , w_2901 , w_2902 , w_2903 , w_2904 , w_2905 , w_2906 , w_2907 , w_2908 , w_2909 , 
		w_2910 , w_2911 , w_2912 , w_2913 , w_2914 , w_2915 , w_2916 , w_2917 , w_2918 , w_2919 , 
		w_2920 , w_2921 , w_2922 , w_2923 , w_2924 , w_2925 , w_2926 , w_2927 , w_2928 , w_2929 , 
		w_2930 , w_2931 , w_2932 , w_2933 , w_2934 , w_2935 , w_2936 , w_2937 , w_2938 , w_2939 , 
		w_2940 , w_2941 , w_2942 , w_2943 , w_2944 , w_2945 , w_2946 , w_2947 , w_2948 , w_2949 , 
		w_2950 , w_2951 , w_2952 , w_2953 , w_2954 , w_2955 , w_2956 , w_2957 , w_2958 , w_2959 , 
		w_2960 , w_2961 , w_2962 , w_2963 , w_2964 , w_2965 , w_2966 , w_2967 , w_2968 , w_2969 , 
		w_2970 , w_2971 , w_2972 , w_2973 , w_2974 , w_2975 , w_2976 , w_2977 , w_2978 , w_2979 , 
		w_2980 , w_2981 , w_2982 , w_2983 , w_2984 , w_2985 , w_2986 , w_2987 , w_2988 , w_2989 , 
		w_2990 , w_2991 , w_2992 , w_2993 , w_2994 , w_2995 , w_2996 , w_2997 , w_2998 , w_2999 , 
		w_3000 , w_3001 , w_3002 , w_3003 , w_3004 , w_3005 , w_3006 , w_3007 , w_3008 , w_3009 , 
		w_3010 , w_3011 , w_3012 , w_3013 , w_3014 , w_3015 , w_3016 , w_3017 , w_3018 , w_3019 , 
		w_3020 , w_3021 , w_3022 , w_3023 , w_3024 , w_3025 , w_3026 , w_3027 , w_3028 , w_3029 , 
		w_3030 , w_3031 , w_3032 , w_3033 , w_3034 , w_3035 , w_3036 , w_3037 , w_3038 , w_3039 , 
		w_3040 , w_3041 , w_3042 , w_3043 , w_3044 , w_3045 , w_3046 , w_3047 , w_3048 , w_3049 , 
		w_3050 , w_3051 , w_3052 , w_3053 , w_3054 , w_3055 , w_3056 , w_3057 , w_3058 , w_3059 , 
		w_3060 , w_3061 , w_3062 , w_3063 , w_3064 , w_3065 , w_3066 , w_3067 , w_3068 , w_3069 , 
		w_3070 , w_3071 , w_3072 , w_3073 , w_3074 , w_3075 , w_3076 , w_3077 , w_3078 , w_3079 , 
		w_3080 , w_3081 , w_3082 , w_3083 , w_3084 , w_3085 , w_3086 , w_3087 , w_3088 , w_3089 , 
		w_3090 , w_3091 , w_3092 , w_3093 , w_3094 , w_3095 , w_3096 , w_3097 , w_3098 , w_3099 , 
		w_3100 , w_3101 , w_3102 , w_3103 , w_3104 , w_3105 , w_3106 , w_3107 , w_3108 , w_3109 , 
		w_3110 , w_3111 , w_3112 , w_3113 , w_3114 , w_3115 , w_3116 , w_3117 , w_3118 , w_3119 , 
		w_3120 , w_3121 , w_3122 , w_3123 , w_3124 , w_3125 , w_3126 , w_3127 , w_3128 , w_3129 , 
		w_3130 , w_3131 , w_3132 , w_3133 , w_3134 , w_3135 , w_3136 , w_3137 , w_3138 , w_3139 , 
		w_3140 , w_3141 , w_3142 , w_3143 , w_3144 , w_3145 , w_3146 , w_3147 , w_3148 , w_3149 , 
		w_3150 , w_3151 , w_3152 , w_3153 , w_3154 , w_3155 , w_3156 , w_3157 , w_3158 , w_3159 , 
		w_3160 , w_3161 , w_3162 , w_3163 , w_3164 , w_3165 , w_3166 , w_3167 , w_3168 , w_3169 , 
		w_3170 , w_3171 , w_3172 , w_3173 , w_3174 , w_3175 , w_3176 , w_3177 , w_3178 , w_3179 , 
		w_3180 , w_3181 , w_3182 , w_3183 , w_3184 , w_3185 , w_3186 , w_3187 , w_3188 , w_3189 , 
		w_3190 , w_3191 , w_3192 , w_3193 , w_3194 , w_3195 , w_3196 , w_3197 , w_3198 , w_3199 , 
		w_3200 , w_3201 , w_3202 , w_3203 , w_3204 , w_3205 , w_3206 , w_3207 , w_3208 , w_3209 , 
		w_3210 , w_3211 , w_3212 , w_3213 , w_3214 , w_3215 , w_3216 , w_3217 , w_3218 , w_3219 , 
		w_3220 , w_3221 , w_3222 , w_3223 , w_3224 , w_3225 , w_3226 , w_3227 , w_3228 , w_3229 , 
		w_3230 , w_3231 , w_3232 , w_3233 , w_3234 , w_3235 , w_3236 , w_3237 , w_3238 , w_3239 , 
		w_3240 , w_3241 , w_3242 , w_3243 , w_3244 , w_3245 , w_3246 , w_3247 , w_3248 , w_3249 , 
		w_3250 , w_3251 , w_3252 , w_3253 , w_3254 , w_3255 , w_3256 , w_3257 , w_3258 , w_3259 , 
		w_3260 , w_3261 , w_3262 , w_3263 , w_3264 , w_3265 , w_3266 , w_3267 , w_3268 , w_3269 , 
		w_3270 , w_3271 , w_3272 , w_3273 , w_3274 , w_3275 , w_3276 , w_3277 , w_3278 , w_3279 , 
		w_3280 , w_3281 , w_3282 , w_3283 , w_3284 , w_3285 , w_3286 , w_3287 , w_3288 , w_3289 , 
		w_3290 , w_3291 , w_3292 , w_3293 , w_3294 , w_3295 , w_3296 , w_3297 , w_3298 , w_3299 , 
		w_3300 , w_3301 , w_3302 , w_3303 , w_3304 , w_3305 , w_3306 , w_3307 , w_3308 , w_3309 , 
		w_3310 , w_3311 , w_3312 , w_3313 , w_3314 , w_3315 , w_3316 , w_3317 , w_3318 , w_3319 , 
		w_3320 , w_3321 , w_3322 , w_3323 , w_3324 , w_3325 , w_3326 , w_3327 , w_3328 , w_3329 , 
		w_3330 , w_3331 , w_3332 , w_3333 , w_3334 , w_3335 , w_3336 , w_3337 , w_3338 , w_3339 , 
		w_3340 , w_3341 , w_3342 , w_3343 , w_3344 , w_3345 , w_3346 , w_3347 , w_3348 , w_3349 , 
		w_3350 , w_3351 , w_3352 , w_3353 , w_3354 , w_3355 , w_3356 , w_3357 , w_3358 , w_3359 , 
		w_3360 , w_3361 , w_3362 , w_3363 , w_3364 , w_3365 , w_3366 , w_3367 , w_3368 , w_3369 , 
		w_3370 , w_3371 , w_3372 , w_3373 , w_3374 , w_3375 , w_3376 , w_3377 , w_3378 , w_3379 , 
		w_3380 , w_3381 , w_3382 , w_3383 , w_3384 , w_3385 , w_3386 , w_3387 , w_3388 , w_3389 , 
		w_3390 , w_3391 , w_3392 , w_3393 , w_3394 , w_3395 , w_3396 , w_3397 , w_3398 , w_3399 , 
		w_3400 , w_3401 , w_3402 , w_3403 , w_3404 , w_3405 , w_3406 , w_3407 , w_3408 , w_3409 , 
		w_3410 , w_3411 , w_3412 , w_3413 , w_3414 , w_3415 , w_3416 , w_3417 , w_3418 , w_3419 , 
		w_3420 , w_3421 , w_3422 , w_3423 , w_3424 , w_3425 , w_3426 , w_3427 , w_3428 , w_3429 , 
		w_3430 , w_3431 , w_3432 , w_3433 , w_3434 , w_3435 , w_3436 , w_3437 , w_3438 , w_3439 , 
		w_3440 , w_3441 , w_3442 , w_3443 , w_3444 , w_3445 , w_3446 , w_3447 , w_3448 , w_3449 , 
		w_3450 , w_3451 , w_3452 , w_3453 , w_3454 , w_3455 , w_3456 , w_3457 , w_3458 , w_3459 , 
		w_3460 , w_3461 , w_3462 , w_3463 , w_3464 , w_3465 , w_3466 , w_3467 , w_3468 , w_3469 , 
		w_3470 , w_3471 , w_3472 , w_3473 , w_3474 , w_3475 , w_3476 , w_3477 , w_3478 , w_3479 , 
		w_3480 , w_3481 , w_3482 , w_3483 , w_3484 , w_3485 , w_3486 , w_3487 , w_3488 , w_3489 , 
		w_3490 , w_3491 , w_3492 , w_3493 , w_3494 , w_3495 , w_3496 , w_3497 , w_3498 , w_3499 , 
		w_3500 , w_3501 , w_3502 , w_3503 , w_3504 , w_3505 , w_3506 , w_3507 , w_3508 , w_3509 , 
		w_3510 , w_3511 , w_3512 , w_3513 , w_3514 , w_3515 , w_3516 , w_3517 , w_3518 , w_3519 , 
		w_3520 , w_3521 , w_3522 , w_3523 , w_3524 , w_3525 , w_3526 , w_3527 , w_3528 , w_3529 , 
		w_3530 , w_3531 , w_3532 , w_3533 , w_3534 , w_3535 , w_3536 , w_3537 , w_3538 , w_3539 , 
		w_3540 , w_3541 , w_3542 , w_3543 , w_3544 , w_3545 , w_3546 , w_3547 , w_3548 , w_3549 , 
		w_3550 , w_3551 , w_3552 , w_3553 , w_3554 , w_3555 , w_3556 , w_3557 , w_3558 , w_3559 , 
		w_3560 , w_3561 , w_3562 , w_3563 , w_3564 , w_3565 , w_3566 , w_3567 , w_3568 , w_3569 , 
		w_3570 , w_3571 , w_3572 , w_3573 , w_3574 , w_3575 , w_3576 , w_3577 , w_3578 , w_3579 , 
		w_3580 , w_3581 , w_3582 , w_3583 , w_3584 , w_3585 , w_3586 , w_3587 , w_3588 , w_3589 , 
		w_3590 , w_3591 , w_3592 , w_3593 , w_3594 , w_3595 , w_3596 , w_3597 , w_3598 , w_3599 , 
		w_3600 , w_3601 , w_3602 , w_3603 , w_3604 , w_3605 , w_3606 , w_3607 , w_3608 , w_3609 , 
		w_3610 , w_3611 , w_3612 , w_3613 , w_3614 , w_3615 , w_3616 , w_3617 , w_3618 , w_3619 , 
		w_3620 , w_3621 , w_3622 , w_3623 , w_3624 , w_3625 , w_3626 , w_3627 , w_3628 , w_3629 , 
		w_3630 , w_3631 , w_3632 , w_3633 , w_3634 , w_3635 , w_3636 , w_3637 , w_3638 , w_3639 , 
		w_3640 , w_3641 , w_3642 , w_3643 , w_3644 , w_3645 , w_3646 , w_3647 , w_3648 , w_3649 , 
		w_3650 , w_3651 , w_3652 , w_3653 , w_3654 , w_3655 , w_3656 , w_3657 , w_3658 , w_3659 , 
		w_3660 , w_3661 , w_3662 , w_3663 , w_3664 , w_3665 , w_3666 , w_3667 , w_3668 , w_3669 , 
		w_3670 , w_3671 , w_3672 , w_3673 , w_3674 , w_3675 , w_3676 , w_3677 , w_3678 , w_3679 , 
		w_3680 , w_3681 , w_3682 , w_3683 , w_3684 , w_3685 , w_3686 , w_3687 , w_3688 , w_3689 , 
		w_3690 , w_3691 , w_3692 , w_3693 , w_3694 , w_3695 , w_3696 , w_3697 , w_3698 , w_3699 , 
		w_3700 , w_3701 , w_3702 , w_3703 , w_3704 , w_3705 , w_3706 , w_3707 , w_3708 , w_3709 , 
		w_3710 , w_3711 , w_3712 , w_3713 , w_3714 , w_3715 , w_3716 , w_3717 , w_3718 , w_3719 , 
		w_3720 , w_3721 , w_3722 , w_3723 , w_3724 , w_3725 , w_3726 , w_3727 , w_3728 , w_3729 , 
		w_3730 , w_3731 , w_3732 , w_3733 , w_3734 , w_3735 , w_3736 , w_3737 , w_3738 , w_3739 , 
		w_3740 , w_3741 , w_3742 , w_3743 , w_3744 , w_3745 , w_3746 , w_3747 , w_3748 , w_3749 , 
		w_3750 , w_3751 , w_3752 , w_3753 , w_3754 , w_3755 , w_3756 , w_3757 , w_3758 , w_3759 , 
		w_3760 , w_3761 , w_3762 , w_3763 , w_3764 , w_3765 , w_3766 , w_3767 , w_3768 , w_3769 , 
		w_3770 , w_3771 , w_3772 , w_3773 , w_3774 , w_3775 , w_3776 , w_3777 , w_3778 , w_3779 , 
		w_3780 , w_3781 , w_3782 , w_3783 , w_3784 , w_3785 , w_3786 , w_3787 , w_3788 , w_3789 , 
		w_3790 , w_3791 , w_3792 , w_3793 , w_3794 , w_3795 , w_3796 , w_3797 , w_3798 , w_3799 , 
		w_3800 , w_3801 , w_3802 , w_3803 , w_3804 , w_3805 , w_3806 , w_3807 , w_3808 , w_3809 , 
		w_3810 , w_3811 , w_3812 , w_3813 , w_3814 , w_3815 , w_3816 , w_3817 , w_3818 , w_3819 , 
		w_3820 , w_3821 , w_3822 , w_3823 , w_3824 , w_3825 , w_3826 , w_3827 , w_3828 , w_3829 , 
		w_3830 , w_3831 , w_3832 , w_3833 , w_3834 , w_3835 , w_3836 , w_3837 , w_3838 , w_3839 , 
		w_3840 , w_3841 , w_3842 , w_3843 , w_3844 , w_3845 , w_3846 , w_3847 , w_3848 , w_3849 , 
		w_3850 , w_3851 , w_3852 , w_3853 , w_3854 , w_3855 , w_3856 , w_3857 , w_3858 , w_3859 , 
		w_3860 , w_3861 , w_3862 , w_3863 , w_3864 , w_3865 , w_3866 , w_3867 , w_3868 , w_3869 , 
		w_3870 , w_3871 , w_3872 , w_3873 , w_3874 , w_3875 , w_3876 , w_3877 , w_3878 , w_3879 , 
		w_3880 , w_3881 , w_3882 , w_3883 , w_3884 , w_3885 , w_3886 , w_3887 , w_3888 , w_3889 , 
		w_3890 , w_3891 , w_3892 , w_3893 , w_3894 , w_3895 , w_3896 , w_3897 , w_3898 , w_3899 , 
		w_3900 , w_3901 , w_3902 , w_3903 , w_3904 , w_3905 , w_3906 , w_3907 , w_3908 , w_3909 , 
		w_3910 , w_3911 , w_3912 , w_3913 , w_3914 , w_3915 , w_3916 , w_3917 , w_3918 , w_3919 , 
		w_3920 , w_3921 , w_3922 , w_3923 , w_3924 , w_3925 , w_3926 , w_3927 , w_3928 , w_3929 , 
		w_3930 , w_3931 , w_3932 , w_3933 , w_3934 , w_3935 , w_3936 , w_3937 , w_3938 , w_3939 , 
		w_3940 , w_3941 , w_3942 , w_3943 , w_3944 , w_3945 , w_3946 , w_3947 , w_3948 , w_3949 , 
		w_3950 , w_3951 , w_3952 , w_3953 , w_3954 , w_3955 , w_3956 , w_3957 , w_3958 , w_3959 , 
		w_3960 , w_3961 , w_3962 , w_3963 , w_3964 , w_3965 , w_3966 , w_3967 , w_3968 , w_3969 , 
		w_3970 , w_3971 , w_3972 , w_3973 , w_3974 , w_3975 , w_3976 , w_3977 , w_3978 , w_3979 , 
		w_3980 , w_3981 , w_3982 , w_3983 , w_3984 , w_3985 , w_3986 , w_3987 , w_3988 , w_3989 , 
		w_3990 , w_3991 , w_3992 , w_3993 , w_3994 , w_3995 , w_3996 , w_3997 , w_3998 , w_3999 , 
		w_4000 , w_4001 , w_4002 , w_4003 , w_4004 , w_4005 , w_4006 , w_4007 , w_4008 , w_4009 , 
		w_4010 , w_4011 , w_4012 , w_4013 , w_4014 , w_4015 , w_4016 , w_4017 , w_4018 , w_4019 , 
		w_4020 , w_4021 , w_4022 , w_4023 , w_4024 , w_4025 , w_4026 , w_4027 , w_4028 , w_4029 , 
		w_4030 , w_4031 , w_4032 , w_4033 , w_4034 , w_4035 , w_4036 , w_4037 , w_4038 , w_4039 , 
		w_4040 , w_4041 , w_4042 , w_4043 , w_4044 , w_4045 , w_4046 , w_4047 , w_4048 , w_4049 , 
		w_4050 , w_4051 , w_4052 , w_4053 , w_4054 , w_4055 , w_4056 , w_4057 , w_4058 , w_4059 , 
		w_4060 , w_4061 , w_4062 , w_4063 , w_4064 , w_4065 , w_4066 , w_4067 , w_4068 , w_4069 , 
		w_4070 , w_4071 , w_4072 , w_4073 , w_4074 , w_4075 , w_4076 , w_4077 , w_4078 , w_4079 , 
		w_4080 , w_4081 , w_4082 , w_4083 , w_4084 , w_4085 , w_4086 , w_4087 , w_4088 , w_4089 , 
		w_4090 , w_4091 , w_4092 , w_4093 , w_4094 , w_4095 , w_4096 , w_4097 , w_4098 , w_4099 , 
		w_4100 , w_4101 , w_4102 , w_4103 , w_4104 , w_4105 , w_4106 , w_4107 , w_4108 , w_4109 , 
		w_4110 , w_4111 , w_4112 , w_4113 , w_4114 , w_4115 , w_4116 , w_4117 , w_4118 , w_4119 , 
		w_4120 , w_4121 , w_4122 , w_4123 , w_4124 , w_4125 , w_4126 , w_4127 , w_4128 , w_4129 , 
		w_4130 , w_4131 , w_4132 , w_4133 , w_4134 , w_4135 , w_4136 , w_4137 , w_4138 , w_4139 , 
		w_4140 , w_4141 , w_4142 , w_4143 , w_4144 , w_4145 , w_4146 , w_4147 , w_4148 , w_4149 , 
		w_4150 , w_4151 , w_4152 , w_4153 , w_4154 , w_4155 , w_4156 , w_4157 , w_4158 , w_4159 , 
		w_4160 , w_4161 , w_4162 , w_4163 , w_4164 , w_4165 , w_4166 , w_4167 , w_4168 , w_4169 , 
		w_4170 , w_4171 , w_4172 , w_4173 , w_4174 , w_4175 , w_4176 , w_4177 , w_4178 , w_4179 , 
		w_4180 , w_4181 , w_4182 , w_4183 , w_4184 , w_4185 , w_4186 , w_4187 , w_4188 , w_4189 , 
		w_4190 , w_4191 , w_4192 , w_4193 , w_4194 , w_4195 , w_4196 , w_4197 , w_4198 , w_4199 , 
		w_4200 , w_4201 , w_4202 , w_4203 , w_4204 , w_4205 , w_4206 , w_4207 , w_4208 , w_4209 , 
		w_4210 , w_4211 , w_4212 , w_4213 , w_4214 , w_4215 , w_4216 , w_4217 , w_4218 , w_4219 , 
		w_4220 , w_4221 , w_4222 , w_4223 , w_4224 , w_4225 , w_4226 , w_4227 , w_4228 , w_4229 , 
		w_4230 , w_4231 , w_4232 , w_4233 , w_4234 , w_4235 , w_4236 , w_4237 , w_4238 , w_4239 , 
		w_4240 , w_4241 , w_4242 , w_4243 , w_4244 , w_4245 , w_4246 , w_4247 , w_4248 , w_4249 , 
		w_4250 , w_4251 , w_4252 , w_4253 , w_4254 , w_4255 , w_4256 , w_4257 , w_4258 , w_4259 , 
		w_4260 , w_4261 , w_4262 , w_4263 , w_4264 , w_4265 , w_4266 , w_4267 , w_4268 , w_4269 , 
		w_4270 , w_4271 , w_4272 , w_4273 , w_4274 , w_4275 , w_4276 , w_4277 , w_4278 , w_4279 , 
		w_4280 , w_4281 , w_4282 , w_4283 , w_4284 , w_4285 , w_4286 , w_4287 , w_4288 , w_4289 , 
		w_4290 , w_4291 , w_4292 , w_4293 , w_4294 , w_4295 , w_4296 , w_4297 , w_4298 , w_4299 , 
		w_4300 , w_4301 , w_4302 , w_4303 , w_4304 , w_4305 , w_4306 , w_4307 , w_4308 , w_4309 , 
		w_4310 , w_4311 , w_4312 , w_4313 , w_4314 , w_4315 , w_4316 , w_4317 , w_4318 , w_4319 , 
		w_4320 , w_4321 , w_4322 , w_4323 , w_4324 , w_4325 , w_4326 , w_4327 , w_4328 , w_4329 , 
		w_4330 , w_4331 , w_4332 , w_4333 , w_4334 , w_4335 , w_4336 , w_4337 , w_4338 , w_4339 , 
		w_4340 , w_4341 , w_4342 , w_4343 , w_4344 , w_4345 , w_4346 , w_4347 , w_4348 , w_4349 , 
		w_4350 , w_4351 , w_4352 , w_4353 , w_4354 , w_4355 , w_4356 , w_4357 , w_4358 , w_4359 , 
		w_4360 , w_4361 , w_4362 , w_4363 , w_4364 , w_4365 , w_4366 , w_4367 , w_4368 , w_4369 , 
		w_4370 , w_4371 , w_4372 , w_4373 , w_4374 , w_4375 , w_4376 , w_4377 , w_4378 , w_4379 , 
		w_4380 , w_4381 , w_4382 , w_4383 , w_4384 , w_4385 , w_4386 , w_4387 , w_4388 , w_4389 , 
		w_4390 , w_4391 , w_4392 , w_4393 , w_4394 , w_4395 , w_4396 , w_4397 , w_4398 , w_4399 , 
		w_4400 , w_4401 , w_4402 , w_4403 , w_4404 , w_4405 , w_4406 , w_4407 , w_4408 , w_4409 , 
		w_4410 , w_4411 , w_4412 , w_4413 , w_4414 , w_4415 , w_4416 , w_4417 , w_4418 , w_4419 , 
		w_4420 , w_4421 , w_4422 , w_4423 , w_4424 , w_4425 , w_4426 , w_4427 , w_4428 , w_4429 , 
		w_4430 , w_4431 , w_4432 , w_4433 , w_4434 , w_4435 , w_4436 , w_4437 , w_4438 , w_4439 , 
		w_4440 , w_4441 , w_4442 , w_4443 , w_4444 , w_4445 , w_4446 , w_4447 , w_4448 , w_4449 , 
		w_4450 , w_4451 , w_4452 , w_4453 , w_4454 , w_4455 , w_4456 , w_4457 , w_4458 , w_4459 , 
		w_4460 , w_4461 , w_4462 , w_4463 , w_4464 , w_4465 , w_4466 , w_4467 , w_4468 , w_4469 , 
		w_4470 , w_4471 , w_4472 , w_4473 , w_4474 , w_4475 , w_4476 , w_4477 , w_4478 , w_4479 , 
		w_4480 , w_4481 , w_4482 , w_4483 , w_4484 , w_4485 , w_4486 , w_4487 , w_4488 , w_4489 , 
		w_4490 , w_4491 , w_4492 , w_4493 , w_4494 , w_4495 , w_4496 , w_4497 , w_4498 , w_4499 , 
		w_4500 , w_4501 , w_4502 , w_4503 , w_4504 , w_4505 , w_4506 , w_4507 , w_4508 , w_4509 , 
		w_4510 , w_4511 , w_4512 , w_4513 , w_4514 , w_4515 , w_4516 , w_4517 , w_4518 , w_4519 , 
		w_4520 , w_4521 , w_4522 , w_4523 , w_4524 , w_4525 , w_4526 , w_4527 , w_4528 , w_4529 , 
		w_4530 , w_4531 , w_4532 , w_4533 , w_4534 , w_4535 , w_4536 , w_4537 , w_4538 , w_4539 , 
		w_4540 , w_4541 , w_4542 , w_4543 , w_4544 , w_4545 , w_4546 , w_4547 , w_4548 , w_4549 , 
		w_4550 , w_4551 , w_4552 , w_4553 , w_4554 , w_4555 , w_4556 , w_4557 , w_4558 , w_4559 , 
		w_4560 , w_4561 , w_4562 , w_4563 , w_4564 , w_4565 , w_4566 , w_4567 , w_4568 , w_4569 , 
		w_4570 , w_4571 , w_4572 , w_4573 , w_4574 , w_4575 , w_4576 , w_4577 , w_4578 , w_4579 , 
		w_4580 , w_4581 , w_4582 , w_4583 , w_4584 , w_4585 , w_4586 , w_4587 , w_4588 , w_4589 , 
		w_4590 , w_4591 , w_4592 , w_4593 , w_4594 , w_4595 , w_4596 , w_4597 , w_4598 , w_4599 , 
		w_4600 , w_4601 , w_4602 , w_4603 , w_4604 , w_4605 , w_4606 , w_4607 , w_4608 , w_4609 , 
		w_4610 , w_4611 , w_4612 , w_4613 , w_4614 , w_4615 , w_4616 , w_4617 , w_4618 , w_4619 , 
		w_4620 , w_4621 , w_4622 , w_4623 , w_4624 , w_4625 , w_4626 , w_4627 , w_4628 , w_4629 , 
		w_4630 , w_4631 , w_4632 , w_4633 , w_4634 , w_4635 , w_4636 , w_4637 , w_4638 , w_4639 , 
		w_4640 , w_4641 , w_4642 , w_4643 , w_4644 , w_4645 , w_4646 , w_4647 , w_4648 , w_4649 , 
		w_4650 , w_4651 , w_4652 , w_4653 , w_4654 , w_4655 , w_4656 , w_4657 , w_4658 , w_4659 , 
		w_4660 , w_4661 , w_4662 , w_4663 , w_4664 , w_4665 , w_4666 , w_4667 , w_4668 , w_4669 , 
		w_4670 , w_4671 , w_4672 , w_4673 , w_4674 , w_4675 , w_4676 , w_4677 , w_4678 , w_4679 , 
		w_4680 , w_4681 , w_4682 , w_4683 , w_4684 , w_4685 , w_4686 , w_4687 , w_4688 , w_4689 , 
		w_4690 , w_4691 , w_4692 , w_4693 , w_4694 , w_4695 , w_4696 , w_4697 , w_4698 , w_4699 , 
		w_4700 , w_4701 , w_4702 , w_4703 , w_4704 , w_4705 , w_4706 , w_4707 , w_4708 , w_4709 , 
		w_4710 , w_4711 , w_4712 , w_4713 , w_4714 , w_4715 , w_4716 , w_4717 , w_4718 , w_4719 , 
		w_4720 , w_4721 , w_4722 , w_4723 , w_4724 , w_4725 , w_4726 , w_4727 , w_4728 , w_4729 , 
		w_4730 , w_4731 , w_4732 , w_4733 , w_4734 , w_4735 , w_4736 , w_4737 , w_4738 , w_4739 , 
		w_4740 , w_4741 , w_4742 , w_4743 , w_4744 , w_4745 , w_4746 , w_4747 , w_4748 , w_4749 , 
		w_4750 , w_4751 , w_4752 , w_4753 , w_4754 , w_4755 , w_4756 , w_4757 , w_4758 , w_4759 , 
		w_4760 , w_4761 , w_4762 , w_4763 , w_4764 , w_4765 , w_4766 , w_4767 , w_4768 , w_4769 , 
		w_4770 , w_4771 , w_4772 , w_4773 , w_4774 , w_4775 , w_4776 , w_4777 , w_4778 , w_4779 , 
		w_4780 , w_4781 , w_4782 , w_4783 , w_4784 , w_4785 , w_4786 , w_4787 , w_4788 , w_4789 , 
		w_4790 , w_4791 , w_4792 , w_4793 , w_4794 , w_4795 , w_4796 , w_4797 , w_4798 , w_4799 , 
		w_4800 , w_4801 , w_4802 , w_4803 , w_4804 , w_4805 , w_4806 , w_4807 , w_4808 , w_4809 , 
		w_4810 , w_4811 , w_4812 , w_4813 , w_4814 , w_4815 , w_4816 , w_4817 , w_4818 , w_4819 , 
		w_4820 , w_4821 , w_4822 , w_4823 , w_4824 , w_4825 , w_4826 , w_4827 , w_4828 , w_4829 , 
		w_4830 , w_4831 , w_4832 , w_4833 , w_4834 , w_4835 , w_4836 , w_4837 , w_4838 , w_4839 , 
		w_4840 , w_4841 , w_4842 , w_4843 , w_4844 , w_4845 , w_4846 , w_4847 , w_4848 , w_4849 , 
		w_4850 , w_4851 , w_4852 , w_4853 , w_4854 , w_4855 , w_4856 , w_4857 , w_4858 , w_4859 , 
		w_4860 , w_4861 , w_4862 , w_4863 , w_4864 , w_4865 , w_4866 , w_4867 , w_4868 , w_4869 , 
		w_4870 , w_4871 , w_4872 , w_4873 , w_4874 , w_4875 , w_4876 , w_4877 , w_4878 , w_4879 , 
		w_4880 , w_4881 , w_4882 , w_4883 , w_4884 , w_4885 , w_4886 , w_4887 , w_4888 , w_4889 , 
		w_4890 , w_4891 , w_4892 , w_4893 , w_4894 , w_4895 , w_4896 , w_4897 , w_4898 , w_4899 , 
		w_4900 , w_4901 , w_4902 , w_4903 , w_4904 , w_4905 , w_4906 , w_4907 , w_4908 , w_4909 , 
		w_4910 , w_4911 , w_4912 , w_4913 , w_4914 , w_4915 , w_4916 , w_4917 , w_4918 , w_4919 , 
		w_4920 , w_4921 , w_4922 , w_4923 , w_4924 , w_4925 , w_4926 , w_4927 , w_4928 , w_4929 , 
		w_4930 , w_4931 , w_4932 , w_4933 , w_4934 , w_4935 , w_4936 , w_4937 , w_4938 , w_4939 , 
		w_4940 , w_4941 , w_4942 , w_4943 , w_4944 , w_4945 , w_4946 , w_4947 , w_4948 , w_4949 , 
		w_4950 , w_4951 , w_4952 , w_4953 , w_4954 , w_4955 , w_4956 , w_4957 , w_4958 , w_4959 , 
		w_4960 , w_4961 , w_4962 , w_4963 , w_4964 , w_4965 , w_4966 , w_4967 , w_4968 , w_4969 , 
		w_4970 , w_4971 , w_4972 , w_4973 , w_4974 , w_4975 , w_4976 , w_4977 , w_4978 , w_4979 , 
		w_4980 , w_4981 , w_4982 , w_4983 , w_4984 , w_4985 , w_4986 , w_4987 , w_4988 , w_4989 , 
		w_4990 , w_4991 , w_4992 , w_4993 , w_4994 , w_4995 , w_4996 , w_4997 , w_4998 , w_4999 , 
		w_5000 , w_5001 , w_5002 , w_5003 , w_5004 , w_5005 , w_5006 , w_5007 , w_5008 , w_5009 , 
		w_5010 , w_5011 , w_5012 , w_5013 , w_5014 , w_5015 , w_5016 , w_5017 , w_5018 , w_5019 , 
		w_5020 , w_5021 , w_5022 , w_5023 , w_5024 , w_5025 , w_5026 , w_5027 , w_5028 , w_5029 , 
		w_5030 , w_5031 , w_5032 , w_5033 , w_5034 , w_5035 , w_5036 , w_5037 , w_5038 , w_5039 , 
		w_5040 , w_5041 , w_5042 , w_5043 , w_5044 , w_5045 , w_5046 , w_5047 , w_5048 , w_5049 , 
		w_5050 , w_5051 , w_5052 , w_5053 , w_5054 , w_5055 , w_5056 , w_5057 , w_5058 , w_5059 , 
		w_5060 , w_5061 , w_5062 , w_5063 , w_5064 , w_5065 , w_5066 , w_5067 , w_5068 , w_5069 , 
		w_5070 , w_5071 , w_5072 , w_5073 , w_5074 , w_5075 , w_5076 , w_5077 , w_5078 , w_5079 , 
		w_5080 , w_5081 , w_5082 , w_5083 , w_5084 , w_5085 , w_5086 , w_5087 , w_5088 , w_5089 , 
		w_5090 , w_5091 , w_5092 , w_5093 , w_5094 , w_5095 , w_5096 , w_5097 , w_5098 , w_5099 , 
		w_5100 , w_5101 , w_5102 , w_5103 , w_5104 , w_5105 , w_5106 , w_5107 , w_5108 , w_5109 , 
		w_5110 , w_5111 , w_5112 , w_5113 , w_5114 , w_5115 , w_5116 , w_5117 , w_5118 , w_5119 , 
		w_5120 , w_5121 , w_5122 , w_5123 , w_5124 , w_5125 , w_5126 , w_5127 , w_5128 , w_5129 , 
		w_5130 , w_5131 , w_5132 , w_5133 , w_5134 , w_5135 , w_5136 , w_5137 , w_5138 , w_5139 , 
		w_5140 , w_5141 , w_5142 , w_5143 , w_5144 , w_5145 , w_5146 , w_5147 , w_5148 , w_5149 , 
		w_5150 , w_5151 , w_5152 , w_5153 , w_5154 , w_5155 , w_5156 , w_5157 , w_5158 , w_5159 , 
		w_5160 , w_5161 , w_5162 , w_5163 , w_5164 , w_5165 , w_5166 , w_5167 , w_5168 , w_5169 , 
		w_5170 , w_5171 , w_5172 , w_5173 , w_5174 , w_5175 , w_5176 , w_5177 , w_5178 , w_5179 , 
		w_5180 , w_5181 , w_5182 , w_5183 , w_5184 , w_5185 , w_5186 , w_5187 , w_5188 , w_5189 , 
		w_5190 , w_5191 , w_5192 , w_5193 , w_5194 , w_5195 , w_5196 , w_5197 , w_5198 , w_5199 , 
		w_5200 , w_5201 , w_5202 , w_5203 , w_5204 , w_5205 , w_5206 , w_5207 , w_5208 , w_5209 , 
		w_5210 , w_5211 , w_5212 , w_5213 , w_5214 , w_5215 , w_5216 , w_5217 , w_5218 , w_5219 , 
		w_5220 , w_5221 , w_5222 , w_5223 , w_5224 , w_5225 , w_5226 , w_5227 , w_5228 , w_5229 , 
		w_5230 , w_5231 , w_5232 , w_5233 , w_5234 , w_5235 , w_5236 , w_5237 , w_5238 , w_5239 , 
		w_5240 , w_5241 , w_5242 , w_5243 , w_5244 , w_5245 , w_5246 , w_5247 , w_5248 , w_5249 , 
		w_5250 , w_5251 , w_5252 , w_5253 , w_5254 , w_5255 , w_5256 , w_5257 , w_5258 , w_5259 , 
		w_5260 , w_5261 , w_5262 , w_5263 , w_5264 , w_5265 , w_5266 , w_5267 , w_5268 , w_5269 , 
		w_5270 , w_5271 , w_5272 , w_5273 , w_5274 , w_5275 , w_5276 , w_5277 , w_5278 , w_5279 , 
		w_5280 , w_5281 , w_5282 , w_5283 , w_5284 , w_5285 , w_5286 , w_5287 , w_5288 , w_5289 , 
		w_5290 , w_5291 , w_5292 , w_5293 , w_5294 , w_5295 , w_5296 , w_5297 , w_5298 , w_5299 , 
		w_5300 , w_5301 , w_5302 , w_5303 , w_5304 , w_5305 , w_5306 , w_5307 , w_5308 , w_5309 , 
		w_5310 , w_5311 , w_5312 , w_5313 , w_5314 , w_5315 , w_5316 , w_5317 , w_5318 , w_5319 , 
		w_5320 , w_5321 , w_5322 , w_5323 , w_5324 , w_5325 , w_5326 , w_5327 , w_5328 , w_5329 , 
		w_5330 , w_5331 , w_5332 , w_5333 , w_5334 , w_5335 , w_5336 , w_5337 , w_5338 , w_5339 , 
		w_5340 , w_5341 , w_5342 , w_5343 , w_5344 , w_5345 , w_5346 , w_5347 , w_5348 , w_5349 , 
		w_5350 , w_5351 , w_5352 , w_5353 , w_5354 , w_5355 , w_5356 , w_5357 , w_5358 , w_5359 , 
		w_5360 , w_5361 , w_5362 , w_5363 , w_5364 , w_5365 , w_5366 , w_5367 , w_5368 , w_5369 , 
		w_5370 , w_5371 , w_5372 , w_5373 , w_5374 , w_5375 , w_5376 , w_5377 , w_5378 , w_5379 , 
		w_5380 , w_5381 , w_5382 , w_5383 , w_5384 , w_5385 , w_5386 , w_5387 , w_5388 , w_5389 , 
		w_5390 , w_5391 , w_5392 , w_5393 , w_5394 , w_5395 , w_5396 , w_5397 , w_5398 , w_5399 , 
		w_5400 , w_5401 , w_5402 , w_5403 , w_5404 , w_5405 , w_5406 , w_5407 , w_5408 , w_5409 , 
		w_5410 , w_5411 , w_5412 , w_5413 , w_5414 , w_5415 , w_5416 , w_5417 , w_5418 , w_5419 , 
		w_5420 , w_5421 , w_5422 , w_5423 , w_5424 , w_5425 , w_5426 , w_5427 , w_5428 , w_5429 , 
		w_5430 , w_5431 , w_5432 , w_5433 , w_5434 , w_5435 , w_5436 , w_5437 , w_5438 , w_5439 , 
		w_5440 , w_5441 , w_5442 , w_5443 , w_5444 , w_5445 , w_5446 , w_5447 , w_5448 , w_5449 , 
		w_5450 , w_5451 , w_5452 , w_5453 , w_5454 , w_5455 , w_5456 , w_5457 , w_5458 , w_5459 , 
		w_5460 , w_5461 , w_5462 , w_5463 , w_5464 , w_5465 , w_5466 , w_5467 , w_5468 , w_5469 , 
		w_5470 , w_5471 , w_5472 , w_5473 , w_5474 , w_5475 , w_5476 , w_5477 , w_5478 , w_5479 , 
		w_5480 , w_5481 , w_5482 , w_5483 , w_5484 , w_5485 , w_5486 , w_5487 , w_5488 , w_5489 , 
		w_5490 , w_5491 , w_5492 , w_5493 , w_5494 , w_5495 , w_5496 , w_5497 , w_5498 , w_5499 , 
		w_5500 , w_5501 , w_5502 , w_5503 , w_5504 , w_5505 , w_5506 , w_5507 , w_5508 , w_5509 , 
		w_5510 , w_5511 , w_5512 , w_5513 , w_5514 , w_5515 , w_5516 , w_5517 , w_5518 , w_5519 , 
		w_5520 , w_5521 , w_5522 , w_5523 , w_5524 , w_5525 , w_5526 , w_5527 , w_5528 , w_5529 , 
		w_5530 , w_5531 , w_5532 , w_5533 , w_5534 , w_5535 , w_5536 , w_5537 , w_5538 , w_5539 , 
		w_5540 , w_5541 , w_5542 , w_5543 , w_5544 , w_5545 , w_5546 , w_5547 , w_5548 , w_5549 , 
		w_5550 , w_5551 , w_5552 , w_5553 , w_5554 , w_5555 , w_5556 , w_5557 , w_5558 , w_5559 , 
		w_5560 , w_5561 , w_5562 , w_5563 , w_5564 , w_5565 , w_5566 , w_5567 , w_5568 , w_5569 , 
		w_5570 , w_5571 , w_5572 , w_5573 , w_5574 , w_5575 , w_5576 , w_5577 , w_5578 , w_5579 , 
		w_5580 , w_5581 , w_5582 , w_5583 , w_5584 , w_5585 , w_5586 , w_5587 , w_5588 , w_5589 , 
		w_5590 , w_5591 , w_5592 , w_5593 , w_5594 , w_5595 , w_5596 , w_5597 , w_5598 , w_5599 , 
		w_5600 , w_5601 , w_5602 , w_5603 , w_5604 , w_5605 , w_5606 , w_5607 , w_5608 , w_5609 , 
		w_5610 , w_5611 , w_5612 , w_5613 , w_5614 , w_5615 , w_5616 , w_5617 , w_5618 , w_5619 , 
		w_5620 , w_5621 , w_5622 , w_5623 , w_5624 , w_5625 , w_5626 , w_5627 , w_5628 , w_5629 , 
		w_5630 , w_5631 , w_5632 , w_5633 , w_5634 , w_5635 , w_5636 , w_5637 , w_5638 , w_5639 , 
		w_5640 , w_5641 , w_5642 , w_5643 , w_5644 , w_5645 , w_5646 , w_5647 , w_5648 , w_5649 , 
		w_5650 , w_5651 , w_5652 , w_5653 , w_5654 , w_5655 , w_5656 , w_5657 , w_5658 , w_5659 , 
		w_5660 , w_5661 , w_5662 , w_5663 , w_5664 , w_5665 , w_5666 , w_5667 , w_5668 , w_5669 , 
		w_5670 , w_5671 , w_5672 , w_5673 , w_5674 , w_5675 , w_5676 , w_5677 , w_5678 , w_5679 , 
		w_5680 , w_5681 , w_5682 , w_5683 , w_5684 , w_5685 , w_5686 , w_5687 , w_5688 , w_5689 , 
		w_5690 , w_5691 , w_5692 , w_5693 , w_5694 , w_5695 , w_5696 , w_5697 , w_5698 , w_5699 , 
		w_5700 , w_5701 , w_5702 , w_5703 , w_5704 , w_5705 , w_5706 , w_5707 , w_5708 , w_5709 , 
		w_5710 , w_5711 , w_5712 , w_5713 , w_5714 , w_5715 , w_5716 , w_5717 , w_5718 , w_5719 , 
		w_5720 , w_5721 , w_5722 , w_5723 , w_5724 , w_5725 , w_5726 , w_5727 , w_5728 , w_5729 , 
		w_5730 , w_5731 , w_5732 , w_5733 , w_5734 , w_5735 , w_5736 , w_5737 , w_5738 , w_5739 , 
		w_5740 , w_5741 , w_5742 , w_5743 , w_5744 , w_5745 , w_5746 , w_5747 , w_5748 , w_5749 , 
		w_5750 , w_5751 , w_5752 , w_5753 , w_5754 , w_5755 , w_5756 , w_5757 , w_5758 , w_5759 , 
		w_5760 , w_5761 , w_5762 , w_5763 , w_5764 , w_5765 , w_5766 , w_5767 , w_5768 , w_5769 , 
		w_5770 , w_5771 , w_5772 , w_5773 , w_5774 , w_5775 , w_5776 , w_5777 , w_5778 , w_5779 , 
		w_5780 , w_5781 , w_5782 , w_5783 , w_5784 , w_5785 , w_5786 , w_5787 , w_5788 , w_5789 , 
		w_5790 , w_5791 , w_5792 , w_5793 , w_5794 , w_5795 , w_5796 , w_5797 , w_5798 , w_5799 , 
		w_5800 , w_5801 , w_5802 , w_5803 , w_5804 , w_5805 , w_5806 , w_5807 , w_5808 , w_5809 , 
		w_5810 , w_5811 , w_5812 , w_5813 , w_5814 , w_5815 , w_5816 , w_5817 , w_5818 , w_5819 , 
		w_5820 , w_5821 , w_5822 , w_5823 , w_5824 , w_5825 , w_5826 , w_5827 , w_5828 , w_5829 , 
		w_5830 , w_5831 , w_5832 , w_5833 , w_5834 , w_5835 , w_5836 , w_5837 , w_5838 , w_5839 , 
		w_5840 , w_5841 , w_5842 , w_5843 , w_5844 , w_5845 , w_5846 , w_5847 , w_5848 , w_5849 , 
		w_5850 , w_5851 , w_5852 , w_5853 , w_5854 , w_5855 , w_5856 , w_5857 , w_5858 , w_5859 , 
		w_5860 , w_5861 , w_5862 , w_5863 , w_5864 , w_5865 , w_5866 , w_5867 , w_5868 , w_5869 , 
		w_5870 , w_5871 , w_5872 , w_5873 , w_5874 , w_5875 , w_5876 , w_5877 , w_5878 , w_5879 , 
		w_5880 , w_5881 , w_5882 , w_5883 , w_5884 , w_5885 , w_5886 , w_5887 , w_5888 , w_5889 , 
		w_5890 , w_5891 , w_5892 , w_5893 , w_5894 , w_5895 , w_5896 , w_5897 , w_5898 , w_5899 , 
		w_5900 , w_5901 , w_5902 , w_5903 , w_5904 , w_5905 , w_5906 , w_5907 , w_5908 , w_5909 , 
		w_5910 , w_5911 , w_5912 , w_5913 , w_5914 , w_5915 , w_5916 , w_5917 , w_5918 , w_5919 , 
		w_5920 , w_5921 , w_5922 , w_5923 , w_5924 , w_5925 , w_5926 , w_5927 , w_5928 , w_5929 , 
		w_5930 , w_5931 , w_5932 , w_5933 , w_5934 , w_5935 , w_5936 , w_5937 , w_5938 , w_5939 , 
		w_5940 , w_5941 , w_5942 , w_5943 , w_5944 , w_5945 , w_5946 , w_5947 , w_5948 , w_5949 , 
		w_5950 , w_5951 , w_5952 , w_5953 , w_5954 , w_5955 , w_5956 , w_5957 , w_5958 , w_5959 , 
		w_5960 , w_5961 , w_5962 , w_5963 , w_5964 , w_5965 , w_5966 , w_5967 , w_5968 , w_5969 , 
		w_5970 , w_5971 , w_5972 , w_5973 , w_5974 , w_5975 , w_5976 , w_5977 , w_5978 , w_5979 , 
		w_5980 , w_5981 , w_5982 , w_5983 , w_5984 , w_5985 , w_5986 , w_5987 , w_5988 , w_5989 , 
		w_5990 , w_5991 , w_5992 , w_5993 , w_5994 , w_5995 , w_5996 , w_5997 , w_5998 , w_5999 , 
		w_6000 , w_6001 , w_6002 , w_6003 , w_6004 , w_6005 , w_6006 , w_6007 , w_6008 , w_6009 , 
		w_6010 , w_6011 , w_6012 , w_6013 , w_6014 , w_6015 , w_6016 , w_6017 , w_6018 , w_6019 , 
		w_6020 , w_6021 , w_6022 , w_6023 , w_6024 , w_6025 , w_6026 , w_6027 , w_6028 , w_6029 , 
		w_6030 , w_6031 , w_6032 , w_6033 , w_6034 , w_6035 , w_6036 , w_6037 , w_6038 , w_6039 , 
		w_6040 , w_6041 , w_6042 , w_6043 , w_6044 , w_6045 , w_6046 , w_6047 , w_6048 , w_6049 , 
		w_6050 , w_6051 , w_6052 , w_6053 , w_6054 , w_6055 , w_6056 , w_6057 , w_6058 , w_6059 , 
		w_6060 , w_6061 , w_6062 , w_6063 , w_6064 , w_6065 , w_6066 , w_6067 , w_6068 , w_6069 , 
		w_6070 , w_6071 , w_6072 , w_6073 , w_6074 , w_6075 , w_6076 , w_6077 , w_6078 , w_6079 , 
		w_6080 , w_6081 , w_6082 , w_6083 , w_6084 , w_6085 , w_6086 , w_6087 , w_6088 , w_6089 , 
		w_6090 , w_6091 , w_6092 , w_6093 , w_6094 , w_6095 , w_6096 , w_6097 , w_6098 , w_6099 , 
		w_6100 , w_6101 , w_6102 , w_6103 , w_6104 , w_6105 , w_6106 , w_6107 , w_6108 , w_6109 , 
		w_6110 , w_6111 , w_6112 , w_6113 , w_6114 , w_6115 , w_6116 , w_6117 , w_6118 , w_6119 , 
		w_6120 , w_6121 , w_6122 , w_6123 , w_6124 , w_6125 , w_6126 , w_6127 , w_6128 , w_6129 , 
		w_6130 , w_6131 , w_6132 , w_6133 , w_6134 , w_6135 , w_6136 , w_6137 , w_6138 , w_6139 , 
		w_6140 , w_6141 , w_6142 , w_6143 , w_6144 , w_6145 , w_6146 , w_6147 , w_6148 , w_6149 , 
		w_6150 , w_6151 , w_6152 , w_6153 , w_6154 , w_6155 , w_6156 , w_6157 , w_6158 , w_6159 , 
		w_6160 , w_6161 , w_6162 , w_6163 , w_6164 , w_6165 , w_6166 , w_6167 , w_6168 , w_6169 , 
		w_6170 , w_6171 , w_6172 , w_6173 , w_6174 , w_6175 , w_6176 , w_6177 , w_6178 , w_6179 , 
		w_6180 , w_6181 , w_6182 , w_6183 , w_6184 , w_6185 , w_6186 , w_6187 , w_6188 , w_6189 , 
		w_6190 , w_6191 , w_6192 , w_6193 , w_6194 , w_6195 , w_6196 , w_6197 , w_6198 , w_6199 , 
		w_6200 , w_6201 , w_6202 , w_6203 , w_6204 , w_6205 , w_6206 , w_6207 , w_6208 , w_6209 , 
		w_6210 , w_6211 , w_6212 , w_6213 , w_6214 , w_6215 , w_6216 , w_6217 , w_6218 , w_6219 , 
		w_6220 , w_6221 , w_6222 , w_6223 , w_6224 , w_6225 , w_6226 , w_6227 , w_6228 , w_6229 , 
		w_6230 , w_6231 , w_6232 , w_6233 , w_6234 , w_6235 , w_6236 , w_6237 , w_6238 , w_6239 , 
		w_6240 , w_6241 , w_6242 , w_6243 , w_6244 , w_6245 , w_6246 , w_6247 , w_6248 , w_6249 , 
		w_6250 , w_6251 , w_6252 , w_6253 , w_6254 , w_6255 , w_6256 , w_6257 , w_6258 , w_6259 , 
		w_6260 , w_6261 , w_6262 , w_6263 , w_6264 , w_6265 , w_6266 , w_6267 , w_6268 , w_6269 , 
		w_6270 , w_6271 , w_6272 , w_6273 , w_6274 , w_6275 , w_6276 , w_6277 , w_6278 , w_6279 , 
		w_6280 , w_6281 , w_6282 , w_6283 , w_6284 , w_6285 , w_6286 , w_6287 , w_6288 , w_6289 , 
		w_6290 , w_6291 , w_6292 , w_6293 , w_6294 , w_6295 , w_6296 , w_6297 , w_6298 , w_6299 , 
		w_6300 , w_6301 , w_6302 , w_6303 , w_6304 , w_6305 , w_6306 , w_6307 , w_6308 , w_6309 , 
		w_6310 , w_6311 , w_6312 , w_6313 , w_6314 , w_6315 , w_6316 , w_6317 , w_6318 , w_6319 , 
		w_6320 , w_6321 , w_6322 , w_6323 , w_6324 , w_6325 , w_6326 , w_6327 , w_6328 , w_6329 , 
		w_6330 , w_6331 , w_6332 , w_6333 , w_6334 , w_6335 , w_6336 , w_6337 , w_6338 , w_6339 , 
		w_6340 , w_6341 , w_6342 , w_6343 , w_6344 , w_6345 , w_6346 , w_6347 , w_6348 , w_6349 , 
		w_6350 , w_6351 , w_6352 , w_6353 , w_6354 , w_6355 , w_6356 , w_6357 , w_6358 , w_6359 , 
		w_6360 , w_6361 , w_6362 , w_6363 , w_6364 , w_6365 , w_6366 , w_6367 , w_6368 , w_6369 , 
		w_6370 , w_6371 , w_6372 , w_6373 , w_6374 , w_6375 , w_6376 , w_6377 , w_6378 , w_6379 , 
		w_6380 , w_6381 , w_6382 , w_6383 , w_6384 , w_6385 , w_6386 , w_6387 , w_6388 , w_6389 , 
		w_6390 , w_6391 , w_6392 , w_6393 , w_6394 , w_6395 , w_6396 , w_6397 , w_6398 , w_6399 , 
		w_6400 , w_6401 , w_6402 , w_6403 , w_6404 , w_6405 , w_6406 , w_6407 , w_6408 , w_6409 , 
		w_6410 , w_6411 , w_6412 , w_6413 , w_6414 , w_6415 , w_6416 , w_6417 , w_6418 , w_6419 , 
		w_6420 , w_6421 , w_6422 , w_6423 , w_6424 , w_6425 , w_6426 , w_6427 , w_6428 , w_6429 , 
		w_6430 , w_6431 , w_6432 , w_6433 , w_6434 , w_6435 , w_6436 , w_6437 , w_6438 , w_6439 , 
		w_6440 , w_6441 , w_6442 , w_6443 , w_6444 , w_6445 , w_6446 , w_6447 , w_6448 , w_6449 , 
		w_6450 , w_6451 , w_6452 , w_6453 , w_6454 , w_6455 , w_6456 , w_6457 , w_6458 , w_6459 , 
		w_6460 , w_6461 , w_6462 , w_6463 , w_6464 , w_6465 , w_6466 , w_6467 , w_6468 , w_6469 , 
		w_6470 , w_6471 , w_6472 , w_6473 , w_6474 , w_6475 , w_6476 , w_6477 , w_6478 , w_6479 , 
		w_6480 , w_6481 , w_6482 , w_6483 , w_6484 , w_6485 , w_6486 , w_6487 , w_6488 , w_6489 , 
		w_6490 , w_6491 , w_6492 , w_6493 , w_6494 , w_6495 , w_6496 , w_6497 , w_6498 , w_6499 , 
		w_6500 , w_6501 , w_6502 , w_6503 , w_6504 , w_6505 , w_6506 , w_6507 , w_6508 , w_6509 , 
		w_6510 , w_6511 , w_6512 , w_6513 , w_6514 , w_6515 , w_6516 , w_6517 , w_6518 , w_6519 , 
		w_6520 , w_6521 , w_6522 , w_6523 , w_6524 , w_6525 , w_6526 , w_6527 , w_6528 , w_6529 , 
		w_6530 , w_6531 , w_6532 , w_6533 , w_6534 , w_6535 , w_6536 , w_6537 , w_6538 , w_6539 , 
		w_6540 , w_6541 , w_6542 , w_6543 , w_6544 , w_6545 , w_6546 , w_6547 , w_6548 , w_6549 , 
		w_6550 , w_6551 , w_6552 , w_6553 , w_6554 , w_6555 , w_6556 , w_6557 , w_6558 , w_6559 , 
		w_6560 , w_6561 , w_6562 , w_6563 , w_6564 , w_6565 , w_6566 , w_6567 , w_6568 , w_6569 , 
		w_6570 , w_6571 , w_6572 , w_6573 , w_6574 , w_6575 , w_6576 , w_6577 , w_6578 , w_6579 , 
		w_6580 , w_6581 , w_6582 , w_6583 , w_6584 , w_6585 , w_6586 , w_6587 , w_6588 , w_6589 , 
		w_6590 , w_6591 , w_6592 , w_6593 , w_6594 , w_6595 , w_6596 , w_6597 , w_6598 , w_6599 , 
		w_6600 , w_6601 , w_6602 , w_6603 , w_6604 , w_6605 , w_6606 , w_6607 , w_6608 , w_6609 , 
		w_6610 , w_6611 , w_6612 , w_6613 , w_6614 , w_6615 , w_6616 , w_6617 , w_6618 , w_6619 , 
		w_6620 , w_6621 , w_6622 , w_6623 , w_6624 , w_6625 , w_6626 , w_6627 , w_6628 , w_6629 , 
		w_6630 , w_6631 , w_6632 , w_6633 , w_6634 , w_6635 , w_6636 , w_6637 , w_6638 , w_6639 , 
		w_6640 , w_6641 , w_6642 , w_6643 , w_6644 , w_6645 , w_6646 , w_6647 , w_6648 , w_6649 , 
		w_6650 , w_6651 , w_6652 , w_6653 , w_6654 , w_6655 , w_6656 , w_6657 , w_6658 , w_6659 , 
		w_6660 , w_6661 , w_6662 , w_6663 , w_6664 , w_6665 , w_6666 , w_6667 , w_6668 , w_6669 , 
		w_6670 , w_6671 , w_6672 , w_6673 , w_6674 , w_6675 , w_6676 , w_6677 , w_6678 , w_6679 , 
		w_6680 , w_6681 , w_6682 , w_6683 , w_6684 , w_6685 , w_6686 , w_6687 , w_6688 , w_6689 , 
		w_6690 , w_6691 , w_6692 , w_6693 , w_6694 , w_6695 , w_6696 , w_6697 , w_6698 , w_6699 , 
		w_6700 , w_6701 , w_6702 , w_6703 , w_6704 , w_6705 , w_6706 , w_6707 , w_6708 , w_6709 , 
		w_6710 , w_6711 , w_6712 , w_6713 , w_6714 , w_6715 , w_6716 , w_6717 , w_6718 , w_6719 , 
		w_6720 , w_6721 , w_6722 , w_6723 , w_6724 , w_6725 , w_6726 , w_6727 , w_6728 , w_6729 , 
		w_6730 , w_6731 , w_6732 , w_6733 , w_6734 , w_6735 , w_6736 , w_6737 , w_6738 , w_6739 , 
		w_6740 , w_6741 , w_6742 , w_6743 , w_6744 , w_6745 , w_6746 , w_6747 , w_6748 , w_6749 , 
		w_6750 , w_6751 , w_6752 , w_6753 , w_6754 , w_6755 , w_6756 , w_6757 , w_6758 , w_6759 , 
		w_6760 , w_6761 , w_6762 , w_6763 , w_6764 , w_6765 , w_6766 , w_6767 , w_6768 , w_6769 , 
		w_6770 , w_6771 , w_6772 , w_6773 , w_6774 , w_6775 , w_6776 , w_6777 , w_6778 , w_6779 , 
		w_6780 , w_6781 , w_6782 , w_6783 , w_6784 , w_6785 , w_6786 , w_6787 , w_6788 , w_6789 , 
		w_6790 , w_6791 , w_6792 , w_6793 , w_6794 , w_6795 , w_6796 , w_6797 , w_6798 , w_6799 , 
		w_6800 , w_6801 , w_6802 , w_6803 , w_6804 , w_6805 , w_6806 , w_6807 , w_6808 , w_6809 , 
		w_6810 , w_6811 , w_6812 , w_6813 , w_6814 , w_6815 , w_6816 , w_6817 , w_6818 , w_6819 , 
		w_6820 , w_6821 , w_6822 , w_6823 , w_6824 , w_6825 , w_6826 , w_6827 , w_6828 , w_6829 , 
		w_6830 , w_6831 , w_6832 , w_6833 , w_6834 , w_6835 , w_6836 , w_6837 , w_6838 , w_6839 , 
		w_6840 , w_6841 , w_6842 , w_6843 , w_6844 , w_6845 , w_6846 , w_6847 , w_6848 , w_6849 , 
		w_6850 , w_6851 , w_6852 , w_6853 , w_6854 , w_6855 , w_6856 , w_6857 , w_6858 , w_6859 , 
		w_6860 , w_6861 , w_6862 , w_6863 , w_6864 , w_6865 , w_6866 , w_6867 , w_6868 , w_6869 , 
		w_6870 , w_6871 , w_6872 , w_6873 , w_6874 , w_6875 , w_6876 , w_6877 , w_6878 , w_6879 , 
		w_6880 , w_6881 , w_6882 , w_6883 , w_6884 , w_6885 , w_6886 , w_6887 , w_6888 , w_6889 , 
		w_6890 , w_6891 , w_6892 , w_6893 , w_6894 , w_6895 , w_6896 , w_6897 , w_6898 , w_6899 , 
		w_6900 , w_6901 , w_6902 , w_6903 , w_6904 , w_6905 , w_6906 , w_6907 , w_6908 , w_6909 , 
		w_6910 , w_6911 , w_6912 , w_6913 , w_6914 , w_6915 , w_6916 , w_6917 , w_6918 , w_6919 , 
		w_6920 , w_6921 , w_6922 , w_6923 , w_6924 , w_6925 , w_6926 , w_6927 , w_6928 , w_6929 , 
		w_6930 , w_6931 , w_6932 , w_6933 , w_6934 , w_6935 , w_6936 , w_6937 , w_6938 , w_6939 , 
		w_6940 , w_6941 , w_6942 , w_6943 , w_6944 , w_6945 , w_6946 , w_6947 , w_6948 , w_6949 , 
		w_6950 , w_6951 , w_6952 , w_6953 , w_6954 , w_6955 , w_6956 , w_6957 , w_6958 , w_6959 , 
		w_6960 , w_6961 , w_6962 , w_6963 , w_6964 , w_6965 , w_6966 , w_6967 , w_6968 , w_6969 , 
		w_6970 , w_6971 , w_6972 , w_6973 , w_6974 , w_6975 , w_6976 , w_6977 , w_6978 , w_6979 , 
		w_6980 , w_6981 , w_6982 , w_6983 , w_6984 , w_6985 , w_6986 , w_6987 , w_6988 , w_6989 , 
		w_6990 , w_6991 , w_6992 , w_6993 , w_6994 , w_6995 , w_6996 , w_6997 , w_6998 , w_6999 , 
		w_7000 , w_7001 , w_7002 , w_7003 , w_7004 , w_7005 , w_7006 , w_7007 , w_7008 , w_7009 , 
		w_7010 , w_7011 , w_7012 , w_7013 , w_7014 , w_7015 , w_7016 , w_7017 , w_7018 , w_7019 , 
		w_7020 , w_7021 , w_7022 , w_7023 , w_7024 , w_7025 , w_7026 , w_7027 , w_7028 , w_7029 , 
		w_7030 , w_7031 , w_7032 , w_7033 , w_7034 , w_7035 , w_7036 , w_7037 , w_7038 , w_7039 , 
		w_7040 , w_7041 , w_7042 , w_7043 , w_7044 , w_7045 , w_7046 , w_7047 , w_7048 , w_7049 , 
		w_7050 , w_7051 , w_7052 , w_7053 , w_7054 , w_7055 , w_7056 , w_7057 , w_7058 , w_7059 , 
		w_7060 , w_7061 , w_7062 , w_7063 , w_7064 , w_7065 , w_7066 , w_7067 , w_7068 , w_7069 , 
		w_7070 , w_7071 , w_7072 , w_7073 , w_7074 , w_7075 , w_7076 , w_7077 , w_7078 , w_7079 , 
		w_7080 , w_7081 , w_7082 , w_7083 , w_7084 , w_7085 , w_7086 , w_7087 , w_7088 , w_7089 , 
		w_7090 , w_7091 , w_7092 , w_7093 , w_7094 , w_7095 , w_7096 , w_7097 , w_7098 , w_7099 , 
		w_7100 , w_7101 , w_7102 , w_7103 , w_7104 , w_7105 , w_7106 , w_7107 , w_7108 , w_7109 , 
		w_7110 , w_7111 , w_7112 , w_7113 , w_7114 , w_7115 , w_7116 , w_7117 , w_7118 , w_7119 , 
		w_7120 , w_7121 , w_7122 , w_7123 , w_7124 , w_7125 , w_7126 , w_7127 , w_7128 , w_7129 , 
		w_7130 , w_7131 , w_7132 , w_7133 , w_7134 , w_7135 , w_7136 , w_7137 , w_7138 , w_7139 , 
		w_7140 , w_7141 , w_7142 , w_7143 , w_7144 , w_7145 , w_7146 , w_7147 , w_7148 , w_7149 , 
		w_7150 , w_7151 , w_7152 , w_7153 , w_7154 , w_7155 , w_7156 , w_7157 , w_7158 , w_7159 , 
		w_7160 , w_7161 , w_7162 , w_7163 , w_7164 , w_7165 , w_7166 , w_7167 , w_7168 , w_7169 , 
		w_7170 , w_7171 , w_7172 , w_7173 , w_7174 , w_7175 , w_7176 , w_7177 , w_7178 , w_7179 , 
		w_7180 , w_7181 , w_7182 , w_7183 , w_7184 , w_7185 , w_7186 , w_7187 , w_7188 , w_7189 , 
		w_7190 , w_7191 , w_7192 , w_7193 , w_7194 , w_7195 , w_7196 , w_7197 , w_7198 , w_7199 , 
		w_7200 , w_7201 , w_7202 , w_7203 , w_7204 , w_7205 , w_7206 , w_7207 , w_7208 , w_7209 , 
		w_7210 , w_7211 , w_7212 , w_7213 , w_7214 , w_7215 , w_7216 , w_7217 , w_7218 , w_7219 , 
		w_7220 , w_7221 , w_7222 , w_7223 , w_7224 , w_7225 , w_7226 , w_7227 , w_7228 , w_7229 , 
		w_7230 , w_7231 , w_7232 , w_7233 , w_7234 , w_7235 , w_7236 , w_7237 , w_7238 , w_7239 , 
		w_7240 , w_7241 , w_7242 , w_7243 , w_7244 , w_7245 , w_7246 , w_7247 , w_7248 , w_7249 , 
		w_7250 , w_7251 , w_7252 , w_7253 , w_7254 , w_7255 , w_7256 , w_7257 , w_7258 , w_7259 , 
		w_7260 , w_7261 , w_7262 , w_7263 , w_7264 , w_7265 , w_7266 , w_7267 , w_7268 , w_7269 , 
		w_7270 , w_7271 , w_7272 , w_7273 , w_7274 , w_7275 , w_7276 , w_7277 , w_7278 , w_7279 , 
		w_7280 , w_7281 , w_7282 , w_7283 , w_7284 , w_7285 , w_7286 , w_7287 , w_7288 , w_7289 , 
		w_7290 , w_7291 , w_7292 , w_7293 , w_7294 , w_7295 , w_7296 , w_7297 , w_7298 , w_7299 , 
		w_7300 , w_7301 , w_7302 , w_7303 , w_7304 , w_7305 , w_7306 , w_7307 , w_7308 , w_7309 , 
		w_7310 , w_7311 , w_7312 , w_7313 , w_7314 , w_7315 , w_7316 , w_7317 , w_7318 , w_7319 , 
		w_7320 , w_7321 , w_7322 , w_7323 , w_7324 , w_7325 , w_7326 , w_7327 , w_7328 , w_7329 , 
		w_7330 , w_7331 , w_7332 , w_7333 , w_7334 , w_7335 , w_7336 , w_7337 , w_7338 , w_7339 , 
		w_7340 , w_7341 , w_7342 , w_7343 , w_7344 , w_7345 , w_7346 , w_7347 , w_7348 , w_7349 , 
		w_7350 , w_7351 , w_7352 , w_7353 , w_7354 , w_7355 , w_7356 , w_7357 , w_7358 , w_7359 , 
		w_7360 , w_7361 , w_7362 , w_7363 , w_7364 , w_7365 , w_7366 , w_7367 , w_7368 , w_7369 , 
		w_7370 , w_7371 , w_7372 , w_7373 , w_7374 , w_7375 , w_7376 , w_7377 , w_7378 , w_7379 , 
		w_7380 , w_7381 , w_7382 , w_7383 , w_7384 , w_7385 , w_7386 , w_7387 , w_7388 , w_7389 , 
		w_7390 , w_7391 , w_7392 , w_7393 , w_7394 , w_7395 , w_7396 , w_7397 , w_7398 , w_7399 , 
		w_7400 , w_7401 , w_7402 , w_7403 , w_7404 , w_7405 , w_7406 , w_7407 , w_7408 , w_7409 , 
		w_7410 , w_7411 , w_7412 , w_7413 , w_7414 , w_7415 , w_7416 , w_7417 , w_7418 , w_7419 , 
		w_7420 , w_7421 , w_7422 , w_7423 , w_7424 , w_7425 , w_7426 , w_7427 , w_7428 , w_7429 , 
		w_7430 , w_7431 , w_7432 , w_7433 , w_7434 , w_7435 , w_7436 , w_7437 , w_7438 , w_7439 , 
		w_7440 , w_7441 , w_7442 , w_7443 , w_7444 , w_7445 , w_7446 , w_7447 , w_7448 , w_7449 , 
		w_7450 , w_7451 , w_7452 , w_7453 , w_7454 , w_7455 , w_7456 , w_7457 , w_7458 , w_7459 , 
		w_7460 , w_7461 , w_7462 , w_7463 , w_7464 , w_7465 , w_7466 , w_7467 , w_7468 , w_7469 , 
		w_7470 , w_7471 , w_7472 , w_7473 , w_7474 , w_7475 , w_7476 , w_7477 , w_7478 , w_7479 , 
		w_7480 , w_7481 , w_7482 , w_7483 , w_7484 , w_7485 , w_7486 , w_7487 , w_7488 , w_7489 , 
		w_7490 , w_7491 , w_7492 , w_7493 , w_7494 , w_7495 , w_7496 , w_7497 , w_7498 , w_7499 , 
		w_7500 , w_7501 , w_7502 , w_7503 , w_7504 , w_7505 , w_7506 , w_7507 , w_7508 , w_7509 , 
		w_7510 , w_7511 , w_7512 , w_7513 , w_7514 , w_7515 , w_7516 , w_7517 , w_7518 , w_7519 , 
		w_7520 , w_7521 , w_7522 , w_7523 , w_7524 , w_7525 , w_7526 , w_7527 , w_7528 , w_7529 , 
		w_7530 , w_7531 , w_7532 , w_7533 , w_7534 , w_7535 , w_7536 , w_7537 , w_7538 , w_7539 , 
		w_7540 , w_7541 , w_7542 , w_7543 , w_7544 , w_7545 , w_7546 , w_7547 , w_7548 , w_7549 , 
		w_7550 , w_7551 , w_7552 , w_7553 , w_7554 , w_7555 , w_7556 , w_7557 , w_7558 , w_7559 , 
		w_7560 , w_7561 , w_7562 , w_7563 , w_7564 , w_7565 , w_7566 , w_7567 , w_7568 , w_7569 , 
		w_7570 , w_7571 , w_7572 , w_7573 , w_7574 , w_7575 , w_7576 , w_7577 , w_7578 , w_7579 , 
		w_7580 , w_7581 , w_7582 , w_7583 , w_7584 , w_7585 , w_7586 , w_7587 , w_7588 , w_7589 , 
		w_7590 , w_7591 , w_7592 , w_7593 , w_7594 , w_7595 , w_7596 , w_7597 , w_7598 , w_7599 , 
		w_7600 , w_7601 , w_7602 , w_7603 , w_7604 , w_7605 , w_7606 , w_7607 , w_7608 , w_7609 , 
		w_7610 , w_7611 , w_7612 , w_7613 , w_7614 , w_7615 , w_7616 , w_7617 , w_7618 , w_7619 , 
		w_7620 , w_7621 , w_7622 , w_7623 , w_7624 , w_7625 , w_7626 , w_7627 , w_7628 , w_7629 , 
		w_7630 , w_7631 , w_7632 , w_7633 , w_7634 , w_7635 , w_7636 , w_7637 , w_7638 , w_7639 , 
		w_7640 , w_7641 , w_7642 , w_7643 , w_7644 , w_7645 , w_7646 , w_7647 , w_7648 , w_7649 , 
		w_7650 , w_7651 , w_7652 , w_7653 , w_7654 , w_7655 , w_7656 , w_7657 , w_7658 , w_7659 , 
		w_7660 , w_7661 , w_7662 , w_7663 , w_7664 , w_7665 , w_7666 , w_7667 , w_7668 , w_7669 , 
		w_7670 , w_7671 , w_7672 , w_7673 , w_7674 , w_7675 , w_7676 , w_7677 , w_7678 , w_7679 , 
		w_7680 , w_7681 , w_7682 , w_7683 , w_7684 , w_7685 , w_7686 , w_7687 , w_7688 , w_7689 , 
		w_7690 , w_7691 , w_7692 , w_7693 , w_7694 , w_7695 , w_7696 , w_7697 , w_7698 , w_7699 , 
		w_7700 , w_7701 , w_7702 , w_7703 , w_7704 , w_7705 , w_7706 , w_7707 , w_7708 , w_7709 , 
		w_7710 , w_7711 , w_7712 , w_7713 , w_7714 , w_7715 , w_7716 , w_7717 , w_7718 , w_7719 , 
		w_7720 , w_7721 , w_7722 , w_7723 , w_7724 , w_7725 , w_7726 , w_7727 , w_7728 , w_7729 , 
		w_7730 , w_7731 , w_7732 , w_7733 , w_7734 , w_7735 , w_7736 , w_7737 , w_7738 , w_7739 , 
		w_7740 , w_7741 , w_7742 , w_7743 , w_7744 , w_7745 , w_7746 , w_7747 , w_7748 , w_7749 , 
		w_7750 , w_7751 , w_7752 , w_7753 , w_7754 , w_7755 , w_7756 , w_7757 , w_7758 , w_7759 , 
		w_7760 , w_7761 , w_7762 , w_7763 , w_7764 , w_7765 , w_7766 , w_7767 , w_7768 , w_7769 , 
		w_7770 , w_7771 , w_7772 , w_7773 , w_7774 , w_7775 , w_7776 , w_7777 , w_7778 , w_7779 , 
		w_7780 , w_7781 , w_7782 , w_7783 , w_7784 , w_7785 , w_7786 , w_7787 , w_7788 , w_7789 , 
		w_7790 , w_7791 , w_7792 , w_7793 , w_7794 , w_7795 , w_7796 , w_7797 , w_7798 , w_7799 , 
		w_7800 , w_7801 , w_7802 , w_7803 , w_7804 , w_7805 , w_7806 , w_7807 , w_7808 , w_7809 , 
		w_7810 , w_7811 , w_7812 , w_7813 , w_7814 , w_7815 , w_7816 , w_7817 , w_7818 , w_7819 , 
		w_7820 , w_7821 , w_7822 , w_7823 , w_7824 , w_7825 , w_7826 , w_7827 , w_7828 , w_7829 , 
		w_7830 , w_7831 , w_7832 , w_7833 , w_7834 , w_7835 , w_7836 , w_7837 , w_7838 , w_7839 , 
		w_7840 , w_7841 , w_7842 , w_7843 , w_7844 , w_7845 , w_7846 , w_7847 , w_7848 , w_7849 , 
		w_7850 , w_7851 , w_7852 , w_7853 , w_7854 , w_7855 , w_7856 , w_7857 , w_7858 , w_7859 , 
		w_7860 , w_7861 , w_7862 , w_7863 , w_7864 , w_7865 , w_7866 , w_7867 , w_7868 , w_7869 , 
		w_7870 , w_7871 , w_7872 , w_7873 , w_7874 , w_7875 , w_7876 , w_7877 , w_7878 , w_7879 , 
		w_7880 , w_7881 , w_7882 , w_7883 , w_7884 , w_7885 , w_7886 , w_7887 , w_7888 , w_7889 , 
		w_7890 , w_7891 , w_7892 , w_7893 , w_7894 , w_7895 , w_7896 , w_7897 , w_7898 , w_7899 , 
		w_7900 , w_7901 , w_7902 , w_7903 , w_7904 , w_7905 , w_7906 , w_7907 , w_7908 , w_7909 , 
		w_7910 , w_7911 , w_7912 , w_7913 , w_7914 , w_7915 , w_7916 , w_7917 , w_7918 , w_7919 , 
		w_7920 , w_7921 , w_7922 , w_7923 , w_7924 , w_7925 , w_7926 , w_7927 , w_7928 , w_7929 , 
		w_7930 , w_7931 , w_7932 , w_7933 , w_7934 , w_7935 , w_7936 , w_7937 , w_7938 , w_7939 , 
		w_7940 , w_7941 , w_7942 , w_7943 , w_7944 , w_7945 , w_7946 , w_7947 , w_7948 , w_7949 , 
		w_7950 , w_7951 , w_7952 , w_7953 , w_7954 , w_7955 , w_7956 , w_7957 , w_7958 , w_7959 , 
		w_7960 , w_7961 , w_7962 , w_7963 , w_7964 , w_7965 , w_7966 , w_7967 , w_7968 , w_7969 , 
		w_7970 , w_7971 , w_7972 , w_7973 , w_7974 , w_7975 , w_7976 , w_7977 , w_7978 , w_7979 , 
		w_7980 , w_7981 , w_7982 , w_7983 , w_7984 , w_7985 , w_7986 , w_7987 , w_7988 , w_7989 , 
		w_7990 , w_7991 , w_7992 , w_7993 , w_7994 , w_7995 , w_7996 , w_7997 , w_7998 , w_7999 , 
		w_8000 , w_8001 , w_8002 , w_8003 , w_8004 , w_8005 , w_8006 , w_8007 , w_8008 , w_8009 , 
		w_8010 , w_8011 , w_8012 , w_8013 , w_8014 , w_8015 , w_8016 , w_8017 , w_8018 , w_8019 , 
		w_8020 , w_8021 , w_8022 , w_8023 , w_8024 , w_8025 , w_8026 , w_8027 , w_8028 , w_8029 , 
		w_8030 , w_8031 , w_8032 , w_8033 , w_8034 , w_8035 , w_8036 , w_8037 , w_8038 , w_8039 , 
		w_8040 , w_8041 , w_8042 , w_8043 , w_8044 , w_8045 , w_8046 , w_8047 , w_8048 , w_8049 , 
		w_8050 , w_8051 , w_8052 , w_8053 , w_8054 , w_8055 , w_8056 , w_8057 , w_8058 , w_8059 , 
		w_8060 , w_8061 , w_8062 , w_8063 , w_8064 , w_8065 , w_8066 , w_8067 , w_8068 , w_8069 , 
		w_8070 , w_8071 , w_8072 , w_8073 , w_8074 , w_8075 , w_8076 , w_8077 , w_8078 , w_8079 , 
		w_8080 , w_8081 , w_8082 , w_8083 , w_8084 , w_8085 , w_8086 , w_8087 , w_8088 , w_8089 , 
		w_8090 , w_8091 , w_8092 , w_8093 , w_8094 , w_8095 , w_8096 , w_8097 , w_8098 , w_8099 , 
		w_8100 , w_8101 , w_8102 , w_8103 , w_8104 , w_8105 , w_8106 , w_8107 , w_8108 , w_8109 , 
		w_8110 , w_8111 , w_8112 , w_8113 , w_8114 , w_8115 , w_8116 , w_8117 , w_8118 , w_8119 , 
		w_8120 , w_8121 , w_8122 , w_8123 , w_8124 , w_8125 , w_8126 , w_8127 , w_8128 , w_8129 , 
		w_8130 , w_8131 , w_8132 , w_8133 , w_8134 , w_8135 , w_8136 , w_8137 , w_8138 , w_8139 , 
		w_8140 , w_8141 , w_8142 , w_8143 , w_8144 , w_8145 , w_8146 , w_8147 , w_8148 , w_8149 , 
		w_8150 , w_8151 , w_8152 , w_8153 , w_8154 , w_8155 , w_8156 , w_8157 , w_8158 , w_8159 , 
		w_8160 , w_8161 , w_8162 , w_8163 , w_8164 , w_8165 , w_8166 , w_8167 , w_8168 , w_8169 , 
		w_8170 , w_8171 , w_8172 , w_8173 , w_8174 , w_8175 , w_8176 , w_8177 , w_8178 , w_8179 , 
		w_8180 , w_8181 , w_8182 , w_8183 , w_8184 , w_8185 , w_8186 , w_8187 , w_8188 , w_8189 , 
		w_8190 , w_8191 , w_8192 , w_8193 , w_8194 , w_8195 , w_8196 , w_8197 , w_8198 , w_8199 , 
		w_8200 , w_8201 , w_8202 , w_8203 , w_8204 , w_8205 , w_8206 , w_8207 , w_8208 , w_8209 , 
		w_8210 , w_8211 , w_8212 , w_8213 , w_8214 , w_8215 , w_8216 , w_8217 , w_8218 , w_8219 , 
		w_8220 , w_8221 , w_8222 , w_8223 , w_8224 , w_8225 , w_8226 , w_8227 , w_8228 , w_8229 , 
		w_8230 , w_8231 , w_8232 , w_8233 , w_8234 , w_8235 , w_8236 , w_8237 , w_8238 , w_8239 , 
		w_8240 , w_8241 , w_8242 , w_8243 , w_8244 , w_8245 , w_8246 , w_8247 , w_8248 , w_8249 , 
		w_8250 , w_8251 , w_8252 , w_8253 , w_8254 , w_8255 , w_8256 , w_8257 , w_8258 , w_8259 , 
		w_8260 , w_8261 , w_8262 , w_8263 , w_8264 , w_8265 , w_8266 , w_8267 , w_8268 , w_8269 , 
		w_8270 , w_8271 , w_8272 , w_8273 , w_8274 , w_8275 , w_8276 , w_8277 , w_8278 , w_8279 , 
		w_8280 , w_8281 , w_8282 , w_8283 , w_8284 , w_8285 , w_8286 , w_8287 , w_8288 , w_8289 , 
		w_8290 , w_8291 , w_8292 , w_8293 , w_8294 , w_8295 , w_8296 , w_8297 , w_8298 , w_8299 , 
		w_8300 , w_8301 , w_8302 , w_8303 , w_8304 , w_8305 , w_8306 , w_8307 , w_8308 , w_8309 , 
		w_8310 , w_8311 , w_8312 , w_8313 , w_8314 , w_8315 , w_8316 , w_8317 , w_8318 , w_8319 , 
		w_8320 , w_8321 , w_8322 , w_8323 , w_8324 , w_8325 , w_8326 , w_8327 , w_8328 , w_8329 , 
		w_8330 , w_8331 , w_8332 , w_8333 , w_8334 , w_8335 , w_8336 , w_8337 , w_8338 , w_8339 , 
		w_8340 , w_8341 , w_8342 , w_8343 , w_8344 , w_8345 , w_8346 , w_8347 , w_8348 , w_8349 , 
		w_8350 , w_8351 , w_8352 , w_8353 , w_8354 , w_8355 , w_8356 , w_8357 , w_8358 , w_8359 , 
		w_8360 , w_8361 , w_8362 , w_8363 , w_8364 , w_8365 , w_8366 , w_8367 , w_8368 , w_8369 , 
		w_8370 , w_8371 , w_8372 , w_8373 , w_8374 , w_8375 , w_8376 , w_8377 , w_8378 , w_8379 , 
		w_8380 , w_8381 , w_8382 , w_8383 , w_8384 , w_8385 , w_8386 , w_8387 , w_8388 , w_8389 , 
		w_8390 , w_8391 , w_8392 , w_8393 , w_8394 , w_8395 , w_8396 , w_8397 , w_8398 , w_8399 , 
		w_8400 , w_8401 , w_8402 , w_8403 , w_8404 , w_8405 , w_8406 , w_8407 , w_8408 , w_8409 , 
		w_8410 , w_8411 , w_8412 , w_8413 , w_8414 , w_8415 , w_8416 , w_8417 , w_8418 , w_8419 , 
		w_8420 , w_8421 , w_8422 , w_8423 , w_8424 , w_8425 , w_8426 , w_8427 , w_8428 , w_8429 , 
		w_8430 , w_8431 , w_8432 , w_8433 , w_8434 , w_8435 , w_8436 , w_8437 , w_8438 , w_8439 , 
		w_8440 , w_8441 , w_8442 , w_8443 , w_8444 , w_8445 , w_8446 , w_8447 , w_8448 , w_8449 , 
		w_8450 , w_8451 , w_8452 , w_8453 , w_8454 , w_8455 , w_8456 , w_8457 , w_8458 , w_8459 , 
		w_8460 , w_8461 , w_8462 , w_8463 , w_8464 , w_8465 , w_8466 , w_8467 , w_8468 , w_8469 , 
		w_8470 , w_8471 , w_8472 , w_8473 , w_8474 , w_8475 , w_8476 , w_8477 , w_8478 , w_8479 , 
		w_8480 , w_8481 , w_8482 , w_8483 , w_8484 , w_8485 , w_8486 , w_8487 , w_8488 , w_8489 , 
		w_8490 , w_8491 , w_8492 , w_8493 , w_8494 , w_8495 , w_8496 , w_8497 , w_8498 , w_8499 , 
		w_8500 , w_8501 , w_8502 , w_8503 , w_8504 , w_8505 , w_8506 , w_8507 , w_8508 , w_8509 , 
		w_8510 , w_8511 , w_8512 , w_8513 , w_8514 , w_8515 , w_8516 , w_8517 , w_8518 , w_8519 , 
		w_8520 , w_8521 , w_8522 , w_8523 , w_8524 , w_8525 , w_8526 , w_8527 , w_8528 , w_8529 , 
		w_8530 , w_8531 , w_8532 , w_8533 , w_8534 , w_8535 , w_8536 , w_8537 , w_8538 , w_8539 , 
		w_8540 , w_8541 , w_8542 , w_8543 , w_8544 , w_8545 , w_8546 , w_8547 , w_8548 , w_8549 , 
		w_8550 , w_8551 , w_8552 , w_8553 , w_8554 , w_8555 , w_8556 , w_8557 , w_8558 , w_8559 , 
		w_8560 , w_8561 , w_8562 , w_8563 , w_8564 , w_8565 , w_8566 , w_8567 , w_8568 , w_8569 , 
		w_8570 , w_8571 , w_8572 , w_8573 , w_8574 , w_8575 , w_8576 , w_8577 , w_8578 , w_8579 , 
		w_8580 , w_8581 , w_8582 , w_8583 , w_8584 , w_8585 , w_8586 , w_8587 , w_8588 , w_8589 , 
		w_8590 , w_8591 , w_8592 , w_8593 , w_8594 , w_8595 , w_8596 , w_8597 , w_8598 , w_8599 , 
		w_8600 , w_8601 , w_8602 , w_8603 , w_8604 , w_8605 , w_8606 , w_8607 , w_8608 , w_8609 , 
		w_8610 , w_8611 , w_8612 , w_8613 , w_8614 , w_8615 , w_8616 , w_8617 , w_8618 , w_8619 , 
		w_8620 , w_8621 , w_8622 , w_8623 , w_8624 , w_8625 , w_8626 , w_8627 , w_8628 , w_8629 , 
		w_8630 , w_8631 , w_8632 , w_8633 , w_8634 , w_8635 , w_8636 , w_8637 , w_8638 , w_8639 , 
		w_8640 , w_8641 , w_8642 , w_8643 , w_8644 , w_8645 , w_8646 , w_8647 , w_8648 , w_8649 , 
		w_8650 , w_8651 , w_8652 , w_8653 , w_8654 , w_8655 , w_8656 , w_8657 , w_8658 , w_8659 , 
		w_8660 , w_8661 , w_8662 , w_8663 , w_8664 , w_8665 , w_8666 , w_8667 , w_8668 , w_8669 , 
		w_8670 , w_8671 , w_8672 , w_8673 , w_8674 , w_8675 , w_8676 , w_8677 , w_8678 , w_8679 , 
		w_8680 , w_8681 , w_8682 , w_8683 , w_8684 , w_8685 , w_8686 , w_8687 , w_8688 , w_8689 , 
		w_8690 , w_8691 , w_8692 , w_8693 , w_8694 , w_8695 , w_8696 , w_8697 , w_8698 , w_8699 , 
		w_8700 , w_8701 , w_8702 , w_8703 , w_8704 , w_8705 , w_8706 , w_8707 , w_8708 , w_8709 , 
		w_8710 , w_8711 , w_8712 , w_8713 , w_8714 , w_8715 , w_8716 , w_8717 , w_8718 , w_8719 , 
		w_8720 , w_8721 , w_8722 , w_8723 , w_8724 , w_8725 , w_8726 , w_8727 , w_8728 , w_8729 , 
		w_8730 , w_8731 , w_8732 , w_8733 , w_8734 , w_8735 , w_8736 , w_8737 , w_8738 , w_8739 , 
		w_8740 , w_8741 , w_8742 , w_8743 , w_8744 , w_8745 , w_8746 , w_8747 , w_8748 , w_8749 , 
		w_8750 , w_8751 , w_8752 , w_8753 , w_8754 , w_8755 , w_8756 , w_8757 , w_8758 , w_8759 , 
		w_8760 , w_8761 , w_8762 , w_8763 , w_8764 , w_8765 , w_8766 , w_8767 , w_8768 , w_8769 , 
		w_8770 , w_8771 , w_8772 , w_8773 , w_8774 , w_8775 , w_8776 , w_8777 , w_8778 , w_8779 , 
		w_8780 , w_8781 , w_8782 , w_8783 , w_8784 , w_8785 , w_8786 , w_8787 , w_8788 , w_8789 , 
		w_8790 , w_8791 , w_8792 , w_8793 , w_8794 , w_8795 , w_8796 , w_8797 , w_8798 , w_8799 , 
		w_8800 , w_8801 , w_8802 , w_8803 , w_8804 , w_8805 , w_8806 , w_8807 , w_8808 , w_8809 , 
		w_8810 , w_8811 , w_8812 , w_8813 , w_8814 , w_8815 , w_8816 , w_8817 , w_8818 , w_8819 , 
		w_8820 , w_8821 , w_8822 , w_8823 , w_8824 , w_8825 , w_8826 , w_8827 , w_8828 , w_8829 , 
		w_8830 , w_8831 , w_8832 , w_8833 , w_8834 , w_8835 , w_8836 , w_8837 , w_8838 , w_8839 , 
		w_8840 , w_8841 , w_8842 , w_8843 , w_8844 , w_8845 , w_8846 , w_8847 , w_8848 , w_8849 , 
		w_8850 , w_8851 , w_8852 , w_8853 , w_8854 , w_8855 , w_8856 , w_8857 , w_8858 , w_8859 , 
		w_8860 , w_8861 , w_8862 , w_8863 , w_8864 , w_8865 , w_8866 , w_8867 , w_8868 , w_8869 , 
		w_8870 , w_8871 , w_8872 , w_8873 , w_8874 , w_8875 , w_8876 , w_8877 , w_8878 , w_8879 , 
		w_8880 , w_8881 , w_8882 , w_8883 , w_8884 , w_8885 , w_8886 , w_8887 , w_8888 , w_8889 , 
		w_8890 , w_8891 , w_8892 , w_8893 , w_8894 , w_8895 , w_8896 , w_8897 , w_8898 , w_8899 , 
		w_8900 , w_8901 , w_8902 , w_8903 , w_8904 , w_8905 , w_8906 , w_8907 , w_8908 , w_8909 , 
		w_8910 , w_8911 , w_8912 , w_8913 , w_8914 , w_8915 , w_8916 , w_8917 , w_8918 , w_8919 , 
		w_8920 , w_8921 , w_8922 , w_8923 , w_8924 , w_8925 , w_8926 , w_8927 , w_8928 , w_8929 , 
		w_8930 , w_8931 , w_8932 , w_8933 , w_8934 , w_8935 , w_8936 , w_8937 , w_8938 , w_8939 , 
		w_8940 , w_8941 , w_8942 , w_8943 , w_8944 , w_8945 , w_8946 , w_8947 , w_8948 , w_8949 , 
		w_8950 , w_8951 , w_8952 , w_8953 , w_8954 , w_8955 , w_8956 , w_8957 , w_8958 , w_8959 , 
		w_8960 , w_8961 , w_8962 , w_8963 , w_8964 , w_8965 , w_8966 , w_8967 , w_8968 , w_8969 , 
		w_8970 , w_8971 , w_8972 , w_8973 , w_8974 , w_8975 , w_8976 , w_8977 , w_8978 , w_8979 , 
		w_8980 , w_8981 , w_8982 , w_8983 , w_8984 , w_8985 , w_8986 , w_8987 , w_8988 , w_8989 , 
		w_8990 , w_8991 , w_8992 , w_8993 , w_8994 , w_8995 , w_8996 , w_8997 , w_8998 , w_8999 , 
		w_9000 , w_9001 , w_9002 , w_9003 , w_9004 , w_9005 , w_9006 , w_9007 , w_9008 , w_9009 , 
		w_9010 , w_9011 , w_9012 , w_9013 , w_9014 , w_9015 , w_9016 , w_9017 , w_9018 , w_9019 , 
		w_9020 , w_9021 , w_9022 , w_9023 , w_9024 , w_9025 , w_9026 , w_9027 , w_9028 , w_9029 , 
		w_9030 , w_9031 , w_9032 , w_9033 , w_9034 , w_9035 , w_9036 , w_9037 , w_9038 , w_9039 , 
		w_9040 , w_9041 , w_9042 , w_9043 , w_9044 , w_9045 , w_9046 , w_9047 , w_9048 , w_9049 , 
		w_9050 , w_9051 , w_9052 , w_9053 , w_9054 , w_9055 , w_9056 , w_9057 , w_9058 , w_9059 , 
		w_9060 , w_9061 , w_9062 , w_9063 , w_9064 , w_9065 , w_9066 , w_9067 , w_9068 , w_9069 , 
		w_9070 , w_9071 , w_9072 , w_9073 , w_9074 , w_9075 , w_9076 , w_9077 , w_9078 , w_9079 , 
		w_9080 , w_9081 , w_9082 , w_9083 , w_9084 , w_9085 , w_9086 , w_9087 , w_9088 , w_9089 , 
		w_9090 , w_9091 , w_9092 , w_9093 , w_9094 , w_9095 , w_9096 , w_9097 , w_9098 , w_9099 , 
		w_9100 , w_9101 , w_9102 , w_9103 , w_9104 , w_9105 , w_9106 , w_9107 , w_9108 , w_9109 , 
		w_9110 , w_9111 , w_9112 , w_9113 , w_9114 , w_9115 , w_9116 , w_9117 , w_9118 , w_9119 , 
		w_9120 , w_9121 , w_9122 , w_9123 , w_9124 , w_9125 , w_9126 , w_9127 , w_9128 , w_9129 , 
		w_9130 , w_9131 , w_9132 , w_9133 , w_9134 , w_9135 , w_9136 , w_9137 , w_9138 , w_9139 , 
		w_9140 , w_9141 , w_9142 , w_9143 , w_9144 , w_9145 , w_9146 , w_9147 , w_9148 , w_9149 , 
		w_9150 , w_9151 , w_9152 , w_9153 , w_9154 , w_9155 , w_9156 , w_9157 , w_9158 , w_9159 , 
		w_9160 , w_9161 , w_9162 , w_9163 , w_9164 , w_9165 , w_9166 , w_9167 , w_9168 , w_9169 , 
		w_9170 , w_9171 , w_9172 , w_9173 , w_9174 , w_9175 , w_9176 , w_9177 , w_9178 , w_9179 , 
		w_9180 , w_9181 , w_9182 , w_9183 , w_9184 , w_9185 , w_9186 , w_9187 , w_9188 , w_9189 , 
		w_9190 , w_9191 , w_9192 , w_9193 , w_9194 , w_9195 , w_9196 , w_9197 , w_9198 , w_9199 , 
		w_9200 , w_9201 , w_9202 , w_9203 , w_9204 , w_9205 , w_9206 , w_9207 , w_9208 , w_9209 , 
		w_9210 , w_9211 , w_9212 , w_9213 , w_9214 , w_9215 , w_9216 , w_9217 , w_9218 , w_9219 , 
		w_9220 , w_9221 , w_9222 , w_9223 , w_9224 , w_9225 , w_9226 , w_9227 , w_9228 , w_9229 , 
		w_9230 , w_9231 , w_9232 , w_9233 , w_9234 , w_9235 , w_9236 , w_9237 , w_9238 , w_9239 , 
		w_9240 , w_9241 , w_9242 , w_9243 , w_9244 , w_9245 , w_9246 , w_9247 , w_9248 , w_9249 , 
		w_9250 , w_9251 , w_9252 , w_9253 , w_9254 , w_9255 , w_9256 , w_9257 , w_9258 , w_9259 , 
		w_9260 , w_9261 , w_9262 , w_9263 , w_9264 , w_9265 , w_9266 , w_9267 , w_9268 , w_9269 , 
		w_9270 , w_9271 , w_9272 , w_9273 , w_9274 , w_9275 , w_9276 , w_9277 , w_9278 , w_9279 , 
		w_9280 , w_9281 , w_9282 , w_9283 , w_9284 , w_9285 , w_9286 , w_9287 , w_9288 , w_9289 , 
		w_9290 , w_9291 , w_9292 , w_9293 , w_9294 , w_9295 , w_9296 , w_9297 , w_9298 , w_9299 , 
		w_9300 , w_9301 , w_9302 , w_9303 , w_9304 , w_9305 , w_9306 , w_9307 , w_9308 , w_9309 , 
		w_9310 , w_9311 , w_9312 , w_9313 , w_9314 , w_9315 , w_9316 , w_9317 , w_9318 , w_9319 , 
		w_9320 , w_9321 , w_9322 , w_9323 , w_9324 , w_9325 , w_9326 , w_9327 , w_9328 , w_9329 , 
		w_9330 , w_9331 , w_9332 , w_9333 , w_9334 , w_9335 , w_9336 , w_9337 , w_9338 , w_9339 , 
		w_9340 , w_9341 , w_9342 , w_9343 , w_9344 , w_9345 , w_9346 , w_9347 , w_9348 , w_9349 , 
		w_9350 , w_9351 , w_9352 , w_9353 , w_9354 , w_9355 , w_9356 , w_9357 , w_9358 , w_9359 , 
		w_9360 , w_9361 , w_9362 , w_9363 , w_9364 , w_9365 , w_9366 , w_9367 , w_9368 , w_9369 , 
		w_9370 , w_9371 , w_9372 , w_9373 , w_9374 , w_9375 , w_9376 , w_9377 , w_9378 , w_9379 , 
		w_9380 , w_9381 , w_9382 , w_9383 , w_9384 , w_9385 , w_9386 , w_9387 , w_9388 , w_9389 , 
		w_9390 , w_9391 , w_9392 , w_9393 , w_9394 , w_9395 , w_9396 , w_9397 , w_9398 , w_9399 , 
		w_9400 , w_9401 , w_9402 , w_9403 , w_9404 , w_9405 , w_9406 , w_9407 , w_9408 , w_9409 , 
		w_9410 , w_9411 , w_9412 , w_9413 , w_9414 , w_9415 , w_9416 , w_9417 , w_9418 , w_9419 , 
		w_9420 , w_9421 , w_9422 , w_9423 , w_9424 , w_9425 , w_9426 , w_9427 , w_9428 , w_9429 , 
		w_9430 , w_9431 , w_9432 , w_9433 , w_9434 , w_9435 , w_9436 , w_9437 , w_9438 , w_9439 , 
		w_9440 , w_9441 , w_9442 , w_9443 , w_9444 , w_9445 , w_9446 , w_9447 , w_9448 , w_9449 , 
		w_9450 , w_9451 , w_9452 , w_9453 , w_9454 , w_9455 , w_9456 , w_9457 , w_9458 , w_9459 , 
		w_9460 , w_9461 , w_9462 , w_9463 , w_9464 , w_9465 , w_9466 , w_9467 , w_9468 , w_9469 , 
		w_9470 , w_9471 , w_9472 , w_9473 , w_9474 , w_9475 , w_9476 , w_9477 , w_9478 , w_9479 , 
		w_9480 , w_9481 , w_9482 , w_9483 , w_9484 , w_9485 , w_9486 , w_9487 , w_9488 , w_9489 , 
		w_9490 , w_9491 , w_9492 , w_9493 , w_9494 , w_9495 , w_9496 , w_9497 , w_9498 , w_9499 , 
		w_9500 , w_9501 , w_9502 , w_9503 , w_9504 , w_9505 , w_9506 , w_9507 , w_9508 , w_9509 , 
		w_9510 , w_9511 , w_9512 , w_9513 , w_9514 , w_9515 , w_9516 , w_9517 , w_9518 , w_9519 , 
		w_9520 , w_9521 , w_9522 , w_9523 , w_9524 , w_9525 , w_9526 , w_9527 , w_9528 , w_9529 , 
		w_9530 , w_9531 , w_9532 , w_9533 , w_9534 , w_9535 , w_9536 , w_9537 , w_9538 , w_9539 , 
		w_9540 , w_9541 , w_9542 , w_9543 , w_9544 , w_9545 , w_9546 , w_9547 , w_9548 , w_9549 , 
		w_9550 , w_9551 , w_9552 , w_9553 , w_9554 , w_9555 , w_9556 , w_9557 , w_9558 , w_9559 , 
		w_9560 , w_9561 , w_9562 , w_9563 , w_9564 , w_9565 , w_9566 , w_9567 , w_9568 , w_9569 , 
		w_9570 , w_9571 , w_9572 , w_9573 , w_9574 , w_9575 , w_9576 , w_9577 , w_9578 , w_9579 , 
		w_9580 , w_9581 , w_9582 , w_9583 , w_9584 , w_9585 , w_9586 , w_9587 , w_9588 , w_9589 , 
		w_9590 , w_9591 , w_9592 , w_9593 , w_9594 , w_9595 , w_9596 , w_9597 , w_9598 , w_9599 , 
		w_9600 , w_9601 , w_9602 , w_9603 , w_9604 , w_9605 , w_9606 , w_9607 , w_9608 , w_9609 , 
		w_9610 , w_9611 , w_9612 , w_9613 , w_9614 , w_9615 , w_9616 , w_9617 , w_9618 , w_9619 , 
		w_9620 , w_9621 , w_9622 , w_9623 , w_9624 , w_9625 , w_9626 , w_9627 , w_9628 , w_9629 , 
		w_9630 , w_9631 , w_9632 , w_9633 , w_9634 , w_9635 , w_9636 , w_9637 , w_9638 , w_9639 , 
		w_9640 , w_9641 , w_9642 , w_9643 , w_9644 , w_9645 , w_9646 , w_9647 , w_9648 , w_9649 , 
		w_9650 , w_9651 , w_9652 , w_9653 , w_9654 , w_9655 , w_9656 , w_9657 , w_9658 , w_9659 , 
		w_9660 , w_9661 , w_9662 , w_9663 , w_9664 , w_9665 , w_9666 , w_9667 , w_9668 , w_9669 , 
		w_9670 , w_9671 , w_9672 , w_9673 , w_9674 , w_9675 , w_9676 , w_9677 , w_9678 , w_9679 , 
		w_9680 , w_9681 , w_9682 , w_9683 , w_9684 , w_9685 , w_9686 , w_9687 , w_9688 , w_9689 , 
		w_9690 , w_9691 , w_9692 , w_9693 , w_9694 , w_9695 , w_9696 , w_9697 , w_9698 , w_9699 , 
		w_9700 , w_9701 , w_9702 , w_9703 , w_9704 , w_9705 , w_9706 , w_9707 , w_9708 , w_9709 , 
		w_9710 , w_9711 , w_9712 , w_9713 , w_9714 , w_9715 , w_9716 , w_9717 , w_9718 , w_9719 , 
		w_9720 , w_9721 , w_9722 , w_9723 , w_9724 , w_9725 , w_9726 , w_9727 , w_9728 , w_9729 , 
		w_9730 , w_9731 , w_9732 , w_9733 , w_9734 , w_9735 , w_9736 , w_9737 , w_9738 , w_9739 , 
		w_9740 , w_9741 , w_9742 , w_9743 , w_9744 , w_9745 , w_9746 , w_9747 , w_9748 , w_9749 , 
		w_9750 , w_9751 , w_9752 , w_9753 , w_9754 , w_9755 , w_9756 , w_9757 , w_9758 , w_9759 , 
		w_9760 , w_9761 , w_9762 , w_9763 , w_9764 , w_9765 , w_9766 , w_9767 , w_9768 , w_9769 , 
		w_9770 , w_9771 , w_9772 , w_9773 , w_9774 , w_9775 , w_9776 , w_9777 , w_9778 , w_9779 , 
		w_9780 , w_9781 , w_9782 , w_9783 , w_9784 , w_9785 , w_9786 , w_9787 , w_9788 , w_9789 , 
		w_9790 , w_9791 , w_9792 , w_9793 , w_9794 , w_9795 , w_9796 , w_9797 , w_9798 , w_9799 , 
		w_9800 , w_9801 , w_9802 , w_9803 , w_9804 , w_9805 , w_9806 , w_9807 , w_9808 , w_9809 , 
		w_9810 , w_9811 , w_9812 , w_9813 , w_9814 , w_9815 , w_9816 , w_9817 , w_9818 , w_9819 , 
		w_9820 , w_9821 , w_9822 , w_9823 , w_9824 , w_9825 , w_9826 , w_9827 , w_9828 , w_9829 , 
		w_9830 , w_9831 , w_9832 , w_9833 , w_9834 , w_9835 , w_9836 , w_9837 , w_9838 , w_9839 , 
		w_9840 , w_9841 , w_9842 , w_9843 , w_9844 , w_9845 , w_9846 , w_9847 , w_9848 , w_9849 , 
		w_9850 , w_9851 , w_9852 , w_9853 , w_9854 , w_9855 , w_9856 , w_9857 , w_9858 , w_9859 , 
		w_9860 , w_9861 , w_9862 , w_9863 , w_9864 , w_9865 , w_9866 , w_9867 , w_9868 , w_9869 , 
		w_9870 , w_9871 , w_9872 , w_9873 , w_9874 , w_9875 , w_9876 , w_9877 , w_9878 , w_9879 , 
		w_9880 , w_9881 , w_9882 , w_9883 , w_9884 , w_9885 , w_9886 , w_9887 , w_9888 , w_9889 , 
		w_9890 , w_9891 , w_9892 , w_9893 , w_9894 , w_9895 , w_9896 , w_9897 , w_9898 , w_9899 , 
		w_9900 , w_9901 , w_9902 , w_9903 , w_9904 , w_9905 , w_9906 , w_9907 , w_9908 , w_9909 , 
		w_9910 , w_9911 , w_9912 , w_9913 , w_9914 , w_9915 , w_9916 , w_9917 , w_9918 , w_9919 , 
		w_9920 , w_9921 , w_9922 , w_9923 , w_9924 , w_9925 , w_9926 , w_9927 , w_9928 , w_9929 , 
		w_9930 , w_9931 , w_9932 , w_9933 , w_9934 , w_9935 , w_9936 , w_9937 , w_9938 , w_9939 , 
		w_9940 , w_9941 , w_9942 , w_9943 , w_9944 , w_9945 , w_9946 , w_9947 , w_9948 , w_9949 , 
		w_9950 , w_9951 , w_9952 , w_9953 , w_9954 , w_9955 , w_9956 , w_9957 , w_9958 , w_9959 , 
		w_9960 , w_9961 , w_9962 , w_9963 , w_9964 , w_9965 , w_9966 , w_9967 , w_9968 , w_9969 , 
		w_9970 , w_9971 , w_9972 , w_9973 , w_9974 , w_9975 , w_9976 , w_9977 , w_9978 , w_9979 , 
		w_9980 , w_9981 , w_9982 , w_9983 , w_9984 , w_9985 , w_9986 , w_9987 , w_9988 , w_9989 , 
		w_9990 , w_9991 , w_9992 , w_9993 , w_9994 , w_9995 , w_9996 , w_9997 , w_9998 , w_9999 , 
		w_10000 , w_10001 , w_10002 , w_10003 , w_10004 , w_10005 , w_10006 , w_10007 , w_10008 , w_10009 , 
		w_10010 , w_10011 , w_10012 , w_10013 , w_10014 , w_10015 , w_10016 , w_10017 , w_10018 , w_10019 , 
		w_10020 , w_10021 , w_10022 , w_10023 , w_10024 , w_10025 , w_10026 , w_10027 , w_10028 , w_10029 , 
		w_10030 , w_10031 , w_10032 , w_10033 , w_10034 , w_10035 , w_10036 , w_10037 , w_10038 , w_10039 , 
		w_10040 , w_10041 , w_10042 , w_10043 , w_10044 , w_10045 , w_10046 , w_10047 , w_10048 , w_10049 , 
		w_10050 , w_10051 , w_10052 , w_10053 , w_10054 , w_10055 , w_10056 , w_10057 , w_10058 , w_10059 , 
		w_10060 , w_10061 , w_10062 , w_10063 , w_10064 , w_10065 , w_10066 , w_10067 , w_10068 , w_10069 , 
		w_10070 , w_10071 , w_10072 , w_10073 , w_10074 , w_10075 , w_10076 , w_10077 , w_10078 , w_10079 , 
		w_10080 , w_10081 , w_10082 , w_10083 , w_10084 , w_10085 , w_10086 , w_10087 , w_10088 , w_10089 , 
		w_10090 , w_10091 , w_10092 , w_10093 , w_10094 , w_10095 , w_10096 , w_10097 , w_10098 , w_10099 , 
		w_10100 , w_10101 , w_10102 , w_10103 , w_10104 , w_10105 , w_10106 , w_10107 , w_10108 , w_10109 , 
		w_10110 , w_10111 , w_10112 , w_10113 , w_10114 , w_10115 , w_10116 , w_10117 , w_10118 , w_10119 , 
		w_10120 , w_10121 , w_10122 , w_10123 , w_10124 , w_10125 , w_10126 , w_10127 , w_10128 , w_10129 , 
		w_10130 , w_10131 , w_10132 , w_10133 , w_10134 , w_10135 , w_10136 , w_10137 , w_10138 , w_10139 , 
		w_10140 , w_10141 , w_10142 , w_10143 , w_10144 , w_10145 , w_10146 , w_10147 , w_10148 , w_10149 , 
		w_10150 , w_10151 , w_10152 , w_10153 , w_10154 , w_10155 , w_10156 , w_10157 , w_10158 , w_10159 , 
		w_10160 , w_10161 , w_10162 , w_10163 , w_10164 , w_10165 , w_10166 , w_10167 , w_10168 , w_10169 , 
		w_10170 , w_10171 , w_10172 , w_10173 , w_10174 , w_10175 , w_10176 , w_10177 , w_10178 , w_10179 , 
		w_10180 , w_10181 , w_10182 , w_10183 , w_10184 , w_10185 , w_10186 , w_10187 , w_10188 , w_10189 , 
		w_10190 , w_10191 , w_10192 , w_10193 , w_10194 , w_10195 , w_10196 , w_10197 , w_10198 , w_10199 , 
		w_10200 , w_10201 , w_10202 , w_10203 , w_10204 , w_10205 , w_10206 , w_10207 , w_10208 , w_10209 , 
		w_10210 , w_10211 , w_10212 , w_10213 , w_10214 , w_10215 , w_10216 , w_10217 , w_10218 , w_10219 , 
		w_10220 , w_10221 , w_10222 , w_10223 , w_10224 , w_10225 , w_10226 , w_10227 , w_10228 , w_10229 , 
		w_10230 , w_10231 , w_10232 , w_10233 , w_10234 , w_10235 , w_10236 , w_10237 , w_10238 , w_10239 , 
		w_10240 , w_10241 , w_10242 , w_10243 , w_10244 , w_10245 , w_10246 , w_10247 , w_10248 , w_10249 , 
		w_10250 , w_10251 , w_10252 , w_10253 , w_10254 , w_10255 , w_10256 , w_10257 , w_10258 , w_10259 , 
		w_10260 , w_10261 , w_10262 , w_10263 , w_10264 , w_10265 , w_10266 , w_10267 , w_10268 , w_10269 , 
		w_10270 , w_10271 , w_10272 , w_10273 , w_10274 , w_10275 , w_10276 , w_10277 , w_10278 , w_10279 , 
		w_10280 , w_10281 , w_10282 , w_10283 , w_10284 , w_10285 , w_10286 , w_10287 , w_10288 , w_10289 , 
		w_10290 , w_10291 , w_10292 , w_10293 , w_10294 , w_10295 , w_10296 , w_10297 , w_10298 , w_10299 , 
		w_10300 , w_10301 , w_10302 , w_10303 , w_10304 , w_10305 , w_10306 , w_10307 , w_10308 , w_10309 , 
		w_10310 , w_10311 , w_10312 , w_10313 , w_10314 , w_10315 , w_10316 , w_10317 , w_10318 , w_10319 , 
		w_10320 , w_10321 , w_10322 , w_10323 , w_10324 , w_10325 , w_10326 , w_10327 , w_10328 , w_10329 , 
		w_10330 , w_10331 , w_10332 , w_10333 , w_10334 , w_10335 , w_10336 , w_10337 , w_10338 , w_10339 , 
		w_10340 , w_10341 , w_10342 , w_10343 , w_10344 , w_10345 , w_10346 , w_10347 , w_10348 , w_10349 , 
		w_10350 , w_10351 , w_10352 , w_10353 , w_10354 , w_10355 , w_10356 , w_10357 , w_10358 , w_10359 , 
		w_10360 , w_10361 , w_10362 , w_10363 , w_10364 , w_10365 , w_10366 , w_10367 , w_10368 , w_10369 , 
		w_10370 , w_10371 , w_10372 , w_10373 , w_10374 , w_10375 , w_10376 , w_10377 , w_10378 , w_10379 , 
		w_10380 , w_10381 , w_10382 , w_10383 , w_10384 , w_10385 , w_10386 , w_10387 , w_10388 , w_10389 , 
		w_10390 , w_10391 , w_10392 , w_10393 , w_10394 , w_10395 , w_10396 , w_10397 , w_10398 , w_10399 , 
		w_10400 , w_10401 , w_10402 , w_10403 , w_10404 , w_10405 , w_10406 , w_10407 , w_10408 , w_10409 , 
		w_10410 , w_10411 , w_10412 , w_10413 , w_10414 , w_10415 , w_10416 , w_10417 , w_10418 , w_10419 , 
		w_10420 , w_10421 , w_10422 , w_10423 , w_10424 , w_10425 , w_10426 , w_10427 , w_10428 , w_10429 , 
		w_10430 , w_10431 , w_10432 , w_10433 , w_10434 , w_10435 , w_10436 , w_10437 , w_10438 , w_10439 , 
		w_10440 , w_10441 , w_10442 , w_10443 , w_10444 , w_10445 , w_10446 , w_10447 , w_10448 , w_10449 , 
		w_10450 , w_10451 , w_10452 , w_10453 , w_10454 , w_10455 , w_10456 , w_10457 , w_10458 , w_10459 , 
		w_10460 , w_10461 , w_10462 , w_10463 , w_10464 , w_10465 , w_10466 , w_10467 , w_10468 , w_10469 , 
		w_10470 , w_10471 , w_10472 , w_10473 , w_10474 , w_10475 , w_10476 , w_10477 , w_10478 , w_10479 , 
		w_10480 , w_10481 , w_10482 , w_10483 , w_10484 , w_10485 , w_10486 , w_10487 , w_10488 , w_10489 , 
		w_10490 , w_10491 , w_10492 , w_10493 , w_10494 , w_10495 , w_10496 , w_10497 , w_10498 , w_10499 , 
		w_10500 , w_10501 , w_10502 , w_10503 , w_10504 , w_10505 , w_10506 , w_10507 , w_10508 , w_10509 , 
		w_10510 , w_10511 , w_10512 , w_10513 , w_10514 , w_10515 , w_10516 , w_10517 , w_10518 , w_10519 , 
		w_10520 , w_10521 , w_10522 , w_10523 , w_10524 , w_10525 , w_10526 , w_10527 , w_10528 , w_10529 , 
		w_10530 , w_10531 , w_10532 , w_10533 , w_10534 , w_10535 , w_10536 , w_10537 , w_10538 , w_10539 , 
		w_10540 , w_10541 , w_10542 , w_10543 , w_10544 , w_10545 , w_10546 , w_10547 , w_10548 , w_10549 , 
		w_10550 , w_10551 , w_10552 , w_10553 , w_10554 , w_10555 , w_10556 , w_10557 , w_10558 , w_10559 , 
		w_10560 , w_10561 , w_10562 , w_10563 , w_10564 , w_10565 , w_10566 , w_10567 , w_10568 , w_10569 , 
		w_10570 , w_10571 , w_10572 , w_10573 , w_10574 , w_10575 , w_10576 , w_10577 , w_10578 , w_10579 , 
		w_10580 , w_10581 , w_10582 , w_10583 , w_10584 , w_10585 , w_10586 , w_10587 , w_10588 , w_10589 , 
		w_10590 , w_10591 , w_10592 , w_10593 , w_10594 , w_10595 , w_10596 , w_10597 , w_10598 , w_10599 , 
		w_10600 , w_10601 , w_10602 , w_10603 , w_10604 , w_10605 , w_10606 , w_10607 , w_10608 , w_10609 , 
		w_10610 , w_10611 , w_10612 , w_10613 , w_10614 , w_10615 , w_10616 , w_10617 , w_10618 , w_10619 , 
		w_10620 , w_10621 , w_10622 , w_10623 , w_10624 , w_10625 , w_10626 , w_10627 , w_10628 , w_10629 , 
		w_10630 , w_10631 , w_10632 , w_10633 , w_10634 , w_10635 , w_10636 , w_10637 , w_10638 , w_10639 , 
		w_10640 , w_10641 , w_10642 , w_10643 , w_10644 , w_10645 , w_10646 , w_10647 , w_10648 , w_10649 , 
		w_10650 , w_10651 , w_10652 , w_10653 , w_10654 , w_10655 , w_10656 , w_10657 , w_10658 , w_10659 , 
		w_10660 , w_10661 , w_10662 , w_10663 , w_10664 , w_10665 , w_10666 , w_10667 , w_10668 , w_10669 , 
		w_10670 , w_10671 , w_10672 , w_10673 , w_10674 , w_10675 , w_10676 , w_10677 , w_10678 , w_10679 , 
		w_10680 , w_10681 , w_10682 , w_10683 , w_10684 , w_10685 , w_10686 , w_10687 , w_10688 , w_10689 , 
		w_10690 , w_10691 , w_10692 , w_10693 , w_10694 , w_10695 , w_10696 , w_10697 , w_10698 , w_10699 , 
		w_10700 , w_10701 , w_10702 , w_10703 , w_10704 , w_10705 , w_10706 , w_10707 , w_10708 , w_10709 , 
		w_10710 , w_10711 , w_10712 , w_10713 , w_10714 , w_10715 , w_10716 , w_10717 , w_10718 , w_10719 , 
		w_10720 , w_10721 , w_10722 , w_10723 , w_10724 , w_10725 , w_10726 , w_10727 , w_10728 , w_10729 , 
		w_10730 , w_10731 , w_10732 , w_10733 , w_10734 , w_10735 , w_10736 , w_10737 , w_10738 , w_10739 , 
		w_10740 , w_10741 , w_10742 , w_10743 , w_10744 , w_10745 , w_10746 , w_10747 , w_10748 , w_10749 , 
		w_10750 , w_10751 , w_10752 , w_10753 , w_10754 , w_10755 , w_10756 , w_10757 , w_10758 , w_10759 , 
		w_10760 , w_10761 , w_10762 , w_10763 , w_10764 , w_10765 , w_10766 , w_10767 , w_10768 , w_10769 , 
		w_10770 , w_10771 , w_10772 , w_10773 , w_10774 , w_10775 , w_10776 , w_10777 , w_10778 , w_10779 , 
		w_10780 , w_10781 , w_10782 , w_10783 , w_10784 , w_10785 , w_10786 , w_10787 , w_10788 , w_10789 , 
		w_10790 , w_10791 , w_10792 , w_10793 , w_10794 , w_10795 , w_10796 , w_10797 , w_10798 , w_10799 , 
		w_10800 , w_10801 , w_10802 , w_10803 , w_10804 , w_10805 , w_10806 , w_10807 , w_10808 , w_10809 , 
		w_10810 , w_10811 , w_10812 , w_10813 , w_10814 , w_10815 , w_10816 , w_10817 , w_10818 , w_10819 , 
		w_10820 , w_10821 , w_10822 , w_10823 , w_10824 , w_10825 , w_10826 , w_10827 , w_10828 , w_10829 , 
		w_10830 , w_10831 , w_10832 , w_10833 , w_10834 , w_10835 , w_10836 , w_10837 , w_10838 , w_10839 , 
		w_10840 , w_10841 , w_10842 , w_10843 , w_10844 , w_10845 , w_10846 , w_10847 , w_10848 , w_10849 , 
		w_10850 , w_10851 , w_10852 , w_10853 , w_10854 , w_10855 , w_10856 , w_10857 , w_10858 , w_10859 , 
		w_10860 , w_10861 , w_10862 , w_10863 , w_10864 , w_10865 , w_10866 , w_10867 , w_10868 , w_10869 , 
		w_10870 , w_10871 , w_10872 , w_10873 , w_10874 , w_10875 , w_10876 , w_10877 , w_10878 , w_10879 , 
		w_10880 , w_10881 , w_10882 , w_10883 , w_10884 , w_10885 , w_10886 , w_10887 , w_10888 , w_10889 , 
		w_10890 , w_10891 , w_10892 , w_10893 , w_10894 , w_10895 , w_10896 , w_10897 , w_10898 , w_10899 , 
		w_10900 , w_10901 , w_10902 , w_10903 , w_10904 , w_10905 , w_10906 , w_10907 , w_10908 , w_10909 , 
		w_10910 , w_10911 , w_10912 , w_10913 , w_10914 , w_10915 , w_10916 , w_10917 , w_10918 , w_10919 , 
		w_10920 , w_10921 , w_10922 , w_10923 , w_10924 , w_10925 , w_10926 , w_10927 , w_10928 , w_10929 , 
		w_10930 , w_10931 , w_10932 , w_10933 , w_10934 , w_10935 , w_10936 , w_10937 , w_10938 , w_10939 , 
		w_10940 , w_10941 , w_10942 , w_10943 , w_10944 , w_10945 , w_10946 , w_10947 , w_10948 , w_10949 , 
		w_10950 , w_10951 , w_10952 , w_10953 , w_10954 , w_10955 , w_10956 , w_10957 , w_10958 , w_10959 , 
		w_10960 , w_10961 , w_10962 , w_10963 , w_10964 , w_10965 , w_10966 , w_10967 , w_10968 , w_10969 , 
		w_10970 , w_10971 , w_10972 , w_10973 , w_10974 , w_10975 , w_10976 , w_10977 , w_10978 , w_10979 , 
		w_10980 , w_10981 , w_10982 , w_10983 , w_10984 , w_10985 , w_10986 , w_10987 , w_10988 , w_10989 , 
		w_10990 , w_10991 , w_10992 , w_10993 , w_10994 , w_10995 , w_10996 , w_10997 , w_10998 , w_10999 , 
		w_11000 , w_11001 , w_11002 , w_11003 , w_11004 , w_11005 , w_11006 , w_11007 , w_11008 , w_11009 , 
		w_11010 , w_11011 , w_11012 , w_11013 , w_11014 , w_11015 , w_11016 , w_11017 , w_11018 , w_11019 , 
		w_11020 , w_11021 , w_11022 , w_11023 , w_11024 , w_11025 , w_11026 , w_11027 , w_11028 , w_11029 , 
		w_11030 , w_11031 , w_11032 , w_11033 , w_11034 , w_11035 , w_11036 , w_11037 , w_11038 , w_11039 , 
		w_11040 , w_11041 , w_11042 , w_11043 , w_11044 , w_11045 , w_11046 , w_11047 , w_11048 , w_11049 , 
		w_11050 , w_11051 , w_11052 , w_11053 , w_11054 , w_11055 , w_11056 , w_11057 , w_11058 , w_11059 , 
		w_11060 , w_11061 , w_11062 , w_11063 , w_11064 , w_11065 , w_11066 , w_11067 , w_11068 , w_11069 , 
		w_11070 , w_11071 , w_11072 , w_11073 , w_11074 , w_11075 , w_11076 , w_11077 , w_11078 , w_11079 , 
		w_11080 , w_11081 , w_11082 , w_11083 , w_11084 , w_11085 , w_11086 , w_11087 , w_11088 , w_11089 , 
		w_11090 , w_11091 , w_11092 , w_11093 , w_11094 , w_11095 , w_11096 , w_11097 , w_11098 , w_11099 , 
		w_11100 , w_11101 , w_11102 , w_11103 , w_11104 , w_11105 , w_11106 , w_11107 , w_11108 , w_11109 , 
		w_11110 , w_11111 , w_11112 , w_11113 , w_11114 , w_11115 , w_11116 , w_11117 , w_11118 , w_11119 , 
		w_11120 , w_11121 , w_11122 , w_11123 , w_11124 , w_11125 , w_11126 , w_11127 , w_11128 , w_11129 , 
		w_11130 , w_11131 , w_11132 , w_11133 , w_11134 , w_11135 , w_11136 , w_11137 , w_11138 , w_11139 , 
		w_11140 , w_11141 , w_11142 , w_11143 , w_11144 , w_11145 , w_11146 , w_11147 , w_11148 , w_11149 , 
		w_11150 , w_11151 , w_11152 , w_11153 , w_11154 , w_11155 , w_11156 , w_11157 , w_11158 , w_11159 , 
		w_11160 , w_11161 , w_11162 , w_11163 , w_11164 , w_11165 , w_11166 , w_11167 , w_11168 , w_11169 , 
		w_11170 , w_11171 , w_11172 , w_11173 , w_11174 , w_11175 , w_11176 , w_11177 , w_11178 , w_11179 , 
		w_11180 , w_11181 , w_11182 , w_11183 , w_11184 , w_11185 , w_11186 , w_11187 , w_11188 , w_11189 , 
		w_11190 , w_11191 , w_11192 , w_11193 , w_11194 , w_11195 , w_11196 , w_11197 , w_11198 , w_11199 , 
		w_11200 , w_11201 , w_11202 , w_11203 , w_11204 , w_11205 , w_11206 , w_11207 , w_11208 , w_11209 , 
		w_11210 , w_11211 , w_11212 , w_11213 , w_11214 , w_11215 , w_11216 , w_11217 , w_11218 , w_11219 , 
		w_11220 , w_11221 , w_11222 , w_11223 , w_11224 , w_11225 , w_11226 , w_11227 , w_11228 , w_11229 , 
		w_11230 , w_11231 , w_11232 , w_11233 , w_11234 , w_11235 , w_11236 , w_11237 , w_11238 , w_11239 , 
		w_11240 , w_11241 , w_11242 , w_11243 , w_11244 , w_11245 , w_11246 , w_11247 , w_11248 , w_11249 , 
		w_11250 , w_11251 , w_11252 , w_11253 , w_11254 , w_11255 , w_11256 , w_11257 , w_11258 , w_11259 , 
		w_11260 , w_11261 , w_11262 , w_11263 , w_11264 , w_11265 , w_11266 , w_11267 , w_11268 , w_11269 , 
		w_11270 , w_11271 , w_11272 , w_11273 , w_11274 , w_11275 , w_11276 , w_11277 , w_11278 , w_11279 , 
		w_11280 , w_11281 , w_11282 , w_11283 , w_11284 , w_11285 , w_11286 , w_11287 , w_11288 , w_11289 , 
		w_11290 , w_11291 , w_11292 , w_11293 , w_11294 , w_11295 , w_11296 , w_11297 , w_11298 , w_11299 , 
		w_11300 , w_11301 , w_11302 , w_11303 , w_11304 , w_11305 , w_11306 , w_11307 , w_11308 , w_11309 , 
		w_11310 , w_11311 , w_11312 , w_11313 , w_11314 , w_11315 , w_11316 , w_11317 , w_11318 , w_11319 , 
		w_11320 , w_11321 , w_11322 , w_11323 , w_11324 , w_11325 , w_11326 , w_11327 , w_11328 , w_11329 , 
		w_11330 , w_11331 , w_11332 , w_11333 , w_11334 , w_11335 , w_11336 , w_11337 , w_11338 , w_11339 , 
		w_11340 , w_11341 , w_11342 , w_11343 , w_11344 , w_11345 , w_11346 , w_11347 , w_11348 , w_11349 , 
		w_11350 , w_11351 , w_11352 , w_11353 , w_11354 , w_11355 , w_11356 , w_11357 , w_11358 , w_11359 , 
		w_11360 , w_11361 , w_11362 , w_11363 , w_11364 , w_11365 , w_11366 , w_11367 , w_11368 , w_11369 , 
		w_11370 , w_11371 , w_11372 , w_11373 , w_11374 , w_11375 , w_11376 , w_11377 , w_11378 , w_11379 , 
		w_11380 , w_11381 , w_11382 , w_11383 , w_11384 , w_11385 , w_11386 , w_11387 , w_11388 , w_11389 , 
		w_11390 , w_11391 , w_11392 , w_11393 , w_11394 , w_11395 , w_11396 , w_11397 , w_11398 , w_11399 , 
		w_11400 , w_11401 , w_11402 , w_11403 , w_11404 , w_11405 , w_11406 , w_11407 , w_11408 , w_11409 , 
		w_11410 , w_11411 , w_11412 , w_11413 , w_11414 , w_11415 , w_11416 , w_11417 , w_11418 , w_11419 , 
		w_11420 , w_11421 , w_11422 , w_11423 , w_11424 , w_11425 , w_11426 , w_11427 , w_11428 , w_11429 , 
		w_11430 , w_11431 , w_11432 , w_11433 , w_11434 , w_11435 , w_11436 , w_11437 , w_11438 , w_11439 , 
		w_11440 , w_11441 , w_11442 , w_11443 , w_11444 , w_11445 , w_11446 , w_11447 , w_11448 , w_11449 , 
		w_11450 , w_11451 , w_11452 , w_11453 , w_11454 , w_11455 , w_11456 , w_11457 , w_11458 , w_11459 , 
		w_11460 , w_11461 , w_11462 , w_11463 , w_11464 , w_11465 , w_11466 , w_11467 , w_11468 , w_11469 , 
		w_11470 , w_11471 , w_11472 , w_11473 , w_11474 , w_11475 , w_11476 , w_11477 , w_11478 , w_11479 , 
		w_11480 , w_11481 , w_11482 , w_11483 , w_11484 , w_11485 , w_11486 , w_11487 , w_11488 , w_11489 , 
		w_11490 , w_11491 , w_11492 , w_11493 , w_11494 , w_11495 , w_11496 , w_11497 , w_11498 , w_11499 , 
		w_11500 , w_11501 , w_11502 , w_11503 , w_11504 , w_11505 , w_11506 , w_11507 , w_11508 , w_11509 , 
		w_11510 , w_11511 , w_11512 , w_11513 , w_11514 , w_11515 , w_11516 , w_11517 , w_11518 , w_11519 , 
		w_11520 , w_11521 , w_11522 , w_11523 , w_11524 , w_11525 , w_11526 , w_11527 , w_11528 , w_11529 , 
		w_11530 , w_11531 , w_11532 , w_11533 , w_11534 , w_11535 , w_11536 , w_11537 , w_11538 , w_11539 , 
		w_11540 , w_11541 , w_11542 , w_11543 , w_11544 , w_11545 , w_11546 , w_11547 , w_11548 , w_11549 , 
		w_11550 , w_11551 , w_11552 , w_11553 , w_11554 , w_11555 , w_11556 , w_11557 , w_11558 , w_11559 , 
		w_11560 , w_11561 , w_11562 , w_11563 , w_11564 , w_11565 , w_11566 , w_11567 , w_11568 , w_11569 , 
		w_11570 , w_11571 , w_11572 , w_11573 , w_11574 , w_11575 , w_11576 , w_11577 , w_11578 , w_11579 , 
		w_11580 , w_11581 , w_11582 , w_11583 , w_11584 , w_11585 , w_11586 , w_11587 , w_11588 , w_11589 , 
		w_11590 , w_11591 , w_11592 , w_11593 , w_11594 , w_11595 , w_11596 , w_11597 , w_11598 , w_11599 , 
		w_11600 , w_11601 , w_11602 , w_11603 , w_11604 , w_11605 , w_11606 , w_11607 , w_11608 , w_11609 , 
		w_11610 , w_11611 , w_11612 , w_11613 , w_11614 , w_11615 , w_11616 , w_11617 , w_11618 , w_11619 , 
		w_11620 , w_11621 , w_11622 , w_11623 , w_11624 , w_11625 , w_11626 , w_11627 , w_11628 , w_11629 , 
		w_11630 , w_11631 , w_11632 , w_11633 , w_11634 , w_11635 , w_11636 , w_11637 , w_11638 , w_11639 , 
		w_11640 , w_11641 , w_11642 , w_11643 , w_11644 , w_11645 , w_11646 , w_11647 , w_11648 , w_11649 , 
		w_11650 , w_11651 , w_11652 , w_11653 , w_11654 , w_11655 , w_11656 , w_11657 , w_11658 , w_11659 , 
		w_11660 , w_11661 , w_11662 , w_11663 , w_11664 , w_11665 , w_11666 , w_11667 , w_11668 , w_11669 , 
		w_11670 , w_11671 , w_11672 , w_11673 , w_11674 , w_11675 , w_11676 , w_11677 , w_11678 , w_11679 , 
		w_11680 , w_11681 , w_11682 , w_11683 , w_11684 , w_11685 , w_11686 , w_11687 , w_11688 , w_11689 , 
		w_11690 , w_11691 , w_11692 , w_11693 , w_11694 , w_11695 , w_11696 , w_11697 , w_11698 , w_11699 , 
		w_11700 , w_11701 , w_11702 , w_11703 , w_11704 , w_11705 , w_11706 , w_11707 , w_11708 , w_11709 , 
		w_11710 , w_11711 , w_11712 , w_11713 , w_11714 , w_11715 , w_11716 , w_11717 , w_11718 , w_11719 , 
		w_11720 , w_11721 , w_11722 , w_11723 , w_11724 , w_11725 , w_11726 , w_11727 , w_11728 , w_11729 , 
		w_11730 , w_11731 , w_11732 , w_11733 , w_11734 , w_11735 , w_11736 , w_11737 , w_11738 , w_11739 , 
		w_11740 , w_11741 , w_11742 , w_11743 , w_11744 , w_11745 , w_11746 , w_11747 , w_11748 , w_11749 , 
		w_11750 , w_11751 , w_11752 , w_11753 , w_11754 , w_11755 , w_11756 , w_11757 , w_11758 , w_11759 , 
		w_11760 , w_11761 , w_11762 , w_11763 , w_11764 , w_11765 , w_11766 , w_11767 , w_11768 , w_11769 , 
		w_11770 , w_11771 , w_11772 , w_11773 , w_11774 , w_11775 , w_11776 , w_11777 , w_11778 , w_11779 , 
		w_11780 , w_11781 , w_11782 , w_11783 , w_11784 , w_11785 , w_11786 , w_11787 , w_11788 , w_11789 , 
		w_11790 , w_11791 , w_11792 , w_11793 , w_11794 , w_11795 , w_11796 , w_11797 , w_11798 , w_11799 , 
		w_11800 , w_11801 , w_11802 , w_11803 , w_11804 , w_11805 , w_11806 , w_11807 , w_11808 , w_11809 , 
		w_11810 , w_11811 , w_11812 , w_11813 , w_11814 , w_11815 , w_11816 , w_11817 , w_11818 , w_11819 , 
		w_11820 , w_11821 , w_11822 , w_11823 , w_11824 , w_11825 , w_11826 , w_11827 , w_11828 , w_11829 , 
		w_11830 , w_11831 , w_11832 , w_11833 , w_11834 , w_11835 , w_11836 , w_11837 , w_11838 , w_11839 , 
		w_11840 , w_11841 , w_11842 , w_11843 , w_11844 , w_11845 , w_11846 , w_11847 , w_11848 , w_11849 , 
		w_11850 , w_11851 , w_11852 , w_11853 , w_11854 , w_11855 , w_11856 , w_11857 , w_11858 , w_11859 , 
		w_11860 , w_11861 , w_11862 , w_11863 , w_11864 , w_11865 , w_11866 , w_11867 , w_11868 , w_11869 , 
		w_11870 , w_11871 , w_11872 , w_11873 , w_11874 , w_11875 , w_11876 , w_11877 , w_11878 , w_11879 , 
		w_11880 , w_11881 , w_11882 , w_11883 , w_11884 , w_11885 , w_11886 , w_11887 , w_11888 , w_11889 , 
		w_11890 , w_11891 , w_11892 , w_11893 , w_11894 , w_11895 , w_11896 , w_11897 , w_11898 , w_11899 , 
		w_11900 , w_11901 , w_11902 , w_11903 , w_11904 , w_11905 , w_11906 , w_11907 , w_11908 , w_11909 , 
		w_11910 , w_11911 , w_11912 , w_11913 , w_11914 , w_11915 , w_11916 , w_11917 , w_11918 , w_11919 , 
		w_11920 , w_11921 , w_11922 , w_11923 , w_11924 , w_11925 , w_11926 , w_11927 , w_11928 , w_11929 , 
		w_11930 , w_11931 , w_11932 , w_11933 , w_11934 , w_11935 , w_11936 , w_11937 , w_11938 , w_11939 , 
		w_11940 , w_11941 , w_11942 , w_11943 , w_11944 , w_11945 , w_11946 , w_11947 , w_11948 , w_11949 , 
		w_11950 , w_11951 , w_11952 , w_11953 , w_11954 , w_11955 , w_11956 , w_11957 , w_11958 , w_11959 , 
		w_11960 , w_11961 , w_11962 , w_11963 , w_11964 , w_11965 , w_11966 , w_11967 , w_11968 , w_11969 , 
		w_11970 , w_11971 , w_11972 , w_11973 , w_11974 , w_11975 , w_11976 , w_11977 , w_11978 , w_11979 , 
		w_11980 , w_11981 , w_11982 , w_11983 , w_11984 , w_11985 , w_11986 , w_11987 , w_11988 , w_11989 , 
		w_11990 , w_11991 , w_11992 , w_11993 , w_11994 , w_11995 , w_11996 , w_11997 , w_11998 , w_11999 , 
		w_12000 , w_12001 , w_12002 , w_12003 , w_12004 , w_12005 , w_12006 , w_12007 , w_12008 , w_12009 , 
		w_12010 , w_12011 , w_12012 , w_12013 , w_12014 , w_12015 , w_12016 , w_12017 , w_12018 , w_12019 , 
		w_12020 , w_12021 , w_12022 , w_12023 , w_12024 , w_12025 , w_12026 , w_12027 , w_12028 , w_12029 , 
		w_12030 , w_12031 , w_12032 , w_12033 , w_12034 , w_12035 , w_12036 , w_12037 , w_12038 , w_12039 , 
		w_12040 , w_12041 , w_12042 , w_12043 , w_12044 , w_12045 , w_12046 , w_12047 , w_12048 , w_12049 , 
		w_12050 , w_12051 , w_12052 , w_12053 , w_12054 , w_12055 , w_12056 , w_12057 , w_12058 , w_12059 , 
		w_12060 , w_12061 , w_12062 , w_12063 , w_12064 , w_12065 , w_12066 , w_12067 , w_12068 , w_12069 , 
		w_12070 , w_12071 , w_12072 , w_12073 , w_12074 , w_12075 , w_12076 , w_12077 , w_12078 , w_12079 , 
		w_12080 , w_12081 , w_12082 , w_12083 , w_12084 , w_12085 , w_12086 , w_12087 , w_12088 , w_12089 , 
		w_12090 , w_12091 , w_12092 , w_12093 , w_12094 , w_12095 , w_12096 , w_12097 , w_12098 , w_12099 , 
		w_12100 , w_12101 , w_12102 , w_12103 , w_12104 , w_12105 , w_12106 , w_12107 , w_12108 , w_12109 , 
		w_12110 , w_12111 , w_12112 , w_12113 , w_12114 , w_12115 , w_12116 , w_12117 , w_12118 , w_12119 , 
		w_12120 , w_12121 , w_12122 , w_12123 , w_12124 , w_12125 , w_12126 , w_12127 , w_12128 , w_12129 , 
		w_12130 , w_12131 , w_12132 , w_12133 , w_12134 , w_12135 , w_12136 , w_12137 , w_12138 , w_12139 , 
		w_12140 , w_12141 , w_12142 , w_12143 , w_12144 , w_12145 , w_12146 , w_12147 , w_12148 , w_12149 , 
		w_12150 , w_12151 , w_12152 , w_12153 , w_12154 , w_12155 , w_12156 , w_12157 , w_12158 , w_12159 , 
		w_12160 , w_12161 , w_12162 , w_12163 , w_12164 , w_12165 , w_12166 , w_12167 , w_12168 , w_12169 , 
		w_12170 , w_12171 , w_12172 , w_12173 , w_12174 , w_12175 , w_12176 , w_12177 , w_12178 , w_12179 , 
		w_12180 , w_12181 , w_12182 , w_12183 , w_12184 , w_12185 , w_12186 , w_12187 , w_12188 , w_12189 , 
		w_12190 , w_12191 , w_12192 , w_12193 , w_12194 , w_12195 , w_12196 , w_12197 , w_12198 , w_12199 , 
		w_12200 , w_12201 , w_12202 , w_12203 , w_12204 , w_12205 , w_12206 , w_12207 , w_12208 , w_12209 , 
		w_12210 , w_12211 , w_12212 , w_12213 , w_12214 , w_12215 , w_12216 , w_12217 , w_12218 , w_12219 , 
		w_12220 , w_12221 , w_12222 , w_12223 , w_12224 , w_12225 , w_12226 , w_12227 , w_12228 , w_12229 , 
		w_12230 , w_12231 , w_12232 , w_12233 , w_12234 , w_12235 , w_12236 , w_12237 , w_12238 , w_12239 , 
		w_12240 , w_12241 , w_12242 , w_12243 , w_12244 , w_12245 , w_12246 , w_12247 , w_12248 , w_12249 , 
		w_12250 , w_12251 , w_12252 , w_12253 , w_12254 , w_12255 , w_12256 , w_12257 , w_12258 , w_12259 , 
		w_12260 , w_12261 , w_12262 , w_12263 , w_12264 , w_12265 , w_12266 , w_12267 , w_12268 , w_12269 , 
		w_12270 , w_12271 , w_12272 , w_12273 , w_12274 , w_12275 , w_12276 , w_12277 , w_12278 , w_12279 , 
		w_12280 , w_12281 , w_12282 , w_12283 , w_12284 , w_12285 , w_12286 , w_12287 , w_12288 , w_12289 , 
		w_12290 , w_12291 , w_12292 , w_12293 , w_12294 , w_12295 , w_12296 , w_12297 , w_12298 , w_12299 , 
		w_12300 , w_12301 , w_12302 , w_12303 , w_12304 , w_12305 , w_12306 , w_12307 , w_12308 , w_12309 , 
		w_12310 , w_12311 , w_12312 , w_12313 , w_12314 , w_12315 , w_12316 , w_12317 , w_12318 , w_12319 , 
		w_12320 , w_12321 , w_12322 , w_12323 , w_12324 , w_12325 , w_12326 , w_12327 , w_12328 , w_12329 , 
		w_12330 , w_12331 , w_12332 , w_12333 , w_12334 , w_12335 , w_12336 , w_12337 , w_12338 , w_12339 , 
		w_12340 , w_12341 , w_12342 , w_12343 , w_12344 , w_12345 , w_12346 , w_12347 , w_12348 , w_12349 , 
		w_12350 , w_12351 , w_12352 , w_12353 , w_12354 , w_12355 , w_12356 , w_12357 , w_12358 , w_12359 , 
		w_12360 , w_12361 , w_12362 , w_12363 , w_12364 , w_12365 , w_12366 , w_12367 , w_12368 , w_12369 , 
		w_12370 , w_12371 , w_12372 , w_12373 , w_12374 , w_12375 , w_12376 , w_12377 , w_12378 , w_12379 , 
		w_12380 , w_12381 , w_12382 , w_12383 , w_12384 , w_12385 , w_12386 , w_12387 , w_12388 , w_12389 , 
		w_12390 , w_12391 , w_12392 , w_12393 , w_12394 , w_12395 , w_12396 , w_12397 , w_12398 , w_12399 , 
		w_12400 , w_12401 , w_12402 , w_12403 , w_12404 , w_12405 , w_12406 , w_12407 , w_12408 , w_12409 , 
		w_12410 , w_12411 , w_12412 , w_12413 , w_12414 , w_12415 , w_12416 , w_12417 , w_12418 , w_12419 , 
		w_12420 , w_12421 , w_12422 , w_12423 , w_12424 , w_12425 , w_12426 , w_12427 , w_12428 , w_12429 , 
		w_12430 , w_12431 , w_12432 , w_12433 , w_12434 , w_12435 , w_12436 , w_12437 , w_12438 , w_12439 , 
		w_12440 , w_12441 , w_12442 , w_12443 , w_12444 , w_12445 , w_12446 , w_12447 , w_12448 , w_12449 , 
		w_12450 , w_12451 , w_12452 , w_12453 , w_12454 , w_12455 , w_12456 , w_12457 , w_12458 , w_12459 , 
		w_12460 , w_12461 , w_12462 , w_12463 , w_12464 , w_12465 , w_12466 , w_12467 , w_12468 , w_12469 , 
		w_12470 , w_12471 , w_12472 , w_12473 , w_12474 , w_12475 , w_12476 , w_12477 , w_12478 , w_12479 , 
		w_12480 , w_12481 , w_12482 , w_12483 , w_12484 , w_12485 , w_12486 , w_12487 , w_12488 , w_12489 , 
		w_12490 , w_12491 , w_12492 , w_12493 , w_12494 , w_12495 , w_12496 , w_12497 , w_12498 , w_12499 , 
		w_12500 , w_12501 , w_12502 , w_12503 , w_12504 , w_12505 , w_12506 , w_12507 , w_12508 , w_12509 , 
		w_12510 , w_12511 , w_12512 , w_12513 , w_12514 , w_12515 , w_12516 , w_12517 , w_12518 , w_12519 , 
		w_12520 , w_12521 , w_12522 , w_12523 , w_12524 , w_12525 , w_12526 , w_12527 , w_12528 , w_12529 , 
		w_12530 , w_12531 , w_12532 , w_12533 , w_12534 , w_12535 , w_12536 , w_12537 , w_12538 , w_12539 , 
		w_12540 , w_12541 , w_12542 , w_12543 , w_12544 , w_12545 , w_12546 , w_12547 , w_12548 , w_12549 , 
		w_12550 , w_12551 , w_12552 , w_12553 , w_12554 , w_12555 , w_12556 , w_12557 , w_12558 , w_12559 , 
		w_12560 , w_12561 , w_12562 , w_12563 , w_12564 , w_12565 , w_12566 , w_12567 , w_12568 , w_12569 , 
		w_12570 , w_12571 , w_12572 , w_12573 , w_12574 , w_12575 , w_12576 , w_12577 , w_12578 , w_12579 , 
		w_12580 , w_12581 , w_12582 , w_12583 , w_12584 , w_12585 , w_12586 , w_12587 , w_12588 , w_12589 , 
		w_12590 , w_12591 , w_12592 , w_12593 , w_12594 , w_12595 , w_12596 , w_12597 , w_12598 , w_12599 , 
		w_12600 , w_12601 , w_12602 , w_12603 , w_12604 , w_12605 , w_12606 , w_12607 , w_12608 , w_12609 , 
		w_12610 , w_12611 , w_12612 , w_12613 , w_12614 , w_12615 , w_12616 , w_12617 , w_12618 , w_12619 , 
		w_12620 , w_12621 , w_12622 , w_12623 , w_12624 , w_12625 , w_12626 , w_12627 , w_12628 , w_12629 , 
		w_12630 , w_12631 , w_12632 , w_12633 , w_12634 , w_12635 , w_12636 , w_12637 , w_12638 , w_12639 , 
		w_12640 , w_12641 , w_12642 , w_12643 , w_12644 , w_12645 , w_12646 , w_12647 , w_12648 , w_12649 , 
		w_12650 , w_12651 , w_12652 , w_12653 , w_12654 , w_12655 , w_12656 , w_12657 , w_12658 , w_12659 , 
		w_12660 , w_12661 , w_12662 , w_12663 , w_12664 , w_12665 , w_12666 , w_12667 , w_12668 , w_12669 , 
		w_12670 , w_12671 , w_12672 , w_12673 , w_12674 , w_12675 , w_12676 , w_12677 , w_12678 , w_12679 , 
		w_12680 , w_12681 , w_12682 , w_12683 , w_12684 , w_12685 , w_12686 , w_12687 , w_12688 , w_12689 , 
		w_12690 , w_12691 , w_12692 , w_12693 , w_12694 , w_12695 , w_12696 , w_12697 , w_12698 , w_12699 , 
		w_12700 , w_12701 , w_12702 , w_12703 , w_12704 , w_12705 , w_12706 , w_12707 , w_12708 , w_12709 , 
		w_12710 , w_12711 , w_12712 , w_12713 , w_12714 , w_12715 , w_12716 , w_12717 , w_12718 , w_12719 , 
		w_12720 , w_12721 , w_12722 , w_12723 , w_12724 , w_12725 , w_12726 , w_12727 , w_12728 , w_12729 , 
		w_12730 , w_12731 , w_12732 , w_12733 , w_12734 , w_12735 , w_12736 , w_12737 , w_12738 , w_12739 , 
		w_12740 , w_12741 , w_12742 , w_12743 , w_12744 , w_12745 , w_12746 , w_12747 , w_12748 , w_12749 , 
		w_12750 , w_12751 , w_12752 , w_12753 , w_12754 , w_12755 , w_12756 , w_12757 , w_12758 , w_12759 , 
		w_12760 , w_12761 , w_12762 , w_12763 , w_12764 , w_12765 , w_12766 , w_12767 , w_12768 , w_12769 , 
		w_12770 , w_12771 , w_12772 , w_12773 , w_12774 , w_12775 , w_12776 , w_12777 , w_12778 , w_12779 , 
		w_12780 , w_12781 , w_12782 , w_12783 , w_12784 , w_12785 , w_12786 , w_12787 , w_12788 , w_12789 , 
		w_12790 , w_12791 , w_12792 , w_12793 , w_12794 , w_12795 , w_12796 , w_12797 , w_12798 , w_12799 , 
		w_12800 , w_12801 , w_12802 , w_12803 , w_12804 , w_12805 , w_12806 , w_12807 , w_12808 , w_12809 , 
		w_12810 , w_12811 , w_12812 , w_12813 , w_12814 , w_12815 , w_12816 , w_12817 , w_12818 , w_12819 , 
		w_12820 , w_12821 , w_12822 , w_12823 , w_12824 , w_12825 , w_12826 , w_12827 , w_12828 , w_12829 , 
		w_12830 , w_12831 , w_12832 , w_12833 , w_12834 , w_12835 , w_12836 , w_12837 , w_12838 , w_12839 , 
		w_12840 , w_12841 , w_12842 , w_12843 , w_12844 , w_12845 , w_12846 , w_12847 , w_12848 , w_12849 , 
		w_12850 , w_12851 , w_12852 , w_12853 , w_12854 , w_12855 , w_12856 , w_12857 , w_12858 , w_12859 , 
		w_12860 , w_12861 , w_12862 , w_12863 , w_12864 , w_12865 , w_12866 , w_12867 , w_12868 , w_12869 , 
		w_12870 , w_12871 , w_12872 , w_12873 , w_12874 , w_12875 , w_12876 , w_12877 , w_12878 , w_12879 , 
		w_12880 , w_12881 , w_12882 , w_12883 , w_12884 , w_12885 , w_12886 , w_12887 , w_12888 , w_12889 , 
		w_12890 , w_12891 , w_12892 , w_12893 , w_12894 , w_12895 , w_12896 , w_12897 , w_12898 , w_12899 , 
		w_12900 , w_12901 , w_12902 , w_12903 , w_12904 , w_12905 , w_12906 , w_12907 , w_12908 , w_12909 , 
		w_12910 , w_12911 , w_12912 , w_12913 , w_12914 , w_12915 , w_12916 , w_12917 , w_12918 , w_12919 , 
		w_12920 , w_12921 , w_12922 , w_12923 , w_12924 , w_12925 , w_12926 , w_12927 , w_12928 , w_12929 , 
		w_12930 , w_12931 , w_12932 , w_12933 , w_12934 , w_12935 , w_12936 , w_12937 , w_12938 , w_12939 , 
		w_12940 , w_12941 , w_12942 , w_12943 , w_12944 , w_12945 , w_12946 , w_12947 , w_12948 , w_12949 , 
		w_12950 , w_12951 , w_12952 , w_12953 , w_12954 , w_12955 , w_12956 , w_12957 , w_12958 , w_12959 , 
		w_12960 , w_12961 , w_12962 , w_12963 , w_12964 , w_12965 , w_12966 , w_12967 , w_12968 , w_12969 , 
		w_12970 , w_12971 , w_12972 , w_12973 , w_12974 , w_12975 , w_12976 , w_12977 , w_12978 , w_12979 , 
		w_12980 , w_12981 , w_12982 , w_12983 , w_12984 , w_12985 , w_12986 , w_12987 , w_12988 , w_12989 , 
		w_12990 , w_12991 , w_12992 , w_12993 , w_12994 , w_12995 , w_12996 , w_12997 , w_12998 , w_12999 , 
		w_13000 , w_13001 , w_13002 , w_13003 , w_13004 , w_13005 , w_13006 , w_13007 , w_13008 , w_13009 , 
		w_13010 , w_13011 , w_13012 , w_13013 , w_13014 , w_13015 , w_13016 , w_13017 , w_13018 , w_13019 , 
		w_13020 , w_13021 , w_13022 , w_13023 , w_13024 , w_13025 , w_13026 , w_13027 , w_13028 , w_13029 , 
		w_13030 , w_13031 , w_13032 , w_13033 , w_13034 , w_13035 , w_13036 , w_13037 , w_13038 , w_13039 , 
		w_13040 , w_13041 , w_13042 , w_13043 , w_13044 , w_13045 , w_13046 , w_13047 , w_13048 , w_13049 , 
		w_13050 , w_13051 , w_13052 , w_13053 , w_13054 , w_13055 , w_13056 , w_13057 , w_13058 , w_13059 , 
		w_13060 , w_13061 , w_13062 , w_13063 , w_13064 , w_13065 , w_13066 , w_13067 , w_13068 , w_13069 , 
		w_13070 , w_13071 , w_13072 , w_13073 , w_13074 , w_13075 , w_13076 , w_13077 , w_13078 , w_13079 , 
		w_13080 , w_13081 , w_13082 , w_13083 , w_13084 , w_13085 , w_13086 , w_13087 , w_13088 , w_13089 , 
		w_13090 , w_13091 , w_13092 , w_13093 , w_13094 , w_13095 , w_13096 , w_13097 , w_13098 , w_13099 , 
		w_13100 , w_13101 , w_13102 , w_13103 , w_13104 , w_13105 , w_13106 , w_13107 , w_13108 , w_13109 , 
		w_13110 , w_13111 , w_13112 , w_13113 , w_13114 , w_13115 , w_13116 , w_13117 , w_13118 , w_13119 , 
		w_13120 , w_13121 , w_13122 , w_13123 , w_13124 , w_13125 , w_13126 , w_13127 , w_13128 , w_13129 , 
		w_13130 , w_13131 , w_13132 , w_13133 , w_13134 , w_13135 , w_13136 , w_13137 , w_13138 , w_13139 , 
		w_13140 , w_13141 , w_13142 , w_13143 , w_13144 , w_13145 , w_13146 , w_13147 , w_13148 , w_13149 , 
		w_13150 , w_13151 , w_13152 , w_13153 , w_13154 , w_13155 , w_13156 , w_13157 , w_13158 , w_13159 , 
		w_13160 , w_13161 , w_13162 , w_13163 , w_13164 , w_13165 , w_13166 , w_13167 , w_13168 , w_13169 , 
		w_13170 , w_13171 , w_13172 , w_13173 , w_13174 , w_13175 , w_13176 , w_13177 , w_13178 , w_13179 , 
		w_13180 , w_13181 , w_13182 , w_13183 , w_13184 , w_13185 , w_13186 , w_13187 , w_13188 , w_13189 , 
		w_13190 , w_13191 , w_13192 , w_13193 , w_13194 , w_13195 , w_13196 , w_13197 , w_13198 , w_13199 , 
		w_13200 , w_13201 , w_13202 , w_13203 , w_13204 , w_13205 , w_13206 , w_13207 , w_13208 , w_13209 , 
		w_13210 , w_13211 , w_13212 , w_13213 , w_13214 , w_13215 , w_13216 , w_13217 , w_13218 , w_13219 , 
		w_13220 , w_13221 , w_13222 , w_13223 , w_13224 , w_13225 , w_13226 , w_13227 , w_13228 , w_13229 , 
		w_13230 , w_13231 , w_13232 , w_13233 , w_13234 , w_13235 , w_13236 , w_13237 , w_13238 , w_13239 , 
		w_13240 , w_13241 , w_13242 , w_13243 , w_13244 , w_13245 , w_13246 , w_13247 , w_13248 , w_13249 , 
		w_13250 , w_13251 , w_13252 , w_13253 , w_13254 , w_13255 , w_13256 , w_13257 , w_13258 , w_13259 , 
		w_13260 , w_13261 , w_13262 , w_13263 , w_13264 , w_13265 , w_13266 , w_13267 , w_13268 , w_13269 , 
		w_13270 , w_13271 , w_13272 , w_13273 , w_13274 , w_13275 , w_13276 , w_13277 , w_13278 , w_13279 , 
		w_13280 , w_13281 , w_13282 , w_13283 , w_13284 , w_13285 , w_13286 , w_13287 , w_13288 , w_13289 , 
		w_13290 , w_13291 , w_13292 , w_13293 , w_13294 , w_13295 , w_13296 , w_13297 , w_13298 , w_13299 , 
		w_13300 , w_13301 , w_13302 , w_13303 , w_13304 , w_13305 , w_13306 , w_13307 , w_13308 , w_13309 , 
		w_13310 , w_13311 , w_13312 , w_13313 , w_13314 , w_13315 , w_13316 , w_13317 , w_13318 , w_13319 , 
		w_13320 , w_13321 , w_13322 , w_13323 , w_13324 , w_13325 , w_13326 , w_13327 , w_13328 , w_13329 , 
		w_13330 , w_13331 , w_13332 , w_13333 , w_13334 , w_13335 , w_13336 , w_13337 , w_13338 , w_13339 , 
		w_13340 , w_13341 , w_13342 , w_13343 , w_13344 , w_13345 , w_13346 , w_13347 , w_13348 , w_13349 , 
		w_13350 , w_13351 , w_13352 , w_13353 , w_13354 , w_13355 , w_13356 , w_13357 , w_13358 , w_13359 , 
		w_13360 , w_13361 , w_13362 , w_13363 , w_13364 , w_13365 , w_13366 , w_13367 , w_13368 , w_13369 , 
		w_13370 , w_13371 , w_13372 , w_13373 , w_13374 , w_13375 , w_13376 , w_13377 , w_13378 , w_13379 , 
		w_13380 , w_13381 , w_13382 , w_13383 , w_13384 , w_13385 , w_13386 , w_13387 , w_13388 , w_13389 , 
		w_13390 , w_13391 , w_13392 , w_13393 , w_13394 , w_13395 , w_13396 , w_13397 , w_13398 , w_13399 , 
		w_13400 , w_13401 , w_13402 , w_13403 , w_13404 , w_13405 , w_13406 , w_13407 , w_13408 , w_13409 , 
		w_13410 , w_13411 , w_13412 , w_13413 , w_13414 , w_13415 , w_13416 , w_13417 , w_13418 , w_13419 , 
		w_13420 , w_13421 , w_13422 , w_13423 , w_13424 , w_13425 , w_13426 , w_13427 , w_13428 , w_13429 , 
		w_13430 , w_13431 , w_13432 , w_13433 , w_13434 , w_13435 , w_13436 , w_13437 , w_13438 , w_13439 , 
		w_13440 , w_13441 , w_13442 , w_13443 , w_13444 , w_13445 , w_13446 , w_13447 , w_13448 , w_13449 , 
		w_13450 , w_13451 , w_13452 , w_13453 , w_13454 , w_13455 , w_13456 , w_13457 , w_13458 , w_13459 , 
		w_13460 , w_13461 , w_13462 , w_13463 , w_13464 , w_13465 , w_13466 , w_13467 , w_13468 , w_13469 , 
		w_13470 , w_13471 , w_13472 , w_13473 , w_13474 , w_13475 , w_13476 , w_13477 , w_13478 , w_13479 , 
		w_13480 , w_13481 , w_13482 , w_13483 , w_13484 , w_13485 , w_13486 , w_13487 , w_13488 , w_13489 , 
		w_13490 , w_13491 , w_13492 , w_13493 , w_13494 , w_13495 , w_13496 , w_13497 , w_13498 , w_13499 , 
		w_13500 , w_13501 , w_13502 , w_13503 , w_13504 , w_13505 , w_13506 , w_13507 , w_13508 , w_13509 , 
		w_13510 , w_13511 , w_13512 , w_13513 , w_13514 , w_13515 , w_13516 , w_13517 , w_13518 , w_13519 , 
		w_13520 , w_13521 , w_13522 , w_13523 , w_13524 , w_13525 , w_13526 , w_13527 , w_13528 , w_13529 , 
		w_13530 , w_13531 , w_13532 , w_13533 , w_13534 , w_13535 , w_13536 , w_13537 , w_13538 , w_13539 , 
		w_13540 , w_13541 , w_13542 , w_13543 , w_13544 , w_13545 , w_13546 , w_13547 , w_13548 , w_13549 , 
		w_13550 , w_13551 , w_13552 , w_13553 , w_13554 , w_13555 , w_13556 , w_13557 , w_13558 , w_13559 , 
		w_13560 , w_13561 , w_13562 , w_13563 , w_13564 , w_13565 , w_13566 , w_13567 , w_13568 , w_13569 , 
		w_13570 , w_13571 , w_13572 , w_13573 , w_13574 , w_13575 , w_13576 , w_13577 , w_13578 , w_13579 , 
		w_13580 , w_13581 , w_13582 , w_13583 , w_13584 , w_13585 , w_13586 , w_13587 , w_13588 , w_13589 , 
		w_13590 , w_13591 , w_13592 , w_13593 , w_13594 , w_13595 , w_13596 , w_13597 , w_13598 , w_13599 , 
		w_13600 , w_13601 , w_13602 , w_13603 , w_13604 , w_13605 , w_13606 , w_13607 , w_13608 , w_13609 , 
		w_13610 , w_13611 , w_13612 , w_13613 , w_13614 , w_13615 , w_13616 , w_13617 , w_13618 , w_13619 , 
		w_13620 , w_13621 , w_13622 , w_13623 , w_13624 , w_13625 , w_13626 , w_13627 , w_13628 , w_13629 , 
		w_13630 , w_13631 , w_13632 , w_13633 , w_13634 , w_13635 , w_13636 , w_13637 , w_13638 , w_13639 , 
		w_13640 , w_13641 , w_13642 , w_13643 , w_13644 , w_13645 , w_13646 , w_13647 , w_13648 , w_13649 , 
		w_13650 , w_13651 , w_13652 , w_13653 , w_13654 , w_13655 , w_13656 , w_13657 , w_13658 , w_13659 , 
		w_13660 , w_13661 , w_13662 , w_13663 , w_13664 , w_13665 , w_13666 , w_13667 , w_13668 , w_13669 , 
		w_13670 , w_13671 , w_13672 , w_13673 , w_13674 , w_13675 , w_13676 , w_13677 , w_13678 , w_13679 , 
		w_13680 , w_13681 , w_13682 , w_13683 , w_13684 , w_13685 , w_13686 , w_13687 , w_13688 , w_13689 , 
		w_13690 , w_13691 , w_13692 , w_13693 , w_13694 , w_13695 , w_13696 , w_13697 , w_13698 , w_13699 , 
		w_13700 , w_13701 , w_13702 , w_13703 , w_13704 , w_13705 , w_13706 , w_13707 , w_13708 , w_13709 , 
		w_13710 , w_13711 , w_13712 , w_13713 , w_13714 , w_13715 , w_13716 , w_13717 , w_13718 , w_13719 , 
		w_13720 , w_13721 , w_13722 , w_13723 , w_13724 , w_13725 , w_13726 , w_13727 , w_13728 , w_13729 , 
		w_13730 , w_13731 , w_13732 , w_13733 , w_13734 , w_13735 , w_13736 , w_13737 , w_13738 , w_13739 , 
		w_13740 , w_13741 , w_13742 , w_13743 , w_13744 , w_13745 , w_13746 , w_13747 , w_13748 , w_13749 , 
		w_13750 , w_13751 , w_13752 , w_13753 , w_13754 , w_13755 , w_13756 , w_13757 , w_13758 , w_13759 , 
		w_13760 , w_13761 , w_13762 , w_13763 , w_13764 , w_13765 , w_13766 , w_13767 , w_13768 , w_13769 , 
		w_13770 , w_13771 , w_13772 , w_13773 , w_13774 , w_13775 , w_13776 , w_13777 , w_13778 , w_13779 , 
		w_13780 , w_13781 , w_13782 , w_13783 , w_13784 , w_13785 , w_13786 , w_13787 , w_13788 , w_13789 , 
		w_13790 , w_13791 , w_13792 , w_13793 , w_13794 , w_13795 , w_13796 , w_13797 , w_13798 , w_13799 , 
		w_13800 , w_13801 , w_13802 , w_13803 , w_13804 , w_13805 , w_13806 , w_13807 , w_13808 , w_13809 , 
		w_13810 , w_13811 , w_13812 , w_13813 , w_13814 , w_13815 , w_13816 , w_13817 , w_13818 , w_13819 , 
		w_13820 , w_13821 , w_13822 , w_13823 , w_13824 , w_13825 , w_13826 , w_13827 , w_13828 , w_13829 , 
		w_13830 , w_13831 , w_13832 , w_13833 , w_13834 , w_13835 , w_13836 , w_13837 , w_13838 , w_13839 , 
		w_13840 , w_13841 , w_13842 , w_13843 , w_13844 , w_13845 , w_13846 , w_13847 , w_13848 , w_13849 , 
		w_13850 , w_13851 , w_13852 , w_13853 , w_13854 , w_13855 , w_13856 , w_13857 , w_13858 , w_13859 , 
		w_13860 , w_13861 , w_13862 , w_13863 , w_13864 , w_13865 , w_13866 , w_13867 , w_13868 , w_13869 , 
		w_13870 , w_13871 , w_13872 , w_13873 , w_13874 , w_13875 , w_13876 , w_13877 , w_13878 , w_13879 , 
		w_13880 , w_13881 , w_13882 , w_13883 , w_13884 , w_13885 , w_13886 , w_13887 , w_13888 , w_13889 , 
		w_13890 , w_13891 , w_13892 , w_13893 , w_13894 , w_13895 , w_13896 , w_13897 , w_13898 , w_13899 , 
		w_13900 , w_13901 , w_13902 , w_13903 , w_13904 , w_13905 , w_13906 , w_13907 , w_13908 , w_13909 , 
		w_13910 , w_13911 , w_13912 , w_13913 , w_13914 , w_13915 , w_13916 , w_13917 , w_13918 , w_13919 , 
		w_13920 , w_13921 , w_13922 , w_13923 , w_13924 , w_13925 , w_13926 , w_13927 , w_13928 , w_13929 , 
		w_13930 , w_13931 , w_13932 , w_13933 , w_13934 , w_13935 , w_13936 , w_13937 , w_13938 , w_13939 , 
		w_13940 , w_13941 , w_13942 , w_13943 , w_13944 , w_13945 , w_13946 , w_13947 , w_13948 , w_13949 , 
		w_13950 , w_13951 , w_13952 , w_13953 , w_13954 , w_13955 , w_13956 , w_13957 , w_13958 , w_13959 , 
		w_13960 , w_13961 , w_13962 , w_13963 , w_13964 , w_13965 , w_13966 , w_13967 , w_13968 , w_13969 , 
		w_13970 , w_13971 , w_13972 , w_13973 , w_13974 , w_13975 , w_13976 , w_13977 , w_13978 , w_13979 , 
		w_13980 , w_13981 , w_13982 , w_13983 , w_13984 , w_13985 , w_13986 , w_13987 , w_13988 , w_13989 , 
		w_13990 , w_13991 , w_13992 , w_13993 , w_13994 , w_13995 , w_13996 , w_13997 , w_13998 , w_13999 , 
		w_14000 , w_14001 , w_14002 , w_14003 , w_14004 , w_14005 , w_14006 , w_14007 , w_14008 , w_14009 , 
		w_14010 , w_14011 , w_14012 , w_14013 , w_14014 , w_14015 , w_14016 , w_14017 , w_14018 , w_14019 , 
		w_14020 , w_14021 , w_14022 , w_14023 , w_14024 , w_14025 , w_14026 , w_14027 , w_14028 , w_14029 , 
		w_14030 , w_14031 , w_14032 , w_14033 , w_14034 , w_14035 , w_14036 , w_14037 , w_14038 , w_14039 , 
		w_14040 , w_14041 , w_14042 , w_14043 , w_14044 , w_14045 , w_14046 , w_14047 , w_14048 , w_14049 , 
		w_14050 , w_14051 , w_14052 , w_14053 , w_14054 , w_14055 , w_14056 , w_14057 , w_14058 , w_14059 , 
		w_14060 , w_14061 , w_14062 , w_14063 , w_14064 , w_14065 , w_14066 , w_14067 , w_14068 , w_14069 , 
		w_14070 , w_14071 , w_14072 , w_14073 , w_14074 , w_14075 , w_14076 , w_14077 , w_14078 , w_14079 , 
		w_14080 , w_14081 , w_14082 , w_14083 , w_14084 , w_14085 , w_14086 , w_14087 , w_14088 , w_14089 , 
		w_14090 , w_14091 , w_14092 , w_14093 , w_14094 , w_14095 , w_14096 , w_14097 , w_14098 , w_14099 , 
		w_14100 , w_14101 , w_14102 , w_14103 , w_14104 , w_14105 , w_14106 , w_14107 , w_14108 , w_14109 , 
		w_14110 , w_14111 , w_14112 , w_14113 , w_14114 , w_14115 , w_14116 , w_14117 , w_14118 , w_14119 , 
		w_14120 , w_14121 , w_14122 , w_14123 , w_14124 , w_14125 , w_14126 , w_14127 , w_14128 , w_14129 , 
		w_14130 , w_14131 , w_14132 , w_14133 , w_14134 , w_14135 , w_14136 , w_14137 , w_14138 , w_14139 , 
		w_14140 , w_14141 , w_14142 , w_14143 , w_14144 , w_14145 , w_14146 , w_14147 , w_14148 , w_14149 , 
		w_14150 , w_14151 , w_14152 , w_14153 , w_14154 , w_14155 , w_14156 , w_14157 , w_14158 , w_14159 , 
		w_14160 , w_14161 , w_14162 , w_14163 , w_14164 , w_14165 , w_14166 , w_14167 , w_14168 , w_14169 , 
		w_14170 , w_14171 , w_14172 , w_14173 , w_14174 , w_14175 , w_14176 , w_14177 , w_14178 , w_14179 , 
		w_14180 , w_14181 , w_14182 , w_14183 , w_14184 , w_14185 , w_14186 , w_14187 , w_14188 , w_14189 , 
		w_14190 , w_14191 , w_14192 , w_14193 , w_14194 , w_14195 , w_14196 , w_14197 , w_14198 , w_14199 , 
		w_14200 , w_14201 , w_14202 , w_14203 , w_14204 , w_14205 , w_14206 , w_14207 , w_14208 , w_14209 , 
		w_14210 , w_14211 , w_14212 , w_14213 , w_14214 , w_14215 , w_14216 , w_14217 , w_14218 , w_14219 , 
		w_14220 , w_14221 , w_14222 , w_14223 , w_14224 , w_14225 , w_14226 , w_14227 , w_14228 , w_14229 , 
		w_14230 , w_14231 , w_14232 , w_14233 , w_14234 , w_14235 , w_14236 , w_14237 , w_14238 , w_14239 , 
		w_14240 , w_14241 , w_14242 , w_14243 , w_14244 , w_14245 , w_14246 , w_14247 , w_14248 , w_14249 , 
		w_14250 , w_14251 , w_14252 , w_14253 , w_14254 , w_14255 , w_14256 , w_14257 , w_14258 , w_14259 , 
		w_14260 , w_14261 , w_14262 , w_14263 , w_14264 , w_14265 , w_14266 , w_14267 , w_14268 , w_14269 , 
		w_14270 , w_14271 , w_14272 , w_14273 , w_14274 , w_14275 , w_14276 , w_14277 , w_14278 , w_14279 , 
		w_14280 , w_14281 , w_14282 , w_14283 , w_14284 , w_14285 , w_14286 , w_14287 , w_14288 , w_14289 , 
		w_14290 , w_14291 , w_14292 , w_14293 , w_14294 , w_14295 , w_14296 , w_14297 , w_14298 , w_14299 , 
		w_14300 , w_14301 , w_14302 , w_14303 , w_14304 , w_14305 , w_14306 , w_14307 , w_14308 , w_14309 , 
		w_14310 , w_14311 , w_14312 , w_14313 , w_14314 , w_14315 , w_14316 , w_14317 , w_14318 , w_14319 , 
		w_14320 , w_14321 , w_14322 , w_14323 , w_14324 , w_14325 , w_14326 , w_14327 , w_14328 , w_14329 , 
		w_14330 , w_14331 , w_14332 , w_14333 , w_14334 , w_14335 , w_14336 , w_14337 , w_14338 , w_14339 , 
		w_14340 , w_14341 , w_14342 , w_14343 , w_14344 , w_14345 , w_14346 , w_14347 , w_14348 , w_14349 , 
		w_14350 , w_14351 , w_14352 , w_14353 , w_14354 , w_14355 , w_14356 , w_14357 , w_14358 , w_14359 , 
		w_14360 , w_14361 , w_14362 , w_14363 , w_14364 , w_14365 , w_14366 , w_14367 , w_14368 , w_14369 , 
		w_14370 , w_14371 , w_14372 , w_14373 , w_14374 , w_14375 , w_14376 , w_14377 , w_14378 , w_14379 , 
		w_14380 , w_14381 , w_14382 , w_14383 , w_14384 , w_14385 , w_14386 , w_14387 , w_14388 , w_14389 , 
		w_14390 , w_14391 , w_14392 , w_14393 , w_14394 , w_14395 , w_14396 , w_14397 , w_14398 , w_14399 , 
		w_14400 , w_14401 , w_14402 , w_14403 , w_14404 , w_14405 , w_14406 , w_14407 , w_14408 , w_14409 , 
		w_14410 , w_14411 , w_14412 , w_14413 , w_14414 , w_14415 , w_14416 , w_14417 , w_14418 , w_14419 , 
		w_14420 , w_14421 , w_14422 , w_14423 , w_14424 , w_14425 , w_14426 , w_14427 , w_14428 , w_14429 , 
		w_14430 , w_14431 , w_14432 , w_14433 , w_14434 , w_14435 , w_14436 , w_14437 , w_14438 , w_14439 , 
		w_14440 , w_14441 , w_14442 , w_14443 , w_14444 , w_14445 , w_14446 , w_14447 , w_14448 , w_14449 , 
		w_14450 , w_14451 , w_14452 , w_14453 , w_14454 , w_14455 , w_14456 , w_14457 , w_14458 , w_14459 , 
		w_14460 , w_14461 , w_14462 , w_14463 , w_14464 , w_14465 , w_14466 , w_14467 , w_14468 , w_14469 , 
		w_14470 , w_14471 , w_14472 , w_14473 , w_14474 , w_14475 , w_14476 , w_14477 , w_14478 , w_14479 , 
		w_14480 , w_14481 , w_14482 , w_14483 , w_14484 , w_14485 , w_14486 , w_14487 , w_14488 , w_14489 , 
		w_14490 , w_14491 , w_14492 , w_14493 , w_14494 , w_14495 , w_14496 , w_14497 , w_14498 , w_14499 , 
		w_14500 , w_14501 , w_14502 , w_14503 , w_14504 , w_14505 , w_14506 , w_14507 , w_14508 , w_14509 , 
		w_14510 , w_14511 , w_14512 , w_14513 , w_14514 , w_14515 , w_14516 , w_14517 , w_14518 , w_14519 , 
		w_14520 , w_14521 , w_14522 , w_14523 , w_14524 , w_14525 , w_14526 , w_14527 , w_14528 , w_14529 , 
		w_14530 , w_14531 , w_14532 , w_14533 , w_14534 , w_14535 , w_14536 , w_14537 , w_14538 , w_14539 , 
		w_14540 , w_14541 , w_14542 , w_14543 , w_14544 , w_14545 , w_14546 , w_14547 , w_14548 , w_14549 , 
		w_14550 , w_14551 , w_14552 , w_14553 , w_14554 , w_14555 , w_14556 , w_14557 , w_14558 , w_14559 , 
		w_14560 , w_14561 , w_14562 , w_14563 , w_14564 , w_14565 , w_14566 , w_14567 , w_14568 , w_14569 , 
		w_14570 , w_14571 , w_14572 , w_14573 , w_14574 , w_14575 , w_14576 , w_14577 , w_14578 , w_14579 , 
		w_14580 , w_14581 , w_14582 , w_14583 , w_14584 , w_14585 , w_14586 , w_14587 , w_14588 , w_14589 , 
		w_14590 , w_14591 , w_14592 , w_14593 , w_14594 , w_14595 , w_14596 , w_14597 , w_14598 , w_14599 , 
		w_14600 , w_14601 , w_14602 , w_14603 , w_14604 , w_14605 , w_14606 , w_14607 , w_14608 , w_14609 , 
		w_14610 , w_14611 , w_14612 , w_14613 , w_14614 , w_14615 , w_14616 , w_14617 , w_14618 , w_14619 , 
		w_14620 , w_14621 , w_14622 , w_14623 , w_14624 , w_14625 , w_14626 , w_14627 , w_14628 , w_14629 , 
		w_14630 , w_14631 , w_14632 , w_14633 , w_14634 , w_14635 , w_14636 , w_14637 , w_14638 , w_14639 , 
		w_14640 , w_14641 , w_14642 , w_14643 , w_14644 , w_14645 , w_14646 , w_14647 , w_14648 , w_14649 , 
		w_14650 , w_14651 , w_14652 , w_14653 , w_14654 , w_14655 , w_14656 , w_14657 , w_14658 , w_14659 , 
		w_14660 , w_14661 , w_14662 , w_14663 , w_14664 , w_14665 , w_14666 , w_14667 , w_14668 , w_14669 , 
		w_14670 , w_14671 , w_14672 , w_14673 , w_14674 , w_14675 , w_14676 , w_14677 , w_14678 , w_14679 , 
		w_14680 , w_14681 , w_14682 , w_14683 , w_14684 , w_14685 , w_14686 , w_14687 , w_14688 , w_14689 , 
		w_14690 , w_14691 , w_14692 , w_14693 , w_14694 , w_14695 , w_14696 , w_14697 , w_14698 , w_14699 , 
		w_14700 , w_14701 , w_14702 , w_14703 , w_14704 , w_14705 , w_14706 , w_14707 , w_14708 , w_14709 , 
		w_14710 , w_14711 , w_14712 , w_14713 , w_14714 , w_14715 , w_14716 , w_14717 , w_14718 , w_14719 , 
		w_14720 , w_14721 , w_14722 , w_14723 , w_14724 , w_14725 , w_14726 , w_14727 , w_14728 , w_14729 , 
		w_14730 , w_14731 , w_14732 , w_14733 , w_14734 , w_14735 , w_14736 , w_14737 , w_14738 , w_14739 , 
		w_14740 , w_14741 , w_14742 , w_14743 , w_14744 , w_14745 , w_14746 , w_14747 , w_14748 , w_14749 , 
		w_14750 , w_14751 , w_14752 , w_14753 , w_14754 , w_14755 , w_14756 , w_14757 , w_14758 , w_14759 , 
		w_14760 , w_14761 , w_14762 , w_14763 , w_14764 , w_14765 , w_14766 , w_14767 , w_14768 , w_14769 , 
		w_14770 , w_14771 , w_14772 , w_14773 , w_14774 , w_14775 , w_14776 , w_14777 , w_14778 , w_14779 , 
		w_14780 , w_14781 , w_14782 , w_14783 , w_14784 , w_14785 , w_14786 , w_14787 , w_14788 , w_14789 , 
		w_14790 , w_14791 , w_14792 , w_14793 , w_14794 , w_14795 , w_14796 , w_14797 , w_14798 , w_14799 , 
		w_14800 , w_14801 , w_14802 , w_14803 , w_14804 , w_14805 , w_14806 , w_14807 , w_14808 , w_14809 , 
		w_14810 , w_14811 , w_14812 , w_14813 , w_14814 , w_14815 , w_14816 , w_14817 , w_14818 , w_14819 , 
		w_14820 , w_14821 , w_14822 , w_14823 , w_14824 , w_14825 , w_14826 , w_14827 , w_14828 , w_14829 , 
		w_14830 , w_14831 , w_14832 , w_14833 , w_14834 , w_14835 , w_14836 , w_14837 , w_14838 , w_14839 , 
		w_14840 , w_14841 , w_14842 , w_14843 , w_14844 , w_14845 , w_14846 , w_14847 , w_14848 , w_14849 , 
		w_14850 , w_14851 , w_14852 , w_14853 , w_14854 , w_14855 , w_14856 , w_14857 , w_14858 , w_14859 , 
		w_14860 , w_14861 , w_14862 , w_14863 , w_14864 , w_14865 , w_14866 , w_14867 , w_14868 , w_14869 , 
		w_14870 , w_14871 , w_14872 , w_14873 , w_14874 , w_14875 , w_14876 , w_14877 , w_14878 , w_14879 , 
		w_14880 , w_14881 , w_14882 , w_14883 , w_14884 , w_14885 , w_14886 , w_14887 , w_14888 , w_14889 , 
		w_14890 , w_14891 , w_14892 , w_14893 , w_14894 , w_14895 , w_14896 , w_14897 , w_14898 , w_14899 , 
		w_14900 , w_14901 , w_14902 , w_14903 , w_14904 , w_14905 , w_14906 , w_14907 , w_14908 , w_14909 , 
		w_14910 , w_14911 , w_14912 , w_14913 , w_14914 , w_14915 , w_14916 , w_14917 , w_14918 , w_14919 , 
		w_14920 , w_14921 , w_14922 , w_14923 , w_14924 , w_14925 , w_14926 , w_14927 , w_14928 , w_14929 , 
		w_14930 , w_14931 , w_14932 , w_14933 , w_14934 , w_14935 , w_14936 , w_14937 , w_14938 , w_14939 , 
		w_14940 , w_14941 , w_14942 , w_14943 , w_14944 , w_14945 , w_14946 , w_14947 , w_14948 , w_14949 , 
		w_14950 , w_14951 , w_14952 , w_14953 , w_14954 , w_14955 , w_14956 , w_14957 , w_14958 , w_14959 , 
		w_14960 , w_14961 , w_14962 , w_14963 , w_14964 , w_14965 , w_14966 , w_14967 , w_14968 , w_14969 , 
		w_14970 , w_14971 , w_14972 , w_14973 , w_14974 , w_14975 , w_14976 , w_14977 , w_14978 , w_14979 , 
		w_14980 , w_14981 , w_14982 , w_14983 , w_14984 , w_14985 , w_14986 , w_14987 , w_14988 , w_14989 , 
		w_14990 , w_14991 , w_14992 , w_14993 , w_14994 , w_14995 , w_14996 , w_14997 , w_14998 , w_14999 , 
		w_15000 , w_15001 , w_15002 , w_15003 , w_15004 , w_15005 , w_15006 , w_15007 , w_15008 , w_15009 , 
		w_15010 , w_15011 , w_15012 , w_15013 , w_15014 , w_15015 , w_15016 , w_15017 , w_15018 , w_15019 , 
		w_15020 , w_15021 , w_15022 , w_15023 , w_15024 , w_15025 , w_15026 , w_15027 , w_15028 , w_15029 , 
		w_15030 , w_15031 , w_15032 , w_15033 , w_15034 , w_15035 , w_15036 , w_15037 , w_15038 , w_15039 , 
		w_15040 , w_15041 , w_15042 , w_15043 , w_15044 , w_15045 , w_15046 , w_15047 , w_15048 , w_15049 , 
		w_15050 , w_15051 , w_15052 , w_15053 , w_15054 , w_15055 , w_15056 , w_15057 , w_15058 , w_15059 , 
		w_15060 , w_15061 , w_15062 , w_15063 , w_15064 , w_15065 , w_15066 , w_15067 , w_15068 , w_15069 , 
		w_15070 , w_15071 , w_15072 , w_15073 , w_15074 , w_15075 , w_15076 , w_15077 , w_15078 , w_15079 , 
		w_15080 , w_15081 , w_15082 , w_15083 , w_15084 , w_15085 , w_15086 , w_15087 , w_15088 , w_15089 , 
		w_15090 , w_15091 , w_15092 , w_15093 , w_15094 , w_15095 , w_15096 , w_15097 , w_15098 , w_15099 , 
		w_15100 , w_15101 , w_15102 , w_15103 , w_15104 , w_15105 , w_15106 , w_15107 , w_15108 , w_15109 , 
		w_15110 , w_15111 , w_15112 , w_15113 , w_15114 , w_15115 , w_15116 , w_15117 , w_15118 , w_15119 , 
		w_15120 , w_15121 , w_15122 , w_15123 , w_15124 , w_15125 , w_15126 , w_15127 , w_15128 , w_15129 , 
		w_15130 , w_15131 , w_15132 , w_15133 , w_15134 , w_15135 , w_15136 , w_15137 , w_15138 , w_15139 , 
		w_15140 , w_15141 , w_15142 , w_15143 , w_15144 , w_15145 , w_15146 , w_15147 , w_15148 , w_15149 , 
		w_15150 , w_15151 , w_15152 , w_15153 , w_15154 , w_15155 , w_15156 , w_15157 , w_15158 , w_15159 , 
		w_15160 , w_15161 , w_15162 , w_15163 , w_15164 , w_15165 , w_15166 , w_15167 , w_15168 , w_15169 , 
		w_15170 , w_15171 , w_15172 , w_15173 , w_15174 , w_15175 , w_15176 , w_15177 , w_15178 , w_15179 , 
		w_15180 , w_15181 , w_15182 , w_15183 , w_15184 , w_15185 , w_15186 , w_15187 , w_15188 , w_15189 , 
		w_15190 , w_15191 , w_15192 , w_15193 , w_15194 , w_15195 , w_15196 , w_15197 , w_15198 , w_15199 , 
		w_15200 , w_15201 , w_15202 , w_15203 , w_15204 , w_15205 , w_15206 , w_15207 , w_15208 , w_15209 , 
		w_15210 , w_15211 , w_15212 , w_15213 , w_15214 , w_15215 , w_15216 , w_15217 , w_15218 , w_15219 , 
		w_15220 , w_15221 , w_15222 , w_15223 , w_15224 , w_15225 , w_15226 , w_15227 , w_15228 , w_15229 , 
		w_15230 , w_15231 , w_15232 , w_15233 , w_15234 , w_15235 , w_15236 , w_15237 , w_15238 , w_15239 , 
		w_15240 , w_15241 , w_15242 , w_15243 , w_15244 , w_15245 , w_15246 , w_15247 , w_15248 , w_15249 , 
		w_15250 , w_15251 , w_15252 , w_15253 , w_15254 , w_15255 , w_15256 , w_15257 , w_15258 , w_15259 , 
		w_15260 , w_15261 , w_15262 , w_15263 , w_15264 , w_15265 , w_15266 , w_15267 , w_15268 , w_15269 , 
		w_15270 , w_15271 , w_15272 , w_15273 , w_15274 , w_15275 , w_15276 , w_15277 , w_15278 , w_15279 , 
		w_15280 , w_15281 , w_15282 , w_15283 , w_15284 , w_15285 , w_15286 , w_15287 , w_15288 , w_15289 , 
		w_15290 , w_15291 , w_15292 , w_15293 , w_15294 , w_15295 , w_15296 , w_15297 , w_15298 , w_15299 , 
		w_15300 , w_15301 , w_15302 , w_15303 , w_15304 , w_15305 , w_15306 , w_15307 , w_15308 , w_15309 , 
		w_15310 , w_15311 , w_15312 , w_15313 , w_15314 , w_15315 , w_15316 , w_15317 , w_15318 , w_15319 , 
		w_15320 , w_15321 , w_15322 , w_15323 , w_15324 , w_15325 , w_15326 , w_15327 , w_15328 , w_15329 , 
		w_15330 , w_15331 , w_15332 , w_15333 , w_15334 , w_15335 , w_15336 , w_15337 , w_15338 , w_15339 , 
		w_15340 , w_15341 , w_15342 , w_15343 , w_15344 , w_15345 , w_15346 , w_15347 , w_15348 , w_15349 , 
		w_15350 , w_15351 , w_15352 , w_15353 , w_15354 , w_15355 , w_15356 , w_15357 , w_15358 , w_15359 , 
		w_15360 , w_15361 , w_15362 , w_15363 , w_15364 , w_15365 , w_15366 , w_15367 , w_15368 , w_15369 , 
		w_15370 , w_15371 , w_15372 , w_15373 , w_15374 , w_15375 , w_15376 , w_15377 , w_15378 , w_15379 , 
		w_15380 , w_15381 , w_15382 , w_15383 , w_15384 , w_15385 , w_15386 , w_15387 , w_15388 , w_15389 , 
		w_15390 , w_15391 , w_15392 , w_15393 , w_15394 , w_15395 , w_15396 , w_15397 , w_15398 , w_15399 , 
		w_15400 , w_15401 , w_15402 , w_15403 , w_15404 , w_15405 , w_15406 , w_15407 , w_15408 , w_15409 , 
		w_15410 , w_15411 , w_15412 , w_15413 , w_15414 , w_15415 , w_15416 , w_15417 , w_15418 , w_15419 , 
		w_15420 , w_15421 , w_15422 , w_15423 , w_15424 , w_15425 , w_15426 , w_15427 , w_15428 , w_15429 , 
		w_15430 , w_15431 , w_15432 , w_15433 , w_15434 , w_15435 , w_15436 , w_15437 , w_15438 , w_15439 , 
		w_15440 , w_15441 , w_15442 , w_15443 , w_15444 , w_15445 , w_15446 , w_15447 , w_15448 , w_15449 , 
		w_15450 , w_15451 , w_15452 , w_15453 , w_15454 , w_15455 , w_15456 , w_15457 , w_15458 , w_15459 , 
		w_15460 , w_15461 , w_15462 , w_15463 , w_15464 , w_15465 , w_15466 , w_15467 , w_15468 , w_15469 , 
		w_15470 , w_15471 , w_15472 , w_15473 , w_15474 , w_15475 , w_15476 , w_15477 , w_15478 , w_15479 , 
		w_15480 , w_15481 , w_15482 , w_15483 , w_15484 , w_15485 , w_15486 , w_15487 , w_15488 , w_15489 , 
		w_15490 , w_15491 , w_15492 , w_15493 , w_15494 , w_15495 , w_15496 , w_15497 , w_15498 , w_15499 , 
		w_15500 , w_15501 , w_15502 , w_15503 , w_15504 , w_15505 , w_15506 , w_15507 , w_15508 , w_15509 , 
		w_15510 , w_15511 , w_15512 , w_15513 , w_15514 , w_15515 , w_15516 , w_15517 , w_15518 , w_15519 , 
		w_15520 , w_15521 , w_15522 , w_15523 , w_15524 , w_15525 , w_15526 , w_15527 , w_15528 , w_15529 , 
		w_15530 , w_15531 , w_15532 , w_15533 , w_15534 , w_15535 , w_15536 , w_15537 , w_15538 , w_15539 , 
		w_15540 , w_15541 , w_15542 , w_15543 , w_15544 , w_15545 , w_15546 , w_15547 , w_15548 , w_15549 , 
		w_15550 , w_15551 , w_15552 , w_15553 , w_15554 , w_15555 , w_15556 , w_15557 , w_15558 , w_15559 , 
		w_15560 , w_15561 , w_15562 , w_15563 , w_15564 , w_15565 , w_15566 , w_15567 , w_15568 , w_15569 , 
		w_15570 , w_15571 , w_15572 , w_15573 , w_15574 , w_15575 , w_15576 , w_15577 , w_15578 , w_15579 , 
		w_15580 , w_15581 , w_15582 , w_15583 , w_15584 , w_15585 , w_15586 , w_15587 , w_15588 , w_15589 , 
		w_15590 , w_15591 , w_15592 , w_15593 , w_15594 , w_15595 , w_15596 , w_15597 , w_15598 , w_15599 , 
		w_15600 , w_15601 , w_15602 , w_15603 , w_15604 , w_15605 , w_15606 , w_15607 , w_15608 , w_15609 , 
		w_15610 , w_15611 , w_15612 , w_15613 , w_15614 , w_15615 , w_15616 , w_15617 , w_15618 , w_15619 , 
		w_15620 , w_15621 , w_15622 , w_15623 , w_15624 , w_15625 , w_15626 , w_15627 , w_15628 , w_15629 , 
		w_15630 , w_15631 , w_15632 , w_15633 , w_15634 , w_15635 , w_15636 , w_15637 , w_15638 , w_15639 , 
		w_15640 , w_15641 , w_15642 , w_15643 , w_15644 , w_15645 , w_15646 , w_15647 , w_15648 , w_15649 , 
		w_15650 , w_15651 , w_15652 , w_15653 , w_15654 , w_15655 , w_15656 , w_15657 , w_15658 , w_15659 , 
		w_15660 , w_15661 , w_15662 , w_15663 , w_15664 , w_15665 , w_15666 , w_15667 , w_15668 , w_15669 , 
		w_15670 , w_15671 , w_15672 , w_15673 , w_15674 , w_15675 , w_15676 , w_15677 , w_15678 , w_15679 , 
		w_15680 , w_15681 , w_15682 , w_15683 , w_15684 , w_15685 , w_15686 , w_15687 , w_15688 , w_15689 , 
		w_15690 , w_15691 , w_15692 , w_15693 , w_15694 , w_15695 , w_15696 , w_15697 , w_15698 , w_15699 , 
		w_15700 , w_15701 , w_15702 , w_15703 , w_15704 , w_15705 , w_15706 , w_15707 , w_15708 , w_15709 , 
		w_15710 , w_15711 , w_15712 , w_15713 , w_15714 , w_15715 , w_15716 , w_15717 , w_15718 , w_15719 , 
		w_15720 , w_15721 , w_15722 , w_15723 , w_15724 , w_15725 , w_15726 , w_15727 , w_15728 , w_15729 , 
		w_15730 , w_15731 , w_15732 , w_15733 , w_15734 , w_15735 , w_15736 , w_15737 , w_15738 , w_15739 , 
		w_15740 , w_15741 , w_15742 , w_15743 , w_15744 , w_15745 , w_15746 , w_15747 , w_15748 , w_15749 , 
		w_15750 , w_15751 , w_15752 , w_15753 , w_15754 , w_15755 , w_15756 , w_15757 , w_15758 , w_15759 , 
		w_15760 , w_15761 , w_15762 , w_15763 , w_15764 , w_15765 , w_15766 , w_15767 , w_15768 , w_15769 , 
		w_15770 , w_15771 , w_15772 , w_15773 , w_15774 , w_15775 , w_15776 , w_15777 , w_15778 , w_15779 , 
		w_15780 , w_15781 , w_15782 , w_15783 , w_15784 , w_15785 , w_15786 , w_15787 , w_15788 , w_15789 , 
		w_15790 , w_15791 , w_15792 , w_15793 , w_15794 , w_15795 , w_15796 , w_15797 , w_15798 , w_15799 , 
		w_15800 , w_15801 , w_15802 , w_15803 , w_15804 , w_15805 , w_15806 , w_15807 , w_15808 , w_15809 , 
		w_15810 , w_15811 , w_15812 , w_15813 , w_15814 , w_15815 , w_15816 , w_15817 , w_15818 , w_15819 , 
		w_15820 , w_15821 , w_15822 , w_15823 , w_15824 , w_15825 , w_15826 , w_15827 , w_15828 , w_15829 , 
		w_15830 , w_15831 , w_15832 , w_15833 , w_15834 , w_15835 , w_15836 , w_15837 , w_15838 , w_15839 , 
		w_15840 , w_15841 , w_15842 , w_15843 , w_15844 , w_15845 , w_15846 , w_15847 , w_15848 , w_15849 , 
		w_15850 , w_15851 , w_15852 , w_15853 , w_15854 , w_15855 , w_15856 , w_15857 , w_15858 , w_15859 , 
		w_15860 , w_15861 , w_15862 , w_15863 , w_15864 , w_15865 , w_15866 , w_15867 , w_15868 , w_15869 , 
		w_15870 , w_15871 , w_15872 , w_15873 , w_15874 , w_15875 , w_15876 , w_15877 , w_15878 , w_15879 , 
		w_15880 , w_15881 , w_15882 , w_15883 , w_15884 , w_15885 , w_15886 , w_15887 , w_15888 , w_15889 , 
		w_15890 , w_15891 , w_15892 , w_15893 , w_15894 , w_15895 , w_15896 , w_15897 , w_15898 , w_15899 , 
		w_15900 , w_15901 , w_15902 , w_15903 , w_15904 , w_15905 , w_15906 , w_15907 , w_15908 , w_15909 , 
		w_15910 , w_15911 , w_15912 , w_15913 , w_15914 , w_15915 , w_15916 , w_15917 , w_15918 , w_15919 , 
		w_15920 , w_15921 , w_15922 , w_15923 , w_15924 , w_15925 , w_15926 , w_15927 , w_15928 , w_15929 , 
		w_15930 , w_15931 , w_15932 , w_15933 , w_15934 , w_15935 , w_15936 , w_15937 , w_15938 , w_15939 , 
		w_15940 , w_15941 , w_15942 , w_15943 , w_15944 , w_15945 , w_15946 , w_15947 , w_15948 , w_15949 , 
		w_15950 , w_15951 , w_15952 , w_15953 , w_15954 , w_15955 , w_15956 , w_15957 , w_15958 , w_15959 , 
		w_15960 , w_15961 , w_15962 , w_15963 , w_15964 , w_15965 , w_15966 , w_15967 , w_15968 , w_15969 , 
		w_15970 , w_15971 , w_15972 , w_15973 , w_15974 , w_15975 , w_15976 , w_15977 , w_15978 , w_15979 , 
		w_15980 , w_15981 , w_15982 , w_15983 , w_15984 , w_15985 , w_15986 , w_15987 , w_15988 , w_15989 , 
		w_15990 , w_15991 , w_15992 , w_15993 , w_15994 , w_15995 , w_15996 , w_15997 , w_15998 , w_15999 , 
		w_16000 , w_16001 , w_16002 , w_16003 , w_16004 , w_16005 , w_16006 , w_16007 , w_16008 , w_16009 , 
		w_16010 , w_16011 , w_16012 , w_16013 , w_16014 , w_16015 , w_16016 , w_16017 , w_16018 , w_16019 , 
		w_16020 , w_16021 , w_16022 , w_16023 , w_16024 , w_16025 , w_16026 , w_16027 , w_16028 , w_16029 , 
		w_16030 , w_16031 , w_16032 , w_16033 , w_16034 , w_16035 , w_16036 , w_16037 , w_16038 , w_16039 , 
		w_16040 , w_16041 , w_16042 , w_16043 , w_16044 , w_16045 , w_16046 , w_16047 , w_16048 , w_16049 , 
		w_16050 , w_16051 , w_16052 , w_16053 , w_16054 , w_16055 , w_16056 , w_16057 , w_16058 , w_16059 , 
		w_16060 , w_16061 , w_16062 , w_16063 , w_16064 , w_16065 , w_16066 , w_16067 , w_16068 , w_16069 , 
		w_16070 , w_16071 , w_16072 , w_16073 , w_16074 , w_16075 , w_16076 , w_16077 , w_16078 , w_16079 , 
		w_16080 , w_16081 , w_16082 , w_16083 , w_16084 , w_16085 , w_16086 , w_16087 , w_16088 , w_16089 , 
		w_16090 , w_16091 , w_16092 , w_16093 , w_16094 , w_16095 , w_16096 , w_16097 , w_16098 , w_16099 , 
		w_16100 , w_16101 , w_16102 , w_16103 , w_16104 , w_16105 , w_16106 , w_16107 , w_16108 , w_16109 , 
		w_16110 , w_16111 , w_16112 , w_16113 , w_16114 , w_16115 , w_16116 , w_16117 , w_16118 , w_16119 , 
		w_16120 , w_16121 , w_16122 , w_16123 , w_16124 , w_16125 , w_16126 , w_16127 , w_16128 , w_16129 , 
		w_16130 , w_16131 , w_16132 , w_16133 , w_16134 , w_16135 , w_16136 , w_16137 , w_16138 , w_16139 , 
		w_16140 , w_16141 , w_16142 , w_16143 , w_16144 , w_16145 , w_16146 , w_16147 , w_16148 , w_16149 , 
		w_16150 , w_16151 , w_16152 , w_16153 , w_16154 , w_16155 , w_16156 , w_16157 , w_16158 , w_16159 , 
		w_16160 , w_16161 , w_16162 , w_16163 , w_16164 , w_16165 , w_16166 , w_16167 , w_16168 , w_16169 , 
		w_16170 , w_16171 , w_16172 , w_16173 , w_16174 , w_16175 , w_16176 , w_16177 , w_16178 , w_16179 , 
		w_16180 , w_16181 , w_16182 , w_16183 , w_16184 , w_16185 , w_16186 , w_16187 , w_16188 , w_16189 , 
		w_16190 , w_16191 , w_16192 , w_16193 , w_16194 , w_16195 , w_16196 , w_16197 , w_16198 , w_16199 , 
		w_16200 , w_16201 , w_16202 , w_16203 , w_16204 , w_16205 , w_16206 , w_16207 , w_16208 , w_16209 , 
		w_16210 , w_16211 , w_16212 , w_16213 , w_16214 , w_16215 , w_16216 , w_16217 , w_16218 , w_16219 , 
		w_16220 , w_16221 , w_16222 , w_16223 , w_16224 , w_16225 , w_16226 , w_16227 , w_16228 , w_16229 , 
		w_16230 , w_16231 , w_16232 , w_16233 , w_16234 , w_16235 , w_16236 , w_16237 , w_16238 , w_16239 , 
		w_16240 , w_16241 , w_16242 , w_16243 , w_16244 , w_16245 , w_16246 , w_16247 , w_16248 , w_16249 , 
		w_16250 , w_16251 , w_16252 , w_16253 , w_16254 , w_16255 , w_16256 , w_16257 , w_16258 , w_16259 , 
		w_16260 , w_16261 , w_16262 , w_16263 , w_16264 , w_16265 , w_16266 , w_16267 , w_16268 , w_16269 , 
		w_16270 , w_16271 , w_16272 , w_16273 , w_16274 , w_16275 , w_16276 , w_16277 , w_16278 , w_16279 , 
		w_16280 , w_16281 , w_16282 , w_16283 , w_16284 , w_16285 , w_16286 , w_16287 , w_16288 , w_16289 , 
		w_16290 , w_16291 , w_16292 , w_16293 , w_16294 , w_16295 , w_16296 , w_16297 , w_16298 , w_16299 , 
		w_16300 , w_16301 , w_16302 , w_16303 , w_16304 , w_16305 , w_16306 , w_16307 , w_16308 , w_16309 , 
		w_16310 , w_16311 , w_16312 , w_16313 , w_16314 , w_16315 , w_16316 , w_16317 , w_16318 , w_16319 , 
		w_16320 , w_16321 , w_16322 , w_16323 , w_16324 , w_16325 , w_16326 , w_16327 , w_16328 , w_16329 , 
		w_16330 , w_16331 , w_16332 , w_16333 , w_16334 , w_16335 , w_16336 , w_16337 , w_16338 , w_16339 , 
		w_16340 , w_16341 , w_16342 , w_16343 , w_16344 , w_16345 , w_16346 , w_16347 , w_16348 , w_16349 , 
		w_16350 , w_16351 , w_16352 , w_16353 , w_16354 , w_16355 , w_16356 , w_16357 , w_16358 , w_16359 , 
		w_16360 , w_16361 , w_16362 , w_16363 , w_16364 , w_16365 , w_16366 , w_16367 , w_16368 , w_16369 , 
		w_16370 , w_16371 , w_16372 , w_16373 , w_16374 , w_16375 , w_16376 , w_16377 , w_16378 , w_16379 , 
		w_16380 , w_16381 , w_16382 , w_16383 , w_16384 , w_16385 , w_16386 , w_16387 , w_16388 , w_16389 , 
		w_16390 , w_16391 , w_16392 , w_16393 , w_16394 , w_16395 , w_16396 , w_16397 , w_16398 , w_16399 , 
		w_16400 , w_16401 , w_16402 , w_16403 , w_16404 , w_16405 , w_16406 , w_16407 , w_16408 , w_16409 , 
		w_16410 , w_16411 , w_16412 , w_16413 , w_16414 , w_16415 , w_16416 , w_16417 , w_16418 , w_16419 , 
		w_16420 , w_16421 , w_16422 , w_16423 , w_16424 , w_16425 , w_16426 , w_16427 , w_16428 , w_16429 , 
		w_16430 , w_16431 , w_16432 , w_16433 , w_16434 , w_16435 , w_16436 , w_16437 , w_16438 , w_16439 , 
		w_16440 , w_16441 , w_16442 , w_16443 , w_16444 , w_16445 , w_16446 , w_16447 , w_16448 , w_16449 , 
		w_16450 , w_16451 , w_16452 , w_16453 , w_16454 , w_16455 , w_16456 , w_16457 , w_16458 , w_16459 , 
		w_16460 , w_16461 , w_16462 , w_16463 , w_16464 , w_16465 , w_16466 , w_16467 , w_16468 , w_16469 , 
		w_16470 , w_16471 , w_16472 , w_16473 , w_16474 , w_16475 , w_16476 , w_16477 , w_16478 , w_16479 , 
		w_16480 , w_16481 , w_16482 , w_16483 , w_16484 , w_16485 , w_16486 , w_16487 , w_16488 , w_16489 , 
		w_16490 , w_16491 , w_16492 , w_16493 , w_16494 , w_16495 , w_16496 , w_16497 , w_16498 , w_16499 , 
		w_16500 , w_16501 , w_16502 , w_16503 , w_16504 , w_16505 , w_16506 , w_16507 , w_16508 , w_16509 , 
		w_16510 , w_16511 , w_16512 , w_16513 , w_16514 , w_16515 , w_16516 , w_16517 , w_16518 , w_16519 , 
		w_16520 , w_16521 , w_16522 , w_16523 , w_16524 , w_16525 , w_16526 , w_16527 , w_16528 , w_16529 , 
		w_16530 , w_16531 , w_16532 , w_16533 , w_16534 , w_16535 , w_16536 , w_16537 , w_16538 , w_16539 , 
		w_16540 , w_16541 , w_16542 , w_16543 , w_16544 , w_16545 , w_16546 , w_16547 , w_16548 , w_16549 , 
		w_16550 , w_16551 , w_16552 , w_16553 , w_16554 , w_16555 , w_16556 , w_16557 , w_16558 , w_16559 , 
		w_16560 , w_16561 , w_16562 , w_16563 , w_16564 , w_16565 , w_16566 , w_16567 , w_16568 , w_16569 , 
		w_16570 , w_16571 , w_16572 , w_16573 , w_16574 , w_16575 , w_16576 , w_16577 , w_16578 , w_16579 , 
		w_16580 , w_16581 , w_16582 , w_16583 , w_16584 , w_16585 , w_16586 , w_16587 , w_16588 , w_16589 , 
		w_16590 , w_16591 , w_16592 , w_16593 , w_16594 , w_16595 , w_16596 , w_16597 , w_16598 , w_16599 , 
		w_16600 , w_16601 , w_16602 , w_16603 , w_16604 , w_16605 , w_16606 , w_16607 , w_16608 , w_16609 , 
		w_16610 , w_16611 , w_16612 , w_16613 , w_16614 , w_16615 , w_16616 , w_16617 , w_16618 , w_16619 , 
		w_16620 , w_16621 , w_16622 , w_16623 , w_16624 , w_16625 , w_16626 , w_16627 , w_16628 , w_16629 , 
		w_16630 , w_16631 , w_16632 , w_16633 , w_16634 , w_16635 , w_16636 , w_16637 , w_16638 , w_16639 , 
		w_16640 , w_16641 , w_16642 , w_16643 , w_16644 , w_16645 , w_16646 , w_16647 , w_16648 , w_16649 , 
		w_16650 , w_16651 , w_16652 , w_16653 , w_16654 , w_16655 , w_16656 , w_16657 , w_16658 , w_16659 , 
		w_16660 , w_16661 , w_16662 , w_16663 , w_16664 , w_16665 , w_16666 , w_16667 , w_16668 , w_16669 , 
		w_16670 , w_16671 , w_16672 , w_16673 , w_16674 , w_16675 , w_16676 , w_16677 , w_16678 , w_16679 , 
		w_16680 , w_16681 , w_16682 , w_16683 , w_16684 , w_16685 , w_16686 , w_16687 , w_16688 , w_16689 , 
		w_16690 , w_16691 , w_16692 , w_16693 , w_16694 , w_16695 , w_16696 , w_16697 , w_16698 , w_16699 , 
		w_16700 , w_16701 , w_16702 , w_16703 , w_16704 , w_16705 , w_16706 , w_16707 , w_16708 , w_16709 , 
		w_16710 , w_16711 , w_16712 , w_16713 , w_16714 , w_16715 , w_16716 , w_16717 , w_16718 , w_16719 , 
		w_16720 , w_16721 , w_16722 , w_16723 , w_16724 , w_16725 , w_16726 , w_16727 , w_16728 , w_16729 , 
		w_16730 , w_16731 , w_16732 , w_16733 , w_16734 , w_16735 , w_16736 , w_16737 , w_16738 , w_16739 , 
		w_16740 , w_16741 , w_16742 , w_16743 , w_16744 , w_16745 , w_16746 , w_16747 , w_16748 , w_16749 , 
		w_16750 , w_16751 , w_16752 , w_16753 , w_16754 , w_16755 , w_16756 , w_16757 , w_16758 , w_16759 , 
		w_16760 , w_16761 , w_16762 , w_16763 , w_16764 , w_16765 , w_16766 , w_16767 , w_16768 , w_16769 , 
		w_16770 , w_16771 , w_16772 , w_16773 , w_16774 , w_16775 , w_16776 , w_16777 , w_16778 , w_16779 , 
		w_16780 , w_16781 , w_16782 , w_16783 , w_16784 , w_16785 , w_16786 , w_16787 , w_16788 , w_16789 , 
		w_16790 , w_16791 , w_16792 , w_16793 , w_16794 , w_16795 , w_16796 , w_16797 , w_16798 , w_16799 , 
		w_16800 , w_16801 , w_16802 , w_16803 , w_16804 , w_16805 , w_16806 , w_16807 , w_16808 , w_16809 , 
		w_16810 , w_16811 , w_16812 , w_16813 , w_16814 , w_16815 , w_16816 , w_16817 , w_16818 , w_16819 , 
		w_16820 , w_16821 , w_16822 , w_16823 , w_16824 , w_16825 , w_16826 , w_16827 , w_16828 , w_16829 , 
		w_16830 , w_16831 , w_16832 , w_16833 , w_16834 , w_16835 , w_16836 , w_16837 , w_16838 , w_16839 , 
		w_16840 , w_16841 , w_16842 , w_16843 , w_16844 , w_16845 , w_16846 , w_16847 , w_16848 , w_16849 , 
		w_16850 , w_16851 , w_16852 , w_16853 , w_16854 , w_16855 , w_16856 , w_16857 , w_16858 , w_16859 , 
		w_16860 , w_16861 , w_16862 , w_16863 , w_16864 , w_16865 , w_16866 , w_16867 , w_16868 , w_16869 , 
		w_16870 , w_16871 , w_16872 , w_16873 , w_16874 , w_16875 , w_16876 , w_16877 , w_16878 , w_16879 , 
		w_16880 , w_16881 , w_16882 , w_16883 , w_16884 , w_16885 , w_16886 , w_16887 , w_16888 , w_16889 , 
		w_16890 , w_16891 , w_16892 , w_16893 , w_16894 , w_16895 , w_16896 , w_16897 , w_16898 , w_16899 , 
		w_16900 , w_16901 , w_16902 , w_16903 , w_16904 , w_16905 , w_16906 , w_16907 , w_16908 , w_16909 , 
		w_16910 , w_16911 , w_16912 , w_16913 , w_16914 , w_16915 , w_16916 , w_16917 , w_16918 , w_16919 , 
		w_16920 , w_16921 , w_16922 , w_16923 , w_16924 , w_16925 , w_16926 , w_16927 , w_16928 , w_16929 , 
		w_16930 , w_16931 , w_16932 , w_16933 , w_16934 , w_16935 , w_16936 , w_16937 , w_16938 , w_16939 , 
		w_16940 , w_16941 , w_16942 , w_16943 , w_16944 , w_16945 , w_16946 , w_16947 , w_16948 , w_16949 , 
		w_16950 , w_16951 , w_16952 , w_16953 , w_16954 , w_16955 , w_16956 , w_16957 , w_16958 , w_16959 , 
		w_16960 , w_16961 , w_16962 , w_16963 , w_16964 , w_16965 , w_16966 , w_16967 , w_16968 , w_16969 , 
		w_16970 , w_16971 , w_16972 , w_16973 , w_16974 , w_16975 , w_16976 , w_16977 , w_16978 , w_16979 , 
		w_16980 , w_16981 , w_16982 , w_16983 , w_16984 , w_16985 , w_16986 , w_16987 , w_16988 , w_16989 , 
		w_16990 , w_16991 , w_16992 , w_16993 , w_16994 , w_16995 , w_16996 , w_16997 , w_16998 , w_16999 , 
		w_17000 , w_17001 , w_17002 , w_17003 , w_17004 , w_17005 , w_17006 , w_17007 , w_17008 , w_17009 , 
		w_17010 , w_17011 , w_17012 , w_17013 , w_17014 , w_17015 , w_17016 , w_17017 , w_17018 , w_17019 , 
		w_17020 , w_17021 , w_17022 , w_17023 , w_17024 , w_17025 , w_17026 , w_17027 , w_17028 , w_17029 , 
		w_17030 , w_17031 , w_17032 , w_17033 , w_17034 , w_17035 , w_17036 , w_17037 , w_17038 , w_17039 , 
		w_17040 , w_17041 , w_17042 , w_17043 , w_17044 , w_17045 , w_17046 , w_17047 , w_17048 , w_17049 , 
		w_17050 , w_17051 , w_17052 , w_17053 , w_17054 , w_17055 , w_17056 , w_17057 , w_17058 , w_17059 , 
		w_17060 , w_17061 , w_17062 , w_17063 , w_17064 , w_17065 , w_17066 , w_17067 , w_17068 , w_17069 , 
		w_17070 , w_17071 , w_17072 , w_17073 , w_17074 , w_17075 , w_17076 , w_17077 , w_17078 , w_17079 , 
		w_17080 , w_17081 , w_17082 , w_17083 , w_17084 , w_17085 , w_17086 , w_17087 , w_17088 , w_17089 , 
		w_17090 , w_17091 , w_17092 , w_17093 , w_17094 , w_17095 , w_17096 , w_17097 , w_17098 , w_17099 , 
		w_17100 , w_17101 , w_17102 , w_17103 , w_17104 , w_17105 , w_17106 , w_17107 , w_17108 , w_17109 , 
		w_17110 , w_17111 , w_17112 , w_17113 , w_17114 , w_17115 , w_17116 , w_17117 , w_17118 , w_17119 , 
		w_17120 , w_17121 , w_17122 , w_17123 , w_17124 , w_17125 , w_17126 , w_17127 , w_17128 , w_17129 , 
		w_17130 , w_17131 , w_17132 , w_17133 , w_17134 , w_17135 , w_17136 , w_17137 , w_17138 , w_17139 , 
		w_17140 , w_17141 , w_17142 , w_17143 , w_17144 , w_17145 , w_17146 , w_17147 , w_17148 , w_17149 , 
		w_17150 , w_17151 , w_17152 , w_17153 , w_17154 , w_17155 , w_17156 , w_17157 , w_17158 , w_17159 , 
		w_17160 , w_17161 , w_17162 , w_17163 , w_17164 , w_17165 , w_17166 , w_17167 , w_17168 , w_17169 , 
		w_17170 , w_17171 , w_17172 , w_17173 , w_17174 , w_17175 , w_17176 , w_17177 , w_17178 , w_17179 , 
		w_17180 , w_17181 , w_17182 , w_17183 , w_17184 , w_17185 , w_17186 , w_17187 , w_17188 , w_17189 , 
		w_17190 , w_17191 , w_17192 , w_17193 , w_17194 , w_17195 , w_17196 , w_17197 , w_17198 , w_17199 , 
		w_17200 , w_17201 , w_17202 , w_17203 , w_17204 , w_17205 , w_17206 , w_17207 , w_17208 , w_17209 , 
		w_17210 , w_17211 , w_17212 , w_17213 , w_17214 , w_17215 , w_17216 , w_17217 , w_17218 , w_17219 , 
		w_17220 , w_17221 , w_17222 , w_17223 , w_17224 , w_17225 , w_17226 , w_17227 , w_17228 , w_17229 , 
		w_17230 , w_17231 , w_17232 , w_17233 , w_17234 , w_17235 , w_17236 , w_17237 , w_17238 , w_17239 , 
		w_17240 , w_17241 , w_17242 , w_17243 , w_17244 , w_17245 , w_17246 , w_17247 , w_17248 , w_17249 , 
		w_17250 , w_17251 , w_17252 , w_17253 , w_17254 , w_17255 , w_17256 , w_17257 , w_17258 , w_17259 , 
		w_17260 , w_17261 , w_17262 , w_17263 , w_17264 , w_17265 , w_17266 , w_17267 , w_17268 , w_17269 , 
		w_17270 , w_17271 , w_17272 , w_17273 , w_17274 , w_17275 , w_17276 , w_17277 , w_17278 , w_17279 , 
		w_17280 , w_17281 , w_17282 , w_17283 , w_17284 , w_17285 , w_17286 , w_17287 , w_17288 , w_17289 , 
		w_17290 , w_17291 , w_17292 , w_17293 , w_17294 , w_17295 , w_17296 , w_17297 , w_17298 , w_17299 , 
		w_17300 , w_17301 , w_17302 , w_17303 , w_17304 , w_17305 , w_17306 , w_17307 , w_17308 , w_17309 , 
		w_17310 , w_17311 , w_17312 , w_17313 , w_17314 , w_17315 , w_17316 , w_17317 , w_17318 , w_17319 , 
		w_17320 , w_17321 , w_17322 , w_17323 , w_17324 , w_17325 , w_17326 , w_17327 , w_17328 , w_17329 , 
		w_17330 , w_17331 , w_17332 , w_17333 , w_17334 , w_17335 , w_17336 , w_17337 , w_17338 , w_17339 , 
		w_17340 , w_17341 , w_17342 , w_17343 , w_17344 , w_17345 , w_17346 , w_17347 , w_17348 , w_17349 , 
		w_17350 , w_17351 , w_17352 , w_17353 , w_17354 , w_17355 , w_17356 , w_17357 , w_17358 , w_17359 , 
		w_17360 , w_17361 , w_17362 , w_17363 , w_17364 , w_17365 , w_17366 , w_17367 , w_17368 , w_17369 , 
		w_17370 , w_17371 , w_17372 , w_17373 , w_17374 , w_17375 , w_17376 , w_17377 , w_17378 , w_17379 , 
		w_17380 , w_17381 , w_17382 , w_17383 , w_17384 , w_17385 , w_17386 , w_17387 , w_17388 , w_17389 , 
		w_17390 , w_17391 , w_17392 , w_17393 , w_17394 , w_17395 , w_17396 , w_17397 , w_17398 , w_17399 , 
		w_17400 , w_17401 , w_17402 , w_17403 , w_17404 , w_17405 , w_17406 , w_17407 , w_17408 , w_17409 , 
		w_17410 , w_17411 , w_17412 , w_17413 , w_17414 , w_17415 , w_17416 , w_17417 , w_17418 , w_17419 , 
		w_17420 , w_17421 , w_17422 , w_17423 , w_17424 , w_17425 , w_17426 , w_17427 , w_17428 , w_17429 , 
		w_17430 , w_17431 , w_17432 , w_17433 , w_17434 , w_17435 , w_17436 , w_17437 , w_17438 , w_17439 , 
		w_17440 , w_17441 , w_17442 , w_17443 , w_17444 , w_17445 , w_17446 , w_17447 , w_17448 , w_17449 , 
		w_17450 , w_17451 , w_17452 , w_17453 , w_17454 , w_17455 , w_17456 , w_17457 , w_17458 , w_17459 , 
		w_17460 , w_17461 , w_17462 , w_17463 , w_17464 , w_17465 , w_17466 , w_17467 , w_17468 , w_17469 , 
		w_17470 , w_17471 , w_17472 , w_17473 , w_17474 , w_17475 , w_17476 , w_17477 , w_17478 , w_17479 , 
		w_17480 , w_17481 , w_17482 , w_17483 , w_17484 , w_17485 , w_17486 , w_17487 , w_17488 , w_17489 , 
		w_17490 , w_17491 , w_17492 , w_17493 , w_17494 , w_17495 , w_17496 , w_17497 , w_17498 , w_17499 , 
		w_17500 , w_17501 , w_17502 , w_17503 , w_17504 , w_17505 , w_17506 , w_17507 , w_17508 , w_17509 , 
		w_17510 , w_17511 , w_17512 , w_17513 , w_17514 , w_17515 , w_17516 , w_17517 , w_17518 , w_17519 , 
		w_17520 , w_17521 , w_17522 , w_17523 , w_17524 , w_17525 , w_17526 , w_17527 , w_17528 , w_17529 , 
		w_17530 , w_17531 , w_17532 , w_17533 , w_17534 , w_17535 , w_17536 , w_17537 , w_17538 , w_17539 , 
		w_17540 , w_17541 , w_17542 , w_17543 , w_17544 , w_17545 , w_17546 , w_17547 , w_17548 , w_17549 , 
		w_17550 , w_17551 , w_17552 , w_17553 , w_17554 , w_17555 , w_17556 , w_17557 , w_17558 , w_17559 , 
		w_17560 , w_17561 , w_17562 , w_17563 , w_17564 , w_17565 , w_17566 , w_17567 , w_17568 , w_17569 , 
		w_17570 , w_17571 , w_17572 , w_17573 , w_17574 , w_17575 , w_17576 , w_17577 , w_17578 , w_17579 , 
		w_17580 , w_17581 , w_17582 , w_17583 , w_17584 , w_17585 , w_17586 , w_17587 , w_17588 , w_17589 , 
		w_17590 , w_17591 , w_17592 , w_17593 , w_17594 , w_17595 , w_17596 , w_17597 , w_17598 , w_17599 , 
		w_17600 , w_17601 , w_17602 , w_17603 , w_17604 , w_17605 , w_17606 , w_17607 , w_17608 , w_17609 , 
		w_17610 , w_17611 , w_17612 , w_17613 , w_17614 , w_17615 , w_17616 , w_17617 , w_17618 , w_17619 , 
		w_17620 , w_17621 , w_17622 , w_17623 , w_17624 , w_17625 , w_17626 , w_17627 , w_17628 , w_17629 , 
		w_17630 , w_17631 , w_17632 , w_17633 , w_17634 , w_17635 , w_17636 , w_17637 , w_17638 , w_17639 , 
		w_17640 , w_17641 , w_17642 , w_17643 , w_17644 , w_17645 , w_17646 , w_17647 , w_17648 , w_17649 , 
		w_17650 , w_17651 , w_17652 , w_17653 , w_17654 , w_17655 , w_17656 , w_17657 , w_17658 , w_17659 , 
		w_17660 , w_17661 , w_17662 , w_17663 , w_17664 , w_17665 , w_17666 , w_17667 , w_17668 , w_17669 , 
		w_17670 , w_17671 , w_17672 , w_17673 , w_17674 , w_17675 , w_17676 , w_17677 , w_17678 , w_17679 , 
		w_17680 , w_17681 , w_17682 , w_17683 , w_17684 , w_17685 , w_17686 , w_17687 , w_17688 , w_17689 , 
		w_17690 , w_17691 , w_17692 , w_17693 , w_17694 , w_17695 , w_17696 , w_17697 , w_17698 , w_17699 , 
		w_17700 , w_17701 , w_17702 , w_17703 , w_17704 , w_17705 , w_17706 , w_17707 , w_17708 , w_17709 , 
		w_17710 , w_17711 , w_17712 , w_17713 , w_17714 , w_17715 , w_17716 , w_17717 , w_17718 , w_17719 , 
		w_17720 , w_17721 , w_17722 , w_17723 , w_17724 , w_17725 , w_17726 , w_17727 , w_17728 , w_17729 , 
		w_17730 , w_17731 , w_17732 , w_17733 , w_17734 , w_17735 , w_17736 , w_17737 , w_17738 , w_17739 , 
		w_17740 , w_17741 , w_17742 , w_17743 , w_17744 , w_17745 , w_17746 , w_17747 , w_17748 , w_17749 , 
		w_17750 , w_17751 , w_17752 , w_17753 , w_17754 , w_17755 , w_17756 , w_17757 , w_17758 , w_17759 , 
		w_17760 , w_17761 , w_17762 , w_17763 , w_17764 , w_17765 , w_17766 , w_17767 , w_17768 , w_17769 , 
		w_17770 , w_17771 , w_17772 , w_17773 , w_17774 , w_17775 , w_17776 , w_17777 , w_17778 , w_17779 , 
		w_17780 , w_17781 , w_17782 , w_17783 , w_17784 , w_17785 , w_17786 , w_17787 , w_17788 , w_17789 , 
		w_17790 , w_17791 , w_17792 , w_17793 , w_17794 , w_17795 , w_17796 , w_17797 , w_17798 , w_17799 , 
		w_17800 , w_17801 , w_17802 , w_17803 , w_17804 , w_17805 , w_17806 , w_17807 , w_17808 , w_17809 , 
		w_17810 , w_17811 , w_17812 , w_17813 , w_17814 , w_17815 , w_17816 , w_17817 , w_17818 , w_17819 , 
		w_17820 , w_17821 , w_17822 , w_17823 , w_17824 , w_17825 , w_17826 , w_17827 , w_17828 , w_17829 , 
		w_17830 , w_17831 , w_17832 , w_17833 , w_17834 , w_17835 , w_17836 , w_17837 , w_17838 , w_17839 , 
		w_17840 , w_17841 , w_17842 , w_17843 , w_17844 , w_17845 , w_17846 , w_17847 , w_17848 , w_17849 , 
		w_17850 , w_17851 , w_17852 , w_17853 , w_17854 , w_17855 , w_17856 , w_17857 , w_17858 , w_17859 , 
		w_17860 , w_17861 , w_17862 , w_17863 , w_17864 , w_17865 , w_17866 , w_17867 , w_17868 , w_17869 , 
		w_17870 , w_17871 , w_17872 , w_17873 , w_17874 , w_17875 , w_17876 , w_17877 , w_17878 , w_17879 , 
		w_17880 , w_17881 , w_17882 , w_17883 , w_17884 , w_17885 , w_17886 , w_17887 , w_17888 , w_17889 , 
		w_17890 , w_17891 , w_17892 , w_17893 , w_17894 , w_17895 , w_17896 , w_17897 , w_17898 , w_17899 , 
		w_17900 , w_17901 , w_17902 , w_17903 , w_17904 , w_17905 , w_17906 , w_17907 , w_17908 , w_17909 , 
		w_17910 , w_17911 , w_17912 , w_17913 , w_17914 , w_17915 , w_17916 , w_17917 , w_17918 , w_17919 , 
		w_17920 , w_17921 , w_17922 , w_17923 , w_17924 , w_17925 , w_17926 , w_17927 , w_17928 , w_17929 , 
		w_17930 , w_17931 , w_17932 , w_17933 , w_17934 , w_17935 , w_17936 , w_17937 , w_17938 , w_17939 , 
		w_17940 , w_17941 , w_17942 , w_17943 , w_17944 , w_17945 , w_17946 , w_17947 , w_17948 , w_17949 , 
		w_17950 , w_17951 , w_17952 , w_17953 , w_17954 , w_17955 , w_17956 , w_17957 , w_17958 , w_17959 , 
		w_17960 , w_17961 , w_17962 , w_17963 , w_17964 , w_17965 , w_17966 , w_17967 , w_17968 , w_17969 , 
		w_17970 , w_17971 , w_17972 , w_17973 , w_17974 , w_17975 , w_17976 , w_17977 , w_17978 , w_17979 , 
		w_17980 , w_17981 , w_17982 , w_17983 , w_17984 , w_17985 , w_17986 , w_17987 , w_17988 , w_17989 , 
		w_17990 , w_17991 , w_17992 , w_17993 , w_17994 , w_17995 , w_17996 , w_17997 , w_17998 , w_17999 , 
		w_18000 , w_18001 , w_18002 , w_18003 , w_18004 , w_18005 , w_18006 , w_18007 , w_18008 , w_18009 , 
		w_18010 , w_18011 , w_18012 , w_18013 , w_18014 , w_18015 , w_18016 , w_18017 , w_18018 , w_18019 , 
		w_18020 , w_18021 , w_18022 , w_18023 , w_18024 , w_18025 , w_18026 , w_18027 , w_18028 , w_18029 , 
		w_18030 , w_18031 , w_18032 , w_18033 , w_18034 , w_18035 , w_18036 , w_18037 , w_18038 , w_18039 , 
		w_18040 , w_18041 , w_18042 , w_18043 , w_18044 , w_18045 , w_18046 , w_18047 , w_18048 , w_18049 , 
		w_18050 , w_18051 , w_18052 , w_18053 , w_18054 , w_18055 , w_18056 , w_18057 , w_18058 , w_18059 , 
		w_18060 , w_18061 , w_18062 , w_18063 , w_18064 , w_18065 , w_18066 , w_18067 , w_18068 , w_18069 , 
		w_18070 , w_18071 , w_18072 , w_18073 , w_18074 , w_18075 , w_18076 , w_18077 , w_18078 , w_18079 , 
		w_18080 , w_18081 , w_18082 , w_18083 , w_18084 , w_18085 , w_18086 , w_18087 , w_18088 , w_18089 , 
		w_18090 , w_18091 , w_18092 , w_18093 , w_18094 , w_18095 , w_18096 , w_18097 , w_18098 , w_18099 , 
		w_18100 , w_18101 , w_18102 , w_18103 , w_18104 , w_18105 , w_18106 , w_18107 , w_18108 , w_18109 , 
		w_18110 , w_18111 , w_18112 , w_18113 , w_18114 , w_18115 , w_18116 , w_18117 , w_18118 , w_18119 , 
		w_18120 , w_18121 , w_18122 , w_18123 , w_18124 , w_18125 , w_18126 , w_18127 , w_18128 , w_18129 , 
		w_18130 , w_18131 , w_18132 , w_18133 , w_18134 , w_18135 , w_18136 , w_18137 , w_18138 , w_18139 , 
		w_18140 , w_18141 , w_18142 , w_18143 , w_18144 , w_18145 , w_18146 , w_18147 , w_18148 , w_18149 , 
		w_18150 , w_18151 , w_18152 , w_18153 , w_18154 , w_18155 , w_18156 , w_18157 , w_18158 , w_18159 , 
		w_18160 , w_18161 , w_18162 , w_18163 , w_18164 , w_18165 , w_18166 , w_18167 , w_18168 , w_18169 , 
		w_18170 , w_18171 , w_18172 , w_18173 , w_18174 , w_18175 , w_18176 , w_18177 , w_18178 , w_18179 , 
		w_18180 , w_18181 , w_18182 , w_18183 , w_18184 , w_18185 , w_18186 , w_18187 , w_18188 , w_18189 , 
		w_18190 , w_18191 , w_18192 , w_18193 , w_18194 , w_18195 , w_18196 , w_18197 , w_18198 , w_18199 , 
		w_18200 , w_18201 , w_18202 , w_18203 , w_18204 , w_18205 , w_18206 , w_18207 , w_18208 , w_18209 , 
		w_18210 , w_18211 , w_18212 , w_18213 , w_18214 , w_18215 , w_18216 , w_18217 , w_18218 , w_18219 , 
		w_18220 , w_18221 , w_18222 , w_18223 , w_18224 , w_18225 , w_18226 , w_18227 , w_18228 , w_18229 , 
		w_18230 , w_18231 , w_18232 , w_18233 , w_18234 , w_18235 , w_18236 , w_18237 , w_18238 , w_18239 , 
		w_18240 , w_18241 , w_18242 , w_18243 , w_18244 , w_18245 , w_18246 , w_18247 , w_18248 , w_18249 , 
		w_18250 , w_18251 , w_18252 , w_18253 , w_18254 , w_18255 , w_18256 , w_18257 , w_18258 , w_18259 , 
		w_18260 , w_18261 , w_18262 , w_18263 , w_18264 , w_18265 , w_18266 , w_18267 , w_18268 , w_18269 , 
		w_18270 , w_18271 , w_18272 , w_18273 , w_18274 , w_18275 , w_18276 , w_18277 , w_18278 , w_18279 , 
		w_18280 , w_18281 , w_18282 , w_18283 , w_18284 , w_18285 , w_18286 , w_18287 , w_18288 , w_18289 , 
		w_18290 , w_18291 , w_18292 , w_18293 , w_18294 , w_18295 , w_18296 , w_18297 , w_18298 , w_18299 , 
		w_18300 , w_18301 , w_18302 , w_18303 , w_18304 , w_18305 , w_18306 , w_18307 , w_18308 , w_18309 , 
		w_18310 , w_18311 , w_18312 , w_18313 , w_18314 , w_18315 , w_18316 , w_18317 , w_18318 , w_18319 , 
		w_18320 , w_18321 , w_18322 , w_18323 , w_18324 , w_18325 , w_18326 , w_18327 , w_18328 , w_18329 , 
		w_18330 , w_18331 , w_18332 , w_18333 , w_18334 , w_18335 , w_18336 , w_18337 , w_18338 , w_18339 , 
		w_18340 , w_18341 , w_18342 , w_18343 , w_18344 , w_18345 , w_18346 , w_18347 , w_18348 , w_18349 , 
		w_18350 , w_18351 , w_18352 , w_18353 , w_18354 , w_18355 , w_18356 , w_18357 , w_18358 , w_18359 , 
		w_18360 , w_18361 , w_18362 , w_18363 , w_18364 , w_18365 , w_18366 , w_18367 , w_18368 , w_18369 , 
		w_18370 , w_18371 , w_18372 , w_18373 , w_18374 , w_18375 , w_18376 , w_18377 , w_18378 , w_18379 , 
		w_18380 , w_18381 , w_18382 , w_18383 , w_18384 , w_18385 , w_18386 , w_18387 , w_18388 , w_18389 , 
		w_18390 , w_18391 , w_18392 , w_18393 , w_18394 , w_18395 , w_18396 , w_18397 , w_18398 , w_18399 , 
		w_18400 , w_18401 , w_18402 , w_18403 , w_18404 , w_18405 , w_18406 , w_18407 , w_18408 , w_18409 , 
		w_18410 , w_18411 , w_18412 , w_18413 , w_18414 , w_18415 , w_18416 , w_18417 , w_18418 , w_18419 , 
		w_18420 , w_18421 , w_18422 , w_18423 , w_18424 , w_18425 , w_18426 , w_18427 , w_18428 , w_18429 , 
		w_18430 , w_18431 , w_18432 , w_18433 , w_18434 , w_18435 , w_18436 , w_18437 , w_18438 , w_18439 , 
		w_18440 , w_18441 , w_18442 , w_18443 , w_18444 , w_18445 , w_18446 , w_18447 , w_18448 , w_18449 , 
		w_18450 , w_18451 , w_18452 , w_18453 , w_18454 , w_18455 , w_18456 , w_18457 , w_18458 , w_18459 , 
		w_18460 , w_18461 , w_18462 , w_18463 , w_18464 , w_18465 , w_18466 , w_18467 , w_18468 , w_18469 , 
		w_18470 , w_18471 , w_18472 , w_18473 , w_18474 , w_18475 , w_18476 , w_18477 , w_18478 , w_18479 , 
		w_18480 , w_18481 , w_18482 , w_18483 , w_18484 , w_18485 , w_18486 , w_18487 , w_18488 , w_18489 , 
		w_18490 , w_18491 , w_18492 , w_18493 , w_18494 , w_18495 , w_18496 , w_18497 , w_18498 , w_18499 , 
		w_18500 , w_18501 , w_18502 , w_18503 , w_18504 , w_18505 , w_18506 , w_18507 , w_18508 , w_18509 , 
		w_18510 , w_18511 , w_18512 , w_18513 , w_18514 , w_18515 , w_18516 , w_18517 , w_18518 , w_18519 , 
		w_18520 , w_18521 , w_18522 , w_18523 , w_18524 , w_18525 , w_18526 , w_18527 , w_18528 , w_18529 , 
		w_18530 , w_18531 , w_18532 , w_18533 , w_18534 , w_18535 , w_18536 , w_18537 , w_18538 , w_18539 , 
		w_18540 , w_18541 , w_18542 , w_18543 , w_18544 , w_18545 , w_18546 , w_18547 , w_18548 , w_18549 , 
		w_18550 , w_18551 , w_18552 , w_18553 , w_18554 , w_18555 , w_18556 , w_18557 , w_18558 , w_18559 , 
		w_18560 , w_18561 , w_18562 , w_18563 , w_18564 , w_18565 , w_18566 , w_18567 , w_18568 , w_18569 , 
		w_18570 , w_18571 , w_18572 , w_18573 , w_18574 , w_18575 , w_18576 , w_18577 , w_18578 , w_18579 , 
		w_18580 , w_18581 , w_18582 , w_18583 , w_18584 , w_18585 , w_18586 , w_18587 , w_18588 , w_18589 , 
		w_18590 , w_18591 , w_18592 , w_18593 , w_18594 , w_18595 , w_18596 , w_18597 , w_18598 , w_18599 , 
		w_18600 , w_18601 , w_18602 , w_18603 , w_18604 , w_18605 , w_18606 , w_18607 , w_18608 , w_18609 , 
		w_18610 , w_18611 , w_18612 , w_18613 , w_18614 , w_18615 , w_18616 , w_18617 , w_18618 , w_18619 , 
		w_18620 , w_18621 , w_18622 , w_18623 , w_18624 , w_18625 , w_18626 , w_18627 , w_18628 , w_18629 , 
		w_18630 , w_18631 , w_18632 , w_18633 , w_18634 , w_18635 , w_18636 , w_18637 , w_18638 , w_18639 , 
		w_18640 , w_18641 , w_18642 , w_18643 , w_18644 , w_18645 , w_18646 , w_18647 , w_18648 , w_18649 , 
		w_18650 , w_18651 , w_18652 , w_18653 , w_18654 , w_18655 , w_18656 , w_18657 , w_18658 , w_18659 , 
		w_18660 , w_18661 , w_18662 , w_18663 , w_18664 , w_18665 , w_18666 , w_18667 , w_18668 , w_18669 , 
		w_18670 , w_18671 , w_18672 , w_18673 , w_18674 , w_18675 , w_18676 , w_18677 , w_18678 , w_18679 , 
		w_18680 , w_18681 , w_18682 , w_18683 , w_18684 , w_18685 , w_18686 , w_18687 , w_18688 , w_18689 , 
		w_18690 , w_18691 , w_18692 , w_18693 , w_18694 , w_18695 , w_18696 , w_18697 , w_18698 , w_18699 , 
		w_18700 , w_18701 , w_18702 , w_18703 , w_18704 , w_18705 , w_18706 , w_18707 , w_18708 , w_18709 , 
		w_18710 , w_18711 , w_18712 , w_18713 , w_18714 , w_18715 , w_18716 , w_18717 , w_18718 , w_18719 , 
		w_18720 , w_18721 , w_18722 , w_18723 , w_18724 , w_18725 , w_18726 , w_18727 , w_18728 , w_18729 , 
		w_18730 , w_18731 , w_18732 , w_18733 , w_18734 , w_18735 , w_18736 , w_18737 , w_18738 , w_18739 , 
		w_18740 , w_18741 , w_18742 , w_18743 , w_18744 , w_18745 , w_18746 , w_18747 , w_18748 , w_18749 , 
		w_18750 , w_18751 , w_18752 , w_18753 , w_18754 , w_18755 , w_18756 , w_18757 , w_18758 , w_18759 , 
		w_18760 , w_18761 , w_18762 , w_18763 , w_18764 , w_18765 , w_18766 , w_18767 , w_18768 , w_18769 , 
		w_18770 , w_18771 , w_18772 , w_18773 , w_18774 , w_18775 , w_18776 , w_18777 , w_18778 , w_18779 , 
		w_18780 , w_18781 , w_18782 , w_18783 , w_18784 , w_18785 , w_18786 , w_18787 , w_18788 , w_18789 , 
		w_18790 , w_18791 , w_18792 , w_18793 , w_18794 , w_18795 , w_18796 , w_18797 , w_18798 , w_18799 , 
		w_18800 , w_18801 , w_18802 , w_18803 , w_18804 , w_18805 , w_18806 , w_18807 , w_18808 , w_18809 , 
		w_18810 , w_18811 , w_18812 , w_18813 , w_18814 , w_18815 , w_18816 , w_18817 , w_18818 , w_18819 , 
		w_18820 , w_18821 , w_18822 , w_18823 , w_18824 , w_18825 , w_18826 , w_18827 , w_18828 , w_18829 , 
		w_18830 , w_18831 , w_18832 , w_18833 , w_18834 , w_18835 , w_18836 , w_18837 , w_18838 , w_18839 , 
		w_18840 , w_18841 , w_18842 , w_18843 , w_18844 , w_18845 , w_18846 , w_18847 , w_18848 , w_18849 , 
		w_18850 , w_18851 , w_18852 , w_18853 , w_18854 , w_18855 , w_18856 , w_18857 , w_18858 , w_18859 , 
		w_18860 , w_18861 , w_18862 , w_18863 , w_18864 , w_18865 , w_18866 , w_18867 , w_18868 , w_18869 , 
		w_18870 , w_18871 , w_18872 , w_18873 , w_18874 , w_18875 , w_18876 , w_18877 , w_18878 , w_18879 , 
		w_18880 , w_18881 , w_18882 , w_18883 , w_18884 , w_18885 , w_18886 , w_18887 , w_18888 , w_18889 , 
		w_18890 , w_18891 , w_18892 , w_18893 , w_18894 , w_18895 , w_18896 , w_18897 , w_18898 , w_18899 , 
		w_18900 , w_18901 , w_18902 , w_18903 , w_18904 , w_18905 , w_18906 , w_18907 , w_18908 , w_18909 , 
		w_18910 , w_18911 , w_18912 , w_18913 , w_18914 , w_18915 , w_18916 , w_18917 , w_18918 , w_18919 , 
		w_18920 , w_18921 , w_18922 , w_18923 , w_18924 , w_18925 , w_18926 , w_18927 , w_18928 , w_18929 , 
		w_18930 , w_18931 , w_18932 , w_18933 , w_18934 , w_18935 , w_18936 , w_18937 , w_18938 , w_18939 , 
		w_18940 , w_18941 , w_18942 , w_18943 , w_18944 , w_18945 , w_18946 , w_18947 , w_18948 , w_18949 , 
		w_18950 , w_18951 , w_18952 , w_18953 , w_18954 , w_18955 , w_18956 , w_18957 , w_18958 , w_18959 , 
		w_18960 , w_18961 , w_18962 , w_18963 , w_18964 , w_18965 , w_18966 , w_18967 , w_18968 , w_18969 , 
		w_18970 , w_18971 , w_18972 , w_18973 , w_18974 , w_18975 , w_18976 , w_18977 , w_18978 , w_18979 , 
		w_18980 , w_18981 , w_18982 , w_18983 , w_18984 , w_18985 , w_18986 , w_18987 , w_18988 , w_18989 , 
		w_18990 , w_18991 , w_18992 , w_18993 , w_18994 , w_18995 , w_18996 , w_18997 , w_18998 , w_18999 , 
		w_19000 , w_19001 , w_19002 , w_19003 , w_19004 , w_19005 , w_19006 , w_19007 , w_19008 , w_19009 , 
		w_19010 , w_19011 , w_19012 , w_19013 , w_19014 , w_19015 , w_19016 , w_19017 , w_19018 , w_19019 , 
		w_19020 , w_19021 , w_19022 , w_19023 , w_19024 , w_19025 , w_19026 , w_19027 , w_19028 , w_19029 , 
		w_19030 , w_19031 , w_19032 , w_19033 , w_19034 , w_19035 , w_19036 , w_19037 , w_19038 , w_19039 , 
		w_19040 , w_19041 , w_19042 , w_19043 , w_19044 , w_19045 , w_19046 , w_19047 , w_19048 , w_19049 , 
		w_19050 , w_19051 , w_19052 , w_19053 , w_19054 , w_19055 , w_19056 , w_19057 , w_19058 , w_19059 , 
		w_19060 , w_19061 , w_19062 , w_19063 , w_19064 , w_19065 , w_19066 , w_19067 , w_19068 , w_19069 , 
		w_19070 , w_19071 , w_19072 , w_19073 , w_19074 , w_19075 , w_19076 , w_19077 , w_19078 , w_19079 , 
		w_19080 , w_19081 , w_19082 , w_19083 , w_19084 , w_19085 , w_19086 , w_19087 , w_19088 , w_19089 , 
		w_19090 , w_19091 , w_19092 , w_19093 , w_19094 , w_19095 , w_19096 , w_19097 , w_19098 , w_19099 , 
		w_19100 , w_19101 , w_19102 , w_19103 , w_19104 , w_19105 , w_19106 , w_19107 , w_19108 , w_19109 , 
		w_19110 , w_19111 , w_19112 , w_19113 , w_19114 , w_19115 , w_19116 , w_19117 , w_19118 , w_19119 , 
		w_19120 , w_19121 , w_19122 , w_19123 , w_19124 , w_19125 , w_19126 , w_19127 , w_19128 , w_19129 , 
		w_19130 , w_19131 , w_19132 , w_19133 , w_19134 , w_19135 , w_19136 , w_19137 , w_19138 , w_19139 , 
		w_19140 , w_19141 , w_19142 , w_19143 , w_19144 , w_19145 , w_19146 , w_19147 , w_19148 , w_19149 , 
		w_19150 , w_19151 , w_19152 , w_19153 , w_19154 , w_19155 , w_19156 , w_19157 , w_19158 , w_19159 , 
		w_19160 , w_19161 , w_19162 , w_19163 , w_19164 , w_19165 , w_19166 , w_19167 , w_19168 , w_19169 , 
		w_19170 , w_19171 , w_19172 , w_19173 , w_19174 , w_19175 , w_19176 , w_19177 , w_19178 , w_19179 , 
		w_19180 , w_19181 , w_19182 , w_19183 , w_19184 , w_19185 , w_19186 , w_19187 , w_19188 , w_19189 , 
		w_19190 , w_19191 , w_19192 , w_19193 , w_19194 , w_19195 , w_19196 , w_19197 , w_19198 , w_19199 , 
		w_19200 , w_19201 , w_19202 , w_19203 , w_19204 , w_19205 , w_19206 , w_19207 , w_19208 , w_19209 , 
		w_19210 , w_19211 , w_19212 , w_19213 , w_19214 , w_19215 , w_19216 , w_19217 , w_19218 , w_19219 , 
		w_19220 , w_19221 , w_19222 , w_19223 , w_19224 , w_19225 , w_19226 , w_19227 , w_19228 , w_19229 , 
		w_19230 , w_19231 , w_19232 , w_19233 , w_19234 , w_19235 , w_19236 , w_19237 , w_19238 , w_19239 , 
		w_19240 , w_19241 , w_19242 , w_19243 , w_19244 , w_19245 , w_19246 , w_19247 , w_19248 , w_19249 , 
		w_19250 , w_19251 , w_19252 , w_19253 , w_19254 , w_19255 , w_19256 , w_19257 , w_19258 , w_19259 , 
		w_19260 , w_19261 , w_19262 , w_19263 , w_19264 , w_19265 , w_19266 , w_19267 , w_19268 , w_19269 , 
		w_19270 , w_19271 , w_19272 , w_19273 , w_19274 , w_19275 , w_19276 , w_19277 , w_19278 , w_19279 , 
		w_19280 , w_19281 , w_19282 , w_19283 , w_19284 , w_19285 , w_19286 , w_19287 , w_19288 , w_19289 , 
		w_19290 , w_19291 , w_19292 , w_19293 , w_19294 , w_19295 , w_19296 , w_19297 , w_19298 , w_19299 , 
		w_19300 , w_19301 , w_19302 , w_19303 , w_19304 , w_19305 , w_19306 , w_19307 , w_19308 , w_19309 , 
		w_19310 , w_19311 , w_19312 , w_19313 , w_19314 , w_19315 , w_19316 , w_19317 , w_19318 , w_19319 , 
		w_19320 , w_19321 , w_19322 , w_19323 , w_19324 , w_19325 , w_19326 , w_19327 , w_19328 , w_19329 , 
		w_19330 , w_19331 , w_19332 , w_19333 , w_19334 , w_19335 , w_19336 , w_19337 , w_19338 , w_19339 , 
		w_19340 , w_19341 , w_19342 , w_19343 , w_19344 , w_19345 , w_19346 , w_19347 , w_19348 , w_19349 , 
		w_19350 , w_19351 , w_19352 , w_19353 , w_19354 , w_19355 , w_19356 , w_19357 , w_19358 , w_19359 , 
		w_19360 , w_19361 , w_19362 , w_19363 , w_19364 , w_19365 , w_19366 , w_19367 , w_19368 , w_19369 , 
		w_19370 , w_19371 , w_19372 , w_19373 , w_19374 , w_19375 , w_19376 , w_19377 , w_19378 , w_19379 , 
		w_19380 , w_19381 , w_19382 , w_19383 , w_19384 , w_19385 , w_19386 , w_19387 , w_19388 , w_19389 , 
		w_19390 , w_19391 , w_19392 , w_19393 , w_19394 , w_19395 , w_19396 , w_19397 , w_19398 , w_19399 , 
		w_19400 , w_19401 , w_19402 , w_19403 , w_19404 , w_19405 , w_19406 , w_19407 , w_19408 , w_19409 , 
		w_19410 , w_19411 , w_19412 , w_19413 , w_19414 , w_19415 , w_19416 , w_19417 , w_19418 , w_19419 , 
		w_19420 , w_19421 , w_19422 , w_19423 , w_19424 , w_19425 , w_19426 , w_19427 , w_19428 , w_19429 , 
		w_19430 , w_19431 , w_19432 , w_19433 , w_19434 , w_19435 , w_19436 , w_19437 , w_19438 , w_19439 , 
		w_19440 , w_19441 , w_19442 , w_19443 , w_19444 , w_19445 , w_19446 , w_19447 , w_19448 , w_19449 , 
		w_19450 , w_19451 , w_19452 , w_19453 , w_19454 , w_19455 , w_19456 , w_19457 , w_19458 , w_19459 , 
		w_19460 , w_19461 , w_19462 , w_19463 , w_19464 , w_19465 , w_19466 , w_19467 , w_19468 , w_19469 , 
		w_19470 , w_19471 , w_19472 , w_19473 , w_19474 , w_19475 , w_19476 , w_19477 , w_19478 , w_19479 , 
		w_19480 , w_19481 , w_19482 , w_19483 , w_19484 , w_19485 , w_19486 , w_19487 , w_19488 , w_19489 , 
		w_19490 , w_19491 , w_19492 , w_19493 , w_19494 , w_19495 , w_19496 , w_19497 , w_19498 , w_19499 , 
		w_19500 , w_19501 , w_19502 , w_19503 , w_19504 , w_19505 , w_19506 , w_19507 , w_19508 , w_19509 , 
		w_19510 , w_19511 , w_19512 , w_19513 , w_19514 , w_19515 , w_19516 , w_19517 , w_19518 , w_19519 , 
		w_19520 , w_19521 , w_19522 , w_19523 , w_19524 , w_19525 , w_19526 , w_19527 , w_19528 , w_19529 , 
		w_19530 , w_19531 , w_19532 , w_19533 , w_19534 , w_19535 , w_19536 , w_19537 , w_19538 , w_19539 , 
		w_19540 , w_19541 , w_19542 , w_19543 , w_19544 , w_19545 , w_19546 , w_19547 , w_19548 , w_19549 , 
		w_19550 , w_19551 , w_19552 , w_19553 , w_19554 , w_19555 , w_19556 , w_19557 , w_19558 , w_19559 , 
		w_19560 , w_19561 , w_19562 , w_19563 , w_19564 , w_19565 , w_19566 , w_19567 , w_19568 , w_19569 , 
		w_19570 , w_19571 , w_19572 , w_19573 , w_19574 , w_19575 , w_19576 , w_19577 , w_19578 , w_19579 , 
		w_19580 , w_19581 , w_19582 , w_19583 , w_19584 , w_19585 , w_19586 , w_19587 , w_19588 , w_19589 , 
		w_19590 , w_19591 , w_19592 , w_19593 , w_19594 , w_19595 , w_19596 , w_19597 , w_19598 , w_19599 , 
		w_19600 , w_19601 , w_19602 , w_19603 , w_19604 , w_19605 , w_19606 , w_19607 , w_19608 , w_19609 , 
		w_19610 , w_19611 , w_19612 , w_19613 , w_19614 , w_19615 , w_19616 , w_19617 , w_19618 , w_19619 , 
		w_19620 , w_19621 , w_19622 , w_19623 , w_19624 , w_19625 , w_19626 , w_19627 , w_19628 , w_19629 , 
		w_19630 , w_19631 , w_19632 , w_19633 , w_19634 , w_19635 , w_19636 , w_19637 , w_19638 , w_19639 , 
		w_19640 , w_19641 , w_19642 , w_19643 , w_19644 , w_19645 , w_19646 , w_19647 , w_19648 , w_19649 , 
		w_19650 , w_19651 , w_19652 , w_19653 , w_19654 , w_19655 , w_19656 , w_19657 , w_19658 , w_19659 , 
		w_19660 , w_19661 , w_19662 , w_19663 , w_19664 , w_19665 , w_19666 , w_19667 , w_19668 , w_19669 , 
		w_19670 , w_19671 , w_19672 , w_19673 , w_19674 , w_19675 , w_19676 , w_19677 , w_19678 , w_19679 , 
		w_19680 , w_19681 , w_19682 , w_19683 , w_19684 , w_19685 , w_19686 , w_19687 , w_19688 , w_19689 , 
		w_19690 , w_19691 , w_19692 , w_19693 , w_19694 , w_19695 , w_19696 , w_19697 , w_19698 , w_19699 , 
		w_19700 , w_19701 , w_19702 , w_19703 , w_19704 , w_19705 , w_19706 , w_19707 , w_19708 , w_19709 , 
		w_19710 , w_19711 , w_19712 , w_19713 , w_19714 , w_19715 , w_19716 , w_19717 , w_19718 , w_19719 , 
		w_19720 , w_19721 , w_19722 , w_19723 , w_19724 , w_19725 , w_19726 , w_19727 , w_19728 , w_19729 , 
		w_19730 , w_19731 , w_19732 , w_19733 , w_19734 , w_19735 , w_19736 , w_19737 , w_19738 , w_19739 , 
		w_19740 , w_19741 , w_19742 , w_19743 , w_19744 , w_19745 , w_19746 , w_19747 , w_19748 , w_19749 , 
		w_19750 , w_19751 , w_19752 , w_19753 , w_19754 , w_19755 , w_19756 , w_19757 , w_19758 , w_19759 , 
		w_19760 , w_19761 , w_19762 , w_19763 , w_19764 , w_19765 , w_19766 , w_19767 , w_19768 , w_19769 , 
		w_19770 , w_19771 , w_19772 , w_19773 , w_19774 , w_19775 , w_19776 , w_19777 , w_19778 , w_19779 , 
		w_19780 , w_19781 , w_19782 , w_19783 , w_19784 , w_19785 , w_19786 , w_19787 , w_19788 , w_19789 , 
		w_19790 , w_19791 , w_19792 , w_19793 , w_19794 , w_19795 , w_19796 , w_19797 , w_19798 , w_19799 , 
		w_19800 , w_19801 , w_19802 , w_19803 , w_19804 , w_19805 , w_19806 , w_19807 , w_19808 , w_19809 , 
		w_19810 , w_19811 , w_19812 , w_19813 , w_19814 , w_19815 , w_19816 , w_19817 , w_19818 , w_19819 , 
		w_19820 , w_19821 , w_19822 , w_19823 , w_19824 , w_19825 , w_19826 , w_19827 , w_19828 , w_19829 , 
		w_19830 , w_19831 , w_19832 , w_19833 , w_19834 , w_19835 , w_19836 , w_19837 , w_19838 , w_19839 , 
		w_19840 , w_19841 , w_19842 , w_19843 , w_19844 , w_19845 , w_19846 , w_19847 , w_19848 , w_19849 , 
		w_19850 , w_19851 , w_19852 , w_19853 , w_19854 , w_19855 , w_19856 , w_19857 , w_19858 , w_19859 , 
		w_19860 , w_19861 , w_19862 , w_19863 , w_19864 , w_19865 , w_19866 , w_19867 , w_19868 , w_19869 , 
		w_19870 , w_19871 , w_19872 , w_19873 , w_19874 , w_19875 , w_19876 , w_19877 , w_19878 , w_19879 , 
		w_19880 , w_19881 , w_19882 , w_19883 , w_19884 , w_19885 , w_19886 , w_19887 , w_19888 , w_19889 , 
		w_19890 , w_19891 , w_19892 , w_19893 , w_19894 , w_19895 , w_19896 , w_19897 , w_19898 , w_19899 , 
		w_19900 , w_19901 , w_19902 , w_19903 , w_19904 , w_19905 , w_19906 , w_19907 , w_19908 , w_19909 , 
		w_19910 , w_19911 , w_19912 , w_19913 , w_19914 , w_19915 , w_19916 , w_19917 , w_19918 , w_19919 , 
		w_19920 , w_19921 , w_19922 , w_19923 , w_19924 , w_19925 , w_19926 , w_19927 , w_19928 , w_19929 , 
		w_19930 , w_19931 , w_19932 , w_19933 , w_19934 , w_19935 , w_19936 , w_19937 , w_19938 , w_19939 , 
		w_19940 , w_19941 , w_19942 , w_19943 , w_19944 , w_19945 , w_19946 , w_19947 , w_19948 , w_19949 , 
		w_19950 , w_19951 , w_19952 , w_19953 , w_19954 , w_19955 , w_19956 , w_19957 , w_19958 , w_19959 , 
		w_19960 , w_19961 , w_19962 , w_19963 , w_19964 , w_19965 , w_19966 , w_19967 , w_19968 , w_19969 , 
		w_19970 , w_19971 , w_19972 , w_19973 , w_19974 , w_19975 , w_19976 , w_19977 , w_19978 , w_19979 , 
		w_19980 , w_19981 , w_19982 , w_19983 , w_19984 , w_19985 , w_19986 , w_19987 , w_19988 , w_19989 , 
		w_19990 , w_19991 , w_19992 , w_19993 , w_19994 , w_19995 , w_19996 , w_19997 , w_19998 , w_19999 , 
		w_20000 , w_20001 , w_20002 , w_20003 , w_20004 , w_20005 , w_20006 , w_20007 , w_20008 , w_20009 , 
		w_20010 , w_20011 , w_20012 , w_20013 , w_20014 , w_20015 , w_20016 , w_20017 , w_20018 , w_20019 , 
		w_20020 , w_20021 , w_20022 , w_20023 , w_20024 , w_20025 , w_20026 , w_20027 , w_20028 , w_20029 , 
		w_20030 , w_20031 , w_20032 , w_20033 , w_20034 , w_20035 , w_20036 , w_20037 , w_20038 , w_20039 , 
		w_20040 , w_20041 , w_20042 , w_20043 , w_20044 , w_20045 , w_20046 , w_20047 , w_20048 , w_20049 , 
		w_20050 , w_20051 , w_20052 , w_20053 , w_20054 , w_20055 , w_20056 , w_20057 , w_20058 , w_20059 , 
		w_20060 , w_20061 , w_20062 , w_20063 , w_20064 , w_20065 , w_20066 , w_20067 , w_20068 , w_20069 , 
		w_20070 , w_20071 , w_20072 , w_20073 , w_20074 , w_20075 , w_20076 , w_20077 , w_20078 , w_20079 , 
		w_20080 , w_20081 , w_20082 , w_20083 , w_20084 , w_20085 , w_20086 , w_20087 , w_20088 , w_20089 , 
		w_20090 , w_20091 , w_20092 , w_20093 , w_20094 , w_20095 , w_20096 , w_20097 , w_20098 , w_20099 , 
		w_20100 , w_20101 , w_20102 , w_20103 , w_20104 , w_20105 , w_20106 , w_20107 , w_20108 , w_20109 , 
		w_20110 , w_20111 , w_20112 , w_20113 , w_20114 , w_20115 , w_20116 , w_20117 , w_20118 , w_20119 , 
		w_20120 , w_20121 , w_20122 , w_20123 , w_20124 , w_20125 , w_20126 , w_20127 , w_20128 , w_20129 , 
		w_20130 , w_20131 , w_20132 , w_20133 , w_20134 , w_20135 , w_20136 , w_20137 , w_20138 , w_20139 , 
		w_20140 , w_20141 , w_20142 , w_20143 , w_20144 , w_20145 , w_20146 , w_20147 , w_20148 , w_20149 , 
		w_20150 , w_20151 , w_20152 , w_20153 , w_20154 , w_20155 , w_20156 , w_20157 , w_20158 , w_20159 , 
		w_20160 , w_20161 , w_20162 , w_20163 , w_20164 , w_20165 , w_20166 , w_20167 , w_20168 , w_20169 , 
		w_20170 , w_20171 , w_20172 , w_20173 , w_20174 , w_20175 , w_20176 , w_20177 , w_20178 , w_20179 , 
		w_20180 , w_20181 , w_20182 , w_20183 , w_20184 , w_20185 , w_20186 , w_20187 , w_20188 , w_20189 , 
		w_20190 , w_20191 , w_20192 , w_20193 , w_20194 , w_20195 , w_20196 , w_20197 , w_20198 , w_20199 , 
		w_20200 , w_20201 , w_20202 , w_20203 , w_20204 , w_20205 , w_20206 , w_20207 , w_20208 , w_20209 , 
		w_20210 , w_20211 , w_20212 , w_20213 , w_20214 , w_20215 , w_20216 , w_20217 , w_20218 , w_20219 , 
		w_20220 , w_20221 , w_20222 , w_20223 , w_20224 , w_20225 , w_20226 , w_20227 , w_20228 , w_20229 , 
		w_20230 , w_20231 , w_20232 , w_20233 , w_20234 , w_20235 , w_20236 , w_20237 , w_20238 , w_20239 , 
		w_20240 , w_20241 , w_20242 , w_20243 , w_20244 , w_20245 , w_20246 , w_20247 , w_20248 , w_20249 , 
		w_20250 , w_20251 , w_20252 , w_20253 , w_20254 , w_20255 , w_20256 , w_20257 , w_20258 , w_20259 , 
		w_20260 , w_20261 , w_20262 , w_20263 , w_20264 , w_20265 , w_20266 , w_20267 , w_20268 , w_20269 , 
		w_20270 , w_20271 , w_20272 , w_20273 , w_20274 , w_20275 , w_20276 , w_20277 , w_20278 , w_20279 , 
		w_20280 , w_20281 , w_20282 , w_20283 , w_20284 , w_20285 , w_20286 , w_20287 , w_20288 , w_20289 , 
		w_20290 , w_20291 , w_20292 , w_20293 , w_20294 , w_20295 , w_20296 , w_20297 , w_20298 , w_20299 , 
		w_20300 , w_20301 , w_20302 , w_20303 , w_20304 , w_20305 , w_20306 , w_20307 , w_20308 , w_20309 , 
		w_20310 , w_20311 , w_20312 , w_20313 , w_20314 , w_20315 , w_20316 , w_20317 , w_20318 , w_20319 , 
		w_20320 , w_20321 , w_20322 , w_20323 , w_20324 , w_20325 , w_20326 , w_20327 , w_20328 , w_20329 , 
		w_20330 , w_20331 , w_20332 , w_20333 , w_20334 , w_20335 , w_20336 , w_20337 , w_20338 , w_20339 , 
		w_20340 , w_20341 , w_20342 , w_20343 , w_20344 , w_20345 , w_20346 , w_20347 , w_20348 , w_20349 , 
		w_20350 , w_20351 , w_20352 , w_20353 , w_20354 , w_20355 , w_20356 , w_20357 , w_20358 , w_20359 , 
		w_20360 , w_20361 , w_20362 , w_20363 , w_20364 , w_20365 , w_20366 , w_20367 , w_20368 , w_20369 , 
		w_20370 , w_20371 , w_20372 , w_20373 , w_20374 , w_20375 , w_20376 , w_20377 , w_20378 , w_20379 , 
		w_20380 , w_20381 , w_20382 , w_20383 , w_20384 , w_20385 , w_20386 , w_20387 , w_20388 , w_20389 , 
		w_20390 , w_20391 , w_20392 , w_20393 , w_20394 , w_20395 , w_20396 , w_20397 , w_20398 , w_20399 , 
		w_20400 , w_20401 , w_20402 , w_20403 , w_20404 , w_20405 , w_20406 , w_20407 , w_20408 , w_20409 , 
		w_20410 , w_20411 , w_20412 , w_20413 , w_20414 , w_20415 , w_20416 , w_20417 , w_20418 , w_20419 , 
		w_20420 , w_20421 , w_20422 , w_20423 , w_20424 , w_20425 , w_20426 , w_20427 , w_20428 , w_20429 , 
		w_20430 , w_20431 , w_20432 , w_20433 , w_20434 , w_20435 , w_20436 , w_20437 , w_20438 , w_20439 , 
		w_20440 , w_20441 , w_20442 , w_20443 , w_20444 , w_20445 , w_20446 , w_20447 , w_20448 , w_20449 , 
		w_20450 , w_20451 , w_20452 , w_20453 , w_20454 , w_20455 , w_20456 , w_20457 , w_20458 , w_20459 , 
		w_20460 , w_20461 , w_20462 , w_20463 , w_20464 , w_20465 , w_20466 , w_20467 , w_20468 , w_20469 , 
		w_20470 , w_20471 , w_20472 , w_20473 , w_20474 , w_20475 , w_20476 , w_20477 , w_20478 , w_20479 , 
		w_20480 , w_20481 , w_20482 , w_20483 , w_20484 , w_20485 , w_20486 , w_20487 , w_20488 , w_20489 , 
		w_20490 , w_20491 , w_20492 , w_20493 , w_20494 , w_20495 , w_20496 , w_20497 , w_20498 , w_20499 , 
		w_20500 , w_20501 , w_20502 , w_20503 , w_20504 , w_20505 , w_20506 , w_20507 , w_20508 , w_20509 , 
		w_20510 , w_20511 , w_20512 , w_20513 , w_20514 , w_20515 , w_20516 , w_20517 , w_20518 , w_20519 , 
		w_20520 , w_20521 , w_20522 , w_20523 , w_20524 , w_20525 , w_20526 , w_20527 , w_20528 , w_20529 , 
		w_20530 , w_20531 , w_20532 , w_20533 , w_20534 , w_20535 , w_20536 , w_20537 , w_20538 , w_20539 , 
		w_20540 , w_20541 , w_20542 , w_20543 , w_20544 , w_20545 , w_20546 , w_20547 , w_20548 , w_20549 , 
		w_20550 , w_20551 , w_20552 , w_20553 , w_20554 , w_20555 , w_20556 , w_20557 , w_20558 , w_20559 , 
		w_20560 , w_20561 , w_20562 , w_20563 , w_20564 , w_20565 , w_20566 , w_20567 , w_20568 , w_20569 , 
		w_20570 , w_20571 , w_20572 , w_20573 , w_20574 , w_20575 , w_20576 , w_20577 , w_20578 , w_20579 , 
		w_20580 , w_20581 , w_20582 , w_20583 , w_20584 , w_20585 , w_20586 , w_20587 , w_20588 , w_20589 , 
		w_20590 , w_20591 , w_20592 , w_20593 , w_20594 , w_20595 , w_20596 , w_20597 , w_20598 , w_20599 , 
		w_20600 , w_20601 , w_20602 , w_20603 , w_20604 , w_20605 , w_20606 , w_20607 , w_20608 , w_20609 , 
		w_20610 , w_20611 , w_20612 , w_20613 , w_20614 , w_20615 , w_20616 , w_20617 , w_20618 , w_20619 , 
		w_20620 , w_20621 , w_20622 , w_20623 , w_20624 , w_20625 , w_20626 , w_20627 , w_20628 , w_20629 , 
		w_20630 , w_20631 , w_20632 , w_20633 , w_20634 , w_20635 , w_20636 , w_20637 , w_20638 , w_20639 , 
		w_20640 , w_20641 , w_20642 , w_20643 , w_20644 , w_20645 , w_20646 , w_20647 , w_20648 , w_20649 , 
		w_20650 , w_20651 , w_20652 , w_20653 , w_20654 , w_20655 , w_20656 , w_20657 , w_20658 , w_20659 , 
		w_20660 , w_20661 , w_20662 , w_20663 , w_20664 , w_20665 , w_20666 , w_20667 , w_20668 , w_20669 , 
		w_20670 , w_20671 , w_20672 , w_20673 , w_20674 , w_20675 , w_20676 , w_20677 , w_20678 , w_20679 , 
		w_20680 , w_20681 , w_20682 , w_20683 , w_20684 , w_20685 , w_20686 , w_20687 , w_20688 , w_20689 , 
		w_20690 , w_20691 , w_20692 , w_20693 , w_20694 , w_20695 , w_20696 , w_20697 , w_20698 , w_20699 , 
		w_20700 , w_20701 , w_20702 , w_20703 , w_20704 , w_20705 , w_20706 , w_20707 , w_20708 , w_20709 , 
		w_20710 , w_20711 , w_20712 , w_20713 , w_20714 , w_20715 , w_20716 , w_20717 , w_20718 , w_20719 , 
		w_20720 , w_20721 , w_20722 , w_20723 , w_20724 , w_20725 , w_20726 , w_20727 , w_20728 , w_20729 , 
		w_20730 , w_20731 , w_20732 , w_20733 , w_20734 , w_20735 , w_20736 , w_20737 , w_20738 , w_20739 , 
		w_20740 , w_20741 , w_20742 , w_20743 , w_20744 , w_20745 , w_20746 , w_20747 , w_20748 , w_20749 , 
		w_20750 , w_20751 , w_20752 , w_20753 , w_20754 , w_20755 , w_20756 , w_20757 , w_20758 , w_20759 , 
		w_20760 , w_20761 , w_20762 , w_20763 , w_20764 , w_20765 , w_20766 , w_20767 , w_20768 , w_20769 , 
		w_20770 , w_20771 , w_20772 , w_20773 , w_20774 , w_20775 , w_20776 , w_20777 , w_20778 , w_20779 , 
		w_20780 , w_20781 , w_20782 , w_20783 , w_20784 , w_20785 , w_20786 , w_20787 , w_20788 , w_20789 , 
		w_20790 , w_20791 , w_20792 , w_20793 , w_20794 , w_20795 , w_20796 , w_20797 , w_20798 , w_20799 , 
		w_20800 , w_20801 , w_20802 , w_20803 , w_20804 , w_20805 , w_20806 , w_20807 , w_20808 , w_20809 , 
		w_20810 , w_20811 , w_20812 , w_20813 , w_20814 , w_20815 , w_20816 , w_20817 , w_20818 , w_20819 , 
		w_20820 , w_20821 , w_20822 , w_20823 , w_20824 , w_20825 , w_20826 , w_20827 , w_20828 , w_20829 , 
		w_20830 , w_20831 , w_20832 , w_20833 , w_20834 , w_20835 , w_20836 , w_20837 , w_20838 , w_20839 , 
		w_20840 , w_20841 , w_20842 , w_20843 , w_20844 , w_20845 , w_20846 , w_20847 , w_20848 , w_20849 , 
		w_20850 , w_20851 , w_20852 , w_20853 , w_20854 , w_20855 , w_20856 , w_20857 , w_20858 , w_20859 , 
		w_20860 , w_20861 , w_20862 , w_20863 , w_20864 , w_20865 , w_20866 , w_20867 , w_20868 , w_20869 , 
		w_20870 , w_20871 , w_20872 , w_20873 , w_20874 , w_20875 , w_20876 , w_20877 , w_20878 , w_20879 , 
		w_20880 , w_20881 , w_20882 , w_20883 , w_20884 , w_20885 , w_20886 , w_20887 , w_20888 , w_20889 , 
		w_20890 , w_20891 , w_20892 , w_20893 , w_20894 , w_20895 , w_20896 , w_20897 , w_20898 , w_20899 , 
		w_20900 , w_20901 , w_20902 , w_20903 , w_20904 , w_20905 , w_20906 , w_20907 , w_20908 , w_20909 , 
		w_20910 , w_20911 , w_20912 , w_20913 , w_20914 , w_20915 , w_20916 , w_20917 , w_20918 , w_20919 , 
		w_20920 , w_20921 , w_20922 , w_20923 , w_20924 , w_20925 , w_20926 , w_20927 , w_20928 , w_20929 , 
		w_20930 , w_20931 , w_20932 , w_20933 , w_20934 , w_20935 , w_20936 , w_20937 , w_20938 , w_20939 , 
		w_20940 , w_20941 , w_20942 , w_20943 , w_20944 , w_20945 , w_20946 , w_20947 , w_20948 , w_20949 , 
		w_20950 , w_20951 , w_20952 , w_20953 , w_20954 , w_20955 , w_20956 , w_20957 , w_20958 , w_20959 , 
		w_20960 , w_20961 , w_20962 , w_20963 , w_20964 , w_20965 , w_20966 , w_20967 , w_20968 , w_20969 , 
		w_20970 , w_20971 , w_20972 , w_20973 , w_20974 , w_20975 , w_20976 , w_20977 , w_20978 , w_20979 , 
		w_20980 , w_20981 , w_20982 , w_20983 , w_20984 , w_20985 , w_20986 , w_20987 , w_20988 , w_20989 , 
		w_20990 , w_20991 , w_20992 , w_20993 , w_20994 , w_20995 , w_20996 , w_20997 , w_20998 , w_20999 , 
		w_21000 , w_21001 , w_21002 , w_21003 , w_21004 , w_21005 , w_21006 , w_21007 , w_21008 , w_21009 , 
		w_21010 , w_21011 , w_21012 , w_21013 , w_21014 , w_21015 , w_21016 , w_21017 , w_21018 , w_21019 , 
		w_21020 , w_21021 , w_21022 , w_21023 , w_21024 , w_21025 , w_21026 , w_21027 , w_21028 , w_21029 , 
		w_21030 , w_21031 , w_21032 , w_21033 , w_21034 , w_21035 , w_21036 , w_21037 , w_21038 , w_21039 , 
		w_21040 , w_21041 , w_21042 , w_21043 , w_21044 , w_21045 , w_21046 , w_21047 , w_21048 , w_21049 , 
		w_21050 , w_21051 , w_21052 , w_21053 , w_21054 , w_21055 , w_21056 , w_21057 , w_21058 , w_21059 , 
		w_21060 , w_21061 , w_21062 , w_21063 , w_21064 , w_21065 , w_21066 , w_21067 , w_21068 , w_21069 , 
		w_21070 , w_21071 , w_21072 , w_21073 , w_21074 , w_21075 , w_21076 , w_21077 , w_21078 , w_21079 , 
		w_21080 , w_21081 , w_21082 , w_21083 , w_21084 , w_21085 , w_21086 , w_21087 , w_21088 , w_21089 , 
		w_21090 , w_21091 , w_21092 , w_21093 , w_21094 , w_21095 , w_21096 , w_21097 , w_21098 , w_21099 , 
		w_21100 , w_21101 , w_21102 , w_21103 , w_21104 , w_21105 , w_21106 , w_21107 , w_21108 , w_21109 , 
		w_21110 , w_21111 , w_21112 , w_21113 , w_21114 , w_21115 , w_21116 , w_21117 , w_21118 , w_21119 , 
		w_21120 , w_21121 , w_21122 , w_21123 , w_21124 , w_21125 , w_21126 , w_21127 , w_21128 , w_21129 , 
		w_21130 , w_21131 , w_21132 , w_21133 , w_21134 , w_21135 , w_21136 , w_21137 , w_21138 , w_21139 , 
		w_21140 , w_21141 , w_21142 , w_21143 , w_21144 , w_21145 , w_21146 , w_21147 , w_21148 , w_21149 , 
		w_21150 , w_21151 , w_21152 , w_21153 , w_21154 , w_21155 , w_21156 , w_21157 , w_21158 , w_21159 , 
		w_21160 , w_21161 , w_21162 , w_21163 , w_21164 , w_21165 , w_21166 , w_21167 , w_21168 , w_21169 , 
		w_21170 , w_21171 , w_21172 , w_21173 , w_21174 , w_21175 , w_21176 , w_21177 , w_21178 , w_21179 , 
		w_21180 , w_21181 , w_21182 , w_21183 , w_21184 , w_21185 , w_21186 , w_21187 , w_21188 , w_21189 , 
		w_21190 , w_21191 , w_21192 , w_21193 , w_21194 , w_21195 , w_21196 , w_21197 , w_21198 , w_21199 , 
		w_21200 , w_21201 , w_21202 , w_21203 , w_21204 , w_21205 , w_21206 , w_21207 , w_21208 , w_21209 , 
		w_21210 , w_21211 , w_21212 , w_21213 , w_21214 , w_21215 , w_21216 , w_21217 , w_21218 , w_21219 , 
		w_21220 , w_21221 , w_21222 , w_21223 , w_21224 , w_21225 , w_21226 , w_21227 , w_21228 , w_21229 , 
		w_21230 , w_21231 , w_21232 , w_21233 , w_21234 , w_21235 , w_21236 , w_21237 , w_21238 , w_21239 , 
		w_21240 , w_21241 , w_21242 , w_21243 , w_21244 , w_21245 , w_21246 , w_21247 , w_21248 , w_21249 , 
		w_21250 , w_21251 , w_21252 , w_21253 , w_21254 , w_21255 , w_21256 , w_21257 , w_21258 , w_21259 , 
		w_21260 , w_21261 , w_21262 , w_21263 , w_21264 , w_21265 , w_21266 , w_21267 , w_21268 , w_21269 , 
		w_21270 , w_21271 , w_21272 , w_21273 , w_21274 , w_21275 , w_21276 , w_21277 , w_21278 , w_21279 , 
		w_21280 , w_21281 , w_21282 , w_21283 , w_21284 , w_21285 , w_21286 , w_21287 , w_21288 , w_21289 , 
		w_21290 , w_21291 , w_21292 , w_21293 , w_21294 , w_21295 , w_21296 , w_21297 , w_21298 , w_21299 , 
		w_21300 , w_21301 , w_21302 , w_21303 , w_21304 , w_21305 , w_21306 , w_21307 , w_21308 , w_21309 , 
		w_21310 , w_21311 , w_21312 , w_21313 , w_21314 , w_21315 , w_21316 , w_21317 , w_21318 , w_21319 , 
		w_21320 , w_21321 , w_21322 , w_21323 , w_21324 , w_21325 , w_21326 , w_21327 , w_21328 , w_21329 , 
		w_21330 , w_21331 , w_21332 , w_21333 , w_21334 , w_21335 , w_21336 , w_21337 , w_21338 , w_21339 , 
		w_21340 , w_21341 , w_21342 , w_21343 , w_21344 , w_21345 , w_21346 , w_21347 , w_21348 , w_21349 , 
		w_21350 , w_21351 , w_21352 , w_21353 , w_21354 , w_21355 , w_21356 , w_21357 , w_21358 , w_21359 , 
		w_21360 , w_21361 , w_21362 , w_21363 , w_21364 , w_21365 , w_21366 , w_21367 , w_21368 , w_21369 , 
		w_21370 , w_21371 , w_21372 , w_21373 , w_21374 , w_21375 , w_21376 , w_21377 , w_21378 , w_21379 , 
		w_21380 , w_21381 , w_21382 , w_21383 , w_21384 , w_21385 , w_21386 , w_21387 , w_21388 , w_21389 , 
		w_21390 , w_21391 , w_21392 , w_21393 , w_21394 , w_21395 , w_21396 , w_21397 , w_21398 , w_21399 , 
		w_21400 , w_21401 , w_21402 , w_21403 , w_21404 , w_21405 , w_21406 , w_21407 , w_21408 , w_21409 , 
		w_21410 , w_21411 , w_21412 , w_21413 , w_21414 , w_21415 , w_21416 , w_21417 , w_21418 , w_21419 , 
		w_21420 , w_21421 , w_21422 , w_21423 , w_21424 , w_21425 , w_21426 , w_21427 , w_21428 , w_21429 , 
		w_21430 , w_21431 , w_21432 , w_21433 , w_21434 , w_21435 , w_21436 , w_21437 , w_21438 , w_21439 , 
		w_21440 , w_21441 , w_21442 , w_21443 , w_21444 , w_21445 , w_21446 , w_21447 , w_21448 , w_21449 , 
		w_21450 , w_21451 , w_21452 , w_21453 , w_21454 , w_21455 , w_21456 , w_21457 , w_21458 , w_21459 , 
		w_21460 , w_21461 , w_21462 , w_21463 , w_21464 , w_21465 , w_21466 , w_21467 , w_21468 , w_21469 , 
		w_21470 , w_21471 , w_21472 , w_21473 , w_21474 , w_21475 , w_21476 , w_21477 , w_21478 , w_21479 , 
		w_21480 , w_21481 , w_21482 , w_21483 , w_21484 , w_21485 , w_21486 , w_21487 , w_21488 , w_21489 , 
		w_21490 , w_21491 , w_21492 , w_21493 , w_21494 , w_21495 , w_21496 , w_21497 , w_21498 , w_21499 , 
		w_21500 , w_21501 , w_21502 , w_21503 , w_21504 , w_21505 , w_21506 , w_21507 , w_21508 , w_21509 , 
		w_21510 , w_21511 , w_21512 , w_21513 , w_21514 , w_21515 , w_21516 , w_21517 , w_21518 , w_21519 , 
		w_21520 , w_21521 , w_21522 , w_21523 , w_21524 , w_21525 , w_21526 , w_21527 , w_21528 , w_21529 , 
		w_21530 , w_21531 , w_21532 , w_21533 , w_21534 , w_21535 , w_21536 , w_21537 , w_21538 , w_21539 , 
		w_21540 , w_21541 , w_21542 , w_21543 , w_21544 , w_21545 , w_21546 , w_21547 , w_21548 , w_21549 , 
		w_21550 , w_21551 , w_21552 , w_21553 , w_21554 , w_21555 , w_21556 , w_21557 , w_21558 , w_21559 , 
		w_21560 , w_21561 , w_21562 , w_21563 , w_21564 , w_21565 , w_21566 , w_21567 , w_21568 , w_21569 , 
		w_21570 , w_21571 , w_21572 , w_21573 , w_21574 , w_21575 , w_21576 , w_21577 , w_21578 , w_21579 , 
		w_21580 , w_21581 , w_21582 , w_21583 , w_21584 , w_21585 , w_21586 , w_21587 , w_21588 , w_21589 , 
		w_21590 , w_21591 , w_21592 , w_21593 , w_21594 , w_21595 , w_21596 , w_21597 , w_21598 , w_21599 , 
		w_21600 , w_21601 , w_21602 , w_21603 , w_21604 , w_21605 , w_21606 , w_21607 , w_21608 , w_21609 , 
		w_21610 , w_21611 , w_21612 , w_21613 , w_21614 , w_21615 , w_21616 , w_21617 , w_21618 , w_21619 , 
		w_21620 , w_21621 , w_21622 , w_21623 , w_21624 , w_21625 , w_21626 , w_21627 , w_21628 , w_21629 , 
		w_21630 , w_21631 , w_21632 , w_21633 , w_21634 , w_21635 , w_21636 , w_21637 , w_21638 , w_21639 , 
		w_21640 , w_21641 , w_21642 , w_21643 , w_21644 , w_21645 , w_21646 , w_21647 , w_21648 , w_21649 , 
		w_21650 , w_21651 , w_21652 , w_21653 , w_21654 , w_21655 , w_21656 , w_21657 , w_21658 , w_21659 , 
		w_21660 , w_21661 , w_21662 , w_21663 , w_21664 , w_21665 , w_21666 , w_21667 , w_21668 , w_21669 , 
		w_21670 , w_21671 , w_21672 , w_21673 , w_21674 , w_21675 , w_21676 , w_21677 , w_21678 , w_21679 , 
		w_21680 , w_21681 , w_21682 , w_21683 , w_21684 , w_21685 , w_21686 , w_21687 , w_21688 , w_21689 , 
		w_21690 , w_21691 , w_21692 , w_21693 , w_21694 , w_21695 , w_21696 , w_21697 , w_21698 , w_21699 , 
		w_21700 , w_21701 , w_21702 , w_21703 , w_21704 , w_21705 , w_21706 , w_21707 , w_21708 , w_21709 , 
		w_21710 , w_21711 , w_21712 , w_21713 , w_21714 , w_21715 , w_21716 , w_21717 , w_21718 , w_21719 , 
		w_21720 , w_21721 , w_21722 , w_21723 , w_21724 , w_21725 , w_21726 , w_21727 , w_21728 , w_21729 , 
		w_21730 , w_21731 , w_21732 , w_21733 , w_21734 , w_21735 , w_21736 , w_21737 , w_21738 , w_21739 , 
		w_21740 , w_21741 , w_21742 , w_21743 , w_21744 , w_21745 , w_21746 , w_21747 , w_21748 , w_21749 , 
		w_21750 , w_21751 , w_21752 , w_21753 , w_21754 , w_21755 , w_21756 , w_21757 , w_21758 , w_21759 , 
		w_21760 , w_21761 , w_21762 , w_21763 , w_21764 , w_21765 , w_21766 , w_21767 , w_21768 , w_21769 , 
		w_21770 , w_21771 , w_21772 , w_21773 , w_21774 , w_21775 , w_21776 , w_21777 , w_21778 , w_21779 , 
		w_21780 , w_21781 , w_21782 , w_21783 , w_21784 , w_21785 , w_21786 , w_21787 , w_21788 , w_21789 , 
		w_21790 , w_21791 , w_21792 , w_21793 , w_21794 , w_21795 , w_21796 , w_21797 , w_21798 , w_21799 , 
		w_21800 , w_21801 , w_21802 , w_21803 , w_21804 , w_21805 , w_21806 , w_21807 , w_21808 , w_21809 , 
		w_21810 , w_21811 , w_21812 , w_21813 , w_21814 , w_21815 , w_21816 , w_21817 , w_21818 , w_21819 , 
		w_21820 , w_21821 , w_21822 , w_21823 , w_21824 , w_21825 , w_21826 , w_21827 , w_21828 , w_21829 , 
		w_21830 , w_21831 , w_21832 , w_21833 , w_21834 , w_21835 , w_21836 , w_21837 , w_21838 , w_21839 , 
		w_21840 , w_21841 , w_21842 , w_21843 , w_21844 , w_21845 , w_21846 , w_21847 , w_21848 , w_21849 , 
		w_21850 , w_21851 , w_21852 , w_21853 , w_21854 , w_21855 , w_21856 , w_21857 , w_21858 , w_21859 , 
		w_21860 , w_21861 , w_21862 , w_21863 , w_21864 , w_21865 , w_21866 , w_21867 , w_21868 , w_21869 , 
		w_21870 , w_21871 , w_21872 , w_21873 , w_21874 , w_21875 , w_21876 , w_21877 , w_21878 , w_21879 , 
		w_21880 , w_21881 , w_21882 , w_21883 , w_21884 , w_21885 , w_21886 , w_21887 , w_21888 , w_21889 , 
		w_21890 , w_21891 , w_21892 , w_21893 , w_21894 , w_21895 , w_21896 , w_21897 , w_21898 , w_21899 , 
		w_21900 , w_21901 , w_21902 , w_21903 , w_21904 , w_21905 , w_21906 , w_21907 , w_21908 , w_21909 , 
		w_21910 , w_21911 , w_21912 , w_21913 , w_21914 , w_21915 , w_21916 , w_21917 , w_21918 , w_21919 , 
		w_21920 , w_21921 , w_21922 , w_21923 , w_21924 , w_21925 , w_21926 , w_21927 , w_21928 , w_21929 , 
		w_21930 , w_21931 , w_21932 , w_21933 , w_21934 , w_21935 , w_21936 , w_21937 , w_21938 , w_21939 , 
		w_21940 , w_21941 , w_21942 , w_21943 , w_21944 , w_21945 , w_21946 , w_21947 , w_21948 , w_21949 , 
		w_21950 , w_21951 , w_21952 , w_21953 , w_21954 , w_21955 , w_21956 , w_21957 , w_21958 , w_21959 , 
		w_21960 , w_21961 , w_21962 , w_21963 , w_21964 , w_21965 , w_21966 , w_21967 , w_21968 , w_21969 , 
		w_21970 , w_21971 , w_21972 , w_21973 , w_21974 , w_21975 , w_21976 , w_21977 , w_21978 , w_21979 , 
		w_21980 , w_21981 , w_21982 , w_21983 , w_21984 , w_21985 , w_21986 , w_21987 , w_21988 , w_21989 , 
		w_21990 , w_21991 , w_21992 , w_21993 , w_21994 , w_21995 , w_21996 , w_21997 , w_21998 , w_21999 , 
		w_22000 , w_22001 , w_22002 , w_22003 , w_22004 , w_22005 , w_22006 , w_22007 , w_22008 , w_22009 , 
		w_22010 , w_22011 , w_22012 , w_22013 , w_22014 , w_22015 , w_22016 , w_22017 , w_22018 , w_22019 , 
		w_22020 , w_22021 , w_22022 , w_22023 , w_22024 , w_22025 , w_22026 , w_22027 , w_22028 , w_22029 , 
		w_22030 , w_22031 , w_22032 , w_22033 , w_22034 , w_22035 , w_22036 , w_22037 , w_22038 , w_22039 , 
		w_22040 , w_22041 , w_22042 , w_22043 , w_22044 , w_22045 , w_22046 , w_22047 , w_22048 , w_22049 , 
		w_22050 , w_22051 , w_22052 , w_22053 , w_22054 , w_22055 , w_22056 , w_22057 , w_22058 , w_22059 , 
		w_22060 , w_22061 , w_22062 , w_22063 , w_22064 , w_22065 , w_22066 , w_22067 , w_22068 , w_22069 , 
		w_22070 , w_22071 , w_22072 , w_22073 , w_22074 , w_22075 , w_22076 , w_22077 , w_22078 , w_22079 , 
		w_22080 , w_22081 , w_22082 , w_22083 , w_22084 , w_22085 , w_22086 , w_22087 , w_22088 , w_22089 , 
		w_22090 , w_22091 , w_22092 , w_22093 , w_22094 , w_22095 , w_22096 , w_22097 , w_22098 , w_22099 , 
		w_22100 , w_22101 , w_22102 , w_22103 , w_22104 , w_22105 , w_22106 , w_22107 , w_22108 , w_22109 , 
		w_22110 , w_22111 , w_22112 , w_22113 , w_22114 , w_22115 , w_22116 , w_22117 , w_22118 , w_22119 , 
		w_22120 , w_22121 , w_22122 , w_22123 , w_22124 , w_22125 , w_22126 , w_22127 , w_22128 , w_22129 , 
		w_22130 , w_22131 , w_22132 , w_22133 , w_22134 , w_22135 , w_22136 , w_22137 , w_22138 , w_22139 , 
		w_22140 , w_22141 , w_22142 , w_22143 , w_22144 , w_22145 , w_22146 , w_22147 , w_22148 , w_22149 , 
		w_22150 , w_22151 , w_22152 , w_22153 , w_22154 , w_22155 , w_22156 , w_22157 , w_22158 , w_22159 , 
		w_22160 , w_22161 , w_22162 , w_22163 , w_22164 , w_22165 , w_22166 , w_22167 , w_22168 , w_22169 , 
		w_22170 , w_22171 , w_22172 , w_22173 , w_22174 , w_22175 , w_22176 , w_22177 , w_22178 , w_22179 , 
		w_22180 , w_22181 , w_22182 , w_22183 , w_22184 , w_22185 , w_22186 , w_22187 , w_22188 , w_22189 , 
		w_22190 , w_22191 , w_22192 , w_22193 , w_22194 , w_22195 , w_22196 , w_22197 , w_22198 , w_22199 , 
		w_22200 , w_22201 , w_22202 , w_22203 , w_22204 , w_22205 , w_22206 , w_22207 , w_22208 , w_22209 , 
		w_22210 , w_22211 , w_22212 , w_22213 , w_22214 , w_22215 , w_22216 , w_22217 , w_22218 , w_22219 , 
		w_22220 , w_22221 , w_22222 , w_22223 , w_22224 , w_22225 , w_22226 , w_22227 , w_22228 , w_22229 , 
		w_22230 , w_22231 , w_22232 , w_22233 , w_22234 , w_22235 , w_22236 , w_22237 , w_22238 , w_22239 , 
		w_22240 , w_22241 , w_22242 , w_22243 , w_22244 , w_22245 , w_22246 , w_22247 , w_22248 , w_22249 , 
		w_22250 , w_22251 , w_22252 , w_22253 , w_22254 , w_22255 , w_22256 , w_22257 , w_22258 , w_22259 , 
		w_22260 , w_22261 , w_22262 , w_22263 , w_22264 , w_22265 , w_22266 , w_22267 , w_22268 , w_22269 , 
		w_22270 , w_22271 , w_22272 , w_22273 , w_22274 , w_22275 , w_22276 , w_22277 , w_22278 , w_22279 , 
		w_22280 , w_22281 , w_22282 , w_22283 , w_22284 , w_22285 , w_22286 , w_22287 , w_22288 , w_22289 , 
		w_22290 , w_22291 , w_22292 , w_22293 , w_22294 , w_22295 , w_22296 , w_22297 , w_22298 , w_22299 , 
		w_22300 , w_22301 , w_22302 , w_22303 , w_22304 , w_22305 , w_22306 , w_22307 , w_22308 , w_22309 , 
		w_22310 , w_22311 , w_22312 , w_22313 , w_22314 , w_22315 , w_22316 , w_22317 , w_22318 , w_22319 , 
		w_22320 , w_22321 , w_22322 , w_22323 , w_22324 , w_22325 , w_22326 , w_22327 , w_22328 , w_22329 , 
		w_22330 , w_22331 , w_22332 , w_22333 , w_22334 , w_22335 , w_22336 , w_22337 , w_22338 , w_22339 , 
		w_22340 , w_22341 , w_22342 , w_22343 , w_22344 , w_22345 , w_22346 , w_22347 , w_22348 , w_22349 , 
		w_22350 , w_22351 , w_22352 , w_22353 , w_22354 , w_22355 , w_22356 , w_22357 , w_22358 , w_22359 , 
		w_22360 , w_22361 , w_22362 , w_22363 , w_22364 , w_22365 , w_22366 , w_22367 , w_22368 , w_22369 , 
		w_22370 , w_22371 , w_22372 , w_22373 , w_22374 , w_22375 , w_22376 , w_22377 , w_22378 , w_22379 , 
		w_22380 , w_22381 , w_22382 , w_22383 , w_22384 , w_22385 , w_22386 , w_22387 , w_22388 , w_22389 , 
		w_22390 , w_22391 , w_22392 , w_22393 , w_22394 , w_22395 , w_22396 , w_22397 , w_22398 , w_22399 , 
		w_22400 , w_22401 , w_22402 , w_22403 , w_22404 , w_22405 , w_22406 , w_22407 , w_22408 , w_22409 , 
		w_22410 , w_22411 , w_22412 , w_22413 , w_22414 , w_22415 , w_22416 , w_22417 , w_22418 , w_22419 , 
		w_22420 , w_22421 , w_22422 , w_22423 , w_22424 , w_22425 , w_22426 , w_22427 , w_22428 , w_22429 , 
		w_22430 , w_22431 , w_22432 , w_22433 , w_22434 , w_22435 , w_22436 , w_22437 , w_22438 , w_22439 , 
		w_22440 , w_22441 , w_22442 , w_22443 , w_22444 , w_22445 , w_22446 , w_22447 , w_22448 , w_22449 , 
		w_22450 , w_22451 , w_22452 , w_22453 , w_22454 , w_22455 , w_22456 , w_22457 , w_22458 , w_22459 , 
		w_22460 , w_22461 , w_22462 , w_22463 , w_22464 , w_22465 , w_22466 , w_22467 , w_22468 , w_22469 , 
		w_22470 , w_22471 , w_22472 , w_22473 , w_22474 , w_22475 , w_22476 , w_22477 , w_22478 , w_22479 , 
		w_22480 , w_22481 , w_22482 , w_22483 , w_22484 , w_22485 , w_22486 , w_22487 , w_22488 , w_22489 , 
		w_22490 , w_22491 , w_22492 , w_22493 , w_22494 , w_22495 , w_22496 , w_22497 , w_22498 , w_22499 , 
		w_22500 , w_22501 , w_22502 , w_22503 , w_22504 , w_22505 , w_22506 , w_22507 , w_22508 , w_22509 , 
		w_22510 , w_22511 , w_22512 , w_22513 , w_22514 , w_22515 , w_22516 , w_22517 , w_22518 , w_22519 , 
		w_22520 , w_22521 , w_22522 , w_22523 , w_22524 , w_22525 , w_22526 , w_22527 , w_22528 , w_22529 , 
		w_22530 , w_22531 , w_22532 , w_22533 , w_22534 , w_22535 , w_22536 , w_22537 , w_22538 , w_22539 , 
		w_22540 , w_22541 , w_22542 , w_22543 , w_22544 , w_22545 , w_22546 , w_22547 , w_22548 , w_22549 , 
		w_22550 , w_22551 , w_22552 , w_22553 , w_22554 , w_22555 , w_22556 , w_22557 , w_22558 , w_22559 , 
		w_22560 , w_22561 , w_22562 , w_22563 , w_22564 , w_22565 , w_22566 , w_22567 , w_22568 , w_22569 , 
		w_22570 , w_22571 , w_22572 , w_22573 , w_22574 , w_22575 , w_22576 , w_22577 , w_22578 , w_22579 , 
		w_22580 , w_22581 , w_22582 , w_22583 , w_22584 , w_22585 , w_22586 , w_22587 , w_22588 , w_22589 , 
		w_22590 , w_22591 , w_22592 , w_22593 , w_22594 , w_22595 , w_22596 , w_22597 , w_22598 , w_22599 , 
		w_22600 , w_22601 , w_22602 , w_22603 , w_22604 , w_22605 , w_22606 , w_22607 , w_22608 , w_22609 , 
		w_22610 , w_22611 , w_22612 , w_22613 , w_22614 , w_22615 , w_22616 , w_22617 , w_22618 , w_22619 , 
		w_22620 , w_22621 , w_22622 , w_22623 , w_22624 , w_22625 , w_22626 , w_22627 , w_22628 , w_22629 , 
		w_22630 , w_22631 , w_22632 , w_22633 , w_22634 , w_22635 , w_22636 , w_22637 , w_22638 , w_22639 , 
		w_22640 , w_22641 , w_22642 , w_22643 , w_22644 , w_22645 , w_22646 , w_22647 , w_22648 , w_22649 , 
		w_22650 , w_22651 , w_22652 , w_22653 , w_22654 , w_22655 , w_22656 , w_22657 , w_22658 , w_22659 , 
		w_22660 , w_22661 , w_22662 , w_22663 , w_22664 , w_22665 , w_22666 , w_22667 , w_22668 , w_22669 , 
		w_22670 , w_22671 , w_22672 , w_22673 , w_22674 , w_22675 , w_22676 , w_22677 , w_22678 , w_22679 , 
		w_22680 , w_22681 , w_22682 , w_22683 , w_22684 , w_22685 , w_22686 , w_22687 , w_22688 , w_22689 , 
		w_22690 , w_22691 , w_22692 , w_22693 , w_22694 , w_22695 , w_22696 , w_22697 , w_22698 , w_22699 , 
		w_22700 , w_22701 , w_22702 , w_22703 , w_22704 , w_22705 , w_22706 , w_22707 , w_22708 , w_22709 , 
		w_22710 , w_22711 , w_22712 , w_22713 , w_22714 , w_22715 , w_22716 , w_22717 , w_22718 , w_22719 , 
		w_22720 , w_22721 , w_22722 , w_22723 , w_22724 , w_22725 , w_22726 , w_22727 , w_22728 , w_22729 , 
		w_22730 , w_22731 , w_22732 , w_22733 , w_22734 , w_22735 , w_22736 , w_22737 , w_22738 , w_22739 , 
		w_22740 , w_22741 , w_22742 , w_22743 , w_22744 , w_22745 , w_22746 , w_22747 , w_22748 , w_22749 , 
		w_22750 , w_22751 , w_22752 , w_22753 , w_22754 , w_22755 , w_22756 , w_22757 , w_22758 , w_22759 , 
		w_22760 , w_22761 , w_22762 , w_22763 , w_22764 , w_22765 , w_22766 , w_22767 , w_22768 , w_22769 , 
		w_22770 , w_22771 , w_22772 , w_22773 , w_22774 , w_22775 , w_22776 , w_22777 , w_22778 , w_22779 , 
		w_22780 , w_22781 , w_22782 , w_22783 , w_22784 , w_22785 , w_22786 , w_22787 , w_22788 , w_22789 , 
		w_22790 , w_22791 , w_22792 , w_22793 , w_22794 , w_22795 , w_22796 , w_22797 , w_22798 , w_22799 , 
		w_22800 , w_22801 , w_22802 , w_22803 , w_22804 , w_22805 , w_22806 , w_22807 , w_22808 , w_22809 , 
		w_22810 , w_22811 , w_22812 , w_22813 , w_22814 , w_22815 , w_22816 , w_22817 , w_22818 , w_22819 , 
		w_22820 , w_22821 , w_22822 , w_22823 , w_22824 , w_22825 , w_22826 , w_22827 , w_22828 , w_22829 , 
		w_22830 , w_22831 , w_22832 , w_22833 , w_22834 , w_22835 , w_22836 , w_22837 , w_22838 , w_22839 , 
		w_22840 , w_22841 , w_22842 , w_22843 , w_22844 , w_22845 , w_22846 , w_22847 , w_22848 , w_22849 , 
		w_22850 , w_22851 , w_22852 , w_22853 , w_22854 , w_22855 , w_22856 , w_22857 , w_22858 , w_22859 , 
		w_22860 , w_22861 , w_22862 , w_22863 , w_22864 , w_22865 , w_22866 , w_22867 , w_22868 , w_22869 , 
		w_22870 , w_22871 , w_22872 , w_22873 , w_22874 , w_22875 , w_22876 , w_22877 , w_22878 , w_22879 , 
		w_22880 , w_22881 , w_22882 , w_22883 , w_22884 , w_22885 , w_22886 , w_22887 , w_22888 , w_22889 , 
		w_22890 , w_22891 , w_22892 , w_22893 , w_22894 , w_22895 , w_22896 , w_22897 , w_22898 , w_22899 , 
		w_22900 , w_22901 , w_22902 , w_22903 , w_22904 , w_22905 , w_22906 , w_22907 , w_22908 , w_22909 , 
		w_22910 , w_22911 , w_22912 , w_22913 , w_22914 , w_22915 , w_22916 , w_22917 , w_22918 , w_22919 , 
		w_22920 , w_22921 , w_22922 , w_22923 , w_22924 , w_22925 , w_22926 , w_22927 , w_22928 , w_22929 , 
		w_22930 , w_22931 , w_22932 , w_22933 , w_22934 , w_22935 , w_22936 , w_22937 , w_22938 , w_22939 , 
		w_22940 , w_22941 , w_22942 , w_22943 , w_22944 , w_22945 , w_22946 , w_22947 , w_22948 , w_22949 , 
		w_22950 , w_22951 , w_22952 , w_22953 , w_22954 , w_22955 , w_22956 , w_22957 , w_22958 , w_22959 , 
		w_22960 , w_22961 , w_22962 , w_22963 , w_22964 , w_22965 , w_22966 , w_22967 , w_22968 , w_22969 , 
		w_22970 , w_22971 , w_22972 , w_22973 , w_22974 , w_22975 , w_22976 , w_22977 , w_22978 , w_22979 , 
		w_22980 , w_22981 , w_22982 , w_22983 , w_22984 , w_22985 , w_22986 , w_22987 , w_22988 , w_22989 , 
		w_22990 , w_22991 , w_22992 , w_22993 , w_22994 , w_22995 , w_22996 , w_22997 , w_22998 , w_22999 , 
		w_23000 , w_23001 , w_23002 , w_23003 , w_23004 , w_23005 , w_23006 , w_23007 , w_23008 , w_23009 , 
		w_23010 , w_23011 , w_23012 , w_23013 , w_23014 , w_23015 , w_23016 , w_23017 , w_23018 , w_23019 , 
		w_23020 , w_23021 , w_23022 , w_23023 , w_23024 , w_23025 , w_23026 , w_23027 , w_23028 , w_23029 , 
		w_23030 , w_23031 , w_23032 , w_23033 , w_23034 , w_23035 , w_23036 , w_23037 , w_23038 , w_23039 , 
		w_23040 , w_23041 , w_23042 , w_23043 , w_23044 , w_23045 , w_23046 , w_23047 , w_23048 , w_23049 , 
		w_23050 , w_23051 , w_23052 , w_23053 , w_23054 , w_23055 , w_23056 , w_23057 , w_23058 , w_23059 , 
		w_23060 , w_23061 , w_23062 , w_23063 , w_23064 , w_23065 , w_23066 , w_23067 , w_23068 , w_23069 , 
		w_23070 , w_23071 , w_23072 , w_23073 , w_23074 , w_23075 , w_23076 , w_23077 , w_23078 , w_23079 , 
		w_23080 , w_23081 , w_23082 , w_23083 , w_23084 , w_23085 , w_23086 , w_23087 , w_23088 , w_23089 , 
		w_23090 , w_23091 , w_23092 , w_23093 , w_23094 , w_23095 , w_23096 , w_23097 , w_23098 , w_23099 , 
		w_23100 , w_23101 , w_23102 , w_23103 , w_23104 , w_23105 , w_23106 , w_23107 , w_23108 , w_23109 , 
		w_23110 , w_23111 , w_23112 , w_23113 , w_23114 , w_23115 , w_23116 , w_23117 , w_23118 , w_23119 , 
		w_23120 , w_23121 , w_23122 , w_23123 , w_23124 , w_23125 , w_23126 , w_23127 , w_23128 , w_23129 , 
		w_23130 , w_23131 , w_23132 , w_23133 , w_23134 , w_23135 , w_23136 , w_23137 , w_23138 , w_23139 , 
		w_23140 , w_23141 , w_23142 , w_23143 , w_23144 , w_23145 , w_23146 , w_23147 , w_23148 , w_23149 , 
		w_23150 , w_23151 , w_23152 , w_23153 , w_23154 , w_23155 , w_23156 , w_23157 , w_23158 , w_23159 , 
		w_23160 , w_23161 , w_23162 , w_23163 , w_23164 , w_23165 , w_23166 , w_23167 , w_23168 , w_23169 , 
		w_23170 , w_23171 , w_23172 , w_23173 , w_23174 , w_23175 , w_23176 , w_23177 , w_23178 , w_23179 , 
		w_23180 , w_23181 , w_23182 , w_23183 , w_23184 , w_23185 , w_23186 , w_23187 , w_23188 , w_23189 , 
		w_23190 , w_23191 , w_23192 , w_23193 , w_23194 , w_23195 , w_23196 , w_23197 , w_23198 , w_23199 , 
		w_23200 , w_23201 , w_23202 , w_23203 , w_23204 , w_23205 , w_23206 , w_23207 , w_23208 , w_23209 , 
		w_23210 , w_23211 , w_23212 , w_23213 , w_23214 , w_23215 , w_23216 , w_23217 , w_23218 , w_23219 , 
		w_23220 , w_23221 , w_23222 , w_23223 , w_23224 , w_23225 , w_23226 , w_23227 , w_23228 , w_23229 , 
		w_23230 , w_23231 , w_23232 , w_23233 , w_23234 , w_23235 , w_23236 , w_23237 , w_23238 , w_23239 , 
		w_23240 , w_23241 , w_23242 , w_23243 , w_23244 , w_23245 , w_23246 , w_23247 , w_23248 , w_23249 , 
		w_23250 , w_23251 , w_23252 , w_23253 , w_23254 , w_23255 , w_23256 , w_23257 , w_23258 , w_23259 , 
		w_23260 , w_23261 , w_23262 , w_23263 , w_23264 , w_23265 , w_23266 , w_23267 , w_23268 , w_23269 , 
		w_23270 , w_23271 , w_23272 , w_23273 , w_23274 , w_23275 , w_23276 , w_23277 , w_23278 , w_23279 , 
		w_23280 , w_23281 , w_23282 , w_23283 , w_23284 , w_23285 , w_23286 , w_23287 , w_23288 , w_23289 , 
		w_23290 , w_23291 , w_23292 , w_23293 , w_23294 , w_23295 , w_23296 , w_23297 , w_23298 , w_23299 , 
		w_23300 , w_23301 , w_23302 , w_23303 , w_23304 , w_23305 , w_23306 , w_23307 , w_23308 , w_23309 , 
		w_23310 , w_23311 , w_23312 , w_23313 , w_23314 , w_23315 , w_23316 , w_23317 , w_23318 , w_23319 , 
		w_23320 , w_23321 , w_23322 , w_23323 , w_23324 , w_23325 , w_23326 , w_23327 , w_23328 , w_23329 , 
		w_23330 , w_23331 , w_23332 , w_23333 , w_23334 , w_23335 , w_23336 , w_23337 , w_23338 , w_23339 , 
		w_23340 , w_23341 , w_23342 , w_23343 , w_23344 , w_23345 , w_23346 , w_23347 , w_23348 , w_23349 , 
		w_23350 , w_23351 , w_23352 , w_23353 , w_23354 , w_23355 , w_23356 , w_23357 , w_23358 , w_23359 , 
		w_23360 , w_23361 , w_23362 , w_23363 , w_23364 , w_23365 , w_23366 , w_23367 , w_23368 , w_23369 , 
		w_23370 , w_23371 , w_23372 , w_23373 , w_23374 , w_23375 , w_23376 , w_23377 , w_23378 , w_23379 , 
		w_23380 , w_23381 , w_23382 , w_23383 , w_23384 , w_23385 , w_23386 , w_23387 , w_23388 , w_23389 , 
		w_23390 , w_23391 , w_23392 , w_23393 , w_23394 , w_23395 , w_23396 , w_23397 , w_23398 , w_23399 , 
		w_23400 , w_23401 , w_23402 , w_23403 , w_23404 , w_23405 , w_23406 , w_23407 , w_23408 , w_23409 , 
		w_23410 , w_23411 , w_23412 , w_23413 , w_23414 , w_23415 , w_23416 , w_23417 , w_23418 , w_23419 , 
		w_23420 , w_23421 , w_23422 , w_23423 , w_23424 , w_23425 , w_23426 , w_23427 , w_23428 , w_23429 , 
		w_23430 , w_23431 , w_23432 , w_23433 , w_23434 , w_23435 , w_23436 , w_23437 , w_23438 , w_23439 , 
		w_23440 , w_23441 , w_23442 , w_23443 , w_23444 , w_23445 , w_23446 , w_23447 , w_23448 , w_23449 , 
		w_23450 , w_23451 , w_23452 , w_23453 , w_23454 , w_23455 , w_23456 , w_23457 , w_23458 , w_23459 , 
		w_23460 , w_23461 , w_23462 , w_23463 , w_23464 , w_23465 , w_23466 , w_23467 , w_23468 , w_23469 , 
		w_23470 , w_23471 , w_23472 , w_23473 , w_23474 , w_23475 , w_23476 , w_23477 , w_23478 , w_23479 , 
		w_23480 , w_23481 , w_23482 , w_23483 , w_23484 , w_23485 , w_23486 , w_23487 , w_23488 , w_23489 , 
		w_23490 , w_23491 , w_23492 , w_23493 , w_23494 , w_23495 , w_23496 , w_23497 , w_23498 , w_23499 , 
		w_23500 , w_23501 , w_23502 , w_23503 , w_23504 , w_23505 , w_23506 , w_23507 , w_23508 , w_23509 , 
		w_23510 , w_23511 , w_23512 , w_23513 , w_23514 , w_23515 , w_23516 , w_23517 , w_23518 , w_23519 , 
		w_23520 , w_23521 , w_23522 , w_23523 , w_23524 , w_23525 , w_23526 , w_23527 , w_23528 , w_23529 , 
		w_23530 , w_23531 , w_23532 , w_23533 , w_23534 , w_23535 , w_23536 , w_23537 , w_23538 , w_23539 , 
		w_23540 , w_23541 , w_23542 , w_23543 , w_23544 , w_23545 , w_23546 , w_23547 , w_23548 , w_23549 , 
		w_23550 , w_23551 , w_23552 , w_23553 , w_23554 , w_23555 , w_23556 , w_23557 , w_23558 , w_23559 , 
		w_23560 , w_23561 , w_23562 , w_23563 , w_23564 , w_23565 , w_23566 , w_23567 , w_23568 , w_23569 , 
		w_23570 , w_23571 , w_23572 , w_23573 , w_23574 , w_23575 , w_23576 , w_23577 , w_23578 , w_23579 , 
		w_23580 , w_23581 , w_23582 , w_23583 , w_23584 , w_23585 , w_23586 , w_23587 , w_23588 , w_23589 , 
		w_23590 , w_23591 , w_23592 , w_23593 , w_23594 , w_23595 , w_23596 , w_23597 , w_23598 , w_23599 , 
		w_23600 , w_23601 , w_23602 , w_23603 , w_23604 , w_23605 , w_23606 , w_23607 , w_23608 , w_23609 , 
		w_23610 , w_23611 , w_23612 , w_23613 , w_23614 , w_23615 , w_23616 , w_23617 , w_23618 , w_23619 , 
		w_23620 , w_23621 , w_23622 , w_23623 , w_23624 , w_23625 , w_23626 , w_23627 , w_23628 , w_23629 , 
		w_23630 , w_23631 , w_23632 , w_23633 , w_23634 , w_23635 , w_23636 , w_23637 , w_23638 , w_23639 , 
		w_23640 , w_23641 , w_23642 , w_23643 , w_23644 , w_23645 , w_23646 , w_23647 , w_23648 , w_23649 , 
		w_23650 , w_23651 , w_23652 , w_23653 , w_23654 , w_23655 , w_23656 , w_23657 , w_23658 , w_23659 , 
		w_23660 , w_23661 , w_23662 , w_23663 , w_23664 , w_23665 , w_23666 , w_23667 , w_23668 , w_23669 , 
		w_23670 , w_23671 , w_23672 , w_23673 , w_23674 , w_23675 , w_23676 , w_23677 , w_23678 , w_23679 , 
		w_23680 , w_23681 , w_23682 , w_23683 , w_23684 , w_23685 , w_23686 , w_23687 , w_23688 , w_23689 , 
		w_23690 , w_23691 , w_23692 , w_23693 , w_23694 , w_23695 , w_23696 , w_23697 , w_23698 , w_23699 , 
		w_23700 , w_23701 , w_23702 , w_23703 , w_23704 , w_23705 , w_23706 , w_23707 , w_23708 , w_23709 , 
		w_23710 , w_23711 , w_23712 , w_23713 , w_23714 , w_23715 , w_23716 , w_23717 , w_23718 , w_23719 , 
		w_23720 , w_23721 , w_23722 , w_23723 , w_23724 , w_23725 , w_23726 , w_23727 , w_23728 , w_23729 , 
		w_23730 , w_23731 , w_23732 , w_23733 , w_23734 , w_23735 , w_23736 , w_23737 , w_23738 , w_23739 , 
		w_23740 , w_23741 , w_23742 , w_23743 , w_23744 , w_23745 , w_23746 , w_23747 , w_23748 , w_23749 , 
		w_23750 , w_23751 , w_23752 , w_23753 , w_23754 , w_23755 , w_23756 , w_23757 , w_23758 , w_23759 , 
		w_23760 , w_23761 , w_23762 , w_23763 , w_23764 , w_23765 , w_23766 , w_23767 , w_23768 , w_23769 , 
		w_23770 , w_23771 , w_23772 , w_23773 , w_23774 , w_23775 , w_23776 , w_23777 , w_23778 , w_23779 , 
		w_23780 , w_23781 , w_23782 , w_23783 , w_23784 , w_23785 , w_23786 , w_23787 , w_23788 , w_23789 , 
		w_23790 , w_23791 , w_23792 , w_23793 , w_23794 , w_23795 , w_23796 , w_23797 , w_23798 , w_23799 , 
		w_23800 , w_23801 , w_23802 , w_23803 , w_23804 , w_23805 , w_23806 , w_23807 , w_23808 , w_23809 , 
		w_23810 , w_23811 , w_23812 , w_23813 , w_23814 , w_23815 , w_23816 , w_23817 , w_23818 , w_23819 , 
		w_23820 , w_23821 , w_23822 , w_23823 , w_23824 , w_23825 , w_23826 , w_23827 , w_23828 , w_23829 , 
		w_23830 , w_23831 , w_23832 , w_23833 , w_23834 , w_23835 , w_23836 , w_23837 , w_23838 , w_23839 , 
		w_23840 , w_23841 , w_23842 , w_23843 , w_23844 , w_23845 , w_23846 , w_23847 , w_23848 , w_23849 , 
		w_23850 , w_23851 , w_23852 , w_23853 , w_23854 , w_23855 , w_23856 , w_23857 , w_23858 , w_23859 , 
		w_23860 , w_23861 , w_23862 , w_23863 , w_23864 , w_23865 , w_23866 , w_23867 , w_23868 , w_23869 , 
		w_23870 , w_23871 , w_23872 , w_23873 , w_23874 , w_23875 ;
buf ( \o[31]_b1 , \6967_b1 );
buf ( \o[31]_b0 , \6967_b0 );
buf ( \o[30]_b1 , \7061_b1 );
buf ( \o[30]_b0 , \7061_b0 );
buf ( \o[29]_b1 , \6979_b1 );
buf ( \o[29]_b0 , \6979_b0 );
buf ( \o[28]_b1 , \6991_b1 );
buf ( \o[28]_b0 , \6991_b0 );
buf ( \o[27]_b1 , \7007_b1 );
buf ( \o[27]_b0 , \7007_b0 );
buf ( \o[26]_b1 , \7020_b1 );
buf ( \o[26]_b0 , \7020_b0 );
buf ( \o[25]_b1 , \7030_b1 );
buf ( \o[25]_b0 , \7030_b0 );
buf ( \o[24]_b1 , \7216_b1 );
buf ( \o[24]_b0 , \7216_b0 );
buf ( \o[23]_b1 , \7046_b1 );
buf ( \o[23]_b0 , \7046_b0 );
buf ( \o[22]_b1 , \7206_b1 );
buf ( \o[22]_b0 , \7206_b0 );
buf ( \o[21]_b1 , \7072_b1 );
buf ( \o[21]_b0 , \7072_b0 );
buf ( \o[20]_b1 , \7078_b1 );
buf ( \o[20]_b0 , \7078_b0 );
buf ( \o[19]_b1 , \7095_b1 );
buf ( \o[19]_b0 , \7095_b0 );
buf ( \o[18]_b1 , \7102_b1 );
buf ( \o[18]_b0 , \7102_b0 );
buf ( \o[17]_b1 , \7112_b1 );
buf ( \o[17]_b0 , \7112_b0 );
buf ( \o[16]_b1 , \7118_b1 );
buf ( \o[16]_b0 , \7118_b0 );
buf ( \o[15]_b1 , \7132_b1 );
buf ( \o[15]_b0 , \7132_b0 );
buf ( \o[14]_b1 , \7138_b1 );
buf ( \o[14]_b0 , \7138_b0 );
buf ( \o[13]_b1 , \7147_b1 );
buf ( \o[13]_b0 , \7147_b0 );
buf ( \o[12]_b1 , \7154_b1 );
buf ( \o[12]_b0 , \7154_b0 );
buf ( \o[11]_b1 , \7171_b1 );
buf ( \o[11]_b0 , \7171_b0 );
buf ( \o[10]_b1 , \7178_b1 );
buf ( \o[10]_b0 , \7178_b0 );
buf ( \o[9]_b1 , \7188_b1 );
buf ( \o[9]_b0 , \7188_b0 );
buf ( \o[8]_b1 , \7194_b1 );
buf ( \o[8]_b0 , \7194_b0 );
buf ( \o[7]_b1 , \7215_b1 );
buf ( \o[7]_b0 , \7215_b0 );
buf ( \o[6]_b1 , \7207_b1 );
buf ( \o[6]_b0 , \7207_b0 );
buf ( \o[5]_b1 , \7210_b1 );
buf ( \o[5]_b0 , \7210_b0 );
buf ( \o[4]_b1 , \7211_b1 );
buf ( \o[4]_b0 , \7211_b0 );
buf ( \o[3]_b1 , \7212_b1 );
buf ( \o[3]_b0 , \7212_b0 );
buf ( \o[2]_b1 , \7213_b1 );
buf ( \o[2]_b0 , \7213_b0 );
buf ( \o[1]_b1 , \7203_b1 );
buf ( \o[1]_b0 , \7203_b0 );
buf ( \o[0]_b1 , \7204_b1 );
buf ( \o[0]_b0 , \7204_b0 );
buf ( \99_b1 , \a[7]_b1 );
not ( \99_b1 , w_0 );
not ( \99_b0 , w_1 );
and ( w_0 , w_1 , \a[7]_b0 );
buf ( \100_b1 , \d[7]_b1 );
not ( \100_b1 , w_2 );
not ( \100_b0 , w_3 );
and ( w_2 , w_3 , \d[7]_b0 );
or ( \101_b1 , \99_b1 , \100_b1 );
not ( \100_b1 , w_4 );
and ( \101_b0 , \99_b0 , w_5 );
and ( w_4 , w_5 , \100_b0 );
or ( \102_b1 , \a[0]_b1 , \b[9]_b1 );
xor ( \102_b0 , \a[0]_b0 , w_6 );
not ( w_6 , w_7 );
and ( w_7 , \b[9]_b1 , \b[9]_b0 );
buf ( \103_b1 , \102_b1 );
not ( \103_b1 , w_8 );
not ( \103_b0 , w_9 );
and ( w_8 , w_9 , \102_b0 );
or ( \104_b1 , \b[8]_b1 , \b[7]_b1 );
xor ( \104_b0 , \b[8]_b0 , w_10 );
not ( w_10 , w_11 );
and ( w_11 , \b[7]_b1 , \b[7]_b0 );
or ( \105_b1 , \b[9]_b1 , w_12 );
xor ( \105_b0 , \b[9]_b0 , w_14 );
not ( w_14 , w_15 );
and ( w_15 , w_12 , w_13 );
buf ( w_12 , \b[8]_b1 );
not ( w_12 , w_16 );
not ( w_13 , w_17 );
and ( w_16 , w_17 , \b[8]_b0 );
or ( \106_b1 , \104_b1 , w_19 );
not ( w_19 , w_20 );
and ( \106_b0 , \104_b0 , w_21 );
and ( w_20 ,  , w_21 );
buf ( w_19 , \105_b1 );
not ( w_19 , w_22 );
not (  , w_23 );
and ( w_22 , w_23 , \105_b0 );
buf ( \107_b1 , \106_b1 );
not ( \107_b1 , w_24 );
not ( \107_b0 , w_25 );
and ( w_24 , w_25 , \106_b0 );
or ( \108_b1 , \103_b1 , w_26 );
or ( \108_b0 , \103_b0 , \107_b0 );
not ( \107_b0 , w_27 );
and ( w_27 , w_26 , \107_b1 );
or ( \109_b1 , \a[1]_b1 , \b[9]_b1 );
xor ( \109_b0 , \a[1]_b0 , w_28 );
not ( w_28 , w_29 );
and ( w_29 , \b[9]_b1 , \b[9]_b0 );
or ( \110_b1 , \104_b1 , w_31 );
not ( w_31 , w_32 );
and ( \110_b0 , \104_b0 , w_33 );
and ( w_32 ,  , w_33 );
buf ( w_31 , \109_b1 );
not ( w_31 , w_34 );
not (  , w_35 );
and ( w_34 , w_35 , \109_b0 );
or ( \111_b1 , \108_b1 , w_37 );
not ( w_37 , w_38 );
and ( \111_b0 , \108_b0 , w_39 );
and ( w_38 ,  , w_39 );
buf ( w_37 , \110_b1 );
not ( w_37 , w_40 );
not (  , w_41 );
and ( w_40 , w_41 , \110_b0 );
or ( \112_b1 , \a[0]_b1 , w_42 );
or ( \112_b0 , \a[0]_b0 , \b[8]_b0 );
not ( \b[8]_b0 , w_43 );
and ( w_43 , w_42 , \b[8]_b1 );
or ( \113_b1 , \112_b1 , w_45 );
not ( w_45 , w_46 );
and ( \113_b0 , \112_b0 , w_47 );
and ( w_46 ,  , w_47 );
buf ( w_45 , \b[7]_b1 );
not ( w_45 , w_48 );
not (  , w_49 );
and ( w_48 , w_49 , \b[7]_b0 );
or ( \114_b1 , \a[0]_b1 , w_51 );
not ( w_51 , w_52 );
and ( \114_b0 , \a[0]_b0 , w_53 );
and ( w_52 ,  , w_53 );
buf ( w_51 , \b[8]_b1 );
not ( w_51 , w_54 );
not (  , w_55 );
and ( w_54 , w_55 , \b[8]_b0 );
or ( \116_b1 , \a[4]_b1 , \b[5]_b1 );
xor ( \116_b0 , \a[4]_b0 , w_56 );
not ( w_56 , w_57 );
and ( w_57 , \b[5]_b1 , \b[5]_b0 );
or ( \117_b1 , \b[5]_b1 , \b[4]_b1 );
xor ( \117_b0 , \b[5]_b0 , w_58 );
not ( w_58 , w_59 );
and ( w_59 , \b[4]_b1 , \b[4]_b0 );
or ( \118_b1 , \116_b1 , w_61 );
not ( w_61 , w_62 );
and ( \118_b0 , \116_b0 , w_63 );
and ( w_62 ,  , w_63 );
buf ( w_61 , \117_b1 );
not ( w_61 , w_64 );
not (  , w_65 );
and ( w_64 , w_65 , \117_b0 );
or ( \119_b1 , \b[4]_b1 , \b[3]_b1 );
xor ( \119_b0 , \b[4]_b0 , w_66 );
not ( w_66 , w_67 );
and ( w_67 , \b[3]_b1 , \b[3]_b0 );
or ( \120_b1 , \118_b1 , w_68 );
or ( \120_b0 , \118_b0 , \119_b0 );
not ( \119_b0 , w_69 );
and ( w_69 , w_68 , \119_b1 );
or ( \121_b1 , \b[4]_b1 , \b[3]_b1 );
xor ( \121_b0 , \b[4]_b0 , w_70 );
not ( w_70 , w_71 );
and ( w_71 , \b[3]_b1 , \b[3]_b0 );
or ( \122_b1 , \a[5]_b1 , \b[5]_b1 );
xor ( \122_b0 , \a[5]_b0 , w_72 );
not ( w_72 , w_73 );
and ( w_73 , \b[5]_b1 , \b[5]_b0 );
or ( \123_b1 , \121_b1 , w_75 );
not ( w_75 , w_76 );
and ( \123_b0 , \121_b0 , w_77 );
and ( w_76 ,  , w_77 );
buf ( w_75 , \122_b1 );
not ( w_75 , w_78 );
not (  , w_79 );
and ( w_78 , w_79 , \122_b0 );
or ( \124_b1 , \120_b1 , w_81 );
not ( w_81 , w_82 );
and ( \124_b0 , \120_b0 , w_83 );
and ( w_82 ,  , w_83 );
buf ( w_81 , \123_b1 );
not ( w_81 , w_84 );
not (  , w_85 );
and ( w_84 , w_85 , \123_b0 );
or ( \125_b1 , \115_b1 , \124_b1 );
xor ( \125_b0 , \115_b0 , w_86 );
not ( w_86 , w_87 );
and ( w_87 , \124_b1 , \124_b0 );
or ( \126_b1 , \111_b1 , \125_b1 );
xor ( \126_b0 , \111_b0 , w_88 );
not ( w_88 , w_89 );
and ( w_89 , \125_b1 , \125_b0 );
or ( \127_b1 , \104_b1 , w_91 );
not ( w_91 , w_92 );
and ( \127_b0 , \104_b0 , w_93 );
and ( w_92 ,  , w_93 );
buf ( w_91 , \a[0]_b1 );
not ( w_91 , w_94 );
not (  , w_95 );
and ( w_94 , w_95 , \a[0]_b0 );
buf ( \128_b1 , \127_b1 );
not ( \128_b1 , w_96 );
not ( \128_b0 , w_97 );
and ( w_96 , w_97 , \127_b0 );
or ( \129_b1 , \a[7]_b1 , \b[1]_b1 );
xor ( \129_b0 , \a[7]_b0 , w_98 );
not ( w_98 , w_99 );
and ( w_99 , \b[1]_b1 , \b[1]_b0 );
buf ( \130_b1 , \129_b1 );
not ( \130_b1 , w_100 );
not ( \130_b0 , w_101 );
and ( w_100 , w_101 , \129_b0 );
buf ( \131_b1 , \b[0]_b1 );
not ( \131_b1 , w_102 );
not ( \131_b0 , w_103 );
and ( w_102 , w_103 , \b[0]_b0 );
or ( \132_b1 , \131_b1 , w_105 );
not ( w_105 , w_106 );
and ( \132_b0 , \131_b0 , w_107 );
and ( w_106 ,  , w_107 );
buf ( w_105 , \b[1]_b1 );
not ( w_105 , w_108 );
not (  , w_109 );
and ( w_108 , w_109 , \b[1]_b0 );
buf ( \133_b1 , \132_b1 );
not ( \133_b1 , w_110 );
not ( \133_b0 , w_111 );
and ( w_110 , w_111 , \132_b0 );
buf ( \134_b1 , \133_b1 );
not ( \134_b1 , w_112 );
not ( \134_b0 , w_113 );
and ( w_112 , w_113 , \133_b0 );
or ( \135_b1 , \130_b1 , w_114 );
or ( \135_b0 , \130_b0 , \134_b0 );
not ( \134_b0 , w_115 );
and ( w_115 , w_114 , \134_b1 );
or ( \136_b1 , \b[1]_b1 , \a[8]_b1 );
xor ( \136_b0 , \b[1]_b0 , w_116 );
not ( w_116 , w_117 );
and ( w_117 , \a[8]_b1 , \a[8]_b0 );
or ( \137_b1 , \136_b1 , w_119 );
not ( w_119 , w_120 );
and ( \137_b0 , \136_b0 , w_121 );
and ( w_120 ,  , w_121 );
buf ( w_119 , \b[0]_b1 );
not ( w_119 , w_122 );
not (  , w_123 );
and ( w_122 , w_123 , \b[0]_b0 );
or ( \138_b1 , \135_b1 , w_125 );
not ( w_125 , w_126 );
and ( \138_b0 , \135_b0 , w_127 );
and ( w_126 ,  , w_127 );
buf ( w_125 , \137_b1 );
not ( w_125 , w_128 );
not (  , w_129 );
and ( w_128 , w_129 , \137_b0 );
or ( \139_b1 , \128_b1 , w_130 );
or ( \139_b0 , \128_b0 , \138_b0 );
not ( \138_b0 , w_131 );
and ( w_131 , w_130 , \138_b1 );
buf ( \140_b1 , \139_b1 );
not ( \140_b1 , w_132 );
not ( \140_b0 , w_133 );
and ( w_132 , w_133 , \139_b0 );
or ( \141_b1 , \a[5]_b1 , \b[3]_b1 );
xor ( \141_b0 , \a[5]_b0 , w_134 );
not ( w_134 , w_135 );
and ( w_135 , \b[3]_b1 , \b[3]_b0 );
buf ( \142_b1 , \141_b1 );
not ( \142_b1 , w_136 );
not ( \142_b0 , w_137 );
and ( w_136 , w_137 , \141_b0 );
or ( \143_b1 , \b[3]_b1 , w_138 );
xor ( \143_b0 , \b[3]_b0 , w_140 );
not ( w_140 , w_141 );
and ( w_141 , w_138 , w_139 );
buf ( w_138 , \b[2]_b1 );
not ( w_138 , w_142 );
not ( w_139 , w_143 );
and ( w_142 , w_143 , \b[2]_b0 );
or ( \144_b1 , \b[2]_b1 , \b[1]_b1 );
xor ( \144_b0 , \b[2]_b0 , w_144 );
not ( w_144 , w_145 );
and ( w_145 , \b[1]_b1 , \b[1]_b0 );
or ( \145_b1 , \143_b1 , w_147 );
not ( w_147 , w_148 );
and ( \145_b0 , \143_b0 , w_149 );
and ( w_148 ,  , w_149 );
buf ( w_147 , \144_b1 );
not ( w_147 , w_150 );
not (  , w_151 );
and ( w_150 , w_151 , \144_b0 );
buf ( \146_b1 , \145_b1 );
not ( \146_b1 , w_152 );
not ( \146_b0 , w_153 );
and ( w_152 , w_153 , \145_b0 );
buf ( \147_b1 , \146_b1 );
not ( \147_b1 , w_154 );
not ( \147_b0 , w_155 );
and ( w_154 , w_155 , \146_b0 );
buf ( \148_b1 , \147_b1 );
not ( \148_b1 , w_156 );
not ( \148_b0 , w_157 );
and ( w_156 , w_157 , \147_b0 );
or ( \149_b1 , \142_b1 , w_158 );
or ( \149_b0 , \142_b0 , \148_b0 );
not ( \148_b0 , w_159 );
and ( w_159 , w_158 , \148_b1 );
or ( \150_b1 , \b[2]_b1 , \b[1]_b1 );
xor ( \150_b0 , \b[2]_b0 , w_160 );
not ( w_160 , w_161 );
and ( w_161 , \b[1]_b1 , \b[1]_b0 );
or ( \151_b1 , \a[6]_b1 , \b[3]_b1 );
xor ( \151_b0 , \a[6]_b0 , w_162 );
not ( w_162 , w_163 );
and ( w_163 , \b[3]_b1 , \b[3]_b0 );
or ( \152_b1 , \150_b1 , w_165 );
not ( w_165 , w_166 );
and ( \152_b0 , \150_b0 , w_167 );
and ( w_166 ,  , w_167 );
buf ( w_165 , \151_b1 );
not ( w_165 , w_168 );
not (  , w_169 );
and ( w_168 , w_169 , \151_b0 );
or ( \153_b1 , \149_b1 , w_171 );
not ( w_171 , w_172 );
and ( \153_b0 , \149_b0 , w_173 );
and ( w_172 ,  , w_173 );
buf ( w_171 , \152_b1 );
not ( w_171 , w_174 );
not (  , w_175 );
and ( w_174 , w_175 , \152_b0 );
buf ( \154_b1 , \153_b1 );
not ( \154_b1 , w_176 );
not ( \154_b0 , w_177 );
and ( w_176 , w_177 , \153_b0 );
or ( \155_b1 , \140_b1 , w_178 );
or ( \155_b0 , \140_b0 , \154_b0 );
not ( \154_b0 , w_179 );
and ( w_179 , w_178 , \154_b1 );
or ( \156_b1 , \138_b1 , w_181 );
not ( w_181 , w_182 );
and ( \156_b0 , \138_b0 , w_183 );
and ( w_182 ,  , w_183 );
buf ( w_181 , \128_b1 );
not ( w_181 , w_184 );
not (  , w_185 );
and ( w_184 , w_185 , \128_b0 );
or ( \157_b1 , \155_b1 , w_187 );
not ( w_187 , w_188 );
and ( \157_b0 , \155_b0 , w_189 );
and ( w_188 ,  , w_189 );
buf ( w_187 , \156_b1 );
not ( w_187 , w_190 );
not (  , w_191 );
and ( w_190 , w_191 , \156_b0 );
or ( \158_b1 , \126_b1 , w_192 );
xor ( \158_b0 , \126_b0 , w_194 );
not ( w_194 , w_195 );
and ( w_195 , w_192 , w_193 );
buf ( w_192 , \157_b1 );
not ( w_192 , w_196 );
not ( w_193 , w_197 );
and ( w_196 , w_197 , \157_b0 );
buf ( \159_b1 , \158_b1 );
not ( \159_b1 , w_198 );
not ( \159_b0 , w_199 );
and ( w_198 , w_199 , \158_b0 );
or ( \160_b1 , \a[9]_b1 , \b[1]_b1 );
xor ( \160_b0 , \a[9]_b0 , w_200 );
not ( w_200 , w_201 );
and ( w_201 , \b[1]_b1 , \b[1]_b0 );
or ( \161_b1 , \160_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_202 );
and ( \161_b0 , \160_b0 , w_203 );
and ( w_202 , w_203 , \b[0]_b0 );
buf ( \162_b1 , \b[1]_b1 );
not ( \162_b1 , w_204 );
not ( \162_b0 , w_205 );
and ( w_204 , w_205 , \b[1]_b0 );
or ( \163_b1 , \162_b1 , w_207 );
not ( w_207 , w_208 );
and ( \163_b0 , \162_b0 , w_209 );
and ( w_208 ,  , w_209 );
buf ( w_207 , \b[0]_b1 );
not ( w_207 , w_210 );
not (  , w_211 );
and ( w_210 , w_211 , \b[0]_b0 );
or ( \164_b1 , \163_b1 , \136_b1 );
not ( \136_b1 , w_212 );
and ( \164_b0 , \163_b0 , w_213 );
and ( w_212 , w_213 , \136_b0 );
or ( \165_b1 , \161_b1 , w_215 );
not ( w_215 , w_216 );
and ( \165_b0 , \161_b0 , w_217 );
and ( w_216 ,  , w_217 );
buf ( w_215 , \164_b1 );
not ( w_215 , w_218 );
not (  , w_219 );
and ( w_218 , w_219 , \164_b0 );
buf ( \166_b1 , \151_b1 );
not ( \166_b1 , w_220 );
not ( \166_b0 , w_221 );
and ( w_220 , w_221 , \151_b0 );
buf ( \167_b1 , \145_b1 );
not ( \167_b1 , w_222 );
not ( \167_b0 , w_223 );
and ( w_222 , w_223 , \145_b0 );
or ( \168_b1 , \166_b1 , w_224 );
or ( \168_b0 , \166_b0 , \167_b0 );
not ( \167_b0 , w_225 );
and ( w_225 , w_224 , \167_b1 );
or ( \169_b1 , \a[7]_b1 , \b[3]_b1 );
xor ( \169_b0 , \a[7]_b0 , w_226 );
not ( w_226 , w_227 );
and ( w_227 , \b[3]_b1 , \b[3]_b0 );
or ( \170_b1 , \150_b1 , w_229 );
not ( w_229 , w_230 );
and ( \170_b0 , \150_b0 , w_231 );
and ( w_230 ,  , w_231 );
buf ( w_229 , \169_b1 );
not ( w_229 , w_232 );
not (  , w_233 );
and ( w_232 , w_233 , \169_b0 );
or ( \171_b1 , \168_b1 , w_235 );
not ( w_235 , w_236 );
and ( \171_b0 , \168_b0 , w_237 );
and ( w_236 ,  , w_237 );
buf ( w_235 , \170_b1 );
not ( w_235 , w_238 );
not (  , w_239 );
and ( w_238 , w_239 , \170_b0 );
or ( \172_b1 , \165_b1 , \171_b1 );
xor ( \172_b0 , \165_b0 , w_240 );
not ( w_240 , w_241 );
and ( w_241 , \171_b1 , \171_b0 );
or ( \173_b1 , \a[2]_b1 , \b[7]_b1 );
xor ( \173_b0 , \a[2]_b0 , w_242 );
not ( w_242 , w_243 );
and ( w_243 , \b[7]_b1 , \b[7]_b0 );
buf ( \174_b1 , \173_b1 );
not ( \174_b1 , w_244 );
not ( \174_b0 , w_245 );
and ( w_244 , w_245 , \173_b0 );
or ( \175_b1 , \b[7]_b1 , \b[6]_b1 );
xor ( \175_b0 , \b[7]_b0 , w_246 );
not ( w_246 , w_247 );
and ( w_247 , \b[6]_b1 , \b[6]_b0 );
buf ( \176_b1 , \175_b1 );
not ( \176_b1 , w_248 );
not ( \176_b0 , w_249 );
and ( w_248 , w_249 , \175_b0 );
or ( \177_b1 , \b[6]_b1 , \b[5]_b1 );
xor ( \177_b0 , \b[6]_b0 , w_250 );
not ( w_250 , w_251 );
and ( w_251 , \b[5]_b1 , \b[5]_b0 );
or ( \178_b1 , \176_b1 , w_253 );
not ( w_253 , w_254 );
and ( \178_b0 , \176_b0 , w_255 );
and ( w_254 ,  , w_255 );
buf ( w_253 , \177_b1 );
not ( w_253 , w_256 );
not (  , w_257 );
and ( w_256 , w_257 , \177_b0 );
buf ( \179_b1 , \178_b1 );
not ( \179_b1 , w_258 );
not ( \179_b0 , w_259 );
and ( w_258 , w_259 , \178_b0 );
or ( \180_b1 , \174_b1 , w_260 );
or ( \180_b0 , \174_b0 , \179_b0 );
not ( \179_b0 , w_261 );
and ( w_261 , w_260 , \179_b1 );
or ( \181_b1 , \a[3]_b1 , \b[7]_b1 );
xor ( \181_b0 , \a[3]_b0 , w_262 );
not ( w_262 , w_263 );
and ( w_263 , \b[7]_b1 , \b[7]_b0 );
or ( \182_b1 , \177_b1 , w_265 );
not ( w_265 , w_266 );
and ( \182_b0 , \177_b0 , w_267 );
and ( w_266 ,  , w_267 );
buf ( w_265 , \181_b1 );
not ( w_265 , w_268 );
not (  , w_269 );
and ( w_268 , w_269 , \181_b0 );
or ( \183_b1 , \180_b1 , w_271 );
not ( w_271 , w_272 );
and ( \183_b0 , \180_b0 , w_273 );
and ( w_272 ,  , w_273 );
buf ( w_271 , \182_b1 );
not ( w_271 , w_274 );
not (  , w_275 );
and ( w_274 , w_275 , \182_b0 );
buf ( \184_b1 , \183_b1 );
not ( \184_b1 , w_276 );
not ( \184_b0 , w_277 );
and ( w_276 , w_277 , \183_b0 );
or ( \185_b1 , \172_b1 , w_278 );
xor ( \185_b0 , \172_b0 , w_280 );
not ( w_280 , w_281 );
and ( w_281 , w_278 , w_279 );
buf ( w_278 , \184_b1 );
not ( w_278 , w_282 );
not ( w_279 , w_283 );
and ( w_282 , w_283 , \184_b0 );
buf ( \186_b1 , \185_b1 );
buf ( \186_b0 , \185_b0 );
buf ( \187_b1 , \186_b1 );
not ( \187_b1 , w_284 );
not ( \187_b0 , w_285 );
and ( w_284 , w_285 , \186_b0 );
or ( \188_b1 , \159_b1 , w_286 );
or ( \188_b0 , \159_b0 , \187_b0 );
not ( \187_b0 , w_287 );
and ( w_287 , w_286 , \187_b1 );
or ( \189_b1 , \a[1]_b1 , \b[7]_b1 );
xor ( \189_b0 , \a[1]_b0 , w_288 );
not ( w_288 , w_289 );
and ( w_289 , \b[7]_b1 , \b[7]_b0 );
buf ( \190_b1 , \189_b1 );
not ( \190_b1 , w_290 );
not ( \190_b0 , w_291 );
and ( w_290 , w_291 , \189_b0 );
buf ( \191_b1 , \178_b1 );
not ( \191_b1 , w_292 );
not ( \191_b0 , w_293 );
and ( w_292 , w_293 , \178_b0 );
or ( \192_b1 , \190_b1 , w_294 );
or ( \192_b0 , \190_b0 , \191_b0 );
not ( \191_b0 , w_295 );
and ( w_295 , w_294 , \191_b1 );
or ( \193_b1 , \173_b1 , w_297 );
not ( w_297 , w_298 );
and ( \193_b0 , \173_b0 , w_299 );
and ( w_298 ,  , w_299 );
buf ( w_297 , \177_b1 );
not ( w_297 , w_300 );
not (  , w_301 );
and ( w_300 , w_301 , \177_b0 );
or ( \194_b1 , \192_b1 , w_303 );
not ( w_303 , w_304 );
and ( \194_b0 , \192_b0 , w_305 );
and ( w_304 ,  , w_305 );
buf ( w_303 , \193_b1 );
not ( w_303 , w_306 );
not (  , w_307 );
and ( w_306 , w_307 , \193_b0 );
or ( \195_b1 , \a[3]_b1 , \b[5]_b1 );
xor ( \195_b0 , \a[3]_b0 , w_308 );
not ( w_308 , w_309 );
and ( w_309 , \b[5]_b1 , \b[5]_b0 );
buf ( \196_b1 , \195_b1 );
not ( \196_b1 , w_310 );
not ( \196_b0 , w_311 );
and ( w_310 , w_311 , \195_b0 );
buf ( \197_b1 , \117_b1 );
not ( \197_b1 , w_312 );
not ( \197_b0 , w_313 );
and ( w_312 , w_313 , \117_b0 );
or ( \198_b1 , \197_b1 , w_315 );
not ( w_315 , w_316 );
and ( \198_b0 , \197_b0 , w_317 );
and ( w_316 ,  , w_317 );
buf ( w_315 , \121_b1 );
not ( w_315 , w_318 );
not (  , w_319 );
and ( w_318 , w_319 , \121_b0 );
buf ( \199_b1 , \198_b1 );
not ( \199_b1 , w_320 );
not ( \199_b0 , w_321 );
and ( w_320 , w_321 , \198_b0 );
or ( \200_b1 , \196_b1 , w_322 );
or ( \200_b0 , \196_b0 , \199_b0 );
not ( \199_b0 , w_323 );
and ( w_323 , w_322 , \199_b1 );
or ( \201_b1 , \121_b1 , w_325 );
not ( w_325 , w_326 );
and ( \201_b0 , \121_b0 , w_327 );
and ( w_326 ,  , w_327 );
buf ( w_325 , \116_b1 );
not ( w_325 , w_328 );
not (  , w_329 );
and ( w_328 , w_329 , \116_b0 );
or ( \202_b1 , \200_b1 , w_331 );
not ( w_331 , w_332 );
and ( \202_b0 , \200_b0 , w_333 );
and ( w_332 ,  , w_333 );
buf ( w_331 , \201_b1 );
not ( w_331 , w_334 );
not (  , w_335 );
and ( w_334 , w_335 , \201_b0 );
or ( \203_b1 , \194_b1 , \202_b1 );
xor ( \203_b0 , \194_b0 , w_336 );
not ( w_336 , w_337 );
and ( w_337 , \202_b1 , \202_b0 );
or ( \204_b1 , \a[0]_b1 , w_338 );
or ( \204_b0 , \a[0]_b0 , \b[6]_b0 );
not ( \b[6]_b0 , w_339 );
and ( w_339 , w_338 , \b[6]_b1 );
or ( \205_b1 , \204_b1 , w_341 );
not ( w_341 , w_342 );
and ( \205_b0 , \204_b0 , w_343 );
and ( w_342 ,  , w_343 );
buf ( w_341 , \b[5]_b1 );
not ( w_341 , w_344 );
not (  , w_345 );
and ( w_344 , w_345 , \b[5]_b0 );
or ( \206_b1 , \a[0]_b1 , w_347 );
not ( w_347 , w_348 );
and ( \206_b0 , \a[0]_b0 , w_349 );
and ( w_348 ,  , w_349 );
buf ( w_347 , \b[6]_b1 );
not ( w_347 , w_350 );
not (  , w_351 );
and ( w_350 , w_351 , \b[6]_b0 );
buf ( \208_b1 , \141_b1 );
not ( \208_b1 , w_352 );
not ( \208_b0 , w_353 );
and ( w_352 , w_353 , \141_b0 );
buf ( \209_b1 , \150_b1 );
not ( \209_b1 , w_354 );
not ( \209_b0 , w_355 );
and ( w_354 , w_355 , \150_b0 );
or ( \210_b1 , \208_b1 , w_356 );
or ( \210_b0 , \208_b0 , \209_b0 );
not ( \209_b0 , w_357 );
and ( w_357 , w_356 , \209_b1 );
buf ( \211_b1 , \144_b1 );
not ( \211_b1 , w_358 );
not ( \211_b0 , w_359 );
and ( w_358 , w_359 , \144_b0 );
or ( \212_b1 , \a[4]_b1 , w_360 );
xor ( \212_b0 , \a[4]_b0 , w_362 );
not ( w_362 , w_363 );
and ( w_363 , w_360 , w_361 );
buf ( w_360 , \b[3]_b1 );
not ( w_360 , w_364 );
not ( w_361 , w_365 );
and ( w_364 , w_365 , \b[3]_b0 );
or ( \213_b1 , \212_b1 , w_367 );
not ( w_367 , w_368 );
and ( \213_b0 , \212_b0 , w_369 );
and ( w_368 ,  , w_369 );
buf ( w_367 , \143_b1 );
not ( w_367 , w_370 );
not (  , w_371 );
and ( w_370 , w_371 , \143_b0 );
or ( \214_b1 , \211_b1 , w_373 );
not ( w_373 , w_374 );
and ( \214_b0 , \211_b0 , w_375 );
and ( w_374 ,  , w_375 );
buf ( w_373 , \213_b1 );
not ( w_373 , w_376 );
not (  , w_377 );
and ( w_376 , w_377 , \213_b0 );
or ( \215_b1 , \210_b1 , w_379 );
not ( w_379 , w_380 );
and ( \215_b0 , \210_b0 , w_381 );
and ( w_380 ,  , w_381 );
buf ( w_379 , \214_b1 );
not ( w_379 , w_382 );
not (  , w_383 );
and ( w_382 , w_383 , \214_b0 );
or ( \216_b1 , \207_b1 , \215_b1 );
not ( \215_b1 , w_384 );
and ( \216_b0 , \207_b0 , w_385 );
and ( w_384 , w_385 , \215_b0 );
or ( \217_b1 , \203_b1 , \216_b1 );
not ( \216_b1 , w_386 );
and ( \217_b0 , \203_b0 , w_387 );
and ( w_386 , w_387 , \216_b0 );
or ( \218_b1 , \194_b1 , \202_b1 );
not ( \202_b1 , w_388 );
and ( \218_b0 , \194_b0 , w_389 );
and ( w_388 , w_389 , \202_b0 );
or ( \219_b1 , \217_b1 , w_390 );
or ( \219_b0 , \217_b0 , \218_b0 );
not ( \218_b0 , w_391 );
and ( w_391 , w_390 , \218_b1 );
buf ( \220_b1 , \219_b1 );
buf ( \220_b0 , \219_b0 );
or ( \221_b1 , \188_b1 , w_393 );
not ( w_393 , w_394 );
and ( \221_b0 , \188_b0 , w_395 );
and ( w_394 ,  , w_395 );
buf ( w_393 , \220_b1 );
not ( w_393 , w_396 );
not (  , w_397 );
and ( w_396 , w_397 , \220_b0 );
buf ( \222_b1 , \186_b1 );
not ( \222_b1 , w_398 );
not ( \222_b0 , w_399 );
and ( w_398 , w_399 , \186_b0 );
buf ( \223_b1 , \158_b1 );
not ( \223_b1 , w_400 );
not ( \223_b0 , w_401 );
and ( w_400 , w_401 , \158_b0 );
or ( \224_b1 , \222_b1 , w_403 );
not ( w_403 , w_404 );
and ( \224_b0 , \222_b0 , w_405 );
and ( w_404 ,  , w_405 );
buf ( w_403 , \223_b1 );
not ( w_403 , w_406 );
not (  , w_407 );
and ( w_406 , w_407 , \223_b0 );
or ( \225_b1 , \221_b1 , w_409 );
not ( w_409 , w_410 );
and ( \225_b0 , \221_b0 , w_411 );
and ( w_410 ,  , w_411 );
buf ( w_409 , \224_b1 );
not ( w_409 , w_412 );
not (  , w_413 );
and ( w_412 , w_413 , \224_b0 );
buf ( \226_b1 , \225_b1 );
not ( \226_b1 , w_414 );
not ( \226_b0 , w_415 );
and ( w_414 , w_415 , \225_b0 );
buf ( \227_b1 , \109_b1 );
not ( \227_b1 , w_416 );
not ( \227_b0 , w_417 );
and ( w_416 , w_417 , \109_b0 );
or ( \228_b1 , \104_b1 , w_419 );
not ( w_419 , w_420 );
and ( \228_b0 , \104_b0 , w_421 );
and ( w_420 ,  , w_421 );
buf ( w_419 , \105_b1 );
not ( w_419 , w_422 );
not (  , w_423 );
and ( w_422 , w_423 , \105_b0 );
buf ( \229_b1 , \228_b1 );
not ( \229_b1 , w_424 );
not ( \229_b0 , w_425 );
and ( w_424 , w_425 , \228_b0 );
or ( \230_b1 , \227_b1 , w_426 );
or ( \230_b0 , \227_b0 , \229_b0 );
not ( \229_b0 , w_427 );
and ( w_427 , w_426 , \229_b1 );
or ( \231_b1 , \a[2]_b1 , \b[9]_b1 );
xor ( \231_b0 , \a[2]_b0 , w_428 );
not ( w_428 , w_429 );
and ( w_429 , \b[9]_b1 , \b[9]_b0 );
or ( \232_b1 , \104_b1 , w_431 );
not ( w_431 , w_432 );
and ( \232_b0 , \104_b0 , w_433 );
and ( w_432 ,  , w_433 );
buf ( w_431 , \231_b1 );
not ( w_431 , w_434 );
not (  , w_435 );
and ( w_434 , w_435 , \231_b0 );
or ( \233_b1 , \230_b1 , w_437 );
not ( w_437 , w_438 );
and ( \233_b0 , \230_b0 , w_439 );
and ( w_438 ,  , w_439 );
buf ( w_437 , \232_b1 );
not ( w_437 , w_440 );
not (  , w_441 );
and ( w_440 , w_441 , \232_b0 );
buf ( \234_b1 , \181_b1 );
not ( \234_b1 , w_442 );
not ( \234_b0 , w_443 );
and ( w_442 , w_443 , \181_b0 );
buf ( \235_b1 , \178_b1 );
not ( \235_b1 , w_444 );
not ( \235_b0 , w_445 );
and ( w_444 , w_445 , \178_b0 );
or ( \236_b1 , \234_b1 , w_446 );
or ( \236_b0 , \234_b0 , \235_b0 );
not ( \235_b0 , w_447 );
and ( w_447 , w_446 , \235_b1 );
or ( \237_b1 , \a[4]_b1 , \b[7]_b1 );
xor ( \237_b0 , \a[4]_b0 , w_448 );
not ( w_448 , w_449 );
and ( w_449 , \b[7]_b1 , \b[7]_b0 );
or ( \238_b1 , \177_b1 , w_451 );
not ( w_451 , w_452 );
and ( \238_b0 , \177_b0 , w_453 );
and ( w_452 ,  , w_453 );
buf ( w_451 , \237_b1 );
not ( w_451 , w_454 );
not (  , w_455 );
and ( w_454 , w_455 , \237_b0 );
or ( \239_b1 , \236_b1 , w_457 );
not ( w_457 , w_458 );
and ( \239_b0 , \236_b0 , w_459 );
and ( w_458 ,  , w_459 );
buf ( w_457 , \238_b1 );
not ( w_457 , w_460 );
not (  , w_461 );
and ( w_460 , w_461 , \238_b0 );
or ( \240_b1 , \233_b1 , \239_b1 );
xor ( \240_b0 , \233_b0 , w_462 );
not ( w_462 , w_463 );
and ( w_463 , \239_b1 , \239_b0 );
buf ( \241_b1 , \169_b1 );
not ( \241_b1 , w_464 );
not ( \241_b0 , w_465 );
and ( w_464 , w_465 , \169_b0 );
buf ( \242_b1 , \146_b1 );
not ( \242_b1 , w_466 );
not ( \242_b0 , w_467 );
and ( w_466 , w_467 , \146_b0 );
buf ( \243_b1 , \242_b1 );
not ( \243_b1 , w_468 );
not ( \243_b0 , w_469 );
and ( w_468 , w_469 , \242_b0 );
or ( \244_b1 , \241_b1 , w_470 );
or ( \244_b0 , \241_b0 , \243_b0 );
not ( \243_b0 , w_471 );
and ( w_471 , w_470 , \243_b1 );
or ( \245_b1 , \a[8]_b1 , \b[3]_b1 );
xor ( \245_b0 , \a[8]_b0 , w_472 );
not ( w_472 , w_473 );
and ( w_473 , \b[3]_b1 , \b[3]_b0 );
or ( \246_b1 , \150_b1 , w_475 );
not ( w_475 , w_476 );
and ( \246_b0 , \150_b0 , w_477 );
and ( w_476 ,  , w_477 );
buf ( w_475 , \245_b1 );
not ( w_475 , w_478 );
not (  , w_479 );
and ( w_478 , w_479 , \245_b0 );
or ( \247_b1 , \244_b1 , w_481 );
not ( w_481 , w_482 );
and ( \247_b0 , \244_b0 , w_483 );
and ( w_482 ,  , w_483 );
buf ( w_481 , \246_b1 );
not ( w_481 , w_484 );
not (  , w_485 );
and ( w_484 , w_485 , \246_b0 );
or ( \248_b1 , \240_b1 , \247_b1 );
xor ( \248_b0 , \240_b0 , w_486 );
not ( w_486 , w_487 );
and ( w_487 , \247_b1 , \247_b0 );
buf ( \249_b1 , \111_b1 );
not ( \249_b1 , w_488 );
not ( \249_b0 , w_489 );
and ( w_488 , w_489 , \111_b0 );
buf ( \250_b1 , \125_b1 );
not ( \250_b1 , w_490 );
not ( \250_b0 , w_491 );
and ( w_490 , w_491 , \125_b0 );
or ( \251_b1 , \249_b1 , w_492 );
or ( \251_b0 , \249_b0 , \250_b0 );
not ( \250_b0 , w_493 );
and ( w_493 , w_492 , \250_b1 );
or ( \252_b1 , \125_b1 , w_494 );
or ( \252_b0 , \125_b0 , \111_b0 );
not ( \111_b0 , w_495 );
and ( w_495 , w_494 , \111_b1 );
or ( \253_b1 , \252_b1 , w_497 );
not ( w_497 , w_498 );
and ( \253_b0 , \252_b0 , w_499 );
and ( w_498 ,  , w_499 );
buf ( w_497 , \157_b1 );
not ( w_497 , w_500 );
not (  , w_501 );
and ( w_500 , w_501 , \157_b0 );
or ( \254_b1 , \251_b1 , w_503 );
not ( w_503 , w_504 );
and ( \254_b0 , \251_b0 , w_505 );
and ( w_504 ,  , w_505 );
buf ( w_503 , \253_b1 );
not ( w_503 , w_506 );
not (  , w_507 );
and ( w_506 , w_507 , \253_b0 );
or ( \255_b1 , \248_b1 , \254_b1 );
xor ( \255_b0 , \248_b0 , w_508 );
not ( w_508 , w_509 );
and ( w_509 , \254_b1 , \254_b0 );
or ( \256_b1 , \115_b1 , \124_b1 );
not ( \124_b1 , w_510 );
and ( \256_b0 , \115_b0 , w_511 );
and ( w_510 , w_511 , \124_b0 );
or ( \257_b1 , \b[10]_b1 , \b[9]_b1 );
xor ( \257_b0 , \b[10]_b0 , w_512 );
not ( w_512 , w_513 );
and ( w_513 , \b[9]_b1 , \b[9]_b0 );
or ( \258_b1 , \257_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_514 );
and ( \258_b0 , \257_b0 , w_515 );
and ( w_514 , w_515 , \a[0]_b0 );
buf ( \259_b1 , \160_b1 );
not ( \259_b1 , w_516 );
not ( \259_b0 , w_517 );
and ( w_516 , w_517 , \160_b0 );
buf ( \260_b1 , \163_b1 );
not ( \260_b1 , w_518 );
not ( \260_b0 , w_519 );
and ( w_518 , w_519 , \163_b0 );
or ( \261_b1 , \259_b1 , w_520 );
or ( \261_b0 , \259_b0 , \260_b0 );
not ( \260_b0 , w_521 );
and ( w_521 , w_520 , \260_b1 );
or ( \262_b1 , \a[10]_b1 , \b[1]_b1 );
xor ( \262_b0 , \a[10]_b0 , w_522 );
not ( w_522 , w_523 );
and ( w_523 , \b[1]_b1 , \b[1]_b0 );
or ( \263_b1 , \b[0]_b1 , w_525 );
not ( w_525 , w_526 );
and ( \263_b0 , \b[0]_b0 , w_527 );
and ( w_526 ,  , w_527 );
buf ( w_525 , \262_b1 );
not ( w_525 , w_528 );
not (  , w_529 );
and ( w_528 , w_529 , \262_b0 );
or ( \264_b1 , \261_b1 , w_531 );
not ( w_531 , w_532 );
and ( \264_b0 , \261_b0 , w_533 );
and ( w_532 ,  , w_533 );
buf ( w_531 , \263_b1 );
not ( w_531 , w_534 );
not (  , w_535 );
and ( w_534 , w_535 , \263_b0 );
or ( \265_b1 , \258_b1 , \264_b1 );
xor ( \265_b0 , \258_b0 , w_536 );
not ( w_536 , w_537 );
and ( w_537 , \264_b1 , \264_b0 );
buf ( \266_b1 , \122_b1 );
not ( \266_b1 , w_538 );
not ( \266_b0 , w_539 );
and ( w_538 , w_539 , \122_b0 );
or ( \267_b1 , \119_b1 , w_541 );
not ( w_541 , w_542 );
and ( \267_b0 , \119_b0 , w_543 );
and ( w_542 ,  , w_543 );
buf ( w_541 , \197_b1 );
not ( w_541 , w_544 );
not (  , w_545 );
and ( w_544 , w_545 , \197_b0 );
buf ( \268_b1 , \267_b1 );
not ( \268_b1 , w_546 );
not ( \268_b0 , w_547 );
and ( w_546 , w_547 , \267_b0 );
or ( \269_b1 , \266_b1 , w_548 );
or ( \269_b0 , \266_b0 , \268_b0 );
not ( \268_b0 , w_549 );
and ( w_549 , w_548 , \268_b1 );
or ( \270_b1 , \a[6]_b1 , \b[5]_b1 );
xor ( \270_b0 , \a[6]_b0 , w_550 );
not ( w_550 , w_551 );
and ( w_551 , \b[5]_b1 , \b[5]_b0 );
or ( \271_b1 , \121_b1 , w_553 );
not ( w_553 , w_554 );
and ( \271_b0 , \121_b0 , w_555 );
and ( w_554 ,  , w_555 );
buf ( w_553 , \270_b1 );
not ( w_553 , w_556 );
not (  , w_557 );
and ( w_556 , w_557 , \270_b0 );
or ( \272_b1 , \269_b1 , w_559 );
not ( w_559 , w_560 );
and ( \272_b0 , \269_b0 , w_561 );
and ( w_560 ,  , w_561 );
buf ( w_559 , \271_b1 );
not ( w_559 , w_562 );
not (  , w_563 );
and ( w_562 , w_563 , \271_b0 );
or ( \273_b1 , \265_b1 , \272_b1 );
xor ( \273_b0 , \265_b0 , w_564 );
not ( w_564 , w_565 );
and ( w_565 , \272_b1 , \272_b0 );
or ( \274_b1 , \256_b1 , \273_b1 );
xor ( \274_b0 , \256_b0 , w_566 );
not ( w_566 , w_567 );
and ( w_567 , \273_b1 , \273_b0 );
buf ( \275_b1 , \165_b1 );
not ( \275_b1 , w_568 );
not ( \275_b0 , w_569 );
and ( w_568 , w_569 , \165_b0 );
buf ( \276_b1 , \184_b1 );
not ( \276_b1 , w_570 );
not ( \276_b0 , w_571 );
and ( w_570 , w_571 , \184_b0 );
or ( \277_b1 , \275_b1 , w_572 );
or ( \277_b0 , \275_b0 , \276_b0 );
not ( \276_b0 , w_573 );
and ( w_573 , w_572 , \276_b1 );
or ( \278_b1 , \277_b1 , w_575 );
not ( w_575 , w_576 );
and ( \278_b0 , \277_b0 , w_577 );
and ( w_576 ,  , w_577 );
buf ( w_575 , \171_b1 );
not ( w_575 , w_578 );
not (  , w_579 );
and ( w_578 , w_579 , \171_b0 );
buf ( \279_b1 , \165_b1 );
not ( \279_b1 , w_580 );
not ( \279_b0 , w_581 );
and ( w_580 , w_581 , \165_b0 );
or ( \280_b1 , \279_b1 , w_583 );
not ( w_583 , w_584 );
and ( \280_b0 , \279_b0 , w_585 );
and ( w_584 ,  , w_585 );
buf ( w_583 , \183_b1 );
not ( w_583 , w_586 );
not (  , w_587 );
and ( w_586 , w_587 , \183_b0 );
or ( \281_b1 , \278_b1 , w_589 );
not ( w_589 , w_590 );
and ( \281_b0 , \278_b0 , w_591 );
and ( w_590 ,  , w_591 );
buf ( w_589 , \280_b1 );
not ( w_589 , w_592 );
not (  , w_593 );
and ( w_592 , w_593 , \280_b0 );
or ( \282_b1 , \274_b1 , \281_b1 );
xor ( \282_b0 , \274_b0 , w_594 );
not ( w_594 , w_595 );
and ( w_595 , \281_b1 , \281_b0 );
or ( \283_b1 , \255_b1 , w_596 );
xor ( \283_b0 , \255_b0 , w_598 );
not ( w_598 , w_599 );
and ( w_599 , w_596 , w_597 );
buf ( w_596 , \282_b1 );
not ( w_596 , w_600 );
not ( w_597 , w_601 );
and ( w_600 , w_601 , \282_b0 );
or ( \284_b1 , \226_b1 , w_603 );
not ( w_603 , w_604 );
and ( \284_b0 , \226_b0 , w_605 );
and ( w_604 ,  , w_605 );
buf ( w_603 , \283_b1 );
not ( w_603 , w_606 );
not (  , w_607 );
and ( w_606 , w_607 , \283_b0 );
buf ( \285_b1 , \284_b1 );
not ( \285_b1 , w_608 );
not ( \285_b0 , w_609 );
and ( w_608 , w_609 , \284_b0 );
buf ( \286_b1 , \219_b1 );
not ( \286_b1 , w_610 );
not ( \286_b0 , w_611 );
and ( w_610 , w_611 , \219_b0 );
buf ( \287_b1 , \185_b1 );
not ( \287_b1 , w_612 );
not ( \287_b0 , w_613 );
and ( w_612 , w_613 , \185_b0 );
or ( \288_b1 , \286_b1 , \287_b1 );
not ( \287_b1 , w_614 );
and ( \288_b0 , \286_b0 , w_615 );
and ( w_614 , w_615 , \287_b0 );
or ( \289_b1 , \219_b1 , \185_b1 );
not ( \185_b1 , w_616 );
and ( \289_b0 , \219_b0 , w_617 );
and ( w_616 , w_617 , \185_b0 );
or ( \290_b1 , \288_b1 , w_619 );
not ( w_619 , w_620 );
and ( \290_b0 , \288_b0 , w_621 );
and ( w_620 ,  , w_621 );
buf ( w_619 , \289_b1 );
not ( w_619 , w_622 );
not (  , w_623 );
and ( w_622 , w_623 , \289_b0 );
or ( \291_b1 , \290_b1 , \158_b1 );
not ( \158_b1 , w_624 );
and ( \291_b0 , \290_b0 , w_625 );
and ( w_624 , w_625 , \158_b0 );
buf ( \292_b1 , \290_b1 );
not ( \292_b1 , w_626 );
not ( \292_b0 , w_627 );
and ( w_626 , w_627 , \290_b0 );
or ( \293_b1 , \292_b1 , \223_b1 );
not ( \223_b1 , w_628 );
and ( \293_b0 , \292_b0 , w_629 );
and ( w_628 , w_629 , \223_b0 );
or ( \294_b1 , \291_b1 , w_631 );
not ( w_631 , w_632 );
and ( \294_b0 , \291_b0 , w_633 );
and ( w_632 ,  , w_633 );
buf ( w_631 , \293_b1 );
not ( w_631 , w_634 );
not (  , w_635 );
and ( w_634 , w_635 , \293_b0 );
buf ( \295_b1 , \294_b1 );
not ( \295_b1 , w_636 );
not ( \295_b0 , w_637 );
and ( w_636 , w_637 , \294_b0 );
buf ( \296_b1 , \132_b1 );
not ( \296_b1 , w_638 );
not ( \296_b0 , w_639 );
and ( w_638 , w_639 , \132_b0 );
buf ( \297_b1 , \296_b1 );
not ( \297_b1 , w_640 );
not ( \297_b0 , w_641 );
and ( w_640 , w_641 , \296_b0 );
or ( \298_b1 , \a[6]_b1 , \b[1]_b1 );
xor ( \298_b0 , \a[6]_b0 , w_642 );
not ( w_642 , w_643 );
and ( w_643 , \b[1]_b1 , \b[1]_b0 );
buf ( \299_b1 , \298_b1 );
not ( \299_b1 , w_644 );
not ( \299_b0 , w_645 );
and ( w_644 , w_645 , \298_b0 );
or ( \300_b1 , \297_b1 , w_646 );
or ( \300_b0 , \297_b0 , \299_b0 );
not ( \299_b0 , w_647 );
and ( w_647 , w_646 , \299_b1 );
or ( \301_b1 , \129_b1 , w_649 );
not ( w_649 , w_650 );
and ( \301_b0 , \129_b0 , w_651 );
and ( w_650 ,  , w_651 );
buf ( w_649 , \b[0]_b1 );
not ( w_649 , w_652 );
not (  , w_653 );
and ( w_652 , w_653 , \b[0]_b0 );
or ( \302_b1 , \300_b1 , w_655 );
not ( w_655 , w_656 );
and ( \302_b0 , \300_b0 , w_657 );
and ( w_656 ,  , w_657 );
buf ( w_655 , \301_b1 );
not ( w_655 , w_658 );
not (  , w_659 );
and ( w_658 , w_659 , \301_b0 );
or ( \303_b1 , \a[0]_b1 , \b[7]_b1 );
xor ( \303_b0 , \a[0]_b0 , w_660 );
not ( w_660 , w_661 );
and ( w_661 , \b[7]_b1 , \b[7]_b0 );
or ( \304_b1 , \303_b1 , w_663 );
not ( w_663 , w_664 );
and ( \304_b0 , \303_b0 , w_665 );
and ( w_664 ,  , w_665 );
buf ( w_663 , \175_b1 );
not ( w_663 , w_666 );
not (  , w_667 );
and ( w_666 , w_667 , \175_b0 );
or ( \305_b1 , \304_b1 , w_668 );
or ( \305_b0 , \304_b0 , \177_b0 );
not ( \177_b0 , w_669 );
and ( w_669 , w_668 , \177_b1 );
or ( \306_b1 , \189_b1 , w_671 );
not ( w_671 , w_672 );
and ( \306_b0 , \189_b0 , w_673 );
and ( w_672 ,  , w_673 );
buf ( w_671 , \177_b1 );
not ( w_671 , w_674 );
not (  , w_675 );
and ( w_674 , w_675 , \177_b0 );
or ( \307_b1 , \305_b1 , w_677 );
not ( w_677 , w_678 );
and ( \307_b0 , \305_b0 , w_679 );
and ( w_678 ,  , w_679 );
buf ( w_677 , \306_b1 );
not ( w_677 , w_680 );
not (  , w_681 );
and ( w_680 , w_681 , \306_b0 );
or ( \308_b1 , \302_b1 , \307_b1 );
xor ( \308_b0 , \302_b0 , w_682 );
not ( w_682 , w_683 );
and ( w_683 , \307_b1 , \307_b0 );
or ( \309_b1 , \a[2]_b1 , \b[5]_b1 );
xor ( \309_b0 , \a[2]_b0 , w_684 );
not ( w_684 , w_685 );
and ( w_685 , \b[5]_b1 , \b[5]_b0 );
buf ( \310_b1 , \309_b1 );
not ( \310_b1 , w_686 );
not ( \310_b0 , w_687 );
and ( w_686 , w_687 , \309_b0 );
buf ( \311_b1 , \267_b1 );
not ( \311_b1 , w_688 );
not ( \311_b0 , w_689 );
and ( w_688 , w_689 , \267_b0 );
or ( \312_b1 , \310_b1 , w_690 );
or ( \312_b0 , \310_b0 , \311_b0 );
not ( \311_b0 , w_691 );
and ( w_691 , w_690 , \311_b1 );
or ( \313_b1 , \121_b1 , w_693 );
not ( w_693 , w_694 );
and ( \313_b0 , \121_b0 , w_695 );
and ( w_694 ,  , w_695 );
buf ( w_693 , \195_b1 );
not ( w_693 , w_696 );
not (  , w_697 );
and ( w_696 , w_697 , \195_b0 );
or ( \314_b1 , \312_b1 , w_699 );
not ( w_699 , w_700 );
and ( \314_b0 , \312_b0 , w_701 );
and ( w_700 ,  , w_701 );
buf ( w_699 , \313_b1 );
not ( w_699 , w_702 );
not (  , w_703 );
and ( w_702 , w_703 , \313_b0 );
or ( \315_b1 , \308_b1 , \314_b1 );
not ( \314_b1 , w_704 );
and ( \315_b0 , \308_b0 , w_705 );
and ( w_704 , w_705 , \314_b0 );
or ( \316_b1 , \302_b1 , \307_b1 );
not ( \307_b1 , w_706 );
and ( \316_b0 , \302_b0 , w_707 );
and ( w_706 , w_707 , \307_b0 );
or ( \317_b1 , \315_b1 , w_708 );
or ( \317_b0 , \315_b0 , \316_b0 );
not ( \316_b0 , w_709 );
and ( w_709 , w_708 , \316_b1 );
or ( \318_b1 , \194_b1 , \202_b1 );
xor ( \318_b0 , \194_b0 , w_710 );
not ( w_710 , w_711 );
and ( w_711 , \202_b1 , \202_b0 );
or ( \319_b1 , \318_b1 , \216_b1 );
xor ( \319_b0 , \318_b0 , w_712 );
not ( w_712 , w_713 );
and ( w_713 , \216_b1 , \216_b0 );
or ( \320_b1 , \317_b1 , \319_b1 );
xor ( \320_b0 , \317_b0 , w_714 );
not ( w_714 , w_715 );
and ( w_715 , \319_b1 , \319_b0 );
or ( \321_b1 , \127_b1 , \138_b1 );
xor ( \321_b0 , \127_b0 , w_716 );
not ( w_716 , w_717 );
and ( w_717 , \138_b1 , \138_b0 );
or ( \322_b1 , \321_b1 , w_718 );
xor ( \322_b0 , \321_b0 , w_720 );
not ( w_720 , w_721 );
and ( w_721 , w_718 , w_719 );
buf ( w_718 , \153_b1 );
not ( w_718 , w_722 );
not ( w_719 , w_723 );
and ( w_722 , w_723 , \153_b0 );
buf ( \323_b1 , \322_b1 );
buf ( \323_b0 , \322_b0 );
or ( \324_b1 , \320_b1 , \323_b1 );
not ( \323_b1 , w_724 );
and ( \324_b0 , \320_b0 , w_725 );
and ( w_724 , w_725 , \323_b0 );
or ( \325_b1 , \317_b1 , \319_b1 );
not ( \319_b1 , w_726 );
and ( \325_b0 , \317_b0 , w_727 );
and ( w_726 , w_727 , \319_b0 );
or ( \326_b1 , \324_b1 , w_728 );
or ( \326_b0 , \324_b0 , \325_b0 );
not ( \325_b0 , w_729 );
and ( w_729 , w_728 , \325_b1 );
buf ( \327_b1 , \326_b1 );
not ( \327_b1 , w_730 );
not ( \327_b0 , w_731 );
and ( w_730 , w_731 , \326_b0 );
or ( \328_b1 , \295_b1 , w_733 );
not ( w_733 , w_734 );
and ( \328_b0 , \295_b0 , w_735 );
and ( w_734 ,  , w_735 );
buf ( w_733 , \327_b1 );
not ( w_733 , w_736 );
not (  , w_737 );
and ( w_736 , w_737 , \327_b0 );
or ( \329_b1 , \a[5]_b1 , \b[1]_b1 );
xor ( \329_b0 , \a[5]_b0 , w_738 );
not ( w_738 , w_739 );
and ( w_739 , \b[1]_b1 , \b[1]_b0 );
buf ( \330_b1 , \329_b1 );
not ( \330_b1 , w_740 );
not ( \330_b0 , w_741 );
and ( w_740 , w_741 , \329_b0 );
buf ( \331_b1 , \133_b1 );
not ( \331_b1 , w_742 );
not ( \331_b0 , w_743 );
and ( w_742 , w_743 , \133_b0 );
or ( \332_b1 , \330_b1 , w_744 );
or ( \332_b0 , \330_b0 , \331_b0 );
not ( \331_b0 , w_745 );
and ( w_745 , w_744 , \331_b1 );
or ( \333_b1 , \298_b1 , w_747 );
not ( w_747 , w_748 );
and ( \333_b0 , \298_b0 , w_749 );
and ( w_748 ,  , w_749 );
buf ( w_747 , \b[0]_b1 );
not ( w_747 , w_750 );
not (  , w_751 );
and ( w_750 , w_751 , \b[0]_b0 );
or ( \334_b1 , \332_b1 , w_753 );
not ( w_753 , w_754 );
and ( \334_b0 , \332_b0 , w_755 );
and ( w_754 ,  , w_755 );
buf ( w_753 , \333_b1 );
not ( w_753 , w_756 );
not (  , w_757 );
and ( w_756 , w_757 , \333_b0 );
buf ( \335_b1 , \334_b1 );
not ( \335_b1 , w_758 );
not ( \335_b0 , w_759 );
and ( w_758 , w_759 , \334_b0 );
buf ( \336_b1 , \335_b1 );
not ( \336_b1 , w_760 );
not ( \336_b0 , w_761 );
and ( w_760 , w_761 , \335_b0 );
or ( \337_b1 , \a[0]_b1 , w_762 );
or ( \337_b0 , \a[0]_b0 , \b[4]_b0 );
not ( \b[4]_b0 , w_763 );
and ( w_763 , w_762 , \b[4]_b1 );
or ( \338_b1 , \337_b1 , w_765 );
not ( w_765 , w_766 );
and ( \338_b0 , \337_b0 , w_767 );
and ( w_766 ,  , w_767 );
buf ( w_765 , \b[3]_b1 );
not ( w_765 , w_768 );
not (  , w_769 );
and ( w_768 , w_769 , \b[3]_b0 );
or ( \339_b1 , \a[0]_b1 , w_771 );
not ( w_771 , w_772 );
and ( \339_b0 , \a[0]_b0 , w_773 );
and ( w_772 ,  , w_773 );
buf ( w_771 , \b[4]_b1 );
not ( w_771 , w_774 );
not (  , w_775 );
and ( w_774 , w_775 , \b[4]_b0 );
buf ( \341_b1 , \340_b1 );
not ( \341_b1 , w_776 );
not ( \341_b0 , w_777 );
and ( w_776 , w_777 , \340_b0 );
or ( \342_b1 , \a[2]_b1 , \b[3]_b1 );
xor ( \342_b0 , \a[2]_b0 , w_778 );
not ( w_778 , w_779 );
and ( w_779 , \b[3]_b1 , \b[3]_b0 );
or ( \343_b1 , \b[3]_b1 , \b[2]_b1 );
xor ( \343_b0 , \b[3]_b0 , w_780 );
not ( w_780 , w_781 );
and ( w_781 , \b[2]_b1 , \b[2]_b0 );
or ( \344_b1 , \342_b1 , w_783 );
not ( w_783 , w_784 );
and ( \344_b0 , \342_b0 , w_785 );
and ( w_784 ,  , w_785 );
buf ( w_783 , \343_b1 );
not ( w_783 , w_786 );
not (  , w_787 );
and ( w_786 , w_787 , \343_b0 );
or ( \345_b1 , \344_b1 , w_788 );
or ( \345_b0 , \344_b0 , \150_b0 );
not ( \150_b0 , w_789 );
and ( w_789 , w_788 , \150_b1 );
or ( \346_b1 , \b[3]_b1 , \a[3]_b1 );
xor ( \346_b0 , \b[3]_b0 , w_790 );
not ( w_790 , w_791 );
and ( w_791 , \a[3]_b1 , \a[3]_b0 );
or ( \347_b1 , \346_b1 , w_793 );
not ( w_793 , w_794 );
and ( \347_b0 , \346_b0 , w_795 );
and ( w_794 ,  , w_795 );
buf ( w_793 , \150_b1 );
not ( w_793 , w_796 );
not (  , w_797 );
and ( w_796 , w_797 , \150_b0 );
or ( \348_b1 , \345_b1 , w_799 );
not ( w_799 , w_800 );
and ( \348_b0 , \345_b0 , w_801 );
and ( w_800 ,  , w_801 );
buf ( w_799 , \347_b1 );
not ( w_799 , w_802 );
not (  , w_803 );
and ( w_802 , w_803 , \347_b0 );
or ( \349_b1 , \341_b1 , w_805 );
not ( w_805 , w_806 );
and ( \349_b0 , \341_b0 , w_807 );
and ( w_806 ,  , w_807 );
buf ( w_805 , \348_b1 );
not ( w_805 , w_808 );
not (  , w_809 );
and ( w_808 , w_809 , \348_b0 );
buf ( \350_b1 , \349_b1 );
not ( \350_b1 , w_810 );
not ( \350_b0 , w_811 );
and ( w_810 , w_811 , \349_b0 );
buf ( \351_b1 , \350_b1 );
not ( \351_b1 , w_812 );
not ( \351_b0 , w_813 );
and ( w_812 , w_813 , \350_b0 );
or ( \352_b1 , \336_b1 , w_814 );
or ( \352_b0 , \336_b0 , \351_b0 );
not ( \351_b0 , w_815 );
and ( w_815 , w_814 , \351_b1 );
or ( \353_b1 , \350_b1 , w_816 );
or ( \353_b0 , \350_b0 , \335_b0 );
not ( \335_b0 , w_817 );
and ( w_817 , w_816 , \335_b1 );
or ( \354_b1 , \352_b1 , w_819 );
not ( w_819 , w_820 );
and ( \354_b0 , \352_b0 , w_821 );
and ( w_820 ,  , w_821 );
buf ( w_819 , \353_b1 );
not ( w_819 , w_822 );
not (  , w_823 );
and ( w_822 , w_823 , \353_b0 );
buf ( \355_b1 , \354_b1 );
not ( \355_b1 , w_824 );
not ( \355_b0 , w_825 );
and ( w_824 , w_825 , \354_b0 );
buf ( \356_b1 , \355_b1 );
not ( \356_b1 , w_826 );
not ( \356_b0 , w_827 );
and ( w_826 , w_827 , \355_b0 );
or ( \357_b1 , \177_b1 , w_829 );
not ( w_829 , w_830 );
and ( \357_b0 , \177_b0 , w_831 );
and ( w_830 ,  , w_831 );
buf ( w_829 , \a[0]_b1 );
not ( w_829 , w_832 );
not (  , w_833 );
and ( w_832 , w_833 , \a[0]_b0 );
buf ( \358_b1 , \357_b1 );
not ( \358_b1 , w_834 );
not ( \358_b0 , w_835 );
and ( w_834 , w_835 , \357_b0 );
or ( \359_b1 , \a[1]_b1 , \b[5]_b1 );
xor ( \359_b0 , \a[1]_b0 , w_836 );
not ( w_836 , w_837 );
and ( w_837 , \b[5]_b1 , \b[5]_b0 );
or ( \360_b1 , \359_b1 , w_839 );
not ( w_839 , w_840 );
and ( \360_b0 , \359_b0 , w_841 );
and ( w_840 ,  , w_841 );
buf ( w_839 , \117_b1 );
not ( w_839 , w_842 );
not (  , w_843 );
and ( w_842 , w_843 , \117_b0 );
or ( \361_b1 , \360_b1 , w_844 );
or ( \361_b0 , \360_b0 , \119_b0 );
not ( \119_b0 , w_845 );
and ( w_845 , w_844 , \119_b1 );
or ( \362_b1 , \309_b1 , w_847 );
not ( w_847 , w_848 );
and ( \362_b0 , \309_b0 , w_849 );
and ( w_848 ,  , w_849 );
buf ( w_847 , \119_b1 );
not ( w_847 , w_850 );
not (  , w_851 );
and ( w_850 , w_851 , \119_b0 );
or ( \363_b1 , \361_b1 , w_853 );
not ( w_853 , w_854 );
and ( \363_b0 , \361_b0 , w_855 );
and ( w_854 ,  , w_855 );
buf ( w_853 , \362_b1 );
not ( w_853 , w_856 );
not (  , w_857 );
and ( w_856 , w_857 , \362_b0 );
or ( \364_b1 , \358_b1 , \363_b1 );
xor ( \364_b0 , \358_b0 , w_858 );
not ( w_858 , w_859 );
and ( w_859 , \363_b1 , \363_b0 );
buf ( \365_b1 , \346_b1 );
not ( \365_b1 , w_860 );
not ( \365_b0 , w_861 );
and ( w_860 , w_861 , \346_b0 );
buf ( \366_b1 , \147_b1 );
not ( \366_b1 , w_862 );
not ( \366_b0 , w_863 );
and ( w_862 , w_863 , \147_b0 );
or ( \367_b1 , \365_b1 , w_864 );
or ( \367_b0 , \365_b0 , \366_b0 );
not ( \366_b0 , w_865 );
and ( w_865 , w_864 , \366_b1 );
buf ( \368_b1 , \212_b1 );
not ( \368_b1 , w_866 );
not ( \368_b0 , w_867 );
and ( w_866 , w_867 , \212_b0 );
or ( \369_b1 , \368_b1 , w_869 );
not ( w_869 , w_870 );
and ( \369_b0 , \368_b0 , w_871 );
and ( w_870 ,  , w_871 );
buf ( w_869 , \150_b1 );
not ( w_869 , w_872 );
not (  , w_873 );
and ( w_872 , w_873 , \150_b0 );
or ( \370_b1 , \367_b1 , w_875 );
not ( w_875 , w_876 );
and ( \370_b0 , \367_b0 , w_877 );
and ( w_876 ,  , w_877 );
buf ( w_875 , \369_b1 );
not ( w_875 , w_878 );
not (  , w_879 );
and ( w_878 , w_879 , \369_b0 );
or ( \371_b1 , \364_b1 , w_880 );
xor ( \371_b0 , \364_b0 , w_882 );
not ( w_882 , w_883 );
and ( w_883 , w_880 , w_881 );
buf ( w_880 , \370_b1 );
not ( w_880 , w_884 );
not ( w_881 , w_885 );
and ( w_884 , w_885 , \370_b0 );
buf ( \372_b1 , \371_b1 );
not ( \372_b1 , w_886 );
not ( \372_b0 , w_887 );
and ( w_886 , w_887 , \371_b0 );
buf ( \373_b1 , \372_b1 );
not ( \373_b1 , w_888 );
not ( \373_b0 , w_889 );
and ( w_888 , w_889 , \372_b0 );
or ( \374_b1 , \356_b1 , w_890 );
or ( \374_b0 , \356_b0 , \373_b0 );
not ( \373_b0 , w_891 );
and ( w_891 , w_890 , \373_b1 );
or ( \375_b1 , \354_b1 , w_893 );
not ( w_893 , w_894 );
and ( \375_b0 , \354_b0 , w_895 );
and ( w_894 ,  , w_895 );
buf ( w_893 , \371_b1 );
not ( w_893 , w_896 );
not (  , w_897 );
and ( w_896 , w_897 , \371_b0 );
or ( \376_b1 , \374_b1 , w_899 );
not ( w_899 , w_900 );
and ( \376_b0 , \374_b0 , w_901 );
and ( w_900 ,  , w_901 );
buf ( w_899 , \375_b1 );
not ( w_899 , w_902 );
not (  , w_903 );
and ( w_902 , w_903 , \375_b0 );
buf ( \377_b1 , \376_b1 );
not ( \377_b1 , w_904 );
not ( \377_b0 , w_905 );
and ( w_904 , w_905 , \376_b0 );
buf ( \378_b1 , \348_b1 );
not ( \378_b1 , w_906 );
not ( \378_b0 , w_907 );
and ( w_906 , w_907 , \348_b0 );
buf ( \379_b1 , \340_b1 );
not ( \379_b1 , w_908 );
not ( \379_b0 , w_909 );
and ( w_908 , w_909 , \340_b0 );
or ( \380_b1 , \378_b1 , \379_b1 );
not ( \379_b1 , w_910 );
and ( \380_b0 , \378_b0 , w_911 );
and ( w_910 , w_911 , \379_b0 );
or ( \381_b1 , \348_b1 , \340_b1 );
not ( \340_b1 , w_912 );
and ( \381_b0 , \348_b0 , w_913 );
and ( w_912 , w_913 , \340_b0 );
or ( \382_b1 , \380_b1 , w_915 );
not ( w_915 , w_916 );
and ( \382_b0 , \380_b0 , w_917 );
and ( w_916 ,  , w_917 );
buf ( w_915 , \381_b1 );
not ( w_915 , w_918 );
not (  , w_919 );
and ( w_918 , w_919 , \381_b0 );
buf ( \383_b1 , \382_b1 );
not ( \383_b1 , w_920 );
not ( \383_b0 , w_921 );
and ( w_920 , w_921 , \382_b0 );
or ( \384_b1 , \b[1]_b1 , \a[4]_b1 );
xor ( \384_b0 , \b[1]_b0 , w_922 );
not ( w_922 , w_923 );
and ( w_923 , \a[4]_b1 , \a[4]_b0 );
buf ( \385_b1 , \384_b1 );
not ( \385_b1 , w_924 );
not ( \385_b0 , w_925 );
and ( w_924 , w_925 , \384_b0 );
buf ( \386_b1 , \133_b1 );
not ( \386_b1 , w_926 );
not ( \386_b0 , w_927 );
and ( w_926 , w_927 , \133_b0 );
or ( \387_b1 , \385_b1 , w_928 );
or ( \387_b0 , \385_b0 , \386_b0 );
not ( \386_b0 , w_929 );
and ( w_929 , w_928 , \386_b1 );
or ( \388_b1 , \329_b1 , w_931 );
not ( w_931 , w_932 );
and ( \388_b0 , \329_b0 , w_933 );
and ( w_932 ,  , w_933 );
buf ( w_931 , \b[0]_b1 );
not ( w_931 , w_934 );
not (  , w_935 );
and ( w_934 , w_935 , \b[0]_b0 );
or ( \389_b1 , \387_b1 , w_937 );
not ( w_937 , w_938 );
and ( \389_b0 , \387_b0 , w_939 );
and ( w_938 ,  , w_939 );
buf ( w_937 , \388_b1 );
not ( w_937 , w_940 );
not (  , w_941 );
and ( w_940 , w_941 , \388_b0 );
or ( \390_b1 , \383_b1 , w_942 );
or ( \390_b0 , \383_b0 , \389_b0 );
not ( \389_b0 , w_943 );
and ( w_943 , w_942 , \389_b1 );
or ( \391_b1 , \a[0]_b1 , \b[5]_b1 );
xor ( \391_b0 , \a[0]_b0 , w_944 );
not ( w_944 , w_945 );
and ( w_945 , \b[5]_b1 , \b[5]_b0 );
buf ( \392_b1 , \391_b1 );
not ( \392_b1 , w_946 );
not ( \392_b0 , w_947 );
and ( w_946 , w_947 , \391_b0 );
buf ( \393_b1 , \198_b1 );
not ( \393_b1 , w_948 );
not ( \393_b0 , w_949 );
and ( w_948 , w_949 , \198_b0 );
or ( \394_b1 , \392_b1 , w_950 );
or ( \394_b0 , \392_b0 , \393_b0 );
not ( \393_b0 , w_951 );
and ( w_951 , w_950 , \393_b1 );
or ( \395_b1 , \121_b1 , w_953 );
not ( w_953 , w_954 );
and ( \395_b0 , \121_b0 , w_955 );
and ( w_954 ,  , w_955 );
buf ( w_953 , \359_b1 );
not ( w_953 , w_956 );
not (  , w_957 );
and ( w_956 , w_957 , \359_b0 );
or ( \396_b1 , \394_b1 , w_959 );
not ( w_959 , w_960 );
and ( \396_b0 , \394_b0 , w_961 );
and ( w_960 ,  , w_961 );
buf ( w_959 , \395_b1 );
not ( w_959 , w_962 );
not (  , w_963 );
and ( w_962 , w_963 , \395_b0 );
or ( \397_b1 , \390_b1 , w_965 );
not ( w_965 , w_966 );
and ( \397_b0 , \390_b0 , w_967 );
and ( w_966 ,  , w_967 );
buf ( w_965 , \396_b1 );
not ( w_965 , w_968 );
not (  , w_969 );
and ( w_968 , w_969 , \396_b0 );
buf ( \398_b1 , \389_b1 );
not ( \398_b1 , w_970 );
not ( \398_b0 , w_971 );
and ( w_970 , w_971 , \389_b0 );
buf ( \399_b1 , \398_b1 );
not ( \399_b1 , w_972 );
not ( \399_b0 , w_973 );
and ( w_972 , w_973 , \398_b0 );
or ( \400_b1 , \399_b1 , w_975 );
not ( w_975 , w_976 );
and ( \400_b0 , \399_b0 , w_977 );
and ( w_976 ,  , w_977 );
buf ( w_975 , \383_b1 );
not ( w_975 , w_978 );
not (  , w_979 );
and ( w_978 , w_979 , \383_b0 );
or ( \401_b1 , \397_b1 , w_981 );
not ( w_981 , w_982 );
and ( \401_b0 , \397_b0 , w_983 );
and ( w_982 ,  , w_983 );
buf ( w_981 , \400_b1 );
not ( w_981 , w_984 );
not (  , w_985 );
and ( w_984 , w_985 , \400_b0 );
buf ( \402_b1 , \401_b1 );
not ( \402_b1 , w_986 );
not ( \402_b0 , w_987 );
and ( w_986 , w_987 , \401_b0 );
or ( \403_b1 , \377_b1 , w_989 );
not ( w_989 , w_990 );
and ( \403_b0 , \377_b0 , w_991 );
and ( w_990 ,  , w_991 );
buf ( w_989 , \402_b1 );
not ( w_989 , w_992 );
not (  , w_993 );
and ( w_992 , w_993 , \402_b0 );
buf ( \404_b1 , \403_b1 );
not ( \404_b1 , w_994 );
not ( \404_b0 , w_995 );
and ( w_994 , w_995 , \403_b0 );
or ( \405_b1 , \207_b1 , \215_b1 );
xor ( \405_b0 , \207_b0 , w_996 );
not ( w_996 , w_997 );
and ( w_997 , \215_b1 , \215_b0 );
or ( \406_b1 , \302_b1 , \307_b1 );
xor ( \406_b0 , \302_b0 , w_998 );
not ( w_998 , w_999 );
and ( w_999 , \307_b1 , \307_b0 );
or ( \407_b1 , \406_b1 , \314_b1 );
xor ( \407_b0 , \406_b0 , w_1000 );
not ( w_1000 , w_1001 );
and ( w_1001 , \314_b1 , \314_b0 );
or ( \408_b1 , \405_b1 , \407_b1 );
xor ( \408_b0 , \405_b0 , w_1002 );
not ( w_1002 , w_1003 );
and ( w_1003 , \407_b1 , \407_b0 );
buf ( \409_b1 , \363_b1 );
not ( \409_b1 , w_1004 );
not ( \409_b0 , w_1005 );
and ( w_1004 , w_1005 , \363_b0 );
or ( \410_b1 , \409_b1 , w_1007 );
not ( w_1007 , w_1008 );
and ( \410_b0 , \409_b0 , w_1009 );
and ( w_1008 ,  , w_1009 );
buf ( w_1007 , \357_b1 );
not ( w_1007 , w_1010 );
not (  , w_1011 );
and ( w_1010 , w_1011 , \357_b0 );
buf ( \411_b1 , \410_b1 );
not ( \411_b1 , w_1012 );
not ( \411_b0 , w_1013 );
and ( w_1012 , w_1013 , \410_b0 );
buf ( \412_b1 , \370_b1 );
not ( \412_b1 , w_1014 );
not ( \412_b0 , w_1015 );
and ( w_1014 , w_1015 , \370_b0 );
or ( \413_b1 , \411_b1 , w_1016 );
or ( \413_b0 , \411_b0 , \412_b0 );
not ( \412_b0 , w_1017 );
and ( w_1017 , w_1016 , \412_b1 );
or ( \414_b1 , \363_b1 , w_1019 );
not ( w_1019 , w_1020 );
and ( \414_b0 , \363_b0 , w_1021 );
and ( w_1020 ,  , w_1021 );
buf ( w_1019 , \358_b1 );
not ( w_1019 , w_1022 );
not (  , w_1023 );
and ( w_1022 , w_1023 , \358_b0 );
or ( \415_b1 , \413_b1 , w_1025 );
not ( w_1025 , w_1026 );
and ( \415_b0 , \413_b0 , w_1027 );
and ( w_1026 ,  , w_1027 );
buf ( w_1025 , \414_b1 );
not ( w_1025 , w_1028 );
not (  , w_1029 );
and ( w_1028 , w_1029 , \414_b0 );
or ( \416_b1 , \408_b1 , \415_b1 );
xor ( \416_b0 , \408_b0 , w_1030 );
not ( w_1030 , w_1031 );
and ( w_1031 , \415_b1 , \415_b0 );
or ( \417_b1 , \349_b1 , w_1033 );
not ( w_1033 , w_1034 );
and ( \417_b0 , \349_b0 , w_1035 );
and ( w_1034 ,  , w_1035 );
buf ( w_1033 , \335_b1 );
not ( w_1033 , w_1036 );
not (  , w_1037 );
and ( w_1036 , w_1037 , \335_b0 );
buf ( \418_b1 , \417_b1 );
not ( \418_b1 , w_1038 );
not ( \418_b0 , w_1039 );
and ( w_1038 , w_1039 , \417_b0 );
buf ( \419_b1 , \372_b1 );
not ( \419_b1 , w_1040 );
not ( \419_b0 , w_1041 );
and ( w_1040 , w_1041 , \372_b0 );
or ( \420_b1 , \418_b1 , w_1042 );
or ( \420_b0 , \418_b0 , \419_b0 );
not ( \419_b0 , w_1043 );
and ( w_1043 , w_1042 , \419_b1 );
or ( \421_b1 , \350_b1 , w_1045 );
not ( w_1045 , w_1046 );
and ( \421_b0 , \350_b0 , w_1047 );
and ( w_1046 ,  , w_1047 );
buf ( w_1045 , \334_b1 );
not ( w_1045 , w_1048 );
not (  , w_1049 );
and ( w_1048 , w_1049 , \334_b0 );
or ( \422_b1 , \420_b1 , w_1051 );
not ( w_1051 , w_1052 );
and ( \422_b0 , \420_b0 , w_1053 );
and ( w_1052 ,  , w_1053 );
buf ( w_1051 , \421_b1 );
not ( w_1051 , w_1054 );
not (  , w_1055 );
and ( w_1054 , w_1055 , \421_b0 );
or ( \423_b1 , \416_b1 , w_1057 );
not ( w_1057 , w_1058 );
and ( \423_b0 , \416_b0 , w_1059 );
and ( w_1058 ,  , w_1059 );
buf ( w_1057 , \422_b1 );
not ( w_1057 , w_1060 );
not (  , w_1061 );
and ( w_1060 , w_1061 , \422_b0 );
or ( \424_b1 , \404_b1 , \423_b1 );
not ( \423_b1 , w_1062 );
and ( \424_b0 , \404_b0 , w_1063 );
and ( w_1062 , w_1063 , \423_b0 );
or ( \425_b1 , \416_b1 , w_1065 );
not ( w_1065 , w_1066 );
and ( \425_b0 , \416_b0 , w_1067 );
and ( w_1066 ,  , w_1067 );
buf ( w_1065 , \422_b1 );
not ( w_1065 , w_1068 );
not (  , w_1069 );
and ( w_1068 , w_1069 , \422_b0 );
or ( \426_b1 , \424_b1 , w_1071 );
not ( w_1071 , w_1072 );
and ( \426_b0 , \424_b0 , w_1073 );
and ( w_1072 ,  , w_1073 );
buf ( w_1071 , \425_b1 );
not ( w_1071 , w_1074 );
not (  , w_1075 );
and ( w_1074 , w_1075 , \425_b0 );
buf ( \427_b1 , \163_b1 );
not ( \427_b1 , w_1076 );
not ( \427_b0 , w_1077 );
and ( w_1076 , w_1077 , \163_b0 );
or ( \428_b1 , \b[1]_b1 , \a[3]_b1 );
xor ( \428_b0 , \b[1]_b0 , w_1078 );
not ( w_1078 , w_1079 );
and ( w_1079 , \a[3]_b1 , \a[3]_b0 );
buf ( \429_b1 , \428_b1 );
not ( \429_b1 , w_1080 );
not ( \429_b0 , w_1081 );
and ( w_1080 , w_1081 , \428_b0 );
or ( \430_b1 , \427_b1 , w_1082 );
or ( \430_b0 , \427_b0 , \429_b0 );
not ( \429_b0 , w_1083 );
and ( w_1083 , w_1082 , \429_b1 );
or ( \431_b1 , \384_b1 , w_1085 );
not ( w_1085 , w_1086 );
and ( \431_b0 , \384_b0 , w_1087 );
and ( w_1086 ,  , w_1087 );
buf ( w_1085 , \b[0]_b1 );
not ( w_1085 , w_1088 );
not (  , w_1089 );
and ( w_1088 , w_1089 , \b[0]_b0 );
or ( \432_b1 , \430_b1 , w_1091 );
not ( w_1091 , w_1092 );
and ( \432_b0 , \430_b0 , w_1093 );
and ( w_1092 ,  , w_1093 );
buf ( w_1091 , \431_b1 );
not ( w_1091 , w_1094 );
not (  , w_1095 );
and ( w_1094 , w_1095 , \431_b0 );
buf ( \433_b1 , \432_b1 );
not ( \433_b1 , w_1096 );
not ( \433_b0 , w_1097 );
and ( w_1096 , w_1097 , \432_b0 );
or ( \434_b1 , \121_b1 , w_1099 );
not ( w_1099 , w_1100 );
and ( \434_b0 , \121_b0 , w_1101 );
and ( w_1100 ,  , w_1101 );
buf ( w_1099 , \a[0]_b1 );
not ( w_1099 , w_1102 );
not (  , w_1103 );
and ( w_1102 , w_1103 , \a[0]_b0 );
or ( \435_b1 , \433_b1 , w_1105 );
not ( w_1105 , w_1106 );
and ( \435_b0 , \433_b0 , w_1107 );
and ( w_1106 ,  , w_1107 );
buf ( w_1105 , \434_b1 );
not ( w_1105 , w_1108 );
not (  , w_1109 );
and ( w_1108 , w_1109 , \434_b0 );
buf ( \436_b1 , \435_b1 );
not ( \436_b1 , w_1110 );
not ( \436_b0 , w_1111 );
and ( w_1110 , w_1111 , \435_b0 );
or ( \437_b1 , \a[1]_b1 , \b[3]_b1 );
xor ( \437_b0 , \a[1]_b0 , w_1112 );
not ( w_1112 , w_1113 );
and ( w_1113 , \b[3]_b1 , \b[3]_b0 );
buf ( \438_b1 , \437_b1 );
not ( \438_b1 , w_1114 );
not ( \438_b0 , w_1115 );
and ( w_1114 , w_1115 , \437_b0 );
buf ( \439_b1 , \242_b1 );
not ( \439_b1 , w_1116 );
not ( \439_b0 , w_1117 );
and ( w_1116 , w_1117 , \242_b0 );
or ( \440_b1 , \438_b1 , w_1118 );
or ( \440_b0 , \438_b0 , \439_b0 );
not ( \439_b0 , w_1119 );
and ( w_1119 , w_1118 , \439_b1 );
or ( \441_b1 , \150_b1 , w_1121 );
not ( w_1121 , w_1122 );
and ( \441_b0 , \150_b0 , w_1123 );
and ( w_1122 ,  , w_1123 );
buf ( w_1121 , \342_b1 );
not ( w_1121 , w_1124 );
not (  , w_1125 );
and ( w_1124 , w_1125 , \342_b0 );
or ( \442_b1 , \440_b1 , w_1127 );
not ( w_1127 , w_1128 );
and ( \442_b0 , \440_b0 , w_1129 );
and ( w_1128 ,  , w_1129 );
buf ( w_1127 , \441_b1 );
not ( w_1127 , w_1130 );
not (  , w_1131 );
and ( w_1130 , w_1131 , \441_b0 );
buf ( \443_b1 , \442_b1 );
not ( \443_b1 , w_1132 );
not ( \443_b0 , w_1133 );
and ( w_1132 , w_1133 , \442_b0 );
or ( \444_b1 , \436_b1 , w_1134 );
or ( \444_b0 , \436_b0 , \443_b0 );
not ( \443_b0 , w_1135 );
and ( w_1135 , w_1134 , \443_b1 );
buf ( \445_b1 , \434_b1 );
not ( \445_b1 , w_1136 );
not ( \445_b0 , w_1137 );
and ( w_1136 , w_1137 , \434_b0 );
or ( \446_b1 , \445_b1 , w_1139 );
not ( w_1139 , w_1140 );
and ( \446_b0 , \445_b0 , w_1141 );
and ( w_1140 ,  , w_1141 );
buf ( w_1139 , \432_b1 );
not ( w_1139 , w_1142 );
not (  , w_1143 );
and ( w_1142 , w_1143 , \432_b0 );
or ( \447_b1 , \444_b1 , w_1145 );
not ( w_1145 , w_1146 );
and ( \447_b0 , \444_b0 , w_1147 );
and ( w_1146 ,  , w_1147 );
buf ( w_1145 , \446_b1 );
not ( w_1145 , w_1148 );
not (  , w_1149 );
and ( w_1148 , w_1149 , \446_b0 );
buf ( \448_b1 , \447_b1 );
not ( \448_b1 , w_1150 );
not ( \448_b0 , w_1151 );
and ( w_1150 , w_1151 , \447_b0 );
buf ( \449_b1 , \398_b1 );
not ( \449_b1 , w_1152 );
not ( \449_b0 , w_1153 );
and ( w_1152 , w_1153 , \398_b0 );
buf ( \450_b1 , \396_b1 );
not ( \450_b1 , w_1154 );
not ( \450_b0 , w_1155 );
and ( w_1154 , w_1155 , \396_b0 );
or ( \451_b1 , \449_b1 , w_1156 );
or ( \451_b0 , \449_b0 , \450_b0 );
not ( \450_b0 , w_1157 );
and ( w_1157 , w_1156 , \450_b1 );
or ( \452_b1 , \396_b1 , w_1158 );
or ( \452_b0 , \396_b0 , \398_b0 );
not ( \398_b0 , w_1159 );
and ( w_1159 , w_1158 , \398_b1 );
or ( \453_b1 , \451_b1 , w_1161 );
not ( w_1161 , w_1162 );
and ( \453_b0 , \451_b0 , w_1163 );
and ( w_1162 ,  , w_1163 );
buf ( w_1161 , \452_b1 );
not ( w_1161 , w_1164 );
not (  , w_1165 );
and ( w_1164 , w_1165 , \452_b0 );
or ( \454_b1 , \453_b1 , \382_b1 );
not ( \382_b1 , w_1166 );
and ( \454_b0 , \453_b0 , w_1167 );
and ( w_1166 , w_1167 , \382_b0 );
buf ( \455_b1 , \453_b1 );
not ( \455_b1 , w_1168 );
not ( \455_b0 , w_1169 );
and ( w_1168 , w_1169 , \453_b0 );
or ( \456_b1 , \455_b1 , \383_b1 );
not ( \383_b1 , w_1170 );
and ( \456_b0 , \455_b0 , w_1171 );
and ( w_1170 , w_1171 , \383_b0 );
or ( \457_b1 , \454_b1 , w_1173 );
not ( w_1173 , w_1174 );
and ( \457_b0 , \454_b0 , w_1175 );
and ( w_1174 ,  , w_1175 );
buf ( w_1173 , \456_b1 );
not ( w_1173 , w_1176 );
not (  , w_1177 );
and ( w_1176 , w_1177 , \456_b0 );
or ( \458_b1 , \448_b1 , w_1179 );
not ( w_1179 , w_1180 );
and ( \458_b0 , \448_b0 , w_1181 );
and ( w_1180 ,  , w_1181 );
buf ( w_1179 , \457_b1 );
not ( w_1179 , w_1182 );
not (  , w_1183 );
and ( w_1182 , w_1183 , \457_b0 );
buf ( \459_b1 , \458_b1 );
not ( \459_b1 , w_1184 );
not ( \459_b0 , w_1185 );
and ( w_1184 , w_1185 , \458_b0 );
or ( \460_b1 , \a[0]_b1 , w_1187 );
not ( w_1187 , w_1188 );
and ( \460_b0 , \a[0]_b0 , w_1189 );
and ( w_1188 ,  , w_1189 );
buf ( w_1187 , \b[2]_b1 );
not ( w_1187 , w_1190 );
not (  , w_1191 );
and ( w_1190 , w_1191 , \b[2]_b0 );
or ( \461_b1 , \460_b1 , \b[3]_b1 );
not ( \b[3]_b1 , w_1192 );
and ( \461_b0 , \460_b0 , w_1193 );
and ( w_1192 , w_1193 , \b[3]_b0 );
or ( \462_b1 , \a[0]_b1 , w_1194 );
or ( \462_b0 , \a[0]_b0 , \b[2]_b0 );
not ( \b[2]_b0 , w_1195 );
and ( w_1195 , w_1194 , \b[2]_b1 );
or ( \463_b1 , \462_b1 , w_1197 );
not ( w_1197 , w_1198 );
and ( \463_b0 , \462_b0 , w_1199 );
and ( w_1198 ,  , w_1199 );
buf ( w_1197 , \b[1]_b1 );
not ( w_1197 , w_1200 );
not (  , w_1201 );
and ( w_1200 , w_1201 , \b[1]_b0 );
or ( \464_b1 , \461_b1 , w_1203 );
not ( w_1203 , w_1204 );
and ( \464_b0 , \461_b0 , w_1205 );
and ( w_1204 ,  , w_1205 );
buf ( w_1203 , \463_b1 );
not ( w_1203 , w_1206 );
not (  , w_1207 );
and ( w_1206 , w_1207 , \463_b0 );
buf ( \465_b1 , \464_b1 );
not ( \465_b1 , w_1208 );
not ( \465_b0 , w_1209 );
and ( w_1208 , w_1209 , \464_b0 );
or ( \466_b1 , \a[2]_b1 , \b[1]_b1 );
xor ( \466_b0 , \a[2]_b0 , w_1210 );
not ( w_1210 , w_1211 );
and ( w_1211 , \b[1]_b1 , \b[1]_b0 );
buf ( \467_b1 , \466_b1 );
not ( \467_b1 , w_1212 );
not ( \467_b0 , w_1213 );
and ( w_1212 , w_1213 , \466_b0 );
buf ( \468_b1 , \163_b1 );
not ( \468_b1 , w_1214 );
not ( \468_b0 , w_1215 );
and ( w_1214 , w_1215 , \163_b0 );
or ( \469_b1 , \467_b1 , w_1216 );
or ( \469_b0 , \467_b0 , \468_b0 );
not ( \468_b0 , w_1217 );
and ( w_1217 , w_1216 , \468_b1 );
or ( \470_b1 , \428_b1 , w_1219 );
not ( w_1219 , w_1220 );
and ( \470_b0 , \428_b0 , w_1221 );
and ( w_1220 ,  , w_1221 );
buf ( w_1219 , \b[0]_b1 );
not ( w_1219 , w_1222 );
not (  , w_1223 );
and ( w_1222 , w_1223 , \b[0]_b0 );
or ( \471_b1 , \469_b1 , w_1225 );
not ( w_1225 , w_1226 );
and ( \471_b0 , \469_b0 , w_1227 );
and ( w_1226 ,  , w_1227 );
buf ( w_1225 , \470_b1 );
not ( w_1225 , w_1228 );
not (  , w_1229 );
and ( w_1228 , w_1229 , \470_b0 );
or ( \472_b1 , \465_b1 , w_1231 );
not ( w_1231 , w_1232 );
and ( \472_b0 , \465_b0 , w_1233 );
and ( w_1232 ,  , w_1233 );
buf ( w_1231 , \471_b1 );
not ( w_1231 , w_1234 );
not (  , w_1235 );
and ( w_1234 , w_1235 , \471_b0 );
buf ( \473_b1 , \472_b1 );
not ( \473_b1 , w_1236 );
not ( \473_b0 , w_1237 );
and ( w_1236 , w_1237 , \472_b0 );
buf ( \474_b1 , \432_b1 );
not ( \474_b1 , w_1238 );
not ( \474_b0 , w_1239 );
and ( w_1238 , w_1239 , \432_b0 );
buf ( \475_b1 , \434_b1 );
not ( \475_b1 , w_1240 );
not ( \475_b0 , w_1241 );
and ( w_1240 , w_1241 , \434_b0 );
or ( \476_b1 , \474_b1 , \475_b1 );
not ( \475_b1 , w_1242 );
and ( \476_b0 , \474_b0 , w_1243 );
and ( w_1242 , w_1243 , \475_b0 );
or ( \477_b1 , \432_b1 , \434_b1 );
not ( \434_b1 , w_1244 );
and ( \477_b0 , \432_b0 , w_1245 );
and ( w_1244 , w_1245 , \434_b0 );
or ( \478_b1 , \476_b1 , w_1247 );
not ( w_1247 , w_1248 );
and ( \478_b0 , \476_b0 , w_1249 );
and ( w_1248 ,  , w_1249 );
buf ( w_1247 , \477_b1 );
not ( w_1247 , w_1250 );
not (  , w_1251 );
and ( w_1250 , w_1251 , \477_b0 );
buf ( \479_b1 , \478_b1 );
not ( \479_b1 , w_1252 );
not ( \479_b0 , w_1253 );
and ( w_1252 , w_1253 , \478_b0 );
buf ( \480_b1 , \442_b1 );
not ( \480_b1 , w_1254 );
not ( \480_b0 , w_1255 );
and ( w_1254 , w_1255 , \442_b0 );
or ( \481_b1 , \479_b1 , \480_b1 );
not ( \480_b1 , w_1256 );
and ( \481_b0 , \479_b0 , w_1257 );
and ( w_1256 , w_1257 , \480_b0 );
or ( \482_b1 , \442_b1 , \478_b1 );
not ( \478_b1 , w_1258 );
and ( \482_b0 , \442_b0 , w_1259 );
and ( w_1258 , w_1259 , \478_b0 );
or ( \483_b1 , \481_b1 , w_1261 );
not ( w_1261 , w_1262 );
and ( \483_b0 , \481_b0 , w_1263 );
and ( w_1262 ,  , w_1263 );
buf ( w_1261 , \482_b1 );
not ( w_1261 , w_1264 );
not (  , w_1265 );
and ( w_1264 , w_1265 , \482_b0 );
buf ( \484_b1 , \483_b1 );
not ( \484_b1 , w_1266 );
not ( \484_b0 , w_1267 );
and ( w_1266 , w_1267 , \483_b0 );
or ( \485_b1 , \473_b1 , w_1268 );
or ( \485_b0 , \473_b0 , \484_b0 );
not ( \484_b0 , w_1269 );
and ( w_1269 , w_1268 , \484_b1 );
or ( \486_b1 , \b[3]_b1 , \a[0]_b1 );
xor ( \486_b0 , \b[3]_b0 , w_1270 );
not ( w_1270 , w_1271 );
and ( w_1271 , \a[0]_b1 , \a[0]_b0 );
buf ( \487_b1 , \486_b1 );
not ( \487_b1 , w_1272 );
not ( \487_b0 , w_1273 );
and ( w_1272 , w_1273 , \486_b0 );
buf ( \488_b1 , \242_b1 );
not ( \488_b1 , w_1274 );
not ( \488_b0 , w_1275 );
and ( w_1274 , w_1275 , \242_b0 );
or ( \489_b1 , \487_b1 , w_1276 );
or ( \489_b0 , \487_b0 , \488_b0 );
not ( \488_b0 , w_1277 );
and ( w_1277 , w_1276 , \488_b1 );
or ( \490_b1 , \150_b1 , w_1279 );
not ( w_1279 , w_1280 );
and ( \490_b0 , \150_b0 , w_1281 );
and ( w_1280 ,  , w_1281 );
buf ( w_1279 , \437_b1 );
not ( w_1279 , w_1282 );
not (  , w_1283 );
and ( w_1282 , w_1283 , \437_b0 );
or ( \491_b1 , \489_b1 , w_1285 );
not ( w_1285 , w_1286 );
and ( \491_b0 , \489_b0 , w_1287 );
and ( w_1286 ,  , w_1287 );
buf ( w_1285 , \490_b1 );
not ( w_1285 , w_1288 );
not (  , w_1289 );
and ( w_1288 , w_1289 , \490_b0 );
buf ( \492_b1 , \491_b1 );
not ( \492_b1 , w_1290 );
not ( \492_b0 , w_1291 );
and ( w_1290 , w_1291 , \491_b0 );
buf ( \493_b1 , \471_b1 );
not ( \493_b1 , w_1292 );
not ( \493_b0 , w_1293 );
and ( w_1292 , w_1293 , \471_b0 );
buf ( \494_b1 , \464_b1 );
not ( \494_b1 , w_1294 );
not ( \494_b0 , w_1295 );
and ( w_1294 , w_1295 , \464_b0 );
or ( \495_b1 , \493_b1 , \494_b1 );
not ( \494_b1 , w_1296 );
and ( \495_b0 , \493_b0 , w_1297 );
and ( w_1296 , w_1297 , \494_b0 );
or ( \496_b1 , \471_b1 , \464_b1 );
not ( \464_b1 , w_1298 );
and ( \496_b0 , \471_b0 , w_1299 );
and ( w_1298 , w_1299 , \464_b0 );
or ( \497_b1 , \495_b1 , w_1301 );
not ( w_1301 , w_1302 );
and ( \497_b0 , \495_b0 , w_1303 );
and ( w_1302 ,  , w_1303 );
buf ( w_1301 , \496_b1 );
not ( w_1301 , w_1304 );
not (  , w_1305 );
and ( w_1304 , w_1305 , \496_b0 );
or ( \498_b1 , \492_b1 , w_1307 );
not ( w_1307 , w_1308 );
and ( \498_b0 , \492_b0 , w_1309 );
and ( w_1308 ,  , w_1309 );
buf ( w_1307 , \497_b1 );
not ( w_1307 , w_1310 );
not (  , w_1311 );
and ( w_1310 , w_1311 , \497_b0 );
or ( \499_b1 , \a[1]_b1 , \b[1]_b1 );
xor ( \499_b0 , \a[1]_b0 , w_1312 );
not ( w_1312 , w_1313 );
and ( w_1313 , \b[1]_b1 , \b[1]_b0 );
buf ( \500_b1 , \499_b1 );
not ( \500_b1 , w_1314 );
not ( \500_b0 , w_1315 );
and ( w_1314 , w_1315 , \499_b0 );
buf ( \501_b1 , \133_b1 );
not ( \501_b1 , w_1316 );
not ( \501_b0 , w_1317 );
and ( w_1316 , w_1317 , \133_b0 );
or ( \502_b1 , \500_b1 , w_1318 );
or ( \502_b0 , \500_b0 , \501_b0 );
not ( \501_b0 , w_1319 );
and ( w_1319 , w_1318 , \501_b1 );
or ( \503_b1 , \466_b1 , w_1321 );
not ( w_1321 , w_1322 );
and ( \503_b0 , \466_b0 , w_1323 );
and ( w_1322 ,  , w_1323 );
buf ( w_1321 , \b[0]_b1 );
not ( w_1321 , w_1324 );
not (  , w_1325 );
and ( w_1324 , w_1325 , \b[0]_b0 );
or ( \504_b1 , \502_b1 , w_1327 );
not ( w_1327 , w_1328 );
and ( \504_b0 , \502_b0 , w_1329 );
and ( w_1328 ,  , w_1329 );
buf ( w_1327 , \503_b1 );
not ( w_1327 , w_1330 );
not (  , w_1331 );
and ( w_1330 , w_1331 , \503_b0 );
or ( \505_b1 , \144_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_1332 );
and ( \505_b0 , \144_b0 , w_1333 );
and ( w_1332 , w_1333 , \a[0]_b0 );
or ( \506_b1 , \504_b1 , w_1335 );
not ( w_1335 , w_1336 );
and ( \506_b0 , \504_b0 , w_1337 );
and ( w_1336 ,  , w_1337 );
buf ( w_1335 , \505_b1 );
not ( w_1335 , w_1338 );
not (  , w_1339 );
and ( w_1338 , w_1339 , \505_b0 );
or ( \507_b1 , \a[0]_b1 , w_1341 );
not ( w_1341 , w_1342 );
and ( \507_b0 , \a[0]_b0 , w_1343 );
and ( w_1342 ,  , w_1343 );
buf ( w_1341 , \b[0]_b1 );
not ( w_1341 , w_1344 );
not (  , w_1345 );
and ( w_1344 , w_1345 , \b[0]_b0 );
or ( \508_b1 , \507_b1 , w_1347 );
not ( w_1347 , w_1348 );
and ( \508_b0 , \507_b0 , w_1349 );
and ( w_1348 ,  , w_1349 );
buf ( w_1347 , \b[1]_b1 );
not ( w_1347 , w_1350 );
not (  , w_1351 );
and ( w_1350 , w_1351 , \b[1]_b0 );
or ( \509_b1 , \508_b1 , w_1353 );
not ( w_1353 , w_1354 );
and ( \509_b0 , \508_b0 , w_1355 );
and ( w_1354 ,  , w_1355 );
buf ( w_1353 , \a[0]_b1 );
not ( w_1353 , w_1356 );
not (  , w_1357 );
and ( w_1356 , w_1357 , \a[0]_b0 );
buf ( \510_b1 , \499_b1 );
not ( \510_b1 , w_1358 );
not ( \510_b0 , w_1359 );
and ( w_1358 , w_1359 , \499_b0 );
or ( \511_b1 , \510_b1 , w_1361 );
not ( w_1361 , w_1362 );
and ( \511_b0 , \510_b0 , w_1363 );
and ( w_1362 ,  , w_1363 );
buf ( w_1361 , \b[0]_b1 );
not ( w_1361 , w_1364 );
not (  , w_1365 );
and ( w_1364 , w_1365 , \b[0]_b0 );
or ( \512_b1 , \509_b1 , w_1367 );
not ( w_1367 , w_1368 );
and ( \512_b0 , \509_b0 , w_1369 );
and ( w_1368 ,  , w_1369 );
buf ( w_1367 , \511_b1 );
not ( w_1367 , w_1370 );
not (  , w_1371 );
and ( w_1370 , w_1371 , \511_b0 );
or ( \513_b1 , \506_b1 , w_1372 );
or ( \513_b0 , \506_b0 , \512_b0 );
not ( \512_b0 , w_1373 );
and ( w_1373 , w_1372 , \512_b1 );
or ( \514_b1 , \504_b1 , w_1375 );
not ( w_1375 , w_1376 );
and ( \514_b0 , \504_b0 , w_1377 );
and ( w_1376 ,  , w_1377 );
buf ( w_1375 , \505_b1 );
not ( w_1375 , w_1378 );
not (  , w_1379 );
and ( w_1378 , w_1379 , \505_b0 );
or ( \515_b1 , \513_b1 , w_1381 );
not ( w_1381 , w_1382 );
and ( \515_b0 , \513_b0 , w_1383 );
and ( w_1382 ,  , w_1383 );
buf ( w_1381 , \514_b1 );
not ( w_1381 , w_1384 );
not (  , w_1385 );
and ( w_1384 , w_1385 , \514_b0 );
or ( \516_b1 , \498_b1 , w_1387 );
not ( w_1387 , w_1388 );
and ( \516_b0 , \498_b0 , w_1389 );
and ( w_1388 ,  , w_1389 );
buf ( w_1387 , \515_b1 );
not ( w_1387 , w_1390 );
not (  , w_1391 );
and ( w_1390 , w_1391 , \515_b0 );
buf ( \517_b1 , \497_b1 );
not ( \517_b1 , w_1392 );
not ( \517_b0 , w_1393 );
and ( w_1392 , w_1393 , \497_b0 );
or ( \518_b1 , \517_b1 , w_1395 );
not ( w_1395 , w_1396 );
and ( \518_b0 , \517_b0 , w_1397 );
and ( w_1396 ,  , w_1397 );
buf ( w_1395 , \491_b1 );
not ( w_1395 , w_1398 );
not (  , w_1399 );
and ( w_1398 , w_1399 , \491_b0 );
or ( \519_b1 , \516_b1 , w_1401 );
not ( w_1401 , w_1402 );
and ( \519_b0 , \516_b0 , w_1403 );
and ( w_1402 ,  , w_1403 );
buf ( w_1401 , \518_b1 );
not ( w_1401 , w_1404 );
not (  , w_1405 );
and ( w_1404 , w_1405 , \518_b0 );
or ( \520_b1 , \485_b1 , w_1407 );
not ( w_1407 , w_1408 );
and ( \520_b0 , \485_b0 , w_1409 );
and ( w_1408 ,  , w_1409 );
buf ( w_1407 , \519_b1 );
not ( w_1407 , w_1410 );
not (  , w_1411 );
and ( w_1410 , w_1411 , \519_b0 );
buf ( \521_b1 , \483_b1 );
not ( \521_b1 , w_1412 );
not ( \521_b0 , w_1413 );
and ( w_1412 , w_1413 , \483_b0 );
buf ( \522_b1 , \472_b1 );
not ( \522_b1 , w_1414 );
not ( \522_b0 , w_1415 );
and ( w_1414 , w_1415 , \472_b0 );
or ( \523_b1 , \521_b1 , w_1417 );
not ( w_1417 , w_1418 );
and ( \523_b0 , \521_b0 , w_1419 );
and ( w_1418 ,  , w_1419 );
buf ( w_1417 , \522_b1 );
not ( w_1417 , w_1420 );
not (  , w_1421 );
and ( w_1420 , w_1421 , \522_b0 );
or ( \524_b1 , \520_b1 , w_1423 );
not ( w_1423 , w_1424 );
and ( \524_b0 , \520_b0 , w_1425 );
and ( w_1424 ,  , w_1425 );
buf ( w_1423 , \523_b1 );
not ( w_1423 , w_1426 );
not (  , w_1427 );
and ( w_1426 , w_1427 , \523_b0 );
buf ( \525_b1 , \524_b1 );
not ( \525_b1 , w_1428 );
not ( \525_b0 , w_1429 );
and ( w_1428 , w_1429 , \524_b0 );
or ( \526_b1 , \459_b1 , w_1430 );
or ( \526_b0 , \459_b0 , \525_b0 );
not ( \525_b0 , w_1431 );
and ( w_1431 , w_1430 , \525_b1 );
buf ( \527_b1 , \457_b1 );
not ( \527_b1 , w_1432 );
not ( \527_b0 , w_1433 );
and ( w_1432 , w_1433 , \457_b0 );
or ( \528_b1 , \527_b1 , w_1435 );
not ( w_1435 , w_1436 );
and ( \528_b0 , \527_b0 , w_1437 );
and ( w_1436 ,  , w_1437 );
buf ( w_1435 , \447_b1 );
not ( w_1435 , w_1438 );
not (  , w_1439 );
and ( w_1438 , w_1439 , \447_b0 );
or ( \529_b1 , \526_b1 , w_1441 );
not ( w_1441 , w_1442 );
and ( \529_b0 , \526_b0 , w_1443 );
and ( w_1442 ,  , w_1443 );
buf ( w_1441 , \528_b1 );
not ( w_1441 , w_1444 );
not (  , w_1445 );
and ( w_1444 , w_1445 , \528_b0 );
buf ( \530_b1 , \529_b1 );
not ( \530_b1 , w_1446 );
not ( \530_b0 , w_1447 );
and ( w_1446 , w_1447 , \529_b0 );
or ( \531_b1 , \376_b1 , w_1449 );
not ( w_1449 , w_1450 );
and ( \531_b0 , \376_b0 , w_1451 );
and ( w_1450 ,  , w_1451 );
buf ( w_1449 , \401_b1 );
not ( w_1449 , w_1452 );
not (  , w_1453 );
and ( w_1452 , w_1453 , \401_b0 );
or ( \533_b1 , \317_b1 , \322_b1 );
xor ( \533_b0 , \317_b0 , w_1454 );
not ( w_1454 , w_1455 );
and ( w_1455 , \322_b1 , \322_b0 );
or ( \534_b1 , \533_b1 , w_1456 );
xor ( \534_b0 , \533_b0 , w_1458 );
not ( w_1458 , w_1459 );
and ( w_1459 , w_1456 , w_1457 );
buf ( w_1456 , \319_b1 );
not ( w_1456 , w_1460 );
not ( w_1457 , w_1461 );
and ( w_1460 , w_1461 , \319_b0 );
or ( \535_b1 , \405_b1 , \407_b1 );
xor ( \535_b0 , \405_b0 , w_1462 );
not ( w_1462 , w_1463 );
and ( w_1463 , \407_b1 , \407_b0 );
or ( \536_b1 , \535_b1 , \415_b1 );
not ( \415_b1 , w_1464 );
and ( \536_b0 , \535_b0 , w_1465 );
and ( w_1464 , w_1465 , \415_b0 );
or ( \537_b1 , \405_b1 , \407_b1 );
not ( \407_b1 , w_1466 );
and ( \537_b0 , \405_b0 , w_1467 );
and ( w_1466 , w_1467 , \407_b0 );
or ( \538_b1 , \536_b1 , w_1468 );
or ( \538_b0 , \536_b0 , \537_b0 );
not ( \537_b0 , w_1469 );
and ( w_1469 , w_1468 , \537_b1 );
buf ( \539_b1 , \538_b1 );
not ( \539_b1 , w_1470 );
not ( \539_b0 , w_1471 );
and ( w_1470 , w_1471 , \538_b0 );
or ( \540_b1 , \534_b1 , w_1473 );
not ( w_1473 , w_1474 );
and ( \540_b0 , \534_b0 , w_1475 );
and ( w_1474 ,  , w_1475 );
buf ( w_1473 , \539_b1 );
not ( w_1473 , w_1476 );
not (  , w_1477 );
and ( w_1476 , w_1477 , \539_b0 );
buf ( \542_b1 , \541_b1 );
not ( \542_b1 , w_1478 );
not ( \542_b0 , w_1479 );
and ( w_1478 , w_1479 , \541_b0 );
or ( \543_b1 , \285_b1 , w_1480 );
or ( \543_b0 , \285_b0 , \542_b0 );
not ( \542_b0 , w_1481 );
and ( w_1481 , w_1480 , \542_b1 );
buf ( \544_b1 , \225_b1 );
not ( \544_b1 , w_1482 );
not ( \544_b0 , w_1483 );
and ( w_1482 , w_1483 , \225_b0 );
or ( \545_b1 , \283_b1 , w_1485 );
not ( w_1485 , w_1486 );
and ( \545_b0 , \283_b0 , w_1487 );
and ( w_1486 ,  , w_1487 );
buf ( w_1485 , \544_b1 );
not ( w_1485 , w_1488 );
not (  , w_1489 );
and ( w_1488 , w_1489 , \544_b0 );
buf ( \546_b1 , \326_b1 );
not ( \546_b1 , w_1490 );
not ( \546_b0 , w_1491 );
and ( w_1490 , w_1491 , \326_b0 );
buf ( \547_b1 , \294_b1 );
not ( \547_b1 , w_1492 );
not ( \547_b0 , w_1493 );
and ( w_1492 , w_1493 , \294_b0 );
or ( \548_b1 , \546_b1 , w_1494 );
or ( \548_b0 , \546_b0 , \547_b0 );
not ( \547_b0 , w_1495 );
and ( w_1495 , w_1494 , \547_b1 );
buf ( \549_b1 , \534_b1 );
not ( \549_b1 , w_1496 );
not ( \549_b0 , w_1497 );
and ( w_1496 , w_1497 , \534_b0 );
or ( \550_b1 , \549_b1 , w_1499 );
not ( w_1499 , w_1500 );
and ( \550_b0 , \549_b0 , w_1501 );
and ( w_1500 ,  , w_1501 );
buf ( w_1499 , \538_b1 );
not ( w_1499 , w_1502 );
not (  , w_1503 );
and ( w_1502 , w_1503 , \538_b0 );
or ( \551_b1 , \548_b1 , w_1505 );
not ( w_1505 , w_1506 );
and ( \551_b0 , \548_b0 , w_1507 );
and ( w_1506 ,  , w_1507 );
buf ( w_1505 , \550_b1 );
not ( w_1505 , w_1508 );
not (  , w_1509 );
and ( w_1508 , w_1509 , \550_b0 );
or ( \552_b1 , \294_b1 , w_1510 );
or ( \552_b0 , \294_b0 , \326_b0 );
not ( \326_b0 , w_1511 );
and ( w_1511 , w_1510 , \326_b1 );
or ( \554_b1 , \283_b1 , w_1513 );
not ( w_1513 , w_1514 );
and ( \554_b0 , \283_b0 , w_1515 );
and ( w_1514 ,  , w_1515 );
buf ( w_1513 , \544_b1 );
not ( w_1513 , w_1516 );
not (  , w_1517 );
and ( w_1516 , w_1517 , \544_b0 );
or ( \555_b1 , \553_b1 , w_1519 );
not ( w_1519 , w_1520 );
and ( \555_b0 , \553_b0 , w_1521 );
and ( w_1520 ,  , w_1521 );
buf ( w_1519 , \554_b1 );
not ( w_1519 , w_1522 );
not (  , w_1523 );
and ( w_1522 , w_1523 , \554_b0 );
or ( \556_b1 , \543_b1 , w_1525 );
not ( w_1525 , w_1526 );
and ( \556_b0 , \543_b0 , w_1527 );
and ( w_1526 ,  , w_1527 );
buf ( w_1525 , \555_b1 );
not ( w_1525 , w_1528 );
not (  , w_1529 );
and ( w_1528 , w_1529 , \555_b0 );
buf ( \557_b1 , \231_b1 );
not ( \557_b1 , w_1530 );
not ( \557_b0 , w_1531 );
and ( w_1530 , w_1531 , \231_b0 );
buf ( \558_b1 , \106_b1 );
not ( \558_b1 , w_1532 );
not ( \558_b0 , w_1533 );
and ( w_1532 , w_1533 , \106_b0 );
or ( \559_b1 , \557_b1 , w_1534 );
or ( \559_b0 , \557_b0 , \558_b0 );
not ( \558_b0 , w_1535 );
and ( w_1535 , w_1534 , \558_b1 );
or ( \560_b1 , \a[3]_b1 , \b[9]_b1 );
xor ( \560_b0 , \a[3]_b0 , w_1536 );
not ( w_1536 , w_1537 );
and ( w_1537 , \b[9]_b1 , \b[9]_b0 );
or ( \561_b1 , \104_b1 , w_1539 );
not ( w_1539 , w_1540 );
and ( \561_b0 , \104_b0 , w_1541 );
and ( w_1540 ,  , w_1541 );
buf ( w_1539 , \560_b1 );
not ( w_1539 , w_1542 );
not (  , w_1543 );
and ( w_1542 , w_1543 , \560_b0 );
or ( \562_b1 , \559_b1 , w_1545 );
not ( w_1545 , w_1546 );
and ( \562_b0 , \559_b0 , w_1547 );
and ( w_1546 ,  , w_1547 );
buf ( w_1545 , \561_b1 );
not ( w_1545 , w_1548 );
not (  , w_1549 );
and ( w_1548 , w_1549 , \561_b0 );
buf ( \563_b1 , \562_b1 );
not ( \563_b1 , w_1550 );
not ( \563_b0 , w_1551 );
and ( w_1550 , w_1551 , \562_b0 );
buf ( \564_b1 , \245_b1 );
not ( \564_b1 , w_1552 );
not ( \564_b0 , w_1553 );
and ( w_1552 , w_1553 , \245_b0 );
buf ( \565_b1 , \242_b1 );
not ( \565_b1 , w_1554 );
not ( \565_b0 , w_1555 );
and ( w_1554 , w_1555 , \242_b0 );
or ( \566_b1 , \564_b1 , w_1556 );
or ( \566_b0 , \564_b0 , \565_b0 );
not ( \565_b0 , w_1557 );
and ( w_1557 , w_1556 , \565_b1 );
buf ( \567_b1 , \b[3]_b1 );
not ( \567_b1 , w_1558 );
not ( \567_b0 , w_1559 );
and ( w_1558 , w_1559 , \b[3]_b0 );
or ( \568_b1 , \567_b1 , w_1561 );
not ( w_1561 , w_1562 );
and ( \568_b0 , \567_b0 , w_1563 );
and ( w_1562 ,  , w_1563 );
buf ( w_1561 , \a[9]_b1 );
not ( w_1561 , w_1564 );
not (  , w_1565 );
and ( w_1564 , w_1565 , \a[9]_b0 );
buf ( \569_b1 , \568_b1 );
not ( \569_b1 , w_1566 );
not ( \569_b0 , w_1567 );
and ( w_1566 , w_1567 , \568_b0 );
buf ( \570_b1 , \a[9]_b1 );
not ( \570_b1 , w_1568 );
not ( \570_b0 , w_1569 );
and ( w_1568 , w_1569 , \a[9]_b0 );
or ( \571_b1 , \570_b1 , w_1571 );
not ( w_1571 , w_1572 );
and ( \571_b0 , \570_b0 , w_1573 );
and ( w_1572 ,  , w_1573 );
buf ( w_1571 , \b[3]_b1 );
not ( w_1571 , w_1574 );
not (  , w_1575 );
and ( w_1574 , w_1575 , \b[3]_b0 );
buf ( \572_b1 , \571_b1 );
not ( \572_b1 , w_1576 );
not ( \572_b0 , w_1577 );
and ( w_1576 , w_1577 , \571_b0 );
or ( \573_b1 , \569_b1 , w_1578 );
or ( \573_b0 , \569_b0 , \572_b0 );
not ( \572_b0 , w_1579 );
and ( w_1579 , w_1578 , \572_b1 );
or ( \574_b1 , \573_b1 , w_1581 );
not ( w_1581 , w_1582 );
and ( \574_b0 , \573_b0 , w_1583 );
and ( w_1582 ,  , w_1583 );
buf ( w_1581 , \150_b1 );
not ( w_1581 , w_1584 );
not (  , w_1585 );
and ( w_1584 , w_1585 , \150_b0 );
or ( \575_b1 , \566_b1 , w_1587 );
not ( w_1587 , w_1588 );
and ( \575_b0 , \566_b0 , w_1589 );
and ( w_1588 ,  , w_1589 );
buf ( w_1587 , \574_b1 );
not ( w_1587 , w_1590 );
not (  , w_1591 );
and ( w_1590 , w_1591 , \574_b0 );
or ( \576_b1 , \563_b1 , \575_b1 );
xor ( \576_b0 , \563_b0 , w_1592 );
not ( w_1592 , w_1593 );
and ( w_1593 , \575_b1 , \575_b0 );
or ( \577_b1 , \b[11]_b1 , \b[10]_b1 );
xor ( \577_b0 , \b[11]_b0 , w_1594 );
not ( w_1594 , w_1595 );
and ( w_1595 , \b[10]_b1 , \b[10]_b0 );
or ( \578_b1 , \a[0]_b1 , \b[11]_b1 );
xor ( \578_b0 , \a[0]_b0 , w_1596 );
not ( w_1596 , w_1597 );
and ( w_1597 , \b[11]_b1 , \b[11]_b0 );
or ( \579_b1 , \577_b1 , w_1599 );
not ( w_1599 , w_1600 );
and ( \579_b0 , \577_b0 , w_1601 );
and ( w_1600 ,  , w_1601 );
buf ( w_1599 , \578_b1 );
not ( w_1599 , w_1602 );
not (  , w_1603 );
and ( w_1602 , w_1603 , \578_b0 );
or ( \580_b1 , \579_b1 , w_1604 );
or ( \580_b0 , \579_b0 , \257_b0 );
not ( \257_b0 , w_1605 );
and ( w_1605 , w_1604 , \257_b1 );
or ( \581_b1 , \a[1]_b1 , \b[11]_b1 );
xor ( \581_b0 , \a[1]_b0 , w_1606 );
not ( w_1606 , w_1607 );
and ( w_1607 , \b[11]_b1 , \b[11]_b0 );
or ( \582_b1 , \257_b1 , w_1609 );
not ( w_1609 , w_1610 );
and ( \582_b0 , \257_b0 , w_1611 );
and ( w_1610 ,  , w_1611 );
buf ( w_1609 , \581_b1 );
not ( w_1609 , w_1612 );
not (  , w_1613 );
and ( w_1612 , w_1613 , \581_b0 );
or ( \583_b1 , \580_b1 , w_1615 );
not ( w_1615 , w_1616 );
and ( \583_b0 , \580_b0 , w_1617 );
and ( w_1616 ,  , w_1617 );
buf ( w_1615 , \582_b1 );
not ( w_1615 , w_1618 );
not (  , w_1619 );
and ( w_1618 , w_1619 , \582_b0 );
or ( \584_b1 , \a[0]_b1 , w_1620 );
or ( \584_b0 , \a[0]_b0 , \b[10]_b0 );
not ( \b[10]_b0 , w_1621 );
and ( w_1621 , w_1620 , \b[10]_b1 );
or ( \585_b1 , \584_b1 , w_1623 );
not ( w_1623 , w_1624 );
and ( \585_b0 , \584_b0 , w_1625 );
and ( w_1624 ,  , w_1625 );
buf ( w_1623 , \b[9]_b1 );
not ( w_1623 , w_1626 );
not (  , w_1627 );
and ( w_1626 , w_1627 , \b[9]_b0 );
or ( \586_b1 , \a[0]_b1 , w_1629 );
not ( w_1629 , w_1630 );
and ( \586_b0 , \a[0]_b0 , w_1631 );
and ( w_1630 ,  , w_1631 );
buf ( w_1629 , \b[10]_b1 );
not ( w_1629 , w_1632 );
not (  , w_1633 );
and ( w_1632 , w_1633 , \b[10]_b0 );
buf ( \588_b1 , \587_b1 );
not ( \588_b1 , w_1634 );
not ( \588_b0 , w_1635 );
and ( w_1634 , w_1635 , \587_b0 );
or ( \589_b1 , \583_b1 , \588_b1 );
not ( \588_b1 , w_1636 );
and ( \589_b0 , \583_b0 , w_1637 );
and ( w_1636 , w_1637 , \588_b0 );
buf ( \590_b1 , \583_b1 );
not ( \590_b1 , w_1638 );
not ( \590_b0 , w_1639 );
and ( w_1638 , w_1639 , \583_b0 );
or ( \591_b1 , \590_b1 , \587_b1 );
not ( \587_b1 , w_1640 );
and ( \591_b0 , \590_b0 , w_1641 );
and ( w_1640 , w_1641 , \587_b0 );
or ( \592_b1 , \589_b1 , w_1643 );
not ( w_1643 , w_1644 );
and ( \592_b0 , \589_b0 , w_1645 );
and ( w_1644 ,  , w_1645 );
buf ( w_1643 , \591_b1 );
not ( w_1643 , w_1646 );
not (  , w_1647 );
and ( w_1646 , w_1647 , \591_b0 );
buf ( \593_b1 , \262_b1 );
not ( \593_b1 , w_1648 );
not ( \593_b0 , w_1649 );
and ( w_1648 , w_1649 , \262_b0 );
buf ( \594_b1 , \133_b1 );
not ( \594_b1 , w_1650 );
not ( \594_b0 , w_1651 );
and ( w_1650 , w_1651 , \133_b0 );
or ( \595_b1 , \593_b1 , w_1652 );
or ( \595_b0 , \593_b0 , \594_b0 );
not ( \594_b0 , w_1653 );
and ( w_1653 , w_1652 , \594_b1 );
or ( \596_b1 , \a[11]_b1 , \b[1]_b1 );
xor ( \596_b0 , \a[11]_b0 , w_1654 );
not ( w_1654 , w_1655 );
and ( w_1655 , \b[1]_b1 , \b[1]_b0 );
or ( \597_b1 , \596_b1 , w_1657 );
not ( w_1657 , w_1658 );
and ( \597_b0 , \596_b0 , w_1659 );
and ( w_1658 ,  , w_1659 );
buf ( w_1657 , \b[0]_b1 );
not ( w_1657 , w_1660 );
not (  , w_1661 );
and ( w_1660 , w_1661 , \b[0]_b0 );
or ( \598_b1 , \595_b1 , w_1663 );
not ( w_1663 , w_1664 );
and ( \598_b0 , \595_b0 , w_1665 );
and ( w_1664 ,  , w_1665 );
buf ( w_1663 , \597_b1 );
not ( w_1663 , w_1666 );
not (  , w_1667 );
and ( w_1666 , w_1667 , \597_b0 );
or ( \599_b1 , \592_b1 , w_1668 );
xor ( \599_b0 , \592_b0 , w_1670 );
not ( w_1670 , w_1671 );
and ( w_1671 , w_1668 , w_1669 );
buf ( w_1668 , \598_b1 );
not ( w_1668 , w_1672 );
not ( w_1669 , w_1673 );
and ( w_1672 , w_1673 , \598_b0 );
or ( \600_b1 , \576_b1 , w_1674 );
xor ( \600_b0 , \576_b0 , w_1676 );
not ( w_1676 , w_1677 );
and ( w_1677 , w_1674 , w_1675 );
buf ( w_1674 , \599_b1 );
not ( w_1674 , w_1678 );
not ( w_1675 , w_1679 );
and ( w_1678 , w_1679 , \599_b0 );
buf ( \601_b1 , \237_b1 );
not ( \601_b1 , w_1680 );
not ( \601_b0 , w_1681 );
and ( w_1680 , w_1681 , \237_b0 );
buf ( \602_b1 , \178_b1 );
not ( \602_b1 , w_1682 );
not ( \602_b0 , w_1683 );
and ( w_1682 , w_1683 , \178_b0 );
or ( \603_b1 , \601_b1 , w_1684 );
or ( \603_b0 , \601_b0 , \602_b0 );
not ( \602_b0 , w_1685 );
and ( w_1685 , w_1684 , \602_b1 );
or ( \604_b1 , \a[5]_b1 , \b[7]_b1 );
xor ( \604_b0 , \a[5]_b0 , w_1686 );
not ( w_1686 , w_1687 );
and ( w_1687 , \b[7]_b1 , \b[7]_b0 );
or ( \605_b1 , \177_b1 , w_1689 );
not ( w_1689 , w_1690 );
and ( \605_b0 , \177_b0 , w_1691 );
and ( w_1690 ,  , w_1691 );
buf ( w_1689 , \604_b1 );
not ( w_1689 , w_1692 );
not (  , w_1693 );
and ( w_1692 , w_1693 , \604_b0 );
or ( \606_b1 , \603_b1 , w_1695 );
not ( w_1695 , w_1696 );
and ( \606_b0 , \603_b0 , w_1697 );
and ( w_1696 ,  , w_1697 );
buf ( w_1695 , \605_b1 );
not ( w_1695 , w_1698 );
not (  , w_1699 );
and ( w_1698 , w_1699 , \605_b0 );
buf ( \607_b1 , \270_b1 );
not ( \607_b1 , w_1700 );
not ( \607_b0 , w_1701 );
and ( w_1700 , w_1701 , \270_b0 );
buf ( \608_b1 , \198_b1 );
not ( \608_b1 , w_1702 );
not ( \608_b0 , w_1703 );
and ( w_1702 , w_1703 , \198_b0 );
or ( \609_b1 , \607_b1 , w_1704 );
or ( \609_b0 , \607_b0 , \608_b0 );
not ( \608_b0 , w_1705 );
and ( w_1705 , w_1704 , \608_b1 );
or ( \610_b1 , \a[7]_b1 , \b[5]_b1 );
xor ( \610_b0 , \a[7]_b0 , w_1706 );
not ( w_1706 , w_1707 );
and ( w_1707 , \b[5]_b1 , \b[5]_b0 );
or ( \611_b1 , \121_b1 , w_1709 );
not ( w_1709 , w_1710 );
and ( \611_b0 , \121_b0 , w_1711 );
and ( w_1710 ,  , w_1711 );
buf ( w_1709 , \610_b1 );
not ( w_1709 , w_1712 );
not (  , w_1713 );
and ( w_1712 , w_1713 , \610_b0 );
or ( \612_b1 , \609_b1 , w_1715 );
not ( w_1715 , w_1716 );
and ( \612_b0 , \609_b0 , w_1717 );
and ( w_1716 ,  , w_1717 );
buf ( w_1715 , \611_b1 );
not ( w_1715 , w_1718 );
not (  , w_1719 );
and ( w_1718 , w_1719 , \611_b0 );
buf ( \613_b1 , \612_b1 );
not ( \613_b1 , w_1720 );
not ( \613_b0 , w_1721 );
and ( w_1720 , w_1721 , \612_b0 );
or ( \614_b1 , \606_b1 , \613_b1 );
xor ( \614_b0 , \606_b0 , w_1722 );
not ( w_1722 , w_1723 );
and ( w_1723 , \613_b1 , \613_b0 );
or ( \615_b1 , \600_b1 , \614_b1 );
not ( \614_b1 , w_1724 );
and ( \615_b0 , \600_b0 , w_1725 );
and ( w_1724 , w_1725 , \614_b0 );
buf ( \616_b1 , \600_b1 );
not ( \616_b1 , w_1726 );
not ( \616_b0 , w_1727 );
and ( w_1726 , w_1727 , \600_b0 );
buf ( \617_b1 , \614_b1 );
not ( \617_b1 , w_1728 );
not ( \617_b0 , w_1729 );
and ( w_1728 , w_1729 , \614_b0 );
or ( \618_b1 , \616_b1 , \617_b1 );
not ( \617_b1 , w_1730 );
and ( \618_b0 , \616_b0 , w_1731 );
and ( w_1730 , w_1731 , \617_b0 );
or ( \619_b1 , \615_b1 , w_1733 );
not ( w_1733 , w_1734 );
and ( \619_b0 , \615_b0 , w_1735 );
and ( w_1734 ,  , w_1735 );
buf ( w_1733 , \618_b1 );
not ( w_1733 , w_1736 );
not (  , w_1737 );
and ( w_1736 , w_1737 , \618_b0 );
or ( \620_b1 , \233_b1 , \239_b1 );
xor ( \620_b0 , \233_b0 , w_1738 );
not ( w_1738 , w_1739 );
and ( w_1739 , \239_b1 , \239_b0 );
or ( \621_b1 , \620_b1 , \247_b1 );
not ( \247_b1 , w_1740 );
and ( \621_b0 , \620_b0 , w_1741 );
and ( w_1740 , w_1741 , \247_b0 );
or ( \622_b1 , \233_b1 , \239_b1 );
not ( \239_b1 , w_1742 );
and ( \622_b0 , \233_b0 , w_1743 );
and ( w_1742 , w_1743 , \239_b0 );
or ( \623_b1 , \621_b1 , w_1744 );
or ( \623_b0 , \621_b0 , \622_b0 );
not ( \622_b0 , w_1745 );
and ( w_1745 , w_1744 , \622_b1 );
or ( \624_b1 , \258_b1 , \264_b1 );
xor ( \624_b0 , \258_b0 , w_1746 );
not ( w_1746 , w_1747 );
and ( w_1747 , \264_b1 , \264_b0 );
or ( \625_b1 , \624_b1 , \272_b1 );
not ( \272_b1 , w_1748 );
and ( \625_b0 , \624_b0 , w_1749 );
and ( w_1748 , w_1749 , \272_b0 );
or ( \626_b1 , \258_b1 , \264_b1 );
not ( \264_b1 , w_1750 );
and ( \626_b0 , \258_b0 , w_1751 );
and ( w_1750 , w_1751 , \264_b0 );
or ( \627_b1 , \625_b1 , w_1752 );
or ( \627_b0 , \625_b0 , \626_b0 );
not ( \626_b0 , w_1753 );
and ( w_1753 , w_1752 , \626_b1 );
or ( \628_b1 , \623_b1 , \627_b1 );
xor ( \628_b0 , \623_b0 , w_1754 );
not ( w_1754 , w_1755 );
and ( w_1755 , \627_b1 , \627_b0 );
or ( \629_b1 , \619_b1 , \628_b1 );
xor ( \629_b0 , \619_b0 , w_1756 );
not ( w_1756 , w_1757 );
and ( w_1757 , \628_b1 , \628_b0 );
or ( \630_b1 , \256_b1 , \273_b1 );
xor ( \630_b0 , \256_b0 , w_1758 );
not ( w_1758 , w_1759 );
and ( w_1759 , \273_b1 , \273_b0 );
or ( \631_b1 , \630_b1 , \281_b1 );
not ( \281_b1 , w_1760 );
and ( \631_b0 , \630_b0 , w_1761 );
and ( w_1760 , w_1761 , \281_b0 );
or ( \632_b1 , \256_b1 , \273_b1 );
not ( \273_b1 , w_1762 );
and ( \632_b0 , \256_b0 , w_1763 );
and ( w_1762 , w_1763 , \273_b0 );
or ( \633_b1 , \631_b1 , w_1764 );
or ( \633_b0 , \631_b0 , \632_b0 );
not ( \632_b0 , w_1765 );
and ( w_1765 , w_1764 , \632_b1 );
or ( \634_b1 , \629_b1 , \633_b1 );
xor ( \634_b0 , \629_b0 , w_1766 );
not ( w_1766 , w_1767 );
and ( w_1767 , \633_b1 , \633_b0 );
buf ( \635_b1 , \248_b1 );
buf ( \635_b0 , \248_b0 );
or ( \636_b1 , \254_b1 , w_1768 );
or ( \636_b0 , \254_b0 , \635_b0 );
not ( \635_b0 , w_1769 );
and ( w_1769 , w_1768 , \635_b1 );
buf ( \637_b1 , \636_b1 );
not ( \637_b1 , w_1770 );
not ( \637_b0 , w_1771 );
and ( w_1770 , w_1771 , \636_b0 );
buf ( \638_b1 , \282_b1 );
not ( \638_b1 , w_1772 );
not ( \638_b0 , w_1773 );
and ( w_1772 , w_1773 , \282_b0 );
or ( \639_b1 , \637_b1 , w_1774 );
or ( \639_b0 , \637_b0 , \638_b0 );
not ( \638_b0 , w_1775 );
and ( w_1775 , w_1774 , \638_b1 );
or ( \640_b1 , \254_b1 , w_1777 );
not ( w_1777 , w_1778 );
and ( \640_b0 , \254_b0 , w_1779 );
and ( w_1778 ,  , w_1779 );
buf ( w_1777 , \635_b1 );
not ( w_1777 , w_1780 );
not (  , w_1781 );
and ( w_1780 , w_1781 , \635_b0 );
or ( \641_b1 , \639_b1 , w_1783 );
not ( w_1783 , w_1784 );
and ( \641_b0 , \639_b0 , w_1785 );
and ( w_1784 ,  , w_1785 );
buf ( w_1783 , \640_b1 );
not ( w_1783 , w_1786 );
not (  , w_1787 );
and ( w_1786 , w_1787 , \640_b0 );
or ( \642_b1 , \634_b1 , \641_b1 );
xor ( \642_b0 , \634_b0 , w_1788 );
not ( w_1788 , w_1789 );
and ( w_1789 , \641_b1 , \641_b0 );
or ( \643_b1 , \556_b1 , \642_b1 );
xor ( \643_b0 , \556_b0 , w_1790 );
not ( w_1790 , w_1791 );
and ( w_1791 , \642_b1 , \642_b0 );
buf ( \644_b1 , \643_b1 );
buf ( \644_b0 , \643_b0 );
buf ( \645_b1 , \644_b1 );
not ( \645_b1 , w_1792 );
not ( \645_b0 , w_1793 );
and ( w_1792 , w_1793 , \644_b0 );
or ( \646_b1 , \101_b1 , w_1795 );
not ( w_1795 , w_1796 );
and ( \646_b0 , \101_b0 , w_1797 );
and ( w_1796 ,  , w_1797 );
buf ( w_1795 , \645_b1 );
not ( w_1795 , w_1798 );
not (  , w_1799 );
and ( w_1798 , w_1799 , \645_b0 );
buf ( \647_b1 , \b[7]_b1 );
not ( \647_b1 , w_1800 );
not ( \647_b0 , w_1801 );
and ( w_1800 , w_1801 , \b[7]_b0 );
buf ( \648_b1 , \a[7]_b1 );
not ( \648_b1 , w_1802 );
not ( \648_b0 , w_1803 );
and ( w_1802 , w_1803 , \a[7]_b0 );
or ( \649_b1 , \647_b1 , w_1805 );
not ( w_1805 , w_1806 );
and ( \649_b0 , \647_b0 , w_1807 );
and ( w_1806 ,  , w_1807 );
buf ( w_1805 , \648_b1 );
not ( w_1805 , w_1808 );
not (  , w_1809 );
and ( w_1808 , w_1809 , \648_b0 );
buf ( \650_b1 , \649_b1 );
not ( \650_b1 , w_1810 );
not ( \650_b0 , w_1811 );
and ( w_1810 , w_1811 , \649_b0 );
buf ( \651_b1 , \540_b1 );
not ( \651_b1 , w_1812 );
not ( \651_b0 , w_1813 );
and ( w_1812 , w_1813 , \540_b0 );
or ( \652_b1 , \416_b1 , w_1814 );
or ( \652_b0 , \416_b0 , \422_b0 );
not ( \422_b0 , w_1815 );
and ( w_1815 , w_1814 , \422_b1 );
buf ( \653_b1 , \652_b1 );
not ( \653_b1 , w_1816 );
not ( \653_b0 , w_1817 );
and ( w_1816 , w_1817 , \652_b0 );
or ( \654_b1 , \423_b1 , w_1819 );
not ( w_1819 , w_1820 );
and ( \654_b0 , \423_b0 , w_1821 );
and ( w_1820 ,  , w_1821 );
buf ( w_1819 , \531_b1 );
not ( w_1819 , w_1822 );
not (  , w_1823 );
and ( w_1822 , w_1823 , \531_b0 );
buf ( \655_b1 , \654_b1 );
not ( \655_b1 , w_1824 );
not ( \655_b0 , w_1825 );
and ( w_1824 , w_1825 , \654_b0 );
or ( \656_b1 , \653_b1 , w_1826 );
or ( \656_b0 , \653_b0 , \655_b0 );
not ( \655_b0 , w_1827 );
and ( w_1827 , w_1826 , \655_b1 );
or ( \658_b1 , \656_b1 , w_1829 );
not ( w_1829 , w_1830 );
and ( \658_b0 , \656_b0 , w_1831 );
and ( w_1830 ,  , w_1831 );
buf ( w_1829 , \657_b1 );
not ( w_1829 , w_1832 );
not (  , w_1833 );
and ( w_1832 , w_1833 , \657_b0 );
buf ( \659_b1 , \658_b1 );
not ( \659_b1 , w_1834 );
not ( \659_b0 , w_1835 );
and ( w_1834 , w_1835 , \658_b0 );
or ( \660_b1 , \651_b1 , w_1836 );
or ( \660_b0 , \651_b0 , \659_b0 );
not ( \659_b0 , w_1837 );
and ( w_1837 , w_1836 , \659_b1 );
or ( \661_b1 , \539_b1 , w_1839 );
not ( w_1839 , w_1840 );
and ( \661_b0 , \539_b0 , w_1841 );
and ( w_1840 ,  , w_1841 );
buf ( w_1839 , \534_b1 );
not ( w_1839 , w_1842 );
not (  , w_1843 );
and ( w_1842 , w_1843 , \534_b0 );
buf ( \662_b1 , \661_b1 );
not ( \662_b1 , w_1844 );
not ( \662_b0 , w_1845 );
and ( w_1844 , w_1845 , \661_b0 );
or ( \663_b1 , \660_b1 , w_1847 );
not ( w_1847 , w_1848 );
and ( \663_b0 , \660_b0 , w_1849 );
and ( w_1848 ,  , w_1849 );
buf ( w_1847 , \662_b1 );
not ( w_1847 , w_1850 );
not (  , w_1851 );
and ( w_1850 , w_1851 , \662_b0 );
or ( \664_b1 , \294_b1 , \326_b1 );
not ( \326_b1 , w_1852 );
and ( \664_b0 , \294_b0 , w_1853 );
and ( w_1852 , w_1853 , \326_b0 );
buf ( \665_b1 , \664_b1 );
not ( \665_b1 , w_1854 );
not ( \665_b0 , w_1855 );
and ( w_1854 , w_1855 , \664_b0 );
or ( \666_b1 , \665_b1 , w_1857 );
not ( w_1857 , w_1858 );
and ( \666_b0 , \665_b0 , w_1859 );
and ( w_1858 ,  , w_1859 );
buf ( w_1857 , \552_b1 );
not ( w_1857 , w_1860 );
not (  , w_1861 );
and ( w_1860 , w_1861 , \552_b0 );
buf ( \667_b1 , \666_b1 );
not ( \667_b1 , w_1862 );
not ( \667_b0 , w_1863 );
and ( w_1862 , w_1863 , \666_b0 );
or ( \668_b1 , \663_b1 , \667_b1 );
not ( \667_b1 , w_1864 );
and ( \668_b0 , \663_b0 , w_1865 );
and ( w_1864 , w_1865 , \667_b0 );
buf ( \669_b1 , \663_b1 );
not ( \669_b1 , w_1866 );
not ( \669_b0 , w_1867 );
and ( w_1866 , w_1867 , \663_b0 );
or ( \670_b1 , \669_b1 , \666_b1 );
not ( \666_b1 , w_1868 );
and ( \670_b0 , \669_b0 , w_1869 );
and ( w_1868 , w_1869 , \666_b0 );
or ( \671_b1 , \668_b1 , w_1871 );
not ( w_1871 , w_1872 );
and ( \671_b0 , \668_b0 , w_1873 );
and ( w_1872 ,  , w_1873 );
buf ( w_1871 , \670_b1 );
not ( w_1871 , w_1874 );
not (  , w_1875 );
and ( w_1874 , w_1875 , \670_b0 );
buf ( \672_b1 , \671_b1 );
buf ( \672_b0 , \671_b0 );
buf ( \673_b1 , \672_b1 );
not ( \673_b1 , w_1876 );
not ( \673_b0 , w_1877 );
and ( w_1876 , w_1877 , \672_b0 );
or ( \674_b1 , \650_b1 , w_1878 );
or ( \674_b0 , \650_b0 , \673_b0 );
not ( \673_b0 , w_1879 );
and ( w_1879 , w_1878 , \673_b1 );
or ( \675_b1 , \b[6]_b1 , \c[1]_b1 );
xor ( \675_b0 , \b[6]_b0 , w_1880 );
not ( w_1880 , w_1881 );
and ( w_1881 , \c[1]_b1 , \c[1]_b0 );
buf ( \676_b1 , \675_b1 );
not ( \676_b1 , w_1882 );
not ( \676_b0 , w_1883 );
and ( w_1882 , w_1883 , \675_b0 );
buf ( \677_b1 , \c[0]_b1 );
not ( \677_b1 , w_1884 );
not ( \677_b0 , w_1885 );
and ( w_1884 , w_1885 , \c[0]_b0 );
or ( \678_b1 , \677_b1 , w_1887 );
not ( w_1887 , w_1888 );
and ( \678_b0 , \677_b0 , w_1889 );
and ( w_1888 ,  , w_1889 );
buf ( w_1887 , \c[1]_b1 );
not ( w_1887 , w_1890 );
not (  , w_1891 );
and ( w_1890 , w_1891 , \c[1]_b0 );
buf ( \679_b1 , \678_b1 );
not ( \679_b1 , w_1892 );
not ( \679_b0 , w_1893 );
and ( w_1892 , w_1893 , \678_b0 );
buf ( \680_b1 , \679_b1 );
not ( \680_b1 , w_1894 );
not ( \680_b0 , w_1895 );
and ( w_1894 , w_1895 , \679_b0 );
or ( \681_b1 , \676_b1 , w_1896 );
or ( \681_b0 , \676_b0 , \680_b0 );
not ( \680_b0 , w_1897 );
and ( w_1897 , w_1896 , \680_b1 );
or ( \682_b1 , \b[7]_b1 , \c[1]_b1 );
xor ( \682_b0 , \b[7]_b0 , w_1898 );
not ( w_1898 , w_1899 );
and ( w_1899 , \c[1]_b1 , \c[1]_b0 );
or ( \683_b1 , \682_b1 , w_1901 );
not ( w_1901 , w_1902 );
and ( \683_b0 , \682_b0 , w_1903 );
and ( w_1902 ,  , w_1903 );
buf ( w_1901 , \c[0]_b1 );
not ( w_1901 , w_1904 );
not (  , w_1905 );
and ( w_1904 , w_1905 , \c[0]_b0 );
or ( \684_b1 , \681_b1 , w_1907 );
not ( w_1907 , w_1908 );
and ( \684_b0 , \681_b0 , w_1909 );
and ( w_1908 ,  , w_1909 );
buf ( w_1907 , \683_b1 );
not ( w_1907 , w_1910 );
not (  , w_1911 );
and ( w_1910 , w_1911 , \683_b0 );
buf ( \685_b1 , \684_b1 );
not ( \685_b1 , w_1912 );
not ( \685_b0 , w_1913 );
and ( w_1912 , w_1913 , \684_b0 );
or ( \686_b1 , \b[0]_b1 , w_1914 );
or ( \686_b0 , \b[0]_b0 , \c[6]_b0 );
not ( \c[6]_b0 , w_1915 );
and ( w_1915 , w_1914 , \c[6]_b1 );
or ( \687_b1 , \686_b1 , w_1917 );
not ( w_1917 , w_1918 );
and ( \687_b0 , \686_b0 , w_1919 );
and ( w_1918 ,  , w_1919 );
buf ( w_1917 , \c[5]_b1 );
not ( w_1917 , w_1920 );
not (  , w_1921 );
and ( w_1920 , w_1921 , \c[5]_b0 );
or ( \688_b1 , \b[0]_b1 , w_1923 );
not ( w_1923 , w_1924 );
and ( \688_b0 , \b[0]_b0 , w_1925 );
and ( w_1924 ,  , w_1925 );
buf ( w_1923 , \c[6]_b1 );
not ( w_1923 , w_1926 );
not (  , w_1927 );
and ( w_1926 , w_1927 , \c[6]_b0 );
buf ( \690_b1 , \689_b1 );
not ( \690_b1 , w_1928 );
not ( \690_b0 , w_1929 );
and ( w_1928 , w_1929 , \689_b0 );
or ( \691_b1 , \685_b1 , \690_b1 );
not ( \690_b1 , w_1930 );
and ( \691_b0 , \685_b0 , w_1931 );
and ( w_1930 , w_1931 , \690_b0 );
or ( \692_b1 , \684_b1 , \689_b1 );
not ( \689_b1 , w_1932 );
and ( \692_b0 , \684_b0 , w_1933 );
and ( w_1932 , w_1933 , \689_b0 );
or ( \693_b1 , \691_b1 , w_1935 );
not ( w_1935 , w_1936 );
and ( \693_b0 , \691_b0 , w_1937 );
and ( w_1936 ,  , w_1937 );
buf ( w_1935 , \692_b1 );
not ( w_1935 , w_1938 );
not (  , w_1939 );
and ( w_1938 , w_1939 , \692_b0 );
or ( \694_b1 , \b[3]_b1 , \c[3]_b1 );
xor ( \694_b0 , \b[3]_b0 , w_1940 );
not ( w_1940 , w_1941 );
and ( w_1941 , \c[3]_b1 , \c[3]_b0 );
buf ( \695_b1 , \694_b1 );
not ( \695_b1 , w_1942 );
not ( \695_b0 , w_1943 );
and ( w_1942 , w_1943 , \694_b0 );
or ( \696_b1 , \c[3]_b1 , \c[2]_b1 );
xor ( \696_b0 , \c[3]_b0 , w_1944 );
not ( w_1944 , w_1945 );
and ( w_1945 , \c[2]_b1 , \c[2]_b0 );
buf ( \697_b1 , \696_b1 );
not ( \697_b1 , w_1946 );
not ( \697_b0 , w_1947 );
and ( w_1946 , w_1947 , \696_b0 );
or ( \698_b1 , \c[2]_b1 , \c[1]_b1 );
xor ( \698_b0 , \c[2]_b0 , w_1948 );
not ( w_1948 , w_1949 );
and ( w_1949 , \c[1]_b1 , \c[1]_b0 );
or ( \699_b1 , \697_b1 , w_1951 );
not ( w_1951 , w_1952 );
and ( \699_b0 , \697_b0 , w_1953 );
and ( w_1952 ,  , w_1953 );
buf ( w_1951 , \698_b1 );
not ( w_1951 , w_1954 );
not (  , w_1955 );
and ( w_1954 , w_1955 , \698_b0 );
buf ( \700_b1 , \699_b1 );
not ( \700_b1 , w_1956 );
not ( \700_b0 , w_1957 );
and ( w_1956 , w_1957 , \699_b0 );
or ( \701_b1 , \695_b1 , w_1958 );
or ( \701_b0 , \695_b0 , \700_b0 );
not ( \700_b0 , w_1959 );
and ( w_1959 , w_1958 , \700_b1 );
buf ( \702_b1 , \698_b1 );
buf ( \702_b0 , \698_b0 );
or ( \703_b1 , \b[4]_b1 , \c[3]_b1 );
xor ( \703_b0 , \b[4]_b0 , w_1960 );
not ( w_1960 , w_1961 );
and ( w_1961 , \c[3]_b1 , \c[3]_b0 );
or ( \704_b1 , \702_b1 , w_1963 );
not ( w_1963 , w_1964 );
and ( \704_b0 , \702_b0 , w_1965 );
and ( w_1964 ,  , w_1965 );
buf ( w_1963 , \703_b1 );
not ( w_1963 , w_1966 );
not (  , w_1967 );
and ( w_1966 , w_1967 , \703_b0 );
or ( \705_b1 , \701_b1 , w_1969 );
not ( w_1969 , w_1970 );
and ( \705_b0 , \701_b0 , w_1971 );
and ( w_1970 ,  , w_1971 );
buf ( w_1969 , \704_b1 );
not ( w_1969 , w_1972 );
not (  , w_1973 );
and ( w_1972 , w_1973 , \704_b0 );
buf ( \706_b1 , \705_b1 );
not ( \706_b1 , w_1974 );
not ( \706_b0 , w_1975 );
and ( w_1974 , w_1975 , \705_b0 );
or ( \707_b1 , \b[5]_b1 , \c[1]_b1 );
xor ( \707_b0 , \b[5]_b0 , w_1976 );
not ( w_1976 , w_1977 );
and ( w_1977 , \c[1]_b1 , \c[1]_b0 );
buf ( \708_b1 , \707_b1 );
not ( \708_b1 , w_1978 );
not ( \708_b0 , w_1979 );
and ( w_1978 , w_1979 , \707_b0 );
buf ( \709_b1 , \679_b1 );
not ( \709_b1 , w_1980 );
not ( \709_b0 , w_1981 );
and ( w_1980 , w_1981 , \679_b0 );
or ( \710_b1 , \708_b1 , w_1982 );
or ( \710_b0 , \708_b0 , \709_b0 );
not ( \709_b0 , w_1983 );
and ( w_1983 , w_1982 , \709_b1 );
or ( \711_b1 , \675_b1 , w_1985 );
not ( w_1985 , w_1986 );
and ( \711_b0 , \675_b0 , w_1987 );
and ( w_1986 ,  , w_1987 );
buf ( w_1985 , \c[0]_b1 );
not ( w_1985 , w_1988 );
not (  , w_1989 );
and ( w_1988 , w_1989 , \c[0]_b0 );
or ( \712_b1 , \710_b1 , w_1991 );
not ( w_1991 , w_1992 );
and ( \712_b0 , \710_b0 , w_1993 );
and ( w_1992 ,  , w_1993 );
buf ( w_1991 , \711_b1 );
not ( w_1991 , w_1994 );
not (  , w_1995 );
and ( w_1994 , w_1995 , \711_b0 );
or ( \713_b1 , \c[6]_b1 , \c[5]_b1 );
xor ( \713_b0 , \c[6]_b0 , w_1996 );
not ( w_1996 , w_1997 );
and ( w_1997 , \c[5]_b1 , \c[5]_b0 );
buf ( \714_b1 , \713_b1 );
buf ( \714_b0 , \713_b0 );
or ( \715_b1 , \714_b1 , w_1999 );
not ( w_1999 , w_2000 );
and ( \715_b0 , \714_b0 , w_2001 );
and ( w_2000 ,  , w_2001 );
buf ( w_1999 , \b[0]_b1 );
not ( w_1999 , w_2002 );
not (  , w_2003 );
and ( w_2002 , w_2003 , \b[0]_b0 );
buf ( \716_b1 , \715_b1 );
not ( \716_b1 , w_2004 );
not ( \716_b0 , w_2005 );
and ( w_2004 , w_2005 , \715_b0 );
or ( \717_b1 , \712_b1 , w_2006 );
or ( \717_b0 , \712_b0 , \716_b0 );
not ( \716_b0 , w_2007 );
and ( w_2007 , w_2006 , \716_b1 );
buf ( \718_b1 , \717_b1 );
not ( \718_b1 , w_2008 );
not ( \718_b0 , w_2009 );
and ( w_2008 , w_2009 , \717_b0 );
or ( \719_b1 , \706_b1 , w_2010 );
or ( \719_b0 , \706_b0 , \718_b0 );
not ( \718_b0 , w_2011 );
and ( w_2011 , w_2010 , \718_b1 );
or ( \720_b1 , \712_b1 , w_2013 );
not ( w_2013 , w_2014 );
and ( \720_b0 , \712_b0 , w_2015 );
and ( w_2014 ,  , w_2015 );
buf ( w_2013 , \716_b1 );
not ( w_2013 , w_2016 );
not (  , w_2017 );
and ( w_2016 , w_2017 , \716_b0 );
or ( \721_b1 , \719_b1 , w_2019 );
not ( w_2019 , w_2020 );
and ( \721_b0 , \719_b0 , w_2021 );
and ( w_2020 ,  , w_2021 );
buf ( w_2019 , \720_b1 );
not ( w_2019 , w_2022 );
not (  , w_2023 );
and ( w_2022 , w_2023 , \720_b0 );
or ( \722_b1 , \693_b1 , \721_b1 );
xor ( \722_b0 , \693_b0 , w_2024 );
not ( w_2024 , w_2025 );
and ( w_2025 , \721_b1 , \721_b0 );
or ( \723_b1 , \b[0]_b1 , \c[7]_b1 );
xor ( \723_b0 , \b[0]_b0 , w_2026 );
not ( w_2026 , w_2027 );
and ( w_2027 , \c[7]_b1 , \c[7]_b0 );
buf ( \724_b1 , \723_b1 );
not ( \724_b1 , w_2028 );
not ( \724_b0 , w_2029 );
and ( w_2028 , w_2029 , \723_b0 );
or ( \725_b1 , \c[7]_b1 , w_2030 );
xor ( \725_b0 , \c[7]_b0 , w_2032 );
not ( w_2032 , w_2033 );
and ( w_2033 , w_2030 , w_2031 );
buf ( w_2030 , \c[6]_b1 );
not ( w_2030 , w_2034 );
not ( w_2031 , w_2035 );
and ( w_2034 , w_2035 , \c[6]_b0 );
or ( \726_b1 , \725_b1 , w_2037 );
not ( w_2037 , w_2038 );
and ( \726_b0 , \725_b0 , w_2039 );
and ( w_2038 ,  , w_2039 );
buf ( w_2037 , \713_b1 );
not ( w_2037 , w_2040 );
not (  , w_2041 );
and ( w_2040 , w_2041 , \713_b0 );
buf ( \727_b1 , \726_b1 );
not ( \727_b1 , w_2042 );
not ( \727_b0 , w_2043 );
and ( w_2042 , w_2043 , \726_b0 );
or ( \728_b1 , \724_b1 , w_2044 );
or ( \728_b0 , \724_b0 , \727_b0 );
not ( \727_b0 , w_2045 );
and ( w_2045 , w_2044 , \727_b1 );
or ( \729_b1 , \b[1]_b1 , \c[7]_b1 );
xor ( \729_b0 , \b[1]_b0 , w_2046 );
not ( w_2046 , w_2047 );
and ( w_2047 , \c[7]_b1 , \c[7]_b0 );
or ( \730_b1 , \714_b1 , w_2049 );
not ( w_2049 , w_2050 );
and ( \730_b0 , \714_b0 , w_2051 );
and ( w_2050 ,  , w_2051 );
buf ( w_2049 , \729_b1 );
not ( w_2049 , w_2052 );
not (  , w_2053 );
and ( w_2052 , w_2053 , \729_b0 );
or ( \731_b1 , \728_b1 , w_2055 );
not ( w_2055 , w_2056 );
and ( \731_b0 , \728_b0 , w_2057 );
and ( w_2056 ,  , w_2057 );
buf ( w_2055 , \730_b1 );
not ( w_2055 , w_2058 );
not (  , w_2059 );
and ( w_2058 , w_2059 , \730_b0 );
or ( \732_b1 , \b[2]_b1 , \c[5]_b1 );
xor ( \732_b0 , \b[2]_b0 , w_2060 );
not ( w_2060 , w_2061 );
and ( w_2061 , \c[5]_b1 , \c[5]_b0 );
buf ( \733_b1 , \732_b1 );
not ( \733_b1 , w_2062 );
not ( \733_b0 , w_2063 );
and ( w_2062 , w_2063 , \732_b0 );
or ( \734_b1 , \c[4]_b1 , \c[3]_b1 );
xor ( \734_b0 , \c[4]_b0 , w_2064 );
not ( w_2064 , w_2065 );
and ( w_2065 , \c[3]_b1 , \c[3]_b0 );
or ( \735_b1 , \c[5]_b1 , w_2066 );
xor ( \735_b0 , \c[5]_b0 , w_2068 );
not ( w_2068 , w_2069 );
and ( w_2069 , w_2066 , w_2067 );
buf ( w_2066 , \c[4]_b1 );
not ( w_2066 , w_2070 );
not ( w_2067 , w_2071 );
and ( w_2070 , w_2071 , \c[4]_b0 );
or ( \736_b1 , \734_b1 , w_2073 );
not ( w_2073 , w_2074 );
and ( \736_b0 , \734_b0 , w_2075 );
and ( w_2074 ,  , w_2075 );
buf ( w_2073 , \735_b1 );
not ( w_2073 , w_2076 );
not (  , w_2077 );
and ( w_2076 , w_2077 , \735_b0 );
buf ( \737_b1 , \736_b1 );
not ( \737_b1 , w_2078 );
not ( \737_b0 , w_2079 );
and ( w_2078 , w_2079 , \736_b0 );
or ( \738_b1 , \733_b1 , w_2080 );
or ( \738_b0 , \733_b0 , \737_b0 );
not ( \737_b0 , w_2081 );
and ( w_2081 , w_2080 , \737_b1 );
or ( \739_b1 , \c[4]_b1 , \c[3]_b1 );
xor ( \739_b0 , \c[4]_b0 , w_2082 );
not ( w_2082 , w_2083 );
and ( w_2083 , \c[3]_b1 , \c[3]_b0 );
or ( \740_b1 , \b[3]_b1 , \c[5]_b1 );
xor ( \740_b0 , \b[3]_b0 , w_2084 );
not ( w_2084 , w_2085 );
and ( w_2085 , \c[5]_b1 , \c[5]_b0 );
or ( \741_b1 , \739_b1 , w_2087 );
not ( w_2087 , w_2088 );
and ( \741_b0 , \739_b0 , w_2089 );
and ( w_2088 ,  , w_2089 );
buf ( w_2087 , \740_b1 );
not ( w_2087 , w_2090 );
not (  , w_2091 );
and ( w_2090 , w_2091 , \740_b0 );
or ( \742_b1 , \738_b1 , w_2093 );
not ( w_2093 , w_2094 );
and ( \742_b0 , \738_b0 , w_2095 );
and ( w_2094 ,  , w_2095 );
buf ( w_2093 , \741_b1 );
not ( w_2093 , w_2096 );
not (  , w_2097 );
and ( w_2096 , w_2097 , \741_b0 );
or ( \743_b1 , \731_b1 , \742_b1 );
xor ( \743_b0 , \731_b0 , w_2098 );
not ( w_2098 , w_2099 );
and ( w_2099 , \742_b1 , \742_b0 );
buf ( \744_b1 , \703_b1 );
not ( \744_b1 , w_2100 );
not ( \744_b0 , w_2101 );
and ( w_2100 , w_2101 , \703_b0 );
buf ( \745_b1 , \696_b1 );
not ( \745_b1 , w_2102 );
not ( \745_b0 , w_2103 );
and ( w_2102 , w_2103 , \696_b0 );
or ( \746_b1 , \745_b1 , w_2105 );
not ( w_2105 , w_2106 );
and ( \746_b0 , \745_b0 , w_2107 );
and ( w_2106 ,  , w_2107 );
buf ( w_2105 , \698_b1 );
not ( w_2105 , w_2108 );
not (  , w_2109 );
and ( w_2108 , w_2109 , \698_b0 );
buf ( \747_b1 , \746_b1 );
not ( \747_b1 , w_2110 );
not ( \747_b0 , w_2111 );
and ( w_2110 , w_2111 , \746_b0 );
or ( \748_b1 , \744_b1 , w_2112 );
or ( \748_b0 , \744_b0 , \747_b0 );
not ( \747_b0 , w_2113 );
and ( w_2113 , w_2112 , \747_b1 );
or ( \749_b1 , \b[5]_b1 , \c[3]_b1 );
xor ( \749_b0 , \b[5]_b0 , w_2114 );
not ( w_2114 , w_2115 );
and ( w_2115 , \c[3]_b1 , \c[3]_b0 );
or ( \750_b1 , \702_b1 , w_2117 );
not ( w_2117 , w_2118 );
and ( \750_b0 , \702_b0 , w_2119 );
and ( w_2118 ,  , w_2119 );
buf ( w_2117 , \749_b1 );
not ( w_2117 , w_2120 );
not (  , w_2121 );
and ( w_2120 , w_2121 , \749_b0 );
or ( \751_b1 , \748_b1 , w_2123 );
not ( w_2123 , w_2124 );
and ( \751_b0 , \748_b0 , w_2125 );
and ( w_2124 ,  , w_2125 );
buf ( w_2123 , \750_b1 );
not ( w_2123 , w_2126 );
not (  , w_2127 );
and ( w_2126 , w_2127 , \750_b0 );
or ( \752_b1 , \743_b1 , \751_b1 );
xor ( \752_b0 , \743_b0 , w_2128 );
not ( w_2128 , w_2129 );
and ( w_2129 , \751_b1 , \751_b0 );
or ( \753_b1 , \722_b1 , w_2130 );
xor ( \753_b0 , \722_b0 , w_2132 );
not ( w_2132 , w_2133 );
and ( w_2133 , w_2130 , w_2131 );
buf ( w_2130 , \752_b1 );
not ( w_2130 , w_2134 );
not ( w_2131 , w_2135 );
and ( w_2134 , w_2135 , \752_b0 );
or ( \754_b1 , \b[4]_b1 , \c[1]_b1 );
xor ( \754_b0 , \b[4]_b0 , w_2136 );
not ( w_2136 , w_2137 );
and ( w_2137 , \c[1]_b1 , \c[1]_b0 );
buf ( \755_b1 , \754_b1 );
not ( \755_b1 , w_2138 );
not ( \755_b0 , w_2139 );
and ( w_2138 , w_2139 , \754_b0 );
buf ( \756_b1 , \679_b1 );
not ( \756_b1 , w_2140 );
not ( \756_b0 , w_2141 );
and ( w_2140 , w_2141 , \679_b0 );
or ( \757_b1 , \755_b1 , w_2142 );
or ( \757_b0 , \755_b0 , \756_b0 );
not ( \756_b0 , w_2143 );
and ( w_2143 , w_2142 , \756_b1 );
or ( \758_b1 , \707_b1 , w_2145 );
not ( w_2145 , w_2146 );
and ( \758_b0 , \707_b0 , w_2147 );
and ( w_2146 ,  , w_2147 );
buf ( w_2145 , \c[0]_b1 );
not ( w_2145 , w_2148 );
not (  , w_2149 );
and ( w_2148 , w_2149 , \c[0]_b0 );
or ( \759_b1 , \757_b1 , w_2151 );
not ( w_2151 , w_2152 );
and ( \759_b0 , \757_b0 , w_2153 );
and ( w_2152 ,  , w_2153 );
buf ( w_2151 , \758_b1 );
not ( w_2151 , w_2154 );
not (  , w_2155 );
and ( w_2154 , w_2155 , \758_b0 );
buf ( \760_b1 , \759_b1 );
not ( \760_b1 , w_2156 );
not ( \760_b0 , w_2157 );
and ( w_2156 , w_2157 , \759_b0 );
or ( \761_b1 , \b[0]_b1 , w_2158 );
or ( \761_b0 , \b[0]_b0 , \c[4]_b0 );
not ( \c[4]_b0 , w_2159 );
and ( w_2159 , w_2158 , \c[4]_b1 );
or ( \762_b1 , \761_b1 , w_2161 );
not ( w_2161 , w_2162 );
and ( \762_b0 , \761_b0 , w_2163 );
and ( w_2162 ,  , w_2163 );
buf ( w_2161 , \c[3]_b1 );
not ( w_2161 , w_2164 );
not (  , w_2165 );
and ( w_2164 , w_2165 , \c[3]_b0 );
or ( \763_b1 , \b[0]_b1 , w_2167 );
not ( w_2167 , w_2168 );
and ( \763_b0 , \b[0]_b0 , w_2169 );
and ( w_2168 ,  , w_2169 );
buf ( w_2167 , \c[4]_b1 );
not ( w_2167 , w_2170 );
not (  , w_2171 );
and ( w_2170 , w_2171 , \c[4]_b0 );
or ( \765_b1 , \760_b1 , w_2173 );
not ( w_2173 , w_2174 );
and ( \765_b0 , \760_b0 , w_2175 );
and ( w_2174 ,  , w_2175 );
buf ( w_2173 , \764_b1 );
not ( w_2173 , w_2176 );
not (  , w_2177 );
and ( w_2176 , w_2177 , \764_b0 );
buf ( \766_b1 , \765_b1 );
not ( \766_b1 , w_2178 );
not ( \766_b0 , w_2179 );
and ( w_2178 , w_2179 , \765_b0 );
or ( \767_b1 , \b[1]_b1 , \c[5]_b1 );
xor ( \767_b0 , \b[1]_b0 , w_2180 );
not ( w_2180 , w_2181 );
and ( w_2181 , \c[5]_b1 , \c[5]_b0 );
buf ( \768_b1 , \767_b1 );
not ( \768_b1 , w_2182 );
not ( \768_b0 , w_2183 );
and ( w_2182 , w_2183 , \767_b0 );
buf ( \769_b1 , \736_b1 );
not ( \769_b1 , w_2184 );
not ( \769_b0 , w_2185 );
and ( w_2184 , w_2185 , \736_b0 );
or ( \770_b1 , \768_b1 , w_2186 );
or ( \770_b0 , \768_b0 , \769_b0 );
not ( \769_b0 , w_2187 );
and ( w_2187 , w_2186 , \769_b1 );
or ( \771_b1 , \734_b1 , w_2189 );
not ( w_2189 , w_2190 );
and ( \771_b0 , \734_b0 , w_2191 );
and ( w_2190 ,  , w_2191 );
buf ( w_2189 , \732_b1 );
not ( w_2189 , w_2192 );
not (  , w_2193 );
and ( w_2192 , w_2193 , \732_b0 );
or ( \772_b1 , \770_b1 , w_2195 );
not ( w_2195 , w_2196 );
and ( \772_b0 , \770_b0 , w_2197 );
and ( w_2196 ,  , w_2197 );
buf ( w_2195 , \771_b1 );
not ( w_2195 , w_2198 );
not (  , w_2199 );
and ( w_2198 , w_2199 , \771_b0 );
buf ( \773_b1 , \772_b1 );
not ( \773_b1 , w_2200 );
not ( \773_b0 , w_2201 );
and ( w_2200 , w_2201 , \772_b0 );
or ( \774_b1 , \766_b1 , w_2203 );
not ( w_2203 , w_2204 );
and ( \774_b0 , \766_b0 , w_2205 );
and ( w_2204 ,  , w_2205 );
buf ( w_2203 , \773_b1 );
not ( w_2203 , w_2206 );
not (  , w_2207 );
and ( w_2206 , w_2207 , \773_b0 );
buf ( \775_b1 , \774_b1 );
not ( \775_b1 , w_2208 );
not ( \775_b0 , w_2209 );
and ( w_2208 , w_2209 , \774_b0 );
or ( \776_b1 , \715_b1 , \712_b1 );
xor ( \776_b0 , \715_b0 , w_2210 );
not ( w_2210 , w_2211 );
and ( w_2211 , \712_b1 , \712_b0 );
or ( \777_b1 , \776_b1 , w_2212 );
xor ( \777_b0 , \776_b0 , w_2214 );
not ( w_2214 , w_2215 );
and ( w_2215 , w_2212 , w_2213 );
buf ( w_2212 , \705_b1 );
not ( w_2212 , w_2216 );
not ( w_2213 , w_2217 );
and ( w_2216 , w_2217 , \705_b0 );
buf ( \778_b1 , \777_b1 );
not ( \778_b1 , w_2218 );
not ( \778_b0 , w_2219 );
and ( w_2218 , w_2219 , \777_b0 );
or ( \779_b1 , \775_b1 , w_2220 );
or ( \779_b0 , \775_b0 , \778_b0 );
not ( \778_b0 , w_2221 );
and ( w_2221 , w_2220 , \778_b1 );
or ( \780_b1 , \772_b1 , w_2223 );
not ( w_2223 , w_2224 );
and ( \780_b0 , \772_b0 , w_2225 );
and ( w_2224 ,  , w_2225 );
buf ( w_2223 , \765_b1 );
not ( w_2223 , w_2226 );
not (  , w_2227 );
and ( w_2226 , w_2227 , \765_b0 );
or ( \781_b1 , \779_b1 , w_2229 );
not ( w_2229 , w_2230 );
and ( \781_b0 , \779_b0 , w_2231 );
and ( w_2230 ,  , w_2231 );
buf ( w_2229 , \780_b1 );
not ( w_2229 , w_2232 );
not (  , w_2233 );
and ( w_2232 , w_2233 , \780_b0 );
or ( \782_b1 , \753_b1 , w_2234 );
or ( \782_b0 , \753_b0 , \781_b0 );
not ( \781_b0 , w_2235 );
and ( w_2235 , w_2234 , \781_b1 );
or ( \783_b1 , \753_b1 , w_2237 );
not ( w_2237 , w_2238 );
and ( \783_b0 , \753_b0 , w_2239 );
and ( w_2238 ,  , w_2239 );
buf ( w_2237 , \781_b1 );
not ( w_2237 , w_2240 );
not (  , w_2241 );
and ( w_2240 , w_2241 , \781_b0 );
or ( \784_b1 , \782_b1 , w_2243 );
not ( w_2243 , w_2244 );
and ( \784_b0 , \782_b0 , w_2245 );
and ( w_2244 ,  , w_2245 );
buf ( w_2243 , \783_b1 );
not ( w_2243 , w_2246 );
not (  , w_2247 );
and ( w_2246 , w_2247 , \783_b0 );
or ( \785_b1 , \b[0]_b1 , \c[5]_b1 );
xor ( \785_b0 , \b[0]_b0 , w_2248 );
not ( w_2248 , w_2249 );
and ( w_2249 , \c[5]_b1 , \c[5]_b0 );
buf ( \786_b1 , \785_b1 );
not ( \786_b1 , w_2250 );
not ( \786_b0 , w_2251 );
and ( w_2250 , w_2251 , \785_b0 );
buf ( \787_b1 , \736_b1 );
not ( \787_b1 , w_2252 );
not ( \787_b0 , w_2253 );
and ( w_2252 , w_2253 , \736_b0 );
or ( \788_b1 , \786_b1 , w_2254 );
or ( \788_b0 , \786_b0 , \787_b0 );
not ( \787_b0 , w_2255 );
and ( w_2255 , w_2254 , \787_b1 );
or ( \789_b1 , \739_b1 , w_2257 );
not ( w_2257 , w_2258 );
and ( \789_b0 , \739_b0 , w_2259 );
and ( w_2258 ,  , w_2259 );
buf ( w_2257 , \767_b1 );
not ( w_2257 , w_2260 );
not (  , w_2261 );
and ( w_2260 , w_2261 , \767_b0 );
or ( \790_b1 , \788_b1 , w_2263 );
not ( w_2263 , w_2264 );
and ( \790_b0 , \788_b0 , w_2265 );
and ( w_2264 ,  , w_2265 );
buf ( w_2263 , \789_b1 );
not ( w_2263 , w_2266 );
not (  , w_2267 );
and ( w_2266 , w_2267 , \789_b0 );
buf ( \791_b1 , \759_b1 );
not ( \791_b1 , w_2268 );
not ( \791_b0 , w_2269 );
and ( w_2268 , w_2269 , \759_b0 );
buf ( \792_b1 , \764_b1 );
not ( \792_b1 , w_2270 );
not ( \792_b0 , w_2271 );
and ( w_2270 , w_2271 , \764_b0 );
or ( \793_b1 , \791_b1 , \792_b1 );
not ( \792_b1 , w_2272 );
and ( \793_b0 , \791_b0 , w_2273 );
and ( w_2272 , w_2273 , \792_b0 );
or ( \794_b1 , \759_b1 , \764_b1 );
not ( \764_b1 , w_2274 );
and ( \794_b0 , \759_b0 , w_2275 );
and ( w_2274 , w_2275 , \764_b0 );
or ( \795_b1 , \793_b1 , w_2277 );
not ( w_2277 , w_2278 );
and ( \795_b0 , \793_b0 , w_2279 );
and ( w_2278 ,  , w_2279 );
buf ( w_2277 , \794_b1 );
not ( w_2277 , w_2280 );
not (  , w_2281 );
and ( w_2280 , w_2281 , \794_b0 );
or ( \796_b1 , \790_b1 , \795_b1 );
xor ( \796_b0 , \790_b0 , w_2282 );
not ( w_2282 , w_2283 );
and ( w_2283 , \795_b1 , \795_b0 );
or ( \797_b1 , \b[2]_b1 , \c[3]_b1 );
xor ( \797_b0 , \b[2]_b0 , w_2284 );
not ( w_2284 , w_2285 );
and ( w_2285 , \c[3]_b1 , \c[3]_b0 );
buf ( \798_b1 , \797_b1 );
not ( \798_b1 , w_2286 );
not ( \798_b0 , w_2287 );
and ( w_2286 , w_2287 , \797_b0 );
buf ( \799_b1 , \746_b1 );
not ( \799_b1 , w_2288 );
not ( \799_b0 , w_2289 );
and ( w_2288 , w_2289 , \746_b0 );
or ( \800_b1 , \798_b1 , w_2290 );
or ( \800_b0 , \798_b0 , \799_b0 );
not ( \799_b0 , w_2291 );
and ( w_2291 , w_2290 , \799_b1 );
or ( \801_b1 , \702_b1 , w_2293 );
not ( w_2293 , w_2294 );
and ( \801_b0 , \702_b0 , w_2295 );
and ( w_2294 ,  , w_2295 );
buf ( w_2293 , \694_b1 );
not ( w_2293 , w_2296 );
not (  , w_2297 );
and ( w_2296 , w_2297 , \694_b0 );
or ( \802_b1 , \800_b1 , w_2299 );
not ( w_2299 , w_2300 );
and ( \802_b0 , \800_b0 , w_2301 );
and ( w_2300 ,  , w_2301 );
buf ( w_2299 , \801_b1 );
not ( w_2299 , w_2302 );
not (  , w_2303 );
and ( w_2302 , w_2303 , \801_b0 );
or ( \803_b1 , \796_b1 , \802_b1 );
xor ( \803_b0 , \796_b0 , w_2304 );
not ( w_2304 , w_2305 );
and ( w_2305 , \802_b1 , \802_b0 );
or ( \804_b1 , \739_b1 , w_2307 );
not ( w_2307 , w_2308 );
and ( \804_b0 , \739_b0 , w_2309 );
and ( w_2308 ,  , w_2309 );
buf ( w_2307 , \b[0]_b1 );
not ( w_2307 , w_2310 );
not (  , w_2311 );
and ( w_2310 , w_2311 , \b[0]_b0 );
or ( \805_b1 , \702_b1 , \797_b1 );
not ( \797_b1 , w_2312 );
and ( \805_b0 , \702_b0 , w_2313 );
and ( w_2312 , w_2313 , \797_b0 );
buf ( \806_b1 , \702_b1 );
not ( \806_b1 , w_2314 );
not ( \806_b0 , w_2315 );
and ( w_2314 , w_2315 , \702_b0 );
or ( \807_b1 , \b[1]_b1 , \c[3]_b1 );
xor ( \807_b0 , \b[1]_b0 , w_2316 );
not ( w_2316 , w_2317 );
and ( w_2317 , \c[3]_b1 , \c[3]_b0 );
or ( \808_b1 , \696_b1 , \807_b1 );
not ( \807_b1 , w_2318 );
and ( \808_b0 , \696_b0 , w_2319 );
and ( w_2318 , w_2319 , \807_b0 );
or ( \809_b1 , \806_b1 , \808_b1 );
not ( \808_b1 , w_2320 );
and ( \809_b0 , \806_b0 , w_2321 );
and ( w_2320 , w_2321 , \808_b0 );
or ( \810_b1 , \805_b1 , w_2323 );
not ( w_2323 , w_2324 );
and ( \810_b0 , \805_b0 , w_2325 );
and ( w_2324 ,  , w_2325 );
buf ( w_2323 , \809_b1 );
not ( w_2323 , w_2326 );
not (  , w_2327 );
and ( w_2326 , w_2327 , \809_b0 );
or ( \811_b1 , \804_b1 , \810_b1 );
xor ( \811_b0 , \804_b0 , w_2328 );
not ( w_2328 , w_2329 );
and ( w_2329 , \810_b1 , \810_b0 );
or ( \812_b1 , \b[3]_b1 , \c[1]_b1 );
xor ( \812_b0 , \b[3]_b0 , w_2330 );
not ( w_2330 , w_2331 );
and ( w_2331 , \c[1]_b1 , \c[1]_b0 );
or ( \813_b1 , \679_b1 , \812_b1 );
not ( \812_b1 , w_2332 );
and ( \813_b0 , \679_b0 , w_2333 );
and ( w_2332 , w_2333 , \812_b0 );
or ( \814_b1 , \754_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_2334 );
and ( \814_b0 , \754_b0 , w_2335 );
and ( w_2334 , w_2335 , \c[0]_b0 );
or ( \815_b1 , \813_b1 , w_2337 );
not ( w_2337 , w_2338 );
and ( \815_b0 , \813_b0 , w_2339 );
and ( w_2338 ,  , w_2339 );
buf ( w_2337 , \814_b1 );
not ( w_2337 , w_2340 );
not (  , w_2341 );
and ( w_2340 , w_2341 , \814_b0 );
or ( \816_b1 , \811_b1 , \815_b1 );
not ( \815_b1 , w_2342 );
and ( \816_b0 , \811_b0 , w_2343 );
and ( w_2342 , w_2343 , \815_b0 );
or ( \817_b1 , \804_b1 , \810_b1 );
not ( \810_b1 , w_2344 );
and ( \817_b0 , \804_b0 , w_2345 );
and ( w_2344 , w_2345 , \810_b0 );
or ( \818_b1 , \816_b1 , w_2346 );
or ( \818_b0 , \816_b0 , \817_b0 );
not ( \817_b0 , w_2347 );
and ( w_2347 , w_2346 , \817_b1 );
or ( \819_b1 , \803_b1 , w_2349 );
not ( w_2349 , w_2350 );
and ( \819_b0 , \803_b0 , w_2351 );
and ( w_2350 ,  , w_2351 );
buf ( w_2349 , \818_b1 );
not ( w_2349 , w_2352 );
not (  , w_2353 );
and ( w_2352 , w_2353 , \818_b0 );
or ( \820_b1 , \b[0]_b1 , \c[3]_b1 );
xor ( \820_b0 , \b[0]_b0 , w_2354 );
not ( w_2354 , w_2355 );
and ( w_2355 , \c[3]_b1 , \c[3]_b0 );
buf ( \821_b1 , \820_b1 );
not ( \821_b1 , w_2356 );
not ( \821_b0 , w_2357 );
and ( w_2356 , w_2357 , \820_b0 );
buf ( \822_b1 , \746_b1 );
not ( \822_b1 , w_2358 );
not ( \822_b0 , w_2359 );
and ( w_2358 , w_2359 , \746_b0 );
or ( \823_b1 , \821_b1 , w_2360 );
or ( \823_b0 , \821_b0 , \822_b0 );
not ( \822_b0 , w_2361 );
and ( w_2361 , w_2360 , \822_b1 );
or ( \824_b1 , \702_b1 , w_2363 );
not ( w_2363 , w_2364 );
and ( \824_b0 , \702_b0 , w_2365 );
and ( w_2364 ,  , w_2365 );
buf ( w_2363 , \807_b1 );
not ( w_2363 , w_2366 );
not (  , w_2367 );
and ( w_2366 , w_2367 , \807_b0 );
or ( \825_b1 , \823_b1 , w_2369 );
not ( w_2369 , w_2370 );
and ( \825_b0 , \823_b0 , w_2371 );
and ( w_2370 ,  , w_2371 );
buf ( w_2369 , \824_b1 );
not ( w_2369 , w_2372 );
not (  , w_2373 );
and ( w_2372 , w_2373 , \824_b0 );
buf ( \826_b1 , \825_b1 );
not ( \826_b1 , w_2374 );
not ( \826_b0 , w_2375 );
and ( w_2374 , w_2375 , \825_b0 );
or ( \827_b1 , \b[2]_b1 , \c[1]_b1 );
xor ( \827_b0 , \b[2]_b0 , w_2376 );
not ( w_2376 , w_2377 );
and ( w_2377 , \c[1]_b1 , \c[1]_b0 );
buf ( \828_b1 , \827_b1 );
not ( \828_b1 , w_2378 );
not ( \828_b0 , w_2379 );
and ( w_2378 , w_2379 , \827_b0 );
buf ( \829_b1 , \679_b1 );
not ( \829_b1 , w_2380 );
not ( \829_b0 , w_2381 );
and ( w_2380 , w_2381 , \679_b0 );
or ( \830_b1 , \828_b1 , w_2382 );
or ( \830_b0 , \828_b0 , \829_b0 );
not ( \829_b0 , w_2383 );
and ( w_2383 , w_2382 , \829_b1 );
or ( \831_b1 , \812_b1 , w_2385 );
not ( w_2385 , w_2386 );
and ( \831_b0 , \812_b0 , w_2387 );
and ( w_2386 ,  , w_2387 );
buf ( w_2385 , \c[0]_b1 );
not ( w_2385 , w_2388 );
not (  , w_2389 );
and ( w_2388 , w_2389 , \c[0]_b0 );
or ( \832_b1 , \830_b1 , w_2391 );
not ( w_2391 , w_2392 );
and ( \832_b0 , \830_b0 , w_2393 );
and ( w_2392 ,  , w_2393 );
buf ( w_2391 , \831_b1 );
not ( w_2391 , w_2394 );
not (  , w_2395 );
and ( w_2394 , w_2395 , \831_b0 );
buf ( \833_b1 , \832_b1 );
not ( \833_b1 , w_2396 );
not ( \833_b0 , w_2397 );
and ( w_2396 , w_2397 , \832_b0 );
or ( \834_b1 , \b[0]_b1 , w_2399 );
not ( w_2399 , w_2400 );
and ( \834_b0 , \b[0]_b0 , w_2401 );
and ( w_2400 ,  , w_2401 );
buf ( w_2399 , \c[2]_b1 );
not ( w_2399 , w_2402 );
not (  , w_2403 );
and ( w_2402 , w_2403 , \c[2]_b0 );
or ( \835_b1 , \b[0]_b1 , w_2404 );
or ( \835_b0 , \b[0]_b0 , \c[2]_b0 );
not ( \c[2]_b0 , w_2405 );
and ( w_2405 , w_2404 , \c[2]_b1 );
or ( \836_b1 , \835_b1 , w_2407 );
not ( w_2407 , w_2408 );
and ( \836_b0 , \835_b0 , w_2409 );
and ( w_2408 ,  , w_2409 );
buf ( w_2407 , \c[1]_b1 );
not ( w_2407 , w_2410 );
not (  , w_2411 );
and ( w_2410 , w_2411 , \c[1]_b0 );
buf ( \838_b1 , \837_b1 );
not ( \838_b1 , w_2412 );
not ( \838_b0 , w_2413 );
and ( w_2412 , w_2413 , \837_b0 );
or ( \839_b1 , \833_b1 , \838_b1 );
not ( \838_b1 , w_2414 );
and ( \839_b0 , \833_b0 , w_2415 );
and ( w_2414 , w_2415 , \838_b0 );
or ( \840_b1 , \832_b1 , \837_b1 );
not ( \837_b1 , w_2416 );
and ( \840_b0 , \832_b0 , w_2417 );
and ( w_2416 , w_2417 , \837_b0 );
or ( \841_b1 , \839_b1 , w_2419 );
not ( w_2419 , w_2420 );
and ( \841_b0 , \839_b0 , w_2421 );
and ( w_2420 ,  , w_2421 );
buf ( w_2419 , \840_b1 );
not ( w_2419 , w_2422 );
not (  , w_2423 );
and ( w_2422 , w_2423 , \840_b0 );
or ( \842_b1 , \826_b1 , w_2425 );
not ( w_2425 , w_2426 );
and ( \842_b0 , \826_b0 , w_2427 );
and ( w_2426 ,  , w_2427 );
buf ( w_2425 , \841_b1 );
not ( w_2425 , w_2428 );
not (  , w_2429 );
and ( w_2428 , w_2429 , \841_b0 );
buf ( \843_b1 , \842_b1 );
not ( \843_b1 , w_2430 );
not ( \843_b0 , w_2431 );
and ( w_2430 , w_2431 , \842_b0 );
or ( \844_b1 , \c[1]_b1 , \b[1]_b1 );
xor ( \844_b0 , \c[1]_b0 , w_2432 );
not ( w_2432 , w_2433 );
and ( w_2433 , \b[1]_b1 , \b[1]_b0 );
buf ( \845_b1 , \844_b1 );
not ( \845_b1 , w_2434 );
not ( \845_b0 , w_2435 );
and ( w_2434 , w_2435 , \844_b0 );
buf ( \846_b1 , \679_b1 );
not ( \846_b1 , w_2436 );
not ( \846_b0 , w_2437 );
and ( w_2436 , w_2437 , \679_b0 );
or ( \847_b1 , \845_b1 , w_2438 );
or ( \847_b0 , \845_b0 , \846_b0 );
not ( \846_b0 , w_2439 );
and ( w_2439 , w_2438 , \846_b1 );
or ( \848_b1 , \827_b1 , w_2441 );
not ( w_2441 , w_2442 );
and ( \848_b0 , \827_b0 , w_2443 );
and ( w_2442 ,  , w_2443 );
buf ( w_2441 , \c[0]_b1 );
not ( w_2441 , w_2444 );
not (  , w_2445 );
and ( w_2444 , w_2445 , \c[0]_b0 );
or ( \849_b1 , \847_b1 , w_2447 );
not ( w_2447 , w_2448 );
and ( \849_b0 , \847_b0 , w_2449 );
and ( w_2448 ,  , w_2449 );
buf ( w_2447 , \848_b1 );
not ( w_2447 , w_2450 );
not (  , w_2451 );
and ( w_2450 , w_2451 , \848_b0 );
or ( \850_b1 , \702_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_2452 );
and ( \850_b0 , \702_b0 , w_2453 );
and ( w_2452 , w_2453 , \b[0]_b0 );
or ( \851_b1 , \849_b1 , w_2455 );
not ( w_2455 , w_2456 );
and ( \851_b0 , \849_b0 , w_2457 );
and ( w_2456 ,  , w_2457 );
buf ( w_2455 , \850_b1 );
not ( w_2455 , w_2458 );
not (  , w_2459 );
and ( w_2458 , w_2459 , \850_b0 );
or ( \852_b1 , \b[0]_b1 , w_2461 );
not ( w_2461 , w_2462 );
and ( \852_b0 , \b[0]_b0 , w_2463 );
and ( w_2462 ,  , w_2463 );
buf ( w_2461 , \c[0]_b1 );
not ( w_2461 , w_2464 );
not (  , w_2465 );
and ( w_2464 , w_2465 , \c[0]_b0 );
or ( \853_b1 , \852_b1 , w_2467 );
not ( w_2467 , w_2468 );
and ( \853_b0 , \852_b0 , w_2469 );
and ( w_2468 ,  , w_2469 );
buf ( w_2467 , \c[1]_b1 );
not ( w_2467 , w_2470 );
not (  , w_2471 );
and ( w_2470 , w_2471 , \c[1]_b0 );
buf ( \854_b1 , \853_b1 );
not ( \854_b1 , w_2472 );
not ( \854_b0 , w_2473 );
and ( w_2472 , w_2473 , \853_b0 );
or ( \855_b1 , \b[0]_b1 , \c[1]_b1 );
xor ( \855_b0 , \b[0]_b0 , w_2474 );
not ( w_2474 , w_2475 );
and ( w_2475 , \c[1]_b1 , \c[1]_b0 );
buf ( \856_b1 , \855_b1 );
not ( \856_b1 , w_2476 );
not ( \856_b0 , w_2477 );
and ( w_2476 , w_2477 , \855_b0 );
buf ( \857_b1 , \679_b1 );
not ( \857_b1 , w_2478 );
not ( \857_b0 , w_2479 );
and ( w_2478 , w_2479 , \679_b0 );
or ( \858_b1 , \856_b1 , w_2480 );
or ( \858_b0 , \856_b0 , \857_b0 );
not ( \857_b0 , w_2481 );
and ( w_2481 , w_2480 , \857_b1 );
or ( \859_b1 , \844_b1 , w_2483 );
not ( w_2483 , w_2484 );
and ( \859_b0 , \844_b0 , w_2485 );
and ( w_2484 ,  , w_2485 );
buf ( w_2483 , \c[0]_b1 );
not ( w_2483 , w_2486 );
not (  , w_2487 );
and ( w_2486 , w_2487 , \c[0]_b0 );
or ( \860_b1 , \858_b1 , w_2489 );
not ( w_2489 , w_2490 );
and ( \860_b0 , \858_b0 , w_2491 );
and ( w_2490 ,  , w_2491 );
buf ( w_2489 , \859_b1 );
not ( w_2489 , w_2492 );
not (  , w_2493 );
and ( w_2492 , w_2493 , \859_b0 );
or ( \861_b1 , \854_b1 , w_2495 );
not ( w_2495 , w_2496 );
and ( \861_b0 , \854_b0 , w_2497 );
and ( w_2496 ,  , w_2497 );
buf ( w_2495 , \860_b1 );
not ( w_2495 , w_2498 );
not (  , w_2499 );
and ( w_2498 , w_2499 , \860_b0 );
or ( \862_b1 , \851_b1 , w_2500 );
or ( \862_b0 , \851_b0 , \861_b0 );
not ( \861_b0 , w_2501 );
and ( w_2501 , w_2500 , \861_b1 );
or ( \863_b1 , \849_b1 , w_2503 );
not ( w_2503 , w_2504 );
and ( \863_b0 , \849_b0 , w_2505 );
and ( w_2504 ,  , w_2505 );
buf ( w_2503 , \850_b1 );
not ( w_2503 , w_2506 );
not (  , w_2507 );
and ( w_2506 , w_2507 , \850_b0 );
or ( \864_b1 , \862_b1 , w_2509 );
not ( w_2509 , w_2510 );
and ( \864_b0 , \862_b0 , w_2511 );
and ( w_2510 ,  , w_2511 );
buf ( w_2509 , \863_b1 );
not ( w_2509 , w_2512 );
not (  , w_2513 );
and ( w_2512 , w_2513 , \863_b0 );
buf ( \865_b1 , \864_b1 );
not ( \865_b1 , w_2514 );
not ( \865_b0 , w_2515 );
and ( w_2514 , w_2515 , \864_b0 );
or ( \866_b1 , \843_b1 , w_2516 );
or ( \866_b0 , \843_b0 , \865_b0 );
not ( \865_b0 , w_2517 );
and ( w_2517 , w_2516 , \865_b1 );
buf ( \867_b1 , \841_b1 );
not ( \867_b1 , w_2518 );
not ( \867_b0 , w_2519 );
and ( w_2518 , w_2519 , \841_b0 );
or ( \868_b1 , \867_b1 , w_2521 );
not ( w_2521 , w_2522 );
and ( \868_b0 , \867_b0 , w_2523 );
and ( w_2522 ,  , w_2523 );
buf ( w_2521 , \825_b1 );
not ( w_2521 , w_2524 );
not (  , w_2525 );
and ( w_2524 , w_2525 , \825_b0 );
or ( \869_b1 , \866_b1 , w_2527 );
not ( w_2527 , w_2528 );
and ( \869_b0 , \866_b0 , w_2529 );
and ( w_2528 ,  , w_2529 );
buf ( w_2527 , \868_b1 );
not ( w_2527 , w_2530 );
not (  , w_2531 );
and ( w_2530 , w_2531 , \868_b0 );
buf ( \870_b1 , \869_b1 );
not ( \870_b1 , w_2532 );
not ( \870_b0 , w_2533 );
and ( w_2532 , w_2533 , \869_b0 );
or ( \871_b1 , \804_b1 , \810_b1 );
xor ( \871_b0 , \804_b0 , w_2534 );
not ( w_2534 , w_2535 );
and ( w_2535 , \810_b1 , \810_b0 );
or ( \872_b1 , \871_b1 , \815_b1 );
xor ( \872_b0 , \871_b0 , w_2536 );
not ( w_2536 , w_2537 );
and ( w_2537 , \815_b1 , \815_b0 );
buf ( \873_b1 , \837_b1 );
not ( \873_b1 , w_2538 );
not ( \873_b0 , w_2539 );
and ( w_2538 , w_2539 , \837_b0 );
or ( \874_b1 , \873_b1 , w_2541 );
not ( w_2541 , w_2542 );
and ( \874_b0 , \873_b0 , w_2543 );
and ( w_2542 ,  , w_2543 );
buf ( w_2541 , \832_b1 );
not ( w_2541 , w_2544 );
not (  , w_2545 );
and ( w_2544 , w_2545 , \832_b0 );
or ( \875_b1 , \872_b1 , w_2547 );
not ( w_2547 , w_2548 );
and ( \875_b0 , \872_b0 , w_2549 );
and ( w_2548 ,  , w_2549 );
buf ( w_2547 , \874_b1 );
not ( w_2547 , w_2550 );
not (  , w_2551 );
and ( w_2550 , w_2551 , \874_b0 );
buf ( \876_b1 , \875_b1 );
not ( \876_b1 , w_2552 );
not ( \876_b0 , w_2553 );
and ( w_2552 , w_2553 , \875_b0 );
or ( \877_b1 , \870_b1 , w_2554 );
or ( \877_b0 , \870_b0 , \876_b0 );
not ( \876_b0 , w_2555 );
and ( w_2555 , w_2554 , \876_b1 );
or ( \878_b1 , \872_b1 , w_2556 );
or ( \878_b0 , \872_b0 , \874_b0 );
not ( \874_b0 , w_2557 );
and ( w_2557 , w_2556 , \874_b1 );
or ( \879_b1 , \877_b1 , w_2559 );
not ( w_2559 , w_2560 );
and ( \879_b0 , \877_b0 , w_2561 );
and ( w_2560 ,  , w_2561 );
buf ( w_2559 , \878_b1 );
not ( w_2559 , w_2562 );
not (  , w_2563 );
and ( w_2562 , w_2563 , \878_b0 );
or ( \880_b1 , \819_b1 , w_2565 );
not ( w_2565 , w_2566 );
and ( \880_b0 , \819_b0 , w_2567 );
and ( w_2566 ,  , w_2567 );
buf ( w_2565 , \879_b1 );
not ( w_2565 , w_2568 );
not (  , w_2569 );
and ( w_2568 , w_2569 , \879_b0 );
buf ( \881_b1 , \765_b1 );
not ( \881_b1 , w_2570 );
not ( \881_b0 , w_2571 );
and ( w_2570 , w_2571 , \765_b0 );
buf ( \882_b1 , \773_b1 );
not ( \882_b1 , w_2572 );
not ( \882_b0 , w_2573 );
and ( w_2572 , w_2573 , \773_b0 );
or ( \883_b1 , \881_b1 , \882_b1 );
not ( \882_b1 , w_2574 );
and ( \883_b0 , \881_b0 , w_2575 );
and ( w_2574 , w_2575 , \882_b0 );
or ( \884_b1 , \765_b1 , \773_b1 );
not ( \773_b1 , w_2576 );
and ( \884_b0 , \765_b0 , w_2577 );
and ( w_2576 , w_2577 , \773_b0 );
or ( \885_b1 , \883_b1 , w_2579 );
not ( w_2579 , w_2580 );
and ( \885_b0 , \883_b0 , w_2581 );
and ( w_2580 ,  , w_2581 );
buf ( w_2579 , \884_b1 );
not ( w_2579 , w_2582 );
not (  , w_2583 );
and ( w_2582 , w_2583 , \884_b0 );
or ( \886_b1 , \777_b1 , w_2584 );
xor ( \886_b0 , \777_b0 , w_2586 );
not ( w_2586 , w_2587 );
and ( w_2587 , w_2584 , w_2585 );
buf ( w_2584 , \885_b1 );
not ( w_2584 , w_2588 );
not ( w_2585 , w_2589 );
and ( w_2588 , w_2589 , \885_b0 );
buf ( \887_b1 , \795_b1 );
not ( \887_b1 , w_2590 );
not ( \887_b0 , w_2591 );
and ( w_2590 , w_2591 , \795_b0 );
or ( \888_b1 , \887_b1 , w_2593 );
not ( w_2593 , w_2594 );
and ( \888_b0 , \887_b0 , w_2595 );
and ( w_2594 ,  , w_2595 );
buf ( w_2593 , \790_b1 );
not ( w_2593 , w_2596 );
not (  , w_2597 );
and ( w_2596 , w_2597 , \790_b0 );
buf ( \889_b1 , \790_b1 );
not ( \889_b1 , w_2598 );
not ( \889_b0 , w_2599 );
and ( w_2598 , w_2599 , \790_b0 );
buf ( \890_b1 , \889_b1 );
not ( \890_b1 , w_2600 );
not ( \890_b0 , w_2601 );
and ( w_2600 , w_2601 , \889_b0 );
buf ( \891_b1 , \795_b1 );
not ( \891_b1 , w_2602 );
not ( \891_b0 , w_2603 );
and ( w_2602 , w_2603 , \795_b0 );
or ( \892_b1 , \890_b1 , w_2604 );
or ( \892_b0 , \890_b0 , \891_b0 );
not ( \891_b0 , w_2605 );
and ( w_2605 , w_2604 , \891_b1 );
or ( \893_b1 , \892_b1 , w_2607 );
not ( w_2607 , w_2608 );
and ( \893_b0 , \892_b0 , w_2609 );
and ( w_2608 ,  , w_2609 );
buf ( w_2607 , \802_b1 );
not ( w_2607 , w_2610 );
not (  , w_2611 );
and ( w_2610 , w_2611 , \802_b0 );
or ( \894_b1 , \888_b1 , w_2613 );
not ( w_2613 , w_2614 );
and ( \894_b0 , \888_b0 , w_2615 );
and ( w_2614 ,  , w_2615 );
buf ( w_2613 , \893_b1 );
not ( w_2613 , w_2616 );
not (  , w_2617 );
and ( w_2616 , w_2617 , \893_b0 );
or ( \895_b1 , \886_b1 , w_2619 );
not ( w_2619 , w_2620 );
and ( \895_b0 , \886_b0 , w_2621 );
and ( w_2620 ,  , w_2621 );
buf ( w_2619 , \894_b1 );
not ( w_2619 , w_2622 );
not (  , w_2623 );
and ( w_2622 , w_2623 , \894_b0 );
or ( \896_b1 , \880_b1 , w_2625 );
not ( w_2625 , w_2626 );
and ( \896_b0 , \880_b0 , w_2627 );
and ( w_2626 ,  , w_2627 );
buf ( w_2625 , \895_b1 );
not ( w_2625 , w_2628 );
not (  , w_2629 );
and ( w_2628 , w_2629 , \895_b0 );
buf ( \897_b1 , \803_b1 );
not ( \897_b1 , w_2630 );
not ( \897_b0 , w_2631 );
and ( w_2630 , w_2631 , \803_b0 );
buf ( \898_b1 , \818_b1 );
not ( \898_b1 , w_2632 );
not ( \898_b0 , w_2633 );
and ( w_2632 , w_2633 , \818_b0 );
or ( \899_b1 , \897_b1 , w_2635 );
not ( w_2635 , w_2636 );
and ( \899_b0 , \897_b0 , w_2637 );
and ( w_2636 ,  , w_2637 );
buf ( w_2635 , \898_b1 );
not ( w_2635 , w_2638 );
not (  , w_2639 );
and ( w_2638 , w_2639 , \898_b0 );
or ( \900_b1 , \895_b1 , w_2640 );
or ( \900_b0 , \895_b0 , \899_b0 );
not ( \899_b0 , w_2641 );
and ( w_2641 , w_2640 , \899_b1 );
or ( \901_b1 , \886_b1 , w_2643 );
not ( w_2643 , w_2644 );
and ( \901_b0 , \886_b0 , w_2645 );
and ( w_2644 ,  , w_2645 );
buf ( w_2643 , \894_b1 );
not ( w_2643 , w_2646 );
not (  , w_2647 );
and ( w_2646 , w_2647 , \894_b0 );
or ( \902_b1 , \900_b1 , w_2649 );
not ( w_2649 , w_2650 );
and ( \902_b0 , \900_b0 , w_2651 );
and ( w_2650 ,  , w_2651 );
buf ( w_2649 , \901_b1 );
not ( w_2649 , w_2652 );
not (  , w_2653 );
and ( w_2652 , w_2653 , \901_b0 );
or ( \903_b1 , \896_b1 , w_2655 );
not ( w_2655 , w_2656 );
and ( \903_b0 , \896_b0 , w_2657 );
and ( w_2656 ,  , w_2657 );
buf ( w_2655 , \902_b1 );
not ( w_2655 , w_2658 );
not (  , w_2659 );
and ( w_2658 , w_2659 , \902_b0 );
buf ( \904_b1 , \903_b1 );
not ( \904_b1 , w_2660 );
not ( \904_b0 , w_2661 );
and ( w_2660 , w_2661 , \903_b0 );
or ( \905_b1 , \784_b1 , \904_b1 );
xor ( \905_b0 , \784_b0 , w_2662 );
not ( w_2662 , w_2663 );
and ( w_2663 , \904_b1 , \904_b0 );
buf ( \906_b1 , \905_b1 );
not ( \906_b1 , w_2664 );
not ( \906_b0 , w_2665 );
and ( w_2664 , w_2665 , \905_b0 );
buf ( \907_b1 , \403_b1 );
not ( \907_b1 , w_2666 );
not ( \907_b0 , w_2667 );
and ( w_2666 , w_2667 , \403_b0 );
buf ( \908_b1 , \529_b1 );
not ( \908_b1 , w_2668 );
not ( \908_b0 , w_2669 );
and ( w_2668 , w_2669 , \529_b0 );
or ( \909_b1 , \907_b1 , w_2670 );
or ( \909_b0 , \907_b0 , \908_b0 );
not ( \908_b0 , w_2671 );
and ( w_2671 , w_2670 , \908_b1 );
or ( \910_b1 , \909_b1 , w_2673 );
not ( w_2673 , w_2674 );
and ( \910_b0 , \909_b0 , w_2675 );
and ( w_2674 ,  , w_2675 );
buf ( w_2673 , \531_b1 );
not ( w_2673 , w_2676 );
not (  , w_2677 );
and ( w_2676 , w_2677 , \531_b0 );
buf ( \911_b1 , \425_b1 );
not ( \911_b1 , w_2678 );
not ( \911_b0 , w_2679 );
and ( w_2678 , w_2679 , \425_b0 );
or ( \912_b1 , \911_b1 , w_2681 );
not ( w_2681 , w_2682 );
and ( \912_b0 , \911_b0 , w_2683 );
and ( w_2682 ,  , w_2683 );
buf ( w_2681 , \423_b1 );
not ( w_2681 , w_2684 );
not (  , w_2685 );
and ( w_2684 , w_2685 , \423_b0 );
or ( \913_b1 , \910_b1 , w_2687 );
not ( w_2687 , w_2688 );
and ( \913_b0 , \910_b0 , w_2689 );
and ( w_2688 ,  , w_2689 );
buf ( w_2687 , \912_b1 );
not ( w_2687 , w_2690 );
not (  , w_2691 );
and ( w_2690 , w_2691 , \912_b0 );
buf ( \914_b1 , \913_b1 );
not ( \914_b1 , w_2692 );
not ( \914_b0 , w_2693 );
and ( w_2692 , w_2693 , \913_b0 );
or ( \915_b1 , \910_b1 , w_2695 );
not ( w_2695 , w_2696 );
and ( \915_b0 , \910_b0 , w_2697 );
and ( w_2696 ,  , w_2697 );
buf ( w_2695 , \912_b1 );
not ( w_2695 , w_2698 );
not (  , w_2699 );
and ( w_2698 , w_2699 , \912_b0 );
or ( \916_b1 , \914_b1 , w_2701 );
not ( w_2701 , w_2702 );
and ( \916_b0 , \914_b0 , w_2703 );
and ( w_2702 ,  , w_2703 );
buf ( w_2701 , \915_b1 );
not ( w_2701 , w_2704 );
not (  , w_2705 );
and ( w_2704 , w_2705 , \915_b0 );
buf ( \917_b1 , \916_b1 );
not ( \917_b1 , w_2706 );
not ( \917_b0 , w_2707 );
and ( w_2706 , w_2707 , \916_b0 );
buf ( \918_b1 , \917_b1 );
not ( \918_b1 , w_2708 );
not ( \918_b0 , w_2709 );
and ( w_2708 , w_2709 , \917_b0 );
or ( \919_b1 , \906_b1 , \918_b1 );
not ( \918_b1 , w_2710 );
and ( \919_b0 , \906_b0 , w_2711 );
and ( w_2710 , w_2711 , \918_b0 );
or ( \920_b1 , \c[7]_b1 , \d[7]_b1 );
xor ( \920_b0 , \c[7]_b0 , w_2712 );
not ( w_2712 , w_2713 );
and ( w_2713 , \d[7]_b1 , \d[7]_b0 );
buf ( \921_b1 , \920_b1 );
not ( \921_b1 , w_2714 );
not ( \921_b0 , w_2715 );
and ( w_2714 , w_2715 , \920_b0 );
buf ( \922_b1 , \661_b1 );
not ( \922_b1 , w_2716 );
not ( \922_b0 , w_2717 );
and ( w_2716 , w_2717 , \661_b0 );
or ( \923_b1 , \922_b1 , w_2719 );
not ( w_2719 , w_2720 );
and ( \923_b0 , \922_b0 , w_2721 );
and ( w_2720 ,  , w_2721 );
buf ( w_2719 , \540_b1 );
not ( w_2719 , w_2722 );
not (  , w_2723 );
and ( w_2722 , w_2723 , \540_b0 );
or ( \924_b1 , \923_b1 , \658_b1 );
xor ( \924_b0 , \923_b0 , w_2724 );
not ( w_2724 , w_2725 );
and ( w_2725 , \658_b1 , \658_b0 );
buf ( \925_b1 , \924_b1 );
not ( \925_b1 , w_2726 );
not ( \925_b0 , w_2727 );
and ( w_2726 , w_2727 , \924_b0 );
buf ( \926_b1 , \925_b1 );
not ( \926_b1 , w_2728 );
not ( \926_b0 , w_2729 );
and ( w_2728 , w_2729 , \925_b0 );
or ( \927_b1 , \921_b1 , w_2730 );
or ( \927_b0 , \921_b0 , \926_b0 );
not ( \926_b0 , w_2731 );
and ( w_2731 , w_2730 , \926_b1 );
or ( \928_b1 , \a[4]_b1 , \d[1]_b1 );
xor ( \928_b0 , \a[4]_b0 , w_2732 );
not ( w_2732 , w_2733 );
and ( w_2733 , \d[1]_b1 , \d[1]_b0 );
buf ( \929_b1 , \928_b1 );
not ( \929_b1 , w_2734 );
not ( \929_b0 , w_2735 );
and ( w_2734 , w_2735 , \928_b0 );
buf ( \930_b1 , \d[0]_b1 );
not ( \930_b1 , w_2736 );
not ( \930_b0 , w_2737 );
and ( w_2736 , w_2737 , \d[0]_b0 );
or ( \931_b1 , \930_b1 , w_2739 );
not ( w_2739 , w_2740 );
and ( \931_b0 , \930_b0 , w_2741 );
and ( w_2740 ,  , w_2741 );
buf ( w_2739 , \d[1]_b1 );
not ( w_2739 , w_2742 );
not (  , w_2743 );
and ( w_2742 , w_2743 , \d[1]_b0 );
buf ( \932_b1 , \931_b1 );
not ( \932_b1 , w_2744 );
not ( \932_b0 , w_2745 );
and ( w_2744 , w_2745 , \931_b0 );
buf ( \933_b1 , \932_b1 );
not ( \933_b1 , w_2746 );
not ( \933_b0 , w_2747 );
and ( w_2746 , w_2747 , \932_b0 );
or ( \934_b1 , \929_b1 , w_2748 );
or ( \934_b0 , \929_b0 , \933_b0 );
not ( \933_b0 , w_2749 );
and ( w_2749 , w_2748 , \933_b1 );
or ( \935_b1 , \a[5]_b1 , \d[1]_b1 );
xor ( \935_b0 , \a[5]_b0 , w_2750 );
not ( w_2750 , w_2751 );
and ( w_2751 , \d[1]_b1 , \d[1]_b0 );
or ( \936_b1 , \935_b1 , w_2753 );
not ( w_2753 , w_2754 );
and ( \936_b0 , \935_b0 , w_2755 );
and ( w_2754 ,  , w_2755 );
buf ( w_2753 , \d[0]_b1 );
not ( w_2753 , w_2756 );
not (  , w_2757 );
and ( w_2756 , w_2757 , \d[0]_b0 );
or ( \937_b1 , \934_b1 , w_2759 );
not ( w_2759 , w_2760 );
and ( \937_b0 , \934_b0 , w_2761 );
and ( w_2760 ,  , w_2761 );
buf ( w_2759 , \936_b1 );
not ( w_2759 , w_2762 );
not (  , w_2763 );
and ( w_2762 , w_2763 , \936_b0 );
buf ( \938_b1 , \937_b1 );
not ( \938_b1 , w_2764 );
not ( \938_b0 , w_2765 );
and ( w_2764 , w_2765 , \937_b0 );
or ( \939_b1 , \a[0]_b1 , w_2766 );
or ( \939_b0 , \a[0]_b0 , \d[4]_b0 );
not ( \d[4]_b0 , w_2767 );
and ( w_2767 , w_2766 , \d[4]_b1 );
or ( \940_b1 , \939_b1 , w_2769 );
not ( w_2769 , w_2770 );
and ( \940_b0 , \939_b0 , w_2771 );
and ( w_2770 ,  , w_2771 );
buf ( w_2769 , \d[3]_b1 );
not ( w_2769 , w_2772 );
not (  , w_2773 );
and ( w_2772 , w_2773 , \d[3]_b0 );
or ( \941_b1 , \a[0]_b1 , w_2775 );
not ( w_2775 , w_2776 );
and ( \941_b0 , \a[0]_b0 , w_2777 );
and ( w_2776 ,  , w_2777 );
buf ( w_2775 , \d[4]_b1 );
not ( w_2775 , w_2778 );
not (  , w_2779 );
and ( w_2778 , w_2779 , \d[4]_b0 );
or ( \943_b1 , \938_b1 , w_2781 );
not ( w_2781 , w_2782 );
and ( \943_b0 , \938_b0 , w_2783 );
and ( w_2782 ,  , w_2783 );
buf ( w_2781 , \942_b1 );
not ( w_2781 , w_2784 );
not (  , w_2785 );
and ( w_2784 , w_2785 , \942_b0 );
or ( \944_b1 , \a[1]_b1 , \d[5]_b1 );
xor ( \944_b0 , \a[1]_b0 , w_2786 );
not ( w_2786 , w_2787 );
and ( w_2787 , \d[5]_b1 , \d[5]_b0 );
buf ( \945_b1 , \944_b1 );
not ( \945_b1 , w_2788 );
not ( \945_b0 , w_2789 );
and ( w_2788 , w_2789 , \944_b0 );
or ( \946_b1 , \d[5]_b1 , w_2790 );
xor ( \946_b0 , \d[5]_b0 , w_2792 );
not ( w_2792 , w_2793 );
and ( w_2793 , w_2790 , w_2791 );
buf ( w_2790 , \d[4]_b1 );
not ( w_2790 , w_2794 );
not ( w_2791 , w_2795 );
and ( w_2794 , w_2795 , \d[4]_b0 );
or ( \947_b1 , \d[4]_b1 , \d[3]_b1 );
xor ( \947_b0 , \d[4]_b0 , w_2796 );
not ( w_2796 , w_2797 );
and ( w_2797 , \d[3]_b1 , \d[3]_b0 );
or ( \948_b1 , \946_b1 , w_2799 );
not ( w_2799 , w_2800 );
and ( \948_b0 , \946_b0 , w_2801 );
and ( w_2800 ,  , w_2801 );
buf ( w_2799 , \947_b1 );
not ( w_2799 , w_2802 );
not (  , w_2803 );
and ( w_2802 , w_2803 , \947_b0 );
buf ( \949_b1 , \948_b1 );
not ( \949_b1 , w_2804 );
not ( \949_b0 , w_2805 );
and ( w_2804 , w_2805 , \948_b0 );
or ( \950_b1 , \945_b1 , w_2806 );
or ( \950_b0 , \945_b0 , \949_b0 );
not ( \949_b0 , w_2807 );
and ( w_2807 , w_2806 , \949_b1 );
buf ( \951_b1 , \947_b1 );
buf ( \951_b0 , \947_b0 );
or ( \952_b1 , \a[2]_b1 , \d[5]_b1 );
xor ( \952_b0 , \a[2]_b0 , w_2808 );
not ( w_2808 , w_2809 );
and ( w_2809 , \d[5]_b1 , \d[5]_b0 );
or ( \953_b1 , \951_b1 , w_2811 );
not ( w_2811 , w_2812 );
and ( \953_b0 , \951_b0 , w_2813 );
and ( w_2812 ,  , w_2813 );
buf ( w_2811 , \952_b1 );
not ( w_2811 , w_2814 );
not (  , w_2815 );
and ( w_2814 , w_2815 , \952_b0 );
or ( \954_b1 , \950_b1 , w_2817 );
not ( w_2817 , w_2818 );
and ( \954_b0 , \950_b0 , w_2819 );
and ( w_2818 ,  , w_2819 );
buf ( w_2817 , \953_b1 );
not ( w_2817 , w_2820 );
not (  , w_2821 );
and ( w_2820 , w_2821 , \953_b0 );
buf ( \955_b1 , \954_b1 );
not ( \955_b1 , w_2822 );
not ( \955_b0 , w_2823 );
and ( w_2822 , w_2823 , \954_b0 );
or ( \956_b1 , \943_b1 , \955_b1 );
xor ( \956_b0 , \943_b0 , w_2824 );
not ( w_2824 , w_2825 );
and ( w_2825 , \955_b1 , \955_b0 );
or ( \957_b1 , \d[6]_b1 , \d[5]_b1 );
xor ( \957_b0 , \d[6]_b0 , w_2826 );
not ( w_2826 , w_2827 );
and ( w_2827 , \d[5]_b1 , \d[5]_b0 );
buf ( \958_b1 , \957_b1 );
buf ( \958_b0 , \957_b0 );
or ( \959_b1 , \958_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_2828 );
and ( \959_b0 , \958_b0 , w_2829 );
and ( w_2828 , w_2829 , \a[0]_b0 );
buf ( \960_b1 , \935_b1 );
not ( \960_b1 , w_2830 );
not ( \960_b0 , w_2831 );
and ( w_2830 , w_2831 , \935_b0 );
buf ( \961_b1 , \932_b1 );
not ( \961_b1 , w_2832 );
not ( \961_b0 , w_2833 );
and ( w_2832 , w_2833 , \932_b0 );
or ( \962_b1 , \960_b1 , w_2834 );
or ( \962_b0 , \960_b0 , \961_b0 );
not ( \961_b0 , w_2835 );
and ( w_2835 , w_2834 , \961_b1 );
or ( \963_b1 , \a[6]_b1 , \d[1]_b1 );
xor ( \963_b0 , \a[6]_b0 , w_2836 );
not ( w_2836 , w_2837 );
and ( w_2837 , \d[1]_b1 , \d[1]_b0 );
or ( \964_b1 , \963_b1 , w_2839 );
not ( w_2839 , w_2840 );
and ( \964_b0 , \963_b0 , w_2841 );
and ( w_2840 ,  , w_2841 );
buf ( w_2839 , \d[0]_b1 );
not ( w_2839 , w_2842 );
not (  , w_2843 );
and ( w_2842 , w_2843 , \d[0]_b0 );
or ( \965_b1 , \962_b1 , w_2845 );
not ( w_2845 , w_2846 );
and ( \965_b0 , \962_b0 , w_2847 );
and ( w_2846 ,  , w_2847 );
buf ( w_2845 , \964_b1 );
not ( w_2845 , w_2848 );
not (  , w_2849 );
and ( w_2848 , w_2849 , \964_b0 );
or ( \966_b1 , \959_b1 , \965_b1 );
xor ( \966_b0 , \959_b0 , w_2850 );
not ( w_2850 , w_2851 );
and ( w_2851 , \965_b1 , \965_b0 );
or ( \967_b1 , \a[3]_b1 , \d[3]_b1 );
xor ( \967_b0 , \a[3]_b0 , w_2852 );
not ( w_2852 , w_2853 );
and ( w_2853 , \d[3]_b1 , \d[3]_b0 );
buf ( \968_b1 , \967_b1 );
not ( \968_b1 , w_2854 );
not ( \968_b0 , w_2855 );
and ( w_2854 , w_2855 , \967_b0 );
or ( \969_b1 , \d[2]_b1 , \d[1]_b1 );
xor ( \969_b0 , \d[2]_b0 , w_2856 );
not ( w_2856 , w_2857 );
and ( w_2857 , \d[1]_b1 , \d[1]_b0 );
buf ( \970_b1 , \969_b1 );
not ( \970_b1 , w_2858 );
not ( \970_b0 , w_2859 );
and ( w_2858 , w_2859 , \969_b0 );
or ( \971_b1 , \d[3]_b1 , \d[2]_b1 );
xor ( \971_b0 , \d[3]_b0 , w_2860 );
not ( w_2860 , w_2861 );
and ( w_2861 , \d[2]_b1 , \d[2]_b0 );
or ( \972_b1 , \970_b1 , w_2863 );
not ( w_2863 , w_2864 );
and ( \972_b0 , \970_b0 , w_2865 );
and ( w_2864 ,  , w_2865 );
buf ( w_2863 , \971_b1 );
not ( w_2863 , w_2866 );
not (  , w_2867 );
and ( w_2866 , w_2867 , \971_b0 );
buf ( \973_b1 , \972_b1 );
not ( \973_b1 , w_2868 );
not ( \973_b0 , w_2869 );
and ( w_2868 , w_2869 , \972_b0 );
buf ( \974_b1 , \973_b1 );
not ( \974_b1 , w_2870 );
not ( \974_b0 , w_2871 );
and ( w_2870 , w_2871 , \973_b0 );
or ( \975_b1 , \968_b1 , w_2872 );
or ( \975_b0 , \968_b0 , \974_b0 );
not ( \974_b0 , w_2873 );
and ( w_2873 , w_2872 , \974_b1 );
buf ( \976_b1 , \969_b1 );
buf ( \976_b0 , \969_b0 );
or ( \977_b1 , \a[4]_b1 , \d[3]_b1 );
xor ( \977_b0 , \a[4]_b0 , w_2874 );
not ( w_2874 , w_2875 );
and ( w_2875 , \d[3]_b1 , \d[3]_b0 );
or ( \978_b1 , \976_b1 , w_2877 );
not ( w_2877 , w_2878 );
and ( \978_b0 , \976_b0 , w_2879 );
and ( w_2878 ,  , w_2879 );
buf ( w_2877 , \977_b1 );
not ( w_2877 , w_2880 );
not (  , w_2881 );
and ( w_2880 , w_2881 , \977_b0 );
or ( \979_b1 , \975_b1 , w_2883 );
not ( w_2883 , w_2884 );
and ( \979_b0 , \975_b0 , w_2885 );
and ( w_2884 ,  , w_2885 );
buf ( w_2883 , \978_b1 );
not ( w_2883 , w_2886 );
not (  , w_2887 );
and ( w_2886 , w_2887 , \978_b0 );
or ( \980_b1 , \966_b1 , \979_b1 );
xor ( \980_b0 , \966_b0 , w_2888 );
not ( w_2888 , w_2889 );
and ( w_2889 , \979_b1 , \979_b0 );
or ( \981_b1 , \956_b1 , w_2890 );
xor ( \981_b0 , \956_b0 , w_2892 );
not ( w_2892 , w_2893 );
and ( w_2893 , w_2890 , w_2891 );
buf ( w_2890 , \980_b1 );
not ( w_2890 , w_2894 );
not ( w_2891 , w_2895 );
and ( w_2894 , w_2895 , \980_b0 );
buf ( \982_b1 , \981_b1 );
not ( \982_b1 , w_2896 );
not ( \982_b0 , w_2897 );
and ( w_2896 , w_2897 , \981_b0 );
or ( \983_b1 , \a[0]_b1 , \d[5]_b1 );
xor ( \983_b0 , \a[0]_b0 , w_2898 );
not ( w_2898 , w_2899 );
and ( w_2899 , \d[5]_b1 , \d[5]_b0 );
buf ( \984_b1 , \983_b1 );
not ( \984_b1 , w_2900 );
not ( \984_b0 , w_2901 );
and ( w_2900 , w_2901 , \983_b0 );
buf ( \985_b1 , \948_b1 );
not ( \985_b1 , w_2902 );
not ( \985_b0 , w_2903 );
and ( w_2902 , w_2903 , \948_b0 );
or ( \986_b1 , \984_b1 , w_2904 );
or ( \986_b0 , \984_b0 , \985_b0 );
not ( \985_b0 , w_2905 );
and ( w_2905 , w_2904 , \985_b1 );
or ( \987_b1 , \951_b1 , w_2907 );
not ( w_2907 , w_2908 );
and ( \987_b0 , \951_b0 , w_2909 );
and ( w_2908 ,  , w_2909 );
buf ( w_2907 , \944_b1 );
not ( w_2907 , w_2910 );
not (  , w_2911 );
and ( w_2910 , w_2911 , \944_b0 );
or ( \988_b1 , \986_b1 , w_2913 );
not ( w_2913 , w_2914 );
and ( \988_b0 , \986_b0 , w_2915 );
and ( w_2914 ,  , w_2915 );
buf ( w_2913 , \987_b1 );
not ( w_2913 , w_2916 );
not (  , w_2917 );
and ( w_2916 , w_2917 , \987_b0 );
buf ( \989_b1 , \988_b1 );
not ( \989_b1 , w_2918 );
not ( \989_b0 , w_2919 );
and ( w_2918 , w_2919 , \988_b0 );
buf ( \990_b1 , \989_b1 );
not ( \990_b1 , w_2920 );
not ( \990_b0 , w_2921 );
and ( w_2920 , w_2921 , \989_b0 );
buf ( \991_b1 , \937_b1 );
not ( \991_b1 , w_2922 );
not ( \991_b0 , w_2923 );
and ( w_2922 , w_2923 , \937_b0 );
buf ( \992_b1 , \942_b1 );
not ( \992_b1 , w_2924 );
not ( \992_b0 , w_2925 );
and ( w_2924 , w_2925 , \942_b0 );
or ( \993_b1 , \991_b1 , \992_b1 );
not ( \992_b1 , w_2926 );
and ( \993_b0 , \991_b0 , w_2927 );
and ( w_2926 , w_2927 , \992_b0 );
or ( \994_b1 , \937_b1 , \942_b1 );
not ( \942_b1 , w_2928 );
and ( \994_b0 , \937_b0 , w_2929 );
and ( w_2928 , w_2929 , \942_b0 );
or ( \995_b1 , \993_b1 , w_2931 );
not ( w_2931 , w_2932 );
and ( \995_b0 , \993_b0 , w_2933 );
and ( w_2932 ,  , w_2933 );
buf ( w_2931 , \994_b1 );
not ( w_2931 , w_2934 );
not (  , w_2935 );
and ( w_2934 , w_2935 , \994_b0 );
buf ( \996_b1 , \995_b1 );
not ( \996_b1 , w_2936 );
not ( \996_b0 , w_2937 );
and ( w_2936 , w_2937 , \995_b0 );
or ( \997_b1 , \990_b1 , w_2938 );
or ( \997_b0 , \990_b0 , \996_b0 );
not ( \996_b0 , w_2939 );
and ( w_2939 , w_2938 , \996_b1 );
or ( \998_b1 , \a[2]_b1 , \d[3]_b1 );
xor ( \998_b0 , \a[2]_b0 , w_2940 );
not ( w_2940 , w_2941 );
and ( w_2941 , \d[3]_b1 , \d[3]_b0 );
buf ( \999_b1 , \998_b1 );
not ( \999_b1 , w_2942 );
not ( \999_b0 , w_2943 );
and ( w_2942 , w_2943 , \998_b0 );
buf ( \1000_b1 , \973_b1 );
not ( \1000_b1 , w_2944 );
not ( \1000_b0 , w_2945 );
and ( w_2944 , w_2945 , \973_b0 );
or ( \1001_b1 , \999_b1 , w_2946 );
or ( \1001_b0 , \999_b0 , \1000_b0 );
not ( \1000_b0 , w_2947 );
and ( w_2947 , w_2946 , \1000_b1 );
or ( \1002_b1 , \976_b1 , w_2949 );
not ( w_2949 , w_2950 );
and ( \1002_b0 , \976_b0 , w_2951 );
and ( w_2950 ,  , w_2951 );
buf ( w_2949 , \967_b1 );
not ( w_2949 , w_2952 );
not (  , w_2953 );
and ( w_2952 , w_2953 , \967_b0 );
or ( \1003_b1 , \1001_b1 , w_2955 );
not ( w_2955 , w_2956 );
and ( \1003_b0 , \1001_b0 , w_2957 );
and ( w_2956 ,  , w_2957 );
buf ( w_2955 , \1002_b1 );
not ( w_2955 , w_2958 );
not (  , w_2959 );
and ( w_2958 , w_2959 , \1002_b0 );
or ( \1004_b1 , \997_b1 , w_2961 );
not ( w_2961 , w_2962 );
and ( \1004_b0 , \997_b0 , w_2963 );
and ( w_2962 ,  , w_2963 );
buf ( w_2961 , \1003_b1 );
not ( w_2961 , w_2964 );
not (  , w_2965 );
and ( w_2964 , w_2965 , \1003_b0 );
or ( \1005_b1 , \995_b1 , w_2966 );
or ( \1005_b0 , \995_b0 , \989_b0 );
not ( \989_b0 , w_2967 );
and ( w_2967 , w_2966 , \989_b1 );
or ( \1006_b1 , \1004_b1 , w_2969 );
not ( w_2969 , w_2970 );
and ( \1006_b0 , \1004_b0 , w_2971 );
and ( w_2970 ,  , w_2971 );
buf ( w_2969 , \1005_b1 );
not ( w_2969 , w_2972 );
not (  , w_2973 );
and ( w_2972 , w_2973 , \1005_b0 );
buf ( \1007_b1 , \1006_b1 );
not ( \1007_b1 , w_2974 );
not ( \1007_b0 , w_2975 );
and ( w_2974 , w_2975 , \1006_b0 );
or ( \1008_b1 , \982_b1 , w_2977 );
not ( w_2977 , w_2978 );
and ( \1008_b0 , \982_b0 , w_2979 );
and ( w_2978 ,  , w_2979 );
buf ( w_2977 , \1007_b1 );
not ( w_2977 , w_2980 );
not (  , w_2981 );
and ( w_2980 , w_2981 , \1007_b0 );
buf ( \1009_b1 , \1008_b1 );
not ( \1009_b1 , w_2982 );
not ( \1009_b0 , w_2983 );
and ( w_2982 , w_2983 , \1008_b0 );
or ( \1010_b1 , \988_b1 , \995_b1 );
xor ( \1010_b0 , \988_b0 , w_2984 );
not ( w_2984 , w_2985 );
and ( w_2985 , \995_b1 , \995_b0 );
or ( \1011_b1 , \1010_b1 , \1003_b1 );
xor ( \1011_b0 , \1010_b0 , w_2986 );
not ( w_2986 , w_2987 );
and ( w_2987 , \1003_b1 , \1003_b0 );
or ( \1012_b1 , \951_b1 , w_2989 );
not ( w_2989 , w_2990 );
and ( \1012_b0 , \951_b0 , w_2991 );
and ( w_2990 ,  , w_2991 );
buf ( w_2989 , \a[0]_b1 );
not ( w_2989 , w_2992 );
not (  , w_2993 );
and ( w_2992 , w_2993 , \a[0]_b0 );
or ( \1013_b1 , \976_b1 , \998_b1 );
not ( \998_b1 , w_2994 );
and ( \1013_b0 , \976_b0 , w_2995 );
and ( w_2994 , w_2995 , \998_b0 );
buf ( \1014_b1 , \976_b1 );
not ( \1014_b1 , w_2996 );
not ( \1014_b0 , w_2997 );
and ( w_2996 , w_2997 , \976_b0 );
or ( \1015_b1 , \a[1]_b1 , \d[3]_b1 );
xor ( \1015_b0 , \a[1]_b0 , w_2998 );
not ( w_2998 , w_2999 );
and ( w_2999 , \d[3]_b1 , \d[3]_b0 );
or ( \1016_b1 , \971_b1 , \1015_b1 );
not ( \1015_b1 , w_3000 );
and ( \1016_b0 , \971_b0 , w_3001 );
and ( w_3000 , w_3001 , \1015_b0 );
or ( \1017_b1 , \1014_b1 , \1016_b1 );
not ( \1016_b1 , w_3002 );
and ( \1017_b0 , \1014_b0 , w_3003 );
and ( w_3002 , w_3003 , \1016_b0 );
or ( \1018_b1 , \1013_b1 , w_3005 );
not ( w_3005 , w_3006 );
and ( \1018_b0 , \1013_b0 , w_3007 );
and ( w_3006 ,  , w_3007 );
buf ( w_3005 , \1017_b1 );
not ( w_3005 , w_3008 );
not (  , w_3009 );
and ( w_3008 , w_3009 , \1017_b0 );
or ( \1019_b1 , \1012_b1 , \1018_b1 );
xor ( \1019_b0 , \1012_b0 , w_3010 );
not ( w_3010 , w_3011 );
and ( w_3011 , \1018_b1 , \1018_b0 );
or ( \1020_b1 , \a[3]_b1 , \d[1]_b1 );
xor ( \1020_b0 , \a[3]_b0 , w_3012 );
not ( w_3012 , w_3013 );
and ( w_3013 , \d[1]_b1 , \d[1]_b0 );
or ( \1021_b1 , \932_b1 , \1020_b1 );
not ( \1020_b1 , w_3014 );
and ( \1021_b0 , \932_b0 , w_3015 );
and ( w_3014 , w_3015 , \1020_b0 );
or ( \1022_b1 , \928_b1 , \d[0]_b1 );
not ( \d[0]_b1 , w_3016 );
and ( \1022_b0 , \928_b0 , w_3017 );
and ( w_3016 , w_3017 , \d[0]_b0 );
or ( \1023_b1 , \1021_b1 , w_3019 );
not ( w_3019 , w_3020 );
and ( \1023_b0 , \1021_b0 , w_3021 );
and ( w_3020 ,  , w_3021 );
buf ( w_3019 , \1022_b1 );
not ( w_3019 , w_3022 );
not (  , w_3023 );
and ( w_3022 , w_3023 , \1022_b0 );
or ( \1024_b1 , \1019_b1 , \1023_b1 );
not ( \1023_b1 , w_3024 );
and ( \1024_b0 , \1019_b0 , w_3025 );
and ( w_3024 , w_3025 , \1023_b0 );
or ( \1025_b1 , \1012_b1 , \1018_b1 );
not ( \1018_b1 , w_3026 );
and ( \1025_b0 , \1012_b0 , w_3027 );
and ( w_3026 , w_3027 , \1018_b0 );
or ( \1026_b1 , \1024_b1 , w_3028 );
or ( \1026_b0 , \1024_b0 , \1025_b0 );
not ( \1025_b0 , w_3029 );
and ( w_3029 , w_3028 , \1025_b1 );
or ( \1027_b1 , \1011_b1 , w_3031 );
not ( w_3031 , w_3032 );
and ( \1027_b0 , \1011_b0 , w_3033 );
and ( w_3032 ,  , w_3033 );
buf ( w_3031 , \1026_b1 );
not ( w_3031 , w_3034 );
not (  , w_3035 );
and ( w_3034 , w_3035 , \1026_b0 );
or ( \1028_b1 , \976_b1 , w_3037 );
not ( w_3037 , w_3038 );
and ( \1028_b0 , \976_b0 , w_3039 );
and ( w_3038 ,  , w_3039 );
buf ( w_3037 , \a[0]_b1 );
not ( w_3037 , w_3040 );
not (  , w_3041 );
and ( w_3040 , w_3041 , \a[0]_b0 );
buf ( \1029_b1 , \1028_b1 );
not ( \1029_b1 , w_3042 );
not ( \1029_b0 , w_3043 );
and ( w_3042 , w_3043 , \1028_b0 );
or ( \1030_b1 , \a[1]_b1 , \d[1]_b1 );
xor ( \1030_b0 , \a[1]_b0 , w_3044 );
not ( w_3044 , w_3045 );
and ( w_3045 , \d[1]_b1 , \d[1]_b0 );
buf ( \1031_b1 , \1030_b1 );
not ( \1031_b1 , w_3046 );
not ( \1031_b0 , w_3047 );
and ( w_3046 , w_3047 , \1030_b0 );
buf ( \1032_b1 , \932_b1 );
not ( \1032_b1 , w_3048 );
not ( \1032_b0 , w_3049 );
and ( w_3048 , w_3049 , \932_b0 );
or ( \1033_b1 , \1031_b1 , w_3050 );
or ( \1033_b0 , \1031_b0 , \1032_b0 );
not ( \1032_b0 , w_3051 );
and ( w_3051 , w_3050 , \1032_b1 );
or ( \1034_b1 , \a[2]_b1 , \d[1]_b1 );
xor ( \1034_b0 , \a[2]_b0 , w_3052 );
not ( w_3052 , w_3053 );
and ( w_3053 , \d[1]_b1 , \d[1]_b0 );
or ( \1035_b1 , \1034_b1 , w_3055 );
not ( w_3055 , w_3056 );
and ( \1035_b0 , \1034_b0 , w_3057 );
and ( w_3056 ,  , w_3057 );
buf ( w_3055 , \d[0]_b1 );
not ( w_3055 , w_3058 );
not (  , w_3059 );
and ( w_3058 , w_3059 , \d[0]_b0 );
or ( \1036_b1 , \1033_b1 , w_3061 );
not ( w_3061 , w_3062 );
and ( \1036_b0 , \1033_b0 , w_3063 );
and ( w_3062 ,  , w_3063 );
buf ( w_3061 , \1035_b1 );
not ( w_3061 , w_3064 );
not (  , w_3065 );
and ( w_3064 , w_3065 , \1035_b0 );
or ( \1037_b1 , \1029_b1 , w_3067 );
not ( w_3067 , w_3068 );
and ( \1037_b0 , \1029_b0 , w_3069 );
and ( w_3068 ,  , w_3069 );
buf ( w_3067 , \1036_b1 );
not ( w_3067 , w_3070 );
not (  , w_3071 );
and ( w_3070 , w_3071 , \1036_b0 );
or ( \1038_b1 , \a[0]_b1 , \d[1]_b1 );
xor ( \1038_b0 , \a[0]_b0 , w_3072 );
not ( w_3072 , w_3073 );
and ( w_3073 , \d[1]_b1 , \d[1]_b0 );
buf ( \1039_b1 , \1038_b1 );
not ( \1039_b1 , w_3074 );
not ( \1039_b0 , w_3075 );
and ( w_3074 , w_3075 , \1038_b0 );
buf ( \1040_b1 , \932_b1 );
not ( \1040_b1 , w_3076 );
not ( \1040_b0 , w_3077 );
and ( w_3076 , w_3077 , \932_b0 );
or ( \1041_b1 , \1039_b1 , w_3078 );
or ( \1041_b0 , \1039_b0 , \1040_b0 );
not ( \1040_b0 , w_3079 );
and ( w_3079 , w_3078 , \1040_b1 );
or ( \1042_b1 , \1030_b1 , w_3081 );
not ( w_3081 , w_3082 );
and ( \1042_b0 , \1030_b0 , w_3083 );
and ( w_3082 ,  , w_3083 );
buf ( w_3081 , \d[0]_b1 );
not ( w_3081 , w_3084 );
not (  , w_3085 );
and ( w_3084 , w_3085 , \d[0]_b0 );
or ( \1043_b1 , \1041_b1 , w_3087 );
not ( w_3087 , w_3088 );
and ( \1043_b0 , \1041_b0 , w_3089 );
and ( w_3088 ,  , w_3089 );
buf ( w_3087 , \1042_b1 );
not ( w_3087 , w_3090 );
not (  , w_3091 );
and ( w_3090 , w_3091 , \1042_b0 );
or ( \1044_b1 , \a[0]_b1 , w_3093 );
not ( w_3093 , w_3094 );
and ( \1044_b0 , \a[0]_b0 , w_3095 );
and ( w_3094 ,  , w_3095 );
buf ( w_3093 , \d[0]_b1 );
not ( w_3093 , w_3096 );
not (  , w_3097 );
and ( w_3096 , w_3097 , \d[0]_b0 );
or ( \1045_b1 , \1044_b1 , \d[1]_b1 );
not ( \d[1]_b1 , w_3098 );
and ( \1045_b0 , \1044_b0 , w_3099 );
and ( w_3098 , w_3099 , \d[1]_b0 );
or ( \1046_b1 , \1043_b1 , w_3101 );
not ( w_3101 , w_3102 );
and ( \1046_b0 , \1043_b0 , w_3103 );
and ( w_3102 ,  , w_3103 );
buf ( w_3101 , \1045_b1 );
not ( w_3101 , w_3104 );
not (  , w_3105 );
and ( w_3104 , w_3105 , \1045_b0 );
or ( \1047_b1 , \1037_b1 , w_3106 );
or ( \1047_b0 , \1037_b0 , \1046_b0 );
not ( \1046_b0 , w_3107 );
and ( w_3107 , w_3106 , \1046_b1 );
buf ( \1048_b1 , \1028_b1 );
not ( \1048_b1 , w_3108 );
not ( \1048_b0 , w_3109 );
and ( w_3108 , w_3109 , \1028_b0 );
or ( \1049_b1 , \1048_b1 , w_3111 );
not ( w_3111 , w_3112 );
and ( \1049_b0 , \1048_b0 , w_3113 );
and ( w_3112 ,  , w_3113 );
buf ( w_3111 , \1036_b1 );
not ( w_3111 , w_3114 );
not (  , w_3115 );
and ( w_3114 , w_3115 , \1036_b0 );
or ( \1050_b1 , \1047_b1 , w_3117 );
not ( w_3117 , w_3118 );
and ( \1050_b0 , \1047_b0 , w_3119 );
and ( w_3118 ,  , w_3119 );
buf ( w_3117 , \1049_b1 );
not ( w_3117 , w_3120 );
not (  , w_3121 );
and ( w_3120 , w_3121 , \1049_b0 );
buf ( \1051_b1 , \1050_b1 );
not ( \1051_b1 , w_3122 );
not ( \1051_b0 , w_3123 );
and ( w_3122 , w_3123 , \1050_b0 );
buf ( \1052_b1 , \1034_b1 );
not ( \1052_b1 , w_3124 );
not ( \1052_b0 , w_3125 );
and ( w_3124 , w_3125 , \1034_b0 );
buf ( \1053_b1 , \932_b1 );
not ( \1053_b1 , w_3126 );
not ( \1053_b0 , w_3127 );
and ( w_3126 , w_3127 , \932_b0 );
or ( \1054_b1 , \1052_b1 , w_3128 );
or ( \1054_b0 , \1052_b0 , \1053_b0 );
not ( \1053_b0 , w_3129 );
and ( w_3129 , w_3128 , \1053_b1 );
or ( \1055_b1 , \d[0]_b1 , w_3131 );
not ( w_3131 , w_3132 );
and ( \1055_b0 , \d[0]_b0 , w_3133 );
and ( w_3132 ,  , w_3133 );
buf ( w_3131 , \1020_b1 );
not ( w_3131 , w_3134 );
not (  , w_3135 );
and ( w_3134 , w_3135 , \1020_b0 );
or ( \1056_b1 , \1054_b1 , w_3137 );
not ( w_3137 , w_3138 );
and ( \1056_b0 , \1054_b0 , w_3139 );
and ( w_3138 ,  , w_3139 );
buf ( w_3137 , \1055_b1 );
not ( w_3137 , w_3140 );
not (  , w_3141 );
and ( w_3140 , w_3141 , \1055_b0 );
buf ( \1057_b1 , \1056_b1 );
not ( \1057_b1 , w_3142 );
not ( \1057_b0 , w_3143 );
and ( w_3142 , w_3143 , \1056_b0 );
or ( \1058_b1 , \a[0]_b1 , w_3145 );
not ( w_3145 , w_3146 );
and ( \1058_b0 , \a[0]_b0 , w_3147 );
and ( w_3146 ,  , w_3147 );
buf ( w_3145 , \d[2]_b1 );
not ( w_3145 , w_3148 );
not (  , w_3149 );
and ( w_3148 , w_3149 , \d[2]_b0 );
or ( \1059_b1 , \1058_b1 , \d[3]_b1 );
not ( \d[3]_b1 , w_3150 );
and ( \1059_b0 , \1058_b0 , w_3151 );
and ( w_3150 , w_3151 , \d[3]_b0 );
or ( \1060_b1 , \a[0]_b1 , w_3152 );
or ( \1060_b0 , \a[0]_b0 , \d[2]_b0 );
not ( \d[2]_b0 , w_3153 );
and ( w_3153 , w_3152 , \d[2]_b1 );
or ( \1061_b1 , \1060_b1 , w_3155 );
not ( w_3155 , w_3156 );
and ( \1061_b0 , \1060_b0 , w_3157 );
and ( w_3156 ,  , w_3157 );
buf ( w_3155 , \d[1]_b1 );
not ( w_3155 , w_3158 );
not (  , w_3159 );
and ( w_3158 , w_3159 , \d[1]_b0 );
or ( \1062_b1 , \1059_b1 , w_3161 );
not ( w_3161 , w_3162 );
and ( \1062_b0 , \1059_b0 , w_3163 );
and ( w_3162 ,  , w_3163 );
buf ( w_3161 , \1061_b1 );
not ( w_3161 , w_3164 );
not (  , w_3165 );
and ( w_3164 , w_3165 , \1061_b0 );
buf ( \1063_b1 , \1062_b1 );
not ( \1063_b1 , w_3166 );
not ( \1063_b0 , w_3167 );
and ( w_3166 , w_3167 , \1062_b0 );
or ( \1064_b1 , \1057_b1 , \1063_b1 );
not ( \1063_b1 , w_3168 );
and ( \1064_b0 , \1057_b0 , w_3169 );
and ( w_3168 , w_3169 , \1063_b0 );
or ( \1065_b1 , \1056_b1 , \1062_b1 );
not ( \1062_b1 , w_3170 );
and ( \1065_b0 , \1056_b0 , w_3171 );
and ( w_3170 , w_3171 , \1062_b0 );
or ( \1066_b1 , \1064_b1 , w_3173 );
not ( w_3173 , w_3174 );
and ( \1066_b0 , \1064_b0 , w_3175 );
and ( w_3174 ,  , w_3175 );
buf ( w_3173 , \1065_b1 );
not ( w_3173 , w_3176 );
not (  , w_3177 );
and ( w_3176 , w_3177 , \1065_b0 );
buf ( \1067_b1 , \973_b1 );
buf ( \1067_b0 , \973_b0 );
or ( \1068_b1 , \a[0]_b1 , \d[3]_b1 );
xor ( \1068_b0 , \a[0]_b0 , w_3178 );
not ( w_3178 , w_3179 );
and ( w_3179 , \d[3]_b1 , \d[3]_b0 );
or ( \1069_b1 , \1067_b1 , w_3181 );
not ( w_3181 , w_3182 );
and ( \1069_b0 , \1067_b0 , w_3183 );
and ( w_3182 ,  , w_3183 );
buf ( w_3181 , \1068_b1 );
not ( w_3181 , w_3184 );
not (  , w_3185 );
and ( w_3184 , w_3185 , \1068_b0 );
or ( \1070_b1 , \976_b1 , w_3187 );
not ( w_3187 , w_3188 );
and ( \1070_b0 , \976_b0 , w_3189 );
and ( w_3188 ,  , w_3189 );
buf ( w_3187 , \1015_b1 );
not ( w_3187 , w_3190 );
not (  , w_3191 );
and ( w_3190 , w_3191 , \1015_b0 );
buf ( \1072_b1 , \1071_b1 );
not ( \1072_b1 , w_3192 );
not ( \1072_b0 , w_3193 );
and ( w_3192 , w_3193 , \1071_b0 );
or ( \1073_b1 , \1051_b1 , w_3194 );
or ( \1073_b0 , \1051_b0 , \1072_b0 );
not ( \1072_b0 , w_3195 );
and ( w_3195 , w_3194 , \1072_b1 );
buf ( \1074_b1 , \1066_b1 );
not ( \1074_b1 , w_3196 );
not ( \1074_b0 , w_3197 );
and ( w_3196 , w_3197 , \1066_b0 );
or ( \1075_b1 , \1069_b1 , w_3199 );
not ( w_3199 , w_3200 );
and ( \1075_b0 , \1069_b0 , w_3201 );
and ( w_3200 ,  , w_3201 );
buf ( w_3199 , \1070_b1 );
not ( w_3199 , w_3202 );
not (  , w_3203 );
and ( w_3202 , w_3203 , \1070_b0 );
or ( \1076_b1 , \1074_b1 , w_3205 );
not ( w_3205 , w_3206 );
and ( \1076_b0 , \1074_b0 , w_3207 );
and ( w_3206 ,  , w_3207 );
buf ( w_3205 , \1075_b1 );
not ( w_3205 , w_3208 );
not (  , w_3209 );
and ( w_3208 , w_3209 , \1075_b0 );
or ( \1077_b1 , \1073_b1 , w_3211 );
not ( w_3211 , w_3212 );
and ( \1077_b0 , \1073_b0 , w_3213 );
and ( w_3212 ,  , w_3213 );
buf ( w_3211 , \1076_b1 );
not ( w_3211 , w_3214 );
not (  , w_3215 );
and ( w_3214 , w_3215 , \1076_b0 );
buf ( \1078_b1 , \1077_b1 );
not ( \1078_b1 , w_3216 );
not ( \1078_b0 , w_3217 );
and ( w_3216 , w_3217 , \1077_b0 );
or ( \1079_b1 , \1012_b1 , \1018_b1 );
xor ( \1079_b0 , \1012_b0 , w_3218 );
not ( w_3218 , w_3219 );
and ( w_3219 , \1018_b1 , \1018_b0 );
or ( \1080_b1 , \1079_b1 , \1023_b1 );
xor ( \1080_b0 , \1079_b0 , w_3220 );
not ( w_3220 , w_3221 );
and ( w_3221 , \1023_b1 , \1023_b0 );
buf ( \1081_b1 , \1062_b1 );
not ( \1081_b1 , w_3222 );
not ( \1081_b0 , w_3223 );
and ( w_3222 , w_3223 , \1062_b0 );
or ( \1082_b1 , \1081_b1 , w_3225 );
not ( w_3225 , w_3226 );
and ( \1082_b0 , \1081_b0 , w_3227 );
and ( w_3226 ,  , w_3227 );
buf ( w_3225 , \1056_b1 );
not ( w_3225 , w_3228 );
not (  , w_3229 );
and ( w_3228 , w_3229 , \1056_b0 );
or ( \1083_b1 , \1080_b1 , w_3231 );
not ( w_3231 , w_3232 );
and ( \1083_b0 , \1080_b0 , w_3233 );
and ( w_3232 ,  , w_3233 );
buf ( w_3231 , \1082_b1 );
not ( w_3231 , w_3234 );
not (  , w_3235 );
and ( w_3234 , w_3235 , \1082_b0 );
buf ( \1084_b1 , \1083_b1 );
not ( \1084_b1 , w_3236 );
not ( \1084_b0 , w_3237 );
and ( w_3236 , w_3237 , \1083_b0 );
or ( \1085_b1 , \1078_b1 , w_3238 );
or ( \1085_b0 , \1078_b0 , \1084_b0 );
not ( \1084_b0 , w_3239 );
and ( w_3239 , w_3238 , \1084_b1 );
buf ( \1086_b1 , \1080_b1 );
not ( \1086_b1 , w_3240 );
not ( \1086_b0 , w_3241 );
and ( w_3240 , w_3241 , \1080_b0 );
buf ( \1087_b1 , \1082_b1 );
not ( \1087_b1 , w_3242 );
not ( \1087_b0 , w_3243 );
and ( w_3242 , w_3243 , \1082_b0 );
or ( \1088_b1 , \1086_b1 , w_3245 );
not ( w_3245 , w_3246 );
and ( \1088_b0 , \1086_b0 , w_3247 );
and ( w_3246 ,  , w_3247 );
buf ( w_3245 , \1087_b1 );
not ( w_3245 , w_3248 );
not (  , w_3249 );
and ( w_3248 , w_3249 , \1087_b0 );
or ( \1089_b1 , \1085_b1 , w_3251 );
not ( w_3251 , w_3252 );
and ( \1089_b0 , \1085_b0 , w_3253 );
and ( w_3252 ,  , w_3253 );
buf ( w_3251 , \1088_b1 );
not ( w_3251 , w_3254 );
not (  , w_3255 );
and ( w_3254 , w_3255 , \1088_b0 );
or ( \1090_b1 , \1027_b1 , \1089_b1 );
not ( \1089_b1 , w_3256 );
and ( \1090_b0 , \1027_b0 , w_3257 );
and ( w_3256 , w_3257 , \1089_b0 );
buf ( \1091_b1 , \1090_b1 );
not ( \1091_b1 , w_3258 );
not ( \1091_b0 , w_3259 );
and ( w_3258 , w_3259 , \1090_b0 );
or ( \1092_b1 , \1009_b1 , w_3260 );
or ( \1092_b0 , \1009_b0 , \1091_b0 );
not ( \1091_b0 , w_3261 );
and ( w_3261 , w_3260 , \1091_b1 );
buf ( \1093_b1 , \1011_b1 );
not ( \1093_b1 , w_3262 );
not ( \1093_b0 , w_3263 );
and ( w_3262 , w_3263 , \1011_b0 );
buf ( \1094_b1 , \1026_b1 );
not ( \1094_b1 , w_3264 );
not ( \1094_b0 , w_3265 );
and ( w_3264 , w_3265 , \1026_b0 );
or ( \1095_b1 , \1093_b1 , w_3267 );
not ( w_3267 , w_3268 );
and ( \1095_b0 , \1093_b0 , w_3269 );
and ( w_3268 ,  , w_3269 );
buf ( w_3267 , \1094_b1 );
not ( w_3267 , w_3270 );
not (  , w_3271 );
and ( w_3270 , w_3271 , \1094_b0 );
buf ( \1096_b1 , \1095_b1 );
not ( \1096_b1 , w_3272 );
not ( \1096_b0 , w_3273 );
and ( w_3272 , w_3273 , \1095_b0 );
or ( \1097_b1 , \981_b1 , w_3275 );
not ( w_3275 , w_3276 );
and ( \1097_b0 , \981_b0 , w_3277 );
and ( w_3276 ,  , w_3277 );
buf ( w_3275 , \1006_b1 );
not ( w_3275 , w_3278 );
not (  , w_3279 );
and ( w_3278 , w_3279 , \1006_b0 );
buf ( \1098_b1 , \1097_b1 );
not ( \1098_b1 , w_3280 );
not ( \1098_b0 , w_3281 );
and ( w_3280 , w_3281 , \1097_b0 );
or ( \1099_b1 , \1096_b1 , w_3282 );
or ( \1099_b0 , \1096_b0 , \1098_b0 );
not ( \1098_b0 , w_3283 );
and ( w_3283 , w_3282 , \1098_b1 );
or ( \1100_b1 , \1099_b1 , w_3285 );
not ( w_3285 , w_3286 );
and ( \1100_b0 , \1099_b0 , w_3287 );
and ( w_3286 ,  , w_3287 );
buf ( w_3285 , \1008_b1 );
not ( w_3285 , w_3288 );
not (  , w_3289 );
and ( w_3288 , w_3289 , \1008_b0 );
or ( \1101_b1 , \1092_b1 , w_3291 );
not ( w_3291 , w_3292 );
and ( \1101_b0 , \1092_b0 , w_3293 );
and ( w_3292 ,  , w_3293 );
buf ( w_3291 , \1100_b1 );
not ( w_3291 , w_3294 );
not (  , w_3295 );
and ( w_3294 , w_3295 , \1100_b0 );
buf ( \1102_b1 , \1101_b1 );
not ( \1102_b1 , w_3296 );
not ( \1102_b0 , w_3297 );
and ( w_3296 , w_3297 , \1101_b0 );
buf ( \1103_b1 , \963_b1 );
not ( \1103_b1 , w_3298 );
not ( \1103_b0 , w_3299 );
and ( w_3298 , w_3299 , \963_b0 );
buf ( \1104_b1 , \932_b1 );
not ( \1104_b1 , w_3300 );
not ( \1104_b0 , w_3301 );
and ( w_3300 , w_3301 , \932_b0 );
or ( \1105_b1 , \1103_b1 , w_3302 );
or ( \1105_b0 , \1103_b0 , \1104_b0 );
not ( \1104_b0 , w_3303 );
and ( w_3303 , w_3302 , \1104_b1 );
or ( \1106_b1 , \a[7]_b1 , \d[1]_b1 );
xor ( \1106_b0 , \a[7]_b0 , w_3304 );
not ( w_3304 , w_3305 );
and ( w_3305 , \d[1]_b1 , \d[1]_b0 );
or ( \1107_b1 , \1106_b1 , w_3307 );
not ( w_3307 , w_3308 );
and ( \1107_b0 , \1106_b0 , w_3309 );
and ( w_3308 ,  , w_3309 );
buf ( w_3307 , \d[0]_b1 );
not ( w_3307 , w_3310 );
not (  , w_3311 );
and ( w_3310 , w_3311 , \d[0]_b0 );
or ( \1108_b1 , \1105_b1 , w_3313 );
not ( w_3313 , w_3314 );
and ( \1108_b0 , \1105_b0 , w_3315 );
and ( w_3314 ,  , w_3315 );
buf ( w_3313 , \1107_b1 );
not ( w_3313 , w_3316 );
not (  , w_3317 );
and ( w_3316 , w_3317 , \1107_b0 );
or ( \1109_b1 , \a[0]_b1 , w_3318 );
or ( \1109_b0 , \a[0]_b0 , \d[6]_b0 );
not ( \d[6]_b0 , w_3319 );
and ( w_3319 , w_3318 , \d[6]_b1 );
or ( \1110_b1 , \1109_b1 , w_3321 );
not ( w_3321 , w_3322 );
and ( \1110_b0 , \1109_b0 , w_3323 );
and ( w_3322 ,  , w_3323 );
buf ( w_3321 , \d[5]_b1 );
not ( w_3321 , w_3324 );
not (  , w_3325 );
and ( w_3324 , w_3325 , \d[5]_b0 );
or ( \1111_b1 , \a[0]_b1 , w_3327 );
not ( w_3327 , w_3328 );
and ( \1111_b0 , \a[0]_b0 , w_3329 );
and ( w_3328 ,  , w_3329 );
buf ( w_3327 , \d[6]_b1 );
not ( w_3327 , w_3330 );
not (  , w_3331 );
and ( w_3330 , w_3331 , \d[6]_b0 );
buf ( \1113_b1 , \1112_b1 );
not ( \1113_b1 , w_3332 );
not ( \1113_b0 , w_3333 );
and ( w_3332 , w_3333 , \1112_b0 );
or ( \1114_b1 , \1108_b1 , \1113_b1 );
not ( \1113_b1 , w_3334 );
and ( \1114_b0 , \1108_b0 , w_3335 );
and ( w_3334 , w_3335 , \1113_b0 );
buf ( \1115_b1 , \1108_b1 );
not ( \1115_b1 , w_3336 );
not ( \1115_b0 , w_3337 );
and ( w_3336 , w_3337 , \1108_b0 );
or ( \1116_b1 , \1115_b1 , \1112_b1 );
not ( \1112_b1 , w_3338 );
and ( \1116_b0 , \1115_b0 , w_3339 );
and ( w_3338 , w_3339 , \1112_b0 );
or ( \1117_b1 , \1114_b1 , w_3341 );
not ( w_3341 , w_3342 );
and ( \1117_b0 , \1114_b0 , w_3343 );
and ( w_3342 ,  , w_3343 );
buf ( w_3341 , \1116_b1 );
not ( w_3341 , w_3344 );
not (  , w_3345 );
and ( w_3344 , w_3345 , \1116_b0 );
or ( \1118_b1 , \959_b1 , \965_b1 );
xor ( \1118_b0 , \959_b0 , w_3346 );
not ( w_3346 , w_3347 );
and ( w_3347 , \965_b1 , \965_b0 );
or ( \1119_b1 , \1118_b1 , \979_b1 );
not ( \979_b1 , w_3348 );
and ( \1119_b0 , \1118_b0 , w_3349 );
and ( w_3348 , w_3349 , \979_b0 );
or ( \1120_b1 , \959_b1 , \965_b1 );
not ( \965_b1 , w_3350 );
and ( \1120_b0 , \959_b0 , w_3351 );
and ( w_3350 , w_3351 , \965_b0 );
or ( \1121_b1 , \1119_b1 , w_3352 );
or ( \1121_b0 , \1119_b0 , \1120_b0 );
not ( \1120_b0 , w_3353 );
and ( w_3353 , w_3352 , \1120_b1 );
or ( \1122_b1 , \1117_b1 , \1121_b1 );
xor ( \1122_b0 , \1117_b0 , w_3354 );
not ( w_3354 , w_3355 );
and ( w_3355 , \1121_b1 , \1121_b0 );
or ( \1123_b1 , \a[0]_b1 , \d[7]_b1 );
xor ( \1123_b0 , \a[0]_b0 , w_3356 );
not ( w_3356 , w_3357 );
and ( w_3357 , \d[7]_b1 , \d[7]_b0 );
buf ( \1124_b1 , \1123_b1 );
not ( \1124_b1 , w_3358 );
not ( \1124_b0 , w_3359 );
and ( w_3358 , w_3359 , \1123_b0 );
or ( \1125_b1 , \d[7]_b1 , \d[6]_b1 );
xor ( \1125_b0 , \d[7]_b0 , w_3360 );
not ( w_3360 , w_3361 );
and ( w_3361 , \d[6]_b1 , \d[6]_b0 );
buf ( \1126_b1 , \1125_b1 );
not ( \1126_b1 , w_3362 );
not ( \1126_b0 , w_3363 );
and ( w_3362 , w_3363 , \1125_b0 );
or ( \1127_b1 , \957_b1 , w_3365 );
not ( w_3365 , w_3366 );
and ( \1127_b0 , \957_b0 , w_3367 );
and ( w_3366 ,  , w_3367 );
buf ( w_3365 , \1126_b1 );
not ( w_3365 , w_3368 );
not (  , w_3369 );
and ( w_3368 , w_3369 , \1126_b0 );
buf ( \1128_b1 , \1127_b1 );
buf ( \1128_b0 , \1127_b0 );
buf ( \1129_b1 , \1128_b1 );
not ( \1129_b1 , w_3370 );
not ( \1129_b0 , w_3371 );
and ( w_3370 , w_3371 , \1128_b0 );
or ( \1130_b1 , \1124_b1 , w_3372 );
or ( \1130_b0 , \1124_b0 , \1129_b0 );
not ( \1129_b0 , w_3373 );
and ( w_3373 , w_3372 , \1129_b1 );
or ( \1131_b1 , \a[1]_b1 , \d[7]_b1 );
xor ( \1131_b0 , \a[1]_b0 , w_3374 );
not ( w_3374 , w_3375 );
and ( w_3375 , \d[7]_b1 , \d[7]_b0 );
or ( \1132_b1 , \958_b1 , w_3377 );
not ( w_3377 , w_3378 );
and ( \1132_b0 , \958_b0 , w_3379 );
and ( w_3378 ,  , w_3379 );
buf ( w_3377 , \1131_b1 );
not ( w_3377 , w_3380 );
not (  , w_3381 );
and ( w_3380 , w_3381 , \1131_b0 );
or ( \1133_b1 , \1130_b1 , w_3383 );
not ( w_3383 , w_3384 );
and ( \1133_b0 , \1130_b0 , w_3385 );
and ( w_3384 ,  , w_3385 );
buf ( w_3383 , \1132_b1 );
not ( w_3383 , w_3386 );
not (  , w_3387 );
and ( w_3386 , w_3387 , \1132_b0 );
buf ( \1134_b1 , \952_b1 );
not ( \1134_b1 , w_3388 );
not ( \1134_b0 , w_3389 );
and ( w_3388 , w_3389 , \952_b0 );
or ( \1135_b1 , \946_b1 , w_3391 );
not ( w_3391 , w_3392 );
and ( \1135_b0 , \946_b0 , w_3393 );
and ( w_3392 ,  , w_3393 );
buf ( w_3391 , \947_b1 );
not ( w_3391 , w_3394 );
not (  , w_3395 );
and ( w_3394 , w_3395 , \947_b0 );
buf ( \1136_b1 , \1135_b1 );
not ( \1136_b1 , w_3396 );
not ( \1136_b0 , w_3397 );
and ( w_3396 , w_3397 , \1135_b0 );
or ( \1137_b1 , \1134_b1 , w_3398 );
or ( \1137_b0 , \1134_b0 , \1136_b0 );
not ( \1136_b0 , w_3399 );
and ( w_3399 , w_3398 , \1136_b1 );
or ( \1138_b1 , \a[3]_b1 , \d[5]_b1 );
xor ( \1138_b0 , \a[3]_b0 , w_3400 );
not ( w_3400 , w_3401 );
and ( w_3401 , \d[5]_b1 , \d[5]_b0 );
or ( \1139_b1 , \951_b1 , w_3403 );
not ( w_3403 , w_3404 );
and ( \1139_b0 , \951_b0 , w_3405 );
and ( w_3404 ,  , w_3405 );
buf ( w_3403 , \1138_b1 );
not ( w_3403 , w_3406 );
not (  , w_3407 );
and ( w_3406 , w_3407 , \1138_b0 );
or ( \1140_b1 , \1137_b1 , w_3409 );
not ( w_3409 , w_3410 );
and ( \1140_b0 , \1137_b0 , w_3411 );
and ( w_3410 ,  , w_3411 );
buf ( w_3409 , \1139_b1 );
not ( w_3409 , w_3412 );
not (  , w_3413 );
and ( w_3412 , w_3413 , \1139_b0 );
or ( \1141_b1 , \1133_b1 , \1140_b1 );
xor ( \1141_b0 , \1133_b0 , w_3414 );
not ( w_3414 , w_3415 );
and ( w_3415 , \1140_b1 , \1140_b0 );
buf ( \1142_b1 , \977_b1 );
not ( \1142_b1 , w_3416 );
not ( \1142_b0 , w_3417 );
and ( w_3416 , w_3417 , \977_b0 );
buf ( \1143_b1 , \1067_b1 );
not ( \1143_b1 , w_3418 );
not ( \1143_b0 , w_3419 );
and ( w_3418 , w_3419 , \1067_b0 );
or ( \1144_b1 , \1142_b1 , w_3420 );
or ( \1144_b0 , \1142_b0 , \1143_b0 );
not ( \1143_b0 , w_3421 );
and ( w_3421 , w_3420 , \1143_b1 );
or ( \1145_b1 , \a[5]_b1 , \d[3]_b1 );
xor ( \1145_b0 , \a[5]_b0 , w_3422 );
not ( w_3422 , w_3423 );
and ( w_3423 , \d[3]_b1 , \d[3]_b0 );
or ( \1146_b1 , \976_b1 , w_3425 );
not ( w_3425 , w_3426 );
and ( \1146_b0 , \976_b0 , w_3427 );
and ( w_3426 ,  , w_3427 );
buf ( w_3425 , \1145_b1 );
not ( w_3425 , w_3428 );
not (  , w_3429 );
and ( w_3428 , w_3429 , \1145_b0 );
or ( \1147_b1 , \1144_b1 , w_3431 );
not ( w_3431 , w_3432 );
and ( \1147_b0 , \1144_b0 , w_3433 );
and ( w_3432 ,  , w_3433 );
buf ( w_3431 , \1146_b1 );
not ( w_3431 , w_3434 );
not (  , w_3435 );
and ( w_3434 , w_3435 , \1146_b0 );
or ( \1148_b1 , \1141_b1 , \1147_b1 );
xor ( \1148_b0 , \1141_b0 , w_3436 );
not ( w_3436 , w_3437 );
and ( w_3437 , \1147_b1 , \1147_b0 );
or ( \1149_b1 , \1122_b1 , \1148_b1 );
xor ( \1149_b0 , \1122_b0 , w_3438 );
not ( w_3438 , w_3439 );
and ( w_3439 , \1148_b1 , \1148_b0 );
buf ( \1150_b1 , \943_b1 );
not ( \1150_b1 , w_3440 );
not ( \1150_b0 , w_3441 );
and ( w_3440 , w_3441 , \943_b0 );
or ( \1151_b1 , \1150_b1 , w_3443 );
not ( w_3443 , w_3444 );
and ( \1151_b0 , \1150_b0 , w_3445 );
and ( w_3444 ,  , w_3445 );
buf ( w_3443 , \955_b1 );
not ( w_3443 , w_3446 );
not (  , w_3447 );
and ( w_3446 , w_3447 , \955_b0 );
buf ( \1152_b1 , \1151_b1 );
not ( \1152_b1 , w_3448 );
not ( \1152_b0 , w_3449 );
and ( w_3448 , w_3449 , \1151_b0 );
buf ( \1153_b1 , \980_b1 );
not ( \1153_b1 , w_3450 );
not ( \1153_b0 , w_3451 );
and ( w_3450 , w_3451 , \980_b0 );
or ( \1154_b1 , \1152_b1 , w_3452 );
or ( \1154_b0 , \1152_b0 , \1153_b0 );
not ( \1153_b0 , w_3453 );
and ( w_3453 , w_3452 , \1153_b1 );
or ( \1155_b1 , \943_b1 , w_3455 );
not ( w_3455 , w_3456 );
and ( \1155_b0 , \943_b0 , w_3457 );
and ( w_3456 ,  , w_3457 );
buf ( w_3455 , \954_b1 );
not ( w_3455 , w_3458 );
not (  , w_3459 );
and ( w_3458 , w_3459 , \954_b0 );
or ( \1156_b1 , \1154_b1 , w_3461 );
not ( w_3461 , w_3462 );
and ( \1156_b0 , \1154_b0 , w_3463 );
and ( w_3462 ,  , w_3463 );
buf ( w_3461 , \1155_b1 );
not ( w_3461 , w_3464 );
not (  , w_3465 );
and ( w_3464 , w_3465 , \1155_b0 );
or ( \1157_b1 , \1149_b1 , w_3466 );
or ( \1157_b0 , \1149_b0 , \1156_b0 );
not ( \1156_b0 , w_3467 );
and ( w_3467 , w_3466 , \1156_b1 );
or ( \1158_b1 , \1149_b1 , w_3469 );
not ( w_3469 , w_3470 );
and ( \1158_b0 , \1149_b0 , w_3471 );
and ( w_3470 ,  , w_3471 );
buf ( w_3469 , \1156_b1 );
not ( w_3469 , w_3472 );
not (  , w_3473 );
and ( w_3472 , w_3473 , \1156_b0 );
or ( \1159_b1 , \1157_b1 , w_3475 );
not ( w_3475 , w_3476 );
and ( \1159_b0 , \1157_b0 , w_3477 );
and ( w_3476 ,  , w_3477 );
buf ( w_3475 , \1158_b1 );
not ( w_3475 , w_3478 );
not (  , w_3479 );
and ( w_3478 , w_3479 , \1158_b0 );
buf ( \1160_b1 , \1159_b1 );
not ( \1160_b1 , w_3480 );
not ( \1160_b0 , w_3481 );
and ( w_3480 , w_3481 , \1159_b0 );
or ( \1161_b1 , \1102_b1 , w_3482 );
or ( \1161_b0 , \1102_b0 , \1160_b0 );
not ( \1160_b0 , w_3483 );
and ( w_3483 , w_3482 , \1160_b1 );
or ( \1162_b1 , \1159_b1 , w_3484 );
or ( \1162_b0 , \1159_b0 , \1101_b0 );
not ( \1101_b0 , w_3485 );
and ( w_3485 , w_3484 , \1101_b1 );
or ( \1163_b1 , \1161_b1 , w_3487 );
not ( w_3487 , w_3488 );
and ( \1163_b0 , \1161_b0 , w_3489 );
and ( w_3488 ,  , w_3489 );
buf ( w_3487 , \1162_b1 );
not ( w_3487 , w_3490 );
not (  , w_3491 );
and ( w_3490 , w_3491 , \1162_b0 );
or ( \1164_b1 , \403_b1 , \531_b1 );
not ( \531_b1 , w_3492 );
and ( \1164_b0 , \403_b0 , w_3493 );
and ( w_3492 , w_3493 , \531_b0 );
buf ( \1165_b1 , \529_b1 );
buf ( \1165_b0 , \529_b0 );
or ( \1166_b1 , \1164_b1 , \1165_b1 );
xor ( \1166_b0 , \1164_b0 , w_3494 );
not ( w_3494 , w_3495 );
and ( w_3495 , \1165_b1 , \1165_b0 );
buf ( \1167_b1 , \1166_b1 );
not ( \1167_b1 , w_3496 );
not ( \1167_b0 , w_3497 );
and ( w_3496 , w_3497 , \1166_b0 );
buf ( \1168_b1 , \1167_b1 );
not ( \1168_b1 , w_3498 );
not ( \1168_b0 , w_3499 );
and ( w_3498 , w_3499 , \1167_b0 );
or ( \1169_b1 , \1163_b1 , \1168_b1 );
not ( \1168_b1 , w_3500 );
and ( \1169_b0 , \1163_b0 , w_3501 );
and ( w_3500 , w_3501 , \1168_b0 );
or ( \1170_b1 , \b[2]_b1 , w_3503 );
not ( w_3503 , w_3504 );
and ( \1170_b0 , \b[2]_b0 , w_3505 );
and ( w_3504 ,  , w_3505 );
buf ( w_3503 , \d[2]_b1 );
not ( w_3503 , w_3506 );
not (  , w_3507 );
and ( w_3506 , w_3507 , \d[2]_b0 );
or ( \1171_b1 , \b[3]_b1 , w_3509 );
not ( w_3509 , w_3510 );
and ( \1171_b0 , \b[3]_b0 , w_3511 );
and ( w_3510 ,  , w_3511 );
buf ( w_3509 , \d[3]_b1 );
not ( w_3509 , w_3512 );
not (  , w_3513 );
and ( w_3512 , w_3513 , \d[3]_b0 );
or ( \1172_b1 , \1170_b1 , w_3515 );
not ( w_3515 , w_3516 );
and ( \1172_b0 , \1170_b0 , w_3517 );
and ( w_3516 ,  , w_3517 );
buf ( w_3515 , \1171_b1 );
not ( w_3515 , w_3518 );
not (  , w_3519 );
and ( w_3518 , w_3519 , \1171_b0 );
buf ( \1173_b1 , \1172_b1 );
not ( \1173_b1 , w_3520 );
not ( \1173_b0 , w_3521 );
and ( w_3520 , w_3521 , \1172_b0 );
or ( \1174_b1 , \b[0]_b1 , w_3523 );
not ( w_3523 , w_3524 );
and ( \1174_b0 , \b[0]_b0 , w_3525 );
and ( w_3524 ,  , w_3525 );
buf ( w_3523 , \d[0]_b1 );
not ( w_3523 , w_3526 );
not (  , w_3527 );
and ( w_3526 , w_3527 , \d[0]_b0 );
buf ( \1175_b1 , \1174_b1 );
not ( \1175_b1 , w_3528 );
not ( \1175_b0 , w_3529 );
and ( w_3528 , w_3529 , \1174_b0 );
buf ( \1176_b1 , \1175_b1 );
not ( \1176_b1 , w_3530 );
not ( \1176_b0 , w_3531 );
and ( w_3530 , w_3531 , \1175_b0 );
or ( \1177_b1 , \b[1]_b1 , w_3532 );
or ( \1177_b0 , \b[1]_b0 , \d[1]_b0 );
not ( \d[1]_b0 , w_3533 );
and ( w_3533 , w_3532 , \d[1]_b1 );
buf ( \1178_b1 , \1177_b1 );
not ( \1178_b1 , w_3534 );
not ( \1178_b0 , w_3535 );
and ( w_3534 , w_3535 , \1177_b0 );
or ( \1179_b1 , \1176_b1 , w_3536 );
or ( \1179_b0 , \1176_b0 , \1178_b0 );
not ( \1178_b0 , w_3537 );
and ( w_3537 , w_3536 , \1178_b1 );
or ( \1180_b1 , \b[1]_b1 , w_3539 );
not ( w_3539 , w_3540 );
and ( \1180_b0 , \b[1]_b0 , w_3541 );
and ( w_3540 ,  , w_3541 );
buf ( w_3539 , \d[1]_b1 );
not ( w_3539 , w_3542 );
not (  , w_3543 );
and ( w_3542 , w_3543 , \d[1]_b0 );
or ( \1181_b1 , \1179_b1 , w_3545 );
not ( w_3545 , w_3546 );
and ( \1181_b0 , \1179_b0 , w_3547 );
and ( w_3546 ,  , w_3547 );
buf ( w_3545 , \1180_b1 );
not ( w_3545 , w_3548 );
not (  , w_3549 );
and ( w_3548 , w_3549 , \1180_b0 );
buf ( \1182_b1 , \1181_b1 );
not ( \1182_b1 , w_3550 );
not ( \1182_b0 , w_3551 );
and ( w_3550 , w_3551 , \1181_b0 );
or ( \1183_b1 , \1173_b1 , w_3552 );
or ( \1183_b0 , \1173_b0 , \1182_b0 );
not ( \1182_b0 , w_3553 );
and ( w_3553 , w_3552 , \1182_b1 );
or ( \1184_b1 , \b[3]_b1 , w_3555 );
not ( w_3555 , w_3556 );
and ( \1184_b0 , \b[3]_b0 , w_3557 );
and ( w_3556 ,  , w_3557 );
buf ( w_3555 , \d[3]_b1 );
not ( w_3555 , w_3558 );
not (  , w_3559 );
and ( w_3558 , w_3559 , \d[3]_b0 );
buf ( \1185_b1 , \1184_b1 );
not ( \1185_b1 , w_3560 );
not ( \1185_b0 , w_3561 );
and ( w_3560 , w_3561 , \1184_b0 );
or ( \1186_b1 , \b[2]_b1 , w_3563 );
not ( w_3563 , w_3564 );
and ( \1186_b0 , \b[2]_b0 , w_3565 );
and ( w_3564 ,  , w_3565 );
buf ( w_3563 , \d[2]_b1 );
not ( w_3563 , w_3566 );
not (  , w_3567 );
and ( w_3566 , w_3567 , \d[2]_b0 );
or ( \1187_b1 , \1171_b1 , w_3569 );
not ( w_3569 , w_3570 );
and ( \1187_b0 , \1171_b0 , w_3571 );
and ( w_3570 ,  , w_3571 );
buf ( w_3569 , \1186_b1 );
not ( w_3569 , w_3572 );
not (  , w_3573 );
and ( w_3572 , w_3573 , \1186_b0 );
or ( \1188_b1 , \1185_b1 , w_3575 );
not ( w_3575 , w_3576 );
and ( \1188_b0 , \1185_b0 , w_3577 );
and ( w_3576 ,  , w_3577 );
buf ( w_3575 , \1187_b1 );
not ( w_3575 , w_3578 );
not (  , w_3579 );
and ( w_3578 , w_3579 , \1187_b0 );
or ( \1189_b1 , \1183_b1 , w_3581 );
not ( w_3581 , w_3582 );
and ( \1189_b0 , \1183_b0 , w_3583 );
and ( w_3582 ,  , w_3583 );
buf ( w_3581 , \1188_b1 );
not ( w_3581 , w_3584 );
not (  , w_3585 );
and ( w_3584 , w_3585 , \1188_b0 );
or ( \1190_b1 , \b[4]_b1 , w_3587 );
not ( w_3587 , w_3588 );
and ( \1190_b0 , \b[4]_b0 , w_3589 );
and ( w_3588 ,  , w_3589 );
buf ( w_3587 , \d[4]_b1 );
not ( w_3587 , w_3590 );
not (  , w_3591 );
and ( w_3590 , w_3591 , \d[4]_b0 );
buf ( \1191_b1 , \1190_b1 );
not ( \1191_b1 , w_3592 );
not ( \1191_b0 , w_3593 );
and ( w_3592 , w_3593 , \1190_b0 );
or ( \1192_b1 , \b[5]_b1 , w_3594 );
or ( \1192_b0 , \b[5]_b0 , \d[5]_b0 );
not ( \d[5]_b0 , w_3595 );
and ( w_3595 , w_3594 , \d[5]_b1 );
or ( \1193_b1 , \1191_b1 , w_3597 );
not ( w_3597 , w_3598 );
and ( \1193_b0 , \1191_b0 , w_3599 );
and ( w_3598 ,  , w_3599 );
buf ( w_3597 , \1192_b1 );
not ( w_3597 , w_3600 );
not (  , w_3601 );
and ( w_3600 , w_3601 , \1192_b0 );
or ( \1194_b1 , \b[6]_b1 , w_3603 );
not ( w_3603 , w_3604 );
and ( \1194_b0 , \b[6]_b0 , w_3605 );
and ( w_3604 ,  , w_3605 );
buf ( w_3603 , \d[6]_b1 );
not ( w_3603 , w_3606 );
not (  , w_3607 );
and ( w_3606 , w_3607 , \d[6]_b0 );
or ( \1195_b1 , \1193_b1 , w_3609 );
not ( w_3609 , w_3610 );
and ( \1195_b0 , \1193_b0 , w_3611 );
and ( w_3610 ,  , w_3611 );
buf ( w_3609 , \1194_b1 );
not ( w_3609 , w_3612 );
not (  , w_3613 );
and ( w_3612 , w_3613 , \1194_b0 );
or ( \1196_b1 , \1189_b1 , w_3615 );
not ( w_3615 , w_3616 );
and ( \1196_b0 , \1189_b0 , w_3617 );
and ( w_3616 ,  , w_3617 );
buf ( w_3615 , \1195_b1 );
not ( w_3615 , w_3618 );
not (  , w_3619 );
and ( w_3618 , w_3619 , \1195_b0 );
or ( \1197_b1 , \b[4]_b1 , w_3621 );
not ( w_3621 , w_3622 );
and ( \1197_b0 , \b[4]_b0 , w_3623 );
and ( w_3622 ,  , w_3623 );
buf ( w_3621 , \d[4]_b1 );
not ( w_3621 , w_3624 );
not (  , w_3625 );
and ( w_3624 , w_3625 , \d[4]_b0 );
buf ( \1198_b1 , \1197_b1 );
not ( \1198_b1 , w_3626 );
not ( \1198_b0 , w_3627 );
and ( w_3626 , w_3627 , \1197_b0 );
or ( \1199_b1 , \1192_b1 , w_3629 );
not ( w_3629 , w_3630 );
and ( \1199_b0 , \1192_b0 , w_3631 );
and ( w_3630 ,  , w_3631 );
buf ( w_3629 , \1198_b1 );
not ( w_3629 , w_3632 );
not (  , w_3633 );
and ( w_3632 , w_3633 , \1198_b0 );
or ( \1200_b1 , \b[5]_b1 , w_3635 );
not ( w_3635 , w_3636 );
and ( \1200_b0 , \b[5]_b0 , w_3637 );
and ( w_3636 ,  , w_3637 );
buf ( w_3635 , \d[5]_b1 );
not ( w_3635 , w_3638 );
not (  , w_3639 );
and ( w_3638 , w_3639 , \d[5]_b0 );
or ( \1201_b1 , \1199_b1 , w_3641 );
not ( w_3641 , w_3642 );
and ( \1201_b0 , \1199_b0 , w_3643 );
and ( w_3642 ,  , w_3643 );
buf ( w_3641 , \1200_b1 );
not ( w_3641 , w_3644 );
not (  , w_3645 );
and ( w_3644 , w_3645 , \1200_b0 );
buf ( \1202_b1 , \1194_b1 );
not ( \1202_b1 , w_3646 );
not ( \1202_b0 , w_3647 );
and ( w_3646 , w_3647 , \1194_b0 );
or ( \1203_b1 , \1201_b1 , \1202_b1 );
not ( \1202_b1 , w_3648 );
and ( \1203_b0 , \1201_b0 , w_3649 );
and ( w_3648 , w_3649 , \1202_b0 );
or ( \1204_b1 , \b[6]_b1 , w_3651 );
not ( w_3651 , w_3652 );
and ( \1204_b0 , \b[6]_b0 , w_3653 );
and ( w_3652 ,  , w_3653 );
buf ( w_3651 , \d[6]_b1 );
not ( w_3651 , w_3654 );
not (  , w_3655 );
and ( w_3654 , w_3655 , \d[6]_b0 );
buf ( \1205_b1 , \1204_b1 );
not ( \1205_b1 , w_3656 );
not ( \1205_b0 , w_3657 );
and ( w_3656 , w_3657 , \1204_b0 );
or ( \1206_b1 , \1203_b1 , w_3659 );
not ( w_3659 , w_3660 );
and ( \1206_b0 , \1203_b0 , w_3661 );
and ( w_3660 ,  , w_3661 );
buf ( w_3659 , \1205_b1 );
not ( w_3659 , w_3662 );
not (  , w_3663 );
and ( w_3662 , w_3663 , \1205_b0 );
or ( \1207_b1 , \1196_b1 , w_3665 );
not ( w_3665 , w_3666 );
and ( \1207_b0 , \1196_b0 , w_3667 );
and ( w_3666 ,  , w_3667 );
buf ( w_3665 , \1206_b1 );
not ( w_3665 , w_3668 );
not (  , w_3669 );
and ( w_3668 , w_3669 , \1206_b0 );
or ( \1208_b1 , \b[7]_b1 , w_3671 );
not ( w_3671 , w_3672 );
and ( \1208_b0 , \b[7]_b0 , w_3673 );
and ( w_3672 ,  , w_3673 );
buf ( w_3671 , \d[7]_b1 );
not ( w_3671 , w_3674 );
not (  , w_3675 );
and ( w_3674 , w_3675 , \d[7]_b0 );
buf ( \1209_b1 , \1208_b1 );
not ( \1209_b1 , w_3676 );
not ( \1209_b0 , w_3677 );
and ( w_3676 , w_3677 , \1208_b0 );
or ( \1210_b1 , \b[7]_b1 , w_3679 );
not ( w_3679 , w_3680 );
and ( \1210_b0 , \b[7]_b0 , w_3681 );
and ( w_3680 ,  , w_3681 );
buf ( w_3679 , \d[7]_b1 );
not ( w_3679 , w_3682 );
not (  , w_3683 );
and ( w_3682 , w_3683 , \d[7]_b0 );
or ( \1211_b1 , \1209_b1 , w_3685 );
not ( w_3685 , w_3686 );
and ( \1211_b0 , \1209_b0 , w_3687 );
and ( w_3686 ,  , w_3687 );
buf ( w_3685 , \1210_b1 );
not ( w_3685 , w_3688 );
not (  , w_3689 );
and ( w_3688 , w_3689 , \1210_b0 );
or ( \1212_b1 , \1207_b1 , w_3690 );
xor ( \1212_b0 , \1207_b0 , w_3692 );
not ( w_3692 , w_3693 );
and ( w_3693 , w_3690 , w_3691 );
buf ( w_3690 , \1211_b1 );
not ( w_3690 , w_3694 );
not ( w_3691 , w_3695 );
and ( w_3694 , w_3695 , \1211_b0 );
buf ( \1213_b1 , \1212_b1 );
not ( \1213_b1 , w_3696 );
not ( \1213_b0 , w_3697 );
and ( w_3696 , w_3697 , \1212_b0 );
buf ( \1214_b1 , \447_b1 );
not ( \1214_b1 , w_3698 );
not ( \1214_b0 , w_3699 );
and ( w_3698 , w_3699 , \447_b0 );
buf ( \1215_b1 , \1214_b1 );
not ( \1215_b1 , w_3700 );
not ( \1215_b0 , w_3701 );
and ( w_3700 , w_3701 , \1214_b0 );
buf ( \1216_b1 , \457_b1 );
not ( \1216_b1 , w_3702 );
not ( \1216_b0 , w_3703 );
and ( w_3702 , w_3703 , \457_b0 );
or ( \1217_b1 , \1215_b1 , w_3704 );
or ( \1217_b0 , \1215_b0 , \1216_b0 );
not ( \1216_b0 , w_3705 );
and ( w_3705 , w_3704 , \1216_b1 );
or ( \1218_b1 , \1217_b1 , w_3707 );
not ( w_3707 , w_3708 );
and ( \1218_b0 , \1217_b0 , w_3709 );
and ( w_3708 ,  , w_3709 );
buf ( w_3707 , \528_b1 );
not ( w_3707 , w_3710 );
not (  , w_3711 );
and ( w_3710 , w_3711 , \528_b0 );
buf ( \1219_b1 , \524_b1 );
buf ( \1219_b0 , \524_b0 );
or ( \1220_b1 , \1218_b1 , w_3712 );
xor ( \1220_b0 , \1218_b0 , w_3714 );
not ( w_3714 , w_3715 );
and ( w_3715 , w_3712 , w_3713 );
buf ( w_3712 , \1219_b1 );
not ( w_3712 , w_3716 );
not ( w_3713 , w_3717 );
and ( w_3716 , w_3717 , \1219_b0 );
buf ( \1221_b1 , \1220_b1 );
not ( \1221_b1 , w_3718 );
not ( \1221_b0 , w_3719 );
and ( w_3718 , w_3719 , \1220_b0 );
or ( \1222_b1 , \1213_b1 , w_3720 );
or ( \1222_b0 , \1213_b0 , \1221_b0 );
not ( \1221_b0 , w_3721 );
and ( w_3721 , w_3720 , \1221_b1 );
buf ( \1223_b1 , \519_b1 );
buf ( \1223_b0 , \519_b0 );
buf ( \1224_b1 , \1223_b1 );
not ( \1224_b1 , w_3722 );
not ( \1224_b0 , w_3723 );
and ( w_3722 , w_3723 , \1223_b0 );
buf ( \1225_b1 , \472_b1 );
not ( \1225_b1 , w_3724 );
not ( \1225_b0 , w_3725 );
and ( w_3724 , w_3725 , \472_b0 );
buf ( \1226_b1 , \483_b1 );
not ( \1226_b1 , w_3726 );
not ( \1226_b0 , w_3727 );
and ( w_3726 , w_3727 , \483_b0 );
or ( \1227_b1 , \1225_b1 , w_3728 );
or ( \1227_b0 , \1225_b0 , \1226_b0 );
not ( \1226_b0 , w_3729 );
and ( w_3729 , w_3728 , \1226_b1 );
or ( \1228_b1 , \1227_b1 , w_3731 );
not ( w_3731 , w_3732 );
and ( \1228_b0 , \1227_b0 , w_3733 );
and ( w_3732 ,  , w_3733 );
buf ( w_3731 , \523_b1 );
not ( w_3731 , w_3734 );
not (  , w_3735 );
and ( w_3734 , w_3735 , \523_b0 );
buf ( \1229_b1 , \1228_b1 );
not ( \1229_b1 , w_3736 );
not ( \1229_b0 , w_3737 );
and ( w_3736 , w_3737 , \1228_b0 );
or ( \1230_b1 , \1224_b1 , w_3738 );
or ( \1230_b0 , \1224_b0 , \1229_b0 );
not ( \1229_b0 , w_3739 );
and ( w_3739 , w_3738 , \1229_b1 );
or ( \1231_b1 , \1228_b1 , w_3740 );
or ( \1231_b0 , \1228_b0 , \1223_b0 );
not ( \1223_b0 , w_3741 );
and ( w_3741 , w_3740 , \1223_b1 );
or ( \1232_b1 , \1230_b1 , w_3743 );
not ( w_3743 , w_3744 );
and ( \1232_b0 , \1230_b0 , w_3745 );
and ( w_3744 ,  , w_3745 );
buf ( w_3743 , \1231_b1 );
not ( w_3743 , w_3746 );
not (  , w_3747 );
and ( w_3746 , w_3747 , \1231_b0 );
or ( \1233_b1 , \a[2]_b1 , w_3749 );
not ( w_3749 , w_3750 );
and ( \1233_b0 , \a[2]_b0 , w_3751 );
and ( w_3750 ,  , w_3751 );
buf ( w_3749 , \c[2]_b1 );
not ( w_3749 , w_3752 );
not (  , w_3753 );
and ( w_3752 , w_3753 , \c[2]_b0 );
or ( \1234_b1 , \a[3]_b1 , w_3755 );
not ( w_3755 , w_3756 );
and ( \1234_b0 , \a[3]_b0 , w_3757 );
and ( w_3756 ,  , w_3757 );
buf ( w_3755 , \c[3]_b1 );
not ( w_3755 , w_3758 );
not (  , w_3759 );
and ( w_3758 , w_3759 , \c[3]_b0 );
or ( \1235_b1 , \1233_b1 , w_3761 );
not ( w_3761 , w_3762 );
and ( \1235_b0 , \1233_b0 , w_3763 );
and ( w_3762 ,  , w_3763 );
buf ( w_3761 , \1234_b1 );
not ( w_3761 , w_3764 );
not (  , w_3765 );
and ( w_3764 , w_3765 , \1234_b0 );
buf ( \1236_b1 , \1235_b1 );
not ( \1236_b1 , w_3766 );
not ( \1236_b0 , w_3767 );
and ( w_3766 , w_3767 , \1235_b0 );
or ( \1237_b1 , \a[0]_b1 , w_3769 );
not ( w_3769 , w_3770 );
and ( \1237_b0 , \a[0]_b0 , w_3771 );
and ( w_3770 ,  , w_3771 );
buf ( w_3769 , \c[0]_b1 );
not ( w_3769 , w_3772 );
not (  , w_3773 );
and ( w_3772 , w_3773 , \c[0]_b0 );
buf ( \1238_b1 , \1237_b1 );
not ( \1238_b1 , w_3774 );
not ( \1238_b0 , w_3775 );
and ( w_3774 , w_3775 , \1237_b0 );
buf ( \1239_b1 , \1238_b1 );
not ( \1239_b1 , w_3776 );
not ( \1239_b0 , w_3777 );
and ( w_3776 , w_3777 , \1238_b0 );
or ( \1240_b1 , \a[1]_b1 , w_3778 );
or ( \1240_b0 , \a[1]_b0 , \c[1]_b0 );
not ( \c[1]_b0 , w_3779 );
and ( w_3779 , w_3778 , \c[1]_b1 );
buf ( \1241_b1 , \1240_b1 );
not ( \1241_b1 , w_3780 );
not ( \1241_b0 , w_3781 );
and ( w_3780 , w_3781 , \1240_b0 );
or ( \1242_b1 , \1239_b1 , w_3782 );
or ( \1242_b0 , \1239_b0 , \1241_b0 );
not ( \1241_b0 , w_3783 );
and ( w_3783 , w_3782 , \1241_b1 );
or ( \1243_b1 , \a[1]_b1 , w_3785 );
not ( w_3785 , w_3786 );
and ( \1243_b0 , \a[1]_b0 , w_3787 );
and ( w_3786 ,  , w_3787 );
buf ( w_3785 , \c[1]_b1 );
not ( w_3785 , w_3788 );
not (  , w_3789 );
and ( w_3788 , w_3789 , \c[1]_b0 );
or ( \1244_b1 , \1242_b1 , w_3791 );
not ( w_3791 , w_3792 );
and ( \1244_b0 , \1242_b0 , w_3793 );
and ( w_3792 ,  , w_3793 );
buf ( w_3791 , \1243_b1 );
not ( w_3791 , w_3794 );
not (  , w_3795 );
and ( w_3794 , w_3795 , \1243_b0 );
buf ( \1245_b1 , \1244_b1 );
not ( \1245_b1 , w_3796 );
not ( \1245_b0 , w_3797 );
and ( w_3796 , w_3797 , \1244_b0 );
or ( \1246_b1 , \1236_b1 , w_3798 );
or ( \1246_b0 , \1236_b0 , \1245_b0 );
not ( \1245_b0 , w_3799 );
and ( w_3799 , w_3798 , \1245_b1 );
or ( \1247_b1 , \a[3]_b1 , w_3801 );
not ( w_3801 , w_3802 );
and ( \1247_b0 , \a[3]_b0 , w_3803 );
and ( w_3802 ,  , w_3803 );
buf ( w_3801 , \c[3]_b1 );
not ( w_3801 , w_3804 );
not (  , w_3805 );
and ( w_3804 , w_3805 , \c[3]_b0 );
buf ( \1248_b1 , \1247_b1 );
not ( \1248_b1 , w_3806 );
not ( \1248_b0 , w_3807 );
and ( w_3806 , w_3807 , \1247_b0 );
or ( \1249_b1 , \a[2]_b1 , w_3809 );
not ( w_3809 , w_3810 );
and ( \1249_b0 , \a[2]_b0 , w_3811 );
and ( w_3810 ,  , w_3811 );
buf ( w_3809 , \c[2]_b1 );
not ( w_3809 , w_3812 );
not (  , w_3813 );
and ( w_3812 , w_3813 , \c[2]_b0 );
or ( \1250_b1 , \1234_b1 , w_3815 );
not ( w_3815 , w_3816 );
and ( \1250_b0 , \1234_b0 , w_3817 );
and ( w_3816 ,  , w_3817 );
buf ( w_3815 , \1249_b1 );
not ( w_3815 , w_3818 );
not (  , w_3819 );
and ( w_3818 , w_3819 , \1249_b0 );
or ( \1251_b1 , \1248_b1 , w_3821 );
not ( w_3821 , w_3822 );
and ( \1251_b0 , \1248_b0 , w_3823 );
and ( w_3822 ,  , w_3823 );
buf ( w_3821 , \1250_b1 );
not ( w_3821 , w_3824 );
not (  , w_3825 );
and ( w_3824 , w_3825 , \1250_b0 );
or ( \1252_b1 , \1246_b1 , w_3827 );
not ( w_3827 , w_3828 );
and ( \1252_b0 , \1246_b0 , w_3829 );
and ( w_3828 ,  , w_3829 );
buf ( w_3827 , \1251_b1 );
not ( w_3827 , w_3830 );
not (  , w_3831 );
and ( w_3830 , w_3831 , \1251_b0 );
or ( \1253_b1 , \a[4]_b1 , w_3833 );
not ( w_3833 , w_3834 );
and ( \1253_b0 , \a[4]_b0 , w_3835 );
and ( w_3834 ,  , w_3835 );
buf ( w_3833 , \c[4]_b1 );
not ( w_3833 , w_3836 );
not (  , w_3837 );
and ( w_3836 , w_3837 , \c[4]_b0 );
buf ( \1254_b1 , \1253_b1 );
not ( \1254_b1 , w_3838 );
not ( \1254_b0 , w_3839 );
and ( w_3838 , w_3839 , \1253_b0 );
or ( \1255_b1 , \a[5]_b1 , w_3840 );
or ( \1255_b0 , \a[5]_b0 , \c[5]_b0 );
not ( \c[5]_b0 , w_3841 );
and ( w_3841 , w_3840 , \c[5]_b1 );
or ( \1256_b1 , \1254_b1 , w_3843 );
not ( w_3843 , w_3844 );
and ( \1256_b0 , \1254_b0 , w_3845 );
and ( w_3844 ,  , w_3845 );
buf ( w_3843 , \1255_b1 );
not ( w_3843 , w_3846 );
not (  , w_3847 );
and ( w_3846 , w_3847 , \1255_b0 );
or ( \1257_b1 , \a[6]_b1 , w_3849 );
not ( w_3849 , w_3850 );
and ( \1257_b0 , \a[6]_b0 , w_3851 );
and ( w_3850 ,  , w_3851 );
buf ( w_3849 , \c[6]_b1 );
not ( w_3849 , w_3852 );
not (  , w_3853 );
and ( w_3852 , w_3853 , \c[6]_b0 );
or ( \1258_b1 , \1256_b1 , w_3855 );
not ( w_3855 , w_3856 );
and ( \1258_b0 , \1256_b0 , w_3857 );
and ( w_3856 ,  , w_3857 );
buf ( w_3855 , \1257_b1 );
not ( w_3855 , w_3858 );
not (  , w_3859 );
and ( w_3858 , w_3859 , \1257_b0 );
or ( \1259_b1 , \1252_b1 , w_3861 );
not ( w_3861 , w_3862 );
and ( \1259_b0 , \1252_b0 , w_3863 );
and ( w_3862 ,  , w_3863 );
buf ( w_3861 , \1258_b1 );
not ( w_3861 , w_3864 );
not (  , w_3865 );
and ( w_3864 , w_3865 , \1258_b0 );
or ( \1260_b1 , \a[4]_b1 , w_3867 );
not ( w_3867 , w_3868 );
and ( \1260_b0 , \a[4]_b0 , w_3869 );
and ( w_3868 ,  , w_3869 );
buf ( w_3867 , \c[4]_b1 );
not ( w_3867 , w_3870 );
not (  , w_3871 );
and ( w_3870 , w_3871 , \c[4]_b0 );
buf ( \1261_b1 , \1260_b1 );
not ( \1261_b1 , w_3872 );
not ( \1261_b0 , w_3873 );
and ( w_3872 , w_3873 , \1260_b0 );
or ( \1262_b1 , \1255_b1 , w_3875 );
not ( w_3875 , w_3876 );
and ( \1262_b0 , \1255_b0 , w_3877 );
and ( w_3876 ,  , w_3877 );
buf ( w_3875 , \1261_b1 );
not ( w_3875 , w_3878 );
not (  , w_3879 );
and ( w_3878 , w_3879 , \1261_b0 );
or ( \1263_b1 , \a[5]_b1 , w_3881 );
not ( w_3881 , w_3882 );
and ( \1263_b0 , \a[5]_b0 , w_3883 );
and ( w_3882 ,  , w_3883 );
buf ( w_3881 , \c[5]_b1 );
not ( w_3881 , w_3884 );
not (  , w_3885 );
and ( w_3884 , w_3885 , \c[5]_b0 );
or ( \1264_b1 , \1262_b1 , w_3887 );
not ( w_3887 , w_3888 );
and ( \1264_b0 , \1262_b0 , w_3889 );
and ( w_3888 ,  , w_3889 );
buf ( w_3887 , \1263_b1 );
not ( w_3887 , w_3890 );
not (  , w_3891 );
and ( w_3890 , w_3891 , \1263_b0 );
buf ( \1265_b1 , \1257_b1 );
not ( \1265_b1 , w_3892 );
not ( \1265_b0 , w_3893 );
and ( w_3892 , w_3893 , \1257_b0 );
or ( \1266_b1 , \1264_b1 , \1265_b1 );
not ( \1265_b1 , w_3894 );
and ( \1266_b0 , \1264_b0 , w_3895 );
and ( w_3894 , w_3895 , \1265_b0 );
or ( \1267_b1 , \a[6]_b1 , w_3897 );
not ( w_3897 , w_3898 );
and ( \1267_b0 , \a[6]_b0 , w_3899 );
and ( w_3898 ,  , w_3899 );
buf ( w_3897 , \c[6]_b1 );
not ( w_3897 , w_3900 );
not (  , w_3901 );
and ( w_3900 , w_3901 , \c[6]_b0 );
buf ( \1268_b1 , \1267_b1 );
not ( \1268_b1 , w_3902 );
not ( \1268_b0 , w_3903 );
and ( w_3902 , w_3903 , \1267_b0 );
or ( \1269_b1 , \1266_b1 , w_3905 );
not ( w_3905 , w_3906 );
and ( \1269_b0 , \1266_b0 , w_3907 );
and ( w_3906 ,  , w_3907 );
buf ( w_3905 , \1268_b1 );
not ( w_3905 , w_3908 );
not (  , w_3909 );
and ( w_3908 , w_3909 , \1268_b0 );
or ( \1270_b1 , \1259_b1 , w_3911 );
not ( w_3911 , w_3912 );
and ( \1270_b0 , \1259_b0 , w_3913 );
and ( w_3912 ,  , w_3913 );
buf ( w_3911 , \1269_b1 );
not ( w_3911 , w_3914 );
not (  , w_3915 );
and ( w_3914 , w_3915 , \1269_b0 );
or ( \1271_b1 , \a[7]_b1 , w_3917 );
not ( w_3917 , w_3918 );
and ( \1271_b0 , \a[7]_b0 , w_3919 );
and ( w_3918 ,  , w_3919 );
buf ( w_3917 , \c[7]_b1 );
not ( w_3917 , w_3920 );
not (  , w_3921 );
and ( w_3920 , w_3921 , \c[7]_b0 );
buf ( \1272_b1 , \1271_b1 );
not ( \1272_b1 , w_3922 );
not ( \1272_b0 , w_3923 );
and ( w_3922 , w_3923 , \1271_b0 );
or ( \1273_b1 , \a[7]_b1 , w_3925 );
not ( w_3925 , w_3926 );
and ( \1273_b0 , \a[7]_b0 , w_3927 );
and ( w_3926 ,  , w_3927 );
buf ( w_3925 , \c[7]_b1 );
not ( w_3925 , w_3928 );
not (  , w_3929 );
and ( w_3928 , w_3929 , \c[7]_b0 );
or ( \1274_b1 , \1272_b1 , w_3931 );
not ( w_3931 , w_3932 );
and ( \1274_b0 , \1272_b0 , w_3933 );
and ( w_3932 ,  , w_3933 );
buf ( w_3931 , \1273_b1 );
not ( w_3931 , w_3934 );
not (  , w_3935 );
and ( w_3934 , w_3935 , \1273_b0 );
or ( \1275_b1 , \1270_b1 , w_3936 );
xor ( \1275_b0 , \1270_b0 , w_3938 );
not ( w_3938 , w_3939 );
and ( w_3939 , w_3936 , w_3937 );
buf ( w_3936 , \1274_b1 );
not ( w_3936 , w_3940 );
not ( w_3937 , w_3941 );
and ( w_3940 , w_3941 , \1274_b0 );
or ( \1276_b1 , \1232_b1 , \1275_b1 );
not ( \1275_b1 , w_3942 );
and ( \1276_b0 , \1232_b0 , w_3943 );
and ( w_3942 , w_3943 , \1275_b0 );
buf ( \1277_b1 , \d[7]_b1 );
not ( \1277_b1 , w_3944 );
not ( \1277_b0 , w_3945 );
and ( w_3944 , w_3945 , \d[7]_b0 );
or ( \1278_b1 , \518_b1 , w_3947 );
not ( w_3947 , w_3948 );
and ( \1278_b0 , \518_b0 , w_3949 );
and ( w_3948 ,  , w_3949 );
buf ( w_3947 , \498_b1 );
not ( w_3947 , w_3950 );
not (  , w_3951 );
and ( w_3950 , w_3951 , \498_b0 );
buf ( \1279_b1 , \515_b1 );
buf ( \1279_b0 , \515_b0 );
or ( \1280_b1 , \1278_b1 , w_3952 );
xor ( \1280_b0 , \1278_b0 , w_3954 );
not ( w_3954 , w_3955 );
and ( w_3955 , w_3952 , w_3953 );
buf ( w_3952 , \1279_b1 );
not ( w_3952 , w_3956 );
not ( w_3953 , w_3957 );
and ( w_3956 , w_3957 , \1279_b0 );
buf ( \1281_b1 , \1280_b1 );
not ( \1281_b1 , w_3958 );
not ( \1281_b0 , w_3959 );
and ( w_3958 , w_3959 , \1280_b0 );
buf ( \1282_b1 , \1281_b1 );
not ( \1282_b1 , w_3960 );
not ( \1282_b0 , w_3961 );
and ( w_3960 , w_3961 , \1281_b0 );
buf ( \1283_b1 , \1282_b1 );
not ( \1283_b1 , w_3962 );
not ( \1283_b0 , w_3963 );
and ( w_3962 , w_3963 , \1282_b0 );
or ( \1284_b1 , \1277_b1 , w_3964 );
or ( \1284_b0 , \1277_b0 , \1283_b0 );
not ( \1283_b0 , w_3965 );
and ( w_3965 , w_3964 , \1283_b1 );
buf ( \1285_b1 , \506_b1 );
not ( \1285_b1 , w_3966 );
not ( \1285_b0 , w_3967 );
and ( w_3966 , w_3967 , \506_b0 );
or ( \1286_b1 , \1285_b1 , w_3969 );
not ( w_3969 , w_3970 );
and ( \1286_b0 , \1285_b0 , w_3971 );
and ( w_3970 ,  , w_3971 );
buf ( w_3969 , \514_b1 );
not ( w_3969 , w_3972 );
not (  , w_3973 );
and ( w_3972 , w_3973 , \514_b0 );
or ( \1287_b1 , \1286_b1 , \512_b1 );
xor ( \1287_b0 , \1286_b0 , w_3974 );
not ( w_3974 , w_3975 );
and ( w_3975 , \512_b1 , \512_b0 );
or ( \1288_b1 , \1287_b1 , \c[7]_b1 );
not ( \c[7]_b1 , w_3976 );
and ( \1288_b0 , \1287_b0 , w_3977 );
and ( w_3976 , w_3977 , \c[7]_b0 );
buf ( \1289_b1 , \b[0]_b1 );
not ( \1289_b1 , w_3978 );
not ( \1289_b0 , w_3979 );
and ( w_3978 , w_3979 , \b[0]_b0 );
buf ( \1290_b1 , \499_b1 );
not ( \1290_b1 , w_3980 );
not ( \1290_b0 , w_3981 );
and ( w_3980 , w_3981 , \499_b0 );
or ( \1291_b1 , \1289_b1 , w_3982 );
or ( \1291_b0 , \1289_b0 , \1290_b0 );
not ( \1290_b0 , w_3983 );
and ( w_3983 , w_3982 , \1290_b1 );
or ( \1292_b1 , \1291_b1 , w_3985 );
not ( w_3985 , w_3986 );
and ( \1292_b0 , \1291_b0 , w_3987 );
and ( w_3986 ,  , w_3987 );
buf ( w_3985 , \508_b1 );
not ( w_3985 , w_3988 );
not (  , w_3989 );
and ( w_3988 , w_3989 , \508_b0 );
or ( \1293_b1 , \512_b1 , \1292_b1 );
not ( \1292_b1 , w_3990 );
and ( \1293_b0 , \512_b0 , w_3991 );
and ( w_3990 , w_3991 , \1292_b0 );
or ( \1294_b1 , \1293_b1 , \b[7]_b1 );
not ( \b[7]_b1 , w_3992 );
and ( \1294_b0 , \1293_b0 , w_3993 );
and ( w_3992 , w_3993 , \b[7]_b0 );
or ( \1295_b1 , \1288_b1 , w_3995 );
not ( w_3995 , w_3996 );
and ( \1295_b0 , \1288_b0 , w_3997 );
and ( w_3996 ,  , w_3997 );
buf ( w_3995 , \1294_b1 );
not ( w_3995 , w_3998 );
not (  , w_3999 );
and ( w_3998 , w_3999 , \1294_b0 );
or ( \1296_b1 , \1284_b1 , w_4001 );
not ( w_4001 , w_4002 );
and ( \1296_b0 , \1284_b0 , w_4003 );
and ( w_4002 ,  , w_4003 );
buf ( w_4001 , \1295_b1 );
not ( w_4001 , w_4004 );
not (  , w_4005 );
and ( w_4004 , w_4005 , \1295_b0 );
or ( \1297_b1 , \1276_b1 , w_4007 );
not ( w_4007 , w_4008 );
and ( \1297_b0 , \1276_b0 , w_4009 );
and ( w_4008 ,  , w_4009 );
buf ( w_4007 , \1296_b1 );
not ( w_4007 , w_4010 );
not (  , w_4011 );
and ( w_4010 , w_4011 , \1296_b0 );
or ( \1298_b1 , \1222_b1 , w_4013 );
not ( w_4013 , w_4014 );
and ( \1298_b0 , \1222_b0 , w_4015 );
and ( w_4014 ,  , w_4015 );
buf ( w_4013 , \1297_b1 );
not ( w_4013 , w_4016 );
not (  , w_4017 );
and ( w_4016 , w_4017 , \1297_b0 );
or ( \1299_b1 , \1169_b1 , w_4019 );
not ( w_4019 , w_4020 );
and ( \1299_b0 , \1169_b0 , w_4021 );
and ( w_4020 ,  , w_4021 );
buf ( w_4019 , \1298_b1 );
not ( w_4019 , w_4022 );
not (  , w_4023 );
and ( w_4022 , w_4023 , \1298_b0 );
or ( \1300_b1 , \927_b1 , w_4025 );
not ( w_4025 , w_4026 );
and ( \1300_b0 , \927_b0 , w_4027 );
and ( w_4026 ,  , w_4027 );
buf ( w_4025 , \1299_b1 );
not ( w_4025 , w_4028 );
not (  , w_4029 );
and ( w_4028 , w_4029 , \1299_b0 );
or ( \1301_b1 , \919_b1 , w_4031 );
not ( w_4031 , w_4032 );
and ( \1301_b0 , \919_b0 , w_4033 );
and ( w_4032 ,  , w_4033 );
buf ( w_4031 , \1300_b1 );
not ( w_4031 , w_4034 );
not (  , w_4035 );
and ( w_4034 , w_4035 , \1300_b0 );
or ( \1302_b1 , \674_b1 , w_4037 );
not ( w_4037 , w_4038 );
and ( \1302_b0 , \674_b0 , w_4039 );
and ( w_4038 ,  , w_4039 );
buf ( w_4037 , \1301_b1 );
not ( w_4037 , w_4040 );
not (  , w_4041 );
and ( w_4040 , w_4041 , \1301_b0 );
buf ( \1303_b1 , \1302_b1 );
not ( \1303_b1 , w_4042 );
not ( \1303_b0 , w_4043 );
and ( w_4042 , w_4043 , \1302_b0 );
or ( \1304_b1 , \551_b1 , w_4045 );
not ( w_4045 , w_4046 );
and ( \1304_b0 , \551_b0 , w_4047 );
and ( w_4046 ,  , w_4047 );
buf ( w_4045 , \328_b1 );
not ( w_4045 , w_4048 );
not (  , w_4049 );
and ( w_4048 , w_4049 , \328_b0 );
buf ( \1305_b1 , \1304_b1 );
not ( \1305_b1 , w_4050 );
not ( \1305_b0 , w_4051 );
and ( w_4050 , w_4051 , \1304_b0 );
or ( \1306_b1 , \1305_b1 , w_4053 );
not ( w_4053 , w_4054 );
and ( \1306_b0 , \1305_b0 , w_4055 );
and ( w_4054 ,  , w_4055 );
buf ( w_4053 , \541_b1 );
not ( w_4053 , w_4056 );
not (  , w_4057 );
and ( w_4056 , w_4057 , \541_b0 );
buf ( \1307_b1 , \544_b1 );
not ( \1307_b1 , w_4058 );
not ( \1307_b0 , w_4059 );
and ( w_4058 , w_4059 , \544_b0 );
buf ( \1308_b1 , \283_b1 );
not ( \1308_b1 , w_4060 );
not ( \1308_b0 , w_4061 );
and ( w_4060 , w_4061 , \283_b0 );
or ( \1309_b1 , \1307_b1 , w_4063 );
not ( w_4063 , w_4064 );
and ( \1309_b0 , \1307_b0 , w_4065 );
and ( w_4064 ,  , w_4065 );
buf ( w_4063 , \1308_b1 );
not ( w_4063 , w_4066 );
not (  , w_4067 );
and ( w_4066 , w_4067 , \1308_b0 );
or ( \1310_b1 , \1309_b1 , w_4069 );
not ( w_4069 , w_4070 );
and ( \1310_b0 , \1309_b0 , w_4071 );
and ( w_4070 ,  , w_4071 );
buf ( w_4069 , \284_b1 );
not ( w_4069 , w_4072 );
not (  , w_4073 );
and ( w_4072 , w_4073 , \284_b0 );
or ( \1311_b1 , \1306_b1 , \1310_b1 );
not ( \1310_b1 , w_4074 );
and ( \1311_b0 , \1306_b0 , w_4075 );
and ( w_4074 , w_4075 , \1310_b0 );
buf ( \1312_b1 , \1306_b1 );
not ( \1312_b1 , w_4076 );
not ( \1312_b0 , w_4077 );
and ( w_4076 , w_4077 , \1306_b0 );
buf ( \1313_b1 , \1310_b1 );
not ( \1313_b1 , w_4078 );
not ( \1313_b0 , w_4079 );
and ( w_4078 , w_4079 , \1310_b0 );
or ( \1314_b1 , \1312_b1 , \1313_b1 );
not ( \1313_b1 , w_4080 );
and ( \1314_b0 , \1312_b0 , w_4081 );
and ( w_4080 , w_4081 , \1313_b0 );
or ( \1315_b1 , \1311_b1 , w_4083 );
not ( w_4083 , w_4084 );
and ( \1315_b0 , \1311_b0 , w_4085 );
and ( w_4084 ,  , w_4085 );
buf ( w_4083 , \1314_b1 );
not ( w_4083 , w_4086 );
not (  , w_4087 );
and ( w_4086 , w_4087 , \1314_b0 );
buf ( \1316_b1 , \1315_b1 );
buf ( \1316_b0 , \1315_b0 );
or ( \1317_b1 , \b[7]_b1 , \c[7]_b1 );
not ( \c[7]_b1 , w_4088 );
and ( \1317_b0 , \b[7]_b0 , w_4089 );
and ( w_4088 , w_4089 , \c[7]_b0 );
or ( \1318_b1 , \1316_b1 , w_4091 );
not ( w_4091 , w_4092 );
and ( \1318_b0 , \1316_b0 , w_4093 );
and ( w_4092 ,  , w_4093 );
buf ( w_4091 , \1317_b1 );
not ( w_4091 , w_4094 );
not (  , w_4095 );
and ( w_4094 , w_4095 , \1317_b0 );
buf ( \1319_b1 , \1316_b1 );
not ( \1319_b1 , w_4096 );
not ( \1319_b0 , w_4097 );
and ( w_4096 , w_4097 , \1316_b0 );
buf ( \1320_b1 , \924_b1 );
not ( \1320_b1 , w_4098 );
not ( \1320_b0 , w_4099 );
and ( w_4098 , w_4099 , \924_b0 );
buf ( \1321_b1 , \1320_b1 );
not ( \1321_b1 , w_4100 );
not ( \1321_b0 , w_4101 );
and ( w_4100 , w_4101 , \1320_b0 );
buf ( \1322_b1 , \1232_b1 );
not ( \1322_b1 , w_4102 );
not ( \1322_b0 , w_4103 );
and ( w_4102 , w_4103 , \1232_b0 );
buf ( \1323_b1 , \1287_b1 );
not ( \1323_b1 , w_4104 );
not ( \1323_b0 , w_4105 );
and ( w_4104 , w_4105 , \1287_b0 );
buf ( \1324_b1 , \1293_b1 );
not ( \1324_b1 , w_4106 );
not ( \1324_b0 , w_4107 );
and ( w_4106 , w_4107 , \1293_b0 );
or ( \1325_b1 , \1323_b1 , w_4109 );
not ( w_4109 , w_4110 );
and ( \1325_b0 , \1323_b0 , w_4111 );
and ( w_4110 ,  , w_4111 );
buf ( w_4109 , \1324_b1 );
not ( w_4109 , w_4112 );
not (  , w_4113 );
and ( w_4112 , w_4113 , \1324_b0 );
or ( \1326_b1 , \1280_b1 , w_4115 );
not ( w_4115 , w_4116 );
and ( \1326_b0 , \1280_b0 , w_4117 );
and ( w_4116 ,  , w_4117 );
buf ( w_4115 , \1325_b1 );
not ( w_4115 , w_4118 );
not (  , w_4119 );
and ( w_4118 , w_4119 , \1325_b0 );
or ( \1327_b1 , \1322_b1 , w_4121 );
not ( w_4121 , w_4122 );
and ( \1327_b0 , \1322_b0 , w_4123 );
and ( w_4122 ,  , w_4123 );
buf ( w_4121 , \1326_b1 );
not ( w_4121 , w_4124 );
not (  , w_4125 );
and ( w_4124 , w_4125 , \1326_b0 );
or ( \1328_b1 , \1220_b1 , w_4127 );
not ( w_4127 , w_4128 );
and ( \1328_b0 , \1220_b0 , w_4129 );
and ( w_4128 ,  , w_4129 );
buf ( w_4127 , \1327_b1 );
not ( w_4127 , w_4130 );
not (  , w_4131 );
and ( w_4130 , w_4131 , \1327_b0 );
or ( \1329_b1 , \1167_b1 , w_4133 );
not ( w_4133 , w_4134 );
and ( \1329_b0 , \1167_b0 , w_4135 );
and ( w_4134 ,  , w_4135 );
buf ( w_4133 , \1328_b1 );
not ( w_4133 , w_4136 );
not (  , w_4137 );
and ( w_4136 , w_4137 , \1328_b0 );
or ( \1330_b1 , \916_b1 , w_4139 );
not ( w_4139 , w_4140 );
and ( \1330_b0 , \916_b0 , w_4141 );
and ( w_4140 ,  , w_4141 );
buf ( w_4139 , \1329_b1 );
not ( w_4139 , w_4142 );
not (  , w_4143 );
and ( w_4142 , w_4143 , \1329_b0 );
or ( \1331_b1 , \1321_b1 , w_4145 );
not ( w_4145 , w_4146 );
and ( \1331_b0 , \1321_b0 , w_4147 );
and ( w_4146 ,  , w_4147 );
buf ( w_4145 , \1330_b1 );
not ( w_4145 , w_4148 );
not (  , w_4149 );
and ( w_4148 , w_4149 , \1330_b0 );
or ( \1332_b1 , \1331_b1 , w_4151 );
not ( w_4151 , w_4152 );
and ( \1332_b0 , \1331_b0 , w_4153 );
and ( w_4152 ,  , w_4153 );
buf ( w_4151 , \648_b1 );
not ( w_4151 , w_4154 );
not (  , w_4155 );
and ( w_4154 , w_4155 , \648_b0 );
or ( \1333_b1 , \1319_b1 , w_4157 );
not ( w_4157 , w_4158 );
and ( \1333_b0 , \1319_b0 , w_4159 );
and ( w_4158 ,  , w_4159 );
buf ( w_4157 , \1332_b1 );
not ( w_4157 , w_4160 );
not (  , w_4161 );
and ( w_4160 , w_4161 , \1332_b0 );
or ( \1335_b1 , \646_b1 , w_4163 );
not ( w_4163 , w_4164 );
and ( \1335_b0 , \646_b0 , w_4165 );
and ( w_4164 ,  , w_4165 );
buf ( w_4163 , \1334_b1 );
not ( w_4163 , w_4166 );
not (  , w_4167 );
and ( w_4166 , w_4167 , \1334_b0 );
buf ( \1336_b1 , \1335_b1 );
not ( \1336_b1 , w_4168 );
not ( \1336_b0 , w_4169 );
and ( w_4168 , w_4169 , \1335_b0 );
buf ( \1337_b1 , \a[1]_b1 );
not ( \1337_b1 , w_4170 );
not ( \1337_b0 , w_4171 );
and ( w_4170 , w_4171 , \a[1]_b0 );
or ( \1338_b1 , \1316_b1 , w_4173 );
not ( w_4173 , w_4174 );
and ( \1338_b0 , \1316_b0 , w_4175 );
and ( w_4174 ,  , w_4175 );
buf ( w_4173 , \1331_b1 );
not ( w_4173 , w_4176 );
not (  , w_4177 );
and ( w_4176 , w_4177 , \1331_b0 );
buf ( \1339_b1 , \1338_b1 );
not ( \1339_b1 , w_4178 );
not ( \1339_b0 , w_4179 );
and ( w_4178 , w_4179 , \1338_b0 );
or ( \1340_b1 , \1337_b1 , w_4180 );
or ( \1340_b0 , \1337_b0 , \1339_b0 );
not ( \1339_b0 , w_4181 );
and ( w_4181 , w_4180 , \1339_b1 );
buf ( \1341_b1 , \643_b1 );
not ( \1341_b1 , w_4182 );
not ( \1341_b0 , w_4183 );
and ( w_4182 , w_4183 , \643_b0 );
buf ( \1342_b1 , \1341_b1 );
not ( \1342_b1 , w_4184 );
not ( \1342_b0 , w_4185 );
and ( w_4184 , w_4185 , \1341_b0 );
or ( \1343_b1 , \a[1]_b1 , w_4186 );
or ( \1343_b0 , \a[1]_b0 , \d[1]_b0 );
not ( \d[1]_b0 , w_4187 );
and ( w_4187 , w_4186 , \d[1]_b1 );
or ( \1344_b1 , \1342_b1 , \1343_b1 );
not ( \1343_b1 , w_4188 );
and ( \1344_b0 , \1342_b0 , w_4189 );
and ( w_4188 , w_4189 , \1343_b0 );
or ( \1345_b1 , \b[1]_b1 , \c[1]_b1 );
not ( \c[1]_b1 , w_4190 );
and ( \1345_b0 , \b[1]_b0 , w_4191 );
and ( w_4190 , w_4191 , \c[1]_b0 );
buf ( \1346_b1 , \1345_b1 );
not ( \1346_b1 , w_4192 );
not ( \1346_b0 , w_4193 );
and ( w_4192 , w_4193 , \1345_b0 );
buf ( \1347_b1 , \1316_b1 );
not ( \1347_b1 , w_4194 );
not ( \1347_b0 , w_4195 );
and ( w_4194 , w_4195 , \1316_b0 );
or ( \1348_b1 , \1346_b1 , w_4196 );
or ( \1348_b0 , \1346_b0 , \1347_b0 );
not ( \1347_b0 , w_4197 );
and ( w_4197 , w_4196 , \1347_b1 );
or ( \1349_b1 , \a[1]_b1 , w_4198 );
or ( \1349_b0 , \a[1]_b0 , \b[1]_b0 );
not ( \b[1]_b0 , w_4199 );
and ( w_4199 , w_4198 , \b[1]_b1 );
buf ( \1350_b1 , \671_b1 );
not ( \1350_b1 , w_4200 );
not ( \1350_b0 , w_4201 );
and ( w_4200 , w_4201 , \671_b0 );
buf ( \1351_b1 , \1350_b1 );
not ( \1351_b1 , w_4202 );
not ( \1351_b0 , w_4203 );
and ( w_4202 , w_4203 , \1350_b0 );
or ( \1352_b1 , \1349_b1 , \1351_b1 );
not ( \1351_b1 , w_4204 );
and ( \1352_b0 , \1349_b0 , w_4205 );
and ( w_4204 , w_4205 , \1351_b0 );
buf ( \1353_b1 , \1167_b1 );
not ( \1353_b1 , w_4206 );
not ( \1353_b0 , w_4207 );
and ( w_4206 , w_4207 , \1167_b0 );
or ( \1354_b1 , \1043_b1 , w_4208 );
or ( \1354_b0 , \1043_b0 , \1045_b0 );
not ( \1045_b0 , w_4209 );
and ( w_4209 , w_4208 , \1045_b1 );
or ( \1355_b1 , \1354_b1 , \1046_b1 );
not ( \1046_b1 , w_4210 );
and ( \1355_b0 , \1354_b0 , w_4211 );
and ( w_4210 , w_4211 , \1046_b0 );
or ( \1356_b1 , \1353_b1 , \1355_b1 );
not ( \1355_b1 , w_4212 );
and ( \1356_b0 , \1353_b0 , w_4213 );
and ( w_4212 , w_4213 , \1355_b0 );
buf ( \1357_b1 , \1175_b1 );
not ( \1357_b1 , w_4214 );
not ( \1357_b0 , w_4215 );
and ( w_4214 , w_4215 , \1175_b0 );
or ( \1358_b1 , \1177_b1 , w_4217 );
not ( w_4217 , w_4218 );
and ( \1358_b0 , \1177_b0 , w_4219 );
and ( w_4218 ,  , w_4219 );
buf ( w_4217 , \1180_b1 );
not ( w_4217 , w_4220 );
not (  , w_4221 );
and ( w_4220 , w_4221 , \1180_b0 );
buf ( \1359_b1 , \1358_b1 );
not ( \1359_b1 , w_4222 );
not ( \1359_b0 , w_4223 );
and ( w_4222 , w_4223 , \1358_b0 );
or ( \1360_b1 , \1357_b1 , w_4224 );
or ( \1360_b0 , \1357_b0 , \1359_b0 );
not ( \1359_b0 , w_4225 );
and ( w_4225 , w_4224 , \1359_b1 );
or ( \1361_b1 , \1358_b1 , w_4226 );
or ( \1361_b0 , \1358_b0 , \1175_b0 );
not ( \1175_b0 , w_4227 );
and ( w_4227 , w_4226 , \1175_b1 );
or ( \1362_b1 , \1360_b1 , w_4229 );
not ( w_4229 , w_4230 );
and ( \1362_b0 , \1360_b0 , w_4231 );
and ( w_4230 ,  , w_4231 );
buf ( w_4229 , \1361_b1 );
not ( w_4229 , w_4232 );
not (  , w_4233 );
and ( w_4232 , w_4233 , \1361_b0 );
buf ( \1363_b1 , \1362_b1 );
not ( \1363_b1 , w_4234 );
not ( \1363_b0 , w_4235 );
and ( w_4234 , w_4235 , \1362_b0 );
buf ( \1364_b1 , \1220_b1 );
not ( \1364_b1 , w_4236 );
not ( \1364_b0 , w_4237 );
and ( w_4236 , w_4237 , \1220_b0 );
or ( \1365_b1 , \1363_b1 , w_4238 );
or ( \1365_b0 , \1363_b0 , \1364_b0 );
not ( \1364_b0 , w_4239 );
and ( w_4239 , w_4238 , \1364_b1 );
buf ( \1366_b1 , \1238_b1 );
not ( \1366_b1 , w_4240 );
not ( \1366_b0 , w_4241 );
and ( w_4240 , w_4241 , \1238_b0 );
or ( \1367_b1 , \1240_b1 , w_4243 );
not ( w_4243 , w_4244 );
and ( \1367_b0 , \1240_b0 , w_4245 );
and ( w_4244 ,  , w_4245 );
buf ( w_4243 , \1243_b1 );
not ( w_4243 , w_4246 );
not (  , w_4247 );
and ( w_4246 , w_4247 , \1243_b0 );
buf ( \1368_b1 , \1367_b1 );
not ( \1368_b1 , w_4248 );
not ( \1368_b0 , w_4249 );
and ( w_4248 , w_4249 , \1367_b0 );
or ( \1369_b1 , \1366_b1 , w_4250 );
or ( \1369_b0 , \1366_b0 , \1368_b0 );
not ( \1368_b0 , w_4251 );
and ( w_4251 , w_4250 , \1368_b1 );
or ( \1370_b1 , \1367_b1 , w_4252 );
or ( \1370_b0 , \1367_b0 , \1238_b0 );
not ( \1238_b0 , w_4253 );
and ( w_4253 , w_4252 , \1238_b1 );
or ( \1371_b1 , \1369_b1 , w_4255 );
not ( w_4255 , w_4256 );
and ( \1371_b0 , \1369_b0 , w_4257 );
and ( w_4256 ,  , w_4257 );
buf ( w_4255 , \1370_b1 );
not ( w_4255 , w_4258 );
not (  , w_4259 );
and ( w_4258 , w_4259 , \1370_b0 );
or ( \1372_b1 , \1232_b1 , \1371_b1 );
not ( \1371_b1 , w_4260 );
and ( \1372_b0 , \1232_b0 , w_4261 );
and ( w_4260 , w_4261 , \1371_b0 );
buf ( \1373_b1 , \d[1]_b1 );
not ( \1373_b1 , w_4262 );
not ( \1373_b0 , w_4263 );
and ( w_4262 , w_4263 , \d[1]_b0 );
buf ( \1374_b1 , \1282_b1 );
not ( \1374_b1 , w_4264 );
not ( \1374_b0 , w_4265 );
and ( w_4264 , w_4265 , \1282_b0 );
or ( \1375_b1 , \1373_b1 , w_4266 );
or ( \1375_b0 , \1373_b0 , \1374_b0 );
not ( \1374_b0 , w_4267 );
and ( w_4267 , w_4266 , \1374_b1 );
or ( \1376_b1 , \1287_b1 , \c[1]_b1 );
not ( \c[1]_b1 , w_4268 );
and ( \1376_b0 , \1287_b0 , w_4269 );
and ( w_4268 , w_4269 , \c[1]_b0 );
or ( \1377_b1 , \1293_b1 , \b[1]_b1 );
not ( \b[1]_b1 , w_4270 );
and ( \1377_b0 , \1293_b0 , w_4271 );
and ( w_4270 , w_4271 , \b[1]_b0 );
or ( \1378_b1 , \1376_b1 , w_4273 );
not ( w_4273 , w_4274 );
and ( \1378_b0 , \1376_b0 , w_4275 );
and ( w_4274 ,  , w_4275 );
buf ( w_4273 , \1377_b1 );
not ( w_4273 , w_4276 );
not (  , w_4277 );
and ( w_4276 , w_4277 , \1377_b0 );
or ( \1379_b1 , \1375_b1 , w_4279 );
not ( w_4279 , w_4280 );
and ( \1379_b0 , \1375_b0 , w_4281 );
and ( w_4280 ,  , w_4281 );
buf ( w_4279 , \1378_b1 );
not ( w_4279 , w_4282 );
not (  , w_4283 );
and ( w_4282 , w_4283 , \1378_b0 );
or ( \1380_b1 , \1372_b1 , w_4285 );
not ( w_4285 , w_4286 );
and ( \1380_b0 , \1372_b0 , w_4287 );
and ( w_4286 ,  , w_4287 );
buf ( w_4285 , \1379_b1 );
not ( w_4285 , w_4288 );
not (  , w_4289 );
and ( w_4288 , w_4289 , \1379_b0 );
or ( \1381_b1 , \1365_b1 , w_4291 );
not ( w_4291 , w_4292 );
and ( \1381_b0 , \1365_b0 , w_4293 );
and ( w_4292 ,  , w_4293 );
buf ( w_4291 , \1380_b1 );
not ( w_4291 , w_4294 );
not (  , w_4295 );
and ( w_4294 , w_4295 , \1380_b0 );
or ( \1382_b1 , \1356_b1 , w_4297 );
not ( w_4297 , w_4298 );
and ( \1382_b0 , \1356_b0 , w_4299 );
and ( w_4298 ,  , w_4299 );
buf ( w_4297 , \1381_b1 );
not ( w_4297 , w_4300 );
not (  , w_4301 );
and ( w_4300 , w_4301 , \1381_b0 );
buf ( \1383_b1 , \924_b1 );
not ( \1383_b1 , w_4302 );
not ( \1383_b0 , w_4303 );
and ( w_4302 , w_4303 , \924_b0 );
or ( \1384_b1 , \c[1]_b1 , \d[1]_b1 );
xor ( \1384_b0 , \c[1]_b0 , w_4304 );
not ( w_4304 , w_4305 );
and ( w_4305 , \d[1]_b1 , \d[1]_b0 );
or ( \1385_b1 , \1383_b1 , w_4307 );
not ( w_4307 , w_4308 );
and ( \1385_b0 , \1383_b0 , w_4309 );
and ( w_4308 ,  , w_4309 );
buf ( w_4307 , \1384_b1 );
not ( w_4307 , w_4310 );
not (  , w_4311 );
and ( w_4310 , w_4311 , \1384_b0 );
buf ( \1386_b1 , \860_b1 );
not ( \1386_b1 , w_4312 );
not ( \1386_b0 , w_4313 );
and ( w_4312 , w_4313 , \860_b0 );
or ( \1387_b1 , \1386_b1 , \853_b1 );
not ( \853_b1 , w_4314 );
and ( \1387_b0 , \1386_b0 , w_4315 );
and ( w_4314 , w_4315 , \853_b0 );
buf ( \1388_b1 , \861_b1 );
not ( \1388_b1 , w_4316 );
not ( \1388_b0 , w_4317 );
and ( w_4316 , w_4317 , \861_b0 );
or ( \1389_b1 , \1387_b1 , w_4319 );
not ( w_4319 , w_4320 );
and ( \1389_b0 , \1387_b0 , w_4321 );
and ( w_4320 ,  , w_4321 );
buf ( w_4319 , \1388_b1 );
not ( w_4319 , w_4322 );
not (  , w_4323 );
and ( w_4322 , w_4323 , \1388_b0 );
or ( \1390_b1 , \916_b1 , w_4325 );
not ( w_4325 , w_4326 );
and ( \1390_b0 , \916_b0 , w_4327 );
and ( w_4326 ,  , w_4327 );
buf ( w_4325 , \1389_b1 );
not ( w_4325 , w_4328 );
not (  , w_4329 );
and ( w_4328 , w_4329 , \1389_b0 );
or ( \1392_b1 , \1352_b1 , w_4331 );
not ( w_4331 , w_4332 );
and ( \1392_b0 , \1352_b0 , w_4333 );
and ( w_4332 ,  , w_4333 );
buf ( w_4331 , \1391_b1 );
not ( w_4331 , w_4334 );
not (  , w_4335 );
and ( w_4334 , w_4335 , \1391_b0 );
or ( \1393_b1 , \1348_b1 , w_4337 );
not ( w_4337 , w_4338 );
and ( \1393_b0 , \1348_b0 , w_4339 );
and ( w_4338 ,  , w_4339 );
buf ( w_4337 , \1392_b1 );
not ( w_4337 , w_4340 );
not (  , w_4341 );
and ( w_4340 , w_4341 , \1392_b0 );
or ( \1394_b1 , \1344_b1 , w_4343 );
not ( w_4343 , w_4344 );
and ( \1394_b0 , \1344_b0 , w_4345 );
and ( w_4344 ,  , w_4345 );
buf ( w_4343 , \1393_b1 );
not ( w_4343 , w_4346 );
not (  , w_4347 );
and ( w_4346 , w_4347 , \1393_b0 );
or ( \1395_b1 , \1340_b1 , w_4349 );
not ( w_4349 , w_4350 );
and ( \1395_b0 , \1340_b0 , w_4351 );
and ( w_4350 ,  , w_4351 );
buf ( w_4349 , \1394_b1 );
not ( w_4349 , w_4352 );
not (  , w_4353 );
and ( w_4352 , w_4353 , \1394_b0 );
buf ( \1396_b1 , \a[4]_b1 );
not ( \1396_b1 , w_4354 );
not ( \1396_b0 , w_4355 );
and ( w_4354 , w_4355 , \a[4]_b0 );
or ( \1397_b1 , \1316_b1 , w_4357 );
not ( w_4357 , w_4358 );
and ( \1397_b0 , \1316_b0 , w_4359 );
and ( w_4358 ,  , w_4359 );
buf ( w_4357 , \1331_b1 );
not ( w_4357 , w_4360 );
not (  , w_4361 );
and ( w_4360 , w_4361 , \1331_b0 );
buf ( \1398_b1 , \1397_b1 );
not ( \1398_b1 , w_4362 );
not ( \1398_b0 , w_4363 );
and ( w_4362 , w_4363 , \1397_b0 );
or ( \1399_b1 , \1396_b1 , w_4364 );
or ( \1399_b0 , \1396_b0 , \1398_b0 );
not ( \1398_b0 , w_4365 );
and ( w_4365 , w_4364 , \1398_b1 );
or ( \1400_b1 , \b[4]_b1 , \c[4]_b1 );
not ( \c[4]_b1 , w_4366 );
and ( \1400_b0 , \b[4]_b0 , w_4367 );
and ( w_4366 , w_4367 , \c[4]_b0 );
or ( \1401_b1 , \1400_b1 , \1316_b1 );
not ( \1316_b1 , w_4368 );
and ( \1401_b0 , \1400_b0 , w_4369 );
and ( w_4368 , w_4369 , \1316_b0 );
or ( \1402_b1 , \a[4]_b1 , w_4370 );
or ( \1402_b0 , \a[4]_b0 , \b[4]_b0 );
not ( \b[4]_b0 , w_4371 );
and ( w_4371 , w_4370 , \b[4]_b1 );
buf ( \1403_b1 , \1402_b1 );
not ( \1403_b1 , w_4372 );
not ( \1403_b0 , w_4373 );
and ( w_4372 , w_4373 , \1402_b0 );
buf ( \1404_b1 , \671_b1 );
not ( \1404_b1 , w_4374 );
not ( \1404_b0 , w_4375 );
and ( w_4374 , w_4375 , \671_b0 );
or ( \1405_b1 , \1403_b1 , w_4376 );
or ( \1405_b0 , \1403_b0 , \1404_b0 );
not ( \1404_b0 , w_4377 );
and ( w_4377 , w_4376 , \1404_b1 );
or ( \1406_b1 , \c[4]_b1 , \d[4]_b1 );
xor ( \1406_b0 , \c[4]_b0 , w_4378 );
not ( w_4378 , w_4379 );
and ( w_4379 , \d[4]_b1 , \d[4]_b0 );
or ( \1407_b1 , \1383_b1 , w_4381 );
not ( w_4381 , w_4382 );
and ( \1407_b0 , \1383_b0 , w_4383 );
and ( w_4382 ,  , w_4383 );
buf ( w_4381 , \1406_b1 );
not ( w_4381 , w_4384 );
not (  , w_4385 );
and ( w_4384 , w_4385 , \1406_b0 );
or ( \1408_b1 , \875_b1 , w_4387 );
not ( w_4387 , w_4388 );
and ( \1408_b0 , \875_b0 , w_4389 );
and ( w_4388 ,  , w_4389 );
buf ( w_4387 , \878_b1 );
not ( w_4387 , w_4390 );
not (  , w_4391 );
and ( w_4390 , w_4391 , \878_b0 );
or ( \1409_b1 , \869_b1 , w_4392 );
xor ( \1409_b0 , \869_b0 , w_4394 );
not ( w_4394 , w_4395 );
and ( w_4395 , w_4392 , w_4393 );
buf ( w_4392 , \1408_b1 );
not ( w_4392 , w_4396 );
not ( w_4393 , w_4397 );
and ( w_4396 , w_4397 , \1408_b0 );
or ( \1410_b1 , \1409_b1 , w_4399 );
not ( w_4399 , w_4400 );
and ( \1410_b0 , \1409_b0 , w_4401 );
and ( w_4400 ,  , w_4401 );
buf ( w_4399 , \916_b1 );
not ( w_4399 , w_4402 );
not (  , w_4403 );
and ( w_4402 , w_4403 , \916_b0 );
or ( \1411_b1 , \1088_b1 , w_4405 );
not ( w_4405 , w_4406 );
and ( \1411_b0 , \1088_b0 , w_4407 );
and ( w_4406 ,  , w_4407 );
buf ( w_4405 , \1083_b1 );
not ( w_4405 , w_4408 );
not (  , w_4409 );
and ( w_4408 , w_4409 , \1083_b0 );
or ( \1412_b1 , \1411_b1 , w_4410 );
xor ( \1412_b0 , \1411_b0 , w_4412 );
not ( w_4412 , w_4413 );
and ( w_4413 , w_4410 , w_4411 );
buf ( w_4410 , \1077_b1 );
not ( w_4410 , w_4414 );
not ( w_4411 , w_4415 );
and ( w_4414 , w_4415 , \1077_b0 );
or ( \1413_b1 , \1168_b1 , \1412_b1 );
not ( \1412_b1 , w_4416 );
and ( \1413_b0 , \1168_b0 , w_4417 );
and ( w_4416 , w_4417 , \1412_b0 );
or ( \1414_b1 , \1198_b1 , w_4419 );
not ( w_4419 , w_4420 );
and ( \1414_b0 , \1198_b0 , w_4421 );
and ( w_4420 ,  , w_4421 );
buf ( w_4419 , \1190_b1 );
not ( w_4419 , w_4422 );
not (  , w_4423 );
and ( w_4422 , w_4423 , \1190_b0 );
buf ( \1415_b1 , \1414_b1 );
not ( \1415_b1 , w_4424 );
not ( \1415_b0 , w_4425 );
and ( w_4424 , w_4425 , \1414_b0 );
buf ( \1416_b1 , \1189_b1 );
not ( \1416_b1 , w_4426 );
not ( \1416_b0 , w_4427 );
and ( w_4426 , w_4427 , \1189_b0 );
buf ( \1417_b1 , \1416_b1 );
not ( \1417_b1 , w_4428 );
not ( \1417_b0 , w_4429 );
and ( w_4428 , w_4429 , \1416_b0 );
or ( \1418_b1 , \1415_b1 , w_4430 );
or ( \1418_b0 , \1415_b0 , \1417_b0 );
not ( \1417_b0 , w_4431 );
and ( w_4431 , w_4430 , \1417_b1 );
or ( \1419_b1 , \1416_b1 , w_4432 );
or ( \1419_b0 , \1416_b0 , \1414_b0 );
not ( \1414_b0 , w_4433 );
and ( w_4433 , w_4432 , \1414_b1 );
or ( \1420_b1 , \1418_b1 , w_4435 );
not ( w_4435 , w_4436 );
and ( \1420_b0 , \1418_b0 , w_4437 );
and ( w_4436 ,  , w_4437 );
buf ( w_4435 , \1419_b1 );
not ( w_4435 , w_4438 );
not (  , w_4439 );
and ( w_4438 , w_4439 , \1419_b0 );
buf ( \1421_b1 , \1420_b1 );
not ( \1421_b1 , w_4440 );
not ( \1421_b0 , w_4441 );
and ( w_4440 , w_4441 , \1420_b0 );
buf ( \1422_b1 , \1220_b1 );
not ( \1422_b1 , w_4442 );
not ( \1422_b0 , w_4443 );
and ( w_4442 , w_4443 , \1220_b0 );
or ( \1423_b1 , \1421_b1 , w_4444 );
or ( \1423_b0 , \1421_b0 , \1422_b0 );
not ( \1422_b0 , w_4445 );
and ( w_4445 , w_4444 , \1422_b1 );
or ( \1424_b1 , \1261_b1 , w_4447 );
not ( w_4447 , w_4448 );
and ( \1424_b0 , \1261_b0 , w_4449 );
and ( w_4448 ,  , w_4449 );
buf ( w_4447 , \1253_b1 );
not ( w_4447 , w_4450 );
not (  , w_4451 );
and ( w_4450 , w_4451 , \1253_b0 );
buf ( \1425_b1 , \1424_b1 );
not ( \1425_b1 , w_4452 );
not ( \1425_b0 , w_4453 );
and ( w_4452 , w_4453 , \1424_b0 );
buf ( \1426_b1 , \1252_b1 );
not ( \1426_b1 , w_4454 );
not ( \1426_b0 , w_4455 );
and ( w_4454 , w_4455 , \1252_b0 );
buf ( \1427_b1 , \1426_b1 );
not ( \1427_b1 , w_4456 );
not ( \1427_b0 , w_4457 );
and ( w_4456 , w_4457 , \1426_b0 );
or ( \1428_b1 , \1425_b1 , w_4458 );
or ( \1428_b0 , \1425_b0 , \1427_b0 );
not ( \1427_b0 , w_4459 );
and ( w_4459 , w_4458 , \1427_b1 );
or ( \1429_b1 , \1426_b1 , w_4460 );
or ( \1429_b0 , \1426_b0 , \1424_b0 );
not ( \1424_b0 , w_4461 );
and ( w_4461 , w_4460 , \1424_b1 );
or ( \1430_b1 , \1428_b1 , w_4463 );
not ( w_4463 , w_4464 );
and ( \1430_b0 , \1428_b0 , w_4465 );
and ( w_4464 ,  , w_4465 );
buf ( w_4463 , \1429_b1 );
not ( w_4463 , w_4466 );
not (  , w_4467 );
and ( w_4466 , w_4467 , \1429_b0 );
or ( \1431_b1 , \1232_b1 , \1430_b1 );
not ( \1430_b1 , w_4468 );
and ( \1431_b0 , \1232_b0 , w_4469 );
and ( w_4468 , w_4469 , \1430_b0 );
buf ( \1432_b1 , \d[4]_b1 );
not ( \1432_b1 , w_4470 );
not ( \1432_b0 , w_4471 );
and ( w_4470 , w_4471 , \d[4]_b0 );
buf ( \1433_b1 , \1280_b1 );
not ( \1433_b1 , w_4472 );
not ( \1433_b0 , w_4473 );
and ( w_4472 , w_4473 , \1280_b0 );
or ( \1434_b1 , \1432_b1 , w_4474 );
or ( \1434_b0 , \1432_b0 , \1433_b0 );
not ( \1433_b0 , w_4475 );
and ( w_4475 , w_4474 , \1433_b1 );
buf ( \1435_b1 , \1323_b1 );
not ( \1435_b1 , w_4476 );
not ( \1435_b0 , w_4477 );
and ( w_4476 , w_4477 , \1323_b0 );
or ( \1436_b1 , \1435_b1 , \c[4]_b1 );
not ( \c[4]_b1 , w_4478 );
and ( \1436_b0 , \1435_b0 , w_4479 );
and ( w_4478 , w_4479 , \c[4]_b0 );
or ( \1437_b1 , \1293_b1 , \b[4]_b1 );
not ( \b[4]_b1 , w_4480 );
and ( \1437_b0 , \1293_b0 , w_4481 );
and ( w_4480 , w_4481 , \b[4]_b0 );
or ( \1438_b1 , \1436_b1 , w_4483 );
not ( w_4483 , w_4484 );
and ( \1438_b0 , \1436_b0 , w_4485 );
and ( w_4484 ,  , w_4485 );
buf ( w_4483 , \1437_b1 );
not ( w_4483 , w_4486 );
not (  , w_4487 );
and ( w_4486 , w_4487 , \1437_b0 );
or ( \1439_b1 , \1434_b1 , w_4489 );
not ( w_4489 , w_4490 );
and ( \1439_b0 , \1434_b0 , w_4491 );
and ( w_4490 ,  , w_4491 );
buf ( w_4489 , \1438_b1 );
not ( w_4489 , w_4492 );
not (  , w_4493 );
and ( w_4492 , w_4493 , \1438_b0 );
or ( \1440_b1 , \1431_b1 , w_4495 );
not ( w_4495 , w_4496 );
and ( \1440_b0 , \1431_b0 , w_4497 );
and ( w_4496 ,  , w_4497 );
buf ( w_4495 , \1439_b1 );
not ( w_4495 , w_4498 );
not (  , w_4499 );
and ( w_4498 , w_4499 , \1439_b0 );
or ( \1441_b1 , \1423_b1 , w_4501 );
not ( w_4501 , w_4502 );
and ( \1441_b0 , \1423_b0 , w_4503 );
and ( w_4502 ,  , w_4503 );
buf ( w_4501 , \1440_b1 );
not ( w_4501 , w_4504 );
not (  , w_4505 );
and ( w_4504 , w_4505 , \1440_b0 );
or ( \1442_b1 , \1413_b1 , w_4507 );
not ( w_4507 , w_4508 );
and ( \1442_b0 , \1413_b0 , w_4509 );
and ( w_4508 ,  , w_4509 );
buf ( w_4507 , \1441_b1 );
not ( w_4507 , w_4510 );
not (  , w_4511 );
and ( w_4510 , w_4511 , \1441_b0 );
or ( \1444_b1 , \1405_b1 , w_4513 );
not ( w_4513 , w_4514 );
and ( \1444_b0 , \1405_b0 , w_4515 );
and ( w_4514 ,  , w_4515 );
buf ( w_4513 , \1443_b1 );
not ( w_4513 , w_4516 );
not (  , w_4517 );
and ( w_4516 , w_4517 , \1443_b0 );
or ( \1445_b1 , \1401_b1 , w_4519 );
not ( w_4519 , w_4520 );
and ( \1445_b0 , \1401_b0 , w_4521 );
and ( w_4520 ,  , w_4521 );
buf ( w_4519 , \1444_b1 );
not ( w_4519 , w_4522 );
not (  , w_4523 );
and ( w_4522 , w_4523 , \1444_b0 );
or ( \1446_b1 , \1399_b1 , w_4525 );
not ( w_4525 , w_4526 );
and ( \1446_b0 , \1399_b0 , w_4527 );
and ( w_4526 ,  , w_4527 );
buf ( w_4525 , \1445_b1 );
not ( w_4525 , w_4528 );
not (  , w_4529 );
and ( w_4528 , w_4529 , \1445_b0 );
buf ( \1447_b1 , \d[4]_b1 );
not ( \1447_b1 , w_4530 );
not ( \1447_b0 , w_4531 );
and ( w_4530 , w_4531 , \d[4]_b0 );
buf ( \1448_b1 , \644_b1 );
not ( \1448_b1 , w_4532 );
not ( \1448_b0 , w_4533 );
and ( w_4532 , w_4533 , \644_b0 );
or ( \1449_b1 , \1447_b1 , w_4534 );
or ( \1449_b0 , \1447_b0 , \1448_b0 );
not ( \1448_b0 , w_4535 );
and ( w_4535 , w_4534 , \1448_b1 );
buf ( \1450_b1 , \1341_b1 );
not ( \1450_b1 , w_4536 );
not ( \1450_b0 , w_4537 );
and ( w_4536 , w_4537 , \1341_b0 );
or ( \1451_b1 , \1450_b1 , w_4539 );
not ( w_4539 , w_4540 );
and ( \1451_b0 , \1450_b0 , w_4541 );
and ( w_4540 ,  , w_4541 );
buf ( w_4539 , \a[4]_b1 );
not ( w_4539 , w_4542 );
not (  , w_4543 );
and ( w_4542 , w_4543 , \a[4]_b0 );
or ( \1452_b1 , \1449_b1 , w_4545 );
not ( w_4545 , w_4546 );
and ( \1452_b0 , \1449_b0 , w_4547 );
and ( w_4546 ,  , w_4547 );
buf ( w_4545 , \1451_b1 );
not ( w_4545 , w_4548 );
not (  , w_4549 );
and ( w_4548 , w_4549 , \1451_b0 );
or ( \1453_b1 , \1446_b1 , w_4551 );
not ( w_4551 , w_4552 );
and ( \1453_b0 , \1446_b0 , w_4553 );
and ( w_4552 ,  , w_4553 );
buf ( w_4551 , \1452_b1 );
not ( w_4551 , w_4554 );
not (  , w_4555 );
and ( w_4554 , w_4555 , \1452_b0 );
buf ( \1454_b1 , \1453_b1 );
not ( \1454_b1 , w_4556 );
not ( \1454_b0 , w_4557 );
and ( w_4556 , w_4557 , \1453_b0 );
or ( \1455_b1 , \a[3]_b1 , w_4558 );
or ( \1455_b0 , \a[3]_b0 , \d[3]_b0 );
not ( \d[3]_b0 , w_4559 );
and ( w_4559 , w_4558 , \d[3]_b1 );
buf ( \1456_b1 , \1455_b1 );
not ( \1456_b1 , w_4560 );
not ( \1456_b0 , w_4561 );
and ( w_4560 , w_4561 , \1455_b0 );
buf ( \1457_b1 , \1341_b1 );
not ( \1457_b1 , w_4562 );
not ( \1457_b0 , w_4563 );
and ( w_4562 , w_4563 , \1341_b0 );
buf ( \1458_b1 , \1457_b1 );
not ( \1458_b1 , w_4564 );
not ( \1458_b0 , w_4565 );
and ( w_4564 , w_4565 , \1457_b0 );
or ( \1459_b1 , \1456_b1 , w_4566 );
or ( \1459_b0 , \1456_b0 , \1458_b0 );
not ( \1458_b0 , w_4567 );
and ( w_4567 , w_4566 , \1458_b1 );
or ( \1460_b1 , \b[3]_b1 , \c[3]_b1 );
not ( \c[3]_b1 , w_4568 );
and ( \1460_b0 , \b[3]_b0 , w_4569 );
and ( w_4568 , w_4569 , \c[3]_b0 );
or ( \1461_b1 , \1316_b1 , \1460_b1 );
not ( \1460_b1 , w_4570 );
and ( \1461_b0 , \1316_b0 , w_4571 );
and ( w_4570 , w_4571 , \1460_b0 );
buf ( \1462_b1 , \a[3]_b1 );
not ( \1462_b1 , w_4572 );
not ( \1462_b0 , w_4573 );
and ( w_4572 , w_4573 , \a[3]_b0 );
buf ( \1463_b1 , \b[3]_b1 );
not ( \1463_b1 , w_4574 );
not ( \1463_b0 , w_4575 );
and ( w_4574 , w_4575 , \b[3]_b0 );
or ( \1464_b1 , \1462_b1 , w_4577 );
not ( w_4577 , w_4578 );
and ( \1464_b0 , \1462_b0 , w_4579 );
and ( w_4578 ,  , w_4579 );
buf ( w_4577 , \1463_b1 );
not ( w_4577 , w_4580 );
not (  , w_4581 );
and ( w_4580 , w_4581 , \1463_b0 );
buf ( \1465_b1 , \1464_b1 );
not ( \1465_b1 , w_4582 );
not ( \1465_b0 , w_4583 );
and ( w_4582 , w_4583 , \1464_b0 );
buf ( \1466_b1 , \1350_b1 );
not ( \1466_b1 , w_4584 );
not ( \1466_b0 , w_4585 );
and ( w_4584 , w_4585 , \1350_b0 );
buf ( \1467_b1 , \1466_b1 );
not ( \1467_b1 , w_4586 );
not ( \1467_b0 , w_4587 );
and ( w_4586 , w_4587 , \1466_b0 );
or ( \1468_b1 , \1465_b1 , w_4588 );
or ( \1468_b0 , \1465_b0 , \1467_b0 );
not ( \1467_b0 , w_4589 );
and ( w_4589 , w_4588 , \1467_b1 );
buf ( \1469_b1 , \917_b1 );
not ( \1469_b1 , w_4590 );
not ( \1469_b0 , w_4591 );
and ( w_4590 , w_4591 , \917_b0 );
or ( \1470_b1 , \868_b1 , w_4593 );
not ( w_4593 , w_4594 );
and ( \1470_b0 , \868_b0 , w_4595 );
and ( w_4594 ,  , w_4595 );
buf ( w_4593 , \842_b1 );
not ( w_4593 , w_4596 );
not (  , w_4597 );
and ( w_4596 , w_4597 , \842_b0 );
or ( \1471_b1 , \864_b1 , \1470_b1 );
xor ( \1471_b0 , \864_b0 , w_4598 );
not ( w_4598 , w_4599 );
and ( w_4599 , \1470_b1 , \1470_b0 );
buf ( \1472_b1 , \1471_b1 );
not ( \1472_b1 , w_4600 );
not ( \1472_b0 , w_4601 );
and ( w_4600 , w_4601 , \1471_b0 );
or ( \1473_b1 , \1469_b1 , \1472_b1 );
not ( \1472_b1 , w_4602 );
and ( \1473_b0 , \1469_b0 , w_4603 );
and ( w_4602 , w_4603 , \1472_b0 );
or ( \1474_b1 , \c[3]_b1 , \d[3]_b1 );
xor ( \1474_b0 , \c[3]_b0 , w_4604 );
not ( w_4604 , w_4605 );
and ( w_4605 , \d[3]_b1 , \d[3]_b0 );
buf ( \1475_b1 , \1474_b1 );
not ( \1475_b1 , w_4606 );
not ( \1475_b0 , w_4607 );
and ( w_4606 , w_4607 , \1474_b0 );
buf ( \1476_b1 , \1320_b1 );
not ( \1476_b1 , w_4608 );
not ( \1476_b0 , w_4609 );
and ( w_4608 , w_4609 , \1320_b0 );
or ( \1477_b1 , \1475_b1 , w_4610 );
or ( \1477_b0 , \1475_b0 , \1476_b0 );
not ( \1476_b0 , w_4611 );
and ( w_4611 , w_4610 , \1476_b1 );
buf ( \1478_b1 , \1167_b1 );
not ( \1478_b1 , w_4612 );
not ( \1478_b0 , w_4613 );
and ( w_4612 , w_4613 , \1167_b0 );
or ( \1479_b1 , \1071_b1 , w_4615 );
not ( w_4615 , w_4616 );
and ( \1479_b0 , \1071_b0 , w_4617 );
and ( w_4616 ,  , w_4617 );
buf ( w_4615 , \1076_b1 );
not ( w_4615 , w_4618 );
not (  , w_4619 );
and ( w_4618 , w_4619 , \1076_b0 );
or ( \1480_b1 , \1479_b1 , w_4620 );
xor ( \1480_b0 , \1479_b0 , w_4622 );
not ( w_4622 , w_4623 );
and ( w_4623 , w_4620 , w_4621 );
buf ( w_4620 , \1050_b1 );
not ( w_4620 , w_4624 );
not ( w_4621 , w_4625 );
and ( w_4624 , w_4625 , \1050_b0 );
or ( \1481_b1 , \1478_b1 , \1480_b1 );
not ( \1480_b1 , w_4626 );
and ( \1481_b0 , \1478_b0 , w_4627 );
and ( w_4626 , w_4627 , \1480_b0 );
buf ( \1482_b1 , \1171_b1 );
not ( \1482_b1 , w_4628 );
not ( \1482_b0 , w_4629 );
and ( w_4628 , w_4629 , \1171_b0 );
or ( \1483_b1 , \1482_b1 , w_4631 );
not ( w_4631 , w_4632 );
and ( \1483_b0 , \1482_b0 , w_4633 );
and ( w_4632 ,  , w_4633 );
buf ( w_4631 , \1184_b1 );
not ( w_4631 , w_4634 );
not (  , w_4635 );
and ( w_4634 , w_4635 , \1184_b0 );
buf ( \1484_b1 , \1483_b1 );
not ( \1484_b1 , w_4636 );
not ( \1484_b0 , w_4637 );
and ( w_4636 , w_4637 , \1483_b0 );
or ( \1485_b1 , \1174_b1 , w_4639 );
not ( w_4639 , w_4640 );
and ( \1485_b0 , \1174_b0 , w_4641 );
and ( w_4640 ,  , w_4641 );
buf ( w_4639 , \1180_b1 );
not ( w_4639 , w_4642 );
not (  , w_4643 );
and ( w_4642 , w_4643 , \1180_b0 );
buf ( \1486_b1 , \1170_b1 );
not ( \1486_b1 , w_4644 );
not ( \1486_b0 , w_4645 );
and ( w_4644 , w_4645 , \1170_b0 );
or ( \1488_b1 , \1487_b1 , w_4647 );
not ( w_4647 , w_4648 );
and ( \1488_b0 , \1487_b0 , w_4649 );
and ( w_4648 ,  , w_4649 );
buf ( w_4647 , \1186_b1 );
not ( w_4647 , w_4650 );
not (  , w_4651 );
and ( w_4650 , w_4651 , \1186_b0 );
buf ( \1489_b1 , \1488_b1 );
not ( \1489_b1 , w_4652 );
not ( \1489_b0 , w_4653 );
and ( w_4652 , w_4653 , \1488_b0 );
or ( \1490_b1 , \1484_b1 , w_4654 );
or ( \1490_b0 , \1484_b0 , \1489_b0 );
not ( \1489_b0 , w_4655 );
and ( w_4655 , w_4654 , \1489_b1 );
or ( \1491_b1 , \1488_b1 , w_4656 );
or ( \1491_b0 , \1488_b0 , \1483_b0 );
not ( \1483_b0 , w_4657 );
and ( w_4657 , w_4656 , \1483_b1 );
or ( \1492_b1 , \1490_b1 , w_4659 );
not ( w_4659 , w_4660 );
and ( \1492_b0 , \1490_b0 , w_4661 );
and ( w_4660 ,  , w_4661 );
buf ( w_4659 , \1491_b1 );
not ( w_4659 , w_4662 );
not (  , w_4663 );
and ( w_4662 , w_4663 , \1491_b0 );
buf ( \1493_b1 , \1492_b1 );
not ( \1493_b1 , w_4664 );
not ( \1493_b0 , w_4665 );
and ( w_4664 , w_4665 , \1492_b0 );
buf ( \1494_b1 , \1220_b1 );
not ( \1494_b1 , w_4666 );
not ( \1494_b0 , w_4667 );
and ( w_4666 , w_4667 , \1220_b0 );
or ( \1495_b1 , \1493_b1 , w_4668 );
or ( \1495_b0 , \1493_b0 , \1494_b0 );
not ( \1494_b0 , w_4669 );
and ( w_4669 , w_4668 , \1494_b1 );
buf ( \1496_b1 , \1234_b1 );
not ( \1496_b1 , w_4670 );
not ( \1496_b0 , w_4671 );
and ( w_4670 , w_4671 , \1234_b0 );
or ( \1497_b1 , \1496_b1 , w_4673 );
not ( w_4673 , w_4674 );
and ( \1497_b0 , \1496_b0 , w_4675 );
and ( w_4674 ,  , w_4675 );
buf ( w_4673 , \1247_b1 );
not ( w_4673 , w_4676 );
not (  , w_4677 );
and ( w_4676 , w_4677 , \1247_b0 );
buf ( \1498_b1 , \1497_b1 );
not ( \1498_b1 , w_4678 );
not ( \1498_b0 , w_4679 );
and ( w_4678 , w_4679 , \1497_b0 );
or ( \1499_b1 , \1237_b1 , w_4681 );
not ( w_4681 , w_4682 );
and ( \1499_b0 , \1237_b0 , w_4683 );
and ( w_4682 ,  , w_4683 );
buf ( w_4681 , \1243_b1 );
not ( w_4681 , w_4684 );
not (  , w_4685 );
and ( w_4684 , w_4685 , \1243_b0 );
buf ( \1500_b1 , \1233_b1 );
not ( \1500_b1 , w_4686 );
not ( \1500_b0 , w_4687 );
and ( w_4686 , w_4687 , \1233_b0 );
or ( \1502_b1 , \1501_b1 , w_4689 );
not ( w_4689 , w_4690 );
and ( \1502_b0 , \1501_b0 , w_4691 );
and ( w_4690 ,  , w_4691 );
buf ( w_4689 , \1249_b1 );
not ( w_4689 , w_4692 );
not (  , w_4693 );
and ( w_4692 , w_4693 , \1249_b0 );
buf ( \1503_b1 , \1502_b1 );
not ( \1503_b1 , w_4694 );
not ( \1503_b0 , w_4695 );
and ( w_4694 , w_4695 , \1502_b0 );
or ( \1504_b1 , \1498_b1 , w_4696 );
or ( \1504_b0 , \1498_b0 , \1503_b0 );
not ( \1503_b0 , w_4697 );
and ( w_4697 , w_4696 , \1503_b1 );
or ( \1505_b1 , \1502_b1 , w_4698 );
or ( \1505_b0 , \1502_b0 , \1497_b0 );
not ( \1497_b0 , w_4699 );
and ( w_4699 , w_4698 , \1497_b1 );
or ( \1506_b1 , \1504_b1 , w_4701 );
not ( w_4701 , w_4702 );
and ( \1506_b0 , \1504_b0 , w_4703 );
and ( w_4702 ,  , w_4703 );
buf ( w_4701 , \1505_b1 );
not ( w_4701 , w_4704 );
not (  , w_4705 );
and ( w_4704 , w_4705 , \1505_b0 );
or ( \1507_b1 , \1232_b1 , \1506_b1 );
not ( \1506_b1 , w_4706 );
and ( \1507_b0 , \1232_b0 , w_4707 );
and ( w_4706 , w_4707 , \1506_b0 );
buf ( \1508_b1 , \d[3]_b1 );
not ( \1508_b1 , w_4708 );
not ( \1508_b0 , w_4709 );
and ( w_4708 , w_4709 , \d[3]_b0 );
buf ( \1509_b1 , \1280_b1 );
not ( \1509_b1 , w_4710 );
not ( \1509_b0 , w_4711 );
and ( w_4710 , w_4711 , \1280_b0 );
or ( \1510_b1 , \1508_b1 , w_4712 );
or ( \1510_b0 , \1508_b0 , \1509_b0 );
not ( \1509_b0 , w_4713 );
and ( w_4713 , w_4712 , \1509_b1 );
buf ( \1511_b1 , \1324_b1 );
not ( \1511_b1 , w_4714 );
not ( \1511_b0 , w_4715 );
and ( w_4714 , w_4715 , \1324_b0 );
buf ( \1512_b1 , \1463_b1 );
not ( \1512_b1 , w_4716 );
not ( \1512_b0 , w_4717 );
and ( w_4716 , w_4717 , \1463_b0 );
or ( \1513_b1 , \1511_b1 , \1512_b1 );
not ( \1512_b1 , w_4718 );
and ( \1513_b0 , \1511_b0 , w_4719 );
and ( w_4718 , w_4719 , \1512_b0 );
buf ( \1514_b1 , \1323_b1 );
not ( \1514_b1 , w_4720 );
not ( \1514_b0 , w_4721 );
and ( w_4720 , w_4721 , \1323_b0 );
or ( \1515_b1 , \1514_b1 , \c[3]_b1 );
not ( \c[3]_b1 , w_4722 );
and ( \1515_b0 , \1514_b0 , w_4723 );
and ( w_4722 , w_4723 , \c[3]_b0 );
or ( \1516_b1 , \1513_b1 , w_4725 );
not ( w_4725 , w_4726 );
and ( \1516_b0 , \1513_b0 , w_4727 );
and ( w_4726 ,  , w_4727 );
buf ( w_4725 , \1515_b1 );
not ( w_4725 , w_4728 );
not (  , w_4729 );
and ( w_4728 , w_4729 , \1515_b0 );
or ( \1517_b1 , \1510_b1 , w_4731 );
not ( w_4731 , w_4732 );
and ( \1517_b0 , \1510_b0 , w_4733 );
and ( w_4732 ,  , w_4733 );
buf ( w_4731 , \1516_b1 );
not ( w_4731 , w_4734 );
not (  , w_4735 );
and ( w_4734 , w_4735 , \1516_b0 );
or ( \1518_b1 , \1507_b1 , w_4737 );
not ( w_4737 , w_4738 );
and ( \1518_b0 , \1507_b0 , w_4739 );
and ( w_4738 ,  , w_4739 );
buf ( w_4737 , \1517_b1 );
not ( w_4737 , w_4740 );
not (  , w_4741 );
and ( w_4740 , w_4741 , \1517_b0 );
or ( \1519_b1 , \1495_b1 , w_4743 );
not ( w_4743 , w_4744 );
and ( \1519_b0 , \1495_b0 , w_4745 );
and ( w_4744 ,  , w_4745 );
buf ( w_4743 , \1518_b1 );
not ( w_4743 , w_4746 );
not (  , w_4747 );
and ( w_4746 , w_4747 , \1518_b0 );
or ( \1520_b1 , \1481_b1 , w_4749 );
not ( w_4749 , w_4750 );
and ( \1520_b0 , \1481_b0 , w_4751 );
and ( w_4750 ,  , w_4751 );
buf ( w_4749 , \1519_b1 );
not ( w_4749 , w_4752 );
not (  , w_4753 );
and ( w_4752 , w_4753 , \1519_b0 );
or ( \1521_b1 , \1477_b1 , w_4755 );
not ( w_4755 , w_4756 );
and ( \1521_b0 , \1477_b0 , w_4757 );
and ( w_4756 ,  , w_4757 );
buf ( w_4755 , \1520_b1 );
not ( w_4755 , w_4758 );
not (  , w_4759 );
and ( w_4758 , w_4759 , \1520_b0 );
or ( \1522_b1 , \1473_b1 , w_4761 );
not ( w_4761 , w_4762 );
and ( \1522_b0 , \1473_b0 , w_4763 );
and ( w_4762 ,  , w_4763 );
buf ( w_4761 , \1521_b1 );
not ( w_4761 , w_4764 );
not (  , w_4765 );
and ( w_4764 , w_4765 , \1521_b0 );
or ( \1523_b1 , \1468_b1 , w_4767 );
not ( w_4767 , w_4768 );
and ( \1523_b0 , \1468_b0 , w_4769 );
and ( w_4768 ,  , w_4769 );
buf ( w_4767 , \1522_b1 );
not ( w_4767 , w_4770 );
not (  , w_4771 );
and ( w_4770 , w_4771 , \1522_b0 );
or ( \1524_b1 , \1461_b1 , w_4773 );
not ( w_4773 , w_4774 );
and ( \1524_b0 , \1461_b0 , w_4775 );
and ( w_4774 ,  , w_4775 );
buf ( w_4773 , \1523_b1 );
not ( w_4773 , w_4776 );
not (  , w_4777 );
and ( w_4776 , w_4777 , \1523_b0 );
or ( \1525_b1 , \1459_b1 , w_4779 );
not ( w_4779 , w_4780 );
and ( \1525_b0 , \1459_b0 , w_4781 );
and ( w_4780 ,  , w_4781 );
buf ( w_4779 , \1524_b1 );
not ( w_4779 , w_4782 );
not (  , w_4783 );
and ( w_4782 , w_4783 , \1524_b0 );
or ( \1526_b1 , \1338_b1 , \a[3]_b1 );
not ( \a[3]_b1 , w_4784 );
and ( \1526_b0 , \1338_b0 , w_4785 );
and ( w_4784 , w_4785 , \a[3]_b0 );
or ( \1527_b1 , \1525_b1 , w_4787 );
not ( w_4787 , w_4788 );
and ( \1527_b0 , \1525_b0 , w_4789 );
and ( w_4788 ,  , w_4789 );
buf ( w_4787 , \1526_b1 );
not ( w_4787 , w_4790 );
not (  , w_4791 );
and ( w_4790 , w_4791 , \1526_b0 );
buf ( \1528_b1 , \1527_b1 );
not ( \1528_b1 , w_4792 );
not ( \1528_b0 , w_4793 );
and ( w_4792 , w_4793 , \1527_b0 );
buf ( \1529_b1 , \1478_b1 );
buf ( \1529_b0 , \1478_b0 );
buf ( \1530_b1 , \1529_b1 );
not ( \1530_b1 , w_4794 );
not ( \1530_b0 , w_4795 );
and ( w_4794 , w_4795 , \1529_b0 );
or ( \1531_b1 , \a[9]_b1 , \d[7]_b1 );
xor ( \1531_b0 , \a[9]_b0 , w_4796 );
not ( w_4796 , w_4797 );
and ( w_4797 , \d[7]_b1 , \d[7]_b0 );
buf ( \1532_b1 , \1531_b1 );
not ( \1532_b1 , w_4798 );
not ( \1532_b0 , w_4799 );
and ( w_4798 , w_4799 , \1531_b0 );
buf ( \1533_b1 , \958_b1 );
not ( \1533_b1 , w_4800 );
not ( \1533_b0 , w_4801 );
and ( w_4800 , w_4801 , \958_b0 );
or ( \1534_b1 , \1532_b1 , w_4802 );
or ( \1534_b0 , \1532_b0 , \1533_b0 );
not ( \1533_b0 , w_4803 );
and ( w_4803 , w_4802 , \1533_b1 );
or ( \1535_b1 , \a[8]_b1 , \d[7]_b1 );
xor ( \1535_b0 , \a[8]_b0 , w_4804 );
not ( w_4804 , w_4805 );
and ( w_4805 , \d[7]_b1 , \d[7]_b0 );
or ( \1536_b1 , \1128_b1 , w_4807 );
not ( w_4807 , w_4808 );
and ( \1536_b0 , \1128_b0 , w_4809 );
and ( w_4808 ,  , w_4809 );
buf ( w_4807 , \1535_b1 );
not ( w_4807 , w_4810 );
not (  , w_4811 );
and ( w_4810 , w_4811 , \1535_b0 );
or ( \1537_b1 , \1534_b1 , w_4813 );
not ( w_4813 , w_4814 );
and ( \1537_b0 , \1534_b0 , w_4815 );
and ( w_4814 ,  , w_4815 );
buf ( w_4813 , \1536_b1 );
not ( w_4813 , w_4816 );
not (  , w_4817 );
and ( w_4816 , w_4817 , \1536_b0 );
or ( \1538_b1 , \a[6]_b1 , \d[9]_b1 );
xor ( \1538_b0 , \a[6]_b0 , w_4818 );
not ( w_4818 , w_4819 );
and ( w_4819 , \d[9]_b1 , \d[9]_b0 );
buf ( \1539_b1 , \1538_b1 );
not ( \1539_b1 , w_4820 );
not ( \1539_b0 , w_4821 );
and ( w_4820 , w_4821 , \1538_b0 );
or ( \1540_b1 , \d[9]_b1 , w_4822 );
xor ( \1540_b0 , \d[9]_b0 , w_4824 );
not ( w_4824 , w_4825 );
and ( w_4825 , w_4822 , w_4823 );
buf ( w_4822 , \d[8]_b1 );
not ( w_4822 , w_4826 );
not ( w_4823 , w_4827 );
and ( w_4826 , w_4827 , \d[8]_b0 );
or ( \1541_b1 , \d[8]_b1 , \d[7]_b1 );
xor ( \1541_b0 , \d[8]_b0 , w_4828 );
not ( w_4828 , w_4829 );
and ( w_4829 , \d[7]_b1 , \d[7]_b0 );
or ( \1542_b1 , \1540_b1 , w_4831 );
not ( w_4831 , w_4832 );
and ( \1542_b0 , \1540_b0 , w_4833 );
and ( w_4832 ,  , w_4833 );
buf ( w_4831 , \1541_b1 );
not ( w_4831 , w_4834 );
not (  , w_4835 );
and ( w_4834 , w_4835 , \1541_b0 );
buf ( \1543_b1 , \1542_b1 );
not ( \1543_b1 , w_4836 );
not ( \1543_b0 , w_4837 );
and ( w_4836 , w_4837 , \1542_b0 );
or ( \1544_b1 , \1539_b1 , w_4838 );
or ( \1544_b0 , \1539_b0 , \1543_b0 );
not ( \1543_b0 , w_4839 );
and ( w_4839 , w_4838 , \1543_b1 );
buf ( \1545_b1 , \1541_b1 );
buf ( \1545_b0 , \1541_b0 );
or ( \1546_b1 , \a[7]_b1 , \d[9]_b1 );
xor ( \1546_b0 , \a[7]_b0 , w_4840 );
not ( w_4840 , w_4841 );
and ( w_4841 , \d[9]_b1 , \d[9]_b0 );
or ( \1547_b1 , \1545_b1 , w_4843 );
not ( w_4843 , w_4844 );
and ( \1547_b0 , \1545_b0 , w_4845 );
and ( w_4844 ,  , w_4845 );
buf ( w_4843 , \1546_b1 );
not ( w_4843 , w_4846 );
not (  , w_4847 );
and ( w_4846 , w_4847 , \1546_b0 );
or ( \1548_b1 , \1544_b1 , w_4849 );
not ( w_4849 , w_4850 );
and ( \1548_b0 , \1544_b0 , w_4851 );
and ( w_4850 ,  , w_4851 );
buf ( w_4849 , \1547_b1 );
not ( w_4849 , w_4852 );
not (  , w_4853 );
and ( w_4852 , w_4853 , \1547_b0 );
or ( \1549_b1 , \1537_b1 , \1548_b1 );
xor ( \1549_b0 , \1537_b0 , w_4854 );
not ( w_4854 , w_4855 );
and ( w_4855 , \1548_b1 , \1548_b0 );
or ( \1550_b1 , \a[2]_b1 , \d[13]_b1 );
xor ( \1550_b0 , \a[2]_b0 , w_4856 );
not ( w_4856 , w_4857 );
and ( w_4857 , \d[13]_b1 , \d[13]_b0 );
buf ( \1551_b1 , \1550_b1 );
not ( \1551_b1 , w_4858 );
not ( \1551_b0 , w_4859 );
and ( w_4858 , w_4859 , \1550_b0 );
or ( \1552_b1 , \d[12]_b1 , \d[11]_b1 );
xor ( \1552_b0 , \d[12]_b0 , w_4860 );
not ( w_4860 , w_4861 );
and ( w_4861 , \d[11]_b1 , \d[11]_b0 );
or ( \1553_b1 , \d[13]_b1 , w_4862 );
xor ( \1553_b0 , \d[13]_b0 , w_4864 );
not ( w_4864 , w_4865 );
and ( w_4865 , w_4862 , w_4863 );
buf ( w_4862 , \d[12]_b1 );
not ( w_4862 , w_4866 );
not ( w_4863 , w_4867 );
and ( w_4866 , w_4867 , \d[12]_b0 );
or ( \1554_b1 , \1552_b1 , w_4869 );
not ( w_4869 , w_4870 );
and ( \1554_b0 , \1552_b0 , w_4871 );
and ( w_4870 ,  , w_4871 );
buf ( w_4869 , \1553_b1 );
not ( w_4869 , w_4872 );
not (  , w_4873 );
and ( w_4872 , w_4873 , \1553_b0 );
buf ( \1555_b1 , \1554_b1 );
not ( \1555_b1 , w_4874 );
not ( \1555_b0 , w_4875 );
and ( w_4874 , w_4875 , \1554_b0 );
or ( \1556_b1 , \1551_b1 , w_4876 );
or ( \1556_b0 , \1551_b0 , \1555_b0 );
not ( \1555_b0 , w_4877 );
and ( w_4877 , w_4876 , \1555_b1 );
or ( \1557_b1 , \a[3]_b1 , \d[13]_b1 );
xor ( \1557_b0 , \a[3]_b0 , w_4878 );
not ( w_4878 , w_4879 );
and ( w_4879 , \d[13]_b1 , \d[13]_b0 );
or ( \1558_b1 , \1552_b1 , w_4881 );
not ( w_4881 , w_4882 );
and ( \1558_b0 , \1552_b0 , w_4883 );
and ( w_4882 ,  , w_4883 );
buf ( w_4881 , \1557_b1 );
not ( w_4881 , w_4884 );
not (  , w_4885 );
and ( w_4884 , w_4885 , \1557_b0 );
or ( \1559_b1 , \1556_b1 , w_4887 );
not ( w_4887 , w_4888 );
and ( \1559_b0 , \1556_b0 , w_4889 );
and ( w_4888 ,  , w_4889 );
buf ( w_4887 , \1558_b1 );
not ( w_4887 , w_4890 );
not (  , w_4891 );
and ( w_4890 , w_4891 , \1558_b0 );
or ( \1560_b1 , \d[15]_b1 , \d[14]_b1 );
xor ( \1560_b0 , \d[15]_b0 , w_4892 );
not ( w_4892 , w_4893 );
and ( w_4893 , \d[14]_b1 , \d[14]_b0 );
or ( \1561_b1 , \a[0]_b1 , \d[15]_b1 );
xor ( \1561_b0 , \a[0]_b0 , w_4894 );
not ( w_4894 , w_4895 );
and ( w_4895 , \d[15]_b1 , \d[15]_b0 );
or ( \1562_b1 , \1560_b1 , w_4897 );
not ( w_4897 , w_4898 );
and ( \1562_b0 , \1560_b0 , w_4899 );
and ( w_4898 ,  , w_4899 );
buf ( w_4897 , \1561_b1 );
not ( w_4897 , w_4900 );
not (  , w_4901 );
and ( w_4900 , w_4901 , \1561_b0 );
or ( \1563_b1 , \d[14]_b1 , \d[13]_b1 );
xor ( \1563_b0 , \d[14]_b0 , w_4902 );
not ( w_4902 , w_4903 );
and ( w_4903 , \d[13]_b1 , \d[13]_b0 );
or ( \1564_b1 , \1562_b1 , w_4904 );
or ( \1564_b0 , \1562_b0 , \1563_b0 );
not ( \1563_b0 , w_4905 );
and ( w_4905 , w_4904 , \1563_b1 );
or ( \1565_b1 , \a[1]_b1 , \d[15]_b1 );
xor ( \1565_b0 , \a[1]_b0 , w_4906 );
not ( w_4906 , w_4907 );
and ( w_4907 , \d[15]_b1 , \d[15]_b0 );
or ( \1566_b1 , \1563_b1 , w_4909 );
not ( w_4909 , w_4910 );
and ( \1566_b0 , \1563_b0 , w_4911 );
and ( w_4910 ,  , w_4911 );
buf ( w_4909 , \1565_b1 );
not ( w_4909 , w_4912 );
not (  , w_4913 );
and ( w_4912 , w_4913 , \1565_b0 );
or ( \1567_b1 , \1564_b1 , w_4915 );
not ( w_4915 , w_4916 );
and ( \1567_b0 , \1564_b0 , w_4917 );
and ( w_4916 ,  , w_4917 );
buf ( w_4915 , \1566_b1 );
not ( w_4915 , w_4918 );
not (  , w_4919 );
and ( w_4918 , w_4919 , \1566_b0 );
or ( \1568_b1 , \1559_b1 , \1567_b1 );
xor ( \1568_b0 , \1559_b0 , w_4920 );
not ( w_4920 , w_4921 );
and ( w_4921 , \1567_b1 , \1567_b0 );
or ( \1569_b1 , \1549_b1 , \1568_b1 );
xor ( \1569_b0 , \1549_b0 , w_4922 );
not ( w_4922 , w_4923 );
and ( w_4923 , \1568_b1 , \1568_b0 );
buf ( \1570_b1 , \1569_b1 );
not ( \1570_b1 , w_4924 );
not ( \1570_b0 , w_4925 );
and ( w_4924 , w_4925 , \1569_b0 );
or ( \1571_b1 , \1563_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_4926 );
and ( \1571_b0 , \1563_b0 , w_4927 );
and ( w_4926 , w_4927 , \a[0]_b0 );
or ( \1572_b1 , \a[13]_b1 , \d[1]_b1 );
xor ( \1572_b0 , \a[13]_b0 , w_4928 );
not ( w_4928 , w_4929 );
and ( w_4929 , \d[1]_b1 , \d[1]_b0 );
buf ( \1573_b1 , \1572_b1 );
not ( \1573_b1 , w_4930 );
not ( \1573_b0 , w_4931 );
and ( w_4930 , w_4931 , \1572_b0 );
buf ( \1574_b1 , \932_b1 );
not ( \1574_b1 , w_4932 );
not ( \1574_b0 , w_4933 );
and ( w_4932 , w_4933 , \932_b0 );
or ( \1575_b1 , \1573_b1 , w_4934 );
or ( \1575_b0 , \1573_b0 , \1574_b0 );
not ( \1574_b0 , w_4935 );
and ( w_4935 , w_4934 , \1574_b1 );
or ( \1576_b1 , \a[14]_b1 , \d[1]_b1 );
xor ( \1576_b0 , \a[14]_b0 , w_4936 );
not ( w_4936 , w_4937 );
and ( w_4937 , \d[1]_b1 , \d[1]_b0 );
or ( \1577_b1 , \1576_b1 , w_4939 );
not ( w_4939 , w_4940 );
and ( \1577_b0 , \1576_b0 , w_4941 );
and ( w_4940 ,  , w_4941 );
buf ( w_4939 , \d[0]_b1 );
not ( w_4939 , w_4942 );
not (  , w_4943 );
and ( w_4942 , w_4943 , \d[0]_b0 );
or ( \1578_b1 , \1575_b1 , w_4945 );
not ( w_4945 , w_4946 );
and ( \1578_b0 , \1575_b0 , w_4947 );
and ( w_4946 ,  , w_4947 );
buf ( w_4945 , \1577_b1 );
not ( w_4945 , w_4948 );
not (  , w_4949 );
and ( w_4948 , w_4949 , \1577_b0 );
or ( \1579_b1 , \1571_b1 , \1578_b1 );
xor ( \1579_b0 , \1571_b0 , w_4950 );
not ( w_4950 , w_4951 );
and ( w_4951 , \1578_b1 , \1578_b0 );
or ( \1580_b1 , \a[11]_b1 , \d[3]_b1 );
xor ( \1580_b0 , \a[11]_b0 , w_4952 );
not ( w_4952 , w_4953 );
and ( w_4953 , \d[3]_b1 , \d[3]_b0 );
buf ( \1581_b1 , \1580_b1 );
not ( \1581_b1 , w_4954 );
not ( \1581_b0 , w_4955 );
and ( w_4954 , w_4955 , \1580_b0 );
buf ( \1582_b1 , \973_b1 );
not ( \1582_b1 , w_4956 );
not ( \1582_b0 , w_4957 );
and ( w_4956 , w_4957 , \973_b0 );
or ( \1583_b1 , \1581_b1 , w_4958 );
or ( \1583_b0 , \1581_b0 , \1582_b0 );
not ( \1582_b0 , w_4959 );
and ( w_4959 , w_4958 , \1582_b1 );
or ( \1584_b1 , \a[12]_b1 , \d[3]_b1 );
xor ( \1584_b0 , \a[12]_b0 , w_4960 );
not ( w_4960 , w_4961 );
and ( w_4961 , \d[3]_b1 , \d[3]_b0 );
or ( \1585_b1 , \976_b1 , w_4963 );
not ( w_4963 , w_4964 );
and ( \1585_b0 , \976_b0 , w_4965 );
and ( w_4964 ,  , w_4965 );
buf ( w_4963 , \1584_b1 );
not ( w_4963 , w_4966 );
not (  , w_4967 );
and ( w_4966 , w_4967 , \1584_b0 );
or ( \1586_b1 , \1583_b1 , w_4969 );
not ( w_4969 , w_4970 );
and ( \1586_b0 , \1583_b0 , w_4971 );
and ( w_4970 ,  , w_4971 );
buf ( w_4969 , \1585_b1 );
not ( w_4969 , w_4972 );
not (  , w_4973 );
and ( w_4972 , w_4973 , \1585_b0 );
or ( \1587_b1 , \1579_b1 , \1586_b1 );
not ( \1586_b1 , w_4974 );
and ( \1587_b0 , \1579_b0 , w_4975 );
and ( w_4974 , w_4975 , \1586_b0 );
or ( \1588_b1 , \1571_b1 , \1578_b1 );
not ( \1578_b1 , w_4976 );
and ( \1588_b0 , \1571_b0 , w_4977 );
and ( w_4976 , w_4977 , \1578_b0 );
or ( \1589_b1 , \1587_b1 , w_4978 );
or ( \1589_b0 , \1587_b0 , \1588_b0 );
not ( \1588_b0 , w_4979 );
and ( w_4979 , w_4978 , \1588_b1 );
buf ( \1590_b1 , \1589_b1 );
not ( \1590_b1 , w_4980 );
not ( \1590_b0 , w_4981 );
and ( w_4980 , w_4981 , \1589_b0 );
buf ( \1591_b1 , \1584_b1 );
not ( \1591_b1 , w_4982 );
not ( \1591_b0 , w_4983 );
and ( w_4982 , w_4983 , \1584_b0 );
buf ( \1592_b1 , \973_b1 );
not ( \1592_b1 , w_4984 );
not ( \1592_b0 , w_4985 );
and ( w_4984 , w_4985 , \973_b0 );
or ( \1593_b1 , \1591_b1 , w_4986 );
or ( \1593_b0 , \1591_b0 , \1592_b0 );
not ( \1592_b0 , w_4987 );
and ( w_4987 , w_4986 , \1592_b1 );
buf ( \1594_b1 , \d[3]_b1 );
not ( \1594_b1 , w_4988 );
not ( \1594_b0 , w_4989 );
and ( w_4988 , w_4989 , \d[3]_b0 );
or ( \1595_b1 , \1594_b1 , w_4991 );
not ( w_4991 , w_4992 );
and ( \1595_b0 , \1594_b0 , w_4993 );
and ( w_4992 ,  , w_4993 );
buf ( w_4991 , \a[13]_b1 );
not ( w_4991 , w_4994 );
not (  , w_4995 );
and ( w_4994 , w_4995 , \a[13]_b0 );
buf ( \1596_b1 , \1595_b1 );
not ( \1596_b1 , w_4996 );
not ( \1596_b0 , w_4997 );
and ( w_4996 , w_4997 , \1595_b0 );
buf ( \1597_b1 , \a[13]_b1 );
not ( \1597_b1 , w_4998 );
not ( \1597_b0 , w_4999 );
and ( w_4998 , w_4999 , \a[13]_b0 );
or ( \1598_b1 , \1597_b1 , w_5001 );
not ( w_5001 , w_5002 );
and ( \1598_b0 , \1597_b0 , w_5003 );
and ( w_5002 ,  , w_5003 );
buf ( w_5001 , \d[3]_b1 );
not ( w_5001 , w_5004 );
not (  , w_5005 );
and ( w_5004 , w_5005 , \d[3]_b0 );
buf ( \1599_b1 , \1598_b1 );
not ( \1599_b1 , w_5006 );
not ( \1599_b0 , w_5007 );
and ( w_5006 , w_5007 , \1598_b0 );
or ( \1600_b1 , \1596_b1 , w_5008 );
or ( \1600_b0 , \1596_b0 , \1599_b0 );
not ( \1599_b0 , w_5009 );
and ( w_5009 , w_5008 , \1599_b1 );
or ( \1601_b1 , \1600_b1 , w_5011 );
not ( w_5011 , w_5012 );
and ( \1601_b0 , \1600_b0 , w_5013 );
and ( w_5012 ,  , w_5013 );
buf ( w_5011 , \976_b1 );
not ( w_5011 , w_5014 );
not (  , w_5015 );
and ( w_5014 , w_5015 , \976_b0 );
or ( \1602_b1 , \1593_b1 , w_5017 );
not ( w_5017 , w_5018 );
and ( \1602_b0 , \1593_b0 , w_5019 );
and ( w_5018 ,  , w_5019 );
buf ( w_5017 , \1601_b1 );
not ( w_5017 , w_5020 );
not (  , w_5021 );
and ( w_5020 , w_5021 , \1601_b0 );
or ( \1603_b1 , \a[10]_b1 , \d[5]_b1 );
xor ( \1603_b0 , \a[10]_b0 , w_5022 );
not ( w_5022 , w_5023 );
and ( w_5023 , \d[5]_b1 , \d[5]_b0 );
buf ( \1604_b1 , \1603_b1 );
not ( \1604_b1 , w_5024 );
not ( \1604_b0 , w_5025 );
and ( w_5024 , w_5025 , \1603_b0 );
buf ( \1605_b1 , \1135_b1 );
not ( \1605_b1 , w_5026 );
not ( \1605_b0 , w_5027 );
and ( w_5026 , w_5027 , \1135_b0 );
or ( \1606_b1 , \1604_b1 , w_5028 );
or ( \1606_b0 , \1604_b0 , \1605_b0 );
not ( \1605_b0 , w_5029 );
and ( w_5029 , w_5028 , \1605_b1 );
buf ( \1607_b1 , \d[5]_b1 );
not ( \1607_b1 , w_5030 );
not ( \1607_b0 , w_5031 );
and ( w_5030 , w_5031 , \d[5]_b0 );
or ( \1608_b1 , \1607_b1 , w_5033 );
not ( w_5033 , w_5034 );
and ( \1608_b0 , \1607_b0 , w_5035 );
and ( w_5034 ,  , w_5035 );
buf ( w_5033 , \a[11]_b1 );
not ( w_5033 , w_5036 );
not (  , w_5037 );
and ( w_5036 , w_5037 , \a[11]_b0 );
buf ( \1609_b1 , \1608_b1 );
not ( \1609_b1 , w_5038 );
not ( \1609_b0 , w_5039 );
and ( w_5038 , w_5039 , \1608_b0 );
buf ( \1610_b1 , \a[11]_b1 );
not ( \1610_b1 , w_5040 );
not ( \1610_b0 , w_5041 );
and ( w_5040 , w_5041 , \a[11]_b0 );
or ( \1611_b1 , \1610_b1 , w_5043 );
not ( w_5043 , w_5044 );
and ( \1611_b0 , \1610_b0 , w_5045 );
and ( w_5044 ,  , w_5045 );
buf ( w_5043 , \d[5]_b1 );
not ( w_5043 , w_5046 );
not (  , w_5047 );
and ( w_5046 , w_5047 , \d[5]_b0 );
buf ( \1612_b1 , \1611_b1 );
not ( \1612_b1 , w_5048 );
not ( \1612_b0 , w_5049 );
and ( w_5048 , w_5049 , \1611_b0 );
or ( \1613_b1 , \1609_b1 , w_5050 );
or ( \1613_b0 , \1609_b0 , \1612_b0 );
not ( \1612_b0 , w_5051 );
and ( w_5051 , w_5050 , \1612_b1 );
or ( \1614_b1 , \1613_b1 , w_5053 );
not ( w_5053 , w_5054 );
and ( \1614_b0 , \1613_b0 , w_5055 );
and ( w_5054 ,  , w_5055 );
buf ( w_5053 , \951_b1 );
not ( w_5053 , w_5056 );
not (  , w_5057 );
and ( w_5056 , w_5057 , \951_b0 );
or ( \1615_b1 , \1606_b1 , w_5059 );
not ( w_5059 , w_5060 );
and ( \1615_b0 , \1606_b0 , w_5061 );
and ( w_5060 ,  , w_5061 );
buf ( w_5059 , \1614_b1 );
not ( w_5059 , w_5062 );
not (  , w_5063 );
and ( w_5062 , w_5063 , \1614_b0 );
buf ( \1616_b1 , \1615_b1 );
not ( \1616_b1 , w_5064 );
not ( \1616_b0 , w_5065 );
and ( w_5064 , w_5065 , \1615_b0 );
or ( \1617_b1 , \1602_b1 , \1616_b1 );
xor ( \1617_b0 , \1602_b0 , w_5066 );
not ( w_5066 , w_5067 );
and ( w_5067 , \1616_b1 , \1616_b0 );
buf ( \1618_b1 , \1617_b1 );
not ( \1618_b1 , w_5068 );
not ( \1618_b0 , w_5069 );
and ( w_5068 , w_5069 , \1617_b0 );
or ( \1619_b1 , \1590_b1 , \1618_b1 );
not ( \1618_b1 , w_5070 );
and ( \1619_b0 , \1590_b0 , w_5071 );
and ( w_5070 , w_5071 , \1618_b0 );
or ( \1620_b1 , \1589_b1 , \1617_b1 );
not ( \1617_b1 , w_5072 );
and ( \1620_b0 , \1589_b0 , w_5073 );
and ( w_5072 , w_5073 , \1617_b0 );
or ( \1621_b1 , \1619_b1 , w_5075 );
not ( w_5075 , w_5076 );
and ( \1621_b0 , \1619_b0 , w_5077 );
and ( w_5076 ,  , w_5077 );
buf ( w_5075 , \1620_b1 );
not ( w_5075 , w_5078 );
not (  , w_5079 );
and ( w_5078 , w_5079 , \1620_b0 );
buf ( \1622_b1 , \1621_b1 );
not ( \1622_b1 , w_5080 );
not ( \1622_b0 , w_5081 );
and ( w_5080 , w_5081 , \1621_b0 );
or ( \1623_b1 , \1570_b1 , w_5082 );
or ( \1623_b0 , \1570_b0 , \1622_b0 );
not ( \1622_b0 , w_5083 );
and ( w_5083 , w_5082 , \1622_b1 );
or ( \1624_b1 , \1569_b1 , w_5084 );
or ( \1624_b0 , \1569_b0 , \1621_b0 );
not ( \1621_b0 , w_5085 );
and ( w_5085 , w_5084 , \1621_b1 );
or ( \1625_b1 , \1623_b1 , w_5087 );
not ( w_5087 , w_5088 );
and ( \1625_b0 , \1623_b0 , w_5089 );
and ( w_5088 ,  , w_5089 );
buf ( w_5087 , \1624_b1 );
not ( w_5087 , w_5090 );
not (  , w_5091 );
and ( w_5090 , w_5091 , \1624_b0 );
buf ( \1626_b1 , \1625_b1 );
not ( \1626_b1 , w_5092 );
not ( \1626_b0 , w_5093 );
and ( w_5092 , w_5093 , \1625_b0 );
or ( \1627_b1 , \a[1]_b1 , \d[13]_b1 );
xor ( \1627_b0 , \a[1]_b0 , w_5094 );
not ( w_5094 , w_5095 );
and ( w_5095 , \d[13]_b1 , \d[13]_b0 );
buf ( \1628_b1 , \1627_b1 );
not ( \1628_b1 , w_5096 );
not ( \1628_b0 , w_5097 );
and ( w_5096 , w_5097 , \1627_b0 );
buf ( \1629_b1 , \1554_b1 );
not ( \1629_b1 , w_5098 );
not ( \1629_b0 , w_5099 );
and ( w_5098 , w_5099 , \1554_b0 );
or ( \1630_b1 , \1628_b1 , w_5100 );
or ( \1630_b0 , \1628_b0 , \1629_b0 );
not ( \1629_b0 , w_5101 );
and ( w_5101 , w_5100 , \1629_b1 );
or ( \1631_b1 , \1552_b1 , w_5103 );
not ( w_5103 , w_5104 );
and ( \1631_b0 , \1552_b0 , w_5105 );
and ( w_5104 ,  , w_5105 );
buf ( w_5103 , \1550_b1 );
not ( w_5103 , w_5106 );
not (  , w_5107 );
and ( w_5106 , w_5107 , \1550_b0 );
or ( \1632_b1 , \1630_b1 , w_5109 );
not ( w_5109 , w_5110 );
and ( \1632_b0 , \1630_b0 , w_5111 );
and ( w_5110 ,  , w_5111 );
buf ( w_5109 , \1631_b1 );
not ( w_5109 , w_5112 );
not (  , w_5113 );
and ( w_5112 , w_5113 , \1631_b0 );
or ( \1633_b1 , \a[3]_b1 , \d[11]_b1 );
xor ( \1633_b0 , \a[3]_b0 , w_5114 );
not ( w_5114 , w_5115 );
and ( w_5115 , \d[11]_b1 , \d[11]_b0 );
buf ( \1634_b1 , \1633_b1 );
not ( \1634_b1 , w_5116 );
not ( \1634_b0 , w_5117 );
and ( w_5116 , w_5117 , \1633_b0 );
or ( \1635_b1 , \d[10]_b1 , \d[9]_b1 );
xor ( \1635_b0 , \d[10]_b0 , w_5118 );
not ( w_5118 , w_5119 );
and ( w_5119 , \d[9]_b1 , \d[9]_b0 );
buf ( \1636_b1 , \d[10]_b1 );
not ( \1636_b1 , w_5120 );
not ( \1636_b0 , w_5121 );
and ( w_5120 , w_5121 , \d[10]_b0 );
or ( \1637_b1 , \d[11]_b1 , \1636_b1 );
xor ( \1637_b0 , \d[11]_b0 , w_5122 );
not ( w_5122 , w_5123 );
and ( w_5123 , \1636_b1 , \1636_b0 );
or ( \1638_b1 , \1635_b1 , w_5125 );
not ( w_5125 , w_5126 );
and ( \1638_b0 , \1635_b0 , w_5127 );
and ( w_5126 ,  , w_5127 );
buf ( w_5125 , \1637_b1 );
not ( w_5125 , w_5128 );
not (  , w_5129 );
and ( w_5128 , w_5129 , \1637_b0 );
buf ( \1639_b1 , \1638_b1 );
not ( \1639_b1 , w_5130 );
not ( \1639_b0 , w_5131 );
and ( w_5130 , w_5131 , \1638_b0 );
or ( \1640_b1 , \1634_b1 , w_5132 );
or ( \1640_b0 , \1634_b0 , \1639_b0 );
not ( \1639_b0 , w_5133 );
and ( w_5133 , w_5132 , \1639_b1 );
or ( \1641_b1 , \d[10]_b1 , \d[9]_b1 );
xor ( \1641_b0 , \d[10]_b0 , w_5134 );
not ( w_5134 , w_5135 );
and ( w_5135 , \d[9]_b1 , \d[9]_b0 );
or ( \1642_b1 , \a[4]_b1 , \d[11]_b1 );
xor ( \1642_b0 , \a[4]_b0 , w_5136 );
not ( w_5136 , w_5137 );
and ( w_5137 , \d[11]_b1 , \d[11]_b0 );
or ( \1643_b1 , \1641_b1 , w_5139 );
not ( w_5139 , w_5140 );
and ( \1643_b0 , \1641_b0 , w_5141 );
and ( w_5140 ,  , w_5141 );
buf ( w_5139 , \1642_b1 );
not ( w_5139 , w_5142 );
not (  , w_5143 );
and ( w_5142 , w_5143 , \1642_b0 );
or ( \1644_b1 , \1640_b1 , w_5145 );
not ( w_5145 , w_5146 );
and ( \1644_b0 , \1640_b0 , w_5147 );
and ( w_5146 ,  , w_5147 );
buf ( w_5145 , \1643_b1 );
not ( w_5145 , w_5148 );
not (  , w_5149 );
and ( w_5148 , w_5149 , \1643_b0 );
or ( \1645_b1 , \1632_b1 , \1644_b1 );
xor ( \1645_b0 , \1632_b0 , w_5150 );
not ( w_5150 , w_5151 );
and ( w_5151 , \1644_b1 , \1644_b0 );
or ( \1646_b1 , \a[0]_b1 , w_5152 );
or ( \1646_b0 , \a[0]_b0 , \d[12]_b0 );
not ( \d[12]_b0 , w_5153 );
and ( w_5153 , w_5152 , \d[12]_b1 );
or ( \1647_b1 , \1646_b1 , w_5155 );
not ( w_5155 , w_5156 );
and ( \1647_b0 , \1646_b0 , w_5157 );
and ( w_5156 ,  , w_5157 );
buf ( w_5155 , \d[11]_b1 );
not ( w_5155 , w_5158 );
not (  , w_5159 );
and ( w_5158 , w_5159 , \d[11]_b0 );
or ( \1648_b1 , \a[0]_b1 , w_5161 );
not ( w_5161 , w_5162 );
and ( \1648_b0 , \a[0]_b0 , w_5163 );
and ( w_5162 ,  , w_5163 );
buf ( w_5161 , \d[12]_b1 );
not ( w_5161 , w_5164 );
not (  , w_5165 );
and ( w_5164 , w_5165 , \d[12]_b0 );
or ( \1650_b1 , \a[12]_b1 , \d[1]_b1 );
xor ( \1650_b0 , \a[12]_b0 , w_5166 );
not ( w_5166 , w_5167 );
and ( w_5167 , \d[1]_b1 , \d[1]_b0 );
buf ( \1651_b1 , \1650_b1 );
not ( \1651_b1 , w_5168 );
not ( \1651_b0 , w_5169 );
and ( w_5168 , w_5169 , \1650_b0 );
buf ( \1652_b1 , \932_b1 );
not ( \1652_b1 , w_5170 );
not ( \1652_b0 , w_5171 );
and ( w_5170 , w_5171 , \932_b0 );
or ( \1653_b1 , \1651_b1 , w_5172 );
or ( \1653_b0 , \1651_b0 , \1652_b0 );
not ( \1652_b0 , w_5173 );
and ( w_5173 , w_5172 , \1652_b1 );
or ( \1654_b1 , \1572_b1 , w_5175 );
not ( w_5175 , w_5176 );
and ( \1654_b0 , \1572_b0 , w_5177 );
and ( w_5176 ,  , w_5177 );
buf ( w_5175 , \d[0]_b1 );
not ( w_5175 , w_5178 );
not (  , w_5179 );
and ( w_5178 , w_5179 , \d[0]_b0 );
or ( \1655_b1 , \1653_b1 , w_5181 );
not ( w_5181 , w_5182 );
and ( \1655_b0 , \1653_b0 , w_5183 );
and ( w_5182 ,  , w_5183 );
buf ( w_5181 , \1654_b1 );
not ( w_5181 , w_5184 );
not (  , w_5185 );
and ( w_5184 , w_5185 , \1654_b0 );
or ( \1656_b1 , \1649_b1 , \1655_b1 );
not ( \1655_b1 , w_5186 );
and ( \1656_b0 , \1649_b0 , w_5187 );
and ( w_5186 , w_5187 , \1655_b0 );
or ( \1657_b1 , \1645_b1 , \1656_b1 );
not ( \1656_b1 , w_5188 );
and ( \1657_b0 , \1645_b0 , w_5189 );
and ( w_5188 , w_5189 , \1656_b0 );
or ( \1658_b1 , \1632_b1 , \1644_b1 );
not ( \1644_b1 , w_5190 );
and ( \1658_b0 , \1632_b0 , w_5191 );
and ( w_5190 , w_5191 , \1644_b0 );
or ( \1659_b1 , \1657_b1 , w_5192 );
or ( \1659_b0 , \1657_b0 , \1658_b0 );
not ( \1658_b0 , w_5193 );
and ( w_5193 , w_5192 , \1658_b1 );
buf ( \1660_b1 , \1576_b1 );
not ( \1660_b1 , w_5194 );
not ( \1660_b0 , w_5195 );
and ( w_5194 , w_5195 , \1576_b0 );
buf ( \1661_b1 , \932_b1 );
not ( \1661_b1 , w_5196 );
not ( \1661_b0 , w_5197 );
and ( w_5196 , w_5197 , \932_b0 );
or ( \1662_b1 , \1660_b1 , w_5198 );
or ( \1662_b0 , \1660_b0 , \1661_b0 );
not ( \1661_b0 , w_5199 );
and ( w_5199 , w_5198 , \1661_b1 );
or ( \1663_b1 , \a[15]_b1 , \d[1]_b1 );
xor ( \1663_b0 , \a[15]_b0 , w_5200 );
not ( w_5200 , w_5201 );
and ( w_5201 , \d[1]_b1 , \d[1]_b0 );
or ( \1664_b1 , \1663_b1 , w_5203 );
not ( w_5203 , w_5204 );
and ( \1664_b0 , \1663_b0 , w_5205 );
and ( w_5204 ,  , w_5205 );
buf ( w_5203 , \d[0]_b1 );
not ( w_5203 , w_5206 );
not (  , w_5207 );
and ( w_5206 , w_5207 , \d[0]_b0 );
or ( \1665_b1 , \1662_b1 , w_5209 );
not ( w_5209 , w_5210 );
and ( \1665_b0 , \1662_b0 , w_5211 );
and ( w_5210 ,  , w_5211 );
buf ( w_5209 , \1664_b1 );
not ( w_5209 , w_5212 );
not (  , w_5213 );
and ( w_5212 , w_5213 , \1664_b0 );
or ( \1666_b1 , \a[0]_b1 , w_5214 );
or ( \1666_b0 , \a[0]_b0 , \d[14]_b0 );
not ( \d[14]_b0 , w_5215 );
and ( w_5215 , w_5214 , \d[14]_b1 );
or ( \1667_b1 , \1666_b1 , w_5217 );
not ( w_5217 , w_5218 );
and ( \1667_b0 , \1666_b0 , w_5219 );
and ( w_5218 ,  , w_5219 );
buf ( w_5217 , \d[13]_b1 );
not ( w_5217 , w_5220 );
not (  , w_5221 );
and ( w_5220 , w_5221 , \d[13]_b0 );
or ( \1668_b1 , \a[0]_b1 , w_5223 );
not ( w_5223 , w_5224 );
and ( \1668_b0 , \a[0]_b0 , w_5225 );
and ( w_5224 ,  , w_5225 );
buf ( w_5223 , \d[14]_b1 );
not ( w_5223 , w_5226 );
not (  , w_5227 );
and ( w_5226 , w_5227 , \d[14]_b0 );
or ( \1670_b1 , \1665_b1 , \1669_b1 );
xor ( \1670_b0 , \1665_b0 , w_5228 );
not ( w_5228 , w_5229 );
and ( w_5229 , \1669_b1 , \1669_b0 );
buf ( \1671_b1 , \1642_b1 );
not ( \1671_b1 , w_5230 );
not ( \1671_b0 , w_5231 );
and ( w_5230 , w_5231 , \1642_b0 );
buf ( \1672_b1 , \1638_b1 );
not ( \1672_b1 , w_5232 );
not ( \1672_b0 , w_5233 );
and ( w_5232 , w_5233 , \1638_b0 );
or ( \1673_b1 , \1671_b1 , w_5234 );
or ( \1673_b0 , \1671_b0 , \1672_b0 );
not ( \1672_b0 , w_5235 );
and ( w_5235 , w_5234 , \1672_b1 );
or ( \1674_b1 , \a[5]_b1 , \d[11]_b1 );
xor ( \1674_b0 , \a[5]_b0 , w_5236 );
not ( w_5236 , w_5237 );
and ( w_5237 , \d[11]_b1 , \d[11]_b0 );
or ( \1675_b1 , \1641_b1 , w_5239 );
not ( w_5239 , w_5240 );
and ( \1675_b0 , \1641_b0 , w_5241 );
and ( w_5240 ,  , w_5241 );
buf ( w_5239 , \1674_b1 );
not ( w_5239 , w_5242 );
not (  , w_5243 );
and ( w_5242 , w_5243 , \1674_b0 );
or ( \1676_b1 , \1673_b1 , w_5245 );
not ( w_5245 , w_5246 );
and ( \1676_b0 , \1673_b0 , w_5247 );
and ( w_5246 ,  , w_5247 );
buf ( w_5245 , \1675_b1 );
not ( w_5245 , w_5248 );
not (  , w_5249 );
and ( w_5248 , w_5249 , \1675_b0 );
or ( \1677_b1 , \1670_b1 , w_5250 );
xor ( \1677_b0 , \1670_b0 , w_5252 );
not ( w_5252 , w_5253 );
and ( w_5253 , w_5250 , w_5251 );
buf ( w_5250 , \1676_b1 );
not ( w_5250 , w_5254 );
not ( w_5251 , w_5255 );
and ( w_5254 , w_5255 , \1676_b0 );
or ( \1678_b1 , \1659_b1 , \1677_b1 );
xor ( \1678_b0 , \1659_b0 , w_5256 );
not ( w_5256 , w_5257 );
and ( w_5257 , \1677_b1 , \1677_b0 );
or ( \1679_b1 , \a[7]_b1 , \d[7]_b1 );
xor ( \1679_b0 , \a[7]_b0 , w_5258 );
not ( w_5258 , w_5259 );
and ( w_5259 , \d[7]_b1 , \d[7]_b0 );
buf ( \1680_b1 , \1679_b1 );
not ( \1680_b1 , w_5260 );
not ( \1680_b0 , w_5261 );
and ( w_5260 , w_5261 , \1679_b0 );
buf ( \1681_b1 , \1127_b1 );
not ( \1681_b1 , w_5262 );
not ( \1681_b0 , w_5263 );
and ( w_5262 , w_5263 , \1127_b0 );
or ( \1682_b1 , \1680_b1 , w_5264 );
or ( \1682_b0 , \1680_b0 , \1681_b0 );
not ( \1681_b0 , w_5265 );
and ( w_5265 , w_5264 , \1681_b1 );
or ( \1683_b1 , \958_b1 , w_5267 );
not ( w_5267 , w_5268 );
and ( \1683_b0 , \958_b0 , w_5269 );
and ( w_5268 ,  , w_5269 );
buf ( w_5267 , \1535_b1 );
not ( w_5267 , w_5270 );
not (  , w_5271 );
and ( w_5270 , w_5271 , \1535_b0 );
or ( \1684_b1 , \1682_b1 , w_5273 );
not ( w_5273 , w_5274 );
and ( \1684_b0 , \1682_b0 , w_5275 );
and ( w_5274 ,  , w_5275 );
buf ( w_5273 , \1683_b1 );
not ( w_5273 , w_5276 );
not (  , w_5277 );
and ( w_5276 , w_5277 , \1683_b0 );
or ( \1685_b1 , \a[5]_b1 , \d[9]_b1 );
xor ( \1685_b0 , \a[5]_b0 , w_5278 );
not ( w_5278 , w_5279 );
and ( w_5279 , \d[9]_b1 , \d[9]_b0 );
buf ( \1686_b1 , \1685_b1 );
not ( \1686_b1 , w_5280 );
not ( \1686_b0 , w_5281 );
and ( w_5280 , w_5281 , \1685_b0 );
buf ( \1687_b1 , \1542_b1 );
not ( \1687_b1 , w_5282 );
not ( \1687_b0 , w_5283 );
and ( w_5282 , w_5283 , \1542_b0 );
or ( \1688_b1 , \1686_b1 , w_5284 );
or ( \1688_b0 , \1686_b0 , \1687_b0 );
not ( \1687_b0 , w_5285 );
and ( w_5285 , w_5284 , \1687_b1 );
or ( \1689_b1 , \1545_b1 , w_5287 );
not ( w_5287 , w_5288 );
and ( \1689_b0 , \1545_b0 , w_5289 );
and ( w_5288 ,  , w_5289 );
buf ( w_5287 , \1538_b1 );
not ( w_5287 , w_5290 );
not (  , w_5291 );
and ( w_5290 , w_5291 , \1538_b0 );
or ( \1690_b1 , \1688_b1 , w_5293 );
not ( w_5293 , w_5294 );
and ( \1690_b0 , \1688_b0 , w_5295 );
and ( w_5294 ,  , w_5295 );
buf ( w_5293 , \1689_b1 );
not ( w_5293 , w_5296 );
not (  , w_5297 );
and ( w_5296 , w_5297 , \1689_b0 );
or ( \1691_b1 , \1684_b1 , \1690_b1 );
xor ( \1691_b0 , \1684_b0 , w_5298 );
not ( w_5298 , w_5299 );
and ( w_5299 , \1690_b1 , \1690_b0 );
or ( \1692_b1 , \a[9]_b1 , \d[5]_b1 );
xor ( \1692_b0 , \a[9]_b0 , w_5300 );
not ( w_5300 , w_5301 );
and ( w_5301 , \d[5]_b1 , \d[5]_b0 );
buf ( \1693_b1 , \1692_b1 );
not ( \1693_b1 , w_5302 );
not ( \1693_b0 , w_5303 );
and ( w_5302 , w_5303 , \1692_b0 );
buf ( \1694_b1 , \1135_b1 );
not ( \1694_b1 , w_5304 );
not ( \1694_b0 , w_5305 );
and ( w_5304 , w_5305 , \1135_b0 );
or ( \1695_b1 , \1693_b1 , w_5306 );
or ( \1695_b0 , \1693_b0 , \1694_b0 );
not ( \1694_b0 , w_5307 );
and ( w_5307 , w_5306 , \1694_b1 );
or ( \1696_b1 , \951_b1 , w_5309 );
not ( w_5309 , w_5310 );
and ( \1696_b0 , \951_b0 , w_5311 );
and ( w_5310 ,  , w_5311 );
buf ( w_5309 , \1603_b1 );
not ( w_5309 , w_5312 );
not (  , w_5313 );
and ( w_5312 , w_5313 , \1603_b0 );
or ( \1697_b1 , \1695_b1 , w_5315 );
not ( w_5315 , w_5316 );
and ( \1697_b0 , \1695_b0 , w_5317 );
and ( w_5316 ,  , w_5317 );
buf ( w_5315 , \1696_b1 );
not ( w_5315 , w_5318 );
not (  , w_5319 );
and ( w_5318 , w_5319 , \1696_b0 );
or ( \1698_b1 , \1691_b1 , \1697_b1 );
not ( \1697_b1 , w_5320 );
and ( \1698_b0 , \1691_b0 , w_5321 );
and ( w_5320 , w_5321 , \1697_b0 );
or ( \1699_b1 , \1684_b1 , \1690_b1 );
not ( \1690_b1 , w_5322 );
and ( \1699_b0 , \1684_b0 , w_5323 );
and ( w_5322 , w_5323 , \1690_b0 );
or ( \1700_b1 , \1698_b1 , w_5324 );
or ( \1700_b0 , \1698_b0 , \1699_b0 );
not ( \1699_b0 , w_5325 );
and ( w_5325 , w_5324 , \1699_b1 );
buf ( \1701_b1 , \1700_b1 );
not ( \1701_b1 , w_5326 );
not ( \1701_b0 , w_5327 );
and ( w_5326 , w_5327 , \1700_b0 );
or ( \1702_b1 , \1678_b1 , \1701_b1 );
not ( \1701_b1 , w_5328 );
and ( \1702_b0 , \1678_b0 , w_5329 );
and ( w_5328 , w_5329 , \1701_b0 );
buf ( \1703_b1 , \1678_b1 );
not ( \1703_b1 , w_5330 );
not ( \1703_b0 , w_5331 );
and ( w_5330 , w_5331 , \1678_b0 );
or ( \1704_b1 , \1703_b1 , \1700_b1 );
not ( \1700_b1 , w_5332 );
and ( \1704_b0 , \1703_b0 , w_5333 );
and ( w_5332 , w_5333 , \1700_b0 );
or ( \1705_b1 , \1702_b1 , w_5335 );
not ( w_5335 , w_5336 );
and ( \1705_b0 , \1702_b0 , w_5337 );
and ( w_5336 ,  , w_5337 );
buf ( w_5335 , \1704_b1 );
not ( w_5335 , w_5338 );
not (  , w_5339 );
and ( w_5338 , w_5339 , \1704_b0 );
buf ( \1706_b1 , \1705_b1 );
not ( \1706_b1 , w_5340 );
not ( \1706_b0 , w_5341 );
and ( w_5340 , w_5341 , \1705_b0 );
or ( \1707_b1 , \1626_b1 , w_5342 );
or ( \1707_b0 , \1626_b0 , \1706_b0 );
not ( \1706_b0 , w_5343 );
and ( w_5343 , w_5342 , \1706_b1 );
or ( \1708_b1 , \1705_b1 , w_5344 );
or ( \1708_b0 , \1705_b0 , \1625_b0 );
not ( \1625_b0 , w_5345 );
and ( w_5345 , w_5344 , \1625_b1 );
or ( \1709_b1 , \1707_b1 , w_5347 );
not ( w_5347 , w_5348 );
and ( \1709_b0 , \1707_b0 , w_5349 );
and ( w_5348 ,  , w_5349 );
buf ( w_5347 , \1708_b1 );
not ( w_5347 , w_5350 );
not (  , w_5351 );
and ( w_5350 , w_5351 , \1708_b0 );
or ( \1710_b1 , \1571_b1 , \1578_b1 );
xor ( \1710_b0 , \1571_b0 , w_5352 );
not ( w_5352 , w_5353 );
and ( w_5353 , \1578_b1 , \1578_b0 );
or ( \1711_b1 , \1710_b1 , \1586_b1 );
xor ( \1711_b0 , \1710_b0 , w_5354 );
not ( w_5354 , w_5355 );
and ( w_5355 , \1586_b1 , \1586_b0 );
or ( \1712_b1 , \a[0]_b1 , \d[13]_b1 );
xor ( \1712_b0 , \a[0]_b0 , w_5356 );
not ( w_5356 , w_5357 );
and ( w_5357 , \d[13]_b1 , \d[13]_b0 );
buf ( \1713_b1 , \1712_b1 );
not ( \1713_b1 , w_5358 );
not ( \1713_b0 , w_5359 );
and ( w_5358 , w_5359 , \1712_b0 );
or ( \1714_b1 , \1552_b1 , w_5361 );
not ( w_5361 , w_5362 );
and ( \1714_b0 , \1552_b0 , w_5363 );
and ( w_5362 ,  , w_5363 );
buf ( w_5361 , \1553_b1 );
not ( w_5361 , w_5364 );
not (  , w_5365 );
and ( w_5364 , w_5365 , \1553_b0 );
buf ( \1715_b1 , \1714_b1 );
not ( \1715_b1 , w_5366 );
not ( \1715_b0 , w_5367 );
and ( w_5366 , w_5367 , \1714_b0 );
or ( \1716_b1 , \1713_b1 , w_5368 );
or ( \1716_b0 , \1713_b0 , \1715_b0 );
not ( \1715_b0 , w_5369 );
and ( w_5369 , w_5368 , \1715_b1 );
or ( \1717_b1 , \1552_b1 , w_5371 );
not ( w_5371 , w_5372 );
and ( \1717_b0 , \1552_b0 , w_5373 );
and ( w_5372 ,  , w_5373 );
buf ( w_5371 , \1627_b1 );
not ( w_5371 , w_5374 );
not (  , w_5375 );
and ( w_5374 , w_5375 , \1627_b0 );
or ( \1718_b1 , \1716_b1 , w_5377 );
not ( w_5377 , w_5378 );
and ( \1718_b0 , \1716_b0 , w_5379 );
and ( w_5378 ,  , w_5379 );
buf ( w_5377 , \1717_b1 );
not ( w_5377 , w_5380 );
not (  , w_5381 );
and ( w_5380 , w_5381 , \1717_b0 );
or ( \1719_b1 , \a[2]_b1 , \d[11]_b1 );
xor ( \1719_b0 , \a[2]_b0 , w_5382 );
not ( w_5382 , w_5383 );
and ( w_5383 , \d[11]_b1 , \d[11]_b0 );
buf ( \1720_b1 , \1719_b1 );
not ( \1720_b1 , w_5384 );
not ( \1720_b0 , w_5385 );
and ( w_5384 , w_5385 , \1719_b0 );
or ( \1721_b1 , \1637_b1 , w_5387 );
not ( w_5387 , w_5388 );
and ( \1721_b0 , \1637_b0 , w_5389 );
and ( w_5388 ,  , w_5389 );
buf ( w_5387 , \1635_b1 );
not ( w_5387 , w_5390 );
not (  , w_5391 );
and ( w_5390 , w_5391 , \1635_b0 );
buf ( \1722_b1 , \1721_b1 );
not ( \1722_b1 , w_5392 );
not ( \1722_b0 , w_5393 );
and ( w_5392 , w_5393 , \1721_b0 );
or ( \1723_b1 , \1720_b1 , w_5394 );
or ( \1723_b0 , \1720_b0 , \1722_b0 );
not ( \1722_b0 , w_5395 );
and ( w_5395 , w_5394 , \1722_b1 );
or ( \1724_b1 , \1641_b1 , w_5397 );
not ( w_5397 , w_5398 );
and ( \1724_b0 , \1641_b0 , w_5399 );
and ( w_5398 ,  , w_5399 );
buf ( w_5397 , \1633_b1 );
not ( w_5397 , w_5400 );
not (  , w_5401 );
and ( w_5400 , w_5401 , \1633_b0 );
or ( \1725_b1 , \1723_b1 , w_5403 );
not ( w_5403 , w_5404 );
and ( \1725_b0 , \1723_b0 , w_5405 );
and ( w_5404 ,  , w_5405 );
buf ( w_5403 , \1724_b1 );
not ( w_5403 , w_5406 );
not (  , w_5407 );
and ( w_5406 , w_5407 , \1724_b0 );
or ( \1726_b1 , \1718_b1 , \1725_b1 );
xor ( \1726_b0 , \1718_b0 , w_5408 );
not ( w_5408 , w_5409 );
and ( w_5409 , \1725_b1 , \1725_b0 );
or ( \1727_b1 , \a[8]_b1 , \d[5]_b1 );
xor ( \1727_b0 , \a[8]_b0 , w_5410 );
not ( w_5410 , w_5411 );
and ( w_5411 , \d[5]_b1 , \d[5]_b0 );
buf ( \1728_b1 , \1727_b1 );
not ( \1728_b1 , w_5412 );
not ( \1728_b0 , w_5413 );
and ( w_5412 , w_5413 , \1727_b0 );
buf ( \1729_b1 , \1135_b1 );
not ( \1729_b1 , w_5414 );
not ( \1729_b0 , w_5415 );
and ( w_5414 , w_5415 , \1135_b0 );
or ( \1730_b1 , \1728_b1 , w_5416 );
or ( \1730_b0 , \1728_b0 , \1729_b0 );
not ( \1729_b0 , w_5417 );
and ( w_5417 , w_5416 , \1729_b1 );
or ( \1731_b1 , \951_b1 , w_5419 );
not ( w_5419 , w_5420 );
and ( \1731_b0 , \951_b0 , w_5421 );
and ( w_5420 ,  , w_5421 );
buf ( w_5419 , \1692_b1 );
not ( w_5419 , w_5422 );
not (  , w_5423 );
and ( w_5422 , w_5423 , \1692_b0 );
or ( \1732_b1 , \1730_b1 , w_5425 );
not ( w_5425 , w_5426 );
and ( \1732_b0 , \1730_b0 , w_5427 );
and ( w_5426 ,  , w_5427 );
buf ( w_5425 , \1731_b1 );
not ( w_5425 , w_5428 );
not (  , w_5429 );
and ( w_5428 , w_5429 , \1731_b0 );
or ( \1733_b1 , \1726_b1 , \1732_b1 );
not ( \1732_b1 , w_5430 );
and ( \1733_b0 , \1726_b0 , w_5431 );
and ( w_5430 , w_5431 , \1732_b0 );
or ( \1734_b1 , \1718_b1 , \1725_b1 );
not ( \1725_b1 , w_5432 );
and ( \1734_b0 , \1718_b0 , w_5433 );
and ( w_5432 , w_5433 , \1725_b0 );
or ( \1735_b1 , \1733_b1 , w_5434 );
or ( \1735_b0 , \1733_b0 , \1734_b0 );
not ( \1734_b0 , w_5435 );
and ( w_5435 , w_5434 , \1734_b1 );
or ( \1736_b1 , \1711_b1 , w_5436 );
or ( \1736_b0 , \1711_b0 , \1735_b0 );
not ( \1735_b0 , w_5437 );
and ( w_5437 , w_5436 , \1735_b1 );
or ( \1737_b1 , \a[4]_b1 , \d[9]_b1 );
xor ( \1737_b0 , \a[4]_b0 , w_5438 );
not ( w_5438 , w_5439 );
and ( w_5439 , \d[9]_b1 , \d[9]_b0 );
buf ( \1738_b1 , \1737_b1 );
not ( \1738_b1 , w_5440 );
not ( \1738_b0 , w_5441 );
and ( w_5440 , w_5441 , \1737_b0 );
buf ( \1739_b1 , \1542_b1 );
not ( \1739_b1 , w_5442 );
not ( \1739_b0 , w_5443 );
and ( w_5442 , w_5443 , \1542_b0 );
or ( \1740_b1 , \1738_b1 , w_5444 );
or ( \1740_b0 , \1738_b0 , \1739_b0 );
not ( \1739_b0 , w_5445 );
and ( w_5445 , w_5444 , \1739_b1 );
or ( \1741_b1 , \1545_b1 , w_5447 );
not ( w_5447 , w_5448 );
and ( \1741_b0 , \1545_b0 , w_5449 );
and ( w_5448 ,  , w_5449 );
buf ( w_5447 , \1685_b1 );
not ( w_5447 , w_5450 );
not (  , w_5451 );
and ( w_5450 , w_5451 , \1685_b0 );
or ( \1742_b1 , \1740_b1 , w_5453 );
not ( w_5453 , w_5454 );
and ( \1742_b0 , \1740_b0 , w_5455 );
and ( w_5454 ,  , w_5455 );
buf ( w_5453 , \1741_b1 );
not ( w_5453 , w_5456 );
not (  , w_5457 );
and ( w_5456 , w_5457 , \1741_b0 );
buf ( \1743_b1 , \1742_b1 );
not ( \1743_b1 , w_5458 );
not ( \1743_b0 , w_5459 );
and ( w_5458 , w_5459 , \1742_b0 );
or ( \1744_b1 , \a[10]_b1 , \d[3]_b1 );
xor ( \1744_b0 , \a[10]_b0 , w_5460 );
not ( w_5460 , w_5461 );
and ( w_5461 , \d[3]_b1 , \d[3]_b0 );
buf ( \1745_b1 , \1744_b1 );
not ( \1745_b1 , w_5462 );
not ( \1745_b0 , w_5463 );
and ( w_5462 , w_5463 , \1744_b0 );
buf ( \1746_b1 , \1067_b1 );
not ( \1746_b1 , w_5464 );
not ( \1746_b0 , w_5465 );
and ( w_5464 , w_5465 , \1067_b0 );
or ( \1747_b1 , \1745_b1 , w_5466 );
or ( \1747_b0 , \1745_b0 , \1746_b0 );
not ( \1746_b0 , w_5467 );
and ( w_5467 , w_5466 , \1746_b1 );
or ( \1748_b1 , \976_b1 , w_5469 );
not ( w_5469 , w_5470 );
and ( \1748_b0 , \976_b0 , w_5471 );
and ( w_5470 ,  , w_5471 );
buf ( w_5469 , \1580_b1 );
not ( w_5469 , w_5472 );
not (  , w_5473 );
and ( w_5472 , w_5473 , \1580_b0 );
or ( \1749_b1 , \1747_b1 , w_5475 );
not ( w_5475 , w_5476 );
and ( \1749_b0 , \1747_b0 , w_5477 );
and ( w_5476 ,  , w_5477 );
buf ( w_5475 , \1748_b1 );
not ( w_5475 , w_5478 );
not (  , w_5479 );
and ( w_5478 , w_5479 , \1748_b0 );
buf ( \1750_b1 , \1749_b1 );
not ( \1750_b1 , w_5480 );
not ( \1750_b0 , w_5481 );
and ( w_5480 , w_5481 , \1749_b0 );
or ( \1751_b1 , \1743_b1 , w_5482 );
or ( \1751_b0 , \1743_b0 , \1750_b0 );
not ( \1750_b0 , w_5483 );
and ( w_5483 , w_5482 , \1750_b1 );
or ( \1752_b1 , \1749_b1 , w_5484 );
or ( \1752_b0 , \1749_b0 , \1742_b0 );
not ( \1742_b0 , w_5485 );
and ( w_5485 , w_5484 , \1742_b1 );
buf ( \1753_b1 , \1679_b1 );
not ( \1753_b1 , w_5486 );
not ( \1753_b0 , w_5487 );
and ( w_5486 , w_5487 , \1679_b0 );
buf ( \1754_b1 , \958_b1 );
not ( \1754_b1 , w_5488 );
not ( \1754_b0 , w_5489 );
and ( w_5488 , w_5489 , \958_b0 );
or ( \1755_b1 , \1753_b1 , w_5490 );
or ( \1755_b0 , \1753_b0 , \1754_b0 );
not ( \1754_b0 , w_5491 );
and ( w_5491 , w_5490 , \1754_b1 );
or ( \1756_b1 , \a[6]_b1 , \d[7]_b1 );
xor ( \1756_b0 , \a[6]_b0 , w_5492 );
not ( w_5492 , w_5493 );
and ( w_5493 , \d[7]_b1 , \d[7]_b0 );
or ( \1757_b1 , \1127_b1 , w_5495 );
not ( w_5495 , w_5496 );
and ( \1757_b0 , \1127_b0 , w_5497 );
and ( w_5496 ,  , w_5497 );
buf ( w_5495 , \1756_b1 );
not ( w_5495 , w_5498 );
not (  , w_5499 );
and ( w_5498 , w_5499 , \1756_b0 );
or ( \1758_b1 , \1755_b1 , w_5501 );
not ( w_5501 , w_5502 );
and ( \1758_b0 , \1755_b0 , w_5503 );
and ( w_5502 ,  , w_5503 );
buf ( w_5501 , \1757_b1 );
not ( w_5501 , w_5504 );
not (  , w_5505 );
and ( w_5504 , w_5505 , \1757_b0 );
or ( \1759_b1 , \1752_b1 , w_5507 );
not ( w_5507 , w_5508 );
and ( \1759_b0 , \1752_b0 , w_5509 );
and ( w_5508 ,  , w_5509 );
buf ( w_5507 , \1758_b1 );
not ( w_5507 , w_5510 );
not (  , w_5511 );
and ( w_5510 , w_5511 , \1758_b0 );
or ( \1760_b1 , \1751_b1 , w_5513 );
not ( w_5513 , w_5514 );
and ( \1760_b0 , \1751_b0 , w_5515 );
and ( w_5514 ,  , w_5515 );
buf ( w_5513 , \1759_b1 );
not ( w_5513 , w_5516 );
not (  , w_5517 );
and ( w_5516 , w_5517 , \1759_b0 );
or ( \1761_b1 , \1736_b1 , w_5519 );
not ( w_5519 , w_5520 );
and ( \1761_b0 , \1736_b0 , w_5521 );
and ( w_5520 ,  , w_5521 );
buf ( w_5519 , \1760_b1 );
not ( w_5519 , w_5522 );
not (  , w_5523 );
and ( w_5522 , w_5523 , \1760_b0 );
or ( \1762_b1 , \1711_b1 , w_5525 );
not ( w_5525 , w_5526 );
and ( \1762_b0 , \1711_b0 , w_5527 );
and ( w_5526 ,  , w_5527 );
buf ( w_5525 , \1735_b1 );
not ( w_5525 , w_5528 );
not (  , w_5529 );
and ( w_5528 , w_5529 , \1735_b0 );
or ( \1763_b1 , \1761_b1 , w_5531 );
not ( w_5531 , w_5532 );
and ( \1763_b0 , \1761_b0 , w_5533 );
and ( w_5532 ,  , w_5533 );
buf ( w_5531 , \1762_b1 );
not ( w_5531 , w_5534 );
not (  , w_5535 );
and ( w_5534 , w_5535 , \1762_b0 );
buf ( \1764_b1 , \1763_b1 );
not ( \1764_b1 , w_5536 );
not ( \1764_b0 , w_5537 );
and ( w_5536 , w_5537 , \1763_b0 );
or ( \1765_b1 , \1709_b1 , \1764_b1 );
not ( \1764_b1 , w_5538 );
and ( \1765_b0 , \1709_b0 , w_5539 );
and ( w_5538 , w_5539 , \1764_b0 );
buf ( \1766_b1 , \1709_b1 );
not ( \1766_b1 , w_5540 );
not ( \1766_b0 , w_5541 );
and ( w_5540 , w_5541 , \1709_b0 );
or ( \1767_b1 , \1766_b1 , \1763_b1 );
not ( \1763_b1 , w_5542 );
and ( \1767_b0 , \1766_b0 , w_5543 );
and ( w_5542 , w_5543 , \1763_b0 );
or ( \1768_b1 , \1765_b1 , w_5545 );
not ( w_5545 , w_5546 );
and ( \1768_b0 , \1765_b0 , w_5547 );
and ( w_5546 ,  , w_5547 );
buf ( w_5545 , \1767_b1 );
not ( w_5545 , w_5548 );
not (  , w_5549 );
and ( w_5548 , w_5549 , \1767_b0 );
or ( \1769_b1 , \1684_b1 , \1690_b1 );
xor ( \1769_b0 , \1684_b0 , w_5550 );
not ( w_5550 , w_5551 );
and ( w_5551 , \1690_b1 , \1690_b0 );
or ( \1770_b1 , \1769_b1 , \1697_b1 );
xor ( \1770_b0 , \1769_b0 , w_5552 );
not ( w_5552 , w_5553 );
and ( w_5553 , \1697_b1 , \1697_b0 );
or ( \1771_b1 , \1632_b1 , \1644_b1 );
xor ( \1771_b0 , \1632_b0 , w_5554 );
not ( w_5554 , w_5555 );
and ( w_5555 , \1644_b1 , \1644_b0 );
or ( \1772_b1 , \1771_b1 , \1656_b1 );
xor ( \1772_b0 , \1771_b0 , w_5556 );
not ( w_5556 , w_5557 );
and ( w_5557 , \1656_b1 , \1656_b0 );
or ( \1773_b1 , \1770_b1 , \1772_b1 );
xor ( \1773_b0 , \1770_b0 , w_5558 );
not ( w_5558 , w_5559 );
and ( w_5559 , \1772_b1 , \1772_b0 );
or ( \1774_b1 , \1552_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_5560 );
and ( \1774_b0 , \1552_b0 , w_5561 );
and ( w_5560 , w_5561 , \a[0]_b0 );
or ( \1775_b1 , \d[7]_b1 , \a[5]_b1 );
xor ( \1775_b0 , \d[7]_b0 , w_5562 );
not ( w_5562 , w_5563 );
and ( w_5563 , \a[5]_b1 , \a[5]_b0 );
buf ( \1776_b1 , \1775_b1 );
not ( \1776_b1 , w_5564 );
not ( \1776_b0 , w_5565 );
and ( w_5564 , w_5565 , \1775_b0 );
buf ( \1777_b1 , \1127_b1 );
not ( \1777_b1 , w_5566 );
not ( \1777_b0 , w_5567 );
and ( w_5566 , w_5567 , \1127_b0 );
or ( \1778_b1 , \1776_b1 , w_5568 );
or ( \1778_b0 , \1776_b0 , \1777_b0 );
not ( \1777_b0 , w_5569 );
and ( w_5569 , w_5568 , \1777_b1 );
or ( \1779_b1 , \958_b1 , w_5571 );
not ( w_5571 , w_5572 );
and ( \1779_b0 , \958_b0 , w_5573 );
and ( w_5572 ,  , w_5573 );
buf ( w_5571 , \1756_b1 );
not ( w_5571 , w_5574 );
not (  , w_5575 );
and ( w_5574 , w_5575 , \1756_b0 );
or ( \1780_b1 , \1778_b1 , w_5577 );
not ( w_5577 , w_5578 );
and ( \1780_b0 , \1778_b0 , w_5579 );
and ( w_5578 ,  , w_5579 );
buf ( w_5577 , \1779_b1 );
not ( w_5577 , w_5580 );
not (  , w_5581 );
and ( w_5580 , w_5581 , \1779_b0 );
or ( \1781_b1 , \1774_b1 , \1780_b1 );
xor ( \1781_b0 , \1774_b0 , w_5582 );
not ( w_5582 , w_5583 );
and ( w_5583 , \1780_b1 , \1780_b0 );
or ( \1782_b1 , \a[9]_b1 , \d[3]_b1 );
xor ( \1782_b0 , \a[9]_b0 , w_5584 );
not ( w_5584 , w_5585 );
and ( w_5585 , \d[3]_b1 , \d[3]_b0 );
buf ( \1783_b1 , \1782_b1 );
not ( \1783_b1 , w_5586 );
not ( \1783_b0 , w_5587 );
and ( w_5586 , w_5587 , \1782_b0 );
buf ( \1784_b1 , \973_b1 );
not ( \1784_b1 , w_5588 );
not ( \1784_b0 , w_5589 );
and ( w_5588 , w_5589 , \973_b0 );
or ( \1785_b1 , \1783_b1 , w_5590 );
or ( \1785_b0 , \1783_b0 , \1784_b0 );
not ( \1784_b0 , w_5591 );
and ( w_5591 , w_5590 , \1784_b1 );
or ( \1786_b1 , \976_b1 , w_5593 );
not ( w_5593 , w_5594 );
and ( \1786_b0 , \976_b0 , w_5595 );
and ( w_5594 ,  , w_5595 );
buf ( w_5593 , \1744_b1 );
not ( w_5593 , w_5596 );
not (  , w_5597 );
and ( w_5596 , w_5597 , \1744_b0 );
or ( \1787_b1 , \1785_b1 , w_5599 );
not ( w_5599 , w_5600 );
and ( \1787_b0 , \1785_b0 , w_5601 );
and ( w_5600 ,  , w_5601 );
buf ( w_5599 , \1786_b1 );
not ( w_5599 , w_5602 );
not (  , w_5603 );
and ( w_5602 , w_5603 , \1786_b0 );
or ( \1788_b1 , \1781_b1 , \1787_b1 );
not ( \1787_b1 , w_5604 );
and ( \1788_b0 , \1781_b0 , w_5605 );
and ( w_5604 , w_5605 , \1787_b0 );
or ( \1789_b1 , \1774_b1 , \1780_b1 );
not ( \1780_b1 , w_5606 );
and ( \1789_b0 , \1774_b0 , w_5607 );
and ( w_5606 , w_5607 , \1780_b0 );
or ( \1790_b1 , \1788_b1 , w_5608 );
or ( \1790_b0 , \1788_b0 , \1789_b0 );
not ( \1789_b0 , w_5609 );
and ( w_5609 , w_5608 , \1789_b1 );
or ( \1791_b1 , \1649_b1 , \1655_b1 );
xor ( \1791_b0 , \1649_b0 , w_5610 );
not ( w_5610 , w_5611 );
and ( w_5611 , \1655_b1 , \1655_b0 );
or ( \1792_b1 , \1790_b1 , w_5612 );
or ( \1792_b0 , \1790_b0 , \1791_b0 );
not ( \1791_b0 , w_5613 );
and ( w_5613 , w_5612 , \1791_b1 );
or ( \1793_b1 , \a[11]_b1 , \d[1]_b1 );
xor ( \1793_b0 , \a[11]_b0 , w_5614 );
not ( w_5614 , w_5615 );
and ( w_5615 , \d[1]_b1 , \d[1]_b0 );
buf ( \1794_b1 , \1793_b1 );
not ( \1794_b1 , w_5616 );
not ( \1794_b0 , w_5617 );
and ( w_5616 , w_5617 , \1793_b0 );
buf ( \1795_b1 , \932_b1 );
not ( \1795_b1 , w_5618 );
not ( \1795_b0 , w_5619 );
and ( w_5618 , w_5619 , \932_b0 );
or ( \1796_b1 , \1794_b1 , w_5620 );
or ( \1796_b0 , \1794_b0 , \1795_b0 );
not ( \1795_b0 , w_5621 );
and ( w_5621 , w_5620 , \1795_b1 );
or ( \1797_b1 , \1650_b1 , w_5623 );
not ( w_5623 , w_5624 );
and ( \1797_b0 , \1650_b0 , w_5625 );
and ( w_5624 ,  , w_5625 );
buf ( w_5623 , \d[0]_b1 );
not ( w_5623 , w_5626 );
not (  , w_5627 );
and ( w_5626 , w_5627 , \d[0]_b0 );
or ( \1798_b1 , \1796_b1 , w_5629 );
not ( w_5629 , w_5630 );
and ( \1798_b0 , \1796_b0 , w_5631 );
and ( w_5630 ,  , w_5631 );
buf ( w_5629 , \1797_b1 );
not ( w_5629 , w_5632 );
not (  , w_5633 );
and ( w_5632 , w_5633 , \1797_b0 );
or ( \1799_b1 , \a[3]_b1 , \d[9]_b1 );
xor ( \1799_b0 , \a[3]_b0 , w_5634 );
not ( w_5634 , w_5635 );
and ( w_5635 , \d[9]_b1 , \d[9]_b0 );
buf ( \1800_b1 , \1799_b1 );
not ( \1800_b1 , w_5636 );
not ( \1800_b0 , w_5637 );
and ( w_5636 , w_5637 , \1799_b0 );
buf ( \1801_b1 , \1542_b1 );
not ( \1801_b1 , w_5638 );
not ( \1801_b0 , w_5639 );
and ( w_5638 , w_5639 , \1542_b0 );
or ( \1802_b1 , \1800_b1 , w_5640 );
or ( \1802_b0 , \1800_b0 , \1801_b0 );
not ( \1801_b0 , w_5641 );
and ( w_5641 , w_5640 , \1801_b1 );
or ( \1803_b1 , \1545_b1 , w_5643 );
not ( w_5643 , w_5644 );
and ( \1803_b0 , \1545_b0 , w_5645 );
and ( w_5644 ,  , w_5645 );
buf ( w_5643 , \1737_b1 );
not ( w_5643 , w_5646 );
not (  , w_5647 );
and ( w_5646 , w_5647 , \1737_b0 );
or ( \1804_b1 , \1802_b1 , w_5649 );
not ( w_5649 , w_5650 );
and ( \1804_b0 , \1802_b0 , w_5651 );
and ( w_5650 ,  , w_5651 );
buf ( w_5649 , \1803_b1 );
not ( w_5649 , w_5652 );
not (  , w_5653 );
and ( w_5652 , w_5653 , \1803_b0 );
or ( \1805_b1 , \1798_b1 , \1804_b1 );
xor ( \1805_b0 , \1798_b0 , w_5654 );
not ( w_5654 , w_5655 );
and ( w_5655 , \1804_b1 , \1804_b0 );
or ( \1806_b1 , \a[1]_b1 , \d[11]_b1 );
xor ( \1806_b0 , \a[1]_b0 , w_5656 );
not ( w_5656 , w_5657 );
and ( w_5657 , \d[11]_b1 , \d[11]_b0 );
buf ( \1807_b1 , \1806_b1 );
not ( \1807_b1 , w_5658 );
not ( \1807_b0 , w_5659 );
and ( w_5658 , w_5659 , \1806_b0 );
buf ( \1808_b1 , \1721_b1 );
not ( \1808_b1 , w_5660 );
not ( \1808_b0 , w_5661 );
and ( w_5660 , w_5661 , \1721_b0 );
or ( \1809_b1 , \1807_b1 , w_5662 );
or ( \1809_b0 , \1807_b0 , \1808_b0 );
not ( \1808_b0 , w_5663 );
and ( w_5663 , w_5662 , \1808_b1 );
or ( \1810_b1 , \1641_b1 , w_5665 );
not ( w_5665 , w_5666 );
and ( \1810_b0 , \1641_b0 , w_5667 );
and ( w_5666 ,  , w_5667 );
buf ( w_5665 , \1719_b1 );
not ( w_5665 , w_5668 );
not (  , w_5669 );
and ( w_5668 , w_5669 , \1719_b0 );
or ( \1811_b1 , \1809_b1 , w_5671 );
not ( w_5671 , w_5672 );
and ( \1811_b0 , \1809_b0 , w_5673 );
and ( w_5672 ,  , w_5673 );
buf ( w_5671 , \1810_b1 );
not ( w_5671 , w_5674 );
not (  , w_5675 );
and ( w_5674 , w_5675 , \1810_b0 );
or ( \1812_b1 , \1805_b1 , \1811_b1 );
not ( \1811_b1 , w_5676 );
and ( \1812_b0 , \1805_b0 , w_5677 );
and ( w_5676 , w_5677 , \1811_b0 );
or ( \1813_b1 , \1798_b1 , \1804_b1 );
not ( \1804_b1 , w_5678 );
and ( \1813_b0 , \1798_b0 , w_5679 );
and ( w_5678 , w_5679 , \1804_b0 );
or ( \1814_b1 , \1812_b1 , w_5680 );
or ( \1814_b0 , \1812_b0 , \1813_b0 );
not ( \1813_b0 , w_5681 );
and ( w_5681 , w_5680 , \1813_b1 );
or ( \1815_b1 , \1792_b1 , w_5683 );
not ( w_5683 , w_5684 );
and ( \1815_b0 , \1792_b0 , w_5685 );
and ( w_5684 ,  , w_5685 );
buf ( w_5683 , \1814_b1 );
not ( w_5683 , w_5686 );
not (  , w_5687 );
and ( w_5686 , w_5687 , \1814_b0 );
or ( \1816_b1 , \1790_b1 , w_5689 );
not ( w_5689 , w_5690 );
and ( \1816_b0 , \1790_b0 , w_5691 );
and ( w_5690 ,  , w_5691 );
buf ( w_5689 , \1791_b1 );
not ( w_5689 , w_5692 );
not (  , w_5693 );
and ( w_5692 , w_5693 , \1791_b0 );
or ( \1817_b1 , \1815_b1 , w_5695 );
not ( w_5695 , w_5696 );
and ( \1817_b0 , \1815_b0 , w_5697 );
and ( w_5696 ,  , w_5697 );
buf ( w_5695 , \1816_b1 );
not ( w_5695 , w_5698 );
not (  , w_5699 );
and ( w_5698 , w_5699 , \1816_b0 );
or ( \1818_b1 , \1773_b1 , \1817_b1 );
not ( \1817_b1 , w_5700 );
and ( \1818_b0 , \1773_b0 , w_5701 );
and ( w_5700 , w_5701 , \1817_b0 );
or ( \1819_b1 , \1770_b1 , \1772_b1 );
not ( \1772_b1 , w_5702 );
and ( \1819_b0 , \1770_b0 , w_5703 );
and ( w_5702 , w_5703 , \1772_b0 );
or ( \1820_b1 , \1818_b1 , w_5704 );
or ( \1820_b0 , \1818_b0 , \1819_b0 );
not ( \1819_b0 , w_5705 );
and ( w_5705 , w_5704 , \1819_b1 );
buf ( \1821_b1 , \1820_b1 );
not ( \1821_b1 , w_5706 );
not ( \1821_b0 , w_5707 );
and ( w_5706 , w_5707 , \1820_b0 );
or ( \1822_b1 , \1768_b1 , \1821_b1 );
not ( \1821_b1 , w_5708 );
and ( \1822_b0 , \1768_b0 , w_5709 );
and ( w_5708 , w_5709 , \1821_b0 );
buf ( \1823_b1 , \1768_b1 );
not ( \1823_b1 , w_5710 );
not ( \1823_b0 , w_5711 );
and ( w_5710 , w_5711 , \1768_b0 );
or ( \1824_b1 , \1823_b1 , \1820_b1 );
not ( \1820_b1 , w_5712 );
and ( \1824_b0 , \1823_b0 , w_5713 );
and ( w_5712 , w_5713 , \1820_b0 );
or ( \1825_b1 , \1822_b1 , w_5715 );
not ( w_5715 , w_5716 );
and ( \1825_b0 , \1822_b0 , w_5717 );
and ( w_5716 ,  , w_5717 );
buf ( w_5715 , \1824_b1 );
not ( w_5715 , w_5718 );
not (  , w_5719 );
and ( w_5718 , w_5719 , \1824_b0 );
or ( \1826_b1 , \1735_b1 , \1711_b1 );
xor ( \1826_b0 , \1735_b0 , w_5720 );
not ( w_5720 , w_5721 );
and ( w_5721 , \1711_b1 , \1711_b0 );
or ( \1827_b1 , \1826_b1 , w_5722 );
xor ( \1827_b0 , \1826_b0 , w_5724 );
not ( w_5724 , w_5725 );
and ( w_5725 , w_5722 , w_5723 );
buf ( w_5722 , \1760_b1 );
not ( w_5722 , w_5726 );
not ( w_5723 , w_5727 );
and ( w_5726 , w_5727 , \1760_b0 );
buf ( \1828_b1 , \1827_b1 );
not ( \1828_b1 , w_5728 );
not ( \1828_b0 , w_5729 );
and ( w_5728 , w_5729 , \1827_b0 );
buf ( \1829_b1 , \1828_b1 );
not ( \1829_b1 , w_5730 );
not ( \1829_b0 , w_5731 );
and ( w_5730 , w_5731 , \1828_b0 );
or ( \1830_b1 , \1770_b1 , \1772_b1 );
xor ( \1830_b0 , \1770_b0 , w_5732 );
not ( w_5732 , w_5733 );
and ( w_5733 , \1772_b1 , \1772_b0 );
or ( \1831_b1 , \1830_b1 , \1817_b1 );
xor ( \1831_b0 , \1830_b0 , w_5734 );
not ( w_5734 , w_5735 );
and ( w_5735 , \1817_b1 , \1817_b0 );
buf ( \1832_b1 , \1831_b1 );
not ( \1832_b1 , w_5736 );
not ( \1832_b0 , w_5737 );
and ( w_5736 , w_5737 , \1831_b0 );
or ( \1833_b1 , \1829_b1 , w_5738 );
or ( \1833_b0 , \1829_b0 , \1832_b0 );
not ( \1832_b0 , w_5739 );
and ( w_5739 , w_5738 , \1832_b1 );
or ( \1834_b1 , \1831_b1 , w_5740 );
or ( \1834_b0 , \1831_b0 , \1828_b0 );
not ( \1828_b0 , w_5741 );
and ( w_5741 , w_5740 , \1828_b1 );
or ( \1835_b1 , \1718_b1 , \1725_b1 );
xor ( \1835_b0 , \1718_b0 , w_5742 );
not ( w_5742 , w_5743 );
and ( w_5743 , \1725_b1 , \1725_b0 );
or ( \1836_b1 , \1835_b1 , \1732_b1 );
xor ( \1836_b0 , \1835_b0 , w_5744 );
not ( w_5744 , w_5745 );
and ( w_5745 , \1732_b1 , \1732_b0 );
buf ( \1837_b1 , \1836_b1 );
not ( \1837_b1 , w_5746 );
not ( \1837_b0 , w_5747 );
and ( w_5746 , w_5747 , \1836_b0 );
or ( \1838_b1 , \1742_b1 , \1758_b1 );
xor ( \1838_b0 , \1742_b0 , w_5748 );
not ( w_5748 , w_5749 );
and ( w_5749 , \1758_b1 , \1758_b0 );
or ( \1839_b1 , \1838_b1 , w_5750 );
xor ( \1839_b0 , \1838_b0 , w_5752 );
not ( w_5752 , w_5753 );
and ( w_5753 , w_5750 , w_5751 );
buf ( w_5750 , \1749_b1 );
not ( w_5750 , w_5754 );
not ( w_5751 , w_5755 );
and ( w_5754 , w_5755 , \1749_b0 );
or ( \1840_b1 , \1837_b1 , w_5757 );
not ( w_5757 , w_5758 );
and ( \1840_b0 , \1837_b0 , w_5759 );
and ( w_5758 ,  , w_5759 );
buf ( w_5757 , \1839_b1 );
not ( w_5757 , w_5760 );
not (  , w_5761 );
and ( w_5760 , w_5761 , \1839_b0 );
buf ( \1841_b1 , \1840_b1 );
not ( \1841_b1 , w_5762 );
not ( \1841_b0 , w_5763 );
and ( w_5762 , w_5763 , \1840_b0 );
or ( \1842_b1 , \a[7]_b1 , \d[5]_b1 );
xor ( \1842_b0 , \a[7]_b0 , w_5764 );
not ( w_5764 , w_5765 );
and ( w_5765 , \d[5]_b1 , \d[5]_b0 );
buf ( \1843_b1 , \1842_b1 );
not ( \1843_b1 , w_5766 );
not ( \1843_b0 , w_5767 );
and ( w_5766 , w_5767 , \1842_b0 );
buf ( \1844_b1 , \1135_b1 );
not ( \1844_b1 , w_5768 );
not ( \1844_b0 , w_5769 );
and ( w_5768 , w_5769 , \1135_b0 );
or ( \1845_b1 , \1843_b1 , w_5770 );
or ( \1845_b0 , \1843_b0 , \1844_b0 );
not ( \1844_b0 , w_5771 );
and ( w_5771 , w_5770 , \1844_b1 );
or ( \1846_b1 , \951_b1 , w_5773 );
not ( w_5773 , w_5774 );
and ( \1846_b0 , \951_b0 , w_5775 );
and ( w_5774 ,  , w_5775 );
buf ( w_5773 , \1727_b1 );
not ( w_5773 , w_5776 );
not (  , w_5777 );
and ( w_5776 , w_5777 , \1727_b0 );
or ( \1847_b1 , \1845_b1 , w_5779 );
not ( w_5779 , w_5780 );
and ( \1847_b0 , \1845_b0 , w_5781 );
and ( w_5780 ,  , w_5781 );
buf ( w_5779 , \1846_b1 );
not ( w_5779 , w_5782 );
not (  , w_5783 );
and ( w_5782 , w_5783 , \1846_b0 );
buf ( \1848_b1 , \1847_b1 );
not ( \1848_b1 , w_5784 );
not ( \1848_b0 , w_5785 );
and ( w_5784 , w_5785 , \1847_b0 );
buf ( \1849_b1 , \1848_b1 );
not ( \1849_b1 , w_5786 );
not ( \1849_b0 , w_5787 );
and ( w_5786 , w_5787 , \1848_b0 );
or ( \1850_b1 , \a[8]_b1 , \d[3]_b1 );
xor ( \1850_b0 , \a[8]_b0 , w_5788 );
not ( w_5788 , w_5789 );
and ( w_5789 , \d[3]_b1 , \d[3]_b0 );
buf ( \1851_b1 , \1850_b1 );
not ( \1851_b1 , w_5790 );
not ( \1851_b0 , w_5791 );
and ( w_5790 , w_5791 , \1850_b0 );
buf ( \1852_b1 , \973_b1 );
not ( \1852_b1 , w_5792 );
not ( \1852_b0 , w_5793 );
and ( w_5792 , w_5793 , \973_b0 );
or ( \1853_b1 , \1851_b1 , w_5794 );
or ( \1853_b0 , \1851_b0 , \1852_b0 );
not ( \1852_b0 , w_5795 );
and ( w_5795 , w_5794 , \1852_b1 );
or ( \1854_b1 , \976_b1 , w_5797 );
not ( w_5797 , w_5798 );
and ( \1854_b0 , \976_b0 , w_5799 );
and ( w_5798 ,  , w_5799 );
buf ( w_5797 , \1782_b1 );
not ( w_5797 , w_5800 );
not (  , w_5801 );
and ( w_5800 , w_5801 , \1782_b0 );
or ( \1855_b1 , \1853_b1 , w_5803 );
not ( w_5803 , w_5804 );
and ( \1855_b0 , \1853_b0 , w_5805 );
and ( w_5804 ,  , w_5805 );
buf ( w_5803 , \1854_b1 );
not ( w_5803 , w_5806 );
not (  , w_5807 );
and ( w_5806 , w_5807 , \1854_b0 );
or ( \1856_b1 , \a[0]_b1 , w_5808 );
or ( \1856_b0 , \a[0]_b0 , \d[10]_b0 );
not ( \d[10]_b0 , w_5809 );
and ( w_5809 , w_5808 , \d[10]_b1 );
or ( \1857_b1 , \1856_b1 , w_5811 );
not ( w_5811 , w_5812 );
and ( \1857_b0 , \1856_b0 , w_5813 );
and ( w_5812 ,  , w_5813 );
buf ( w_5811 , \d[9]_b1 );
not ( w_5811 , w_5814 );
not (  , w_5815 );
and ( w_5814 , w_5815 , \d[9]_b0 );
or ( \1858_b1 , \a[0]_b1 , w_5817 );
not ( w_5817 , w_5818 );
and ( \1858_b0 , \a[0]_b0 , w_5819 );
and ( w_5818 ,  , w_5819 );
buf ( w_5817 , \d[10]_b1 );
not ( w_5817 , w_5820 );
not (  , w_5821 );
and ( w_5820 , w_5821 , \d[10]_b0 );
buf ( \1860_b1 , \1859_b1 );
not ( \1860_b1 , w_5822 );
not ( \1860_b0 , w_5823 );
and ( w_5822 , w_5823 , \1859_b0 );
or ( \1861_b1 , \1855_b1 , w_5825 );
not ( w_5825 , w_5826 );
and ( \1861_b0 , \1855_b0 , w_5827 );
and ( w_5826 ,  , w_5827 );
buf ( w_5825 , \1860_b1 );
not ( w_5825 , w_5828 );
not (  , w_5829 );
and ( w_5828 , w_5829 , \1860_b0 );
buf ( \1862_b1 , \1861_b1 );
not ( \1862_b1 , w_5830 );
not ( \1862_b0 , w_5831 );
and ( w_5830 , w_5831 , \1861_b0 );
or ( \1863_b1 , \1849_b1 , w_5832 );
or ( \1863_b0 , \1849_b0 , \1862_b0 );
not ( \1862_b0 , w_5833 );
and ( w_5833 , w_5832 , \1862_b1 );
or ( \1864_b1 , \a[10]_b1 , \d[1]_b1 );
xor ( \1864_b0 , \a[10]_b0 , w_5834 );
not ( w_5834 , w_5835 );
and ( w_5835 , \d[1]_b1 , \d[1]_b0 );
buf ( \1865_b1 , \1864_b1 );
not ( \1865_b1 , w_5836 );
not ( \1865_b0 , w_5837 );
and ( w_5836 , w_5837 , \1864_b0 );
buf ( \1866_b1 , \932_b1 );
not ( \1866_b1 , w_5838 );
not ( \1866_b0 , w_5839 );
and ( w_5838 , w_5839 , \932_b0 );
or ( \1867_b1 , \1865_b1 , w_5840 );
or ( \1867_b0 , \1865_b0 , \1866_b0 );
not ( \1866_b0 , w_5841 );
and ( w_5841 , w_5840 , \1866_b1 );
or ( \1868_b1 , \1793_b1 , w_5843 );
not ( w_5843 , w_5844 );
and ( \1868_b0 , \1793_b0 , w_5845 );
and ( w_5844 ,  , w_5845 );
buf ( w_5843 , \d[0]_b1 );
not ( w_5843 , w_5846 );
not (  , w_5847 );
and ( w_5846 , w_5847 , \d[0]_b0 );
or ( \1869_b1 , \1867_b1 , w_5849 );
not ( w_5849 , w_5850 );
and ( \1869_b0 , \1867_b0 , w_5851 );
and ( w_5850 ,  , w_5851 );
buf ( w_5849 , \1868_b1 );
not ( w_5849 , w_5852 );
not (  , w_5853 );
and ( w_5852 , w_5853 , \1868_b0 );
buf ( \1870_b1 , \1869_b1 );
not ( \1870_b1 , w_5854 );
not ( \1870_b0 , w_5855 );
and ( w_5854 , w_5855 , \1869_b0 );
or ( \1871_b1 , \d[9]_b1 , \a[2]_b1 );
xor ( \1871_b0 , \d[9]_b0 , w_5856 );
not ( w_5856 , w_5857 );
and ( w_5857 , \a[2]_b1 , \a[2]_b0 );
buf ( \1872_b1 , \1871_b1 );
not ( \1872_b1 , w_5858 );
not ( \1872_b0 , w_5859 );
and ( w_5858 , w_5859 , \1871_b0 );
buf ( \1873_b1 , \1542_b1 );
not ( \1873_b1 , w_5860 );
not ( \1873_b0 , w_5861 );
and ( w_5860 , w_5861 , \1542_b0 );
or ( \1874_b1 , \1872_b1 , w_5862 );
or ( \1874_b0 , \1872_b0 , \1873_b0 );
not ( \1873_b0 , w_5863 );
and ( w_5863 , w_5862 , \1873_b1 );
or ( \1875_b1 , \1545_b1 , w_5865 );
not ( w_5865 , w_5866 );
and ( \1875_b0 , \1545_b0 , w_5867 );
and ( w_5866 ,  , w_5867 );
buf ( w_5865 , \1799_b1 );
not ( w_5865 , w_5868 );
not (  , w_5869 );
and ( w_5868 , w_5869 , \1799_b0 );
or ( \1876_b1 , \1874_b1 , w_5871 );
not ( w_5871 , w_5872 );
and ( \1876_b0 , \1874_b0 , w_5873 );
and ( w_5872 ,  , w_5873 );
buf ( w_5871 , \1875_b1 );
not ( w_5871 , w_5874 );
not (  , w_5875 );
and ( w_5874 , w_5875 , \1875_b0 );
buf ( \1877_b1 , \1876_b1 );
not ( \1877_b1 , w_5876 );
not ( \1877_b0 , w_5877 );
and ( w_5876 , w_5877 , \1876_b0 );
or ( \1878_b1 , \1870_b1 , w_5878 );
or ( \1878_b0 , \1870_b0 , \1877_b0 );
not ( \1877_b0 , w_5879 );
and ( w_5879 , w_5878 , \1877_b1 );
or ( \1879_b1 , \1876_b1 , w_5880 );
or ( \1879_b0 , \1876_b0 , \1869_b0 );
not ( \1869_b0 , w_5881 );
and ( w_5881 , w_5880 , \1869_b1 );
or ( \1880_b1 , \d[7]_b1 , \a[4]_b1 );
xor ( \1880_b0 , \d[7]_b0 , w_5882 );
not ( w_5882 , w_5883 );
and ( w_5883 , \a[4]_b1 , \a[4]_b0 );
buf ( \1881_b1 , \1880_b1 );
not ( \1881_b1 , w_5884 );
not ( \1881_b0 , w_5885 );
and ( w_5884 , w_5885 , \1880_b0 );
or ( \1882_b1 , \d[7]_b1 , w_5886 );
xor ( \1882_b0 , \d[7]_b0 , w_5888 );
not ( w_5888 , w_5889 );
and ( w_5889 , w_5886 , w_5887 );
buf ( w_5886 , \d[6]_b1 );
not ( w_5886 , w_5890 );
not ( w_5887 , w_5891 );
and ( w_5890 , w_5891 , \d[6]_b0 );
or ( \1883_b1 , \1882_b1 , w_5893 );
not ( w_5893 , w_5894 );
and ( \1883_b0 , \1882_b0 , w_5895 );
and ( w_5894 ,  , w_5895 );
buf ( w_5893 , \957_b1 );
not ( w_5893 , w_5896 );
not (  , w_5897 );
and ( w_5896 , w_5897 , \957_b0 );
buf ( \1884_b1 , \1883_b1 );
not ( \1884_b1 , w_5898 );
not ( \1884_b0 , w_5899 );
and ( w_5898 , w_5899 , \1883_b0 );
or ( \1885_b1 , \1881_b1 , w_5900 );
or ( \1885_b0 , \1881_b0 , \1884_b0 );
not ( \1884_b0 , w_5901 );
and ( w_5901 , w_5900 , \1884_b1 );
or ( \1886_b1 , \1775_b1 , w_5903 );
not ( w_5903 , w_5904 );
and ( \1886_b0 , \1775_b0 , w_5905 );
and ( w_5904 ,  , w_5905 );
buf ( w_5903 , \957_b1 );
not ( w_5903 , w_5906 );
not (  , w_5907 );
and ( w_5906 , w_5907 , \957_b0 );
or ( \1887_b1 , \1885_b1 , w_5909 );
not ( w_5909 , w_5910 );
and ( \1887_b0 , \1885_b0 , w_5911 );
and ( w_5910 ,  , w_5911 );
buf ( w_5909 , \1886_b1 );
not ( w_5909 , w_5912 );
not (  , w_5913 );
and ( w_5912 , w_5913 , \1886_b0 );
or ( \1888_b1 , \1879_b1 , w_5915 );
not ( w_5915 , w_5916 );
and ( \1888_b0 , \1879_b0 , w_5917 );
and ( w_5916 ,  , w_5917 );
buf ( w_5915 , \1887_b1 );
not ( w_5915 , w_5918 );
not (  , w_5919 );
and ( w_5918 , w_5919 , \1887_b0 );
or ( \1889_b1 , \1878_b1 , w_5921 );
not ( w_5921 , w_5922 );
and ( \1889_b0 , \1878_b0 , w_5923 );
and ( w_5922 ,  , w_5923 );
buf ( w_5921 , \1888_b1 );
not ( w_5921 , w_5924 );
not (  , w_5925 );
and ( w_5924 , w_5925 , \1888_b0 );
or ( \1890_b1 , \1863_b1 , w_5927 );
not ( w_5927 , w_5928 );
and ( \1890_b0 , \1863_b0 , w_5929 );
and ( w_5928 ,  , w_5929 );
buf ( w_5927 , \1889_b1 );
not ( w_5927 , w_5930 );
not (  , w_5931 );
and ( w_5930 , w_5931 , \1889_b0 );
buf ( \1891_b1 , \1861_b1 );
not ( \1891_b1 , w_5932 );
not ( \1891_b0 , w_5933 );
and ( w_5932 , w_5933 , \1861_b0 );
or ( \1892_b1 , \1891_b1 , w_5935 );
not ( w_5935 , w_5936 );
and ( \1892_b0 , \1891_b0 , w_5937 );
and ( w_5936 ,  , w_5937 );
buf ( w_5935 , \1847_b1 );
not ( w_5935 , w_5938 );
not (  , w_5939 );
and ( w_5938 , w_5939 , \1847_b0 );
or ( \1893_b1 , \1890_b1 , w_5941 );
not ( w_5941 , w_5942 );
and ( \1893_b0 , \1890_b0 , w_5943 );
and ( w_5942 ,  , w_5943 );
buf ( w_5941 , \1892_b1 );
not ( w_5941 , w_5944 );
not (  , w_5945 );
and ( w_5944 , w_5945 , \1892_b0 );
buf ( \1894_b1 , \1893_b1 );
not ( \1894_b1 , w_5946 );
not ( \1894_b0 , w_5947 );
and ( w_5946 , w_5947 , \1893_b0 );
or ( \1895_b1 , \1841_b1 , w_5948 );
or ( \1895_b0 , \1841_b0 , \1894_b0 );
not ( \1894_b0 , w_5949 );
and ( w_5949 , w_5948 , \1894_b1 );
buf ( \1896_b1 , \1839_b1 );
not ( \1896_b1 , w_5950 );
not ( \1896_b0 , w_5951 );
and ( w_5950 , w_5951 , \1839_b0 );
or ( \1897_b1 , \1896_b1 , w_5953 );
not ( w_5953 , w_5954 );
and ( \1897_b0 , \1896_b0 , w_5955 );
and ( w_5954 ,  , w_5955 );
buf ( w_5953 , \1836_b1 );
not ( w_5953 , w_5956 );
not (  , w_5957 );
and ( w_5956 , w_5957 , \1836_b0 );
or ( \1898_b1 , \1895_b1 , w_5959 );
not ( w_5959 , w_5960 );
and ( \1898_b0 , \1895_b0 , w_5961 );
and ( w_5960 ,  , w_5961 );
buf ( w_5959 , \1897_b1 );
not ( w_5959 , w_5962 );
not (  , w_5963 );
and ( w_5962 , w_5963 , \1897_b0 );
or ( \1899_b1 , \1834_b1 , w_5965 );
not ( w_5965 , w_5966 );
and ( \1899_b0 , \1834_b0 , w_5967 );
and ( w_5966 ,  , w_5967 );
buf ( w_5965 , \1898_b1 );
not ( w_5965 , w_5968 );
not (  , w_5969 );
and ( w_5968 , w_5969 , \1898_b0 );
or ( \1900_b1 , \1833_b1 , w_5971 );
not ( w_5971 , w_5972 );
and ( \1900_b0 , \1833_b0 , w_5973 );
and ( w_5972 ,  , w_5973 );
buf ( w_5971 , \1899_b1 );
not ( w_5971 , w_5974 );
not (  , w_5975 );
and ( w_5974 , w_5975 , \1899_b0 );
or ( \1901_b1 , \1825_b1 , w_5976 );
xor ( \1901_b0 , \1825_b0 , w_5978 );
not ( w_5978 , w_5979 );
and ( w_5979 , w_5976 , w_5977 );
buf ( w_5976 , \1900_b1 );
not ( w_5976 , w_5980 );
not ( w_5977 , w_5981 );
and ( w_5980 , w_5981 , \1900_b0 );
buf ( \1902_b1 , \1901_b1 );
not ( \1902_b1 , w_5982 );
not ( \1902_b0 , w_5983 );
and ( w_5982 , w_5983 , \1901_b0 );
or ( \1903_b1 , \1831_b1 , w_5984 );
xor ( \1903_b0 , \1831_b0 , w_5986 );
not ( w_5986 , w_5987 );
and ( w_5987 , w_5984 , w_5985 );
buf ( w_5984 , \1827_b1 );
not ( w_5984 , w_5988 );
not ( w_5985 , w_5989 );
and ( w_5988 , w_5989 , \1827_b0 );
buf ( \1904_b1 , \1898_b1 );
not ( \1904_b1 , w_5990 );
not ( \1904_b0 , w_5991 );
and ( w_5990 , w_5991 , \1898_b0 );
or ( \1905_b1 , \1903_b1 , \1904_b1 );
not ( \1904_b1 , w_5992 );
and ( \1905_b0 , \1903_b0 , w_5993 );
and ( w_5992 , w_5993 , \1904_b0 );
buf ( \1906_b1 , \1903_b1 );
not ( \1906_b1 , w_5994 );
not ( \1906_b0 , w_5995 );
and ( w_5994 , w_5995 , \1903_b0 );
or ( \1907_b1 , \1906_b1 , \1898_b1 );
not ( \1898_b1 , w_5996 );
and ( \1907_b0 , \1906_b0 , w_5997 );
and ( w_5996 , w_5997 , \1898_b0 );
or ( \1908_b1 , \1905_b1 , w_5999 );
not ( w_5999 , w_6000 );
and ( \1908_b0 , \1905_b0 , w_6001 );
and ( w_6000 ,  , w_6001 );
buf ( w_5999 , \1907_b1 );
not ( w_5999 , w_6002 );
not (  , w_6003 );
and ( w_6002 , w_6003 , \1907_b0 );
or ( \1909_b1 , \1791_b1 , \1790_b1 );
xor ( \1909_b0 , \1791_b0 , w_6004 );
not ( w_6004 , w_6005 );
and ( w_6005 , \1790_b1 , \1790_b0 );
or ( \1910_b1 , \1909_b1 , w_6006 );
xor ( \1910_b0 , \1909_b0 , w_6008 );
not ( w_6008 , w_6009 );
and ( w_6009 , w_6006 , w_6007 );
buf ( w_6006 , \1814_b1 );
not ( w_6006 , w_6010 );
not ( w_6007 , w_6011 );
and ( w_6010 , w_6011 , \1814_b0 );
buf ( \1911_b1 , \1910_b1 );
not ( \1911_b1 , w_6012 );
not ( \1911_b0 , w_6013 );
and ( w_6012 , w_6013 , \1910_b0 );
buf ( \1912_b1 , \1911_b1 );
not ( \1912_b1 , w_6014 );
not ( \1912_b0 , w_6015 );
and ( w_6014 , w_6015 , \1911_b0 );
or ( \1913_b1 , \1836_b1 , \1839_b1 );
xor ( \1913_b0 , \1836_b0 , w_6016 );
not ( w_6016 , w_6017 );
and ( w_6017 , \1839_b1 , \1839_b0 );
or ( \1914_b1 , \1913_b1 , \1893_b1 );
xor ( \1914_b0 , \1913_b0 , w_6018 );
not ( w_6018 , w_6019 );
and ( w_6019 , \1893_b1 , \1893_b0 );
or ( \1915_b1 , \1912_b1 , w_6021 );
not ( w_6021 , w_6022 );
and ( \1915_b0 , \1912_b0 , w_6023 );
and ( w_6022 ,  , w_6023 );
buf ( w_6021 , \1914_b1 );
not ( w_6021 , w_6024 );
not (  , w_6025 );
and ( w_6024 , w_6025 , \1914_b0 );
or ( \1916_b1 , \1774_b1 , \1780_b1 );
xor ( \1916_b0 , \1774_b0 , w_6026 );
not ( w_6026 , w_6027 );
and ( w_6027 , \1780_b1 , \1780_b0 );
or ( \1917_b1 , \1916_b1 , \1787_b1 );
xor ( \1917_b0 , \1916_b0 , w_6028 );
not ( w_6028 , w_6029 );
and ( w_6029 , \1787_b1 , \1787_b0 );
buf ( \1918_b1 , \1917_b1 );
not ( \1918_b1 , w_6030 );
not ( \1918_b0 , w_6031 );
and ( w_6030 , w_6031 , \1917_b0 );
or ( \1919_b1 , \1798_b1 , \1804_b1 );
xor ( \1919_b0 , \1798_b0 , w_6032 );
not ( w_6032 , w_6033 );
and ( w_6033 , \1804_b1 , \1804_b0 );
or ( \1920_b1 , \1919_b1 , \1811_b1 );
xor ( \1920_b0 , \1919_b0 , w_6034 );
not ( w_6034 , w_6035 );
and ( w_6035 , \1811_b1 , \1811_b0 );
buf ( \1921_b1 , \1920_b1 );
not ( \1921_b1 , w_6036 );
not ( \1921_b0 , w_6037 );
and ( w_6036 , w_6037 , \1920_b0 );
or ( \1922_b1 , \1918_b1 , w_6039 );
not ( w_6039 , w_6040 );
and ( \1922_b0 , \1918_b0 , w_6041 );
and ( w_6040 ,  , w_6041 );
buf ( w_6039 , \1921_b1 );
not ( w_6039 , w_6042 );
not (  , w_6043 );
and ( w_6042 , w_6043 , \1921_b0 );
buf ( \1923_b1 , \1922_b1 );
not ( \1923_b1 , w_6044 );
not ( \1923_b0 , w_6045 );
and ( w_6044 , w_6045 , \1922_b0 );
or ( \1924_b1 , \a[0]_b1 , \d[11]_b1 );
xor ( \1924_b0 , \a[0]_b0 , w_6046 );
not ( w_6046 , w_6047 );
and ( w_6047 , \d[11]_b1 , \d[11]_b0 );
buf ( \1925_b1 , \1924_b1 );
not ( \1925_b1 , w_6048 );
not ( \1925_b0 , w_6049 );
and ( w_6048 , w_6049 , \1924_b0 );
buf ( \1926_b1 , \1638_b1 );
not ( \1926_b1 , w_6050 );
not ( \1926_b0 , w_6051 );
and ( w_6050 , w_6051 , \1638_b0 );
or ( \1927_b1 , \1925_b1 , w_6052 );
or ( \1927_b0 , \1925_b0 , \1926_b0 );
not ( \1926_b0 , w_6053 );
and ( w_6053 , w_6052 , \1926_b1 );
or ( \1928_b1 , \1641_b1 , w_6055 );
not ( w_6055 , w_6056 );
and ( \1928_b0 , \1641_b0 , w_6057 );
and ( w_6056 ,  , w_6057 );
buf ( w_6055 , \1806_b1 );
not ( w_6055 , w_6058 );
not (  , w_6059 );
and ( w_6058 , w_6059 , \1806_b0 );
or ( \1929_b1 , \1927_b1 , w_6061 );
not ( w_6061 , w_6062 );
and ( \1929_b0 , \1927_b0 , w_6063 );
and ( w_6062 ,  , w_6063 );
buf ( w_6061 , \1928_b1 );
not ( w_6061 , w_6064 );
not (  , w_6065 );
and ( w_6064 , w_6065 , \1928_b0 );
buf ( \1930_b1 , \1929_b1 );
not ( \1930_b1 , w_6066 );
not ( \1930_b0 , w_6067 );
and ( w_6066 , w_6067 , \1929_b0 );
or ( \1931_b1 , \a[6]_b1 , \d[5]_b1 );
xor ( \1931_b0 , \a[6]_b0 , w_6068 );
not ( w_6068 , w_6069 );
and ( w_6069 , \d[5]_b1 , \d[5]_b0 );
buf ( \1932_b1 , \1931_b1 );
not ( \1932_b1 , w_6070 );
not ( \1932_b0 , w_6071 );
and ( w_6070 , w_6071 , \1931_b0 );
buf ( \1933_b1 , \1135_b1 );
not ( \1933_b1 , w_6072 );
not ( \1933_b0 , w_6073 );
and ( w_6072 , w_6073 , \1135_b0 );
or ( \1934_b1 , \1932_b1 , w_6074 );
or ( \1934_b0 , \1932_b0 , \1933_b0 );
not ( \1933_b0 , w_6075 );
and ( w_6075 , w_6074 , \1933_b1 );
or ( \1935_b1 , \951_b1 , w_6077 );
not ( w_6077 , w_6078 );
and ( \1935_b0 , \951_b0 , w_6079 );
and ( w_6078 ,  , w_6079 );
buf ( w_6077 , \1842_b1 );
not ( w_6077 , w_6080 );
not (  , w_6081 );
and ( w_6080 , w_6081 , \1842_b0 );
or ( \1936_b1 , \1934_b1 , w_6083 );
not ( w_6083 , w_6084 );
and ( \1936_b0 , \1934_b0 , w_6085 );
and ( w_6084 ,  , w_6085 );
buf ( w_6083 , \1935_b1 );
not ( w_6083 , w_6086 );
not (  , w_6087 );
and ( w_6086 , w_6087 , \1935_b0 );
buf ( \1937_b1 , \1936_b1 );
not ( \1937_b1 , w_6088 );
not ( \1937_b0 , w_6089 );
and ( w_6088 , w_6089 , \1936_b0 );
or ( \1938_b1 , \1930_b1 , w_6090 );
or ( \1938_b0 , \1930_b0 , \1937_b0 );
not ( \1937_b0 , w_6091 );
and ( w_6091 , w_6090 , \1937_b1 );
or ( \1939_b1 , \1936_b1 , w_6092 );
or ( \1939_b0 , \1936_b0 , \1929_b0 );
not ( \1929_b0 , w_6093 );
and ( w_6093 , w_6092 , \1929_b1 );
or ( \1940_b1 , \1855_b1 , \1860_b1 );
not ( \1860_b1 , w_6094 );
and ( \1940_b0 , \1855_b0 , w_6095 );
and ( w_6094 , w_6095 , \1860_b0 );
buf ( \1941_b1 , \1855_b1 );
not ( \1941_b1 , w_6096 );
not ( \1941_b0 , w_6097 );
and ( w_6096 , w_6097 , \1855_b0 );
or ( \1942_b1 , \1941_b1 , \1859_b1 );
not ( \1859_b1 , w_6098 );
and ( \1942_b0 , \1941_b0 , w_6099 );
and ( w_6098 , w_6099 , \1859_b0 );
or ( \1943_b1 , \1940_b1 , w_6101 );
not ( w_6101 , w_6102 );
and ( \1943_b0 , \1940_b0 , w_6103 );
and ( w_6102 ,  , w_6103 );
buf ( w_6101 , \1942_b1 );
not ( w_6101 , w_6104 );
not (  , w_6105 );
and ( w_6104 , w_6105 , \1942_b0 );
or ( \1944_b1 , \1939_b1 , w_6107 );
not ( w_6107 , w_6108 );
and ( \1944_b0 , \1939_b0 , w_6109 );
and ( w_6108 ,  , w_6109 );
buf ( w_6107 , \1943_b1 );
not ( w_6107 , w_6110 );
not (  , w_6111 );
and ( w_6110 , w_6111 , \1943_b0 );
or ( \1945_b1 , \1938_b1 , w_6113 );
not ( w_6113 , w_6114 );
and ( \1945_b0 , \1938_b0 , w_6115 );
and ( w_6114 ,  , w_6115 );
buf ( w_6113 , \1944_b1 );
not ( w_6113 , w_6116 );
not (  , w_6117 );
and ( w_6116 , w_6117 , \1944_b0 );
buf ( \1946_b1 , \1945_b1 );
not ( \1946_b1 , w_6118 );
not ( \1946_b0 , w_6119 );
and ( w_6118 , w_6119 , \1945_b0 );
or ( \1947_b1 , \1923_b1 , w_6120 );
or ( \1947_b0 , \1923_b0 , \1946_b0 );
not ( \1946_b0 , w_6121 );
and ( w_6121 , w_6120 , \1946_b1 );
buf ( \1948_b1 , \1921_b1 );
not ( \1948_b1 , w_6122 );
not ( \1948_b0 , w_6123 );
and ( w_6122 , w_6123 , \1921_b0 );
or ( \1949_b1 , \1948_b1 , w_6125 );
not ( w_6125 , w_6126 );
and ( \1949_b0 , \1948_b0 , w_6127 );
and ( w_6126 ,  , w_6127 );
buf ( w_6125 , \1917_b1 );
not ( w_6125 , w_6128 );
not (  , w_6129 );
and ( w_6128 , w_6129 , \1917_b0 );
or ( \1950_b1 , \1947_b1 , w_6131 );
not ( w_6131 , w_6132 );
and ( \1950_b0 , \1947_b0 , w_6133 );
and ( w_6132 ,  , w_6133 );
buf ( w_6131 , \1949_b1 );
not ( w_6131 , w_6134 );
not (  , w_6135 );
and ( w_6134 , w_6135 , \1949_b0 );
or ( \1951_b1 , \1915_b1 , \1950_b1 );
not ( \1950_b1 , w_6136 );
and ( \1951_b0 , \1915_b0 , w_6137 );
and ( w_6136 , w_6137 , \1950_b0 );
or ( \1952_b1 , \1914_b1 , w_6139 );
not ( w_6139 , w_6140 );
and ( \1952_b0 , \1914_b0 , w_6141 );
and ( w_6140 ,  , w_6141 );
buf ( w_6139 , \1910_b1 );
not ( w_6139 , w_6142 );
not (  , w_6143 );
and ( w_6142 , w_6143 , \1910_b0 );
or ( \1953_b1 , \1951_b1 , w_6145 );
not ( w_6145 , w_6146 );
and ( \1953_b0 , \1951_b0 , w_6147 );
and ( w_6146 ,  , w_6147 );
buf ( w_6145 , \1952_b1 );
not ( w_6145 , w_6148 );
not (  , w_6149 );
and ( w_6148 , w_6149 , \1952_b0 );
or ( \1954_b1 , \1908_b1 , w_6151 );
not ( w_6151 , w_6152 );
and ( \1954_b0 , \1908_b0 , w_6153 );
and ( w_6152 ,  , w_6153 );
buf ( w_6151 , \1953_b1 );
not ( w_6151 , w_6154 );
not (  , w_6155 );
and ( w_6154 , w_6155 , \1953_b0 );
buf ( \1955_b1 , \1954_b1 );
not ( \1955_b1 , w_6156 );
not ( \1955_b0 , w_6157 );
and ( w_6156 , w_6157 , \1954_b0 );
buf ( \1956_b1 , \1911_b1 );
not ( \1956_b1 , w_6158 );
not ( \1956_b0 , w_6159 );
and ( w_6158 , w_6159 , \1911_b0 );
buf ( \1957_b1 , \1950_b1 );
not ( \1957_b1 , w_6160 );
not ( \1957_b0 , w_6161 );
and ( w_6160 , w_6161 , \1950_b0 );
buf ( \1958_b1 , \1957_b1 );
not ( \1958_b1 , w_6162 );
not ( \1958_b0 , w_6163 );
and ( w_6162 , w_6163 , \1957_b0 );
or ( \1959_b1 , \1956_b1 , w_6164 );
or ( \1959_b0 , \1956_b0 , \1958_b0 );
not ( \1958_b0 , w_6165 );
and ( w_6165 , w_6164 , \1958_b1 );
or ( \1960_b1 , \1950_b1 , w_6167 );
not ( w_6167 , w_6168 );
and ( \1960_b0 , \1950_b0 , w_6169 );
and ( w_6168 ,  , w_6169 );
buf ( w_6167 , \1910_b1 );
not ( w_6167 , w_6170 );
not (  , w_6171 );
and ( w_6170 , w_6171 , \1910_b0 );
or ( \1961_b1 , \1959_b1 , w_6173 );
not ( w_6173 , w_6174 );
and ( \1961_b0 , \1959_b0 , w_6175 );
and ( w_6174 ,  , w_6175 );
buf ( w_6173 , \1960_b1 );
not ( w_6173 , w_6176 );
not (  , w_6177 );
and ( w_6176 , w_6177 , \1960_b0 );
or ( \1962_b1 , \1914_b1 , \1961_b1 );
xor ( \1962_b0 , \1914_b0 , w_6178 );
not ( w_6178 , w_6179 );
and ( w_6179 , \1961_b1 , \1961_b0 );
or ( \1963_b1 , \1848_b1 , \1861_b1 );
xor ( \1963_b0 , \1848_b0 , w_6180 );
not ( w_6180 , w_6181 );
and ( w_6181 , \1861_b1 , \1861_b0 );
or ( \1964_b1 , \1963_b1 , w_6182 );
xor ( \1964_b0 , \1963_b0 , w_6184 );
not ( w_6184 , w_6185 );
and ( w_6185 , w_6182 , w_6183 );
buf ( w_6182 , \1889_b1 );
not ( w_6182 , w_6186 );
not ( w_6183 , w_6187 );
and ( w_6186 , w_6187 , \1889_b0 );
or ( \1965_b1 , \a[9]_b1 , \d[1]_b1 );
xor ( \1965_b0 , \a[9]_b0 , w_6188 );
not ( w_6188 , w_6189 );
and ( w_6189 , \d[1]_b1 , \d[1]_b0 );
buf ( \1966_b1 , \1965_b1 );
not ( \1966_b1 , w_6190 );
not ( \1966_b0 , w_6191 );
and ( w_6190 , w_6191 , \1965_b0 );
buf ( \1967_b1 , \932_b1 );
not ( \1967_b1 , w_6192 );
not ( \1967_b0 , w_6193 );
and ( w_6192 , w_6193 , \932_b0 );
or ( \1968_b1 , \1966_b1 , w_6194 );
or ( \1968_b0 , \1966_b0 , \1967_b0 );
not ( \1967_b0 , w_6195 );
and ( w_6195 , w_6194 , \1967_b1 );
or ( \1969_b1 , \1864_b1 , w_6197 );
not ( w_6197 , w_6198 );
and ( \1969_b0 , \1864_b0 , w_6199 );
and ( w_6198 ,  , w_6199 );
buf ( w_6197 , \d[0]_b1 );
not ( w_6197 , w_6200 );
not (  , w_6201 );
and ( w_6200 , w_6201 , \d[0]_b0 );
or ( \1970_b1 , \1968_b1 , w_6203 );
not ( w_6203 , w_6204 );
and ( \1970_b0 , \1968_b0 , w_6205 );
and ( w_6204 ,  , w_6205 );
buf ( w_6203 , \1969_b1 );
not ( w_6203 , w_6206 );
not (  , w_6207 );
and ( w_6206 , w_6207 , \1969_b0 );
or ( \1971_b1 , \a[1]_b1 , \d[9]_b1 );
xor ( \1971_b0 , \a[1]_b0 , w_6208 );
not ( w_6208 , w_6209 );
and ( w_6209 , \d[9]_b1 , \d[9]_b0 );
buf ( \1972_b1 , \1971_b1 );
not ( \1972_b1 , w_6210 );
not ( \1972_b0 , w_6211 );
and ( w_6210 , w_6211 , \1971_b0 );
buf ( \1973_b1 , \1542_b1 );
not ( \1973_b1 , w_6212 );
not ( \1973_b0 , w_6213 );
and ( w_6212 , w_6213 , \1542_b0 );
or ( \1974_b1 , \1972_b1 , w_6214 );
or ( \1974_b0 , \1972_b0 , \1973_b0 );
not ( \1973_b0 , w_6215 );
and ( w_6215 , w_6214 , \1973_b1 );
or ( \1975_b1 , \1541_b1 , w_6217 );
not ( w_6217 , w_6218 );
and ( \1975_b0 , \1541_b0 , w_6219 );
and ( w_6218 ,  , w_6219 );
buf ( w_6217 , \1871_b1 );
not ( w_6217 , w_6220 );
not (  , w_6221 );
and ( w_6220 , w_6221 , \1871_b0 );
or ( \1976_b1 , \1974_b1 , w_6223 );
not ( w_6223 , w_6224 );
and ( \1976_b0 , \1974_b0 , w_6225 );
and ( w_6224 ,  , w_6225 );
buf ( w_6223 , \1975_b1 );
not ( w_6223 , w_6226 );
not (  , w_6227 );
and ( w_6226 , w_6227 , \1975_b0 );
or ( \1977_b1 , \1970_b1 , w_6228 );
or ( \1977_b0 , \1970_b0 , \1976_b0 );
not ( \1976_b0 , w_6229 );
and ( w_6229 , w_6228 , \1976_b1 );
or ( \1978_b1 , \a[5]_b1 , \d[5]_b1 );
xor ( \1978_b0 , \a[5]_b0 , w_6230 );
not ( w_6230 , w_6231 );
and ( w_6231 , \d[5]_b1 , \d[5]_b0 );
buf ( \1979_b1 , \1978_b1 );
not ( \1979_b1 , w_6232 );
not ( \1979_b0 , w_6233 );
and ( w_6232 , w_6233 , \1978_b0 );
buf ( \1980_b1 , \948_b1 );
not ( \1980_b1 , w_6234 );
not ( \1980_b0 , w_6235 );
and ( w_6234 , w_6235 , \948_b0 );
or ( \1981_b1 , \1979_b1 , w_6236 );
or ( \1981_b0 , \1979_b0 , \1980_b0 );
not ( \1980_b0 , w_6237 );
and ( w_6237 , w_6236 , \1980_b1 );
or ( \1982_b1 , \951_b1 , w_6239 );
not ( w_6239 , w_6240 );
and ( \1982_b0 , \951_b0 , w_6241 );
and ( w_6240 ,  , w_6241 );
buf ( w_6239 , \1931_b1 );
not ( w_6239 , w_6242 );
not (  , w_6243 );
and ( w_6242 , w_6243 , \1931_b0 );
or ( \1983_b1 , \1981_b1 , w_6245 );
not ( w_6245 , w_6246 );
and ( \1983_b0 , \1981_b0 , w_6247 );
and ( w_6246 ,  , w_6247 );
buf ( w_6245 , \1982_b1 );
not ( w_6245 , w_6248 );
not (  , w_6249 );
and ( w_6248 , w_6249 , \1982_b0 );
or ( \1984_b1 , \1977_b1 , w_6251 );
not ( w_6251 , w_6252 );
and ( \1984_b0 , \1977_b0 , w_6253 );
and ( w_6252 ,  , w_6253 );
buf ( w_6251 , \1983_b1 );
not ( w_6251 , w_6254 );
not (  , w_6255 );
and ( w_6254 , w_6255 , \1983_b0 );
or ( \1985_b1 , \1976_b1 , w_6257 );
not ( w_6257 , w_6258 );
and ( \1985_b0 , \1976_b0 , w_6259 );
and ( w_6258 ,  , w_6259 );
buf ( w_6257 , \1970_b1 );
not ( w_6257 , w_6260 );
not (  , w_6261 );
and ( w_6260 , w_6261 , \1970_b0 );
or ( \1986_b1 , \1984_b1 , w_6263 );
not ( w_6263 , w_6264 );
and ( \1986_b0 , \1984_b0 , w_6265 );
and ( w_6264 ,  , w_6265 );
buf ( w_6263 , \1985_b1 );
not ( w_6263 , w_6266 );
not (  , w_6267 );
and ( w_6266 , w_6267 , \1985_b0 );
buf ( \1987_b1 , \1986_b1 );
not ( \1987_b1 , w_6268 );
not ( \1987_b0 , w_6269 );
and ( w_6268 , w_6269 , \1986_b0 );
buf ( \1988_b1 , \1987_b1 );
not ( \1988_b1 , w_6270 );
not ( \1988_b0 , w_6271 );
and ( w_6270 , w_6271 , \1987_b0 );
buf ( \1989_b1 , \1887_b1 );
not ( \1989_b1 , w_6272 );
not ( \1989_b0 , w_6273 );
and ( w_6272 , w_6273 , \1887_b0 );
buf ( \1990_b1 , \1869_b1 );
not ( \1990_b1 , w_6274 );
not ( \1990_b0 , w_6275 );
and ( w_6274 , w_6275 , \1869_b0 );
buf ( \1991_b1 , \1990_b1 );
not ( \1991_b1 , w_6276 );
not ( \1991_b0 , w_6277 );
and ( w_6276 , w_6277 , \1990_b0 );
or ( \1992_b1 , \1989_b1 , w_6278 );
or ( \1992_b0 , \1989_b0 , \1991_b0 );
not ( \1991_b0 , w_6279 );
and ( w_6279 , w_6278 , \1991_b1 );
buf ( \1993_b1 , \1887_b1 );
not ( \1993_b1 , w_6280 );
not ( \1993_b0 , w_6281 );
and ( w_6280 , w_6281 , \1887_b0 );
or ( \1994_b1 , \1993_b1 , w_6283 );
not ( w_6283 , w_6284 );
and ( \1994_b0 , \1993_b0 , w_6285 );
and ( w_6284 ,  , w_6285 );
buf ( w_6283 , \1869_b1 );
not ( w_6283 , w_6286 );
not (  , w_6287 );
and ( w_6286 , w_6287 , \1869_b0 );
or ( \1995_b1 , \1992_b1 , w_6289 );
not ( w_6289 , w_6290 );
and ( \1995_b0 , \1992_b0 , w_6291 );
and ( w_6290 ,  , w_6291 );
buf ( w_6289 , \1994_b1 );
not ( w_6289 , w_6292 );
not (  , w_6293 );
and ( w_6292 , w_6293 , \1994_b0 );
buf ( \1996_b1 , \1876_b1 );
not ( \1996_b1 , w_6294 );
not ( \1996_b0 , w_6295 );
and ( w_6294 , w_6295 , \1876_b0 );
or ( \1997_b1 , \1995_b1 , \1996_b1 );
not ( \1996_b1 , w_6296 );
and ( \1997_b0 , \1995_b0 , w_6297 );
and ( w_6296 , w_6297 , \1996_b0 );
buf ( \1998_b1 , \1995_b1 );
not ( \1998_b1 , w_6298 );
not ( \1998_b0 , w_6299 );
and ( w_6298 , w_6299 , \1995_b0 );
or ( \1999_b1 , \1998_b1 , \1876_b1 );
not ( \1876_b1 , w_6300 );
and ( \1999_b0 , \1998_b0 , w_6301 );
and ( w_6300 , w_6301 , \1876_b0 );
or ( \2000_b1 , \1997_b1 , w_6303 );
not ( w_6303 , w_6304 );
and ( \2000_b0 , \1997_b0 , w_6305 );
and ( w_6304 ,  , w_6305 );
buf ( w_6303 , \1999_b1 );
not ( w_6303 , w_6306 );
not (  , w_6307 );
and ( w_6306 , w_6307 , \1999_b0 );
buf ( \2001_b1 , \2000_b1 );
not ( \2001_b1 , w_6308 );
not ( \2001_b0 , w_6309 );
and ( w_6308 , w_6309 , \2000_b0 );
or ( \2002_b1 , \1988_b1 , w_6310 );
or ( \2002_b0 , \1988_b0 , \2001_b0 );
not ( \2001_b0 , w_6311 );
and ( w_6311 , w_6310 , \2001_b1 );
or ( \2003_b1 , \d[3]_b1 , \a[7]_b1 );
xor ( \2003_b0 , \d[3]_b0 , w_6312 );
not ( w_6312 , w_6313 );
and ( w_6313 , \a[7]_b1 , \a[7]_b0 );
buf ( \2004_b1 , \2003_b1 );
not ( \2004_b1 , w_6314 );
not ( \2004_b0 , w_6315 );
and ( w_6314 , w_6315 , \2003_b0 );
buf ( \2005_b1 , \973_b1 );
not ( \2005_b1 , w_6316 );
not ( \2005_b0 , w_6317 );
and ( w_6316 , w_6317 , \973_b0 );
or ( \2006_b1 , \2004_b1 , w_6318 );
or ( \2006_b0 , \2004_b0 , \2005_b0 );
not ( \2005_b0 , w_6319 );
and ( w_6319 , w_6318 , \2005_b1 );
or ( \2007_b1 , \976_b1 , w_6321 );
not ( w_6321 , w_6322 );
and ( \2007_b0 , \976_b0 , w_6323 );
and ( w_6322 ,  , w_6323 );
buf ( w_6321 , \1850_b1 );
not ( w_6321 , w_6324 );
not (  , w_6325 );
and ( w_6324 , w_6325 , \1850_b0 );
or ( \2008_b1 , \2006_b1 , w_6327 );
not ( w_6327 , w_6328 );
and ( \2008_b0 , \2006_b0 , w_6329 );
and ( w_6328 ,  , w_6329 );
buf ( w_6327 , \2007_b1 );
not ( w_6327 , w_6330 );
not (  , w_6331 );
and ( w_6330 , w_6331 , \2007_b0 );
or ( \2009_b1 , \1641_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_6332 );
and ( \2009_b0 , \1641_b0 , w_6333 );
and ( w_6332 , w_6333 , \a[0]_b0 );
or ( \2010_b1 , \2008_b1 , w_6334 );
or ( \2010_b0 , \2008_b0 , \2009_b0 );
not ( \2009_b0 , w_6335 );
and ( w_6335 , w_6334 , \2009_b1 );
or ( \2011_b1 , \a[3]_b1 , \d[7]_b1 );
xor ( \2011_b0 , \a[3]_b0 , w_6336 );
not ( w_6336 , w_6337 );
and ( w_6337 , \d[7]_b1 , \d[7]_b0 );
buf ( \2012_b1 , \2011_b1 );
not ( \2012_b1 , w_6338 );
not ( \2012_b0 , w_6339 );
and ( w_6338 , w_6339 , \2011_b0 );
buf ( \2013_b1 , \1127_b1 );
not ( \2013_b1 , w_6340 );
not ( \2013_b0 , w_6341 );
and ( w_6340 , w_6341 , \1127_b0 );
or ( \2014_b1 , \2012_b1 , w_6342 );
or ( \2014_b0 , \2012_b0 , \2013_b0 );
not ( \2013_b0 , w_6343 );
and ( w_6343 , w_6342 , \2013_b1 );
or ( \2015_b1 , \958_b1 , w_6345 );
not ( w_6345 , w_6346 );
and ( \2015_b0 , \958_b0 , w_6347 );
and ( w_6346 ,  , w_6347 );
buf ( w_6345 , \1880_b1 );
not ( w_6345 , w_6348 );
not (  , w_6349 );
and ( w_6348 , w_6349 , \1880_b0 );
or ( \2016_b1 , \2014_b1 , w_6351 );
not ( w_6351 , w_6352 );
and ( \2016_b0 , \2014_b0 , w_6353 );
and ( w_6352 ,  , w_6353 );
buf ( w_6351 , \2015_b1 );
not ( w_6351 , w_6354 );
not (  , w_6355 );
and ( w_6354 , w_6355 , \2015_b0 );
or ( \2017_b1 , \2010_b1 , \2016_b1 );
not ( \2016_b1 , w_6356 );
and ( \2017_b0 , \2010_b0 , w_6357 );
and ( w_6356 , w_6357 , \2016_b0 );
or ( \2018_b1 , \2008_b1 , \2009_b1 );
not ( \2009_b1 , w_6358 );
and ( \2018_b0 , \2008_b0 , w_6359 );
and ( w_6358 , w_6359 , \2009_b0 );
or ( \2019_b1 , \2017_b1 , w_6361 );
not ( w_6361 , w_6362 );
and ( \2019_b0 , \2017_b0 , w_6363 );
and ( w_6362 ,  , w_6363 );
buf ( w_6361 , \2018_b1 );
not ( w_6361 , w_6364 );
not (  , w_6365 );
and ( w_6364 , w_6365 , \2018_b0 );
buf ( \2020_b1 , \2019_b1 );
not ( \2020_b1 , w_6366 );
not ( \2020_b0 , w_6367 );
and ( w_6366 , w_6367 , \2019_b0 );
or ( \2021_b1 , \2002_b1 , w_6369 );
not ( w_6369 , w_6370 );
and ( \2021_b0 , \2002_b0 , w_6371 );
and ( w_6370 ,  , w_6371 );
buf ( w_6369 , \2020_b1 );
not ( w_6369 , w_6372 );
not (  , w_6373 );
and ( w_6372 , w_6373 , \2020_b0 );
buf ( \2022_b1 , \2000_b1 );
not ( \2022_b1 , w_6374 );
not ( \2022_b0 , w_6375 );
and ( w_6374 , w_6375 , \2000_b0 );
or ( \2023_b1 , \2022_b1 , w_6377 );
not ( w_6377 , w_6378 );
and ( \2023_b0 , \2022_b0 , w_6379 );
and ( w_6378 ,  , w_6379 );
buf ( w_6377 , \1986_b1 );
not ( w_6377 , w_6380 );
not (  , w_6381 );
and ( w_6380 , w_6381 , \1986_b0 );
or ( \2024_b1 , \2021_b1 , \2023_b1 );
not ( \2023_b1 , w_6382 );
and ( \2024_b0 , \2021_b0 , w_6383 );
and ( w_6382 , w_6383 , \2023_b0 );
or ( \2025_b1 , \1964_b1 , \2024_b1 );
xor ( \2025_b0 , \1964_b0 , w_6384 );
not ( w_6384 , w_6385 );
and ( w_6385 , \2024_b1 , \2024_b0 );
or ( \2026_b1 , \1917_b1 , \1920_b1 );
xor ( \2026_b0 , \1917_b0 , w_6386 );
not ( w_6386 , w_6387 );
and ( w_6387 , \1920_b1 , \1920_b0 );
or ( \2027_b1 , \2026_b1 , w_6388 );
xor ( \2027_b0 , \2026_b0 , w_6390 );
not ( w_6390 , w_6391 );
and ( w_6391 , w_6388 , w_6389 );
buf ( w_6388 , \1945_b1 );
not ( w_6388 , w_6392 );
not ( w_6389 , w_6393 );
and ( w_6392 , w_6393 , \1945_b0 );
or ( \2028_b1 , \2025_b1 , \2027_b1 );
not ( \2027_b1 , w_6394 );
and ( \2028_b0 , \2025_b0 , w_6395 );
and ( w_6394 , w_6395 , \2027_b0 );
or ( \2029_b1 , \1964_b1 , \2024_b1 );
not ( \2024_b1 , w_6396 );
and ( \2029_b0 , \1964_b0 , w_6397 );
and ( w_6396 , w_6397 , \2024_b0 );
or ( \2030_b1 , \2028_b1 , w_6398 );
or ( \2030_b0 , \2028_b0 , \2029_b0 );
not ( \2029_b0 , w_6399 );
and ( w_6399 , w_6398 , \2029_b1 );
or ( \2031_b1 , \1962_b1 , w_6401 );
not ( w_6401 , w_6402 );
and ( \2031_b0 , \1962_b0 , w_6403 );
and ( w_6402 ,  , w_6403 );
buf ( w_6401 , \2030_b1 );
not ( w_6401 , w_6404 );
not (  , w_6405 );
and ( w_6404 , w_6405 , \2030_b0 );
or ( \2032_b1 , \a[0]_b1 , w_6406 );
or ( \2032_b0 , \a[0]_b0 , \d[8]_b0 );
not ( \d[8]_b0 , w_6407 );
and ( w_6407 , w_6406 , \d[8]_b1 );
or ( \2033_b1 , \2032_b1 , w_6409 );
not ( w_6409 , w_6410 );
and ( \2033_b0 , \2032_b0 , w_6411 );
and ( w_6410 ,  , w_6411 );
buf ( w_6409 , \d[7]_b1 );
not ( w_6409 , w_6412 );
not (  , w_6413 );
and ( w_6412 , w_6413 , \d[7]_b0 );
or ( \2034_b1 , \a[0]_b1 , w_6415 );
not ( w_6415 , w_6416 );
and ( \2034_b0 , \a[0]_b0 , w_6417 );
and ( w_6416 ,  , w_6417 );
buf ( w_6415 , \d[8]_b1 );
not ( w_6415 , w_6418 );
not (  , w_6419 );
and ( w_6418 , w_6419 , \d[8]_b0 );
or ( \2036_b1 , \a[6]_b1 , \d[3]_b1 );
xor ( \2036_b0 , \a[6]_b0 , w_6420 );
not ( w_6420 , w_6421 );
and ( w_6421 , \d[3]_b1 , \d[3]_b0 );
buf ( \2037_b1 , \2036_b1 );
not ( \2037_b1 , w_6422 );
not ( \2037_b0 , w_6423 );
and ( w_6422 , w_6423 , \2036_b0 );
buf ( \2038_b1 , \973_b1 );
not ( \2038_b1 , w_6424 );
not ( \2038_b0 , w_6425 );
and ( w_6424 , w_6425 , \973_b0 );
or ( \2039_b1 , \2037_b1 , w_6426 );
or ( \2039_b0 , \2037_b0 , \2038_b0 );
not ( \2038_b0 , w_6427 );
and ( w_6427 , w_6426 , \2038_b1 );
or ( \2040_b1 , \976_b1 , w_6429 );
not ( w_6429 , w_6430 );
and ( \2040_b0 , \976_b0 , w_6431 );
and ( w_6430 ,  , w_6431 );
buf ( w_6429 , \2003_b1 );
not ( w_6429 , w_6432 );
not (  , w_6433 );
and ( w_6432 , w_6433 , \2003_b0 );
or ( \2041_b1 , \2039_b1 , w_6435 );
not ( w_6435 , w_6436 );
and ( \2041_b0 , \2039_b0 , w_6437 );
and ( w_6436 ,  , w_6437 );
buf ( w_6435 , \2040_b1 );
not ( w_6435 , w_6438 );
not (  , w_6439 );
and ( w_6438 , w_6439 , \2040_b0 );
or ( \2042_b1 , \2035_b1 , \2041_b1 );
not ( \2041_b1 , w_6440 );
and ( \2042_b0 , \2035_b0 , w_6441 );
and ( w_6440 , w_6441 , \2041_b0 );
or ( \2043_b1 , \a[8]_b1 , \d[1]_b1 );
xor ( \2043_b0 , \a[8]_b0 , w_6442 );
not ( w_6442 , w_6443 );
and ( w_6443 , \d[1]_b1 , \d[1]_b0 );
buf ( \2044_b1 , \2043_b1 );
not ( \2044_b1 , w_6444 );
not ( \2044_b0 , w_6445 );
and ( w_6444 , w_6445 , \2043_b0 );
buf ( \2045_b1 , \932_b1 );
not ( \2045_b1 , w_6446 );
not ( \2045_b0 , w_6447 );
and ( w_6446 , w_6447 , \932_b0 );
or ( \2046_b1 , \2044_b1 , w_6448 );
or ( \2046_b0 , \2044_b0 , \2045_b0 );
not ( \2045_b0 , w_6449 );
and ( w_6449 , w_6448 , \2045_b1 );
or ( \2047_b1 , \1965_b1 , w_6451 );
not ( w_6451 , w_6452 );
and ( \2047_b0 , \1965_b0 , w_6453 );
and ( w_6452 ,  , w_6453 );
buf ( w_6451 , \d[0]_b1 );
not ( w_6451 , w_6454 );
not (  , w_6455 );
and ( w_6454 , w_6455 , \d[0]_b0 );
or ( \2048_b1 , \2046_b1 , w_6457 );
not ( w_6457 , w_6458 );
and ( \2048_b0 , \2046_b0 , w_6459 );
and ( w_6458 ,  , w_6459 );
buf ( w_6457 , \2047_b1 );
not ( w_6457 , w_6460 );
not (  , w_6461 );
and ( w_6460 , w_6461 , \2047_b0 );
or ( \2049_b1 , \a[0]_b1 , \d[9]_b1 );
xor ( \2049_b0 , \a[0]_b0 , w_6462 );
not ( w_6462 , w_6463 );
and ( w_6463 , \d[9]_b1 , \d[9]_b0 );
buf ( \2050_b1 , \2049_b1 );
not ( \2050_b1 , w_6464 );
not ( \2050_b0 , w_6465 );
and ( w_6464 , w_6465 , \2049_b0 );
buf ( \2051_b1 , \1542_b1 );
not ( \2051_b1 , w_6466 );
not ( \2051_b0 , w_6467 );
and ( w_6466 , w_6467 , \1542_b0 );
or ( \2052_b1 , \2050_b1 , w_6468 );
or ( \2052_b0 , \2050_b0 , \2051_b0 );
not ( \2051_b0 , w_6469 );
and ( w_6469 , w_6468 , \2051_b1 );
or ( \2053_b1 , \1545_b1 , w_6471 );
not ( w_6471 , w_6472 );
and ( \2053_b0 , \1545_b0 , w_6473 );
and ( w_6472 ,  , w_6473 );
buf ( w_6471 , \1971_b1 );
not ( w_6471 , w_6474 );
not (  , w_6475 );
and ( w_6474 , w_6475 , \1971_b0 );
or ( \2054_b1 , \2052_b1 , w_6477 );
not ( w_6477 , w_6478 );
and ( \2054_b0 , \2052_b0 , w_6479 );
and ( w_6478 ,  , w_6479 );
buf ( w_6477 , \2053_b1 );
not ( w_6477 , w_6480 );
not (  , w_6481 );
and ( w_6480 , w_6481 , \2053_b0 );
or ( \2055_b1 , \2048_b1 , w_6482 );
or ( \2055_b0 , \2048_b0 , \2054_b0 );
not ( \2054_b0 , w_6483 );
and ( w_6483 , w_6482 , \2054_b1 );
or ( \2056_b1 , \a[2]_b1 , \d[7]_b1 );
xor ( \2056_b0 , \a[2]_b0 , w_6484 );
not ( w_6484 , w_6485 );
and ( w_6485 , \d[7]_b1 , \d[7]_b0 );
buf ( \2057_b1 , \2056_b1 );
not ( \2057_b1 , w_6486 );
not ( \2057_b0 , w_6487 );
and ( w_6486 , w_6487 , \2056_b0 );
buf ( \2058_b1 , \1883_b1 );
not ( \2058_b1 , w_6488 );
not ( \2058_b0 , w_6489 );
and ( w_6488 , w_6489 , \1883_b0 );
or ( \2059_b1 , \2057_b1 , w_6490 );
or ( \2059_b0 , \2057_b0 , \2058_b0 );
not ( \2058_b0 , w_6491 );
and ( w_6491 , w_6490 , \2058_b1 );
or ( \2060_b1 , \958_b1 , w_6493 );
not ( w_6493 , w_6494 );
and ( \2060_b0 , \958_b0 , w_6495 );
and ( w_6494 ,  , w_6495 );
buf ( w_6493 , \2011_b1 );
not ( w_6493 , w_6496 );
not (  , w_6497 );
and ( w_6496 , w_6497 , \2011_b0 );
or ( \2061_b1 , \2059_b1 , w_6499 );
not ( w_6499 , w_6500 );
and ( \2061_b0 , \2059_b0 , w_6501 );
and ( w_6500 ,  , w_6501 );
buf ( w_6499 , \2060_b1 );
not ( w_6499 , w_6502 );
not (  , w_6503 );
and ( w_6502 , w_6503 , \2060_b0 );
or ( \2062_b1 , \2055_b1 , w_6505 );
not ( w_6505 , w_6506 );
and ( \2062_b0 , \2055_b0 , w_6507 );
and ( w_6506 ,  , w_6507 );
buf ( w_6505 , \2061_b1 );
not ( w_6505 , w_6508 );
not (  , w_6509 );
and ( w_6508 , w_6509 , \2061_b0 );
or ( \2063_b1 , \2048_b1 , w_6511 );
not ( w_6511 , w_6512 );
and ( \2063_b0 , \2048_b0 , w_6513 );
and ( w_6512 ,  , w_6513 );
buf ( w_6511 , \2054_b1 );
not ( w_6511 , w_6514 );
not (  , w_6515 );
and ( w_6514 , w_6515 , \2054_b0 );
or ( \2064_b1 , \2062_b1 , w_6517 );
not ( w_6517 , w_6518 );
and ( \2064_b0 , \2062_b0 , w_6519 );
and ( w_6518 ,  , w_6519 );
buf ( w_6517 , \2063_b1 );
not ( w_6517 , w_6520 );
not (  , w_6521 );
and ( w_6520 , w_6521 , \2063_b0 );
or ( \2065_b1 , \2042_b1 , \2064_b1 );
xor ( \2065_b0 , \2042_b0 , w_6522 );
not ( w_6522 , w_6523 );
and ( w_6523 , \2064_b1 , \2064_b0 );
or ( \2066_b1 , \2009_b1 , \2016_b1 );
xor ( \2066_b0 , \2009_b0 , w_6524 );
not ( w_6524 , w_6525 );
and ( w_6525 , \2016_b1 , \2016_b0 );
or ( \2067_b1 , \2066_b1 , \2008_b1 );
xor ( \2067_b0 , \2066_b0 , w_6526 );
not ( w_6526 , w_6527 );
and ( w_6527 , \2008_b1 , \2008_b0 );
or ( \2068_b1 , \2065_b1 , \2067_b1 );
xor ( \2068_b0 , \2065_b0 , w_6528 );
not ( w_6528 , w_6529 );
and ( w_6529 , \2067_b1 , \2067_b0 );
or ( \2069_b1 , \1976_b1 , \1970_b1 );
xor ( \2069_b0 , \1976_b0 , w_6530 );
not ( w_6530 , w_6531 );
and ( w_6531 , \1970_b1 , \1970_b0 );
or ( \2070_b1 , \2069_b1 , \1983_b1 );
xor ( \2070_b0 , \2069_b0 , w_6532 );
not ( w_6532 , w_6533 );
and ( w_6533 , \1983_b1 , \1983_b0 );
or ( \2071_b1 , \2068_b1 , w_6534 );
or ( \2071_b0 , \2068_b0 , \2070_b0 );
not ( \2070_b0 , w_6535 );
and ( w_6535 , w_6534 , \2070_b1 );
or ( \2072_b1 , \a[4]_b1 , \d[5]_b1 );
xor ( \2072_b0 , \a[4]_b0 , w_6536 );
not ( w_6536 , w_6537 );
and ( w_6537 , \d[5]_b1 , \d[5]_b0 );
buf ( \2073_b1 , \2072_b1 );
not ( \2073_b1 , w_6538 );
not ( \2073_b0 , w_6539 );
and ( w_6538 , w_6539 , \2072_b0 );
buf ( \2074_b1 , \1135_b1 );
not ( \2074_b1 , w_6540 );
not ( \2074_b0 , w_6541 );
and ( w_6540 , w_6541 , \1135_b0 );
or ( \2075_b1 , \2073_b1 , w_6542 );
or ( \2075_b0 , \2073_b0 , \2074_b0 );
not ( \2074_b0 , w_6543 );
and ( w_6543 , w_6542 , \2074_b1 );
or ( \2076_b1 , \951_b1 , w_6545 );
not ( w_6545 , w_6546 );
and ( \2076_b0 , \951_b0 , w_6547 );
and ( w_6546 ,  , w_6547 );
buf ( w_6545 , \1978_b1 );
not ( w_6545 , w_6548 );
not (  , w_6549 );
and ( w_6548 , w_6549 , \1978_b0 );
or ( \2077_b1 , \2075_b1 , w_6551 );
not ( w_6551 , w_6552 );
and ( \2077_b0 , \2075_b0 , w_6553 );
and ( w_6552 ,  , w_6553 );
buf ( w_6551 , \2076_b1 );
not ( w_6551 , w_6554 );
not (  , w_6555 );
and ( w_6554 , w_6555 , \2076_b0 );
or ( \2078_b1 , \1541_b1 , \a[0]_b1 );
not ( \a[0]_b1 , w_6556 );
and ( \2078_b0 , \1541_b0 , w_6557 );
and ( w_6556 , w_6557 , \a[0]_b0 );
buf ( \2079_b1 , \1131_b1 );
not ( \2079_b1 , w_6558 );
not ( \2079_b0 , w_6559 );
and ( w_6558 , w_6559 , \1131_b0 );
buf ( \2080_b1 , \1127_b1 );
not ( \2080_b1 , w_6560 );
not ( \2080_b0 , w_6561 );
and ( w_6560 , w_6561 , \1127_b0 );
or ( \2081_b1 , \2079_b1 , w_6562 );
or ( \2081_b0 , \2079_b0 , \2080_b0 );
not ( \2080_b0 , w_6563 );
and ( w_6563 , w_6562 , \2080_b1 );
or ( \2082_b1 , \958_b1 , w_6565 );
not ( w_6565 , w_6566 );
and ( \2082_b0 , \958_b0 , w_6567 );
and ( w_6566 ,  , w_6567 );
buf ( w_6565 , \2056_b1 );
not ( w_6565 , w_6568 );
not (  , w_6569 );
and ( w_6568 , w_6569 , \2056_b0 );
or ( \2083_b1 , \2081_b1 , w_6571 );
not ( w_6571 , w_6572 );
and ( \2083_b0 , \2081_b0 , w_6573 );
and ( w_6572 ,  , w_6573 );
buf ( w_6571 , \2082_b1 );
not ( w_6571 , w_6574 );
not (  , w_6575 );
and ( w_6574 , w_6575 , \2082_b0 );
or ( \2084_b1 , \2078_b1 , \2083_b1 );
xor ( \2084_b0 , \2078_b0 , w_6576 );
not ( w_6576 , w_6577 );
and ( w_6577 , \2083_b1 , \2083_b0 );
buf ( \2085_b1 , \1106_b1 );
not ( \2085_b1 , w_6578 );
not ( \2085_b0 , w_6579 );
and ( w_6578 , w_6579 , \1106_b0 );
buf ( \2086_b1 , \932_b1 );
not ( \2086_b1 , w_6580 );
not ( \2086_b0 , w_6581 );
and ( w_6580 , w_6581 , \932_b0 );
or ( \2087_b1 , \2085_b1 , w_6582 );
or ( \2087_b0 , \2085_b0 , \2086_b0 );
not ( \2086_b0 , w_6583 );
and ( w_6583 , w_6582 , \2086_b1 );
or ( \2088_b1 , \2043_b1 , w_6585 );
not ( w_6585 , w_6586 );
and ( \2088_b0 , \2043_b0 , w_6587 );
and ( w_6586 ,  , w_6587 );
buf ( w_6585 , \d[0]_b1 );
not ( w_6585 , w_6588 );
not (  , w_6589 );
and ( w_6588 , w_6589 , \d[0]_b0 );
or ( \2089_b1 , \2087_b1 , w_6591 );
not ( w_6591 , w_6592 );
and ( \2089_b0 , \2087_b0 , w_6593 );
and ( w_6592 ,  , w_6593 );
buf ( w_6591 , \2088_b1 );
not ( w_6591 , w_6594 );
not (  , w_6595 );
and ( w_6594 , w_6595 , \2088_b0 );
or ( \2090_b1 , \2084_b1 , \2089_b1 );
not ( \2089_b1 , w_6596 );
and ( \2090_b0 , \2084_b0 , w_6597 );
and ( w_6596 , w_6597 , \2089_b0 );
or ( \2091_b1 , \2078_b1 , \2083_b1 );
not ( \2083_b1 , w_6598 );
and ( \2091_b0 , \2078_b0 , w_6599 );
and ( w_6598 , w_6599 , \2083_b0 );
or ( \2092_b1 , \2090_b1 , w_6600 );
or ( \2092_b0 , \2090_b0 , \2091_b0 );
not ( \2091_b0 , w_6601 );
and ( w_6601 , w_6600 , \2091_b1 );
or ( \2093_b1 , \2077_b1 , \2092_b1 );
xor ( \2093_b0 , \2077_b0 , w_6602 );
not ( w_6602 , w_6603 );
and ( w_6603 , \2092_b1 , \2092_b0 );
or ( \2094_b1 , \2035_b1 , \2041_b1 );
xor ( \2094_b0 , \2035_b0 , w_6604 );
not ( w_6604 , w_6605 );
and ( w_6605 , \2041_b1 , \2041_b0 );
or ( \2095_b1 , \2093_b1 , \2094_b1 );
not ( \2094_b1 , w_6606 );
and ( \2095_b0 , \2093_b0 , w_6607 );
and ( w_6606 , w_6607 , \2094_b0 );
or ( \2096_b1 , \2077_b1 , \2092_b1 );
not ( \2092_b1 , w_6608 );
and ( \2096_b0 , \2077_b0 , w_6609 );
and ( w_6608 , w_6609 , \2092_b0 );
or ( \2097_b1 , \2095_b1 , w_6610 );
or ( \2097_b0 , \2095_b0 , \2096_b0 );
not ( \2096_b0 , w_6611 );
and ( w_6611 , w_6610 , \2096_b1 );
or ( \2098_b1 , \2071_b1 , w_6613 );
not ( w_6613 , w_6614 );
and ( \2098_b0 , \2071_b0 , w_6615 );
and ( w_6614 ,  , w_6615 );
buf ( w_6613 , \2097_b1 );
not ( w_6613 , w_6616 );
not (  , w_6617 );
and ( w_6616 , w_6617 , \2097_b0 );
or ( \2099_b1 , \2068_b1 , w_6619 );
not ( w_6619 , w_6620 );
and ( \2099_b0 , \2068_b0 , w_6621 );
and ( w_6620 ,  , w_6621 );
buf ( w_6619 , \2070_b1 );
not ( w_6619 , w_6622 );
not (  , w_6623 );
and ( w_6622 , w_6623 , \2070_b0 );
or ( \2100_b1 , \2098_b1 , w_6625 );
not ( w_6625 , w_6626 );
and ( \2100_b0 , \2098_b0 , w_6627 );
and ( w_6626 ,  , w_6627 );
buf ( w_6625 , \2099_b1 );
not ( w_6625 , w_6628 );
not (  , w_6629 );
and ( w_6628 , w_6629 , \2099_b0 );
buf ( \2101_b1 , \2100_b1 );
not ( \2101_b1 , w_6630 );
not ( \2101_b0 , w_6631 );
and ( w_6630 , w_6631 , \2100_b0 );
or ( \2102_b1 , \1929_b1 , \1936_b1 );
xor ( \2102_b0 , \1929_b0 , w_6632 );
not ( w_6632 , w_6633 );
and ( w_6633 , \1936_b1 , \1936_b0 );
or ( \2103_b1 , \2102_b1 , \1943_b1 );
xor ( \2103_b0 , \2102_b0 , w_6634 );
not ( w_6634 , w_6635 );
and ( w_6635 , \1943_b1 , \1943_b0 );
or ( \2104_b1 , \1986_b1 , \2000_b1 );
xor ( \2104_b0 , \1986_b0 , w_6636 );
not ( w_6636 , w_6637 );
and ( w_6637 , \2000_b1 , \2000_b0 );
or ( \2105_b1 , \2104_b1 , w_6638 );
xor ( \2105_b0 , \2104_b0 , w_6640 );
not ( w_6640 , w_6641 );
and ( w_6641 , w_6638 , w_6639 );
buf ( w_6638 , \2019_b1 );
not ( w_6638 , w_6642 );
not ( w_6639 , w_6643 );
and ( w_6642 , w_6643 , \2019_b0 );
or ( \2106_b1 , \2103_b1 , \2105_b1 );
xor ( \2106_b0 , \2103_b0 , w_6644 );
not ( w_6644 , w_6645 );
and ( w_6645 , \2105_b1 , \2105_b0 );
or ( \2107_b1 , \2042_b1 , \2064_b1 );
xor ( \2107_b0 , \2042_b0 , w_6646 );
not ( w_6646 , w_6647 );
and ( w_6647 , \2064_b1 , \2064_b0 );
or ( \2108_b1 , \2107_b1 , \2067_b1 );
not ( \2067_b1 , w_6648 );
and ( \2108_b0 , \2107_b0 , w_6649 );
and ( w_6648 , w_6649 , \2067_b0 );
or ( \2109_b1 , \2042_b1 , \2064_b1 );
not ( \2064_b1 , w_6650 );
and ( \2109_b0 , \2042_b0 , w_6651 );
and ( w_6650 , w_6651 , \2064_b0 );
or ( \2110_b1 , \2108_b1 , w_6652 );
or ( \2110_b0 , \2108_b0 , \2109_b0 );
not ( \2109_b0 , w_6653 );
and ( w_6653 , w_6652 , \2109_b1 );
or ( \2111_b1 , \2106_b1 , \2110_b1 );
xor ( \2111_b0 , \2106_b0 , w_6654 );
not ( w_6654 , w_6655 );
and ( w_6655 , \2110_b1 , \2110_b0 );
or ( \2112_b1 , \2101_b1 , w_6657 );
not ( w_6657 , w_6658 );
and ( \2112_b0 , \2101_b0 , w_6659 );
and ( w_6658 ,  , w_6659 );
buf ( w_6657 , \2111_b1 );
not ( w_6657 , w_6660 );
not (  , w_6661 );
and ( w_6660 , w_6661 , \2111_b0 );
or ( \2113_b1 , \2031_b1 , w_6663 );
not ( w_6663 , w_6664 );
and ( \2113_b0 , \2031_b0 , w_6665 );
and ( w_6664 ,  , w_6665 );
buf ( w_6663 , \2112_b1 );
not ( w_6663 , w_6666 );
not (  , w_6667 );
and ( w_6666 , w_6667 , \2112_b0 );
or ( \2114_b1 , \1955_b1 , w_6669 );
not ( w_6669 , w_6670 );
and ( \2114_b0 , \1955_b0 , w_6671 );
and ( w_6670 ,  , w_6671 );
buf ( w_6669 , \2113_b1 );
not ( w_6669 , w_6672 );
not (  , w_6673 );
and ( w_6672 , w_6673 , \2113_b0 );
buf ( \2115_b1 , \2114_b1 );
not ( \2115_b1 , w_6674 );
not ( \2115_b0 , w_6675 );
and ( w_6674 , w_6675 , \2114_b0 );
or ( \2116_b1 , \1149_b1 , w_6676 );
or ( \2116_b0 , \1149_b0 , \1156_b0 );
not ( \1156_b0 , w_6677 );
and ( w_6677 , w_6676 , \1156_b1 );
buf ( \2117_b1 , \2116_b1 );
not ( \2117_b1 , w_6678 );
not ( \2117_b0 , w_6679 );
and ( w_6678 , w_6679 , \2116_b0 );
buf ( \2118_b1 , \1101_b1 );
not ( \2118_b1 , w_6680 );
not ( \2118_b0 , w_6681 );
and ( w_6680 , w_6681 , \1101_b0 );
or ( \2119_b1 , \2117_b1 , w_6682 );
or ( \2119_b0 , \2117_b0 , \2118_b0 );
not ( \2118_b0 , w_6683 );
and ( w_6683 , w_6682 , \2118_b1 );
or ( \2120_b1 , \2119_b1 , w_6685 );
not ( w_6685 , w_6686 );
and ( \2120_b0 , \2119_b0 , w_6687 );
and ( w_6686 ,  , w_6687 );
buf ( w_6685 , \1158_b1 );
not ( w_6685 , w_6688 );
not (  , w_6689 );
and ( w_6688 , w_6689 , \1158_b0 );
buf ( \2121_b1 , \2120_b1 );
not ( \2121_b1 , w_6690 );
not ( \2121_b0 , w_6691 );
and ( w_6690 , w_6691 , \2120_b0 );
buf ( \2122_b1 , \1138_b1 );
not ( \2122_b1 , w_6692 );
not ( \2122_b0 , w_6693 );
and ( w_6692 , w_6693 , \1138_b0 );
buf ( \2123_b1 , \948_b1 );
not ( \2123_b1 , w_6694 );
not ( \2123_b0 , w_6695 );
and ( w_6694 , w_6695 , \948_b0 );
or ( \2124_b1 , \2122_b1 , w_6696 );
or ( \2124_b0 , \2122_b0 , \2123_b0 );
not ( \2123_b0 , w_6697 );
and ( w_6697 , w_6696 , \2123_b1 );
or ( \2125_b1 , \951_b1 , w_6699 );
not ( w_6699 , w_6700 );
and ( \2125_b0 , \951_b0 , w_6701 );
and ( w_6700 ,  , w_6701 );
buf ( w_6699 , \2072_b1 );
not ( w_6699 , w_6702 );
not (  , w_6703 );
and ( w_6702 , w_6703 , \2072_b0 );
or ( \2126_b1 , \2124_b1 , w_6705 );
not ( w_6705 , w_6706 );
and ( \2126_b0 , \2124_b0 , w_6707 );
and ( w_6706 ,  , w_6707 );
buf ( w_6705 , \2125_b1 );
not ( w_6705 , w_6708 );
not (  , w_6709 );
and ( w_6708 , w_6709 , \2125_b0 );
buf ( \2127_b1 , \2126_b1 );
not ( \2127_b1 , w_6710 );
not ( \2127_b0 , w_6711 );
and ( w_6710 , w_6711 , \2126_b0 );
or ( \2128_b1 , \1108_b1 , w_6713 );
not ( w_6713 , w_6714 );
and ( \2128_b0 , \1108_b0 , w_6715 );
and ( w_6714 ,  , w_6715 );
buf ( w_6713 , \1113_b1 );
not ( w_6713 , w_6716 );
not (  , w_6717 );
and ( w_6716 , w_6717 , \1113_b0 );
buf ( \2129_b1 , \2128_b1 );
not ( \2129_b1 , w_6718 );
not ( \2129_b0 , w_6719 );
and ( w_6718 , w_6719 , \2128_b0 );
buf ( \2130_b1 , \2129_b1 );
not ( \2130_b1 , w_6720 );
not ( \2130_b0 , w_6721 );
and ( w_6720 , w_6721 , \2129_b0 );
or ( \2131_b1 , \2127_b1 , w_6722 );
or ( \2131_b0 , \2127_b0 , \2130_b0 );
not ( \2130_b0 , w_6723 );
and ( w_6723 , w_6722 , \2130_b1 );
buf ( \2132_b1 , \2126_b1 );
not ( \2132_b1 , w_6724 );
not ( \2132_b0 , w_6725 );
and ( w_6724 , w_6725 , \2126_b0 );
buf ( \2133_b1 , \2132_b1 );
not ( \2133_b1 , w_6726 );
not ( \2133_b0 , w_6727 );
and ( w_6726 , w_6727 , \2132_b0 );
buf ( \2134_b1 , \2128_b1 );
not ( \2134_b1 , w_6728 );
not ( \2134_b0 , w_6729 );
and ( w_6728 , w_6729 , \2128_b0 );
or ( \2135_b1 , \2133_b1 , w_6730 );
or ( \2135_b0 , \2133_b0 , \2134_b0 );
not ( \2134_b0 , w_6731 );
and ( w_6731 , w_6730 , \2134_b1 );
buf ( \2136_b1 , \1145_b1 );
not ( \2136_b1 , w_6732 );
not ( \2136_b0 , w_6733 );
and ( w_6732 , w_6733 , \1145_b0 );
buf ( \2137_b1 , \1067_b1 );
not ( \2137_b1 , w_6734 );
not ( \2137_b0 , w_6735 );
and ( w_6734 , w_6735 , \1067_b0 );
or ( \2138_b1 , \2136_b1 , w_6736 );
or ( \2138_b0 , \2136_b0 , \2137_b0 );
not ( \2137_b0 , w_6737 );
and ( w_6737 , w_6736 , \2137_b1 );
or ( \2139_b1 , \976_b1 , w_6739 );
not ( w_6739 , w_6740 );
and ( \2139_b0 , \976_b0 , w_6741 );
and ( w_6740 ,  , w_6741 );
buf ( w_6739 , \2036_b1 );
not ( w_6739 , w_6742 );
not (  , w_6743 );
and ( w_6742 , w_6743 , \2036_b0 );
or ( \2140_b1 , \2138_b1 , w_6745 );
not ( w_6745 , w_6746 );
and ( \2140_b0 , \2138_b0 , w_6747 );
and ( w_6746 ,  , w_6747 );
buf ( w_6745 , \2139_b1 );
not ( w_6745 , w_6748 );
not (  , w_6749 );
and ( w_6748 , w_6749 , \2139_b0 );
or ( \2141_b1 , \2135_b1 , w_6751 );
not ( w_6751 , w_6752 );
and ( \2141_b0 , \2135_b0 , w_6753 );
and ( w_6752 ,  , w_6753 );
buf ( w_6751 , \2140_b1 );
not ( w_6751 , w_6754 );
not (  , w_6755 );
and ( w_6754 , w_6755 , \2140_b0 );
or ( \2142_b1 , \2131_b1 , w_6757 );
not ( w_6757 , w_6758 );
and ( \2142_b0 , \2131_b0 , w_6759 );
and ( w_6758 ,  , w_6759 );
buf ( w_6757 , \2141_b1 );
not ( w_6757 , w_6760 );
not (  , w_6761 );
and ( w_6760 , w_6761 , \2141_b0 );
buf ( \2143_b1 , \2142_b1 );
not ( \2143_b1 , w_6762 );
not ( \2143_b0 , w_6763 );
and ( w_6762 , w_6763 , \2142_b0 );
or ( \2144_b1 , \2061_b1 , \2048_b1 );
xor ( \2144_b0 , \2061_b0 , w_6764 );
not ( w_6764 , w_6765 );
and ( w_6765 , \2048_b1 , \2048_b0 );
or ( \2145_b1 , \2144_b1 , w_6766 );
xor ( \2145_b0 , \2144_b0 , w_6768 );
not ( w_6768 , w_6769 );
and ( w_6769 , w_6766 , w_6767 );
buf ( w_6766 , \2054_b1 );
not ( w_6766 , w_6770 );
not ( w_6767 , w_6771 );
and ( w_6770 , w_6771 , \2054_b0 );
buf ( \2146_b1 , \2145_b1 );
not ( \2146_b1 , w_6772 );
not ( \2146_b0 , w_6773 );
and ( w_6772 , w_6773 , \2145_b0 );
or ( \2147_b1 , \2143_b1 , w_6774 );
or ( \2147_b0 , \2143_b0 , \2146_b0 );
not ( \2146_b0 , w_6775 );
and ( w_6775 , w_6774 , \2146_b1 );
or ( \2148_b1 , \2142_b1 , w_6776 );
or ( \2148_b0 , \2142_b0 , \2145_b0 );
not ( \2145_b0 , w_6777 );
and ( w_6777 , w_6776 , \2145_b1 );
or ( \2149_b1 , \2147_b1 , w_6779 );
not ( w_6779 , w_6780 );
and ( \2149_b0 , \2147_b0 , w_6781 );
and ( w_6780 ,  , w_6781 );
buf ( w_6779 , \2148_b1 );
not ( w_6779 , w_6782 );
not (  , w_6783 );
and ( w_6782 , w_6783 , \2148_b0 );
or ( \2150_b1 , \2077_b1 , \2092_b1 );
xor ( \2150_b0 , \2077_b0 , w_6784 );
not ( w_6784 , w_6785 );
and ( w_6785 , \2092_b1 , \2092_b0 );
or ( \2151_b1 , \2150_b1 , \2094_b1 );
xor ( \2151_b0 , \2150_b0 , w_6786 );
not ( w_6786 , w_6787 );
and ( w_6787 , \2094_b1 , \2094_b0 );
or ( \2152_b1 , \2149_b1 , \2151_b1 );
xor ( \2152_b0 , \2149_b0 , w_6788 );
not ( w_6788 , w_6789 );
and ( w_6789 , \2151_b1 , \2151_b0 );
or ( \2153_b1 , \2078_b1 , \2083_b1 );
xor ( \2153_b0 , \2078_b0 , w_6790 );
not ( w_6790 , w_6791 );
and ( w_6791 , \2083_b1 , \2083_b0 );
or ( \2154_b1 , \2153_b1 , \2089_b1 );
xor ( \2154_b0 , \2153_b0 , w_6792 );
not ( w_6792 , w_6793 );
and ( w_6793 , \2089_b1 , \2089_b0 );
or ( \2155_b1 , \1133_b1 , \1140_b1 );
xor ( \2155_b0 , \1133_b0 , w_6794 );
not ( w_6794 , w_6795 );
and ( w_6795 , \1140_b1 , \1140_b0 );
or ( \2156_b1 , \2155_b1 , \1147_b1 );
not ( \1147_b1 , w_6796 );
and ( \2156_b0 , \2155_b0 , w_6797 );
and ( w_6796 , w_6797 , \1147_b0 );
or ( \2157_b1 , \1133_b1 , \1140_b1 );
not ( \1140_b1 , w_6798 );
and ( \2157_b0 , \1133_b0 , w_6799 );
and ( w_6798 , w_6799 , \1140_b0 );
or ( \2158_b1 , \2156_b1 , w_6800 );
or ( \2158_b0 , \2156_b0 , \2157_b0 );
not ( \2157_b0 , w_6801 );
and ( w_6801 , w_6800 , \2157_b1 );
or ( \2159_b1 , \2154_b1 , \2158_b1 );
xor ( \2159_b0 , \2154_b0 , w_6802 );
not ( w_6802 , w_6803 );
and ( w_6803 , \2158_b1 , \2158_b0 );
or ( \2160_b1 , \2126_b1 , \2128_b1 );
xor ( \2160_b0 , \2126_b0 , w_6804 );
not ( w_6804 , w_6805 );
and ( w_6805 , \2128_b1 , \2128_b0 );
or ( \2161_b1 , \2160_b1 , w_6806 );
xor ( \2161_b0 , \2160_b0 , w_6808 );
not ( w_6808 , w_6809 );
and ( w_6809 , w_6806 , w_6807 );
buf ( w_6806 , \2140_b1 );
not ( w_6806 , w_6810 );
not ( w_6807 , w_6811 );
and ( w_6810 , w_6811 , \2140_b0 );
or ( \2162_b1 , \2159_b1 , \2161_b1 );
not ( \2161_b1 , w_6812 );
and ( \2162_b0 , \2159_b0 , w_6813 );
and ( w_6812 , w_6813 , \2161_b0 );
or ( \2163_b1 , \2154_b1 , \2158_b1 );
not ( \2158_b1 , w_6814 );
and ( \2163_b0 , \2154_b0 , w_6815 );
and ( w_6814 , w_6815 , \2158_b0 );
or ( \2164_b1 , \2162_b1 , w_6816 );
or ( \2164_b0 , \2162_b0 , \2163_b0 );
not ( \2163_b0 , w_6817 );
and ( w_6817 , w_6816 , \2163_b1 );
or ( \2165_b1 , \2152_b1 , w_6819 );
not ( w_6819 , w_6820 );
and ( \2165_b0 , \2152_b0 , w_6821 );
and ( w_6820 ,  , w_6821 );
buf ( w_6819 , \2164_b1 );
not ( w_6819 , w_6822 );
not (  , w_6823 );
and ( w_6822 , w_6823 , \2164_b0 );
or ( \2166_b1 , \1117_b1 , \1121_b1 );
xor ( \2166_b0 , \1117_b0 , w_6824 );
not ( w_6824 , w_6825 );
and ( w_6825 , \1121_b1 , \1121_b0 );
or ( \2167_b1 , \2166_b1 , \1148_b1 );
not ( \1148_b1 , w_6826 );
and ( \2167_b0 , \2166_b0 , w_6827 );
and ( w_6826 , w_6827 , \1148_b0 );
or ( \2168_b1 , \1117_b1 , \1121_b1 );
not ( \1121_b1 , w_6828 );
and ( \2168_b0 , \1117_b0 , w_6829 );
and ( w_6828 , w_6829 , \1121_b0 );
or ( \2169_b1 , \2167_b1 , w_6830 );
or ( \2169_b0 , \2167_b0 , \2168_b0 );
not ( \2168_b0 , w_6831 );
and ( w_6831 , w_6830 , \2168_b1 );
or ( \2170_b1 , \2154_b1 , \2158_b1 );
xor ( \2170_b0 , \2154_b0 , w_6832 );
not ( w_6832 , w_6833 );
and ( w_6833 , \2158_b1 , \2158_b0 );
or ( \2171_b1 , \2170_b1 , \2161_b1 );
xor ( \2171_b0 , \2170_b0 , w_6834 );
not ( w_6834 , w_6835 );
and ( w_6835 , \2161_b1 , \2161_b0 );
or ( \2172_b1 , \2169_b1 , w_6837 );
not ( w_6837 , w_6838 );
and ( \2172_b0 , \2169_b0 , w_6839 );
and ( w_6838 ,  , w_6839 );
buf ( w_6837 , \2171_b1 );
not ( w_6837 , w_6840 );
not (  , w_6841 );
and ( w_6840 , w_6841 , \2171_b0 );
or ( \2173_b1 , \2165_b1 , w_6843 );
not ( w_6843 , w_6844 );
and ( \2173_b0 , \2165_b0 , w_6845 );
and ( w_6844 ,  , w_6845 );
buf ( w_6843 , \2172_b1 );
not ( w_6843 , w_6846 );
not (  , w_6847 );
and ( w_6846 , w_6847 , \2172_b0 );
buf ( \2174_b1 , \2173_b1 );
not ( \2174_b1 , w_6848 );
not ( \2174_b0 , w_6849 );
and ( w_6848 , w_6849 , \2173_b0 );
or ( \2175_b1 , \2121_b1 , w_6850 );
or ( \2175_b0 , \2121_b0 , \2174_b0 );
not ( \2174_b0 , w_6851 );
and ( w_6851 , w_6850 , \2174_b1 );
or ( \2176_b1 , \2070_b1 , \2097_b1 );
xor ( \2176_b0 , \2070_b0 , w_6852 );
not ( w_6852 , w_6853 );
and ( w_6853 , \2097_b1 , \2097_b0 );
or ( \2177_b1 , \2176_b1 , w_6854 );
xor ( \2177_b0 , \2176_b0 , w_6856 );
not ( w_6856 , w_6857 );
and ( w_6857 , w_6854 , w_6855 );
buf ( w_6854 , \2068_b1 );
not ( w_6854 , w_6858 );
not ( w_6855 , w_6859 );
and ( w_6858 , w_6859 , \2068_b0 );
buf ( \2178_b1 , \2142_b1 );
not ( \2178_b1 , w_6860 );
not ( \2178_b0 , w_6861 );
and ( w_6860 , w_6861 , \2142_b0 );
or ( \2179_b1 , \2178_b1 , w_6863 );
not ( w_6863 , w_6864 );
and ( \2179_b0 , \2178_b0 , w_6865 );
and ( w_6864 ,  , w_6865 );
buf ( w_6863 , \2145_b1 );
not ( w_6863 , w_6866 );
not (  , w_6867 );
and ( w_6866 , w_6867 , \2145_b0 );
buf ( \2180_b1 , \2179_b1 );
not ( \2180_b1 , w_6868 );
not ( \2180_b0 , w_6869 );
and ( w_6868 , w_6869 , \2179_b0 );
buf ( \2181_b1 , \2151_b1 );
not ( \2181_b1 , w_6870 );
not ( \2181_b0 , w_6871 );
and ( w_6870 , w_6871 , \2151_b0 );
or ( \2182_b1 , \2180_b1 , w_6872 );
or ( \2182_b0 , \2180_b0 , \2181_b0 );
not ( \2181_b0 , w_6873 );
and ( w_6873 , w_6872 , \2181_b1 );
buf ( \2183_b1 , \2145_b1 );
not ( \2183_b1 , w_6874 );
not ( \2183_b0 , w_6875 );
and ( w_6874 , w_6875 , \2145_b0 );
or ( \2184_b1 , \2183_b1 , w_6877 );
not ( w_6877 , w_6878 );
and ( \2184_b0 , \2183_b0 , w_6879 );
and ( w_6878 ,  , w_6879 );
buf ( w_6877 , \2142_b1 );
not ( w_6877 , w_6880 );
not (  , w_6881 );
and ( w_6880 , w_6881 , \2142_b0 );
or ( \2185_b1 , \2182_b1 , w_6883 );
not ( w_6883 , w_6884 );
and ( \2185_b0 , \2182_b0 , w_6885 );
and ( w_6884 ,  , w_6885 );
buf ( w_6883 , \2184_b1 );
not ( w_6883 , w_6886 );
not (  , w_6887 );
and ( w_6886 , w_6887 , \2184_b0 );
buf ( \2186_b1 , \2185_b1 );
not ( \2186_b1 , w_6888 );
not ( \2186_b0 , w_6889 );
and ( w_6888 , w_6889 , \2185_b0 );
or ( \2187_b1 , \2177_b1 , w_6891 );
not ( w_6891 , w_6892 );
and ( \2187_b0 , \2177_b0 , w_6893 );
and ( w_6892 ,  , w_6893 );
buf ( w_6891 , \2186_b1 );
not ( w_6891 , w_6894 );
not (  , w_6895 );
and ( w_6894 , w_6895 , \2186_b0 );
or ( \2188_b1 , \2171_b1 , w_6897 );
not ( w_6897 , w_6898 );
and ( \2188_b0 , \2171_b0 , w_6899 );
and ( w_6898 ,  , w_6899 );
buf ( w_6897 , \2169_b1 );
not ( w_6897 , w_6900 );
not (  , w_6901 );
and ( w_6900 , w_6901 , \2169_b0 );
or ( \2189_b1 , \2165_b1 , w_6902 );
or ( \2189_b0 , \2165_b0 , \2188_b0 );
not ( \2188_b0 , w_6903 );
and ( w_6903 , w_6902 , \2188_b1 );
or ( \2190_b1 , \2152_b1 , w_6905 );
not ( w_6905 , w_6906 );
and ( \2190_b0 , \2152_b0 , w_6907 );
and ( w_6906 ,  , w_6907 );
buf ( w_6905 , \2164_b1 );
not ( w_6905 , w_6908 );
not (  , w_6909 );
and ( w_6908 , w_6909 , \2164_b0 );
or ( \2191_b1 , \2189_b1 , w_6911 );
not ( w_6911 , w_6912 );
and ( \2191_b0 , \2189_b0 , w_6913 );
and ( w_6912 ,  , w_6913 );
buf ( w_6911 , \2190_b1 );
not ( w_6911 , w_6914 );
not (  , w_6915 );
and ( w_6914 , w_6915 , \2190_b0 );
or ( \2192_b1 , \2187_b1 , w_6917 );
not ( w_6917 , w_6918 );
and ( \2192_b0 , \2187_b0 , w_6919 );
and ( w_6918 ,  , w_6919 );
buf ( w_6917 , \2191_b1 );
not ( w_6917 , w_6920 );
not (  , w_6921 );
and ( w_6920 , w_6921 , \2191_b0 );
or ( \2193_b1 , \2175_b1 , w_6923 );
not ( w_6923 , w_6924 );
and ( \2193_b0 , \2175_b0 , w_6925 );
and ( w_6924 ,  , w_6925 );
buf ( w_6923 , \2192_b1 );
not ( w_6923 , w_6926 );
not (  , w_6927 );
and ( w_6926 , w_6927 , \2192_b0 );
buf ( \2194_b1 , \2193_b1 );
not ( \2194_b1 , w_6928 );
not ( \2194_b0 , w_6929 );
and ( w_6928 , w_6929 , \2193_b0 );
or ( \2195_b1 , \1964_b1 , \2024_b1 );
xor ( \2195_b0 , \1964_b0 , w_6930 );
not ( w_6930 , w_6931 );
and ( w_6931 , \2024_b1 , \2024_b0 );
or ( \2196_b1 , \2195_b1 , \2027_b1 );
xor ( \2196_b0 , \2195_b0 , w_6932 );
not ( w_6932 , w_6933 );
and ( w_6933 , \2027_b1 , \2027_b0 );
or ( \2197_b1 , \2110_b1 , w_6935 );
not ( w_6935 , w_6936 );
and ( \2197_b0 , \2110_b0 , w_6937 );
and ( w_6936 ,  , w_6937 );
buf ( w_6935 , \2103_b1 );
not ( w_6935 , w_6938 );
not (  , w_6939 );
and ( w_6938 , w_6939 , \2103_b0 );
buf ( \2198_b1 , \2197_b1 );
not ( \2198_b1 , w_6940 );
not ( \2198_b0 , w_6941 );
and ( w_6940 , w_6941 , \2197_b0 );
buf ( \2199_b1 , \2110_b1 );
not ( \2199_b1 , w_6942 );
not ( \2199_b0 , w_6943 );
and ( w_6942 , w_6943 , \2110_b0 );
buf ( \2200_b1 , \2103_b1 );
not ( \2200_b1 , w_6944 );
not ( \2200_b0 , w_6945 );
and ( w_6944 , w_6945 , \2103_b0 );
or ( \2201_b1 , \2199_b1 , \2200_b1 );
not ( \2200_b1 , w_6946 );
and ( \2201_b0 , \2199_b0 , w_6947 );
and ( w_6946 , w_6947 , \2200_b0 );
buf ( \2202_b1 , \2105_b1 );
buf ( \2202_b0 , \2105_b0 );
or ( \2203_b1 , \2201_b1 , w_6949 );
not ( w_6949 , w_6950 );
and ( \2203_b0 , \2201_b0 , w_6951 );
and ( w_6950 ,  , w_6951 );
buf ( w_6949 , \2202_b1 );
not ( w_6949 , w_6952 );
not (  , w_6953 );
and ( w_6952 , w_6953 , \2202_b0 );
or ( \2204_b1 , \2198_b1 , w_6955 );
not ( w_6955 , w_6956 );
and ( \2204_b0 , \2198_b0 , w_6957 );
and ( w_6956 ,  , w_6957 );
buf ( w_6955 , \2203_b1 );
not ( w_6955 , w_6958 );
not (  , w_6959 );
and ( w_6958 , w_6959 , \2203_b0 );
or ( \2205_b1 , \2196_b1 , w_6961 );
not ( w_6961 , w_6962 );
and ( \2205_b0 , \2196_b0 , w_6963 );
and ( w_6962 ,  , w_6963 );
buf ( w_6961 , \2204_b1 );
not ( w_6961 , w_6964 );
not (  , w_6965 );
and ( w_6964 , w_6965 , \2204_b0 );
or ( \2206_b1 , \2177_b1 , w_6967 );
not ( w_6967 , w_6968 );
and ( \2206_b0 , \2177_b0 , w_6969 );
and ( w_6968 ,  , w_6969 );
buf ( w_6967 , \2186_b1 );
not ( w_6967 , w_6970 );
not (  , w_6971 );
and ( w_6970 , w_6971 , \2186_b0 );
or ( \2207_b1 , \2205_b1 , \2206_b1 );
not ( \2206_b1 , w_6972 );
and ( \2207_b0 , \2205_b0 , w_6973 );
and ( w_6972 , w_6973 , \2206_b0 );
buf ( \2208_b1 , \2207_b1 );
not ( \2208_b1 , w_6974 );
not ( \2208_b0 , w_6975 );
and ( w_6974 , w_6975 , \2207_b0 );
or ( \2209_b1 , \2194_b1 , w_6976 );
or ( \2209_b0 , \2194_b0 , \2208_b0 );
not ( \2208_b0 , w_6977 );
and ( w_6977 , w_6976 , \2208_b1 );
buf ( \2210_b1 , \2100_b1 );
not ( \2210_b1 , w_6978 );
not ( \2210_b0 , w_6979 );
and ( w_6978 , w_6979 , \2100_b0 );
or ( \2211_b1 , \2210_b1 , w_6981 );
not ( w_6981 , w_6982 );
and ( \2211_b0 , \2210_b0 , w_6983 );
and ( w_6982 ,  , w_6983 );
buf ( w_6981 , \2111_b1 );
not ( w_6981 , w_6984 );
not (  , w_6985 );
and ( w_6984 , w_6985 , \2111_b0 );
or ( \2212_b1 , \2205_b1 , w_6987 );
not ( w_6987 , w_6988 );
and ( \2212_b0 , \2205_b0 , w_6989 );
and ( w_6988 ,  , w_6989 );
buf ( w_6987 , \2211_b1 );
not ( w_6987 , w_6990 );
not (  , w_6991 );
and ( w_6990 , w_6991 , \2211_b0 );
or ( \2213_b1 , \2209_b1 , w_6993 );
not ( w_6993 , w_6994 );
and ( \2213_b0 , \2209_b0 , w_6995 );
and ( w_6994 ,  , w_6995 );
buf ( w_6993 , \2212_b1 );
not ( w_6993 , w_6996 );
not (  , w_6997 );
and ( w_6996 , w_6997 , \2212_b0 );
buf ( \2214_b1 , \2213_b1 );
not ( \2214_b1 , w_6998 );
not ( \2214_b0 , w_6999 );
and ( w_6998 , w_6999 , \2213_b0 );
or ( \2215_b1 , \2115_b1 , w_7000 );
or ( \2215_b0 , \2115_b0 , \2214_b0 );
not ( \2214_b0 , w_7001 );
and ( w_7001 , w_7000 , \2214_b1 );
buf ( \2216_b1 , \2030_b1 );
not ( \2216_b1 , w_7002 );
not ( \2216_b0 , w_7003 );
and ( w_7002 , w_7003 , \2030_b0 );
buf ( \2217_b1 , \2216_b1 );
not ( \2217_b1 , w_7004 );
not ( \2217_b0 , w_7005 );
and ( w_7004 , w_7005 , \2216_b0 );
buf ( \2218_b1 , \1962_b1 );
not ( \2218_b1 , w_7006 );
not ( \2218_b0 , w_7007 );
and ( w_7006 , w_7007 , \1962_b0 );
buf ( \2219_b1 , \2218_b1 );
not ( \2219_b1 , w_7008 );
not ( \2219_b0 , w_7009 );
and ( w_7008 , w_7009 , \2218_b0 );
or ( \2220_b1 , \2217_b1 , w_7010 );
or ( \2220_b0 , \2217_b0 , \2219_b0 );
not ( \2219_b0 , w_7011 );
and ( w_7011 , w_7010 , \2219_b1 );
or ( \2221_b1 , \2196_b1 , w_7013 );
not ( w_7013 , w_7014 );
and ( \2221_b0 , \2196_b0 , w_7015 );
and ( w_7014 ,  , w_7015 );
buf ( w_7013 , \2204_b1 );
not ( w_7013 , w_7016 );
not (  , w_7017 );
and ( w_7016 , w_7017 , \2204_b0 );
buf ( \2222_b1 , \2221_b1 );
not ( \2222_b1 , w_7018 );
not ( \2222_b0 , w_7019 );
and ( w_7018 , w_7019 , \2221_b0 );
or ( \2223_b1 , \2220_b1 , w_7021 );
not ( w_7021 , w_7022 );
and ( \2223_b0 , \2220_b0 , w_7023 );
and ( w_7022 ,  , w_7023 );
buf ( w_7021 , \2222_b1 );
not ( w_7021 , w_7024 );
not (  , w_7025 );
and ( w_7024 , w_7025 , \2222_b0 );
or ( \2225_b1 , \1908_b1 , w_7027 );
not ( w_7027 , w_7028 );
and ( \2225_b0 , \1908_b0 , w_7029 );
and ( w_7028 ,  , w_7029 );
buf ( w_7027 , \1953_b1 );
not ( w_7027 , w_7030 );
not (  , w_7031 );
and ( w_7030 , w_7031 , \1953_b0 );
or ( \2226_b1 , \2224_b1 , w_7033 );
not ( w_7033 , w_7034 );
and ( \2226_b0 , \2224_b0 , w_7035 );
and ( w_7034 ,  , w_7035 );
buf ( w_7033 , \2225_b1 );
not ( w_7033 , w_7036 );
not (  , w_7037 );
and ( w_7036 , w_7037 , \2225_b0 );
or ( \2227_b1 , \2215_b1 , w_7039 );
not ( w_7039 , w_7040 );
and ( \2227_b0 , \2215_b0 , w_7041 );
and ( w_7040 ,  , w_7041 );
buf ( w_7039 , \2226_b1 );
not ( w_7039 , w_7042 );
not (  , w_7043 );
and ( w_7042 , w_7043 , \2226_b0 );
buf ( \2228_b1 , \2227_b1 );
not ( \2228_b1 , w_7044 );
not ( \2228_b0 , w_7045 );
and ( w_7044 , w_7045 , \2227_b0 );
or ( \2229_b1 , \1902_b1 , w_7046 );
or ( \2229_b0 , \1902_b0 , \2228_b0 );
not ( \2228_b0 , w_7047 );
and ( w_7047 , w_7046 , \2228_b1 );
or ( \2230_b1 , \1901_b1 , w_7048 );
or ( \2230_b0 , \1901_b0 , \2227_b0 );
not ( \2227_b0 , w_7049 );
and ( w_7049 , w_7048 , \2227_b1 );
or ( \2231_b1 , \2229_b1 , w_7051 );
not ( w_7051 , w_7052 );
and ( \2231_b0 , \2229_b0 , w_7053 );
and ( w_7052 ,  , w_7053 );
buf ( w_7051 , \2230_b1 );
not ( w_7051 , w_7054 );
not (  , w_7055 );
and ( w_7054 , w_7055 , \2230_b0 );
buf ( \2232_b1 , \2231_b1 );
not ( \2232_b1 , w_7056 );
not ( \2232_b0 , w_7057 );
and ( w_7056 , w_7057 , \2231_b0 );
or ( \2233_b1 , \1530_b1 , w_7058 );
or ( \2233_b0 , \1530_b0 , \2232_b0 );
not ( \2232_b0 , w_7059 );
and ( w_7059 , w_7058 , \2232_b1 );
or ( \2234_b1 , \b[2]_b1 , \c[11]_b1 );
xor ( \2234_b0 , \b[2]_b0 , w_7060 );
not ( w_7060 , w_7061 );
and ( w_7061 , \c[11]_b1 , \c[11]_b0 );
buf ( \2235_b1 , \2234_b1 );
not ( \2235_b1 , w_7062 );
not ( \2235_b0 , w_7063 );
and ( w_7062 , w_7063 , \2234_b0 );
or ( \2236_b1 , \c[10]_b1 , \c[9]_b1 );
xor ( \2236_b0 , \c[10]_b0 , w_7064 );
not ( w_7064 , w_7065 );
and ( w_7065 , \c[9]_b1 , \c[9]_b0 );
or ( \2237_b1 , \c[11]_b1 , w_7066 );
xor ( \2237_b0 , \c[11]_b0 , w_7068 );
not ( w_7068 , w_7069 );
and ( w_7069 , w_7066 , w_7067 );
buf ( w_7066 , \c[10]_b1 );
not ( w_7066 , w_7070 );
not ( w_7067 , w_7071 );
and ( w_7070 , w_7071 , \c[10]_b0 );
or ( \2238_b1 , \2236_b1 , w_7073 );
not ( w_7073 , w_7074 );
and ( \2238_b0 , \2236_b0 , w_7075 );
and ( w_7074 ,  , w_7075 );
buf ( w_7073 , \2237_b1 );
not ( w_7073 , w_7076 );
not (  , w_7077 );
and ( w_7076 , w_7077 , \2237_b0 );
buf ( \2239_b1 , \2238_b1 );
not ( \2239_b1 , w_7078 );
not ( \2239_b0 , w_7079 );
and ( w_7078 , w_7079 , \2238_b0 );
or ( \2240_b1 , \2235_b1 , w_7080 );
or ( \2240_b0 , \2235_b0 , \2239_b0 );
not ( \2239_b0 , w_7081 );
and ( w_7081 , w_7080 , \2239_b1 );
or ( \2241_b1 , \c[11]_b1 , \b[3]_b1 );
xor ( \2241_b0 , \c[11]_b0 , w_7082 );
not ( w_7082 , w_7083 );
and ( w_7083 , \b[3]_b1 , \b[3]_b0 );
or ( \2242_b1 , \2236_b1 , w_7085 );
not ( w_7085 , w_7086 );
and ( \2242_b0 , \2236_b0 , w_7087 );
and ( w_7086 ,  , w_7087 );
buf ( w_7085 , \2241_b1 );
not ( w_7085 , w_7088 );
not (  , w_7089 );
and ( w_7088 , w_7089 , \2241_b0 );
or ( \2243_b1 , \2240_b1 , w_7091 );
not ( w_7091 , w_7092 );
and ( \2243_b0 , \2240_b0 , w_7093 );
and ( w_7092 ,  , w_7093 );
buf ( w_7091 , \2242_b1 );
not ( w_7091 , w_7094 );
not (  , w_7095 );
and ( w_7094 , w_7095 , \2242_b0 );
or ( \2244_b1 , \c[13]_b1 , \b[0]_b1 );
xor ( \2244_b0 , \c[13]_b0 , w_7096 );
not ( w_7096 , w_7097 );
and ( w_7097 , \b[0]_b1 , \b[0]_b0 );
buf ( \2245_b1 , \2244_b1 );
not ( \2245_b1 , w_7098 );
not ( \2245_b0 , w_7099 );
and ( w_7098 , w_7099 , \2244_b0 );
or ( \2246_b1 , \c[12]_b1 , \c[11]_b1 );
xor ( \2246_b0 , \c[12]_b0 , w_7100 );
not ( w_7100 , w_7101 );
and ( w_7101 , \c[11]_b1 , \c[11]_b0 );
buf ( \2247_b1 , \c[12]_b1 );
not ( \2247_b1 , w_7102 );
not ( \2247_b0 , w_7103 );
and ( w_7102 , w_7103 , \c[12]_b0 );
buf ( \2248_b1 , \c[13]_b1 );
not ( \2248_b1 , w_7104 );
not ( \2248_b0 , w_7105 );
and ( w_7104 , w_7105 , \c[13]_b0 );
or ( \2249_b1 , \2247_b1 , w_7106 );
or ( \2249_b0 , \2247_b0 , \2248_b0 );
not ( \2248_b0 , w_7107 );
and ( w_7107 , w_7106 , \2248_b1 );
or ( \2250_b1 , \c[13]_b1 , w_7108 );
or ( \2250_b0 , \c[13]_b0 , \c[12]_b0 );
not ( \c[12]_b0 , w_7109 );
and ( w_7109 , w_7108 , \c[12]_b1 );
or ( \2251_b1 , \2249_b1 , w_7111 );
not ( w_7111 , w_7112 );
and ( \2251_b0 , \2249_b0 , w_7113 );
and ( w_7112 ,  , w_7113 );
buf ( w_7111 , \2250_b1 );
not ( w_7111 , w_7114 );
not (  , w_7115 );
and ( w_7114 , w_7115 , \2250_b0 );
or ( \2252_b1 , \2246_b1 , w_7117 );
not ( w_7117 , w_7118 );
and ( \2252_b0 , \2246_b0 , w_7119 );
and ( w_7118 ,  , w_7119 );
buf ( w_7117 , \2251_b1 );
not ( w_7117 , w_7120 );
not (  , w_7121 );
and ( w_7120 , w_7121 , \2251_b0 );
buf ( \2253_b1 , \2252_b1 );
not ( \2253_b1 , w_7122 );
not ( \2253_b0 , w_7123 );
and ( w_7122 , w_7123 , \2252_b0 );
or ( \2254_b1 , \2245_b1 , w_7124 );
or ( \2254_b0 , \2245_b0 , \2253_b0 );
not ( \2253_b0 , w_7125 );
and ( w_7125 , w_7124 , \2253_b1 );
or ( \2255_b1 , \c[13]_b1 , \b[1]_b1 );
xor ( \2255_b0 , \c[13]_b0 , w_7126 );
not ( w_7126 , w_7127 );
and ( w_7127 , \b[1]_b1 , \b[1]_b0 );
or ( \2256_b1 , \2246_b1 , w_7129 );
not ( w_7129 , w_7130 );
and ( \2256_b0 , \2246_b0 , w_7131 );
and ( w_7130 ,  , w_7131 );
buf ( w_7129 , \2255_b1 );
not ( w_7129 , w_7132 );
not (  , w_7133 );
and ( w_7132 , w_7133 , \2255_b0 );
or ( \2257_b1 , \2254_b1 , w_7135 );
not ( w_7135 , w_7136 );
and ( \2257_b0 , \2254_b0 , w_7137 );
and ( w_7136 ,  , w_7137 );
buf ( w_7135 , \2256_b1 );
not ( w_7135 , w_7138 );
not (  , w_7139 );
and ( w_7138 , w_7139 , \2256_b0 );
buf ( \2258_b1 , \2257_b1 );
not ( \2258_b1 , w_7140 );
not ( \2258_b0 , w_7141 );
and ( w_7140 , w_7141 , \2257_b0 );
or ( \2259_b1 , \2243_b1 , \2258_b1 );
not ( \2258_b1 , w_7142 );
and ( \2259_b0 , \2243_b0 , w_7143 );
and ( w_7142 , w_7143 , \2258_b0 );
buf ( \2260_b1 , \2243_b1 );
not ( \2260_b1 , w_7144 );
not ( \2260_b0 , w_7145 );
and ( w_7144 , w_7145 , \2243_b0 );
or ( \2261_b1 , \2260_b1 , \2257_b1 );
not ( \2257_b1 , w_7146 );
and ( \2261_b0 , \2260_b0 , w_7147 );
and ( w_7146 , w_7147 , \2257_b0 );
or ( \2262_b1 , \2259_b1 , w_7148 );
or ( \2262_b0 , \2259_b0 , \2261_b0 );
not ( \2261_b0 , w_7149 );
and ( w_7149 , w_7148 , \2261_b1 );
or ( \2263_b1 , \b[8]_b1 , \c[5]_b1 );
xor ( \2263_b0 , \b[8]_b0 , w_7150 );
not ( w_7150 , w_7151 );
and ( w_7151 , \c[5]_b1 , \c[5]_b0 );
buf ( \2264_b1 , \2263_b1 );
not ( \2264_b1 , w_7152 );
not ( \2264_b0 , w_7153 );
and ( w_7152 , w_7153 , \2263_b0 );
buf ( \2265_b1 , \736_b1 );
buf ( \2265_b0 , \736_b0 );
buf ( \2266_b1 , \2265_b1 );
not ( \2266_b1 , w_7154 );
not ( \2266_b0 , w_7155 );
and ( w_7154 , w_7155 , \2265_b0 );
or ( \2267_b1 , \2264_b1 , w_7156 );
or ( \2267_b0 , \2264_b0 , \2266_b0 );
not ( \2266_b0 , w_7157 );
and ( w_7157 , w_7156 , \2266_b1 );
or ( \2268_b1 , \b[9]_b1 , \c[5]_b1 );
xor ( \2268_b0 , \b[9]_b0 , w_7158 );
not ( w_7158 , w_7159 );
and ( w_7159 , \c[5]_b1 , \c[5]_b0 );
or ( \2269_b1 , \739_b1 , w_7161 );
not ( w_7161 , w_7162 );
and ( \2269_b0 , \739_b0 , w_7163 );
and ( w_7162 ,  , w_7163 );
buf ( w_7161 , \2268_b1 );
not ( w_7161 , w_7164 );
not (  , w_7165 );
and ( w_7164 , w_7165 , \2268_b0 );
or ( \2270_b1 , \2267_b1 , w_7167 );
not ( w_7167 , w_7168 );
and ( \2270_b0 , \2267_b0 , w_7169 );
and ( w_7168 ,  , w_7169 );
buf ( w_7167 , \2269_b1 );
not ( w_7167 , w_7170 );
not (  , w_7171 );
and ( w_7170 , w_7171 , \2269_b0 );
buf ( \2271_b1 , \2270_b1 );
not ( \2271_b1 , w_7172 );
not ( \2271_b0 , w_7173 );
and ( w_7172 , w_7173 , \2270_b0 );
or ( \2272_b1 , \2262_b1 , \2271_b1 );
not ( \2271_b1 , w_7174 );
and ( \2272_b0 , \2262_b0 , w_7175 );
and ( w_7174 , w_7175 , \2271_b0 );
buf ( \2273_b1 , \2262_b1 );
not ( \2273_b1 , w_7176 );
not ( \2273_b0 , w_7177 );
and ( w_7176 , w_7177 , \2262_b0 );
or ( \2274_b1 , \2273_b1 , \2270_b1 );
not ( \2270_b1 , w_7178 );
and ( \2274_b0 , \2273_b0 , w_7179 );
and ( w_7178 , w_7179 , \2270_b0 );
or ( \2275_b1 , \2272_b1 , w_7181 );
not ( w_7181 , w_7182 );
and ( \2275_b0 , \2272_b0 , w_7183 );
and ( w_7182 ,  , w_7183 );
buf ( w_7181 , \2274_b1 );
not ( w_7181 , w_7184 );
not (  , w_7185 );
and ( w_7184 , w_7185 , \2274_b0 );
buf ( \2276_b1 , \2275_b1 );
not ( \2276_b1 , w_7186 );
not ( \2276_b0 , w_7187 );
and ( w_7186 , w_7187 , \2275_b0 );
or ( \2277_b1 , \b[4]_b1 , \c[9]_b1 );
xor ( \2277_b0 , \b[4]_b0 , w_7188 );
not ( w_7188 , w_7189 );
and ( w_7189 , \c[9]_b1 , \c[9]_b0 );
buf ( \2278_b1 , \2277_b1 );
not ( \2278_b1 , w_7190 );
not ( \2278_b0 , w_7191 );
and ( w_7190 , w_7191 , \2277_b0 );
or ( \2279_b1 , \c[9]_b1 , w_7192 );
xor ( \2279_b0 , \c[9]_b0 , w_7194 );
not ( w_7194 , w_7195 );
and ( w_7195 , w_7192 , w_7193 );
buf ( w_7192 , \c[8]_b1 );
not ( w_7192 , w_7196 );
not ( w_7193 , w_7197 );
and ( w_7196 , w_7197 , \c[8]_b0 );
or ( \2280_b1 , \c[8]_b1 , \c[7]_b1 );
xor ( \2280_b0 , \c[8]_b0 , w_7198 );
not ( w_7198 , w_7199 );
and ( w_7199 , \c[7]_b1 , \c[7]_b0 );
or ( \2281_b1 , \2279_b1 , w_7201 );
not ( w_7201 , w_7202 );
and ( \2281_b0 , \2279_b0 , w_7203 );
and ( w_7202 ,  , w_7203 );
buf ( w_7201 , \2280_b1 );
not ( w_7201 , w_7204 );
not (  , w_7205 );
and ( w_7204 , w_7205 , \2280_b0 );
buf ( \2282_b1 , \2281_b1 );
not ( \2282_b1 , w_7206 );
not ( \2282_b0 , w_7207 );
and ( w_7206 , w_7207 , \2281_b0 );
or ( \2283_b1 , \2278_b1 , w_7208 );
or ( \2283_b0 , \2278_b0 , \2282_b0 );
not ( \2282_b0 , w_7209 );
and ( w_7209 , w_7208 , \2282_b1 );
buf ( \2284_b1 , \2280_b1 );
buf ( \2284_b0 , \2280_b0 );
or ( \2285_b1 , \b[5]_b1 , \c[9]_b1 );
xor ( \2285_b0 , \b[5]_b0 , w_7210 );
not ( w_7210 , w_7211 );
and ( w_7211 , \c[9]_b1 , \c[9]_b0 );
or ( \2286_b1 , \2284_b1 , w_7213 );
not ( w_7213 , w_7214 );
and ( \2286_b0 , \2284_b0 , w_7215 );
and ( w_7214 ,  , w_7215 );
buf ( w_7213 , \2285_b1 );
not ( w_7213 , w_7216 );
not (  , w_7217 );
and ( w_7216 , w_7217 , \2285_b0 );
or ( \2287_b1 , \2283_b1 , w_7219 );
not ( w_7219 , w_7220 );
and ( \2287_b0 , \2283_b0 , w_7221 );
and ( w_7220 ,  , w_7221 );
buf ( w_7219 , \2286_b1 );
not ( w_7219 , w_7222 );
not (  , w_7223 );
and ( w_7222 , w_7223 , \2286_b0 );
or ( \2288_b1 , \b[7]_b1 , \c[7]_b1 );
xor ( \2288_b0 , \b[7]_b0 , w_7224 );
not ( w_7224 , w_7225 );
and ( w_7225 , \c[7]_b1 , \c[7]_b0 );
buf ( \2289_b1 , \2288_b1 );
not ( \2289_b1 , w_7226 );
not ( \2289_b0 , w_7227 );
and ( w_7226 , w_7227 , \2288_b0 );
buf ( \2290_b1 , \714_b1 );
not ( \2290_b1 , w_7228 );
not ( \2290_b0 , w_7229 );
and ( w_7228 , w_7229 , \714_b0 );
or ( \2291_b1 , \2289_b1 , w_7230 );
or ( \2291_b0 , \2289_b0 , \2290_b0 );
not ( \2290_b0 , w_7231 );
and ( w_7231 , w_7230 , \2290_b1 );
or ( \2292_b1 , \725_b1 , w_7233 );
not ( w_7233 , w_7234 );
and ( \2292_b0 , \725_b0 , w_7235 );
and ( w_7234 ,  , w_7235 );
buf ( w_7233 , \713_b1 );
not ( w_7233 , w_7236 );
not (  , w_7237 );
and ( w_7236 , w_7237 , \713_b0 );
or ( \2293_b1 , \b[6]_b1 , \c[7]_b1 );
xor ( \2293_b0 , \b[6]_b0 , w_7238 );
not ( w_7238 , w_7239 );
and ( w_7239 , \c[7]_b1 , \c[7]_b0 );
or ( \2294_b1 , \2292_b1 , w_7241 );
not ( w_7241 , w_7242 );
and ( \2294_b0 , \2292_b0 , w_7243 );
and ( w_7242 ,  , w_7243 );
buf ( w_7241 , \2293_b1 );
not ( w_7241 , w_7244 );
not (  , w_7245 );
and ( w_7244 , w_7245 , \2293_b0 );
or ( \2295_b1 , \2291_b1 , w_7247 );
not ( w_7247 , w_7248 );
and ( \2295_b0 , \2291_b0 , w_7249 );
and ( w_7248 ,  , w_7249 );
buf ( w_7247 , \2294_b1 );
not ( w_7247 , w_7250 );
not (  , w_7251 );
and ( w_7250 , w_7251 , \2294_b0 );
or ( \2296_b1 , \2287_b1 , \2295_b1 );
xor ( \2296_b0 , \2287_b0 , w_7252 );
not ( w_7252 , w_7253 );
and ( w_7253 , \2295_b1 , \2295_b0 );
or ( \2297_b1 , \b[10]_b1 , \c[3]_b1 );
xor ( \2297_b0 , \b[10]_b0 , w_7254 );
not ( w_7254 , w_7255 );
and ( w_7255 , \c[3]_b1 , \c[3]_b0 );
buf ( \2298_b1 , \2297_b1 );
not ( \2298_b1 , w_7256 );
not ( \2298_b0 , w_7257 );
and ( w_7256 , w_7257 , \2297_b0 );
buf ( \2299_b1 , \746_b1 );
not ( \2299_b1 , w_7258 );
not ( \2299_b0 , w_7259 );
and ( w_7258 , w_7259 , \746_b0 );
or ( \2300_b1 , \2298_b1 , w_7260 );
or ( \2300_b0 , \2298_b0 , \2299_b0 );
not ( \2299_b0 , w_7261 );
and ( w_7261 , w_7260 , \2299_b1 );
or ( \2301_b1 , \b[11]_b1 , \c[3]_b1 );
xor ( \2301_b0 , \b[11]_b0 , w_7262 );
not ( w_7262 , w_7263 );
and ( w_7263 , \c[3]_b1 , \c[3]_b0 );
or ( \2302_b1 , \702_b1 , w_7265 );
not ( w_7265 , w_7266 );
and ( \2302_b0 , \702_b0 , w_7267 );
and ( w_7266 ,  , w_7267 );
buf ( w_7265 , \2301_b1 );
not ( w_7265 , w_7268 );
not (  , w_7269 );
and ( w_7268 , w_7269 , \2301_b0 );
or ( \2303_b1 , \2300_b1 , w_7271 );
not ( w_7271 , w_7272 );
and ( \2303_b0 , \2300_b0 , w_7273 );
and ( w_7272 ,  , w_7273 );
buf ( w_7271 , \2302_b1 );
not ( w_7271 , w_7274 );
not (  , w_7275 );
and ( w_7274 , w_7275 , \2302_b0 );
or ( \2304_b1 , \2296_b1 , w_7276 );
xor ( \2304_b0 , \2296_b0 , w_7278 );
not ( w_7278 , w_7279 );
and ( w_7279 , w_7276 , w_7277 );
buf ( w_7276 , \2303_b1 );
not ( w_7276 , w_7280 );
not ( w_7277 , w_7281 );
and ( w_7280 , w_7281 , \2303_b0 );
buf ( \2305_b1 , \2304_b1 );
not ( \2305_b1 , w_7282 );
not ( \2305_b0 , w_7283 );
and ( w_7282 , w_7283 , \2304_b0 );
or ( \2306_b1 , \2276_b1 , w_7284 );
or ( \2306_b0 , \2276_b0 , \2305_b0 );
not ( \2305_b0 , w_7285 );
and ( w_7285 , w_7284 , \2305_b1 );
or ( \2307_b1 , \b[7]_b1 , \c[5]_b1 );
xor ( \2307_b0 , \b[7]_b0 , w_7286 );
not ( w_7286 , w_7287 );
and ( w_7287 , \c[5]_b1 , \c[5]_b0 );
buf ( \2308_b1 , \2307_b1 );
not ( \2308_b1 , w_7288 );
not ( \2308_b0 , w_7289 );
and ( w_7288 , w_7289 , \2307_b0 );
buf ( \2309_b1 , \2265_b1 );
not ( \2309_b1 , w_7290 );
not ( \2309_b0 , w_7291 );
and ( w_7290 , w_7291 , \2265_b0 );
or ( \2310_b1 , \2308_b1 , w_7292 );
or ( \2310_b0 , \2308_b0 , \2309_b0 );
not ( \2309_b0 , w_7293 );
and ( w_7293 , w_7292 , \2309_b1 );
or ( \2311_b1 , \739_b1 , w_7295 );
not ( w_7295 , w_7296 );
and ( \2311_b0 , \739_b0 , w_7297 );
and ( w_7296 ,  , w_7297 );
buf ( w_7295 , \2263_b1 );
not ( w_7295 , w_7298 );
not (  , w_7299 );
and ( w_7298 , w_7299 , \2263_b0 );
or ( \2312_b1 , \2310_b1 , w_7301 );
not ( w_7301 , w_7302 );
and ( \2312_b0 , \2310_b0 , w_7303 );
and ( w_7302 ,  , w_7303 );
buf ( w_7301 , \2311_b1 );
not ( w_7301 , w_7304 );
not (  , w_7305 );
and ( w_7304 , w_7305 , \2311_b0 );
buf ( \2313_b1 , \2312_b1 );
not ( \2313_b1 , w_7306 );
not ( \2313_b0 , w_7307 );
and ( w_7306 , w_7307 , \2312_b0 );
or ( \2314_b1 , \b[8]_b1 , \c[3]_b1 );
xor ( \2314_b0 , \b[8]_b0 , w_7308 );
not ( w_7308 , w_7309 );
and ( w_7309 , \c[3]_b1 , \c[3]_b0 );
buf ( \2315_b1 , \2314_b1 );
not ( \2315_b1 , w_7310 );
not ( \2315_b0 , w_7311 );
and ( w_7310 , w_7311 , \2314_b0 );
buf ( \2316_b1 , \746_b1 );
not ( \2316_b1 , w_7312 );
not ( \2316_b0 , w_7313 );
and ( w_7312 , w_7313 , \746_b0 );
or ( \2317_b1 , \2315_b1 , w_7314 );
or ( \2317_b0 , \2315_b0 , \2316_b0 );
not ( \2316_b0 , w_7315 );
and ( w_7315 , w_7314 , \2316_b1 );
or ( \2318_b1 , \b[9]_b1 , \c[3]_b1 );
xor ( \2318_b0 , \b[9]_b0 , w_7316 );
not ( w_7316 , w_7317 );
and ( w_7317 , \c[3]_b1 , \c[3]_b0 );
or ( \2319_b1 , \702_b1 , w_7319 );
not ( w_7319 , w_7320 );
and ( \2319_b0 , \702_b0 , w_7321 );
and ( w_7320 ,  , w_7321 );
buf ( w_7319 , \2318_b1 );
not ( w_7319 , w_7322 );
not (  , w_7323 );
and ( w_7322 , w_7323 , \2318_b0 );
or ( \2320_b1 , \2317_b1 , w_7325 );
not ( w_7325 , w_7326 );
and ( \2320_b0 , \2317_b0 , w_7327 );
and ( w_7326 ,  , w_7327 );
buf ( w_7325 , \2319_b1 );
not ( w_7325 , w_7328 );
not (  , w_7329 );
and ( w_7328 , w_7329 , \2319_b0 );
or ( \2321_b1 , \b[0]_b1 , w_7330 );
or ( \2321_b0 , \b[0]_b0 , \c[10]_b0 );
not ( \c[10]_b0 , w_7331 );
and ( w_7331 , w_7330 , \c[10]_b1 );
or ( \2322_b1 , \2321_b1 , w_7333 );
not ( w_7333 , w_7334 );
and ( \2322_b0 , \2321_b0 , w_7335 );
and ( w_7334 ,  , w_7335 );
buf ( w_7333 , \c[9]_b1 );
not ( w_7333 , w_7336 );
not (  , w_7337 );
and ( w_7336 , w_7337 , \c[9]_b0 );
or ( \2323_b1 , \b[0]_b1 , w_7339 );
not ( w_7339 , w_7340 );
and ( \2323_b0 , \b[0]_b0 , w_7341 );
and ( w_7340 ,  , w_7341 );
buf ( w_7339 , \c[10]_b1 );
not ( w_7339 , w_7342 );
not (  , w_7343 );
and ( w_7342 , w_7343 , \c[10]_b0 );
buf ( \2325_b1 , \2324_b1 );
not ( \2325_b1 , w_7344 );
not ( \2325_b0 , w_7345 );
and ( w_7344 , w_7345 , \2324_b0 );
or ( \2326_b1 , \2320_b1 , \2325_b1 );
not ( \2325_b1 , w_7346 );
and ( \2326_b0 , \2320_b0 , w_7347 );
and ( w_7346 , w_7347 , \2325_b0 );
buf ( \2327_b1 , \2326_b1 );
not ( \2327_b1 , w_7348 );
not ( \2327_b0 , w_7349 );
and ( w_7348 , w_7349 , \2326_b0 );
or ( \2328_b1 , \2313_b1 , w_7350 );
or ( \2328_b0 , \2313_b0 , \2327_b0 );
not ( \2327_b0 , w_7351 );
and ( w_7351 , w_7350 , \2327_b1 );
or ( \2329_b1 , \2312_b1 , w_7352 );
or ( \2329_b0 , \2312_b0 , \2326_b0 );
not ( \2326_b0 , w_7353 );
and ( w_7353 , w_7352 , \2326_b1 );
or ( \2330_b1 , \b[10]_b1 , \c[1]_b1 );
xor ( \2330_b0 , \b[10]_b0 , w_7354 );
not ( w_7354 , w_7355 );
and ( w_7355 , \c[1]_b1 , \c[1]_b0 );
buf ( \2331_b1 , \2330_b1 );
not ( \2331_b1 , w_7356 );
not ( \2331_b0 , w_7357 );
and ( w_7356 , w_7357 , \2330_b0 );
buf ( \2332_b1 , \679_b1 );
not ( \2332_b1 , w_7358 );
not ( \2332_b0 , w_7359 );
and ( w_7358 , w_7359 , \679_b0 );
or ( \2333_b1 , \2331_b1 , w_7360 );
or ( \2333_b0 , \2331_b0 , \2332_b0 );
not ( \2332_b0 , w_7361 );
and ( w_7361 , w_7360 , \2332_b1 );
or ( \2334_b1 , \b[11]_b1 , \c[1]_b1 );
xor ( \2334_b0 , \b[11]_b0 , w_7362 );
not ( w_7362 , w_7363 );
and ( w_7363 , \c[1]_b1 , \c[1]_b0 );
or ( \2335_b1 , \2334_b1 , w_7365 );
not ( w_7365 , w_7366 );
and ( \2335_b0 , \2334_b0 , w_7367 );
and ( w_7366 ,  , w_7367 );
buf ( w_7365 , \c[0]_b1 );
not ( w_7365 , w_7368 );
not (  , w_7369 );
and ( w_7368 , w_7369 , \c[0]_b0 );
or ( \2336_b1 , \2333_b1 , w_7371 );
not ( w_7371 , w_7372 );
and ( \2336_b0 , \2333_b0 , w_7373 );
and ( w_7372 ,  , w_7373 );
buf ( w_7371 , \2335_b1 );
not ( w_7371 , w_7374 );
not (  , w_7375 );
and ( w_7374 , w_7375 , \2335_b0 );
buf ( \2337_b1 , \2336_b1 );
not ( \2337_b1 , w_7376 );
not ( \2337_b0 , w_7377 );
and ( w_7376 , w_7377 , \2336_b0 );
or ( \2338_b1 , \b[2]_b1 , \c[9]_b1 );
xor ( \2338_b0 , \b[2]_b0 , w_7378 );
not ( w_7378 , w_7379 );
and ( w_7379 , \c[9]_b1 , \c[9]_b0 );
buf ( \2339_b1 , \2338_b1 );
not ( \2339_b1 , w_7380 );
not ( \2339_b0 , w_7381 );
and ( w_7380 , w_7381 , \2338_b0 );
buf ( \2340_b1 , \2281_b1 );
not ( \2340_b1 , w_7382 );
not ( \2340_b0 , w_7383 );
and ( w_7382 , w_7383 , \2281_b0 );
or ( \2341_b1 , \2339_b1 , w_7384 );
or ( \2341_b0 , \2339_b0 , \2340_b0 );
not ( \2340_b0 , w_7385 );
and ( w_7385 , w_7384 , \2340_b1 );
or ( \2342_b1 , \b[3]_b1 , \c[9]_b1 );
xor ( \2342_b0 , \b[3]_b0 , w_7386 );
not ( w_7386 , w_7387 );
and ( w_7387 , \c[9]_b1 , \c[9]_b0 );
or ( \2343_b1 , \2284_b1 , w_7389 );
not ( w_7389 , w_7390 );
and ( \2343_b0 , \2284_b0 , w_7391 );
and ( w_7390 ,  , w_7391 );
buf ( w_7389 , \2342_b1 );
not ( w_7389 , w_7392 );
not (  , w_7393 );
and ( w_7392 , w_7393 , \2342_b0 );
or ( \2344_b1 , \2341_b1 , w_7395 );
not ( w_7395 , w_7396 );
and ( \2344_b0 , \2341_b0 , w_7397 );
and ( w_7396 ,  , w_7397 );
buf ( w_7395 , \2343_b1 );
not ( w_7395 , w_7398 );
not (  , w_7399 );
and ( w_7398 , w_7399 , \2343_b0 );
buf ( \2345_b1 , \2344_b1 );
not ( \2345_b1 , w_7400 );
not ( \2345_b0 , w_7401 );
and ( w_7400 , w_7401 , \2344_b0 );
or ( \2346_b1 , \2337_b1 , w_7402 );
or ( \2346_b0 , \2337_b0 , \2345_b0 );
not ( \2345_b0 , w_7403 );
and ( w_7403 , w_7402 , \2345_b1 );
or ( \2347_b1 , \2344_b1 , w_7404 );
or ( \2347_b0 , \2344_b0 , \2336_b0 );
not ( \2336_b0 , w_7405 );
and ( w_7405 , w_7404 , \2336_b1 );
or ( \2348_b1 , \b[4]_b1 , \c[7]_b1 );
xor ( \2348_b0 , \b[4]_b0 , w_7406 );
not ( w_7406 , w_7407 );
and ( w_7407 , \c[7]_b1 , \c[7]_b0 );
buf ( \2349_b1 , \2348_b1 );
not ( \2349_b1 , w_7408 );
not ( \2349_b0 , w_7409 );
and ( w_7408 , w_7409 , \2348_b0 );
buf ( \2350_b1 , \2292_b1 );
not ( \2350_b1 , w_7410 );
not ( \2350_b0 , w_7411 );
and ( w_7410 , w_7411 , \2292_b0 );
or ( \2351_b1 , \2349_b1 , w_7412 );
or ( \2351_b0 , \2349_b0 , \2350_b0 );
not ( \2350_b0 , w_7413 );
and ( w_7413 , w_7412 , \2350_b1 );
or ( \2352_b1 , \b[5]_b1 , \c[7]_b1 );
xor ( \2352_b0 , \b[5]_b0 , w_7414 );
not ( w_7414 , w_7415 );
and ( w_7415 , \c[7]_b1 , \c[7]_b0 );
or ( \2353_b1 , \714_b1 , w_7417 );
not ( w_7417 , w_7418 );
and ( \2353_b0 , \714_b0 , w_7419 );
and ( w_7418 ,  , w_7419 );
buf ( w_7417 , \2352_b1 );
not ( w_7417 , w_7420 );
not (  , w_7421 );
and ( w_7420 , w_7421 , \2352_b0 );
or ( \2354_b1 , \2351_b1 , w_7423 );
not ( w_7423 , w_7424 );
and ( \2354_b0 , \2351_b0 , w_7425 );
and ( w_7424 ,  , w_7425 );
buf ( w_7423 , \2353_b1 );
not ( w_7423 , w_7426 );
not (  , w_7427 );
and ( w_7426 , w_7427 , \2353_b0 );
or ( \2355_b1 , \2347_b1 , w_7429 );
not ( w_7429 , w_7430 );
and ( \2355_b0 , \2347_b0 , w_7431 );
and ( w_7430 ,  , w_7431 );
buf ( w_7429 , \2354_b1 );
not ( w_7429 , w_7432 );
not (  , w_7433 );
and ( w_7432 , w_7433 , \2354_b0 );
or ( \2356_b1 , \2346_b1 , w_7435 );
not ( w_7435 , w_7436 );
and ( \2356_b0 , \2346_b0 , w_7437 );
and ( w_7436 ,  , w_7437 );
buf ( w_7435 , \2355_b1 );
not ( w_7435 , w_7438 );
not (  , w_7439 );
and ( w_7438 , w_7439 , \2355_b0 );
or ( \2357_b1 , \2329_b1 , w_7441 );
not ( w_7441 , w_7442 );
and ( \2357_b0 , \2329_b0 , w_7443 );
and ( w_7442 ,  , w_7443 );
buf ( w_7441 , \2356_b1 );
not ( w_7441 , w_7444 );
not (  , w_7445 );
and ( w_7444 , w_7445 , \2356_b0 );
or ( \2358_b1 , \2328_b1 , w_7447 );
not ( w_7447 , w_7448 );
and ( \2358_b0 , \2328_b0 , w_7449 );
and ( w_7448 ,  , w_7449 );
buf ( w_7447 , \2357_b1 );
not ( w_7447 , w_7450 );
not (  , w_7451 );
and ( w_7450 , w_7451 , \2357_b0 );
or ( \2359_b1 , \2306_b1 , w_7453 );
not ( w_7453 , w_7454 );
and ( \2359_b0 , \2306_b0 , w_7455 );
and ( w_7454 ,  , w_7455 );
buf ( w_7453 , \2358_b1 );
not ( w_7453 , w_7456 );
not (  , w_7457 );
and ( w_7456 , w_7457 , \2358_b0 );
buf ( \2360_b1 , \2304_b1 );
not ( \2360_b1 , w_7458 );
not ( \2360_b0 , w_7459 );
and ( w_7458 , w_7459 , \2304_b0 );
buf ( \2361_b1 , \2275_b1 );
not ( \2361_b1 , w_7460 );
not ( \2361_b0 , w_7461 );
and ( w_7460 , w_7461 , \2275_b0 );
or ( \2362_b1 , \2360_b1 , w_7463 );
not ( w_7463 , w_7464 );
and ( \2362_b0 , \2360_b0 , w_7465 );
and ( w_7464 ,  , w_7465 );
buf ( w_7463 , \2361_b1 );
not ( w_7463 , w_7466 );
not (  , w_7467 );
and ( w_7466 , w_7467 , \2361_b0 );
or ( \2363_b1 , \2359_b1 , w_7469 );
not ( w_7469 , w_7470 );
and ( \2363_b0 , \2359_b0 , w_7471 );
and ( w_7470 ,  , w_7471 );
buf ( w_7469 , \2362_b1 );
not ( w_7469 , w_7472 );
not (  , w_7473 );
and ( w_7472 , w_7473 , \2362_b0 );
or ( \2364_b1 , \c[14]_b1 , \c[13]_b1 );
xor ( \2364_b0 , \c[14]_b0 , w_7474 );
not ( w_7474 , w_7475 );
and ( w_7475 , \c[13]_b1 , \c[13]_b0 );
or ( \2365_b1 , \2364_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_7476 );
and ( \2365_b0 , \2364_b0 , w_7477 );
and ( w_7476 , w_7477 , \b[0]_b0 );
or ( \2366_b1 , \b[13]_b1 , \c[1]_b1 );
xor ( \2366_b0 , \b[13]_b0 , w_7478 );
not ( w_7478 , w_7479 );
and ( w_7479 , \c[1]_b1 , \c[1]_b0 );
buf ( \2367_b1 , \2366_b1 );
not ( \2367_b1 , w_7480 );
not ( \2367_b0 , w_7481 );
and ( w_7480 , w_7481 , \2366_b0 );
buf ( \2368_b1 , \679_b1 );
not ( \2368_b1 , w_7482 );
not ( \2368_b0 , w_7483 );
and ( w_7482 , w_7483 , \679_b0 );
or ( \2369_b1 , \2367_b1 , w_7484 );
or ( \2369_b0 , \2367_b0 , \2368_b0 );
not ( \2368_b0 , w_7485 );
and ( w_7485 , w_7484 , \2368_b1 );
or ( \2370_b1 , \b[14]_b1 , \c[1]_b1 );
xor ( \2370_b0 , \b[14]_b0 , w_7486 );
not ( w_7486 , w_7487 );
and ( w_7487 , \c[1]_b1 , \c[1]_b0 );
or ( \2371_b1 , \2370_b1 , w_7489 );
not ( w_7489 , w_7490 );
and ( \2371_b0 , \2370_b0 , w_7491 );
and ( w_7490 ,  , w_7491 );
buf ( w_7489 , \c[0]_b1 );
not ( w_7489 , w_7492 );
not (  , w_7493 );
and ( w_7492 , w_7493 , \c[0]_b0 );
or ( \2372_b1 , \2369_b1 , w_7495 );
not ( w_7495 , w_7496 );
and ( \2372_b0 , \2369_b0 , w_7497 );
and ( w_7496 ,  , w_7497 );
buf ( w_7495 , \2371_b1 );
not ( w_7495 , w_7498 );
not (  , w_7499 );
and ( w_7498 , w_7499 , \2371_b0 );
or ( \2373_b1 , \2365_b1 , \2372_b1 );
xor ( \2373_b0 , \2365_b0 , w_7500 );
not ( w_7500 , w_7501 );
and ( w_7501 , \2372_b1 , \2372_b0 );
buf ( \2374_b1 , \2301_b1 );
not ( \2374_b1 , w_7502 );
not ( \2374_b0 , w_7503 );
and ( w_7502 , w_7503 , \2301_b0 );
buf ( \2375_b1 , \746_b1 );
not ( \2375_b1 , w_7504 );
not ( \2375_b0 , w_7505 );
and ( w_7504 , w_7505 , \746_b0 );
or ( \2376_b1 , \2374_b1 , w_7506 );
or ( \2376_b0 , \2374_b0 , \2375_b0 );
not ( \2375_b0 , w_7507 );
and ( w_7507 , w_7506 , \2375_b1 );
or ( \2377_b1 , \b[12]_b1 , \c[3]_b1 );
xor ( \2377_b0 , \b[12]_b0 , w_7508 );
not ( w_7508 , w_7509 );
and ( w_7509 , \c[3]_b1 , \c[3]_b0 );
or ( \2378_b1 , \702_b1 , w_7511 );
not ( w_7511 , w_7512 );
and ( \2378_b0 , \702_b0 , w_7513 );
and ( w_7512 ,  , w_7513 );
buf ( w_7511 , \2377_b1 );
not ( w_7511 , w_7514 );
not (  , w_7515 );
and ( w_7514 , w_7515 , \2377_b0 );
or ( \2379_b1 , \2376_b1 , w_7517 );
not ( w_7517 , w_7518 );
and ( \2379_b0 , \2376_b0 , w_7519 );
and ( w_7518 ,  , w_7519 );
buf ( w_7517 , \2378_b1 );
not ( w_7517 , w_7520 );
not (  , w_7521 );
and ( w_7520 , w_7521 , \2378_b0 );
or ( \2380_b1 , \2373_b1 , \2379_b1 );
xor ( \2380_b0 , \2373_b0 , w_7522 );
not ( w_7522 , w_7523 );
and ( w_7523 , \2379_b1 , \2379_b0 );
buf ( \2381_b1 , \2287_b1 );
not ( \2381_b1 , w_7524 );
not ( \2381_b0 , w_7525 );
and ( w_7524 , w_7525 , \2287_b0 );
buf ( \2382_b1 , \2303_b1 );
not ( \2382_b1 , w_7526 );
not ( \2382_b0 , w_7527 );
and ( w_7526 , w_7527 , \2303_b0 );
or ( \2383_b1 , \2381_b1 , w_7528 );
or ( \2383_b0 , \2381_b0 , \2382_b0 );
not ( \2382_b0 , w_7529 );
and ( w_7529 , w_7528 , \2382_b1 );
or ( \2384_b1 , \2303_b1 , w_7530 );
or ( \2384_b0 , \2303_b0 , \2287_b0 );
not ( \2287_b0 , w_7531 );
and ( w_7531 , w_7530 , \2287_b1 );
or ( \2385_b1 , \2384_b1 , w_7533 );
not ( w_7533 , w_7534 );
and ( \2385_b0 , \2384_b0 , w_7535 );
and ( w_7534 ,  , w_7535 );
buf ( w_7533 , \2295_b1 );
not ( w_7533 , w_7536 );
not (  , w_7537 );
and ( w_7536 , w_7537 , \2295_b0 );
or ( \2386_b1 , \2383_b1 , w_7539 );
not ( w_7539 , w_7540 );
and ( \2386_b0 , \2383_b0 , w_7541 );
and ( w_7540 ,  , w_7541 );
buf ( w_7539 , \2385_b1 );
not ( w_7539 , w_7542 );
not (  , w_7543 );
and ( w_7542 , w_7543 , \2385_b0 );
or ( \2387_b1 , \2380_b1 , \2386_b1 );
xor ( \2387_b0 , \2380_b0 , w_7544 );
not ( w_7544 , w_7545 );
and ( w_7545 , \2386_b1 , \2386_b0 );
buf ( \2388_b1 , \2258_b1 );
not ( \2388_b1 , w_7546 );
not ( \2388_b0 , w_7547 );
and ( w_7546 , w_7547 , \2258_b0 );
buf ( \2389_b1 , \2271_b1 );
not ( \2389_b1 , w_7548 );
not ( \2389_b0 , w_7549 );
and ( w_7548 , w_7549 , \2271_b0 );
or ( \2390_b1 , \2388_b1 , w_7550 );
or ( \2390_b0 , \2388_b0 , \2389_b0 );
not ( \2389_b0 , w_7551 );
and ( w_7551 , w_7550 , \2389_b1 );
or ( \2391_b1 , \2390_b1 , w_7553 );
not ( w_7553 , w_7554 );
and ( \2391_b0 , \2390_b0 , w_7555 );
and ( w_7554 ,  , w_7555 );
buf ( w_7553 , \2243_b1 );
not ( w_7553 , w_7556 );
not (  , w_7557 );
and ( w_7556 , w_7557 , \2243_b0 );
or ( \2392_b1 , \2270_b1 , w_7559 );
not ( w_7559 , w_7560 );
and ( \2392_b0 , \2270_b0 , w_7561 );
and ( w_7560 ,  , w_7561 );
buf ( w_7559 , \2257_b1 );
not ( w_7559 , w_7562 );
not (  , w_7563 );
and ( w_7562 , w_7563 , \2257_b0 );
or ( \2393_b1 , \2391_b1 , w_7565 );
not ( w_7565 , w_7566 );
and ( \2393_b0 , \2391_b0 , w_7567 );
and ( w_7566 ,  , w_7567 );
buf ( w_7565 , \2392_b1 );
not ( w_7565 , w_7568 );
not (  , w_7569 );
and ( w_7568 , w_7569 , \2392_b0 );
or ( \2394_b1 , \2387_b1 , \2393_b1 );
xor ( \2394_b0 , \2387_b0 , w_7570 );
not ( w_7570 , w_7571 );
and ( w_7571 , \2393_b1 , \2393_b0 );
or ( \2395_b1 , \2363_b1 , \2394_b1 );
xor ( \2395_b0 , \2363_b0 , w_7572 );
not ( w_7572 , w_7573 );
and ( w_7573 , \2394_b1 , \2394_b0 );
buf ( \2396_b1 , \2288_b1 );
not ( \2396_b1 , w_7574 );
not ( \2396_b0 , w_7575 );
and ( w_7574 , w_7575 , \2288_b0 );
buf ( \2397_b1 , \2292_b1 );
not ( \2397_b1 , w_7576 );
not ( \2397_b0 , w_7577 );
and ( w_7576 , w_7577 , \2292_b0 );
or ( \2398_b1 , \2396_b1 , w_7578 );
or ( \2398_b0 , \2396_b0 , \2397_b0 );
not ( \2397_b0 , w_7579 );
and ( w_7579 , w_7578 , \2397_b1 );
or ( \2399_b1 , \b[8]_b1 , \c[7]_b1 );
xor ( \2399_b0 , \b[8]_b0 , w_7580 );
not ( w_7580 , w_7581 );
and ( w_7581 , \c[7]_b1 , \c[7]_b0 );
or ( \2400_b1 , \714_b1 , w_7583 );
not ( w_7583 , w_7584 );
and ( \2400_b0 , \714_b0 , w_7585 );
and ( w_7584 ,  , w_7585 );
buf ( w_7583 , \2399_b1 );
not ( w_7583 , w_7586 );
not (  , w_7587 );
and ( w_7586 , w_7587 , \2399_b0 );
or ( \2401_b1 , \2398_b1 , w_7589 );
not ( w_7589 , w_7590 );
and ( \2401_b0 , \2398_b0 , w_7591 );
and ( w_7590 ,  , w_7591 );
buf ( w_7589 , \2400_b1 );
not ( w_7589 , w_7592 );
not (  , w_7593 );
and ( w_7592 , w_7593 , \2400_b0 );
buf ( \2402_b1 , \2285_b1 );
not ( \2402_b1 , w_7594 );
not ( \2402_b0 , w_7595 );
and ( w_7594 , w_7595 , \2285_b0 );
buf ( \2403_b1 , \2281_b1 );
not ( \2403_b1 , w_7596 );
not ( \2403_b0 , w_7597 );
and ( w_7596 , w_7597 , \2281_b0 );
or ( \2404_b1 , \2402_b1 , w_7598 );
or ( \2404_b0 , \2402_b0 , \2403_b0 );
not ( \2403_b0 , w_7599 );
and ( w_7599 , w_7598 , \2403_b1 );
or ( \2405_b1 , \b[6]_b1 , \c[9]_b1 );
xor ( \2405_b0 , \b[6]_b0 , w_7600 );
not ( w_7600 , w_7601 );
and ( w_7601 , \c[9]_b1 , \c[9]_b0 );
or ( \2406_b1 , \2284_b1 , w_7603 );
not ( w_7603 , w_7604 );
and ( \2406_b0 , \2284_b0 , w_7605 );
and ( w_7604 ,  , w_7605 );
buf ( w_7603 , \2405_b1 );
not ( w_7603 , w_7606 );
not (  , w_7607 );
and ( w_7606 , w_7607 , \2405_b0 );
or ( \2407_b1 , \2404_b1 , w_7609 );
not ( w_7609 , w_7610 );
and ( \2407_b0 , \2404_b0 , w_7611 );
and ( w_7610 ,  , w_7611 );
buf ( w_7609 , \2406_b1 );
not ( w_7609 , w_7612 );
not (  , w_7613 );
and ( w_7612 , w_7613 , \2406_b0 );
or ( \2408_b1 , \2401_b1 , \2407_b1 );
xor ( \2408_b0 , \2401_b0 , w_7614 );
not ( w_7614 , w_7615 );
and ( w_7615 , \2407_b1 , \2407_b0 );
buf ( \2409_b1 , \2268_b1 );
not ( \2409_b1 , w_7616 );
not ( \2409_b0 , w_7617 );
and ( w_7616 , w_7617 , \2268_b0 );
buf ( \2410_b1 , \2265_b1 );
not ( \2410_b1 , w_7618 );
not ( \2410_b0 , w_7619 );
and ( w_7618 , w_7619 , \2265_b0 );
or ( \2411_b1 , \2409_b1 , w_7620 );
or ( \2411_b0 , \2409_b0 , \2410_b0 );
not ( \2410_b0 , w_7621 );
and ( w_7621 , w_7620 , \2410_b1 );
or ( \2412_b1 , \b[10]_b1 , \c[5]_b1 );
xor ( \2412_b0 , \b[10]_b0 , w_7622 );
not ( w_7622 , w_7623 );
and ( w_7623 , \c[5]_b1 , \c[5]_b0 );
or ( \2413_b1 , \739_b1 , w_7625 );
not ( w_7625 , w_7626 );
and ( \2413_b0 , \739_b0 , w_7627 );
and ( w_7626 ,  , w_7627 );
buf ( w_7625 , \2412_b1 );
not ( w_7625 , w_7628 );
not (  , w_7629 );
and ( w_7628 , w_7629 , \2412_b0 );
or ( \2414_b1 , \2411_b1 , w_7631 );
not ( w_7631 , w_7632 );
and ( \2414_b0 , \2411_b0 , w_7633 );
and ( w_7632 ,  , w_7633 );
buf ( w_7631 , \2413_b1 );
not ( w_7631 , w_7634 );
not (  , w_7635 );
and ( w_7634 , w_7635 , \2413_b0 );
or ( \2415_b1 , \2408_b1 , \2414_b1 );
xor ( \2415_b0 , \2408_b0 , w_7636 );
not ( w_7636 , w_7637 );
and ( w_7637 , \2414_b1 , \2414_b0 );
buf ( \2416_b1 , \2255_b1 );
not ( \2416_b1 , w_7638 );
not ( \2416_b0 , w_7639 );
and ( w_7638 , w_7639 , \2255_b0 );
buf ( \2417_b1 , \2252_b1 );
not ( \2417_b1 , w_7640 );
not ( \2417_b0 , w_7641 );
and ( w_7640 , w_7641 , \2252_b0 );
or ( \2418_b1 , \2416_b1 , w_7642 );
or ( \2418_b0 , \2416_b0 , \2417_b0 );
not ( \2417_b0 , w_7643 );
and ( w_7643 , w_7642 , \2417_b1 );
or ( \2419_b1 , \b[2]_b1 , \c[13]_b1 );
xor ( \2419_b0 , \b[2]_b0 , w_7644 );
not ( w_7644 , w_7645 );
and ( w_7645 , \c[13]_b1 , \c[13]_b0 );
or ( \2420_b1 , \2246_b1 , w_7647 );
not ( w_7647 , w_7648 );
and ( \2420_b0 , \2246_b0 , w_7649 );
and ( w_7648 ,  , w_7649 );
buf ( w_7647 , \2419_b1 );
not ( w_7647 , w_7650 );
not (  , w_7651 );
and ( w_7650 , w_7651 , \2419_b0 );
or ( \2421_b1 , \2418_b1 , w_7653 );
not ( w_7653 , w_7654 );
and ( \2421_b0 , \2418_b0 , w_7655 );
and ( w_7654 ,  , w_7655 );
buf ( w_7653 , \2420_b1 );
not ( w_7653 , w_7656 );
not (  , w_7657 );
and ( w_7656 , w_7657 , \2420_b0 );
buf ( \2422_b1 , \2241_b1 );
not ( \2422_b1 , w_7658 );
not ( \2422_b0 , w_7659 );
and ( w_7658 , w_7659 , \2241_b0 );
buf ( \2423_b1 , \2238_b1 );
not ( \2423_b1 , w_7660 );
not ( \2423_b0 , w_7661 );
and ( w_7660 , w_7661 , \2238_b0 );
or ( \2424_b1 , \2422_b1 , w_7662 );
or ( \2424_b0 , \2422_b0 , \2423_b0 );
not ( \2423_b0 , w_7663 );
and ( w_7663 , w_7662 , \2423_b1 );
or ( \2425_b1 , \b[4]_b1 , \c[11]_b1 );
xor ( \2425_b0 , \b[4]_b0 , w_7664 );
not ( w_7664 , w_7665 );
and ( w_7665 , \c[11]_b1 , \c[11]_b0 );
or ( \2426_b1 , \2236_b1 , w_7667 );
not ( w_7667 , w_7668 );
and ( \2426_b0 , \2236_b0 , w_7669 );
and ( w_7668 ,  , w_7669 );
buf ( w_7667 , \2425_b1 );
not ( w_7667 , w_7670 );
not (  , w_7671 );
and ( w_7670 , w_7671 , \2425_b0 );
or ( \2427_b1 , \2424_b1 , w_7673 );
not ( w_7673 , w_7674 );
and ( \2427_b0 , \2424_b0 , w_7675 );
and ( w_7674 ,  , w_7675 );
buf ( w_7673 , \2426_b1 );
not ( w_7673 , w_7676 );
not (  , w_7677 );
and ( w_7676 , w_7677 , \2426_b0 );
or ( \2428_b1 , \2421_b1 , \2427_b1 );
xor ( \2428_b0 , \2421_b0 , w_7678 );
not ( w_7678 , w_7679 );
and ( w_7679 , \2427_b1 , \2427_b0 );
or ( \2429_b1 , \b[0]_b1 , w_7680 );
or ( \2429_b0 , \b[0]_b0 , \c[12]_b0 );
not ( \c[12]_b0 , w_7681 );
and ( w_7681 , w_7680 , \c[12]_b1 );
or ( \2430_b1 , \2429_b1 , w_7683 );
not ( w_7683 , w_7684 );
and ( \2430_b0 , \2429_b0 , w_7685 );
and ( w_7684 ,  , w_7685 );
buf ( w_7683 , \c[11]_b1 );
not ( w_7683 , w_7686 );
not (  , w_7687 );
and ( w_7686 , w_7687 , \c[11]_b0 );
or ( \2431_b1 , \b[0]_b1 , w_7689 );
not ( w_7689 , w_7690 );
and ( \2431_b0 , \b[0]_b0 , w_7691 );
and ( w_7690 ,  , w_7691 );
buf ( w_7689 , \c[12]_b1 );
not ( w_7689 , w_7692 );
not (  , w_7693 );
and ( w_7692 , w_7693 , \c[12]_b0 );
or ( \2433_b1 , \b[12]_b1 , \c[1]_b1 );
xor ( \2433_b0 , \b[12]_b0 , w_7694 );
not ( w_7694 , w_7695 );
and ( w_7695 , \c[1]_b1 , \c[1]_b0 );
buf ( \2434_b1 , \2433_b1 );
not ( \2434_b1 , w_7696 );
not ( \2434_b0 , w_7697 );
and ( w_7696 , w_7697 , \2433_b0 );
buf ( \2435_b1 , \679_b1 );
not ( \2435_b1 , w_7698 );
not ( \2435_b0 , w_7699 );
and ( w_7698 , w_7699 , \679_b0 );
or ( \2436_b1 , \2434_b1 , w_7700 );
or ( \2436_b0 , \2434_b0 , \2435_b0 );
not ( \2435_b0 , w_7701 );
and ( w_7701 , w_7700 , \2435_b1 );
or ( \2437_b1 , \2366_b1 , w_7703 );
not ( w_7703 , w_7704 );
and ( \2437_b0 , \2366_b0 , w_7705 );
and ( w_7704 ,  , w_7705 );
buf ( w_7703 , \c[0]_b1 );
not ( w_7703 , w_7706 );
not (  , w_7707 );
and ( w_7706 , w_7707 , \c[0]_b0 );
or ( \2438_b1 , \2436_b1 , w_7709 );
not ( w_7709 , w_7710 );
and ( \2438_b0 , \2436_b0 , w_7711 );
and ( w_7710 ,  , w_7711 );
buf ( w_7709 , \2437_b1 );
not ( w_7709 , w_7712 );
not (  , w_7713 );
and ( w_7712 , w_7713 , \2437_b0 );
or ( \2439_b1 , \2432_b1 , \2438_b1 );
not ( \2438_b1 , w_7714 );
and ( \2439_b0 , \2432_b0 , w_7715 );
and ( w_7714 , w_7715 , \2438_b0 );
or ( \2440_b1 , \2428_b1 , \2439_b1 );
xor ( \2440_b0 , \2428_b0 , w_7716 );
not ( w_7716 , w_7717 );
and ( w_7717 , \2439_b1 , \2439_b0 );
or ( \2441_b1 , \2415_b1 , \2440_b1 );
xor ( \2441_b0 , \2415_b0 , w_7718 );
not ( w_7718 , w_7719 );
and ( w_7719 , \2440_b1 , \2440_b0 );
buf ( \2442_b1 , \2334_b1 );
not ( \2442_b1 , w_7720 );
not ( \2442_b0 , w_7721 );
and ( w_7720 , w_7721 , \2334_b0 );
buf ( \2443_b1 , \679_b1 );
not ( \2443_b1 , w_7722 );
not ( \2443_b0 , w_7723 );
and ( w_7722 , w_7723 , \679_b0 );
or ( \2444_b1 , \2442_b1 , w_7724 );
or ( \2444_b0 , \2442_b0 , \2443_b0 );
not ( \2443_b0 , w_7725 );
and ( w_7725 , w_7724 , \2443_b1 );
or ( \2445_b1 , \2433_b1 , w_7727 );
not ( w_7727 , w_7728 );
and ( \2445_b0 , \2433_b0 , w_7729 );
and ( w_7728 ,  , w_7729 );
buf ( w_7727 , \c[0]_b1 );
not ( w_7727 , w_7730 );
not (  , w_7731 );
and ( w_7730 , w_7731 , \c[0]_b0 );
or ( \2446_b1 , \2444_b1 , w_7733 );
not ( w_7733 , w_7734 );
and ( \2446_b0 , \2444_b0 , w_7735 );
and ( w_7734 ,  , w_7735 );
buf ( w_7733 , \2445_b1 );
not ( w_7733 , w_7736 );
not (  , w_7737 );
and ( w_7736 , w_7737 , \2445_b0 );
buf ( \2447_b1 , \2342_b1 );
not ( \2447_b1 , w_7738 );
not ( \2447_b0 , w_7739 );
and ( w_7738 , w_7739 , \2342_b0 );
or ( \2448_b1 , \2279_b1 , w_7741 );
not ( w_7741 , w_7742 );
and ( \2448_b0 , \2279_b0 , w_7743 );
and ( w_7742 ,  , w_7743 );
buf ( w_7741 , \2280_b1 );
not ( w_7741 , w_7744 );
not (  , w_7745 );
and ( w_7744 , w_7745 , \2280_b0 );
buf ( \2449_b1 , \2448_b1 );
not ( \2449_b1 , w_7746 );
not ( \2449_b0 , w_7747 );
and ( w_7746 , w_7747 , \2448_b0 );
or ( \2450_b1 , \2447_b1 , w_7748 );
or ( \2450_b0 , \2447_b0 , \2449_b0 );
not ( \2449_b0 , w_7749 );
and ( w_7749 , w_7748 , \2449_b1 );
or ( \2451_b1 , \2284_b1 , w_7751 );
not ( w_7751 , w_7752 );
and ( \2451_b0 , \2284_b0 , w_7753 );
and ( w_7752 ,  , w_7753 );
buf ( w_7751 , \2277_b1 );
not ( w_7751 , w_7754 );
not (  , w_7755 );
and ( w_7754 , w_7755 , \2277_b0 );
or ( \2452_b1 , \2450_b1 , w_7757 );
not ( w_7757 , w_7758 );
and ( \2452_b0 , \2450_b0 , w_7759 );
and ( w_7758 ,  , w_7759 );
buf ( w_7757 , \2451_b1 );
not ( w_7757 , w_7760 );
not (  , w_7761 );
and ( w_7760 , w_7761 , \2451_b0 );
or ( \2453_b1 , \2446_b1 , \2452_b1 );
xor ( \2453_b0 , \2446_b0 , w_7762 );
not ( w_7762 , w_7763 );
and ( w_7763 , \2452_b1 , \2452_b0 );
or ( \2454_b1 , \b[1]_b1 , \c[11]_b1 );
xor ( \2454_b0 , \b[1]_b0 , w_7764 );
not ( w_7764 , w_7765 );
and ( w_7765 , \c[11]_b1 , \c[11]_b0 );
buf ( \2455_b1 , \2454_b1 );
not ( \2455_b1 , w_7766 );
not ( \2455_b0 , w_7767 );
and ( w_7766 , w_7767 , \2454_b0 );
buf ( \2456_b1 , \2238_b1 );
not ( \2456_b1 , w_7768 );
not ( \2456_b0 , w_7769 );
and ( w_7768 , w_7769 , \2238_b0 );
or ( \2457_b1 , \2455_b1 , w_7770 );
or ( \2457_b0 , \2455_b0 , \2456_b0 );
not ( \2456_b0 , w_7771 );
and ( w_7771 , w_7770 , \2456_b1 );
or ( \2458_b1 , \2236_b1 , w_7773 );
not ( w_7773 , w_7774 );
and ( \2458_b0 , \2236_b0 , w_7775 );
and ( w_7774 ,  , w_7775 );
buf ( w_7773 , \2234_b1 );
not ( w_7773 , w_7776 );
not (  , w_7777 );
and ( w_7776 , w_7777 , \2234_b0 );
or ( \2459_b1 , \2457_b1 , w_7779 );
not ( w_7779 , w_7780 );
and ( \2459_b0 , \2457_b0 , w_7781 );
and ( w_7780 ,  , w_7781 );
buf ( w_7779 , \2458_b1 );
not ( w_7779 , w_7782 );
not (  , w_7783 );
and ( w_7782 , w_7783 , \2458_b0 );
or ( \2460_b1 , \2453_b1 , \2459_b1 );
not ( \2459_b1 , w_7784 );
and ( \2460_b0 , \2453_b0 , w_7785 );
and ( w_7784 , w_7785 , \2459_b0 );
or ( \2461_b1 , \2446_b1 , \2452_b1 );
not ( \2452_b1 , w_7786 );
and ( \2461_b0 , \2446_b0 , w_7787 );
and ( w_7786 , w_7787 , \2452_b0 );
or ( \2462_b1 , \2460_b1 , w_7788 );
or ( \2462_b0 , \2460_b0 , \2461_b0 );
not ( \2461_b0 , w_7789 );
and ( w_7789 , w_7788 , \2461_b1 );
or ( \2463_b1 , \2432_b1 , \2438_b1 );
xor ( \2463_b0 , \2432_b0 , w_7790 );
not ( w_7790 , w_7791 );
and ( w_7791 , \2438_b1 , \2438_b0 );
or ( \2464_b1 , \2462_b1 , w_7792 );
or ( \2464_b0 , \2462_b0 , \2463_b0 );
not ( \2463_b0 , w_7793 );
and ( w_7793 , w_7792 , \2463_b1 );
or ( \2465_b1 , \2246_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_7794 );
and ( \2465_b0 , \2246_b0 , w_7795 );
and ( w_7794 , w_7795 , \b[0]_b0 );
buf ( \2466_b1 , \2352_b1 );
not ( \2466_b1 , w_7796 );
not ( \2466_b0 , w_7797 );
and ( w_7796 , w_7797 , \2352_b0 );
buf ( \2467_b1 , \726_b1 );
not ( \2467_b1 , w_7798 );
not ( \2467_b0 , w_7799 );
and ( w_7798 , w_7799 , \726_b0 );
or ( \2468_b1 , \2466_b1 , w_7800 );
or ( \2468_b0 , \2466_b0 , \2467_b0 );
not ( \2467_b0 , w_7801 );
and ( w_7801 , w_7800 , \2467_b1 );
or ( \2469_b1 , \714_b1 , w_7803 );
not ( w_7803 , w_7804 );
and ( \2469_b0 , \714_b0 , w_7805 );
and ( w_7804 ,  , w_7805 );
buf ( w_7803 , \2293_b1 );
not ( w_7803 , w_7806 );
not (  , w_7807 );
and ( w_7806 , w_7807 , \2293_b0 );
or ( \2470_b1 , \2468_b1 , w_7809 );
not ( w_7809 , w_7810 );
and ( \2470_b0 , \2468_b0 , w_7811 );
and ( w_7810 ,  , w_7811 );
buf ( w_7809 , \2469_b1 );
not ( w_7809 , w_7812 );
not (  , w_7813 );
and ( w_7812 , w_7813 , \2469_b0 );
or ( \2471_b1 , \2465_b1 , \2470_b1 );
xor ( \2471_b0 , \2465_b0 , w_7814 );
not ( w_7814 , w_7815 );
and ( w_7815 , \2470_b1 , \2470_b0 );
buf ( \2472_b1 , \2318_b1 );
not ( \2472_b1 , w_7816 );
not ( \2472_b0 , w_7817 );
and ( w_7816 , w_7817 , \2318_b0 );
buf ( \2473_b1 , \699_b1 );
not ( \2473_b1 , w_7818 );
not ( \2473_b0 , w_7819 );
and ( w_7818 , w_7819 , \699_b0 );
or ( \2474_b1 , \2472_b1 , w_7820 );
or ( \2474_b0 , \2472_b0 , \2473_b0 );
not ( \2473_b0 , w_7821 );
and ( w_7821 , w_7820 , \2473_b1 );
or ( \2475_b1 , \702_b1 , w_7823 );
not ( w_7823 , w_7824 );
and ( \2475_b0 , \702_b0 , w_7825 );
and ( w_7824 ,  , w_7825 );
buf ( w_7823 , \2297_b1 );
not ( w_7823 , w_7826 );
not (  , w_7827 );
and ( w_7826 , w_7827 , \2297_b0 );
or ( \2476_b1 , \2474_b1 , w_7829 );
not ( w_7829 , w_7830 );
and ( \2476_b0 , \2474_b0 , w_7831 );
and ( w_7830 ,  , w_7831 );
buf ( w_7829 , \2475_b1 );
not ( w_7829 , w_7832 );
not (  , w_7833 );
and ( w_7832 , w_7833 , \2475_b0 );
or ( \2477_b1 , \2471_b1 , \2476_b1 );
not ( \2476_b1 , w_7834 );
and ( \2477_b0 , \2471_b0 , w_7835 );
and ( w_7834 , w_7835 , \2476_b0 );
or ( \2478_b1 , \2465_b1 , \2470_b1 );
not ( \2470_b1 , w_7836 );
and ( \2478_b0 , \2465_b0 , w_7837 );
and ( w_7836 , w_7837 , \2470_b0 );
or ( \2479_b1 , \2477_b1 , w_7838 );
or ( \2479_b0 , \2477_b0 , \2478_b0 );
not ( \2478_b0 , w_7839 );
and ( w_7839 , w_7838 , \2478_b1 );
or ( \2480_b1 , \2464_b1 , w_7841 );
not ( w_7841 , w_7842 );
and ( \2480_b0 , \2464_b0 , w_7843 );
and ( w_7842 ,  , w_7843 );
buf ( w_7841 , \2479_b1 );
not ( w_7841 , w_7844 );
not (  , w_7845 );
and ( w_7844 , w_7845 , \2479_b0 );
or ( \2481_b1 , \2462_b1 , w_7847 );
not ( w_7847 , w_7848 );
and ( \2481_b0 , \2462_b0 , w_7849 );
and ( w_7848 ,  , w_7849 );
buf ( w_7847 , \2463_b1 );
not ( w_7847 , w_7850 );
not (  , w_7851 );
and ( w_7850 , w_7851 , \2463_b0 );
or ( \2482_b1 , \2480_b1 , w_7853 );
not ( w_7853 , w_7854 );
and ( \2482_b0 , \2480_b0 , w_7855 );
and ( w_7854 ,  , w_7855 );
buf ( w_7853 , \2481_b1 );
not ( w_7853 , w_7856 );
not (  , w_7857 );
and ( w_7856 , w_7857 , \2481_b0 );
or ( \2483_b1 , \2441_b1 , \2482_b1 );
xor ( \2483_b0 , \2441_b0 , w_7858 );
not ( w_7858 , w_7859 );
and ( w_7859 , \2482_b1 , \2482_b0 );
or ( \2484_b1 , \2395_b1 , \2483_b1 );
not ( \2483_b1 , w_7860 );
and ( \2484_b0 , \2395_b0 , w_7861 );
and ( w_7860 , w_7861 , \2483_b0 );
or ( \2485_b1 , \2363_b1 , \2394_b1 );
not ( \2394_b1 , w_7862 );
and ( \2485_b0 , \2363_b0 , w_7863 );
and ( w_7862 , w_7863 , \2394_b0 );
or ( \2486_b1 , \2484_b1 , w_7864 );
or ( \2486_b0 , \2484_b0 , \2485_b0 );
not ( \2485_b0 , w_7865 );
and ( w_7865 , w_7864 , \2485_b1 );
or ( \2487_b1 , \2415_b1 , \2440_b1 );
xor ( \2487_b0 , \2415_b0 , w_7866 );
not ( w_7866 , w_7867 );
and ( w_7867 , \2440_b1 , \2440_b0 );
or ( \2488_b1 , \2487_b1 , \2482_b1 );
not ( \2482_b1 , w_7868 );
and ( \2488_b0 , \2487_b0 , w_7869 );
and ( w_7868 , w_7869 , \2482_b0 );
or ( \2489_b1 , \2415_b1 , \2440_b1 );
not ( \2440_b1 , w_7870 );
and ( \2489_b0 , \2415_b0 , w_7871 );
and ( w_7870 , w_7871 , \2440_b0 );
or ( \2490_b1 , \2488_b1 , w_7872 );
or ( \2490_b0 , \2488_b0 , \2489_b0 );
not ( \2489_b0 , w_7873 );
and ( w_7873 , w_7872 , \2489_b1 );
buf ( \2491_b1 , \2490_b1 );
not ( \2491_b1 , w_7874 );
not ( \2491_b0 , w_7875 );
and ( w_7874 , w_7875 , \2490_b0 );
or ( \2492_b1 , \2380_b1 , \2386_b1 );
xor ( \2492_b0 , \2380_b0 , w_7876 );
not ( w_7876 , w_7877 );
and ( w_7877 , \2386_b1 , \2386_b0 );
or ( \2493_b1 , \2492_b1 , \2393_b1 );
not ( \2393_b1 , w_7878 );
and ( \2493_b0 , \2492_b0 , w_7879 );
and ( w_7878 , w_7879 , \2393_b0 );
or ( \2494_b1 , \2380_b1 , \2386_b1 );
not ( \2386_b1 , w_7880 );
and ( \2494_b0 , \2380_b0 , w_7881 );
and ( w_7880 , w_7881 , \2386_b0 );
or ( \2495_b1 , \2493_b1 , w_7882 );
or ( \2495_b0 , \2493_b0 , \2494_b0 );
not ( \2494_b0 , w_7883 );
and ( w_7883 , w_7882 , \2494_b1 );
buf ( \2496_b1 , \2495_b1 );
not ( \2496_b1 , w_7884 );
not ( \2496_b0 , w_7885 );
and ( w_7884 , w_7885 , \2495_b0 );
buf ( \2497_b1 , \2496_b1 );
not ( \2497_b1 , w_7886 );
not ( \2497_b0 , w_7887 );
and ( w_7886 , w_7887 , \2496_b0 );
or ( \2498_b1 , \2491_b1 , \2497_b1 );
not ( \2497_b1 , w_7888 );
and ( \2498_b0 , \2491_b0 , w_7889 );
and ( w_7888 , w_7889 , \2497_b0 );
or ( \2499_b1 , \2490_b1 , \2496_b1 );
not ( \2496_b1 , w_7890 );
and ( \2499_b0 , \2490_b0 , w_7891 );
and ( w_7890 , w_7891 , \2496_b0 );
or ( \2500_b1 , \2498_b1 , w_7893 );
not ( w_7893 , w_7894 );
and ( \2500_b0 , \2498_b0 , w_7895 );
and ( w_7894 ,  , w_7895 );
buf ( w_7893 , \2499_b1 );
not ( w_7893 , w_7896 );
not (  , w_7897 );
and ( w_7896 , w_7897 , \2499_b0 );
buf ( \2501_b1 , \2377_b1 );
not ( \2501_b1 , w_7898 );
not ( \2501_b0 , w_7899 );
and ( w_7898 , w_7899 , \2377_b0 );
buf ( \2502_b1 , \746_b1 );
not ( \2502_b1 , w_7900 );
not ( \2502_b0 , w_7901 );
and ( w_7900 , w_7901 , \746_b0 );
or ( \2503_b1 , \2501_b1 , w_7902 );
or ( \2503_b0 , \2501_b0 , \2502_b0 );
not ( \2502_b0 , w_7903 );
and ( w_7903 , w_7902 , \2502_b1 );
or ( \2504_b1 , \b[13]_b1 , \c[3]_b1 );
xor ( \2504_b0 , \b[13]_b0 , w_7904 );
not ( w_7904 , w_7905 );
and ( w_7905 , \c[3]_b1 , \c[3]_b0 );
or ( \2505_b1 , \702_b1 , w_7907 );
not ( w_7907 , w_7908 );
and ( \2505_b0 , \702_b0 , w_7909 );
and ( w_7908 ,  , w_7909 );
buf ( w_7907 , \2504_b1 );
not ( w_7907 , w_7910 );
not (  , w_7911 );
and ( w_7910 , w_7911 , \2504_b0 );
or ( \2506_b1 , \2503_b1 , w_7913 );
not ( w_7913 , w_7914 );
and ( \2506_b0 , \2503_b0 , w_7915 );
and ( w_7914 ,  , w_7915 );
buf ( w_7913 , \2505_b1 );
not ( w_7913 , w_7916 );
not (  , w_7917 );
and ( w_7916 , w_7917 , \2505_b0 );
buf ( \2507_b1 , \2412_b1 );
not ( \2507_b1 , w_7918 );
not ( \2507_b0 , w_7919 );
and ( w_7918 , w_7919 , \2412_b0 );
buf ( \2508_b1 , \2265_b1 );
not ( \2508_b1 , w_7920 );
not ( \2508_b0 , w_7921 );
and ( w_7920 , w_7921 , \2265_b0 );
or ( \2509_b1 , \2507_b1 , w_7922 );
or ( \2509_b0 , \2507_b0 , \2508_b0 );
not ( \2508_b0 , w_7923 );
and ( w_7923 , w_7922 , \2508_b1 );
or ( \2510_b1 , \b[11]_b1 , \c[5]_b1 );
xor ( \2510_b0 , \b[11]_b0 , w_7924 );
not ( w_7924 , w_7925 );
and ( w_7925 , \c[5]_b1 , \c[5]_b0 );
or ( \2511_b1 , \739_b1 , w_7927 );
not ( w_7927 , w_7928 );
and ( \2511_b0 , \739_b0 , w_7929 );
and ( w_7928 ,  , w_7929 );
buf ( w_7927 , \2510_b1 );
not ( w_7927 , w_7930 );
not (  , w_7931 );
and ( w_7930 , w_7931 , \2510_b0 );
or ( \2512_b1 , \2509_b1 , w_7933 );
not ( w_7933 , w_7934 );
and ( \2512_b0 , \2509_b0 , w_7935 );
and ( w_7934 ,  , w_7935 );
buf ( w_7933 , \2511_b1 );
not ( w_7933 , w_7936 );
not (  , w_7937 );
and ( w_7936 , w_7937 , \2511_b0 );
or ( \2513_b1 , \2506_b1 , \2512_b1 );
xor ( \2513_b0 , \2506_b0 , w_7938 );
not ( w_7938 , w_7939 );
and ( w_7939 , \2512_b1 , \2512_b0 );
or ( \2514_b1 , \2365_b1 , \2372_b1 );
xor ( \2514_b0 , \2365_b0 , w_7940 );
not ( w_7940 , w_7941 );
and ( w_7941 , \2372_b1 , \2372_b0 );
or ( \2515_b1 , \2514_b1 , \2379_b1 );
not ( \2379_b1 , w_7942 );
and ( \2515_b0 , \2514_b0 , w_7943 );
and ( w_7942 , w_7943 , \2379_b0 );
or ( \2516_b1 , \2365_b1 , \2372_b1 );
not ( \2372_b1 , w_7944 );
and ( \2516_b0 , \2365_b0 , w_7945 );
and ( w_7944 , w_7945 , \2372_b0 );
or ( \2517_b1 , \2515_b1 , w_7946 );
or ( \2517_b0 , \2515_b0 , \2516_b0 );
not ( \2516_b0 , w_7947 );
and ( w_7947 , w_7946 , \2516_b1 );
or ( \2518_b1 , \2513_b1 , \2517_b1 );
xor ( \2518_b0 , \2513_b0 , w_7948 );
not ( w_7948 , w_7949 );
and ( w_7949 , \2517_b1 , \2517_b0 );
buf ( \2519_b1 , \2399_b1 );
not ( \2519_b1 , w_7950 );
not ( \2519_b0 , w_7951 );
and ( w_7950 , w_7951 , \2399_b0 );
buf ( \2520_b1 , \2292_b1 );
not ( \2520_b1 , w_7952 );
not ( \2520_b0 , w_7953 );
and ( w_7952 , w_7953 , \2292_b0 );
or ( \2521_b1 , \2519_b1 , w_7954 );
or ( \2521_b0 , \2519_b0 , \2520_b0 );
not ( \2520_b0 , w_7955 );
and ( w_7955 , w_7954 , \2520_b1 );
buf ( \2522_b1 , \c[7]_b1 );
not ( \2522_b1 , w_7956 );
not ( \2522_b0 , w_7957 );
and ( w_7956 , w_7957 , \c[7]_b0 );
or ( \2523_b1 , \2522_b1 , w_7959 );
not ( w_7959 , w_7960 );
and ( \2523_b0 , \2522_b0 , w_7961 );
and ( w_7960 ,  , w_7961 );
buf ( w_7959 , \b[9]_b1 );
not ( w_7959 , w_7962 );
not (  , w_7963 );
and ( w_7962 , w_7963 , \b[9]_b0 );
buf ( \2524_b1 , \2523_b1 );
not ( \2524_b1 , w_7964 );
not ( \2524_b0 , w_7965 );
and ( w_7964 , w_7965 , \2523_b0 );
buf ( \2525_b1 , \b[9]_b1 );
not ( \2525_b1 , w_7966 );
not ( \2525_b0 , w_7967 );
and ( w_7966 , w_7967 , \b[9]_b0 );
or ( \2526_b1 , \2525_b1 , w_7969 );
not ( w_7969 , w_7970 );
and ( \2526_b0 , \2525_b0 , w_7971 );
and ( w_7970 ,  , w_7971 );
buf ( w_7969 , \c[7]_b1 );
not ( w_7969 , w_7972 );
not (  , w_7973 );
and ( w_7972 , w_7973 , \c[7]_b0 );
buf ( \2527_b1 , \2526_b1 );
not ( \2527_b1 , w_7974 );
not ( \2527_b0 , w_7975 );
and ( w_7974 , w_7975 , \2526_b0 );
or ( \2528_b1 , \2524_b1 , w_7976 );
or ( \2528_b0 , \2524_b0 , \2527_b0 );
not ( \2527_b0 , w_7977 );
and ( w_7977 , w_7976 , \2527_b1 );
or ( \2529_b1 , \2528_b1 , w_7979 );
not ( w_7979 , w_7980 );
and ( \2529_b0 , \2528_b0 , w_7981 );
and ( w_7980 ,  , w_7981 );
buf ( w_7979 , \714_b1 );
not ( w_7979 , w_7982 );
not (  , w_7983 );
and ( w_7982 , w_7983 , \714_b0 );
or ( \2530_b1 , \2521_b1 , w_7985 );
not ( w_7985 , w_7986 );
and ( \2530_b0 , \2521_b0 , w_7987 );
and ( w_7986 ,  , w_7987 );
buf ( w_7985 , \2529_b1 );
not ( w_7985 , w_7988 );
not (  , w_7989 );
and ( w_7988 , w_7989 , \2529_b0 );
buf ( \2531_b1 , \2405_b1 );
not ( \2531_b1 , w_7990 );
not ( \2531_b0 , w_7991 );
and ( w_7990 , w_7991 , \2405_b0 );
buf ( \2532_b1 , \2281_b1 );
not ( \2532_b1 , w_7992 );
not ( \2532_b0 , w_7993 );
and ( w_7992 , w_7993 , \2281_b0 );
or ( \2533_b1 , \2531_b1 , w_7994 );
or ( \2533_b0 , \2531_b0 , \2532_b0 );
not ( \2532_b0 , w_7995 );
and ( w_7995 , w_7994 , \2532_b1 );
or ( \2534_b1 , \b[7]_b1 , \c[9]_b1 );
xor ( \2534_b0 , \b[7]_b0 , w_7996 );
not ( w_7996 , w_7997 );
and ( w_7997 , \c[9]_b1 , \c[9]_b0 );
or ( \2535_b1 , \2284_b1 , w_7999 );
not ( w_7999 , w_8000 );
and ( \2535_b0 , \2284_b0 , w_8001 );
and ( w_8000 ,  , w_8001 );
buf ( w_7999 , \2534_b1 );
not ( w_7999 , w_8002 );
not (  , w_8003 );
and ( w_8002 , w_8003 , \2534_b0 );
or ( \2536_b1 , \2533_b1 , w_8005 );
not ( w_8005 , w_8006 );
and ( \2536_b0 , \2533_b0 , w_8007 );
and ( w_8006 ,  , w_8007 );
buf ( w_8005 , \2535_b1 );
not ( w_8005 , w_8008 );
not (  , w_8009 );
and ( w_8008 , w_8009 , \2535_b0 );
or ( \2537_b1 , \2530_b1 , \2536_b1 );
xor ( \2537_b0 , \2530_b0 , w_8010 );
not ( w_8010 , w_8011 );
and ( w_8011 , \2536_b1 , \2536_b0 );
buf ( \2538_b1 , \2419_b1 );
not ( \2538_b1 , w_8012 );
not ( \2538_b0 , w_8013 );
and ( w_8012 , w_8013 , \2419_b0 );
buf ( \2539_b1 , \2252_b1 );
not ( \2539_b1 , w_8014 );
not ( \2539_b0 , w_8015 );
and ( w_8014 , w_8015 , \2252_b0 );
or ( \2540_b1 , \2538_b1 , w_8016 );
or ( \2540_b0 , \2538_b0 , \2539_b0 );
not ( \2539_b0 , w_8017 );
and ( w_8017 , w_8016 , \2539_b1 );
or ( \2541_b1 , \b[3]_b1 , \c[13]_b1 );
xor ( \2541_b0 , \b[3]_b0 , w_8018 );
not ( w_8018 , w_8019 );
and ( w_8019 , \c[13]_b1 , \c[13]_b0 );
or ( \2542_b1 , \2246_b1 , w_8021 );
not ( w_8021 , w_8022 );
and ( \2542_b0 , \2246_b0 , w_8023 );
and ( w_8022 ,  , w_8023 );
buf ( w_8021 , \2541_b1 );
not ( w_8021 , w_8024 );
not (  , w_8025 );
and ( w_8024 , w_8025 , \2541_b0 );
or ( \2543_b1 , \2540_b1 , w_8027 );
not ( w_8027 , w_8028 );
and ( \2543_b0 , \2540_b0 , w_8029 );
and ( w_8028 ,  , w_8029 );
buf ( w_8027 , \2542_b1 );
not ( w_8027 , w_8030 );
not (  , w_8031 );
and ( w_8030 , w_8031 , \2542_b0 );
buf ( \2544_b1 , \2543_b1 );
not ( \2544_b1 , w_8032 );
not ( \2544_b0 , w_8033 );
and ( w_8032 , w_8033 , \2543_b0 );
or ( \2545_b1 , \b[1]_b1 , w_8034 );
xor ( \2545_b0 , \b[1]_b0 , w_8036 );
not ( w_8036 , w_8037 );
and ( w_8037 , w_8034 , w_8035 );
buf ( w_8034 , \c[15]_b1 );
not ( w_8034 , w_8038 );
not ( w_8035 , w_8039 );
and ( w_8038 , w_8039 , \c[15]_b0 );
or ( \2546_b1 , \2364_b1 , \2545_b1 );
not ( \2545_b1 , w_8040 );
and ( \2546_b0 , \2364_b0 , w_8041 );
and ( w_8040 , w_8041 , \2545_b0 );
buf ( \2547_b1 , \2364_b1 );
not ( \2547_b1 , w_8042 );
not ( \2547_b0 , w_8043 );
and ( w_8042 , w_8043 , \2364_b0 );
or ( \2548_b1 , \c[15]_b1 , \c[14]_b1 );
xor ( \2548_b0 , \c[15]_b0 , w_8044 );
not ( w_8044 , w_8045 );
and ( w_8045 , \c[14]_b1 , \c[14]_b0 );
or ( \2549_b1 , \b[0]_b1 , \c[15]_b1 );
xor ( \2549_b0 , \b[0]_b0 , w_8046 );
not ( w_8046 , w_8047 );
and ( w_8047 , \c[15]_b1 , \c[15]_b0 );
or ( \2550_b1 , \2548_b1 , w_8049 );
not ( w_8049 , w_8050 );
and ( \2550_b0 , \2548_b0 , w_8051 );
and ( w_8050 ,  , w_8051 );
buf ( w_8049 , \2549_b1 );
not ( w_8049 , w_8052 );
not (  , w_8053 );
and ( w_8052 , w_8053 , \2549_b0 );
or ( \2551_b1 , \2547_b1 , \2550_b1 );
not ( \2550_b1 , w_8054 );
and ( \2551_b0 , \2547_b0 , w_8055 );
and ( w_8054 , w_8055 , \2550_b0 );
or ( \2552_b1 , \2546_b1 , w_8056 );
or ( \2552_b0 , \2546_b0 , \2551_b0 );
not ( \2551_b0 , w_8057 );
and ( w_8057 , w_8056 , \2551_b1 );
buf ( \2553_b1 , \2552_b1 );
not ( \2553_b1 , w_8058 );
not ( \2553_b0 , w_8059 );
and ( w_8058 , w_8059 , \2552_b0 );
or ( \2554_b1 , \2544_b1 , \2553_b1 );
not ( \2553_b1 , w_8060 );
and ( \2554_b0 , \2544_b0 , w_8061 );
and ( w_8060 , w_8061 , \2553_b0 );
or ( \2555_b1 , \2543_b1 , \2552_b1 );
not ( \2552_b1 , w_8062 );
and ( \2555_b0 , \2543_b0 , w_8063 );
and ( w_8062 , w_8063 , \2552_b0 );
or ( \2556_b1 , \2554_b1 , w_8065 );
not ( w_8065 , w_8066 );
and ( \2556_b0 , \2554_b0 , w_8067 );
and ( w_8066 ,  , w_8067 );
buf ( w_8065 , \2555_b1 );
not ( w_8065 , w_8068 );
not (  , w_8069 );
and ( w_8068 , w_8069 , \2555_b0 );
or ( \2557_b1 , \2537_b1 , \2556_b1 );
xor ( \2557_b0 , \2537_b0 , w_8070 );
not ( w_8070 , w_8071 );
and ( w_8071 , \2556_b1 , \2556_b0 );
or ( \2558_b1 , \2518_b1 , w_8072 );
xor ( \2558_b0 , \2518_b0 , w_8074 );
not ( w_8074 , w_8075 );
and ( w_8075 , w_8072 , w_8073 );
buf ( w_8072 , \2557_b1 );
not ( w_8072 , w_8076 );
not ( w_8073 , w_8077 );
and ( w_8076 , w_8077 , \2557_b0 );
buf ( \2559_b1 , \2558_b1 );
not ( \2559_b1 , w_8078 );
not ( \2559_b0 , w_8079 );
and ( w_8078 , w_8079 , \2558_b0 );
or ( \2560_b1 , \2421_b1 , \2427_b1 );
xor ( \2560_b0 , \2421_b0 , w_8080 );
not ( w_8080 , w_8081 );
and ( w_8081 , \2427_b1 , \2427_b0 );
or ( \2561_b1 , \2560_b1 , \2439_b1 );
not ( \2439_b1 , w_8082 );
and ( \2561_b0 , \2560_b0 , w_8083 );
and ( w_8082 , w_8083 , \2439_b0 );
or ( \2562_b1 , \2421_b1 , \2427_b1 );
not ( \2427_b1 , w_8084 );
and ( \2562_b0 , \2421_b0 , w_8085 );
and ( w_8084 , w_8085 , \2427_b0 );
or ( \2563_b1 , \2561_b1 , w_8086 );
or ( \2563_b0 , \2561_b0 , \2562_b0 );
not ( \2562_b0 , w_8087 );
and ( w_8087 , w_8086 , \2562_b1 );
buf ( \2564_b1 , \2563_b1 );
not ( \2564_b1 , w_8088 );
not ( \2564_b0 , w_8089 );
and ( w_8088 , w_8089 , \2563_b0 );
buf ( \2565_b1 , \2370_b1 );
not ( \2565_b1 , w_8090 );
not ( \2565_b0 , w_8091 );
and ( w_8090 , w_8091 , \2370_b0 );
buf ( \2566_b1 , \679_b1 );
not ( \2566_b1 , w_8092 );
not ( \2566_b0 , w_8093 );
and ( w_8092 , w_8093 , \679_b0 );
or ( \2567_b1 , \2565_b1 , w_8094 );
or ( \2567_b0 , \2565_b0 , \2566_b0 );
not ( \2566_b0 , w_8095 );
and ( w_8095 , w_8094 , \2566_b1 );
or ( \2568_b1 , \b[15]_b1 , \c[1]_b1 );
xor ( \2568_b0 , \b[15]_b0 , w_8096 );
not ( w_8096 , w_8097 );
and ( w_8097 , \c[1]_b1 , \c[1]_b0 );
or ( \2569_b1 , \2568_b1 , w_8099 );
not ( w_8099 , w_8100 );
and ( \2569_b0 , \2568_b0 , w_8101 );
and ( w_8100 ,  , w_8101 );
buf ( w_8099 , \c[0]_b1 );
not ( w_8099 , w_8102 );
not (  , w_8103 );
and ( w_8102 , w_8103 , \c[0]_b0 );
or ( \2570_b1 , \2567_b1 , w_8105 );
not ( w_8105 , w_8106 );
and ( \2570_b0 , \2567_b0 , w_8107 );
and ( w_8106 ,  , w_8107 );
buf ( w_8105 , \2569_b1 );
not ( w_8105 , w_8108 );
not (  , w_8109 );
and ( w_8108 , w_8109 , \2569_b0 );
or ( \2571_b1 , \b[0]_b1 , w_8110 );
or ( \2571_b0 , \b[0]_b0 , \c[14]_b0 );
not ( \c[14]_b0 , w_8111 );
and ( w_8111 , w_8110 , \c[14]_b1 );
or ( \2572_b1 , \2571_b1 , w_8113 );
not ( w_8113 , w_8114 );
and ( \2572_b0 , \2571_b0 , w_8115 );
and ( w_8114 ,  , w_8115 );
buf ( w_8113 , \c[13]_b1 );
not ( w_8113 , w_8116 );
not (  , w_8117 );
and ( w_8116 , w_8117 , \c[13]_b0 );
or ( \2573_b1 , \b[0]_b1 , w_8119 );
not ( w_8119 , w_8120 );
and ( \2573_b0 , \b[0]_b0 , w_8121 );
and ( w_8120 ,  , w_8121 );
buf ( w_8119 , \c[14]_b1 );
not ( w_8119 , w_8122 );
not (  , w_8123 );
and ( w_8122 , w_8123 , \c[14]_b0 );
or ( \2575_b1 , \2570_b1 , \2574_b1 );
xor ( \2575_b0 , \2570_b0 , w_8124 );
not ( w_8124 , w_8125 );
and ( w_8125 , \2574_b1 , \2574_b0 );
buf ( \2576_b1 , \2425_b1 );
not ( \2576_b1 , w_8126 );
not ( \2576_b0 , w_8127 );
and ( w_8126 , w_8127 , \2425_b0 );
buf ( \2577_b1 , \2238_b1 );
not ( \2577_b1 , w_8128 );
not ( \2577_b0 , w_8129 );
and ( w_8128 , w_8129 , \2238_b0 );
or ( \2578_b1 , \2576_b1 , w_8130 );
or ( \2578_b0 , \2576_b0 , \2577_b0 );
not ( \2577_b0 , w_8131 );
and ( w_8131 , w_8130 , \2577_b1 );
or ( \2579_b1 , \b[5]_b1 , \c[11]_b1 );
xor ( \2579_b0 , \b[5]_b0 , w_8132 );
not ( w_8132 , w_8133 );
and ( w_8133 , \c[11]_b1 , \c[11]_b0 );
or ( \2580_b1 , \2236_b1 , w_8135 );
not ( w_8135 , w_8136 );
and ( \2580_b0 , \2236_b0 , w_8137 );
and ( w_8136 ,  , w_8137 );
buf ( w_8135 , \2579_b1 );
not ( w_8135 , w_8138 );
not (  , w_8139 );
and ( w_8138 , w_8139 , \2579_b0 );
or ( \2581_b1 , \2578_b1 , w_8141 );
not ( w_8141 , w_8142 );
and ( \2581_b0 , \2578_b0 , w_8143 );
and ( w_8142 ,  , w_8143 );
buf ( w_8141 , \2580_b1 );
not ( w_8141 , w_8144 );
not (  , w_8145 );
and ( w_8144 , w_8145 , \2580_b0 );
or ( \2582_b1 , \2575_b1 , \2581_b1 );
xor ( \2582_b0 , \2575_b0 , w_8146 );
not ( w_8146 , w_8147 );
and ( w_8147 , \2581_b1 , \2581_b0 );
buf ( \2583_b1 , \2582_b1 );
not ( \2583_b1 , w_8148 );
not ( \2583_b0 , w_8149 );
and ( w_8148 , w_8149 , \2582_b0 );
or ( \2584_b1 , \2564_b1 , \2583_b1 );
not ( \2583_b1 , w_8150 );
and ( \2584_b0 , \2564_b0 , w_8151 );
and ( w_8150 , w_8151 , \2583_b0 );
or ( \2585_b1 , \2563_b1 , \2582_b1 );
not ( \2582_b1 , w_8152 );
and ( \2585_b0 , \2563_b0 , w_8153 );
and ( w_8152 , w_8153 , \2582_b0 );
or ( \2586_b1 , \2584_b1 , w_8155 );
not ( w_8155 , w_8156 );
and ( \2586_b0 , \2584_b0 , w_8157 );
and ( w_8156 ,  , w_8157 );
buf ( w_8155 , \2585_b1 );
not ( w_8155 , w_8158 );
not (  , w_8159 );
and ( w_8158 , w_8159 , \2585_b0 );
or ( \2587_b1 , \2401_b1 , \2407_b1 );
xor ( \2587_b0 , \2401_b0 , w_8160 );
not ( w_8160 , w_8161 );
and ( w_8161 , \2407_b1 , \2407_b0 );
or ( \2588_b1 , \2587_b1 , \2414_b1 );
not ( \2414_b1 , w_8162 );
and ( \2588_b0 , \2587_b0 , w_8163 );
and ( w_8162 , w_8163 , \2414_b0 );
or ( \2589_b1 , \2401_b1 , \2407_b1 );
not ( \2407_b1 , w_8164 );
and ( \2589_b0 , \2401_b0 , w_8165 );
and ( w_8164 , w_8165 , \2407_b0 );
or ( \2590_b1 , \2588_b1 , w_8166 );
or ( \2590_b0 , \2588_b0 , \2589_b0 );
not ( \2589_b0 , w_8167 );
and ( w_8167 , w_8166 , \2589_b1 );
or ( \2591_b1 , \2586_b1 , \2590_b1 );
xor ( \2591_b0 , \2586_b0 , w_8168 );
not ( w_8168 , w_8169 );
and ( w_8169 , \2590_b1 , \2590_b0 );
buf ( \2592_b1 , \2591_b1 );
not ( \2592_b1 , w_8170 );
not ( \2592_b0 , w_8171 );
and ( w_8170 , w_8171 , \2591_b0 );
or ( \2593_b1 , \2559_b1 , w_8172 );
or ( \2593_b0 , \2559_b0 , \2592_b0 );
not ( \2592_b0 , w_8173 );
and ( w_8173 , w_8172 , \2592_b1 );
or ( \2594_b1 , \2591_b1 , w_8174 );
or ( \2594_b0 , \2591_b0 , \2558_b0 );
not ( \2558_b0 , w_8175 );
and ( w_8175 , w_8174 , \2558_b1 );
or ( \2595_b1 , \2593_b1 , w_8177 );
not ( w_8177 , w_8178 );
and ( \2595_b0 , \2593_b0 , w_8179 );
and ( w_8178 ,  , w_8179 );
buf ( w_8177 , \2594_b1 );
not ( w_8177 , w_8180 );
not (  , w_8181 );
and ( w_8180 , w_8181 , \2594_b0 );
or ( \2596_b1 , \2500_b1 , \2595_b1 );
xor ( \2596_b0 , \2500_b0 , w_8182 );
not ( w_8182 , w_8183 );
and ( w_8183 , \2595_b1 , \2595_b0 );
or ( \2597_b1 , \2486_b1 , \2596_b1 );
xor ( \2597_b0 , \2486_b0 , w_8184 );
not ( w_8184 , w_8185 );
and ( w_8185 , \2596_b1 , \2596_b0 );
buf ( \2598_b1 , \2597_b1 );
not ( \2598_b1 , w_8186 );
not ( \2598_b0 , w_8187 );
and ( w_8186 , w_8187 , \2597_b0 );
or ( \2599_b1 , \2363_b1 , \2394_b1 );
xor ( \2599_b0 , \2363_b0 , w_8188 );
not ( w_8188 , w_8189 );
and ( w_8189 , \2394_b1 , \2394_b0 );
or ( \2600_b1 , \2599_b1 , \2483_b1 );
xor ( \2600_b0 , \2599_b0 , w_8190 );
not ( w_8190 , w_8191 );
and ( w_8191 , \2483_b1 , \2483_b0 );
buf ( \2601_b1 , \2600_b1 );
not ( \2601_b1 , w_8192 );
not ( \2601_b0 , w_8193 );
and ( w_8192 , w_8193 , \2600_b0 );
or ( \2602_b1 , \2463_b1 , \2479_b1 );
xor ( \2602_b0 , \2463_b0 , w_8194 );
not ( w_8194 , w_8195 );
and ( w_8195 , \2479_b1 , \2479_b0 );
or ( \2603_b1 , \2602_b1 , w_8196 );
xor ( \2603_b0 , \2602_b0 , w_8198 );
not ( w_8198 , w_8199 );
and ( w_8199 , w_8196 , w_8197 );
buf ( w_8196 , \2462_b1 );
not ( w_8196 , w_8200 );
not ( w_8197 , w_8201 );
and ( w_8200 , w_8201 , \2462_b0 );
buf ( \2604_b1 , \2603_b1 );
not ( \2604_b1 , w_8202 );
not ( \2604_b0 , w_8203 );
and ( w_8202 , w_8203 , \2603_b0 );
buf ( \2605_b1 , \2604_b1 );
not ( \2605_b1 , w_8204 );
not ( \2605_b0 , w_8205 );
and ( w_8204 , w_8205 , \2604_b0 );
buf ( \2606_b1 , \2275_b1 );
not ( \2606_b1 , w_8206 );
not ( \2606_b0 , w_8207 );
and ( w_8206 , w_8207 , \2275_b0 );
buf ( \2607_b1 , \2304_b1 );
not ( \2607_b1 , w_8208 );
not ( \2607_b0 , w_8209 );
and ( w_8208 , w_8209 , \2304_b0 );
buf ( \2608_b1 , \2607_b1 );
not ( \2608_b1 , w_8210 );
not ( \2608_b0 , w_8211 );
and ( w_8210 , w_8211 , \2607_b0 );
or ( \2609_b1 , \2606_b1 , w_8212 );
or ( \2609_b0 , \2606_b0 , \2608_b0 );
not ( \2608_b0 , w_8213 );
and ( w_8213 , w_8212 , \2608_b1 );
or ( \2610_b1 , \2361_b1 , w_8215 );
not ( w_8215 , w_8216 );
and ( \2610_b0 , \2361_b0 , w_8217 );
and ( w_8216 ,  , w_8217 );
buf ( w_8215 , \2304_b1 );
not ( w_8215 , w_8218 );
not (  , w_8219 );
and ( w_8218 , w_8219 , \2304_b0 );
or ( \2611_b1 , \2609_b1 , w_8221 );
not ( w_8221 , w_8222 );
and ( \2611_b0 , \2609_b0 , w_8223 );
and ( w_8222 ,  , w_8223 );
buf ( w_8221 , \2610_b1 );
not ( w_8221 , w_8224 );
not (  , w_8225 );
and ( w_8224 , w_8225 , \2610_b0 );
or ( \2612_b1 , \2611_b1 , \2358_b1 );
not ( \2358_b1 , w_8226 );
and ( \2612_b0 , \2611_b0 , w_8227 );
and ( w_8226 , w_8227 , \2358_b0 );
buf ( \2613_b1 , \2611_b1 );
not ( \2613_b1 , w_8228 );
not ( \2613_b0 , w_8229 );
and ( w_8228 , w_8229 , \2611_b0 );
buf ( \2614_b1 , \2358_b1 );
not ( \2614_b1 , w_8230 );
not ( \2614_b0 , w_8231 );
and ( w_8230 , w_8231 , \2358_b0 );
or ( \2615_b1 , \2613_b1 , \2614_b1 );
not ( \2614_b1 , w_8232 );
and ( \2615_b0 , \2613_b0 , w_8233 );
and ( w_8232 , w_8233 , \2614_b0 );
or ( \2616_b1 , \2612_b1 , w_8235 );
not ( w_8235 , w_8236 );
and ( \2616_b0 , \2612_b0 , w_8237 );
and ( w_8236 ,  , w_8237 );
buf ( w_8235 , \2615_b1 );
not ( w_8235 , w_8238 );
not (  , w_8239 );
and ( w_8238 , w_8239 , \2615_b0 );
buf ( \2617_b1 , \2616_b1 );
not ( \2617_b1 , w_8240 );
not ( \2617_b0 , w_8241 );
and ( w_8240 , w_8241 , \2616_b0 );
or ( \2618_b1 , \2605_b1 , w_8242 );
or ( \2618_b0 , \2605_b0 , \2617_b0 );
not ( \2617_b0 , w_8243 );
and ( w_8243 , w_8242 , \2617_b1 );
buf ( \2619_b1 , \2603_b1 );
not ( \2619_b1 , w_8244 );
not ( \2619_b0 , w_8245 );
and ( w_8244 , w_8245 , \2603_b0 );
buf ( \2620_b1 , \2616_b1 );
not ( \2620_b1 , w_8246 );
not ( \2620_b0 , w_8247 );
and ( w_8246 , w_8247 , \2616_b0 );
buf ( \2621_b1 , \2620_b1 );
not ( \2621_b1 , w_8248 );
not ( \2621_b0 , w_8249 );
and ( w_8248 , w_8249 , \2620_b0 );
or ( \2622_b1 , \2619_b1 , w_8250 );
or ( \2622_b0 , \2619_b0 , \2621_b0 );
not ( \2621_b0 , w_8251 );
and ( w_8251 , w_8250 , \2621_b1 );
or ( \2623_b1 , \2465_b1 , \2470_b1 );
xor ( \2623_b0 , \2465_b0 , w_8252 );
not ( w_8252 , w_8253 );
and ( w_8253 , \2470_b1 , \2470_b0 );
or ( \2624_b1 , \2623_b1 , \2476_b1 );
xor ( \2624_b0 , \2623_b0 , w_8254 );
not ( w_8254 , w_8255 );
and ( w_8255 , \2476_b1 , \2476_b0 );
buf ( \2625_b1 , \2624_b1 );
not ( \2625_b1 , w_8256 );
not ( \2625_b0 , w_8257 );
and ( w_8256 , w_8257 , \2624_b0 );
or ( \2626_b1 , \2446_b1 , \2452_b1 );
xor ( \2626_b0 , \2446_b0 , w_8258 );
not ( w_8258 , w_8259 );
and ( w_8259 , \2452_b1 , \2452_b0 );
or ( \2627_b1 , \2626_b1 , \2459_b1 );
xor ( \2627_b0 , \2626_b0 , w_8260 );
not ( w_8260 , w_8261 );
and ( w_8261 , \2459_b1 , \2459_b0 );
buf ( \2628_b1 , \2627_b1 );
not ( \2628_b1 , w_8262 );
not ( \2628_b0 , w_8263 );
and ( w_8262 , w_8263 , \2627_b0 );
or ( \2629_b1 , \2625_b1 , w_8264 );
or ( \2629_b0 , \2625_b0 , \2628_b0 );
not ( \2628_b0 , w_8265 );
and ( w_8265 , w_8264 , \2628_b1 );
or ( \2630_b1 , \2627_b1 , w_8266 );
or ( \2630_b0 , \2627_b0 , \2624_b0 );
not ( \2624_b0 , w_8267 );
and ( w_8267 , w_8266 , \2624_b1 );
or ( \2631_b1 , \c[11]_b1 , \b[0]_b1 );
xor ( \2631_b0 , \c[11]_b0 , w_8268 );
not ( w_8268 , w_8269 );
and ( w_8269 , \b[0]_b1 , \b[0]_b0 );
buf ( \2632_b1 , \2631_b1 );
not ( \2632_b1 , w_8270 );
not ( \2632_b0 , w_8271 );
and ( w_8270 , w_8271 , \2631_b0 );
buf ( \2633_b1 , \2238_b1 );
not ( \2633_b1 , w_8272 );
not ( \2633_b0 , w_8273 );
and ( w_8272 , w_8273 , \2238_b0 );
or ( \2634_b1 , \2632_b1 , w_8274 );
or ( \2634_b0 , \2632_b0 , \2633_b0 );
not ( \2633_b0 , w_8275 );
and ( w_8275 , w_8274 , \2633_b1 );
or ( \2635_b1 , \2236_b1 , w_8277 );
not ( w_8277 , w_8278 );
and ( \2635_b0 , \2236_b0 , w_8279 );
and ( w_8278 ,  , w_8279 );
buf ( w_8277 , \2454_b1 );
not ( w_8277 , w_8280 );
not (  , w_8281 );
and ( w_8280 , w_8281 , \2454_b0 );
or ( \2636_b1 , \2634_b1 , w_8283 );
not ( w_8283 , w_8284 );
and ( \2636_b0 , \2634_b0 , w_8285 );
and ( w_8284 ,  , w_8285 );
buf ( w_8283 , \2635_b1 );
not ( w_8283 , w_8286 );
not (  , w_8287 );
and ( w_8286 , w_8287 , \2635_b0 );
buf ( \2637_b1 , \2636_b1 );
not ( \2637_b1 , w_8288 );
not ( \2637_b0 , w_8289 );
and ( w_8288 , w_8289 , \2636_b0 );
or ( \2638_b1 , \b[6]_b1 , \c[5]_b1 );
xor ( \2638_b0 , \b[6]_b0 , w_8290 );
not ( w_8290 , w_8291 );
and ( w_8291 , \c[5]_b1 , \c[5]_b0 );
buf ( \2639_b1 , \2638_b1 );
not ( \2639_b1 , w_8292 );
not ( \2639_b0 , w_8293 );
and ( w_8292 , w_8293 , \2638_b0 );
buf ( \2640_b1 , \2265_b1 );
not ( \2640_b1 , w_8294 );
not ( \2640_b0 , w_8295 );
and ( w_8294 , w_8295 , \2265_b0 );
or ( \2641_b1 , \2639_b1 , w_8296 );
or ( \2641_b0 , \2639_b0 , \2640_b0 );
not ( \2640_b0 , w_8297 );
and ( w_8297 , w_8296 , \2640_b1 );
or ( \2642_b1 , \739_b1 , w_8299 );
not ( w_8299 , w_8300 );
and ( \2642_b0 , \739_b0 , w_8301 );
and ( w_8300 ,  , w_8301 );
buf ( w_8299 , \2307_b1 );
not ( w_8299 , w_8302 );
not (  , w_8303 );
and ( w_8302 , w_8303 , \2307_b0 );
or ( \2643_b1 , \2641_b1 , w_8305 );
not ( w_8305 , w_8306 );
and ( \2643_b0 , \2641_b0 , w_8307 );
and ( w_8306 ,  , w_8307 );
buf ( w_8305 , \2642_b1 );
not ( w_8305 , w_8308 );
not (  , w_8309 );
and ( w_8308 , w_8309 , \2642_b0 );
buf ( \2644_b1 , \2643_b1 );
not ( \2644_b1 , w_8310 );
not ( \2644_b0 , w_8311 );
and ( w_8310 , w_8311 , \2643_b0 );
or ( \2645_b1 , \2637_b1 , w_8313 );
not ( w_8313 , w_8314 );
and ( \2645_b0 , \2637_b0 , w_8315 );
and ( w_8314 ,  , w_8315 );
buf ( w_8313 , \2644_b1 );
not ( w_8313 , w_8316 );
not (  , w_8317 );
and ( w_8316 , w_8317 , \2644_b0 );
buf ( \2646_b1 , \2645_b1 );
not ( \2646_b1 , w_8318 );
not ( \2646_b0 , w_8319 );
and ( w_8318 , w_8319 , \2645_b0 );
or ( \2647_b1 , \2320_b1 , \2325_b1 );
not ( \2325_b1 , w_8320 );
and ( \2647_b0 , \2320_b0 , w_8321 );
and ( w_8320 , w_8321 , \2325_b0 );
buf ( \2648_b1 , \2320_b1 );
not ( \2648_b1 , w_8322 );
not ( \2648_b0 , w_8323 );
and ( w_8322 , w_8323 , \2320_b0 );
or ( \2649_b1 , \2648_b1 , \2324_b1 );
not ( \2324_b1 , w_8324 );
and ( \2649_b0 , \2648_b0 , w_8325 );
and ( w_8324 , w_8325 , \2324_b0 );
or ( \2650_b1 , \2647_b1 , w_8327 );
not ( w_8327 , w_8328 );
and ( \2650_b0 , \2647_b0 , w_8329 );
and ( w_8328 ,  , w_8329 );
buf ( w_8327 , \2649_b1 );
not ( w_8327 , w_8330 );
not (  , w_8331 );
and ( w_8330 , w_8331 , \2649_b0 );
buf ( \2651_b1 , \2650_b1 );
not ( \2651_b1 , w_8332 );
not ( \2651_b0 , w_8333 );
and ( w_8332 , w_8333 , \2650_b0 );
or ( \2652_b1 , \2646_b1 , w_8334 );
or ( \2652_b0 , \2646_b0 , \2651_b0 );
not ( \2651_b0 , w_8335 );
and ( w_8335 , w_8334 , \2651_b1 );
or ( \2653_b1 , \2643_b1 , w_8337 );
not ( w_8337 , w_8338 );
and ( \2653_b0 , \2643_b0 , w_8339 );
and ( w_8338 ,  , w_8339 );
buf ( w_8337 , \2636_b1 );
not ( w_8337 , w_8340 );
not (  , w_8341 );
and ( w_8340 , w_8341 , \2636_b0 );
or ( \2654_b1 , \2652_b1 , w_8343 );
not ( w_8343 , w_8344 );
and ( \2654_b0 , \2652_b0 , w_8345 );
and ( w_8344 ,  , w_8345 );
buf ( w_8343 , \2653_b1 );
not ( w_8343 , w_8346 );
not (  , w_8347 );
and ( w_8346 , w_8347 , \2653_b0 );
or ( \2655_b1 , \2630_b1 , w_8349 );
not ( w_8349 , w_8350 );
and ( \2655_b0 , \2630_b0 , w_8351 );
and ( w_8350 ,  , w_8351 );
buf ( w_8349 , \2654_b1 );
not ( w_8349 , w_8352 );
not (  , w_8353 );
and ( w_8352 , w_8353 , \2654_b0 );
or ( \2656_b1 , \2629_b1 , w_8355 );
not ( w_8355 , w_8356 );
and ( \2656_b0 , \2629_b0 , w_8357 );
and ( w_8356 ,  , w_8357 );
buf ( w_8355 , \2655_b1 );
not ( w_8355 , w_8358 );
not (  , w_8359 );
and ( w_8358 , w_8359 , \2655_b0 );
or ( \2657_b1 , \2622_b1 , w_8361 );
not ( w_8361 , w_8362 );
and ( \2657_b0 , \2622_b0 , w_8363 );
and ( w_8362 ,  , w_8363 );
buf ( w_8361 , \2656_b1 );
not ( w_8361 , w_8364 );
not (  , w_8365 );
and ( w_8364 , w_8365 , \2656_b0 );
or ( \2658_b1 , \2618_b1 , w_8367 );
not ( w_8367 , w_8368 );
and ( \2658_b0 , \2618_b0 , w_8369 );
and ( w_8368 ,  , w_8369 );
buf ( w_8367 , \2657_b1 );
not ( w_8367 , w_8370 );
not (  , w_8371 );
and ( w_8370 , w_8371 , \2657_b0 );
buf ( \2659_b1 , \2658_b1 );
not ( \2659_b1 , w_8372 );
not ( \2659_b0 , w_8373 );
and ( w_8372 , w_8373 , \2658_b0 );
or ( \2660_b1 , \2601_b1 , \2659_b1 );
not ( \2659_b1 , w_8374 );
and ( \2660_b0 , \2601_b0 , w_8375 );
and ( w_8374 , w_8375 , \2659_b0 );
buf ( \2661_b1 , \2603_b1 );
not ( \2661_b1 , w_8376 );
not ( \2661_b0 , w_8377 );
and ( w_8376 , w_8377 , \2603_b0 );
buf ( \2662_b1 , \2656_b1 );
not ( \2662_b1 , w_8378 );
not ( \2662_b0 , w_8379 );
and ( w_8378 , w_8379 , \2656_b0 );
or ( \2663_b1 , \2661_b1 , w_8380 );
or ( \2663_b0 , \2661_b0 , \2662_b0 );
not ( \2662_b0 , w_8381 );
and ( w_8381 , w_8380 , \2662_b1 );
or ( \2664_b1 , \2603_b1 , w_8382 );
or ( \2664_b0 , \2603_b0 , \2656_b0 );
not ( \2656_b0 , w_8383 );
and ( w_8383 , w_8382 , \2656_b1 );
or ( \2665_b1 , \2663_b1 , w_8385 );
not ( w_8385 , w_8386 );
and ( \2665_b0 , \2663_b0 , w_8387 );
and ( w_8386 ,  , w_8387 );
buf ( w_8385 , \2664_b1 );
not ( w_8385 , w_8388 );
not (  , w_8389 );
and ( w_8388 , w_8389 , \2664_b0 );
or ( \2666_b1 , \2665_b1 , \2620_b1 );
not ( \2620_b1 , w_8390 );
and ( \2666_b0 , \2665_b0 , w_8391 );
and ( w_8390 , w_8391 , \2620_b0 );
buf ( \2667_b1 , \2665_b1 );
not ( \2667_b1 , w_8392 );
not ( \2667_b0 , w_8393 );
and ( w_8392 , w_8393 , \2665_b0 );
or ( \2668_b1 , \2667_b1 , \2616_b1 );
not ( \2616_b1 , w_8394 );
and ( \2668_b0 , \2667_b0 , w_8395 );
and ( w_8394 , w_8395 , \2616_b0 );
or ( \2669_b1 , \2666_b1 , w_8397 );
not ( w_8397 , w_8398 );
and ( \2669_b0 , \2666_b0 , w_8399 );
and ( w_8398 ,  , w_8399 );
buf ( w_8397 , \2668_b1 );
not ( w_8397 , w_8400 );
not (  , w_8401 );
and ( w_8400 , w_8401 , \2668_b0 );
or ( \2670_b1 , \2312_b1 , \2326_b1 );
xor ( \2670_b0 , \2312_b0 , w_8402 );
not ( w_8402 , w_8403 );
and ( w_8403 , \2326_b1 , \2326_b0 );
or ( \2671_b1 , \2670_b1 , w_8404 );
xor ( \2671_b0 , \2670_b0 , w_8406 );
not ( w_8406 , w_8407 );
and ( w_8407 , w_8404 , w_8405 );
buf ( w_8404 , \2356_b1 );
not ( w_8404 , w_8408 );
not ( w_8405 , w_8409 );
and ( w_8408 , w_8409 , \2356_b0 );
buf ( \2672_b1 , \2671_b1 );
not ( \2672_b1 , w_8410 );
not ( \2672_b0 , w_8411 );
and ( w_8410 , w_8411 , \2671_b0 );
or ( \2673_b1 , \2624_b1 , \2627_b1 );
xor ( \2673_b0 , \2624_b0 , w_8412 );
not ( w_8412 , w_8413 );
and ( w_8413 , \2627_b1 , \2627_b0 );
or ( \2674_b1 , \2673_b1 , w_8414 );
xor ( \2674_b0 , \2673_b0 , w_8416 );
not ( w_8416 , w_8417 );
and ( w_8417 , w_8414 , w_8415 );
buf ( w_8414 , \2654_b1 );
not ( w_8414 , w_8418 );
not ( w_8415 , w_8419 );
and ( w_8418 , w_8419 , \2654_b0 );
buf ( \2675_b1 , \2674_b1 );
not ( \2675_b1 , w_8420 );
not ( \2675_b0 , w_8421 );
and ( w_8420 , w_8421 , \2674_b0 );
or ( \2676_b1 , \2672_b1 , w_8422 );
or ( \2676_b0 , \2672_b0 , \2675_b0 );
not ( \2675_b0 , w_8423 );
and ( w_8423 , w_8422 , \2675_b1 );
or ( \2677_b1 , \2236_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_8424 );
and ( \2677_b0 , \2236_b0 , w_8425 );
and ( w_8424 , w_8425 , \b[0]_b0 );
or ( \2678_b1 , \b[3]_b1 , \c[7]_b1 );
xor ( \2678_b0 , \b[3]_b0 , w_8426 );
not ( w_8426 , w_8427 );
and ( w_8427 , \c[7]_b1 , \c[7]_b0 );
buf ( \2679_b1 , \2678_b1 );
not ( \2679_b1 , w_8428 );
not ( \2679_b0 , w_8429 );
and ( w_8428 , w_8429 , \2678_b0 );
buf ( \2680_b1 , \726_b1 );
not ( \2680_b1 , w_8430 );
not ( \2680_b0 , w_8431 );
and ( w_8430 , w_8431 , \726_b0 );
or ( \2681_b1 , \2679_b1 , w_8432 );
or ( \2681_b0 , \2679_b0 , \2680_b0 );
not ( \2680_b0 , w_8433 );
and ( w_8433 , w_8432 , \2680_b1 );
or ( \2682_b1 , \714_b1 , w_8435 );
not ( w_8435 , w_8436 );
and ( \2682_b0 , \714_b0 , w_8437 );
and ( w_8436 ,  , w_8437 );
buf ( w_8435 , \2348_b1 );
not ( w_8435 , w_8438 );
not (  , w_8439 );
and ( w_8438 , w_8439 , \2348_b0 );
or ( \2683_b1 , \2681_b1 , w_8441 );
not ( w_8441 , w_8442 );
and ( \2683_b0 , \2681_b0 , w_8443 );
and ( w_8442 ,  , w_8443 );
buf ( w_8441 , \2682_b1 );
not ( w_8441 , w_8444 );
not (  , w_8445 );
and ( w_8444 , w_8445 , \2682_b0 );
or ( \2684_b1 , \2677_b1 , \2683_b1 );
xor ( \2684_b0 , \2677_b0 , w_8446 );
not ( w_8446 , w_8447 );
and ( w_8447 , \2683_b1 , \2683_b0 );
or ( \2685_b1 , \b[7]_b1 , \c[3]_b1 );
xor ( \2685_b0 , \b[7]_b0 , w_8448 );
not ( w_8448 , w_8449 );
and ( w_8449 , \c[3]_b1 , \c[3]_b0 );
buf ( \2686_b1 , \2685_b1 );
not ( \2686_b1 , w_8450 );
not ( \2686_b0 , w_8451 );
and ( w_8450 , w_8451 , \2685_b0 );
buf ( \2687_b1 , \699_b1 );
not ( \2687_b1 , w_8452 );
not ( \2687_b0 , w_8453 );
and ( w_8452 , w_8453 , \699_b0 );
or ( \2688_b1 , \2686_b1 , w_8454 );
or ( \2688_b0 , \2686_b0 , \2687_b0 );
not ( \2687_b0 , w_8455 );
and ( w_8455 , w_8454 , \2687_b1 );
or ( \2689_b1 , \702_b1 , w_8457 );
not ( w_8457 , w_8458 );
and ( \2689_b0 , \702_b0 , w_8459 );
and ( w_8458 ,  , w_8459 );
buf ( w_8457 , \2314_b1 );
not ( w_8457 , w_8460 );
not (  , w_8461 );
and ( w_8460 , w_8461 , \2314_b0 );
or ( \2690_b1 , \2688_b1 , w_8463 );
not ( w_8463 , w_8464 );
and ( \2690_b0 , \2688_b0 , w_8465 );
and ( w_8464 ,  , w_8465 );
buf ( w_8463 , \2689_b1 );
not ( w_8463 , w_8466 );
not (  , w_8467 );
and ( w_8466 , w_8467 , \2689_b0 );
or ( \2691_b1 , \2684_b1 , \2690_b1 );
not ( \2690_b1 , w_8468 );
and ( \2691_b0 , \2684_b0 , w_8469 );
and ( w_8468 , w_8469 , \2690_b0 );
or ( \2692_b1 , \2677_b1 , \2683_b1 );
not ( \2683_b1 , w_8470 );
and ( \2692_b0 , \2677_b0 , w_8471 );
and ( w_8470 , w_8471 , \2683_b0 );
or ( \2693_b1 , \2691_b1 , w_8472 );
or ( \2693_b0 , \2691_b0 , \2692_b0 );
not ( \2692_b0 , w_8473 );
and ( w_8473 , w_8472 , \2692_b1 );
or ( \2694_b1 , \b[1]_b1 , \c[9]_b1 );
xor ( \2694_b0 , \b[1]_b0 , w_8474 );
not ( w_8474 , w_8475 );
and ( w_8475 , \c[9]_b1 , \c[9]_b0 );
buf ( \2695_b1 , \2694_b1 );
not ( \2695_b1 , w_8476 );
not ( \2695_b0 , w_8477 );
and ( w_8476 , w_8477 , \2694_b0 );
buf ( \2696_b1 , \2448_b1 );
not ( \2696_b1 , w_8478 );
not ( \2696_b0 , w_8479 );
and ( w_8478 , w_8479 , \2448_b0 );
or ( \2697_b1 , \2695_b1 , w_8480 );
or ( \2697_b0 , \2695_b0 , \2696_b0 );
not ( \2696_b0 , w_8481 );
and ( w_8481 , w_8480 , \2696_b1 );
or ( \2698_b1 , \2280_b1 , w_8483 );
not ( w_8483 , w_8484 );
and ( \2698_b0 , \2280_b0 , w_8485 );
and ( w_8484 ,  , w_8485 );
buf ( w_8483 , \2338_b1 );
not ( w_8483 , w_8486 );
not (  , w_8487 );
and ( w_8486 , w_8487 , \2338_b0 );
or ( \2699_b1 , \2697_b1 , w_8489 );
not ( w_8489 , w_8490 );
and ( \2699_b0 , \2697_b0 , w_8491 );
and ( w_8490 ,  , w_8491 );
buf ( w_8489 , \2698_b1 );
not ( w_8489 , w_8492 );
not (  , w_8493 );
and ( w_8492 , w_8493 , \2698_b0 );
or ( \2700_b1 , \b[9]_b1 , \c[1]_b1 );
xor ( \2700_b0 , \b[9]_b0 , w_8494 );
not ( w_8494 , w_8495 );
and ( w_8495 , \c[1]_b1 , \c[1]_b0 );
buf ( \2701_b1 , \2700_b1 );
not ( \2701_b1 , w_8496 );
not ( \2701_b0 , w_8497 );
and ( w_8496 , w_8497 , \2700_b0 );
buf ( \2702_b1 , \679_b1 );
not ( \2702_b1 , w_8498 );
not ( \2702_b0 , w_8499 );
and ( w_8498 , w_8499 , \679_b0 );
or ( \2703_b1 , \2701_b1 , w_8500 );
or ( \2703_b0 , \2701_b0 , \2702_b0 );
not ( \2702_b0 , w_8501 );
and ( w_8501 , w_8500 , \2702_b1 );
or ( \2704_b1 , \2330_b1 , w_8503 );
not ( w_8503 , w_8504 );
and ( \2704_b0 , \2330_b0 , w_8505 );
and ( w_8504 ,  , w_8505 );
buf ( w_8503 , \c[0]_b1 );
not ( w_8503 , w_8506 );
not (  , w_8507 );
and ( w_8506 , w_8507 , \c[0]_b0 );
or ( \2705_b1 , \2703_b1 , w_8509 );
not ( w_8509 , w_8510 );
and ( \2705_b0 , \2703_b0 , w_8511 );
and ( w_8510 ,  , w_8511 );
buf ( w_8509 , \2704_b1 );
not ( w_8509 , w_8512 );
not (  , w_8513 );
and ( w_8512 , w_8513 , \2704_b0 );
or ( \2706_b1 , \2699_b1 , w_8514 );
or ( \2706_b0 , \2699_b0 , \2705_b0 );
not ( \2705_b0 , w_8515 );
and ( w_8515 , w_8514 , \2705_b1 );
or ( \2707_b1 , \b[5]_b1 , \c[5]_b1 );
xor ( \2707_b0 , \b[5]_b0 , w_8516 );
not ( w_8516 , w_8517 );
and ( w_8517 , \c[5]_b1 , \c[5]_b0 );
buf ( \2708_b1 , \2707_b1 );
not ( \2708_b1 , w_8518 );
not ( \2708_b0 , w_8519 );
and ( w_8518 , w_8519 , \2707_b0 );
buf ( \2709_b1 , \736_b1 );
not ( \2709_b1 , w_8520 );
not ( \2709_b0 , w_8521 );
and ( w_8520 , w_8521 , \736_b0 );
or ( \2710_b1 , \2708_b1 , w_8522 );
or ( \2710_b0 , \2708_b0 , \2709_b0 );
not ( \2709_b0 , w_8523 );
and ( w_8523 , w_8522 , \2709_b1 );
or ( \2711_b1 , \739_b1 , w_8525 );
not ( w_8525 , w_8526 );
and ( \2711_b0 , \739_b0 , w_8527 );
and ( w_8526 ,  , w_8527 );
buf ( w_8525 , \2638_b1 );
not ( w_8525 , w_8528 );
not (  , w_8529 );
and ( w_8528 , w_8529 , \2638_b0 );
or ( \2712_b1 , \2710_b1 , w_8531 );
not ( w_8531 , w_8532 );
and ( \2712_b0 , \2710_b0 , w_8533 );
and ( w_8532 ,  , w_8533 );
buf ( w_8531 , \2711_b1 );
not ( w_8531 , w_8534 );
not (  , w_8535 );
and ( w_8534 , w_8535 , \2711_b0 );
or ( \2713_b1 , \2706_b1 , w_8537 );
not ( w_8537 , w_8538 );
and ( \2713_b0 , \2706_b0 , w_8539 );
and ( w_8538 ,  , w_8539 );
buf ( w_8537 , \2712_b1 );
not ( w_8537 , w_8540 );
not (  , w_8541 );
and ( w_8540 , w_8541 , \2712_b0 );
or ( \2714_b1 , \2699_b1 , w_8543 );
not ( w_8543 , w_8544 );
and ( \2714_b0 , \2699_b0 , w_8545 );
and ( w_8544 ,  , w_8545 );
buf ( w_8543 , \2705_b1 );
not ( w_8543 , w_8546 );
not (  , w_8547 );
and ( w_8546 , w_8547 , \2705_b0 );
or ( \2715_b1 , \2713_b1 , w_8549 );
not ( w_8549 , w_8550 );
and ( \2715_b0 , \2713_b0 , w_8551 );
and ( w_8550 ,  , w_8551 );
buf ( w_8549 , \2714_b1 );
not ( w_8549 , w_8552 );
not (  , w_8553 );
and ( w_8552 , w_8553 , \2714_b0 );
or ( \2716_b1 , \2693_b1 , w_8555 );
not ( w_8555 , w_8556 );
and ( \2716_b0 , \2693_b0 , w_8557 );
and ( w_8556 ,  , w_8557 );
buf ( w_8555 , \2715_b1 );
not ( w_8555 , w_8558 );
not (  , w_8559 );
and ( w_8558 , w_8559 , \2715_b0 );
or ( \2717_b1 , \2354_b1 , \2336_b1 );
xor ( \2717_b0 , \2354_b0 , w_8560 );
not ( w_8560 , w_8561 );
and ( w_8561 , \2336_b1 , \2336_b0 );
or ( \2718_b1 , \2717_b1 , w_8562 );
xor ( \2718_b0 , \2717_b0 , w_8564 );
not ( w_8564 , w_8565 );
and ( w_8565 , w_8562 , w_8563 );
buf ( w_8562 , \2344_b1 );
not ( w_8562 , w_8566 );
not ( w_8563 , w_8567 );
and ( w_8566 , w_8567 , \2344_b0 );
or ( \2719_b1 , \2716_b1 , w_8568 );
or ( \2719_b0 , \2716_b0 , \2718_b0 );
not ( \2718_b0 , w_8569 );
and ( w_8569 , w_8568 , \2718_b1 );
or ( \2720_b1 , \2693_b1 , w_8571 );
not ( w_8571 , w_8572 );
and ( \2720_b0 , \2693_b0 , w_8573 );
and ( w_8572 ,  , w_8573 );
buf ( w_8571 , \2715_b1 );
not ( w_8571 , w_8574 );
not (  , w_8575 );
and ( w_8574 , w_8575 , \2715_b0 );
or ( \2721_b1 , \2719_b1 , w_8577 );
not ( w_8577 , w_8578 );
and ( \2721_b0 , \2719_b0 , w_8579 );
and ( w_8578 ,  , w_8579 );
buf ( w_8577 , \2720_b1 );
not ( w_8577 , w_8580 );
not (  , w_8581 );
and ( w_8580 , w_8581 , \2720_b0 );
or ( \2722_b1 , \2676_b1 , w_8583 );
not ( w_8583 , w_8584 );
and ( \2722_b0 , \2676_b0 , w_8585 );
and ( w_8584 ,  , w_8585 );
buf ( w_8583 , \2721_b1 );
not ( w_8583 , w_8586 );
not (  , w_8587 );
and ( w_8586 , w_8587 , \2721_b0 );
buf ( \2723_b1 , \2671_b1 );
not ( \2723_b1 , w_8588 );
not ( \2723_b0 , w_8589 );
and ( w_8588 , w_8589 , \2671_b0 );
buf ( \2724_b1 , \2674_b1 );
not ( \2724_b1 , w_8590 );
not ( \2724_b0 , w_8591 );
and ( w_8590 , w_8591 , \2674_b0 );
or ( \2725_b1 , \2723_b1 , w_8593 );
not ( w_8593 , w_8594 );
and ( \2725_b0 , \2723_b0 , w_8595 );
and ( w_8594 ,  , w_8595 );
buf ( w_8593 , \2724_b1 );
not ( w_8593 , w_8596 );
not (  , w_8597 );
and ( w_8596 , w_8597 , \2724_b0 );
or ( \2726_b1 , \2722_b1 , w_8599 );
not ( w_8599 , w_8600 );
and ( \2726_b0 , \2722_b0 , w_8601 );
and ( w_8600 ,  , w_8601 );
buf ( w_8599 , \2725_b1 );
not ( w_8599 , w_8602 );
not (  , w_8603 );
and ( w_8602 , w_8603 , \2725_b0 );
buf ( \2727_b1 , \2726_b1 );
not ( \2727_b1 , w_8604 );
not ( \2727_b0 , w_8605 );
and ( w_8604 , w_8605 , \2726_b0 );
or ( \2728_b1 , \2669_b1 , w_8607 );
not ( w_8607 , w_8608 );
and ( \2728_b0 , \2669_b0 , w_8609 );
and ( w_8608 ,  , w_8609 );
buf ( w_8607 , \2727_b1 );
not ( w_8607 , w_8610 );
not (  , w_8611 );
and ( w_8610 , w_8611 , \2727_b0 );
buf ( \2729_b1 , \2644_b1 );
not ( \2729_b1 , w_8612 );
not ( \2729_b0 , w_8613 );
and ( w_8612 , w_8613 , \2644_b0 );
buf ( \2730_b1 , \2636_b1 );
not ( \2730_b1 , w_8614 );
not ( \2730_b0 , w_8615 );
and ( w_8614 , w_8615 , \2636_b0 );
or ( \2731_b1 , \2729_b1 , w_8616 );
or ( \2731_b0 , \2729_b0 , \2730_b0 );
not ( \2730_b0 , w_8617 );
and ( w_8617 , w_8616 , \2730_b1 );
buf ( \2732_b1 , \2636_b1 );
not ( \2732_b1 , w_8618 );
not ( \2732_b0 , w_8619 );
and ( w_8618 , w_8619 , \2636_b0 );
or ( \2733_b1 , \2732_b1 , w_8621 );
not ( w_8621 , w_8622 );
and ( \2733_b0 , \2732_b0 , w_8623 );
and ( w_8622 ,  , w_8623 );
buf ( w_8621 , \2643_b1 );
not ( w_8621 , w_8624 );
not (  , w_8625 );
and ( w_8624 , w_8625 , \2643_b0 );
or ( \2734_b1 , \2731_b1 , w_8627 );
not ( w_8627 , w_8628 );
and ( \2734_b0 , \2731_b0 , w_8629 );
and ( w_8628 ,  , w_8629 );
buf ( w_8627 , \2733_b1 );
not ( w_8627 , w_8630 );
not (  , w_8631 );
and ( w_8630 , w_8631 , \2733_b0 );
or ( \2735_b1 , \2734_b1 , w_8632 );
xor ( \2735_b0 , \2734_b0 , w_8634 );
not ( w_8634 , w_8635 );
and ( w_8635 , w_8632 , w_8633 );
buf ( w_8632 , \2650_b1 );
not ( w_8632 , w_8636 );
not ( w_8633 , w_8637 );
and ( w_8636 , w_8637 , \2650_b0 );
or ( \2736_b1 , \b[0]_b1 , w_8638 );
or ( \2736_b0 , \b[0]_b0 , \c[8]_b0 );
not ( \c[8]_b0 , w_8639 );
and ( w_8639 , w_8638 , \c[8]_b1 );
or ( \2737_b1 , \2736_b1 , w_8641 );
not ( w_8641 , w_8642 );
and ( \2737_b0 , \2736_b0 , w_8643 );
and ( w_8642 ,  , w_8643 );
buf ( w_8641 , \c[7]_b1 );
not ( w_8641 , w_8644 );
not (  , w_8645 );
and ( w_8644 , w_8645 , \c[7]_b0 );
or ( \2738_b1 , \b[0]_b1 , w_8647 );
not ( w_8647 , w_8648 );
and ( \2738_b0 , \b[0]_b0 , w_8649 );
and ( w_8648 ,  , w_8649 );
buf ( w_8647 , \c[8]_b1 );
not ( w_8647 , w_8650 );
not (  , w_8651 );
and ( w_8650 , w_8651 , \c[8]_b0 );
or ( \2740_b1 , \b[6]_b1 , \c[3]_b1 );
xor ( \2740_b0 , \b[6]_b0 , w_8652 );
not ( w_8652 , w_8653 );
and ( w_8653 , \c[3]_b1 , \c[3]_b0 );
buf ( \2741_b1 , \2740_b1 );
not ( \2741_b1 , w_8654 );
not ( \2741_b0 , w_8655 );
and ( w_8654 , w_8655 , \2740_b0 );
buf ( \2742_b1 , \699_b1 );
not ( \2742_b1 , w_8656 );
not ( \2742_b0 , w_8657 );
and ( w_8656 , w_8657 , \699_b0 );
or ( \2743_b1 , \2741_b1 , w_8658 );
or ( \2743_b0 , \2741_b0 , \2742_b0 );
not ( \2742_b0 , w_8659 );
and ( w_8659 , w_8658 , \2742_b1 );
or ( \2744_b1 , \702_b1 , w_8661 );
not ( w_8661 , w_8662 );
and ( \2744_b0 , \702_b0 , w_8663 );
and ( w_8662 ,  , w_8663 );
buf ( w_8661 , \2685_b1 );
not ( w_8661 , w_8664 );
not (  , w_8665 );
and ( w_8664 , w_8665 , \2685_b0 );
or ( \2745_b1 , \2743_b1 , w_8667 );
not ( w_8667 , w_8668 );
and ( \2745_b0 , \2743_b0 , w_8669 );
and ( w_8668 ,  , w_8669 );
buf ( w_8667 , \2744_b1 );
not ( w_8667 , w_8670 );
not (  , w_8671 );
and ( w_8670 , w_8671 , \2744_b0 );
or ( \2746_b1 , \2739_b1 , \2745_b1 );
not ( \2745_b1 , w_8672 );
and ( \2746_b0 , \2739_b0 , w_8673 );
and ( w_8672 , w_8673 , \2745_b0 );
or ( \2747_b1 , \2677_b1 , \2683_b1 );
xor ( \2747_b0 , \2677_b0 , w_8674 );
not ( w_8674 , w_8675 );
and ( w_8675 , \2683_b1 , \2683_b0 );
or ( \2748_b1 , \2747_b1 , \2690_b1 );
xor ( \2748_b0 , \2747_b0 , w_8676 );
not ( w_8676 , w_8677 );
and ( w_8677 , \2690_b1 , \2690_b0 );
or ( \2749_b1 , \2746_b1 , \2748_b1 );
xor ( \2749_b0 , \2746_b0 , w_8678 );
not ( w_8678 , w_8679 );
and ( w_8679 , \2748_b1 , \2748_b0 );
or ( \2750_b1 , \c[9]_b1 , \b[0]_b1 );
xor ( \2750_b0 , \c[9]_b0 , w_8680 );
not ( w_8680 , w_8681 );
and ( w_8681 , \b[0]_b1 , \b[0]_b0 );
buf ( \2751_b1 , \2750_b1 );
not ( \2751_b1 , w_8682 );
not ( \2751_b0 , w_8683 );
and ( w_8682 , w_8683 , \2750_b0 );
buf ( \2752_b1 , \2281_b1 );
not ( \2752_b1 , w_8684 );
not ( \2752_b0 , w_8685 );
and ( w_8684 , w_8685 , \2281_b0 );
or ( \2753_b1 , \2751_b1 , w_8686 );
or ( \2753_b0 , \2751_b0 , \2752_b0 );
not ( \2752_b0 , w_8687 );
and ( w_8687 , w_8686 , \2752_b1 );
or ( \2754_b1 , \2284_b1 , w_8689 );
not ( w_8689 , w_8690 );
and ( \2754_b0 , \2284_b0 , w_8691 );
and ( w_8690 ,  , w_8691 );
buf ( w_8689 , \2694_b1 );
not ( w_8689 , w_8692 );
not (  , w_8693 );
and ( w_8692 , w_8693 , \2694_b0 );
or ( \2755_b1 , \2753_b1 , w_8695 );
not ( w_8695 , w_8696 );
and ( \2755_b0 , \2753_b0 , w_8697 );
and ( w_8696 ,  , w_8697 );
buf ( w_8695 , \2754_b1 );
not ( w_8695 , w_8698 );
not (  , w_8699 );
and ( w_8698 , w_8699 , \2754_b0 );
or ( \2756_b1 , \c[1]_b1 , \b[8]_b1 );
xor ( \2756_b0 , \c[1]_b0 , w_8700 );
not ( w_8700 , w_8701 );
and ( w_8701 , \b[8]_b1 , \b[8]_b0 );
buf ( \2757_b1 , \2756_b1 );
not ( \2757_b1 , w_8702 );
not ( \2757_b0 , w_8703 );
and ( w_8702 , w_8703 , \2756_b0 );
buf ( \2758_b1 , \679_b1 );
not ( \2758_b1 , w_8704 );
not ( \2758_b0 , w_8705 );
and ( w_8704 , w_8705 , \679_b0 );
or ( \2759_b1 , \2757_b1 , w_8706 );
or ( \2759_b0 , \2757_b0 , \2758_b0 );
not ( \2758_b0 , w_8707 );
and ( w_8707 , w_8706 , \2758_b1 );
or ( \2760_b1 , \2700_b1 , w_8709 );
not ( w_8709 , w_8710 );
and ( \2760_b0 , \2700_b0 , w_8711 );
and ( w_8710 ,  , w_8711 );
buf ( w_8709 , \c[0]_b1 );
not ( w_8709 , w_8712 );
not (  , w_8713 );
and ( w_8712 , w_8713 , \c[0]_b0 );
or ( \2761_b1 , \2759_b1 , w_8715 );
not ( w_8715 , w_8716 );
and ( \2761_b0 , \2759_b0 , w_8717 );
and ( w_8716 ,  , w_8717 );
buf ( w_8715 , \2760_b1 );
not ( w_8715 , w_8718 );
not (  , w_8719 );
and ( w_8718 , w_8719 , \2760_b0 );
or ( \2762_b1 , \2755_b1 , w_8720 );
or ( \2762_b0 , \2755_b0 , \2761_b0 );
not ( \2761_b0 , w_8721 );
and ( w_8721 , w_8720 , \2761_b1 );
or ( \2763_b1 , \b[2]_b1 , \c[7]_b1 );
xor ( \2763_b0 , \b[2]_b0 , w_8722 );
not ( w_8722 , w_8723 );
and ( w_8723 , \c[7]_b1 , \c[7]_b0 );
buf ( \2764_b1 , \2763_b1 );
not ( \2764_b1 , w_8724 );
not ( \2764_b0 , w_8725 );
and ( w_8724 , w_8725 , \2763_b0 );
buf ( \2765_b1 , \726_b1 );
not ( \2765_b1 , w_8726 );
not ( \2765_b0 , w_8727 );
and ( w_8726 , w_8727 , \726_b0 );
or ( \2766_b1 , \2764_b1 , w_8728 );
or ( \2766_b0 , \2764_b0 , \2765_b0 );
not ( \2765_b0 , w_8729 );
and ( w_8729 , w_8728 , \2765_b1 );
or ( \2767_b1 , \714_b1 , w_8731 );
not ( w_8731 , w_8732 );
and ( \2767_b0 , \714_b0 , w_8733 );
and ( w_8732 ,  , w_8733 );
buf ( w_8731 , \2678_b1 );
not ( w_8731 , w_8734 );
not (  , w_8735 );
and ( w_8734 , w_8735 , \2678_b0 );
or ( \2768_b1 , \2766_b1 , w_8737 );
not ( w_8737 , w_8738 );
and ( \2768_b0 , \2766_b0 , w_8739 );
and ( w_8738 ,  , w_8739 );
buf ( w_8737 , \2767_b1 );
not ( w_8737 , w_8740 );
not (  , w_8741 );
and ( w_8740 , w_8741 , \2767_b0 );
or ( \2769_b1 , \2762_b1 , w_8743 );
not ( w_8743 , w_8744 );
and ( \2769_b0 , \2762_b0 , w_8745 );
and ( w_8744 ,  , w_8745 );
buf ( w_8743 , \2768_b1 );
not ( w_8743 , w_8746 );
not (  , w_8747 );
and ( w_8746 , w_8747 , \2768_b0 );
or ( \2770_b1 , \2755_b1 , w_8749 );
not ( w_8749 , w_8750 );
and ( \2770_b0 , \2755_b0 , w_8751 );
and ( w_8750 ,  , w_8751 );
buf ( w_8749 , \2761_b1 );
not ( w_8749 , w_8752 );
not (  , w_8753 );
and ( w_8752 , w_8753 , \2761_b0 );
or ( \2771_b1 , \2769_b1 , w_8755 );
not ( w_8755 , w_8756 );
and ( \2771_b0 , \2769_b0 , w_8757 );
and ( w_8756 ,  , w_8757 );
buf ( w_8755 , \2770_b1 );
not ( w_8755 , w_8758 );
not (  , w_8759 );
and ( w_8758 , w_8759 , \2770_b0 );
or ( \2772_b1 , \2749_b1 , \2771_b1 );
not ( \2771_b1 , w_8760 );
and ( \2772_b0 , \2749_b0 , w_8761 );
and ( w_8760 , w_8761 , \2771_b0 );
or ( \2773_b1 , \2746_b1 , \2748_b1 );
not ( \2748_b1 , w_8762 );
and ( \2773_b0 , \2746_b0 , w_8763 );
and ( w_8762 , w_8763 , \2748_b0 );
or ( \2774_b1 , \2772_b1 , w_8764 );
or ( \2774_b0 , \2772_b0 , \2773_b0 );
not ( \2773_b0 , w_8765 );
and ( w_8765 , w_8764 , \2773_b1 );
buf ( \2775_b1 , \2774_b1 );
not ( \2775_b1 , w_8766 );
not ( \2775_b0 , w_8767 );
and ( w_8766 , w_8767 , \2774_b0 );
or ( \2776_b1 , \2735_b1 , \2775_b1 );
xor ( \2776_b0 , \2735_b0 , w_8768 );
not ( w_8768 , w_8769 );
and ( w_8769 , \2775_b1 , \2775_b0 );
or ( \2777_b1 , \2715_b1 , \2693_b1 );
xor ( \2777_b0 , \2715_b0 , w_8770 );
not ( w_8770 , w_8771 );
and ( w_8771 , \2693_b1 , \2693_b0 );
or ( \2778_b1 , \2777_b1 , \2718_b1 );
xor ( \2778_b0 , \2777_b0 , w_8772 );
not ( w_8772 , w_8773 );
and ( w_8773 , \2718_b1 , \2718_b0 );
or ( \2779_b1 , \2776_b1 , \2778_b1 );
xor ( \2779_b0 , \2776_b0 , w_8774 );
not ( w_8774 , w_8775 );
and ( w_8775 , \2778_b1 , \2778_b0 );
or ( \2780_b1 , \2705_b1 , \2699_b1 );
xor ( \2780_b0 , \2705_b0 , w_8776 );
not ( w_8776 , w_8777 );
and ( w_8777 , \2699_b1 , \2699_b0 );
or ( \2781_b1 , \2780_b1 , \2712_b1 );
xor ( \2781_b0 , \2780_b0 , w_8778 );
not ( w_8778 , w_8779 );
and ( w_8779 , \2712_b1 , \2712_b0 );
or ( \2782_b1 , \2746_b1 , \2748_b1 );
xor ( \2782_b0 , \2746_b0 , w_8780 );
not ( w_8780 , w_8781 );
and ( w_8781 , \2748_b1 , \2748_b0 );
or ( \2783_b1 , \2782_b1 , \2771_b1 );
xor ( \2783_b0 , \2782_b0 , w_8782 );
not ( w_8782 , w_8783 );
and ( w_8783 , \2771_b1 , \2771_b0 );
or ( \2784_b1 , \2781_b1 , w_8784 );
or ( \2784_b0 , \2781_b0 , \2783_b0 );
not ( \2783_b0 , w_8785 );
and ( w_8785 , w_8784 , \2783_b1 );
or ( \2785_b1 , \b[4]_b1 , \c[5]_b1 );
xor ( \2785_b0 , \b[4]_b0 , w_8786 );
not ( w_8786 , w_8787 );
and ( w_8787 , \c[5]_b1 , \c[5]_b0 );
buf ( \2786_b1 , \2785_b1 );
not ( \2786_b1 , w_8788 );
not ( \2786_b0 , w_8789 );
and ( w_8788 , w_8789 , \2785_b0 );
buf ( \2787_b1 , \2265_b1 );
not ( \2787_b1 , w_8790 );
not ( \2787_b0 , w_8791 );
and ( w_8790 , w_8791 , \2265_b0 );
or ( \2788_b1 , \2786_b1 , w_8792 );
or ( \2788_b0 , \2786_b0 , \2787_b0 );
not ( \2787_b0 , w_8793 );
and ( w_8793 , w_8792 , \2787_b1 );
or ( \2789_b1 , \739_b1 , w_8795 );
not ( w_8795 , w_8796 );
and ( \2789_b0 , \739_b0 , w_8797 );
and ( w_8796 ,  , w_8797 );
buf ( w_8795 , \2707_b1 );
not ( w_8795 , w_8798 );
not (  , w_8799 );
and ( w_8798 , w_8799 , \2707_b0 );
or ( \2790_b1 , \2788_b1 , w_8801 );
not ( w_8801 , w_8802 );
and ( \2790_b0 , \2788_b0 , w_8803 );
and ( w_8802 ,  , w_8803 );
buf ( w_8801 , \2789_b1 );
not ( w_8801 , w_8804 );
not (  , w_8805 );
and ( w_8804 , w_8805 , \2789_b0 );
or ( \2791_b1 , \2739_b1 , \2745_b1 );
xor ( \2791_b0 , \2739_b0 , w_8806 );
not ( w_8806 , w_8807 );
and ( w_8807 , \2745_b1 , \2745_b0 );
or ( \2792_b1 , \2790_b1 , \2791_b1 );
xor ( \2792_b0 , \2790_b0 , w_8808 );
not ( w_8808 , w_8809 );
and ( w_8809 , \2791_b1 , \2791_b0 );
buf ( \2793_b1 , \682_b1 );
not ( \2793_b1 , w_8810 );
not ( \2793_b0 , w_8811 );
and ( w_8810 , w_8811 , \682_b0 );
buf ( \2794_b1 , \679_b1 );
not ( \2794_b1 , w_8812 );
not ( \2794_b0 , w_8813 );
and ( w_8812 , w_8813 , \679_b0 );
or ( \2795_b1 , \2793_b1 , w_8814 );
or ( \2795_b0 , \2793_b0 , \2794_b0 );
not ( \2794_b0 , w_8815 );
and ( w_8815 , w_8814 , \2794_b1 );
or ( \2796_b1 , \2756_b1 , w_8817 );
not ( w_8817 , w_8818 );
and ( \2796_b0 , \2756_b0 , w_8819 );
and ( w_8818 ,  , w_8819 );
buf ( w_8817 , \c[0]_b1 );
not ( w_8817 , w_8820 );
not (  , w_8821 );
and ( w_8820 , w_8821 , \c[0]_b0 );
or ( \2797_b1 , \2795_b1 , w_8823 );
not ( w_8823 , w_8824 );
and ( \2797_b0 , \2795_b0 , w_8825 );
and ( w_8824 ,  , w_8825 );
buf ( w_8823 , \2796_b1 );
not ( w_8823 , w_8826 );
not (  , w_8827 );
and ( w_8826 , w_8827 , \2796_b0 );
or ( \2798_b1 , \2280_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_8828 );
and ( \2798_b0 , \2280_b0 , w_8829 );
and ( w_8828 , w_8829 , \b[0]_b0 );
or ( \2799_b1 , \2797_b1 , w_8830 );
or ( \2799_b0 , \2797_b0 , \2798_b0 );
not ( \2798_b0 , w_8831 );
and ( w_8831 , w_8830 , \2798_b1 );
buf ( \2800_b1 , \729_b1 );
not ( \2800_b1 , w_8832 );
not ( \2800_b0 , w_8833 );
and ( w_8832 , w_8833 , \729_b0 );
buf ( \2801_b1 , \2292_b1 );
not ( \2801_b1 , w_8834 );
not ( \2801_b0 , w_8835 );
and ( w_8834 , w_8835 , \2292_b0 );
or ( \2802_b1 , \2800_b1 , w_8836 );
or ( \2802_b0 , \2800_b0 , \2801_b0 );
not ( \2801_b0 , w_8837 );
and ( w_8837 , w_8836 , \2801_b1 );
or ( \2803_b1 , \714_b1 , w_8839 );
not ( w_8839 , w_8840 );
and ( \2803_b0 , \714_b0 , w_8841 );
and ( w_8840 ,  , w_8841 );
buf ( w_8839 , \2763_b1 );
not ( w_8839 , w_8842 );
not (  , w_8843 );
and ( w_8842 , w_8843 , \2763_b0 );
or ( \2804_b1 , \2802_b1 , w_8845 );
not ( w_8845 , w_8846 );
and ( \2804_b0 , \2802_b0 , w_8847 );
and ( w_8846 ,  , w_8847 );
buf ( w_8845 , \2803_b1 );
not ( w_8845 , w_8848 );
not (  , w_8849 );
and ( w_8848 , w_8849 , \2803_b0 );
or ( \2805_b1 , \2799_b1 , w_8851 );
not ( w_8851 , w_8852 );
and ( \2805_b0 , \2799_b0 , w_8853 );
and ( w_8852 ,  , w_8853 );
buf ( w_8851 , \2804_b1 );
not ( w_8851 , w_8854 );
not (  , w_8855 );
and ( w_8854 , w_8855 , \2804_b0 );
or ( \2806_b1 , \2797_b1 , w_8857 );
not ( w_8857 , w_8858 );
and ( \2806_b0 , \2797_b0 , w_8859 );
and ( w_8858 ,  , w_8859 );
buf ( w_8857 , \2798_b1 );
not ( w_8857 , w_8860 );
not (  , w_8861 );
and ( w_8860 , w_8861 , \2798_b0 );
or ( \2807_b1 , \2805_b1 , w_8863 );
not ( w_8863 , w_8864 );
and ( \2807_b0 , \2805_b0 , w_8865 );
and ( w_8864 ,  , w_8865 );
buf ( w_8863 , \2806_b1 );
not ( w_8863 , w_8866 );
not (  , w_8867 );
and ( w_8866 , w_8867 , \2806_b0 );
or ( \2808_b1 , \2792_b1 , \2807_b1 );
not ( \2807_b1 , w_8868 );
and ( \2808_b0 , \2792_b0 , w_8869 );
and ( w_8868 , w_8869 , \2807_b0 );
or ( \2809_b1 , \2790_b1 , \2791_b1 );
not ( \2791_b1 , w_8870 );
and ( \2809_b0 , \2790_b0 , w_8871 );
and ( w_8870 , w_8871 , \2791_b0 );
or ( \2810_b1 , \2808_b1 , w_8872 );
or ( \2810_b0 , \2808_b0 , \2809_b0 );
not ( \2809_b0 , w_8873 );
and ( w_8873 , w_8872 , \2809_b1 );
or ( \2811_b1 , \2784_b1 , w_8875 );
not ( w_8875 , w_8876 );
and ( \2811_b0 , \2784_b0 , w_8877 );
and ( w_8876 ,  , w_8877 );
buf ( w_8875 , \2810_b1 );
not ( w_8875 , w_8878 );
not (  , w_8879 );
and ( w_8878 , w_8879 , \2810_b0 );
or ( \2812_b1 , \2783_b1 , w_8881 );
not ( w_8881 , w_8882 );
and ( \2812_b0 , \2783_b0 , w_8883 );
and ( w_8882 ,  , w_8883 );
buf ( w_8881 , \2781_b1 );
not ( w_8881 , w_8884 );
not (  , w_8885 );
and ( w_8884 , w_8885 , \2781_b0 );
or ( \2813_b1 , \2811_b1 , \2812_b1 );
not ( \2812_b1 , w_8886 );
and ( \2813_b0 , \2811_b0 , w_8887 );
and ( w_8886 , w_8887 , \2812_b0 );
or ( \2814_b1 , \2779_b1 , w_8889 );
not ( w_8889 , w_8890 );
and ( \2814_b0 , \2779_b0 , w_8891 );
and ( w_8890 ,  , w_8891 );
buf ( w_8889 , \2813_b1 );
not ( w_8889 , w_8892 );
not (  , w_8893 );
and ( w_8892 , w_8893 , \2813_b0 );
or ( \2815_b1 , \2728_b1 , w_8895 );
not ( w_8895 , w_8896 );
and ( \2815_b0 , \2728_b0 , w_8897 );
and ( w_8896 ,  , w_8897 );
buf ( w_8895 , \2814_b1 );
not ( w_8895 , w_8898 );
not (  , w_8899 );
and ( w_8898 , w_8899 , \2814_b0 );
or ( \2816_b1 , \2660_b1 , w_8901 );
not ( w_8901 , w_8902 );
and ( \2816_b0 , \2660_b0 , w_8903 );
and ( w_8902 ,  , w_8903 );
buf ( w_8901 , \2815_b1 );
not ( w_8901 , w_8904 );
not (  , w_8905 );
and ( w_8904 , w_8905 , \2815_b0 );
buf ( \2817_b1 , \2816_b1 );
not ( \2817_b1 , w_8906 );
not ( \2817_b0 , w_8907 );
and ( w_8906 , w_8907 , \2816_b0 );
buf ( \2818_b1 , \2721_b1 );
not ( \2818_b1 , w_8908 );
not ( \2818_b0 , w_8909 );
and ( w_8908 , w_8909 , \2721_b0 );
buf ( \2819_b1 , \2671_b1 );
not ( \2819_b1 , w_8910 );
not ( \2819_b0 , w_8911 );
and ( w_8910 , w_8911 , \2671_b0 );
or ( \2820_b1 , \2818_b1 , w_8912 );
or ( \2820_b0 , \2818_b0 , \2819_b0 );
not ( \2819_b0 , w_8913 );
and ( w_8913 , w_8912 , \2819_b1 );
or ( \2821_b1 , \2671_b1 , w_8914 );
or ( \2821_b0 , \2671_b0 , \2721_b0 );
not ( \2721_b0 , w_8915 );
and ( w_8915 , w_8914 , \2721_b1 );
or ( \2822_b1 , \2820_b1 , w_8917 );
not ( w_8917 , w_8918 );
and ( \2822_b0 , \2820_b0 , w_8919 );
and ( w_8918 ,  , w_8919 );
buf ( w_8917 , \2821_b1 );
not ( w_8917 , w_8920 );
not (  , w_8921 );
and ( w_8920 , w_8921 , \2821_b0 );
or ( \2823_b1 , \2822_b1 , \2674_b1 );
not ( \2674_b1 , w_8922 );
and ( \2823_b0 , \2822_b0 , w_8923 );
and ( w_8922 , w_8923 , \2674_b0 );
buf ( \2824_b1 , \2822_b1 );
not ( \2824_b1 , w_8924 );
not ( \2824_b0 , w_8925 );
and ( w_8924 , w_8925 , \2822_b0 );
or ( \2825_b1 , \2824_b1 , \2724_b1 );
not ( \2724_b1 , w_8926 );
and ( \2825_b0 , \2824_b0 , w_8927 );
and ( w_8926 , w_8927 , \2724_b0 );
or ( \2826_b1 , \2823_b1 , w_8929 );
not ( w_8929 , w_8930 );
and ( \2826_b0 , \2823_b0 , w_8931 );
and ( w_8930 ,  , w_8931 );
buf ( w_8929 , \2825_b1 );
not ( w_8929 , w_8932 );
not (  , w_8933 );
and ( w_8932 , w_8933 , \2825_b0 );
or ( \2827_b1 , \2735_b1 , \2775_b1 );
xor ( \2827_b0 , \2735_b0 , w_8934 );
not ( w_8934 , w_8935 );
and ( w_8935 , \2775_b1 , \2775_b0 );
or ( \2828_b1 , \2827_b1 , \2778_b1 );
not ( \2778_b1 , w_8936 );
and ( \2828_b0 , \2827_b0 , w_8937 );
and ( w_8936 , w_8937 , \2778_b0 );
or ( \2829_b1 , \2735_b1 , \2775_b1 );
not ( \2775_b1 , w_8938 );
and ( \2829_b0 , \2735_b0 , w_8939 );
and ( w_8938 , w_8939 , \2775_b0 );
or ( \2830_b1 , \2828_b1 , w_8940 );
or ( \2830_b0 , \2828_b0 , \2829_b0 );
not ( \2829_b0 , w_8941 );
and ( w_8941 , w_8940 , \2829_b1 );
or ( \2831_b1 , \2826_b1 , w_8943 );
not ( w_8943 , w_8944 );
and ( \2831_b0 , \2826_b0 , w_8945 );
and ( w_8944 ,  , w_8945 );
buf ( w_8943 , \2830_b1 );
not ( w_8943 , w_8946 );
not (  , w_8947 );
and ( w_8946 , w_8947 , \2830_b0 );
or ( \2832_b1 , \2781_b1 , \2810_b1 );
xor ( \2832_b0 , \2781_b0 , w_8948 );
not ( w_8948 , w_8949 );
and ( w_8949 , \2810_b1 , \2810_b0 );
or ( \2833_b1 , \2832_b1 , w_8950 );
xor ( \2833_b0 , \2832_b0 , w_8952 );
not ( w_8952 , w_8953 );
and ( w_8953 , w_8950 , w_8951 );
buf ( w_8950 , \2783_b1 );
not ( w_8950 , w_8954 );
not ( w_8951 , w_8955 );
and ( w_8954 , w_8955 , \2783_b0 );
buf ( \2834_b1 , \740_b1 );
not ( \2834_b1 , w_8956 );
not ( \2834_b0 , w_8957 );
and ( w_8956 , w_8957 , \740_b0 );
buf ( \2835_b1 , \736_b1 );
not ( \2835_b1 , w_8958 );
not ( \2835_b0 , w_8959 );
and ( w_8958 , w_8959 , \736_b0 );
or ( \2836_b1 , \2834_b1 , w_8960 );
or ( \2836_b0 , \2834_b0 , \2835_b0 );
not ( \2835_b0 , w_8961 );
and ( w_8961 , w_8960 , \2835_b1 );
or ( \2837_b1 , \739_b1 , w_8963 );
not ( w_8963 , w_8964 );
and ( \2837_b0 , \739_b0 , w_8965 );
and ( w_8964 ,  , w_8965 );
buf ( w_8963 , \2785_b1 );
not ( w_8963 , w_8966 );
not (  , w_8967 );
and ( w_8966 , w_8967 , \2785_b0 );
or ( \2838_b1 , \2836_b1 , w_8969 );
not ( w_8969 , w_8970 );
and ( \2838_b0 , \2836_b0 , w_8971 );
and ( w_8970 ,  , w_8971 );
buf ( w_8969 , \2837_b1 );
not ( w_8969 , w_8972 );
not (  , w_8973 );
and ( w_8972 , w_8973 , \2837_b0 );
buf ( \2839_b1 , \2838_b1 );
not ( \2839_b1 , w_8974 );
not ( \2839_b0 , w_8975 );
and ( w_8974 , w_8975 , \2838_b0 );
buf ( \2840_b1 , \2839_b1 );
not ( \2840_b1 , w_8976 );
not ( \2840_b0 , w_8977 );
and ( w_8976 , w_8977 , \2839_b0 );
buf ( \2841_b1 , \689_b1 );
not ( \2841_b1 , w_8978 );
not ( \2841_b0 , w_8979 );
and ( w_8978 , w_8979 , \689_b0 );
or ( \2842_b1 , \2841_b1 , w_8981 );
not ( w_8981 , w_8982 );
and ( \2842_b0 , \2841_b0 , w_8983 );
and ( w_8982 ,  , w_8983 );
buf ( w_8981 , \684_b1 );
not ( w_8981 , w_8984 );
not (  , w_8985 );
and ( w_8984 , w_8985 , \684_b0 );
buf ( \2843_b1 , \2842_b1 );
not ( \2843_b1 , w_8986 );
not ( \2843_b0 , w_8987 );
and ( w_8986 , w_8987 , \2842_b0 );
or ( \2844_b1 , \2840_b1 , w_8988 );
or ( \2844_b0 , \2840_b0 , \2843_b0 );
not ( \2843_b0 , w_8989 );
and ( w_8989 , w_8988 , \2843_b1 );
buf ( \2845_b1 , \749_b1 );
not ( \2845_b1 , w_8990 );
not ( \2845_b0 , w_8991 );
and ( w_8990 , w_8991 , \749_b0 );
buf ( \2846_b1 , \746_b1 );
not ( \2846_b1 , w_8992 );
not ( \2846_b0 , w_8993 );
and ( w_8992 , w_8993 , \746_b0 );
or ( \2847_b1 , \2845_b1 , w_8994 );
or ( \2847_b0 , \2845_b0 , \2846_b0 );
not ( \2846_b0 , w_8995 );
and ( w_8995 , w_8994 , \2846_b1 );
or ( \2848_b1 , \702_b1 , w_8997 );
not ( w_8997 , w_8998 );
and ( \2848_b0 , \702_b0 , w_8999 );
and ( w_8998 ,  , w_8999 );
buf ( w_8997 , \2740_b1 );
not ( w_8997 , w_9000 );
not (  , w_9001 );
and ( w_9000 , w_9001 , \2740_b0 );
or ( \2849_b1 , \2847_b1 , w_9003 );
not ( w_9003 , w_9004 );
and ( \2849_b0 , \2847_b0 , w_9005 );
and ( w_9004 ,  , w_9005 );
buf ( w_9003 , \2848_b1 );
not ( w_9003 , w_9006 );
not (  , w_9007 );
and ( w_9006 , w_9007 , \2848_b0 );
or ( \2850_b1 , \2844_b1 , w_9009 );
not ( w_9009 , w_9010 );
and ( \2850_b0 , \2844_b0 , w_9011 );
and ( w_9010 ,  , w_9011 );
buf ( w_9009 , \2849_b1 );
not ( w_9009 , w_9012 );
not (  , w_9013 );
and ( w_9012 , w_9013 , \2849_b0 );
buf ( \2851_b1 , \2842_b1 );
not ( \2851_b1 , w_9014 );
not ( \2851_b0 , w_9015 );
and ( w_9014 , w_9015 , \2842_b0 );
or ( \2852_b1 , \2851_b1 , w_9017 );
not ( w_9017 , w_9018 );
and ( \2852_b0 , \2851_b0 , w_9019 );
and ( w_9018 ,  , w_9019 );
buf ( w_9017 , \2838_b1 );
not ( w_9017 , w_9020 );
not (  , w_9021 );
and ( w_9020 , w_9021 , \2838_b0 );
or ( \2853_b1 , \2850_b1 , w_9023 );
not ( w_9023 , w_9024 );
and ( \2853_b0 , \2850_b0 , w_9025 );
and ( w_9024 ,  , w_9025 );
buf ( w_9023 , \2852_b1 );
not ( w_9023 , w_9026 );
not (  , w_9027 );
and ( w_9026 , w_9027 , \2852_b0 );
buf ( \2854_b1 , \2853_b1 );
not ( \2854_b1 , w_9028 );
not ( \2854_b0 , w_9029 );
and ( w_9028 , w_9029 , \2853_b0 );
buf ( \2855_b1 , \2854_b1 );
not ( \2855_b1 , w_9030 );
not ( \2855_b0 , w_9031 );
and ( w_9030 , w_9031 , \2854_b0 );
or ( \2856_b1 , \2761_b1 , \2768_b1 );
xor ( \2856_b0 , \2761_b0 , w_9032 );
not ( w_9032 , w_9033 );
and ( w_9033 , \2768_b1 , \2768_b0 );
or ( \2857_b1 , \2856_b1 , w_9034 );
xor ( \2857_b0 , \2856_b0 , w_9036 );
not ( w_9036 , w_9037 );
and ( w_9037 , w_9034 , w_9035 );
buf ( w_9034 , \2755_b1 );
not ( w_9034 , w_9038 );
not ( w_9035 , w_9039 );
and ( w_9038 , w_9039 , \2755_b0 );
buf ( \2858_b1 , \2857_b1 );
not ( \2858_b1 , w_9040 );
not ( \2858_b0 , w_9041 );
and ( w_9040 , w_9041 , \2857_b0 );
or ( \2859_b1 , \2855_b1 , w_9042 );
or ( \2859_b0 , \2855_b0 , \2858_b0 );
not ( \2858_b0 , w_9043 );
and ( w_9043 , w_9042 , \2858_b1 );
or ( \2860_b1 , \2790_b1 , \2791_b1 );
xor ( \2860_b0 , \2790_b0 , w_9044 );
not ( w_9044 , w_9045 );
and ( w_9045 , \2791_b1 , \2791_b0 );
or ( \2861_b1 , \2860_b1 , \2807_b1 );
xor ( \2861_b0 , \2860_b0 , w_9046 );
not ( w_9046 , w_9047 );
and ( w_9047 , \2807_b1 , \2807_b0 );
or ( \2862_b1 , \2859_b1 , w_9049 );
not ( w_9049 , w_9050 );
and ( \2862_b0 , \2859_b0 , w_9051 );
and ( w_9050 ,  , w_9051 );
buf ( w_9049 , \2861_b1 );
not ( w_9049 , w_9052 );
not (  , w_9053 );
and ( w_9052 , w_9053 , \2861_b0 );
buf ( \2863_b1 , \2857_b1 );
not ( \2863_b1 , w_9054 );
not ( \2863_b0 , w_9055 );
and ( w_9054 , w_9055 , \2857_b0 );
or ( \2864_b1 , \2863_b1 , w_9057 );
not ( w_9057 , w_9058 );
and ( \2864_b0 , \2863_b0 , w_9059 );
and ( w_9058 ,  , w_9059 );
buf ( w_9057 , \2853_b1 );
not ( w_9057 , w_9060 );
not (  , w_9061 );
and ( w_9060 , w_9061 , \2853_b0 );
or ( \2865_b1 , \2862_b1 , \2864_b1 );
not ( \2864_b1 , w_9062 );
and ( \2865_b0 , \2862_b0 , w_9063 );
and ( w_9062 , w_9063 , \2864_b0 );
or ( \2866_b1 , \2833_b1 , w_9065 );
not ( w_9065 , w_9066 );
and ( \2866_b0 , \2833_b0 , w_9067 );
and ( w_9066 ,  , w_9067 );
buf ( w_9065 , \2865_b1 );
not ( w_9065 , w_9068 );
not (  , w_9069 );
and ( w_9068 , w_9069 , \2865_b0 );
or ( \2867_b1 , \2831_b1 , \2866_b1 );
not ( \2866_b1 , w_9070 );
and ( \2867_b0 , \2831_b0 , w_9071 );
and ( w_9070 , w_9071 , \2866_b0 );
buf ( \2868_b1 , \2867_b1 );
not ( \2868_b1 , w_9072 );
not ( \2868_b0 , w_9073 );
and ( w_9072 , w_9073 , \2867_b0 );
or ( \2869_b1 , \903_b1 , w_9075 );
not ( w_9075 , w_9076 );
and ( \2869_b0 , \903_b0 , w_9077 );
and ( w_9076 ,  , w_9077 );
buf ( w_9075 , \783_b1 );
not ( w_9075 , w_9078 );
not (  , w_9079 );
and ( w_9078 , w_9079 , \783_b0 );
or ( \2870_b1 , \2854_b1 , \2863_b1 );
not ( \2863_b1 , w_9080 );
and ( \2870_b0 , \2854_b0 , w_9081 );
and ( w_9080 , w_9081 , \2863_b0 );
buf ( \2871_b1 , \2854_b1 );
not ( \2871_b1 , w_9082 );
not ( \2871_b0 , w_9083 );
and ( w_9082 , w_9083 , \2854_b0 );
or ( \2872_b1 , \2871_b1 , \2857_b1 );
not ( \2857_b1 , w_9084 );
and ( \2872_b0 , \2871_b0 , w_9085 );
and ( w_9084 , w_9085 , \2857_b0 );
or ( \2873_b1 , \2870_b1 , w_9087 );
not ( w_9087 , w_9088 );
and ( \2873_b0 , \2870_b0 , w_9089 );
and ( w_9088 ,  , w_9089 );
buf ( w_9087 , \2872_b1 );
not ( w_9087 , w_9090 );
not (  , w_9091 );
and ( w_9090 , w_9091 , \2872_b0 );
buf ( \2874_b1 , \2873_b1 );
not ( \2874_b1 , w_9092 );
not ( \2874_b0 , w_9093 );
and ( w_9092 , w_9093 , \2873_b0 );
buf ( \2875_b1 , \2861_b1 );
not ( \2875_b1 , w_9094 );
not ( \2875_b0 , w_9095 );
and ( w_9094 , w_9095 , \2861_b0 );
or ( \2876_b1 , \2874_b1 , \2875_b1 );
not ( \2875_b1 , w_9096 );
and ( \2876_b0 , \2874_b0 , w_9097 );
and ( w_9096 , w_9097 , \2875_b0 );
or ( \2877_b1 , \2861_b1 , \2873_b1 );
not ( \2873_b1 , w_9098 );
and ( \2877_b0 , \2861_b0 , w_9099 );
and ( w_9098 , w_9099 , \2873_b0 );
or ( \2878_b1 , \2876_b1 , w_9101 );
not ( w_9101 , w_9102 );
and ( \2878_b0 , \2876_b0 , w_9103 );
and ( w_9102 ,  , w_9103 );
buf ( w_9101 , \2877_b1 );
not ( w_9101 , w_9104 );
not (  , w_9105 );
and ( w_9104 , w_9105 , \2877_b0 );
or ( \2879_b1 , \2798_b1 , \2797_b1 );
xor ( \2879_b0 , \2798_b0 , w_9106 );
not ( w_9106 , w_9107 );
and ( w_9107 , \2797_b1 , \2797_b0 );
or ( \2880_b1 , \2879_b1 , w_9108 );
xor ( \2880_b0 , \2879_b0 , w_9110 );
not ( w_9110 , w_9111 );
and ( w_9111 , w_9108 , w_9109 );
buf ( w_9108 , \2804_b1 );
not ( w_9108 , w_9112 );
not ( w_9109 , w_9113 );
and ( w_9112 , w_9113 , \2804_b0 );
or ( \2881_b1 , \731_b1 , \742_b1 );
xor ( \2881_b0 , \731_b0 , w_9114 );
not ( w_9114 , w_9115 );
and ( w_9115 , \742_b1 , \742_b0 );
or ( \2882_b1 , \2881_b1 , \751_b1 );
not ( \751_b1 , w_9116 );
and ( \2882_b0 , \2881_b0 , w_9117 );
and ( w_9116 , w_9117 , \751_b0 );
or ( \2883_b1 , \731_b1 , \742_b1 );
not ( \742_b1 , w_9118 );
and ( \2883_b0 , \731_b0 , w_9119 );
and ( w_9118 , w_9119 , \742_b0 );
or ( \2884_b1 , \2882_b1 , w_9120 );
or ( \2884_b0 , \2882_b0 , \2883_b0 );
not ( \2883_b0 , w_9121 );
and ( w_9121 , w_9120 , \2883_b1 );
buf ( \2885_b1 , \2884_b1 );
not ( \2885_b1 , w_9122 );
not ( \2885_b0 , w_9123 );
and ( w_9122 , w_9123 , \2884_b0 );
or ( \2886_b1 , \2880_b1 , \2885_b1 );
xor ( \2886_b0 , \2880_b0 , w_9124 );
not ( w_9124 , w_9125 );
and ( w_9125 , \2885_b1 , \2885_b0 );
or ( \2887_b1 , \2838_b1 , \2849_b1 );
xor ( \2887_b0 , \2838_b0 , w_9126 );
not ( w_9126 , w_9127 );
and ( w_9127 , \2849_b1 , \2849_b0 );
or ( \2888_b1 , \2887_b1 , \2842_b1 );
xor ( \2888_b0 , \2887_b0 , w_9128 );
not ( w_9128 , w_9129 );
and ( w_9129 , \2842_b1 , \2842_b0 );
or ( \2889_b1 , \2886_b1 , \2888_b1 );
not ( \2888_b1 , w_9130 );
and ( \2889_b0 , \2886_b0 , w_9131 );
and ( w_9130 , w_9131 , \2888_b0 );
or ( \2890_b1 , \2880_b1 , \2885_b1 );
not ( \2885_b1 , w_9132 );
and ( \2890_b0 , \2880_b0 , w_9133 );
and ( w_9132 , w_9133 , \2885_b0 );
or ( \2891_b1 , \2889_b1 , w_9134 );
or ( \2891_b0 , \2889_b0 , \2890_b0 );
not ( \2890_b0 , w_9135 );
and ( w_9135 , w_9134 , \2890_b1 );
or ( \2892_b1 , \2878_b1 , w_9137 );
not ( w_9137 , w_9138 );
and ( \2892_b0 , \2878_b0 , w_9139 );
and ( w_9138 ,  , w_9139 );
buf ( w_9137 , \2891_b1 );
not ( w_9137 , w_9140 );
not (  , w_9141 );
and ( w_9140 , w_9141 , \2891_b0 );
or ( \2893_b1 , \2880_b1 , \2885_b1 );
xor ( \2893_b0 , \2880_b0 , w_9142 );
not ( w_9142 , w_9143 );
and ( w_9143 , \2885_b1 , \2885_b0 );
or ( \2894_b1 , \2893_b1 , \2888_b1 );
xor ( \2894_b0 , \2893_b0 , w_9144 );
not ( w_9144 , w_9145 );
and ( w_9145 , \2888_b1 , \2888_b0 );
buf ( \2895_b1 , \693_b1 );
not ( \2895_b1 , w_9146 );
not ( \2895_b0 , w_9147 );
and ( w_9146 , w_9147 , \693_b0 );
or ( \2896_b1 , \752_b1 , w_9148 );
or ( \2896_b0 , \752_b0 , \2895_b0 );
not ( \2895_b0 , w_9149 );
and ( w_9149 , w_9148 , \2895_b1 );
or ( \2897_b1 , \2896_b1 , w_9151 );
not ( w_9151 , w_9152 );
and ( \2897_b0 , \2896_b0 , w_9153 );
and ( w_9152 ,  , w_9153 );
buf ( w_9151 , \721_b1 );
not ( w_9151 , w_9154 );
not (  , w_9155 );
and ( w_9154 , w_9155 , \721_b0 );
or ( \2898_b1 , \752_b1 , w_9157 );
not ( w_9157 , w_9158 );
and ( \2898_b0 , \752_b0 , w_9159 );
and ( w_9158 ,  , w_9159 );
buf ( w_9157 , \2895_b1 );
not ( w_9157 , w_9160 );
not (  , w_9161 );
and ( w_9160 , w_9161 , \2895_b0 );
or ( \2899_b1 , \2897_b1 , \2898_b1 );
not ( \2898_b1 , w_9162 );
and ( \2899_b0 , \2897_b0 , w_9163 );
and ( w_9162 , w_9163 , \2898_b0 );
or ( \2900_b1 , \2894_b1 , w_9165 );
not ( w_9165 , w_9166 );
and ( \2900_b0 , \2894_b0 , w_9167 );
and ( w_9166 ,  , w_9167 );
buf ( w_9165 , \2899_b1 );
not ( w_9165 , w_9168 );
not (  , w_9169 );
and ( w_9168 , w_9169 , \2899_b0 );
buf ( \2902_b1 , \2892_b1 );
not ( \2902_b1 , w_9170 );
not ( \2902_b0 , w_9171 );
and ( w_9170 , w_9171 , \2892_b0 );
or ( \2903_b1 , \2894_b1 , w_9173 );
not ( w_9173 , w_9174 );
and ( \2903_b0 , \2894_b0 , w_9175 );
and ( w_9174 ,  , w_9175 );
buf ( w_9173 , \2899_b1 );
not ( w_9173 , w_9176 );
not (  , w_9177 );
and ( w_9176 , w_9177 , \2899_b0 );
buf ( \2904_b1 , \2903_b1 );
not ( \2904_b1 , w_9178 );
not ( \2904_b0 , w_9179 );
and ( w_9178 , w_9179 , \2903_b0 );
or ( \2905_b1 , \2902_b1 , w_9180 );
or ( \2905_b0 , \2902_b0 , \2904_b0 );
not ( \2904_b0 , w_9181 );
and ( w_9181 , w_9180 , \2904_b1 );
or ( \2906_b1 , \2878_b1 , w_9182 );
or ( \2906_b0 , \2878_b0 , \2891_b0 );
not ( \2891_b0 , w_9183 );
and ( w_9183 , w_9182 , \2891_b1 );
or ( \2907_b1 , \2905_b1 , w_9185 );
not ( w_9185 , w_9186 );
and ( \2907_b0 , \2905_b0 , w_9187 );
and ( w_9186 ,  , w_9187 );
buf ( w_9185 , \2906_b1 );
not ( w_9185 , w_9188 );
not (  , w_9189 );
and ( w_9188 , w_9189 , \2906_b0 );
or ( \2908_b1 , \2833_b1 , w_9191 );
not ( w_9191 , w_9192 );
and ( \2908_b0 , \2833_b0 , w_9193 );
and ( w_9192 ,  , w_9193 );
buf ( w_9191 , \2865_b1 );
not ( w_9191 , w_9194 );
not (  , w_9195 );
and ( w_9194 , w_9195 , \2865_b0 );
or ( \2909_b1 , \2907_b1 , w_9197 );
not ( w_9197 , w_9198 );
and ( \2909_b0 , \2907_b0 , w_9199 );
and ( w_9198 ,  , w_9199 );
buf ( w_9197 , \2908_b1 );
not ( w_9197 , w_9200 );
not (  , w_9201 );
and ( w_9200 , w_9201 , \2908_b0 );
or ( \2910_b1 , \2901_b1 , w_9203 );
not ( w_9203 , w_9204 );
and ( \2910_b0 , \2901_b0 , w_9205 );
and ( w_9204 ,  , w_9205 );
buf ( w_9203 , \2909_b1 );
not ( w_9203 , w_9206 );
not (  , w_9207 );
and ( w_9206 , w_9207 , \2909_b0 );
buf ( \2911_b1 , \2910_b1 );
not ( \2911_b1 , w_9208 );
not ( \2911_b0 , w_9209 );
and ( w_9208 , w_9209 , \2910_b0 );
or ( \2912_b1 , \2868_b1 , w_9210 );
or ( \2912_b0 , \2868_b0 , \2911_b0 );
not ( \2911_b0 , w_9211 );
and ( w_9211 , w_9210 , \2911_b1 );
buf ( \2913_b1 , \2831_b1 );
buf ( \2913_b0 , \2831_b0 );
or ( \2914_b1 , \2779_b1 , w_9213 );
not ( w_9213 , w_9214 );
and ( \2914_b0 , \2779_b0 , w_9215 );
and ( w_9214 ,  , w_9215 );
buf ( w_9213 , \2813_b1 );
not ( w_9213 , w_9216 );
not (  , w_9217 );
and ( w_9216 , w_9217 , \2813_b0 );
or ( \2915_b1 , \2913_b1 , w_9219 );
not ( w_9219 , w_9220 );
and ( \2915_b0 , \2913_b0 , w_9221 );
and ( w_9220 ,  , w_9221 );
buf ( w_9219 , \2914_b1 );
not ( w_9219 , w_9222 );
not (  , w_9223 );
and ( w_9222 , w_9223 , \2914_b0 );
or ( \2916_b1 , \2912_b1 , w_9225 );
not ( w_9225 , w_9226 );
and ( \2916_b0 , \2912_b0 , w_9227 );
and ( w_9226 ,  , w_9227 );
buf ( w_9225 , \2915_b1 );
not ( w_9225 , w_9228 );
not (  , w_9229 );
and ( w_9228 , w_9229 , \2915_b0 );
buf ( \2917_b1 , \2916_b1 );
not ( \2917_b1 , w_9230 );
not ( \2917_b0 , w_9231 );
and ( w_9230 , w_9231 , \2916_b0 );
or ( \2918_b1 , \2817_b1 , w_9232 );
or ( \2918_b0 , \2817_b0 , \2917_b0 );
not ( \2917_b0 , w_9233 );
and ( w_9233 , w_9232 , \2917_b1 );
buf ( \2919_b1 , \2600_b1 );
not ( \2919_b1 , w_9234 );
not ( \2919_b0 , w_9235 );
and ( w_9234 , w_9235 , \2600_b0 );
buf ( \2920_b1 , \2658_b1 );
not ( \2920_b1 , w_9236 );
not ( \2920_b0 , w_9237 );
and ( w_9236 , w_9237 , \2658_b0 );
or ( \2921_b1 , \2919_b1 , w_9239 );
not ( w_9239 , w_9240 );
and ( \2921_b0 , \2919_b0 , w_9241 );
and ( w_9240 ,  , w_9241 );
buf ( w_9239 , \2920_b1 );
not ( w_9239 , w_9242 );
not (  , w_9243 );
and ( w_9242 , w_9243 , \2920_b0 );
buf ( \2922_b1 , \2726_b1 );
not ( \2922_b1 , w_9244 );
not ( \2922_b0 , w_9245 );
and ( w_9244 , w_9245 , \2726_b0 );
buf ( \2923_b1 , \2669_b1 );
not ( \2923_b1 , w_9246 );
not ( \2923_b0 , w_9247 );
and ( w_9246 , w_9247 , \2669_b0 );
buf ( \2924_b1 , \2923_b1 );
not ( \2924_b1 , w_9248 );
not ( \2924_b0 , w_9249 );
and ( w_9248 , w_9249 , \2923_b0 );
or ( \2925_b1 , \2922_b1 , w_9250 );
or ( \2925_b0 , \2922_b0 , \2924_b0 );
not ( \2924_b0 , w_9251 );
and ( w_9251 , w_9250 , \2924_b1 );
or ( \2926_b1 , \2826_b1 , w_9252 );
or ( \2926_b0 , \2826_b0 , \2830_b0 );
not ( \2830_b0 , w_9253 );
and ( w_9253 , w_9252 , \2830_b1 );
or ( \2927_b1 , \2925_b1 , w_9255 );
not ( w_9255 , w_9256 );
and ( \2927_b0 , \2925_b0 , w_9257 );
and ( w_9256 ,  , w_9257 );
buf ( w_9255 , \2926_b1 );
not ( w_9255 , w_9258 );
not (  , w_9259 );
and ( w_9258 , w_9259 , \2926_b0 );
or ( \2929_b1 , \2920_b1 , w_9261 );
not ( w_9261 , w_9262 );
and ( \2929_b0 , \2920_b0 , w_9263 );
and ( w_9262 ,  , w_9263 );
buf ( w_9261 , \2919_b1 );
not ( w_9261 , w_9264 );
not (  , w_9265 );
and ( w_9264 , w_9265 , \2919_b0 );
or ( \2930_b1 , \2928_b1 , w_9267 );
not ( w_9267 , w_9268 );
and ( \2930_b0 , \2928_b0 , w_9269 );
and ( w_9268 ,  , w_9269 );
buf ( w_9267 , \2929_b1 );
not ( w_9267 , w_9270 );
not (  , w_9271 );
and ( w_9270 , w_9271 , \2929_b0 );
or ( \2931_b1 , \2918_b1 , w_9273 );
not ( w_9273 , w_9274 );
and ( \2931_b0 , \2918_b0 , w_9275 );
and ( w_9274 ,  , w_9275 );
buf ( w_9273 , \2930_b1 );
not ( w_9273 , w_9276 );
not (  , w_9277 );
and ( w_9276 , w_9277 , \2930_b0 );
buf ( \2932_b1 , \2931_b1 );
not ( \2932_b1 , w_9278 );
not ( \2932_b0 , w_9279 );
and ( w_9278 , w_9279 , \2931_b0 );
or ( \2933_b1 , \2598_b1 , w_9280 );
or ( \2933_b0 , \2598_b0 , \2932_b0 );
not ( \2932_b0 , w_9281 );
and ( w_9281 , w_9280 , \2932_b1 );
or ( \2934_b1 , \2931_b1 , w_9282 );
or ( \2934_b0 , \2931_b0 , \2597_b0 );
not ( \2597_b0 , w_9283 );
and ( w_9283 , w_9282 , \2597_b1 );
or ( \2935_b1 , \2933_b1 , w_9285 );
not ( w_9285 , w_9286 );
and ( \2935_b0 , \2933_b0 , w_9287 );
and ( w_9286 ,  , w_9287 );
buf ( w_9285 , \2934_b1 );
not ( w_9285 , w_9288 );
not (  , w_9289 );
and ( w_9288 , w_9289 , \2934_b0 );
buf ( \2936_b1 , \917_b1 );
not ( \2936_b1 , w_9290 );
not ( \2936_b0 , w_9291 );
and ( w_9290 , w_9291 , \917_b0 );
or ( \2937_b1 , \2935_b1 , w_9293 );
not ( w_9293 , w_9294 );
and ( \2937_b0 , \2935_b0 , w_9295 );
and ( w_9294 ,  , w_9295 );
buf ( w_9293 , \2936_b1 );
not ( w_9293 , w_9296 );
not (  , w_9297 );
and ( w_9296 , w_9297 , \2936_b0 );
or ( \2938_b1 , \2233_b1 , w_9299 );
not ( w_9299 , w_9300 );
and ( \2938_b0 , \2233_b0 , w_9301 );
and ( w_9300 ,  , w_9301 );
buf ( w_9299 , \2937_b1 );
not ( w_9299 , w_9302 );
not (  , w_9303 );
and ( w_9302 , w_9303 , \2937_b0 );
buf ( \2939_b1 , \a[15]_b1 );
not ( \2939_b1 , w_9304 );
not ( \2939_b0 , w_9305 );
and ( w_9304 , w_9305 , \a[15]_b0 );
buf ( \2940_b1 , \1331_b1 );
not ( \2940_b1 , w_9306 );
not ( \2940_b0 , w_9307 );
and ( w_9306 , w_9307 , \1331_b0 );
buf ( \2941_b1 , \2940_b1 );
not ( \2941_b1 , w_9308 );
not ( \2941_b0 , w_9309 );
and ( w_9308 , w_9309 , \2940_b0 );
buf ( \2942_b1 , \1316_b1 );
not ( \2942_b1 , w_9310 );
not ( \2942_b0 , w_9311 );
and ( w_9310 , w_9311 , \1316_b0 );
buf ( \2943_b1 , \2942_b1 );
not ( \2943_b1 , w_9312 );
not ( \2943_b0 , w_9313 );
and ( w_9312 , w_9313 , \2942_b0 );
or ( \2944_b1 , \2941_b1 , w_9314 );
or ( \2944_b0 , \2941_b0 , \2943_b0 );
not ( \2943_b0 , w_9315 );
and ( w_9315 , w_9314 , \2943_b1 );
buf ( \2945_b1 , \644_b1 );
not ( \2945_b1 , w_9316 );
not ( \2945_b0 , w_9317 );
and ( w_9316 , w_9317 , \644_b0 );
or ( \2946_b1 , \2944_b1 , w_9319 );
not ( w_9319 , w_9320 );
and ( \2946_b0 , \2944_b0 , w_9321 );
and ( w_9320 ,  , w_9321 );
buf ( w_9319 , \2945_b1 );
not ( w_9319 , w_9322 );
not (  , w_9323 );
and ( w_9322 , w_9323 , \2945_b0 );
buf ( \2947_b1 , \2946_b1 );
not ( \2947_b1 , w_9324 );
not ( \2947_b0 , w_9325 );
and ( w_9324 , w_9325 , \2946_b0 );
or ( \2948_b1 , \2939_b1 , w_9326 );
or ( \2948_b0 , \2939_b0 , \2947_b0 );
not ( \2947_b0 , w_9327 );
and ( w_9327 , w_9326 , \2947_b1 );
buf ( \2949_b1 , \b[15]_b1 );
not ( \2949_b1 , w_9328 );
not ( \2949_b0 , w_9329 );
and ( w_9328 , w_9329 , \b[15]_b0 );
buf ( \2950_b1 , \672_b1 );
not ( \2950_b1 , w_9330 );
not ( \2950_b0 , w_9331 );
and ( w_9330 , w_9331 , \672_b0 );
or ( \2951_b1 , \2950_b1 , w_9333 );
not ( w_9333 , w_9334 );
and ( \2951_b0 , \2950_b0 , w_9335 );
and ( w_9334 ,  , w_9335 );
buf ( w_9333 , \1324_b1 );
not ( w_9333 , w_9336 );
not (  , w_9337 );
and ( w_9336 , w_9337 , \1324_b0 );
buf ( \2952_b1 , \2951_b1 );
not ( \2952_b1 , w_9338 );
not ( \2952_b0 , w_9339 );
and ( w_9338 , w_9339 , \2951_b0 );
or ( \2953_b1 , \2949_b1 , w_9340 );
or ( \2953_b0 , \2949_b0 , \2952_b0 );
not ( \2952_b0 , w_9341 );
and ( w_9341 , w_9340 , \2952_b1 );
buf ( \2954_b1 , \1466_b1 );
buf ( \2954_b0 , \1466_b0 );
or ( \2955_b1 , \2954_b1 , \a[15]_b1 );
not ( \a[15]_b1 , w_9342 );
and ( \2955_b0 , \2954_b0 , w_9343 );
and ( w_9342 , w_9343 , \a[15]_b0 );
or ( \2956_b1 , \c[15]_b1 , \d[15]_b1 );
xor ( \2956_b0 , \c[15]_b0 , w_9344 );
not ( w_9344 , w_9345 );
and ( w_9345 , \d[15]_b1 , \d[15]_b0 );
buf ( \2957_b1 , \2956_b1 );
not ( \2957_b1 , w_9346 );
not ( \2957_b0 , w_9347 );
and ( w_9346 , w_9347 , \2956_b0 );
buf ( \2958_b1 , \925_b1 );
not ( \2958_b1 , w_9348 );
not ( \2958_b0 , w_9349 );
and ( w_9348 , w_9349 , \925_b0 );
or ( \2959_b1 , \2957_b1 , w_9350 );
or ( \2959_b0 , \2957_b0 , \2958_b0 );
not ( \2958_b0 , w_9351 );
and ( w_9351 , w_9350 , \2958_b1 );
buf ( \2960_b1 , \1220_b1 );
not ( \2960_b1 , w_9352 );
not ( \2960_b0 , w_9353 );
and ( w_9352 , w_9353 , \1220_b0 );
buf ( \2961_b1 , \2960_b1 );
not ( \2961_b1 , w_9354 );
not ( \2961_b0 , w_9355 );
and ( w_9354 , w_9355 , \2960_b0 );
or ( \2962_b1 , \b[15]_b1 , \d[15]_b1 );
not ( \d[15]_b1 , w_9356 );
and ( \2962_b0 , \b[15]_b0 , w_9357 );
and ( w_9356 , w_9357 , \d[15]_b0 );
or ( \2963_b1 , \b[15]_b1 , w_9359 );
not ( w_9359 , w_9360 );
and ( \2963_b0 , \b[15]_b0 , w_9361 );
and ( w_9360 ,  , w_9361 );
buf ( w_9359 , \d[15]_b1 );
not ( w_9359 , w_9362 );
not (  , w_9363 );
and ( w_9362 , w_9363 , \d[15]_b0 );
or ( \2964_b1 , \2962_b1 , w_9365 );
not ( w_9365 , w_9366 );
and ( \2964_b0 , \2962_b0 , w_9367 );
and ( w_9366 ,  , w_9367 );
buf ( w_9365 , \2963_b1 );
not ( w_9365 , w_9368 );
not (  , w_9369 );
and ( w_9368 , w_9369 , \2963_b0 );
buf ( \2965_b1 , \2964_b1 );
not ( \2965_b1 , w_9370 );
not ( \2965_b0 , w_9371 );
and ( w_9370 , w_9371 , \2964_b0 );
buf ( \2967_b1 , \2966_b1 );
not ( \2967_b1 , w_9372 );
not ( \2967_b0 , w_9373 );
and ( w_9372 , w_9373 , \2966_b0 );
or ( \2969_b1 , \1193_b1 , w_9375 );
not ( w_9375 , w_9376 );
and ( \2969_b0 , \1193_b0 , w_9377 );
and ( w_9376 ,  , w_9377 );
buf ( w_9375 , \2968_b1 );
not ( w_9375 , w_9378 );
not (  , w_9379 );
and ( w_9378 , w_9379 , \2968_b0 );
buf ( \2970_b1 , \2969_b1 );
not ( \2970_b1 , w_9380 );
not ( \2970_b0 , w_9381 );
and ( w_9380 , w_9381 , \2969_b0 );
or ( \2971_b1 , \2967_b1 , w_9382 );
or ( \2971_b0 , \2967_b0 , \2970_b0 );
not ( \2970_b0 , w_9383 );
and ( w_9383 , w_9382 , \2970_b1 );
buf ( \2973_b1 , \2972_b1 );
not ( \2973_b1 , w_9384 );
not ( \2973_b0 , w_9385 );
and ( w_9384 , w_9385 , \2972_b0 );
buf ( \2974_b1 , \1199_b1 );
not ( \2974_b1 , w_9386 );
not ( \2974_b0 , w_9387 );
and ( w_9386 , w_9387 , \1199_b0 );
or ( \2975_b1 , \2973_b1 , w_9388 );
or ( \2975_b0 , \2973_b0 , \2974_b0 );
not ( \2974_b0 , w_9389 );
and ( w_9389 , w_9388 , \2974_b1 );
or ( \2976_b1 , \1208_b1 , w_9390 );
or ( \2976_b0 , \1208_b0 , \1194_b0 );
not ( \1194_b0 , w_9391 );
and ( w_9391 , w_9390 , \1194_b1 );
or ( \2977_b1 , \2976_b1 , w_9393 );
not ( w_9393 , w_9394 );
and ( \2977_b0 , \2976_b0 , w_9395 );
and ( w_9394 ,  , w_9395 );
buf ( w_9393 , \1210_b1 );
not ( w_9393 , w_9396 );
not (  , w_9397 );
and ( w_9396 , w_9397 , \1210_b0 );
or ( \2978_b1 , \2975_b1 , w_9399 );
not ( w_9399 , w_9400 );
and ( \2978_b0 , \2975_b0 , w_9401 );
and ( w_9400 ,  , w_9401 );
buf ( w_9399 , \2977_b1 );
not ( w_9399 , w_9402 );
not (  , w_9403 );
and ( w_9402 , w_9403 , \2977_b0 );
or ( \2979_b1 , \2971_b1 , w_9405 );
not ( w_9405 , w_9406 );
and ( \2979_b0 , \2971_b0 , w_9407 );
and ( w_9406 ,  , w_9407 );
buf ( w_9405 , \2978_b1 );
not ( w_9405 , w_9408 );
not (  , w_9409 );
and ( w_9408 , w_9409 , \2978_b0 );
or ( \2980_b1 , \b[13]_b1 , w_9411 );
not ( w_9411 , w_9412 );
and ( \2980_b0 , \b[13]_b0 , w_9413 );
and ( w_9412 ,  , w_9413 );
buf ( w_9411 , \d[13]_b1 );
not ( w_9411 , w_9414 );
not (  , w_9415 );
and ( w_9414 , w_9415 , \d[13]_b0 );
or ( \2981_b1 , \b[12]_b1 , w_9417 );
not ( w_9417 , w_9418 );
and ( \2981_b0 , \b[12]_b0 , w_9419 );
and ( w_9418 ,  , w_9419 );
buf ( w_9417 , \d[12]_b1 );
not ( w_9417 , w_9420 );
not (  , w_9421 );
and ( w_9420 , w_9421 , \d[12]_b0 );
or ( \2982_b1 , \2980_b1 , w_9423 );
not ( w_9423 , w_9424 );
and ( \2982_b0 , \2980_b0 , w_9425 );
and ( w_9424 ,  , w_9425 );
buf ( w_9423 , \2981_b1 );
not ( w_9423 , w_9426 );
not (  , w_9427 );
and ( w_9426 , w_9427 , \2981_b0 );
or ( \2983_b1 , \b[14]_b1 , w_9428 );
or ( \2983_b0 , \b[14]_b0 , \d[14]_b0 );
not ( \d[14]_b0 , w_9429 );
and ( w_9429 , w_9428 , \d[14]_b1 );
or ( \2984_b1 , \2982_b1 , w_9431 );
not ( w_9431 , w_9432 );
and ( \2984_b0 , \2982_b0 , w_9433 );
and ( w_9432 ,  , w_9433 );
buf ( w_9431 , \2983_b1 );
not ( w_9431 , w_9434 );
not (  , w_9435 );
and ( w_9434 , w_9435 , \2983_b0 );
buf ( \2985_b1 , \2984_b1 );
not ( \2985_b1 , w_9436 );
not ( \2985_b0 , w_9437 );
and ( w_9436 , w_9437 , \2984_b0 );
or ( \2986_b1 , \b[11]_b1 , w_9439 );
not ( w_9439 , w_9440 );
and ( \2986_b0 , \b[11]_b0 , w_9441 );
and ( w_9440 ,  , w_9441 );
buf ( w_9439 , \d[11]_b1 );
not ( w_9439 , w_9442 );
not (  , w_9443 );
and ( w_9442 , w_9443 , \d[11]_b0 );
or ( \2987_b1 , \b[10]_b1 , w_9445 );
not ( w_9445 , w_9446 );
and ( \2987_b0 , \b[10]_b0 , w_9447 );
and ( w_9446 ,  , w_9447 );
buf ( w_9445 , \d[10]_b1 );
not ( w_9445 , w_9448 );
not (  , w_9449 );
and ( w_9448 , w_9449 , \d[10]_b0 );
or ( \2988_b1 , \2986_b1 , w_9451 );
not ( w_9451 , w_9452 );
and ( \2988_b0 , \2986_b0 , w_9453 );
and ( w_9452 ,  , w_9453 );
buf ( w_9451 , \2987_b1 );
not ( w_9451 , w_9454 );
not (  , w_9455 );
and ( w_9454 , w_9455 , \2987_b0 );
or ( \2989_b1 , \b[8]_b1 , w_9457 );
not ( w_9457 , w_9458 );
and ( \2989_b0 , \b[8]_b0 , w_9459 );
and ( w_9458 ,  , w_9459 );
buf ( w_9457 , \d[8]_b1 );
not ( w_9457 , w_9460 );
not (  , w_9461 );
and ( w_9460 , w_9461 , \d[8]_b0 );
or ( \2990_b1 , \b[9]_b1 , w_9463 );
not ( w_9463 , w_9464 );
and ( \2990_b0 , \b[9]_b0 , w_9465 );
and ( w_9464 ,  , w_9465 );
buf ( w_9463 , \d[9]_b1 );
not ( w_9463 , w_9466 );
not (  , w_9467 );
and ( w_9466 , w_9467 , \d[9]_b0 );
or ( \2991_b1 , \2989_b1 , w_9469 );
not ( w_9469 , w_9470 );
and ( \2991_b0 , \2989_b0 , w_9471 );
and ( w_9470 ,  , w_9471 );
buf ( w_9469 , \2990_b1 );
not ( w_9469 , w_9472 );
not (  , w_9473 );
and ( w_9472 , w_9473 , \2990_b0 );
or ( \2992_b1 , \2988_b1 , \2991_b1 );
not ( \2991_b1 , w_9474 );
and ( \2992_b0 , \2988_b0 , w_9475 );
and ( w_9474 , w_9475 , \2991_b0 );
or ( \2994_b1 , \b[8]_b1 , w_9477 );
not ( w_9477 , w_9478 );
and ( \2994_b0 , \b[8]_b0 , w_9479 );
and ( w_9478 ,  , w_9479 );
buf ( w_9477 , \d[8]_b1 );
not ( w_9477 , w_9480 );
not (  , w_9481 );
and ( w_9480 , w_9481 , \d[8]_b0 );
or ( \2995_b1 , \2990_b1 , w_9482 );
or ( \2995_b0 , \2990_b0 , \2994_b0 );
not ( \2994_b0 , w_9483 );
and ( w_9483 , w_9482 , \2994_b1 );
or ( \2996_b1 , \b[9]_b1 , w_9485 );
not ( w_9485 , w_9486 );
and ( \2996_b0 , \b[9]_b0 , w_9487 );
and ( w_9486 ,  , w_9487 );
buf ( w_9485 , \d[9]_b1 );
not ( w_9485 , w_9488 );
not (  , w_9489 );
and ( w_9488 , w_9489 , \d[9]_b0 );
or ( \2997_b1 , \2995_b1 , w_9491 );
not ( w_9491 , w_9492 );
and ( \2997_b0 , \2995_b0 , w_9493 );
and ( w_9492 ,  , w_9493 );
buf ( w_9491 , \2996_b1 );
not ( w_9491 , w_9494 );
not (  , w_9495 );
and ( w_9494 , w_9495 , \2996_b0 );
buf ( \2998_b1 , \2997_b1 );
not ( \2998_b1 , w_9496 );
not ( \2998_b0 , w_9497 );
and ( w_9496 , w_9497 , \2997_b0 );
buf ( \2999_b1 , \2988_b1 );
not ( \2999_b1 , w_9498 );
not ( \2999_b0 , w_9499 );
and ( w_9498 , w_9499 , \2988_b0 );
or ( \3000_b1 , \2998_b1 , w_9500 );
or ( \3000_b0 , \2998_b0 , \2999_b0 );
not ( \2999_b0 , w_9501 );
and ( w_9501 , w_9500 , \2999_b1 );
buf ( \3001_b1 , \2986_b1 );
not ( \3001_b1 , w_9502 );
not ( \3001_b0 , w_9503 );
and ( w_9502 , w_9503 , \2986_b0 );
or ( \3002_b1 , \b[10]_b1 , w_9505 );
not ( w_9505 , w_9506 );
and ( \3002_b0 , \b[10]_b0 , w_9507 );
and ( w_9506 ,  , w_9507 );
buf ( w_9505 , \d[10]_b1 );
not ( w_9505 , w_9508 );
not (  , w_9509 );
and ( w_9508 , w_9509 , \d[10]_b0 );
buf ( \3003_b1 , \3002_b1 );
not ( \3003_b1 , w_9510 );
not ( \3003_b0 , w_9511 );
and ( w_9510 , w_9511 , \3002_b0 );
or ( \3004_b1 , \3001_b1 , \3003_b1 );
not ( \3003_b1 , w_9512 );
and ( \3004_b0 , \3001_b0 , w_9513 );
and ( w_9512 , w_9513 , \3003_b0 );
or ( \3005_b1 , \b[11]_b1 , \d[11]_b1 );
not ( \d[11]_b1 , w_9514 );
and ( \3005_b0 , \b[11]_b0 , w_9515 );
and ( w_9514 , w_9515 , \d[11]_b0 );
or ( \3006_b1 , \3004_b1 , w_9517 );
not ( w_9517 , w_9518 );
and ( \3006_b0 , \3004_b0 , w_9519 );
and ( w_9518 ,  , w_9519 );
buf ( w_9517 , \3005_b1 );
not ( w_9517 , w_9520 );
not (  , w_9521 );
and ( w_9520 , w_9521 , \3005_b0 );
or ( \3007_b1 , \3000_b1 , w_9523 );
not ( w_9523 , w_9524 );
and ( \3007_b0 , \3000_b0 , w_9525 );
and ( w_9524 ,  , w_9525 );
buf ( w_9523 , \3006_b1 );
not ( w_9523 , w_9526 );
not (  , w_9527 );
and ( w_9526 , w_9527 , \3006_b0 );
buf ( \3008_b1 , \3007_b1 );
not ( \3008_b1 , w_9528 );
not ( \3008_b0 , w_9529 );
and ( w_9528 , w_9529 , \3007_b0 );
or ( \3009_b1 , \3008_b1 , w_9530 );
or ( \3009_b0 , \3008_b0 , \2984_b0 );
not ( \2984_b0 , w_9531 );
and ( w_9531 , w_9530 , \2984_b1 );
or ( \3010_b1 , \b[12]_b1 , w_9533 );
not ( w_9533 , w_9534 );
and ( \3010_b0 , \b[12]_b0 , w_9535 );
and ( w_9534 ,  , w_9535 );
buf ( w_9533 , \d[12]_b1 );
not ( w_9533 , w_9536 );
not (  , w_9537 );
and ( w_9536 , w_9537 , \d[12]_b0 );
or ( \3011_b1 , \2980_b1 , w_9538 );
or ( \3011_b0 , \2980_b0 , \3010_b0 );
not ( \3010_b0 , w_9539 );
and ( w_9539 , w_9538 , \3010_b1 );
or ( \3012_b1 , \b[13]_b1 , w_9541 );
not ( w_9541 , w_9542 );
and ( \3012_b0 , \b[13]_b0 , w_9543 );
and ( w_9542 ,  , w_9543 );
buf ( w_9541 , \d[13]_b1 );
not ( w_9541 , w_9544 );
not (  , w_9545 );
and ( w_9544 , w_9545 , \d[13]_b0 );
or ( \3013_b1 , \3011_b1 , w_9547 );
not ( w_9547 , w_9548 );
and ( \3013_b0 , \3011_b0 , w_9549 );
and ( w_9548 ,  , w_9549 );
buf ( w_9547 , \3012_b1 );
not ( w_9547 , w_9550 );
not (  , w_9551 );
and ( w_9550 , w_9551 , \3012_b0 );
or ( \3014_b1 , \3013_b1 , \2983_b1 );
not ( \2983_b1 , w_9552 );
and ( \3014_b0 , \3013_b0 , w_9553 );
and ( w_9552 , w_9553 , \2983_b0 );
or ( \3015_b1 , \b[14]_b1 , \d[14]_b1 );
not ( \d[14]_b1 , w_9554 );
and ( \3015_b0 , \b[14]_b0 , w_9555 );
and ( w_9554 , w_9555 , \d[14]_b0 );
or ( \3016_b1 , \3014_b1 , w_9557 );
not ( w_9557 , w_9558 );
and ( \3016_b0 , \3014_b0 , w_9559 );
and ( w_9558 ,  , w_9559 );
buf ( w_9557 , \3015_b1 );
not ( w_9557 , w_9560 );
not (  , w_9561 );
and ( w_9560 , w_9561 , \3015_b0 );
or ( \3017_b1 , \3009_b1 , w_9563 );
not ( w_9563 , w_9564 );
and ( \3017_b0 , \3009_b0 , w_9565 );
and ( w_9564 ,  , w_9565 );
buf ( w_9563 , \3016_b1 );
not ( w_9563 , w_9566 );
not (  , w_9567 );
and ( w_9566 , w_9567 , \3016_b0 );
or ( \3018_b1 , \2993_b1 , w_9569 );
not ( w_9569 , w_9570 );
and ( \3018_b0 , \2993_b0 , w_9571 );
and ( w_9570 ,  , w_9571 );
buf ( w_9569 , \3017_b1 );
not ( w_9569 , w_9572 );
not (  , w_9573 );
and ( w_9572 , w_9573 , \3017_b0 );
buf ( \3019_b1 , \3018_b1 );
not ( \3019_b1 , w_9574 );
not ( \3019_b0 , w_9575 );
and ( w_9574 , w_9575 , \3018_b0 );
or ( \3020_b1 , \2965_b1 , w_9576 );
or ( \3020_b0 , \2965_b0 , \3019_b0 );
not ( \3019_b0 , w_9577 );
and ( w_9577 , w_9576 , \3019_b1 );
or ( \3021_b1 , \3018_b1 , w_9578 );
or ( \3021_b0 , \3018_b0 , \2964_b0 );
not ( \2964_b0 , w_9579 );
and ( w_9579 , w_9578 , \2964_b1 );
or ( \3022_b1 , \3020_b1 , w_9581 );
not ( w_9581 , w_9582 );
and ( \3022_b0 , \3020_b0 , w_9583 );
and ( w_9582 ,  , w_9583 );
buf ( w_9581 , \3021_b1 );
not ( w_9581 , w_9584 );
not (  , w_9585 );
and ( w_9584 , w_9585 , \3021_b0 );
or ( \3023_b1 , \2961_b1 , \3022_b1 );
not ( \3022_b1 , w_9586 );
and ( \3023_b0 , \2961_b0 , w_9587 );
and ( w_9586 , w_9587 , \3022_b0 );
or ( \3024_b1 , \a[15]_b1 , \c[15]_b1 );
not ( \c[15]_b1 , w_9588 );
and ( \3024_b0 , \a[15]_b0 , w_9589 );
and ( w_9588 , w_9589 , \c[15]_b0 );
or ( \3025_b1 , \a[15]_b1 , w_9591 );
not ( w_9591 , w_9592 );
and ( \3025_b0 , \a[15]_b0 , w_9593 );
and ( w_9592 ,  , w_9593 );
buf ( w_9591 , \c[15]_b1 );
not ( w_9591 , w_9594 );
not (  , w_9595 );
and ( w_9594 , w_9595 , \c[15]_b0 );
or ( \3026_b1 , \3024_b1 , w_9597 );
not ( w_9597 , w_9598 );
and ( \3026_b0 , \3024_b0 , w_9599 );
and ( w_9598 ,  , w_9599 );
buf ( w_9597 , \3025_b1 );
not ( w_9597 , w_9600 );
not (  , w_9601 );
and ( w_9600 , w_9601 , \3025_b0 );
buf ( \3027_b1 , \3026_b1 );
not ( \3027_b1 , w_9602 );
not ( \3027_b0 , w_9603 );
and ( w_9602 , w_9603 , \3026_b0 );
buf ( \3029_b1 , \3028_b1 );
not ( \3029_b1 , w_9604 );
not ( \3029_b0 , w_9605 );
and ( w_9604 , w_9605 , \3028_b0 );
or ( \3031_b1 , \1256_b1 , w_9607 );
not ( w_9607 , w_9608 );
and ( \3031_b0 , \1256_b0 , w_9609 );
and ( w_9608 ,  , w_9609 );
buf ( w_9607 , \3030_b1 );
not ( w_9607 , w_9610 );
not (  , w_9611 );
and ( w_9610 , w_9611 , \3030_b0 );
buf ( \3032_b1 , \3031_b1 );
not ( \3032_b1 , w_9612 );
not ( \3032_b0 , w_9613 );
and ( w_9612 , w_9613 , \3031_b0 );
or ( \3033_b1 , \3029_b1 , w_9614 );
or ( \3033_b0 , \3029_b0 , \3032_b0 );
not ( \3032_b0 , w_9615 );
and ( w_9615 , w_9614 , \3032_b1 );
buf ( \3035_b1 , \3034_b1 );
not ( \3035_b1 , w_9616 );
not ( \3035_b0 , w_9617 );
and ( w_9616 , w_9617 , \3034_b0 );
buf ( \3036_b1 , \1262_b1 );
not ( \3036_b1 , w_9618 );
not ( \3036_b0 , w_9619 );
and ( w_9618 , w_9619 , \1262_b0 );
or ( \3037_b1 , \3035_b1 , w_9620 );
or ( \3037_b0 , \3035_b0 , \3036_b0 );
not ( \3036_b0 , w_9621 );
and ( w_9621 , w_9620 , \3036_b1 );
or ( \3038_b1 , \1271_b1 , w_9622 );
or ( \3038_b0 , \1271_b0 , \1257_b0 );
not ( \1257_b0 , w_9623 );
and ( w_9623 , w_9622 , \1257_b1 );
or ( \3039_b1 , \3038_b1 , w_9625 );
not ( w_9625 , w_9626 );
and ( \3039_b0 , \3038_b0 , w_9627 );
and ( w_9626 ,  , w_9627 );
buf ( w_9625 , \1273_b1 );
not ( w_9625 , w_9628 );
not (  , w_9629 );
and ( w_9628 , w_9629 , \1273_b0 );
or ( \3040_b1 , \3037_b1 , w_9631 );
not ( w_9631 , w_9632 );
and ( \3040_b0 , \3037_b0 , w_9633 );
and ( w_9632 ,  , w_9633 );
buf ( w_9631 , \3039_b1 );
not ( w_9631 , w_9634 );
not (  , w_9635 );
and ( w_9634 , w_9635 , \3039_b0 );
or ( \3041_b1 , \3033_b1 , w_9637 );
not ( w_9637 , w_9638 );
and ( \3041_b0 , \3033_b0 , w_9639 );
and ( w_9638 ,  , w_9639 );
buf ( w_9637 , \3040_b1 );
not ( w_9637 , w_9640 );
not (  , w_9641 );
and ( w_9640 , w_9641 , \3040_b0 );
or ( \3042_b1 , \a[13]_b1 , w_9643 );
not ( w_9643 , w_9644 );
and ( \3042_b0 , \a[13]_b0 , w_9645 );
and ( w_9644 ,  , w_9645 );
buf ( w_9643 , \c[13]_b1 );
not ( w_9643 , w_9646 );
not (  , w_9647 );
and ( w_9646 , w_9647 , \c[13]_b0 );
or ( \3043_b1 , \a[12]_b1 , w_9649 );
not ( w_9649 , w_9650 );
and ( \3043_b0 , \a[12]_b0 , w_9651 );
and ( w_9650 ,  , w_9651 );
buf ( w_9649 , \c[12]_b1 );
not ( w_9649 , w_9652 );
not (  , w_9653 );
and ( w_9652 , w_9653 , \c[12]_b0 );
or ( \3044_b1 , \3042_b1 , w_9655 );
not ( w_9655 , w_9656 );
and ( \3044_b0 , \3042_b0 , w_9657 );
and ( w_9656 ,  , w_9657 );
buf ( w_9655 , \3043_b1 );
not ( w_9655 , w_9658 );
not (  , w_9659 );
and ( w_9658 , w_9659 , \3043_b0 );
or ( \3045_b1 , \a[14]_b1 , w_9660 );
or ( \3045_b0 , \a[14]_b0 , \c[14]_b0 );
not ( \c[14]_b0 , w_9661 );
and ( w_9661 , w_9660 , \c[14]_b1 );
or ( \3046_b1 , \3044_b1 , w_9663 );
not ( w_9663 , w_9664 );
and ( \3046_b0 , \3044_b0 , w_9665 );
and ( w_9664 ,  , w_9665 );
buf ( w_9663 , \3045_b1 );
not ( w_9663 , w_9666 );
not (  , w_9667 );
and ( w_9666 , w_9667 , \3045_b0 );
buf ( \3047_b1 , \3046_b1 );
not ( \3047_b1 , w_9668 );
not ( \3047_b0 , w_9669 );
and ( w_9668 , w_9669 , \3046_b0 );
or ( \3048_b1 , \a[11]_b1 , w_9671 );
not ( w_9671 , w_9672 );
and ( \3048_b0 , \a[11]_b0 , w_9673 );
and ( w_9672 ,  , w_9673 );
buf ( w_9671 , \c[11]_b1 );
not ( w_9671 , w_9674 );
not (  , w_9675 );
and ( w_9674 , w_9675 , \c[11]_b0 );
or ( \3049_b1 , \a[10]_b1 , w_9677 );
not ( w_9677 , w_9678 );
and ( \3049_b0 , \a[10]_b0 , w_9679 );
and ( w_9678 ,  , w_9679 );
buf ( w_9677 , \c[10]_b1 );
not ( w_9677 , w_9680 );
not (  , w_9681 );
and ( w_9680 , w_9681 , \c[10]_b0 );
or ( \3050_b1 , \3048_b1 , w_9683 );
not ( w_9683 , w_9684 );
and ( \3050_b0 , \3048_b0 , w_9685 );
and ( w_9684 ,  , w_9685 );
buf ( w_9683 , \3049_b1 );
not ( w_9683 , w_9686 );
not (  , w_9687 );
and ( w_9686 , w_9687 , \3049_b0 );
or ( \3051_b1 , \a[8]_b1 , w_9689 );
not ( w_9689 , w_9690 );
and ( \3051_b0 , \a[8]_b0 , w_9691 );
and ( w_9690 ,  , w_9691 );
buf ( w_9689 , \c[8]_b1 );
not ( w_9689 , w_9692 );
not (  , w_9693 );
and ( w_9692 , w_9693 , \c[8]_b0 );
or ( \3052_b1 , \a[9]_b1 , w_9695 );
not ( w_9695 , w_9696 );
and ( \3052_b0 , \a[9]_b0 , w_9697 );
and ( w_9696 ,  , w_9697 );
buf ( w_9695 , \c[9]_b1 );
not ( w_9695 , w_9698 );
not (  , w_9699 );
and ( w_9698 , w_9699 , \c[9]_b0 );
or ( \3053_b1 , \3051_b1 , w_9701 );
not ( w_9701 , w_9702 );
and ( \3053_b0 , \3051_b0 , w_9703 );
and ( w_9702 ,  , w_9703 );
buf ( w_9701 , \3052_b1 );
not ( w_9701 , w_9704 );
not (  , w_9705 );
and ( w_9704 , w_9705 , \3052_b0 );
or ( \3054_b1 , \3050_b1 , \3053_b1 );
not ( \3053_b1 , w_9706 );
and ( \3054_b0 , \3050_b0 , w_9707 );
and ( w_9706 , w_9707 , \3053_b0 );
or ( \3056_b1 , \a[8]_b1 , w_9709 );
not ( w_9709 , w_9710 );
and ( \3056_b0 , \a[8]_b0 , w_9711 );
and ( w_9710 ,  , w_9711 );
buf ( w_9709 , \c[8]_b1 );
not ( w_9709 , w_9712 );
not (  , w_9713 );
and ( w_9712 , w_9713 , \c[8]_b0 );
or ( \3057_b1 , \3052_b1 , w_9714 );
or ( \3057_b0 , \3052_b0 , \3056_b0 );
not ( \3056_b0 , w_9715 );
and ( w_9715 , w_9714 , \3056_b1 );
or ( \3058_b1 , \a[9]_b1 , w_9717 );
not ( w_9717 , w_9718 );
and ( \3058_b0 , \a[9]_b0 , w_9719 );
and ( w_9718 ,  , w_9719 );
buf ( w_9717 , \c[9]_b1 );
not ( w_9717 , w_9720 );
not (  , w_9721 );
and ( w_9720 , w_9721 , \c[9]_b0 );
or ( \3059_b1 , \3057_b1 , w_9723 );
not ( w_9723 , w_9724 );
and ( \3059_b0 , \3057_b0 , w_9725 );
and ( w_9724 ,  , w_9725 );
buf ( w_9723 , \3058_b1 );
not ( w_9723 , w_9726 );
not (  , w_9727 );
and ( w_9726 , w_9727 , \3058_b0 );
buf ( \3060_b1 , \3059_b1 );
not ( \3060_b1 , w_9728 );
not ( \3060_b0 , w_9729 );
and ( w_9728 , w_9729 , \3059_b0 );
buf ( \3061_b1 , \3050_b1 );
not ( \3061_b1 , w_9730 );
not ( \3061_b0 , w_9731 );
and ( w_9730 , w_9731 , \3050_b0 );
or ( \3062_b1 , \3060_b1 , w_9732 );
or ( \3062_b0 , \3060_b0 , \3061_b0 );
not ( \3061_b0 , w_9733 );
and ( w_9733 , w_9732 , \3061_b1 );
buf ( \3063_b1 , \3048_b1 );
not ( \3063_b1 , w_9734 );
not ( \3063_b0 , w_9735 );
and ( w_9734 , w_9735 , \3048_b0 );
or ( \3064_b1 , \a[10]_b1 , w_9737 );
not ( w_9737 , w_9738 );
and ( \3064_b0 , \a[10]_b0 , w_9739 );
and ( w_9738 ,  , w_9739 );
buf ( w_9737 , \c[10]_b1 );
not ( w_9737 , w_9740 );
not (  , w_9741 );
and ( w_9740 , w_9741 , \c[10]_b0 );
buf ( \3065_b1 , \3064_b1 );
not ( \3065_b1 , w_9742 );
not ( \3065_b0 , w_9743 );
and ( w_9742 , w_9743 , \3064_b0 );
or ( \3066_b1 , \3063_b1 , \3065_b1 );
not ( \3065_b1 , w_9744 );
and ( \3066_b0 , \3063_b0 , w_9745 );
and ( w_9744 , w_9745 , \3065_b0 );
or ( \3067_b1 , \a[11]_b1 , \c[11]_b1 );
not ( \c[11]_b1 , w_9746 );
and ( \3067_b0 , \a[11]_b0 , w_9747 );
and ( w_9746 , w_9747 , \c[11]_b0 );
or ( \3068_b1 , \3066_b1 , w_9749 );
not ( w_9749 , w_9750 );
and ( \3068_b0 , \3066_b0 , w_9751 );
and ( w_9750 ,  , w_9751 );
buf ( w_9749 , \3067_b1 );
not ( w_9749 , w_9752 );
not (  , w_9753 );
and ( w_9752 , w_9753 , \3067_b0 );
or ( \3069_b1 , \3062_b1 , w_9755 );
not ( w_9755 , w_9756 );
and ( \3069_b0 , \3062_b0 , w_9757 );
and ( w_9756 ,  , w_9757 );
buf ( w_9755 , \3068_b1 );
not ( w_9755 , w_9758 );
not (  , w_9759 );
and ( w_9758 , w_9759 , \3068_b0 );
buf ( \3070_b1 , \3069_b1 );
not ( \3070_b1 , w_9760 );
not ( \3070_b0 , w_9761 );
and ( w_9760 , w_9761 , \3069_b0 );
or ( \3071_b1 , \3070_b1 , w_9762 );
or ( \3071_b0 , \3070_b0 , \3046_b0 );
not ( \3046_b0 , w_9763 );
and ( w_9763 , w_9762 , \3046_b1 );
or ( \3072_b1 , \a[12]_b1 , w_9765 );
not ( w_9765 , w_9766 );
and ( \3072_b0 , \a[12]_b0 , w_9767 );
and ( w_9766 ,  , w_9767 );
buf ( w_9765 , \c[12]_b1 );
not ( w_9765 , w_9768 );
not (  , w_9769 );
and ( w_9768 , w_9769 , \c[12]_b0 );
or ( \3073_b1 , \3042_b1 , w_9770 );
or ( \3073_b0 , \3042_b0 , \3072_b0 );
not ( \3072_b0 , w_9771 );
and ( w_9771 , w_9770 , \3072_b1 );
or ( \3074_b1 , \a[13]_b1 , w_9773 );
not ( w_9773 , w_9774 );
and ( \3074_b0 , \a[13]_b0 , w_9775 );
and ( w_9774 ,  , w_9775 );
buf ( w_9773 , \c[13]_b1 );
not ( w_9773 , w_9776 );
not (  , w_9777 );
and ( w_9776 , w_9777 , \c[13]_b0 );
or ( \3075_b1 , \3073_b1 , w_9779 );
not ( w_9779 , w_9780 );
and ( \3075_b0 , \3073_b0 , w_9781 );
and ( w_9780 ,  , w_9781 );
buf ( w_9779 , \3074_b1 );
not ( w_9779 , w_9782 );
not (  , w_9783 );
and ( w_9782 , w_9783 , \3074_b0 );
or ( \3076_b1 , \3075_b1 , \3045_b1 );
not ( \3045_b1 , w_9784 );
and ( \3076_b0 , \3075_b0 , w_9785 );
and ( w_9784 , w_9785 , \3045_b0 );
or ( \3077_b1 , \a[14]_b1 , \c[14]_b1 );
not ( \c[14]_b1 , w_9786 );
and ( \3077_b0 , \a[14]_b0 , w_9787 );
and ( w_9786 , w_9787 , \c[14]_b0 );
or ( \3078_b1 , \3076_b1 , w_9789 );
not ( w_9789 , w_9790 );
and ( \3078_b0 , \3076_b0 , w_9791 );
and ( w_9790 ,  , w_9791 );
buf ( w_9789 , \3077_b1 );
not ( w_9789 , w_9792 );
not (  , w_9793 );
and ( w_9792 , w_9793 , \3077_b0 );
or ( \3079_b1 , \3071_b1 , w_9795 );
not ( w_9795 , w_9796 );
and ( \3079_b0 , \3071_b0 , w_9797 );
and ( w_9796 ,  , w_9797 );
buf ( w_9795 , \3078_b1 );
not ( w_9795 , w_9798 );
not (  , w_9799 );
and ( w_9798 , w_9799 , \3078_b0 );
or ( \3080_b1 , \3055_b1 , w_9801 );
not ( w_9801 , w_9802 );
and ( \3080_b0 , \3055_b0 , w_9803 );
and ( w_9802 ,  , w_9803 );
buf ( w_9801 , \3079_b1 );
not ( w_9801 , w_9804 );
not (  , w_9805 );
and ( w_9804 , w_9805 , \3079_b0 );
buf ( \3081_b1 , \3080_b1 );
not ( \3081_b1 , w_9806 );
not ( \3081_b0 , w_9807 );
and ( w_9806 , w_9807 , \3080_b0 );
or ( \3082_b1 , \3027_b1 , w_9808 );
or ( \3082_b0 , \3027_b0 , \3081_b0 );
not ( \3081_b0 , w_9809 );
and ( w_9809 , w_9808 , \3081_b1 );
or ( \3083_b1 , \3080_b1 , w_9810 );
or ( \3083_b0 , \3080_b0 , \3026_b0 );
not ( \3026_b0 , w_9811 );
and ( w_9811 , w_9810 , \3026_b1 );
or ( \3084_b1 , \3082_b1 , w_9813 );
not ( w_9813 , w_9814 );
and ( \3084_b0 , \3082_b0 , w_9815 );
and ( w_9814 ,  , w_9815 );
buf ( w_9813 , \3083_b1 );
not ( w_9813 , w_9816 );
not (  , w_9817 );
and ( w_9816 , w_9817 , \3083_b0 );
buf ( \3085_b1 , \3084_b1 );
not ( \3085_b1 , w_9818 );
not ( \3085_b0 , w_9819 );
and ( w_9818 , w_9819 , \3084_b0 );
buf ( \3086_b1 , \1232_b1 );
not ( \3086_b1 , w_9820 );
not ( \3086_b0 , w_9821 );
and ( w_9820 , w_9821 , \1232_b0 );
buf ( \3087_b1 , \3086_b1 );
not ( \3087_b1 , w_9822 );
not ( \3087_b0 , w_9823 );
and ( w_9822 , w_9823 , \3086_b0 );
buf ( \3088_b1 , \3087_b1 );
not ( \3088_b1 , w_9824 );
not ( \3088_b0 , w_9825 );
and ( w_9824 , w_9825 , \3087_b0 );
or ( \3089_b1 , \3085_b1 , w_9826 );
or ( \3089_b0 , \3085_b0 , \3088_b0 );
not ( \3088_b0 , w_9827 );
and ( w_9827 , w_9826 , \3088_b1 );
or ( \3090_b1 , \1282_b1 , \d[15]_b1 );
not ( \d[15]_b1 , w_9828 );
and ( \3090_b0 , \1282_b0 , w_9829 );
and ( w_9828 , w_9829 , \d[15]_b0 );
or ( \3091_b1 , \1435_b1 , \c[15]_b1 );
not ( \c[15]_b1 , w_9830 );
and ( \3091_b0 , \1435_b0 , w_9831 );
and ( w_9830 , w_9831 , \c[15]_b0 );
or ( \3092_b1 , \3090_b1 , w_9833 );
not ( w_9833 , w_9834 );
and ( \3092_b0 , \3090_b0 , w_9835 );
and ( w_9834 ,  , w_9835 );
buf ( w_9833 , \3091_b1 );
not ( w_9833 , w_9836 );
not (  , w_9837 );
and ( w_9836 , w_9837 , \3091_b0 );
or ( \3093_b1 , \3089_b1 , w_9839 );
not ( w_9839 , w_9840 );
and ( \3093_b0 , \3089_b0 , w_9841 );
and ( w_9840 ,  , w_9841 );
buf ( w_9839 , \3092_b1 );
not ( w_9839 , w_9842 );
not (  , w_9843 );
and ( w_9842 , w_9843 , \3092_b0 );
or ( \3094_b1 , \3023_b1 , w_9845 );
not ( w_9845 , w_9846 );
and ( \3094_b0 , \3023_b0 , w_9847 );
and ( w_9846 ,  , w_9847 );
buf ( w_9845 , \3093_b1 );
not ( w_9845 , w_9848 );
not (  , w_9849 );
and ( w_9848 , w_9849 , \3093_b0 );
or ( \3095_b1 , \2959_b1 , w_9851 );
not ( w_9851 , w_9852 );
and ( \3095_b0 , \2959_b0 , w_9853 );
and ( w_9852 ,  , w_9853 );
buf ( w_9851 , \3094_b1 );
not ( w_9851 , w_9854 );
not (  , w_9855 );
and ( w_9854 , w_9855 , \3094_b0 );
or ( \3096_b1 , \2955_b1 , w_9857 );
not ( w_9857 , w_9858 );
and ( \3096_b0 , \2955_b0 , w_9859 );
and ( w_9858 ,  , w_9859 );
buf ( w_9857 , \3095_b1 );
not ( w_9857 , w_9860 );
not (  , w_9861 );
and ( w_9860 , w_9861 , \3095_b0 );
or ( \3097_b1 , \2953_b1 , w_9863 );
not ( w_9863 , w_9864 );
and ( \3097_b0 , \2953_b0 , w_9865 );
and ( w_9864 ,  , w_9865 );
buf ( w_9863 , \3096_b1 );
not ( w_9863 , w_9866 );
not (  , w_9867 );
and ( w_9866 , w_9867 , \3096_b0 );
buf ( \3098_b1 , \d[15]_b1 );
not ( \3098_b1 , w_9868 );
not ( \3098_b0 , w_9869 );
and ( w_9868 , w_9869 , \d[15]_b0 );
buf ( \3099_b1 , \1457_b1 );
not ( \3099_b1 , w_9870 );
not ( \3099_b0 , w_9871 );
and ( w_9870 , w_9871 , \1457_b0 );
or ( \3100_b1 , \3098_b1 , w_9872 );
or ( \3100_b0 , \3098_b0 , \3099_b0 );
not ( \3099_b0 , w_9873 );
and ( w_9873 , w_9872 , \3099_b1 );
buf ( \3101_b1 , \1316_b1 );
not ( \3101_b1 , w_9874 );
not ( \3101_b0 , w_9875 );
and ( w_9874 , w_9875 , \1316_b0 );
buf ( \3102_b1 , \3101_b1 );
not ( \3102_b1 , w_9876 );
not ( \3102_b0 , w_9877 );
and ( w_9876 , w_9877 , \3101_b0 );
or ( \3104_b1 , \3100_b1 , w_9879 );
not ( w_9879 , w_9880 );
and ( \3104_b0 , \3100_b0 , w_9881 );
and ( w_9880 ,  , w_9881 );
buf ( w_9879 , \3103_b1 );
not ( w_9879 , w_9882 );
not (  , w_9883 );
and ( w_9882 , w_9883 , \3103_b0 );
or ( \3105_b1 , \3097_b1 , w_9885 );
not ( w_9885 , w_9886 );
and ( \3105_b0 , \3097_b0 , w_9887 );
and ( w_9886 ,  , w_9887 );
buf ( w_9885 , \3104_b1 );
not ( w_9885 , w_9888 );
not (  , w_9889 );
and ( w_9888 , w_9889 , \3104_b0 );
or ( \3106_b1 , \2948_b1 , w_9891 );
not ( w_9891 , w_9892 );
and ( \3106_b0 , \2948_b0 , w_9893 );
and ( w_9892 ,  , w_9893 );
buf ( w_9891 , \3105_b1 );
not ( w_9891 , w_9894 );
not (  , w_9895 );
and ( w_9894 , w_9895 , \3105_b0 );
or ( \3107_b1 , \2938_b1 , w_9897 );
not ( w_9897 , w_9898 );
and ( \3107_b0 , \2938_b0 , w_9899 );
and ( w_9898 ,  , w_9899 );
buf ( w_9897 , \3106_b1 );
not ( w_9897 , w_9900 );
not (  , w_9901 );
and ( w_9900 , w_9901 , \3106_b0 );
buf ( \3108_b1 , \3107_b1 );
not ( \3108_b1 , w_9902 );
not ( \3108_b0 , w_9903 );
and ( w_9902 , w_9903 , \3107_b0 );
buf ( \3109_b1 , \a[11]_b1 );
not ( \3109_b1 , w_9904 );
not ( \3109_b0 , w_9905 );
and ( w_9904 , w_9905 , \a[11]_b0 );
buf ( \3110_b1 , \2940_b1 );
not ( \3110_b1 , w_9906 );
not ( \3110_b0 , w_9907 );
and ( w_9906 , w_9907 , \2940_b0 );
buf ( \3111_b1 , \3101_b1 );
not ( \3111_b1 , w_9908 );
not ( \3111_b0 , w_9909 );
and ( w_9908 , w_9909 , \3101_b0 );
or ( \3112_b1 , \3110_b1 , w_9910 );
or ( \3112_b0 , \3110_b0 , \3111_b0 );
not ( \3111_b0 , w_9911 );
and ( w_9911 , w_9910 , \3111_b1 );
buf ( \3113_b1 , \644_b1 );
not ( \3113_b1 , w_9912 );
not ( \3113_b0 , w_9913 );
and ( w_9912 , w_9913 , \644_b0 );
or ( \3114_b1 , \3112_b1 , w_9915 );
not ( w_9915 , w_9916 );
and ( \3114_b0 , \3112_b0 , w_9917 );
and ( w_9916 ,  , w_9917 );
buf ( w_9915 , \3113_b1 );
not ( w_9915 , w_9918 );
not (  , w_9919 );
and ( w_9918 , w_9919 , \3113_b0 );
buf ( \3115_b1 , \3114_b1 );
not ( \3115_b1 , w_9920 );
not ( \3115_b0 , w_9921 );
and ( w_9920 , w_9921 , \3114_b0 );
or ( \3116_b1 , \3109_b1 , w_9922 );
or ( \3116_b0 , \3109_b0 , \3115_b0 );
not ( \3115_b0 , w_9923 );
and ( w_9923 , w_9922 , \3115_b1 );
buf ( \3117_b1 , \d[11]_b1 );
not ( \3117_b1 , w_9924 );
not ( \3117_b0 , w_9925 );
and ( w_9924 , w_9925 , \d[11]_b0 );
buf ( \3118_b1 , \1450_b1 );
not ( \3118_b1 , w_9926 );
not ( \3118_b0 , w_9927 );
and ( w_9926 , w_9927 , \1450_b0 );
or ( \3119_b1 , \3117_b1 , w_9928 );
or ( \3119_b0 , \3117_b0 , \3118_b0 );
not ( \3118_b0 , w_9929 );
and ( w_9929 , w_9928 , \3118_b1 );
or ( \3121_b1 , \3119_b1 , w_9931 );
not ( w_9931 , w_9932 );
and ( \3121_b0 , \3119_b0 , w_9933 );
and ( w_9932 ,  , w_9933 );
buf ( w_9931 , \3120_b1 );
not ( w_9931 , w_9934 );
not (  , w_9935 );
and ( w_9934 , w_9935 , \3120_b0 );
buf ( \3122_b1 , \b[11]_b1 );
not ( \3122_b1 , w_9936 );
not ( \3122_b0 , w_9937 );
and ( w_9936 , w_9937 , \b[11]_b0 );
buf ( \3123_b1 , \671_b1 );
not ( \3123_b1 , w_9938 );
not ( \3123_b0 , w_9939 );
and ( w_9938 , w_9939 , \671_b0 );
or ( \3124_b1 , \3123_b1 , w_9941 );
not ( w_9941 , w_9942 );
and ( \3124_b0 , \3123_b0 , w_9943 );
and ( w_9942 ,  , w_9943 );
buf ( w_9941 , \1324_b1 );
not ( w_9941 , w_9944 );
not (  , w_9945 );
and ( w_9944 , w_9945 , \1324_b0 );
buf ( \3125_b1 , \3124_b1 );
not ( \3125_b1 , w_9946 );
not ( \3125_b0 , w_9947 );
and ( w_9946 , w_9947 , \3124_b0 );
or ( \3126_b1 , \3122_b1 , w_9948 );
or ( \3126_b0 , \3122_b0 , \3125_b0 );
not ( \3125_b0 , w_9949 );
and ( w_9949 , w_9948 , \3125_b1 );
buf ( \3127_b1 , \a[11]_b1 );
not ( \3127_b1 , w_9950 );
not ( \3127_b0 , w_9951 );
and ( w_9950 , w_9951 , \a[11]_b0 );
buf ( \3128_b1 , \672_b1 );
not ( \3128_b1 , w_9952 );
not ( \3128_b0 , w_9953 );
and ( w_9952 , w_9953 , \672_b0 );
or ( \3129_b1 , \3127_b1 , w_9954 );
or ( \3129_b0 , \3127_b0 , \3128_b0 );
not ( \3128_b0 , w_9955 );
and ( w_9955 , w_9954 , \3128_b1 );
or ( \3130_b1 , \c[11]_b1 , \d[11]_b1 );
xor ( \3130_b0 , \c[11]_b0 , w_9956 );
not ( w_9956 , w_9957 );
and ( w_9957 , \d[11]_b1 , \d[11]_b0 );
or ( \3131_b1 , \3130_b1 , \925_b1 );
not ( \925_b1 , w_9958 );
and ( \3131_b0 , \3130_b0 , w_9959 );
and ( w_9958 , w_9959 , \925_b0 );
or ( \3132_b1 , \2986_b1 , w_9961 );
not ( w_9961 , w_9962 );
and ( \3132_b0 , \2986_b0 , w_9963 );
and ( w_9962 ,  , w_9963 );
buf ( w_9961 , \3005_b1 );
not ( w_9961 , w_9964 );
not (  , w_9965 );
and ( w_9964 , w_9965 , \3005_b0 );
buf ( \3133_b1 , \3132_b1 );
not ( \3133_b1 , w_9966 );
not ( \3133_b0 , w_9967 );
and ( w_9966 , w_9967 , \3132_b0 );
buf ( \3134_b1 , \2987_b1 );
not ( \3134_b1 , w_9968 );
not ( \3134_b0 , w_9969 );
and ( w_9968 , w_9969 , \2987_b0 );
buf ( \3136_b1 , \3134_b1 );
not ( \3136_b1 , w_9970 );
not ( \3136_b0 , w_9971 );
and ( w_9970 , w_9971 , \3134_b0 );
buf ( \3137_b1 , \2997_b1 );
not ( \3137_b1 , w_9972 );
not ( \3137_b0 , w_9973 );
and ( w_9972 , w_9973 , \2997_b0 );
or ( \3138_b1 , \3136_b1 , w_9974 );
or ( \3138_b0 , \3136_b0 , \3137_b0 );
not ( \3137_b0 , w_9975 );
and ( w_9975 , w_9974 , \3137_b1 );
or ( \3139_b1 , \3138_b1 , w_9977 );
not ( w_9977 , w_9978 );
and ( \3139_b0 , \3138_b0 , w_9979 );
and ( w_9978 ,  , w_9979 );
buf ( w_9977 , \3002_b1 );
not ( w_9977 , w_9980 );
not (  , w_9981 );
and ( w_9980 , w_9981 , \3002_b0 );
or ( \3140_b1 , \3135_b1 , w_9983 );
not ( w_9983 , w_9984 );
and ( \3140_b0 , \3135_b0 , w_9985 );
and ( w_9984 ,  , w_9985 );
buf ( w_9983 , \3139_b1 );
not ( w_9983 , w_9986 );
not (  , w_9987 );
and ( w_9986 , w_9987 , \3139_b0 );
buf ( \3141_b1 , \3140_b1 );
not ( \3141_b1 , w_9988 );
not ( \3141_b0 , w_9989 );
and ( w_9988 , w_9989 , \3140_b0 );
or ( \3142_b1 , \3133_b1 , w_9990 );
or ( \3142_b0 , \3133_b0 , \3141_b0 );
not ( \3141_b0 , w_9991 );
and ( w_9991 , w_9990 , \3141_b1 );
or ( \3143_b1 , \3140_b1 , w_9992 );
or ( \3143_b0 , \3140_b0 , \3132_b0 );
not ( \3132_b0 , w_9993 );
and ( w_9993 , w_9992 , \3132_b1 );
or ( \3144_b1 , \3142_b1 , w_9995 );
not ( w_9995 , w_9996 );
and ( \3144_b0 , \3142_b0 , w_9997 );
and ( w_9996 ,  , w_9997 );
buf ( w_9995 , \3143_b1 );
not ( w_9995 , w_9998 );
not (  , w_9999 );
and ( w_9998 , w_9999 , \3143_b0 );
buf ( \3145_b1 , \3144_b1 );
not ( \3145_b1 , w_10000 );
not ( \3145_b0 , w_10001 );
and ( w_10000 , w_10001 , \3144_b0 );
buf ( \3146_b1 , \2961_b1 );
not ( \3146_b1 , w_10002 );
not ( \3146_b0 , w_10003 );
and ( w_10002 , w_10003 , \2961_b0 );
or ( \3147_b1 , \3145_b1 , w_10004 );
or ( \3147_b0 , \3145_b0 , \3146_b0 );
not ( \3146_b0 , w_10005 );
and ( w_10005 , w_10004 , \3146_b1 );
or ( \3148_b1 , \3048_b1 , w_10007 );
not ( w_10007 , w_10008 );
and ( \3148_b0 , \3048_b0 , w_10009 );
and ( w_10008 ,  , w_10009 );
buf ( w_10007 , \3067_b1 );
not ( w_10007 , w_10010 );
not (  , w_10011 );
and ( w_10010 , w_10011 , \3067_b0 );
buf ( \3149_b1 , \3148_b1 );
not ( \3149_b1 , w_10012 );
not ( \3149_b0 , w_10013 );
and ( w_10012 , w_10013 , \3148_b0 );
buf ( \3150_b1 , \3049_b1 );
not ( \3150_b1 , w_10014 );
not ( \3150_b0 , w_10015 );
and ( w_10014 , w_10015 , \3049_b0 );
buf ( \3152_b1 , \3150_b1 );
not ( \3152_b1 , w_10016 );
not ( \3152_b0 , w_10017 );
and ( w_10016 , w_10017 , \3150_b0 );
buf ( \3153_b1 , \3059_b1 );
not ( \3153_b1 , w_10018 );
not ( \3153_b0 , w_10019 );
and ( w_10018 , w_10019 , \3059_b0 );
or ( \3154_b1 , \3152_b1 , w_10020 );
or ( \3154_b0 , \3152_b0 , \3153_b0 );
not ( \3153_b0 , w_10021 );
and ( w_10021 , w_10020 , \3153_b1 );
or ( \3155_b1 , \3154_b1 , w_10023 );
not ( w_10023 , w_10024 );
and ( \3155_b0 , \3154_b0 , w_10025 );
and ( w_10024 ,  , w_10025 );
buf ( w_10023 , \3064_b1 );
not ( w_10023 , w_10026 );
not (  , w_10027 );
and ( w_10026 , w_10027 , \3064_b0 );
or ( \3156_b1 , \3151_b1 , w_10029 );
not ( w_10029 , w_10030 );
and ( \3156_b0 , \3151_b0 , w_10031 );
and ( w_10030 ,  , w_10031 );
buf ( w_10029 , \3155_b1 );
not ( w_10029 , w_10032 );
not (  , w_10033 );
and ( w_10032 , w_10033 , \3155_b0 );
buf ( \3157_b1 , \3156_b1 );
not ( \3157_b1 , w_10034 );
not ( \3157_b0 , w_10035 );
and ( w_10034 , w_10035 , \3156_b0 );
or ( \3158_b1 , \3149_b1 , w_10036 );
or ( \3158_b0 , \3149_b0 , \3157_b0 );
not ( \3157_b0 , w_10037 );
and ( w_10037 , w_10036 , \3157_b1 );
or ( \3159_b1 , \3156_b1 , w_10038 );
or ( \3159_b0 , \3156_b0 , \3148_b0 );
not ( \3148_b0 , w_10039 );
and ( w_10039 , w_10038 , \3148_b1 );
or ( \3160_b1 , \3158_b1 , w_10041 );
not ( w_10041 , w_10042 );
and ( \3160_b0 , \3158_b0 , w_10043 );
and ( w_10042 ,  , w_10043 );
buf ( w_10041 , \3159_b1 );
not ( w_10041 , w_10044 );
not (  , w_10045 );
and ( w_10044 , w_10045 , \3159_b0 );
or ( \3161_b1 , \3087_b1 , \3160_b1 );
not ( \3160_b1 , w_10046 );
and ( \3161_b0 , \3087_b0 , w_10047 );
and ( w_10046 , w_10047 , \3160_b0 );
buf ( \3162_b1 , \d[11]_b1 );
not ( \3162_b1 , w_10048 );
not ( \3162_b0 , w_10049 );
and ( w_10048 , w_10049 , \d[11]_b0 );
buf ( \3163_b1 , \1282_b1 );
not ( \3163_b1 , w_10050 );
not ( \3163_b0 , w_10051 );
and ( w_10050 , w_10051 , \1282_b0 );
or ( \3164_b1 , \3162_b1 , w_10052 );
or ( \3164_b0 , \3162_b0 , \3163_b0 );
not ( \3163_b0 , w_10053 );
and ( w_10053 , w_10052 , \3163_b1 );
or ( \3165_b1 , \1435_b1 , w_10055 );
not ( w_10055 , w_10056 );
and ( \3165_b0 , \1435_b0 , w_10057 );
and ( w_10056 ,  , w_10057 );
buf ( w_10055 , \c[11]_b1 );
not ( w_10055 , w_10058 );
not (  , w_10059 );
and ( w_10058 , w_10059 , \c[11]_b0 );
or ( \3166_b1 , \3164_b1 , w_10061 );
not ( w_10061 , w_10062 );
and ( \3166_b0 , \3164_b0 , w_10063 );
and ( w_10062 ,  , w_10063 );
buf ( w_10061 , \3165_b1 );
not ( w_10061 , w_10064 );
not (  , w_10065 );
and ( w_10064 , w_10065 , \3165_b0 );
or ( \3167_b1 , \3161_b1 , w_10067 );
not ( w_10067 , w_10068 );
and ( \3167_b0 , \3161_b0 , w_10069 );
and ( w_10068 ,  , w_10069 );
buf ( w_10067 , \3166_b1 );
not ( w_10067 , w_10070 );
not (  , w_10071 );
and ( w_10070 , w_10071 , \3166_b0 );
or ( \3168_b1 , \3147_b1 , w_10073 );
not ( w_10073 , w_10074 );
and ( \3168_b0 , \3147_b0 , w_10075 );
and ( w_10074 ,  , w_10075 );
buf ( w_10073 , \3167_b1 );
not ( w_10073 , w_10076 );
not (  , w_10077 );
and ( w_10076 , w_10077 , \3167_b0 );
or ( \3169_b1 , \3131_b1 , w_10079 );
not ( w_10079 , w_10080 );
and ( \3169_b0 , \3131_b0 , w_10081 );
and ( w_10080 ,  , w_10081 );
buf ( w_10079 , \3168_b1 );
not ( w_10079 , w_10082 );
not (  , w_10083 );
and ( w_10082 , w_10083 , \3168_b0 );
or ( \3170_b1 , \3129_b1 , w_10085 );
not ( w_10085 , w_10086 );
and ( \3170_b0 , \3129_b0 , w_10087 );
and ( w_10086 ,  , w_10087 );
buf ( w_10085 , \3169_b1 );
not ( w_10085 , w_10088 );
not (  , w_10089 );
and ( w_10088 , w_10089 , \3169_b0 );
buf ( \3171_b1 , \3170_b1 );
not ( \3171_b1 , w_10090 );
not ( \3171_b0 , w_10091 );
and ( w_10090 , w_10091 , \3170_b0 );
or ( \3172_b1 , \3126_b1 , w_10093 );
not ( w_10093 , w_10094 );
and ( \3172_b0 , \3126_b0 , w_10095 );
and ( w_10094 ,  , w_10095 );
buf ( w_10093 , \3171_b1 );
not ( w_10093 , w_10096 );
not (  , w_10097 );
and ( w_10096 , w_10097 , \3171_b0 );
or ( \3173_b1 , \3121_b1 , w_10099 );
not ( w_10099 , w_10100 );
and ( \3173_b0 , \3121_b0 , w_10101 );
and ( w_10100 ,  , w_10101 );
buf ( w_10099 , \3172_b1 );
not ( w_10099 , w_10102 );
not (  , w_10103 );
and ( w_10102 , w_10103 , \3172_b0 );
or ( \3174_b1 , \3116_b1 , w_10105 );
not ( w_10105 , w_10106 );
and ( \3174_b0 , \3116_b0 , w_10107 );
and ( w_10106 ,  , w_10107 );
buf ( w_10105 , \3173_b1 );
not ( w_10105 , w_10108 );
not (  , w_10109 );
and ( w_10108 , w_10109 , \3173_b0 );
buf ( \3175_b1 , \1529_b1 );
not ( \3175_b1 , w_10110 );
not ( \3175_b0 , w_10111 );
and ( w_10110 , w_10111 , \1529_b0 );
buf ( \3176_b1 , \2211_b1 );
not ( \3176_b1 , w_10112 );
not ( \3176_b0 , w_10113 );
and ( w_10112 , w_10113 , \2211_b0 );
or ( \3177_b1 , \3176_b1 , w_10115 );
not ( w_10115 , w_10116 );
and ( \3177_b0 , \3176_b0 , w_10117 );
and ( w_10116 ,  , w_10117 );
buf ( w_10115 , \2112_b1 );
not ( w_10115 , w_10118 );
not (  , w_10119 );
and ( w_10118 , w_10119 , \2112_b0 );
buf ( \3178_b1 , \3177_b1 );
not ( \3178_b1 , w_10120 );
not ( \3178_b0 , w_10121 );
and ( w_10120 , w_10121 , \3177_b0 );
buf ( \3179_b1 , \2206_b1 );
not ( \3179_b1 , w_10122 );
not ( \3179_b0 , w_10123 );
and ( w_10122 , w_10123 , \2206_b0 );
buf ( \3180_b1 , \2173_b1 );
not ( \3180_b1 , w_10124 );
not ( \3180_b0 , w_10125 );
and ( w_10124 , w_10125 , \2173_b0 );
buf ( \3181_b1 , \2120_b1 );
not ( \3181_b1 , w_10126 );
not ( \3181_b0 , w_10127 );
and ( w_10126 , w_10127 , \2120_b0 );
or ( \3182_b1 , \3180_b1 , w_10128 );
or ( \3182_b0 , \3180_b0 , \3181_b0 );
not ( \3181_b0 , w_10129 );
and ( w_10129 , w_10128 , \3181_b1 );
buf ( \3183_b1 , \2191_b1 );
not ( \3183_b1 , w_10130 );
not ( \3183_b0 , w_10131 );
and ( w_10130 , w_10131 , \2191_b0 );
or ( \3184_b1 , \3182_b1 , w_10133 );
not ( w_10133 , w_10134 );
and ( \3184_b0 , \3182_b0 , w_10135 );
and ( w_10134 ,  , w_10135 );
buf ( w_10133 , \3183_b1 );
not ( w_10133 , w_10136 );
not (  , w_10137 );
and ( w_10136 , w_10137 , \3183_b0 );
buf ( \3185_b1 , \3184_b1 );
not ( \3185_b1 , w_10138 );
not ( \3185_b0 , w_10139 );
and ( w_10138 , w_10139 , \3184_b0 );
or ( \3186_b1 , \3179_b1 , w_10140 );
or ( \3186_b0 , \3179_b0 , \3185_b0 );
not ( \3185_b0 , w_10141 );
and ( w_10141 , w_10140 , \3185_b1 );
buf ( \3187_b1 , \2187_b1 );
not ( \3187_b1 , w_10142 );
not ( \3187_b0 , w_10143 );
and ( w_10142 , w_10143 , \2187_b0 );
or ( \3188_b1 , \3186_b1 , w_10145 );
not ( w_10145 , w_10146 );
and ( \3188_b0 , \3186_b0 , w_10147 );
and ( w_10146 ,  , w_10147 );
buf ( w_10145 , \3187_b1 );
not ( w_10145 , w_10148 );
not (  , w_10149 );
and ( w_10148 , w_10149 , \3187_b0 );
buf ( \3189_b1 , \3188_b1 );
not ( \3189_b1 , w_10150 );
not ( \3189_b0 , w_10151 );
and ( w_10150 , w_10151 , \3188_b0 );
or ( \3190_b1 , \3178_b1 , w_10152 );
or ( \3190_b0 , \3178_b0 , \3189_b0 );
not ( \3189_b0 , w_10153 );
and ( w_10153 , w_10152 , \3189_b1 );
or ( \3191_b1 , \3188_b1 , w_10154 );
or ( \3191_b0 , \3188_b0 , \3177_b0 );
not ( \3177_b0 , w_10155 );
and ( w_10155 , w_10154 , \3177_b1 );
or ( \3192_b1 , \3190_b1 , w_10157 );
not ( w_10157 , w_10158 );
and ( \3192_b0 , \3190_b0 , w_10159 );
and ( w_10158 ,  , w_10159 );
buf ( w_10157 , \3191_b1 );
not ( w_10157 , w_10160 );
not (  , w_10161 );
and ( w_10160 , w_10161 , \3191_b0 );
buf ( \3193_b1 , \3192_b1 );
not ( \3193_b1 , w_10162 );
not ( \3193_b0 , w_10163 );
and ( w_10162 , w_10163 , \3192_b0 );
or ( \3194_b1 , \3175_b1 , w_10164 );
or ( \3194_b0 , \3175_b0 , \3193_b0 );
not ( \3193_b0 , w_10165 );
and ( w_10165 , w_10164 , \3193_b1 );
buf ( \3195_b1 , \2814_b1 );
not ( \3195_b1 , w_10166 );
not ( \3195_b0 , w_10167 );
and ( w_10166 , w_10167 , \2814_b0 );
or ( \3196_b1 , \3195_b1 , w_10169 );
not ( w_10169 , w_10170 );
and ( \3196_b0 , \3195_b0 , w_10171 );
and ( w_10170 ,  , w_10171 );
buf ( w_10169 , \2914_b1 );
not ( w_10169 , w_10172 );
not (  , w_10173 );
and ( w_10172 , w_10173 , \2914_b0 );
buf ( \3197_b1 , \2866_b1 );
not ( \3197_b1 , w_10174 );
not ( \3197_b0 , w_10175 );
and ( w_10174 , w_10175 , \2866_b0 );
buf ( \3198_b1 , \2907_b1 );
not ( \3198_b1 , w_10176 );
not ( \3198_b0 , w_10177 );
and ( w_10176 , w_10177 , \2907_b0 );
or ( \3199_b1 , \3198_b1 , w_10179 );
not ( w_10179 , w_10180 );
and ( \3199_b0 , \3198_b0 , w_10181 );
and ( w_10180 ,  , w_10181 );
buf ( w_10179 , \2901_b1 );
not ( w_10179 , w_10182 );
not (  , w_10183 );
and ( w_10182 , w_10183 , \2901_b0 );
buf ( \3200_b1 , \3199_b1 );
not ( \3200_b1 , w_10184 );
not ( \3200_b0 , w_10185 );
and ( w_10184 , w_10185 , \3199_b0 );
or ( \3201_b1 , \3197_b1 , w_10186 );
or ( \3201_b0 , \3197_b0 , \3200_b0 );
not ( \3200_b0 , w_10187 );
and ( w_10187 , w_10186 , \3200_b1 );
buf ( \3202_b1 , \2908_b1 );
not ( \3202_b1 , w_10188 );
not ( \3202_b0 , w_10189 );
and ( w_10188 , w_10189 , \2908_b0 );
or ( \3203_b1 , \3201_b1 , w_10191 );
not ( w_10191 , w_10192 );
and ( \3203_b0 , \3201_b0 , w_10193 );
and ( w_10192 ,  , w_10193 );
buf ( w_10191 , \3202_b1 );
not ( w_10191 , w_10194 );
not (  , w_10195 );
and ( w_10194 , w_10195 , \3202_b0 );
or ( \3204_b1 , \3196_b1 , \3203_b1 );
xor ( \3204_b0 , \3196_b0 , w_10196 );
not ( w_10196 , w_10197 );
and ( w_10197 , \3203_b1 , \3203_b0 );
or ( \3205_b1 , \3204_b1 , w_10199 );
not ( w_10199 , w_10200 );
and ( \3205_b0 , \3204_b0 , w_10201 );
and ( w_10200 ,  , w_10201 );
buf ( w_10199 , \2936_b1 );
not ( w_10199 , w_10202 );
not (  , w_10203 );
and ( w_10202 , w_10203 , \2936_b0 );
or ( \3206_b1 , \3194_b1 , w_10205 );
not ( w_10205 , w_10206 );
and ( \3206_b0 , \3194_b0 , w_10207 );
and ( w_10206 ,  , w_10207 );
buf ( w_10205 , \3205_b1 );
not ( w_10205 , w_10208 );
not (  , w_10209 );
and ( w_10208 , w_10209 , \3205_b0 );
or ( \3207_b1 , \3174_b1 , w_10211 );
not ( w_10211 , w_10212 );
and ( \3207_b0 , \3174_b0 , w_10213 );
and ( w_10212 ,  , w_10213 );
buf ( w_10211 , \3206_b1 );
not ( w_10211 , w_10214 );
not (  , w_10215 );
and ( w_10214 , w_10215 , \3206_b0 );
buf ( \3208_b1 , \3207_b1 );
not ( \3208_b1 , w_10216 );
not ( \3208_b0 , w_10217 );
and ( w_10216 , w_10217 , \3207_b0 );
buf ( \3209_b1 , \a[6]_b1 );
not ( \3209_b1 , w_10218 );
not ( \3209_b0 , w_10219 );
and ( w_10218 , w_10219 , \a[6]_b0 );
buf ( \3210_b1 , \3114_b1 );
not ( \3210_b1 , w_10220 );
not ( \3210_b0 , w_10221 );
and ( w_10220 , w_10221 , \3114_b0 );
or ( \3211_b1 , \3209_b1 , w_10222 );
or ( \3211_b0 , \3209_b0 , \3210_b0 );
not ( \3210_b0 , w_10223 );
and ( w_10223 , w_10222 , \3210_b1 );
or ( \3212_b1 , \d[6]_b1 , \1342_b1 );
not ( \1342_b1 , w_10224 );
and ( \3212_b0 , \d[6]_b0 , w_10225 );
and ( w_10224 , w_10225 , \1342_b0 );
or ( \3214_b1 , \a[6]_b1 , w_10226 );
or ( \3214_b0 , \a[6]_b0 , \b[6]_b0 );
not ( \b[6]_b0 , w_10227 );
and ( w_10227 , w_10226 , \b[6]_b1 );
or ( \3215_b1 , \3214_b1 , w_10229 );
not ( w_10229 , w_10230 );
and ( \3215_b0 , \3214_b0 , w_10231 );
and ( w_10230 ,  , w_10231 );
buf ( w_10229 , \672_b1 );
not ( w_10229 , w_10232 );
not (  , w_10233 );
and ( w_10232 , w_10233 , \672_b0 );
or ( \3216_b1 , \c[6]_b1 , \d[6]_b1 );
xor ( \3216_b0 , \c[6]_b0 , w_10234 );
not ( w_10234 , w_10235 );
and ( w_10235 , \d[6]_b1 , \d[6]_b0 );
buf ( \3217_b1 , \3216_b1 );
not ( \3217_b1 , w_10236 );
not ( \3217_b0 , w_10237 );
and ( w_10236 , w_10237 , \3216_b0 );
buf ( \3218_b1 , \1320_b1 );
not ( \3218_b1 , w_10238 );
not ( \3218_b0 , w_10239 );
and ( w_10238 , w_10239 , \1320_b0 );
or ( \3219_b1 , \3217_b1 , w_10240 );
or ( \3219_b0 , \3217_b0 , \3218_b0 );
not ( \3218_b0 , w_10241 );
and ( w_10241 , w_10240 , \3218_b1 );
buf ( \3220_b1 , \1090_b1 );
not ( \3220_b1 , w_10242 );
not ( \3220_b0 , w_10243 );
and ( w_10242 , w_10243 , \1090_b0 );
or ( \3221_b1 , \3220_b1 , w_10245 );
not ( w_10245 , w_10246 );
and ( \3221_b0 , \3220_b0 , w_10247 );
and ( w_10246 ,  , w_10247 );
buf ( w_10245 , \1095_b1 );
not ( w_10245 , w_10248 );
not (  , w_10249 );
and ( w_10248 , w_10249 , \1095_b0 );
buf ( \3222_b1 , \3221_b1 );
not ( \3222_b1 , w_10250 );
not ( \3222_b0 , w_10251 );
and ( w_10250 , w_10251 , \3221_b0 );
or ( \3223_b1 , \1097_b1 , w_10253 );
not ( w_10253 , w_10254 );
and ( \3223_b0 , \1097_b0 , w_10255 );
and ( w_10254 ,  , w_10255 );
buf ( w_10253 , \1008_b1 );
not ( w_10253 , w_10256 );
not (  , w_10257 );
and ( w_10256 , w_10257 , \1008_b0 );
buf ( \3224_b1 , \3223_b1 );
not ( \3224_b1 , w_10258 );
not ( \3224_b0 , w_10259 );
and ( w_10258 , w_10259 , \3223_b0 );
or ( \3225_b1 , \3222_b1 , w_10260 );
or ( \3225_b0 , \3222_b0 , \3224_b0 );
not ( \3224_b0 , w_10261 );
and ( w_10261 , w_10260 , \3224_b1 );
or ( \3226_b1 , \3223_b1 , w_10262 );
or ( \3226_b0 , \3223_b0 , \3221_b0 );
not ( \3221_b0 , w_10263 );
and ( w_10263 , w_10262 , \3221_b1 );
or ( \3227_b1 , \3225_b1 , w_10265 );
not ( w_10265 , w_10266 );
and ( \3227_b0 , \3225_b0 , w_10267 );
and ( w_10266 ,  , w_10267 );
buf ( w_10265 , \3226_b1 );
not ( w_10265 , w_10268 );
not (  , w_10269 );
and ( w_10268 , w_10269 , \3226_b0 );
or ( \3228_b1 , \3227_b1 , \1353_b1 );
not ( \1353_b1 , w_10270 );
and ( \3228_b0 , \3227_b0 , w_10271 );
and ( w_10270 , w_10271 , \1353_b0 );
buf ( \3229_b1 , \1193_b1 );
not ( \3229_b1 , w_10272 );
not ( \3229_b0 , w_10273 );
and ( w_10272 , w_10273 , \1193_b0 );
buf ( \3230_b1 , \3229_b1 );
not ( \3230_b1 , w_10274 );
not ( \3230_b0 , w_10275 );
and ( w_10274 , w_10275 , \3229_b0 );
buf ( \3231_b1 , \1189_b1 );
not ( \3231_b1 , w_10276 );
not ( \3231_b0 , w_10277 );
and ( w_10276 , w_10277 , \1189_b0 );
or ( \3232_b1 , \3230_b1 , w_10278 );
or ( \3232_b0 , \3230_b0 , \3231_b0 );
not ( \3231_b0 , w_10279 );
and ( w_10279 , w_10278 , \3231_b1 );
buf ( \3233_b1 , \1201_b1 );
not ( \3233_b1 , w_10280 );
not ( \3233_b0 , w_10281 );
and ( w_10280 , w_10281 , \1201_b0 );
or ( \3234_b1 , \3232_b1 , w_10283 );
not ( w_10283 , w_10284 );
and ( \3234_b0 , \3232_b0 , w_10285 );
and ( w_10284 ,  , w_10285 );
buf ( w_10283 , \3233_b1 );
not ( w_10283 , w_10286 );
not (  , w_10287 );
and ( w_10286 , w_10287 , \3233_b0 );
or ( \3235_b1 , \1202_b1 , w_10289 );
not ( w_10289 , w_10290 );
and ( \3235_b0 , \1202_b0 , w_10291 );
and ( w_10290 ,  , w_10291 );
buf ( w_10289 , \1204_b1 );
not ( w_10289 , w_10292 );
not (  , w_10293 );
and ( w_10292 , w_10293 , \1204_b0 );
or ( \3236_b1 , \3234_b1 , w_10294 );
xor ( \3236_b0 , \3234_b0 , w_10296 );
not ( w_10296 , w_10297 );
and ( w_10297 , w_10294 , w_10295 );
buf ( w_10294 , \3235_b1 );
not ( w_10294 , w_10298 );
not ( w_10295 , w_10299 );
and ( w_10298 , w_10299 , \3235_b0 );
buf ( \3237_b1 , \3236_b1 );
not ( \3237_b1 , w_10300 );
not ( \3237_b0 , w_10301 );
and ( w_10300 , w_10301 , \3236_b0 );
buf ( \3238_b1 , \1220_b1 );
not ( \3238_b1 , w_10302 );
not ( \3238_b0 , w_10303 );
and ( w_10302 , w_10303 , \1220_b0 );
or ( \3239_b1 , \3237_b1 , w_10304 );
or ( \3239_b0 , \3237_b0 , \3238_b0 );
not ( \3238_b0 , w_10305 );
and ( w_10305 , w_10304 , \3238_b1 );
buf ( \3240_b1 , \1256_b1 );
not ( \3240_b1 , w_10306 );
not ( \3240_b0 , w_10307 );
and ( w_10306 , w_10307 , \1256_b0 );
buf ( \3241_b1 , \3240_b1 );
not ( \3241_b1 , w_10308 );
not ( \3241_b0 , w_10309 );
and ( w_10308 , w_10309 , \3240_b0 );
buf ( \3242_b1 , \1252_b1 );
not ( \3242_b1 , w_10310 );
not ( \3242_b0 , w_10311 );
and ( w_10310 , w_10311 , \1252_b0 );
or ( \3243_b1 , \3241_b1 , w_10312 );
or ( \3243_b0 , \3241_b0 , \3242_b0 );
not ( \3242_b0 , w_10313 );
and ( w_10313 , w_10312 , \3242_b1 );
buf ( \3244_b1 , \1264_b1 );
not ( \3244_b1 , w_10314 );
not ( \3244_b0 , w_10315 );
and ( w_10314 , w_10315 , \1264_b0 );
or ( \3245_b1 , \3243_b1 , w_10317 );
not ( w_10317 , w_10318 );
and ( \3245_b0 , \3243_b0 , w_10319 );
and ( w_10318 ,  , w_10319 );
buf ( w_10317 , \3244_b1 );
not ( w_10317 , w_10320 );
not (  , w_10321 );
and ( w_10320 , w_10321 , \3244_b0 );
or ( \3246_b1 , \1265_b1 , w_10323 );
not ( w_10323 , w_10324 );
and ( \3246_b0 , \1265_b0 , w_10325 );
and ( w_10324 ,  , w_10325 );
buf ( w_10323 , \1267_b1 );
not ( w_10323 , w_10326 );
not (  , w_10327 );
and ( w_10326 , w_10327 , \1267_b0 );
or ( \3247_b1 , \3245_b1 , w_10328 );
xor ( \3247_b0 , \3245_b0 , w_10330 );
not ( w_10330 , w_10331 );
and ( w_10331 , w_10328 , w_10329 );
buf ( w_10328 , \3246_b1 );
not ( w_10328 , w_10332 );
not ( w_10329 , w_10333 );
and ( w_10332 , w_10333 , \3246_b0 );
buf ( \3248_b1 , \3247_b1 );
not ( \3248_b1 , w_10334 );
not ( \3248_b0 , w_10335 );
and ( w_10334 , w_10335 , \3247_b0 );
buf ( \3249_b1 , \1232_b1 );
not ( \3249_b1 , w_10336 );
not ( \3249_b0 , w_10337 );
and ( w_10336 , w_10337 , \1232_b0 );
or ( \3250_b1 , \3248_b1 , w_10338 );
or ( \3250_b0 , \3248_b0 , \3249_b0 );
not ( \3249_b0 , w_10339 );
and ( w_10339 , w_10338 , \3249_b1 );
or ( \3251_b1 , \1280_b1 , \d[6]_b1 );
not ( \d[6]_b1 , w_10340 );
and ( \3251_b0 , \1280_b0 , w_10341 );
and ( w_10340 , w_10341 , \d[6]_b0 );
buf ( \3252_b1 , \c[6]_b1 );
not ( \3252_b1 , w_10342 );
not ( \3252_b0 , w_10343 );
and ( w_10342 , w_10343 , \c[6]_b0 );
buf ( \3253_b1 , \1287_b1 );
not ( \3253_b1 , w_10344 );
not ( \3253_b0 , w_10345 );
and ( w_10344 , w_10345 , \1287_b0 );
or ( \3254_b1 , \3252_b1 , w_10346 );
or ( \3254_b0 , \3252_b0 , \3253_b0 );
not ( \3253_b0 , w_10347 );
and ( w_10347 , w_10346 , \3253_b1 );
or ( \3255_b1 , \1293_b1 , w_10349 );
not ( w_10349 , w_10350 );
and ( \3255_b0 , \1293_b0 , w_10351 );
and ( w_10350 ,  , w_10351 );
buf ( w_10349 , \b[6]_b1 );
not ( w_10349 , w_10352 );
not (  , w_10353 );
and ( w_10352 , w_10353 , \b[6]_b0 );
or ( \3256_b1 , \3254_b1 , w_10355 );
not ( w_10355 , w_10356 );
and ( \3256_b0 , \3254_b0 , w_10357 );
and ( w_10356 ,  , w_10357 );
buf ( w_10355 , \3255_b1 );
not ( w_10355 , w_10358 );
not (  , w_10359 );
and ( w_10358 , w_10359 , \3255_b0 );
or ( \3257_b1 , \3251_b1 , w_10361 );
not ( w_10361 , w_10362 );
and ( \3257_b0 , \3251_b0 , w_10363 );
and ( w_10362 ,  , w_10363 );
buf ( w_10361 , \3256_b1 );
not ( w_10361 , w_10364 );
not (  , w_10365 );
and ( w_10364 , w_10365 , \3256_b0 );
or ( \3258_b1 , \3250_b1 , w_10367 );
not ( w_10367 , w_10368 );
and ( \3258_b0 , \3250_b0 , w_10369 );
and ( w_10368 ,  , w_10369 );
buf ( w_10367 , \3257_b1 );
not ( w_10367 , w_10370 );
not (  , w_10371 );
and ( w_10370 , w_10371 , \3257_b0 );
buf ( \3259_b1 , \3258_b1 );
not ( \3259_b1 , w_10372 );
not ( \3259_b0 , w_10373 );
and ( w_10372 , w_10373 , \3258_b0 );
or ( \3260_b1 , \3239_b1 , w_10375 );
not ( w_10375 , w_10376 );
and ( \3260_b0 , \3239_b0 , w_10377 );
and ( w_10376 ,  , w_10377 );
buf ( w_10375 , \3259_b1 );
not ( w_10375 , w_10378 );
not (  , w_10379 );
and ( w_10378 , w_10379 , \3259_b0 );
or ( \3261_b1 , \3228_b1 , w_10381 );
not ( w_10381 , w_10382 );
and ( \3261_b0 , \3228_b0 , w_10383 );
and ( w_10382 ,  , w_10383 );
buf ( w_10381 , \3260_b1 );
not ( w_10381 , w_10384 );
not (  , w_10385 );
and ( w_10384 , w_10385 , \3260_b0 );
or ( \3262_b1 , \3219_b1 , w_10387 );
not ( w_10387 , w_10388 );
and ( \3262_b0 , \3219_b0 , w_10389 );
and ( w_10388 ,  , w_10389 );
buf ( w_10387 , \3261_b1 );
not ( w_10387 , w_10390 );
not (  , w_10391 );
and ( w_10390 , w_10391 , \3261_b0 );
buf ( \3263_b1 , \916_b1 );
not ( \3263_b1 , w_10392 );
not ( \3263_b0 , w_10393 );
and ( w_10392 , w_10393 , \916_b0 );
buf ( \3264_b1 , \895_b1 );
not ( \3264_b1 , w_10394 );
not ( \3264_b0 , w_10395 );
and ( w_10394 , w_10395 , \895_b0 );
or ( \3265_b1 , \3264_b1 , w_10397 );
not ( w_10397 , w_10398 );
and ( \3265_b0 , \3264_b0 , w_10399 );
and ( w_10398 ,  , w_10399 );
buf ( w_10397 , \901_b1 );
not ( w_10397 , w_10400 );
not (  , w_10401 );
and ( w_10400 , w_10401 , \901_b0 );
or ( \3266_b1 , \880_b1 , w_10403 );
not ( w_10403 , w_10404 );
and ( \3266_b0 , \880_b0 , w_10405 );
and ( w_10404 ,  , w_10405 );
buf ( w_10403 , \899_b1 );
not ( w_10403 , w_10406 );
not (  , w_10407 );
and ( w_10406 , w_10407 , \899_b0 );
or ( \3267_b1 , \3265_b1 , \3266_b1 );
xor ( \3267_b0 , \3265_b0 , w_10408 );
not ( w_10408 , w_10409 );
and ( w_10409 , \3266_b1 , \3266_b0 );
or ( \3268_b1 , \3263_b1 , w_10411 );
not ( w_10411 , w_10412 );
and ( \3268_b0 , \3263_b0 , w_10413 );
and ( w_10412 ,  , w_10413 );
buf ( w_10411 , \3267_b1 );
not ( w_10411 , w_10414 );
not (  , w_10415 );
and ( w_10414 , w_10415 , \3267_b0 );
or ( \3269_b1 , \3262_b1 , w_10417 );
not ( w_10417 , w_10418 );
and ( \3269_b0 , \3262_b0 , w_10419 );
and ( w_10418 ,  , w_10419 );
buf ( w_10417 , \3268_b1 );
not ( w_10417 , w_10420 );
not (  , w_10421 );
and ( w_10420 , w_10421 , \3268_b0 );
or ( \3271_b1 , \3212_b1 , w_10423 );
not ( w_10423 , w_10424 );
and ( \3271_b0 , \3212_b0 , w_10425 );
and ( w_10424 ,  , w_10425 );
buf ( w_10423 , \3270_b1 );
not ( w_10423 , w_10426 );
not (  , w_10427 );
and ( w_10426 , w_10427 , \3270_b0 );
or ( \3272_b1 , \3211_b1 , w_10429 );
not ( w_10429 , w_10430 );
and ( \3272_b0 , \3211_b0 , w_10431 );
and ( w_10430 ,  , w_10431 );
buf ( w_10429 , \3271_b1 );
not ( w_10429 , w_10432 );
not (  , w_10433 );
and ( w_10432 , w_10433 , \3271_b0 );
buf ( \3273_b1 , \2929_b1 );
not ( \3273_b1 , w_10434 );
not ( \3273_b0 , w_10435 );
and ( w_10434 , w_10435 , \2929_b0 );
or ( \3274_b1 , \3273_b1 , w_10437 );
not ( w_10437 , w_10438 );
and ( \3274_b0 , \3273_b0 , w_10439 );
and ( w_10438 ,  , w_10439 );
buf ( w_10437 , \2921_b1 );
not ( w_10437 , w_10440 );
not (  , w_10441 );
and ( w_10440 , w_10441 , \2921_b0 );
buf ( \3275_b1 , \3274_b1 );
not ( \3275_b1 , w_10442 );
not ( \3275_b0 , w_10443 );
and ( w_10442 , w_10443 , \3274_b0 );
buf ( \3276_b1 , \2815_b1 );
not ( \3276_b1 , w_10444 );
not ( \3276_b0 , w_10445 );
and ( w_10444 , w_10445 , \2815_b0 );
buf ( \3277_b1 , \3276_b1 );
not ( \3277_b1 , w_10446 );
not ( \3277_b0 , w_10447 );
and ( w_10446 , w_10447 , \3276_b0 );
buf ( \3278_b1 , \2916_b1 );
not ( \3278_b1 , w_10448 );
not ( \3278_b0 , w_10449 );
and ( w_10448 , w_10449 , \2916_b0 );
or ( \3279_b1 , \3277_b1 , w_10450 );
or ( \3279_b0 , \3277_b0 , \3278_b0 );
not ( \3278_b0 , w_10451 );
and ( w_10451 , w_10450 , \3278_b1 );
buf ( \3280_b1 , \2728_b1 );
buf ( \3280_b0 , \2728_b0 );
or ( \3281_b1 , \2927_b1 , w_10453 );
not ( w_10453 , w_10454 );
and ( \3281_b0 , \2927_b0 , w_10455 );
and ( w_10454 ,  , w_10455 );
buf ( w_10453 , \3280_b1 );
not ( w_10453 , w_10456 );
not (  , w_10457 );
and ( w_10456 , w_10457 , \3280_b0 );
or ( \3282_b1 , \3279_b1 , w_10459 );
not ( w_10459 , w_10460 );
and ( \3282_b0 , \3279_b0 , w_10461 );
and ( w_10460 ,  , w_10461 );
buf ( w_10459 , \3281_b1 );
not ( w_10459 , w_10462 );
not (  , w_10463 );
and ( w_10462 , w_10463 , \3281_b0 );
buf ( \3283_b1 , \3282_b1 );
not ( \3283_b1 , w_10464 );
not ( \3283_b0 , w_10465 );
and ( w_10464 , w_10465 , \3282_b0 );
or ( \3284_b1 , \3275_b1 , w_10466 );
or ( \3284_b0 , \3275_b0 , \3283_b0 );
not ( \3283_b0 , w_10467 );
and ( w_10467 , w_10466 , \3283_b1 );
or ( \3285_b1 , \3282_b1 , w_10468 );
or ( \3285_b0 , \3282_b0 , \3274_b0 );
not ( \3274_b0 , w_10469 );
and ( w_10469 , w_10468 , \3274_b1 );
or ( \3286_b1 , \3284_b1 , w_10471 );
not ( w_10471 , w_10472 );
and ( \3286_b0 , \3284_b0 , w_10473 );
and ( w_10472 ,  , w_10473 );
buf ( w_10471 , \3285_b1 );
not ( w_10471 , w_10474 );
not (  , w_10475 );
and ( w_10474 , w_10475 , \3285_b0 );
or ( \3287_b1 , \3286_b1 , w_10477 );
not ( w_10477 , w_10478 );
and ( \3287_b0 , \3286_b0 , w_10479 );
and ( w_10478 ,  , w_10479 );
buf ( w_10477 , \2936_b1 );
not ( w_10477 , w_10480 );
not (  , w_10481 );
and ( w_10480 , w_10481 , \2936_b0 );
or ( \3288_b1 , \a[14]_b1 , w_10483 );
not ( w_10483 , w_10484 );
and ( \3288_b0 , \a[14]_b0 , w_10485 );
and ( w_10484 ,  , w_10485 );
buf ( w_10483 , \1338_b1 );
not ( w_10483 , w_10486 );
not (  , w_10487 );
and ( w_10486 , w_10487 , \1338_b0 );
or ( \3289_b1 , \a[14]_b1 , w_10488 );
or ( \3289_b0 , \a[14]_b0 , \d[14]_b0 );
not ( \d[14]_b0 , w_10489 );
and ( w_10489 , w_10488 , \d[14]_b1 );
buf ( \3290_b1 , \3289_b1 );
not ( \3290_b1 , w_10490 );
not ( \3290_b0 , w_10491 );
and ( w_10490 , w_10491 , \3289_b0 );
buf ( \3291_b1 , \1457_b1 );
not ( \3291_b1 , w_10492 );
not ( \3291_b0 , w_10493 );
and ( w_10492 , w_10493 , \1457_b0 );
or ( \3292_b1 , \3290_b1 , w_10494 );
or ( \3292_b0 , \3290_b0 , \3291_b0 );
not ( \3291_b0 , w_10495 );
and ( w_10495 , w_10494 , \3291_b1 );
or ( \3294_b1 , \3292_b1 , w_10497 );
not ( w_10497 , w_10498 );
and ( \3294_b0 , \3292_b0 , w_10499 );
and ( w_10498 ,  , w_10499 );
buf ( w_10497 , \3293_b1 );
not ( w_10497 , w_10500 );
not (  , w_10501 );
and ( w_10500 , w_10501 , \3293_b0 );
buf ( \3295_b1 , \b[14]_b1 );
not ( \3295_b1 , w_10502 );
not ( \3295_b0 , w_10503 );
and ( w_10502 , w_10503 , \b[14]_b0 );
buf ( \3296_b1 , \2951_b1 );
not ( \3296_b1 , w_10504 );
not ( \3296_b0 , w_10505 );
and ( w_10504 , w_10505 , \2951_b0 );
or ( \3297_b1 , \3295_b1 , w_10506 );
or ( \3297_b0 , \3295_b0 , \3296_b0 );
not ( \3296_b0 , w_10507 );
and ( w_10507 , w_10506 , \3296_b1 );
or ( \3298_b1 , \a[14]_b1 , \1351_b1 );
not ( \1351_b1 , w_10508 );
and ( \3298_b0 , \a[14]_b0 , w_10509 );
and ( w_10508 , w_10509 , \1351_b0 );
or ( \3299_b1 , \d[14]_b1 , \c[14]_b1 );
not ( \c[14]_b1 , w_10510 );
and ( \3299_b0 , \d[14]_b0 , w_10511 );
and ( w_10510 , w_10511 , \c[14]_b0 );
buf ( \3300_b1 , \d[14]_b1 );
not ( \3300_b1 , w_10512 );
not ( \3300_b0 , w_10513 );
and ( w_10512 , w_10513 , \d[14]_b0 );
buf ( \3301_b1 , \c[14]_b1 );
not ( \3301_b1 , w_10514 );
not ( \3301_b0 , w_10515 );
and ( w_10514 , w_10515 , \c[14]_b0 );
or ( \3302_b1 , \3300_b1 , \3301_b1 );
not ( \3301_b1 , w_10516 );
and ( \3302_b0 , \3300_b0 , w_10517 );
and ( w_10516 , w_10517 , \3301_b0 );
or ( \3303_b1 , \3299_b1 , w_10519 );
not ( w_10519 , w_10520 );
and ( \3303_b0 , \3299_b0 , w_10521 );
and ( w_10520 ,  , w_10521 );
buf ( w_10519 , \3302_b1 );
not ( w_10519 , w_10522 );
not (  , w_10523 );
and ( w_10522 , w_10523 , \3302_b0 );
buf ( \3304_b1 , \3303_b1 );
not ( \3304_b1 , w_10524 );
not ( \3304_b0 , w_10525 );
and ( w_10524 , w_10525 , \3303_b0 );
buf ( \3305_b1 , \1320_b1 );
buf ( \3305_b0 , \1320_b0 );
buf ( \3306_b1 , \3305_b1 );
not ( \3306_b1 , w_10526 );
not ( \3306_b0 , w_10527 );
and ( w_10526 , w_10527 , \3305_b0 );
or ( \3307_b1 , \3304_b1 , w_10528 );
or ( \3307_b0 , \3304_b0 , \3306_b0 );
not ( \3306_b0 , w_10529 );
and ( w_10529 , w_10528 , \3306_b1 );
buf ( \3308_b1 , \2983_b1 );
not ( \3308_b1 , w_10530 );
not ( \3308_b0 , w_10531 );
and ( w_10530 , w_10531 , \2983_b0 );
or ( \3309_b1 , \3308_b1 , w_10533 );
not ( w_10533 , w_10534 );
and ( \3309_b0 , \3308_b0 , w_10535 );
and ( w_10534 ,  , w_10535 );
buf ( w_10533 , \3015_b1 );
not ( w_10533 , w_10536 );
not (  , w_10537 );
and ( w_10536 , w_10537 , \3015_b0 );
buf ( \3310_b1 , \3309_b1 );
not ( \3310_b1 , w_10538 );
not ( \3310_b0 , w_10539 );
and ( w_10538 , w_10539 , \3309_b0 );
buf ( \3312_b1 , \3013_b1 );
not ( \3312_b1 , w_10540 );
not ( \3312_b0 , w_10541 );
and ( w_10540 , w_10541 , \3013_b0 );
or ( \3313_b1 , \3007_b1 , w_10543 );
not ( w_10543 , w_10544 );
and ( \3313_b0 , \3007_b0 , w_10545 );
and ( w_10544 ,  , w_10545 );
buf ( w_10543 , \2982_b1 );
not ( w_10543 , w_10546 );
not (  , w_10547 );
and ( w_10546 , w_10547 , \2982_b0 );
or ( \3314_b1 , \3312_b1 , w_10549 );
not ( w_10549 , w_10550 );
and ( \3314_b0 , \3312_b0 , w_10551 );
and ( w_10550 ,  , w_10551 );
buf ( w_10549 , \3313_b1 );
not ( w_10549 , w_10552 );
not (  , w_10553 );
and ( w_10552 , w_10553 , \3313_b0 );
or ( \3315_b1 , \3311_b1 , w_10555 );
not ( w_10555 , w_10556 );
and ( \3315_b0 , \3311_b0 , w_10557 );
and ( w_10556 ,  , w_10557 );
buf ( w_10555 , \3314_b1 );
not ( w_10555 , w_10558 );
not (  , w_10559 );
and ( w_10558 , w_10559 , \3314_b0 );
buf ( \3316_b1 , \3315_b1 );
not ( \3316_b1 , w_10560 );
not ( \3316_b0 , w_10561 );
and ( w_10560 , w_10561 , \3315_b0 );
or ( \3317_b1 , \3310_b1 , w_10562 );
or ( \3317_b0 , \3310_b0 , \3316_b0 );
not ( \3316_b0 , w_10563 );
and ( w_10563 , w_10562 , \3316_b1 );
or ( \3318_b1 , \3315_b1 , w_10564 );
or ( \3318_b0 , \3315_b0 , \3309_b0 );
not ( \3309_b0 , w_10565 );
and ( w_10565 , w_10564 , \3309_b1 );
or ( \3319_b1 , \3317_b1 , w_10567 );
not ( w_10567 , w_10568 );
and ( \3319_b0 , \3317_b0 , w_10569 );
and ( w_10568 ,  , w_10569 );
buf ( w_10567 , \3318_b1 );
not ( w_10567 , w_10570 );
not (  , w_10571 );
and ( w_10570 , w_10571 , \3318_b0 );
or ( \3320_b1 , \2961_b1 , \3319_b1 );
not ( \3319_b1 , w_10572 );
and ( \3320_b0 , \2961_b0 , w_10573 );
and ( w_10572 , w_10573 , \3319_b0 );
buf ( \3321_b1 , \3045_b1 );
not ( \3321_b1 , w_10574 );
not ( \3321_b0 , w_10575 );
and ( w_10574 , w_10575 , \3045_b0 );
or ( \3322_b1 , \3321_b1 , w_10577 );
not ( w_10577 , w_10578 );
and ( \3322_b0 , \3321_b0 , w_10579 );
and ( w_10578 ,  , w_10579 );
buf ( w_10577 , \3077_b1 );
not ( w_10577 , w_10580 );
not (  , w_10581 );
and ( w_10580 , w_10581 , \3077_b0 );
buf ( \3323_b1 , \3322_b1 );
not ( \3323_b1 , w_10582 );
not ( \3323_b0 , w_10583 );
and ( w_10582 , w_10583 , \3322_b0 );
buf ( \3325_b1 , \3075_b1 );
not ( \3325_b1 , w_10584 );
not ( \3325_b0 , w_10585 );
and ( w_10584 , w_10585 , \3075_b0 );
or ( \3326_b1 , \3069_b1 , w_10587 );
not ( w_10587 , w_10588 );
and ( \3326_b0 , \3069_b0 , w_10589 );
and ( w_10588 ,  , w_10589 );
buf ( w_10587 , \3044_b1 );
not ( w_10587 , w_10590 );
not (  , w_10591 );
and ( w_10590 , w_10591 , \3044_b0 );
or ( \3327_b1 , \3325_b1 , w_10593 );
not ( w_10593 , w_10594 );
and ( \3327_b0 , \3325_b0 , w_10595 );
and ( w_10594 ,  , w_10595 );
buf ( w_10593 , \3326_b1 );
not ( w_10593 , w_10596 );
not (  , w_10597 );
and ( w_10596 , w_10597 , \3326_b0 );
or ( \3328_b1 , \3324_b1 , w_10599 );
not ( w_10599 , w_10600 );
and ( \3328_b0 , \3324_b0 , w_10601 );
and ( w_10600 ,  , w_10601 );
buf ( w_10599 , \3327_b1 );
not ( w_10599 , w_10602 );
not (  , w_10603 );
and ( w_10602 , w_10603 , \3327_b0 );
buf ( \3329_b1 , \3328_b1 );
not ( \3329_b1 , w_10604 );
not ( \3329_b0 , w_10605 );
and ( w_10604 , w_10605 , \3328_b0 );
or ( \3330_b1 , \3323_b1 , w_10606 );
or ( \3330_b0 , \3323_b0 , \3329_b0 );
not ( \3329_b0 , w_10607 );
and ( w_10607 , w_10606 , \3329_b1 );
or ( \3331_b1 , \3328_b1 , w_10608 );
or ( \3331_b0 , \3328_b0 , \3322_b0 );
not ( \3322_b0 , w_10609 );
and ( w_10609 , w_10608 , \3322_b1 );
or ( \3332_b1 , \3330_b1 , w_10611 );
not ( w_10611 , w_10612 );
and ( \3332_b0 , \3330_b0 , w_10613 );
and ( w_10612 ,  , w_10613 );
buf ( w_10611 , \3331_b1 );
not ( w_10611 , w_10614 );
not (  , w_10615 );
and ( w_10614 , w_10615 , \3331_b0 );
buf ( \3333_b1 , \3332_b1 );
not ( \3333_b1 , w_10616 );
not ( \3333_b0 , w_10617 );
and ( w_10616 , w_10617 , \3332_b0 );
buf ( \3334_b1 , \3087_b1 );
not ( \3334_b1 , w_10618 );
not ( \3334_b0 , w_10619 );
and ( w_10618 , w_10619 , \3087_b0 );
or ( \3335_b1 , \3333_b1 , w_10620 );
or ( \3335_b0 , \3333_b0 , \3334_b0 );
not ( \3334_b0 , w_10621 );
and ( w_10621 , w_10620 , \3334_b1 );
buf ( \3336_b1 , \1323_b1 );
not ( \3336_b1 , w_10622 );
not ( \3336_b0 , w_10623 );
and ( w_10622 , w_10623 , \1323_b0 );
buf ( \3337_b1 , \3301_b1 );
not ( \3337_b1 , w_10624 );
not ( \3337_b0 , w_10625 );
and ( w_10624 , w_10625 , \3301_b0 );
or ( \3338_b1 , \3336_b1 , \3337_b1 );
not ( \3337_b1 , w_10626 );
and ( \3338_b0 , \3336_b0 , w_10627 );
and ( w_10626 , w_10627 , \3337_b0 );
or ( \3339_b1 , \1282_b1 , \d[14]_b1 );
not ( \d[14]_b1 , w_10628 );
and ( \3339_b0 , \1282_b0 , w_10629 );
and ( w_10628 , w_10629 , \d[14]_b0 );
or ( \3340_b1 , \3338_b1 , w_10631 );
not ( w_10631 , w_10632 );
and ( \3340_b0 , \3338_b0 , w_10633 );
and ( w_10632 ,  , w_10633 );
buf ( w_10631 , \3339_b1 );
not ( w_10631 , w_10634 );
not (  , w_10635 );
and ( w_10634 , w_10635 , \3339_b0 );
or ( \3341_b1 , \3335_b1 , w_10637 );
not ( w_10637 , w_10638 );
and ( \3341_b0 , \3335_b0 , w_10639 );
and ( w_10638 ,  , w_10639 );
buf ( w_10637 , \3340_b1 );
not ( w_10637 , w_10640 );
not (  , w_10641 );
and ( w_10640 , w_10641 , \3340_b0 );
or ( \3342_b1 , \3320_b1 , w_10643 );
not ( w_10643 , w_10644 );
and ( \3342_b0 , \3320_b0 , w_10645 );
and ( w_10644 ,  , w_10645 );
buf ( w_10643 , \3341_b1 );
not ( w_10643 , w_10646 );
not (  , w_10647 );
and ( w_10646 , w_10647 , \3341_b0 );
or ( \3343_b1 , \3307_b1 , w_10649 );
not ( w_10649 , w_10650 );
and ( \3343_b0 , \3307_b0 , w_10651 );
and ( w_10650 ,  , w_10651 );
buf ( w_10649 , \3342_b1 );
not ( w_10649 , w_10652 );
not (  , w_10653 );
and ( w_10652 , w_10653 , \3342_b0 );
or ( \3344_b1 , \3298_b1 , w_10655 );
not ( w_10655 , w_10656 );
and ( \3344_b0 , \3298_b0 , w_10657 );
and ( w_10656 ,  , w_10657 );
buf ( w_10655 , \3343_b1 );
not ( w_10655 , w_10658 );
not (  , w_10659 );
and ( w_10658 , w_10659 , \3343_b0 );
or ( \3345_b1 , \3297_b1 , w_10661 );
not ( w_10661 , w_10662 );
and ( \3345_b0 , \3297_b0 , w_10663 );
and ( w_10662 ,  , w_10663 );
buf ( w_10661 , \3344_b1 );
not ( w_10661 , w_10664 );
not (  , w_10665 );
and ( w_10664 , w_10665 , \3344_b0 );
or ( \3346_b1 , \3294_b1 , w_10667 );
not ( w_10667 , w_10668 );
and ( \3346_b0 , \3294_b0 , w_10669 );
and ( w_10668 ,  , w_10669 );
buf ( w_10667 , \3345_b1 );
not ( w_10667 , w_10670 );
not (  , w_10671 );
and ( w_10670 , w_10671 , \3345_b0 );
buf ( \3347_b1 , \1953_b1 );
not ( \3347_b1 , w_10672 );
not ( \3347_b0 , w_10673 );
and ( w_10672 , w_10673 , \1953_b0 );
buf ( \3348_b1 , \3347_b1 );
not ( \3348_b1 , w_10674 );
not ( \3348_b0 , w_10675 );
and ( w_10674 , w_10675 , \3347_b0 );
buf ( \3349_b1 , \1908_b1 );
not ( \3349_b1 , w_10676 );
not ( \3349_b0 , w_10677 );
and ( w_10676 , w_10677 , \1908_b0 );
buf ( \3350_b1 , \3349_b1 );
not ( \3350_b1 , w_10678 );
not ( \3350_b0 , w_10679 );
and ( w_10678 , w_10679 , \3349_b0 );
or ( \3351_b1 , \3348_b1 , w_10680 );
or ( \3351_b0 , \3348_b0 , \3350_b0 );
not ( \3350_b0 , w_10681 );
and ( w_10681 , w_10680 , \3350_b1 );
or ( \3352_b1 , \3349_b1 , w_10682 );
or ( \3352_b0 , \3349_b0 , \3347_b0 );
not ( \3347_b0 , w_10683 );
and ( w_10683 , w_10682 , \3347_b1 );
or ( \3353_b1 , \3351_b1 , w_10685 );
not ( w_10685 , w_10686 );
and ( \3353_b0 , \3351_b0 , w_10687 );
and ( w_10686 ,  , w_10687 );
buf ( w_10685 , \3352_b1 );
not ( w_10685 , w_10688 );
not (  , w_10689 );
and ( w_10688 , w_10689 , \3352_b0 );
buf ( \3354_b1 , \3353_b1 );
not ( \3354_b1 , w_10690 );
not ( \3354_b0 , w_10691 );
and ( w_10690 , w_10691 , \3353_b0 );
buf ( \3355_b1 , \2113_b1 );
not ( \3355_b1 , w_10692 );
not ( \3355_b0 , w_10693 );
and ( w_10692 , w_10693 , \2113_b0 );
buf ( \3356_b1 , \3355_b1 );
not ( \3356_b1 , w_10694 );
not ( \3356_b0 , w_10695 );
and ( w_10694 , w_10695 , \3355_b0 );
buf ( \3357_b1 , \2213_b1 );
not ( \3357_b1 , w_10696 );
not ( \3357_b0 , w_10697 );
and ( w_10696 , w_10697 , \2213_b0 );
or ( \3358_b1 , \3356_b1 , w_10698 );
or ( \3358_b0 , \3356_b0 , \3357_b0 );
not ( \3357_b0 , w_10699 );
and ( w_10699 , w_10698 , \3357_b1 );
or ( \3359_b1 , \2223_b1 , w_10701 );
not ( w_10701 , w_10702 );
and ( \3359_b0 , \2223_b0 , w_10703 );
and ( w_10702 ,  , w_10703 );
buf ( w_10701 , \2031_b1 );
not ( w_10701 , w_10704 );
not (  , w_10705 );
and ( w_10704 , w_10705 , \2031_b0 );
or ( \3360_b1 , \3358_b1 , w_10707 );
not ( w_10707 , w_10708 );
and ( \3360_b0 , \3358_b0 , w_10709 );
and ( w_10708 ,  , w_10709 );
buf ( w_10707 , \3359_b1 );
not ( w_10707 , w_10710 );
not (  , w_10711 );
and ( w_10710 , w_10711 , \3359_b0 );
buf ( \3361_b1 , \3360_b1 );
not ( \3361_b1 , w_10712 );
not ( \3361_b0 , w_10713 );
and ( w_10712 , w_10713 , \3360_b0 );
or ( \3362_b1 , \3354_b1 , w_10714 );
or ( \3362_b0 , \3354_b0 , \3361_b0 );
not ( \3361_b0 , w_10715 );
and ( w_10715 , w_10714 , \3361_b1 );
or ( \3363_b1 , \3353_b1 , w_10716 );
or ( \3363_b0 , \3353_b0 , \3360_b0 );
not ( \3360_b0 , w_10717 );
and ( w_10717 , w_10716 , \3360_b1 );
or ( \3364_b1 , \3362_b1 , w_10719 );
not ( w_10719 , w_10720 );
and ( \3364_b0 , \3362_b0 , w_10721 );
and ( w_10720 ,  , w_10721 );
buf ( w_10719 , \3363_b1 );
not ( w_10719 , w_10722 );
not (  , w_10723 );
and ( w_10722 , w_10723 , \3363_b0 );
or ( \3365_b1 , \3364_b1 , w_10725 );
not ( w_10725 , w_10726 );
and ( \3365_b0 , \3364_b0 , w_10727 );
and ( w_10726 ,  , w_10727 );
buf ( w_10725 , \1529_b1 );
not ( w_10725 , w_10728 );
not (  , w_10729 );
and ( w_10728 , w_10729 , \1529_b0 );
buf ( \3367_b1 , \a[2]_b1 );
not ( \3367_b1 , w_10730 );
not ( \3367_b0 , w_10731 );
and ( w_10730 , w_10731 , \a[2]_b0 );
buf ( \3368_b1 , \3114_b1 );
not ( \3368_b1 , w_10732 );
not ( \3368_b0 , w_10733 );
and ( w_10732 , w_10733 , \3114_b0 );
or ( \3369_b1 , \3367_b1 , w_10734 );
or ( \3369_b0 , \3367_b0 , \3368_b0 );
not ( \3368_b0 , w_10735 );
and ( w_10735 , w_10734 , \3368_b1 );
buf ( \3370_b1 , \d[2]_b1 );
not ( \3370_b1 , w_10736 );
not ( \3370_b0 , w_10737 );
and ( w_10736 , w_10737 , \d[2]_b0 );
buf ( \3371_b1 , \1457_b1 );
not ( \3371_b1 , w_10738 );
not ( \3371_b0 , w_10739 );
and ( w_10738 , w_10739 , \1457_b0 );
or ( \3372_b1 , \3370_b1 , w_10740 );
or ( \3372_b0 , \3370_b0 , \3371_b0 );
not ( \3371_b0 , w_10741 );
and ( w_10741 , w_10740 , \3371_b1 );
buf ( \3373_b1 , \2942_b1 );
not ( \3373_b1 , w_10742 );
not ( \3373_b0 , w_10743 );
and ( w_10742 , w_10743 , \2942_b0 );
or ( \3374_b1 , \b[2]_b1 , \c[2]_b1 );
not ( \c[2]_b1 , w_10744 );
and ( \3374_b0 , \b[2]_b0 , w_10745 );
and ( w_10744 , w_10745 , \c[2]_b0 );
or ( \3375_b1 , \3373_b1 , \3374_b1 );
not ( \3374_b1 , w_10746 );
and ( \3375_b0 , \3373_b0 , w_10747 );
and ( w_10746 , w_10747 , \3374_b0 );
or ( \3376_b1 , \a[2]_b1 , w_10748 );
or ( \3376_b0 , \a[2]_b0 , \b[2]_b0 );
not ( \b[2]_b0 , w_10749 );
and ( w_10749 , w_10748 , \b[2]_b1 );
buf ( \3377_b1 , \3376_b1 );
not ( \3377_b1 , w_10750 );
not ( \3377_b0 , w_10751 );
and ( w_10750 , w_10751 , \3376_b0 );
buf ( \3378_b1 , \1351_b1 );
not ( \3378_b1 , w_10752 );
not ( \3378_b0 , w_10753 );
and ( w_10752 , w_10753 , \1351_b0 );
or ( \3379_b1 , \3377_b1 , w_10754 );
or ( \3379_b0 , \3377_b0 , \3378_b0 );
not ( \3378_b0 , w_10755 );
and ( w_10755 , w_10754 , \3378_b1 );
or ( \3380_b1 , \c[2]_b1 , \d[2]_b1 );
xor ( \3380_b0 , \c[2]_b0 , w_10756 );
not ( w_10756 , w_10757 );
and ( w_10757 , \d[2]_b1 , \d[2]_b0 );
buf ( \3381_b1 , \3380_b1 );
not ( \3381_b1 , w_10758 );
not ( \3381_b0 , w_10759 );
and ( w_10758 , w_10759 , \3380_b0 );
buf ( \3382_b1 , \1383_b1 );
not ( \3382_b1 , w_10760 );
not ( \3382_b0 , w_10761 );
and ( w_10760 , w_10761 , \1383_b0 );
or ( \3383_b1 , \3381_b1 , w_10762 );
or ( \3383_b0 , \3381_b0 , \3382_b0 );
not ( \3382_b0 , w_10763 );
and ( w_10763 , w_10762 , \3382_b1 );
buf ( \3384_b1 , \1046_b1 );
not ( \3384_b1 , w_10764 );
not ( \3384_b0 , w_10765 );
and ( w_10764 , w_10765 , \1046_b0 );
buf ( \3385_b1 , \1049_b1 );
not ( \3385_b1 , w_10766 );
not ( \3385_b0 , w_10767 );
and ( w_10766 , w_10767 , \1049_b0 );
or ( \3386_b1 , \3385_b1 , w_10769 );
not ( w_10769 , w_10770 );
and ( \3386_b0 , \3385_b0 , w_10771 );
and ( w_10770 ,  , w_10771 );
buf ( w_10769 , \1037_b1 );
not ( w_10769 , w_10772 );
not (  , w_10773 );
and ( w_10772 , w_10773 , \1037_b0 );
buf ( \3387_b1 , \3386_b1 );
not ( \3387_b1 , w_10774 );
not ( \3387_b0 , w_10775 );
and ( w_10774 , w_10775 , \3386_b0 );
or ( \3388_b1 , \3384_b1 , w_10776 );
or ( \3388_b0 , \3384_b0 , \3387_b0 );
not ( \3387_b0 , w_10777 );
and ( w_10777 , w_10776 , \3387_b1 );
or ( \3389_b1 , \3386_b1 , w_10778 );
or ( \3389_b0 , \3386_b0 , \1046_b0 );
not ( \1046_b0 , w_10779 );
and ( w_10779 , w_10778 , \1046_b1 );
or ( \3390_b1 , \3388_b1 , w_10781 );
not ( w_10781 , w_10782 );
and ( \3390_b0 , \3388_b0 , w_10783 );
and ( w_10782 ,  , w_10783 );
buf ( w_10781 , \3389_b1 );
not ( w_10781 , w_10784 );
not (  , w_10785 );
and ( w_10784 , w_10785 , \3389_b0 );
or ( \3391_b1 , \1478_b1 , \3390_b1 );
not ( \3390_b1 , w_10786 );
and ( \3391_b0 , \1478_b0 , w_10787 );
and ( w_10786 , w_10787 , \3390_b0 );
or ( \3392_b1 , \1486_b1 , w_10789 );
not ( w_10789 , w_10790 );
and ( \3392_b0 , \1486_b0 , w_10791 );
and ( w_10790 ,  , w_10791 );
buf ( w_10789 , \1186_b1 );
not ( w_10789 , w_10792 );
not (  , w_10793 );
and ( w_10792 , w_10793 , \1186_b0 );
buf ( \3393_b1 , \3392_b1 );
not ( \3393_b1 , w_10794 );
not ( \3393_b0 , w_10795 );
and ( w_10794 , w_10795 , \3392_b0 );
buf ( \3394_b1 , \1181_b1 );
not ( \3394_b1 , w_10796 );
not ( \3394_b0 , w_10797 );
and ( w_10796 , w_10797 , \1181_b0 );
or ( \3395_b1 , \3393_b1 , w_10798 );
or ( \3395_b0 , \3393_b0 , \3394_b0 );
not ( \3394_b0 , w_10799 );
and ( w_10799 , w_10798 , \3394_b1 );
or ( \3396_b1 , \1181_b1 , w_10800 );
or ( \3396_b0 , \1181_b0 , \3392_b0 );
not ( \3392_b0 , w_10801 );
and ( w_10801 , w_10800 , \3392_b1 );
or ( \3397_b1 , \3395_b1 , w_10803 );
not ( w_10803 , w_10804 );
and ( \3397_b0 , \3395_b0 , w_10805 );
and ( w_10804 ,  , w_10805 );
buf ( w_10803 , \3396_b1 );
not ( w_10803 , w_10806 );
not (  , w_10807 );
and ( w_10806 , w_10807 , \3396_b0 );
buf ( \3398_b1 , \3397_b1 );
not ( \3398_b1 , w_10808 );
not ( \3398_b0 , w_10809 );
and ( w_10808 , w_10809 , \3397_b0 );
buf ( \3399_b1 , \1220_b1 );
not ( \3399_b1 , w_10810 );
not ( \3399_b0 , w_10811 );
and ( w_10810 , w_10811 , \1220_b0 );
or ( \3400_b1 , \3398_b1 , w_10812 );
or ( \3400_b0 , \3398_b0 , \3399_b0 );
not ( \3399_b0 , w_10813 );
and ( w_10813 , w_10812 , \3399_b1 );
or ( \3401_b1 , \1500_b1 , w_10815 );
not ( w_10815 , w_10816 );
and ( \3401_b0 , \1500_b0 , w_10817 );
and ( w_10816 ,  , w_10817 );
buf ( w_10815 , \1249_b1 );
not ( w_10815 , w_10818 );
not (  , w_10819 );
and ( w_10818 , w_10819 , \1249_b0 );
buf ( \3402_b1 , \3401_b1 );
not ( \3402_b1 , w_10820 );
not ( \3402_b0 , w_10821 );
and ( w_10820 , w_10821 , \3401_b0 );
buf ( \3403_b1 , \1244_b1 );
not ( \3403_b1 , w_10822 );
not ( \3403_b0 , w_10823 );
and ( w_10822 , w_10823 , \1244_b0 );
or ( \3404_b1 , \3402_b1 , w_10824 );
or ( \3404_b0 , \3402_b0 , \3403_b0 );
not ( \3403_b0 , w_10825 );
and ( w_10825 , w_10824 , \3403_b1 );
or ( \3405_b1 , \1244_b1 , w_10826 );
or ( \3405_b0 , \1244_b0 , \3401_b0 );
not ( \3401_b0 , w_10827 );
and ( w_10827 , w_10826 , \3401_b1 );
or ( \3406_b1 , \3404_b1 , w_10829 );
not ( w_10829 , w_10830 );
and ( \3406_b0 , \3404_b0 , w_10831 );
and ( w_10830 ,  , w_10831 );
buf ( w_10829 , \3405_b1 );
not ( w_10829 , w_10832 );
not (  , w_10833 );
and ( w_10832 , w_10833 , \3405_b0 );
buf ( \3407_b1 , \3406_b1 );
not ( \3407_b1 , w_10834 );
not ( \3407_b0 , w_10835 );
and ( w_10834 , w_10835 , \3406_b0 );
buf ( \3408_b1 , \1232_b1 );
not ( \3408_b1 , w_10836 );
not ( \3408_b0 , w_10837 );
and ( w_10836 , w_10837 , \1232_b0 );
or ( \3409_b1 , \3407_b1 , w_10838 );
or ( \3409_b0 , \3407_b0 , \3408_b0 );
not ( \3408_b0 , w_10839 );
and ( w_10839 , w_10838 , \3408_b1 );
or ( \3410_b1 , \1282_b1 , \d[2]_b1 );
not ( \d[2]_b1 , w_10840 );
and ( \3410_b0 , \1282_b0 , w_10841 );
and ( w_10840 , w_10841 , \d[2]_b0 );
buf ( \3411_b1 , \c[2]_b1 );
not ( \3411_b1 , w_10842 );
not ( \3411_b0 , w_10843 );
and ( w_10842 , w_10843 , \c[2]_b0 );
buf ( \3412_b1 , \1287_b1 );
not ( \3412_b1 , w_10844 );
not ( \3412_b0 , w_10845 );
and ( w_10844 , w_10845 , \1287_b0 );
or ( \3413_b1 , \3411_b1 , w_10846 );
or ( \3413_b0 , \3411_b0 , \3412_b0 );
not ( \3412_b0 , w_10847 );
and ( w_10847 , w_10846 , \3412_b1 );
or ( \3414_b1 , \1293_b1 , w_10849 );
not ( w_10849 , w_10850 );
and ( \3414_b0 , \1293_b0 , w_10851 );
and ( w_10850 ,  , w_10851 );
buf ( w_10849 , \b[2]_b1 );
not ( w_10849 , w_10852 );
not (  , w_10853 );
and ( w_10852 , w_10853 , \b[2]_b0 );
or ( \3415_b1 , \3413_b1 , w_10855 );
not ( w_10855 , w_10856 );
and ( \3415_b0 , \3413_b0 , w_10857 );
and ( w_10856 ,  , w_10857 );
buf ( w_10855 , \3414_b1 );
not ( w_10855 , w_10858 );
not (  , w_10859 );
and ( w_10858 , w_10859 , \3414_b0 );
or ( \3416_b1 , \3410_b1 , w_10861 );
not ( w_10861 , w_10862 );
and ( \3416_b0 , \3410_b0 , w_10863 );
and ( w_10862 ,  , w_10863 );
buf ( w_10861 , \3415_b1 );
not ( w_10861 , w_10864 );
not (  , w_10865 );
and ( w_10864 , w_10865 , \3415_b0 );
or ( \3417_b1 , \3409_b1 , w_10867 );
not ( w_10867 , w_10868 );
and ( \3417_b0 , \3409_b0 , w_10869 );
and ( w_10868 ,  , w_10869 );
buf ( w_10867 , \3416_b1 );
not ( w_10867 , w_10870 );
not (  , w_10871 );
and ( w_10870 , w_10871 , \3416_b0 );
buf ( \3418_b1 , \3417_b1 );
not ( \3418_b1 , w_10872 );
not ( \3418_b0 , w_10873 );
and ( w_10872 , w_10873 , \3417_b0 );
or ( \3419_b1 , \3400_b1 , w_10875 );
not ( w_10875 , w_10876 );
and ( \3419_b0 , \3400_b0 , w_10877 );
and ( w_10876 ,  , w_10877 );
buf ( w_10875 , \3418_b1 );
not ( w_10875 , w_10878 );
not (  , w_10879 );
and ( w_10878 , w_10879 , \3418_b0 );
or ( \3420_b1 , \3391_b1 , w_10881 );
not ( w_10881 , w_10882 );
and ( \3420_b0 , \3391_b0 , w_10883 );
and ( w_10882 ,  , w_10883 );
buf ( w_10881 , \3419_b1 );
not ( w_10881 , w_10884 );
not (  , w_10885 );
and ( w_10884 , w_10885 , \3419_b0 );
or ( \3421_b1 , \3383_b1 , w_10887 );
not ( w_10887 , w_10888 );
and ( \3421_b0 , \3383_b0 , w_10889 );
and ( w_10888 ,  , w_10889 );
buf ( w_10887 , \3420_b1 );
not ( w_10887 , w_10890 );
not (  , w_10891 );
and ( w_10890 , w_10891 , \3420_b0 );
buf ( \3422_b1 , \916_b1 );
not ( \3422_b1 , w_10892 );
not ( \3422_b0 , w_10893 );
and ( w_10892 , w_10893 , \916_b0 );
buf ( \3423_b1 , \863_b1 );
not ( \3423_b1 , w_10894 );
not ( \3423_b0 , w_10895 );
and ( w_10894 , w_10895 , \863_b0 );
or ( \3424_b1 , \3423_b1 , w_10897 );
not ( w_10897 , w_10898 );
and ( \3424_b0 , \3423_b0 , w_10899 );
and ( w_10898 ,  , w_10899 );
buf ( w_10897 , \851_b1 );
not ( w_10897 , w_10900 );
not (  , w_10901 );
and ( w_10900 , w_10901 , \851_b0 );
or ( \3425_b1 , \861_b1 , \3424_b1 );
xor ( \3425_b0 , \861_b0 , w_10902 );
not ( w_10902 , w_10903 );
and ( w_10903 , \3424_b1 , \3424_b0 );
or ( \3426_b1 , \3422_b1 , w_10905 );
not ( w_10905 , w_10906 );
and ( \3426_b0 , \3422_b0 , w_10907 );
and ( w_10906 ,  , w_10907 );
buf ( w_10905 , \3425_b1 );
not ( w_10905 , w_10908 );
not (  , w_10909 );
and ( w_10908 , w_10909 , \3425_b0 );
or ( \3427_b1 , \3421_b1 , w_10911 );
not ( w_10911 , w_10912 );
and ( \3427_b0 , \3421_b0 , w_10913 );
and ( w_10912 ,  , w_10913 );
buf ( w_10911 , \3426_b1 );
not ( w_10911 , w_10914 );
not (  , w_10915 );
and ( w_10914 , w_10915 , \3426_b0 );
or ( \3428_b1 , \3379_b1 , w_10917 );
not ( w_10917 , w_10918 );
and ( \3428_b0 , \3379_b0 , w_10919 );
and ( w_10918 ,  , w_10919 );
buf ( w_10917 , \3427_b1 );
not ( w_10917 , w_10920 );
not (  , w_10921 );
and ( w_10920 , w_10921 , \3427_b0 );
or ( \3429_b1 , \3375_b1 , w_10923 );
not ( w_10923 , w_10924 );
and ( \3429_b0 , \3375_b0 , w_10925 );
and ( w_10924 ,  , w_10925 );
buf ( w_10923 , \3428_b1 );
not ( w_10923 , w_10926 );
not (  , w_10927 );
and ( w_10926 , w_10927 , \3428_b0 );
or ( \3430_b1 , \3372_b1 , w_10929 );
not ( w_10929 , w_10930 );
and ( \3430_b0 , \3372_b0 , w_10931 );
and ( w_10930 ,  , w_10931 );
buf ( w_10929 , \3429_b1 );
not ( w_10929 , w_10932 );
not (  , w_10933 );
and ( w_10932 , w_10933 , \3429_b0 );
buf ( \3431_b1 , \3430_b1 );
not ( \3431_b1 , w_10934 );
not ( \3431_b0 , w_10935 );
and ( w_10934 , w_10935 , \3430_b0 );
or ( \3432_b1 , \3369_b1 , w_10937 );
not ( w_10937 , w_10938 );
and ( \3432_b0 , \3369_b0 , w_10939 );
and ( w_10938 ,  , w_10939 );
buf ( w_10937 , \3431_b1 );
not ( w_10937 , w_10940 );
not (  , w_10941 );
and ( w_10940 , w_10941 , \3431_b0 );
buf ( \3433_b1 , \a[10]_b1 );
not ( \3433_b1 , w_10942 );
not ( \3433_b0 , w_10943 );
and ( w_10942 , w_10943 , \a[10]_b0 );
buf ( \3434_b1 , \2946_b1 );
not ( \3434_b1 , w_10944 );
not ( \3434_b0 , w_10945 );
and ( w_10944 , w_10945 , \2946_b0 );
or ( \3435_b1 , \3433_b1 , w_10946 );
or ( \3435_b0 , \3433_b0 , \3434_b0 );
not ( \3434_b0 , w_10947 );
and ( w_10947 , w_10946 , \3434_b1 );
buf ( \3436_b1 , \a[10]_b1 );
not ( \3436_b1 , w_10948 );
not ( \3436_b0 , w_10949 );
and ( w_10948 , w_10949 , \a[10]_b0 );
buf ( \3437_b1 , \1466_b1 );
not ( \3437_b1 , w_10950 );
not ( \3437_b0 , w_10951 );
and ( w_10950 , w_10951 , \1466_b0 );
or ( \3438_b1 , \3436_b1 , w_10952 );
or ( \3438_b0 , \3436_b0 , \3437_b0 );
not ( \3437_b0 , w_10953 );
and ( w_10953 , w_10952 , \3437_b1 );
or ( \3439_b1 , \c[10]_b1 , \d[10]_b1 );
xor ( \3439_b0 , \c[10]_b0 , w_10954 );
not ( w_10954 , w_10955 );
and ( w_10955 , \d[10]_b1 , \d[10]_b0 );
or ( \3440_b1 , \3305_b1 , \3439_b1 );
not ( \3439_b1 , w_10956 );
and ( \3440_b0 , \3305_b0 , w_10957 );
and ( w_10956 , w_10957 , \3439_b0 );
or ( \3441_b1 , \3134_b1 , \3002_b1 );
not ( \3002_b1 , w_10958 );
and ( \3441_b0 , \3134_b0 , w_10959 );
and ( w_10958 , w_10959 , \3002_b0 );
buf ( \3442_b1 , \3441_b1 );
not ( \3442_b1 , w_10960 );
not ( \3442_b0 , w_10961 );
and ( w_10960 , w_10961 , \3441_b0 );
or ( \3443_b1 , \2979_b1 , \2991_b1 );
not ( \2991_b1 , w_10962 );
and ( \3443_b0 , \2979_b0 , w_10963 );
and ( w_10962 , w_10963 , \2991_b0 );
or ( \3444_b1 , \3443_b1 , w_10965 );
not ( w_10965 , w_10966 );
and ( \3444_b0 , \3443_b0 , w_10967 );
and ( w_10966 ,  , w_10967 );
buf ( w_10965 , \2997_b1 );
not ( w_10965 , w_10968 );
not (  , w_10969 );
and ( w_10968 , w_10969 , \2997_b0 );
buf ( \3445_b1 , \3444_b1 );
not ( \3445_b1 , w_10970 );
not ( \3445_b0 , w_10971 );
and ( w_10970 , w_10971 , \3444_b0 );
or ( \3446_b1 , \3442_b1 , w_10972 );
or ( \3446_b0 , \3442_b0 , \3445_b0 );
not ( \3445_b0 , w_10973 );
and ( w_10973 , w_10972 , \3445_b1 );
or ( \3447_b1 , \3444_b1 , w_10974 );
or ( \3447_b0 , \3444_b0 , \3441_b0 );
not ( \3441_b0 , w_10975 );
and ( w_10975 , w_10974 , \3441_b1 );
or ( \3448_b1 , \3446_b1 , w_10977 );
not ( w_10977 , w_10978 );
and ( \3448_b0 , \3446_b0 , w_10979 );
and ( w_10978 ,  , w_10979 );
buf ( w_10977 , \3447_b1 );
not ( w_10977 , w_10980 );
not (  , w_10981 );
and ( w_10980 , w_10981 , \3447_b0 );
buf ( \3449_b1 , \3448_b1 );
not ( \3449_b1 , w_10982 );
not ( \3449_b0 , w_10983 );
and ( w_10982 , w_10983 , \3448_b0 );
buf ( \3450_b1 , \2961_b1 );
not ( \3450_b1 , w_10984 );
not ( \3450_b0 , w_10985 );
and ( w_10984 , w_10985 , \2961_b0 );
or ( \3451_b1 , \3449_b1 , w_10986 );
or ( \3451_b0 , \3449_b0 , \3450_b0 );
not ( \3450_b0 , w_10987 );
and ( w_10987 , w_10986 , \3450_b1 );
or ( \3452_b1 , \3150_b1 , \3064_b1 );
not ( \3064_b1 , w_10988 );
and ( \3452_b0 , \3150_b0 , w_10989 );
and ( w_10988 , w_10989 , \3064_b0 );
buf ( \3453_b1 , \3452_b1 );
not ( \3453_b1 , w_10990 );
not ( \3453_b0 , w_10991 );
and ( w_10990 , w_10991 , \3452_b0 );
or ( \3454_b1 , \3041_b1 , \3053_b1 );
not ( \3053_b1 , w_10992 );
and ( \3454_b0 , \3041_b0 , w_10993 );
and ( w_10992 , w_10993 , \3053_b0 );
or ( \3455_b1 , \3454_b1 , w_10995 );
not ( w_10995 , w_10996 );
and ( \3455_b0 , \3454_b0 , w_10997 );
and ( w_10996 ,  , w_10997 );
buf ( w_10995 , \3059_b1 );
not ( w_10995 , w_10998 );
not (  , w_10999 );
and ( w_10998 , w_10999 , \3059_b0 );
buf ( \3456_b1 , \3455_b1 );
not ( \3456_b1 , w_11000 );
not ( \3456_b0 , w_11001 );
and ( w_11000 , w_11001 , \3455_b0 );
or ( \3457_b1 , \3453_b1 , w_11002 );
or ( \3457_b0 , \3453_b0 , \3456_b0 );
not ( \3456_b0 , w_11003 );
and ( w_11003 , w_11002 , \3456_b1 );
or ( \3458_b1 , \3455_b1 , w_11004 );
or ( \3458_b0 , \3455_b0 , \3452_b0 );
not ( \3452_b0 , w_11005 );
and ( w_11005 , w_11004 , \3452_b1 );
or ( \3459_b1 , \3457_b1 , w_11007 );
not ( w_11007 , w_11008 );
and ( \3459_b0 , \3457_b0 , w_11009 );
and ( w_11008 ,  , w_11009 );
buf ( w_11007 , \3458_b1 );
not ( w_11007 , w_11010 );
not (  , w_11011 );
and ( w_11010 , w_11011 , \3458_b0 );
or ( \3460_b1 , \3087_b1 , \3459_b1 );
not ( \3459_b1 , w_11012 );
and ( \3460_b0 , \3087_b0 , w_11013 );
and ( w_11012 , w_11013 , \3459_b0 );
buf ( \3461_b1 , \d[10]_b1 );
not ( \3461_b1 , w_11014 );
not ( \3461_b0 , w_11015 );
and ( w_11014 , w_11015 , \d[10]_b0 );
buf ( \3462_b1 , \1282_b1 );
not ( \3462_b1 , w_11016 );
not ( \3462_b0 , w_11017 );
and ( w_11016 , w_11017 , \1282_b0 );
or ( \3463_b1 , \3461_b1 , w_11018 );
or ( \3463_b0 , \3461_b0 , \3462_b0 );
not ( \3462_b0 , w_11019 );
and ( w_11019 , w_11018 , \3462_b1 );
or ( \3464_b1 , \1435_b1 , w_11021 );
not ( w_11021 , w_11022 );
and ( \3464_b0 , \1435_b0 , w_11023 );
and ( w_11022 ,  , w_11023 );
buf ( w_11021 , \c[10]_b1 );
not ( w_11021 , w_11024 );
not (  , w_11025 );
and ( w_11024 , w_11025 , \c[10]_b0 );
or ( \3465_b1 , \3463_b1 , w_11027 );
not ( w_11027 , w_11028 );
and ( \3465_b0 , \3463_b0 , w_11029 );
and ( w_11028 ,  , w_11029 );
buf ( w_11027 , \3464_b1 );
not ( w_11027 , w_11030 );
not (  , w_11031 );
and ( w_11030 , w_11031 , \3464_b0 );
or ( \3466_b1 , \3460_b1 , w_11033 );
not ( w_11033 , w_11034 );
and ( \3466_b0 , \3460_b0 , w_11035 );
and ( w_11034 ,  , w_11035 );
buf ( w_11033 , \3465_b1 );
not ( w_11033 , w_11036 );
not (  , w_11037 );
and ( w_11036 , w_11037 , \3465_b0 );
or ( \3467_b1 , \3451_b1 , w_11039 );
not ( w_11039 , w_11040 );
and ( \3467_b0 , \3451_b0 , w_11041 );
and ( w_11040 ,  , w_11041 );
buf ( w_11039 , \3466_b1 );
not ( w_11039 , w_11042 );
not (  , w_11043 );
and ( w_11042 , w_11043 , \3466_b0 );
or ( \3468_b1 , \3440_b1 , w_11045 );
not ( w_11045 , w_11046 );
and ( \3468_b0 , \3440_b0 , w_11047 );
and ( w_11046 ,  , w_11047 );
buf ( w_11045 , \3467_b1 );
not ( w_11045 , w_11048 );
not (  , w_11049 );
and ( w_11048 , w_11049 , \3467_b0 );
or ( \3469_b1 , \3438_b1 , w_11051 );
not ( w_11051 , w_11052 );
and ( \3469_b0 , \3438_b0 , w_11053 );
and ( w_11052 ,  , w_11053 );
buf ( w_11051 , \3468_b1 );
not ( w_11051 , w_11054 );
not (  , w_11055 );
and ( w_11054 , w_11055 , \3468_b0 );
buf ( \3470_b1 , \3469_b1 );
not ( \3470_b1 , w_11056 );
not ( \3470_b0 , w_11057 );
and ( w_11056 , w_11057 , \3469_b0 );
buf ( \3471_b1 , \2908_b1 );
not ( \3471_b1 , w_11058 );
not ( \3471_b0 , w_11059 );
and ( w_11058 , w_11059 , \2908_b0 );
or ( \3472_b1 , \3471_b1 , w_11061 );
not ( w_11061 , w_11062 );
and ( \3472_b0 , \3471_b0 , w_11063 );
and ( w_11062 ,  , w_11063 );
buf ( w_11061 , \2866_b1 );
not ( w_11061 , w_11064 );
not (  , w_11065 );
and ( w_11064 , w_11065 , \2866_b0 );
or ( \3473_b1 , \3472_b1 , w_11066 );
xor ( \3473_b0 , \3472_b0 , w_11068 );
not ( w_11068 , w_11069 );
and ( w_11069 , w_11066 , w_11067 );
buf ( w_11066 , \3199_b1 );
not ( w_11066 , w_11070 );
not ( w_11067 , w_11071 );
and ( w_11070 , w_11071 , \3199_b0 );
or ( \3474_b1 , \3473_b1 , \2936_b1 );
not ( \2936_b1 , w_11072 );
and ( \3474_b0 , \3473_b0 , w_11073 );
and ( w_11072 , w_11073 , \2936_b0 );
or ( \3475_b1 , \3187_b1 , w_11075 );
not ( w_11075 , w_11076 );
and ( \3475_b0 , \3187_b0 , w_11077 );
and ( w_11076 ,  , w_11077 );
buf ( w_11075 , \2206_b1 );
not ( w_11075 , w_11078 );
not (  , w_11079 );
and ( w_11078 , w_11079 , \2206_b0 );
or ( \3476_b1 , \3184_b1 , w_11080 );
xor ( \3476_b0 , \3184_b0 , w_11082 );
not ( w_11082 , w_11083 );
and ( w_11083 , w_11080 , w_11081 );
buf ( w_11080 , \3475_b1 );
not ( w_11080 , w_11084 );
not ( w_11081 , w_11085 );
and ( w_11084 , w_11085 , \3475_b0 );
or ( \3477_b1 , \3476_b1 , \1529_b1 );
not ( \1529_b1 , w_11086 );
and ( \3477_b0 , \3476_b0 , w_11087 );
and ( w_11086 , w_11087 , \1529_b0 );
or ( \3478_b1 , \3474_b1 , w_11089 );
not ( w_11089 , w_11090 );
and ( \3478_b0 , \3474_b0 , w_11091 );
and ( w_11090 ,  , w_11091 );
buf ( w_11089 , \3477_b1 );
not ( w_11089 , w_11092 );
not (  , w_11093 );
and ( w_11092 , w_11093 , \3477_b0 );
buf ( \3481_b1 , \d[10]_b1 );
not ( \3481_b1 , w_11094 );
not ( \3481_b0 , w_11095 );
and ( w_11094 , w_11095 , \d[10]_b0 );
buf ( \3482_b1 , \1342_b1 );
not ( \3482_b1 , w_11096 );
not ( \3482_b0 , w_11097 );
and ( w_11096 , w_11097 , \1342_b0 );
or ( \3483_b1 , \3481_b1 , w_11098 );
or ( \3483_b0 , \3481_b0 , \3482_b0 );
not ( \3482_b0 , w_11099 );
and ( w_11099 , w_11098 , \3482_b1 );
or ( \3484_b1 , \2951_b1 , w_11101 );
not ( w_11101 , w_11102 );
and ( \3484_b0 , \2951_b0 , w_11103 );
and ( w_11102 ,  , w_11103 );
buf ( w_11101 , \b[10]_b1 );
not ( w_11101 , w_11104 );
not (  , w_11105 );
and ( w_11104 , w_11105 , \b[10]_b0 );
or ( \3485_b1 , \3483_b1 , w_11107 );
not ( w_11107 , w_11108 );
and ( \3485_b0 , \3483_b0 , w_11109 );
and ( w_11108 ,  , w_11109 );
buf ( w_11107 , \3484_b1 );
not ( w_11107 , w_11110 );
not (  , w_11111 );
and ( w_11110 , w_11111 , \3484_b0 );
or ( \3486_b1 , \3480_b1 , w_11113 );
not ( w_11113 , w_11114 );
and ( \3486_b0 , \3480_b0 , w_11115 );
and ( w_11114 ,  , w_11115 );
buf ( w_11113 , \3485_b1 );
not ( w_11113 , w_11116 );
not (  , w_11117 );
and ( w_11116 , w_11117 , \3485_b0 );
or ( \3487_b1 , \3435_b1 , w_11119 );
not ( w_11119 , w_11120 );
and ( \3487_b0 , \3435_b0 , w_11121 );
and ( w_11120 ,  , w_11121 );
buf ( w_11119 , \3486_b1 );
not ( w_11119 , w_11122 );
not (  , w_11123 );
and ( w_11122 , w_11123 , \3486_b0 );
or ( \3488_b1 , \2030_b1 , w_11125 );
not ( w_11125 , w_11126 );
and ( \3488_b0 , \2030_b0 , w_11127 );
and ( w_11126 ,  , w_11127 );
buf ( w_11125 , \1962_b1 );
not ( w_11125 , w_11128 );
not (  , w_11129 );
and ( w_11128 , w_11129 , \1962_b0 );
buf ( \3489_b1 , \3488_b1 );
not ( \3489_b1 , w_11130 );
not ( \3489_b0 , w_11131 );
and ( w_11130 , w_11131 , \3488_b0 );
or ( \3490_b1 , \3489_b1 , w_11133 );
not ( w_11133 , w_11134 );
and ( \3490_b0 , \3489_b0 , w_11135 );
and ( w_11134 ,  , w_11135 );
buf ( w_11133 , \2031_b1 );
not ( w_11133 , w_11136 );
not (  , w_11137 );
and ( w_11136 , w_11137 , \2031_b0 );
buf ( \3491_b1 , \3490_b1 );
not ( \3491_b1 , w_11138 );
not ( \3491_b0 , w_11139 );
and ( w_11138 , w_11139 , \3490_b0 );
buf ( \3492_b1 , \2193_b1 );
not ( \3492_b1 , w_11140 );
not ( \3492_b0 , w_11141 );
and ( w_11140 , w_11141 , \2193_b0 );
buf ( \3494_b1 , \3493_b1 );
not ( \3494_b1 , w_11142 );
not ( \3494_b0 , w_11143 );
and ( w_11142 , w_11143 , \3493_b0 );
or ( \3495_b1 , \3492_b1 , w_11144 );
or ( \3495_b0 , \3492_b0 , \3494_b0 );
not ( \3494_b0 , w_11145 );
and ( w_11145 , w_11144 , \3494_b1 );
or ( \3496_b1 , \2205_b1 , \2211_b1 );
not ( \2211_b1 , w_11146 );
and ( \3496_b0 , \2205_b0 , w_11147 );
and ( w_11146 , w_11147 , \2211_b0 );
or ( \3497_b1 , \3496_b1 , w_11149 );
not ( w_11149 , w_11150 );
and ( \3497_b0 , \3496_b0 , w_11151 );
and ( w_11150 ,  , w_11151 );
buf ( w_11149 , \2221_b1 );
not ( w_11149 , w_11152 );
not (  , w_11153 );
and ( w_11152 , w_11153 , \2221_b0 );
or ( \3498_b1 , \3495_b1 , w_11155 );
not ( w_11155 , w_11156 );
and ( \3498_b0 , \3495_b0 , w_11157 );
and ( w_11156 ,  , w_11157 );
buf ( w_11155 , \3497_b1 );
not ( w_11155 , w_11158 );
not (  , w_11159 );
and ( w_11158 , w_11159 , \3497_b0 );
buf ( \3499_b1 , \3498_b1 );
not ( \3499_b1 , w_11160 );
not ( \3499_b0 , w_11161 );
and ( w_11160 , w_11161 , \3498_b0 );
or ( \3500_b1 , \3491_b1 , w_11162 );
or ( \3500_b0 , \3491_b0 , \3499_b0 );
not ( \3499_b0 , w_11163 );
and ( w_11163 , w_11162 , \3499_b1 );
or ( \3501_b1 , \3490_b1 , w_11164 );
or ( \3501_b0 , \3490_b0 , \3498_b0 );
not ( \3498_b0 , w_11165 );
and ( w_11165 , w_11164 , \3498_b1 );
or ( \3502_b1 , \3500_b1 , w_11167 );
not ( w_11167 , w_11168 );
and ( \3502_b0 , \3500_b0 , w_11169 );
and ( w_11168 ,  , w_11169 );
buf ( w_11167 , \3501_b1 );
not ( w_11167 , w_11170 );
not (  , w_11171 );
and ( w_11170 , w_11171 , \3501_b0 );
or ( \3503_b1 , \3502_b1 , w_11173 );
not ( w_11173 , w_11174 );
and ( \3503_b0 , \3502_b0 , w_11175 );
and ( w_11174 ,  , w_11175 );
buf ( w_11173 , \1529_b1 );
not ( w_11173 , w_11176 );
not (  , w_11177 );
and ( w_11176 , w_11177 , \1529_b0 );
or ( \3504_b1 , \2669_b1 , w_11179 );
not ( w_11179 , w_11180 );
and ( \3504_b0 , \2669_b0 , w_11181 );
and ( w_11180 ,  , w_11181 );
buf ( w_11179 , \2727_b1 );
not ( w_11179 , w_11182 );
not (  , w_11183 );
and ( w_11182 , w_11183 , \2727_b0 );
buf ( \3505_b1 , \3504_b1 );
not ( \3505_b1 , w_11184 );
not ( \3505_b0 , w_11185 );
and ( w_11184 , w_11185 , \3504_b0 );
or ( \3506_b1 , \3505_b1 , w_11187 );
not ( w_11187 , w_11188 );
and ( \3506_b0 , \3505_b0 , w_11189 );
and ( w_11188 ,  , w_11189 );
buf ( w_11187 , \3280_b1 );
not ( w_11187 , w_11190 );
not (  , w_11191 );
and ( w_11190 , w_11191 , \3280_b0 );
buf ( \3507_b1 , \3506_b1 );
not ( \3507_b1 , w_11192 );
not ( \3507_b0 , w_11193 );
and ( w_11192 , w_11193 , \3506_b0 );
or ( \3508_b1 , \2913_b1 , w_11195 );
not ( w_11195 , w_11196 );
and ( \3508_b0 , \2913_b0 , w_11197 );
and ( w_11196 ,  , w_11197 );
buf ( w_11195 , \2914_b1 );
not ( w_11195 , w_11198 );
not (  , w_11199 );
and ( w_11198 , w_11199 , \2914_b0 );
buf ( \3509_b1 , \2826_b1 );
not ( \3509_b1 , w_11200 );
not ( \3509_b0 , w_11201 );
and ( w_11200 , w_11201 , \2826_b0 );
buf ( \3510_b1 , \2830_b1 );
not ( \3510_b1 , w_11202 );
not ( \3510_b0 , w_11203 );
and ( w_11202 , w_11203 , \2830_b0 );
or ( \3511_b1 , \3509_b1 , w_11204 );
or ( \3511_b0 , \3509_b0 , \3510_b0 );
not ( \3510_b0 , w_11205 );
and ( w_11205 , w_11204 , \3510_b1 );
or ( \3512_b1 , \3511_b1 , w_11207 );
not ( w_11207 , w_11208 );
and ( \3512_b0 , \3511_b0 , w_11209 );
and ( w_11208 ,  , w_11209 );
buf ( w_11207 , \2866_b1 );
not ( w_11207 , w_11210 );
not (  , w_11211 );
and ( w_11210 , w_11211 , \2866_b0 );
buf ( \3513_b1 , \3512_b1 );
not ( \3513_b1 , w_11212 );
not ( \3513_b0 , w_11213 );
and ( w_11212 , w_11213 , \3512_b0 );
buf ( \3516_b1 , \3515_b1 );
not ( \3516_b1 , w_11214 );
not ( \3516_b0 , w_11215 );
and ( w_11214 , w_11215 , \3515_b0 );
or ( \3517_b1 , \3507_b1 , w_11216 );
or ( \3517_b0 , \3507_b0 , \3516_b0 );
not ( \3516_b0 , w_11217 );
and ( w_11217 , w_11216 , \3516_b1 );
or ( \3518_b1 , \3515_b1 , w_11218 );
or ( \3518_b0 , \3515_b0 , \3506_b0 );
not ( \3506_b0 , w_11219 );
and ( w_11219 , w_11218 , \3506_b1 );
or ( \3519_b1 , \3517_b1 , w_11221 );
not ( w_11221 , w_11222 );
and ( \3519_b0 , \3517_b0 , w_11223 );
and ( w_11222 ,  , w_11223 );
buf ( w_11221 , \3518_b1 );
not ( w_11221 , w_11224 );
not (  , w_11225 );
and ( w_11224 , w_11225 , \3518_b0 );
or ( \3520_b1 , \3519_b1 , w_11227 );
not ( w_11227 , w_11228 );
and ( \3520_b0 , \3519_b0 , w_11229 );
and ( w_11228 ,  , w_11229 );
buf ( w_11227 , \2936_b1 );
not ( w_11227 , w_11230 );
not (  , w_11231 );
and ( w_11230 , w_11231 , \2936_b0 );
or ( \3521_b1 , \3503_b1 , w_11233 );
not ( w_11233 , w_11234 );
and ( \3521_b0 , \3503_b0 , w_11235 );
and ( w_11234 ,  , w_11235 );
buf ( w_11233 , \3520_b1 );
not ( w_11233 , w_11236 );
not (  , w_11237 );
and ( w_11236 , w_11237 , \3520_b0 );
buf ( \3522_b1 , \b[13]_b1 );
not ( \3522_b1 , w_11238 );
not ( \3522_b0 , w_11239 );
and ( w_11238 , w_11239 , \b[13]_b0 );
buf ( \3523_b1 , \3124_b1 );
not ( \3523_b1 , w_11240 );
not ( \3523_b0 , w_11241 );
and ( w_11240 , w_11241 , \3124_b0 );
or ( \3524_b1 , \3522_b1 , w_11242 );
or ( \3524_b0 , \3522_b0 , \3523_b0 );
not ( \3523_b0 , w_11243 );
and ( w_11243 , w_11242 , \3523_b1 );
or ( \3525_b1 , \a[13]_b1 , \1466_b1 );
not ( \1466_b1 , w_11244 );
and ( \3525_b0 , \a[13]_b0 , w_11245 );
and ( w_11244 , w_11245 , \1466_b0 );
or ( \3526_b1 , \c[13]_b1 , \d[13]_b1 );
xor ( \3526_b0 , \c[13]_b0 , w_11246 );
not ( w_11246 , w_11247 );
and ( w_11247 , \d[13]_b1 , \d[13]_b0 );
buf ( \3527_b1 , \3526_b1 );
not ( \3527_b1 , w_11248 );
not ( \3527_b0 , w_11249 );
and ( w_11248 , w_11249 , \3526_b0 );
buf ( \3528_b1 , \1383_b1 );
not ( \3528_b1 , w_11250 );
not ( \3528_b0 , w_11251 );
and ( w_11250 , w_11251 , \1383_b0 );
or ( \3529_b1 , \3527_b1 , w_11252 );
or ( \3529_b0 , \3527_b0 , \3528_b0 );
not ( \3528_b0 , w_11253 );
and ( w_11253 , w_11252 , \3528_b1 );
buf ( \3530_b1 , \3012_b1 );
not ( \3530_b1 , w_11254 );
not ( \3530_b0 , w_11255 );
and ( w_11254 , w_11255 , \3012_b0 );
or ( \3531_b1 , \3530_b1 , w_11257 );
not ( w_11257 , w_11258 );
and ( \3531_b0 , \3530_b0 , w_11259 );
and ( w_11258 ,  , w_11259 );
buf ( w_11257 , \2980_b1 );
not ( w_11257 , w_11260 );
not (  , w_11261 );
and ( w_11260 , w_11261 , \2980_b0 );
buf ( \3532_b1 , \3531_b1 );
not ( \3532_b1 , w_11262 );
not ( \3532_b0 , w_11263 );
and ( w_11262 , w_11263 , \3531_b0 );
buf ( \3533_b1 , \2981_b1 );
not ( \3533_b1 , w_11264 );
not ( \3533_b0 , w_11265 );
and ( w_11264 , w_11265 , \2981_b0 );
or ( \3535_b1 , \3007_b1 , w_11267 );
not ( w_11267 , w_11268 );
and ( \3535_b0 , \3007_b0 , w_11269 );
and ( w_11268 ,  , w_11269 );
buf ( w_11267 , \3533_b1 );
not ( w_11267 , w_11270 );
not (  , w_11271 );
and ( w_11270 , w_11271 , \3533_b0 );
or ( \3536_b1 , \3535_b1 , w_11273 );
not ( w_11273 , w_11274 );
and ( \3536_b0 , \3535_b0 , w_11275 );
and ( w_11274 ,  , w_11275 );
buf ( w_11273 , \3010_b1 );
not ( w_11273 , w_11276 );
not (  , w_11277 );
and ( w_11276 , w_11277 , \3010_b0 );
or ( \3537_b1 , \3534_b1 , w_11279 );
not ( w_11279 , w_11280 );
and ( \3537_b0 , \3534_b0 , w_11281 );
and ( w_11280 ,  , w_11281 );
buf ( w_11279 , \3536_b1 );
not ( w_11279 , w_11282 );
not (  , w_11283 );
and ( w_11282 , w_11283 , \3536_b0 );
buf ( \3538_b1 , \3537_b1 );
not ( \3538_b1 , w_11284 );
not ( \3538_b0 , w_11285 );
and ( w_11284 , w_11285 , \3537_b0 );
or ( \3539_b1 , \3532_b1 , w_11286 );
or ( \3539_b0 , \3532_b0 , \3538_b0 );
not ( \3538_b0 , w_11287 );
and ( w_11287 , w_11286 , \3538_b1 );
or ( \3540_b1 , \3537_b1 , w_11288 );
or ( \3540_b0 , \3537_b0 , \3531_b0 );
not ( \3531_b0 , w_11289 );
and ( w_11289 , w_11288 , \3531_b1 );
or ( \3541_b1 , \3539_b1 , w_11291 );
not ( w_11291 , w_11292 );
and ( \3541_b0 , \3539_b0 , w_11293 );
and ( w_11292 ,  , w_11293 );
buf ( w_11291 , \3540_b1 );
not ( w_11291 , w_11294 );
not (  , w_11295 );
and ( w_11294 , w_11295 , \3540_b0 );
or ( \3542_b1 , \2961_b1 , \3541_b1 );
not ( \3541_b1 , w_11296 );
and ( \3542_b0 , \2961_b0 , w_11297 );
and ( w_11296 , w_11297 , \3541_b0 );
buf ( \3543_b1 , \3074_b1 );
not ( \3543_b1 , w_11298 );
not ( \3543_b0 , w_11299 );
and ( w_11298 , w_11299 , \3074_b0 );
or ( \3544_b1 , \3543_b1 , w_11301 );
not ( w_11301 , w_11302 );
and ( \3544_b0 , \3543_b0 , w_11303 );
and ( w_11302 ,  , w_11303 );
buf ( w_11301 , \3042_b1 );
not ( w_11301 , w_11304 );
not (  , w_11305 );
and ( w_11304 , w_11305 , \3042_b0 );
buf ( \3545_b1 , \3544_b1 );
not ( \3545_b1 , w_11306 );
not ( \3545_b0 , w_11307 );
and ( w_11306 , w_11307 , \3544_b0 );
buf ( \3546_b1 , \3043_b1 );
not ( \3546_b1 , w_11308 );
not ( \3546_b0 , w_11309 );
and ( w_11308 , w_11309 , \3043_b0 );
or ( \3548_b1 , \3069_b1 , w_11311 );
not ( w_11311 , w_11312 );
and ( \3548_b0 , \3069_b0 , w_11313 );
and ( w_11312 ,  , w_11313 );
buf ( w_11311 , \3546_b1 );
not ( w_11311 , w_11314 );
not (  , w_11315 );
and ( w_11314 , w_11315 , \3546_b0 );
or ( \3549_b1 , \3548_b1 , w_11317 );
not ( w_11317 , w_11318 );
and ( \3549_b0 , \3548_b0 , w_11319 );
and ( w_11318 ,  , w_11319 );
buf ( w_11317 , \3072_b1 );
not ( w_11317 , w_11320 );
not (  , w_11321 );
and ( w_11320 , w_11321 , \3072_b0 );
or ( \3550_b1 , \3547_b1 , w_11323 );
not ( w_11323 , w_11324 );
and ( \3550_b0 , \3547_b0 , w_11325 );
and ( w_11324 ,  , w_11325 );
buf ( w_11323 , \3549_b1 );
not ( w_11323 , w_11326 );
not (  , w_11327 );
and ( w_11326 , w_11327 , \3549_b0 );
buf ( \3551_b1 , \3550_b1 );
not ( \3551_b1 , w_11328 );
not ( \3551_b0 , w_11329 );
and ( w_11328 , w_11329 , \3550_b0 );
or ( \3552_b1 , \3545_b1 , w_11330 );
or ( \3552_b0 , \3545_b0 , \3551_b0 );
not ( \3551_b0 , w_11331 );
and ( w_11331 , w_11330 , \3551_b1 );
or ( \3553_b1 , \3550_b1 , w_11332 );
or ( \3553_b0 , \3550_b0 , \3544_b0 );
not ( \3544_b0 , w_11333 );
and ( w_11333 , w_11332 , \3544_b1 );
or ( \3554_b1 , \3552_b1 , w_11335 );
not ( w_11335 , w_11336 );
and ( \3554_b0 , \3552_b0 , w_11337 );
and ( w_11336 ,  , w_11337 );
buf ( w_11335 , \3553_b1 );
not ( w_11335 , w_11338 );
not (  , w_11339 );
and ( w_11338 , w_11339 , \3553_b0 );
buf ( \3555_b1 , \3554_b1 );
not ( \3555_b1 , w_11340 );
not ( \3555_b0 , w_11341 );
and ( w_11340 , w_11341 , \3554_b0 );
buf ( \3556_b1 , \3087_b1 );
not ( \3556_b1 , w_11342 );
not ( \3556_b0 , w_11343 );
and ( w_11342 , w_11343 , \3087_b0 );
or ( \3557_b1 , \3555_b1 , w_11344 );
or ( \3557_b0 , \3555_b0 , \3556_b0 );
not ( \3556_b0 , w_11345 );
and ( w_11345 , w_11344 , \3556_b1 );
or ( \3558_b1 , \1282_b1 , \d[13]_b1 );
not ( \d[13]_b1 , w_11346 );
and ( \3558_b0 , \1282_b0 , w_11347 );
and ( w_11346 , w_11347 , \d[13]_b0 );
or ( \3559_b1 , \1514_b1 , \c[13]_b1 );
not ( \c[13]_b1 , w_11348 );
and ( \3559_b0 , \1514_b0 , w_11349 );
and ( w_11348 , w_11349 , \c[13]_b0 );
or ( \3560_b1 , \3558_b1 , w_11351 );
not ( w_11351 , w_11352 );
and ( \3560_b0 , \3558_b0 , w_11353 );
and ( w_11352 ,  , w_11353 );
buf ( w_11351 , \3559_b1 );
not ( w_11351 , w_11354 );
not (  , w_11355 );
and ( w_11354 , w_11355 , \3559_b0 );
or ( \3561_b1 , \3557_b1 , w_11357 );
not ( w_11357 , w_11358 );
and ( \3561_b0 , \3557_b0 , w_11359 );
and ( w_11358 ,  , w_11359 );
buf ( w_11357 , \3560_b1 );
not ( w_11357 , w_11360 );
not (  , w_11361 );
and ( w_11360 , w_11361 , \3560_b0 );
or ( \3562_b1 , \3542_b1 , w_11363 );
not ( w_11363 , w_11364 );
and ( \3562_b0 , \3542_b0 , w_11365 );
and ( w_11364 ,  , w_11365 );
buf ( w_11363 , \3561_b1 );
not ( w_11363 , w_11366 );
not (  , w_11367 );
and ( w_11366 , w_11367 , \3561_b0 );
or ( \3563_b1 , \3529_b1 , w_11369 );
not ( w_11369 , w_11370 );
and ( \3563_b0 , \3529_b0 , w_11371 );
and ( w_11370 ,  , w_11371 );
buf ( w_11369 , \3562_b1 );
not ( w_11369 , w_11372 );
not (  , w_11373 );
and ( w_11372 , w_11373 , \3562_b0 );
or ( \3564_b1 , \3525_b1 , w_11375 );
not ( w_11375 , w_11376 );
and ( \3564_b0 , \3525_b0 , w_11377 );
and ( w_11376 ,  , w_11377 );
buf ( w_11375 , \3563_b1 );
not ( w_11375 , w_11378 );
not (  , w_11379 );
and ( w_11378 , w_11379 , \3563_b0 );
or ( \3565_b1 , \3524_b1 , w_11381 );
not ( w_11381 , w_11382 );
and ( \3565_b0 , \3524_b0 , w_11383 );
and ( w_11382 ,  , w_11383 );
buf ( w_11381 , \3564_b1 );
not ( w_11381 , w_11384 );
not (  , w_11385 );
and ( w_11384 , w_11385 , \3564_b0 );
buf ( \3566_b1 , \3565_b1 );
not ( \3566_b1 , w_11386 );
not ( \3566_b0 , w_11387 );
and ( w_11386 , w_11387 , \3565_b0 );
or ( \3567_b1 , \1338_b1 , w_11389 );
not ( w_11389 , w_11390 );
and ( \3567_b0 , \1338_b0 , w_11391 );
and ( w_11390 ,  , w_11391 );
buf ( w_11389 , \a[13]_b1 );
not ( w_11389 , w_11392 );
not (  , w_11393 );
and ( w_11392 , w_11393 , \a[13]_b0 );
buf ( \3568_b1 , \3101_b1 );
not ( \3568_b1 , w_11394 );
not ( \3568_b0 , w_11395 );
and ( w_11394 , w_11395 , \3101_b0 );
or ( \3569_b1 , \b[13]_b1 , w_11397 );
not ( w_11397 , w_11398 );
and ( \3569_b0 , \b[13]_b0 , w_11399 );
and ( w_11398 ,  , w_11399 );
buf ( w_11397 , \c[13]_b1 );
not ( w_11397 , w_11400 );
not (  , w_11401 );
and ( w_11400 , w_11401 , \c[13]_b0 );
buf ( \3570_b1 , \3569_b1 );
not ( \3570_b1 , w_11402 );
not ( \3570_b0 , w_11403 );
and ( w_11402 , w_11403 , \3569_b0 );
or ( \3571_b1 , \3568_b1 , \3570_b1 );
not ( \3570_b1 , w_11404 );
and ( \3571_b0 , \3568_b0 , w_11405 );
and ( w_11404 , w_11405 , \3570_b0 );
or ( \3572_b1 , \a[13]_b1 , w_11406 );
or ( \3572_b0 , \a[13]_b0 , \d[13]_b0 );
not ( \d[13]_b0 , w_11407 );
and ( w_11407 , w_11406 , \d[13]_b1 );
or ( \3573_b1 , \1457_b1 , \3572_b1 );
not ( \3572_b1 , w_11408 );
and ( \3573_b0 , \1457_b0 , w_11409 );
and ( w_11408 , w_11409 , \3572_b0 );
or ( \3574_b1 , \3571_b1 , w_11411 );
not ( w_11411 , w_11412 );
and ( \3574_b0 , \3571_b0 , w_11413 );
and ( w_11412 ,  , w_11413 );
buf ( w_11411 , \3573_b1 );
not ( w_11411 , w_11414 );
not (  , w_11415 );
and ( w_11414 , w_11415 , \3573_b0 );
or ( \3576_b1 , \3521_b1 , w_11417 );
not ( w_11417 , w_11418 );
and ( \3576_b0 , \3521_b0 , w_11419 );
and ( w_11418 ,  , w_11419 );
buf ( w_11417 , \3575_b1 );
not ( w_11417 , w_11420 );
not (  , w_11421 );
and ( w_11420 , w_11421 , \3575_b0 );
buf ( \3577_b1 , \3576_b1 );
not ( \3577_b1 , w_11422 );
not ( \3577_b0 , w_11423 );
and ( w_11422 , w_11423 , \3576_b0 );
buf ( \3578_b1 , \a[0]_b1 );
not ( \3578_b1 , w_11424 );
not ( \3578_b0 , w_11425 );
and ( w_11424 , w_11425 , \a[0]_b0 );
buf ( \3579_b1 , \2946_b1 );
not ( \3579_b1 , w_11426 );
not ( \3579_b0 , w_11427 );
and ( w_11426 , w_11427 , \2946_b0 );
or ( \3580_b1 , \3578_b1 , w_11428 );
or ( \3580_b0 , \3578_b0 , \3579_b0 );
not ( \3579_b0 , w_11429 );
and ( w_11429 , w_11428 , \3579_b1 );
buf ( \3581_b1 , \d[0]_b1 );
not ( \3581_b1 , w_11430 );
not ( \3581_b0 , w_11431 );
and ( w_11430 , w_11431 , \d[0]_b0 );
buf ( \3582_b1 , \1457_b1 );
not ( \3582_b1 , w_11432 );
not ( \3582_b0 , w_11433 );
and ( w_11432 , w_11433 , \1457_b0 );
or ( \3583_b1 , \3581_b1 , w_11434 );
or ( \3583_b0 , \3581_b0 , \3582_b0 );
not ( \3582_b0 , w_11435 );
and ( w_11435 , w_11434 , \3582_b1 );
or ( \3584_b1 , \c[0]_b1 , \d[0]_b1 );
xor ( \3584_b0 , \c[0]_b0 , w_11436 );
not ( w_11436 , w_11437 );
and ( w_11437 , \d[0]_b1 , \d[0]_b0 );
or ( \3585_b1 , \3305_b1 , \3584_b1 );
not ( \3584_b1 , w_11438 );
and ( \3585_b0 , \3305_b0 , w_11439 );
and ( w_11438 , w_11439 , \3584_b0 );
buf ( \3586_b1 , \1044_b1 );
not ( \3586_b1 , w_11440 );
not ( \3586_b0 , w_11441 );
and ( w_11440 , w_11441 , \1044_b0 );
buf ( \3587_b1 , \3586_b1 );
not ( \3587_b1 , w_11442 );
not ( \3587_b0 , w_11443 );
and ( w_11442 , w_11443 , \3586_b0 );
buf ( \3588_b1 , \1529_b1 );
not ( \3588_b1 , w_11444 );
not ( \3588_b0 , w_11445 );
and ( w_11444 , w_11445 , \1529_b0 );
or ( \3589_b1 , \3587_b1 , w_11446 );
or ( \3589_b0 , \3587_b0 , \3588_b0 );
not ( \3588_b0 , w_11447 );
and ( w_11447 , w_11446 , \3588_b1 );
or ( \3590_b1 , \b[0]_b1 , \d[0]_b1 );
xor ( \3590_b0 , \b[0]_b0 , w_11448 );
not ( w_11448 , w_11449 );
and ( w_11449 , \d[0]_b1 , \d[0]_b0 );
or ( \3591_b1 , \2961_b1 , \3590_b1 );
not ( \3590_b1 , w_11450 );
and ( \3591_b0 , \2961_b0 , w_11451 );
and ( w_11450 , w_11451 , \3590_b0 );
or ( \3592_b1 , \a[0]_b1 , \c[0]_b1 );
xor ( \3592_b0 , \a[0]_b0 , w_11452 );
not ( w_11452 , w_11453 );
and ( w_11453 , \c[0]_b1 , \c[0]_b0 );
buf ( \3593_b1 , \3592_b1 );
not ( \3593_b1 , w_11454 );
not ( \3593_b0 , w_11455 );
and ( w_11454 , w_11455 , \3592_b0 );
buf ( \3594_b1 , \3087_b1 );
not ( \3594_b1 , w_11456 );
not ( \3594_b0 , w_11457 );
and ( w_11456 , w_11457 , \3087_b0 );
or ( \3595_b1 , \3593_b1 , w_11458 );
or ( \3595_b0 , \3593_b0 , \3594_b0 );
not ( \3594_b0 , w_11459 );
and ( w_11459 , w_11458 , \3594_b1 );
or ( \3596_b1 , \1282_b1 , w_11461 );
not ( w_11461 , w_11462 );
and ( \3596_b0 , \1282_b0 , w_11463 );
and ( w_11462 ,  , w_11463 );
buf ( w_11461 , \d[0]_b1 );
not ( w_11461 , w_11464 );
not (  , w_11465 );
and ( w_11464 , w_11465 , \d[0]_b0 );
or ( \3597_b1 , \1293_b1 , \b[0]_b1 );
not ( \b[0]_b1 , w_11466 );
and ( \3597_b0 , \1293_b0 , w_11467 );
and ( w_11466 , w_11467 , \b[0]_b0 );
or ( \3598_b1 , \1435_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_11468 );
and ( \3598_b0 , \1435_b0 , w_11469 );
and ( w_11468 , w_11469 , \c[0]_b0 );
or ( \3599_b1 , \3597_b1 , w_11471 );
not ( w_11471 , w_11472 );
and ( \3599_b0 , \3597_b0 , w_11473 );
and ( w_11472 ,  , w_11473 );
buf ( w_11471 , \3598_b1 );
not ( w_11471 , w_11474 );
not (  , w_11475 );
and ( w_11474 , w_11475 , \3598_b0 );
or ( \3600_b1 , \3596_b1 , \3599_b1 );
not ( \3599_b1 , w_11476 );
and ( \3600_b0 , \3596_b0 , w_11477 );
and ( w_11476 , w_11477 , \3599_b0 );
or ( \3601_b1 , \3595_b1 , w_11479 );
not ( w_11479 , w_11480 );
and ( \3601_b0 , \3595_b0 , w_11481 );
and ( w_11480 ,  , w_11481 );
buf ( w_11479 , \3600_b1 );
not ( w_11479 , w_11482 );
not (  , w_11483 );
and ( w_11482 , w_11483 , \3600_b0 );
or ( \3602_b1 , \3591_b1 , w_11485 );
not ( w_11485 , w_11486 );
and ( \3602_b0 , \3591_b0 , w_11487 );
and ( w_11486 ,  , w_11487 );
buf ( w_11485 , \3601_b1 );
not ( w_11485 , w_11488 );
not (  , w_11489 );
and ( w_11488 , w_11489 , \3601_b0 );
or ( \3603_b1 , \3589_b1 , w_11491 );
not ( w_11491 , w_11492 );
and ( \3603_b0 , \3589_b0 , w_11493 );
and ( w_11492 ,  , w_11493 );
buf ( w_11491 , \3602_b1 );
not ( w_11491 , w_11494 );
not (  , w_11495 );
and ( w_11494 , w_11495 , \3602_b0 );
or ( \3604_b1 , \3585_b1 , w_11497 );
not ( w_11497 , w_11498 );
and ( \3604_b0 , \3585_b0 , w_11499 );
and ( w_11498 ,  , w_11499 );
buf ( w_11497 , \3603_b1 );
not ( w_11497 , w_11500 );
not (  , w_11501 );
and ( w_11500 , w_11501 , \3603_b0 );
or ( \3605_b1 , \3583_b1 , w_11503 );
not ( w_11503 , w_11504 );
and ( \3605_b0 , \3583_b0 , w_11505 );
and ( w_11504 ,  , w_11505 );
buf ( w_11503 , \3604_b1 );
not ( w_11503 , w_11506 );
not (  , w_11507 );
and ( w_11506 , w_11507 , \3604_b0 );
or ( \3606_b1 , \b[0]_b1 , \c[0]_b1 );
not ( \c[0]_b1 , w_11508 );
and ( \3606_b0 , \b[0]_b0 , w_11509 );
and ( w_11508 , w_11509 , \c[0]_b0 );
buf ( \3607_b1 , \3606_b1 );
not ( \3607_b1 , w_11510 );
not ( \3607_b0 , w_11511 );
and ( w_11510 , w_11511 , \3606_b0 );
buf ( \3608_b1 , \3102_b1 );
not ( \3608_b1 , w_11512 );
not ( \3608_b0 , w_11513 );
and ( w_11512 , w_11513 , \3102_b0 );
or ( \3609_b1 , \3607_b1 , w_11514 );
or ( \3609_b0 , \3607_b0 , \3608_b0 );
not ( \3608_b0 , w_11515 );
and ( w_11515 , w_11514 , \3608_b1 );
or ( \3610_b1 , \a[0]_b1 , w_11516 );
or ( \3610_b0 , \a[0]_b0 , \b[0]_b0 );
not ( \b[0]_b0 , w_11517 );
and ( w_11517 , w_11516 , \b[0]_b1 );
or ( \3611_b1 , \2954_b1 , \3610_b1 );
not ( \3610_b1 , w_11518 );
and ( \3611_b0 , \2954_b0 , w_11519 );
and ( w_11518 , w_11519 , \3610_b0 );
buf ( \3612_b1 , \852_b1 );
not ( \3612_b1 , w_11520 );
not ( \3612_b0 , w_11521 );
and ( w_11520 , w_11521 , \852_b0 );
or ( \3613_b1 , \2936_b1 , \3612_b1 );
not ( \3612_b1 , w_11522 );
and ( \3613_b0 , \2936_b0 , w_11523 );
and ( w_11522 , w_11523 , \3612_b0 );
or ( \3614_b1 , \3611_b1 , w_11525 );
not ( w_11525 , w_11526 );
and ( \3614_b0 , \3611_b0 , w_11527 );
and ( w_11526 ,  , w_11527 );
buf ( w_11525 , \3613_b1 );
not ( w_11525 , w_11528 );
not (  , w_11529 );
and ( w_11528 , w_11529 , \3613_b0 );
or ( \3615_b1 , \3609_b1 , w_11531 );
not ( w_11531 , w_11532 );
and ( \3615_b0 , \3609_b0 , w_11533 );
and ( w_11532 ,  , w_11533 );
buf ( w_11531 , \3614_b1 );
not ( w_11531 , w_11534 );
not (  , w_11535 );
and ( w_11534 , w_11535 , \3614_b0 );
or ( \3616_b1 , \3605_b1 , w_11537 );
not ( w_11537 , w_11538 );
and ( \3616_b0 , \3605_b0 , w_11539 );
and ( w_11538 ,  , w_11539 );
buf ( w_11537 , \3615_b1 );
not ( w_11537 , w_11540 );
not (  , w_11541 );
and ( w_11540 , w_11541 , \3615_b0 );
or ( \3617_b1 , \3580_b1 , w_11543 );
not ( w_11543 , w_11544 );
and ( \3617_b0 , \3580_b0 , w_11545 );
and ( w_11544 ,  , w_11545 );
buf ( w_11543 , \3616_b1 );
not ( w_11543 , w_11546 );
not (  , w_11547 );
and ( w_11546 , w_11547 , \3616_b0 );
buf ( \3618_b1 , \a[8]_b1 );
not ( \3618_b1 , w_11548 );
not ( \3618_b0 , w_11549 );
and ( w_11548 , w_11549 , \a[8]_b0 );
buf ( \3619_b1 , \2946_b1 );
not ( \3619_b1 , w_11550 );
not ( \3619_b0 , w_11551 );
and ( w_11550 , w_11551 , \2946_b0 );
or ( \3620_b1 , \3618_b1 , w_11552 );
or ( \3620_b0 , \3618_b0 , \3619_b0 );
not ( \3619_b0 , w_11553 );
and ( w_11553 , w_11552 , \3619_b1 );
buf ( \3621_b1 , \645_b1 );
not ( \3621_b1 , w_11554 );
not ( \3621_b0 , w_11555 );
and ( w_11554 , w_11555 , \645_b0 );
or ( \3622_b1 , \3621_b1 , \d[8]_b1 );
not ( \d[8]_b1 , w_11556 );
and ( \3622_b0 , \3621_b0 , w_11557 );
and ( w_11556 , w_11557 , \d[8]_b0 );
buf ( \3623_b1 , \782_b1 );
not ( \3623_b1 , w_11558 );
not ( \3623_b0 , w_11559 );
and ( w_11558 , w_11559 , \782_b0 );
buf ( \3624_b1 , \904_b1 );
not ( \3624_b1 , w_11560 );
not ( \3624_b0 , w_11561 );
and ( w_11560 , w_11561 , \904_b0 );
or ( \3625_b1 , \3623_b1 , w_11562 );
or ( \3625_b0 , \3623_b0 , \3624_b0 );
not ( \3624_b0 , w_11563 );
and ( w_11563 , w_11562 , \3624_b1 );
or ( \3626_b1 , \3625_b1 , w_11565 );
not ( w_11565 , w_11566 );
and ( \3626_b0 , \3625_b0 , w_11567 );
and ( w_11566 ,  , w_11567 );
buf ( w_11565 , \783_b1 );
not ( w_11565 , w_11568 );
not (  , w_11569 );
and ( w_11568 , w_11569 , \783_b0 );
buf ( \3627_b1 , \2903_b1 );
not ( \3627_b1 , w_11570 );
not ( \3627_b0 , w_11571 );
and ( w_11570 , w_11571 , \2903_b0 );
or ( \3628_b1 , \3627_b1 , w_11573 );
not ( w_11573 , w_11574 );
and ( \3628_b0 , \3627_b0 , w_11575 );
and ( w_11574 ,  , w_11575 );
buf ( w_11573 , \2900_b1 );
not ( w_11573 , w_11576 );
not (  , w_11577 );
and ( w_11576 , w_11577 , \2900_b0 );
or ( \3629_b1 , \3626_b1 , w_11578 );
xor ( \3629_b0 , \3626_b0 , w_11580 );
not ( w_11580 , w_11581 );
and ( w_11581 , w_11578 , w_11579 );
buf ( w_11578 , \3628_b1 );
not ( w_11578 , w_11582 );
not ( w_11579 , w_11583 );
and ( w_11582 , w_11583 , \3628_b0 );
buf ( \3630_b1 , \3629_b1 );
not ( \3630_b1 , w_11584 );
not ( \3630_b0 , w_11585 );
and ( w_11584 , w_11585 , \3629_b0 );
buf ( \3631_b1 , \916_b1 );
not ( \3631_b1 , w_11586 );
not ( \3631_b0 , w_11587 );
and ( w_11586 , w_11587 , \916_b0 );
or ( \3632_b1 , \3630_b1 , w_11588 );
or ( \3632_b0 , \3630_b0 , \3631_b0 );
not ( \3631_b0 , w_11589 );
and ( w_11589 , w_11588 , \3631_b1 );
buf ( \3633_b1 , \2172_b1 );
not ( \3633_b1 , w_11590 );
not ( \3633_b0 , w_11591 );
and ( w_11590 , w_11591 , \2172_b0 );
or ( \3634_b1 , \3633_b1 , w_11593 );
not ( w_11593 , w_11594 );
and ( \3634_b0 , \3633_b0 , w_11595 );
and ( w_11594 ,  , w_11595 );
buf ( w_11593 , \2188_b1 );
not ( w_11593 , w_11596 );
not (  , w_11597 );
and ( w_11596 , w_11597 , \2188_b0 );
buf ( \3635_b1 , \3634_b1 );
not ( \3635_b1 , w_11598 );
not ( \3635_b0 , w_11599 );
and ( w_11598 , w_11599 , \3634_b0 );
buf ( \3636_b1 , \2120_b1 );
not ( \3636_b1 , w_11600 );
not ( \3636_b0 , w_11601 );
and ( w_11600 , w_11601 , \2120_b0 );
or ( \3637_b1 , \3635_b1 , w_11602 );
or ( \3637_b0 , \3635_b0 , \3636_b0 );
not ( \3636_b0 , w_11603 );
and ( w_11603 , w_11602 , \3636_b1 );
or ( \3638_b1 , \2120_b1 , w_11604 );
or ( \3638_b0 , \2120_b0 , \3634_b0 );
not ( \3634_b0 , w_11605 );
and ( w_11605 , w_11604 , \3634_b1 );
or ( \3639_b1 , \3637_b1 , w_11607 );
not ( w_11607 , w_11608 );
and ( \3639_b0 , \3637_b0 , w_11609 );
and ( w_11608 ,  , w_11609 );
buf ( w_11607 , \3638_b1 );
not ( w_11607 , w_11610 );
not (  , w_11611 );
and ( w_11610 , w_11611 , \3638_b0 );
or ( \3640_b1 , \3639_b1 , w_11613 );
not ( w_11613 , w_11614 );
and ( \3640_b0 , \3639_b0 , w_11615 );
and ( w_11614 ,  , w_11615 );
buf ( w_11613 , \1478_b1 );
not ( w_11613 , w_11616 );
not (  , w_11617 );
and ( w_11616 , w_11617 , \1478_b0 );
or ( \3641_b1 , \3632_b1 , w_11619 );
not ( w_11619 , w_11620 );
and ( \3641_b0 , \3632_b0 , w_11621 );
and ( w_11620 ,  , w_11621 );
buf ( w_11619 , \3640_b1 );
not ( w_11619 , w_11622 );
not (  , w_11623 );
and ( w_11622 , w_11623 , \3640_b0 );
or ( \3642_b1 , \c[8]_b1 , \d[8]_b1 );
xor ( \3642_b0 , \c[8]_b0 , w_11624 );
not ( w_11624 , w_11625 );
and ( w_11625 , \d[8]_b1 , \d[8]_b0 );
buf ( \3643_b1 , \3642_b1 );
not ( \3643_b1 , w_11626 );
not ( \3643_b0 , w_11627 );
and ( w_11626 , w_11627 , \3642_b0 );
buf ( \3644_b1 , \1320_b1 );
not ( \3644_b1 , w_11628 );
not ( \3644_b0 , w_11629 );
and ( w_11628 , w_11629 , \1320_b0 );
or ( \3645_b1 , \3643_b1 , w_11630 );
or ( \3645_b0 , \3643_b0 , \3644_b0 );
not ( \3644_b0 , w_11631 );
and ( w_11631 , w_11630 , \3644_b1 );
buf ( \3646_b1 , \2989_b1 );
not ( \3646_b1 , w_11632 );
not ( \3646_b0 , w_11633 );
and ( w_11632 , w_11633 , \2989_b0 );
or ( \3647_b1 , \3646_b1 , w_11635 );
not ( w_11635 , w_11636 );
and ( \3647_b0 , \3646_b0 , w_11637 );
and ( w_11636 ,  , w_11637 );
buf ( w_11635 , \2994_b1 );
not ( w_11635 , w_11638 );
not (  , w_11639 );
and ( w_11638 , w_11639 , \2994_b0 );
buf ( \3648_b1 , \3647_b1 );
not ( \3648_b1 , w_11640 );
not ( \3648_b0 , w_11641 );
and ( w_11640 , w_11641 , \3647_b0 );
buf ( \3649_b1 , \2979_b1 );
not ( \3649_b1 , w_11642 );
not ( \3649_b0 , w_11643 );
and ( w_11642 , w_11643 , \2979_b0 );
or ( \3650_b1 , \3648_b1 , w_11644 );
or ( \3650_b0 , \3648_b0 , \3649_b0 );
not ( \3649_b0 , w_11645 );
and ( w_11645 , w_11644 , \3649_b1 );
or ( \3651_b1 , \2979_b1 , w_11646 );
or ( \3651_b0 , \2979_b0 , \3647_b0 );
not ( \3647_b0 , w_11647 );
and ( w_11647 , w_11646 , \3647_b1 );
or ( \3652_b1 , \3650_b1 , w_11649 );
not ( w_11649 , w_11650 );
and ( \3652_b0 , \3650_b0 , w_11651 );
and ( w_11650 ,  , w_11651 );
buf ( w_11649 , \3651_b1 );
not ( w_11649 , w_11652 );
not (  , w_11653 );
and ( w_11652 , w_11653 , \3651_b0 );
or ( \3653_b1 , \2961_b1 , \3652_b1 );
not ( \3652_b1 , w_11654 );
and ( \3653_b0 , \2961_b0 , w_11655 );
and ( w_11654 , w_11655 , \3652_b0 );
buf ( \3654_b1 , \3051_b1 );
not ( \3654_b1 , w_11656 );
not ( \3654_b0 , w_11657 );
and ( w_11656 , w_11657 , \3051_b0 );
or ( \3655_b1 , \3654_b1 , w_11659 );
not ( w_11659 , w_11660 );
and ( \3655_b0 , \3654_b0 , w_11661 );
and ( w_11660 ,  , w_11661 );
buf ( w_11659 , \3056_b1 );
not ( w_11659 , w_11662 );
not (  , w_11663 );
and ( w_11662 , w_11663 , \3056_b0 );
buf ( \3656_b1 , \3655_b1 );
not ( \3656_b1 , w_11664 );
not ( \3656_b0 , w_11665 );
and ( w_11664 , w_11665 , \3655_b0 );
buf ( \3657_b1 , \3041_b1 );
not ( \3657_b1 , w_11666 );
not ( \3657_b0 , w_11667 );
and ( w_11666 , w_11667 , \3041_b0 );
or ( \3658_b1 , \3656_b1 , w_11668 );
or ( \3658_b0 , \3656_b0 , \3657_b0 );
not ( \3657_b0 , w_11669 );
and ( w_11669 , w_11668 , \3657_b1 );
or ( \3659_b1 , \3041_b1 , w_11670 );
or ( \3659_b0 , \3041_b0 , \3655_b0 );
not ( \3655_b0 , w_11671 );
and ( w_11671 , w_11670 , \3655_b1 );
or ( \3660_b1 , \3658_b1 , w_11673 );
not ( w_11673 , w_11674 );
and ( \3660_b0 , \3658_b0 , w_11675 );
and ( w_11674 ,  , w_11675 );
buf ( w_11673 , \3659_b1 );
not ( w_11673 , w_11676 );
not (  , w_11677 );
and ( w_11676 , w_11677 , \3659_b0 );
buf ( \3661_b1 , \3660_b1 );
not ( \3661_b1 , w_11678 );
not ( \3661_b0 , w_11679 );
and ( w_11678 , w_11679 , \3660_b0 );
buf ( \3662_b1 , \3087_b1 );
not ( \3662_b1 , w_11680 );
not ( \3662_b0 , w_11681 );
and ( w_11680 , w_11681 , \3087_b0 );
or ( \3663_b1 , \3661_b1 , w_11682 );
or ( \3663_b0 , \3661_b0 , \3662_b0 );
not ( \3662_b0 , w_11683 );
and ( w_11683 , w_11682 , \3662_b1 );
or ( \3664_b1 , \1282_b1 , \d[8]_b1 );
not ( \d[8]_b1 , w_11684 );
and ( \3664_b0 , \1282_b0 , w_11685 );
and ( w_11684 , w_11685 , \d[8]_b0 );
or ( \3665_b1 , \c[8]_b1 , \1514_b1 );
not ( \1514_b1 , w_11686 );
and ( \3665_b0 , \c[8]_b0 , w_11687 );
and ( w_11686 , w_11687 , \1514_b0 );
or ( \3666_b1 , \1293_b1 , \b[8]_b1 );
not ( \b[8]_b1 , w_11688 );
and ( \3666_b0 , \1293_b0 , w_11689 );
and ( w_11688 , w_11689 , \b[8]_b0 );
or ( \3668_b1 , \3663_b1 , w_11691 );
not ( w_11691 , w_11692 );
and ( \3668_b0 , \3663_b0 , w_11693 );
and ( w_11692 ,  , w_11693 );
buf ( w_11691 , \3667_b1 );
not ( w_11691 , w_11694 );
not (  , w_11695 );
and ( w_11694 , w_11695 , \3667_b0 );
or ( \3669_b1 , \3653_b1 , w_11697 );
not ( w_11697 , w_11698 );
and ( \3669_b0 , \3653_b0 , w_11699 );
and ( w_11698 ,  , w_11699 );
buf ( w_11697 , \3668_b1 );
not ( w_11697 , w_11700 );
not (  , w_11701 );
and ( w_11700 , w_11701 , \3668_b0 );
or ( \3670_b1 , \3645_b1 , w_11703 );
not ( w_11703 , w_11704 );
and ( \3670_b0 , \3645_b0 , w_11705 );
and ( w_11704 ,  , w_11705 );
buf ( w_11703 , \3669_b1 );
not ( w_11703 , w_11706 );
not (  , w_11707 );
and ( w_11706 , w_11707 , \3669_b0 );
or ( \3671_b1 , \3641_b1 , w_11709 );
not ( w_11709 , w_11710 );
and ( \3671_b0 , \3641_b0 , w_11711 );
and ( w_11710 ,  , w_11711 );
buf ( w_11709 , \3670_b1 );
not ( w_11709 , w_11712 );
not (  , w_11713 );
and ( w_11712 , w_11713 , \3670_b0 );
or ( \3672_b1 , \a[8]_b1 , w_11714 );
or ( \3672_b0 , \a[8]_b0 , \b[8]_b0 );
not ( \b[8]_b0 , w_11715 );
and ( w_11715 , w_11714 , \b[8]_b1 );
or ( \3673_b1 , \3672_b1 , w_11717 );
not ( w_11717 , w_11718 );
and ( \3673_b0 , \3672_b0 , w_11719 );
and ( w_11718 ,  , w_11719 );
buf ( w_11717 , \1351_b1 );
not ( w_11717 , w_11720 );
not (  , w_11721 );
and ( w_11720 , w_11721 , \1351_b0 );
or ( \3674_b1 , \b[8]_b1 , \c[8]_b1 );
not ( \c[8]_b1 , w_11722 );
and ( \3674_b0 , \b[8]_b0 , w_11723 );
and ( w_11722 , w_11723 , \c[8]_b0 );
or ( \3675_b1 , \1316_b1 , w_11725 );
not ( w_11725 , w_11726 );
and ( \3675_b0 , \1316_b0 , w_11727 );
and ( w_11726 ,  , w_11727 );
buf ( w_11725 , \3674_b1 );
not ( w_11725 , w_11728 );
not (  , w_11729 );
and ( w_11728 , w_11729 , \3674_b0 );
or ( \3677_b1 , \3622_b1 , w_11731 );
not ( w_11731 , w_11732 );
and ( \3677_b0 , \3622_b0 , w_11733 );
and ( w_11732 ,  , w_11733 );
buf ( w_11731 , \3676_b1 );
not ( w_11731 , w_11734 );
not (  , w_11735 );
and ( w_11734 , w_11735 , \3676_b0 );
or ( \3678_b1 , \3620_b1 , w_11737 );
not ( w_11737 , w_11738 );
and ( \3678_b0 , \3620_b0 , w_11739 );
and ( w_11738 ,  , w_11739 );
buf ( w_11737 , \3677_b1 );
not ( w_11737 , w_11740 );
not (  , w_11741 );
and ( w_11740 , w_11741 , \3677_b0 );
buf ( \3679_b1 , \a[9]_b1 );
not ( \3679_b1 , w_11742 );
not ( \3679_b0 , w_11743 );
and ( w_11742 , w_11743 , \a[9]_b0 );
buf ( \3680_b1 , \3114_b1 );
not ( \3680_b1 , w_11744 );
not ( \3680_b0 , w_11745 );
and ( w_11744 , w_11745 , \3114_b0 );
or ( \3681_b1 , \3679_b1 , w_11746 );
or ( \3681_b0 , \3679_b0 , \3680_b0 );
not ( \3680_b0 , w_11747 );
and ( w_11747 , w_11746 , \3680_b1 );
or ( \3682_b1 , \644_b1 , \d[9]_b1 );
not ( \d[9]_b1 , w_11748 );
and ( \3682_b0 , \644_b0 , w_11749 );
and ( w_11748 , w_11749 , \d[9]_b0 );
or ( \3683_b1 , \2906_b1 , w_11751 );
not ( w_11751 , w_11752 );
and ( \3683_b0 , \2906_b0 , w_11753 );
and ( w_11752 ,  , w_11753 );
buf ( w_11751 , \2892_b1 );
not ( w_11751 , w_11754 );
not (  , w_11755 );
and ( w_11754 , w_11755 , \2892_b0 );
buf ( \3684_b1 , \3683_b1 );
not ( \3684_b1 , w_11756 );
not ( \3684_b0 , w_11757 );
and ( w_11756 , w_11757 , \3683_b0 );
buf ( \3685_b1 , \2900_b1 );
not ( \3685_b1 , w_11758 );
not ( \3685_b0 , w_11759 );
and ( w_11758 , w_11759 , \2900_b0 );
buf ( \3686_b1 , \3626_b1 );
not ( \3686_b1 , w_11760 );
not ( \3686_b0 , w_11761 );
and ( w_11760 , w_11761 , \3626_b0 );
or ( \3687_b1 , \3685_b1 , w_11762 );
or ( \3687_b0 , \3685_b0 , \3686_b0 );
not ( \3686_b0 , w_11763 );
and ( w_11763 , w_11762 , \3686_b1 );
buf ( \3688_b1 , \2903_b1 );
not ( \3688_b1 , w_11764 );
not ( \3688_b0 , w_11765 );
and ( w_11764 , w_11765 , \2903_b0 );
or ( \3689_b1 , \3687_b1 , w_11767 );
not ( w_11767 , w_11768 );
and ( \3689_b0 , \3687_b0 , w_11769 );
and ( w_11768 ,  , w_11769 );
buf ( w_11767 , \3688_b1 );
not ( w_11767 , w_11770 );
not (  , w_11771 );
and ( w_11770 , w_11771 , \3688_b0 );
buf ( \3690_b1 , \3689_b1 );
not ( \3690_b1 , w_11772 );
not ( \3690_b0 , w_11773 );
and ( w_11772 , w_11773 , \3689_b0 );
or ( \3691_b1 , \3684_b1 , w_11774 );
or ( \3691_b0 , \3684_b0 , \3690_b0 );
not ( \3690_b0 , w_11775 );
and ( w_11775 , w_11774 , \3690_b1 );
or ( \3692_b1 , \3689_b1 , w_11776 );
or ( \3692_b0 , \3689_b0 , \3683_b0 );
not ( \3683_b0 , w_11777 );
and ( w_11777 , w_11776 , \3683_b1 );
or ( \3693_b1 , \3691_b1 , w_11779 );
not ( w_11779 , w_11780 );
and ( \3693_b0 , \3691_b0 , w_11781 );
and ( w_11780 ,  , w_11781 );
buf ( w_11779 , \3692_b1 );
not ( w_11779 , w_11782 );
not (  , w_11783 );
and ( w_11782 , w_11783 , \3692_b0 );
or ( \3694_b1 , \3693_b1 , \2936_b1 );
not ( \2936_b1 , w_11784 );
and ( \3694_b0 , \3693_b0 , w_11785 );
and ( w_11784 , w_11785 , \2936_b0 );
buf ( \3695_b1 , \2165_b1 );
not ( \3695_b1 , w_11786 );
not ( \3695_b0 , w_11787 );
and ( w_11786 , w_11787 , \2165_b0 );
or ( \3696_b1 , \3695_b1 , w_11789 );
not ( w_11789 , w_11790 );
and ( \3696_b0 , \3695_b0 , w_11791 );
and ( w_11790 ,  , w_11791 );
buf ( w_11789 , \2190_b1 );
not ( w_11789 , w_11792 );
not (  , w_11793 );
and ( w_11792 , w_11793 , \2190_b0 );
buf ( \3697_b1 , \3696_b1 );
not ( \3697_b1 , w_11794 );
not ( \3697_b0 , w_11795 );
and ( w_11794 , w_11795 , \3696_b0 );
buf ( \3698_b1 , \2172_b1 );
not ( \3698_b1 , w_11796 );
not ( \3698_b0 , w_11797 );
and ( w_11796 , w_11797 , \2172_b0 );
buf ( \3699_b1 , \3698_b1 );
not ( \3699_b1 , w_11798 );
not ( \3699_b0 , w_11799 );
and ( w_11798 , w_11799 , \3698_b0 );
buf ( \3700_b1 , \2120_b1 );
not ( \3700_b1 , w_11800 );
not ( \3700_b0 , w_11801 );
and ( w_11800 , w_11801 , \2120_b0 );
or ( \3701_b1 , \3699_b1 , w_11802 );
or ( \3701_b0 , \3699_b0 , \3700_b0 );
not ( \3700_b0 , w_11803 );
and ( w_11803 , w_11802 , \3700_b1 );
or ( \3702_b1 , \3701_b1 , w_11805 );
not ( w_11805 , w_11806 );
and ( \3702_b0 , \3701_b0 , w_11807 );
and ( w_11806 ,  , w_11807 );
buf ( w_11805 , \2188_b1 );
not ( w_11805 , w_11808 );
not (  , w_11809 );
and ( w_11808 , w_11809 , \2188_b0 );
buf ( \3703_b1 , \3702_b1 );
not ( \3703_b1 , w_11810 );
not ( \3703_b0 , w_11811 );
and ( w_11810 , w_11811 , \3702_b0 );
or ( \3704_b1 , \3697_b1 , w_11812 );
or ( \3704_b0 , \3697_b0 , \3703_b0 );
not ( \3703_b0 , w_11813 );
and ( w_11813 , w_11812 , \3703_b1 );
or ( \3705_b1 , \3702_b1 , w_11814 );
or ( \3705_b0 , \3702_b0 , \3696_b0 );
not ( \3696_b0 , w_11815 );
and ( w_11815 , w_11814 , \3696_b1 );
or ( \3706_b1 , \3704_b1 , w_11817 );
not ( w_11817 , w_11818 );
and ( \3706_b0 , \3704_b0 , w_11819 );
and ( w_11818 ,  , w_11819 );
buf ( w_11817 , \3705_b1 );
not ( w_11817 , w_11820 );
not (  , w_11821 );
and ( w_11820 , w_11821 , \3705_b0 );
or ( \3707_b1 , \3706_b1 , \1478_b1 );
not ( \1478_b1 , w_11822 );
and ( \3707_b0 , \3706_b0 , w_11823 );
and ( w_11822 , w_11823 , \1478_b0 );
or ( \3708_b1 , \3694_b1 , w_11825 );
not ( w_11825 , w_11826 );
and ( \3708_b0 , \3694_b0 , w_11827 );
and ( w_11826 ,  , w_11827 );
buf ( w_11825 , \3707_b1 );
not ( w_11825 , w_11828 );
not (  , w_11829 );
and ( w_11828 , w_11829 , \3707_b0 );
or ( \3709_b1 , \b[9]_b1 , \c[9]_b1 );
not ( \c[9]_b1 , w_11830 );
and ( \3709_b0 , \b[9]_b0 , w_11831 );
and ( w_11830 , w_11831 , \c[9]_b0 );
or ( \3710_b1 , \1316_b1 , w_11833 );
not ( w_11833 , w_11834 );
and ( \3710_b0 , \1316_b0 , w_11835 );
and ( w_11834 ,  , w_11835 );
buf ( w_11833 , \3709_b1 );
not ( w_11833 , w_11836 );
not (  , w_11837 );
and ( w_11836 , w_11837 , \3709_b0 );
or ( \3711_b1 , \a[9]_b1 , w_11838 );
or ( \3711_b0 , \a[9]_b0 , \b[9]_b0 );
not ( \b[9]_b0 , w_11839 );
and ( w_11839 , w_11838 , \b[9]_b1 );
or ( \3712_b1 , \672_b1 , \3711_b1 );
not ( \3711_b1 , w_11840 );
and ( \3712_b0 , \672_b0 , w_11841 );
and ( w_11840 , w_11841 , \3711_b0 );
or ( \3713_b1 , \c[9]_b1 , \d[9]_b1 );
xor ( \3713_b0 , \c[9]_b0 , w_11842 );
not ( w_11842 , w_11843 );
and ( w_11843 , \d[9]_b1 , \d[9]_b0 );
buf ( \3714_b1 , \3713_b1 );
not ( \3714_b1 , w_11844 );
not ( \3714_b0 , w_11845 );
and ( w_11844 , w_11845 , \3713_b0 );
buf ( \3715_b1 , \925_b1 );
not ( \3715_b1 , w_11846 );
not ( \3715_b0 , w_11847 );
and ( w_11846 , w_11847 , \925_b0 );
or ( \3716_b1 , \3714_b1 , w_11848 );
or ( \3716_b0 , \3714_b0 , \3715_b0 );
not ( \3715_b0 , w_11849 );
and ( w_11849 , w_11848 , \3715_b1 );
buf ( \3717_b1 , \3646_b1 );
not ( \3717_b1 , w_11850 );
not ( \3717_b0 , w_11851 );
and ( w_11850 , w_11851 , \3646_b0 );
buf ( \3718_b1 , \2979_b1 );
not ( \3718_b1 , w_11852 );
not ( \3718_b0 , w_11853 );
and ( w_11852 , w_11853 , \2979_b0 );
or ( \3719_b1 , \3717_b1 , w_11854 );
or ( \3719_b0 , \3717_b0 , \3718_b0 );
not ( \3718_b0 , w_11855 );
and ( w_11855 , w_11854 , \3718_b1 );
or ( \3720_b1 , \3719_b1 , w_11857 );
not ( w_11857 , w_11858 );
and ( \3720_b0 , \3719_b0 , w_11859 );
and ( w_11858 ,  , w_11859 );
buf ( w_11857 , \2994_b1 );
not ( w_11857 , w_11860 );
not (  , w_11861 );
and ( w_11860 , w_11861 , \2994_b0 );
buf ( \3721_b1 , \2990_b1 );
not ( \3721_b1 , w_11862 );
not ( \3721_b0 , w_11863 );
and ( w_11862 , w_11863 , \2990_b0 );
or ( \3722_b1 , \3721_b1 , w_11865 );
not ( w_11865 , w_11866 );
and ( \3722_b0 , \3721_b0 , w_11867 );
and ( w_11866 ,  , w_11867 );
buf ( w_11865 , \2996_b1 );
not ( w_11865 , w_11868 );
not (  , w_11869 );
and ( w_11868 , w_11869 , \2996_b0 );
or ( \3723_b1 , \3720_b1 , w_11870 );
xor ( \3723_b0 , \3720_b0 , w_11872 );
not ( w_11872 , w_11873 );
and ( w_11873 , w_11870 , w_11871 );
buf ( w_11870 , \3722_b1 );
not ( w_11870 , w_11874 );
not ( w_11871 , w_11875 );
and ( w_11874 , w_11875 , \3722_b0 );
or ( \3724_b1 , \2961_b1 , \3723_b1 );
not ( \3723_b1 , w_11876 );
and ( \3724_b0 , \2961_b0 , w_11877 );
and ( w_11876 , w_11877 , \3723_b0 );
buf ( \3725_b1 , \3654_b1 );
not ( \3725_b1 , w_11878 );
not ( \3725_b0 , w_11879 );
and ( w_11878 , w_11879 , \3654_b0 );
buf ( \3726_b1 , \3041_b1 );
not ( \3726_b1 , w_11880 );
not ( \3726_b0 , w_11881 );
and ( w_11880 , w_11881 , \3041_b0 );
or ( \3727_b1 , \3725_b1 , w_11882 );
or ( \3727_b0 , \3725_b0 , \3726_b0 );
not ( \3726_b0 , w_11883 );
and ( w_11883 , w_11882 , \3726_b1 );
or ( \3728_b1 , \3727_b1 , w_11885 );
not ( w_11885 , w_11886 );
and ( \3728_b0 , \3727_b0 , w_11887 );
and ( w_11886 ,  , w_11887 );
buf ( w_11885 , \3056_b1 );
not ( w_11885 , w_11888 );
not (  , w_11889 );
and ( w_11888 , w_11889 , \3056_b0 );
buf ( \3729_b1 , \3052_b1 );
not ( \3729_b1 , w_11890 );
not ( \3729_b0 , w_11891 );
and ( w_11890 , w_11891 , \3052_b0 );
or ( \3730_b1 , \3729_b1 , w_11893 );
not ( w_11893 , w_11894 );
and ( \3730_b0 , \3729_b0 , w_11895 );
and ( w_11894 ,  , w_11895 );
buf ( w_11893 , \3058_b1 );
not ( w_11893 , w_11896 );
not (  , w_11897 );
and ( w_11896 , w_11897 , \3058_b0 );
or ( \3731_b1 , \3728_b1 , w_11898 );
xor ( \3731_b0 , \3728_b0 , w_11900 );
not ( w_11900 , w_11901 );
and ( w_11901 , w_11898 , w_11899 );
buf ( w_11898 , \3730_b1 );
not ( w_11898 , w_11902 );
not ( w_11899 , w_11903 );
and ( w_11902 , w_11903 , \3730_b0 );
buf ( \3732_b1 , \3731_b1 );
not ( \3732_b1 , w_11904 );
not ( \3732_b0 , w_11905 );
and ( w_11904 , w_11905 , \3731_b0 );
buf ( \3733_b1 , \3087_b1 );
not ( \3733_b1 , w_11906 );
not ( \3733_b0 , w_11907 );
and ( w_11906 , w_11907 , \3087_b0 );
or ( \3734_b1 , \3732_b1 , w_11908 );
or ( \3734_b0 , \3732_b0 , \3733_b0 );
not ( \3733_b0 , w_11909 );
and ( w_11909 , w_11908 , \3733_b1 );
or ( \3735_b1 , \1282_b1 , \d[9]_b1 );
not ( \d[9]_b1 , w_11910 );
and ( \3735_b0 , \1282_b0 , w_11911 );
and ( w_11910 , w_11911 , \d[9]_b0 );
or ( \3736_b1 , \c[9]_b1 , \1435_b1 );
not ( \1435_b1 , w_11912 );
and ( \3736_b0 , \c[9]_b0 , w_11913 );
and ( w_11912 , w_11913 , \1435_b0 );
or ( \3737_b1 , \1293_b1 , \b[9]_b1 );
not ( \b[9]_b1 , w_11914 );
and ( \3737_b0 , \1293_b0 , w_11915 );
and ( w_11914 , w_11915 , \b[9]_b0 );
or ( \3739_b1 , \3734_b1 , w_11917 );
not ( w_11917 , w_11918 );
and ( \3739_b0 , \3734_b0 , w_11919 );
and ( w_11918 ,  , w_11919 );
buf ( w_11917 , \3738_b1 );
not ( w_11917 , w_11920 );
not (  , w_11921 );
and ( w_11920 , w_11921 , \3738_b0 );
or ( \3740_b1 , \3724_b1 , w_11923 );
not ( w_11923 , w_11924 );
and ( \3740_b0 , \3724_b0 , w_11925 );
and ( w_11924 ,  , w_11925 );
buf ( w_11923 , \3739_b1 );
not ( w_11923 , w_11926 );
not (  , w_11927 );
and ( w_11926 , w_11927 , \3739_b0 );
or ( \3741_b1 , \3716_b1 , w_11929 );
not ( w_11929 , w_11930 );
and ( \3741_b0 , \3716_b0 , w_11931 );
and ( w_11930 ,  , w_11931 );
buf ( w_11929 , \3740_b1 );
not ( w_11929 , w_11932 );
not (  , w_11933 );
and ( w_11932 , w_11933 , \3740_b0 );
or ( \3742_b1 , \3712_b1 , w_11935 );
not ( w_11935 , w_11936 );
and ( \3742_b0 , \3712_b0 , w_11937 );
and ( w_11936 ,  , w_11937 );
buf ( w_11935 , \3741_b1 );
not ( w_11935 , w_11938 );
not (  , w_11939 );
and ( w_11938 , w_11939 , \3741_b0 );
or ( \3744_b1 , \3682_b1 , w_11941 );
not ( w_11941 , w_11942 );
and ( \3744_b0 , \3682_b0 , w_11943 );
and ( w_11942 ,  , w_11943 );
buf ( w_11941 , \3743_b1 );
not ( w_11941 , w_11944 );
not (  , w_11945 );
and ( w_11944 , w_11945 , \3743_b0 );
or ( \3745_b1 , \3681_b1 , w_11947 );
not ( w_11947 , w_11948 );
and ( \3745_b0 , \3681_b0 , w_11949 );
and ( w_11948 ,  , w_11949 );
buf ( w_11947 , \3744_b1 );
not ( w_11947 , w_11950 );
not (  , w_11951 );
and ( w_11950 , w_11951 , \3744_b0 );
buf ( \3746_b1 , \2866_b1 );
not ( \3746_b1 , w_11952 );
not ( \3746_b0 , w_11953 );
and ( w_11952 , w_11953 , \2866_b0 );
buf ( \3747_b1 , \2910_b1 );
not ( \3747_b1 , w_11954 );
not ( \3747_b0 , w_11955 );
and ( w_11954 , w_11955 , \2910_b0 );
or ( \3748_b1 , \3746_b1 , w_11956 );
or ( \3748_b0 , \3746_b0 , \3747_b0 );
not ( \3747_b0 , w_11957 );
and ( w_11957 , w_11956 , \3747_b1 );
buf ( \3749_b1 , \2914_b1 );
not ( \3749_b1 , w_11958 );
not ( \3749_b0 , w_11959 );
and ( w_11958 , w_11959 , \2914_b0 );
or ( \3750_b1 , \3748_b1 , w_11961 );
not ( w_11961 , w_11962 );
and ( \3750_b0 , \3748_b0 , w_11963 );
and ( w_11962 ,  , w_11963 );
buf ( w_11961 , \3749_b1 );
not ( w_11961 , w_11964 );
not (  , w_11965 );
and ( w_11964 , w_11965 , \3749_b0 );
or ( \3751_b1 , \3750_b1 , w_11967 );
not ( w_11967 , w_11968 );
and ( \3751_b0 , \3750_b0 , w_11969 );
and ( w_11968 ,  , w_11969 );
buf ( w_11967 , \2814_b1 );
not ( w_11967 , w_11970 );
not (  , w_11971 );
and ( w_11970 , w_11971 , \2814_b0 );
or ( \3752_b1 , \2926_b1 , w_11973 );
not ( w_11973 , w_11974 );
and ( \3752_b0 , \2926_b0 , w_11975 );
and ( w_11974 ,  , w_11975 );
buf ( w_11973 , \2913_b1 );
not ( w_11973 , w_11976 );
not (  , w_11977 );
and ( w_11976 , w_11977 , \2913_b0 );
or ( \3753_b1 , \3751_b1 , \3752_b1 );
xor ( \3753_b0 , \3751_b0 , w_11978 );
not ( w_11978 , w_11979 );
and ( w_11979 , \3752_b1 , \3752_b0 );
or ( \3754_b1 , \3753_b1 , \2936_b1 );
not ( \2936_b1 , w_11980 );
and ( \3754_b0 , \3753_b0 , w_11981 );
and ( w_11980 , w_11981 , \2936_b0 );
buf ( \3755_b1 , \2206_b1 );
not ( \3755_b1 , w_11982 );
not ( \3755_b0 , w_11983 );
and ( w_11982 , w_11983 , \2206_b0 );
buf ( \3756_b1 , \2193_b1 );
not ( \3756_b1 , w_11984 );
not ( \3756_b0 , w_11985 );
and ( w_11984 , w_11985 , \2193_b0 );
or ( \3757_b1 , \3755_b1 , w_11986 );
or ( \3757_b0 , \3755_b0 , \3756_b0 );
not ( \3756_b0 , w_11987 );
and ( w_11987 , w_11986 , \3756_b1 );
buf ( \3758_b1 , \2211_b1 );
not ( \3758_b1 , w_11988 );
not ( \3758_b0 , w_11989 );
and ( w_11988 , w_11989 , \2211_b0 );
or ( \3759_b1 , \3757_b1 , w_11991 );
not ( w_11991 , w_11992 );
and ( \3759_b0 , \3757_b0 , w_11993 );
and ( w_11992 ,  , w_11993 );
buf ( w_11991 , \3758_b1 );
not ( w_11991 , w_11994 );
not (  , w_11995 );
and ( w_11994 , w_11995 , \3758_b0 );
or ( \3760_b1 , \3759_b1 , w_11997 );
not ( w_11997 , w_11998 );
and ( \3760_b0 , \3759_b0 , w_11999 );
and ( w_11998 ,  , w_11999 );
buf ( w_11997 , \2112_b1 );
not ( w_11997 , w_12000 );
not (  , w_12001 );
and ( w_12000 , w_12001 , \2112_b0 );
buf ( \3761_b1 , \2221_b1 );
not ( \3761_b1 , w_12002 );
not ( \3761_b0 , w_12003 );
and ( w_12002 , w_12003 , \2221_b0 );
or ( \3762_b1 , \3761_b1 , w_12005 );
not ( w_12005 , w_12006 );
and ( \3762_b0 , \3761_b0 , w_12007 );
and ( w_12006 ,  , w_12007 );
buf ( w_12005 , \2205_b1 );
not ( w_12005 , w_12008 );
not (  , w_12009 );
and ( w_12008 , w_12009 , \2205_b0 );
or ( \3763_b1 , \3760_b1 , \3762_b1 );
not ( \3762_b1 , w_12010 );
and ( \3763_b0 , \3760_b0 , w_12011 );
and ( w_12010 , w_12011 , \3762_b0 );
buf ( \3764_b1 , \3760_b1 );
not ( \3764_b1 , w_12012 );
not ( \3764_b0 , w_12013 );
and ( w_12012 , w_12013 , \3760_b0 );
buf ( \3765_b1 , \3762_b1 );
not ( \3765_b1 , w_12014 );
not ( \3765_b0 , w_12015 );
and ( w_12014 , w_12015 , \3762_b0 );
or ( \3766_b1 , \3764_b1 , \3765_b1 );
not ( \3765_b1 , w_12016 );
and ( \3766_b0 , \3764_b0 , w_12017 );
and ( w_12016 , w_12017 , \3765_b0 );
or ( \3767_b1 , \3763_b1 , w_12019 );
not ( w_12019 , w_12020 );
and ( \3767_b0 , \3763_b0 , w_12021 );
and ( w_12020 ,  , w_12021 );
buf ( w_12019 , \3766_b1 );
not ( w_12019 , w_12022 );
not (  , w_12023 );
and ( w_12022 , w_12023 , \3766_b0 );
or ( \3768_b1 , \3767_b1 , \1529_b1 );
not ( \1529_b1 , w_12024 );
and ( \3768_b0 , \3767_b0 , w_12025 );
and ( w_12024 , w_12025 , \1529_b0 );
or ( \3769_b1 , \3754_b1 , w_12027 );
not ( w_12027 , w_12028 );
and ( \3769_b0 , \3754_b0 , w_12029 );
and ( w_12028 ,  , w_12029 );
buf ( w_12027 , \3768_b1 );
not ( w_12027 , w_12030 );
not (  , w_12031 );
and ( w_12030 , w_12031 , \3768_b0 );
or ( \3770_b1 , \2946_b1 , w_12033 );
not ( w_12033 , w_12034 );
and ( \3770_b0 , \2946_b0 , w_12035 );
and ( w_12034 ,  , w_12035 );
buf ( w_12033 , \a[12]_b1 );
not ( w_12033 , w_12036 );
not (  , w_12037 );
and ( w_12036 , w_12037 , \a[12]_b0 );
buf ( \3771_b1 , \d[12]_b1 );
not ( \3771_b1 , w_12038 );
not ( \3771_b0 , w_12039 );
and ( w_12038 , w_12039 , \d[12]_b0 );
buf ( \3772_b1 , \1457_b1 );
not ( \3772_b1 , w_12040 );
not ( \3772_b0 , w_12041 );
and ( w_12040 , w_12041 , \1457_b0 );
or ( \3773_b1 , \3771_b1 , w_12042 );
or ( \3773_b0 , \3771_b0 , \3772_b0 );
not ( \3772_b0 , w_12043 );
and ( w_12043 , w_12042 , \3772_b1 );
or ( \3774_b1 , \b[12]_b1 , \c[12]_b1 );
not ( \c[12]_b1 , w_12044 );
and ( \3774_b0 , \b[12]_b0 , w_12045 );
and ( w_12044 , w_12045 , \c[12]_b0 );
or ( \3775_b1 , \1316_b1 , w_12047 );
not ( w_12047 , w_12048 );
and ( \3775_b0 , \1316_b0 , w_12049 );
and ( w_12048 ,  , w_12049 );
buf ( w_12047 , \3774_b1 );
not ( w_12047 , w_12050 );
not (  , w_12051 );
and ( w_12050 , w_12051 , \3774_b0 );
or ( \3776_b1 , \3773_b1 , w_12053 );
not ( w_12053 , w_12054 );
and ( \3776_b0 , \3773_b0 , w_12055 );
and ( w_12054 ,  , w_12055 );
buf ( w_12053 , \3775_b1 );
not ( w_12053 , w_12056 );
not (  , w_12057 );
and ( w_12056 , w_12057 , \3775_b0 );
buf ( \3777_b1 , \b[12]_b1 );
not ( \3777_b1 , w_12058 );
not ( \3777_b0 , w_12059 );
and ( w_12058 , w_12059 , \b[12]_b0 );
buf ( \3778_b1 , \3124_b1 );
not ( \3778_b1 , w_12060 );
not ( \3778_b0 , w_12061 );
and ( w_12060 , w_12061 , \3124_b0 );
or ( \3779_b1 , \3777_b1 , w_12062 );
or ( \3779_b0 , \3777_b0 , \3778_b0 );
not ( \3778_b0 , w_12063 );
and ( w_12063 , w_12062 , \3778_b1 );
or ( \3780_b1 , \1351_b1 , \a[12]_b1 );
not ( \a[12]_b1 , w_12064 );
and ( \3780_b0 , \1351_b0 , w_12065 );
and ( w_12064 , w_12065 , \a[12]_b0 );
or ( \3781_b1 , \c[12]_b1 , \d[12]_b1 );
xor ( \3781_b0 , \c[12]_b0 , w_12066 );
not ( w_12066 , w_12067 );
and ( w_12067 , \d[12]_b1 , \d[12]_b0 );
buf ( \3782_b1 , \3781_b1 );
not ( \3782_b1 , w_12068 );
not ( \3782_b0 , w_12069 );
and ( w_12068 , w_12069 , \3781_b0 );
buf ( \3783_b1 , \3305_b1 );
not ( \3783_b1 , w_12070 );
not ( \3783_b0 , w_12071 );
and ( w_12070 , w_12071 , \3305_b0 );
or ( \3784_b1 , \3782_b1 , w_12072 );
or ( \3784_b0 , \3782_b0 , \3783_b0 );
not ( \3783_b0 , w_12073 );
and ( w_12073 , w_12072 , \3783_b1 );
or ( \3785_b1 , \3533_b1 , w_12075 );
not ( w_12075 , w_12076 );
and ( \3785_b0 , \3533_b0 , w_12077 );
and ( w_12076 ,  , w_12077 );
buf ( w_12075 , \3010_b1 );
not ( w_12075 , w_12078 );
not (  , w_12079 );
and ( w_12078 , w_12079 , \3010_b0 );
buf ( \3786_b1 , \3785_b1 );
not ( \3786_b1 , w_12080 );
not ( \3786_b0 , w_12081 );
and ( w_12080 , w_12081 , \3785_b0 );
buf ( \3787_b1 , \2992_b1 );
not ( \3787_b1 , w_12082 );
not ( \3787_b0 , w_12083 );
and ( w_12082 , w_12083 , \2992_b0 );
buf ( \3788_b1 , \2979_b1 );
not ( \3788_b1 , w_12084 );
not ( \3788_b0 , w_12085 );
and ( w_12084 , w_12085 , \2979_b0 );
or ( \3789_b1 , \3787_b1 , w_12086 );
or ( \3789_b0 , \3787_b0 , \3788_b0 );
not ( \3788_b0 , w_12087 );
and ( w_12087 , w_12086 , \3788_b1 );
or ( \3790_b1 , \3789_b1 , w_12089 );
not ( w_12089 , w_12090 );
and ( \3790_b0 , \3789_b0 , w_12091 );
and ( w_12090 ,  , w_12091 );
buf ( w_12089 , \3008_b1 );
not ( w_12089 , w_12092 );
not (  , w_12093 );
and ( w_12092 , w_12093 , \3008_b0 );
buf ( \3791_b1 , \3790_b1 );
not ( \3791_b1 , w_12094 );
not ( \3791_b0 , w_12095 );
and ( w_12094 , w_12095 , \3790_b0 );
or ( \3792_b1 , \3786_b1 , w_12096 );
or ( \3792_b0 , \3786_b0 , \3791_b0 );
not ( \3791_b0 , w_12097 );
and ( w_12097 , w_12096 , \3791_b1 );
or ( \3793_b1 , \3790_b1 , w_12098 );
or ( \3793_b0 , \3790_b0 , \3785_b0 );
not ( \3785_b0 , w_12099 );
and ( w_12099 , w_12098 , \3785_b1 );
or ( \3794_b1 , \3792_b1 , w_12101 );
not ( w_12101 , w_12102 );
and ( \3794_b0 , \3792_b0 , w_12103 );
and ( w_12102 ,  , w_12103 );
buf ( w_12101 , \3793_b1 );
not ( w_12101 , w_12104 );
not (  , w_12105 );
and ( w_12104 , w_12105 , \3793_b0 );
or ( \3795_b1 , \3794_b1 , \2961_b1 );
not ( \2961_b1 , w_12106 );
and ( \3795_b0 , \3794_b0 , w_12107 );
and ( w_12106 , w_12107 , \2961_b0 );
or ( \3796_b1 , \3546_b1 , w_12109 );
not ( w_12109 , w_12110 );
and ( \3796_b0 , \3546_b0 , w_12111 );
and ( w_12110 ,  , w_12111 );
buf ( w_12109 , \3072_b1 );
not ( w_12109 , w_12112 );
not (  , w_12113 );
and ( w_12112 , w_12113 , \3072_b0 );
buf ( \3797_b1 , \3796_b1 );
not ( \3797_b1 , w_12114 );
not ( \3797_b0 , w_12115 );
and ( w_12114 , w_12115 , \3796_b0 );
buf ( \3798_b1 , \3054_b1 );
not ( \3798_b1 , w_12116 );
not ( \3798_b0 , w_12117 );
and ( w_12116 , w_12117 , \3054_b0 );
buf ( \3799_b1 , \3041_b1 );
not ( \3799_b1 , w_12118 );
not ( \3799_b0 , w_12119 );
and ( w_12118 , w_12119 , \3041_b0 );
or ( \3800_b1 , \3798_b1 , w_12120 );
or ( \3800_b0 , \3798_b0 , \3799_b0 );
not ( \3799_b0 , w_12121 );
and ( w_12121 , w_12120 , \3799_b1 );
or ( \3801_b1 , \3800_b1 , w_12123 );
not ( w_12123 , w_12124 );
and ( \3801_b0 , \3800_b0 , w_12125 );
and ( w_12124 ,  , w_12125 );
buf ( w_12123 , \3070_b1 );
not ( w_12123 , w_12126 );
not (  , w_12127 );
and ( w_12126 , w_12127 , \3070_b0 );
buf ( \3802_b1 , \3801_b1 );
not ( \3802_b1 , w_12128 );
not ( \3802_b0 , w_12129 );
and ( w_12128 , w_12129 , \3801_b0 );
or ( \3803_b1 , \3797_b1 , w_12130 );
or ( \3803_b0 , \3797_b0 , \3802_b0 );
not ( \3802_b0 , w_12131 );
and ( w_12131 , w_12130 , \3802_b1 );
or ( \3804_b1 , \3801_b1 , w_12132 );
or ( \3804_b0 , \3801_b0 , \3796_b0 );
not ( \3796_b0 , w_12133 );
and ( w_12133 , w_12132 , \3796_b1 );
or ( \3805_b1 , \3803_b1 , w_12135 );
not ( w_12135 , w_12136 );
and ( \3805_b0 , \3803_b0 , w_12137 );
and ( w_12136 ,  , w_12137 );
buf ( w_12135 , \3804_b1 );
not ( w_12135 , w_12138 );
not (  , w_12139 );
and ( w_12138 , w_12139 , \3804_b0 );
buf ( \3806_b1 , \3805_b1 );
not ( \3806_b1 , w_12140 );
not ( \3806_b0 , w_12141 );
and ( w_12140 , w_12141 , \3805_b0 );
buf ( \3807_b1 , \3087_b1 );
not ( \3807_b1 , w_12142 );
not ( \3807_b0 , w_12143 );
and ( w_12142 , w_12143 , \3087_b0 );
or ( \3808_b1 , \3806_b1 , w_12144 );
or ( \3808_b0 , \3806_b0 , \3807_b0 );
not ( \3807_b0 , w_12145 );
and ( w_12145 , w_12144 , \3807_b1 );
or ( \3809_b1 , \1282_b1 , \d[12]_b1 );
not ( \d[12]_b1 , w_12146 );
and ( \3809_b0 , \1282_b0 , w_12147 );
and ( w_12146 , w_12147 , \d[12]_b0 );
or ( \3810_b1 , \1435_b1 , \c[12]_b1 );
not ( \c[12]_b1 , w_12148 );
and ( \3810_b0 , \1435_b0 , w_12149 );
and ( w_12148 , w_12149 , \c[12]_b0 );
or ( \3811_b1 , \3809_b1 , w_12151 );
not ( w_12151 , w_12152 );
and ( \3811_b0 , \3809_b0 , w_12153 );
and ( w_12152 ,  , w_12153 );
buf ( w_12151 , \3810_b1 );
not ( w_12151 , w_12154 );
not (  , w_12155 );
and ( w_12154 , w_12155 , \3810_b0 );
or ( \3812_b1 , \3808_b1 , w_12157 );
not ( w_12157 , w_12158 );
and ( \3812_b0 , \3808_b0 , w_12159 );
and ( w_12158 ,  , w_12159 );
buf ( w_12157 , \3811_b1 );
not ( w_12157 , w_12160 );
not (  , w_12161 );
and ( w_12160 , w_12161 , \3811_b0 );
or ( \3813_b1 , \3795_b1 , w_12163 );
not ( w_12163 , w_12164 );
and ( \3813_b0 , \3795_b0 , w_12165 );
and ( w_12164 ,  , w_12165 );
buf ( w_12163 , \3812_b1 );
not ( w_12163 , w_12166 );
not (  , w_12167 );
and ( w_12166 , w_12167 , \3812_b0 );
or ( \3814_b1 , \3784_b1 , w_12169 );
not ( w_12169 , w_12170 );
and ( \3814_b0 , \3784_b0 , w_12171 );
and ( w_12170 ,  , w_12171 );
buf ( w_12169 , \3813_b1 );
not ( w_12169 , w_12172 );
not (  , w_12173 );
and ( w_12172 , w_12173 , \3813_b0 );
or ( \3815_b1 , \3780_b1 , w_12175 );
not ( w_12175 , w_12176 );
and ( \3815_b0 , \3780_b0 , w_12177 );
and ( w_12176 ,  , w_12177 );
buf ( w_12175 , \3814_b1 );
not ( w_12175 , w_12178 );
not (  , w_12179 );
and ( w_12178 , w_12179 , \3814_b0 );
or ( \3816_b1 , \3779_b1 , w_12181 );
not ( w_12181 , w_12182 );
and ( \3816_b0 , \3779_b0 , w_12183 );
and ( w_12182 ,  , w_12183 );
buf ( w_12181 , \3815_b1 );
not ( w_12181 , w_12184 );
not (  , w_12185 );
and ( w_12184 , w_12185 , \3815_b0 );
or ( \3817_b1 , \3776_b1 , w_12187 );
not ( w_12187 , w_12188 );
and ( \3817_b0 , \3776_b0 , w_12189 );
and ( w_12188 ,  , w_12189 );
buf ( w_12187 , \3816_b1 );
not ( w_12187 , w_12190 );
not (  , w_12191 );
and ( w_12190 , w_12191 , \3816_b0 );
buf ( \3819_b1 , \a[5]_b1 );
not ( \3819_b1 , w_12192 );
not ( \3819_b0 , w_12193 );
and ( w_12192 , w_12193 , \a[5]_b0 );
buf ( \3820_b1 , \1338_b1 );
not ( \3820_b1 , w_12194 );
not ( \3820_b0 , w_12195 );
and ( w_12194 , w_12195 , \1338_b0 );
or ( \3821_b1 , \3819_b1 , w_12196 );
or ( \3821_b0 , \3819_b0 , \3820_b0 );
not ( \3820_b0 , w_12197 );
and ( w_12197 , w_12196 , \3820_b1 );
or ( \3822_b1 , \a[5]_b1 , w_12198 );
or ( \3822_b0 , \a[5]_b0 , \d[5]_b0 );
not ( \d[5]_b0 , w_12199 );
and ( w_12199 , w_12198 , \d[5]_b1 );
buf ( \3823_b1 , \3822_b1 );
not ( \3823_b1 , w_12200 );
not ( \3823_b0 , w_12201 );
and ( w_12200 , w_12201 , \3822_b0 );
buf ( \3824_b1 , \644_b1 );
not ( \3824_b1 , w_12202 );
not ( \3824_b0 , w_12203 );
and ( w_12202 , w_12203 , \644_b0 );
or ( \3825_b1 , \3823_b1 , w_12204 );
or ( \3825_b0 , \3823_b0 , \3824_b0 );
not ( \3824_b0 , w_12205 );
and ( w_12205 , w_12204 , \3824_b1 );
buf ( \3826_b1 , \917_b1 );
not ( \3826_b1 , w_12206 );
not ( \3826_b0 , w_12207 );
and ( w_12206 , w_12207 , \917_b0 );
or ( \3827_b1 , \899_b1 , w_12209 );
not ( w_12209 , w_12210 );
and ( \3827_b0 , \899_b0 , w_12211 );
and ( w_12210 ,  , w_12211 );
buf ( w_12209 , \819_b1 );
not ( w_12209 , w_12212 );
not (  , w_12213 );
and ( w_12212 , w_12213 , \819_b0 );
or ( \3828_b1 , \3827_b1 , \879_b1 );
xor ( \3828_b0 , \3827_b0 , w_12214 );
not ( w_12214 , w_12215 );
and ( w_12215 , \879_b1 , \879_b0 );
buf ( \3829_b1 , \3828_b1 );
not ( \3829_b1 , w_12216 );
not ( \3829_b0 , w_12217 );
and ( w_12216 , w_12217 , \3828_b0 );
or ( \3830_b1 , \3826_b1 , \3829_b1 );
not ( \3829_b1 , w_12218 );
and ( \3830_b0 , \3826_b0 , w_12219 );
and ( w_12218 , w_12219 , \3829_b0 );
or ( \3831_b1 , \a[5]_b1 , w_12220 );
or ( \3831_b0 , \a[5]_b0 , \b[5]_b0 );
not ( \b[5]_b0 , w_12221 );
and ( w_12221 , w_12220 , \b[5]_b1 );
or ( \3832_b1 , \672_b1 , \3831_b1 );
not ( \3831_b1 , w_12222 );
and ( \3832_b0 , \672_b0 , w_12223 );
and ( w_12222 , w_12223 , \3831_b0 );
or ( \3833_b1 , \3830_b1 , w_12225 );
not ( w_12225 , w_12226 );
and ( \3833_b0 , \3830_b0 , w_12227 );
and ( w_12226 ,  , w_12227 );
buf ( w_12225 , \3832_b1 );
not ( w_12225 , w_12228 );
not (  , w_12229 );
and ( w_12228 , w_12229 , \3832_b0 );
or ( \3834_b1 , \3825_b1 , w_12231 );
not ( w_12231 , w_12232 );
and ( \3834_b0 , \3825_b0 , w_12233 );
and ( w_12232 ,  , w_12233 );
buf ( w_12231 , \3833_b1 );
not ( w_12231 , w_12234 );
not (  , w_12235 );
and ( w_12234 , w_12235 , \3833_b0 );
or ( \3835_b1 , \b[5]_b1 , \c[5]_b1 );
not ( \c[5]_b1 , w_12236 );
and ( \3835_b0 , \b[5]_b0 , w_12237 );
and ( w_12236 , w_12237 , \c[5]_b0 );
buf ( \3836_b1 , \3835_b1 );
not ( \3836_b1 , w_12238 );
not ( \3836_b0 , w_12239 );
and ( w_12238 , w_12239 , \3835_b0 );
buf ( \3837_b1 , \1316_b1 );
not ( \3837_b1 , w_12240 );
not ( \3837_b0 , w_12241 );
and ( w_12240 , w_12241 , \1316_b0 );
or ( \3838_b1 , \3836_b1 , w_12242 );
or ( \3838_b0 , \3836_b0 , \3837_b0 );
not ( \3837_b0 , w_12243 );
and ( w_12243 , w_12242 , \3837_b1 );
or ( \3839_b1 , \c[5]_b1 , \d[5]_b1 );
xor ( \3839_b0 , \c[5]_b0 , w_12244 );
not ( w_12244 , w_12245 );
and ( w_12245 , \d[5]_b1 , \d[5]_b0 );
or ( \3840_b1 , \3305_b1 , \3839_b1 );
not ( \3839_b1 , w_12246 );
and ( \3840_b0 , \3305_b0 , w_12247 );
and ( w_12246 , w_12247 , \3839_b0 );
buf ( \3841_b1 , \1089_b1 );
not ( \3841_b1 , w_12248 );
not ( \3841_b0 , w_12249 );
and ( w_12248 , w_12249 , \1089_b0 );
or ( \3842_b1 , \1095_b1 , w_12251 );
not ( w_12251 , w_12252 );
and ( \3842_b0 , \1095_b0 , w_12253 );
and ( w_12252 ,  , w_12253 );
buf ( w_12251 , \1027_b1 );
not ( w_12251 , w_12254 );
not (  , w_12255 );
and ( w_12254 , w_12255 , \1027_b0 );
buf ( \3843_b1 , \3842_b1 );
not ( \3843_b1 , w_12256 );
not ( \3843_b0 , w_12257 );
and ( w_12256 , w_12257 , \3842_b0 );
or ( \3844_b1 , \3841_b1 , w_12258 );
or ( \3844_b0 , \3841_b0 , \3843_b0 );
not ( \3843_b0 , w_12259 );
and ( w_12259 , w_12258 , \3843_b1 );
or ( \3845_b1 , \3842_b1 , w_12260 );
or ( \3845_b0 , \3842_b0 , \1089_b0 );
not ( \1089_b0 , w_12261 );
and ( w_12261 , w_12260 , \1089_b1 );
or ( \3846_b1 , \3844_b1 , w_12263 );
not ( w_12263 , w_12264 );
and ( \3846_b0 , \3844_b0 , w_12265 );
and ( w_12264 ,  , w_12265 );
buf ( w_12263 , \3845_b1 );
not ( w_12263 , w_12266 );
not (  , w_12267 );
and ( w_12266 , w_12267 , \3845_b0 );
buf ( \3847_b1 , \3846_b1 );
not ( \3847_b1 , w_12268 );
not ( \3847_b0 , w_12269 );
and ( w_12268 , w_12269 , \3846_b0 );
buf ( \3848_b1 , \1478_b1 );
not ( \3848_b1 , w_12270 );
not ( \3848_b0 , w_12271 );
and ( w_12270 , w_12271 , \1478_b0 );
or ( \3849_b1 , \3847_b1 , w_12272 );
or ( \3849_b0 , \3847_b0 , \3848_b0 );
not ( \3848_b0 , w_12273 );
and ( w_12273 , w_12272 , \3848_b1 );
or ( \3850_b1 , \1192_b1 , w_12275 );
not ( w_12275 , w_12276 );
and ( \3850_b0 , \1192_b0 , w_12277 );
and ( w_12276 ,  , w_12277 );
buf ( w_12275 , \1200_b1 );
not ( w_12275 , w_12278 );
not (  , w_12279 );
and ( w_12278 , w_12279 , \1200_b0 );
buf ( \3851_b1 , \3850_b1 );
not ( \3851_b1 , w_12280 );
not ( \3851_b0 , w_12281 );
and ( w_12280 , w_12281 , \3850_b0 );
or ( \3852_b1 , \1416_b1 , w_12282 );
or ( \3852_b0 , \1416_b0 , \1190_b0 );
not ( \1190_b0 , w_12283 );
and ( w_12283 , w_12282 , \1190_b1 );
or ( \3853_b1 , \3852_b1 , w_12285 );
not ( w_12285 , w_12286 );
and ( \3853_b0 , \3852_b0 , w_12287 );
and ( w_12286 ,  , w_12287 );
buf ( w_12285 , \1197_b1 );
not ( w_12285 , w_12288 );
not (  , w_12289 );
and ( w_12288 , w_12289 , \1197_b0 );
buf ( \3854_b1 , \3853_b1 );
not ( \3854_b1 , w_12290 );
not ( \3854_b0 , w_12291 );
and ( w_12290 , w_12291 , \3853_b0 );
or ( \3855_b1 , \3851_b1 , w_12292 );
or ( \3855_b0 , \3851_b0 , \3854_b0 );
not ( \3854_b0 , w_12293 );
and ( w_12293 , w_12292 , \3854_b1 );
or ( \3856_b1 , \3853_b1 , w_12294 );
or ( \3856_b0 , \3853_b0 , \3850_b0 );
not ( \3850_b0 , w_12295 );
and ( w_12295 , w_12294 , \3850_b1 );
or ( \3857_b1 , \3855_b1 , w_12297 );
not ( w_12297 , w_12298 );
and ( \3857_b0 , \3855_b0 , w_12299 );
and ( w_12298 ,  , w_12299 );
buf ( w_12297 , \3856_b1 );
not ( w_12297 , w_12300 );
not (  , w_12301 );
and ( w_12300 , w_12301 , \3856_b0 );
or ( \3858_b1 , \2961_b1 , \3857_b1 );
not ( \3857_b1 , w_12302 );
and ( \3858_b0 , \2961_b0 , w_12303 );
and ( w_12302 , w_12303 , \3857_b0 );
or ( \3859_b1 , \1255_b1 , w_12305 );
not ( w_12305 , w_12306 );
and ( \3859_b0 , \1255_b0 , w_12307 );
and ( w_12306 ,  , w_12307 );
buf ( w_12305 , \1263_b1 );
not ( w_12305 , w_12308 );
not (  , w_12309 );
and ( w_12308 , w_12309 , \1263_b0 );
buf ( \3860_b1 , \3859_b1 );
not ( \3860_b1 , w_12310 );
not ( \3860_b0 , w_12311 );
and ( w_12310 , w_12311 , \3859_b0 );
or ( \3861_b1 , \1426_b1 , w_12312 );
or ( \3861_b0 , \1426_b0 , \1253_b0 );
not ( \1253_b0 , w_12313 );
and ( w_12313 , w_12312 , \1253_b1 );
or ( \3862_b1 , \3861_b1 , w_12315 );
not ( w_12315 , w_12316 );
and ( \3862_b0 , \3861_b0 , w_12317 );
and ( w_12316 ,  , w_12317 );
buf ( w_12315 , \1260_b1 );
not ( w_12315 , w_12318 );
not (  , w_12319 );
and ( w_12318 , w_12319 , \1260_b0 );
buf ( \3863_b1 , \3862_b1 );
not ( \3863_b1 , w_12320 );
not ( \3863_b0 , w_12321 );
and ( w_12320 , w_12321 , \3862_b0 );
or ( \3864_b1 , \3860_b1 , w_12322 );
or ( \3864_b0 , \3860_b0 , \3863_b0 );
not ( \3863_b0 , w_12323 );
and ( w_12323 , w_12322 , \3863_b1 );
or ( \3865_b1 , \3862_b1 , w_12324 );
or ( \3865_b0 , \3862_b0 , \3859_b0 );
not ( \3859_b0 , w_12325 );
and ( w_12325 , w_12324 , \3859_b1 );
or ( \3866_b1 , \3864_b1 , w_12327 );
not ( w_12327 , w_12328 );
and ( \3866_b0 , \3864_b0 , w_12329 );
and ( w_12328 ,  , w_12329 );
buf ( w_12327 , \3865_b1 );
not ( w_12327 , w_12330 );
not (  , w_12331 );
and ( w_12330 , w_12331 , \3865_b0 );
buf ( \3867_b1 , \3866_b1 );
not ( \3867_b1 , w_12332 );
not ( \3867_b0 , w_12333 );
and ( w_12332 , w_12333 , \3866_b0 );
buf ( \3868_b1 , \3087_b1 );
not ( \3868_b1 , w_12334 );
not ( \3868_b0 , w_12335 );
and ( w_12334 , w_12335 , \3087_b0 );
or ( \3869_b1 , \3867_b1 , w_12336 );
or ( \3869_b0 , \3867_b0 , \3868_b0 );
not ( \3868_b0 , w_12337 );
and ( w_12337 , w_12336 , \3868_b1 );
or ( \3870_b1 , \1282_b1 , \d[5]_b1 );
not ( \d[5]_b1 , w_12338 );
and ( \3870_b0 , \1282_b0 , w_12339 );
and ( w_12338 , w_12339 , \d[5]_b0 );
or ( \3871_b1 , \c[5]_b1 , \1514_b1 );
not ( \1514_b1 , w_12340 );
and ( \3871_b0 , \c[5]_b0 , w_12341 );
and ( w_12340 , w_12341 , \1514_b0 );
or ( \3872_b1 , \1293_b1 , \b[5]_b1 );
not ( \b[5]_b1 , w_12342 );
and ( \3872_b0 , \1293_b0 , w_12343 );
and ( w_12342 , w_12343 , \b[5]_b0 );
or ( \3874_b1 , \3869_b1 , w_12345 );
not ( w_12345 , w_12346 );
and ( \3874_b0 , \3869_b0 , w_12347 );
and ( w_12346 ,  , w_12347 );
buf ( w_12345 , \3873_b1 );
not ( w_12345 , w_12348 );
not (  , w_12349 );
and ( w_12348 , w_12349 , \3873_b0 );
or ( \3875_b1 , \3858_b1 , w_12351 );
not ( w_12351 , w_12352 );
and ( \3875_b0 , \3858_b0 , w_12353 );
and ( w_12352 ,  , w_12353 );
buf ( w_12351 , \3874_b1 );
not ( w_12351 , w_12354 );
not (  , w_12355 );
and ( w_12354 , w_12355 , \3874_b0 );
or ( \3876_b1 , \3849_b1 , w_12357 );
not ( w_12357 , w_12358 );
and ( \3876_b0 , \3849_b0 , w_12359 );
and ( w_12358 ,  , w_12359 );
buf ( w_12357 , \3875_b1 );
not ( w_12357 , w_12360 );
not (  , w_12361 );
and ( w_12360 , w_12361 , \3875_b0 );
or ( \3877_b1 , \3840_b1 , w_12363 );
not ( w_12363 , w_12364 );
and ( \3877_b0 , \3840_b0 , w_12365 );
and ( w_12364 ,  , w_12365 );
buf ( w_12363 , \3876_b1 );
not ( w_12363 , w_12366 );
not (  , w_12367 );
and ( w_12366 , w_12367 , \3876_b0 );
or ( \3878_b1 , \3838_b1 , w_12369 );
not ( w_12369 , w_12370 );
and ( \3878_b0 , \3838_b0 , w_12371 );
and ( w_12370 ,  , w_12371 );
buf ( w_12369 , \3877_b1 );
not ( w_12369 , w_12372 );
not (  , w_12373 );
and ( w_12372 , w_12373 , \3877_b0 );
or ( \3879_b1 , \3834_b1 , w_12375 );
not ( w_12375 , w_12376 );
and ( \3879_b0 , \3834_b0 , w_12377 );
and ( w_12376 ,  , w_12377 );
buf ( w_12375 , \3878_b1 );
not ( w_12375 , w_12378 );
not (  , w_12379 );
and ( w_12378 , w_12379 , \3878_b0 );
or ( \3880_b1 , \3821_b1 , w_12381 );
not ( w_12381 , w_12382 );
and ( \3880_b0 , \3821_b0 , w_12383 );
and ( w_12382 ,  , w_12383 );
buf ( w_12381 , \3879_b1 );
not ( w_12381 , w_12384 );
not (  , w_12385 );
and ( w_12384 , w_12385 , \3879_b0 );
or ( \3881_b1 , \c[14]_b1 , w_12387 );
not ( w_12387 , w_12388 );
and ( \3881_b0 , \c[14]_b0 , w_12389 );
and ( w_12388 ,  , w_12389 );
buf ( w_12387 , \d[14]_b1 );
not ( w_12387 , w_12390 );
not (  , w_12391 );
and ( w_12390 , w_12391 , \d[14]_b0 );
buf ( \3882_b1 , \3881_b1 );
not ( \3882_b1 , w_12392 );
not ( \3882_b0 , w_12393 );
and ( w_12392 , w_12393 , \3881_b0 );
or ( \3883_b1 , \c[14]_b1 , w_12395 );
not ( w_12395 , w_12396 );
and ( \3883_b0 , \c[14]_b0 , w_12397 );
and ( w_12396 ,  , w_12397 );
buf ( w_12395 , \d[14]_b1 );
not ( w_12395 , w_12398 );
not (  , w_12399 );
and ( w_12398 , w_12399 , \d[14]_b0 );
or ( \3884_b1 , \3882_b1 , w_12401 );
not ( w_12401 , w_12402 );
and ( \3884_b0 , \3882_b0 , w_12403 );
and ( w_12402 ,  , w_12403 );
buf ( w_12401 , \3883_b1 );
not ( w_12401 , w_12404 );
not (  , w_12405 );
and ( w_12404 , w_12405 , \3883_b0 );
or ( \3885_b1 , \c[1]_b1 , w_12407 );
not ( w_12407 , w_12408 );
and ( \3885_b0 , \c[1]_b0 , w_12409 );
and ( w_12408 ,  , w_12409 );
buf ( w_12407 , \d[1]_b1 );
not ( w_12407 , w_12410 );
not (  , w_12411 );
and ( w_12410 , w_12411 , \d[1]_b0 );
or ( \3886_b1 , \c[0]_b1 , w_12413 );
not ( w_12413 , w_12414 );
and ( \3886_b0 , \c[0]_b0 , w_12415 );
and ( w_12414 ,  , w_12415 );
buf ( w_12413 , \d[0]_b1 );
not ( w_12413 , w_12416 );
not (  , w_12417 );
and ( w_12416 , w_12417 , \d[0]_b0 );
or ( \3887_b1 , \3885_b1 , \3886_b1 );
not ( \3886_b1 , w_12418 );
and ( \3887_b0 , \3885_b0 , w_12419 );
and ( w_12418 , w_12419 , \3886_b0 );
or ( \3888_b1 , \c[1]_b1 , w_12421 );
not ( w_12421 , w_12422 );
and ( \3888_b0 , \c[1]_b0 , w_12423 );
and ( w_12422 ,  , w_12423 );
buf ( w_12421 , \d[1]_b1 );
not ( w_12421 , w_12424 );
not (  , w_12425 );
and ( w_12424 , w_12425 , \d[1]_b0 );
or ( \3889_b1 , \c[2]_b1 , w_12427 );
not ( w_12427 , w_12428 );
and ( \3889_b0 , \c[2]_b0 , w_12429 );
and ( w_12428 ,  , w_12429 );
buf ( w_12427 , \d[2]_b1 );
not ( w_12427 , w_12430 );
not (  , w_12431 );
and ( w_12430 , w_12431 , \d[2]_b0 );
buf ( \3891_b1 , \3890_b1 );
not ( \3891_b1 , w_12432 );
not ( \3891_b0 , w_12433 );
and ( w_12432 , w_12433 , \3890_b0 );
or ( \3892_b1 , \c[3]_b1 , w_12435 );
not ( w_12435 , w_12436 );
and ( \3892_b0 , \c[3]_b0 , w_12437 );
and ( w_12436 ,  , w_12437 );
buf ( w_12435 , \d[3]_b1 );
not ( w_12435 , w_12438 );
not (  , w_12439 );
and ( w_12438 , w_12439 , \d[3]_b0 );
or ( \3893_b1 , \c[2]_b1 , w_12441 );
not ( w_12441 , w_12442 );
and ( \3893_b0 , \c[2]_b0 , w_12443 );
and ( w_12442 ,  , w_12443 );
buf ( w_12441 , \d[2]_b1 );
not ( w_12441 , w_12444 );
not (  , w_12445 );
and ( w_12444 , w_12445 , \d[2]_b0 );
or ( \3895_b1 , \c[5]_b1 , w_12447 );
not ( w_12447 , w_12448 );
and ( \3895_b0 , \c[5]_b0 , w_12449 );
and ( w_12448 ,  , w_12449 );
buf ( w_12447 , \d[5]_b1 );
not ( w_12447 , w_12450 );
not (  , w_12451 );
and ( w_12450 , w_12451 , \d[5]_b0 );
or ( \3896_b1 , \c[4]_b1 , w_12453 );
not ( w_12453 , w_12454 );
and ( \3896_b0 , \c[4]_b0 , w_12455 );
and ( w_12454 ,  , w_12455 );
buf ( w_12453 , \d[4]_b1 );
not ( w_12453 , w_12456 );
not (  , w_12457 );
and ( w_12456 , w_12457 , \d[4]_b0 );
or ( \3897_b1 , \3895_b1 , w_12459 );
not ( w_12459 , w_12460 );
and ( \3897_b0 , \3895_b0 , w_12461 );
and ( w_12460 ,  , w_12461 );
buf ( w_12459 , \3896_b1 );
not ( w_12459 , w_12462 );
not (  , w_12463 );
and ( w_12462 , w_12463 , \3896_b0 );
or ( \3898_b1 , \c[7]_b1 , w_12465 );
not ( w_12465 , w_12466 );
and ( \3898_b0 , \c[7]_b0 , w_12467 );
and ( w_12466 ,  , w_12467 );
buf ( w_12465 , \d[7]_b1 );
not ( w_12465 , w_12468 );
not (  , w_12469 );
and ( w_12468 , w_12469 , \d[7]_b0 );
or ( \3899_b1 , \c[6]_b1 , w_12471 );
not ( w_12471 , w_12472 );
and ( \3899_b0 , \c[6]_b0 , w_12473 );
and ( w_12472 ,  , w_12473 );
buf ( w_12471 , \d[6]_b1 );
not ( w_12471 , w_12474 );
not (  , w_12475 );
and ( w_12474 , w_12475 , \d[6]_b0 );
or ( \3900_b1 , \3898_b1 , w_12477 );
not ( w_12477 , w_12478 );
and ( \3900_b0 , \3898_b0 , w_12479 );
and ( w_12478 ,  , w_12479 );
buf ( w_12477 , \3899_b1 );
not ( w_12477 , w_12480 );
not (  , w_12481 );
and ( w_12480 , w_12481 , \3899_b0 );
or ( \3901_b1 , \c[3]_b1 , w_12483 );
not ( w_12483 , w_12484 );
and ( \3901_b0 , \c[3]_b0 , w_12485 );
and ( w_12484 ,  , w_12485 );
buf ( w_12483 , \d[3]_b1 );
not ( w_12483 , w_12486 );
not (  , w_12487 );
and ( w_12486 , w_12487 , \d[3]_b0 );
buf ( \3902_b1 , \3901_b1 );
not ( \3902_b1 , w_12488 );
not ( \3902_b0 , w_12489 );
and ( w_12488 , w_12489 , \3901_b0 );
or ( \3904_b1 , \c[4]_b1 , w_12491 );
not ( w_12491 , w_12492 );
and ( \3904_b0 , \c[4]_b0 , w_12493 );
and ( w_12492 ,  , w_12493 );
buf ( w_12491 , \d[4]_b1 );
not ( w_12491 , w_12494 );
not (  , w_12495 );
and ( w_12494 , w_12495 , \d[4]_b0 );
or ( \3905_b1 , \3895_b1 , w_12497 );
not ( w_12497 , w_12498 );
and ( \3905_b0 , \3895_b0 , w_12499 );
and ( w_12498 ,  , w_12499 );
buf ( w_12497 , \3904_b1 );
not ( w_12497 , w_12500 );
not (  , w_12501 );
and ( w_12500 , w_12501 , \3904_b0 );
or ( \3906_b1 , \c[6]_b1 , w_12503 );
not ( w_12503 , w_12504 );
and ( \3906_b0 , \c[6]_b0 , w_12505 );
and ( w_12504 ,  , w_12505 );
buf ( w_12503 , \d[6]_b1 );
not ( w_12503 , w_12506 );
not (  , w_12507 );
and ( w_12506 , w_12507 , \d[6]_b0 );
or ( \3907_b1 , \c[7]_b1 , w_12509 );
not ( w_12509 , w_12510 );
and ( \3907_b0 , \c[7]_b0 , w_12511 );
and ( w_12510 ,  , w_12511 );
buf ( w_12509 , \d[7]_b1 );
not ( w_12509 , w_12512 );
not (  , w_12513 );
and ( w_12512 , w_12513 , \d[7]_b0 );
or ( \3908_b1 , \c[5]_b1 , w_12515 );
not ( w_12515 , w_12516 );
and ( \3908_b0 , \c[5]_b0 , w_12517 );
and ( w_12516 ,  , w_12517 );
buf ( w_12515 , \d[5]_b1 );
not ( w_12515 , w_12518 );
not (  , w_12519 );
and ( w_12518 , w_12519 , \d[5]_b0 );
or ( \3910_b1 , \3905_b1 , w_12520 );
or ( \3910_b0 , \3905_b0 , \3909_b0 );
not ( \3909_b0 , w_12521 );
and ( w_12521 , w_12520 , \3909_b1 );
buf ( \3911_b1 , \3907_b1 );
not ( \3911_b1 , w_12522 );
not ( \3911_b0 , w_12523 );
and ( w_12522 , w_12523 , \3907_b0 );
or ( \3912_b1 , \3900_b1 , w_12524 );
or ( \3912_b0 , \3900_b0 , \3911_b0 );
not ( \3911_b0 , w_12525 );
and ( w_12525 , w_12524 , \3911_b1 );
or ( \3913_b1 , \3910_b1 , w_12527 );
not ( w_12527 , w_12528 );
and ( \3913_b0 , \3910_b0 , w_12529 );
and ( w_12528 ,  , w_12529 );
buf ( w_12527 , \3912_b1 );
not ( w_12527 , w_12530 );
not (  , w_12531 );
and ( w_12530 , w_12531 , \3912_b0 );
or ( \3914_b1 , \3903_b1 , w_12533 );
not ( w_12533 , w_12534 );
and ( \3914_b0 , \3903_b0 , w_12535 );
and ( w_12534 ,  , w_12535 );
buf ( w_12533 , \3913_b1 );
not ( w_12533 , w_12536 );
not (  , w_12537 );
and ( w_12536 , w_12537 , \3913_b0 );
or ( \3915_b1 , \c[11]_b1 , w_12539 );
not ( w_12539 , w_12540 );
and ( \3915_b0 , \c[11]_b0 , w_12541 );
and ( w_12540 ,  , w_12541 );
buf ( w_12539 , \d[11]_b1 );
not ( w_12539 , w_12542 );
not (  , w_12543 );
and ( w_12542 , w_12543 , \d[11]_b0 );
or ( \3916_b1 , \c[10]_b1 , w_12545 );
not ( w_12545 , w_12546 );
and ( \3916_b0 , \c[10]_b0 , w_12547 );
and ( w_12546 ,  , w_12547 );
buf ( w_12545 , \d[10]_b1 );
not ( w_12545 , w_12548 );
not (  , w_12549 );
and ( w_12548 , w_12549 , \d[10]_b0 );
or ( \3917_b1 , \3915_b1 , w_12551 );
not ( w_12551 , w_12552 );
and ( \3917_b0 , \3915_b0 , w_12553 );
and ( w_12552 ,  , w_12553 );
buf ( w_12551 , \3916_b1 );
not ( w_12551 , w_12554 );
not (  , w_12555 );
and ( w_12554 , w_12555 , \3916_b0 );
or ( \3918_b1 , \c[9]_b1 , w_12557 );
not ( w_12557 , w_12558 );
and ( \3918_b0 , \c[9]_b0 , w_12559 );
and ( w_12558 ,  , w_12559 );
buf ( w_12557 , \d[9]_b1 );
not ( w_12557 , w_12560 );
not (  , w_12561 );
and ( w_12560 , w_12561 , \d[9]_b0 );
or ( \3919_b1 , \c[8]_b1 , w_12563 );
not ( w_12563 , w_12564 );
and ( \3919_b0 , \c[8]_b0 , w_12565 );
and ( w_12564 ,  , w_12565 );
buf ( w_12563 , \d[8]_b1 );
not ( w_12563 , w_12566 );
not (  , w_12567 );
and ( w_12566 , w_12567 , \d[8]_b0 );
or ( \3920_b1 , \3918_b1 , w_12569 );
not ( w_12569 , w_12570 );
and ( \3920_b0 , \3918_b0 , w_12571 );
and ( w_12570 ,  , w_12571 );
buf ( w_12569 , \3919_b1 );
not ( w_12569 , w_12572 );
not (  , w_12573 );
and ( w_12572 , w_12573 , \3919_b0 );
or ( \3921_b1 , \3917_b1 , \3920_b1 );
not ( \3920_b1 , w_12574 );
and ( \3921_b0 , \3917_b0 , w_12575 );
and ( w_12574 , w_12575 , \3920_b0 );
or ( \3922_b1 , \c[13]_b1 , w_12577 );
not ( w_12577 , w_12578 );
and ( \3922_b0 , \c[13]_b0 , w_12579 );
and ( w_12578 ,  , w_12579 );
buf ( w_12577 , \d[13]_b1 );
not ( w_12577 , w_12580 );
not (  , w_12581 );
and ( w_12580 , w_12581 , \d[13]_b0 );
or ( \3923_b1 , \c[12]_b1 , w_12583 );
not ( w_12583 , w_12584 );
and ( \3923_b0 , \c[12]_b0 , w_12585 );
and ( w_12584 ,  , w_12585 );
buf ( w_12583 , \d[12]_b1 );
not ( w_12583 , w_12586 );
not (  , w_12587 );
and ( w_12586 , w_12587 , \d[12]_b0 );
or ( \3924_b1 , \3922_b1 , w_12589 );
not ( w_12589 , w_12590 );
and ( \3924_b0 , \3922_b0 , w_12591 );
and ( w_12590 ,  , w_12591 );
buf ( w_12589 , \3923_b1 );
not ( w_12589 , w_12592 );
not (  , w_12593 );
and ( w_12592 , w_12593 , \3923_b0 );
or ( \3926_b1 , \c[12]_b1 , w_12595 );
not ( w_12595 , w_12596 );
and ( \3926_b0 , \c[12]_b0 , w_12597 );
and ( w_12596 ,  , w_12597 );
buf ( w_12595 , \d[12]_b1 );
not ( w_12595 , w_12598 );
not (  , w_12599 );
and ( w_12598 , w_12599 , \d[12]_b0 );
or ( \3927_b1 , \3922_b1 , w_12600 );
or ( \3927_b0 , \3922_b0 , \3926_b0 );
not ( \3926_b0 , w_12601 );
and ( w_12601 , w_12600 , \3926_b1 );
or ( \3928_b1 , \c[13]_b1 , w_12603 );
not ( w_12603 , w_12604 );
and ( \3928_b0 , \c[13]_b0 , w_12605 );
and ( w_12604 ,  , w_12605 );
buf ( w_12603 , \d[13]_b1 );
not ( w_12603 , w_12606 );
not (  , w_12607 );
and ( w_12606 , w_12607 , \d[13]_b0 );
or ( \3929_b1 , \3927_b1 , w_12609 );
not ( w_12609 , w_12610 );
and ( \3929_b0 , \3927_b0 , w_12611 );
and ( w_12610 ,  , w_12611 );
buf ( w_12609 , \3928_b1 );
not ( w_12609 , w_12612 );
not (  , w_12613 );
and ( w_12612 , w_12613 , \3928_b0 );
buf ( \3930_b1 , \3929_b1 );
not ( \3930_b1 , w_12614 );
not ( \3930_b0 , w_12615 );
and ( w_12614 , w_12615 , \3929_b0 );
or ( \3931_b1 , \c[10]_b1 , w_12617 );
not ( w_12617 , w_12618 );
and ( \3931_b0 , \c[10]_b0 , w_12619 );
and ( w_12618 ,  , w_12619 );
buf ( w_12617 , \d[10]_b1 );
not ( w_12617 , w_12620 );
not (  , w_12621 );
and ( w_12620 , w_12621 , \d[10]_b0 );
or ( \3932_b1 , \3915_b1 , w_12622 );
or ( \3932_b0 , \3915_b0 , \3931_b0 );
not ( \3931_b0 , w_12623 );
and ( w_12623 , w_12622 , \3931_b1 );
or ( \3933_b1 , \c[8]_b1 , w_12625 );
not ( w_12625 , w_12626 );
and ( \3933_b0 , \c[8]_b0 , w_12627 );
and ( w_12626 ,  , w_12627 );
buf ( w_12625 , \d[8]_b1 );
not ( w_12625 , w_12628 );
not (  , w_12629 );
and ( w_12628 , w_12629 , \d[8]_b0 );
or ( \3934_b1 , \3918_b1 , w_12630 );
or ( \3934_b0 , \3918_b0 , \3933_b0 );
not ( \3933_b0 , w_12631 );
and ( w_12631 , w_12630 , \3933_b1 );
or ( \3935_b1 , \c[9]_b1 , w_12633 );
not ( w_12633 , w_12634 );
and ( \3935_b0 , \c[9]_b0 , w_12635 );
and ( w_12634 ,  , w_12635 );
buf ( w_12633 , \d[9]_b1 );
not ( w_12633 , w_12636 );
not (  , w_12637 );
and ( w_12636 , w_12637 , \d[9]_b0 );
or ( \3936_b1 , \3934_b1 , w_12639 );
not ( w_12639 , w_12640 );
and ( \3936_b0 , \3934_b0 , w_12641 );
and ( w_12640 ,  , w_12641 );
buf ( w_12639 , \3935_b1 );
not ( w_12639 , w_12642 );
not (  , w_12643 );
and ( w_12642 , w_12643 , \3935_b0 );
or ( \3937_b1 , \3917_b1 , w_12645 );
not ( w_12645 , w_12646 );
and ( \3937_b0 , \3917_b0 , w_12647 );
and ( w_12646 ,  , w_12647 );
buf ( w_12645 , \3936_b1 );
not ( w_12645 , w_12648 );
not (  , w_12649 );
and ( w_12648 , w_12649 , \3936_b0 );
or ( \3938_b1 , \c[11]_b1 , w_12651 );
not ( w_12651 , w_12652 );
and ( \3938_b0 , \c[11]_b0 , w_12653 );
and ( w_12652 ,  , w_12653 );
buf ( w_12651 , \d[11]_b1 );
not ( w_12651 , w_12654 );
not (  , w_12655 );
and ( w_12654 , w_12655 , \d[11]_b0 );
or ( \3940_b1 , \3939_b1 , w_12657 );
not ( w_12657 , w_12658 );
and ( \3940_b0 , \3939_b0 , w_12659 );
and ( w_12658 ,  , w_12659 );
buf ( w_12657 , \3924_b1 );
not ( w_12657 , w_12660 );
not (  , w_12661 );
and ( w_12660 , w_12661 , \3924_b0 );
or ( \3941_b1 , \3930_b1 , w_12663 );
not ( w_12663 , w_12664 );
and ( \3941_b0 , \3930_b0 , w_12665 );
and ( w_12664 ,  , w_12665 );
buf ( w_12663 , \3940_b1 );
not ( w_12663 , w_12666 );
not (  , w_12667 );
and ( w_12666 , w_12667 , \3940_b0 );
or ( \3942_b1 , \3925_b1 , w_12669 );
not ( w_12669 , w_12670 );
and ( \3942_b0 , \3925_b0 , w_12671 );
and ( w_12670 ,  , w_12671 );
buf ( w_12669 , \3941_b1 );
not ( w_12669 , w_12672 );
not (  , w_12673 );
and ( w_12672 , w_12673 , \3941_b0 );
or ( \3943_b1 , \3884_b1 , \3942_b1 );
xor ( \3943_b0 , \3884_b0 , w_12674 );
not ( w_12674 , w_12675 );
and ( w_12675 , \3942_b1 , \3942_b0 );
buf ( \3944_b1 , \3899_b1 );
not ( \3944_b1 , w_12676 );
not ( \3944_b0 , w_12677 );
and ( w_12676 , w_12677 , \3899_b0 );
or ( \3945_b1 , \3944_b1 , w_12679 );
not ( w_12679 , w_12680 );
and ( \3945_b0 , \3944_b0 , w_12681 );
and ( w_12680 ,  , w_12681 );
buf ( w_12679 , \3906_b1 );
not ( w_12679 , w_12682 );
not (  , w_12683 );
and ( w_12682 , w_12683 , \3906_b0 );
or ( \3946_b1 , \3888_b1 , w_12684 );
or ( \3946_b0 , \3888_b0 , \3886_b0 );
not ( \3886_b0 , w_12685 );
and ( w_12685 , w_12684 , \3886_b1 );
or ( \3947_b1 , \3946_b1 , w_12687 );
not ( w_12687 , w_12688 );
and ( \3947_b0 , \3946_b0 , w_12689 );
and ( w_12688 ,  , w_12689 );
buf ( w_12687 , \3885_b1 );
not ( w_12687 , w_12690 );
not (  , w_12691 );
and ( w_12690 , w_12691 , \3885_b0 );
or ( \3948_b1 , \3901_b1 , w_12693 );
not ( w_12693 , w_12694 );
and ( \3948_b0 , \3901_b0 , w_12695 );
and ( w_12694 ,  , w_12695 );
buf ( w_12693 , \3889_b1 );
not ( w_12693 , w_12696 );
not (  , w_12697 );
and ( w_12696 , w_12697 , \3889_b0 );
or ( \3949_b1 , \3947_b1 , \3948_b1 );
not ( \3948_b1 , w_12698 );
and ( \3949_b0 , \3947_b0 , w_12699 );
and ( w_12698 , w_12699 , \3948_b0 );
or ( \3950_b1 , \3901_b1 , w_12700 );
or ( \3950_b0 , \3901_b0 , \3893_b0 );
not ( \3893_b0 , w_12701 );
and ( w_12701 , w_12700 , \3893_b1 );
or ( \3951_b1 , \3950_b1 , w_12703 );
not ( w_12703 , w_12704 );
and ( \3951_b0 , \3950_b0 , w_12705 );
and ( w_12704 ,  , w_12705 );
buf ( w_12703 , \3892_b1 );
not ( w_12703 , w_12706 );
not (  , w_12707 );
and ( w_12706 , w_12707 , \3892_b0 );
or ( \3952_b1 , \3949_b1 , w_12709 );
not ( w_12709 , w_12710 );
and ( \3952_b0 , \3949_b0 , w_12711 );
and ( w_12710 ,  , w_12711 );
buf ( w_12709 , \3951_b1 );
not ( w_12709 , w_12712 );
not (  , w_12713 );
and ( w_12712 , w_12713 , \3951_b0 );
buf ( \3953_b1 , \3952_b1 );
not ( \3953_b1 , w_12714 );
not ( \3953_b0 , w_12715 );
and ( w_12714 , w_12715 , \3952_b0 );
or ( \3954_b1 , \3953_b1 , w_12717 );
not ( w_12717 , w_12718 );
and ( \3954_b0 , \3953_b0 , w_12719 );
and ( w_12718 ,  , w_12719 );
buf ( w_12717 , \3897_b1 );
not ( w_12717 , w_12720 );
not (  , w_12721 );
and ( w_12720 , w_12721 , \3897_b0 );
buf ( \3955_b1 , \3908_b1 );
not ( \3955_b1 , w_12722 );
not ( \3955_b0 , w_12723 );
and ( w_12722 , w_12723 , \3908_b0 );
or ( \3956_b1 , \3955_b1 , w_12725 );
not ( w_12725 , w_12726 );
and ( \3956_b0 , \3955_b0 , w_12727 );
and ( w_12726 ,  , w_12727 );
buf ( w_12725 , \3905_b1 );
not ( w_12725 , w_12728 );
not (  , w_12729 );
and ( w_12728 , w_12729 , \3905_b0 );
or ( \3957_b1 , \3954_b1 , \3956_b1 );
not ( \3956_b1 , w_12730 );
and ( \3957_b0 , \3954_b0 , w_12731 );
and ( w_12730 , w_12731 , \3956_b0 );
or ( \3958_b1 , \3945_b1 , \3957_b1 );
xor ( \3958_b0 , \3945_b0 , w_12732 );
not ( w_12732 , w_12733 );
and ( w_12733 , \3957_b1 , \3957_b0 );
buf ( \3959_b1 , \3908_b1 );
not ( \3959_b1 , w_12734 );
not ( \3959_b0 , w_12735 );
and ( w_12734 , w_12735 , \3908_b0 );
or ( \3960_b1 , \3959_b1 , w_12737 );
not ( w_12737 , w_12738 );
and ( \3960_b0 , \3959_b0 , w_12739 );
and ( w_12738 ,  , w_12739 );
buf ( w_12737 , \3895_b1 );
not ( w_12737 , w_12740 );
not (  , w_12741 );
and ( w_12740 , w_12741 , \3895_b0 );
or ( \3961_b1 , \3952_b1 , w_12742 );
or ( \3961_b0 , \3952_b0 , \3896_b0 );
not ( \3896_b0 , w_12743 );
and ( w_12743 , w_12742 , \3896_b1 );
or ( \3962_b1 , \3961_b1 , w_12745 );
not ( w_12745 , w_12746 );
and ( \3962_b0 , \3961_b0 , w_12747 );
and ( w_12746 ,  , w_12747 );
buf ( w_12745 , \3904_b1 );
not ( w_12745 , w_12748 );
not (  , w_12749 );
and ( w_12748 , w_12749 , \3904_b0 );
or ( \3963_b1 , \3960_b1 , \3962_b1 );
xor ( \3963_b0 , \3960_b0 , w_12750 );
not ( w_12750 , w_12751 );
and ( w_12751 , \3962_b1 , \3962_b0 );
or ( \3964_b1 , \3914_b1 , \3920_b1 );
not ( \3920_b1 , w_12752 );
and ( \3964_b0 , \3914_b0 , w_12753 );
and ( w_12752 , w_12753 , \3920_b0 );
or ( \3965_b1 , \3964_b1 , w_12755 );
not ( w_12755 , w_12756 );
and ( \3965_b0 , \3964_b0 , w_12757 );
and ( w_12756 ,  , w_12757 );
buf ( w_12755 , \3936_b1 );
not ( w_12755 , w_12758 );
not (  , w_12759 );
and ( w_12758 , w_12759 , \3936_b0 );
buf ( \3966_b1 , \3923_b1 );
not ( \3966_b1 , w_12760 );
not ( \3966_b0 , w_12761 );
and ( w_12760 , w_12761 , \3923_b0 );
buf ( \3968_b1 , \3939_b1 );
not ( \3968_b1 , w_12762 );
not ( \3968_b0 , w_12763 );
and ( w_12762 , w_12763 , \3939_b0 );
or ( \3969_b1 , \3968_b1 , w_12764 );
or ( \3969_b0 , \3968_b0 , \3923_b0 );
not ( \3923_b0 , w_12765 );
and ( w_12765 , w_12764 , \3923_b1 );
or ( \3970_b1 , \3969_b1 , w_12767 );
not ( w_12767 , w_12768 );
and ( \3970_b0 , \3969_b0 , w_12769 );
and ( w_12768 ,  , w_12769 );
buf ( w_12767 , \3926_b1 );
not ( w_12767 , w_12770 );
not (  , w_12771 );
and ( w_12770 , w_12771 , \3926_b0 );
or ( \3971_b1 , \3967_b1 , w_12773 );
not ( w_12773 , w_12774 );
and ( \3971_b0 , \3967_b0 , w_12775 );
and ( w_12774 ,  , w_12775 );
buf ( w_12773 , \3970_b1 );
not ( w_12773 , w_12776 );
not (  , w_12777 );
and ( w_12776 , w_12777 , \3970_b0 );
buf ( \3972_b1 , \3914_b1 );
not ( \3972_b1 , w_12778 );
not ( \3972_b0 , w_12779 );
and ( w_12778 , w_12779 , \3914_b0 );
or ( \3973_b1 , \3972_b1 , w_12780 );
or ( \3973_b0 , \3972_b0 , \3919_b0 );
not ( \3919_b0 , w_12781 );
and ( w_12781 , w_12780 , \3919_b1 );
or ( \3974_b1 , \3973_b1 , w_12783 );
not ( w_12783 , w_12784 );
and ( \3974_b0 , \3973_b0 , w_12785 );
and ( w_12784 ,  , w_12785 );
buf ( w_12783 , \3933_b1 );
not ( w_12783 , w_12786 );
not (  , w_12787 );
and ( w_12786 , w_12787 , \3933_b0 );
buf ( \3975_b1 , \3924_b1 );
not ( \3975_b1 , w_12788 );
not ( \3975_b0 , w_12789 );
and ( w_12788 , w_12789 , \3924_b0 );
or ( \3976_b1 , \3975_b1 , w_12791 );
not ( w_12791 , w_12792 );
and ( \3976_b0 , \3975_b0 , w_12793 );
and ( w_12792 ,  , w_12793 );
buf ( w_12791 , \3881_b1 );
not ( w_12791 , w_12794 );
not (  , w_12795 );
and ( w_12794 , w_12795 , \3881_b0 );
or ( \3978_b1 , \3939_b1 , w_12797 );
not ( w_12797 , w_12798 );
and ( \3978_b0 , \3939_b0 , w_12799 );
and ( w_12798 ,  , w_12799 );
buf ( w_12797 , \3976_b1 );
not ( w_12797 , w_12800 );
not (  , w_12801 );
and ( w_12800 , w_12801 , \3976_b0 );
buf ( \3979_b1 , \3881_b1 );
not ( \3979_b1 , w_12802 );
not ( \3979_b0 , w_12803 );
and ( w_12802 , w_12803 , \3881_b0 );
or ( \3980_b1 , \3979_b1 , w_12805 );
not ( w_12805 , w_12806 );
and ( \3980_b0 , \3979_b0 , w_12807 );
and ( w_12806 ,  , w_12807 );
buf ( w_12805 , \3929_b1 );
not ( w_12805 , w_12808 );
not (  , w_12809 );
and ( w_12808 , w_12809 , \3929_b0 );
or ( \3982_b1 , \3977_b1 , w_12811 );
not ( w_12811 , w_12812 );
and ( \3982_b0 , \3977_b0 , w_12813 );
and ( w_12812 ,  , w_12813 );
buf ( w_12811 , \3981_b1 );
not ( w_12811 , w_12814 );
not (  , w_12815 );
and ( w_12814 , w_12815 , \3981_b0 );
buf ( \3983_b1 , \3921_b1 );
not ( \3983_b1 , w_12816 );
not ( \3983_b0 , w_12817 );
and ( w_12816 , w_12817 , \3921_b0 );
or ( \3984_b1 , \c[15]_b1 , w_12819 );
not ( w_12819 , w_12820 );
and ( \3984_b0 , \c[15]_b0 , w_12821 );
and ( w_12820 ,  , w_12821 );
buf ( w_12819 , \d[15]_b1 );
not ( w_12819 , w_12822 );
not (  , w_12823 );
and ( w_12822 , w_12823 , \d[15]_b0 );
or ( \3985_b1 , \3881_b1 , w_12825 );
not ( w_12825 , w_12826 );
and ( \3985_b0 , \3881_b0 , w_12827 );
and ( w_12826 ,  , w_12827 );
buf ( w_12825 , \3984_b1 );
not ( w_12825 , w_12828 );
not (  , w_12829 );
and ( w_12828 , w_12829 , \3984_b0 );
or ( \3986_b1 , \3985_b1 , w_12831 );
not ( w_12831 , w_12832 );
and ( \3986_b0 , \3985_b0 , w_12833 );
and ( w_12832 ,  , w_12833 );
buf ( w_12831 , \3924_b1 );
not ( w_12831 , w_12834 );
not (  , w_12835 );
and ( w_12834 , w_12835 , \3924_b0 );
or ( \3988_b1 , \3929_b1 , \3985_b1 );
not ( \3985_b1 , w_12836 );
and ( \3988_b0 , \3929_b0 , w_12837 );
and ( w_12836 , w_12837 , \3985_b0 );
or ( \3989_b1 , \3968_b1 , w_12839 );
not ( w_12839 , w_12840 );
and ( \3989_b0 , \3968_b0 , w_12841 );
and ( w_12840 ,  , w_12841 );
buf ( w_12839 , \3986_b1 );
not ( w_12839 , w_12842 );
not (  , w_12843 );
and ( w_12842 , w_12843 , \3986_b0 );
or ( \3990_b1 , \3984_b1 , w_12844 );
or ( \3990_b0 , \3984_b0 , \3883_b0 );
not ( \3883_b0 , w_12845 );
and ( w_12845 , w_12844 , \3883_b1 );
or ( \3991_b1 , \c[15]_b1 , w_12847 );
not ( w_12847 , w_12848 );
and ( \3991_b0 , \c[15]_b0 , w_12849 );
and ( w_12848 ,  , w_12849 );
buf ( w_12847 , \d[15]_b1 );
not ( w_12847 , w_12850 );
not (  , w_12851 );
and ( w_12850 , w_12851 , \d[15]_b0 );
or ( \3992_b1 , \3990_b1 , w_12853 );
not ( w_12853 , w_12854 );
and ( \3992_b0 , \3990_b0 , w_12855 );
and ( w_12854 ,  , w_12855 );
buf ( w_12853 , \3991_b1 );
not ( w_12853 , w_12856 );
not (  , w_12857 );
and ( w_12856 , w_12857 , \3991_b0 );
or ( \3994_b1 , \3987_b1 , w_12859 );
not ( w_12859 , w_12860 );
and ( \3994_b0 , \3987_b0 , w_12861 );
and ( w_12860 ,  , w_12861 );
buf ( w_12859 , \3993_b1 );
not ( w_12859 , w_12862 );
not (  , w_12863 );
and ( w_12862 , w_12863 , \3993_b0 );
buf ( \3995_b1 , \3916_b1 );
not ( \3995_b1 , w_12864 );
not ( \3995_b0 , w_12865 );
and ( w_12864 , w_12865 , \3916_b0 );
buf ( \3997_b1 , \3995_b1 );
not ( \3997_b1 , w_12866 );
not ( \3997_b0 , w_12867 );
and ( w_12866 , w_12867 , \3995_b0 );
buf ( \3998_b1 , \3936_b1 );
not ( \3998_b1 , w_12868 );
not ( \3998_b0 , w_12869 );
and ( w_12868 , w_12869 , \3936_b0 );
or ( \3999_b1 , \3997_b1 , w_12870 );
or ( \3999_b0 , \3997_b0 , \3998_b0 );
not ( \3998_b0 , w_12871 );
and ( w_12871 , w_12870 , \3998_b1 );
or ( \4000_b1 , \3999_b1 , w_12873 );
not ( w_12873 , w_12874 );
and ( \4000_b0 , \3999_b0 , w_12875 );
and ( w_12874 ,  , w_12875 );
buf ( w_12873 , \3931_b1 );
not ( w_12873 , w_12876 );
not (  , w_12877 );
and ( w_12876 , w_12877 , \3931_b0 );
or ( \4001_b1 , \3996_b1 , w_12879 );
not ( w_12879 , w_12880 );
and ( \4001_b0 , \3996_b0 , w_12881 );
and ( w_12880 ,  , w_12881 );
buf ( w_12879 , \4000_b1 );
not ( w_12879 , w_12882 );
not (  , w_12883 );
and ( w_12882 , w_12883 , \4000_b0 );
buf ( \4002_b1 , \3921_b1 );
not ( \4002_b1 , w_12884 );
not ( \4002_b0 , w_12885 );
and ( w_12884 , w_12885 , \3921_b0 );
buf ( \4003_b1 , \3914_b1 );
not ( \4003_b1 , w_12886 );
not ( \4003_b0 , w_12887 );
and ( w_12886 , w_12887 , \3914_b0 );
or ( \4004_b1 , \4002_b1 , w_12888 );
or ( \4004_b0 , \4002_b0 , \4003_b0 );
not ( \4003_b0 , w_12889 );
and ( w_12889 , w_12888 , \4003_b1 );
or ( \4005_b1 , \4004_b1 , w_12891 );
not ( w_12891 , w_12892 );
and ( \4005_b0 , \4004_b0 , w_12893 );
and ( w_12892 ,  , w_12893 );
buf ( w_12891 , \3968_b1 );
not ( w_12891 , w_12894 );
not (  , w_12895 );
and ( w_12894 , w_12895 , \3968_b0 );
buf ( \4006_b1 , \3919_b1 );
not ( \4006_b1 , w_12896 );
not ( \4006_b0 , w_12897 );
and ( w_12896 , w_12897 , \3919_b0 );
or ( \4007_b1 , \4006_b1 , w_12899 );
not ( w_12899 , w_12900 );
and ( \4007_b0 , \4006_b0 , w_12901 );
and ( w_12900 ,  , w_12901 );
buf ( w_12899 , \3933_b1 );
not ( w_12899 , w_12902 );
not (  , w_12903 );
and ( w_12902 , w_12903 , \3933_b0 );
or ( \4008_b1 , \4007_b1 , \3914_b1 );
not ( \3914_b1 , w_12904 );
and ( \4008_b0 , \4007_b0 , w_12905 );
and ( w_12904 , w_12905 , \3914_b0 );
buf ( \4009_b1 , \4007_b1 );
not ( \4009_b1 , w_12906 );
not ( \4009_b0 , w_12907 );
and ( w_12906 , w_12907 , \4007_b0 );
or ( \4010_b1 , \4009_b1 , \3972_b1 );
not ( \3972_b1 , w_12908 );
and ( \4010_b0 , \4009_b0 , w_12909 );
and ( w_12908 , w_12909 , \3972_b0 );
or ( \4011_b1 , \4008_b1 , w_12910 );
or ( \4011_b0 , \4008_b0 , \4010_b0 );
not ( \4010_b0 , w_12911 );
and ( w_12911 , w_12910 , \4010_b1 );
buf ( \4012_b1 , \3899_b1 );
not ( \4012_b1 , w_12912 );
not ( \4012_b0 , w_12913 );
and ( w_12912 , w_12913 , \3899_b0 );
or ( \4013_b1 , \4012_b1 , w_12915 );
not ( w_12915 , w_12916 );
and ( \4013_b0 , \4012_b0 , w_12917 );
and ( w_12916 ,  , w_12917 );
buf ( w_12915 , \3897_b1 );
not ( w_12915 , w_12918 );
not (  , w_12919 );
and ( w_12918 , w_12919 , \3897_b0 );
or ( \4014_b1 , \3952_b1 , w_12920 );
or ( \4014_b0 , \3952_b0 , \4013_b0 );
not ( \4013_b0 , w_12921 );
and ( w_12921 , w_12920 , \4013_b1 );
or ( \4015_b1 , \3899_b1 , w_12922 );
or ( \4015_b0 , \3899_b0 , \3956_b0 );
not ( \3956_b0 , w_12923 );
and ( w_12923 , w_12922 , \3956_b1 );
buf ( \4017_b1 , \3896_b1 );
not ( \4017_b1 , w_12924 );
not ( \4017_b0 , w_12925 );
and ( w_12924 , w_12925 , \3896_b0 );
or ( \4018_b1 , \4017_b1 , w_12927 );
not ( w_12927 , w_12928 );
and ( \4018_b0 , \4017_b0 , w_12929 );
and ( w_12928 ,  , w_12929 );
buf ( w_12927 , \3904_b1 );
not ( w_12927 , w_12930 );
not (  , w_12931 );
and ( w_12930 , w_12931 , \3904_b0 );
or ( \4019_b1 , \4018_b1 , \3952_b1 );
xor ( \4019_b0 , \4018_b0 , w_12932 );
not ( w_12932 , w_12933 );
and ( w_12933 , \3952_b1 , \3952_b0 );
or ( \4020_b1 , \3902_b1 , \3892_b1 );
not ( \3892_b1 , w_12934 );
and ( \4020_b0 , \3902_b0 , w_12935 );
and ( w_12934 , w_12935 , \3892_b0 );
buf ( \4021_b1 , \3890_b1 );
not ( \4021_b1 , w_12936 );
not ( \4021_b0 , w_12937 );
and ( w_12936 , w_12937 , \3890_b0 );
or ( \4022_b1 , \4021_b1 , w_12939 );
not ( w_12939 , w_12940 );
and ( \4022_b0 , \4021_b0 , w_12941 );
and ( w_12940 ,  , w_12941 );
buf ( w_12939 , \3893_b1 );
not ( w_12939 , w_12942 );
not (  , w_12943 );
and ( w_12942 , w_12943 , \3893_b0 );
or ( \4023_b1 , \4020_b1 , \4022_b1 );
xor ( \4023_b0 , \4020_b0 , w_12944 );
not ( w_12944 , w_12945 );
and ( w_12945 , \4022_b1 , \4022_b0 );
buf ( \4024_b1 , \3893_b1 );
not ( \4024_b1 , w_12946 );
not ( \4024_b0 , w_12947 );
and ( w_12946 , w_12947 , \3893_b0 );
or ( \4025_b1 , \4024_b1 , w_12949 );
not ( w_12949 , w_12950 );
and ( \4025_b0 , \4024_b0 , w_12951 );
and ( w_12950 ,  , w_12951 );
buf ( w_12949 , \3889_b1 );
not ( w_12949 , w_12952 );
not (  , w_12953 );
and ( w_12952 , w_12953 , \3889_b0 );
or ( \4026_b1 , \4025_b1 , \3947_b1 );
xor ( \4026_b0 , \4025_b0 , w_12954 );
not ( w_12954 , w_12955 );
and ( w_12955 , \3947_b1 , \3947_b0 );
buf ( \4027_b1 , \3888_b1 );
not ( \4027_b1 , w_12956 );
not ( \4027_b0 , w_12957 );
and ( w_12956 , w_12957 , \3888_b0 );
or ( \4028_b1 , \4027_b1 , w_12959 );
not ( w_12959 , w_12960 );
and ( \4028_b0 , \4027_b0 , w_12961 );
and ( w_12960 ,  , w_12961 );
buf ( w_12959 , \3885_b1 );
not ( w_12959 , w_12962 );
not (  , w_12963 );
and ( w_12962 , w_12963 , \3885_b0 );
or ( \4029_b1 , \3886_b1 , \4028_b1 );
xor ( \4029_b0 , \3886_b0 , w_12964 );
not ( w_12964 , w_12965 );
and ( w_12965 , \4028_b1 , \4028_b0 );
or ( \4030_b1 , \3966_b1 , w_12967 );
not ( w_12967 , w_12968 );
and ( \4030_b0 , \3966_b0 , w_12969 );
and ( w_12968 ,  , w_12969 );
buf ( w_12967 , \3926_b1 );
not ( w_12967 , w_12970 );
not (  , w_12971 );
and ( w_12970 , w_12971 , \3926_b0 );
buf ( \4031_b1 , \3915_b1 );
not ( \4031_b1 , w_12972 );
not ( \4031_b0 , w_12973 );
and ( w_12972 , w_12973 , \3915_b0 );
or ( \4032_b1 , \4031_b1 , w_12975 );
not ( w_12975 , w_12976 );
and ( \4032_b0 , \4031_b0 , w_12977 );
and ( w_12976 ,  , w_12977 );
buf ( w_12975 , \3938_b1 );
not ( w_12975 , w_12978 );
not (  , w_12979 );
and ( w_12978 , w_12979 , \3938_b0 );
or ( \4033_b1 , \3995_b1 , \3931_b1 );
not ( \3931_b1 , w_12980 );
and ( \4033_b0 , \3995_b0 , w_12981 );
and ( w_12980 , w_12981 , \3931_b0 );
buf ( \4034_b1 , \3935_b1 );
not ( \4034_b1 , w_12982 );
not ( \4034_b0 , w_12983 );
and ( w_12982 , w_12983 , \3935_b0 );
or ( \4035_b1 , \4034_b1 , w_12985 );
not ( w_12985 , w_12986 );
and ( \4035_b0 , \4034_b0 , w_12987 );
and ( w_12986 ,  , w_12987 );
buf ( w_12985 , \3918_b1 );
not ( w_12985 , w_12988 );
not (  , w_12989 );
and ( w_12988 , w_12989 , \3918_b0 );
or ( \4036_b1 , \3911_b1 , w_12990 );
or ( \4036_b0 , \3911_b0 , \3898_b0 );
not ( \3898_b0 , w_12991 );
and ( w_12991 , w_12990 , \3898_b1 );
buf ( \4037_b1 , \3991_b1 );
not ( \4037_b1 , w_12992 );
not ( \4037_b0 , w_12993 );
and ( w_12992 , w_12993 , \3991_b0 );
or ( \4038_b1 , \4037_b1 , w_12995 );
not ( w_12995 , w_12996 );
and ( \4038_b0 , \4037_b0 , w_12997 );
and ( w_12996 ,  , w_12997 );
buf ( w_12995 , \3984_b1 );
not ( w_12995 , w_12998 );
not (  , w_12999 );
and ( w_12998 , w_12999 , \3984_b0 );
buf ( \4039_b1 , \3922_b1 );
not ( \4039_b1 , w_13000 );
not ( \4039_b0 , w_13001 );
and ( w_13000 , w_13001 , \3922_b0 );
or ( \4040_b1 , \4039_b1 , w_13003 );
not ( w_13003 , w_13004 );
and ( \4040_b0 , \4039_b0 , w_13005 );
and ( w_13004 ,  , w_13005 );
buf ( w_13003 , \3928_b1 );
not ( w_13003 , w_13006 );
not (  , w_13007 );
and ( w_13006 , w_13007 , \3928_b0 );
or ( \4041_b1 , \4033_b1 , w_13008 );
xor ( \4041_b0 , \4033_b0 , w_13010 );
not ( w_13010 , w_13011 );
and ( w_13011 , w_13008 , w_13009 );
buf ( w_13008 , \3965_b1 );
not ( w_13008 , w_13012 );
not ( w_13009 , w_13013 );
and ( w_13012 , w_13013 , \3965_b0 );
or ( \4042_b1 , \4040_b1 , \3971_b1 );
xor ( \4042_b0 , \4040_b0 , w_13014 );
not ( w_13014 , w_13015 );
and ( w_13015 , \3971_b1 , \3971_b0 );
or ( \4043_b1 , \4035_b1 , \3974_b1 );
xor ( \4043_b0 , \4035_b0 , w_13016 );
not ( w_13016 , w_13017 );
and ( w_13017 , \3974_b1 , \3974_b0 );
or ( \4044_b1 , \4038_b1 , w_13018 );
xor ( \4044_b0 , \4038_b0 , w_13020 );
not ( w_13020 , w_13021 );
and ( w_13021 , w_13018 , w_13019 );
buf ( w_13018 , \3982_b1 );
not ( w_13018 , w_13022 );
not ( w_13019 , w_13023 );
and ( w_13022 , w_13023 , \3982_b0 );
or ( \4045_b1 , \4032_b1 , \4001_b1 );
xor ( \4045_b0 , \4032_b0 , w_13024 );
not ( w_13024 , w_13025 );
and ( w_13025 , \4001_b1 , \4001_b0 );
or ( \4046_b1 , \4036_b1 , w_13026 );
xor ( \4046_b0 , \4036_b0 , w_13028 );
not ( w_13028 , w_13029 );
and ( w_13029 , w_13026 , w_13027 );
buf ( w_13026 , \4016_b1 );
not ( w_13026 , w_13030 );
not ( w_13027 , w_13031 );
and ( w_13030 , w_13031 , \4016_b0 );
or ( \4047_b1 , \4005_b1 , w_13032 );
xor ( \4047_b0 , \4005_b0 , w_13034 );
not ( w_13034 , w_13035 );
and ( w_13035 , w_13032 , w_13033 );
buf ( w_13032 , \4030_b1 );
not ( w_13032 , w_13036 );
not ( w_13033 , w_13037 );
and ( w_13036 , w_13037 , \4030_b0 );
or ( \4048_b1 , \d[0]_b1 , \c[0]_b1 );
xor ( \4048_b0 , \d[0]_b0 , w_13038 );
not ( w_13038 , w_13039 );
and ( w_13039 , \c[0]_b1 , \c[0]_b0 );
buf ( \4049_b1 , \1454_b1 );
not ( \4049_b1 , w_13040 );
not ( \4049_b0 , w_13041 );
and ( w_13040 , w_13041 , \1454_b0 );
or ( \4050_b1 , \1528_b1 , \4049_b1 );
not ( \4049_b1 , w_13042 );
and ( \4050_b0 , \1528_b0 , w_13043 );
and ( w_13042 , w_13043 , \4049_b0 );
buf ( \4051_b1 , \1528_b1 );
not ( \4051_b1 , w_13044 );
not ( \4051_b0 , w_13045 );
and ( w_13044 , w_13045 , \1528_b0 );
or ( \4052_b1 , \4051_b1 , \1454_b1 );
not ( \1454_b1 , w_13046 );
and ( \4052_b0 , \4051_b0 , w_13047 );
and ( w_13046 , w_13047 , \1454_b0 );
or ( \4053_b1 , \4050_b1 , w_13049 );
not ( w_13049 , w_13050 );
and ( \4053_b0 , \4050_b0 , w_13051 );
and ( w_13050 ,  , w_13051 );
buf ( w_13049 , \4052_b1 );
not ( w_13049 , w_13052 );
not (  , w_13053 );
and ( w_13052 , w_13053 , \4052_b0 );
buf ( \4054_b1 , \4053_b1 );
not ( \4054_b1 , w_13054 );
not ( \4054_b0 , w_13055 );
and ( w_13054 , w_13055 , \4053_b0 );
buf ( \4055_b1 , \4054_b1 );
buf ( \4055_b0 , \4054_b0 );
buf ( \4056_b1 , \4055_b1 );
not ( \4056_b1 , w_13056 );
not ( \4056_b0 , w_13057 );
and ( w_13056 , w_13057 , \4055_b0 );
buf ( \4057_b1 , \4056_b1 );
not ( \4057_b1 , w_13058 );
not ( \4057_b0 , w_13059 );
and ( w_13058 , w_13059 , \4056_b0 );
buf ( \4058_b1 , \4049_b1 );
not ( \4058_b1 , w_13060 );
not ( \4058_b0 , w_13061 );
and ( w_13060 , w_13061 , \4049_b0 );
buf ( \4059_b1 , \3880_b1 );
not ( \4059_b1 , w_13062 );
not ( \4059_b0 , w_13063 );
and ( w_13062 , w_13063 , \3880_b0 );
or ( \4060_b1 , \4058_b1 , w_13064 );
or ( \4060_b0 , \4058_b0 , \4059_b0 );
not ( \4059_b0 , w_13065 );
and ( w_13065 , w_13064 , \4059_b1 );
buf ( \4061_b1 , \3880_b1 );
not ( \4061_b1 , w_13066 );
not ( \4061_b0 , w_13067 );
and ( w_13066 , w_13067 , \3880_b0 );
or ( \4062_b1 , \4061_b1 , w_13069 );
not ( w_13069 , w_13070 );
and ( \4062_b0 , \4061_b0 , w_13071 );
and ( w_13070 ,  , w_13071 );
buf ( w_13069 , \1454_b1 );
not ( w_13069 , w_13072 );
not (  , w_13073 );
and ( w_13072 , w_13073 , \1454_b0 );
or ( \4063_b1 , \4060_b1 , w_13075 );
not ( w_13075 , w_13076 );
and ( \4063_b0 , \4060_b0 , w_13077 );
and ( w_13076 ,  , w_13077 );
buf ( w_13075 , \4062_b1 );
not ( w_13075 , w_13078 );
not (  , w_13079 );
and ( w_13078 , w_13079 , \4062_b0 );
or ( \4064_b1 , \4053_b1 , w_13081 );
not ( w_13081 , w_13082 );
and ( \4064_b0 , \4053_b0 , w_13083 );
and ( w_13082 ,  , w_13083 );
buf ( w_13081 , \4063_b1 );
not ( w_13081 , w_13084 );
not (  , w_13085 );
and ( w_13084 , w_13085 , \4063_b0 );
buf ( \4065_b1 , \4064_b1 );
not ( \4065_b1 , w_13086 );
not ( \4065_b0 , w_13087 );
and ( w_13086 , w_13087 , \4064_b0 );
buf ( \4066_b1 , \4065_b1 );
not ( \4066_b1 , w_13088 );
not ( \4066_b0 , w_13089 );
and ( w_13088 , w_13089 , \4065_b0 );
buf ( \4067_b1 , \4066_b1 );
not ( \4067_b1 , w_13090 );
not ( \4067_b0 , w_13091 );
and ( w_13090 , w_13091 , \4066_b0 );
or ( \4068_b1 , \4057_b1 , w_13092 );
or ( \4068_b0 , \4057_b0 , \4067_b0 );
not ( \4067_b0 , w_13093 );
and ( w_13093 , w_13092 , \4067_b1 );
buf ( \4069_b1 , \4061_b1 );
buf ( \4069_b0 , \4061_b0 );
buf ( \4070_b1 , \4069_b1 );
not ( \4070_b1 , w_13094 );
not ( \4070_b0 , w_13095 );
and ( w_13094 , w_13095 , \4069_b0 );
or ( \4071_b1 , \4068_b1 , w_13097 );
not ( w_13097 , w_13098 );
and ( \4071_b0 , \4068_b0 , w_13099 );
and ( w_13098 ,  , w_13099 );
buf ( w_13097 , \4070_b1 );
not ( w_13097 , w_13100 );
not (  , w_13101 );
and ( w_13100 , w_13101 , \4070_b0 );
buf ( \4072_b1 , \4071_b1 );
not ( \4072_b1 , w_13102 );
not ( \4072_b0 , w_13103 );
and ( w_13102 , w_13103 , \4071_b0 );
buf ( \4073_b1 , \4072_b1 );
not ( \4073_b1 , w_13104 );
not ( \4073_b0 , w_13105 );
and ( w_13104 , w_13105 , \4072_b0 );
or ( \4074_b1 , \4061_b1 , \3272_b1 );
not ( \3272_b1 , w_13106 );
and ( \4074_b0 , \4061_b0 , w_13107 );
and ( w_13106 , w_13107 , \3272_b0 );
buf ( \4075_b1 , \4061_b1 );
not ( \4075_b1 , w_13108 );
not ( \4075_b0 , w_13109 );
and ( w_13108 , w_13109 , \4061_b0 );
buf ( \4076_b1 , \3272_b1 );
not ( \4076_b1 , w_13110 );
not ( \4076_b0 , w_13111 );
and ( w_13110 , w_13111 , \3272_b0 );
or ( \4077_b1 , \4075_b1 , \4076_b1 );
not ( \4076_b1 , w_13112 );
and ( \4077_b0 , \4075_b0 , w_13113 );
and ( w_13112 , w_13113 , \4076_b0 );
or ( \4078_b1 , \4074_b1 , w_13115 );
not ( w_13115 , w_13116 );
and ( \4078_b0 , \4074_b0 , w_13117 );
and ( w_13116 ,  , w_13117 );
buf ( w_13115 , \4077_b1 );
not ( w_13115 , w_13118 );
not (  , w_13119 );
and ( w_13118 , w_13119 , \4077_b0 );
buf ( \4079_b1 , \1336_b1 );
not ( \4079_b1 , w_13120 );
not ( \4079_b0 , w_13121 );
and ( w_13120 , w_13121 , \1336_b0 );
buf ( \4080_b1 , \4076_b1 );
not ( \4080_b1 , w_13122 );
not ( \4080_b0 , w_13123 );
and ( w_13122 , w_13123 , \4076_b0 );
or ( \4081_b1 , \4079_b1 , w_13124 );
or ( \4081_b0 , \4079_b0 , \4080_b0 );
not ( \4080_b0 , w_13125 );
and ( w_13125 , w_13124 , \4080_b1 );
buf ( \4082_b1 , \1336_b1 );
not ( \4082_b1 , w_13126 );
not ( \4082_b0 , w_13127 );
and ( w_13126 , w_13127 , \1336_b0 );
or ( \4083_b1 , \4082_b1 , w_13129 );
not ( w_13129 , w_13130 );
and ( \4083_b0 , \4082_b0 , w_13131 );
and ( w_13130 ,  , w_13131 );
buf ( w_13129 , \3272_b1 );
not ( w_13129 , w_13132 );
not (  , w_13133 );
and ( w_13132 , w_13133 , \3272_b0 );
or ( \4084_b1 , \4081_b1 , w_13135 );
not ( w_13135 , w_13136 );
and ( \4084_b0 , \4081_b0 , w_13137 );
and ( w_13136 ,  , w_13137 );
buf ( w_13135 , \4083_b1 );
not ( w_13135 , w_13138 );
not (  , w_13139 );
and ( w_13138 , w_13139 , \4083_b0 );
or ( \4085_b1 , \4078_b1 , \4084_b1 );
not ( \4084_b1 , w_13140 );
and ( \4085_b0 , \4078_b0 , w_13141 );
and ( w_13140 , w_13141 , \4084_b0 );
buf ( \4086_b1 , \4085_b1 );
buf ( \4086_b0 , \4085_b0 );
buf ( \4087_b1 , \4044_b1 );
not ( \4087_b1 , w_13142 );
not ( \4087_b0 , w_13143 );
and ( w_13142 , w_13143 , \4044_b0 );
buf ( \4088_b1 , \1336_b1 );
buf ( \4088_b0 , \1336_b0 );
buf ( \4089_b1 , \4088_b1 );
not ( \4089_b1 , w_13144 );
not ( \4089_b0 , w_13145 );
and ( w_13144 , w_13145 , \4088_b0 );
buf ( \4090_b1 , \4089_b1 );
not ( \4090_b1 , w_13146 );
not ( \4090_b0 , w_13147 );
and ( w_13146 , w_13147 , \4089_b0 );
or ( \4091_b1 , \4087_b1 , w_13148 );
or ( \4091_b0 , \4087_b0 , \4090_b0 );
not ( \4090_b0 , w_13149 );
and ( w_13149 , w_13148 , \4090_b1 );
buf ( \4092_b1 , \4044_b1 );
not ( \4092_b1 , w_13150 );
not ( \4092_b0 , w_13151 );
and ( w_13150 , w_13151 , \4044_b0 );
or ( \4093_b1 , \4088_b1 , w_13153 );
not ( w_13153 , w_13154 );
and ( \4093_b0 , \4088_b0 , w_13155 );
and ( w_13154 ,  , w_13155 );
buf ( w_13153 , \4092_b1 );
not ( w_13153 , w_13156 );
not (  , w_13157 );
and ( w_13156 , w_13157 , \4092_b0 );
or ( \4094_b1 , \4091_b1 , w_13159 );
not ( w_13159 , w_13160 );
and ( \4094_b0 , \4091_b0 , w_13161 );
and ( w_13160 ,  , w_13161 );
buf ( w_13159 , \4093_b1 );
not ( w_13159 , w_13162 );
not (  , w_13163 );
and ( w_13162 , w_13163 , \4093_b0 );
or ( \4095_b1 , \4086_b1 , \4094_b1 );
not ( \4094_b1 , w_13164 );
and ( \4095_b0 , \4086_b0 , w_13165 );
and ( w_13164 , w_13165 , \4094_b0 );
buf ( \4096_b1 , \3994_b1 );
not ( \4096_b1 , w_13166 );
not ( \4096_b0 , w_13167 );
and ( w_13166 , w_13167 , \3994_b0 );
buf ( \4097_b1 , \4089_b1 );
not ( \4097_b1 , w_13168 );
not ( \4097_b0 , w_13169 );
and ( w_13168 , w_13169 , \4089_b0 );
or ( \4098_b1 , \4096_b1 , w_13170 );
or ( \4098_b0 , \4096_b0 , \4097_b0 );
not ( \4097_b0 , w_13171 );
and ( w_13171 , w_13170 , \4097_b1 );
buf ( \4099_b1 , \3994_b1 );
not ( \4099_b1 , w_13172 );
not ( \4099_b0 , w_13173 );
and ( w_13172 , w_13173 , \3994_b0 );
or ( \4100_b1 , \4088_b1 , w_13175 );
not ( w_13175 , w_13176 );
and ( \4100_b0 , \4088_b0 , w_13177 );
and ( w_13176 ,  , w_13177 );
buf ( w_13175 , \4099_b1 );
not ( w_13175 , w_13178 );
not (  , w_13179 );
and ( w_13178 , w_13179 , \4099_b0 );
or ( \4101_b1 , \4098_b1 , w_13181 );
not ( w_13181 , w_13182 );
and ( \4101_b0 , \4098_b0 , w_13183 );
and ( w_13182 ,  , w_13183 );
buf ( w_13181 , \4100_b1 );
not ( w_13181 , w_13184 );
not (  , w_13185 );
and ( w_13184 , w_13185 , \4100_b0 );
buf ( \4102_b1 , \4101_b1 );
not ( \4102_b1 , w_13186 );
not ( \4102_b0 , w_13187 );
and ( w_13186 , w_13187 , \4101_b0 );
buf ( \4103_b1 , \4078_b1 );
buf ( \4103_b0 , \4078_b0 );
or ( \4104_b1 , \4102_b1 , w_13189 );
not ( w_13189 , w_13190 );
and ( \4104_b0 , \4102_b0 , w_13191 );
and ( w_13190 ,  , w_13191 );
buf ( w_13189 , \4103_b1 );
not ( w_13189 , w_13192 );
not (  , w_13193 );
and ( w_13192 , w_13193 , \4103_b0 );
or ( \4105_b1 , \4095_b1 , w_13195 );
not ( w_13195 , w_13196 );
and ( \4105_b0 , \4095_b0 , w_13197 );
and ( w_13196 ,  , w_13197 );
buf ( w_13195 , \4104_b1 );
not ( w_13195 , w_13198 );
not (  , w_13199 );
and ( w_13198 , w_13199 , \4104_b0 );
buf ( \4106_b1 , \4105_b1 );
not ( \4106_b1 , w_13200 );
not ( \4106_b0 , w_13201 );
and ( w_13200 , w_13201 , \4105_b0 );
or ( \4107_b1 , \4073_b1 , w_13202 );
or ( \4107_b0 , \4073_b0 , \4106_b0 );
not ( \4106_b0 , w_13203 );
and ( w_13203 , w_13202 , \4106_b1 );
buf ( \4108_b1 , \4042_b1 );
not ( \4108_b1 , w_13204 );
not ( \4108_b0 , w_13205 );
and ( w_13204 , w_13205 , \4042_b0 );
buf ( \4109_b1 , \3745_b1 );
buf ( \4109_b0 , \3745_b0 );
buf ( \4110_b1 , \4109_b1 );
not ( \4110_b1 , w_13206 );
not ( \4110_b0 , w_13207 );
and ( w_13206 , w_13207 , \4109_b0 );
buf ( \4111_b1 , \4110_b1 );
not ( \4111_b1 , w_13208 );
not ( \4111_b0 , w_13209 );
and ( w_13208 , w_13209 , \4110_b0 );
or ( \4112_b1 , \4108_b1 , w_13210 );
or ( \4112_b0 , \4108_b0 , \4111_b0 );
not ( \4111_b0 , w_13211 );
and ( w_13211 , w_13210 , \4111_b1 );
buf ( \4113_b1 , \3745_b1 );
buf ( \4113_b0 , \3745_b0 );
buf ( \4114_b1 , \4113_b1 );
not ( \4114_b1 , w_13212 );
not ( \4114_b0 , w_13213 );
and ( w_13212 , w_13213 , \4113_b0 );
buf ( \4115_b1 , \4114_b1 );
not ( \4115_b1 , w_13214 );
not ( \4115_b0 , w_13215 );
and ( w_13214 , w_13215 , \4114_b0 );
buf ( \4116_b1 , \4042_b1 );
not ( \4116_b1 , w_13216 );
not ( \4116_b0 , w_13217 );
and ( w_13216 , w_13217 , \4042_b0 );
or ( \4117_b1 , \4115_b1 , w_13219 );
not ( w_13219 , w_13220 );
and ( \4117_b0 , \4115_b0 , w_13221 );
and ( w_13220 ,  , w_13221 );
buf ( w_13219 , \4116_b1 );
not ( w_13219 , w_13222 );
not (  , w_13223 );
and ( w_13222 , w_13223 , \4116_b0 );
or ( \4118_b1 , \4112_b1 , w_13225 );
not ( w_13225 , w_13226 );
and ( \4118_b0 , \4112_b0 , w_13227 );
and ( w_13226 ,  , w_13227 );
buf ( w_13225 , \4117_b1 );
not ( w_13225 , w_13228 );
not (  , w_13229 );
and ( w_13228 , w_13229 , \4117_b0 );
buf ( \4119_b1 , \4118_b1 );
not ( \4119_b1 , w_13230 );
not ( \4119_b0 , w_13231 );
and ( w_13230 , w_13231 , \4118_b0 );
buf ( \4120_b1 , \1336_b1 );
not ( \4120_b1 , w_13232 );
not ( \4120_b0 , w_13233 );
and ( w_13232 , w_13233 , \1336_b0 );
buf ( \4121_b1 , \3678_b1 );
not ( \4121_b1 , w_13234 );
not ( \4121_b0 , w_13235 );
and ( w_13234 , w_13235 , \3678_b0 );
buf ( \4122_b1 , \4121_b1 );
not ( \4122_b1 , w_13236 );
not ( \4122_b0 , w_13237 );
and ( w_13236 , w_13237 , \4121_b0 );
or ( \4123_b1 , \4120_b1 , w_13238 );
or ( \4123_b0 , \4120_b0 , \4122_b0 );
not ( \4122_b0 , w_13239 );
and ( w_13239 , w_13238 , \4122_b1 );
buf ( \4124_b1 , \1336_b1 );
not ( \4124_b1 , w_13240 );
not ( \4124_b0 , w_13241 );
and ( w_13240 , w_13241 , \1336_b0 );
or ( \4125_b1 , \4124_b1 , w_13243 );
not ( w_13243 , w_13244 );
and ( \4125_b0 , \4124_b0 , w_13245 );
and ( w_13244 ,  , w_13245 );
buf ( w_13243 , \3678_b1 );
not ( w_13243 , w_13246 );
not (  , w_13247 );
and ( w_13246 , w_13247 , \3678_b0 );
or ( \4126_b1 , \4123_b1 , w_13249 );
not ( w_13249 , w_13250 );
and ( \4126_b0 , \4123_b0 , w_13251 );
and ( w_13250 ,  , w_13251 );
buf ( w_13249 , \4125_b1 );
not ( w_13249 , w_13252 );
not (  , w_13253 );
and ( w_13252 , w_13253 , \4125_b0 );
buf ( \4127_b1 , \4126_b1 );
not ( \4127_b1 , w_13254 );
not ( \4127_b0 , w_13255 );
and ( w_13254 , w_13255 , \4126_b0 );
buf ( \4128_b1 , \3678_b1 );
not ( \4128_b1 , w_13256 );
not ( \4128_b0 , w_13257 );
and ( w_13256 , w_13257 , \3678_b0 );
buf ( \4129_b1 , \4128_b1 );
not ( \4129_b1 , w_13258 );
not ( \4129_b0 , w_13259 );
and ( w_13258 , w_13259 , \4128_b0 );
buf ( \4130_b1 , \3745_b1 );
not ( \4130_b1 , w_13260 );
not ( \4130_b0 , w_13261 );
and ( w_13260 , w_13261 , \3745_b0 );
or ( \4131_b1 , \4129_b1 , w_13262 );
or ( \4131_b0 , \4129_b0 , \4130_b0 );
not ( \4130_b0 , w_13263 );
and ( w_13263 , w_13262 , \4130_b1 );
buf ( \4132_b1 , \3745_b1 );
not ( \4132_b1 , w_13264 );
not ( \4132_b0 , w_13265 );
and ( w_13264 , w_13265 , \3745_b0 );
or ( \4133_b1 , \4132_b1 , w_13267 );
not ( w_13267 , w_13268 );
and ( \4133_b0 , \4132_b0 , w_13269 );
and ( w_13268 ,  , w_13269 );
buf ( w_13267 , \3678_b1 );
not ( w_13267 , w_13270 );
not (  , w_13271 );
and ( w_13270 , w_13271 , \3678_b0 );
or ( \4134_b1 , \4131_b1 , w_13273 );
not ( w_13273 , w_13274 );
and ( \4134_b0 , \4131_b0 , w_13275 );
and ( w_13274 ,  , w_13275 );
buf ( w_13273 , \4133_b1 );
not ( w_13273 , w_13276 );
not (  , w_13277 );
and ( w_13276 , w_13277 , \4133_b0 );
or ( \4135_b1 , \4127_b1 , w_13279 );
not ( w_13279 , w_13280 );
and ( \4135_b0 , \4127_b0 , w_13281 );
and ( w_13280 ,  , w_13281 );
buf ( w_13279 , \4134_b1 );
not ( w_13279 , w_13282 );
not (  , w_13283 );
and ( w_13282 , w_13283 , \4134_b0 );
buf ( \4136_b1 , \4135_b1 );
not ( \4136_b1 , w_13284 );
not ( \4136_b0 , w_13285 );
and ( w_13284 , w_13285 , \4135_b0 );
buf ( \4137_b1 , \4136_b1 );
not ( \4137_b1 , w_13286 );
not ( \4137_b0 , w_13287 );
and ( w_13286 , w_13287 , \4136_b0 );
or ( \4138_b1 , \4119_b1 , w_13288 );
or ( \4138_b0 , \4119_b0 , \4137_b0 );
not ( \4137_b0 , w_13289 );
and ( w_13289 , w_13288 , \4137_b1 );
buf ( \4139_b1 , \4126_b1 );
buf ( \4139_b0 , \4126_b0 );
buf ( \4140_b1 , \4139_b1 );
buf ( \4140_b0 , \4139_b0 );
buf ( \4141_b1 , \3943_b1 );
not ( \4141_b1 , w_13290 );
not ( \4141_b0 , w_13291 );
and ( w_13290 , w_13291 , \3943_b0 );
buf ( \4142_b1 , \4113_b1 );
not ( \4142_b1 , w_13292 );
not ( \4142_b0 , w_13293 );
and ( w_13292 , w_13293 , \4113_b0 );
buf ( \4143_b1 , \4142_b1 );
not ( \4143_b1 , w_13294 );
not ( \4143_b0 , w_13295 );
and ( w_13294 , w_13295 , \4142_b0 );
or ( \4144_b1 , \4141_b1 , w_13296 );
or ( \4144_b0 , \4141_b0 , \4143_b0 );
not ( \4143_b0 , w_13297 );
and ( w_13297 , w_13296 , \4143_b1 );
buf ( \4145_b1 , \4113_b1 );
not ( \4145_b1 , w_13298 );
not ( \4145_b0 , w_13299 );
and ( w_13298 , w_13299 , \4113_b0 );
buf ( \4146_b1 , \4145_b1 );
not ( \4146_b1 , w_13300 );
not ( \4146_b0 , w_13301 );
and ( w_13300 , w_13301 , \4145_b0 );
buf ( \4147_b1 , \3943_b1 );
not ( \4147_b1 , w_13302 );
not ( \4147_b0 , w_13303 );
and ( w_13302 , w_13303 , \3943_b0 );
or ( \4148_b1 , \4146_b1 , w_13305 );
not ( w_13305 , w_13306 );
and ( \4148_b0 , \4146_b0 , w_13307 );
and ( w_13306 ,  , w_13307 );
buf ( w_13305 , \4147_b1 );
not ( w_13305 , w_13308 );
not (  , w_13309 );
and ( w_13308 , w_13309 , \4147_b0 );
or ( \4149_b1 , \4144_b1 , w_13311 );
not ( w_13311 , w_13312 );
and ( \4149_b0 , \4144_b0 , w_13313 );
and ( w_13312 ,  , w_13313 );
buf ( w_13311 , \4148_b1 );
not ( w_13311 , w_13314 );
not (  , w_13315 );
and ( w_13314 , w_13315 , \4148_b0 );
or ( \4150_b1 , \4140_b1 , w_13317 );
not ( w_13317 , w_13318 );
and ( \4150_b0 , \4140_b0 , w_13319 );
and ( w_13318 ,  , w_13319 );
buf ( w_13317 , \4149_b1 );
not ( w_13317 , w_13320 );
not (  , w_13321 );
and ( w_13320 , w_13321 , \4149_b0 );
or ( \4151_b1 , \4138_b1 , w_13323 );
not ( w_13323 , w_13324 );
and ( \4151_b0 , \4138_b0 , w_13325 );
and ( w_13324 ,  , w_13325 );
buf ( w_13323 , \4150_b1 );
not ( w_13323 , w_13326 );
not (  , w_13327 );
and ( w_13326 , w_13327 , \4150_b0 );
or ( \4152_b1 , \4107_b1 , w_13329 );
not ( w_13329 , w_13330 );
and ( \4152_b0 , \4107_b0 , w_13331 );
and ( w_13330 ,  , w_13331 );
buf ( w_13329 , \4151_b1 );
not ( w_13329 , w_13332 );
not (  , w_13333 );
and ( w_13332 , w_13333 , \4151_b0 );
buf ( \4153_b1 , \4105_b1 );
not ( \4153_b1 , w_13334 );
not ( \4153_b0 , w_13335 );
and ( w_13334 , w_13335 , \4105_b0 );
or ( \4154_b1 , \4153_b1 , w_13337 );
not ( w_13337 , w_13338 );
and ( \4154_b0 , \4153_b0 , w_13339 );
and ( w_13338 ,  , w_13339 );
buf ( w_13337 , \4071_b1 );
not ( w_13337 , w_13340 );
not (  , w_13341 );
and ( w_13340 , w_13341 , \4071_b0 );
or ( \4155_b1 , \4152_b1 , w_13343 );
not ( w_13343 , w_13344 );
and ( \4155_b0 , \4152_b0 , w_13345 );
and ( w_13344 ,  , w_13345 );
buf ( w_13343 , \4154_b1 );
not ( w_13343 , w_13346 );
not (  , w_13347 );
and ( w_13346 , w_13347 , \4154_b0 );
buf ( \4156_b1 , \3108_b1 );
buf ( \4156_b0 , \3108_b0 );
or ( \4157_b1 , \4156_b1 , w_13349 );
not ( w_13349 , w_13350 );
and ( \4157_b0 , \4156_b0 , w_13351 );
and ( w_13350 ,  , w_13351 );
buf ( w_13349 , \4046_b1 );
not ( w_13349 , w_13352 );
not (  , w_13353 );
and ( w_13352 , w_13353 , \4046_b0 );
buf ( \4158_b1 , \4136_b1 );
not ( \4158_b1 , w_13354 );
not ( \4158_b0 , w_13355 );
and ( w_13354 , w_13355 , \4136_b0 );
buf ( \4159_b1 , \4149_b1 );
not ( \4159_b1 , w_13356 );
not ( \4159_b0 , w_13357 );
and ( w_13356 , w_13357 , \4149_b0 );
or ( \4160_b1 , \4158_b1 , w_13358 );
or ( \4160_b0 , \4158_b0 , \4159_b0 );
not ( \4159_b0 , w_13359 );
and ( w_13359 , w_13358 , \4159_b1 );
buf ( \4161_b1 , \4044_b1 );
not ( \4161_b1 , w_13360 );
not ( \4161_b0 , w_13361 );
and ( w_13360 , w_13361 , \4044_b0 );
buf ( \4162_b1 , \4110_b1 );
not ( \4162_b1 , w_13362 );
not ( \4162_b0 , w_13363 );
and ( w_13362 , w_13363 , \4110_b0 );
or ( \4163_b1 , \4161_b1 , w_13364 );
or ( \4163_b0 , \4161_b0 , \4162_b0 );
not ( \4162_b0 , w_13365 );
and ( w_13365 , w_13364 , \4162_b1 );
or ( \4164_b1 , \4109_b1 , w_13367 );
not ( w_13367 , w_13368 );
and ( \4164_b0 , \4109_b0 , w_13369 );
and ( w_13368 ,  , w_13369 );
buf ( w_13367 , \4092_b1 );
not ( w_13367 , w_13370 );
not (  , w_13371 );
and ( w_13370 , w_13371 , \4092_b0 );
or ( \4165_b1 , \4163_b1 , w_13373 );
not ( w_13373 , w_13374 );
and ( \4165_b0 , \4163_b0 , w_13375 );
and ( w_13374 ,  , w_13375 );
buf ( w_13373 , \4164_b1 );
not ( w_13373 , w_13376 );
not (  , w_13377 );
and ( w_13376 , w_13377 , \4164_b0 );
or ( \4166_b1 , \4140_b1 , w_13379 );
not ( w_13379 , w_13380 );
and ( \4166_b0 , \4140_b0 , w_13381 );
and ( w_13380 ,  , w_13381 );
buf ( w_13379 , \4165_b1 );
not ( w_13379 , w_13382 );
not (  , w_13383 );
and ( w_13382 , w_13383 , \4165_b0 );
or ( \4167_b1 , \4160_b1 , w_13385 );
not ( w_13385 , w_13386 );
and ( \4167_b0 , \4160_b0 , w_13387 );
and ( w_13386 ,  , w_13387 );
buf ( w_13385 , \4166_b1 );
not ( w_13385 , w_13388 );
not (  , w_13389 );
and ( w_13388 , w_13389 , \4166_b0 );
buf ( \4168_b1 , \4167_b1 );
not ( \4168_b1 , w_13390 );
not ( \4168_b0 , w_13391 );
and ( w_13390 , w_13391 , \4167_b0 );
or ( \4169_b1 , \4157_b1 , \4168_b1 );
xor ( \4169_b0 , \4157_b0 , w_13392 );
not ( w_13392 , w_13393 );
and ( w_13393 , \4168_b1 , \4168_b0 );
buf ( \4170_b1 , \4047_b1 );
not ( \4170_b1 , w_13394 );
not ( \4170_b0 , w_13395 );
and ( w_13394 , w_13395 , \4047_b0 );
buf ( \4171_b1 , \3208_b1 );
buf ( \4171_b0 , \3208_b0 );
buf ( \4172_b1 , \4171_b1 );
buf ( \4172_b0 , \4171_b0 );
buf ( \4173_b1 , \4172_b1 );
not ( \4173_b1 , w_13396 );
not ( \4173_b0 , w_13397 );
and ( w_13396 , w_13397 , \4172_b0 );
buf ( \4174_b1 , \4173_b1 );
not ( \4174_b1 , w_13398 );
not ( \4174_b0 , w_13399 );
and ( w_13398 , w_13399 , \4173_b0 );
or ( \4175_b1 , \4170_b1 , w_13400 );
or ( \4175_b0 , \4170_b0 , \4174_b0 );
not ( \4174_b0 , w_13401 );
and ( w_13401 , w_13400 , \4174_b1 );
buf ( \4176_b1 , \4171_b1 );
not ( \4176_b1 , w_13402 );
not ( \4176_b0 , w_13403 );
and ( w_13402 , w_13403 , \4171_b0 );
buf ( \4177_b1 , \4176_b1 );
not ( \4177_b1 , w_13404 );
not ( \4177_b0 , w_13405 );
and ( w_13404 , w_13405 , \4176_b0 );
buf ( \4178_b1 , \4047_b1 );
not ( \4178_b1 , w_13406 );
not ( \4178_b0 , w_13407 );
and ( w_13406 , w_13407 , \4047_b0 );
or ( \4179_b1 , \4177_b1 , w_13409 );
not ( w_13409 , w_13410 );
and ( \4179_b0 , \4177_b0 , w_13411 );
and ( w_13410 ,  , w_13411 );
buf ( w_13409 , \4178_b1 );
not ( w_13409 , w_13412 );
not (  , w_13413 );
and ( w_13412 , w_13413 , \4178_b0 );
or ( \4180_b1 , \4175_b1 , w_13415 );
not ( w_13415 , w_13416 );
and ( \4180_b0 , \4175_b0 , w_13417 );
and ( w_13416 ,  , w_13417 );
buf ( w_13415 , \4179_b1 );
not ( w_13415 , w_13418 );
not (  , w_13419 );
and ( w_13418 , w_13419 , \4179_b0 );
buf ( \4181_b1 , \4180_b1 );
not ( \4181_b1 , w_13420 );
not ( \4181_b0 , w_13421 );
and ( w_13420 , w_13421 , \4180_b0 );
or ( \4182_b1 , \3487_b1 , \4171_b1 );
not ( \4171_b1 , w_13422 );
and ( \4182_b0 , \3487_b0 , w_13423 );
and ( w_13422 , w_13423 , \4171_b0 );
buf ( \4183_b1 , \3487_b1 );
not ( \4183_b1 , w_13424 );
not ( \4183_b0 , w_13425 );
and ( w_13424 , w_13425 , \3487_b0 );
buf ( \4184_b1 , \4171_b1 );
not ( \4184_b1 , w_13426 );
not ( \4184_b0 , w_13427 );
and ( w_13426 , w_13427 , \4171_b0 );
or ( \4185_b1 , \4183_b1 , \4184_b1 );
not ( \4184_b1 , w_13428 );
and ( \4185_b0 , \4183_b0 , w_13429 );
and ( w_13428 , w_13429 , \4184_b0 );
or ( \4186_b1 , \4182_b1 , w_13431 );
not ( w_13431 , w_13432 );
and ( \4186_b0 , \4182_b0 , w_13433 );
and ( w_13432 ,  , w_13433 );
buf ( w_13431 , \4185_b1 );
not ( w_13431 , w_13434 );
not (  , w_13435 );
and ( w_13434 , w_13435 , \4185_b0 );
buf ( \4187_b1 , \3745_b1 );
not ( \4187_b1 , w_13436 );
not ( \4187_b0 , w_13437 );
and ( w_13436 , w_13437 , \3745_b0 );
or ( \4188_b1 , \4187_b1 , \3487_b1 );
not ( \3487_b1 , w_13438 );
and ( \4188_b0 , \4187_b0 , w_13439 );
and ( w_13438 , w_13439 , \3487_b0 );
buf ( \4189_b1 , \4187_b1 );
not ( \4189_b1 , w_13440 );
not ( \4189_b0 , w_13441 );
and ( w_13440 , w_13441 , \4187_b0 );
buf ( \4190_b1 , \3487_b1 );
not ( \4190_b1 , w_13442 );
not ( \4190_b0 , w_13443 );
and ( w_13442 , w_13443 , \3487_b0 );
or ( \4191_b1 , \4189_b1 , \4190_b1 );
not ( \4190_b1 , w_13444 );
and ( \4191_b0 , \4189_b0 , w_13445 );
and ( w_13444 , w_13445 , \4190_b0 );
or ( \4192_b1 , \4188_b1 , w_13447 );
not ( w_13447 , w_13448 );
and ( \4192_b0 , \4188_b0 , w_13449 );
and ( w_13448 ,  , w_13449 );
buf ( w_13447 , \4191_b1 );
not ( w_13447 , w_13450 );
not (  , w_13451 );
and ( w_13450 , w_13451 , \4191_b0 );
or ( \4193_b1 , \4186_b1 , w_13453 );
not ( w_13453 , w_13454 );
and ( \4193_b0 , \4186_b0 , w_13455 );
and ( w_13454 ,  , w_13455 );
buf ( w_13453 , \4192_b1 );
not ( w_13453 , w_13456 );
not (  , w_13457 );
and ( w_13456 , w_13457 , \4192_b0 );
buf ( \4194_b1 , \4193_b1 );
not ( \4194_b1 , w_13458 );
not ( \4194_b0 , w_13459 );
and ( w_13458 , w_13459 , \4193_b0 );
buf ( \4195_b1 , \4194_b1 );
buf ( \4195_b0 , \4194_b0 );
buf ( \4196_b1 , \4195_b1 );
not ( \4196_b1 , w_13460 );
not ( \4196_b0 , w_13461 );
and ( w_13460 , w_13461 , \4195_b0 );
or ( \4197_b1 , \4181_b1 , w_13462 );
or ( \4197_b0 , \4181_b0 , \4196_b0 );
not ( \4196_b0 , w_13463 );
and ( w_13463 , w_13462 , \4196_b1 );
or ( \4198_b1 , \4116_b1 , \4172_b1 );
not ( \4172_b1 , w_13464 );
and ( \4198_b0 , \4116_b0 , w_13465 );
and ( w_13464 , w_13465 , \4172_b0 );
buf ( \4199_b1 , \4116_b1 );
not ( \4199_b1 , w_13466 );
not ( \4199_b0 , w_13467 );
and ( w_13466 , w_13467 , \4116_b0 );
or ( \4200_b1 , \4199_b1 , \4173_b1 );
not ( \4173_b1 , w_13468 );
and ( \4200_b0 , \4199_b0 , w_13469 );
and ( w_13468 , w_13469 , \4173_b0 );
or ( \4201_b1 , \4198_b1 , w_13471 );
not ( w_13471 , w_13472 );
and ( \4201_b0 , \4198_b0 , w_13473 );
and ( w_13472 ,  , w_13473 );
buf ( w_13471 , \4200_b1 );
not ( w_13471 , w_13474 );
not (  , w_13475 );
and ( w_13474 , w_13475 , \4200_b0 );
buf ( \4202_b1 , \4201_b1 );
not ( \4202_b1 , w_13476 );
not ( \4202_b0 , w_13477 );
and ( w_13476 , w_13477 , \4201_b0 );
buf ( \4203_b1 , \4192_b1 );
buf ( \4203_b0 , \4192_b0 );
buf ( \4204_b1 , \4203_b1 );
not ( \4204_b1 , w_13478 );
not ( \4204_b0 , w_13479 );
and ( w_13478 , w_13479 , \4203_b0 );
buf ( \4205_b1 , \4204_b1 );
buf ( \4205_b0 , \4204_b0 );
or ( \4206_b1 , \4202_b1 , w_13481 );
not ( w_13481 , w_13482 );
and ( \4206_b0 , \4202_b0 , w_13483 );
and ( w_13482 ,  , w_13483 );
buf ( w_13481 , \4205_b1 );
not ( w_13481 , w_13484 );
not (  , w_13485 );
and ( w_13484 , w_13485 , \4205_b0 );
or ( \4207_b1 , \4197_b1 , w_13487 );
not ( w_13487 , w_13488 );
and ( \4207_b0 , \4197_b0 , w_13489 );
and ( w_13488 ,  , w_13489 );
buf ( w_13487 , \4206_b1 );
not ( w_13487 , w_13490 );
not (  , w_13491 );
and ( w_13490 , w_13491 , \4206_b0 );
or ( \4208_b1 , \4169_b1 , w_13492 );
xor ( \4208_b0 , \4169_b0 , w_13494 );
not ( w_13494 , w_13495 );
and ( w_13495 , w_13492 , w_13493 );
buf ( w_13492 , \4207_b1 );
not ( w_13492 , w_13496 );
not ( w_13493 , w_13497 );
and ( w_13496 , w_13497 , \4207_b0 );
or ( \4209_b1 , \4155_b1 , \4208_b1 );
xor ( \4209_b0 , \4155_b0 , w_13498 );
not ( w_13498 , w_13499 );
and ( w_13499 , \4208_b1 , \4208_b0 );
buf ( \4210_b1 , \4043_b1 );
not ( \4210_b1 , w_13500 );
not ( \4210_b0 , w_13501 );
and ( w_13500 , w_13501 , \4043_b0 );
buf ( \4211_b1 , \3577_b1 );
not ( \4211_b1 , w_13502 );
not ( \4211_b0 , w_13503 );
and ( w_13502 , w_13503 , \3577_b0 );
buf ( \4212_b1 , \4211_b1 );
buf ( \4212_b0 , \4211_b0 );
buf ( \4213_b1 , \4212_b1 );
buf ( \4213_b0 , \4212_b0 );
buf ( \4214_b1 , \4213_b1 );
not ( \4214_b1 , w_13504 );
not ( \4214_b0 , w_13505 );
and ( w_13504 , w_13505 , \4213_b0 );
or ( \4215_b1 , \4210_b1 , w_13506 );
or ( \4215_b0 , \4210_b0 , \4214_b0 );
not ( \4214_b0 , w_13507 );
and ( w_13507 , w_13506 , \4214_b1 );
buf ( \4216_b1 , \4212_b1 );
not ( \4216_b1 , w_13508 );
not ( \4216_b0 , w_13509 );
and ( w_13508 , w_13509 , \4212_b0 );
buf ( \4217_b1 , \4043_b1 );
not ( \4217_b1 , w_13510 );
not ( \4217_b0 , w_13511 );
and ( w_13510 , w_13511 , \4043_b0 );
or ( \4218_b1 , \4216_b1 , w_13513 );
not ( w_13513 , w_13514 );
and ( \4218_b0 , \4216_b0 , w_13515 );
and ( w_13514 ,  , w_13515 );
buf ( w_13513 , \4217_b1 );
not ( w_13513 , w_13516 );
not (  , w_13517 );
and ( w_13516 , w_13517 , \4217_b0 );
or ( \4219_b1 , \4215_b1 , w_13519 );
not ( w_13519 , w_13520 );
and ( \4219_b0 , \4215_b0 , w_13521 );
and ( w_13520 ,  , w_13521 );
buf ( w_13519 , \4218_b1 );
not ( w_13519 , w_13522 );
not (  , w_13523 );
and ( w_13522 , w_13523 , \4218_b0 );
buf ( \4220_b1 , \4219_b1 );
not ( \4220_b1 , w_13524 );
not ( \4220_b0 , w_13525 );
and ( w_13524 , w_13525 , \4219_b0 );
or ( \4221_b1 , \3208_b1 , \3818_b1 );
xor ( \4221_b0 , \3208_b0 , w_13526 );
not ( w_13526 , w_13527 );
and ( w_13527 , \3818_b1 , \3818_b0 );
buf ( \4222_b1 , \4221_b1 );
not ( \4222_b1 , w_13528 );
not ( \4222_b0 , w_13529 );
and ( w_13528 , w_13529 , \4221_b0 );
buf ( \4223_b1 , \3577_b1 );
not ( \4223_b1 , w_13530 );
not ( \4223_b0 , w_13531 );
and ( w_13530 , w_13531 , \3577_b0 );
buf ( \4224_b1 , \3818_b1 );
not ( \4224_b1 , w_13532 );
not ( \4224_b0 , w_13533 );
and ( w_13532 , w_13533 , \3818_b0 );
buf ( \4225_b1 , \4224_b1 );
not ( \4225_b1 , w_13534 );
not ( \4225_b0 , w_13535 );
and ( w_13534 , w_13535 , \4224_b0 );
or ( \4226_b1 , \4223_b1 , w_13536 );
or ( \4226_b0 , \4223_b0 , \4225_b0 );
not ( \4225_b0 , w_13537 );
and ( w_13537 , w_13536 , \4225_b1 );
buf ( \4227_b1 , \3577_b1 );
not ( \4227_b1 , w_13538 );
not ( \4227_b0 , w_13539 );
and ( w_13538 , w_13539 , \3577_b0 );
or ( \4228_b1 , \4227_b1 , w_13541 );
not ( w_13541 , w_13542 );
and ( \4228_b0 , \4227_b0 , w_13543 );
and ( w_13542 ,  , w_13543 );
buf ( w_13541 , \3818_b1 );
not ( w_13541 , w_13544 );
not (  , w_13545 );
and ( w_13544 , w_13545 , \3818_b0 );
or ( \4229_b1 , \4226_b1 , w_13547 );
not ( w_13547 , w_13548 );
and ( \4229_b0 , \4226_b0 , w_13549 );
and ( w_13548 ,  , w_13549 );
buf ( w_13547 , \4228_b1 );
not ( w_13547 , w_13550 );
not (  , w_13551 );
and ( w_13550 , w_13551 , \4228_b0 );
or ( \4230_b1 , \4222_b1 , w_13553 );
not ( w_13553 , w_13554 );
and ( \4230_b0 , \4222_b0 , w_13555 );
and ( w_13554 ,  , w_13555 );
buf ( w_13553 , \4229_b1 );
not ( w_13553 , w_13556 );
not (  , w_13557 );
and ( w_13556 , w_13557 , \4229_b0 );
buf ( \4231_b1 , \4230_b1 );
not ( \4231_b1 , w_13558 );
not ( \4231_b0 , w_13559 );
and ( w_13558 , w_13559 , \4230_b0 );
buf ( \4232_b1 , \4231_b1 );
not ( \4232_b1 , w_13560 );
not ( \4232_b0 , w_13561 );
and ( w_13560 , w_13561 , \4231_b0 );
or ( \4233_b1 , \4220_b1 , w_13562 );
or ( \4233_b0 , \4220_b0 , \4232_b0 );
not ( \4232_b0 , w_13563 );
and ( w_13563 , w_13562 , \4232_b1 );
buf ( \4234_b1 , \4221_b1 );
buf ( \4234_b0 , \4221_b0 );
buf ( \4235_b1 , \4041_b1 );
not ( \4235_b1 , w_13564 );
not ( \4235_b0 , w_13565 );
and ( w_13564 , w_13565 , \4041_b0 );
buf ( \4236_b1 , \4213_b1 );
not ( \4236_b1 , w_13566 );
not ( \4236_b0 , w_13567 );
and ( w_13566 , w_13567 , \4213_b0 );
or ( \4237_b1 , \4235_b1 , w_13568 );
or ( \4237_b0 , \4235_b0 , \4236_b0 );
not ( \4236_b0 , w_13569 );
and ( w_13569 , w_13568 , \4236_b1 );
buf ( \4238_b1 , \4041_b1 );
not ( \4238_b1 , w_13570 );
not ( \4238_b0 , w_13571 );
and ( w_13570 , w_13571 , \4041_b0 );
or ( \4239_b1 , \4216_b1 , w_13573 );
not ( w_13573 , w_13574 );
and ( \4239_b0 , \4216_b0 , w_13575 );
and ( w_13574 ,  , w_13575 );
buf ( w_13573 , \4238_b1 );
not ( w_13573 , w_13576 );
not (  , w_13577 );
and ( w_13576 , w_13577 , \4238_b0 );
or ( \4240_b1 , \4237_b1 , w_13579 );
not ( w_13579 , w_13580 );
and ( \4240_b0 , \4237_b0 , w_13581 );
and ( w_13580 ,  , w_13581 );
buf ( w_13579 , \4239_b1 );
not ( w_13579 , w_13582 );
not (  , w_13583 );
and ( w_13582 , w_13583 , \4239_b0 );
or ( \4241_b1 , \4234_b1 , w_13585 );
not ( w_13585 , w_13586 );
and ( \4241_b0 , \4234_b0 , w_13587 );
and ( w_13586 ,  , w_13587 );
buf ( w_13585 , \4240_b1 );
not ( w_13585 , w_13588 );
not (  , w_13589 );
and ( w_13588 , w_13589 , \4240_b0 );
or ( \4242_b1 , \4233_b1 , w_13591 );
not ( w_13591 , w_13592 );
and ( \4242_b0 , \4233_b0 , w_13593 );
and ( w_13592 ,  , w_13593 );
buf ( w_13591 , \4241_b1 );
not ( w_13591 , w_13594 );
not (  , w_13595 );
and ( w_13594 , w_13595 , \4241_b0 );
buf ( \4243_b1 , \4242_b1 );
not ( \4243_b1 , w_13596 );
not ( \4243_b0 , w_13597 );
and ( w_13596 , w_13597 , \4242_b0 );
buf ( \4244_b1 , \3366_b1 );
not ( \4244_b1 , w_13598 );
not ( \4244_b0 , w_13599 );
and ( w_13598 , w_13599 , \3366_b0 );
buf ( \4245_b1 , \4244_b1 );
not ( \4245_b1 , w_13600 );
not ( \4245_b0 , w_13601 );
and ( w_13600 , w_13601 , \4244_b0 );
buf ( \4246_b1 , \4245_b1 );
not ( \4246_b1 , w_13602 );
not ( \4246_b0 , w_13603 );
and ( w_13602 , w_13603 , \4245_b0 );
buf ( \4247_b1 , \3108_b1 );
not ( \4247_b1 , w_13604 );
not ( \4247_b0 , w_13605 );
and ( w_13604 , w_13605 , \3108_b0 );
buf ( \4248_b1 , \4247_b1 );
not ( \4248_b1 , w_13606 );
not ( \4248_b0 , w_13607 );
and ( w_13606 , w_13607 , \4247_b0 );
or ( \4249_b1 , \4246_b1 , w_13608 );
or ( \4249_b0 , \4246_b0 , \4248_b0 );
not ( \4248_b0 , w_13609 );
and ( w_13609 , w_13608 , \4248_b1 );
or ( \4250_b1 , \3108_b1 , w_13611 );
not ( w_13611 , w_13612 );
and ( \4250_b0 , \3108_b0 , w_13613 );
and ( w_13612 ,  , w_13613 );
buf ( w_13611 , \4244_b1 );
not ( w_13611 , w_13614 );
not (  , w_13615 );
and ( w_13614 , w_13615 , \4244_b0 );
or ( \4251_b1 , \4249_b1 , w_13617 );
not ( w_13617 , w_13618 );
and ( \4251_b0 , \4249_b0 , w_13619 );
and ( w_13618 ,  , w_13619 );
buf ( w_13617 , \4250_b1 );
not ( w_13617 , w_13620 );
not (  , w_13621 );
and ( w_13620 , w_13621 , \4250_b0 );
or ( \4252_b1 , \3577_b1 , w_13622 );
xor ( \4252_b0 , \3577_b0 , w_13624 );
not ( w_13624 , w_13625 );
and ( w_13625 , w_13622 , w_13623 );
buf ( w_13622 , \3366_b1 );
not ( w_13622 , w_13626 );
not ( w_13623 , w_13627 );
and ( w_13626 , w_13627 , \3366_b0 );
or ( \4253_b1 , \4251_b1 , \4252_b1 );
not ( \4252_b1 , w_13628 );
and ( \4253_b0 , \4251_b0 , w_13629 );
and ( w_13628 , w_13629 , \4252_b0 );
buf ( \4254_b1 , \4253_b1 );
not ( \4254_b1 , w_13630 );
not ( \4254_b0 , w_13631 );
and ( w_13630 , w_13631 , \4253_b0 );
buf ( \4255_b1 , \4254_b1 );
not ( \4255_b1 , w_13632 );
not ( \4255_b0 , w_13633 );
and ( w_13632 , w_13633 , \4254_b0 );
buf ( \4256_b1 , \4046_b1 );
not ( \4256_b1 , w_13634 );
not ( \4256_b0 , w_13635 );
and ( w_13634 , w_13635 , \4046_b0 );
buf ( \4257_b1 , \4256_b1 );
not ( \4257_b1 , w_13636 );
not ( \4257_b0 , w_13637 );
and ( w_13636 , w_13637 , \4256_b0 );
buf ( \4258_b1 , \4156_b1 );
not ( \4258_b1 , w_13638 );
not ( \4258_b0 , w_13639 );
and ( w_13638 , w_13639 , \4156_b0 );
or ( \4259_b1 , \4257_b1 , w_13640 );
or ( \4259_b0 , \4257_b0 , \4258_b0 );
not ( \4258_b0 , w_13641 );
and ( w_13641 , w_13640 , \4258_b1 );
buf ( \4260_b1 , \3108_b1 );
not ( \4260_b1 , w_13642 );
not ( \4260_b0 , w_13643 );
and ( w_13642 , w_13643 , \3108_b0 );
or ( \4261_b1 , \4260_b1 , w_13645 );
not ( w_13645 , w_13646 );
and ( \4261_b0 , \4260_b0 , w_13647 );
and ( w_13646 ,  , w_13647 );
buf ( w_13645 , \4046_b1 );
not ( w_13645 , w_13648 );
not (  , w_13649 );
and ( w_13648 , w_13649 , \4046_b0 );
or ( \4262_b1 , \4259_b1 , w_13651 );
not ( w_13651 , w_13652 );
and ( \4262_b0 , \4259_b0 , w_13653 );
and ( w_13652 ,  , w_13653 );
buf ( w_13651 , \4261_b1 );
not ( w_13651 , w_13654 );
not (  , w_13655 );
and ( w_13654 , w_13655 , \4261_b0 );
buf ( \4263_b1 , \4262_b1 );
not ( \4263_b1 , w_13656 );
not ( \4263_b0 , w_13657 );
and ( w_13656 , w_13657 , \4262_b0 );
buf ( \4264_b1 , \4263_b1 );
not ( \4264_b1 , w_13658 );
not ( \4264_b0 , w_13659 );
and ( w_13658 , w_13659 , \4263_b0 );
or ( \4265_b1 , \4255_b1 , \4264_b1 );
not ( \4264_b1 , w_13660 );
and ( \4265_b0 , \4255_b0 , w_13661 );
and ( w_13660 , w_13661 , \4264_b0 );
buf ( \4266_b1 , \4011_b1 );
not ( \4266_b1 , w_13662 );
not ( \4266_b0 , w_13663 );
and ( w_13662 , w_13663 , \4011_b0 );
buf ( \4267_b1 , \4156_b1 );
not ( \4267_b1 , w_13664 );
not ( \4267_b0 , w_13665 );
and ( w_13664 , w_13665 , \4156_b0 );
buf ( \4268_b1 , \4267_b1 );
not ( \4268_b1 , w_13666 );
not ( \4268_b0 , w_13667 );
and ( w_13666 , w_13667 , \4267_b0 );
or ( \4269_b1 , \4266_b1 , w_13668 );
or ( \4269_b0 , \4266_b0 , \4268_b0 );
not ( \4268_b0 , w_13669 );
and ( w_13669 , w_13668 , \4268_b1 );
buf ( \4270_b1 , \4011_b1 );
not ( \4270_b1 , w_13670 );
not ( \4270_b0 , w_13671 );
and ( w_13670 , w_13671 , \4011_b0 );
or ( \4271_b1 , \4156_b1 , w_13673 );
not ( w_13673 , w_13674 );
and ( \4271_b0 , \4156_b0 , w_13675 );
and ( w_13674 ,  , w_13675 );
buf ( w_13673 , \4270_b1 );
not ( w_13673 , w_13676 );
not (  , w_13677 );
and ( w_13676 , w_13677 , \4270_b0 );
or ( \4272_b1 , \4269_b1 , w_13679 );
not ( w_13679 , w_13680 );
and ( \4272_b0 , \4269_b0 , w_13681 );
and ( w_13680 ,  , w_13681 );
buf ( w_13679 , \4271_b1 );
not ( w_13679 , w_13682 );
not (  , w_13683 );
and ( w_13682 , w_13683 , \4271_b0 );
buf ( \4273_b1 , \4252_b1 );
not ( \4273_b1 , w_13684 );
not ( \4273_b0 , w_13685 );
and ( w_13684 , w_13685 , \4252_b0 );
buf ( \4274_b1 , \4273_b1 );
buf ( \4274_b0 , \4273_b0 );
or ( \4275_b1 , \4272_b1 , \4274_b1 );
not ( \4274_b1 , w_13686 );
and ( \4275_b0 , \4272_b0 , w_13687 );
and ( w_13686 , w_13687 , \4274_b0 );
or ( \4276_b1 , \4265_b1 , w_13689 );
not ( w_13689 , w_13690 );
and ( \4276_b0 , \4265_b0 , w_13691 );
and ( w_13690 ,  , w_13691 );
buf ( w_13689 , \4275_b1 );
not ( w_13689 , w_13692 );
not (  , w_13693 );
and ( w_13692 , w_13693 , \4275_b0 );
buf ( \4277_b1 , \4276_b1 );
not ( \4277_b1 , w_13694 );
not ( \4277_b0 , w_13695 );
and ( w_13694 , w_13695 , \4276_b0 );
buf ( \4278_b1 , \4277_b1 );
not ( \4278_b1 , w_13696 );
not ( \4278_b0 , w_13697 );
and ( w_13696 , w_13697 , \4277_b0 );
or ( \4279_b1 , \4243_b1 , w_13698 );
or ( \4279_b0 , \4243_b0 , \4278_b0 );
not ( \4278_b0 , w_13699 );
and ( w_13699 , w_13698 , \4278_b1 );
or ( \4280_b1 , \4277_b1 , w_13700 );
or ( \4280_b0 , \4277_b0 , \4242_b0 );
not ( \4242_b0 , w_13701 );
and ( w_13701 , w_13700 , \4242_b1 );
buf ( \4281_b1 , \4045_b1 );
not ( \4281_b1 , w_13702 );
not ( \4281_b0 , w_13703 );
and ( w_13702 , w_13703 , \4045_b0 );
buf ( \4282_b1 , \4176_b1 );
not ( \4282_b1 , w_13704 );
not ( \4282_b0 , w_13705 );
and ( w_13704 , w_13705 , \4176_b0 );
or ( \4283_b1 , \4281_b1 , w_13706 );
or ( \4283_b0 , \4281_b0 , \4282_b0 );
not ( \4282_b0 , w_13707 );
and ( w_13707 , w_13706 , \4282_b1 );
buf ( \4284_b1 , \4171_b1 );
not ( \4284_b1 , w_13708 );
not ( \4284_b0 , w_13709 );
and ( w_13708 , w_13709 , \4171_b0 );
buf ( \4285_b1 , \4284_b1 );
not ( \4285_b1 , w_13710 );
not ( \4285_b0 , w_13711 );
and ( w_13710 , w_13711 , \4284_b0 );
buf ( \4286_b1 , \4045_b1 );
not ( \4286_b1 , w_13712 );
not ( \4286_b0 , w_13713 );
and ( w_13712 , w_13713 , \4045_b0 );
or ( \4287_b1 , \4285_b1 , w_13715 );
not ( w_13715 , w_13716 );
and ( \4287_b0 , \4285_b0 , w_13717 );
and ( w_13716 ,  , w_13717 );
buf ( w_13715 , \4286_b1 );
not ( w_13715 , w_13718 );
not (  , w_13719 );
and ( w_13718 , w_13719 , \4286_b0 );
or ( \4288_b1 , \4283_b1 , w_13721 );
not ( w_13721 , w_13722 );
and ( \4288_b0 , \4283_b0 , w_13723 );
and ( w_13722 ,  , w_13723 );
buf ( w_13721 , \4287_b1 );
not ( w_13721 , w_13724 );
not (  , w_13725 );
and ( w_13724 , w_13725 , \4287_b0 );
buf ( \4289_b1 , \4288_b1 );
not ( \4289_b1 , w_13726 );
not ( \4289_b0 , w_13727 );
and ( w_13726 , w_13727 , \4288_b0 );
buf ( \4290_b1 , \4195_b1 );
not ( \4290_b1 , w_13728 );
not ( \4290_b0 , w_13729 );
and ( w_13728 , w_13729 , \4195_b0 );
or ( \4291_b1 , \4289_b1 , w_13730 );
or ( \4291_b0 , \4289_b0 , \4290_b0 );
not ( \4290_b0 , w_13731 );
and ( w_13731 , w_13730 , \4290_b1 );
or ( \4292_b1 , \4205_b1 , w_13733 );
not ( w_13733 , w_13734 );
and ( \4292_b0 , \4205_b0 , w_13735 );
and ( w_13734 ,  , w_13735 );
buf ( w_13733 , \4180_b1 );
not ( w_13733 , w_13736 );
not (  , w_13737 );
and ( w_13736 , w_13737 , \4180_b0 );
or ( \4293_b1 , \4291_b1 , w_13739 );
not ( w_13739 , w_13740 );
and ( \4293_b0 , \4291_b0 , w_13741 );
and ( w_13740 ,  , w_13741 );
buf ( w_13739 , \4292_b1 );
not ( w_13739 , w_13742 );
not (  , w_13743 );
and ( w_13742 , w_13743 , \4292_b0 );
or ( \4294_b1 , \4280_b1 , w_13745 );
not ( w_13745 , w_13746 );
and ( \4294_b0 , \4280_b0 , w_13747 );
and ( w_13746 ,  , w_13747 );
buf ( w_13745 , \4293_b1 );
not ( w_13745 , w_13748 );
not (  , w_13749 );
and ( w_13748 , w_13749 , \4293_b0 );
or ( \4295_b1 , \4279_b1 , w_13751 );
not ( w_13751 , w_13752 );
and ( \4295_b0 , \4279_b0 , w_13753 );
and ( w_13752 ,  , w_13753 );
buf ( w_13751 , \4294_b1 );
not ( w_13751 , w_13754 );
not (  , w_13755 );
and ( w_13754 , w_13755 , \4294_b0 );
or ( \4296_b1 , \4209_b1 , \4295_b1 );
not ( \4295_b1 , w_13756 );
and ( \4296_b0 , \4209_b0 , w_13757 );
and ( w_13756 , w_13757 , \4295_b0 );
or ( \4297_b1 , \4155_b1 , \4208_b1 );
not ( \4208_b1 , w_13758 );
and ( \4297_b0 , \4155_b0 , w_13759 );
and ( w_13758 , w_13759 , \4208_b0 );
or ( \4298_b1 , \4296_b1 , w_13760 );
or ( \4298_b0 , \4296_b0 , \4297_b0 );
not ( \4297_b0 , w_13761 );
and ( w_13761 , w_13760 , \4297_b1 );
buf ( \4299_b1 , \4157_b1 );
not ( \4299_b1 , w_13762 );
not ( \4299_b0 , w_13763 );
and ( w_13762 , w_13763 , \4157_b0 );
buf ( \4300_b1 , \4167_b1 );
not ( \4300_b1 , w_13764 );
not ( \4300_b0 , w_13765 );
and ( w_13764 , w_13765 , \4167_b0 );
or ( \4301_b1 , \4299_b1 , w_13766 );
or ( \4301_b0 , \4299_b0 , \4300_b0 );
not ( \4300_b0 , w_13767 );
and ( w_13767 , w_13766 , \4300_b1 );
or ( \4302_b1 , \4301_b1 , w_13769 );
not ( w_13769 , w_13770 );
and ( \4302_b0 , \4301_b0 , w_13771 );
and ( w_13770 ,  , w_13771 );
buf ( w_13769 , \4207_b1 );
not ( w_13769 , w_13772 );
not (  , w_13773 );
and ( w_13772 , w_13773 , \4207_b0 );
buf ( \4303_b1 , \4157_b1 );
not ( \4303_b1 , w_13774 );
not ( \4303_b0 , w_13775 );
and ( w_13774 , w_13775 , \4157_b0 );
or ( \4304_b1 , \4303_b1 , w_13777 );
not ( w_13777 , w_13778 );
and ( \4304_b0 , \4303_b0 , w_13779 );
and ( w_13778 ,  , w_13779 );
buf ( w_13777 , \4168_b1 );
not ( w_13777 , w_13780 );
not (  , w_13781 );
and ( w_13780 , w_13781 , \4168_b0 );
or ( \4305_b1 , \4302_b1 , w_13783 );
not ( w_13783 , w_13784 );
and ( \4305_b0 , \4302_b0 , w_13785 );
and ( w_13784 ,  , w_13785 );
buf ( w_13783 , \4304_b1 );
not ( w_13783 , w_13786 );
not (  , w_13787 );
and ( w_13786 , w_13787 , \4304_b0 );
buf ( \4306_b1 , \4305_b1 );
not ( \4306_b1 , w_13788 );
not ( \4306_b0 , w_13789 );
and ( w_13788 , w_13789 , \4305_b0 );
or ( \4307_b1 , \4156_b1 , \4011_b1 );
not ( \4011_b1 , w_13790 );
and ( \4307_b0 , \4156_b0 , w_13791 );
and ( w_13790 , w_13791 , \4011_b0 );
buf ( \4308_b1 , \4260_b1 );
not ( \4308_b1 , w_13792 );
not ( \4308_b0 , w_13793 );
and ( w_13792 , w_13793 , \4260_b0 );
or ( \4309_b1 , \4043_b1 , \4308_b1 );
xor ( \4309_b0 , \4043_b0 , w_13794 );
not ( w_13794 , w_13795 );
and ( w_13795 , \4308_b1 , \4308_b0 );
buf ( \4310_b1 , \4309_b1 );
not ( \4310_b1 , w_13796 );
not ( \4310_b0 , w_13797 );
and ( w_13796 , w_13797 , \4309_b0 );
buf ( \4311_b1 , \4253_b1 );
not ( \4311_b1 , w_13798 );
not ( \4311_b0 , w_13799 );
and ( w_13798 , w_13799 , \4253_b0 );
or ( \4312_b1 , \4310_b1 , w_13800 );
or ( \4312_b0 , \4310_b0 , \4311_b0 );
not ( \4311_b0 , w_13801 );
and ( w_13801 , w_13800 , \4311_b1 );
or ( \4313_b1 , \4041_b1 , \4156_b1 );
xor ( \4313_b0 , \4041_b0 , w_13802 );
not ( w_13802 , w_13803 );
and ( w_13803 , \4156_b1 , \4156_b0 );
or ( \4314_b1 , \4313_b1 , w_13805 );
not ( w_13805 , w_13806 );
and ( \4314_b0 , \4313_b0 , w_13807 );
and ( w_13806 ,  , w_13807 );
buf ( w_13805 , \4274_b1 );
not ( w_13805 , w_13808 );
not (  , w_13809 );
and ( w_13808 , w_13809 , \4274_b0 );
or ( \4315_b1 , \4312_b1 , w_13811 );
not ( w_13811 , w_13812 );
and ( \4315_b0 , \4312_b0 , w_13813 );
and ( w_13812 ,  , w_13813 );
buf ( w_13811 , \4314_b1 );
not ( w_13811 , w_13814 );
not (  , w_13815 );
and ( w_13814 , w_13815 , \4314_b0 );
or ( \4316_b1 , \4307_b1 , \4315_b1 );
xor ( \4316_b0 , \4307_b0 , w_13816 );
not ( w_13816 , w_13817 );
and ( w_13817 , \4315_b1 , \4315_b0 );
buf ( \4317_b1 , \4195_b1 );
not ( \4317_b1 , w_13818 );
not ( \4317_b0 , w_13819 );
and ( w_13818 , w_13819 , \4195_b0 );
or ( \4318_b1 , \4317_b1 , w_13820 );
or ( \4318_b0 , \4317_b0 , \4201_b0 );
not ( \4201_b0 , w_13821 );
and ( w_13821 , w_13820 , \4201_b1 );
buf ( \4319_b1 , \4205_b1 );
not ( \4319_b1 , w_13822 );
not ( \4319_b0 , w_13823 );
and ( w_13822 , w_13823 , \4205_b0 );
or ( \4320_b1 , \4147_b1 , \4172_b1 );
not ( \4172_b1 , w_13824 );
and ( \4320_b0 , \4147_b0 , w_13825 );
and ( w_13824 , w_13825 , \4172_b0 );
buf ( \4321_b1 , \4147_b1 );
not ( \4321_b1 , w_13826 );
not ( \4321_b0 , w_13827 );
and ( w_13826 , w_13827 , \4147_b0 );
or ( \4322_b1 , \4321_b1 , \4173_b1 );
not ( \4173_b1 , w_13828 );
and ( \4322_b0 , \4321_b0 , w_13829 );
and ( w_13828 , w_13829 , \4173_b0 );
or ( \4323_b1 , \4320_b1 , w_13831 );
not ( w_13831 , w_13832 );
and ( \4323_b0 , \4320_b0 , w_13833 );
and ( w_13832 ,  , w_13833 );
buf ( w_13831 , \4322_b1 );
not ( w_13831 , w_13834 );
not (  , w_13835 );
and ( w_13834 , w_13835 , \4322_b0 );
or ( \4324_b1 , \4319_b1 , w_13836 );
or ( \4324_b0 , \4319_b0 , \4323_b0 );
not ( \4323_b0 , w_13837 );
and ( w_13837 , w_13836 , \4323_b1 );
or ( \4325_b1 , \4318_b1 , w_13839 );
not ( w_13839 , w_13840 );
and ( \4325_b0 , \4318_b0 , w_13841 );
and ( w_13840 ,  , w_13841 );
buf ( w_13839 , \4324_b1 );
not ( w_13839 , w_13842 );
not (  , w_13843 );
and ( w_13842 , w_13843 , \4324_b0 );
or ( \4326_b1 , \4316_b1 , \4325_b1 );
xor ( \4326_b0 , \4316_b0 , w_13844 );
not ( w_13844 , w_13845 );
and ( w_13845 , \4325_b1 , \4325_b0 );
or ( \4327_b1 , \4306_b1 , \4326_b1 );
xor ( \4327_b0 , \4306_b0 , w_13846 );
not ( w_13846 , w_13847 );
and ( w_13847 , \4326_b1 , \4326_b0 );
buf ( \4328_b1 , \4101_b1 );
not ( \4328_b1 , w_13848 );
not ( \4328_b0 , w_13849 );
and ( w_13848 , w_13849 , \4101_b0 );
buf ( \4329_b1 , \4086_b1 );
not ( \4329_b1 , w_13850 );
not ( \4329_b0 , w_13851 );
and ( w_13850 , w_13851 , \4086_b0 );
or ( \4330_b1 , \4328_b1 , w_13852 );
or ( \4330_b0 , \4328_b0 , \4329_b0 );
not ( \4329_b0 , w_13853 );
and ( w_13853 , w_13852 , \4329_b1 );
buf ( \4331_b1 , \4103_b1 );
not ( \4331_b1 , w_13854 );
not ( \4331_b0 , w_13855 );
and ( w_13854 , w_13855 , \4103_b0 );
or ( \4332_b1 , \4331_b1 , w_13857 );
not ( w_13857 , w_13858 );
and ( \4332_b0 , \4331_b0 , w_13859 );
and ( w_13858 ,  , w_13859 );
buf ( w_13857 , \4088_b1 );
not ( w_13857 , w_13860 );
not (  , w_13861 );
and ( w_13860 , w_13861 , \4088_b0 );
or ( \4333_b1 , \4330_b1 , w_13863 );
not ( w_13863 , w_13864 );
and ( \4333_b0 , \4330_b0 , w_13865 );
and ( w_13864 ,  , w_13865 );
buf ( w_13863 , \4332_b1 );
not ( w_13863 , w_13866 );
not (  , w_13867 );
and ( w_13866 , w_13867 , \4332_b0 );
buf ( \4334_b1 , \4333_b1 );
not ( \4334_b1 , w_13868 );
not ( \4334_b0 , w_13869 );
and ( w_13868 , w_13869 , \4333_b0 );
buf ( \4335_b1 , \4240_b1 );
not ( \4335_b1 , w_13870 );
not ( \4335_b0 , w_13871 );
and ( w_13870 , w_13871 , \4240_b0 );
buf ( \4336_b1 , \4231_b1 );
not ( \4336_b1 , w_13872 );
not ( \4336_b0 , w_13873 );
and ( w_13872 , w_13873 , \4231_b0 );
or ( \4337_b1 , \4335_b1 , w_13874 );
or ( \4337_b0 , \4335_b0 , \4336_b0 );
not ( \4336_b0 , w_13875 );
and ( w_13875 , w_13874 , \4336_b1 );
buf ( \4338_b1 , \4045_b1 );
not ( \4338_b1 , w_13876 );
not ( \4338_b0 , w_13877 );
and ( w_13876 , w_13877 , \4045_b0 );
buf ( \4339_b1 , \4212_b1 );
not ( \4339_b1 , w_13878 );
not ( \4339_b0 , w_13879 );
and ( w_13878 , w_13879 , \4212_b0 );
or ( \4340_b1 , \4338_b1 , w_13880 );
or ( \4340_b0 , \4338_b0 , \4339_b0 );
not ( \4339_b0 , w_13881 );
and ( w_13881 , w_13880 , \4339_b1 );
or ( \4341_b1 , \4216_b1 , w_13883 );
not ( w_13883 , w_13884 );
and ( \4341_b0 , \4216_b0 , w_13885 );
and ( w_13884 ,  , w_13885 );
buf ( w_13883 , \4286_b1 );
not ( w_13883 , w_13886 );
not (  , w_13887 );
and ( w_13886 , w_13887 , \4286_b0 );
or ( \4342_b1 , \4340_b1 , w_13889 );
not ( w_13889 , w_13890 );
and ( \4342_b0 , \4340_b0 , w_13891 );
and ( w_13890 ,  , w_13891 );
buf ( w_13889 , \4341_b1 );
not ( w_13889 , w_13892 );
not (  , w_13893 );
and ( w_13892 , w_13893 , \4341_b0 );
or ( \4343_b1 , \4234_b1 , w_13895 );
not ( w_13895 , w_13896 );
and ( \4343_b0 , \4234_b0 , w_13897 );
and ( w_13896 ,  , w_13897 );
buf ( w_13895 , \4342_b1 );
not ( w_13895 , w_13898 );
not (  , w_13899 );
and ( w_13898 , w_13899 , \4342_b0 );
or ( \4344_b1 , \4337_b1 , w_13901 );
not ( w_13901 , w_13902 );
and ( \4344_b0 , \4337_b0 , w_13903 );
and ( w_13902 ,  , w_13903 );
buf ( w_13901 , \4343_b1 );
not ( w_13901 , w_13904 );
not (  , w_13905 );
and ( w_13904 , w_13905 , \4343_b0 );
buf ( \4345_b1 , \4344_b1 );
not ( \4345_b1 , w_13906 );
not ( \4345_b0 , w_13907 );
and ( w_13906 , w_13907 , \4344_b0 );
or ( \4346_b1 , \4334_b1 , w_13908 );
or ( \4346_b0 , \4334_b0 , \4345_b0 );
not ( \4345_b0 , w_13909 );
and ( w_13909 , w_13908 , \4345_b1 );
or ( \4347_b1 , \4344_b1 , w_13910 );
or ( \4347_b0 , \4344_b0 , \4333_b0 );
not ( \4333_b0 , w_13911 );
and ( w_13911 , w_13910 , \4333_b1 );
buf ( \4348_b1 , \4272_b1 );
not ( \4348_b1 , w_13912 );
not ( \4348_b0 , w_13913 );
and ( w_13912 , w_13913 , \4272_b0 );
buf ( \4349_b1 , \4253_b1 );
not ( \4349_b1 , w_13914 );
not ( \4349_b0 , w_13915 );
and ( w_13914 , w_13915 , \4253_b0 );
or ( \4350_b1 , \4348_b1 , w_13916 );
or ( \4350_b0 , \4348_b0 , \4349_b0 );
not ( \4349_b0 , w_13917 );
and ( w_13917 , w_13916 , \4349_b1 );
or ( \4351_b1 , \4274_b1 , w_13919 );
not ( w_13919 , w_13920 );
and ( \4351_b0 , \4274_b0 , w_13921 );
and ( w_13920 ,  , w_13921 );
buf ( w_13919 , \4309_b1 );
not ( w_13919 , w_13922 );
not (  , w_13923 );
and ( w_13922 , w_13923 , \4309_b0 );
or ( \4352_b1 , \4350_b1 , w_13925 );
not ( w_13925 , w_13926 );
and ( \4352_b0 , \4350_b0 , w_13927 );
and ( w_13926 ,  , w_13927 );
buf ( w_13925 , \4351_b1 );
not ( w_13925 , w_13928 );
not (  , w_13929 );
and ( w_13928 , w_13929 , \4351_b0 );
or ( \4353_b1 , \4347_b1 , w_13931 );
not ( w_13931 , w_13932 );
and ( \4353_b0 , \4347_b0 , w_13933 );
and ( w_13932 ,  , w_13933 );
buf ( w_13931 , \4352_b1 );
not ( w_13931 , w_13934 );
not (  , w_13935 );
and ( w_13934 , w_13935 , \4352_b0 );
or ( \4354_b1 , \4346_b1 , w_13937 );
not ( w_13937 , w_13938 );
and ( \4354_b0 , \4346_b0 , w_13939 );
and ( w_13938 ,  , w_13939 );
buf ( w_13937 , \4353_b1 );
not ( w_13937 , w_13940 );
not (  , w_13941 );
and ( w_13940 , w_13941 , \4353_b0 );
or ( \4355_b1 , \4168_b1 , \4354_b1 );
xor ( \4355_b0 , \4168_b0 , w_13942 );
not ( w_13942 , w_13943 );
and ( w_13943 , \4354_b1 , \4354_b0 );
buf ( \4356_b1 , \4084_b1 );
not ( \4356_b1 , w_13944 );
not ( \4356_b0 , w_13945 );
and ( w_13944 , w_13945 , \4084_b0 );
buf ( \4357_b1 , \4356_b1 );
not ( \4357_b1 , w_13946 );
not ( \4357_b0 , w_13947 );
and ( w_13946 , w_13947 , \4356_b0 );
buf ( \4358_b1 , \4103_b1 );
not ( \4358_b1 , w_13948 );
not ( \4358_b0 , w_13949 );
and ( w_13948 , w_13949 , \4103_b0 );
or ( \4359_b1 , \4357_b1 , w_13950 );
or ( \4359_b0 , \4357_b0 , \4358_b0 );
not ( \4358_b0 , w_13951 );
and ( w_13951 , w_13950 , \4358_b1 );
or ( \4360_b1 , \4359_b1 , w_13953 );
not ( w_13953 , w_13954 );
and ( \4360_b0 , \4359_b0 , w_13955 );
and ( w_13954 ,  , w_13955 );
buf ( w_13953 , \4088_b1 );
not ( w_13953 , w_13956 );
not (  , w_13957 );
and ( w_13956 , w_13957 , \4088_b0 );
buf ( \4361_b1 , \4360_b1 );
not ( \4361_b1 , w_13958 );
not ( \4361_b0 , w_13959 );
and ( w_13958 , w_13959 , \4360_b0 );
buf ( \4362_b1 , \4165_b1 );
not ( \4362_b1 , w_13960 );
not ( \4362_b0 , w_13961 );
and ( w_13960 , w_13961 , \4165_b0 );
buf ( \4363_b1 , \4136_b1 );
not ( \4363_b1 , w_13962 );
not ( \4363_b0 , w_13963 );
and ( w_13962 , w_13963 , \4136_b0 );
or ( \4364_b1 , \4362_b1 , w_13964 );
or ( \4364_b0 , \4362_b0 , \4363_b0 );
not ( \4363_b0 , w_13965 );
and ( w_13965 , w_13964 , \4363_b1 );
buf ( \4365_b1 , \3994_b1 );
not ( \4365_b1 , w_13966 );
not ( \4365_b0 , w_13967 );
and ( w_13966 , w_13967 , \3994_b0 );
buf ( \4366_b1 , \4142_b1 );
not ( \4366_b1 , w_13968 );
not ( \4366_b0 , w_13969 );
and ( w_13968 , w_13969 , \4142_b0 );
or ( \4367_b1 , \4365_b1 , w_13970 );
or ( \4367_b0 , \4365_b0 , \4366_b0 );
not ( \4366_b0 , w_13971 );
and ( w_13971 , w_13970 , \4366_b1 );
buf ( \4368_b1 , \4142_b1 );
not ( \4368_b1 , w_13972 );
not ( \4368_b0 , w_13973 );
and ( w_13972 , w_13973 , \4142_b0 );
or ( \4369_b1 , \4368_b1 , w_13975 );
not ( w_13975 , w_13976 );
and ( \4369_b0 , \4368_b0 , w_13977 );
and ( w_13976 ,  , w_13977 );
buf ( w_13975 , \4099_b1 );
not ( w_13975 , w_13978 );
not (  , w_13979 );
and ( w_13978 , w_13979 , \4099_b0 );
or ( \4370_b1 , \4367_b1 , w_13981 );
not ( w_13981 , w_13982 );
and ( \4370_b0 , \4367_b0 , w_13983 );
and ( w_13982 ,  , w_13983 );
buf ( w_13981 , \4369_b1 );
not ( w_13981 , w_13984 );
not (  , w_13985 );
and ( w_13984 , w_13985 , \4369_b0 );
or ( \4371_b1 , \4140_b1 , w_13987 );
not ( w_13987 , w_13988 );
and ( \4371_b0 , \4140_b0 , w_13989 );
and ( w_13988 ,  , w_13989 );
buf ( w_13987 , \4370_b1 );
not ( w_13987 , w_13990 );
not (  , w_13991 );
and ( w_13990 , w_13991 , \4370_b0 );
or ( \4372_b1 , \4364_b1 , w_13993 );
not ( w_13993 , w_13994 );
and ( \4372_b0 , \4364_b0 , w_13995 );
and ( w_13994 ,  , w_13995 );
buf ( w_13993 , \4371_b1 );
not ( w_13993 , w_13996 );
not (  , w_13997 );
and ( w_13996 , w_13997 , \4371_b0 );
or ( \4373_b1 , \4361_b1 , \4372_b1 );
xor ( \4373_b0 , \4361_b0 , w_13998 );
not ( w_13998 , w_13999 );
and ( w_13999 , \4372_b1 , \4372_b0 );
buf ( \4374_b1 , \4342_b1 );
not ( \4374_b1 , w_14000 );
not ( \4374_b0 , w_14001 );
and ( w_14000 , w_14001 , \4342_b0 );
buf ( \4375_b1 , \4231_b1 );
not ( \4375_b1 , w_14002 );
not ( \4375_b0 , w_14003 );
and ( w_14002 , w_14003 , \4231_b0 );
or ( \4376_b1 , \4374_b1 , w_14004 );
or ( \4376_b0 , \4374_b0 , \4375_b0 );
not ( \4375_b0 , w_14005 );
and ( w_14005 , w_14004 , \4375_b1 );
buf ( \4377_b1 , \4234_b1 );
buf ( \4377_b0 , \4234_b0 );
buf ( \4378_b1 , \4047_b1 );
not ( \4378_b1 , w_14006 );
not ( \4378_b0 , w_14007 );
and ( w_14006 , w_14007 , \4047_b0 );
buf ( \4379_b1 , \4212_b1 );
not ( \4379_b1 , w_14008 );
not ( \4379_b0 , w_14009 );
and ( w_14008 , w_14009 , \4212_b0 );
or ( \4380_b1 , \4378_b1 , w_14010 );
or ( \4380_b0 , \4378_b0 , \4379_b0 );
not ( \4379_b0 , w_14011 );
and ( w_14011 , w_14010 , \4379_b1 );
or ( \4381_b1 , \4216_b1 , w_14013 );
not ( w_14013 , w_14014 );
and ( \4381_b0 , \4216_b0 , w_14015 );
and ( w_14014 ,  , w_14015 );
buf ( w_14013 , \4178_b1 );
not ( w_14013 , w_14016 );
not (  , w_14017 );
and ( w_14016 , w_14017 , \4178_b0 );
or ( \4382_b1 , \4380_b1 , w_14019 );
not ( w_14019 , w_14020 );
and ( \4382_b0 , \4380_b0 , w_14021 );
and ( w_14020 ,  , w_14021 );
buf ( w_14019 , \4381_b1 );
not ( w_14019 , w_14022 );
not (  , w_14023 );
and ( w_14022 , w_14023 , \4381_b0 );
or ( \4383_b1 , \4377_b1 , w_14025 );
not ( w_14025 , w_14026 );
and ( \4383_b0 , \4377_b0 , w_14027 );
and ( w_14026 ,  , w_14027 );
buf ( w_14025 , \4382_b1 );
not ( w_14025 , w_14028 );
not (  , w_14029 );
and ( w_14028 , w_14029 , \4382_b0 );
or ( \4384_b1 , \4376_b1 , w_14031 );
not ( w_14031 , w_14032 );
and ( \4384_b0 , \4376_b0 , w_14033 );
and ( w_14032 ,  , w_14033 );
buf ( w_14031 , \4383_b1 );
not ( w_14031 , w_14034 );
not (  , w_14035 );
and ( w_14034 , w_14035 , \4383_b0 );
or ( \4385_b1 , \4373_b1 , w_14036 );
xor ( \4385_b0 , \4373_b0 , w_14038 );
not ( w_14038 , w_14039 );
and ( w_14039 , w_14036 , w_14037 );
buf ( w_14036 , \4384_b1 );
not ( w_14036 , w_14040 );
not ( w_14037 , w_14041 );
and ( w_14040 , w_14041 , \4384_b0 );
or ( \4386_b1 , \4355_b1 , w_14042 );
xor ( \4386_b0 , \4355_b0 , w_14044 );
not ( w_14044 , w_14045 );
and ( w_14045 , w_14042 , w_14043 );
buf ( w_14042 , \4385_b1 );
not ( w_14042 , w_14046 );
not ( w_14043 , w_14047 );
and ( w_14046 , w_14047 , \4385_b0 );
or ( \4387_b1 , \4327_b1 , w_14048 );
xor ( \4387_b0 , \4327_b0 , w_14050 );
not ( w_14050 , w_14051 );
and ( w_14051 , w_14048 , w_14049 );
buf ( w_14048 , \4386_b1 );
not ( w_14048 , w_14052 );
not ( w_14049 , w_14053 );
and ( w_14052 , w_14053 , \4386_b0 );
or ( \4388_b1 , \4298_b1 , \4387_b1 );
xor ( \4388_b0 , \4298_b0 , w_14054 );
not ( w_14054 , w_14055 );
and ( w_14055 , \4387_b1 , \4387_b0 );
or ( \4389_b1 , \4352_b1 , \4333_b1 );
not ( \4333_b1 , w_14056 );
and ( \4389_b0 , \4352_b0 , w_14057 );
and ( w_14056 , w_14057 , \4333_b0 );
buf ( \4390_b1 , \4352_b1 );
not ( \4390_b1 , w_14058 );
not ( \4390_b0 , w_14059 );
and ( w_14058 , w_14059 , \4352_b0 );
buf ( \4391_b1 , \4333_b1 );
not ( \4391_b1 , w_14060 );
not ( \4391_b0 , w_14061 );
and ( w_14060 , w_14061 , \4333_b0 );
or ( \4392_b1 , \4390_b1 , \4391_b1 );
not ( \4391_b1 , w_14062 );
and ( \4392_b0 , \4390_b0 , w_14063 );
and ( w_14062 , w_14063 , \4391_b0 );
or ( \4393_b1 , \4389_b1 , w_14065 );
not ( w_14065 , w_14066 );
and ( \4393_b0 , \4389_b0 , w_14067 );
and ( w_14066 ,  , w_14067 );
buf ( w_14065 , \4392_b1 );
not ( w_14065 , w_14068 );
not (  , w_14069 );
and ( w_14068 , w_14069 , \4392_b0 );
buf ( \4394_b1 , \4344_b1 );
buf ( \4394_b0 , \4344_b0 );
or ( \4395_b1 , \4393_b1 , w_14070 );
xor ( \4395_b0 , \4393_b0 , w_14072 );
not ( w_14072 , w_14073 );
and ( w_14073 , w_14070 , w_14071 );
buf ( w_14070 , \4394_b1 );
not ( w_14070 , w_14074 );
not ( w_14071 , w_14075 );
and ( w_14074 , w_14075 , \4394_b0 );
buf ( \4396_b1 , \4395_b1 );
not ( \4396_b1 , w_14076 );
not ( \4396_b0 , w_14077 );
and ( w_14076 , w_14077 , \4395_b0 );
buf ( \4397_b1 , \4396_b1 );
not ( \4397_b1 , w_14078 );
not ( \4397_b0 , w_14079 );
and ( w_14078 , w_14079 , \4396_b0 );
buf ( \4398_b1 , \4056_b1 );
not ( \4398_b1 , w_14080 );
not ( \4398_b0 , w_14081 );
and ( w_14080 , w_14081 , \4056_b0 );
buf ( \4399_b1 , \4070_b1 );
not ( \4399_b1 , w_14082 );
not ( \4399_b0 , w_14083 );
and ( w_14082 , w_14083 , \4070_b0 );
buf ( \4400_b1 , \4399_b1 );
not ( \4400_b1 , w_14084 );
not ( \4400_b0 , w_14085 );
and ( w_14084 , w_14085 , \4399_b0 );
or ( \4401_b1 , \4398_b1 , \4400_b1 );
not ( \4400_b1 , w_14086 );
and ( \4401_b0 , \4398_b0 , w_14087 );
and ( w_14086 , w_14087 , \4400_b0 );
buf ( \4402_b1 , \3994_b1 );
not ( \4402_b1 , w_14088 );
not ( \4402_b0 , w_14089 );
and ( w_14088 , w_14089 , \3994_b0 );
buf ( \4403_b1 , \3880_b1 );
buf ( \4403_b0 , \3880_b0 );
buf ( \4404_b1 , \4403_b1 );
not ( \4404_b1 , w_14090 );
not ( \4404_b0 , w_14091 );
and ( w_14090 , w_14091 , \4403_b0 );
buf ( \4405_b1 , \4404_b1 );
not ( \4405_b1 , w_14092 );
not ( \4405_b0 , w_14093 );
and ( w_14092 , w_14093 , \4404_b0 );
or ( \4406_b1 , \4402_b1 , w_14094 );
or ( \4406_b0 , \4402_b0 , \4405_b0 );
not ( \4405_b0 , w_14095 );
and ( w_14095 , w_14094 , \4405_b1 );
buf ( \4407_b1 , \4069_b1 );
not ( \4407_b1 , w_14096 );
not ( \4407_b0 , w_14097 );
and ( w_14096 , w_14097 , \4069_b0 );
or ( \4408_b1 , \4407_b1 , w_14099 );
not ( w_14099 , w_14100 );
and ( \4408_b0 , \4407_b0 , w_14101 );
and ( w_14100 ,  , w_14101 );
buf ( w_14099 , \4099_b1 );
not ( w_14099 , w_14102 );
not (  , w_14103 );
and ( w_14102 , w_14103 , \4099_b0 );
or ( \4409_b1 , \4406_b1 , w_14105 );
not ( w_14105 , w_14106 );
and ( \4409_b0 , \4406_b0 , w_14107 );
and ( w_14106 ,  , w_14107 );
buf ( w_14105 , \4408_b1 );
not ( w_14105 , w_14108 );
not (  , w_14109 );
and ( w_14108 , w_14109 , \4408_b0 );
buf ( \4410_b1 , \4409_b1 );
not ( \4410_b1 , w_14110 );
not ( \4410_b0 , w_14111 );
and ( w_14110 , w_14111 , \4409_b0 );
buf ( \4411_b1 , \4065_b1 );
not ( \4411_b1 , w_14112 );
not ( \4411_b0 , w_14113 );
and ( w_14112 , w_14113 , \4065_b0 );
or ( \4412_b1 , \4410_b1 , w_14115 );
not ( w_14115 , w_14116 );
and ( \4412_b0 , \4410_b0 , w_14117 );
and ( w_14116 ,  , w_14117 );
buf ( w_14115 , \4411_b1 );
not ( w_14115 , w_14118 );
not (  , w_14119 );
and ( w_14118 , w_14119 , \4411_b0 );
or ( \4413_b1 , \4401_b1 , w_14121 );
not ( w_14121 , w_14122 );
and ( \4413_b0 , \4401_b0 , w_14123 );
and ( w_14122 ,  , w_14123 );
buf ( w_14121 , \4412_b1 );
not ( w_14121 , w_14124 );
not (  , w_14125 );
and ( w_14124 , w_14125 , \4412_b0 );
buf ( \4414_b1 , \4413_b1 );
not ( \4414_b1 , w_14126 );
not ( \4414_b0 , w_14127 );
and ( w_14126 , w_14127 , \4413_b0 );
buf ( \4415_b1 , \4414_b1 );
not ( \4415_b1 , w_14128 );
not ( \4415_b0 , w_14129 );
and ( w_14128 , w_14129 , \4414_b0 );
or ( \4416_b1 , \4156_b1 , w_14131 );
not ( w_14131 , w_14132 );
and ( \4416_b0 , \4156_b0 , w_14133 );
and ( w_14132 ,  , w_14133 );
buf ( w_14131 , \3958_b1 );
not ( w_14131 , w_14134 );
not (  , w_14135 );
and ( w_14134 , w_14135 , \3958_b0 );
or ( \4417_b1 , \4415_b1 , w_14137 );
not ( w_14137 , w_14138 );
and ( \4417_b0 , \4415_b0 , w_14139 );
and ( w_14138 ,  , w_14139 );
buf ( w_14137 , \4416_b1 );
not ( w_14137 , w_14140 );
not (  , w_14141 );
and ( w_14140 , w_14141 , \4416_b0 );
buf ( \4418_b1 , \4417_b1 );
not ( \4418_b1 , w_14142 );
not ( \4418_b0 , w_14143 );
and ( w_14142 , w_14143 , \4417_b0 );
buf ( \4419_b1 , \4047_b1 );
not ( \4419_b1 , w_14144 );
not ( \4419_b0 , w_14145 );
and ( w_14144 , w_14145 , \4047_b0 );
buf ( \4420_b1 , \4110_b1 );
not ( \4420_b1 , w_14146 );
not ( \4420_b0 , w_14147 );
and ( w_14146 , w_14147 , \4110_b0 );
or ( \4421_b1 , \4419_b1 , w_14148 );
or ( \4421_b0 , \4419_b0 , \4420_b0 );
not ( \4420_b0 , w_14149 );
and ( w_14149 , w_14148 , \4420_b1 );
or ( \4422_b1 , \4109_b1 , w_14151 );
not ( w_14151 , w_14152 );
and ( \4422_b0 , \4109_b0 , w_14153 );
and ( w_14152 ,  , w_14153 );
buf ( w_14151 , \4178_b1 );
not ( w_14151 , w_14154 );
not (  , w_14155 );
and ( w_14154 , w_14155 , \4178_b0 );
or ( \4423_b1 , \4421_b1 , w_14157 );
not ( w_14157 , w_14158 );
and ( \4423_b0 , \4421_b0 , w_14159 );
and ( w_14158 ,  , w_14159 );
buf ( w_14157 , \4422_b1 );
not ( w_14157 , w_14160 );
not (  , w_14161 );
and ( w_14160 , w_14161 , \4422_b0 );
buf ( \4424_b1 , \4423_b1 );
not ( \4424_b1 , w_14162 );
not ( \4424_b0 , w_14163 );
and ( w_14162 , w_14163 , \4423_b0 );
buf ( \4425_b1 , \4135_b1 );
not ( \4425_b1 , w_14164 );
not ( \4425_b0 , w_14165 );
and ( w_14164 , w_14165 , \4135_b0 );
buf ( \4426_b1 , \4425_b1 );
not ( \4426_b1 , w_14166 );
not ( \4426_b0 , w_14167 );
and ( w_14166 , w_14167 , \4425_b0 );
or ( \4427_b1 , \4424_b1 , w_14168 );
or ( \4427_b0 , \4424_b0 , \4426_b0 );
not ( \4426_b0 , w_14169 );
and ( w_14169 , w_14168 , \4426_b1 );
buf ( \4428_b1 , \4139_b1 );
not ( \4428_b1 , w_14170 );
not ( \4428_b0 , w_14171 );
and ( w_14170 , w_14171 , \4139_b0 );
buf ( \4429_b1 , \4428_b1 );
not ( \4429_b1 , w_14172 );
not ( \4429_b0 , w_14173 );
and ( w_14172 , w_14173 , \4428_b0 );
or ( \4430_b1 , \4118_b1 , w_14175 );
not ( w_14175 , w_14176 );
and ( \4430_b0 , \4118_b0 , w_14177 );
and ( w_14176 ,  , w_14177 );
buf ( w_14175 , \4429_b1 );
not ( w_14175 , w_14178 );
not (  , w_14179 );
and ( w_14178 , w_14179 , \4429_b0 );
or ( \4431_b1 , \4427_b1 , w_14181 );
not ( w_14181 , w_14182 );
and ( \4431_b0 , \4427_b0 , w_14183 );
and ( w_14182 ,  , w_14183 );
buf ( w_14181 , \4430_b1 );
not ( w_14181 , w_14184 );
not (  , w_14185 );
and ( w_14184 , w_14185 , \4430_b0 );
or ( \4432_b1 , \3943_b1 , \4088_b1 );
not ( \4088_b1 , w_14186 );
and ( \4432_b0 , \3943_b0 , w_14187 );
and ( w_14186 , w_14187 , \4088_b0 );
buf ( \4433_b1 , \3943_b1 );
not ( \4433_b1 , w_14188 );
not ( \4433_b0 , w_14189 );
and ( w_14188 , w_14189 , \3943_b0 );
or ( \4434_b1 , \4433_b1 , \4089_b1 );
not ( \4089_b1 , w_14190 );
and ( \4434_b0 , \4433_b0 , w_14191 );
and ( w_14190 , w_14191 , \4089_b0 );
or ( \4435_b1 , \4432_b1 , w_14193 );
not ( w_14193 , w_14194 );
and ( \4435_b0 , \4432_b0 , w_14195 );
and ( w_14194 ,  , w_14195 );
buf ( w_14193 , \4434_b1 );
not ( w_14193 , w_14196 );
not (  , w_14197 );
and ( w_14196 , w_14197 , \4434_b0 );
buf ( \4436_b1 , \4435_b1 );
not ( \4436_b1 , w_14198 );
not ( \4436_b0 , w_14199 );
and ( w_14198 , w_14199 , \4435_b0 );
buf ( \4437_b1 , \4085_b1 );
buf ( \4437_b0 , \4085_b0 );
buf ( \4438_b1 , \4437_b1 );
not ( \4438_b1 , w_14200 );
not ( \4438_b0 , w_14201 );
and ( w_14200 , w_14201 , \4437_b0 );
or ( \4439_b1 , \4436_b1 , w_14202 );
or ( \4439_b0 , \4436_b0 , \4438_b0 );
not ( \4438_b0 , w_14203 );
and ( w_14203 , w_14202 , \4438_b1 );
or ( \4440_b1 , \4331_b1 , w_14205 );
not ( w_14205 , w_14206 );
and ( \4440_b0 , \4331_b0 , w_14207 );
and ( w_14206 ,  , w_14207 );
buf ( w_14205 , \4094_b1 );
not ( w_14205 , w_14208 );
not (  , w_14209 );
and ( w_14208 , w_14209 , \4094_b0 );
or ( \4441_b1 , \4439_b1 , w_14211 );
not ( w_14211 , w_14212 );
and ( \4441_b0 , \4439_b0 , w_14213 );
and ( w_14212 ,  , w_14213 );
buf ( w_14211 , \4440_b1 );
not ( w_14211 , w_14214 );
not (  , w_14215 );
and ( w_14214 , w_14215 , \4440_b0 );
or ( \4442_b1 , \4431_b1 , \4441_b1 );
xor ( \4442_b0 , \4431_b0 , w_14216 );
not ( w_14216 , w_14217 );
and ( w_14217 , \4441_b1 , \4441_b0 );
or ( \4443_b1 , \4041_b1 , \4285_b1 );
not ( \4285_b1 , w_14218 );
and ( \4443_b0 , \4041_b0 , w_14219 );
and ( w_14218 , w_14219 , \4285_b0 );
buf ( \4444_b1 , \4041_b1 );
not ( \4444_b1 , w_14220 );
not ( \4444_b0 , w_14221 );
and ( w_14220 , w_14221 , \4041_b0 );
or ( \4445_b1 , \4444_b1 , \4176_b1 );
not ( \4176_b1 , w_14222 );
and ( \4445_b0 , \4444_b0 , w_14223 );
and ( w_14222 , w_14223 , \4176_b0 );
or ( \4446_b1 , \4443_b1 , w_14225 );
not ( w_14225 , w_14226 );
and ( \4446_b0 , \4443_b0 , w_14227 );
and ( w_14226 ,  , w_14227 );
buf ( w_14225 , \4445_b1 );
not ( w_14225 , w_14228 );
not (  , w_14229 );
and ( w_14228 , w_14229 , \4445_b0 );
buf ( \4447_b1 , \4446_b1 );
not ( \4447_b1 , w_14230 );
not ( \4447_b0 , w_14231 );
and ( w_14230 , w_14231 , \4446_b0 );
buf ( \4448_b1 , \4195_b1 );
not ( \4448_b1 , w_14232 );
not ( \4448_b0 , w_14233 );
and ( w_14232 , w_14233 , \4195_b0 );
or ( \4449_b1 , \4447_b1 , w_14234 );
or ( \4449_b0 , \4447_b0 , \4448_b0 );
not ( \4448_b0 , w_14235 );
and ( w_14235 , w_14234 , \4448_b1 );
or ( \4450_b1 , \4205_b1 , w_14237 );
not ( w_14237 , w_14238 );
and ( \4450_b0 , \4205_b0 , w_14239 );
and ( w_14238 ,  , w_14239 );
buf ( w_14237 , \4288_b1 );
not ( w_14237 , w_14240 );
not (  , w_14241 );
and ( w_14240 , w_14241 , \4288_b0 );
or ( \4451_b1 , \4449_b1 , w_14243 );
not ( w_14243 , w_14244 );
and ( \4451_b0 , \4449_b0 , w_14245 );
and ( w_14244 ,  , w_14245 );
buf ( w_14243 , \4450_b1 );
not ( w_14243 , w_14246 );
not (  , w_14247 );
and ( w_14246 , w_14247 , \4450_b0 );
or ( \4452_b1 , \4442_b1 , \4451_b1 );
not ( \4451_b1 , w_14248 );
and ( \4452_b0 , \4442_b0 , w_14249 );
and ( w_14248 , w_14249 , \4451_b0 );
or ( \4453_b1 , \4431_b1 , \4441_b1 );
not ( \4441_b1 , w_14250 );
and ( \4453_b0 , \4431_b0 , w_14251 );
and ( w_14250 , w_14251 , \4441_b0 );
or ( \4454_b1 , \4452_b1 , w_14252 );
or ( \4454_b0 , \4452_b0 , \4453_b0 );
not ( \4453_b0 , w_14253 );
and ( w_14253 , w_14252 , \4453_b1 );
buf ( \4455_b1 , \4454_b1 );
not ( \4455_b1 , w_14254 );
not ( \4455_b0 , w_14255 );
and ( w_14254 , w_14255 , \4454_b0 );
or ( \4456_b1 , \4418_b1 , w_14256 );
or ( \4456_b0 , \4418_b0 , \4455_b0 );
not ( \4455_b0 , w_14257 );
and ( w_14257 , w_14256 , \4455_b1 );
buf ( \4457_b1 , \4416_b1 );
not ( \4457_b1 , w_14258 );
not ( \4457_b0 , w_14259 );
and ( w_14258 , w_14259 , \4416_b0 );
or ( \4458_b1 , \4457_b1 , w_14261 );
not ( w_14261 , w_14262 );
and ( \4458_b0 , \4457_b0 , w_14263 );
and ( w_14262 ,  , w_14263 );
buf ( w_14261 , \4414_b1 );
not ( w_14261 , w_14264 );
not (  , w_14265 );
and ( w_14264 , w_14265 , \4414_b0 );
or ( \4459_b1 , \4456_b1 , w_14267 );
not ( w_14267 , w_14268 );
and ( \4459_b0 , \4456_b0 , w_14269 );
and ( w_14268 ,  , w_14269 );
buf ( w_14267 , \4458_b1 );
not ( w_14267 , w_14270 );
not (  , w_14271 );
and ( w_14270 , w_14271 , \4458_b0 );
buf ( \4460_b1 , \4459_b1 );
not ( \4460_b1 , w_14272 );
not ( \4460_b0 , w_14273 );
and ( w_14272 , w_14273 , \4459_b0 );
or ( \4461_b1 , \4397_b1 , w_14274 );
or ( \4461_b0 , \4397_b0 , \4460_b0 );
not ( \4460_b0 , w_14275 );
and ( w_14275 , w_14274 , \4460_b1 );
buf ( \4462_b1 , \4242_b1 );
not ( \4462_b1 , w_14276 );
not ( \4462_b0 , w_14277 );
and ( w_14276 , w_14277 , \4242_b0 );
or ( \4463_b1 , \4293_b1 , \4462_b1 );
xor ( \4463_b0 , \4293_b0 , w_14278 );
not ( w_14278 , w_14279 );
and ( w_14279 , \4462_b1 , \4462_b0 );
or ( \4464_b1 , \4463_b1 , \4276_b1 );
xor ( \4464_b0 , \4463_b0 , w_14280 );
not ( w_14280 , w_14281 );
and ( w_14281 , \4276_b1 , \4276_b0 );
or ( \4465_b1 , \4151_b1 , \4072_b1 );
not ( \4072_b1 , w_14282 );
and ( \4465_b0 , \4151_b0 , w_14283 );
and ( w_14282 , w_14283 , \4072_b0 );
buf ( \4466_b1 , \4151_b1 );
not ( \4466_b1 , w_14284 );
not ( \4466_b0 , w_14285 );
and ( w_14284 , w_14285 , \4151_b0 );
or ( \4467_b1 , \4466_b1 , \4071_b1 );
not ( \4071_b1 , w_14286 );
and ( \4467_b0 , \4466_b0 , w_14287 );
and ( w_14286 , w_14287 , \4071_b0 );
or ( \4468_b1 , \4465_b1 , w_14288 );
or ( \4468_b0 , \4465_b0 , \4467_b0 );
not ( \4467_b0 , w_14289 );
and ( w_14289 , w_14288 , \4467_b1 );
or ( \4469_b1 , \4468_b1 , \4105_b1 );
not ( \4105_b1 , w_14290 );
and ( \4469_b0 , \4468_b0 , w_14291 );
and ( w_14290 , w_14291 , \4105_b0 );
buf ( \4470_b1 , \4468_b1 );
not ( \4470_b1 , w_14292 );
not ( \4470_b0 , w_14293 );
and ( w_14292 , w_14293 , \4468_b0 );
or ( \4471_b1 , \4470_b1 , \4153_b1 );
not ( \4153_b1 , w_14294 );
and ( \4471_b0 , \4470_b0 , w_14295 );
and ( w_14294 , w_14295 , \4153_b0 );
or ( \4472_b1 , \4469_b1 , w_14297 );
not ( w_14297 , w_14298 );
and ( \4472_b0 , \4469_b0 , w_14299 );
and ( w_14298 ,  , w_14299 );
buf ( w_14297 , \4471_b1 );
not ( w_14297 , w_14300 );
not (  , w_14301 );
and ( w_14300 , w_14301 , \4471_b0 );
buf ( \4473_b1 , \3958_b1 );
not ( \4473_b1 , w_14302 );
not ( \4473_b0 , w_14303 );
and ( w_14302 , w_14303 , \3958_b0 );
buf ( \4474_b1 , \4473_b1 );
not ( \4474_b1 , w_14304 );
not ( \4474_b0 , w_14305 );
and ( w_14304 , w_14305 , \4473_b0 );
buf ( \4475_b1 , \4156_b1 );
not ( \4475_b1 , w_14306 );
not ( \4475_b0 , w_14307 );
and ( w_14306 , w_14307 , \4156_b0 );
or ( \4476_b1 , \4474_b1 , w_14308 );
or ( \4476_b0 , \4474_b0 , \4475_b0 );
not ( \4475_b0 , w_14309 );
and ( w_14309 , w_14308 , \4475_b1 );
or ( \4477_b1 , \4267_b1 , w_14311 );
not ( w_14311 , w_14312 );
and ( \4477_b0 , \4267_b0 , w_14313 );
and ( w_14312 ,  , w_14313 );
buf ( w_14311 , \3958_b1 );
not ( w_14311 , w_14314 );
not (  , w_14315 );
and ( w_14314 , w_14315 , \3958_b0 );
or ( \4478_b1 , \4476_b1 , w_14317 );
not ( w_14317 , w_14318 );
and ( \4478_b0 , \4476_b0 , w_14319 );
and ( w_14318 ,  , w_14319 );
buf ( w_14317 , \4477_b1 );
not ( w_14317 , w_14320 );
not (  , w_14321 );
and ( w_14320 , w_14321 , \4477_b0 );
buf ( \4479_b1 , \4478_b1 );
not ( \4479_b1 , w_14322 );
not ( \4479_b0 , w_14323 );
and ( w_14322 , w_14323 , \4478_b0 );
or ( \4480_b1 , \4251_b1 , \4252_b1 );
not ( \4252_b1 , w_14324 );
and ( \4480_b0 , \4251_b0 , w_14325 );
and ( w_14324 , w_14325 , \4252_b0 );
buf ( \4481_b1 , \4480_b1 );
not ( \4481_b1 , w_14326 );
not ( \4481_b0 , w_14327 );
and ( w_14326 , w_14327 , \4480_b0 );
or ( \4482_b1 , \4479_b1 , w_14328 );
or ( \4482_b0 , \4479_b0 , \4481_b0 );
not ( \4481_b0 , w_14329 );
and ( w_14329 , w_14328 , \4481_b1 );
or ( \4483_b1 , \4262_b1 , w_14331 );
not ( w_14331 , w_14332 );
and ( \4483_b0 , \4262_b0 , w_14333 );
and ( w_14332 ,  , w_14333 );
buf ( w_14331 , \4273_b1 );
not ( w_14331 , w_14334 );
not (  , w_14335 );
and ( w_14334 , w_14335 , \4273_b0 );
or ( \4484_b1 , \4482_b1 , w_14337 );
not ( w_14337 , w_14338 );
and ( \4484_b0 , \4482_b0 , w_14339 );
and ( w_14338 ,  , w_14339 );
buf ( w_14337 , \4483_b1 );
not ( w_14337 , w_14340 );
not (  , w_14341 );
and ( w_14340 , w_14341 , \4483_b0 );
buf ( \4485_b1 , \4156_b1 );
not ( \4485_b1 , w_14342 );
not ( \4485_b0 , w_14343 );
and ( w_14342 , w_14343 , \4156_b0 );
buf ( \4486_b1 , \3963_b1 );
not ( \4486_b1 , w_14344 );
not ( \4486_b0 , w_14345 );
and ( w_14344 , w_14345 , \3963_b0 );
or ( \4487_b1 , \4485_b1 , w_14347 );
not ( w_14347 , w_14348 );
and ( \4487_b0 , \4485_b0 , w_14349 );
and ( w_14348 ,  , w_14349 );
buf ( w_14347 , \4486_b1 );
not ( w_14347 , w_14350 );
not (  , w_14351 );
and ( w_14350 , w_14351 , \4486_b0 );
or ( \4488_b1 , \4484_b1 , w_14353 );
not ( w_14353 , w_14354 );
and ( \4488_b0 , \4484_b0 , w_14355 );
and ( w_14354 ,  , w_14355 );
buf ( w_14353 , \4487_b1 );
not ( w_14353 , w_14356 );
not (  , w_14357 );
and ( w_14356 , w_14357 , \4487_b0 );
buf ( \4489_b1 , \4011_b1 );
not ( \4489_b1 , w_14358 );
not ( \4489_b0 , w_14359 );
and ( w_14358 , w_14359 , \4011_b0 );
buf ( \4490_b1 , \4212_b1 );
not ( \4490_b1 , w_14360 );
not ( \4490_b0 , w_14361 );
and ( w_14360 , w_14361 , \4212_b0 );
or ( \4491_b1 , \4489_b1 , w_14362 );
or ( \4491_b0 , \4489_b0 , \4490_b0 );
not ( \4490_b0 , w_14363 );
and ( w_14363 , w_14362 , \4490_b1 );
buf ( \4492_b1 , \3577_b1 );
buf ( \4492_b0 , \3577_b0 );
or ( \4493_b1 , \4492_b1 , w_14365 );
not ( w_14365 , w_14366 );
and ( \4493_b0 , \4492_b0 , w_14367 );
and ( w_14366 ,  , w_14367 );
buf ( w_14365 , \4270_b1 );
not ( w_14365 , w_14368 );
not (  , w_14369 );
and ( w_14368 , w_14369 , \4270_b0 );
or ( \4494_b1 , \4491_b1 , w_14371 );
not ( w_14371 , w_14372 );
and ( \4494_b0 , \4491_b0 , w_14373 );
and ( w_14372 ,  , w_14373 );
buf ( w_14371 , \4493_b1 );
not ( w_14371 , w_14374 );
not (  , w_14375 );
and ( w_14374 , w_14375 , \4493_b0 );
buf ( \4495_b1 , \4494_b1 );
not ( \4495_b1 , w_14376 );
not ( \4495_b0 , w_14377 );
and ( w_14376 , w_14377 , \4494_b0 );
buf ( \4496_b1 , \4231_b1 );
buf ( \4496_b0 , \4231_b0 );
buf ( \4497_b1 , \4496_b1 );
not ( \4497_b1 , w_14378 );
not ( \4497_b0 , w_14379 );
and ( w_14378 , w_14379 , \4496_b0 );
or ( \4498_b1 , \4495_b1 , w_14380 );
or ( \4498_b0 , \4495_b0 , \4497_b0 );
not ( \4497_b0 , w_14381 );
and ( w_14381 , w_14380 , \4497_b1 );
or ( \4499_b1 , \4377_b1 , w_14383 );
not ( w_14383 , w_14384 );
and ( \4499_b0 , \4377_b0 , w_14385 );
and ( w_14384 ,  , w_14385 );
buf ( w_14383 , \4219_b1 );
not ( w_14383 , w_14386 );
not (  , w_14387 );
and ( w_14386 , w_14387 , \4219_b0 );
or ( \4500_b1 , \4498_b1 , w_14389 );
not ( w_14389 , w_14390 );
and ( \4500_b0 , \4498_b0 , w_14391 );
and ( w_14390 ,  , w_14391 );
buf ( w_14389 , \4499_b1 );
not ( w_14389 , w_14392 );
not (  , w_14393 );
and ( w_14392 , w_14393 , \4499_b0 );
buf ( \4501_b1 , \4500_b1 );
not ( \4501_b1 , w_14394 );
not ( \4501_b0 , w_14395 );
and ( w_14394 , w_14395 , \4500_b0 );
or ( \4502_b1 , \4488_b1 , w_14396 );
or ( \4502_b0 , \4488_b0 , \4501_b0 );
not ( \4501_b0 , w_14397 );
and ( w_14397 , w_14396 , \4501_b1 );
or ( \4503_b1 , \4484_b1 , w_14399 );
not ( w_14399 , w_14400 );
and ( \4503_b0 , \4484_b0 , w_14401 );
and ( w_14400 ,  , w_14401 );
buf ( w_14399 , \4487_b1 );
not ( w_14399 , w_14402 );
not (  , w_14403 );
and ( w_14402 , w_14403 , \4487_b0 );
or ( \4504_b1 , \4502_b1 , w_14405 );
not ( w_14405 , w_14406 );
and ( \4504_b0 , \4502_b0 , w_14407 );
and ( w_14406 ,  , w_14407 );
buf ( w_14405 , \4503_b1 );
not ( w_14405 , w_14408 );
not (  , w_14409 );
and ( w_14408 , w_14409 , \4503_b0 );
buf ( \4505_b1 , \4504_b1 );
not ( \4505_b1 , w_14410 );
not ( \4505_b0 , w_14411 );
and ( w_14410 , w_14411 , \4504_b0 );
or ( \4506_b1 , \4472_b1 , w_14413 );
not ( w_14413 , w_14414 );
and ( \4506_b0 , \4472_b0 , w_14415 );
and ( w_14414 ,  , w_14415 );
buf ( w_14413 , \4505_b1 );
not ( w_14413 , w_14416 );
not (  , w_14417 );
and ( w_14416 , w_14417 , \4505_b0 );
or ( \4507_b1 , \4464_b1 , \4506_b1 );
not ( \4506_b1 , w_14418 );
and ( \4507_b0 , \4464_b0 , w_14419 );
and ( w_14418 , w_14419 , \4506_b0 );
or ( \4508_b1 , \4472_b1 , w_14421 );
not ( w_14421 , w_14422 );
and ( \4508_b0 , \4472_b0 , w_14423 );
and ( w_14422 ,  , w_14423 );
buf ( w_14421 , \4505_b1 );
not ( w_14421 , w_14424 );
not (  , w_14425 );
and ( w_14424 , w_14425 , \4505_b0 );
or ( \4509_b1 , \4507_b1 , w_14427 );
not ( w_14427 , w_14428 );
and ( \4509_b0 , \4507_b0 , w_14429 );
and ( w_14428 ,  , w_14429 );
buf ( w_14427 , \4508_b1 );
not ( w_14427 , w_14430 );
not (  , w_14431 );
and ( w_14430 , w_14431 , \4508_b0 );
buf ( \4510_b1 , \4509_b1 );
not ( \4510_b1 , w_14432 );
not ( \4510_b0 , w_14433 );
and ( w_14432 , w_14433 , \4509_b0 );
buf ( \4511_b1 , \4459_b1 );
not ( \4511_b1 , w_14434 );
not ( \4511_b0 , w_14435 );
and ( w_14434 , w_14435 , \4459_b0 );
or ( \4512_b1 , \4511_b1 , w_14437 );
not ( w_14437 , w_14438 );
and ( \4512_b0 , \4511_b0 , w_14439 );
and ( w_14438 ,  , w_14439 );
buf ( w_14437 , \4395_b1 );
not ( w_14437 , w_14440 );
not (  , w_14441 );
and ( w_14440 , w_14441 , \4395_b0 );
or ( \4513_b1 , \4510_b1 , w_14443 );
not ( w_14443 , w_14444 );
and ( \4513_b0 , \4510_b0 , w_14445 );
and ( w_14444 ,  , w_14445 );
buf ( w_14443 , \4512_b1 );
not ( w_14443 , w_14446 );
not (  , w_14447 );
and ( w_14446 , w_14447 , \4512_b0 );
or ( \4514_b1 , \4461_b1 , w_14449 );
not ( w_14449 , w_14450 );
and ( \4514_b0 , \4461_b0 , w_14451 );
and ( w_14450 ,  , w_14451 );
buf ( w_14449 , \4513_b1 );
not ( w_14449 , w_14452 );
not (  , w_14453 );
and ( w_14452 , w_14453 , \4513_b0 );
or ( \4515_b1 , \4388_b1 , \4514_b1 );
xor ( \4515_b0 , \4388_b0 , w_14454 );
not ( w_14454 , w_14455 );
and ( w_14455 , \4514_b1 , \4514_b0 );
buf ( \4516_b1 , \4515_b1 );
not ( \4516_b1 , w_14456 );
not ( \4516_b0 , w_14457 );
and ( w_14456 , w_14457 , \4515_b0 );
or ( \4517_b1 , \4155_b1 , \4208_b1 );
xor ( \4517_b0 , \4155_b0 , w_14458 );
not ( w_14458 , w_14459 );
and ( w_14459 , \4208_b1 , \4208_b0 );
or ( \4518_b1 , \4517_b1 , \4295_b1 );
xor ( \4518_b0 , \4517_b0 , w_14460 );
not ( w_14460 , w_14461 );
and ( w_14461 , \4295_b1 , \4295_b0 );
buf ( \4519_b1 , \4518_b1 );
not ( \4519_b1 , w_14462 );
not ( \4519_b0 , w_14463 );
and ( w_14462 , w_14463 , \4518_b0 );
buf ( \4520_b1 , \4510_b1 );
not ( \4520_b1 , w_14464 );
not ( \4520_b0 , w_14465 );
and ( w_14464 , w_14465 , \4510_b0 );
buf ( \4521_b1 , \4395_b1 );
not ( \4521_b1 , w_14466 );
not ( \4521_b0 , w_14467 );
and ( w_14466 , w_14467 , \4395_b0 );
buf ( \4522_b1 , \4459_b1 );
not ( \4522_b1 , w_14468 );
not ( \4522_b0 , w_14469 );
and ( w_14468 , w_14469 , \4459_b0 );
or ( \4523_b1 , \4521_b1 , w_14470 );
or ( \4523_b0 , \4521_b0 , \4522_b0 );
not ( \4522_b0 , w_14471 );
and ( w_14471 , w_14470 , \4522_b1 );
or ( \4524_b1 , \4459_b1 , w_14472 );
or ( \4524_b0 , \4459_b0 , \4395_b0 );
not ( \4395_b0 , w_14473 );
and ( w_14473 , w_14472 , \4395_b1 );
or ( \4525_b1 , \4523_b1 , w_14475 );
not ( w_14475 , w_14476 );
and ( \4525_b0 , \4523_b0 , w_14477 );
and ( w_14476 ,  , w_14477 );
buf ( w_14475 , \4524_b1 );
not ( w_14475 , w_14478 );
not (  , w_14479 );
and ( w_14478 , w_14479 , \4524_b0 );
buf ( \4526_b1 , \4525_b1 );
not ( \4526_b1 , w_14480 );
not ( \4526_b0 , w_14481 );
and ( w_14480 , w_14481 , \4525_b0 );
buf ( \4527_b1 , \4526_b1 );
not ( \4527_b1 , w_14482 );
not ( \4527_b0 , w_14483 );
and ( w_14482 , w_14483 , \4526_b0 );
or ( \4528_b1 , \4520_b1 , w_14484 );
or ( \4528_b0 , \4520_b0 , \4527_b0 );
not ( \4527_b0 , w_14485 );
and ( w_14485 , w_14484 , \4527_b1 );
or ( \4529_b1 , \4525_b1 , w_14487 );
not ( w_14487 , w_14488 );
and ( \4529_b0 , \4525_b0 , w_14489 );
and ( w_14488 ,  , w_14489 );
buf ( w_14487 , \4509_b1 );
not ( w_14487 , w_14490 );
not (  , w_14491 );
and ( w_14490 , w_14491 , \4509_b0 );
or ( \4530_b1 , \4528_b1 , w_14493 );
not ( w_14493 , w_14494 );
and ( \4530_b0 , \4528_b0 , w_14495 );
and ( w_14494 ,  , w_14495 );
buf ( w_14493 , \4529_b1 );
not ( w_14493 , w_14496 );
not (  , w_14497 );
and ( w_14496 , w_14497 , \4529_b0 );
buf ( \4531_b1 , \4530_b1 );
not ( \4531_b1 , w_14498 );
not ( \4531_b0 , w_14499 );
and ( w_14498 , w_14499 , \4530_b0 );
or ( \4532_b1 , \4519_b1 , w_14500 );
or ( \4532_b0 , \4519_b0 , \4531_b0 );
not ( \4531_b0 , w_14501 );
and ( w_14501 , w_14500 , \4531_b1 );
or ( \4533_b1 , \4530_b1 , w_14502 );
or ( \4533_b0 , \4530_b0 , \4518_b0 );
not ( \4518_b0 , w_14503 );
and ( w_14503 , w_14502 , \4518_b1 );
buf ( \4534_b1 , \1528_b1 );
not ( \4534_b1 , w_14504 );
not ( \4534_b0 , w_14505 );
and ( w_14504 , w_14505 , \1528_b0 );
buf ( \4535_b1 , \3432_b1 );
not ( \4535_b1 , w_14506 );
not ( \4535_b0 , w_14507 );
and ( w_14506 , w_14507 , \3432_b0 );
buf ( \4536_b1 , \4535_b1 );
not ( \4536_b1 , w_14508 );
not ( \4536_b0 , w_14509 );
and ( w_14508 , w_14509 , \4535_b0 );
or ( \4537_b1 , \4534_b1 , w_14510 );
or ( \4537_b0 , \4534_b0 , \4536_b0 );
not ( \4536_b0 , w_14511 );
and ( w_14511 , w_14510 , \4536_b1 );
buf ( \4538_b1 , \1528_b1 );
not ( \4538_b1 , w_14512 );
not ( \4538_b0 , w_14513 );
and ( w_14512 , w_14513 , \1528_b0 );
or ( \4539_b1 , \4538_b1 , w_14515 );
not ( w_14515 , w_14516 );
and ( \4539_b0 , \4538_b0 , w_14517 );
and ( w_14516 ,  , w_14517 );
buf ( w_14515 , \3432_b1 );
not ( w_14515 , w_14518 );
not (  , w_14519 );
and ( w_14518 , w_14519 , \3432_b0 );
or ( \4540_b1 , \4537_b1 , w_14521 );
not ( w_14521 , w_14522 );
and ( \4540_b0 , \4537_b0 , w_14523 );
and ( w_14522 ,  , w_14523 );
buf ( w_14521 , \4539_b1 );
not ( w_14521 , w_14524 );
not (  , w_14525 );
and ( w_14524 , w_14525 , \4539_b0 );
buf ( \4541_b1 , \4540_b1 );
buf ( \4541_b0 , \4540_b0 );
buf ( \4542_b1 , \4541_b1 );
not ( \4542_b1 , w_14526 );
not ( \4542_b0 , w_14527 );
and ( w_14526 , w_14527 , \4541_b0 );
buf ( \4543_b1 , \4542_b1 );
not ( \4543_b1 , w_14528 );
not ( \4543_b0 , w_14529 );
and ( w_14528 , w_14529 , \4542_b0 );
or ( \4544_b1 , \1395_b1 , w_14530 );
xor ( \4544_b0 , \1395_b0 , w_14532 );
not ( w_14532 , w_14533 );
and ( w_14533 , w_14530 , w_14531 );
buf ( w_14530 , \3432_b1 );
not ( w_14530 , w_14534 );
not ( w_14531 , w_14535 );
and ( w_14534 , w_14535 , \3432_b0 );
buf ( \4545_b1 , \4544_b1 );
buf ( \4545_b0 , \4544_b0 );
buf ( \4546_b1 , \4545_b1 );
not ( \4546_b1 , w_14536 );
not ( \4546_b0 , w_14537 );
and ( w_14536 , w_14537 , \4545_b0 );
or ( \4547_b1 , \4543_b1 , w_14538 );
or ( \4547_b0 , \4543_b0 , \4546_b0 );
not ( \4546_b0 , w_14539 );
and ( w_14539 , w_14538 , \4546_b1 );
buf ( \4548_b1 , \1528_b1 );
buf ( \4548_b0 , \1528_b0 );
or ( \4549_b1 , \4547_b1 , w_14541 );
not ( w_14541 , w_14542 );
and ( \4549_b0 , \4547_b0 , w_14543 );
and ( w_14542 ,  , w_14543 );
buf ( w_14541 , \4548_b1 );
not ( w_14541 , w_14544 );
not (  , w_14545 );
and ( w_14544 , w_14545 , \4548_b0 );
buf ( \4550_b1 , \4549_b1 );
buf ( \4550_b0 , \4549_b0 );
buf ( \4551_b1 , \4550_b1 );
not ( \4551_b1 , w_14546 );
not ( \4551_b0 , w_14547 );
and ( w_14546 , w_14547 , \4550_b0 );
buf ( \4552_b1 , \4044_b1 );
not ( \4552_b1 , w_14548 );
not ( \4552_b0 , w_14549 );
and ( w_14548 , w_14549 , \4044_b0 );
buf ( \4553_b1 , \4069_b1 );
not ( \4553_b1 , w_14550 );
not ( \4553_b0 , w_14551 );
and ( w_14550 , w_14551 , \4069_b0 );
or ( \4554_b1 , \4552_b1 , w_14552 );
or ( \4554_b0 , \4552_b0 , \4553_b0 );
not ( \4553_b0 , w_14553 );
and ( w_14553 , w_14552 , \4553_b1 );
or ( \4555_b1 , \4407_b1 , w_14555 );
not ( w_14555 , w_14556 );
and ( \4555_b0 , \4407_b0 , w_14557 );
and ( w_14556 ,  , w_14557 );
buf ( w_14555 , \4092_b1 );
not ( w_14555 , w_14558 );
not (  , w_14559 );
and ( w_14558 , w_14559 , \4092_b0 );
or ( \4556_b1 , \4554_b1 , w_14561 );
not ( w_14561 , w_14562 );
and ( \4556_b0 , \4554_b0 , w_14563 );
and ( w_14562 ,  , w_14563 );
buf ( w_14561 , \4555_b1 );
not ( w_14561 , w_14564 );
not (  , w_14565 );
and ( w_14564 , w_14565 , \4555_b0 );
buf ( \4557_b1 , \4556_b1 );
not ( \4557_b1 , w_14566 );
not ( \4557_b0 , w_14567 );
and ( w_14566 , w_14567 , \4556_b0 );
or ( \4558_b1 , \4063_b1 , \4053_b1 );
not ( \4053_b1 , w_14568 );
and ( \4558_b0 , \4063_b0 , w_14569 );
and ( w_14568 , w_14569 , \4053_b0 );
buf ( \4559_b1 , \4558_b1 );
not ( \4559_b1 , w_14570 );
not ( \4559_b0 , w_14571 );
and ( w_14570 , w_14571 , \4558_b0 );
or ( \4560_b1 , \4557_b1 , w_14572 );
or ( \4560_b0 , \4557_b0 , \4559_b0 );
not ( \4559_b0 , w_14573 );
and ( w_14573 , w_14572 , \4559_b1 );
buf ( \4561_b1 , \4053_b1 );
buf ( \4561_b0 , \4053_b0 );
buf ( \4562_b1 , \4561_b1 );
not ( \4562_b1 , w_14574 );
not ( \4562_b0 , w_14575 );
and ( w_14574 , w_14575 , \4561_b0 );
or ( \4563_b1 , \4562_b1 , w_14577 );
not ( w_14577 , w_14578 );
and ( \4563_b0 , \4562_b0 , w_14579 );
and ( w_14578 ,  , w_14579 );
buf ( w_14577 , \4409_b1 );
not ( w_14577 , w_14580 );
not (  , w_14581 );
and ( w_14580 , w_14581 , \4409_b0 );
or ( \4564_b1 , \4560_b1 , w_14583 );
not ( w_14583 , w_14584 );
and ( \4564_b0 , \4560_b0 , w_14585 );
and ( w_14584 ,  , w_14585 );
buf ( w_14583 , \4563_b1 );
not ( w_14583 , w_14586 );
not (  , w_14587 );
and ( w_14586 , w_14587 , \4563_b0 );
buf ( \4565_b1 , \4564_b1 );
not ( \4565_b1 , w_14588 );
not ( \4565_b0 , w_14589 );
and ( w_14588 , w_14589 , \4564_b0 );
or ( \4566_b1 , \4551_b1 , w_14590 );
or ( \4566_b0 , \4551_b0 , \4565_b0 );
not ( \4565_b0 , w_14591 );
and ( w_14591 , w_14590 , \4565_b1 );
or ( \4567_b1 , \4550_b1 , w_14592 );
or ( \4567_b0 , \4550_b0 , \4564_b0 );
not ( \4564_b0 , w_14593 );
and ( w_14593 , w_14592 , \4564_b1 );
buf ( \4568_b1 , \4045_b1 );
not ( \4568_b1 , w_14594 );
not ( \4568_b0 , w_14595 );
and ( w_14594 , w_14595 , \4045_b0 );
buf ( \4569_b1 , \4109_b1 );
not ( \4569_b1 , w_14596 );
not ( \4569_b0 , w_14597 );
and ( w_14596 , w_14597 , \4109_b0 );
buf ( \4570_b1 , \4569_b1 );
not ( \4570_b1 , w_14598 );
not ( \4570_b0 , w_14599 );
and ( w_14598 , w_14599 , \4569_b0 );
or ( \4571_b1 , \4568_b1 , w_14600 );
or ( \4571_b0 , \4568_b0 , \4570_b0 );
not ( \4570_b0 , w_14601 );
and ( w_14601 , w_14600 , \4570_b1 );
or ( \4572_b1 , \4109_b1 , w_14603 );
not ( w_14603 , w_14604 );
and ( \4572_b0 , \4109_b0 , w_14605 );
and ( w_14604 ,  , w_14605 );
buf ( w_14603 , \4286_b1 );
not ( w_14603 , w_14606 );
not (  , w_14607 );
and ( w_14606 , w_14607 , \4286_b0 );
or ( \4573_b1 , \4571_b1 , w_14609 );
not ( w_14609 , w_14610 );
and ( \4573_b0 , \4571_b0 , w_14611 );
and ( w_14610 ,  , w_14611 );
buf ( w_14609 , \4572_b1 );
not ( w_14609 , w_14612 );
not (  , w_14613 );
and ( w_14612 , w_14613 , \4572_b0 );
buf ( \4574_b1 , \4573_b1 );
not ( \4574_b1 , w_14614 );
not ( \4574_b0 , w_14615 );
and ( w_14614 , w_14615 , \4573_b0 );
buf ( \4575_b1 , \4136_b1 );
not ( \4575_b1 , w_14616 );
not ( \4575_b0 , w_14617 );
and ( w_14616 , w_14617 , \4136_b0 );
or ( \4576_b1 , \4574_b1 , w_14618 );
or ( \4576_b0 , \4574_b0 , \4575_b0 );
not ( \4575_b0 , w_14619 );
and ( w_14619 , w_14618 , \4575_b1 );
or ( \4577_b1 , \4429_b1 , w_14621 );
not ( w_14621 , w_14622 );
and ( \4577_b0 , \4429_b0 , w_14623 );
and ( w_14622 ,  , w_14623 );
buf ( w_14621 , \4423_b1 );
not ( w_14621 , w_14624 );
not (  , w_14625 );
and ( w_14624 , w_14625 , \4423_b0 );
or ( \4578_b1 , \4576_b1 , w_14627 );
not ( w_14627 , w_14628 );
and ( \4578_b0 , \4576_b0 , w_14629 );
and ( w_14628 ,  , w_14629 );
buf ( w_14627 , \4577_b1 );
not ( w_14627 , w_14630 );
not (  , w_14631 );
and ( w_14630 , w_14631 , \4577_b0 );
or ( \4579_b1 , \4567_b1 , w_14633 );
not ( w_14633 , w_14634 );
and ( \4579_b0 , \4567_b0 , w_14635 );
and ( w_14634 ,  , w_14635 );
buf ( w_14633 , \4578_b1 );
not ( w_14633 , w_14636 );
not (  , w_14637 );
and ( w_14636 , w_14637 , \4578_b0 );
or ( \4580_b1 , \4566_b1 , w_14639 );
not ( w_14639 , w_14640 );
and ( \4580_b0 , \4566_b0 , w_14641 );
and ( w_14640 ,  , w_14641 );
buf ( w_14639 , \4579_b1 );
not ( w_14639 , w_14642 );
not (  , w_14643 );
and ( w_14642 , w_14643 , \4579_b0 );
buf ( \4581_b1 , \4580_b1 );
not ( \4581_b1 , w_14644 );
not ( \4581_b0 , w_14645 );
and ( w_14644 , w_14645 , \4580_b0 );
or ( \4582_b1 , \4581_b1 , w_14647 );
not ( w_14647 , w_14648 );
and ( \4582_b0 , \4581_b0 , w_14649 );
and ( w_14648 ,  , w_14649 );
buf ( w_14647 , \4414_b1 );
not ( w_14647 , w_14650 );
not (  , w_14651 );
and ( w_14650 , w_14651 , \4414_b0 );
buf ( \4583_b1 , \4582_b1 );
not ( \4583_b1 , w_14652 );
not ( \4583_b0 , w_14653 );
and ( w_14652 , w_14653 , \4582_b0 );
buf ( \4584_b1 , \4156_b1 );
not ( \4584_b1 , w_14654 );
not ( \4584_b0 , w_14655 );
and ( w_14654 , w_14655 , \4156_b0 );
buf ( \4585_b1 , \4019_b1 );
not ( \4585_b1 , w_14656 );
not ( \4585_b0 , w_14657 );
and ( w_14656 , w_14657 , \4019_b0 );
or ( \4586_b1 , \4584_b1 , w_14659 );
not ( w_14659 , w_14660 );
and ( \4586_b0 , \4584_b0 , w_14661 );
and ( w_14660 ,  , w_14661 );
buf ( w_14659 , \4585_b1 );
not ( w_14659 , w_14662 );
not (  , w_14663 );
and ( w_14662 , w_14663 , \4585_b0 );
buf ( \4587_b1 , \4586_b1 );
not ( \4587_b1 , w_14664 );
not ( \4587_b0 , w_14665 );
and ( w_14664 , w_14665 , \4586_b0 );
buf ( \4588_b1 , \4042_b1 );
not ( \4588_b1 , w_14666 );
not ( \4588_b0 , w_14667 );
and ( w_14666 , w_14667 , \4042_b0 );
buf ( \4589_b1 , \4089_b1 );
not ( \4589_b1 , w_14668 );
not ( \4589_b0 , w_14669 );
and ( w_14668 , w_14669 , \4089_b0 );
or ( \4590_b1 , \4588_b1 , w_14670 );
or ( \4590_b0 , \4588_b0 , \4589_b0 );
not ( \4589_b0 , w_14671 );
and ( w_14671 , w_14670 , \4589_b1 );
or ( \4591_b1 , \4088_b1 , w_14673 );
not ( w_14673 , w_14674 );
and ( \4591_b0 , \4088_b0 , w_14675 );
and ( w_14674 ,  , w_14675 );
buf ( w_14673 , \4116_b1 );
not ( w_14673 , w_14676 );
not (  , w_14677 );
and ( w_14676 , w_14677 , \4116_b0 );
or ( \4592_b1 , \4590_b1 , w_14679 );
not ( w_14679 , w_14680 );
and ( \4592_b0 , \4590_b0 , w_14681 );
and ( w_14680 ,  , w_14681 );
buf ( w_14679 , \4591_b1 );
not ( w_14679 , w_14682 );
not (  , w_14683 );
and ( w_14682 , w_14683 , \4591_b0 );
buf ( \4593_b1 , \4592_b1 );
not ( \4593_b1 , w_14684 );
not ( \4593_b0 , w_14685 );
and ( w_14684 , w_14685 , \4592_b0 );
buf ( \4594_b1 , \4437_b1 );
not ( \4594_b1 , w_14686 );
not ( \4594_b0 , w_14687 );
and ( w_14686 , w_14687 , \4437_b0 );
or ( \4595_b1 , \4593_b1 , w_14688 );
or ( \4595_b0 , \4593_b0 , \4594_b0 );
not ( \4594_b0 , w_14689 );
and ( w_14689 , w_14688 , \4594_b1 );
buf ( \4596_b1 , \4103_b1 );
not ( \4596_b1 , w_14690 );
not ( \4596_b0 , w_14691 );
and ( w_14690 , w_14691 , \4103_b0 );
or ( \4597_b1 , \4596_b1 , w_14693 );
not ( w_14693 , w_14694 );
and ( \4597_b0 , \4596_b0 , w_14695 );
and ( w_14694 ,  , w_14695 );
buf ( w_14693 , \4435_b1 );
not ( w_14693 , w_14696 );
not (  , w_14697 );
and ( w_14696 , w_14697 , \4435_b0 );
or ( \4598_b1 , \4595_b1 , w_14699 );
not ( w_14699 , w_14700 );
and ( \4598_b0 , \4595_b0 , w_14701 );
and ( w_14700 ,  , w_14701 );
buf ( w_14699 , \4597_b1 );
not ( w_14699 , w_14702 );
not (  , w_14703 );
and ( w_14702 , w_14703 , \4597_b0 );
buf ( \4599_b1 , \4598_b1 );
not ( \4599_b1 , w_14704 );
not ( \4599_b0 , w_14705 );
and ( w_14704 , w_14705 , \4598_b0 );
or ( \4600_b1 , \4587_b1 , w_14706 );
or ( \4600_b0 , \4587_b0 , \4599_b0 );
not ( \4599_b0 , w_14707 );
and ( w_14707 , w_14706 , \4599_b1 );
or ( \4601_b1 , \4598_b1 , w_14708 );
or ( \4601_b0 , \4598_b0 , \4586_b0 );
not ( \4586_b0 , w_14709 );
and ( w_14709 , w_14708 , \4586_b1 );
or ( \4602_b1 , \4043_b1 , \4172_b1 );
not ( \4172_b1 , w_14710 );
and ( \4602_b0 , \4043_b0 , w_14711 );
and ( w_14710 , w_14711 , \4172_b0 );
buf ( \4603_b1 , \4043_b1 );
not ( \4603_b1 , w_14712 );
not ( \4603_b0 , w_14713 );
and ( w_14712 , w_14713 , \4043_b0 );
or ( \4604_b1 , \4603_b1 , \4173_b1 );
not ( \4173_b1 , w_14714 );
and ( \4604_b0 , \4603_b0 , w_14715 );
and ( w_14714 , w_14715 , \4173_b0 );
or ( \4605_b1 , \4602_b1 , w_14717 );
not ( w_14717 , w_14718 );
and ( \4605_b0 , \4602_b0 , w_14719 );
and ( w_14718 ,  , w_14719 );
buf ( w_14717 , \4604_b1 );
not ( w_14717 , w_14720 );
not (  , w_14721 );
and ( w_14720 , w_14721 , \4604_b0 );
buf ( \4606_b1 , \4605_b1 );
not ( \4606_b1 , w_14722 );
not ( \4606_b0 , w_14723 );
and ( w_14722 , w_14723 , \4605_b0 );
buf ( \4607_b1 , \4195_b1 );
not ( \4607_b1 , w_14724 );
not ( \4607_b0 , w_14725 );
and ( w_14724 , w_14725 , \4195_b0 );
or ( \4608_b1 , \4606_b1 , w_14726 );
or ( \4608_b0 , \4606_b0 , \4607_b0 );
not ( \4607_b0 , w_14727 );
and ( w_14727 , w_14726 , \4607_b1 );
or ( \4609_b1 , \4205_b1 , w_14729 );
not ( w_14729 , w_14730 );
and ( \4609_b0 , \4205_b0 , w_14731 );
and ( w_14730 ,  , w_14731 );
buf ( w_14729 , \4446_b1 );
not ( w_14729 , w_14732 );
not (  , w_14733 );
and ( w_14732 , w_14733 , \4446_b0 );
or ( \4610_b1 , \4608_b1 , w_14735 );
not ( w_14735 , w_14736 );
and ( \4610_b0 , \4608_b0 , w_14737 );
and ( w_14736 ,  , w_14737 );
buf ( w_14735 , \4609_b1 );
not ( w_14735 , w_14738 );
not (  , w_14739 );
and ( w_14738 , w_14739 , \4609_b0 );
or ( \4611_b1 , \4601_b1 , w_14741 );
not ( w_14741 , w_14742 );
and ( \4611_b0 , \4601_b0 , w_14743 );
and ( w_14742 ,  , w_14743 );
buf ( w_14741 , \4610_b1 );
not ( w_14741 , w_14744 );
not (  , w_14745 );
and ( w_14744 , w_14745 , \4610_b0 );
or ( \4612_b1 , \4600_b1 , w_14747 );
not ( w_14747 , w_14748 );
and ( \4612_b0 , \4600_b0 , w_14749 );
and ( w_14748 ,  , w_14749 );
buf ( w_14747 , \4611_b1 );
not ( w_14747 , w_14750 );
not (  , w_14751 );
and ( w_14750 , w_14751 , \4611_b0 );
buf ( \4613_b1 , \4612_b1 );
not ( \4613_b1 , w_14752 );
not ( \4613_b0 , w_14753 );
and ( w_14752 , w_14753 , \4612_b0 );
or ( \4614_b1 , \4583_b1 , w_14754 );
or ( \4614_b0 , \4583_b0 , \4613_b0 );
not ( \4613_b0 , w_14755 );
and ( w_14755 , w_14754 , \4613_b1 );
buf ( \4615_b1 , \4414_b1 );
not ( \4615_b1 , w_14756 );
not ( \4615_b0 , w_14757 );
and ( w_14756 , w_14757 , \4414_b0 );
or ( \4616_b1 , \4615_b1 , w_14759 );
not ( w_14759 , w_14760 );
and ( \4616_b0 , \4615_b0 , w_14761 );
and ( w_14760 ,  , w_14761 );
buf ( w_14759 , \4580_b1 );
not ( w_14759 , w_14762 );
not (  , w_14763 );
and ( w_14762 , w_14763 , \4580_b0 );
or ( \4617_b1 , \4614_b1 , w_14765 );
not ( w_14765 , w_14766 );
and ( \4617_b0 , \4614_b0 , w_14767 );
and ( w_14766 ,  , w_14767 );
buf ( w_14765 , \4616_b1 );
not ( w_14765 , w_14768 );
not (  , w_14769 );
and ( w_14768 , w_14769 , \4616_b0 );
buf ( \4618_b1 , \4617_b1 );
not ( \4618_b1 , w_14770 );
not ( \4618_b0 , w_14771 );
and ( w_14770 , w_14771 , \4617_b0 );
buf ( \4619_b1 , \4454_b1 );
not ( \4619_b1 , w_14772 );
not ( \4619_b0 , w_14773 );
and ( w_14772 , w_14773 , \4454_b0 );
or ( \4620_b1 , \4416_b1 , \4414_b1 );
not ( \4414_b1 , w_14774 );
and ( \4620_b0 , \4416_b0 , w_14775 );
and ( w_14774 , w_14775 , \4414_b0 );
buf ( \4621_b1 , \4416_b1 );
not ( \4621_b1 , w_14776 );
not ( \4621_b0 , w_14777 );
and ( w_14776 , w_14777 , \4416_b0 );
or ( \4622_b1 , \4621_b1 , \4413_b1 );
not ( \4413_b1 , w_14778 );
and ( \4622_b0 , \4621_b0 , w_14779 );
and ( w_14778 , w_14779 , \4413_b0 );
or ( \4623_b1 , \4620_b1 , w_14781 );
not ( w_14781 , w_14782 );
and ( \4623_b0 , \4620_b0 , w_14783 );
and ( w_14782 ,  , w_14783 );
buf ( w_14781 , \4622_b1 );
not ( w_14781 , w_14784 );
not (  , w_14785 );
and ( w_14784 , w_14785 , \4622_b0 );
buf ( \4624_b1 , \4623_b1 );
not ( \4624_b1 , w_14786 );
not ( \4624_b0 , w_14787 );
and ( w_14786 , w_14787 , \4623_b0 );
or ( \4625_b1 , \4619_b1 , \4624_b1 );
not ( \4624_b1 , w_14788 );
and ( \4625_b0 , \4619_b0 , w_14789 );
and ( w_14788 , w_14789 , \4624_b0 );
or ( \4626_b1 , \4454_b1 , \4623_b1 );
not ( \4623_b1 , w_14790 );
and ( \4626_b0 , \4454_b0 , w_14791 );
and ( w_14790 , w_14791 , \4623_b0 );
or ( \4627_b1 , \4625_b1 , w_14793 );
not ( w_14793 , w_14794 );
and ( \4627_b0 , \4625_b0 , w_14795 );
and ( w_14794 ,  , w_14795 );
buf ( w_14793 , \4626_b1 );
not ( w_14793 , w_14796 );
not (  , w_14797 );
and ( w_14796 , w_14797 , \4626_b0 );
or ( \4628_b1 , \4618_b1 , w_14799 );
not ( w_14799 , w_14800 );
and ( \4628_b0 , \4618_b0 , w_14801 );
and ( w_14800 ,  , w_14801 );
buf ( w_14799 , \4627_b1 );
not ( w_14799 , w_14802 );
not (  , w_14803 );
and ( w_14802 , w_14803 , \4627_b0 );
buf ( \4629_b1 , \4628_b1 );
not ( \4629_b1 , w_14804 );
not ( \4629_b0 , w_14805 );
and ( w_14804 , w_14805 , \4628_b0 );
or ( \4630_b1 , \4431_b1 , \4441_b1 );
xor ( \4630_b0 , \4431_b0 , w_14806 );
not ( w_14806 , w_14807 );
and ( w_14807 , \4441_b1 , \4441_b0 );
or ( \4631_b1 , \4630_b1 , \4451_b1 );
xor ( \4631_b0 , \4630_b0 , w_14808 );
not ( w_14808 , w_14809 );
and ( w_14809 , \4451_b1 , \4451_b0 );
buf ( \4632_b1 , \4631_b1 );
not ( \4632_b1 , w_14810 );
not ( \4632_b0 , w_14811 );
and ( w_14810 , w_14811 , \4631_b0 );
buf ( \4633_b1 , \4488_b1 );
not ( \4633_b1 , w_14812 );
not ( \4633_b0 , w_14813 );
and ( w_14812 , w_14813 , \4488_b0 );
or ( \4634_b1 , \4633_b1 , w_14815 );
not ( w_14815 , w_14816 );
and ( \4634_b0 , \4633_b0 , w_14817 );
and ( w_14816 ,  , w_14817 );
buf ( w_14815 , \4503_b1 );
not ( w_14815 , w_14818 );
not (  , w_14819 );
and ( w_14818 , w_14819 , \4503_b0 );
or ( \4635_b1 , \4634_b1 , \4500_b1 );
not ( \4500_b1 , w_14820 );
and ( \4635_b0 , \4634_b0 , w_14821 );
and ( w_14820 , w_14821 , \4500_b0 );
buf ( \4636_b1 , \4634_b1 );
not ( \4636_b1 , w_14822 );
not ( \4636_b0 , w_14823 );
and ( w_14822 , w_14823 , \4634_b0 );
or ( \4637_b1 , \4636_b1 , \4501_b1 );
not ( \4501_b1 , w_14824 );
and ( \4637_b0 , \4636_b0 , w_14825 );
and ( w_14824 , w_14825 , \4501_b0 );
or ( \4638_b1 , \4635_b1 , w_14827 );
not ( w_14827 , w_14828 );
and ( \4638_b0 , \4635_b0 , w_14829 );
and ( w_14828 ,  , w_14829 );
buf ( w_14827 , \4637_b1 );
not ( w_14827 , w_14830 );
not (  , w_14831 );
and ( w_14830 , w_14831 , \4637_b0 );
or ( \4639_b1 , \4632_b1 , w_14833 );
not ( w_14833 , w_14834 );
and ( \4639_b0 , \4632_b0 , w_14835 );
and ( w_14834 ,  , w_14835 );
buf ( w_14833 , \4638_b1 );
not ( w_14833 , w_14836 );
not (  , w_14837 );
and ( w_14836 , w_14837 , \4638_b0 );
buf ( \4640_b1 , \3963_b1 );
not ( \4640_b1 , w_14838 );
not ( \4640_b0 , w_14839 );
and ( w_14838 , w_14839 , \3963_b0 );
buf ( \4641_b1 , \4260_b1 );
not ( \4641_b1 , w_14840 );
not ( \4641_b0 , w_14841 );
and ( w_14840 , w_14841 , \4260_b0 );
or ( \4642_b1 , \4640_b1 , w_14842 );
or ( \4642_b0 , \4640_b0 , \4641_b0 );
not ( \4641_b0 , w_14843 );
and ( w_14843 , w_14842 , \4641_b1 );
or ( \4643_b1 , \4156_b1 , w_14845 );
not ( w_14845 , w_14846 );
and ( \4643_b0 , \4156_b0 , w_14847 );
and ( w_14846 ,  , w_14847 );
buf ( w_14845 , \4486_b1 );
not ( w_14845 , w_14848 );
not (  , w_14849 );
and ( w_14848 , w_14849 , \4486_b0 );
or ( \4644_b1 , \4642_b1 , w_14851 );
not ( w_14851 , w_14852 );
and ( \4644_b0 , \4642_b0 , w_14853 );
and ( w_14852 ,  , w_14853 );
buf ( w_14851 , \4643_b1 );
not ( w_14851 , w_14854 );
not (  , w_14855 );
and ( w_14854 , w_14855 , \4643_b0 );
buf ( \4645_b1 , \4644_b1 );
not ( \4645_b1 , w_14856 );
not ( \4645_b0 , w_14857 );
and ( w_14856 , w_14857 , \4644_b0 );
buf ( \4646_b1 , \4253_b1 );
not ( \4646_b1 , w_14858 );
not ( \4646_b0 , w_14859 );
and ( w_14858 , w_14859 , \4253_b0 );
or ( \4647_b1 , \4645_b1 , w_14860 );
or ( \4647_b0 , \4645_b0 , \4646_b0 );
not ( \4646_b0 , w_14861 );
and ( w_14861 , w_14860 , \4646_b1 );
or ( \4648_b1 , \4273_b1 , w_14863 );
not ( w_14863 , w_14864 );
and ( \4648_b0 , \4273_b0 , w_14865 );
and ( w_14864 ,  , w_14865 );
buf ( w_14863 , \4478_b1 );
not ( w_14863 , w_14866 );
not (  , w_14867 );
and ( w_14866 , w_14867 , \4478_b0 );
or ( \4649_b1 , \4647_b1 , w_14869 );
not ( w_14869 , w_14870 );
and ( \4649_b0 , \4647_b0 , w_14871 );
and ( w_14870 ,  , w_14871 );
buf ( w_14869 , \4648_b1 );
not ( w_14869 , w_14872 );
not (  , w_14873 );
and ( w_14872 , w_14873 , \4648_b0 );
buf ( \4650_b1 , \4046_b1 );
not ( \4650_b1 , w_14874 );
not ( \4650_b0 , w_14875 );
and ( w_14874 , w_14875 , \4046_b0 );
buf ( \4651_b1 , \4212_b1 );
not ( \4651_b1 , w_14876 );
not ( \4651_b0 , w_14877 );
and ( w_14876 , w_14877 , \4212_b0 );
or ( \4652_b1 , \4650_b1 , w_14878 );
or ( \4652_b0 , \4650_b0 , \4651_b0 );
not ( \4651_b0 , w_14879 );
and ( w_14879 , w_14878 , \4651_b1 );
or ( \4653_b1 , \4492_b1 , w_14881 );
not ( w_14881 , w_14882 );
and ( \4653_b0 , \4492_b0 , w_14883 );
and ( w_14882 ,  , w_14883 );
buf ( w_14881 , \4256_b1 );
not ( w_14881 , w_14884 );
not (  , w_14885 );
and ( w_14884 , w_14885 , \4256_b0 );
or ( \4654_b1 , \4652_b1 , w_14887 );
not ( w_14887 , w_14888 );
and ( \4654_b0 , \4652_b0 , w_14889 );
and ( w_14888 ,  , w_14889 );
buf ( w_14887 , \4653_b1 );
not ( w_14887 , w_14890 );
not (  , w_14891 );
and ( w_14890 , w_14891 , \4653_b0 );
buf ( \4655_b1 , \4654_b1 );
not ( \4655_b1 , w_14892 );
not ( \4655_b0 , w_14893 );
and ( w_14892 , w_14893 , \4654_b0 );
buf ( \4656_b1 , \4231_b1 );
not ( \4656_b1 , w_14894 );
not ( \4656_b0 , w_14895 );
and ( w_14894 , w_14895 , \4231_b0 );
or ( \4657_b1 , \4655_b1 , w_14896 );
or ( \4657_b0 , \4655_b0 , \4656_b0 );
not ( \4656_b0 , w_14897 );
and ( w_14897 , w_14896 , \4656_b1 );
or ( \4658_b1 , \4234_b1 , w_14899 );
not ( w_14899 , w_14900 );
and ( \4658_b0 , \4234_b0 , w_14901 );
and ( w_14900 ,  , w_14901 );
buf ( w_14899 , \4494_b1 );
not ( w_14899 , w_14902 );
not (  , w_14903 );
and ( w_14902 , w_14903 , \4494_b0 );
or ( \4659_b1 , \4657_b1 , w_14905 );
not ( w_14905 , w_14906 );
and ( \4659_b0 , \4657_b0 , w_14907 );
and ( w_14906 ,  , w_14907 );
buf ( w_14905 , \4658_b1 );
not ( w_14905 , w_14908 );
not (  , w_14909 );
and ( w_14908 , w_14909 , \4658_b0 );
or ( \4660_b1 , \4649_b1 , w_14910 );
or ( \4660_b0 , \4649_b0 , \4659_b0 );
not ( \4659_b0 , w_14911 );
and ( w_14911 , w_14910 , \4659_b1 );
or ( \4661_b1 , \4540_b1 , \4544_b1 );
not ( \4544_b1 , w_14912 );
and ( \4661_b0 , \4540_b0 , w_14913 );
and ( w_14912 , w_14913 , \4544_b0 );
buf ( \4662_b1 , \4661_b1 );
buf ( \4662_b0 , \4661_b0 );
buf ( \4663_b1 , \4662_b1 );
not ( \4663_b1 , w_14914 );
not ( \4663_b0 , w_14915 );
and ( w_14914 , w_14915 , \4662_b0 );
buf ( \4664_b1 , \4663_b1 );
not ( \4664_b1 , w_14916 );
not ( \4664_b0 , w_14917 );
and ( w_14916 , w_14917 , \4663_b0 );
buf ( \4665_b1 , \1528_b1 );
buf ( \4665_b0 , \1528_b0 );
buf ( \4666_b1 , \4665_b1 );
not ( \4666_b1 , w_14918 );
not ( \4666_b0 , w_14919 );
and ( w_14918 , w_14919 , \4665_b0 );
or ( \4667_b1 , \4666_b1 , \3994_b1 );
not ( \3994_b1 , w_14920 );
and ( \4667_b0 , \4666_b0 , w_14921 );
and ( w_14920 , w_14921 , \3994_b0 );
or ( \4668_b1 , \4548_b1 , \4099_b1 );
not ( \4099_b1 , w_14922 );
and ( \4668_b0 , \4548_b0 , w_14923 );
and ( w_14922 , w_14923 , \4099_b0 );
or ( \4669_b1 , \4667_b1 , w_14925 );
not ( w_14925 , w_14926 );
and ( \4669_b0 , \4667_b0 , w_14927 );
and ( w_14926 ,  , w_14927 );
buf ( w_14925 , \4668_b1 );
not ( w_14925 , w_14928 );
not (  , w_14929 );
and ( w_14928 , w_14929 , \4668_b0 );
buf ( \4670_b1 , \4669_b1 );
not ( \4670_b1 , w_14930 );
not ( \4670_b0 , w_14931 );
and ( w_14930 , w_14931 , \4669_b0 );
or ( \4671_b1 , \4664_b1 , \4670_b1 );
not ( \4670_b1 , w_14932 );
and ( \4671_b0 , \4664_b0 , w_14933 );
and ( w_14932 , w_14933 , \4670_b0 );
buf ( \4672_b1 , \4545_b1 );
not ( \4672_b1 , w_14934 );
not ( \4672_b0 , w_14935 );
and ( w_14934 , w_14935 , \4545_b0 );
buf ( \4673_b1 , \4672_b1 );
not ( \4673_b1 , w_14936 );
not ( \4673_b0 , w_14937 );
and ( w_14936 , w_14937 , \4672_b0 );
or ( \4674_b1 , \4673_b1 , w_14939 );
not ( w_14939 , w_14940 );
and ( \4674_b0 , \4673_b0 , w_14941 );
and ( w_14940 ,  , w_14941 );
buf ( w_14939 , \4666_b1 );
not ( w_14939 , w_14942 );
not (  , w_14943 );
and ( w_14942 , w_14943 , \4666_b0 );
or ( \4675_b1 , \4671_b1 , w_14945 );
not ( w_14945 , w_14946 );
and ( \4675_b0 , \4671_b0 , w_14947 );
and ( w_14946 ,  , w_14947 );
buf ( w_14945 , \4674_b1 );
not ( w_14945 , w_14948 );
not (  , w_14949 );
and ( w_14948 , w_14949 , \4674_b0 );
buf ( \4676_b1 , \4675_b1 );
not ( \4676_b1 , w_14950 );
not ( \4676_b0 , w_14951 );
and ( w_14950 , w_14951 , \4675_b0 );
or ( \4677_b1 , \4660_b1 , w_14953 );
not ( w_14953 , w_14954 );
and ( \4677_b0 , \4660_b0 , w_14955 );
and ( w_14954 ,  , w_14955 );
buf ( w_14953 , \4676_b1 );
not ( w_14953 , w_14956 );
not (  , w_14957 );
and ( w_14956 , w_14957 , \4676_b0 );
or ( \4678_b1 , \4659_b1 , w_14959 );
not ( w_14959 , w_14960 );
and ( \4678_b0 , \4659_b0 , w_14961 );
and ( w_14960 ,  , w_14961 );
buf ( w_14959 , \4649_b1 );
not ( w_14959 , w_14962 );
not (  , w_14963 );
and ( w_14962 , w_14963 , \4649_b0 );
or ( \4679_b1 , \4677_b1 , \4678_b1 );
not ( \4678_b1 , w_14964 );
and ( \4679_b0 , \4677_b0 , w_14965 );
and ( w_14964 , w_14965 , \4678_b0 );
buf ( \4680_b1 , \4679_b1 );
not ( \4680_b1 , w_14966 );
not ( \4680_b0 , w_14967 );
and ( w_14966 , w_14967 , \4679_b0 );
or ( \4681_b1 , \4639_b1 , \4680_b1 );
not ( \4680_b1 , w_14968 );
and ( \4681_b0 , \4639_b0 , w_14969 );
and ( w_14968 , w_14969 , \4680_b0 );
buf ( \4682_b1 , \4631_b1 );
not ( \4682_b1 , w_14970 );
not ( \4682_b0 , w_14971 );
and ( w_14970 , w_14971 , \4631_b0 );
or ( \4683_b1 , \4638_b1 , w_14973 );
not ( w_14973 , w_14974 );
and ( \4683_b0 , \4638_b0 , w_14975 );
and ( w_14974 ,  , w_14975 );
buf ( w_14973 , \4682_b1 );
not ( w_14973 , w_14976 );
not (  , w_14977 );
and ( w_14976 , w_14977 , \4682_b0 );
or ( \4684_b1 , \4681_b1 , w_14979 );
not ( w_14979 , w_14980 );
and ( \4684_b0 , \4681_b0 , w_14981 );
and ( w_14980 ,  , w_14981 );
buf ( w_14979 , \4683_b1 );
not ( w_14979 , w_14982 );
not (  , w_14983 );
and ( w_14982 , w_14983 , \4683_b0 );
buf ( \4685_b1 , \4684_b1 );
not ( \4685_b1 , w_14984 );
not ( \4685_b0 , w_14985 );
and ( w_14984 , w_14985 , \4684_b0 );
buf ( \4686_b1 , \4685_b1 );
not ( \4686_b1 , w_14986 );
not ( \4686_b0 , w_14987 );
and ( w_14986 , w_14987 , \4685_b0 );
or ( \4687_b1 , \4629_b1 , w_14988 );
or ( \4687_b0 , \4629_b0 , \4686_b0 );
not ( \4686_b0 , w_14989 );
and ( w_14989 , w_14988 , \4686_b1 );
buf ( \4688_b1 , \4627_b1 );
not ( \4688_b1 , w_14990 );
not ( \4688_b0 , w_14991 );
and ( w_14990 , w_14991 , \4627_b0 );
or ( \4689_b1 , \4688_b1 , w_14993 );
not ( w_14993 , w_14994 );
and ( \4689_b0 , \4688_b0 , w_14995 );
and ( w_14994 ,  , w_14995 );
buf ( w_14993 , \4617_b1 );
not ( w_14993 , w_14996 );
not (  , w_14997 );
and ( w_14996 , w_14997 , \4617_b0 );
or ( \4690_b1 , \4687_b1 , w_14999 );
not ( w_14999 , w_15000 );
and ( \4690_b0 , \4687_b0 , w_15001 );
and ( w_15000 ,  , w_15001 );
buf ( w_14999 , \4689_b1 );
not ( w_14999 , w_15002 );
not (  , w_15003 );
and ( w_15002 , w_15003 , \4689_b0 );
or ( \4691_b1 , \4533_b1 , w_15005 );
not ( w_15005 , w_15006 );
and ( \4691_b0 , \4533_b0 , w_15007 );
and ( w_15006 ,  , w_15007 );
buf ( w_15005 , \4690_b1 );
not ( w_15005 , w_15008 );
not (  , w_15009 );
and ( w_15008 , w_15009 , \4690_b0 );
or ( \4692_b1 , \4532_b1 , w_15011 );
not ( w_15011 , w_15012 );
and ( \4692_b0 , \4532_b0 , w_15013 );
and ( w_15012 ,  , w_15013 );
buf ( w_15011 , \4691_b1 );
not ( w_15011 , w_15014 );
not (  , w_15015 );
and ( w_15014 , w_15015 , \4691_b0 );
buf ( \4693_b1 , \4692_b1 );
not ( \4693_b1 , w_15016 );
not ( \4693_b0 , w_15017 );
and ( w_15016 , w_15017 , \4692_b0 );
or ( \4694_b1 , \4516_b1 , w_15019 );
not ( w_15019 , w_15020 );
and ( \4694_b0 , \4516_b0 , w_15021 );
and ( w_15020 ,  , w_15021 );
buf ( w_15019 , \4693_b1 );
not ( w_15019 , w_15022 );
not (  , w_15023 );
and ( w_15022 , w_15023 , \4693_b0 );
or ( \4695_b1 , \4298_b1 , \4387_b1 );
xor ( \4695_b0 , \4298_b0 , w_15024 );
not ( w_15024 , w_15025 );
and ( w_15025 , \4387_b1 , \4387_b0 );
or ( \4696_b1 , \4695_b1 , \4514_b1 );
not ( \4514_b1 , w_15026 );
and ( \4696_b0 , \4695_b0 , w_15027 );
and ( w_15026 , w_15027 , \4514_b0 );
or ( \4697_b1 , \4298_b1 , \4387_b1 );
not ( \4387_b1 , w_15028 );
and ( \4697_b0 , \4298_b0 , w_15029 );
and ( w_15028 , w_15029 , \4387_b0 );
or ( \4698_b1 , \4696_b1 , w_15030 );
or ( \4698_b0 , \4696_b0 , \4697_b0 );
not ( \4697_b0 , w_15031 );
and ( w_15031 , w_15030 , \4697_b1 );
buf ( \4699_b1 , \4698_b1 );
not ( \4699_b1 , w_15032 );
not ( \4699_b0 , w_15033 );
and ( w_15032 , w_15033 , \4698_b0 );
buf ( \4700_b1 , \4382_b1 );
not ( \4700_b1 , w_15034 );
not ( \4700_b0 , w_15035 );
and ( w_15034 , w_15035 , \4382_b0 );
buf ( \4701_b1 , \4496_b1 );
not ( \4701_b1 , w_15036 );
not ( \4701_b0 , w_15037 );
and ( w_15036 , w_15037 , \4496_b0 );
or ( \4702_b1 , \4700_b1 , w_15038 );
or ( \4702_b0 , \4700_b0 , \4701_b0 );
not ( \4701_b0 , w_15039 );
and ( w_15039 , w_15038 , \4701_b1 );
buf ( \4703_b1 , \4042_b1 );
not ( \4703_b1 , w_15040 );
not ( \4703_b0 , w_15041 );
and ( w_15040 , w_15041 , \4042_b0 );
buf ( \4704_b1 , \4212_b1 );
not ( \4704_b1 , w_15042 );
not ( \4704_b0 , w_15043 );
and ( w_15042 , w_15043 , \4212_b0 );
or ( \4705_b1 , \4703_b1 , w_15044 );
or ( \4705_b0 , \4703_b0 , \4704_b0 );
not ( \4704_b0 , w_15045 );
and ( w_15045 , w_15044 , \4704_b1 );
or ( \4706_b1 , \4216_b1 , w_15047 );
not ( w_15047 , w_15048 );
and ( \4706_b0 , \4216_b0 , w_15049 );
and ( w_15048 ,  , w_15049 );
buf ( w_15047 , \4116_b1 );
not ( w_15047 , w_15050 );
not (  , w_15051 );
and ( w_15050 , w_15051 , \4116_b0 );
or ( \4707_b1 , \4705_b1 , w_15053 );
not ( w_15053 , w_15054 );
and ( \4707_b0 , \4705_b0 , w_15055 );
and ( w_15054 ,  , w_15055 );
buf ( w_15053 , \4706_b1 );
not ( w_15053 , w_15056 );
not (  , w_15057 );
and ( w_15056 , w_15057 , \4706_b0 );
or ( \4708_b1 , \4377_b1 , w_15059 );
not ( w_15059 , w_15060 );
and ( \4708_b0 , \4377_b0 , w_15061 );
and ( w_15060 ,  , w_15061 );
buf ( w_15059 , \4707_b1 );
not ( w_15059 , w_15062 );
not (  , w_15063 );
and ( w_15062 , w_15063 , \4707_b0 );
or ( \4709_b1 , \4702_b1 , w_15065 );
not ( w_15065 , w_15066 );
and ( \4709_b0 , \4702_b0 , w_15067 );
and ( w_15066 ,  , w_15067 );
buf ( w_15065 , \4708_b1 );
not ( w_15065 , w_15068 );
not (  , w_15069 );
and ( w_15068 , w_15069 , \4708_b0 );
buf ( \4710_b1 , \4370_b1 );
not ( \4710_b1 , w_15070 );
not ( \4710_b0 , w_15071 );
and ( w_15070 , w_15071 , \4370_b0 );
buf ( \4711_b1 , \4136_b1 );
not ( \4711_b1 , w_15072 );
not ( \4711_b0 , w_15073 );
and ( w_15072 , w_15073 , \4136_b0 );
or ( \4712_b1 , \4710_b1 , w_15074 );
or ( \4712_b0 , \4710_b0 , \4711_b0 );
not ( \4711_b0 , w_15075 );
and ( w_15075 , w_15074 , \4711_b1 );
buf ( \4713_b1 , \4110_b1 );
not ( \4713_b1 , w_15076 );
not ( \4713_b0 , w_15077 );
and ( w_15076 , w_15077 , \4110_b0 );
or ( \4714_b1 , \4713_b1 , w_15079 );
not ( w_15079 , w_15080 );
and ( \4714_b0 , \4713_b0 , w_15081 );
and ( w_15080 ,  , w_15081 );
buf ( w_15079 , \4140_b1 );
not ( w_15079 , w_15082 );
not (  , w_15083 );
and ( w_15082 , w_15083 , \4140_b0 );
or ( \4715_b1 , \4712_b1 , w_15085 );
not ( w_15085 , w_15086 );
and ( \4715_b0 , \4712_b0 , w_15087 );
and ( w_15086 ,  , w_15087 );
buf ( w_15085 , \4714_b1 );
not ( w_15085 , w_15088 );
not (  , w_15089 );
and ( w_15088 , w_15089 , \4714_b0 );
buf ( \4716_b1 , \4715_b1 );
not ( \4716_b1 , w_15090 );
not ( \4716_b0 , w_15091 );
and ( w_15090 , w_15091 , \4715_b0 );
or ( \4717_b1 , \4709_b1 , \4716_b1 );
xor ( \4717_b0 , \4709_b0 , w_15092 );
not ( w_15092 , w_15093 );
and ( w_15093 , \4716_b1 , \4716_b0 );
or ( \4718_b1 , \4307_b1 , \4315_b1 );
xor ( \4718_b0 , \4307_b0 , w_15094 );
not ( w_15094 , w_15095 );
and ( w_15095 , \4315_b1 , \4315_b0 );
or ( \4719_b1 , \4718_b1 , \4325_b1 );
not ( \4325_b1 , w_15096 );
and ( \4719_b0 , \4718_b0 , w_15097 );
and ( w_15096 , w_15097 , \4325_b0 );
or ( \4720_b1 , \4307_b1 , \4315_b1 );
not ( \4315_b1 , w_15098 );
and ( \4720_b0 , \4307_b0 , w_15099 );
and ( w_15098 , w_15099 , \4315_b0 );
or ( \4721_b1 , \4719_b1 , w_15100 );
or ( \4721_b0 , \4719_b0 , \4720_b0 );
not ( \4720_b0 , w_15101 );
and ( w_15101 , w_15100 , \4720_b1 );
or ( \4722_b1 , \4717_b1 , \4721_b1 );
xor ( \4722_b0 , \4717_b0 , w_15102 );
not ( w_15102 , w_15103 );
and ( w_15103 , \4721_b1 , \4721_b0 );
buf ( \4723_b1 , \4386_b1 );
not ( \4723_b1 , w_15104 );
not ( \4723_b0 , w_15105 );
and ( w_15104 , w_15105 , \4386_b0 );
buf ( \4724_b1 , \4326_b1 );
not ( \4724_b1 , w_15106 );
not ( \4724_b0 , w_15107 );
and ( w_15106 , w_15107 , \4326_b0 );
or ( \4725_b1 , \4724_b1 , w_15109 );
not ( w_15109 , w_15110 );
and ( \4725_b0 , \4724_b0 , w_15111 );
and ( w_15110 ,  , w_15111 );
buf ( w_15109 , \4306_b1 );
not ( w_15109 , w_15112 );
not (  , w_15113 );
and ( w_15112 , w_15113 , \4306_b0 );
buf ( \4726_b1 , \4725_b1 );
not ( \4726_b1 , w_15114 );
not ( \4726_b0 , w_15115 );
and ( w_15114 , w_15115 , \4725_b0 );
or ( \4727_b1 , \4723_b1 , w_15116 );
or ( \4727_b0 , \4723_b0 , \4726_b0 );
not ( \4726_b0 , w_15117 );
and ( w_15117 , w_15116 , \4726_b1 );
or ( \4728_b1 , \4326_b1 , w_15119 );
not ( w_15119 , w_15120 );
and ( \4728_b0 , \4326_b0 , w_15121 );
and ( w_15120 ,  , w_15121 );
buf ( w_15119 , \4305_b1 );
not ( w_15119 , w_15122 );
not (  , w_15123 );
and ( w_15122 , w_15123 , \4305_b0 );
or ( \4729_b1 , \4727_b1 , w_15125 );
not ( w_15125 , w_15126 );
and ( \4729_b0 , \4727_b0 , w_15127 );
and ( w_15126 ,  , w_15127 );
buf ( w_15125 , \4728_b1 );
not ( w_15125 , w_15128 );
not (  , w_15129 );
and ( w_15128 , w_15129 , \4728_b0 );
or ( \4730_b1 , \4722_b1 , \4729_b1 );
xor ( \4730_b0 , \4722_b0 , w_15130 );
not ( w_15130 , w_15131 );
and ( w_15131 , \4729_b1 , \4729_b0 );
buf ( \4731_b1 , \4372_b1 );
not ( \4731_b1 , w_15132 );
not ( \4731_b0 , w_15133 );
and ( w_15132 , w_15133 , \4372_b0 );
or ( \4732_b1 , \4731_b1 , w_15135 );
not ( w_15135 , w_15136 );
and ( \4732_b0 , \4731_b0 , w_15137 );
and ( w_15136 ,  , w_15137 );
buf ( w_15135 , \4361_b1 );
not ( w_15135 , w_15138 );
not (  , w_15139 );
and ( w_15138 , w_15139 , \4361_b0 );
or ( \4733_b1 , \4732_b1 , w_15141 );
not ( w_15141 , w_15142 );
and ( \4733_b0 , \4732_b0 , w_15143 );
and ( w_15142 ,  , w_15143 );
buf ( w_15141 , \4384_b1 );
not ( w_15141 , w_15144 );
not (  , w_15145 );
and ( w_15144 , w_15145 , \4384_b0 );
buf ( \4734_b1 , \4361_b1 );
not ( \4734_b1 , w_15146 );
not ( \4734_b0 , w_15147 );
and ( w_15146 , w_15147 , \4361_b0 );
or ( \4735_b1 , \4734_b1 , w_15149 );
not ( w_15149 , w_15150 );
and ( \4735_b0 , \4734_b0 , w_15151 );
and ( w_15150 ,  , w_15151 );
buf ( w_15149 , \4372_b1 );
not ( w_15149 , w_15152 );
not (  , w_15153 );
and ( w_15152 , w_15153 , \4372_b0 );
or ( \4736_b1 , \4733_b1 , \4735_b1 );
not ( \4735_b1 , w_15154 );
and ( \4736_b0 , \4733_b0 , w_15155 );
and ( w_15154 , w_15155 , \4735_b0 );
or ( \4737_b1 , \4043_b1 , \4308_b1 );
not ( \4308_b1 , w_15156 );
and ( \4737_b0 , \4043_b0 , w_15157 );
and ( w_15156 , w_15157 , \4308_b0 );
buf ( \4738_b1 , \4313_b1 );
not ( \4738_b1 , w_15158 );
not ( \4738_b0 , w_15159 );
and ( w_15158 , w_15159 , \4313_b0 );
buf ( \4739_b1 , \4253_b1 );
not ( \4739_b1 , w_15160 );
not ( \4739_b0 , w_15161 );
and ( w_15160 , w_15161 , \4253_b0 );
or ( \4740_b1 , \4738_b1 , w_15162 );
or ( \4740_b0 , \4738_b0 , \4739_b0 );
not ( \4739_b0 , w_15163 );
and ( w_15163 , w_15162 , \4739_b1 );
or ( \4741_b1 , \4045_b1 , \4156_b1 );
xor ( \4741_b0 , \4045_b0 , w_15164 );
not ( w_15164 , w_15165 );
and ( w_15165 , \4156_b1 , \4156_b0 );
buf ( \4742_b1 , \4273_b1 );
buf ( \4742_b0 , \4273_b0 );
or ( \4743_b1 , \4741_b1 , w_15167 );
not ( w_15167 , w_15168 );
and ( \4743_b0 , \4741_b0 , w_15169 );
and ( w_15168 ,  , w_15169 );
buf ( w_15167 , \4742_b1 );
not ( w_15167 , w_15170 );
not (  , w_15171 );
and ( w_15170 , w_15171 , \4742_b0 );
or ( \4744_b1 , \4740_b1 , w_15173 );
not ( w_15173 , w_15174 );
and ( \4744_b0 , \4740_b0 , w_15175 );
and ( w_15174 ,  , w_15175 );
buf ( w_15173 , \4743_b1 );
not ( w_15173 , w_15176 );
not (  , w_15177 );
and ( w_15176 , w_15177 , \4743_b0 );
or ( \4745_b1 , \4737_b1 , \4744_b1 );
xor ( \4745_b0 , \4737_b0 , w_15178 );
not ( w_15178 , w_15179 );
and ( w_15179 , \4744_b1 , \4744_b0 );
buf ( \4746_b1 , \4323_b1 );
not ( \4746_b1 , w_15180 );
not ( \4746_b0 , w_15181 );
and ( w_15180 , w_15181 , \4323_b0 );
buf ( \4747_b1 , \4746_b1 );
not ( \4747_b1 , w_15182 );
not ( \4747_b0 , w_15183 );
and ( w_15182 , w_15183 , \4746_b0 );
buf ( \4748_b1 , \4195_b1 );
not ( \4748_b1 , w_15184 );
not ( \4748_b0 , w_15185 );
and ( w_15184 , w_15185 , \4195_b0 );
or ( \4749_b1 , \4747_b1 , w_15186 );
or ( \4749_b0 , \4747_b0 , \4748_b0 );
not ( \4748_b0 , w_15187 );
and ( w_15187 , w_15186 , \4748_b1 );
buf ( \4750_b1 , \4044_b1 );
not ( \4750_b1 , w_15188 );
not ( \4750_b0 , w_15189 );
and ( w_15188 , w_15189 , \4044_b0 );
buf ( \4751_b1 , \4173_b1 );
not ( \4751_b1 , w_15190 );
not ( \4751_b0 , w_15191 );
and ( w_15190 , w_15191 , \4173_b0 );
or ( \4752_b1 , \4750_b1 , w_15192 );
or ( \4752_b0 , \4750_b0 , \4751_b0 );
not ( \4751_b0 , w_15193 );
and ( w_15193 , w_15192 , \4751_b1 );
or ( \4753_b1 , \4172_b1 , w_15195 );
not ( w_15195 , w_15196 );
and ( \4753_b0 , \4172_b0 , w_15197 );
and ( w_15196 ,  , w_15197 );
buf ( w_15195 , \4092_b1 );
not ( w_15195 , w_15198 );
not (  , w_15199 );
and ( w_15198 , w_15199 , \4092_b0 );
or ( \4754_b1 , \4752_b1 , w_15201 );
not ( w_15201 , w_15202 );
and ( \4754_b0 , \4752_b0 , w_15203 );
and ( w_15202 ,  , w_15203 );
buf ( w_15201 , \4753_b1 );
not ( w_15201 , w_15204 );
not (  , w_15205 );
and ( w_15204 , w_15205 , \4753_b0 );
or ( \4755_b1 , \4205_b1 , w_15207 );
not ( w_15207 , w_15208 );
and ( \4755_b0 , \4205_b0 , w_15209 );
and ( w_15208 ,  , w_15209 );
buf ( w_15207 , \4754_b1 );
not ( w_15207 , w_15210 );
not (  , w_15211 );
and ( w_15210 , w_15211 , \4754_b0 );
or ( \4756_b1 , \4749_b1 , w_15213 );
not ( w_15213 , w_15214 );
and ( \4756_b0 , \4749_b0 , w_15215 );
and ( w_15214 ,  , w_15215 );
buf ( w_15213 , \4755_b1 );
not ( w_15213 , w_15216 );
not (  , w_15217 );
and ( w_15216 , w_15217 , \4755_b0 );
or ( \4757_b1 , \4745_b1 , \4756_b1 );
xor ( \4757_b0 , \4745_b0 , w_15218 );
not ( w_15218 , w_15219 );
and ( w_15219 , \4756_b1 , \4756_b0 );
or ( \4758_b1 , \4736_b1 , \4757_b1 );
xor ( \4758_b0 , \4736_b0 , w_15220 );
not ( w_15220 , w_15221 );
and ( w_15221 , \4757_b1 , \4757_b0 );
or ( \4759_b1 , \4385_b1 , w_15222 );
or ( \4759_b0 , \4385_b0 , \4167_b0 );
not ( \4167_b0 , w_15223 );
and ( w_15223 , w_15222 , \4167_b1 );
or ( \4760_b1 , \4759_b1 , w_15225 );
not ( w_15225 , w_15226 );
and ( \4760_b0 , \4759_b0 , w_15227 );
and ( w_15226 ,  , w_15227 );
buf ( w_15225 , \4354_b1 );
not ( w_15225 , w_15228 );
not (  , w_15229 );
and ( w_15228 , w_15229 , \4354_b0 );
or ( \4761_b1 , \4385_b1 , w_15231 );
not ( w_15231 , w_15232 );
and ( \4761_b0 , \4385_b0 , w_15233 );
and ( w_15232 ,  , w_15233 );
buf ( w_15231 , \4167_b1 );
not ( w_15231 , w_15234 );
not (  , w_15235 );
and ( w_15234 , w_15235 , \4167_b0 );
or ( \4762_b1 , \4760_b1 , w_15237 );
not ( w_15237 , w_15238 );
and ( \4762_b0 , \4760_b0 , w_15239 );
and ( w_15238 ,  , w_15239 );
buf ( w_15237 , \4761_b1 );
not ( w_15237 , w_15240 );
not (  , w_15241 );
and ( w_15240 , w_15241 , \4761_b0 );
or ( \4763_b1 , \4758_b1 , w_15242 );
xor ( \4763_b0 , \4758_b0 , w_15244 );
not ( w_15244 , w_15245 );
and ( w_15245 , w_15242 , w_15243 );
buf ( w_15242 , \4762_b1 );
not ( w_15242 , w_15246 );
not ( w_15243 , w_15247 );
and ( w_15246 , w_15247 , \4762_b0 );
or ( \4764_b1 , \4730_b1 , \4763_b1 );
xor ( \4764_b0 , \4730_b0 , w_15248 );
not ( w_15248 , w_15249 );
and ( w_15249 , \4763_b1 , \4763_b0 );
buf ( \4765_b1 , \4764_b1 );
not ( \4765_b1 , w_15250 );
not ( \4765_b0 , w_15251 );
and ( w_15250 , w_15251 , \4764_b0 );
or ( \4766_b1 , \4699_b1 , w_15253 );
not ( w_15253 , w_15254 );
and ( \4766_b0 , \4699_b0 , w_15255 );
and ( w_15254 ,  , w_15255 );
buf ( w_15253 , \4765_b1 );
not ( w_15253 , w_15256 );
not (  , w_15257 );
and ( w_15256 , w_15257 , \4765_b0 );
or ( \4767_b1 , \4694_b1 , w_15259 );
not ( w_15259 , w_15260 );
and ( \4767_b0 , \4694_b0 , w_15261 );
and ( w_15260 ,  , w_15261 );
buf ( w_15259 , \4766_b1 );
not ( w_15259 , w_15262 );
not (  , w_15263 );
and ( w_15262 , w_15263 , \4766_b0 );
or ( \4768_b1 , \4722_b1 , \4729_b1 );
xor ( \4768_b0 , \4722_b0 , w_15264 );
not ( w_15264 , w_15265 );
and ( w_15265 , \4729_b1 , \4729_b0 );
or ( \4769_b1 , \4768_b1 , \4763_b1 );
not ( \4763_b1 , w_15266 );
and ( \4769_b0 , \4768_b0 , w_15267 );
and ( w_15266 , w_15267 , \4763_b0 );
or ( \4770_b1 , \4722_b1 , \4729_b1 );
not ( \4729_b1 , w_15268 );
and ( \4770_b0 , \4722_b0 , w_15269 );
and ( w_15268 , w_15269 , \4729_b0 );
or ( \4771_b1 , \4769_b1 , w_15270 );
or ( \4771_b0 , \4769_b0 , \4770_b0 );
not ( \4770_b0 , w_15271 );
and ( w_15271 , w_15270 , \4770_b1 );
buf ( \4772_b1 , \4771_b1 );
not ( \4772_b1 , w_15272 );
not ( \4772_b0 , w_15273 );
and ( w_15272 , w_15273 , \4771_b0 );
or ( \4773_b1 , \4709_b1 , \4716_b1 );
xor ( \4773_b0 , \4709_b0 , w_15274 );
not ( w_15274 , w_15275 );
and ( w_15275 , \4716_b1 , \4716_b0 );
or ( \4774_b1 , \4773_b1 , \4721_b1 );
not ( \4721_b1 , w_15276 );
and ( \4774_b0 , \4773_b0 , w_15277 );
and ( w_15276 , w_15277 , \4721_b0 );
or ( \4775_b1 , \4709_b1 , \4716_b1 );
not ( \4716_b1 , w_15278 );
and ( \4775_b0 , \4709_b0 , w_15279 );
and ( w_15278 , w_15279 , \4716_b0 );
or ( \4776_b1 , \4774_b1 , w_15280 );
or ( \4776_b0 , \4774_b0 , \4775_b0 );
not ( \4775_b0 , w_15281 );
and ( w_15281 , w_15280 , \4775_b1 );
or ( \4777_b1 , \4041_b1 , \4156_b1 );
not ( \4156_b1 , w_15282 );
and ( \4777_b0 , \4041_b0 , w_15283 );
and ( w_15282 , w_15283 , \4156_b0 );
or ( \4778_b1 , \4777_b1 , \4715_b1 );
xor ( \4778_b0 , \4777_b0 , w_15284 );
not ( w_15284 , w_15285 );
and ( w_15285 , \4715_b1 , \4715_b0 );
buf ( \4779_b1 , \4707_b1 );
not ( \4779_b1 , w_15286 );
not ( \4779_b0 , w_15287 );
and ( w_15286 , w_15287 , \4707_b0 );
buf ( \4780_b1 , \4496_b1 );
not ( \4780_b1 , w_15288 );
not ( \4780_b0 , w_15289 );
and ( w_15288 , w_15289 , \4496_b0 );
or ( \4781_b1 , \4779_b1 , w_15290 );
or ( \4781_b0 , \4779_b0 , \4780_b0 );
not ( \4780_b0 , w_15291 );
and ( w_15291 , w_15290 , \4780_b1 );
buf ( \4782_b1 , \3943_b1 );
not ( \4782_b1 , w_15292 );
not ( \4782_b0 , w_15293 );
and ( w_15292 , w_15293 , \3943_b0 );
buf ( \4783_b1 , \4212_b1 );
not ( \4783_b1 , w_15294 );
not ( \4783_b0 , w_15295 );
and ( w_15294 , w_15295 , \4212_b0 );
or ( \4784_b1 , \4782_b1 , w_15296 );
or ( \4784_b0 , \4782_b0 , \4783_b0 );
not ( \4783_b0 , w_15297 );
and ( w_15297 , w_15296 , \4783_b1 );
or ( \4785_b1 , \4216_b1 , w_15299 );
not ( w_15299 , w_15300 );
and ( \4785_b0 , \4216_b0 , w_15301 );
and ( w_15300 ,  , w_15301 );
buf ( w_15299 , \4147_b1 );
not ( w_15299 , w_15302 );
not (  , w_15303 );
and ( w_15302 , w_15303 , \4147_b0 );
or ( \4786_b1 , \4784_b1 , w_15305 );
not ( w_15305 , w_15306 );
and ( \4786_b0 , \4784_b0 , w_15307 );
and ( w_15306 ,  , w_15307 );
buf ( w_15305 , \4785_b1 );
not ( w_15305 , w_15308 );
not (  , w_15309 );
and ( w_15308 , w_15309 , \4785_b0 );
or ( \4787_b1 , \4377_b1 , w_15311 );
not ( w_15311 , w_15312 );
and ( \4787_b0 , \4377_b0 , w_15313 );
and ( w_15312 ,  , w_15313 );
buf ( w_15311 , \4786_b1 );
not ( w_15311 , w_15314 );
not (  , w_15315 );
and ( w_15314 , w_15315 , \4786_b0 );
or ( \4788_b1 , \4781_b1 , w_15317 );
not ( w_15317 , w_15318 );
and ( \4788_b0 , \4781_b0 , w_15319 );
and ( w_15318 ,  , w_15319 );
buf ( w_15317 , \4787_b1 );
not ( w_15317 , w_15320 );
not (  , w_15321 );
and ( w_15320 , w_15321 , \4787_b0 );
or ( \4789_b1 , \4778_b1 , \4788_b1 );
xor ( \4789_b0 , \4778_b0 , w_15322 );
not ( w_15322 , w_15323 );
and ( w_15323 , \4788_b1 , \4788_b0 );
or ( \4790_b1 , \4737_b1 , \4744_b1 );
xor ( \4790_b0 , \4737_b0 , w_15324 );
not ( w_15324 , w_15325 );
and ( w_15325 , \4744_b1 , \4744_b0 );
or ( \4791_b1 , \4790_b1 , \4756_b1 );
not ( \4756_b1 , w_15326 );
and ( \4791_b0 , \4790_b0 , w_15327 );
and ( w_15326 , w_15327 , \4756_b0 );
or ( \4792_b1 , \4737_b1 , \4744_b1 );
not ( \4744_b1 , w_15328 );
and ( \4792_b0 , \4737_b0 , w_15329 );
and ( w_15328 , w_15329 , \4744_b0 );
or ( \4793_b1 , \4791_b1 , w_15330 );
or ( \4793_b0 , \4791_b0 , \4792_b0 );
not ( \4792_b0 , w_15331 );
and ( w_15331 , w_15330 , \4792_b1 );
or ( \4794_b1 , \4789_b1 , \4793_b1 );
xor ( \4794_b0 , \4789_b0 , w_15332 );
not ( w_15332 , w_15333 );
and ( w_15333 , \4793_b1 , \4793_b0 );
buf ( \4795_b1 , \4754_b1 );
not ( \4795_b1 , w_15334 );
not ( \4795_b0 , w_15335 );
and ( w_15334 , w_15335 , \4754_b0 );
buf ( \4796_b1 , \4195_b1 );
not ( \4796_b1 , w_15336 );
not ( \4796_b0 , w_15337 );
and ( w_15336 , w_15337 , \4195_b0 );
or ( \4797_b1 , \4795_b1 , w_15338 );
or ( \4797_b0 , \4795_b0 , \4796_b0 );
not ( \4796_b0 , w_15339 );
and ( w_15339 , w_15338 , \4796_b1 );
buf ( \4798_b1 , \3994_b1 );
not ( \4798_b1 , w_15340 );
not ( \4798_b0 , w_15341 );
and ( w_15340 , w_15341 , \3994_b0 );
buf ( \4799_b1 , \4173_b1 );
not ( \4799_b1 , w_15342 );
not ( \4799_b0 , w_15343 );
and ( w_15342 , w_15343 , \4173_b0 );
or ( \4800_b1 , \4798_b1 , w_15344 );
or ( \4800_b0 , \4798_b0 , \4799_b0 );
not ( \4799_b0 , w_15345 );
and ( w_15345 , w_15344 , \4799_b1 );
or ( \4801_b1 , \4172_b1 , w_15347 );
not ( w_15347 , w_15348 );
and ( \4801_b0 , \4172_b0 , w_15349 );
and ( w_15348 ,  , w_15349 );
buf ( w_15347 , \4099_b1 );
not ( w_15347 , w_15350 );
not (  , w_15351 );
and ( w_15350 , w_15351 , \4099_b0 );
or ( \4802_b1 , \4800_b1 , w_15353 );
not ( w_15353 , w_15354 );
and ( \4802_b0 , \4800_b0 , w_15355 );
and ( w_15354 ,  , w_15355 );
buf ( w_15353 , \4801_b1 );
not ( w_15353 , w_15356 );
not (  , w_15357 );
and ( w_15356 , w_15357 , \4801_b0 );
or ( \4803_b1 , \4802_b1 , w_15359 );
not ( w_15359 , w_15360 );
and ( \4803_b0 , \4802_b0 , w_15361 );
and ( w_15360 ,  , w_15361 );
buf ( w_15359 , \4205_b1 );
not ( w_15359 , w_15362 );
not (  , w_15363 );
and ( w_15362 , w_15363 , \4205_b0 );
or ( \4804_b1 , \4797_b1 , w_15365 );
not ( w_15365 , w_15366 );
and ( \4804_b0 , \4797_b0 , w_15367 );
and ( w_15366 ,  , w_15367 );
buf ( w_15365 , \4803_b1 );
not ( w_15365 , w_15368 );
not (  , w_15369 );
and ( w_15368 , w_15369 , \4803_b0 );
buf ( \4805_b1 , \4136_b1 );
not ( \4805_b1 , w_15370 );
not ( \4805_b0 , w_15371 );
and ( w_15370 , w_15371 , \4136_b0 );
buf ( \4806_b1 , \4140_b1 );
not ( \4806_b1 , w_15372 );
not ( \4806_b0 , w_15373 );
and ( w_15372 , w_15373 , \4140_b0 );
or ( \4807_b1 , \4805_b1 , \4806_b1 );
not ( \4806_b1 , w_15374 );
and ( \4807_b0 , \4805_b0 , w_15375 );
and ( w_15374 , w_15375 , \4806_b0 );
or ( \4808_b1 , \4807_b1 , w_15377 );
not ( w_15377 , w_15378 );
and ( \4808_b0 , \4807_b0 , w_15379 );
and ( w_15378 ,  , w_15379 );
buf ( w_15377 , \4110_b1 );
not ( w_15377 , w_15380 );
not (  , w_15381 );
and ( w_15380 , w_15381 , \4110_b0 );
buf ( \4809_b1 , \4808_b1 );
not ( \4809_b1 , w_15382 );
not ( \4809_b0 , w_15383 );
and ( w_15382 , w_15383 , \4808_b0 );
or ( \4810_b1 , \4804_b1 , \4809_b1 );
not ( \4809_b1 , w_15384 );
and ( \4810_b0 , \4804_b0 , w_15385 );
and ( w_15384 , w_15385 , \4809_b0 );
buf ( \4811_b1 , \4804_b1 );
not ( \4811_b1 , w_15386 );
not ( \4811_b0 , w_15387 );
and ( w_15386 , w_15387 , \4804_b0 );
or ( \4812_b1 , \4811_b1 , \4808_b1 );
not ( \4808_b1 , w_15388 );
and ( \4812_b0 , \4811_b0 , w_15389 );
and ( w_15388 , w_15389 , \4808_b0 );
or ( \4813_b1 , \4810_b1 , w_15391 );
not ( w_15391 , w_15392 );
and ( \4813_b0 , \4810_b0 , w_15393 );
and ( w_15392 ,  , w_15393 );
buf ( w_15391 , \4812_b1 );
not ( w_15391 , w_15394 );
not (  , w_15395 );
and ( w_15394 , w_15395 , \4812_b0 );
buf ( \4814_b1 , \4741_b1 );
not ( \4814_b1 , w_15396 );
not ( \4814_b0 , w_15397 );
and ( w_15396 , w_15397 , \4741_b0 );
buf ( \4815_b1 , \4254_b1 );
not ( \4815_b1 , w_15398 );
not ( \4815_b0 , w_15399 );
and ( w_15398 , w_15399 , \4254_b0 );
buf ( \4816_b1 , \4815_b1 );
not ( \4816_b1 , w_15400 );
not ( \4816_b0 , w_15401 );
and ( w_15400 , w_15401 , \4815_b0 );
or ( \4817_b1 , \4814_b1 , w_15402 );
or ( \4817_b0 , \4814_b0 , \4816_b0 );
not ( \4816_b0 , w_15403 );
and ( w_15403 , w_15402 , \4816_b1 );
or ( \4818_b1 , \4047_b1 , \4156_b1 );
xor ( \4818_b0 , \4047_b0 , w_15404 );
not ( w_15404 , w_15405 );
and ( w_15405 , \4156_b1 , \4156_b0 );
or ( \4819_b1 , \4818_b1 , w_15407 );
not ( w_15407 , w_15408 );
and ( \4819_b0 , \4818_b0 , w_15409 );
and ( w_15408 ,  , w_15409 );
buf ( w_15407 , \4742_b1 );
not ( w_15407 , w_15410 );
not (  , w_15411 );
and ( w_15410 , w_15411 , \4742_b0 );
or ( \4820_b1 , \4817_b1 , w_15413 );
not ( w_15413 , w_15414 );
and ( \4820_b0 , \4817_b0 , w_15415 );
and ( w_15414 ,  , w_15415 );
buf ( w_15413 , \4819_b1 );
not ( w_15413 , w_15416 );
not (  , w_15417 );
and ( w_15416 , w_15417 , \4819_b0 );
or ( \4821_b1 , \4813_b1 , \4820_b1 );
xor ( \4821_b0 , \4813_b0 , w_15418 );
not ( w_15418 , w_15419 );
and ( w_15419 , \4820_b1 , \4820_b0 );
or ( \4822_b1 , \4794_b1 , \4821_b1 );
xor ( \4822_b0 , \4794_b0 , w_15420 );
not ( w_15420 , w_15421 );
and ( w_15421 , \4821_b1 , \4821_b0 );
or ( \4823_b1 , \4776_b1 , \4822_b1 );
xor ( \4823_b0 , \4776_b0 , w_15422 );
not ( w_15422 , w_15423 );
and ( w_15423 , \4822_b1 , \4822_b0 );
buf ( \4824_b1 , \4757_b1 );
not ( \4824_b1 , w_15424 );
not ( \4824_b0 , w_15425 );
and ( w_15424 , w_15425 , \4757_b0 );
or ( \4825_b1 , \4824_b1 , w_15427 );
not ( w_15427 , w_15428 );
and ( \4825_b0 , \4824_b0 , w_15429 );
and ( w_15428 ,  , w_15429 );
buf ( w_15427 , \4736_b1 );
not ( w_15427 , w_15430 );
not (  , w_15431 );
and ( w_15430 , w_15431 , \4736_b0 );
buf ( \4826_b1 , \4825_b1 );
not ( \4826_b1 , w_15432 );
not ( \4826_b0 , w_15433 );
and ( w_15432 , w_15433 , \4825_b0 );
buf ( \4827_b1 , \4762_b1 );
not ( \4827_b1 , w_15434 );
not ( \4827_b0 , w_15435 );
and ( w_15434 , w_15435 , \4762_b0 );
or ( \4828_b1 , \4826_b1 , w_15436 );
or ( \4828_b0 , \4826_b0 , \4827_b0 );
not ( \4827_b0 , w_15437 );
and ( w_15437 , w_15436 , \4827_b1 );
buf ( \4829_b1 , \4736_b1 );
not ( \4829_b1 , w_15438 );
not ( \4829_b0 , w_15439 );
and ( w_15438 , w_15439 , \4736_b0 );
or ( \4830_b1 , \4829_b1 , w_15441 );
not ( w_15441 , w_15442 );
and ( \4830_b0 , \4829_b0 , w_15443 );
and ( w_15442 ,  , w_15443 );
buf ( w_15441 , \4757_b1 );
not ( w_15441 , w_15444 );
not (  , w_15445 );
and ( w_15444 , w_15445 , \4757_b0 );
or ( \4831_b1 , \4828_b1 , w_15447 );
not ( w_15447 , w_15448 );
and ( \4831_b0 , \4828_b0 , w_15449 );
and ( w_15448 ,  , w_15449 );
buf ( w_15447 , \4830_b1 );
not ( w_15447 , w_15450 );
not (  , w_15451 );
and ( w_15450 , w_15451 , \4830_b0 );
or ( \4832_b1 , \4823_b1 , \4831_b1 );
xor ( \4832_b0 , \4823_b0 , w_15452 );
not ( w_15452 , w_15453 );
and ( w_15453 , \4831_b1 , \4831_b0 );
buf ( \4833_b1 , \4832_b1 );
not ( \4833_b1 , w_15454 );
not ( \4833_b0 , w_15455 );
and ( w_15454 , w_15455 , \4832_b0 );
or ( \4834_b1 , \4772_b1 , w_15457 );
not ( w_15457 , w_15458 );
and ( \4834_b0 , \4772_b0 , w_15459 );
and ( w_15458 ,  , w_15459 );
buf ( w_15457 , \4833_b1 );
not ( w_15457 , w_15460 );
not (  , w_15461 );
and ( w_15460 , w_15461 , \4833_b0 );
buf ( \4835_b1 , \4834_b1 );
not ( \4835_b1 , w_15462 );
not ( \4835_b0 , w_15463 );
and ( w_15462 , w_15463 , \4834_b0 );
or ( \4836_b1 , \4767_b1 , w_15465 );
not ( w_15465 , w_15466 );
and ( \4836_b0 , \4767_b0 , w_15467 );
and ( w_15466 ,  , w_15467 );
buf ( w_15465 , \4835_b1 );
not ( w_15465 , w_15468 );
not (  , w_15469 );
and ( w_15468 , w_15469 , \4835_b0 );
or ( \4837_b1 , \4776_b1 , \4822_b1 );
xor ( \4837_b0 , \4776_b0 , w_15470 );
not ( w_15470 , w_15471 );
and ( w_15471 , \4822_b1 , \4822_b0 );
or ( \4838_b1 , \4837_b1 , \4831_b1 );
not ( \4831_b1 , w_15472 );
and ( \4838_b0 , \4837_b0 , w_15473 );
and ( w_15472 , w_15473 , \4831_b0 );
or ( \4839_b1 , \4776_b1 , \4822_b1 );
not ( \4822_b1 , w_15474 );
and ( \4839_b0 , \4776_b0 , w_15475 );
and ( w_15474 , w_15475 , \4822_b0 );
or ( \4840_b1 , \4838_b1 , w_15476 );
or ( \4840_b0 , \4838_b0 , \4839_b0 );
not ( \4839_b0 , w_15477 );
and ( w_15477 , w_15476 , \4839_b1 );
buf ( \4841_b1 , \4840_b1 );
not ( \4841_b1 , w_15478 );
not ( \4841_b0 , w_15479 );
and ( w_15478 , w_15479 , \4840_b0 );
or ( \4842_b1 , \4045_b1 , \4156_b1 );
not ( \4156_b1 , w_15480 );
and ( \4842_b0 , \4045_b0 , w_15481 );
and ( w_15480 , w_15481 , \4156_b0 );
buf ( \4843_b1 , \4786_b1 );
not ( \4843_b1 , w_15482 );
not ( \4843_b0 , w_15483 );
and ( w_15482 , w_15483 , \4786_b0 );
buf ( \4844_b1 , \4496_b1 );
not ( \4844_b1 , w_15484 );
not ( \4844_b0 , w_15485 );
and ( w_15484 , w_15485 , \4496_b0 );
or ( \4845_b1 , \4843_b1 , w_15486 );
or ( \4845_b0 , \4843_b0 , \4844_b0 );
not ( \4844_b0 , w_15487 );
and ( w_15487 , w_15486 , \4844_b1 );
buf ( \4846_b1 , \4044_b1 );
not ( \4846_b1 , w_15488 );
not ( \4846_b0 , w_15489 );
and ( w_15488 , w_15489 , \4044_b0 );
buf ( \4847_b1 , \4213_b1 );
not ( \4847_b1 , w_15490 );
not ( \4847_b0 , w_15491 );
and ( w_15490 , w_15491 , \4213_b0 );
or ( \4848_b1 , \4846_b1 , w_15492 );
or ( \4848_b0 , \4846_b0 , \4847_b0 );
not ( \4847_b0 , w_15493 );
and ( w_15493 , w_15492 , \4847_b1 );
buf ( \4849_b1 , \4213_b1 );
not ( \4849_b1 , w_15494 );
not ( \4849_b0 , w_15495 );
and ( w_15494 , w_15495 , \4213_b0 );
or ( \4850_b1 , \4849_b1 , w_15497 );
not ( w_15497 , w_15498 );
and ( \4850_b0 , \4849_b0 , w_15499 );
and ( w_15498 ,  , w_15499 );
buf ( w_15497 , \4092_b1 );
not ( w_15497 , w_15500 );
not (  , w_15501 );
and ( w_15500 , w_15501 , \4092_b0 );
or ( \4851_b1 , \4848_b1 , w_15503 );
not ( w_15503 , w_15504 );
and ( \4851_b0 , \4848_b0 , w_15505 );
and ( w_15504 ,  , w_15505 );
buf ( w_15503 , \4850_b1 );
not ( w_15503 , w_15506 );
not (  , w_15507 );
and ( w_15506 , w_15507 , \4850_b0 );
or ( \4852_b1 , \4377_b1 , w_15509 );
not ( w_15509 , w_15510 );
and ( \4852_b0 , \4377_b0 , w_15511 );
and ( w_15510 ,  , w_15511 );
buf ( w_15509 , \4851_b1 );
not ( w_15509 , w_15512 );
not (  , w_15513 );
and ( w_15512 , w_15513 , \4851_b0 );
or ( \4853_b1 , \4845_b1 , w_15515 );
not ( w_15515 , w_15516 );
and ( \4853_b0 , \4845_b0 , w_15517 );
and ( w_15516 ,  , w_15517 );
buf ( w_15515 , \4852_b1 );
not ( w_15515 , w_15518 );
not (  , w_15519 );
and ( w_15518 , w_15519 , \4852_b0 );
or ( \4854_b1 , \4842_b1 , \4853_b1 );
xor ( \4854_b0 , \4842_b0 , w_15520 );
not ( w_15520 , w_15521 );
and ( w_15521 , \4853_b1 , \4853_b0 );
buf ( \4855_b1 , \4818_b1 );
not ( \4855_b1 , w_15522 );
not ( \4855_b0 , w_15523 );
and ( w_15522 , w_15523 , \4818_b0 );
buf ( \4856_b1 , \4815_b1 );
not ( \4856_b1 , w_15524 );
not ( \4856_b0 , w_15525 );
and ( w_15524 , w_15525 , \4815_b0 );
or ( \4857_b1 , \4855_b1 , w_15526 );
or ( \4857_b0 , \4855_b0 , \4856_b0 );
not ( \4856_b0 , w_15527 );
and ( w_15527 , w_15526 , \4856_b1 );
or ( \4858_b1 , \4042_b1 , \4156_b1 );
xor ( \4858_b0 , \4042_b0 , w_15528 );
not ( w_15528 , w_15529 );
and ( w_15529 , \4156_b1 , \4156_b0 );
buf ( \4859_b1 , \4742_b1 );
buf ( \4859_b0 , \4742_b0 );
or ( \4860_b1 , \4858_b1 , w_15531 );
not ( w_15531 , w_15532 );
and ( \4860_b0 , \4858_b0 , w_15533 );
and ( w_15532 ,  , w_15533 );
buf ( w_15531 , \4859_b1 );
not ( w_15531 , w_15534 );
not (  , w_15535 );
and ( w_15534 , w_15535 , \4859_b0 );
or ( \4861_b1 , \4857_b1 , w_15537 );
not ( w_15537 , w_15538 );
and ( \4861_b0 , \4857_b0 , w_15539 );
and ( w_15538 ,  , w_15539 );
buf ( w_15537 , \4860_b1 );
not ( w_15537 , w_15540 );
not (  , w_15541 );
and ( w_15540 , w_15541 , \4860_b0 );
or ( \4862_b1 , \4854_b1 , \4861_b1 );
xor ( \4862_b0 , \4854_b0 , w_15542 );
not ( w_15542 , w_15543 );
and ( w_15543 , \4861_b1 , \4861_b0 );
or ( \4863_b1 , \4195_b1 , \4802_b1 );
not ( \4802_b1 , w_15544 );
and ( \4863_b0 , \4195_b0 , w_15545 );
and ( w_15544 , w_15545 , \4802_b0 );
or ( \4864_b1 , \4205_b1 , \4172_b1 );
not ( \4172_b1 , w_15546 );
and ( \4864_b0 , \4205_b0 , w_15547 );
and ( w_15546 , w_15547 , \4172_b0 );
or ( \4865_b1 , \4863_b1 , w_15549 );
not ( w_15549 , w_15550 );
and ( \4865_b0 , \4863_b0 , w_15551 );
and ( w_15550 ,  , w_15551 );
buf ( w_15549 , \4864_b1 );
not ( w_15549 , w_15552 );
not (  , w_15553 );
and ( w_15552 , w_15553 , \4864_b0 );
or ( \4866_b1 , \4777_b1 , \4715_b1 );
xor ( \4866_b0 , \4777_b0 , w_15554 );
not ( w_15554 , w_15555 );
and ( w_15555 , \4715_b1 , \4715_b0 );
or ( \4867_b1 , \4866_b1 , \4788_b1 );
not ( \4788_b1 , w_15556 );
and ( \4867_b0 , \4866_b0 , w_15557 );
and ( w_15556 , w_15557 , \4788_b0 );
or ( \4868_b1 , \4777_b1 , \4715_b1 );
not ( \4715_b1 , w_15558 );
and ( \4868_b0 , \4777_b0 , w_15559 );
and ( w_15558 , w_15559 , \4715_b0 );
or ( \4869_b1 , \4867_b1 , w_15560 );
or ( \4869_b0 , \4867_b0 , \4868_b0 );
not ( \4868_b0 , w_15561 );
and ( w_15561 , w_15560 , \4868_b1 );
or ( \4870_b1 , \4865_b1 , \4869_b1 );
xor ( \4870_b0 , \4865_b0 , w_15562 );
not ( w_15562 , w_15563 );
and ( w_15563 , \4869_b1 , \4869_b0 );
buf ( \4871_b1 , \4809_b1 );
not ( \4871_b1 , w_15564 );
not ( \4871_b0 , w_15565 );
and ( w_15564 , w_15565 , \4809_b0 );
buf ( \4872_b1 , \4820_b1 );
not ( \4872_b1 , w_15566 );
not ( \4872_b0 , w_15567 );
and ( w_15566 , w_15567 , \4820_b0 );
or ( \4873_b1 , \4871_b1 , w_15568 );
or ( \4873_b0 , \4871_b0 , \4872_b0 );
not ( \4872_b0 , w_15569 );
and ( w_15569 , w_15568 , \4872_b1 );
or ( \4874_b1 , \4820_b1 , w_15570 );
or ( \4874_b0 , \4820_b0 , \4809_b0 );
not ( \4809_b0 , w_15571 );
and ( w_15571 , w_15570 , \4809_b1 );
or ( \4875_b1 , \4874_b1 , w_15573 );
not ( w_15573 , w_15574 );
and ( \4875_b0 , \4874_b0 , w_15575 );
and ( w_15574 ,  , w_15575 );
buf ( w_15573 , \4804_b1 );
not ( w_15573 , w_15576 );
not (  , w_15577 );
and ( w_15576 , w_15577 , \4804_b0 );
or ( \4876_b1 , \4873_b1 , w_15579 );
not ( w_15579 , w_15580 );
and ( \4876_b0 , \4873_b0 , w_15581 );
and ( w_15580 ,  , w_15581 );
buf ( w_15579 , \4875_b1 );
not ( w_15579 , w_15582 );
not (  , w_15583 );
and ( w_15582 , w_15583 , \4875_b0 );
or ( \4877_b1 , \4870_b1 , \4876_b1 );
xor ( \4877_b0 , \4870_b0 , w_15584 );
not ( w_15584 , w_15585 );
and ( w_15585 , \4876_b1 , \4876_b0 );
or ( \4878_b1 , \4862_b1 , \4877_b1 );
xor ( \4878_b0 , \4862_b0 , w_15586 );
not ( w_15586 , w_15587 );
and ( w_15587 , \4877_b1 , \4877_b0 );
or ( \4879_b1 , \4789_b1 , \4793_b1 );
xor ( \4879_b0 , \4789_b0 , w_15588 );
not ( w_15588 , w_15589 );
and ( w_15589 , \4793_b1 , \4793_b0 );
or ( \4880_b1 , \4879_b1 , \4821_b1 );
not ( \4821_b1 , w_15590 );
and ( \4880_b0 , \4879_b0 , w_15591 );
and ( w_15590 , w_15591 , \4821_b0 );
or ( \4881_b1 , \4789_b1 , \4793_b1 );
not ( \4793_b1 , w_15592 );
and ( \4881_b0 , \4789_b0 , w_15593 );
and ( w_15592 , w_15593 , \4793_b0 );
or ( \4882_b1 , \4880_b1 , w_15594 );
or ( \4882_b0 , \4880_b0 , \4881_b0 );
not ( \4881_b0 , w_15595 );
and ( w_15595 , w_15594 , \4881_b1 );
or ( \4883_b1 , \4878_b1 , \4882_b1 );
xor ( \4883_b0 , \4878_b0 , w_15596 );
not ( w_15596 , w_15597 );
and ( w_15597 , \4882_b1 , \4882_b0 );
buf ( \4884_b1 , \4883_b1 );
not ( \4884_b1 , w_15598 );
not ( \4884_b0 , w_15599 );
and ( w_15598 , w_15599 , \4883_b0 );
or ( \4885_b1 , \4841_b1 , w_15601 );
not ( w_15601 , w_15602 );
and ( \4885_b0 , \4841_b0 , w_15603 );
and ( w_15602 ,  , w_15603 );
buf ( w_15601 , \4884_b1 );
not ( w_15601 , w_15604 );
not (  , w_15605 );
and ( w_15604 , w_15605 , \4884_b0 );
or ( \4886_b1 , \4047_b1 , \4156_b1 );
not ( \4156_b1 , w_15606 );
and ( \4886_b0 , \4047_b0 , w_15607 );
and ( w_15606 , w_15607 , \4156_b0 );
buf ( \4887_b1 , \4851_b1 );
not ( \4887_b1 , w_15608 );
not ( \4887_b0 , w_15609 );
and ( w_15608 , w_15609 , \4851_b0 );
buf ( \4888_b1 , \4496_b1 );
not ( \4888_b1 , w_15610 );
not ( \4888_b0 , w_15611 );
and ( w_15610 , w_15611 , \4496_b0 );
or ( \4889_b1 , \4887_b1 , w_15612 );
or ( \4889_b0 , \4887_b0 , \4888_b0 );
not ( \4888_b0 , w_15613 );
and ( w_15613 , w_15612 , \4888_b1 );
or ( \4890_b1 , \4213_b1 , \3994_b1 );
not ( \3994_b1 , w_15614 );
and ( \4890_b0 , \4213_b0 , w_15615 );
and ( w_15614 , w_15615 , \3994_b0 );
or ( \4891_b1 , \4849_b1 , \4099_b1 );
not ( \4099_b1 , w_15616 );
and ( \4891_b0 , \4849_b0 , w_15617 );
and ( w_15616 , w_15617 , \4099_b0 );
or ( \4892_b1 , \4890_b1 , w_15619 );
not ( w_15619 , w_15620 );
and ( \4892_b0 , \4890_b0 , w_15621 );
and ( w_15620 ,  , w_15621 );
buf ( w_15619 , \4891_b1 );
not ( w_15619 , w_15622 );
not (  , w_15623 );
and ( w_15622 , w_15623 , \4891_b0 );
buf ( \4893_b1 , \4892_b1 );
not ( \4893_b1 , w_15624 );
not ( \4893_b0 , w_15625 );
and ( w_15624 , w_15625 , \4892_b0 );
or ( \4894_b1 , \4893_b1 , w_15627 );
not ( w_15627 , w_15628 );
and ( \4894_b0 , \4893_b0 , w_15629 );
and ( w_15628 ,  , w_15629 );
buf ( w_15627 , \4377_b1 );
not ( w_15627 , w_15630 );
not (  , w_15631 );
and ( w_15630 , w_15631 , \4377_b0 );
or ( \4895_b1 , \4889_b1 , w_15633 );
not ( w_15633 , w_15634 );
and ( \4895_b0 , \4889_b0 , w_15635 );
and ( w_15634 ,  , w_15635 );
buf ( w_15633 , \4894_b1 );
not ( w_15633 , w_15636 );
not (  , w_15637 );
and ( w_15636 , w_15637 , \4894_b0 );
or ( \4896_b1 , \4886_b1 , \4895_b1 );
xor ( \4896_b0 , \4886_b0 , w_15638 );
not ( w_15638 , w_15639 );
and ( w_15639 , \4895_b1 , \4895_b0 );
buf ( \4897_b1 , \4319_b1 );
not ( \4897_b1 , w_15640 );
not ( \4897_b0 , w_15641 );
and ( w_15640 , w_15641 , \4319_b0 );
buf ( \4898_b1 , \4317_b1 );
not ( \4898_b1 , w_15642 );
not ( \4898_b0 , w_15643 );
and ( w_15642 , w_15643 , \4317_b0 );
or ( \4899_b1 , \4897_b1 , w_15644 );
or ( \4899_b0 , \4897_b0 , \4898_b0 );
not ( \4898_b0 , w_15645 );
and ( w_15645 , w_15644 , \4898_b1 );
or ( \4900_b1 , \4899_b1 , w_15647 );
not ( w_15647 , w_15648 );
and ( \4900_b0 , \4899_b0 , w_15649 );
and ( w_15648 ,  , w_15649 );
buf ( w_15647 , \4172_b1 );
not ( w_15647 , w_15650 );
not (  , w_15651 );
and ( w_15650 , w_15651 , \4172_b0 );
or ( \4901_b1 , \4896_b1 , \4900_b1 );
xor ( \4901_b0 , \4896_b0 , w_15652 );
not ( w_15652 , w_15653 );
and ( w_15653 , \4900_b1 , \4900_b0 );
buf ( \4902_b1 , \4865_b1 );
not ( \4902_b1 , w_15654 );
not ( \4902_b0 , w_15655 );
and ( w_15654 , w_15655 , \4865_b0 );
buf ( \4903_b1 , \4858_b1 );
not ( \4903_b1 , w_15656 );
not ( \4903_b0 , w_15657 );
and ( w_15656 , w_15657 , \4858_b0 );
buf ( \4904_b1 , \4815_b1 );
not ( \4904_b1 , w_15658 );
not ( \4904_b0 , w_15659 );
and ( w_15658 , w_15659 , \4815_b0 );
or ( \4905_b1 , \4903_b1 , w_15660 );
or ( \4905_b0 , \4903_b0 , \4904_b0 );
not ( \4904_b0 , w_15661 );
and ( w_15661 , w_15660 , \4904_b1 );
or ( \4906_b1 , \3943_b1 , \4156_b1 );
xor ( \4906_b0 , \3943_b0 , w_15662 );
not ( w_15662 , w_15663 );
and ( w_15663 , \4156_b1 , \4156_b0 );
or ( \4907_b1 , \4906_b1 , w_15665 );
not ( w_15665 , w_15666 );
and ( \4907_b0 , \4906_b0 , w_15667 );
and ( w_15666 ,  , w_15667 );
buf ( w_15665 , \4859_b1 );
not ( w_15665 , w_15668 );
not (  , w_15669 );
and ( w_15668 , w_15669 , \4859_b0 );
or ( \4908_b1 , \4905_b1 , w_15671 );
not ( w_15671 , w_15672 );
and ( \4908_b0 , \4905_b0 , w_15673 );
and ( w_15672 ,  , w_15673 );
buf ( w_15671 , \4907_b1 );
not ( w_15671 , w_15674 );
not (  , w_15675 );
and ( w_15674 , w_15675 , \4907_b0 );
or ( \4909_b1 , \4902_b1 , \4908_b1 );
xor ( \4909_b0 , \4902_b0 , w_15676 );
not ( w_15676 , w_15677 );
and ( w_15677 , \4908_b1 , \4908_b0 );
or ( \4910_b1 , \4842_b1 , \4853_b1 );
xor ( \4910_b0 , \4842_b0 , w_15678 );
not ( w_15678 , w_15679 );
and ( w_15679 , \4853_b1 , \4853_b0 );
or ( \4911_b1 , \4910_b1 , \4861_b1 );
not ( \4861_b1 , w_15680 );
and ( \4911_b0 , \4910_b0 , w_15681 );
and ( w_15680 , w_15681 , \4861_b0 );
or ( \4912_b1 , \4842_b1 , \4853_b1 );
not ( \4853_b1 , w_15682 );
and ( \4912_b0 , \4842_b0 , w_15683 );
and ( w_15682 , w_15683 , \4853_b0 );
or ( \4913_b1 , \4911_b1 , w_15684 );
or ( \4913_b0 , \4911_b0 , \4912_b0 );
not ( \4912_b0 , w_15685 );
and ( w_15685 , w_15684 , \4912_b1 );
or ( \4914_b1 , \4909_b1 , \4913_b1 );
xor ( \4914_b0 , \4909_b0 , w_15686 );
not ( w_15686 , w_15687 );
and ( w_15687 , \4913_b1 , \4913_b0 );
or ( \4915_b1 , \4901_b1 , \4914_b1 );
xor ( \4915_b0 , \4901_b0 , w_15688 );
not ( w_15688 , w_15689 );
and ( w_15689 , \4914_b1 , \4914_b0 );
or ( \4916_b1 , \4865_b1 , \4869_b1 );
xor ( \4916_b0 , \4865_b0 , w_15690 );
not ( w_15690 , w_15691 );
and ( w_15691 , \4869_b1 , \4869_b0 );
or ( \4917_b1 , \4916_b1 , \4876_b1 );
not ( \4876_b1 , w_15692 );
and ( \4917_b0 , \4916_b0 , w_15693 );
and ( w_15692 , w_15693 , \4876_b0 );
or ( \4918_b1 , \4865_b1 , \4869_b1 );
not ( \4869_b1 , w_15694 );
and ( \4918_b0 , \4865_b0 , w_15695 );
and ( w_15694 , w_15695 , \4869_b0 );
or ( \4919_b1 , \4917_b1 , w_15696 );
or ( \4919_b0 , \4917_b0 , \4918_b0 );
not ( \4918_b0 , w_15697 );
and ( w_15697 , w_15696 , \4918_b1 );
or ( \4920_b1 , \4915_b1 , w_15698 );
xor ( \4920_b0 , \4915_b0 , w_15700 );
not ( w_15700 , w_15701 );
and ( w_15701 , w_15698 , w_15699 );
buf ( w_15698 , \4919_b1 );
not ( w_15698 , w_15702 );
not ( w_15699 , w_15703 );
and ( w_15702 , w_15703 , \4919_b0 );
buf ( \4921_b1 , \4877_b1 );
not ( \4921_b1 , w_15704 );
not ( \4921_b0 , w_15705 );
and ( w_15704 , w_15705 , \4877_b0 );
buf ( \4922_b1 , \4862_b1 );
not ( \4922_b1 , w_15706 );
not ( \4922_b0 , w_15707 );
and ( w_15706 , w_15707 , \4862_b0 );
or ( \4923_b1 , \4921_b1 , w_15709 );
not ( w_15709 , w_15710 );
and ( \4923_b0 , \4921_b0 , w_15711 );
and ( w_15710 ,  , w_15711 );
buf ( w_15709 , \4922_b1 );
not ( w_15709 , w_15712 );
not (  , w_15713 );
and ( w_15712 , w_15713 , \4922_b0 );
or ( \4924_b1 , \4923_b1 , \4882_b1 );
not ( \4882_b1 , w_15714 );
and ( \4924_b0 , \4923_b0 , w_15715 );
and ( w_15714 , w_15715 , \4882_b0 );
or ( \4925_b1 , \4921_b1 , w_15717 );
not ( w_15717 , w_15718 );
and ( \4925_b0 , \4921_b0 , w_15719 );
and ( w_15718 ,  , w_15719 );
buf ( w_15717 , \4922_b1 );
not ( w_15717 , w_15720 );
not (  , w_15721 );
and ( w_15720 , w_15721 , \4922_b0 );
or ( \4926_b1 , \4924_b1 , w_15723 );
not ( w_15723 , w_15724 );
and ( \4926_b0 , \4924_b0 , w_15725 );
and ( w_15724 ,  , w_15725 );
buf ( w_15723 , \4925_b1 );
not ( w_15723 , w_15726 );
not (  , w_15727 );
and ( w_15726 , w_15727 , \4925_b0 );
or ( \4927_b1 , \4920_b1 , w_15729 );
not ( w_15729 , w_15730 );
and ( \4927_b0 , \4920_b0 , w_15731 );
and ( w_15730 ,  , w_15731 );
buf ( w_15729 , \4926_b1 );
not ( w_15729 , w_15732 );
not (  , w_15733 );
and ( w_15732 , w_15733 , \4926_b0 );
or ( \4929_b1 , \4901_b1 , w_15734 );
or ( \4929_b0 , \4901_b0 , \4914_b0 );
not ( \4914_b0 , w_15735 );
and ( w_15735 , w_15734 , \4914_b1 );
or ( \4930_b1 , \4929_b1 , w_15737 );
not ( w_15737 , w_15738 );
and ( \4930_b0 , \4929_b0 , w_15739 );
and ( w_15738 ,  , w_15739 );
buf ( w_15737 , \4919_b1 );
not ( w_15737 , w_15740 );
not (  , w_15741 );
and ( w_15740 , w_15741 , \4919_b0 );
or ( \4931_b1 , \4914_b1 , w_15743 );
not ( w_15743 , w_15744 );
and ( \4931_b0 , \4914_b0 , w_15745 );
and ( w_15744 ,  , w_15745 );
buf ( w_15743 , \4901_b1 );
not ( w_15743 , w_15746 );
not (  , w_15747 );
and ( w_15746 , w_15747 , \4901_b0 );
or ( \4932_b1 , \4930_b1 , w_15749 );
not ( w_15749 , w_15750 );
and ( \4932_b0 , \4930_b0 , w_15751 );
and ( w_15750 ,  , w_15751 );
buf ( w_15749 , \4931_b1 );
not ( w_15749 , w_15752 );
not (  , w_15753 );
and ( w_15752 , w_15753 , \4931_b0 );
or ( \4933_b1 , \4886_b1 , \4895_b1 );
xor ( \4933_b0 , \4886_b0 , w_15754 );
not ( w_15754 , w_15755 );
and ( w_15755 , \4895_b1 , \4895_b0 );
or ( \4934_b1 , \4933_b1 , \4900_b1 );
not ( \4900_b1 , w_15756 );
and ( \4934_b0 , \4933_b0 , w_15757 );
and ( w_15756 , w_15757 , \4900_b0 );
or ( \4935_b1 , \4886_b1 , \4895_b1 );
not ( \4895_b1 , w_15758 );
and ( \4935_b0 , \4886_b0 , w_15759 );
and ( w_15758 , w_15759 , \4895_b0 );
or ( \4936_b1 , \4934_b1 , w_15760 );
or ( \4936_b0 , \4934_b0 , \4935_b0 );
not ( \4935_b0 , w_15761 );
and ( w_15761 , w_15760 , \4935_b1 );
or ( \4937_b1 , \4042_b1 , \4156_b1 );
not ( \4156_b1 , w_15762 );
and ( \4937_b0 , \4042_b0 , w_15763 );
and ( w_15762 , w_15763 , \4156_b0 );
buf ( \4938_b1 , \4892_b1 );
not ( \4938_b1 , w_15764 );
not ( \4938_b0 , w_15765 );
and ( w_15764 , w_15765 , \4892_b0 );
buf ( \4939_b1 , \4496_b1 );
not ( \4939_b1 , w_15766 );
not ( \4939_b0 , w_15767 );
and ( w_15766 , w_15767 , \4496_b0 );
buf ( \4940_b1 , \4939_b1 );
not ( \4940_b1 , w_15768 );
not ( \4940_b0 , w_15769 );
and ( w_15768 , w_15769 , \4939_b0 );
or ( \4941_b1 , \4938_b1 , \4940_b1 );
not ( \4940_b1 , w_15770 );
and ( \4941_b0 , \4938_b0 , w_15771 );
and ( w_15770 , w_15771 , \4940_b0 );
or ( \4942_b1 , \4377_b1 , \4849_b1 );
not ( \4849_b1 , w_15772 );
and ( \4942_b0 , \4377_b0 , w_15773 );
and ( w_15772 , w_15773 , \4849_b0 );
or ( \4943_b1 , \4941_b1 , w_15775 );
not ( w_15775 , w_15776 );
and ( \4943_b0 , \4941_b0 , w_15777 );
and ( w_15776 ,  , w_15777 );
buf ( w_15775 , \4942_b1 );
not ( w_15775 , w_15778 );
not (  , w_15779 );
and ( w_15778 , w_15779 , \4942_b0 );
or ( \4944_b1 , \4937_b1 , \4943_b1 );
xor ( \4944_b0 , \4937_b0 , w_15780 );
not ( w_15780 , w_15781 );
and ( w_15781 , \4943_b1 , \4943_b0 );
buf ( \4945_b1 , \4906_b1 );
not ( \4945_b1 , w_15782 );
not ( \4945_b0 , w_15783 );
and ( w_15782 , w_15783 , \4906_b0 );
or ( \4946_b1 , \4254_b1 , w_15784 );
or ( \4946_b0 , \4254_b0 , \4945_b0 );
not ( \4945_b0 , w_15785 );
and ( w_15785 , w_15784 , \4945_b1 );
or ( \4947_b1 , \4267_b1 , \4044_b1 );
not ( \4044_b1 , w_15786 );
and ( \4947_b0 , \4267_b0 , w_15787 );
and ( w_15786 , w_15787 , \4044_b0 );
or ( \4948_b1 , \4156_b1 , \4092_b1 );
not ( \4092_b1 , w_15788 );
and ( \4948_b0 , \4156_b0 , w_15789 );
and ( w_15788 , w_15789 , \4092_b0 );
or ( \4949_b1 , \4947_b1 , w_15791 );
not ( w_15791 , w_15792 );
and ( \4949_b0 , \4947_b0 , w_15793 );
and ( w_15792 ,  , w_15793 );
buf ( w_15791 , \4948_b1 );
not ( w_15791 , w_15794 );
not (  , w_15795 );
and ( w_15794 , w_15795 , \4948_b0 );
buf ( \4950_b1 , \4859_b1 );
not ( \4950_b1 , w_15796 );
not ( \4950_b0 , w_15797 );
and ( w_15796 , w_15797 , \4859_b0 );
or ( \4951_b1 , \4949_b1 , w_15798 );
or ( \4951_b0 , \4949_b0 , \4950_b0 );
not ( \4950_b0 , w_15799 );
and ( w_15799 , w_15798 , \4950_b1 );
or ( \4952_b1 , \4946_b1 , w_15801 );
not ( w_15801 , w_15802 );
and ( \4952_b0 , \4946_b0 , w_15803 );
and ( w_15802 ,  , w_15803 );
buf ( w_15801 , \4951_b1 );
not ( w_15801 , w_15804 );
not (  , w_15805 );
and ( w_15804 , w_15805 , \4951_b0 );
or ( \4953_b1 , \4944_b1 , \4952_b1 );
xor ( \4953_b0 , \4944_b0 , w_15806 );
not ( w_15806 , w_15807 );
and ( w_15807 , \4952_b1 , \4952_b0 );
or ( \4954_b1 , \4936_b1 , \4953_b1 );
xor ( \4954_b0 , \4936_b0 , w_15808 );
not ( w_15808 , w_15809 );
and ( w_15809 , \4953_b1 , \4953_b0 );
or ( \4955_b1 , \4902_b1 , \4908_b1 );
xor ( \4955_b0 , \4902_b0 , w_15810 );
not ( w_15810 , w_15811 );
and ( w_15811 , \4908_b1 , \4908_b0 );
or ( \4956_b1 , \4955_b1 , \4913_b1 );
not ( \4913_b1 , w_15812 );
and ( \4956_b0 , \4955_b0 , w_15813 );
and ( w_15812 , w_15813 , \4913_b0 );
or ( \4957_b1 , \4902_b1 , \4908_b1 );
not ( \4908_b1 , w_15814 );
and ( \4957_b0 , \4902_b0 , w_15815 );
and ( w_15814 , w_15815 , \4908_b0 );
or ( \4958_b1 , \4956_b1 , w_15816 );
or ( \4958_b0 , \4956_b0 , \4957_b0 );
not ( \4957_b0 , w_15817 );
and ( w_15817 , w_15816 , \4957_b1 );
or ( \4959_b1 , \4954_b1 , \4958_b1 );
xor ( \4959_b0 , \4954_b0 , w_15818 );
not ( w_15818 , w_15819 );
and ( w_15819 , \4958_b1 , \4958_b0 );
or ( \4960_b1 , \4932_b1 , w_15821 );
not ( w_15821 , w_15822 );
and ( \4960_b0 , \4932_b0 , w_15823 );
and ( w_15822 ,  , w_15823 );
buf ( w_15821 , \4959_b1 );
not ( w_15821 , w_15824 );
not (  , w_15825 );
and ( w_15824 , w_15825 , \4959_b0 );
or ( \4961_b1 , \4936_b1 , \4953_b1 );
xor ( \4961_b0 , \4936_b0 , w_15826 );
not ( w_15826 , w_15827 );
and ( w_15827 , \4953_b1 , \4953_b0 );
or ( \4962_b1 , \4961_b1 , \4958_b1 );
not ( \4958_b1 , w_15828 );
and ( \4962_b0 , \4961_b0 , w_15829 );
and ( w_15828 , w_15829 , \4958_b0 );
or ( \4963_b1 , \4936_b1 , \4953_b1 );
not ( \4953_b1 , w_15830 );
and ( \4963_b0 , \4936_b0 , w_15831 );
and ( w_15830 , w_15831 , \4953_b0 );
or ( \4964_b1 , \4962_b1 , w_15832 );
or ( \4964_b0 , \4962_b0 , \4963_b0 );
not ( \4963_b0 , w_15833 );
and ( w_15833 , w_15832 , \4963_b1 );
or ( \4965_b1 , \4937_b1 , \4943_b1 );
xor ( \4965_b0 , \4937_b0 , w_15834 );
not ( w_15834 , w_15835 );
and ( w_15835 , \4943_b1 , \4943_b0 );
or ( \4966_b1 , \4965_b1 , \4952_b1 );
not ( \4952_b1 , w_15836 );
and ( \4966_b0 , \4965_b0 , w_15837 );
and ( w_15836 , w_15837 , \4952_b0 );
or ( \4967_b1 , \4937_b1 , \4943_b1 );
not ( \4943_b1 , w_15838 );
and ( \4967_b0 , \4937_b0 , w_15839 );
and ( w_15838 , w_15839 , \4943_b0 );
or ( \4968_b1 , \4966_b1 , w_15840 );
or ( \4968_b0 , \4966_b0 , \4967_b0 );
not ( \4967_b0 , w_15841 );
and ( w_15841 , w_15840 , \4967_b1 );
buf ( \4969_b1 , \4943_b1 );
not ( \4969_b1 , w_15842 );
not ( \4969_b0 , w_15843 );
and ( w_15842 , w_15843 , \4943_b0 );
or ( \4970_b1 , \4968_b1 , \4969_b1 );
xor ( \4970_b0 , \4968_b0 , w_15844 );
not ( w_15844 , w_15845 );
and ( w_15845 , \4969_b1 , \4969_b0 );
or ( \4971_b1 , \4496_b1 , w_15846 );
or ( \4971_b0 , \4496_b0 , \4377_b0 );
not ( \4377_b0 , w_15847 );
and ( w_15847 , w_15846 , \4377_b1 );
or ( \4972_b1 , \4971_b1 , w_15849 );
not ( w_15849 , w_15850 );
and ( \4972_b0 , \4971_b0 , w_15851 );
and ( w_15850 ,  , w_15851 );
buf ( w_15849 , \4849_b1 );
not ( w_15849 , w_15852 );
not (  , w_15853 );
and ( w_15852 , w_15853 , \4849_b0 );
or ( \4973_b1 , \3943_b1 , \4156_b1 );
not ( \4156_b1 , w_15854 );
and ( \4973_b0 , \3943_b0 , w_15855 );
and ( w_15854 , w_15855 , \4156_b0 );
or ( \4974_b1 , \4972_b1 , \4973_b1 );
xor ( \4974_b0 , \4972_b0 , w_15856 );
not ( w_15856 , w_15857 );
and ( w_15857 , \4973_b1 , \4973_b0 );
or ( \4975_b1 , \4254_b1 , w_15858 );
or ( \4975_b0 , \4254_b0 , \4949_b0 );
not ( \4949_b0 , w_15859 );
and ( w_15859 , w_15858 , \4949_b1 );
or ( \4976_b1 , \4267_b1 , \3994_b1 );
not ( \3994_b1 , w_15860 );
and ( \4976_b0 , \4267_b0 , w_15861 );
and ( w_15860 , w_15861 , \3994_b0 );
or ( \4977_b1 , \4156_b1 , \4099_b1 );
not ( \4099_b1 , w_15862 );
and ( \4977_b0 , \4156_b0 , w_15863 );
and ( w_15862 , w_15863 , \4099_b0 );
or ( \4978_b1 , \4976_b1 , w_15865 );
not ( w_15865 , w_15866 );
and ( \4978_b0 , \4976_b0 , w_15867 );
and ( w_15866 ,  , w_15867 );
buf ( w_15865 , \4977_b1 );
not ( w_15865 , w_15868 );
not (  , w_15869 );
and ( w_15868 , w_15869 , \4977_b0 );
or ( \4979_b1 , \4978_b1 , w_15870 );
or ( \4979_b0 , \4978_b0 , \4950_b0 );
not ( \4950_b0 , w_15871 );
and ( w_15871 , w_15870 , \4950_b1 );
or ( \4980_b1 , \4975_b1 , w_15873 );
not ( w_15873 , w_15874 );
and ( \4980_b0 , \4975_b0 , w_15875 );
and ( w_15874 ,  , w_15875 );
buf ( w_15873 , \4979_b1 );
not ( w_15873 , w_15876 );
not (  , w_15877 );
and ( w_15876 , w_15877 , \4979_b0 );
or ( \4981_b1 , \4974_b1 , \4980_b1 );
xor ( \4981_b0 , \4974_b0 , w_15878 );
not ( w_15878 , w_15879 );
and ( w_15879 , \4980_b1 , \4980_b0 );
or ( \4982_b1 , \4970_b1 , \4981_b1 );
xor ( \4982_b0 , \4970_b0 , w_15880 );
not ( w_15880 , w_15881 );
and ( w_15881 , \4981_b1 , \4981_b0 );
or ( \4983_b1 , \4964_b1 , w_15883 );
not ( w_15883 , w_15884 );
and ( \4983_b0 , \4964_b0 , w_15885 );
and ( w_15884 ,  , w_15885 );
buf ( w_15883 , \4982_b1 );
not ( w_15883 , w_15886 );
not (  , w_15887 );
and ( w_15886 , w_15887 , \4982_b0 );
buf ( \4985_b1 , \4984_b1 );
not ( \4985_b1 , w_15888 );
not ( \4985_b0 , w_15889 );
and ( w_15888 , w_15889 , \4984_b0 );
or ( \4986_b1 , \4586_b1 , \4598_b1 );
xor ( \4986_b0 , \4586_b0 , w_15890 );
not ( w_15890 , w_15891 );
and ( w_15891 , \4598_b1 , \4598_b0 );
or ( \4987_b1 , \4986_b1 , w_15892 );
xor ( \4987_b0 , \4986_b0 , w_15894 );
not ( w_15894 , w_15895 );
and ( w_15895 , w_15892 , w_15893 );
buf ( w_15892 , \4610_b1 );
not ( w_15892 , w_15896 );
not ( w_15893 , w_15897 );
and ( w_15896 , w_15897 , \4610_b0 );
buf ( \4988_b1 , \4676_b1 );
not ( \4988_b1 , w_15898 );
not ( \4988_b0 , w_15899 );
and ( w_15898 , w_15899 , \4676_b0 );
buf ( \4989_b1 , \4659_b1 );
not ( \4989_b1 , w_15900 );
not ( \4989_b0 , w_15901 );
and ( w_15900 , w_15901 , \4659_b0 );
buf ( \4990_b1 , \4989_b1 );
not ( \4990_b1 , w_15902 );
not ( \4990_b0 , w_15903 );
and ( w_15902 , w_15903 , \4989_b0 );
or ( \4991_b1 , \4988_b1 , w_15904 );
or ( \4991_b0 , \4988_b0 , \4990_b0 );
not ( \4990_b0 , w_15905 );
and ( w_15905 , w_15904 , \4990_b1 );
or ( \4992_b1 , \4675_b1 , w_15907 );
not ( w_15907 , w_15908 );
and ( \4992_b0 , \4675_b0 , w_15909 );
and ( w_15908 ,  , w_15909 );
buf ( w_15907 , \4659_b1 );
not ( w_15907 , w_15910 );
not (  , w_15911 );
and ( w_15910 , w_15911 , \4659_b0 );
or ( \4993_b1 , \4991_b1 , w_15913 );
not ( w_15913 , w_15914 );
and ( \4993_b0 , \4991_b0 , w_15915 );
and ( w_15914 ,  , w_15915 );
buf ( w_15913 , \4992_b1 );
not ( w_15913 , w_15916 );
not (  , w_15917 );
and ( w_15916 , w_15917 , \4992_b0 );
buf ( \4994_b1 , \4993_b1 );
not ( \4994_b1 , w_15918 );
not ( \4994_b0 , w_15919 );
and ( w_15918 , w_15919 , \4993_b0 );
buf ( \4995_b1 , \4649_b1 );
not ( \4995_b1 , w_15920 );
not ( \4995_b0 , w_15921 );
and ( w_15920 , w_15921 , \4649_b0 );
buf ( \4996_b1 , \4995_b1 );
not ( \4996_b1 , w_15922 );
not ( \4996_b0 , w_15923 );
and ( w_15922 , w_15923 , \4995_b0 );
or ( \4997_b1 , \4994_b1 , \4996_b1 );
not ( \4996_b1 , w_15924 );
and ( \4997_b0 , \4994_b0 , w_15925 );
and ( w_15924 , w_15925 , \4996_b0 );
or ( \4998_b1 , \4993_b1 , \4995_b1 );
not ( \4995_b1 , w_15926 );
and ( \4998_b0 , \4993_b0 , w_15927 );
and ( w_15926 , w_15927 , \4995_b0 );
or ( \4999_b1 , \4997_b1 , w_15929 );
not ( w_15929 , w_15930 );
and ( \4999_b0 , \4997_b0 , w_15931 );
and ( w_15930 ,  , w_15931 );
buf ( w_15929 , \4998_b1 );
not ( w_15929 , w_15932 );
not (  , w_15933 );
and ( w_15932 , w_15933 , \4998_b0 );
or ( \5000_b1 , \4987_b1 , \4999_b1 );
xor ( \5000_b0 , \4987_b0 , w_15934 );
not ( w_15934 , w_15935 );
and ( w_15935 , \4999_b1 , \4999_b0 );
buf ( \5001_b1 , \4045_b1 );
not ( \5001_b1 , w_15936 );
not ( \5001_b0 , w_15937 );
and ( w_15936 , w_15937 , \4045_b0 );
buf ( \5002_b1 , \4089_b1 );
not ( \5002_b1 , w_15938 );
not ( \5002_b0 , w_15939 );
and ( w_15938 , w_15939 , \4089_b0 );
or ( \5003_b1 , \5001_b1 , w_15940 );
or ( \5003_b0 , \5001_b0 , \5002_b0 );
not ( \5002_b0 , w_15941 );
and ( w_15941 , w_15940 , \5002_b1 );
or ( \5004_b1 , \4088_b1 , w_15943 );
not ( w_15943 , w_15944 );
and ( \5004_b0 , \4088_b0 , w_15945 );
and ( w_15944 ,  , w_15945 );
buf ( w_15943 , \4286_b1 );
not ( w_15943 , w_15946 );
not (  , w_15947 );
and ( w_15946 , w_15947 , \4286_b0 );
or ( \5005_b1 , \5003_b1 , w_15949 );
not ( w_15949 , w_15950 );
and ( \5005_b0 , \5003_b0 , w_15951 );
and ( w_15950 ,  , w_15951 );
buf ( w_15949 , \5004_b1 );
not ( w_15949 , w_15952 );
not (  , w_15953 );
and ( w_15952 , w_15953 , \5004_b0 );
buf ( \5006_b1 , \5005_b1 );
not ( \5006_b1 , w_15954 );
not ( \5006_b0 , w_15955 );
and ( w_15954 , w_15955 , \5005_b0 );
buf ( \5007_b1 , \4437_b1 );
not ( \5007_b1 , w_15956 );
not ( \5007_b0 , w_15957 );
and ( w_15956 , w_15957 , \4437_b0 );
or ( \5008_b1 , \5006_b1 , w_15958 );
or ( \5008_b0 , \5006_b0 , \5007_b0 );
not ( \5007_b0 , w_15959 );
and ( w_15959 , w_15958 , \5007_b1 );
buf ( \5009_b1 , \4047_b1 );
not ( \5009_b1 , w_15960 );
not ( \5009_b0 , w_15961 );
and ( w_15960 , w_15961 , \4047_b0 );
buf ( \5010_b1 , \4089_b1 );
not ( \5010_b1 , w_15962 );
not ( \5010_b0 , w_15963 );
and ( w_15962 , w_15963 , \4089_b0 );
or ( \5011_b1 , \5009_b1 , w_15964 );
or ( \5011_b0 , \5009_b0 , \5010_b0 );
not ( \5010_b0 , w_15965 );
and ( w_15965 , w_15964 , \5010_b1 );
or ( \5012_b1 , \4088_b1 , w_15967 );
not ( w_15967 , w_15968 );
and ( \5012_b0 , \4088_b0 , w_15969 );
and ( w_15968 ,  , w_15969 );
buf ( w_15967 , \4178_b1 );
not ( w_15967 , w_15970 );
not (  , w_15971 );
and ( w_15970 , w_15971 , \4178_b0 );
or ( \5013_b1 , \5011_b1 , w_15973 );
not ( w_15973 , w_15974 );
and ( \5013_b0 , \5011_b0 , w_15975 );
and ( w_15974 ,  , w_15975 );
buf ( w_15973 , \5012_b1 );
not ( w_15973 , w_15976 );
not (  , w_15977 );
and ( w_15976 , w_15977 , \5012_b0 );
or ( \5014_b1 , \4596_b1 , w_15979 );
not ( w_15979 , w_15980 );
and ( \5014_b0 , \4596_b0 , w_15981 );
and ( w_15980 ,  , w_15981 );
buf ( w_15979 , \5013_b1 );
not ( w_15979 , w_15982 );
not (  , w_15983 );
and ( w_15982 , w_15983 , \5013_b0 );
or ( \5015_b1 , \5008_b1 , w_15985 );
not ( w_15985 , w_15986 );
and ( \5015_b0 , \5008_b0 , w_15987 );
and ( w_15986 ,  , w_15987 );
buf ( w_15985 , \5014_b1 );
not ( w_15985 , w_15988 );
not (  , w_15989 );
and ( w_15988 , w_15989 , \5014_b0 );
buf ( \5016_b1 , \1395_b1 );
buf ( \5016_b0 , \1395_b0 );
buf ( \5017_b1 , \5016_b1 );
not ( \5017_b1 , w_15990 );
not ( \5017_b0 , w_15991 );
and ( w_15990 , w_15991 , \5016_b0 );
or ( \5018_b1 , \5017_b1 , w_15993 );
not ( w_15993 , w_15994 );
and ( \5018_b0 , \5017_b0 , w_15995 );
and ( w_15994 ,  , w_15995 );
buf ( w_15993 , \3617_b1 );
not ( w_15993 , w_15996 );
not (  , w_15997 );
and ( w_15996 , w_15997 , \3617_b0 );
buf ( \5019_b1 , \5018_b1 );
buf ( \5019_b0 , \5018_b0 );
buf ( \5020_b1 , \5019_b1 );
buf ( \5020_b0 , \5019_b0 );
buf ( \5021_b1 , \3617_b1 );
buf ( \5021_b0 , \3617_b0 );
or ( \5022_b1 , \5020_b1 , w_15998 );
or ( \5022_b0 , \5020_b0 , \5021_b0 );
not ( \5021_b0 , w_15999 );
and ( w_15999 , w_15998 , \5021_b1 );
buf ( \5023_b1 , \5016_b1 );
not ( \5023_b1 , w_16000 );
not ( \5023_b0 , w_16001 );
and ( w_16000 , w_16001 , \5016_b0 );
buf ( \5024_b1 , \5023_b1 );
not ( \5024_b1 , w_16002 );
not ( \5024_b0 , w_16003 );
and ( w_16002 , w_16003 , \5023_b0 );
or ( \5025_b1 , \5022_b1 , w_16005 );
not ( w_16005 , w_16006 );
and ( \5025_b0 , \5022_b0 , w_16007 );
and ( w_16006 ,  , w_16007 );
buf ( w_16005 , \5024_b1 );
not ( w_16005 , w_16008 );
not (  , w_16009 );
and ( w_16008 , w_16009 , \5024_b0 );
or ( \5026_b1 , \5015_b1 , w_16011 );
not ( w_16011 , w_16012 );
and ( \5026_b0 , \5015_b0 , w_16013 );
and ( w_16012 ,  , w_16013 );
buf ( w_16011 , \5025_b1 );
not ( w_16011 , w_16014 );
not (  , w_16015 );
and ( w_16014 , w_16015 , \5025_b0 );
buf ( \5027_b1 , \4019_b1 );
not ( \5027_b1 , w_16016 );
not ( \5027_b0 , w_16017 );
and ( w_16016 , w_16017 , \4019_b0 );
buf ( \5028_b1 , \4267_b1 );
not ( \5028_b1 , w_16018 );
not ( \5028_b0 , w_16019 );
and ( w_16018 , w_16019 , \4267_b0 );
or ( \5029_b1 , \5027_b1 , w_16020 );
or ( \5029_b0 , \5027_b0 , \5028_b0 );
not ( \5028_b0 , w_16021 );
and ( w_16021 , w_16020 , \5028_b1 );
or ( \5030_b1 , \4308_b1 , w_16023 );
not ( w_16023 , w_16024 );
and ( \5030_b0 , \4308_b0 , w_16025 );
and ( w_16024 ,  , w_16025 );
buf ( w_16023 , \4585_b1 );
not ( w_16023 , w_16026 );
not (  , w_16027 );
and ( w_16026 , w_16027 , \4585_b0 );
or ( \5031_b1 , \5029_b1 , w_16029 );
not ( w_16029 , w_16030 );
and ( \5031_b0 , \5029_b0 , w_16031 );
and ( w_16030 ,  , w_16031 );
buf ( w_16029 , \5030_b1 );
not ( w_16029 , w_16032 );
not (  , w_16033 );
and ( w_16032 , w_16033 , \5030_b0 );
buf ( \5032_b1 , \5031_b1 );
not ( \5032_b1 , w_16034 );
not ( \5032_b0 , w_16035 );
and ( w_16034 , w_16035 , \5031_b0 );
buf ( \5033_b1 , \4253_b1 );
not ( \5033_b1 , w_16036 );
not ( \5033_b0 , w_16037 );
and ( w_16036 , w_16037 , \4253_b0 );
or ( \5034_b1 , \5032_b1 , w_16038 );
or ( \5034_b0 , \5032_b0 , \5033_b0 );
not ( \5033_b0 , w_16039 );
and ( w_16039 , w_16038 , \5033_b1 );
or ( \5035_b1 , \4644_b1 , w_16041 );
not ( w_16041 , w_16042 );
and ( \5035_b0 , \4644_b0 , w_16043 );
and ( w_16042 ,  , w_16043 );
buf ( w_16041 , \4742_b1 );
not ( w_16041 , w_16044 );
not (  , w_16045 );
and ( w_16044 , w_16045 , \4742_b0 );
or ( \5036_b1 , \5034_b1 , w_16047 );
not ( w_16047 , w_16048 );
and ( \5036_b0 , \5034_b0 , w_16049 );
and ( w_16048 ,  , w_16049 );
buf ( w_16047 , \5035_b1 );
not ( w_16047 , w_16050 );
not (  , w_16051 );
and ( w_16050 , w_16051 , \5035_b0 );
buf ( \5037_b1 , \5036_b1 );
not ( \5037_b1 , w_16052 );
not ( \5037_b0 , w_16053 );
and ( w_16052 , w_16053 , \5036_b0 );
or ( \5038_b1 , \5026_b1 , \5037_b1 );
xor ( \5038_b0 , \5026_b0 , w_16054 );
not ( w_16054 , w_16055 );
and ( w_16055 , \5037_b1 , \5037_b0 );
or ( \5039_b1 , \5038_b1 , \4676_b1 );
not ( \4676_b1 , w_16056 );
and ( \5039_b0 , \5038_b0 , w_16057 );
and ( w_16056 , w_16057 , \4676_b0 );
or ( \5040_b1 , \5026_b1 , \5037_b1 );
not ( \5037_b1 , w_16058 );
and ( \5040_b0 , \5026_b0 , w_16059 );
and ( w_16058 , w_16059 , \5037_b0 );
or ( \5041_b1 , \5039_b1 , w_16060 );
or ( \5041_b0 , \5039_b0 , \5040_b0 );
not ( \5040_b0 , w_16061 );
and ( w_16061 , w_16060 , \5040_b1 );
or ( \5042_b1 , \5000_b1 , \5041_b1 );
not ( \5041_b1 , w_16062 );
and ( \5042_b0 , \5000_b0 , w_16063 );
and ( w_16062 , w_16063 , \5041_b0 );
or ( \5043_b1 , \4987_b1 , \4999_b1 );
not ( \4999_b1 , w_16064 );
and ( \5043_b0 , \4987_b0 , w_16065 );
and ( w_16064 , w_16065 , \4999_b0 );
or ( \5044_b1 , \5042_b1 , w_16066 );
or ( \5044_b0 , \5042_b0 , \5043_b0 );
not ( \5043_b0 , w_16067 );
and ( w_16067 , w_16066 , \5043_b1 );
or ( \5045_b1 , \4413_b1 , \4580_b1 );
xor ( \5045_b0 , \4413_b0 , w_16068 );
not ( w_16068 , w_16069 );
and ( w_16069 , \4580_b1 , \4580_b0 );
or ( \5046_b1 , \5045_b1 , w_16070 );
xor ( \5046_b0 , \5045_b0 , w_16072 );
not ( w_16072 , w_16073 );
and ( w_16073 , w_16070 , w_16071 );
buf ( w_16070 , \4612_b1 );
not ( w_16070 , w_16074 );
not ( w_16071 , w_16075 );
and ( w_16074 , w_16075 , \4612_b0 );
or ( \5047_b1 , \4549_b1 , \4564_b1 );
xor ( \5047_b0 , \4549_b0 , w_16076 );
not ( w_16076 , w_16077 );
and ( w_16077 , \4564_b1 , \4564_b0 );
or ( \5048_b1 , \5047_b1 , w_16078 );
xor ( \5048_b0 , \5047_b0 , w_16080 );
not ( w_16080 , w_16081 );
and ( w_16081 , w_16078 , w_16079 );
buf ( w_16078 , \4578_b1 );
not ( w_16078 , w_16082 );
not ( w_16079 , w_16083 );
and ( w_16082 , w_16083 , \4578_b0 );
buf ( \5049_b1 , \5048_b1 );
not ( \5049_b1 , w_16084 );
not ( \5049_b0 , w_16085 );
and ( w_16084 , w_16085 , \5048_b0 );
buf ( \5050_b1 , \5049_b1 );
not ( \5050_b1 , w_16086 );
not ( \5050_b0 , w_16087 );
and ( w_16086 , w_16087 , \5049_b0 );
buf ( \5051_b1 , \5013_b1 );
not ( \5051_b1 , w_16088 );
not ( \5051_b0 , w_16089 );
and ( w_16088 , w_16089 , \5013_b0 );
buf ( \5052_b1 , \4437_b1 );
not ( \5052_b1 , w_16090 );
not ( \5052_b0 , w_16091 );
and ( w_16090 , w_16091 , \4437_b0 );
or ( \5053_b1 , \5051_b1 , w_16092 );
or ( \5053_b0 , \5051_b0 , \5052_b0 );
not ( \5052_b0 , w_16093 );
and ( w_16093 , w_16092 , \5052_b1 );
or ( \5054_b1 , \4331_b1 , w_16095 );
not ( w_16095 , w_16096 );
and ( \5054_b0 , \4331_b0 , w_16097 );
and ( w_16096 ,  , w_16097 );
buf ( w_16095 , \4592_b1 );
not ( w_16095 , w_16098 );
not (  , w_16099 );
and ( w_16098 , w_16099 , \4592_b0 );
or ( \5055_b1 , \5053_b1 , w_16101 );
not ( w_16101 , w_16102 );
and ( \5055_b0 , \5053_b0 , w_16103 );
and ( w_16102 ,  , w_16103 );
buf ( w_16101 , \5054_b1 );
not ( w_16101 , w_16104 );
not (  , w_16105 );
and ( w_16104 , w_16105 , \5054_b0 );
buf ( \5056_b1 , \5055_b1 );
not ( \5056_b1 , w_16106 );
not ( \5056_b0 , w_16107 );
and ( w_16106 , w_16107 , \5055_b0 );
buf ( \5057_b1 , \3943_b1 );
not ( \5057_b1 , w_16108 );
not ( \5057_b0 , w_16109 );
and ( w_16108 , w_16109 , \3943_b0 );
buf ( \5058_b1 , \4069_b1 );
not ( \5058_b1 , w_16110 );
not ( \5058_b0 , w_16111 );
and ( w_16110 , w_16111 , \4069_b0 );
or ( \5059_b1 , \5057_b1 , w_16112 );
or ( \5059_b0 , \5057_b0 , \5058_b0 );
not ( \5058_b0 , w_16113 );
and ( w_16113 , w_16112 , \5058_b1 );
buf ( \5060_b1 , \4069_b1 );
not ( \5060_b1 , w_16114 );
not ( \5060_b0 , w_16115 );
and ( w_16114 , w_16115 , \4069_b0 );
or ( \5061_b1 , \5060_b1 , w_16117 );
not ( w_16117 , w_16118 );
and ( \5061_b0 , \5060_b0 , w_16119 );
and ( w_16118 ,  , w_16119 );
buf ( w_16117 , \4147_b1 );
not ( w_16117 , w_16120 );
not (  , w_16121 );
and ( w_16120 , w_16121 , \4147_b0 );
or ( \5062_b1 , \5059_b1 , w_16123 );
not ( w_16123 , w_16124 );
and ( \5062_b0 , \5059_b0 , w_16125 );
and ( w_16124 ,  , w_16125 );
buf ( w_16123 , \5061_b1 );
not ( w_16123 , w_16126 );
not (  , w_16127 );
and ( w_16126 , w_16127 , \5061_b0 );
buf ( \5063_b1 , \5062_b1 );
not ( \5063_b1 , w_16128 );
not ( \5063_b0 , w_16129 );
and ( w_16128 , w_16129 , \5062_b0 );
buf ( \5064_b1 , \4065_b1 );
not ( \5064_b1 , w_16130 );
not ( \5064_b0 , w_16131 );
and ( w_16130 , w_16131 , \4065_b0 );
or ( \5065_b1 , \5063_b1 , w_16132 );
or ( \5065_b0 , \5063_b0 , \5064_b0 );
not ( \5064_b0 , w_16133 );
and ( w_16133 , w_16132 , \5064_b1 );
or ( \5066_b1 , \4055_b1 , w_16135 );
not ( w_16135 , w_16136 );
and ( \5066_b0 , \4055_b0 , w_16137 );
and ( w_16136 ,  , w_16137 );
buf ( w_16135 , \4556_b1 );
not ( w_16135 , w_16138 );
not (  , w_16139 );
and ( w_16138 , w_16139 , \4556_b0 );
or ( \5067_b1 , \5065_b1 , w_16141 );
not ( w_16141 , w_16142 );
and ( \5067_b0 , \5065_b0 , w_16143 );
and ( w_16142 ,  , w_16143 );
buf ( w_16141 , \5066_b1 );
not ( w_16141 , w_16144 );
not (  , w_16145 );
and ( w_16144 , w_16145 , \5066_b0 );
buf ( \5068_b1 , \5067_b1 );
not ( \5068_b1 , w_16146 );
not ( \5068_b0 , w_16147 );
and ( w_16146 , w_16147 , \5067_b0 );
or ( \5069_b1 , \5056_b1 , w_16148 );
or ( \5069_b0 , \5056_b0 , \5068_b0 );
not ( \5068_b0 , w_16149 );
and ( w_16149 , w_16148 , \5068_b1 );
or ( \5070_b1 , \5067_b1 , w_16150 );
or ( \5070_b0 , \5067_b0 , \5055_b0 );
not ( \5055_b0 , w_16151 );
and ( w_16151 , w_16150 , \5055_b1 );
buf ( \5071_b1 , \4041_b1 );
not ( \5071_b1 , w_16152 );
not ( \5071_b0 , w_16153 );
and ( w_16152 , w_16153 , \4041_b0 );
buf ( \5072_b1 , \4142_b1 );
not ( \5072_b1 , w_16154 );
not ( \5072_b0 , w_16155 );
and ( w_16154 , w_16155 , \4142_b0 );
or ( \5073_b1 , \5071_b1 , w_16156 );
or ( \5073_b0 , \5071_b0 , \5072_b0 );
not ( \5072_b0 , w_16157 );
and ( w_16157 , w_16156 , \5072_b1 );
or ( \5074_b1 , \4109_b1 , w_16159 );
not ( w_16159 , w_16160 );
and ( \5074_b0 , \4109_b0 , w_16161 );
and ( w_16160 ,  , w_16161 );
buf ( w_16159 , \4238_b1 );
not ( w_16159 , w_16162 );
not (  , w_16163 );
and ( w_16162 , w_16163 , \4238_b0 );
or ( \5075_b1 , \5073_b1 , w_16165 );
not ( w_16165 , w_16166 );
and ( \5075_b0 , \5073_b0 , w_16167 );
and ( w_16166 ,  , w_16167 );
buf ( w_16165 , \5074_b1 );
not ( w_16165 , w_16168 );
not (  , w_16169 );
and ( w_16168 , w_16169 , \5074_b0 );
buf ( \5076_b1 , \5075_b1 );
not ( \5076_b1 , w_16170 );
not ( \5076_b0 , w_16171 );
and ( w_16170 , w_16171 , \5075_b0 );
buf ( \5077_b1 , \4136_b1 );
not ( \5077_b1 , w_16172 );
not ( \5077_b0 , w_16173 );
and ( w_16172 , w_16173 , \4136_b0 );
or ( \5078_b1 , \5076_b1 , w_16174 );
or ( \5078_b0 , \5076_b0 , \5077_b0 );
not ( \5077_b0 , w_16175 );
and ( w_16175 , w_16174 , \5077_b1 );
or ( \5079_b1 , \4140_b1 , w_16177 );
not ( w_16177 , w_16178 );
and ( \5079_b0 , \4140_b0 , w_16179 );
and ( w_16178 ,  , w_16179 );
buf ( w_16177 , \4573_b1 );
not ( w_16177 , w_16180 );
not (  , w_16181 );
and ( w_16180 , w_16181 , \4573_b0 );
or ( \5080_b1 , \5078_b1 , w_16183 );
not ( w_16183 , w_16184 );
and ( \5080_b0 , \5078_b0 , w_16185 );
and ( w_16184 ,  , w_16185 );
buf ( w_16183 , \5079_b1 );
not ( w_16183 , w_16186 );
not (  , w_16187 );
and ( w_16186 , w_16187 , \5079_b0 );
or ( \5081_b1 , \5070_b1 , w_16189 );
not ( w_16189 , w_16190 );
and ( \5081_b0 , \5070_b0 , w_16191 );
and ( w_16190 ,  , w_16191 );
buf ( w_16189 , \5080_b1 );
not ( w_16189 , w_16192 );
not (  , w_16193 );
and ( w_16192 , w_16193 , \5080_b0 );
or ( \5082_b1 , \5069_b1 , w_16195 );
not ( w_16195 , w_16196 );
and ( \5082_b0 , \5069_b0 , w_16197 );
and ( w_16196 ,  , w_16197 );
buf ( w_16195 , \5081_b1 );
not ( w_16195 , w_16198 );
not (  , w_16199 );
and ( w_16198 , w_16199 , \5081_b0 );
buf ( \5083_b1 , \5082_b1 );
not ( \5083_b1 , w_16200 );
not ( \5083_b0 , w_16201 );
and ( w_16200 , w_16201 , \5082_b0 );
or ( \5084_b1 , \5050_b1 , w_16202 );
or ( \5084_b0 , \5050_b0 , \5083_b0 );
not ( \5083_b0 , w_16203 );
and ( w_16203 , w_16202 , \5083_b1 );
buf ( \5085_b1 , \5082_b1 );
not ( \5085_b1 , w_16204 );
not ( \5085_b0 , w_16205 );
and ( w_16204 , w_16205 , \5082_b0 );
buf ( \5086_b1 , \5085_b1 );
not ( \5086_b1 , w_16206 );
not ( \5086_b0 , w_16207 );
and ( w_16206 , w_16207 , \5085_b0 );
buf ( \5087_b1 , \5048_b1 );
not ( \5087_b1 , w_16208 );
not ( \5087_b0 , w_16209 );
and ( w_16208 , w_16209 , \5048_b0 );
or ( \5088_b1 , \5086_b1 , w_16210 );
or ( \5088_b0 , \5086_b0 , \5087_b0 );
not ( \5087_b0 , w_16211 );
and ( w_16211 , w_16210 , \5087_b1 );
or ( \5089_b1 , \4156_b1 , \4023_b1 );
not ( \4023_b1 , w_16212 );
and ( \5089_b0 , \4156_b0 , w_16213 );
and ( w_16212 , w_16213 , \4023_b0 );
buf ( \5090_b1 , \5089_b1 );
not ( \5090_b1 , w_16214 );
not ( \5090_b0 , w_16215 );
and ( w_16214 , w_16215 , \5089_b0 );
or ( \5091_b1 , \3958_b1 , \4216_b1 );
not ( \4216_b1 , w_16216 );
and ( \5091_b0 , \3958_b0 , w_16217 );
and ( w_16216 , w_16217 , \4216_b0 );
buf ( \5092_b1 , \3958_b1 );
not ( \5092_b1 , w_16218 );
not ( \5092_b0 , w_16219 );
and ( w_16218 , w_16219 , \3958_b0 );
or ( \5093_b1 , \5092_b1 , \4213_b1 );
not ( \4213_b1 , w_16220 );
and ( \5093_b0 , \5092_b0 , w_16221 );
and ( w_16220 , w_16221 , \4213_b0 );
or ( \5094_b1 , \5091_b1 , w_16223 );
not ( w_16223 , w_16224 );
and ( \5094_b0 , \5091_b0 , w_16225 );
and ( w_16224 ,  , w_16225 );
buf ( w_16223 , \5093_b1 );
not ( w_16223 , w_16226 );
not (  , w_16227 );
and ( w_16226 , w_16227 , \5093_b0 );
buf ( \5095_b1 , \5094_b1 );
not ( \5095_b1 , w_16228 );
not ( \5095_b0 , w_16229 );
and ( w_16228 , w_16229 , \5094_b0 );
buf ( \5096_b1 , \4231_b1 );
not ( \5096_b1 , w_16230 );
not ( \5096_b0 , w_16231 );
and ( w_16230 , w_16231 , \4231_b0 );
or ( \5097_b1 , \5095_b1 , w_16232 );
or ( \5097_b0 , \5095_b0 , \5096_b0 );
not ( \5096_b0 , w_16233 );
and ( w_16233 , w_16232 , \5096_b1 );
or ( \5098_b1 , \4234_b1 , w_16235 );
not ( w_16235 , w_16236 );
and ( \5098_b0 , \4234_b0 , w_16237 );
and ( w_16236 ,  , w_16237 );
buf ( w_16235 , \4654_b1 );
not ( w_16235 , w_16238 );
not (  , w_16239 );
and ( w_16238 , w_16239 , \4654_b0 );
or ( \5099_b1 , \5097_b1 , w_16241 );
not ( w_16241 , w_16242 );
and ( \5099_b0 , \5097_b0 , w_16243 );
and ( w_16242 ,  , w_16243 );
buf ( w_16241 , \5098_b1 );
not ( w_16241 , w_16244 );
not (  , w_16245 );
and ( w_16244 , w_16245 , \5098_b0 );
buf ( \5100_b1 , \5099_b1 );
not ( \5100_b1 , w_16246 );
not ( \5100_b0 , w_16247 );
and ( w_16246 , w_16247 , \5099_b0 );
or ( \5101_b1 , \5090_b1 , w_16248 );
or ( \5101_b0 , \5090_b0 , \5100_b0 );
not ( \5100_b0 , w_16249 );
and ( w_16249 , w_16248 , \5100_b1 );
or ( \5102_b1 , \5099_b1 , w_16250 );
or ( \5102_b0 , \5099_b0 , \5089_b0 );
not ( \5089_b0 , w_16251 );
and ( w_16251 , w_16250 , \5089_b1 );
buf ( \5103_b1 , \4011_b1 );
not ( \5103_b1 , w_16252 );
not ( \5103_b0 , w_16253 );
and ( w_16252 , w_16253 , \4011_b0 );
buf ( \5104_b1 , \4176_b1 );
not ( \5104_b1 , w_16254 );
not ( \5104_b0 , w_16255 );
and ( w_16254 , w_16255 , \4176_b0 );
or ( \5105_b1 , \5103_b1 , w_16256 );
or ( \5105_b0 , \5103_b0 , \5104_b0 );
not ( \5104_b0 , w_16257 );
and ( w_16257 , w_16256 , \5104_b1 );
or ( \5106_b1 , \4172_b1 , w_16259 );
not ( w_16259 , w_16260 );
and ( \5106_b0 , \4172_b0 , w_16261 );
and ( w_16260 ,  , w_16261 );
buf ( w_16259 , \4270_b1 );
not ( w_16259 , w_16262 );
not (  , w_16263 );
and ( w_16262 , w_16263 , \4270_b0 );
or ( \5107_b1 , \5105_b1 , w_16265 );
not ( w_16265 , w_16266 );
and ( \5107_b0 , \5105_b0 , w_16267 );
and ( w_16266 ,  , w_16267 );
buf ( w_16265 , \5106_b1 );
not ( w_16265 , w_16268 );
not (  , w_16269 );
and ( w_16268 , w_16269 , \5106_b0 );
buf ( \5108_b1 , \5107_b1 );
not ( \5108_b1 , w_16270 );
not ( \5108_b0 , w_16271 );
and ( w_16270 , w_16271 , \5107_b0 );
buf ( \5109_b1 , \4194_b1 );
not ( \5109_b1 , w_16272 );
not ( \5109_b0 , w_16273 );
and ( w_16272 , w_16273 , \4194_b0 );
or ( \5110_b1 , \5108_b1 , w_16274 );
or ( \5110_b0 , \5108_b0 , \5109_b0 );
not ( \5109_b0 , w_16275 );
and ( w_16275 , w_16274 , \5109_b1 );
buf ( \5111_b1 , \4203_b1 );
not ( \5111_b1 , w_16276 );
not ( \5111_b0 , w_16277 );
and ( w_16276 , w_16277 , \4203_b0 );
or ( \5112_b1 , \4605_b1 , w_16279 );
not ( w_16279 , w_16280 );
and ( \5112_b0 , \4605_b0 , w_16281 );
and ( w_16280 ,  , w_16281 );
buf ( w_16279 , \5111_b1 );
not ( w_16279 , w_16282 );
not (  , w_16283 );
and ( w_16282 , w_16283 , \5111_b0 );
or ( \5113_b1 , \5110_b1 , w_16285 );
not ( w_16285 , w_16286 );
and ( \5113_b0 , \5110_b0 , w_16287 );
and ( w_16286 ,  , w_16287 );
buf ( w_16285 , \5112_b1 );
not ( w_16285 , w_16288 );
not (  , w_16289 );
and ( w_16288 , w_16289 , \5112_b0 );
or ( \5114_b1 , \5102_b1 , w_16291 );
not ( w_16291 , w_16292 );
and ( \5114_b0 , \5102_b0 , w_16293 );
and ( w_16292 ,  , w_16293 );
buf ( w_16291 , \5113_b1 );
not ( w_16291 , w_16294 );
not (  , w_16295 );
and ( w_16294 , w_16295 , \5113_b0 );
or ( \5115_b1 , \5101_b1 , w_16297 );
not ( w_16297 , w_16298 );
and ( \5115_b0 , \5101_b0 , w_16299 );
and ( w_16298 ,  , w_16299 );
buf ( w_16297 , \5114_b1 );
not ( w_16297 , w_16300 );
not (  , w_16301 );
and ( w_16300 , w_16301 , \5114_b0 );
or ( \5116_b1 , \5088_b1 , w_16303 );
not ( w_16303 , w_16304 );
and ( \5116_b0 , \5088_b0 , w_16305 );
and ( w_16304 ,  , w_16305 );
buf ( w_16303 , \5115_b1 );
not ( w_16303 , w_16306 );
not (  , w_16307 );
and ( w_16306 , w_16307 , \5115_b0 );
or ( \5117_b1 , \5084_b1 , w_16309 );
not ( w_16309 , w_16310 );
and ( \5117_b0 , \5084_b0 , w_16311 );
and ( w_16310 ,  , w_16311 );
buf ( w_16309 , \5116_b1 );
not ( w_16309 , w_16312 );
not (  , w_16313 );
and ( w_16312 , w_16313 , \5116_b0 );
or ( \5118_b1 , \5046_b1 , \5117_b1 );
xor ( \5118_b0 , \5046_b0 , w_16314 );
not ( w_16314 , w_16315 );
and ( w_16315 , \5117_b1 , \5117_b0 );
or ( \5119_b1 , \4679_b1 , \4631_b1 );
xor ( \5119_b0 , \4679_b0 , w_16316 );
not ( w_16316 , w_16317 );
and ( w_16317 , \4631_b1 , \4631_b0 );
buf ( \5120_b1 , \4638_b1 );
not ( \5120_b1 , w_16318 );
not ( \5120_b0 , w_16319 );
and ( w_16318 , w_16319 , \4638_b0 );
or ( \5121_b1 , \5119_b1 , \5120_b1 );
not ( \5120_b1 , w_16320 );
and ( \5121_b0 , \5119_b0 , w_16321 );
and ( w_16320 , w_16321 , \5120_b0 );
buf ( \5122_b1 , \5119_b1 );
not ( \5122_b1 , w_16322 );
not ( \5122_b0 , w_16323 );
and ( w_16322 , w_16323 , \5119_b0 );
or ( \5123_b1 , \5122_b1 , \4638_b1 );
not ( \4638_b1 , w_16324 );
and ( \5123_b0 , \5122_b0 , w_16325 );
and ( w_16324 , w_16325 , \4638_b0 );
or ( \5124_b1 , \5121_b1 , w_16327 );
not ( w_16327 , w_16328 );
and ( \5124_b0 , \5121_b0 , w_16329 );
and ( w_16328 ,  , w_16329 );
buf ( w_16327 , \5123_b1 );
not ( w_16327 , w_16330 );
not (  , w_16331 );
and ( w_16330 , w_16331 , \5123_b0 );
or ( \5125_b1 , \5118_b1 , w_16332 );
xor ( \5125_b0 , \5118_b0 , w_16334 );
not ( w_16334 , w_16335 );
and ( w_16335 , w_16332 , w_16333 );
buf ( w_16332 , \5124_b1 );
not ( w_16332 , w_16336 );
not ( w_16333 , w_16337 );
and ( w_16336 , w_16337 , \5124_b0 );
or ( \5126_b1 , \5044_b1 , \5125_b1 );
xor ( \5126_b0 , \5044_b0 , w_16338 );
not ( w_16338 , w_16339 );
and ( w_16339 , \5125_b1 , \5125_b0 );
buf ( \5127_b1 , \4480_b1 );
not ( \5127_b1 , w_16340 );
not ( \5127_b0 , w_16341 );
and ( w_16340 , w_16341 , \4480_b0 );
buf ( \5128_b1 , \4023_b1 );
not ( \5128_b1 , w_16342 );
not ( \5128_b0 , w_16343 );
and ( w_16342 , w_16343 , \4023_b0 );
buf ( \5129_b1 , \4267_b1 );
not ( \5129_b1 , w_16344 );
not ( \5129_b0 , w_16345 );
and ( w_16344 , w_16345 , \4267_b0 );
or ( \5130_b1 , \5128_b1 , w_16346 );
or ( \5130_b0 , \5128_b0 , \5129_b0 );
not ( \5129_b0 , w_16347 );
and ( w_16347 , w_16346 , \5129_b1 );
buf ( \5131_b1 , \4023_b1 );
not ( \5131_b1 , w_16348 );
not ( \5131_b0 , w_16349 );
and ( w_16348 , w_16349 , \4023_b0 );
or ( \5132_b1 , \4156_b1 , w_16351 );
not ( w_16351 , w_16352 );
and ( \5132_b0 , \4156_b0 , w_16353 );
and ( w_16352 ,  , w_16353 );
buf ( w_16351 , \5131_b1 );
not ( w_16351 , w_16354 );
not (  , w_16355 );
and ( w_16354 , w_16355 , \5131_b0 );
or ( \5133_b1 , \5130_b1 , w_16357 );
not ( w_16357 , w_16358 );
and ( \5133_b0 , \5130_b0 , w_16359 );
and ( w_16358 ,  , w_16359 );
buf ( w_16357 , \5132_b1 );
not ( w_16357 , w_16360 );
not (  , w_16361 );
and ( w_16360 , w_16361 , \5132_b0 );
buf ( \5134_b1 , \5133_b1 );
not ( \5134_b1 , w_16362 );
not ( \5134_b0 , w_16363 );
and ( w_16362 , w_16363 , \5133_b0 );
or ( \5135_b1 , \5127_b1 , w_16364 );
or ( \5135_b0 , \5127_b0 , \5134_b0 );
not ( \5134_b0 , w_16365 );
and ( w_16365 , w_16364 , \5134_b1 );
or ( \5136_b1 , \5031_b1 , w_16367 );
not ( w_16367 , w_16368 );
and ( \5136_b0 , \5031_b0 , w_16369 );
and ( w_16368 ,  , w_16369 );
buf ( w_16367 , \4273_b1 );
not ( w_16367 , w_16370 );
not (  , w_16371 );
and ( w_16370 , w_16371 , \4273_b0 );
or ( \5137_b1 , \5135_b1 , w_16373 );
not ( w_16373 , w_16374 );
and ( \5137_b0 , \5135_b0 , w_16375 );
and ( w_16374 ,  , w_16375 );
buf ( w_16373 , \5136_b1 );
not ( w_16373 , w_16376 );
not (  , w_16377 );
and ( w_16376 , w_16377 , \5136_b0 );
or ( \5138_b1 , \4156_b1 , \4026_b1 );
not ( \4026_b1 , w_16378 );
and ( \5138_b0 , \4156_b0 , w_16379 );
and ( w_16378 , w_16379 , \4026_b0 );
or ( \5139_b1 , \5137_b1 , w_16380 );
or ( \5139_b0 , \5137_b0 , \5138_b0 );
not ( \5138_b0 , w_16381 );
and ( w_16381 , w_16380 , \5138_b1 );
buf ( \5140_b1 , \4046_b1 );
not ( \5140_b1 , w_16382 );
not ( \5140_b0 , w_16383 );
and ( w_16382 , w_16383 , \4046_b0 );
buf ( \5141_b1 , \4284_b1 );
not ( \5141_b1 , w_16384 );
not ( \5141_b0 , w_16385 );
and ( w_16384 , w_16385 , \4284_b0 );
or ( \5142_b1 , \5140_b1 , w_16386 );
or ( \5142_b0 , \5140_b0 , \5141_b0 );
not ( \5141_b0 , w_16387 );
and ( w_16387 , w_16386 , \5141_b1 );
or ( \5143_b1 , \4177_b1 , w_16389 );
not ( w_16389 , w_16390 );
and ( \5143_b0 , \4177_b0 , w_16391 );
and ( w_16390 ,  , w_16391 );
buf ( w_16389 , \4256_b1 );
not ( w_16389 , w_16392 );
not (  , w_16393 );
and ( w_16392 , w_16393 , \4256_b0 );
or ( \5144_b1 , \5142_b1 , w_16395 );
not ( w_16395 , w_16396 );
and ( \5144_b0 , \5142_b0 , w_16397 );
and ( w_16396 ,  , w_16397 );
buf ( w_16395 , \5143_b1 );
not ( w_16395 , w_16398 );
not (  , w_16399 );
and ( w_16398 , w_16399 , \5143_b0 );
buf ( \5145_b1 , \5144_b1 );
not ( \5145_b1 , w_16400 );
not ( \5145_b0 , w_16401 );
and ( w_16400 , w_16401 , \5144_b0 );
buf ( \5146_b1 , \4194_b1 );
not ( \5146_b1 , w_16402 );
not ( \5146_b0 , w_16403 );
and ( w_16402 , w_16403 , \4194_b0 );
or ( \5147_b1 , \5145_b1 , w_16404 );
or ( \5147_b0 , \5145_b0 , \5146_b0 );
not ( \5146_b0 , w_16405 );
and ( w_16405 , w_16404 , \5146_b1 );
or ( \5148_b1 , \5107_b1 , w_16407 );
not ( w_16407 , w_16408 );
and ( \5148_b0 , \5107_b0 , w_16409 );
and ( w_16408 ,  , w_16409 );
buf ( w_16407 , \4204_b1 );
not ( w_16407 , w_16410 );
not (  , w_16411 );
and ( w_16410 , w_16411 , \4204_b0 );
or ( \5149_b1 , \5147_b1 , w_16413 );
not ( w_16413 , w_16414 );
and ( \5149_b0 , \5147_b0 , w_16415 );
and ( w_16414 ,  , w_16415 );
buf ( w_16413 , \5148_b1 );
not ( w_16413 , w_16416 );
not (  , w_16417 );
and ( w_16416 , w_16417 , \5148_b0 );
or ( \5150_b1 , \5139_b1 , w_16419 );
not ( w_16419 , w_16420 );
and ( \5150_b0 , \5139_b0 , w_16421 );
and ( w_16420 ,  , w_16421 );
buf ( w_16419 , \5149_b1 );
not ( w_16419 , w_16422 );
not (  , w_16423 );
and ( w_16422 , w_16423 , \5149_b0 );
or ( \5151_b1 , \5137_b1 , w_16425 );
not ( w_16425 , w_16426 );
and ( \5151_b0 , \5137_b0 , w_16427 );
and ( w_16426 ,  , w_16427 );
buf ( w_16425 , \5138_b1 );
not ( w_16425 , w_16428 );
not (  , w_16429 );
and ( w_16428 , w_16429 , \5138_b0 );
or ( \5152_b1 , \5150_b1 , w_16431 );
not ( w_16431 , w_16432 );
and ( \5152_b0 , \5150_b0 , w_16433 );
and ( w_16432 ,  , w_16433 );
buf ( w_16431 , \5151_b1 );
not ( w_16431 , w_16434 );
not (  , w_16435 );
and ( w_16434 , w_16435 , \5151_b0 );
buf ( \5153_b1 , \4042_b1 );
not ( \5153_b1 , w_16436 );
not ( \5153_b0 , w_16437 );
and ( w_16436 , w_16437 , \4042_b0 );
buf ( \5154_b1 , \4069_b1 );
not ( \5154_b1 , w_16438 );
not ( \5154_b0 , w_16439 );
and ( w_16438 , w_16439 , \4069_b0 );
or ( \5155_b1 , \5153_b1 , w_16440 );
or ( \5155_b0 , \5153_b0 , \5154_b0 );
not ( \5154_b0 , w_16441 );
and ( w_16441 , w_16440 , \5154_b1 );
or ( \5156_b1 , \5060_b1 , w_16443 );
not ( w_16443 , w_16444 );
and ( \5156_b0 , \5060_b0 , w_16445 );
and ( w_16444 ,  , w_16445 );
buf ( w_16443 , \4116_b1 );
not ( w_16443 , w_16446 );
not (  , w_16447 );
and ( w_16446 , w_16447 , \4116_b0 );
or ( \5157_b1 , \5155_b1 , w_16449 );
not ( w_16449 , w_16450 );
and ( \5157_b0 , \5155_b0 , w_16451 );
and ( w_16450 ,  , w_16451 );
buf ( w_16449 , \5156_b1 );
not ( w_16449 , w_16452 );
not (  , w_16453 );
and ( w_16452 , w_16453 , \5156_b0 );
buf ( \5158_b1 , \5157_b1 );
not ( \5158_b1 , w_16454 );
not ( \5158_b0 , w_16455 );
and ( w_16454 , w_16455 , \5157_b0 );
buf ( \5159_b1 , \4558_b1 );
not ( \5159_b1 , w_16456 );
not ( \5159_b0 , w_16457 );
and ( w_16456 , w_16457 , \4558_b0 );
or ( \5160_b1 , \5158_b1 , w_16458 );
or ( \5160_b0 , \5158_b0 , \5159_b0 );
not ( \5159_b0 , w_16459 );
and ( w_16459 , w_16458 , \5159_b1 );
or ( \5161_b1 , \4054_b1 , w_16461 );
not ( w_16461 , w_16462 );
and ( \5161_b0 , \4054_b0 , w_16463 );
and ( w_16462 ,  , w_16463 );
buf ( w_16461 , \5062_b1 );
not ( w_16461 , w_16464 );
not (  , w_16465 );
and ( w_16464 , w_16465 , \5062_b0 );
or ( \5162_b1 , \5160_b1 , w_16467 );
not ( w_16467 , w_16468 );
and ( \5162_b0 , \5160_b0 , w_16469 );
and ( w_16468 ,  , w_16469 );
buf ( w_16467 , \5161_b1 );
not ( w_16467 , w_16470 );
not (  , w_16471 );
and ( w_16470 , w_16471 , \5161_b0 );
buf ( \5163_b1 , \5162_b1 );
not ( \5163_b1 , w_16472 );
not ( \5163_b0 , w_16473 );
and ( w_16472 , w_16473 , \5162_b0 );
buf ( \5164_b1 , \4140_b1 );
not ( \5164_b1 , w_16474 );
not ( \5164_b0 , w_16475 );
and ( w_16474 , w_16475 , \4140_b0 );
buf ( \5165_b1 , \5075_b1 );
not ( \5165_b1 , w_16476 );
not ( \5165_b0 , w_16477 );
and ( w_16476 , w_16477 , \5075_b0 );
or ( \5166_b1 , \5164_b1 , w_16478 );
or ( \5166_b0 , \5164_b0 , \5165_b0 );
not ( \5165_b0 , w_16479 );
and ( w_16479 , w_16478 , \5165_b1 );
or ( \5167_b1 , \4217_b1 , \4109_b1 );
not ( \4109_b1 , w_16480 );
and ( \5167_b0 , \4217_b0 , w_16481 );
and ( w_16480 , w_16481 , \4109_b0 );
buf ( \5168_b1 , \4217_b1 );
not ( \5168_b1 , w_16482 );
not ( \5168_b0 , w_16483 );
and ( w_16482 , w_16483 , \4217_b0 );
or ( \5169_b1 , \5168_b1 , \4569_b1 );
not ( \4569_b1 , w_16484 );
and ( \5169_b0 , \5168_b0 , w_16485 );
and ( w_16484 , w_16485 , \4569_b0 );
or ( \5170_b1 , \5167_b1 , w_16487 );
not ( w_16487 , w_16488 );
and ( \5170_b0 , \5167_b0 , w_16489 );
and ( w_16488 ,  , w_16489 );
buf ( w_16487 , \5169_b1 );
not ( w_16487 , w_16490 );
not (  , w_16491 );
and ( w_16490 , w_16491 , \5169_b0 );
buf ( \5171_b1 , \5170_b1 );
not ( \5171_b1 , w_16492 );
not ( \5171_b0 , w_16493 );
and ( w_16492 , w_16493 , \5170_b0 );
or ( \5172_b1 , \5171_b1 , w_16495 );
not ( w_16495 , w_16496 );
and ( \5172_b0 , \5171_b0 , w_16497 );
and ( w_16496 ,  , w_16497 );
buf ( w_16495 , \4136_b1 );
not ( w_16495 , w_16498 );
not (  , w_16499 );
and ( w_16498 , w_16499 , \4136_b0 );
or ( \5173_b1 , \5166_b1 , w_16501 );
not ( w_16501 , w_16502 );
and ( \5173_b0 , \5166_b0 , w_16503 );
and ( w_16502 ,  , w_16503 );
buf ( w_16501 , \5172_b1 );
not ( w_16501 , w_16504 );
not (  , w_16505 );
and ( w_16504 , w_16505 , \5172_b0 );
buf ( \5174_b1 , \5173_b1 );
not ( \5174_b1 , w_16506 );
not ( \5174_b0 , w_16507 );
and ( w_16506 , w_16507 , \5173_b0 );
or ( \5175_b1 , \5163_b1 , w_16508 );
or ( \5175_b0 , \5163_b0 , \5174_b0 );
not ( \5174_b0 , w_16509 );
and ( w_16509 , w_16508 , \5174_b1 );
or ( \5176_b1 , \5173_b1 , w_16510 );
or ( \5176_b0 , \5173_b0 , \5162_b0 );
not ( \5162_b0 , w_16511 );
and ( w_16511 , w_16510 , \5162_b1 );
buf ( \5177_b1 , \4044_b1 );
not ( \5177_b1 , w_16512 );
not ( \5177_b0 , w_16513 );
and ( w_16512 , w_16513 , \4044_b0 );
buf ( \5178_b1 , \4548_b1 );
not ( \5178_b1 , w_16514 );
not ( \5178_b0 , w_16515 );
and ( w_16514 , w_16515 , \4548_b0 );
buf ( \5179_b1 , \5178_b1 );
not ( \5179_b1 , w_16516 );
not ( \5179_b0 , w_16517 );
and ( w_16516 , w_16517 , \5178_b0 );
or ( \5180_b1 , \5177_b1 , w_16518 );
or ( \5180_b0 , \5177_b0 , \5179_b0 );
not ( \5179_b0 , w_16519 );
and ( w_16519 , w_16518 , \5179_b1 );
or ( \5181_b1 , \4548_b1 , w_16521 );
not ( w_16521 , w_16522 );
and ( \5181_b0 , \4548_b0 , w_16523 );
and ( w_16522 ,  , w_16523 );
buf ( w_16521 , \4092_b1 );
not ( w_16521 , w_16524 );
not (  , w_16525 );
and ( w_16524 , w_16525 , \4092_b0 );
or ( \5182_b1 , \5180_b1 , w_16527 );
not ( w_16527 , w_16528 );
and ( \5182_b0 , \5180_b0 , w_16529 );
and ( w_16528 ,  , w_16529 );
buf ( w_16527 , \5181_b1 );
not ( w_16527 , w_16530 );
not (  , w_16531 );
and ( w_16530 , w_16531 , \5181_b0 );
buf ( \5183_b1 , \5182_b1 );
not ( \5183_b1 , w_16532 );
not ( \5183_b0 , w_16533 );
and ( w_16532 , w_16533 , \5182_b0 );
buf ( \5184_b1 , \4661_b1 );
not ( \5184_b1 , w_16534 );
not ( \5184_b0 , w_16535 );
and ( w_16534 , w_16535 , \4661_b0 );
or ( \5185_b1 , \5183_b1 , w_16536 );
or ( \5185_b0 , \5183_b0 , \5184_b0 );
not ( \5184_b0 , w_16537 );
and ( w_16537 , w_16536 , \5184_b1 );
buf ( \5186_b1 , \4669_b1 );
not ( \5186_b1 , w_16538 );
not ( \5186_b0 , w_16539 );
and ( w_16538 , w_16539 , \4669_b0 );
buf ( \5187_b1 , \4545_b1 );
not ( \5187_b1 , w_16540 );
not ( \5187_b0 , w_16541 );
and ( w_16540 , w_16541 , \4545_b0 );
or ( \5188_b1 , \5186_b1 , w_16543 );
not ( w_16543 , w_16544 );
and ( \5188_b0 , \5186_b0 , w_16545 );
and ( w_16544 ,  , w_16545 );
buf ( w_16543 , \5187_b1 );
not ( w_16543 , w_16546 );
not (  , w_16547 );
and ( w_16546 , w_16547 , \5187_b0 );
or ( \5189_b1 , \5185_b1 , w_16549 );
not ( w_16549 , w_16550 );
and ( \5189_b0 , \5185_b0 , w_16551 );
and ( w_16550 ,  , w_16551 );
buf ( w_16549 , \5188_b1 );
not ( w_16549 , w_16552 );
not (  , w_16553 );
and ( w_16552 , w_16553 , \5188_b0 );
or ( \5190_b1 , \5176_b1 , w_16555 );
not ( w_16555 , w_16556 );
and ( \5190_b0 , \5176_b0 , w_16557 );
and ( w_16556 ,  , w_16557 );
buf ( w_16555 , \5189_b1 );
not ( w_16555 , w_16558 );
not (  , w_16559 );
and ( w_16558 , w_16559 , \5189_b0 );
or ( \5191_b1 , \5175_b1 , w_16561 );
not ( w_16561 , w_16562 );
and ( \5191_b0 , \5175_b0 , w_16563 );
and ( w_16562 ,  , w_16563 );
buf ( w_16561 , \5190_b1 );
not ( w_16561 , w_16564 );
not (  , w_16565 );
and ( w_16564 , w_16565 , \5190_b0 );
or ( \5192_b1 , \5152_b1 , w_16566 );
or ( \5192_b0 , \5152_b0 , \5191_b0 );
not ( \5191_b0 , w_16567 );
and ( w_16567 , w_16566 , \5191_b1 );
or ( \5193_b1 , \5067_b1 , \5080_b1 );
xor ( \5193_b0 , \5067_b0 , w_16568 );
not ( w_16568 , w_16569 );
and ( w_16569 , \5080_b1 , \5080_b0 );
or ( \5194_b1 , \5193_b1 , \5055_b1 );
xor ( \5194_b0 , \5193_b0 , w_16570 );
not ( w_16570 , w_16571 );
and ( w_16571 , \5055_b1 , \5055_b0 );
or ( \5195_b1 , \5192_b1 , \5194_b1 );
not ( \5194_b1 , w_16572 );
and ( \5195_b0 , \5192_b0 , w_16573 );
and ( w_16572 , w_16573 , \5194_b0 );
or ( \5196_b1 , \5152_b1 , \5191_b1 );
not ( \5191_b1 , w_16574 );
and ( \5196_b0 , \5152_b0 , w_16575 );
and ( w_16574 , w_16575 , \5191_b0 );
or ( \5197_b1 , \5195_b1 , w_16577 );
not ( w_16577 , w_16578 );
and ( \5197_b0 , \5195_b0 , w_16579 );
and ( w_16578 ,  , w_16579 );
buf ( w_16577 , \5196_b1 );
not ( w_16577 , w_16580 );
not (  , w_16581 );
and ( w_16580 , w_16581 , \5196_b0 );
or ( \5198_b1 , \5082_b1 , \5048_b1 );
xor ( \5198_b0 , \5082_b0 , w_16582 );
not ( w_16582 , w_16583 );
and ( w_16583 , \5048_b1 , \5048_b0 );
or ( \5199_b1 , \5198_b1 , \5115_b1 );
xor ( \5199_b0 , \5198_b0 , w_16584 );
not ( w_16584 , w_16585 );
and ( w_16585 , \5115_b1 , \5115_b0 );
or ( \5200_b1 , \5197_b1 , \5199_b1 );
xor ( \5200_b0 , \5197_b0 , w_16586 );
not ( w_16586 , w_16587 );
and ( w_16587 , \5199_b1 , \5199_b0 );
or ( \5201_b1 , \4987_b1 , \4999_b1 );
xor ( \5201_b0 , \4987_b0 , w_16588 );
not ( w_16588 , w_16589 );
and ( w_16589 , \4999_b1 , \4999_b0 );
or ( \5202_b1 , \5201_b1 , \5041_b1 );
xor ( \5202_b0 , \5201_b0 , w_16590 );
not ( w_16590 , w_16591 );
and ( w_16591 , \5041_b1 , \5041_b0 );
or ( \5203_b1 , \5200_b1 , \5202_b1 );
not ( \5202_b1 , w_16592 );
and ( \5203_b0 , \5200_b0 , w_16593 );
and ( w_16592 , w_16593 , \5202_b0 );
or ( \5204_b1 , \5197_b1 , \5199_b1 );
not ( \5199_b1 , w_16594 );
and ( \5204_b0 , \5197_b0 , w_16595 );
and ( w_16594 , w_16595 , \5199_b0 );
or ( \5205_b1 , \5203_b1 , w_16596 );
or ( \5205_b0 , \5203_b0 , \5204_b0 );
not ( \5204_b0 , w_16597 );
and ( w_16597 , w_16596 , \5204_b1 );
or ( \5206_b1 , \5126_b1 , \5205_b1 );
xor ( \5206_b0 , \5126_b0 , w_16598 );
not ( w_16598 , w_16599 );
and ( w_16599 , \5205_b1 , \5205_b0 );
or ( \5207_b1 , \5089_b1 , \5113_b1 );
xor ( \5207_b0 , \5089_b0 , w_16600 );
not ( w_16600 , w_16601 );
and ( w_16601 , \5113_b1 , \5113_b0 );
or ( \5208_b1 , \5207_b1 , w_16602 );
xor ( \5208_b0 , \5207_b0 , w_16604 );
not ( w_16604 , w_16605 );
and ( w_16605 , w_16602 , w_16603 );
buf ( w_16602 , \5099_b1 );
not ( w_16602 , w_16606 );
not ( w_16603 , w_16607 );
and ( w_16606 , w_16607 , \5099_b0 );
or ( \5209_b1 , \4127_b1 , w_16609 );
not ( w_16609 , w_16610 );
and ( \5209_b0 , \4127_b0 , w_16611 );
and ( w_16610 ,  , w_16611 );
buf ( w_16609 , \4134_b1 );
not ( w_16609 , w_16612 );
not (  , w_16613 );
and ( w_16612 , w_16613 , \4134_b0 );
buf ( \5210_b1 , \5209_b1 );
not ( \5210_b1 , w_16614 );
not ( \5210_b0 , w_16615 );
and ( w_16614 , w_16615 , \5209_b0 );
buf ( \5211_b1 , \4011_b1 );
not ( \5211_b1 , w_16616 );
not ( \5211_b0 , w_16617 );
and ( w_16616 , w_16617 , \4011_b0 );
buf ( \5212_b1 , \4145_b1 );
not ( \5212_b1 , w_16618 );
not ( \5212_b0 , w_16619 );
and ( w_16618 , w_16619 , \4145_b0 );
or ( \5213_b1 , \5211_b1 , w_16620 );
or ( \5213_b0 , \5211_b0 , \5212_b0 );
not ( \5212_b0 , w_16621 );
and ( w_16621 , w_16620 , \5212_b1 );
or ( \5214_b1 , \4109_b1 , w_16623 );
not ( w_16623 , w_16624 );
and ( \5214_b0 , \4109_b0 , w_16625 );
and ( w_16624 ,  , w_16625 );
buf ( w_16623 , \4270_b1 );
not ( w_16623 , w_16626 );
not (  , w_16627 );
and ( w_16626 , w_16627 , \4270_b0 );
or ( \5215_b1 , \5213_b1 , w_16629 );
not ( w_16629 , w_16630 );
and ( \5215_b0 , \5213_b0 , w_16631 );
and ( w_16630 ,  , w_16631 );
buf ( w_16629 , \5214_b1 );
not ( w_16629 , w_16632 );
not (  , w_16633 );
and ( w_16632 , w_16633 , \5214_b0 );
buf ( \5216_b1 , \5215_b1 );
not ( \5216_b1 , w_16634 );
not ( \5216_b0 , w_16635 );
and ( w_16634 , w_16635 , \5215_b0 );
buf ( \5217_b1 , \5216_b1 );
not ( \5217_b1 , w_16636 );
not ( \5217_b0 , w_16637 );
and ( w_16636 , w_16637 , \5216_b0 );
or ( \5218_b1 , \5210_b1 , \5217_b1 );
not ( \5217_b1 , w_16638 );
and ( \5218_b0 , \5210_b0 , w_16639 );
and ( w_16638 , w_16639 , \5217_b0 );
or ( \5219_b1 , \5170_b1 , w_16641 );
not ( w_16641 , w_16642 );
and ( \5219_b0 , \5170_b0 , w_16643 );
and ( w_16642 ,  , w_16643 );
buf ( w_16641 , \4428_b1 );
not ( w_16641 , w_16644 );
not (  , w_16645 );
and ( w_16644 , w_16645 , \4428_b0 );
or ( \5220_b1 , \5218_b1 , w_16647 );
not ( w_16647 , w_16648 );
and ( \5220_b0 , \5218_b0 , w_16649 );
and ( w_16648 ,  , w_16649 );
buf ( w_16647 , \5219_b1 );
not ( w_16647 , w_16650 );
not (  , w_16651 );
and ( w_16650 , w_16651 , \5219_b0 );
buf ( \5221_b1 , \3943_b1 );
not ( \5221_b1 , w_16652 );
not ( \5221_b0 , w_16653 );
and ( w_16652 , w_16653 , \3943_b0 );
buf ( \5222_b1 , \5178_b1 );
not ( \5222_b1 , w_16654 );
not ( \5222_b0 , w_16655 );
and ( w_16654 , w_16655 , \5178_b0 );
or ( \5223_b1 , \5221_b1 , w_16656 );
or ( \5223_b0 , \5221_b0 , \5222_b0 );
not ( \5222_b0 , w_16657 );
and ( w_16657 , w_16656 , \5222_b1 );
or ( \5224_b1 , \4665_b1 , w_16659 );
not ( w_16659 , w_16660 );
and ( \5224_b0 , \4665_b0 , w_16661 );
and ( w_16660 ,  , w_16661 );
buf ( w_16659 , \4147_b1 );
not ( w_16659 , w_16662 );
not (  , w_16663 );
and ( w_16662 , w_16663 , \4147_b0 );
or ( \5225_b1 , \5223_b1 , w_16665 );
not ( w_16665 , w_16666 );
and ( \5225_b0 , \5223_b0 , w_16667 );
and ( w_16666 ,  , w_16667 );
buf ( w_16665 , \5224_b1 );
not ( w_16665 , w_16668 );
not (  , w_16669 );
and ( w_16668 , w_16669 , \5224_b0 );
buf ( \5226_b1 , \5225_b1 );
not ( \5226_b1 , w_16670 );
not ( \5226_b0 , w_16671 );
and ( w_16670 , w_16671 , \5225_b0 );
buf ( \5227_b1 , \4662_b1 );
not ( \5227_b1 , w_16672 );
not ( \5227_b0 , w_16673 );
and ( w_16672 , w_16673 , \4662_b0 );
or ( \5228_b1 , \5226_b1 , w_16674 );
or ( \5228_b0 , \5226_b0 , \5227_b0 );
not ( \5227_b0 , w_16675 );
and ( w_16675 , w_16674 , \5227_b1 );
or ( \5229_b1 , \4672_b1 , w_16677 );
not ( w_16677 , w_16678 );
and ( \5229_b0 , \4672_b0 , w_16679 );
and ( w_16678 ,  , w_16679 );
buf ( w_16677 , \5182_b1 );
not ( w_16677 , w_16680 );
not (  , w_16681 );
and ( w_16680 , w_16681 , \5182_b0 );
or ( \5230_b1 , \5228_b1 , w_16683 );
not ( w_16683 , w_16684 );
and ( \5230_b0 , \5228_b0 , w_16685 );
and ( w_16684 ,  , w_16685 );
buf ( w_16683 , \5229_b1 );
not ( w_16683 , w_16686 );
not (  , w_16687 );
and ( w_16686 , w_16687 , \5229_b0 );
buf ( \5231_b1 , \5230_b1 );
not ( \5231_b1 , w_16688 );
not ( \5231_b0 , w_16689 );
and ( w_16688 , w_16689 , \5230_b0 );
or ( \5232_b1 , \5220_b1 , \5231_b1 );
xor ( \5232_b0 , \5220_b0 , w_16690 );
not ( w_16690 , w_16691 );
and ( w_16691 , \5231_b1 , \5231_b0 );
buf ( \5233_b1 , \4041_b1 );
not ( \5233_b1 , w_16692 );
not ( \5233_b0 , w_16693 );
and ( w_16692 , w_16693 , \4041_b0 );
buf ( \5234_b1 , \4088_b1 );
not ( \5234_b1 , w_16694 );
not ( \5234_b0 , w_16695 );
and ( w_16694 , w_16695 , \4088_b0 );
buf ( \5235_b1 , \5234_b1 );
not ( \5235_b1 , w_16696 );
not ( \5235_b0 , w_16697 );
and ( w_16696 , w_16697 , \5234_b0 );
or ( \5236_b1 , \5233_b1 , w_16698 );
or ( \5236_b0 , \5233_b0 , \5235_b0 );
not ( \5235_b0 , w_16699 );
and ( w_16699 , w_16698 , \5235_b1 );
or ( \5237_b1 , \4088_b1 , w_16701 );
not ( w_16701 , w_16702 );
and ( \5237_b0 , \4088_b0 , w_16703 );
and ( w_16702 ,  , w_16703 );
buf ( w_16701 , \4238_b1 );
not ( w_16701 , w_16704 );
not (  , w_16705 );
and ( w_16704 , w_16705 , \4238_b0 );
or ( \5238_b1 , \5236_b1 , w_16707 );
not ( w_16707 , w_16708 );
and ( \5238_b0 , \5236_b0 , w_16709 );
and ( w_16708 ,  , w_16709 );
buf ( w_16707 , \5237_b1 );
not ( w_16707 , w_16710 );
not (  , w_16711 );
and ( w_16710 , w_16711 , \5237_b0 );
or ( \5239_b1 , \4437_b1 , \5238_b1 );
not ( \5238_b1 , w_16712 );
and ( \5239_b0 , \4437_b0 , w_16713 );
and ( w_16712 , w_16713 , \5238_b0 );
buf ( \5240_b1 , \5005_b1 );
not ( \5240_b1 , w_16714 );
not ( \5240_b0 , w_16715 );
and ( w_16714 , w_16715 , \5005_b0 );
buf ( \5241_b1 , \4103_b1 );
buf ( \5241_b0 , \4103_b0 );
or ( \5242_b1 , \5240_b1 , w_16717 );
not ( w_16717 , w_16718 );
and ( \5242_b0 , \5240_b0 , w_16719 );
and ( w_16718 ,  , w_16719 );
buf ( w_16717 , \5241_b1 );
not ( w_16717 , w_16720 );
not (  , w_16721 );
and ( w_16720 , w_16721 , \5241_b0 );
or ( \5243_b1 , \5239_b1 , w_16723 );
not ( w_16723 , w_16724 );
and ( \5243_b0 , \5239_b0 , w_16725 );
and ( w_16724 ,  , w_16725 );
buf ( w_16723 , \5242_b1 );
not ( w_16723 , w_16726 );
not (  , w_16727 );
and ( w_16726 , w_16727 , \5242_b0 );
or ( \5244_b1 , \5232_b1 , \5243_b1 );
not ( \5243_b1 , w_16728 );
and ( \5244_b0 , \5232_b0 , w_16729 );
and ( w_16728 , w_16729 , \5243_b0 );
or ( \5245_b1 , \5220_b1 , \5231_b1 );
not ( \5231_b1 , w_16730 );
and ( \5245_b0 , \5220_b0 , w_16731 );
and ( w_16730 , w_16731 , \5231_b0 );
or ( \5246_b1 , \5244_b1 , w_16732 );
or ( \5246_b0 , \5244_b0 , \5245_b0 );
not ( \5245_b0 , w_16733 );
and ( w_16733 , w_16732 , \5245_b1 );
buf ( \5247_b1 , \5246_b1 );
not ( \5247_b1 , w_16734 );
not ( \5247_b0 , w_16735 );
and ( w_16734 , w_16735 , \5246_b0 );
buf ( \5248_b1 , \3963_b1 );
not ( \5248_b1 , w_16736 );
not ( \5248_b0 , w_16737 );
and ( w_16736 , w_16737 , \3963_b0 );
buf ( \5249_b1 , \4212_b1 );
not ( \5249_b1 , w_16738 );
not ( \5249_b0 , w_16739 );
and ( w_16738 , w_16739 , \4212_b0 );
or ( \5250_b1 , \5248_b1 , w_16740 );
or ( \5250_b0 , \5248_b0 , \5249_b0 );
not ( \5249_b0 , w_16741 );
and ( w_16741 , w_16740 , \5249_b1 );
or ( \5251_b1 , \4492_b1 , w_16743 );
not ( w_16743 , w_16744 );
and ( \5251_b0 , \4492_b0 , w_16745 );
and ( w_16744 ,  , w_16745 );
buf ( w_16743 , \4486_b1 );
not ( w_16743 , w_16746 );
not (  , w_16747 );
and ( w_16746 , w_16747 , \4486_b0 );
or ( \5252_b1 , \5250_b1 , w_16749 );
not ( w_16749 , w_16750 );
and ( \5252_b0 , \5250_b0 , w_16751 );
and ( w_16750 ,  , w_16751 );
buf ( w_16749 , \5251_b1 );
not ( w_16749 , w_16752 );
not (  , w_16753 );
and ( w_16752 , w_16753 , \5251_b0 );
buf ( \5253_b1 , \5252_b1 );
not ( \5253_b1 , w_16754 );
not ( \5253_b0 , w_16755 );
and ( w_16754 , w_16755 , \5252_b0 );
buf ( \5254_b1 , \4496_b1 );
not ( \5254_b1 , w_16756 );
not ( \5254_b0 , w_16757 );
and ( w_16756 , w_16757 , \4496_b0 );
or ( \5255_b1 , \5253_b1 , w_16758 );
or ( \5255_b0 , \5253_b0 , \5254_b0 );
not ( \5254_b0 , w_16759 );
and ( w_16759 , w_16758 , \5254_b1 );
or ( \5256_b1 , \4377_b1 , w_16761 );
not ( w_16761 , w_16762 );
and ( \5256_b0 , \4377_b0 , w_16763 );
and ( w_16762 ,  , w_16763 );
buf ( w_16761 , \5094_b1 );
not ( w_16761 , w_16764 );
not (  , w_16765 );
and ( w_16764 , w_16765 , \5094_b0 );
or ( \5257_b1 , \5255_b1 , w_16767 );
not ( w_16767 , w_16768 );
and ( \5257_b0 , \5255_b0 , w_16769 );
and ( w_16768 ,  , w_16769 );
buf ( w_16767 , \5256_b1 );
not ( w_16767 , w_16770 );
not (  , w_16771 );
and ( w_16770 , w_16771 , \5256_b0 );
or ( \5258_b1 , \5247_b1 , w_16773 );
not ( w_16773 , w_16774 );
and ( \5258_b0 , \5247_b0 , w_16775 );
and ( w_16774 ,  , w_16775 );
buf ( w_16773 , \5257_b1 );
not ( w_16773 , w_16776 );
not (  , w_16777 );
and ( w_16776 , w_16777 , \5257_b0 );
or ( \5259_b1 , \5208_b1 , \5258_b1 );
xor ( \5259_b0 , \5208_b0 , w_16778 );
not ( w_16778 , w_16779 );
and ( w_16779 , \5258_b1 , \5258_b0 );
or ( \5260_b1 , \5026_b1 , \5037_b1 );
xor ( \5260_b0 , \5026_b0 , w_16780 );
not ( w_16780 , w_16781 );
and ( w_16781 , \5037_b1 , \5037_b0 );
or ( \5261_b1 , \5260_b1 , \4676_b1 );
xor ( \5261_b0 , \5260_b0 , w_16782 );
not ( w_16782 , w_16783 );
and ( w_16783 , \4676_b1 , \4676_b0 );
or ( \5262_b1 , \5259_b1 , \5261_b1 );
not ( \5261_b1 , w_16784 );
and ( \5262_b0 , \5259_b0 , w_16785 );
and ( w_16784 , w_16785 , \5261_b0 );
or ( \5263_b1 , \5208_b1 , \5258_b1 );
not ( \5258_b1 , w_16786 );
and ( \5263_b0 , \5208_b0 , w_16787 );
and ( w_16786 , w_16787 , \5258_b0 );
or ( \5264_b1 , \5262_b1 , w_16788 );
or ( \5264_b0 , \5262_b0 , \5263_b0 );
not ( \5263_b0 , w_16789 );
and ( w_16789 , w_16788 , \5263_b1 );
buf ( \5265_b1 , \5021_b1 );
not ( \5265_b1 , w_16790 );
not ( \5265_b0 , w_16791 );
and ( w_16790 , w_16791 , \5021_b0 );
buf ( \5266_b1 , \5265_b1 );
not ( \5266_b1 , w_16792 );
not ( \5266_b0 , w_16793 );
and ( w_16792 , w_16793 , \5265_b0 );
buf ( \5267_b1 , \5023_b1 );
not ( \5267_b1 , w_16794 );
not ( \5267_b0 , w_16795 );
and ( w_16794 , w_16795 , \5023_b0 );
or ( \5268_b1 , \5266_b1 , \5267_b1 );
not ( \5267_b1 , w_16796 );
and ( \5268_b0 , \5266_b0 , w_16797 );
and ( w_16796 , w_16797 , \5267_b0 );
buf ( \5269_b1 , \3994_b1 );
not ( \5269_b1 , w_16798 );
not ( \5269_b0 , w_16799 );
and ( w_16798 , w_16799 , \3994_b0 );
buf ( \5270_b1 , \1395_b1 );
not ( \5270_b1 , w_16800 );
not ( \5270_b0 , w_16801 );
and ( w_16800 , w_16801 , \1395_b0 );
buf ( \5271_b1 , \5270_b1 );
not ( \5271_b1 , w_16802 );
not ( \5271_b0 , w_16803 );
and ( w_16802 , w_16803 , \5270_b0 );
or ( \5272_b1 , \5269_b1 , w_16804 );
or ( \5272_b0 , \5269_b0 , \5271_b0 );
not ( \5271_b0 , w_16805 );
and ( w_16805 , w_16804 , \5271_b1 );
buf ( \5273_b1 , \1395_b1 );
buf ( \5273_b0 , \1395_b0 );
or ( \5274_b1 , \5273_b1 , w_16807 );
not ( w_16807 , w_16808 );
and ( \5274_b0 , \5273_b0 , w_16809 );
and ( w_16808 ,  , w_16809 );
buf ( w_16807 , \4099_b1 );
not ( w_16807 , w_16810 );
not (  , w_16811 );
and ( w_16810 , w_16811 , \4099_b0 );
or ( \5275_b1 , \5272_b1 , w_16813 );
not ( w_16813 , w_16814 );
and ( \5275_b0 , \5272_b0 , w_16815 );
and ( w_16814 ,  , w_16815 );
buf ( w_16813 , \5274_b1 );
not ( w_16813 , w_16816 );
not (  , w_16817 );
and ( w_16816 , w_16817 , \5274_b0 );
or ( \5276_b1 , \5019_b1 , \5275_b1 );
not ( \5275_b1 , w_16818 );
and ( \5276_b0 , \5019_b0 , w_16819 );
and ( w_16818 , w_16819 , \5275_b0 );
or ( \5277_b1 , \5268_b1 , w_16821 );
not ( w_16821 , w_16822 );
and ( \5277_b0 , \5268_b0 , w_16823 );
and ( w_16822 ,  , w_16823 );
buf ( w_16821 , \5276_b1 );
not ( w_16821 , w_16824 );
not (  , w_16825 );
and ( w_16824 , w_16825 , \5276_b0 );
buf ( \5278_b1 , \5277_b1 );
not ( \5278_b1 , w_16826 );
not ( \5278_b0 , w_16827 );
and ( w_16826 , w_16827 , \5277_b0 );
buf ( \5279_b1 , \4019_b1 );
not ( \5279_b1 , w_16828 );
not ( \5279_b0 , w_16829 );
and ( w_16828 , w_16829 , \4019_b0 );
buf ( \5280_b1 , \4211_b1 );
not ( \5280_b1 , w_16830 );
not ( \5280_b0 , w_16831 );
and ( w_16830 , w_16831 , \4211_b0 );
or ( \5281_b1 , \5279_b1 , w_16832 );
or ( \5281_b0 , \5279_b0 , \5280_b0 );
not ( \5280_b0 , w_16833 );
and ( w_16833 , w_16832 , \5280_b1 );
or ( \5282_b1 , \4585_b1 , w_16835 );
not ( w_16835 , w_16836 );
and ( \5282_b0 , \4585_b0 , w_16837 );
and ( w_16836 ,  , w_16837 );
buf ( w_16835 , \3577_b1 );
not ( w_16835 , w_16838 );
not (  , w_16839 );
and ( w_16838 , w_16839 , \3577_b0 );
or ( \5283_b1 , \5281_b1 , w_16841 );
not ( w_16841 , w_16842 );
and ( \5283_b0 , \5281_b0 , w_16843 );
and ( w_16842 ,  , w_16843 );
buf ( w_16841 , \5282_b1 );
not ( w_16841 , w_16844 );
not (  , w_16845 );
and ( w_16844 , w_16845 , \5282_b0 );
buf ( \5284_b1 , \5283_b1 );
not ( \5284_b1 , w_16846 );
not ( \5284_b0 , w_16847 );
and ( w_16846 , w_16847 , \5283_b0 );
buf ( \5285_b1 , \4231_b1 );
not ( \5285_b1 , w_16848 );
not ( \5285_b0 , w_16849 );
and ( w_16848 , w_16849 , \4231_b0 );
or ( \5286_b1 , \5284_b1 , w_16850 );
or ( \5286_b0 , \5284_b0 , \5285_b0 );
not ( \5285_b0 , w_16851 );
and ( w_16851 , w_16850 , \5285_b1 );
or ( \5287_b1 , \4234_b1 , w_16853 );
not ( w_16853 , w_16854 );
and ( \5287_b0 , \4234_b0 , w_16855 );
and ( w_16854 ,  , w_16855 );
buf ( w_16853 , \5252_b1 );
not ( w_16853 , w_16856 );
not (  , w_16857 );
and ( w_16856 , w_16857 , \5252_b0 );
or ( \5288_b1 , \5286_b1 , w_16859 );
not ( w_16859 , w_16860 );
and ( \5288_b0 , \5286_b0 , w_16861 );
and ( w_16860 ,  , w_16861 );
buf ( w_16859 , \5287_b1 );
not ( w_16859 , w_16862 );
not (  , w_16863 );
and ( w_16862 , w_16863 , \5287_b0 );
buf ( \5289_b1 , \5288_b1 );
not ( \5289_b1 , w_16864 );
not ( \5289_b0 , w_16865 );
and ( w_16864 , w_16865 , \5288_b0 );
buf ( \5290_b1 , \5289_b1 );
not ( \5290_b1 , w_16866 );
not ( \5290_b0 , w_16867 );
and ( w_16866 , w_16867 , \5289_b0 );
or ( \5291_b1 , \5278_b1 , w_16868 );
or ( \5291_b0 , \5278_b0 , \5290_b0 );
not ( \5290_b0 , w_16869 );
and ( w_16869 , w_16868 , \5290_b1 );
buf ( \5292_b1 , \3958_b1 );
not ( \5292_b1 , w_16870 );
not ( \5292_b0 , w_16871 );
and ( w_16870 , w_16871 , \3958_b0 );
buf ( \5293_b1 , \4176_b1 );
not ( \5293_b1 , w_16872 );
not ( \5293_b0 , w_16873 );
and ( w_16872 , w_16873 , \4176_b0 );
or ( \5294_b1 , \5292_b1 , w_16874 );
or ( \5294_b0 , \5292_b0 , \5293_b0 );
not ( \5293_b0 , w_16875 );
and ( w_16875 , w_16874 , \5293_b1 );
or ( \5295_b1 , \4172_b1 , w_16877 );
not ( w_16877 , w_16878 );
and ( \5295_b0 , \4172_b0 , w_16879 );
and ( w_16878 ,  , w_16879 );
buf ( w_16877 , \4473_b1 );
not ( w_16877 , w_16880 );
not (  , w_16881 );
and ( w_16880 , w_16881 , \4473_b0 );
or ( \5296_b1 , \5294_b1 , w_16883 );
not ( w_16883 , w_16884 );
and ( \5296_b0 , \5294_b0 , w_16885 );
and ( w_16884 ,  , w_16885 );
buf ( w_16883 , \5295_b1 );
not ( w_16883 , w_16886 );
not (  , w_16887 );
and ( w_16886 , w_16887 , \5295_b0 );
buf ( \5297_b1 , \5296_b1 );
not ( \5297_b1 , w_16888 );
not ( \5297_b0 , w_16889 );
and ( w_16888 , w_16889 , \5296_b0 );
buf ( \5298_b1 , \4194_b1 );
not ( \5298_b1 , w_16890 );
not ( \5298_b0 , w_16891 );
and ( w_16890 , w_16891 , \4194_b0 );
or ( \5299_b1 , \5297_b1 , w_16892 );
or ( \5299_b0 , \5297_b0 , \5298_b0 );
not ( \5298_b0 , w_16893 );
and ( w_16893 , w_16892 , \5298_b1 );
or ( \5300_b1 , \5144_b1 , w_16895 );
not ( w_16895 , w_16896 );
and ( \5300_b0 , \5144_b0 , w_16897 );
and ( w_16896 ,  , w_16897 );
buf ( w_16895 , \4204_b1 );
not ( w_16895 , w_16898 );
not (  , w_16899 );
and ( w_16898 , w_16899 , \4204_b0 );
or ( \5301_b1 , \5299_b1 , w_16901 );
not ( w_16901 , w_16902 );
and ( \5301_b0 , \5299_b0 , w_16903 );
and ( w_16902 ,  , w_16903 );
buf ( w_16901 , \5300_b1 );
not ( w_16901 , w_16904 );
not (  , w_16905 );
and ( w_16904 , w_16905 , \5300_b0 );
or ( \5302_b1 , \5291_b1 , w_16907 );
not ( w_16907 , w_16908 );
and ( \5302_b0 , \5291_b0 , w_16909 );
and ( w_16908 ,  , w_16909 );
buf ( w_16907 , \5301_b1 );
not ( w_16907 , w_16910 );
not (  , w_16911 );
and ( w_16910 , w_16911 , \5301_b0 );
buf ( \5303_b1 , \5277_b1 );
not ( \5303_b1 , w_16912 );
not ( \5303_b0 , w_16913 );
and ( w_16912 , w_16913 , \5277_b0 );
or ( \5304_b1 , \5303_b1 , w_16915 );
not ( w_16915 , w_16916 );
and ( \5304_b0 , \5303_b0 , w_16917 );
and ( w_16916 ,  , w_16917 );
buf ( w_16915 , \5288_b1 );
not ( w_16915 , w_16918 );
not (  , w_16919 );
and ( w_16918 , w_16919 , \5288_b0 );
or ( \5305_b1 , \5302_b1 , w_16921 );
not ( w_16921 , w_16922 );
and ( \5305_b0 , \5302_b0 , w_16923 );
and ( w_16922 ,  , w_16923 );
buf ( w_16921 , \5304_b1 );
not ( w_16921 , w_16924 );
not (  , w_16925 );
and ( w_16924 , w_16925 , \5304_b0 );
buf ( \5306_b1 , \5305_b1 );
not ( \5306_b1 , w_16926 );
not ( \5306_b0 , w_16927 );
and ( w_16926 , w_16927 , \5305_b0 );
or ( \5307_b1 , \5138_b1 , \5149_b1 );
xor ( \5307_b0 , \5138_b0 , w_16928 );
not ( w_16928 , w_16929 );
and ( w_16929 , \5149_b1 , \5149_b0 );
or ( \5308_b1 , \5307_b1 , w_16930 );
xor ( \5308_b0 , \5307_b0 , w_16932 );
not ( w_16932 , w_16933 );
and ( w_16933 , w_16930 , w_16931 );
buf ( w_16930 , \5137_b1 );
not ( w_16930 , w_16934 );
not ( w_16931 , w_16935 );
and ( w_16934 , w_16935 , \5137_b0 );
or ( \5309_b1 , \5306_b1 , w_16937 );
not ( w_16937 , w_16938 );
and ( \5309_b0 , \5306_b0 , w_16939 );
and ( w_16938 ,  , w_16939 );
buf ( w_16937 , \5308_b1 );
not ( w_16937 , w_16940 );
not (  , w_16941 );
and ( w_16940 , w_16941 , \5308_b0 );
buf ( \5310_b1 , \5257_b1 );
not ( \5310_b1 , w_16942 );
not ( \5310_b0 , w_16943 );
and ( w_16942 , w_16943 , \5257_b0 );
buf ( \5311_b1 , \5246_b1 );
not ( \5311_b1 , w_16944 );
not ( \5311_b0 , w_16945 );
and ( w_16944 , w_16945 , \5246_b0 );
or ( \5312_b1 , \5310_b1 , w_16946 );
or ( \5312_b0 , \5310_b0 , \5311_b0 );
not ( \5311_b0 , w_16947 );
and ( w_16947 , w_16946 , \5311_b1 );
or ( \5313_b1 , \5246_b1 , w_16948 );
or ( \5313_b0 , \5246_b0 , \5257_b0 );
not ( \5257_b0 , w_16949 );
and ( w_16949 , w_16948 , \5257_b1 );
or ( \5314_b1 , \5312_b1 , w_16951 );
not ( w_16951 , w_16952 );
and ( \5314_b0 , \5312_b0 , w_16953 );
and ( w_16952 ,  , w_16953 );
buf ( w_16951 , \5313_b1 );
not ( w_16951 , w_16954 );
not (  , w_16955 );
and ( w_16954 , w_16955 , \5313_b0 );
or ( \5315_b1 , \5309_b1 , \5314_b1 );
not ( \5314_b1 , w_16956 );
and ( \5315_b0 , \5309_b0 , w_16957 );
and ( w_16956 , w_16957 , \5314_b0 );
or ( \5316_b1 , \5306_b1 , w_16959 );
not ( w_16959 , w_16960 );
and ( \5316_b0 , \5306_b0 , w_16961 );
and ( w_16960 ,  , w_16961 );
buf ( w_16959 , \5308_b1 );
not ( w_16959 , w_16962 );
not (  , w_16963 );
and ( w_16962 , w_16963 , \5308_b0 );
or ( \5317_b1 , \5315_b1 , w_16965 );
not ( w_16965 , w_16966 );
and ( \5317_b0 , \5315_b0 , w_16967 );
and ( w_16966 ,  , w_16967 );
buf ( w_16965 , \5316_b1 );
not ( w_16965 , w_16968 );
not (  , w_16969 );
and ( w_16968 , w_16969 , \5316_b0 );
buf ( \5318_b1 , \5317_b1 );
not ( \5318_b1 , w_16970 );
not ( \5318_b0 , w_16971 );
and ( w_16970 , w_16971 , \5317_b0 );
or ( \5319_b1 , \5152_b1 , \5191_b1 );
xor ( \5319_b0 , \5152_b0 , w_16972 );
not ( w_16972 , w_16973 );
and ( w_16973 , \5191_b1 , \5191_b0 );
or ( \5320_b1 , \5319_b1 , \5194_b1 );
not ( \5194_b1 , w_16974 );
and ( \5320_b0 , \5319_b0 , w_16975 );
and ( w_16974 , w_16975 , \5194_b0 );
buf ( \5321_b1 , \5319_b1 );
not ( \5321_b1 , w_16976 );
not ( \5321_b0 , w_16977 );
and ( w_16976 , w_16977 , \5319_b0 );
buf ( \5322_b1 , \5194_b1 );
not ( \5322_b1 , w_16978 );
not ( \5322_b0 , w_16979 );
and ( w_16978 , w_16979 , \5194_b0 );
or ( \5323_b1 , \5321_b1 , \5322_b1 );
not ( \5322_b1 , w_16980 );
and ( \5323_b0 , \5321_b0 , w_16981 );
and ( w_16980 , w_16981 , \5322_b0 );
or ( \5324_b1 , \5320_b1 , w_16983 );
not ( w_16983 , w_16984 );
and ( \5324_b0 , \5320_b0 , w_16985 );
and ( w_16984 ,  , w_16985 );
buf ( w_16983 , \5323_b1 );
not ( w_16983 , w_16986 );
not (  , w_16987 );
and ( w_16986 , w_16987 , \5323_b0 );
buf ( \5325_b1 , \5324_b1 );
not ( \5325_b1 , w_16988 );
not ( \5325_b0 , w_16989 );
and ( w_16988 , w_16989 , \5324_b0 );
buf ( \5326_b1 , \5325_b1 );
not ( \5326_b1 , w_16990 );
not ( \5326_b0 , w_16991 );
and ( w_16990 , w_16991 , \5325_b0 );
or ( \5327_b1 , \5318_b1 , w_16992 );
or ( \5327_b0 , \5318_b0 , \5326_b0 );
not ( \5326_b0 , w_16993 );
and ( w_16993 , w_16992 , \5326_b1 );
buf ( \5328_b1 , \5026_b1 );
not ( \5328_b1 , w_16994 );
not ( \5328_b0 , w_16995 );
and ( w_16994 , w_16995 , \5026_b0 );
or ( \5329_b1 , \5015_b1 , w_16997 );
not ( w_16997 , w_16998 );
and ( \5329_b0 , \5015_b0 , w_16999 );
and ( w_16998 ,  , w_16999 );
buf ( w_16997 , \5025_b1 );
not ( w_16997 , w_17000 );
not (  , w_17001 );
and ( w_17000 , w_17001 , \5025_b0 );
or ( \5330_b1 , \5328_b1 , w_17003 );
not ( w_17003 , w_17004 );
and ( \5330_b0 , \5328_b0 , w_17005 );
and ( w_17004 ,  , w_17005 );
buf ( w_17003 , \5329_b1 );
not ( w_17003 , w_17006 );
not (  , w_17007 );
and ( w_17006 , w_17007 , \5329_b0 );
buf ( \5331_b1 , \5330_b1 );
not ( \5331_b1 , w_17008 );
not ( \5331_b0 , w_17009 );
and ( w_17008 , w_17009 , \5330_b0 );
or ( \5332_b1 , \5162_b1 , \5189_b1 );
xor ( \5332_b0 , \5162_b0 , w_17010 );
not ( w_17010 , w_17011 );
and ( w_17011 , \5189_b1 , \5189_b0 );
buf ( \5333_b1 , \5173_b1 );
not ( \5333_b1 , w_17012 );
not ( \5333_b0 , w_17013 );
and ( w_17012 , w_17013 , \5173_b0 );
or ( \5334_b1 , \5332_b1 , \5333_b1 );
not ( \5333_b1 , w_17014 );
and ( \5334_b0 , \5332_b0 , w_17015 );
and ( w_17014 , w_17015 , \5333_b0 );
buf ( \5335_b1 , \5332_b1 );
not ( \5335_b1 , w_17016 );
not ( \5335_b0 , w_17017 );
and ( w_17016 , w_17017 , \5332_b0 );
or ( \5336_b1 , \5335_b1 , \5173_b1 );
not ( \5173_b1 , w_17018 );
and ( \5336_b0 , \5335_b0 , w_17019 );
and ( w_17018 , w_17019 , \5173_b0 );
or ( \5337_b1 , \5334_b1 , w_17021 );
not ( w_17021 , w_17022 );
and ( \5337_b0 , \5334_b0 , w_17023 );
and ( w_17022 ,  , w_17023 );
buf ( w_17021 , \5336_b1 );
not ( w_17021 , w_17024 );
not (  , w_17025 );
and ( w_17024 , w_17025 , \5336_b0 );
or ( \5338_b1 , \5331_b1 , w_17027 );
not ( w_17027 , w_17028 );
and ( \5338_b0 , \5331_b0 , w_17029 );
and ( w_17028 ,  , w_17029 );
buf ( w_17027 , \5337_b1 );
not ( w_17027 , w_17030 );
not (  , w_17031 );
and ( w_17030 , w_17031 , \5337_b0 );
buf ( \5339_b1 , \4029_b1 );
not ( \5339_b1 , w_17032 );
not ( \5339_b0 , w_17033 );
and ( w_17032 , w_17033 , \4029_b0 );
or ( \5340_b1 , \4267_b1 , w_17035 );
not ( w_17035 , w_17036 );
and ( \5340_b0 , \4267_b0 , w_17037 );
and ( w_17036 ,  , w_17037 );
buf ( w_17035 , \5339_b1 );
not ( w_17035 , w_17038 );
not (  , w_17039 );
and ( w_17038 , w_17039 , \5339_b0 );
or ( \5341_b1 , \4260_b1 , \4026_b1 );
not ( \4026_b1 , w_17040 );
and ( \5341_b0 , \4260_b0 , w_17041 );
and ( w_17040 , w_17041 , \4026_b0 );
buf ( \5342_b1 , \3108_b1 );
not ( \5342_b1 , w_17042 );
not ( \5342_b0 , w_17043 );
and ( w_17042 , w_17043 , \3108_b0 );
buf ( \5343_b1 , \5342_b1 );
not ( \5343_b1 , w_17044 );
not ( \5343_b0 , w_17045 );
and ( w_17044 , w_17045 , \5342_b0 );
buf ( \5344_b1 , \4026_b1 );
not ( \5344_b1 , w_17046 );
not ( \5344_b0 , w_17047 );
and ( w_17046 , w_17047 , \4026_b0 );
or ( \5345_b1 , \5343_b1 , \5344_b1 );
not ( \5344_b1 , w_17048 );
and ( \5345_b0 , \5343_b0 , w_17049 );
and ( w_17048 , w_17049 , \5344_b0 );
or ( \5346_b1 , \5341_b1 , w_17051 );
not ( w_17051 , w_17052 );
and ( \5346_b0 , \5341_b0 , w_17053 );
and ( w_17052 ,  , w_17053 );
buf ( w_17051 , \5345_b1 );
not ( w_17051 , w_17054 );
not (  , w_17055 );
and ( w_17054 , w_17055 , \5345_b0 );
buf ( \5347_b1 , \5346_b1 );
not ( \5347_b1 , w_17056 );
not ( \5347_b0 , w_17057 );
and ( w_17056 , w_17057 , \5346_b0 );
buf ( \5348_b1 , \5347_b1 );
not ( \5348_b1 , w_17058 );
not ( \5348_b0 , w_17059 );
and ( w_17058 , w_17059 , \5347_b0 );
buf ( \5349_b1 , \4480_b1 );
not ( \5349_b1 , w_17060 );
not ( \5349_b0 , w_17061 );
and ( w_17060 , w_17061 , \4480_b0 );
or ( \5350_b1 , \5348_b1 , w_17062 );
or ( \5350_b0 , \5348_b0 , \5349_b0 );
not ( \5349_b0 , w_17063 );
and ( w_17063 , w_17062 , \5349_b1 );
or ( \5351_b1 , \5133_b1 , w_17065 );
not ( w_17065 , w_17066 );
and ( \5351_b0 , \5133_b0 , w_17067 );
and ( w_17066 ,  , w_17067 );
buf ( w_17065 , \4273_b1 );
not ( w_17065 , w_17068 );
not (  , w_17069 );
and ( w_17068 , w_17069 , \4273_b0 );
or ( \5352_b1 , \5350_b1 , w_17071 );
not ( w_17071 , w_17072 );
and ( \5352_b0 , \5350_b0 , w_17073 );
and ( w_17072 ,  , w_17073 );
buf ( w_17071 , \5351_b1 );
not ( w_17071 , w_17074 );
not (  , w_17075 );
and ( w_17074 , w_17075 , \5351_b0 );
or ( \5353_b1 , \5340_b1 , \5352_b1 );
xor ( \5353_b0 , \5340_b0 , w_17076 );
not ( w_17076 , w_17077 );
and ( w_17077 , \5352_b1 , \5352_b0 );
buf ( \5354_b1 , \4047_b1 );
not ( \5354_b1 , w_17078 );
not ( \5354_b0 , w_17079 );
and ( w_17078 , w_17079 , \4047_b0 );
buf ( \5355_b1 , \4404_b1 );
not ( \5355_b1 , w_17080 );
not ( \5355_b0 , w_17081 );
and ( w_17080 , w_17081 , \4404_b0 );
or ( \5356_b1 , \5354_b1 , w_17082 );
or ( \5356_b0 , \5354_b0 , \5355_b0 );
not ( \5355_b0 , w_17083 );
and ( w_17083 , w_17082 , \5355_b1 );
buf ( \5357_b1 , \4061_b1 );
not ( \5357_b1 , w_17084 );
not ( \5357_b0 , w_17085 );
and ( w_17084 , w_17085 , \4061_b0 );
or ( \5358_b1 , \5357_b1 , w_17087 );
not ( w_17087 , w_17088 );
and ( \5358_b0 , \5357_b0 , w_17089 );
and ( w_17088 ,  , w_17089 );
buf ( w_17087 , \4178_b1 );
not ( w_17087 , w_17090 );
not (  , w_17091 );
and ( w_17090 , w_17091 , \4178_b0 );
or ( \5359_b1 , \5356_b1 , w_17093 );
not ( w_17093 , w_17094 );
and ( \5359_b0 , \5356_b0 , w_17095 );
and ( w_17094 ,  , w_17095 );
buf ( w_17093 , \5358_b1 );
not ( w_17093 , w_17096 );
not (  , w_17097 );
and ( w_17096 , w_17097 , \5358_b0 );
buf ( \5360_b1 , \5359_b1 );
not ( \5360_b1 , w_17098 );
not ( \5360_b0 , w_17099 );
and ( w_17098 , w_17099 , \5359_b0 );
buf ( \5361_b1 , \4066_b1 );
not ( \5361_b1 , w_17100 );
not ( \5361_b0 , w_17101 );
and ( w_17100 , w_17101 , \4066_b0 );
buf ( \5362_b1 , \5361_b1 );
not ( \5362_b1 , w_17102 );
not ( \5362_b0 , w_17103 );
and ( w_17102 , w_17103 , \5361_b0 );
or ( \5363_b1 , \5360_b1 , w_17104 );
or ( \5363_b0 , \5360_b0 , \5362_b0 );
not ( \5362_b0 , w_17105 );
and ( w_17105 , w_17104 , \5362_b1 );
or ( \5364_b1 , \4562_b1 , w_17107 );
not ( w_17107 , w_17108 );
and ( \5364_b0 , \4562_b0 , w_17109 );
and ( w_17108 ,  , w_17109 );
buf ( w_17107 , \5157_b1 );
not ( w_17107 , w_17110 );
not (  , w_17111 );
and ( w_17110 , w_17111 , \5157_b0 );
or ( \5365_b1 , \5363_b1 , w_17113 );
not ( w_17113 , w_17114 );
and ( \5365_b0 , \5363_b0 , w_17115 );
and ( w_17114 ,  , w_17115 );
buf ( w_17113 , \5364_b1 );
not ( w_17113 , w_17116 );
not (  , w_17117 );
and ( w_17116 , w_17117 , \5364_b0 );
or ( \5366_b1 , \5353_b1 , \5365_b1 );
not ( \5365_b1 , w_17118 );
and ( \5366_b0 , \5353_b0 , w_17119 );
and ( w_17118 , w_17119 , \5365_b0 );
or ( \5367_b1 , \5340_b1 , \5352_b1 );
not ( \5352_b1 , w_17120 );
and ( \5367_b0 , \5340_b0 , w_17121 );
and ( w_17120 , w_17121 , \5352_b0 );
or ( \5368_b1 , \5366_b1 , w_17122 );
or ( \5368_b0 , \5366_b0 , \5367_b0 );
not ( \5367_b0 , w_17123 );
and ( w_17123 , w_17122 , \5367_b1 );
or ( \5369_b1 , \5338_b1 , \5368_b1 );
not ( \5368_b1 , w_17124 );
and ( \5369_b0 , \5338_b0 , w_17125 );
and ( w_17124 , w_17125 , \5368_b0 );
buf ( \5370_b1 , \5330_b1 );
not ( \5370_b1 , w_17126 );
not ( \5370_b0 , w_17127 );
and ( w_17126 , w_17127 , \5330_b0 );
or ( \5371_b1 , \5370_b1 , w_17129 );
not ( w_17129 , w_17130 );
and ( \5371_b0 , \5370_b0 , w_17131 );
and ( w_17130 ,  , w_17131 );
buf ( w_17129 , \5337_b1 );
not ( w_17129 , w_17132 );
not (  , w_17133 );
and ( w_17132 , w_17133 , \5337_b0 );
or ( \5372_b1 , \5369_b1 , w_17135 );
not ( w_17135 , w_17136 );
and ( \5372_b0 , \5369_b0 , w_17137 );
and ( w_17136 ,  , w_17137 );
buf ( w_17135 , \5371_b1 );
not ( w_17135 , w_17138 );
not (  , w_17139 );
and ( w_17138 , w_17139 , \5371_b0 );
buf ( \5373_b1 , \5372_b1 );
not ( \5373_b1 , w_17140 );
not ( \5373_b0 , w_17141 );
and ( w_17140 , w_17141 , \5372_b0 );
or ( \5374_b1 , \5327_b1 , w_17143 );
not ( w_17143 , w_17144 );
and ( \5374_b0 , \5327_b0 , w_17145 );
and ( w_17144 ,  , w_17145 );
buf ( w_17143 , \5373_b1 );
not ( w_17143 , w_17146 );
not (  , w_17147 );
and ( w_17146 , w_17147 , \5373_b0 );
or ( \5375_b1 , \5325_b1 , w_17148 );
or ( \5375_b0 , \5325_b0 , \5317_b0 );
not ( \5317_b0 , w_17149 );
and ( w_17149 , w_17148 , \5317_b1 );
or ( \5376_b1 , \5374_b1 , \5375_b1 );
not ( \5375_b1 , w_17150 );
and ( \5376_b0 , \5374_b0 , w_17151 );
and ( w_17150 , w_17151 , \5375_b0 );
or ( \5377_b1 , \5264_b1 , \5376_b1 );
xor ( \5377_b0 , \5264_b0 , w_17152 );
not ( w_17152 , w_17153 );
and ( w_17153 , \5376_b1 , \5376_b0 );
or ( \5378_b1 , \5197_b1 , \5199_b1 );
xor ( \5378_b0 , \5197_b0 , w_17154 );
not ( w_17154 , w_17155 );
and ( w_17155 , \5199_b1 , \5199_b0 );
or ( \5379_b1 , \5378_b1 , \5202_b1 );
xor ( \5379_b0 , \5378_b0 , w_17156 );
not ( w_17156 , w_17157 );
and ( w_17157 , \5202_b1 , \5202_b0 );
or ( \5380_b1 , \5377_b1 , \5379_b1 );
not ( \5379_b1 , w_17158 );
and ( \5380_b0 , \5377_b0 , w_17159 );
and ( w_17158 , w_17159 , \5379_b0 );
or ( \5381_b1 , \5264_b1 , \5376_b1 );
not ( \5376_b1 , w_17160 );
and ( \5381_b0 , \5264_b0 , w_17161 );
and ( w_17160 , w_17161 , \5376_b0 );
or ( \5382_b1 , \5380_b1 , w_17162 );
or ( \5382_b0 , \5380_b0 , \5381_b0 );
not ( \5381_b0 , w_17163 );
and ( w_17163 , w_17162 , \5381_b1 );
or ( \5383_b1 , \5206_b1 , w_17165 );
not ( w_17165 , w_17166 );
and ( \5383_b0 , \5206_b0 , w_17167 );
and ( w_17166 ,  , w_17167 );
buf ( w_17165 , \5382_b1 );
not ( w_17165 , w_17168 );
not (  , w_17169 );
and ( w_17168 , w_17169 , \5382_b0 );
or ( \5384_b1 , \5264_b1 , \5376_b1 );
xor ( \5384_b0 , \5264_b0 , w_17170 );
not ( w_17170 , w_17171 );
and ( w_17171 , \5376_b1 , \5376_b0 );
or ( \5385_b1 , \5384_b1 , \5379_b1 );
xor ( \5385_b0 , \5384_b0 , w_17172 );
not ( w_17172 , w_17173 );
and ( w_17173 , \5379_b1 , \5379_b0 );
or ( \5386_b1 , \5208_b1 , \5258_b1 );
xor ( \5386_b0 , \5208_b0 , w_17174 );
not ( w_17174 , w_17175 );
and ( w_17175 , \5258_b1 , \5258_b0 );
or ( \5387_b1 , \5386_b1 , \5261_b1 );
xor ( \5387_b0 , \5386_b0 , w_17176 );
not ( w_17176 , w_17177 );
and ( w_17177 , \5261_b1 , \5261_b0 );
buf ( \5388_b1 , \4048_b1 );
not ( \5388_b1 , w_17178 );
not ( \5388_b0 , w_17179 );
and ( w_17178 , w_17179 , \4048_b0 );
or ( \5389_b1 , \5342_b1 , w_17181 );
not ( w_17181 , w_17182 );
and ( \5389_b0 , \5342_b0 , w_17183 );
and ( w_17182 ,  , w_17183 );
buf ( w_17181 , \5388_b1 );
not ( w_17181 , w_17184 );
not (  , w_17185 );
and ( w_17184 , w_17185 , \5388_b0 );
or ( \5390_b1 , \3617_b1 , w_17187 );
not ( w_17187 , w_17188 );
and ( \5390_b0 , \3617_b0 , w_17189 );
and ( w_17188 ,  , w_17189 );
buf ( w_17187 , \5270_b1 );
not ( w_17187 , w_17190 );
not (  , w_17191 );
and ( w_17190 , w_17191 , \5270_b0 );
buf ( \5391_b1 , \5390_b1 );
not ( \5391_b1 , w_17192 );
not ( \5391_b0 , w_17193 );
and ( w_17192 , w_17193 , \5390_b0 );
buf ( \5392_b1 , \4044_b1 );
not ( \5392_b1 , w_17194 );
not ( \5392_b0 , w_17195 );
and ( w_17194 , w_17195 , \4044_b0 );
buf ( \5393_b1 , \5270_b1 );
not ( \5393_b1 , w_17196 );
not ( \5393_b0 , w_17197 );
and ( w_17196 , w_17197 , \5270_b0 );
or ( \5394_b1 , \5392_b1 , w_17198 );
or ( \5394_b0 , \5392_b0 , \5393_b0 );
not ( \5393_b0 , w_17199 );
and ( w_17199 , w_17198 , \5393_b1 );
or ( \5395_b1 , \5273_b1 , w_17201 );
not ( w_17201 , w_17202 );
and ( \5395_b0 , \5273_b0 , w_17203 );
and ( w_17202 ,  , w_17203 );
buf ( w_17201 , \4092_b1 );
not ( w_17201 , w_17204 );
not (  , w_17205 );
and ( w_17204 , w_17205 , \4092_b0 );
or ( \5396_b1 , \5394_b1 , w_17207 );
not ( w_17207 , w_17208 );
and ( \5396_b0 , \5394_b0 , w_17209 );
and ( w_17208 ,  , w_17209 );
buf ( w_17207 , \5395_b1 );
not ( w_17207 , w_17210 );
not (  , w_17211 );
and ( w_17210 , w_17211 , \5395_b0 );
buf ( \5397_b1 , \5396_b1 );
not ( \5397_b1 , w_17212 );
not ( \5397_b0 , w_17213 );
and ( w_17212 , w_17213 , \5396_b0 );
or ( \5398_b1 , \5391_b1 , w_17214 );
or ( \5398_b0 , \5391_b0 , \5397_b0 );
not ( \5397_b0 , w_17215 );
and ( w_17215 , w_17214 , \5397_b1 );
or ( \5399_b1 , \5275_b1 , w_17217 );
not ( w_17217 , w_17218 );
and ( \5399_b0 , \5275_b0 , w_17219 );
and ( w_17218 ,  , w_17219 );
buf ( w_17217 , \5021_b1 );
not ( w_17217 , w_17220 );
not (  , w_17221 );
and ( w_17220 , w_17221 , \5021_b0 );
or ( \5400_b1 , \5398_b1 , w_17223 );
not ( w_17223 , w_17224 );
and ( \5400_b0 , \5398_b0 , w_17225 );
and ( w_17224 ,  , w_17225 );
buf ( w_17223 , \5399_b1 );
not ( w_17223 , w_17226 );
not (  , w_17227 );
and ( w_17226 , w_17227 , \5399_b0 );
or ( \5401_b1 , \5389_b1 , \5400_b1 );
xor ( \5401_b0 , \5389_b0 , w_17228 );
not ( w_17228 , w_17229 );
and ( w_17229 , \5400_b1 , \5400_b0 );
buf ( \5402_b1 , \4042_b1 );
not ( \5402_b1 , w_17230 );
not ( \5402_b0 , w_17231 );
and ( w_17230 , w_17231 , \4042_b0 );
buf ( \5403_b1 , \5178_b1 );
not ( \5403_b1 , w_17232 );
not ( \5403_b0 , w_17233 );
and ( w_17232 , w_17233 , \5178_b0 );
or ( \5404_b1 , \5402_b1 , w_17234 );
or ( \5404_b0 , \5402_b0 , \5403_b0 );
not ( \5403_b0 , w_17235 );
and ( w_17235 , w_17234 , \5403_b1 );
or ( \5405_b1 , \4665_b1 , w_17237 );
not ( w_17237 , w_17238 );
and ( \5405_b0 , \4665_b0 , w_17239 );
and ( w_17238 ,  , w_17239 );
buf ( w_17237 , \4116_b1 );
not ( w_17237 , w_17240 );
not (  , w_17241 );
and ( w_17240 , w_17241 , \4116_b0 );
or ( \5406_b1 , \5404_b1 , w_17243 );
not ( w_17243 , w_17244 );
and ( \5406_b0 , \5404_b0 , w_17245 );
and ( w_17244 ,  , w_17245 );
buf ( w_17243 , \5405_b1 );
not ( w_17243 , w_17246 );
not (  , w_17247 );
and ( w_17246 , w_17247 , \5405_b0 );
buf ( \5407_b1 , \5406_b1 );
not ( \5407_b1 , w_17248 );
not ( \5407_b0 , w_17249 );
and ( w_17248 , w_17249 , \5406_b0 );
buf ( \5408_b1 , \4661_b1 );
not ( \5408_b1 , w_17250 );
not ( \5408_b0 , w_17251 );
and ( w_17250 , w_17251 , \4661_b0 );
or ( \5409_b1 , \5407_b1 , w_17252 );
or ( \5409_b0 , \5407_b0 , \5408_b0 );
not ( \5408_b0 , w_17253 );
and ( w_17253 , w_17252 , \5408_b1 );
or ( \5410_b1 , \5225_b1 , w_17255 );
not ( w_17255 , w_17256 );
and ( \5410_b0 , \5225_b0 , w_17257 );
and ( w_17256 ,  , w_17257 );
buf ( w_17255 , \5187_b1 );
not ( w_17255 , w_17258 );
not (  , w_17259 );
and ( w_17258 , w_17259 , \5187_b0 );
or ( \5411_b1 , \5409_b1 , w_17261 );
not ( w_17261 , w_17262 );
and ( \5411_b0 , \5409_b0 , w_17263 );
and ( w_17262 ,  , w_17263 );
buf ( w_17261 , \5410_b1 );
not ( w_17261 , w_17264 );
not (  , w_17265 );
and ( w_17264 , w_17265 , \5410_b0 );
or ( \5412_b1 , \5401_b1 , \5411_b1 );
not ( \5411_b1 , w_17266 );
and ( \5412_b0 , \5401_b0 , w_17267 );
and ( w_17266 , w_17267 , \5411_b0 );
or ( \5413_b1 , \5389_b1 , \5400_b1 );
not ( \5400_b1 , w_17268 );
and ( \5413_b0 , \5389_b0 , w_17269 );
and ( w_17268 , w_17269 , \5400_b0 );
or ( \5414_b1 , \5412_b1 , w_17270 );
or ( \5414_b0 , \5412_b0 , \5413_b0 );
not ( \5413_b0 , w_17271 );
and ( w_17271 , w_17270 , \5413_b1 );
buf ( \5415_b1 , \4054_b1 );
not ( \5415_b1 , w_17272 );
not ( \5415_b0 , w_17273 );
and ( w_17272 , w_17273 , \4054_b0 );
buf ( \5416_b1 , \5359_b1 );
not ( \5416_b1 , w_17274 );
not ( \5416_b0 , w_17275 );
and ( w_17274 , w_17275 , \5359_b0 );
or ( \5417_b1 , \5415_b1 , w_17276 );
or ( \5417_b0 , \5415_b0 , \5416_b0 );
not ( \5416_b0 , w_17277 );
and ( w_17277 , w_17276 , \5416_b1 );
or ( \5418_b1 , \4045_b1 , \4403_b1 );
not ( \4403_b1 , w_17278 );
and ( \5418_b0 , \4045_b0 , w_17279 );
and ( w_17278 , w_17279 , \4403_b0 );
buf ( \5419_b1 , \4045_b1 );
not ( \5419_b1 , w_17280 );
not ( \5419_b0 , w_17281 );
and ( w_17280 , w_17281 , \4045_b0 );
buf ( \5420_b1 , \5357_b1 );
not ( \5420_b1 , w_17282 );
not ( \5420_b0 , w_17283 );
and ( w_17282 , w_17283 , \5357_b0 );
or ( \5421_b1 , \5419_b1 , \5420_b1 );
not ( \5420_b1 , w_17284 );
and ( \5421_b0 , \5419_b0 , w_17285 );
and ( w_17284 , w_17285 , \5420_b0 );
or ( \5422_b1 , \5418_b1 , w_17287 );
not ( w_17287 , w_17288 );
and ( \5422_b0 , \5418_b0 , w_17289 );
and ( w_17288 ,  , w_17289 );
buf ( w_17287 , \5421_b1 );
not ( w_17287 , w_17290 );
not (  , w_17291 );
and ( w_17290 , w_17291 , \5421_b0 );
or ( \5424_b1 , \5417_b1 , w_17293 );
not ( w_17293 , w_17294 );
and ( \5424_b0 , \5417_b0 , w_17295 );
and ( w_17294 ,  , w_17295 );
buf ( w_17293 , \5423_b1 );
not ( w_17293 , w_17296 );
not (  , w_17297 );
and ( w_17296 , w_17297 , \5423_b0 );
buf ( \5425_b1 , \4046_b1 );
not ( \5425_b1 , w_17298 );
not ( \5425_b0 , w_17299 );
and ( w_17298 , w_17299 , \4046_b0 );
buf ( \5426_b1 , \4145_b1 );
not ( \5426_b1 , w_17300 );
not ( \5426_b0 , w_17301 );
and ( w_17300 , w_17301 , \4145_b0 );
or ( \5427_b1 , \5425_b1 , w_17302 );
or ( \5427_b0 , \5425_b0 , \5426_b0 );
not ( \5426_b0 , w_17303 );
and ( w_17303 , w_17302 , \5426_b1 );
or ( \5428_b1 , \4109_b1 , w_17305 );
not ( w_17305 , w_17306 );
and ( \5428_b0 , \4109_b0 , w_17307 );
and ( w_17306 ,  , w_17307 );
buf ( w_17305 , \4256_b1 );
not ( w_17305 , w_17308 );
not (  , w_17309 );
and ( w_17308 , w_17309 , \4256_b0 );
or ( \5429_b1 , \5427_b1 , w_17311 );
not ( w_17311 , w_17312 );
and ( \5429_b0 , \5427_b0 , w_17313 );
and ( w_17312 ,  , w_17313 );
buf ( w_17311 , \5428_b1 );
not ( w_17311 , w_17314 );
not (  , w_17315 );
and ( w_17314 , w_17315 , \5428_b0 );
buf ( \5430_b1 , \5429_b1 );
not ( \5430_b1 , w_17316 );
not ( \5430_b0 , w_17317 );
and ( w_17316 , w_17317 , \5429_b0 );
buf ( \5431_b1 , \5209_b1 );
not ( \5431_b1 , w_17318 );
not ( \5431_b0 , w_17319 );
and ( w_17318 , w_17319 , \5209_b0 );
buf ( \5432_b1 , \5431_b1 );
not ( \5432_b1 , w_17320 );
not ( \5432_b0 , w_17321 );
and ( w_17320 , w_17321 , \5431_b0 );
or ( \5433_b1 , \5430_b1 , w_17322 );
or ( \5433_b0 , \5430_b0 , \5432_b0 );
not ( \5432_b0 , w_17323 );
and ( w_17323 , w_17322 , \5432_b1 );
or ( \5434_b1 , \4139_b1 , w_17325 );
not ( w_17325 , w_17326 );
and ( \5434_b0 , \4139_b0 , w_17327 );
and ( w_17326 ,  , w_17327 );
buf ( w_17325 , \5215_b1 );
not ( w_17325 , w_17328 );
not (  , w_17329 );
and ( w_17328 , w_17329 , \5215_b0 );
or ( \5435_b1 , \5433_b1 , w_17331 );
not ( w_17331 , w_17332 );
and ( \5435_b0 , \5433_b0 , w_17333 );
and ( w_17332 ,  , w_17333 );
buf ( w_17331 , \5434_b1 );
not ( w_17331 , w_17334 );
not (  , w_17335 );
and ( w_17334 , w_17335 , \5434_b0 );
or ( \5436_b1 , \5424_b1 , \5435_b1 );
xor ( \5436_b0 , \5424_b0 , w_17336 );
not ( w_17336 , w_17337 );
and ( w_17337 , \5435_b1 , \5435_b0 );
buf ( \5437_b1 , \4043_b1 );
not ( \5437_b1 , w_17338 );
not ( \5437_b0 , w_17339 );
and ( w_17338 , w_17339 , \4043_b0 );
buf ( \5438_b1 , \4089_b1 );
not ( \5438_b1 , w_17340 );
not ( \5438_b0 , w_17341 );
and ( w_17340 , w_17341 , \4089_b0 );
or ( \5439_b1 , \5437_b1 , w_17342 );
or ( \5439_b0 , \5437_b0 , \5438_b0 );
not ( \5438_b0 , w_17343 );
and ( w_17343 , w_17342 , \5438_b1 );
or ( \5440_b1 , \4088_b1 , w_17345 );
not ( w_17345 , w_17346 );
and ( \5440_b0 , \4088_b0 , w_17347 );
and ( w_17346 ,  , w_17347 );
buf ( w_17345 , \4217_b1 );
not ( w_17345 , w_17348 );
not (  , w_17349 );
and ( w_17348 , w_17349 , \4217_b0 );
or ( \5441_b1 , \5439_b1 , w_17351 );
not ( w_17351 , w_17352 );
and ( \5441_b0 , \5439_b0 , w_17353 );
and ( w_17352 ,  , w_17353 );
buf ( w_17351 , \5440_b1 );
not ( w_17351 , w_17354 );
not (  , w_17355 );
and ( w_17354 , w_17355 , \5440_b0 );
buf ( \5442_b1 , \5441_b1 );
not ( \5442_b1 , w_17356 );
not ( \5442_b0 , w_17357 );
and ( w_17356 , w_17357 , \5441_b0 );
buf ( \5443_b1 , \4085_b1 );
not ( \5443_b1 , w_17358 );
not ( \5443_b0 , w_17359 );
and ( w_17358 , w_17359 , \4085_b0 );
or ( \5444_b1 , \5442_b1 , w_17360 );
or ( \5444_b0 , \5442_b0 , \5443_b0 );
not ( \5443_b0 , w_17361 );
and ( w_17361 , w_17360 , \5443_b1 );
or ( \5445_b1 , \4331_b1 , w_17363 );
not ( w_17363 , w_17364 );
and ( \5445_b0 , \4331_b0 , w_17365 );
and ( w_17364 ,  , w_17365 );
buf ( w_17363 , \5238_b1 );
not ( w_17363 , w_17366 );
not (  , w_17367 );
and ( w_17366 , w_17367 , \5238_b0 );
or ( \5446_b1 , \5444_b1 , w_17369 );
not ( w_17369 , w_17370 );
and ( \5446_b0 , \5444_b0 , w_17371 );
and ( w_17370 ,  , w_17371 );
buf ( w_17369 , \5445_b1 );
not ( w_17369 , w_17372 );
not (  , w_17373 );
and ( w_17372 , w_17373 , \5445_b0 );
or ( \5447_b1 , \5436_b1 , \5446_b1 );
not ( \5446_b1 , w_17374 );
and ( \5447_b0 , \5436_b0 , w_17375 );
and ( w_17374 , w_17375 , \5446_b0 );
or ( \5448_b1 , \5424_b1 , \5435_b1 );
not ( \5435_b1 , w_17376 );
and ( \5448_b0 , \5424_b0 , w_17377 );
and ( w_17376 , w_17377 , \5435_b0 );
or ( \5449_b1 , \5447_b1 , w_17378 );
or ( \5449_b0 , \5447_b0 , \5448_b0 );
not ( \5448_b0 , w_17379 );
and ( w_17379 , w_17378 , \5448_b1 );
or ( \5450_b1 , \5414_b1 , \5449_b1 );
xor ( \5450_b0 , \5414_b0 , w_17380 );
not ( w_17380 , w_17381 );
and ( w_17381 , \5449_b1 , \5449_b0 );
or ( \5451_b1 , \4023_b1 , \3577_b1 );
xor ( \5451_b0 , \4023_b0 , w_17382 );
not ( w_17382 , w_17383 );
and ( w_17383 , \3577_b1 , \3577_b0 );
or ( \5452_b1 , \4229_b1 , w_17385 );
not ( w_17385 , w_17386 );
and ( \5452_b0 , \4229_b0 , w_17387 );
and ( w_17386 ,  , w_17387 );
buf ( w_17385 , \5451_b1 );
not ( w_17385 , w_17388 );
not (  , w_17389 );
and ( w_17388 , w_17389 , \5451_b0 );
or ( \5453_b1 , \5452_b1 , w_17390 );
or ( \5453_b0 , \5452_b0 , \4221_b0 );
not ( \4221_b0 , w_17391 );
and ( w_17391 , w_17390 , \4221_b1 );
or ( \5454_b1 , \4221_b1 , w_17393 );
not ( w_17393 , w_17394 );
and ( \5454_b0 , \4221_b0 , w_17395 );
and ( w_17394 ,  , w_17395 );
buf ( w_17393 , \5283_b1 );
not ( w_17393 , w_17396 );
not (  , w_17397 );
and ( w_17396 , w_17397 , \5283_b0 );
or ( \5455_b1 , \5453_b1 , w_17399 );
not ( w_17399 , w_17400 );
and ( \5455_b0 , \5453_b0 , w_17401 );
and ( w_17400 ,  , w_17401 );
buf ( w_17399 , \5454_b1 );
not ( w_17399 , w_17402 );
not (  , w_17403 );
and ( w_17402 , w_17403 , \5454_b0 );
or ( \5456_b1 , \5346_b1 , w_17404 );
or ( \5456_b0 , \5346_b0 , \4252_b0 );
not ( \4252_b0 , w_17405 );
and ( w_17405 , w_17404 , \4252_b1 );
or ( \5457_b1 , \3108_b1 , \5339_b1 );
not ( \5339_b1 , w_17406 );
and ( \5457_b0 , \3108_b0 , w_17407 );
and ( w_17406 , w_17407 , \5339_b0 );
buf ( \5458_b1 , \3108_b1 );
not ( \5458_b1 , w_17408 );
not ( \5458_b0 , w_17409 );
and ( w_17408 , w_17409 , \3108_b0 );
or ( \5459_b1 , \5458_b1 , \4029_b1 );
not ( \4029_b1 , w_17410 );
and ( \5459_b0 , \5458_b0 , w_17411 );
and ( w_17410 , w_17411 , \4029_b0 );
or ( \5460_b1 , \5457_b1 , w_17412 );
or ( \5460_b0 , \5457_b0 , \5459_b0 );
not ( \5459_b0 , w_17413 );
and ( w_17413 , w_17412 , \5459_b1 );
or ( \5462_b1 , \5456_b1 , w_17415 );
not ( w_17415 , w_17416 );
and ( \5462_b0 , \5456_b0 , w_17417 );
and ( w_17416 ,  , w_17417 );
buf ( w_17415 , \5461_b1 );
not ( w_17415 , w_17418 );
not (  , w_17419 );
and ( w_17418 , w_17419 , \5461_b0 );
or ( \5463_b1 , \5455_b1 , \5462_b1 );
xor ( \5463_b0 , \5455_b0 , w_17420 );
not ( w_17420 , w_17421 );
and ( w_17421 , \5462_b1 , \5462_b0 );
buf ( \5464_b1 , \3963_b1 );
not ( \5464_b1 , w_17422 );
not ( \5464_b0 , w_17423 );
and ( w_17422 , w_17423 , \3963_b0 );
buf ( \5465_b1 , \4176_b1 );
not ( \5465_b1 , w_17424 );
not ( \5465_b0 , w_17425 );
and ( w_17424 , w_17425 , \4176_b0 );
or ( \5466_b1 , \5464_b1 , w_17426 );
or ( \5466_b0 , \5464_b0 , \5465_b0 );
not ( \5465_b0 , w_17427 );
and ( w_17427 , w_17426 , \5465_b1 );
or ( \5467_b1 , \4171_b1 , w_17429 );
not ( w_17429 , w_17430 );
and ( \5467_b0 , \4171_b0 , w_17431 );
and ( w_17430 ,  , w_17431 );
buf ( w_17429 , \4486_b1 );
not ( w_17429 , w_17432 );
not (  , w_17433 );
and ( w_17432 , w_17433 , \4486_b0 );
or ( \5468_b1 , \5466_b1 , w_17435 );
not ( w_17435 , w_17436 );
and ( \5468_b0 , \5466_b0 , w_17437 );
and ( w_17436 ,  , w_17437 );
buf ( w_17435 , \5467_b1 );
not ( w_17435 , w_17438 );
not (  , w_17439 );
and ( w_17438 , w_17439 , \5467_b0 );
buf ( \5469_b1 , \5468_b1 );
not ( \5469_b1 , w_17440 );
not ( \5469_b0 , w_17441 );
and ( w_17440 , w_17441 , \5468_b0 );
buf ( \5470_b1 , \4194_b1 );
not ( \5470_b1 , w_17442 );
not ( \5470_b0 , w_17443 );
and ( w_17442 , w_17443 , \4194_b0 );
or ( \5471_b1 , \5469_b1 , w_17444 );
or ( \5471_b0 , \5469_b0 , \5470_b0 );
not ( \5470_b0 , w_17445 );
and ( w_17445 , w_17444 , \5470_b1 );
or ( \5472_b1 , \4204_b1 , w_17447 );
not ( w_17447 , w_17448 );
and ( \5472_b0 , \4204_b0 , w_17449 );
and ( w_17448 ,  , w_17449 );
buf ( w_17447 , \5296_b1 );
not ( w_17447 , w_17450 );
not (  , w_17451 );
and ( w_17450 , w_17451 , \5296_b0 );
or ( \5473_b1 , \5471_b1 , w_17453 );
not ( w_17453 , w_17454 );
and ( \5473_b0 , \5471_b0 , w_17455 );
and ( w_17454 ,  , w_17455 );
buf ( w_17453 , \5472_b1 );
not ( w_17453 , w_17456 );
not (  , w_17457 );
and ( w_17456 , w_17457 , \5472_b0 );
or ( \5474_b1 , \5463_b1 , \5473_b1 );
not ( \5473_b1 , w_17458 );
and ( \5474_b0 , \5463_b0 , w_17459 );
and ( w_17458 , w_17459 , \5473_b0 );
or ( \5475_b1 , \5455_b1 , \5462_b1 );
not ( \5462_b1 , w_17460 );
and ( \5475_b0 , \5455_b0 , w_17461 );
and ( w_17460 , w_17461 , \5462_b0 );
or ( \5476_b1 , \5474_b1 , w_17462 );
or ( \5476_b0 , \5474_b0 , \5475_b0 );
not ( \5475_b0 , w_17463 );
and ( w_17463 , w_17462 , \5475_b1 );
or ( \5477_b1 , \5450_b1 , \5476_b1 );
not ( \5476_b1 , w_17464 );
and ( \5477_b0 , \5450_b0 , w_17465 );
and ( w_17464 , w_17465 , \5476_b0 );
or ( \5478_b1 , \5414_b1 , \5449_b1 );
not ( \5449_b1 , w_17466 );
and ( \5478_b0 , \5414_b0 , w_17467 );
and ( w_17466 , w_17467 , \5449_b0 );
or ( \5479_b1 , \5477_b1 , w_17468 );
or ( \5479_b0 , \5477_b0 , \5478_b0 );
not ( \5478_b0 , w_17469 );
and ( w_17469 , w_17468 , \5478_b1 );
buf ( \5480_b1 , \5479_b1 );
not ( \5480_b1 , w_17470 );
not ( \5480_b0 , w_17471 );
and ( w_17470 , w_17471 , \5479_b0 );
buf ( \5481_b1 , \5480_b1 );
not ( \5481_b1 , w_17472 );
not ( \5481_b0 , w_17473 );
and ( w_17472 , w_17473 , \5480_b0 );
or ( \5482_b1 , \5277_b1 , \5301_b1 );
xor ( \5482_b0 , \5277_b0 , w_17474 );
not ( w_17474 , w_17475 );
and ( w_17475 , \5301_b1 , \5301_b0 );
or ( \5483_b1 , \5482_b1 , w_17476 );
xor ( \5483_b0 , \5482_b0 , w_17478 );
not ( w_17478 , w_17479 );
and ( w_17479 , w_17476 , w_17477 );
buf ( w_17476 , \5288_b1 );
not ( w_17476 , w_17480 );
not ( w_17477 , w_17481 );
and ( w_17480 , w_17481 , \5288_b0 );
buf ( \5484_b1 , \5483_b1 );
not ( \5484_b1 , w_17482 );
not ( \5484_b0 , w_17483 );
and ( w_17482 , w_17483 , \5483_b0 );
or ( \5485_b1 , \5220_b1 , \5231_b1 );
xor ( \5485_b0 , \5220_b0 , w_17484 );
not ( w_17484 , w_17485 );
and ( w_17485 , \5231_b1 , \5231_b0 );
or ( \5486_b1 , \5485_b1 , \5243_b1 );
xor ( \5486_b0 , \5485_b0 , w_17486 );
not ( w_17486 , w_17487 );
and ( w_17487 , \5243_b1 , \5243_b0 );
buf ( \5487_b1 , \5486_b1 );
not ( \5487_b1 , w_17488 );
not ( \5487_b0 , w_17489 );
and ( w_17488 , w_17489 , \5486_b0 );
buf ( \5488_b1 , \5487_b1 );
not ( \5488_b1 , w_17490 );
not ( \5488_b0 , w_17491 );
and ( w_17490 , w_17491 , \5487_b0 );
or ( \5489_b1 , \5484_b1 , w_17492 );
or ( \5489_b0 , \5484_b0 , \5488_b0 );
not ( \5488_b0 , w_17493 );
and ( w_17493 , w_17492 , \5488_b1 );
or ( \5490_b1 , \5487_b1 , w_17494 );
or ( \5490_b0 , \5487_b0 , \5483_b0 );
not ( \5483_b0 , w_17495 );
and ( w_17495 , w_17494 , \5483_b1 );
or ( \5491_b1 , \5340_b1 , \5352_b1 );
xor ( \5491_b0 , \5340_b0 , w_17496 );
not ( w_17496 , w_17497 );
and ( w_17497 , \5352_b1 , \5352_b0 );
or ( \5492_b1 , \5491_b1 , \5365_b1 );
xor ( \5492_b0 , \5491_b0 , w_17498 );
not ( w_17498 , w_17499 );
and ( w_17499 , \5365_b1 , \5365_b0 );
or ( \5493_b1 , \5490_b1 , w_17501 );
not ( w_17501 , w_17502 );
and ( \5493_b0 , \5490_b0 , w_17503 );
and ( w_17502 ,  , w_17503 );
buf ( w_17501 , \5492_b1 );
not ( w_17501 , w_17504 );
not (  , w_17505 );
and ( w_17504 , w_17505 , \5492_b0 );
or ( \5494_b1 , \5489_b1 , w_17507 );
not ( w_17507 , w_17508 );
and ( \5494_b0 , \5489_b0 , w_17509 );
and ( w_17508 ,  , w_17509 );
buf ( w_17507 , \5493_b1 );
not ( w_17507 , w_17510 );
not (  , w_17511 );
and ( w_17510 , w_17511 , \5493_b0 );
buf ( \5495_b1 , \5494_b1 );
not ( \5495_b1 , w_17512 );
not ( \5495_b0 , w_17513 );
and ( w_17512 , w_17513 , \5494_b0 );
buf ( \5496_b1 , \5495_b1 );
not ( \5496_b1 , w_17514 );
not ( \5496_b0 , w_17515 );
and ( w_17514 , w_17515 , \5495_b0 );
or ( \5497_b1 , \5481_b1 , w_17516 );
or ( \5497_b0 , \5481_b0 , \5496_b0 );
not ( \5496_b0 , w_17517 );
and ( w_17517 , w_17516 , \5496_b1 );
or ( \5498_b1 , \5330_b1 , \5337_b1 );
xor ( \5498_b0 , \5330_b0 , w_17518 );
not ( w_17518 , w_17519 );
and ( w_17519 , \5337_b1 , \5337_b0 );
or ( \5499_b1 , \5498_b1 , w_17520 );
xor ( \5499_b0 , \5498_b0 , w_17522 );
not ( w_17522 , w_17523 );
and ( w_17523 , w_17520 , w_17521 );
buf ( w_17520 , \5368_b1 );
not ( w_17520 , w_17524 );
not ( w_17521 , w_17525 );
and ( w_17524 , w_17525 , \5368_b0 );
or ( \5500_b1 , \5497_b1 , w_17527 );
not ( w_17527 , w_17528 );
and ( \5500_b0 , \5497_b0 , w_17529 );
and ( w_17528 ,  , w_17529 );
buf ( w_17527 , \5499_b1 );
not ( w_17527 , w_17530 );
not (  , w_17531 );
and ( w_17530 , w_17531 , \5499_b0 );
buf ( \5501_b1 , \5495_b1 );
not ( \5501_b1 , w_17532 );
not ( \5501_b0 , w_17533 );
and ( w_17532 , w_17533 , \5495_b0 );
or ( \5502_b1 , \5501_b1 , w_17535 );
not ( w_17535 , w_17536 );
and ( \5502_b0 , \5501_b0 , w_17537 );
and ( w_17536 ,  , w_17537 );
buf ( w_17535 , \5479_b1 );
not ( w_17535 , w_17538 );
not (  , w_17539 );
and ( w_17538 , w_17539 , \5479_b0 );
or ( \5503_b1 , \5500_b1 , \5502_b1 );
not ( \5502_b1 , w_17540 );
and ( \5503_b0 , \5500_b0 , w_17541 );
and ( w_17540 , w_17541 , \5502_b0 );
or ( \5504_b1 , \5387_b1 , \5503_b1 );
xor ( \5504_b0 , \5387_b0 , w_17542 );
not ( w_17542 , w_17543 );
and ( w_17543 , \5503_b1 , \5503_b0 );
or ( \5505_b1 , \5372_b1 , \5324_b1 );
xor ( \5505_b0 , \5372_b0 , w_17544 );
not ( w_17544 , w_17545 );
and ( w_17545 , \5324_b1 , \5324_b0 );
or ( \5506_b1 , \5505_b1 , w_17546 );
xor ( \5506_b0 , \5505_b0 , w_17548 );
not ( w_17548 , w_17549 );
and ( w_17549 , w_17546 , w_17547 );
buf ( w_17546 , \5317_b1 );
not ( w_17546 , w_17550 );
not ( w_17547 , w_17551 );
and ( w_17550 , w_17551 , \5317_b0 );
or ( \5507_b1 , \5504_b1 , \5506_b1 );
not ( \5506_b1 , w_17552 );
and ( \5507_b0 , \5504_b0 , w_17553 );
and ( w_17552 , w_17553 , \5506_b0 );
or ( \5508_b1 , \5387_b1 , \5503_b1 );
not ( \5503_b1 , w_17554 );
and ( \5508_b0 , \5387_b0 , w_17555 );
and ( w_17554 , w_17555 , \5503_b0 );
or ( \5509_b1 , \5507_b1 , w_17556 );
or ( \5509_b0 , \5507_b0 , \5508_b0 );
not ( \5508_b0 , w_17557 );
and ( w_17557 , w_17556 , \5508_b1 );
or ( \5510_b1 , \5385_b1 , w_17559 );
not ( w_17559 , w_17560 );
and ( \5510_b0 , \5385_b0 , w_17561 );
and ( w_17560 ,  , w_17561 );
buf ( w_17559 , \5509_b1 );
not ( w_17559 , w_17562 );
not (  , w_17563 );
and ( w_17562 , w_17563 , \5509_b0 );
or ( \5511_b1 , \5383_b1 , \5510_b1 );
not ( \5510_b1 , w_17564 );
and ( \5511_b0 , \5383_b0 , w_17565 );
and ( w_17564 , w_17565 , \5510_b0 );
or ( \5512_b1 , \4472_b1 , \4504_b1 );
not ( \4504_b1 , w_17566 );
and ( \5512_b0 , \4472_b0 , w_17567 );
and ( w_17566 , w_17567 , \4504_b0 );
buf ( \5513_b1 , \4472_b1 );
not ( \5513_b1 , w_17568 );
not ( \5513_b0 , w_17569 );
and ( w_17568 , w_17569 , \4472_b0 );
or ( \5514_b1 , \5513_b1 , \4505_b1 );
not ( \4505_b1 , w_17570 );
and ( \5514_b0 , \5513_b0 , w_17571 );
and ( w_17570 , w_17571 , \4505_b0 );
or ( \5515_b1 , \5512_b1 , w_17572 );
or ( \5515_b0 , \5512_b0 , \5514_b0 );
not ( \5514_b0 , w_17573 );
and ( w_17573 , w_17572 , \5514_b1 );
or ( \5516_b1 , \5515_b1 , \4464_b1 );
not ( \4464_b1 , w_17574 );
and ( \5516_b0 , \5515_b0 , w_17575 );
and ( w_17574 , w_17575 , \4464_b0 );
buf ( \5517_b1 , \5515_b1 );
not ( \5517_b1 , w_17576 );
not ( \5517_b0 , w_17577 );
and ( w_17576 , w_17577 , \5515_b0 );
buf ( \5518_b1 , \4464_b1 );
not ( \5518_b1 , w_17578 );
not ( \5518_b0 , w_17579 );
and ( w_17578 , w_17579 , \4464_b0 );
or ( \5519_b1 , \5517_b1 , \5518_b1 );
not ( \5518_b1 , w_17580 );
and ( \5519_b0 , \5517_b0 , w_17581 );
and ( w_17580 , w_17581 , \5518_b0 );
or ( \5520_b1 , \5516_b1 , w_17583 );
not ( w_17583 , w_17584 );
and ( \5520_b0 , \5516_b0 , w_17585 );
and ( w_17584 ,  , w_17585 );
buf ( w_17583 , \5519_b1 );
not ( w_17583 , w_17586 );
not (  , w_17587 );
and ( w_17586 , w_17587 , \5519_b0 );
buf ( \5521_b1 , \4617_b1 );
not ( \5521_b1 , w_17588 );
not ( \5521_b0 , w_17589 );
and ( w_17588 , w_17589 , \4617_b0 );
buf ( \5522_b1 , \4627_b1 );
not ( \5522_b1 , w_17590 );
not ( \5522_b0 , w_17591 );
and ( w_17590 , w_17591 , \4627_b0 );
or ( \5523_b1 , \5521_b1 , w_17592 );
or ( \5523_b0 , \5521_b0 , \5522_b0 );
not ( \5522_b0 , w_17593 );
and ( w_17593 , w_17592 , \5522_b1 );
or ( \5524_b1 , \4617_b1 , w_17594 );
or ( \5524_b0 , \4617_b0 , \4627_b0 );
not ( \4627_b0 , w_17595 );
and ( w_17595 , w_17594 , \4627_b1 );
or ( \5525_b1 , \5523_b1 , w_17597 );
not ( w_17597 , w_17598 );
and ( \5525_b0 , \5523_b0 , w_17599 );
and ( w_17598 ,  , w_17599 );
buf ( w_17597 , \5524_b1 );
not ( w_17597 , w_17600 );
not (  , w_17601 );
and ( w_17600 , w_17601 , \5524_b0 );
or ( \5526_b1 , \4684_b1 , \5525_b1 );
not ( \5525_b1 , w_17602 );
and ( \5526_b0 , \4684_b0 , w_17603 );
and ( w_17602 , w_17603 , \5525_b0 );
buf ( \5527_b1 , \4684_b1 );
not ( \5527_b1 , w_17604 );
not ( \5527_b0 , w_17605 );
and ( w_17604 , w_17605 , \4684_b0 );
buf ( \5528_b1 , \5525_b1 );
not ( \5528_b1 , w_17606 );
not ( \5528_b0 , w_17607 );
and ( w_17606 , w_17607 , \5525_b0 );
or ( \5529_b1 , \5527_b1 , \5528_b1 );
not ( \5528_b1 , w_17608 );
and ( \5529_b0 , \5527_b0 , w_17609 );
and ( w_17608 , w_17609 , \5528_b0 );
or ( \5530_b1 , \5526_b1 , w_17611 );
not ( w_17611 , w_17612 );
and ( \5530_b0 , \5526_b0 , w_17613 );
and ( w_17612 ,  , w_17613 );
buf ( w_17611 , \5529_b1 );
not ( w_17611 , w_17614 );
not (  , w_17615 );
and ( w_17614 , w_17615 , \5529_b0 );
or ( \5531_b1 , \5520_b1 , \5530_b1 );
xor ( \5531_b0 , \5520_b0 , w_17616 );
not ( w_17616 , w_17617 );
and ( w_17617 , \5530_b1 , \5530_b0 );
buf ( \5532_b1 , \5124_b1 );
not ( \5532_b1 , w_17618 );
not ( \5532_b0 , w_17619 );
and ( w_17618 , w_17619 , \5124_b0 );
buf ( \5533_b1 , \5046_b1 );
not ( \5533_b1 , w_17620 );
not ( \5533_b0 , w_17621 );
and ( w_17620 , w_17621 , \5046_b0 );
or ( \5534_b1 , \5532_b1 , w_17622 );
or ( \5534_b0 , \5532_b0 , \5533_b0 );
not ( \5533_b0 , w_17623 );
and ( w_17623 , w_17622 , \5533_b1 );
or ( \5535_b1 , \5534_b1 , w_17625 );
not ( w_17625 , w_17626 );
and ( \5535_b0 , \5534_b0 , w_17627 );
and ( w_17626 ,  , w_17627 );
buf ( w_17625 , \5117_b1 );
not ( w_17625 , w_17628 );
not (  , w_17629 );
and ( w_17628 , w_17629 , \5117_b0 );
or ( \5536_b1 , \5124_b1 , w_17630 );
or ( \5536_b0 , \5124_b0 , \5046_b0 );
not ( \5046_b0 , w_17631 );
and ( w_17631 , w_17630 , \5046_b1 );
or ( \5537_b1 , \5535_b1 , w_17633 );
not ( w_17633 , w_17634 );
and ( \5537_b0 , \5535_b0 , w_17635 );
and ( w_17634 ,  , w_17635 );
buf ( w_17633 , \5536_b1 );
not ( w_17633 , w_17636 );
not (  , w_17637 );
and ( w_17636 , w_17637 , \5536_b0 );
or ( \5538_b1 , \5531_b1 , \5537_b1 );
xor ( \5538_b0 , \5531_b0 , w_17638 );
not ( w_17638 , w_17639 );
and ( w_17639 , \5537_b1 , \5537_b0 );
or ( \5539_b1 , \5044_b1 , \5125_b1 );
xor ( \5539_b0 , \5044_b0 , w_17640 );
not ( w_17640 , w_17641 );
and ( w_17641 , \5125_b1 , \5125_b0 );
or ( \5540_b1 , \5539_b1 , \5205_b1 );
not ( \5205_b1 , w_17642 );
and ( \5540_b0 , \5539_b0 , w_17643 );
and ( w_17642 , w_17643 , \5205_b0 );
or ( \5541_b1 , \5044_b1 , \5125_b1 );
not ( \5125_b1 , w_17644 );
and ( \5541_b0 , \5044_b0 , w_17645 );
and ( w_17644 , w_17645 , \5125_b0 );
or ( \5542_b1 , \5540_b1 , w_17646 );
or ( \5542_b0 , \5540_b0 , \5541_b0 );
not ( \5541_b0 , w_17647 );
and ( w_17647 , w_17646 , \5541_b1 );
or ( \5543_b1 , \5538_b1 , w_17649 );
not ( w_17649 , w_17650 );
and ( \5543_b0 , \5538_b0 , w_17651 );
and ( w_17650 ,  , w_17651 );
buf ( w_17649 , \5542_b1 );
not ( w_17649 , w_17652 );
not (  , w_17653 );
and ( w_17652 , w_17653 , \5542_b0 );
buf ( \5544_b1 , \5520_b1 );
not ( \5544_b1 , w_17654 );
not ( \5544_b0 , w_17655 );
and ( w_17654 , w_17655 , \5520_b0 );
buf ( \5545_b1 , \5530_b1 );
not ( \5545_b1 , w_17656 );
not ( \5545_b0 , w_17657 );
and ( w_17656 , w_17657 , \5530_b0 );
buf ( \5546_b1 , \5545_b1 );
not ( \5546_b1 , w_17658 );
not ( \5546_b0 , w_17659 );
and ( w_17658 , w_17659 , \5545_b0 );
or ( \5547_b1 , \5544_b1 , w_17660 );
or ( \5547_b0 , \5544_b0 , \5546_b0 );
not ( \5546_b0 , w_17661 );
and ( w_17661 , w_17660 , \5546_b1 );
buf ( \5548_b1 , \5520_b1 );
not ( \5548_b1 , w_17662 );
not ( \5548_b0 , w_17663 );
and ( w_17662 , w_17663 , \5520_b0 );
buf ( \5549_b1 , \5548_b1 );
not ( \5549_b1 , w_17664 );
not ( \5549_b0 , w_17665 );
and ( w_17664 , w_17665 , \5548_b0 );
buf ( \5550_b1 , \5530_b1 );
not ( \5550_b1 , w_17666 );
not ( \5550_b0 , w_17667 );
and ( w_17666 , w_17667 , \5530_b0 );
or ( \5551_b1 , \5549_b1 , w_17668 );
or ( \5551_b0 , \5549_b0 , \5550_b0 );
not ( \5550_b0 , w_17669 );
and ( w_17669 , w_17668 , \5550_b1 );
or ( \5552_b1 , \5551_b1 , w_17671 );
not ( w_17671 , w_17672 );
and ( \5552_b0 , \5551_b0 , w_17673 );
and ( w_17672 ,  , w_17673 );
buf ( w_17671 , \5537_b1 );
not ( w_17671 , w_17674 );
not (  , w_17675 );
and ( w_17674 , w_17675 , \5537_b0 );
or ( \5553_b1 , \5547_b1 , w_17677 );
not ( w_17677 , w_17678 );
and ( \5553_b0 , \5547_b0 , w_17679 );
and ( w_17678 ,  , w_17679 );
buf ( w_17677 , \5552_b1 );
not ( w_17677 , w_17680 );
not (  , w_17681 );
and ( w_17680 , w_17681 , \5552_b0 );
buf ( \5554_b1 , \5553_b1 );
not ( \5554_b1 , w_17682 );
not ( \5554_b0 , w_17683 );
and ( w_17682 , w_17683 , \5553_b0 );
or ( \5555_b1 , \4518_b1 , \4530_b1 );
xor ( \5555_b0 , \4518_b0 , w_17684 );
not ( w_17684 , w_17685 );
and ( w_17685 , \4530_b1 , \4530_b0 );
or ( \5556_b1 , \5555_b1 , w_17686 );
xor ( \5556_b0 , \5555_b0 , w_17688 );
not ( w_17688 , w_17689 );
and ( w_17689 , w_17686 , w_17687 );
buf ( w_17686 , \4690_b1 );
not ( w_17686 , w_17690 );
not ( w_17687 , w_17691 );
and ( w_17690 , w_17691 , \4690_b0 );
or ( \5557_b1 , \5554_b1 , w_17693 );
not ( w_17693 , w_17694 );
and ( \5557_b0 , \5554_b0 , w_17695 );
and ( w_17694 ,  , w_17695 );
buf ( w_17693 , \5556_b1 );
not ( w_17693 , w_17696 );
not (  , w_17697 );
and ( w_17696 , w_17697 , \5556_b0 );
or ( \5558_b1 , \5543_b1 , w_17699 );
not ( w_17699 , w_17700 );
and ( \5558_b0 , \5543_b0 , w_17701 );
and ( w_17700 ,  , w_17701 );
buf ( w_17699 , \5557_b1 );
not ( w_17699 , w_17702 );
not (  , w_17703 );
and ( w_17702 , w_17703 , \5557_b0 );
buf ( \5559_b1 , \5558_b1 );
not ( \5559_b1 , w_17704 );
not ( \5559_b0 , w_17705 );
and ( w_17704 , w_17705 , \5558_b0 );
or ( \5560_b1 , \5511_b1 , \5559_b1 );
not ( \5559_b1 , w_17706 );
and ( \5560_b0 , \5511_b0 , w_17707 );
and ( w_17706 , w_17707 , \5559_b0 );
buf ( \5561_b1 , \5560_b1 );
not ( \5561_b1 , w_17708 );
not ( \5561_b0 , w_17709 );
and ( w_17708 , w_17709 , \5560_b0 );
or ( \5562_b1 , \5387_b1 , \5503_b1 );
xor ( \5562_b0 , \5387_b0 , w_17710 );
not ( w_17710 , w_17711 );
and ( w_17711 , \5503_b1 , \5503_b0 );
or ( \5563_b1 , \5562_b1 , \5506_b1 );
xor ( \5563_b0 , \5562_b0 , w_17712 );
not ( w_17712 , w_17713 );
and ( w_17713 , \5506_b1 , \5506_b0 );
or ( \5564_b1 , \5308_b1 , \5305_b1 );
not ( \5305_b1 , w_17714 );
and ( \5564_b0 , \5308_b0 , w_17715 );
and ( w_17714 , w_17715 , \5305_b0 );
buf ( \5565_b1 , \5308_b1 );
not ( \5565_b1 , w_17716 );
not ( \5565_b0 , w_17717 );
and ( w_17716 , w_17717 , \5308_b0 );
or ( \5566_b1 , \5565_b1 , \5306_b1 );
not ( \5306_b1 , w_17718 );
and ( \5566_b0 , \5565_b0 , w_17719 );
and ( w_17718 , w_17719 , \5306_b0 );
or ( \5567_b1 , \5564_b1 , w_17720 );
or ( \5567_b0 , \5564_b0 , \5566_b0 );
not ( \5566_b0 , w_17721 );
and ( w_17721 , w_17720 , \5566_b1 );
or ( \5568_b1 , \5567_b1 , w_17722 );
xor ( \5568_b0 , \5567_b0 , w_17724 );
not ( w_17724 , w_17725 );
and ( w_17725 , w_17722 , w_17723 );
buf ( w_17722 , \5314_b1 );
not ( w_17722 , w_17726 );
not ( w_17723 , w_17727 );
and ( w_17726 , w_17727 , \5314_b0 );
buf ( \5569_b1 , \5388_b1 );
not ( \5569_b1 , w_17728 );
not ( \5569_b0 , w_17729 );
and ( w_17728 , w_17729 , \5388_b0 );
buf ( \5570_b1 , \4244_b1 );
not ( \5570_b1 , w_17730 );
not ( \5570_b0 , w_17731 );
and ( w_17730 , w_17731 , \4244_b0 );
or ( \5571_b1 , \5569_b1 , w_17732 );
or ( \5571_b0 , \5569_b0 , \5570_b0 );
not ( \5570_b0 , w_17733 );
and ( w_17733 , w_17732 , \5570_b1 );
or ( \5572_b1 , \5571_b1 , w_17735 );
not ( w_17735 , w_17736 );
and ( \5572_b0 , \5571_b0 , w_17737 );
and ( w_17736 ,  , w_17737 );
buf ( w_17735 , \4492_b1 );
not ( w_17735 , w_17738 );
not (  , w_17739 );
and ( w_17738 , w_17739 , \4492_b0 );
or ( \5573_b1 , \4245_b1 , w_17741 );
not ( w_17741 , w_17742 );
and ( \5573_b0 , \4245_b0 , w_17743 );
and ( w_17742 ,  , w_17743 );
buf ( w_17741 , \4048_b1 );
not ( w_17741 , w_17744 );
not (  , w_17745 );
and ( w_17744 , w_17745 , \4048_b0 );
buf ( \5575_b1 , \3943_b1 );
not ( \5575_b1 , w_17746 );
not ( \5575_b0 , w_17747 );
and ( w_17746 , w_17747 , \3943_b0 );
buf ( \5576_b1 , \5016_b1 );
not ( \5576_b1 , w_17748 );
not ( \5576_b0 , w_17749 );
and ( w_17748 , w_17749 , \5016_b0 );
buf ( \5577_b1 , \5576_b1 );
not ( \5577_b1 , w_17750 );
not ( \5577_b0 , w_17751 );
and ( w_17750 , w_17751 , \5576_b0 );
or ( \5578_b1 , \5575_b1 , w_17752 );
or ( \5578_b0 , \5575_b0 , \5577_b0 );
not ( \5577_b0 , w_17753 );
and ( w_17753 , w_17752 , \5577_b1 );
or ( \5579_b1 , \5016_b1 , w_17755 );
not ( w_17755 , w_17756 );
and ( \5579_b0 , \5016_b0 , w_17757 );
and ( w_17756 ,  , w_17757 );
buf ( w_17755 , \4147_b1 );
not ( w_17755 , w_17758 );
not (  , w_17759 );
and ( w_17758 , w_17759 , \4147_b0 );
or ( \5580_b1 , \5578_b1 , w_17761 );
not ( w_17761 , w_17762 );
and ( \5580_b0 , \5578_b0 , w_17763 );
and ( w_17762 ,  , w_17763 );
buf ( w_17761 , \5579_b1 );
not ( w_17761 , w_17764 );
not (  , w_17765 );
and ( w_17764 , w_17765 , \5579_b0 );
buf ( \5581_b1 , \5580_b1 );
not ( \5581_b1 , w_17766 );
not ( \5581_b0 , w_17767 );
and ( w_17766 , w_17767 , \5580_b0 );
buf ( \5582_b1 , \5019_b1 );
not ( \5582_b1 , w_17768 );
not ( \5582_b0 , w_17769 );
and ( w_17768 , w_17769 , \5019_b0 );
or ( \5583_b1 , \5581_b1 , w_17770 );
or ( \5583_b0 , \5581_b0 , \5582_b0 );
not ( \5582_b0 , w_17771 );
and ( w_17771 , w_17770 , \5582_b1 );
or ( \5584_b1 , \5396_b1 , w_17773 );
not ( w_17773 , w_17774 );
and ( \5584_b0 , \5396_b0 , w_17775 );
and ( w_17774 ,  , w_17775 );
buf ( w_17773 , \5021_b1 );
not ( w_17773 , w_17776 );
not (  , w_17777 );
and ( w_17776 , w_17777 , \5021_b0 );
or ( \5585_b1 , \5583_b1 , w_17779 );
not ( w_17779 , w_17780 );
and ( \5585_b0 , \5583_b0 , w_17781 );
and ( w_17780 ,  , w_17781 );
buf ( w_17779 , \5584_b1 );
not ( w_17779 , w_17782 );
not (  , w_17783 );
and ( w_17782 , w_17783 , \5584_b0 );
or ( \5586_b1 , \5574_b1 , \5585_b1 );
not ( \5585_b1 , w_17784 );
and ( \5586_b0 , \5574_b0 , w_17785 );
and ( w_17784 , w_17785 , \5585_b0 );
or ( \5587_b1 , \5389_b1 , \5400_b1 );
xor ( \5587_b0 , \5389_b0 , w_17786 );
not ( w_17786 , w_17787 );
and ( w_17787 , \5400_b1 , \5400_b0 );
or ( \5588_b1 , \5587_b1 , \5411_b1 );
xor ( \5588_b0 , \5587_b0 , w_17788 );
not ( w_17788 , w_17789 );
and ( w_17789 , \5411_b1 , \5411_b0 );
or ( \5589_b1 , \5586_b1 , \5588_b1 );
xor ( \5589_b0 , \5586_b0 , w_17790 );
not ( w_17790 , w_17791 );
and ( w_17791 , \5588_b1 , \5588_b0 );
buf ( \5590_b1 , \4011_b1 );
not ( \5590_b1 , w_17792 );
not ( \5590_b0 , w_17793 );
and ( w_17792 , w_17793 , \4011_b0 );
buf ( \5591_b1 , \5234_b1 );
not ( \5591_b1 , w_17794 );
not ( \5591_b0 , w_17795 );
and ( w_17794 , w_17795 , \5234_b0 );
or ( \5592_b1 , \5590_b1 , w_17796 );
or ( \5592_b0 , \5590_b0 , \5591_b0 );
not ( \5591_b0 , w_17797 );
and ( w_17797 , w_17796 , \5591_b1 );
or ( \5593_b1 , \4088_b1 , w_17799 );
not ( w_17799 , w_17800 );
and ( \5593_b0 , \4088_b0 , w_17801 );
and ( w_17800 ,  , w_17801 );
buf ( w_17799 , \4270_b1 );
not ( w_17799 , w_17802 );
not (  , w_17803 );
and ( w_17802 , w_17803 , \4270_b0 );
or ( \5594_b1 , \5592_b1 , w_17805 );
not ( w_17805 , w_17806 );
and ( \5594_b0 , \5592_b0 , w_17807 );
and ( w_17806 ,  , w_17807 );
buf ( w_17805 , \5593_b1 );
not ( w_17805 , w_17808 );
not (  , w_17809 );
and ( w_17808 , w_17809 , \5593_b0 );
buf ( \5595_b1 , \5594_b1 );
not ( \5595_b1 , w_17810 );
not ( \5595_b0 , w_17811 );
and ( w_17810 , w_17811 , \5594_b0 );
buf ( \5596_b1 , \4437_b1 );
not ( \5596_b1 , w_17812 );
not ( \5596_b0 , w_17813 );
and ( w_17812 , w_17813 , \4437_b0 );
or ( \5597_b1 , \5595_b1 , w_17814 );
or ( \5597_b0 , \5595_b0 , \5596_b0 );
not ( \5596_b0 , w_17815 );
and ( w_17815 , w_17814 , \5596_b1 );
or ( \5598_b1 , \4596_b1 , w_17817 );
not ( w_17817 , w_17818 );
and ( \5598_b0 , \4596_b0 , w_17819 );
and ( w_17818 ,  , w_17819 );
buf ( w_17817 , \5441_b1 );
not ( w_17817 , w_17820 );
not (  , w_17821 );
and ( w_17820 , w_17821 , \5441_b0 );
or ( \5599_b1 , \5597_b1 , w_17823 );
not ( w_17823 , w_17824 );
and ( \5599_b0 , \5597_b0 , w_17825 );
and ( w_17824 ,  , w_17825 );
buf ( w_17823 , \5598_b1 );
not ( w_17823 , w_17826 );
not (  , w_17827 );
and ( w_17826 , w_17827 , \5598_b0 );
buf ( \5600_b1 , \3958_b1 );
not ( \5600_b1 , w_17828 );
not ( \5600_b0 , w_17829 );
and ( w_17828 , w_17829 , \3958_b0 );
buf ( \5601_b1 , \4142_b1 );
not ( \5601_b1 , w_17830 );
not ( \5601_b0 , w_17831 );
and ( w_17830 , w_17831 , \4142_b0 );
or ( \5602_b1 , \5600_b1 , w_17832 );
or ( \5602_b0 , \5600_b0 , \5601_b0 );
not ( \5601_b0 , w_17833 );
and ( w_17833 , w_17832 , \5601_b1 );
or ( \5603_b1 , \4109_b1 , w_17835 );
not ( w_17835 , w_17836 );
and ( \5603_b0 , \4109_b0 , w_17837 );
and ( w_17836 ,  , w_17837 );
buf ( w_17835 , \4473_b1 );
not ( w_17835 , w_17838 );
not (  , w_17839 );
and ( w_17838 , w_17839 , \4473_b0 );
or ( \5604_b1 , \5602_b1 , w_17841 );
not ( w_17841 , w_17842 );
and ( \5604_b0 , \5602_b0 , w_17843 );
and ( w_17842 ,  , w_17843 );
buf ( w_17841 , \5603_b1 );
not ( w_17841 , w_17844 );
not (  , w_17845 );
and ( w_17844 , w_17845 , \5603_b0 );
buf ( \5605_b1 , \5604_b1 );
not ( \5605_b1 , w_17846 );
not ( \5605_b0 , w_17847 );
and ( w_17846 , w_17847 , \5604_b0 );
buf ( \5606_b1 , \4425_b1 );
not ( \5606_b1 , w_17848 );
not ( \5606_b0 , w_17849 );
and ( w_17848 , w_17849 , \4425_b0 );
or ( \5607_b1 , \5605_b1 , w_17850 );
or ( \5607_b0 , \5605_b0 , \5606_b0 );
not ( \5606_b0 , w_17851 );
and ( w_17851 , w_17850 , \5606_b1 );
or ( \5608_b1 , \4139_b1 , w_17853 );
not ( w_17853 , w_17854 );
and ( \5608_b0 , \4139_b0 , w_17855 );
and ( w_17854 ,  , w_17855 );
buf ( w_17853 , \5429_b1 );
not ( w_17853 , w_17856 );
not (  , w_17857 );
and ( w_17856 , w_17857 , \5429_b0 );
or ( \5609_b1 , \5607_b1 , w_17859 );
not ( w_17859 , w_17860 );
and ( \5609_b0 , \5607_b0 , w_17861 );
and ( w_17860 ,  , w_17861 );
buf ( w_17859 , \5608_b1 );
not ( w_17859 , w_17862 );
not (  , w_17863 );
and ( w_17862 , w_17863 , \5608_b0 );
or ( \5610_b1 , \5599_b1 , w_17865 );
not ( w_17865 , w_17866 );
and ( \5610_b0 , \5599_b0 , w_17867 );
and ( w_17866 ,  , w_17867 );
buf ( w_17865 , \5609_b1 );
not ( w_17865 , w_17868 );
not (  , w_17869 );
and ( w_17868 , w_17869 , \5609_b0 );
buf ( \5611_b1 , \4047_b1 );
not ( \5611_b1 , w_17870 );
not ( \5611_b0 , w_17871 );
and ( w_17870 , w_17871 , \4047_b0 );
buf ( \5612_b1 , \4666_b1 );
not ( \5612_b1 , w_17872 );
not ( \5612_b0 , w_17873 );
and ( w_17872 , w_17873 , \4666_b0 );
or ( \5613_b1 , \5611_b1 , w_17874 );
or ( \5613_b0 , \5611_b0 , \5612_b0 );
not ( \5612_b0 , w_17875 );
and ( w_17875 , w_17874 , \5612_b1 );
or ( \5614_b1 , \4548_b1 , w_17877 );
not ( w_17877 , w_17878 );
and ( \5614_b0 , \4548_b0 , w_17879 );
and ( w_17878 ,  , w_17879 );
buf ( w_17877 , \4178_b1 );
not ( w_17877 , w_17880 );
not (  , w_17881 );
and ( w_17880 , w_17881 , \4178_b0 );
or ( \5615_b1 , \5613_b1 , w_17883 );
not ( w_17883 , w_17884 );
and ( \5615_b0 , \5613_b0 , w_17885 );
and ( w_17884 ,  , w_17885 );
buf ( w_17883 , \5614_b1 );
not ( w_17883 , w_17886 );
not (  , w_17887 );
and ( w_17886 , w_17887 , \5614_b0 );
buf ( \5616_b1 , \5615_b1 );
not ( \5616_b1 , w_17888 );
not ( \5616_b0 , w_17889 );
and ( w_17888 , w_17889 , \5615_b0 );
buf ( \5617_b1 , \4661_b1 );
not ( \5617_b1 , w_17890 );
not ( \5617_b0 , w_17891 );
and ( w_17890 , w_17891 , \4661_b0 );
or ( \5618_b1 , \5616_b1 , w_17892 );
or ( \5618_b0 , \5616_b0 , \5617_b0 );
not ( \5617_b0 , w_17893 );
and ( w_17893 , w_17892 , \5617_b1 );
or ( \5619_b1 , \4672_b1 , w_17895 );
not ( w_17895 , w_17896 );
and ( \5619_b0 , \4672_b0 , w_17897 );
and ( w_17896 ,  , w_17897 );
buf ( w_17895 , \5406_b1 );
not ( w_17895 , w_17898 );
not (  , w_17899 );
and ( w_17898 , w_17899 , \5406_b0 );
or ( \5620_b1 , \5618_b1 , w_17901 );
not ( w_17901 , w_17902 );
and ( \5620_b0 , \5618_b0 , w_17903 );
and ( w_17902 ,  , w_17903 );
buf ( w_17901 , \5619_b1 );
not ( w_17901 , w_17904 );
not (  , w_17905 );
and ( w_17904 , w_17905 , \5619_b0 );
buf ( \5621_b1 , \5620_b1 );
not ( \5621_b1 , w_17906 );
not ( \5621_b0 , w_17907 );
and ( w_17906 , w_17907 , \5620_b0 );
or ( \5622_b1 , \5610_b1 , w_17908 );
or ( \5622_b0 , \5610_b0 , \5621_b0 );
not ( \5621_b0 , w_17909 );
and ( w_17909 , w_17908 , \5621_b1 );
or ( \5623_b1 , \5599_b1 , w_17911 );
not ( w_17911 , w_17912 );
and ( \5623_b0 , \5599_b0 , w_17913 );
and ( w_17912 ,  , w_17913 );
buf ( w_17911 , \5609_b1 );
not ( w_17911 , w_17914 );
not (  , w_17915 );
and ( w_17914 , w_17915 , \5609_b0 );
or ( \5624_b1 , \5622_b1 , w_17917 );
not ( w_17917 , w_17918 );
and ( \5624_b0 , \5622_b0 , w_17919 );
and ( w_17918 ,  , w_17919 );
buf ( w_17917 , \5623_b1 );
not ( w_17917 , w_17920 );
not (  , w_17921 );
and ( w_17920 , w_17921 , \5623_b0 );
or ( \5625_b1 , \5589_b1 , \5624_b1 );
not ( \5624_b1 , w_17922 );
and ( \5625_b0 , \5589_b0 , w_17923 );
and ( w_17922 , w_17923 , \5624_b0 );
or ( \5626_b1 , \5586_b1 , \5588_b1 );
not ( \5588_b1 , w_17924 );
and ( \5626_b0 , \5586_b0 , w_17925 );
and ( w_17924 , w_17925 , \5588_b0 );
or ( \5627_b1 , \5625_b1 , w_17926 );
or ( \5627_b0 , \5625_b0 , \5626_b0 );
not ( \5626_b0 , w_17927 );
and ( w_17927 , w_17926 , \5626_b1 );
or ( \5628_b1 , \5414_b1 , \5449_b1 );
xor ( \5628_b0 , \5414_b0 , w_17928 );
not ( w_17928 , w_17929 );
and ( w_17929 , \5449_b1 , \5449_b0 );
or ( \5629_b1 , \5628_b1 , \5476_b1 );
xor ( \5629_b0 , \5628_b0 , w_17930 );
not ( w_17930 , w_17931 );
and ( w_17931 , \5476_b1 , \5476_b0 );
or ( \5630_b1 , \5627_b1 , \5629_b1 );
xor ( \5630_b0 , \5627_b0 , w_17932 );
not ( w_17932 , w_17933 );
and ( w_17933 , \5629_b1 , \5629_b0 );
or ( \5631_b1 , \5424_b1 , \5435_b1 );
xor ( \5631_b0 , \5424_b0 , w_17934 );
not ( w_17934 , w_17935 );
and ( w_17935 , \5435_b1 , \5435_b0 );
or ( \5632_b1 , \5631_b1 , \5446_b1 );
xor ( \5632_b0 , \5631_b0 , w_17936 );
not ( w_17936 , w_17937 );
and ( w_17937 , \5446_b1 , \5446_b0 );
or ( \5633_b1 , \5455_b1 , \5462_b1 );
xor ( \5633_b0 , \5455_b0 , w_17938 );
not ( w_17938 , w_17939 );
and ( w_17939 , \5462_b1 , \5462_b0 );
or ( \5634_b1 , \5633_b1 , \5473_b1 );
xor ( \5634_b0 , \5633_b0 , w_17940 );
not ( w_17940 , w_17941 );
and ( w_17941 , \5473_b1 , \5473_b0 );
or ( \5635_b1 , \5632_b1 , \5634_b1 );
xor ( \5635_b0 , \5632_b0 , w_17942 );
not ( w_17942 , w_17943 );
and ( w_17943 , \5634_b1 , \5634_b0 );
buf ( \5636_b1 , \4041_b1 );
not ( \5636_b1 , w_17944 );
not ( \5636_b0 , w_17945 );
and ( w_17944 , w_17945 , \4041_b0 );
buf ( \5637_b1 , \4069_b1 );
not ( \5637_b1 , w_17946 );
not ( \5637_b0 , w_17947 );
and ( w_17946 , w_17947 , \4069_b0 );
or ( \5638_b1 , \5636_b1 , w_17948 );
or ( \5638_b0 , \5636_b0 , \5637_b0 );
not ( \5637_b0 , w_17949 );
and ( w_17949 , w_17948 , \5637_b1 );
or ( \5639_b1 , \5060_b1 , w_17951 );
not ( w_17951 , w_17952 );
and ( \5639_b0 , \5060_b0 , w_17953 );
and ( w_17952 ,  , w_17953 );
buf ( w_17951 , \4238_b1 );
not ( w_17951 , w_17954 );
not (  , w_17955 );
and ( w_17954 , w_17955 , \4238_b0 );
or ( \5640_b1 , \5638_b1 , w_17957 );
not ( w_17957 , w_17958 );
and ( \5640_b0 , \5638_b0 , w_17959 );
and ( w_17958 ,  , w_17959 );
buf ( w_17957 , \5639_b1 );
not ( w_17957 , w_17960 );
not (  , w_17961 );
and ( w_17960 , w_17961 , \5639_b0 );
buf ( \5641_b1 , \5640_b1 );
not ( \5641_b1 , w_17962 );
not ( \5641_b0 , w_17963 );
and ( w_17962 , w_17963 , \5640_b0 );
buf ( \5642_b1 , \4065_b1 );
not ( \5642_b1 , w_17964 );
not ( \5642_b0 , w_17965 );
and ( w_17964 , w_17965 , \4065_b0 );
or ( \5643_b1 , \5641_b1 , w_17966 );
or ( \5643_b0 , \5641_b0 , \5642_b0 );
not ( \5642_b0 , w_17967 );
and ( w_17967 , w_17966 , \5642_b1 );
or ( \5644_b1 , \5422_b1 , w_17969 );
not ( w_17969 , w_17970 );
and ( \5644_b0 , \5422_b0 , w_17971 );
and ( w_17970 ,  , w_17971 );
buf ( w_17969 , \4055_b1 );
not ( w_17969 , w_17972 );
not (  , w_17973 );
and ( w_17972 , w_17973 , \4055_b0 );
or ( \5645_b1 , \5643_b1 , w_17975 );
not ( w_17975 , w_17976 );
and ( \5645_b0 , \5643_b0 , w_17977 );
and ( w_17976 ,  , w_17977 );
buf ( w_17975 , \5644_b1 );
not ( w_17975 , w_17978 );
not (  , w_17979 );
and ( w_17978 , w_17979 , \5644_b0 );
buf ( \5646_b1 , \4585_b1 );
not ( \5646_b1 , w_17980 );
not ( \5646_b0 , w_17981 );
and ( w_17980 , w_17981 , \4585_b0 );
buf ( \5647_b1 , \4171_b1 );
not ( \5647_b1 , w_17982 );
not ( \5647_b0 , w_17983 );
and ( w_17982 , w_17983 , \4171_b0 );
or ( \5648_b1 , \5646_b1 , w_17984 );
or ( \5648_b0 , \5646_b0 , \5647_b0 );
not ( \5647_b0 , w_17985 );
and ( w_17985 , w_17984 , \5647_b1 );
or ( \5649_b1 , \4284_b1 , w_17987 );
not ( w_17987 , w_17988 );
and ( \5649_b0 , \4284_b0 , w_17989 );
and ( w_17988 ,  , w_17989 );
buf ( w_17987 , \4019_b1 );
not ( w_17987 , w_17990 );
not (  , w_17991 );
and ( w_17990 , w_17991 , \4019_b0 );
or ( \5650_b1 , \5648_b1 , w_17993 );
not ( w_17993 , w_17994 );
and ( \5650_b0 , \5648_b0 , w_17995 );
and ( w_17994 ,  , w_17995 );
buf ( w_17993 , \5649_b1 );
not ( w_17993 , w_17996 );
not (  , w_17997 );
and ( w_17996 , w_17997 , \5649_b0 );
buf ( \5651_b1 , \5650_b1 );
not ( \5651_b1 , w_17998 );
not ( \5651_b0 , w_17999 );
and ( w_17998 , w_17999 , \5650_b0 );
buf ( \5652_b1 , \4194_b1 );
not ( \5652_b1 , w_18000 );
not ( \5652_b0 , w_18001 );
and ( w_18000 , w_18001 , \4194_b0 );
or ( \5653_b1 , \5651_b1 , w_18002 );
or ( \5653_b0 , \5651_b0 , \5652_b0 );
not ( \5652_b0 , w_18003 );
and ( w_18003 , w_18002 , \5652_b1 );
or ( \5654_b1 , \5111_b1 , w_18005 );
not ( w_18005 , w_18006 );
and ( \5654_b0 , \5111_b0 , w_18007 );
and ( w_18006 ,  , w_18007 );
buf ( w_18005 , \5468_b1 );
not ( w_18005 , w_18008 );
not (  , w_18009 );
and ( w_18008 , w_18009 , \5468_b0 );
or ( \5655_b1 , \5653_b1 , w_18011 );
not ( w_18011 , w_18012 );
and ( \5655_b0 , \5653_b0 , w_18013 );
and ( w_18012 ,  , w_18013 );
buf ( w_18011 , \5654_b1 );
not ( w_18011 , w_18014 );
not (  , w_18015 );
and ( w_18014 , w_18015 , \5654_b0 );
or ( \5656_b1 , \5645_b1 , \5655_b1 );
xor ( \5656_b0 , \5645_b0 , w_18016 );
not ( w_18016 , w_18017 );
and ( w_18017 , \5655_b1 , \5655_b0 );
or ( \5657_b1 , \5388_b1 , \4267_b1 );
not ( \4267_b1 , w_18018 );
and ( \5657_b0 , \5388_b0 , w_18019 );
and ( w_18018 , w_18019 , \4267_b0 );
buf ( \5658_b1 , \5388_b1 );
not ( \5658_b1 , w_18020 );
not ( \5658_b0 , w_18021 );
and ( w_18020 , w_18021 , \5388_b0 );
or ( \5659_b1 , \5658_b1 , \4156_b1 );
not ( \4156_b1 , w_18022 );
and ( \5659_b0 , \5658_b0 , w_18023 );
and ( w_18022 , w_18023 , \4156_b0 );
or ( \5660_b1 , \5657_b1 , w_18025 );
not ( w_18025 , w_18026 );
and ( \5660_b0 , \5657_b0 , w_18027 );
and ( w_18026 ,  , w_18027 );
buf ( w_18025 , \5659_b1 );
not ( w_18025 , w_18028 );
not (  , w_18029 );
and ( w_18028 , w_18029 , \5659_b0 );
buf ( \5661_b1 , \5660_b1 );
not ( \5661_b1 , w_18030 );
not ( \5661_b0 , w_18031 );
and ( w_18030 , w_18031 , \5660_b0 );
buf ( \5662_b1 , \4253_b1 );
not ( \5662_b1 , w_18032 );
not ( \5662_b0 , w_18033 );
and ( w_18032 , w_18033 , \4253_b0 );
or ( \5663_b1 , \5661_b1 , w_18034 );
or ( \5663_b0 , \5661_b0 , \5662_b0 );
not ( \5662_b0 , w_18035 );
and ( w_18035 , w_18034 , \5662_b1 );
or ( \5664_b1 , \4273_b1 , w_18037 );
not ( w_18037 , w_18038 );
and ( \5664_b0 , \4273_b0 , w_18039 );
and ( w_18038 ,  , w_18039 );
buf ( w_18037 , \5460_b1 );
not ( w_18037 , w_18040 );
not (  , w_18041 );
and ( w_18040 , w_18041 , \5460_b0 );
or ( \5665_b1 , \5663_b1 , w_18043 );
not ( w_18043 , w_18044 );
and ( \5665_b0 , \5663_b0 , w_18045 );
and ( w_18044 ,  , w_18045 );
buf ( w_18043 , \5664_b1 );
not ( w_18043 , w_18046 );
not (  , w_18047 );
and ( w_18046 , w_18047 , \5664_b0 );
or ( \5666_b1 , \5656_b1 , \5665_b1 );
not ( \5665_b1 , w_18048 );
and ( \5666_b0 , \5656_b0 , w_18049 );
and ( w_18048 , w_18049 , \5665_b0 );
or ( \5667_b1 , \5645_b1 , \5655_b1 );
not ( \5655_b1 , w_18050 );
and ( \5667_b0 , \5645_b0 , w_18051 );
and ( w_18050 , w_18051 , \5655_b0 );
or ( \5668_b1 , \5666_b1 , w_18052 );
or ( \5668_b0 , \5666_b0 , \5667_b0 );
not ( \5667_b0 , w_18053 );
and ( w_18053 , w_18052 , \5667_b1 );
or ( \5669_b1 , \5635_b1 , \5668_b1 );
not ( \5668_b1 , w_18054 );
and ( \5669_b0 , \5635_b0 , w_18055 );
and ( w_18054 , w_18055 , \5668_b0 );
or ( \5670_b1 , \5632_b1 , \5634_b1 );
not ( \5634_b1 , w_18056 );
and ( \5670_b0 , \5632_b0 , w_18057 );
and ( w_18056 , w_18057 , \5634_b0 );
or ( \5671_b1 , \5669_b1 , w_18058 );
or ( \5671_b0 , \5669_b0 , \5670_b0 );
not ( \5670_b0 , w_18059 );
and ( w_18059 , w_18058 , \5670_b1 );
or ( \5672_b1 , \5630_b1 , \5671_b1 );
not ( \5671_b1 , w_18060 );
and ( \5672_b0 , \5630_b0 , w_18061 );
and ( w_18060 , w_18061 , \5671_b0 );
or ( \5673_b1 , \5627_b1 , \5629_b1 );
not ( \5629_b1 , w_18062 );
and ( \5673_b0 , \5627_b0 , w_18063 );
and ( w_18062 , w_18063 , \5629_b0 );
or ( \5674_b1 , \5672_b1 , w_18064 );
or ( \5674_b0 , \5672_b0 , \5673_b0 );
not ( \5673_b0 , w_18065 );
and ( w_18065 , w_18064 , \5673_b1 );
buf ( \5675_b1 , \5674_b1 );
not ( \5675_b1 , w_18066 );
not ( \5675_b0 , w_18067 );
and ( w_18066 , w_18067 , \5674_b0 );
or ( \5676_b1 , \5568_b1 , \5675_b1 );
xor ( \5676_b0 , \5568_b0 , w_18068 );
not ( w_18068 , w_18069 );
and ( w_18069 , \5675_b1 , \5675_b0 );
or ( \5677_b1 , \5479_b1 , \5494_b1 );
xor ( \5677_b0 , \5479_b0 , w_18070 );
not ( w_18070 , w_18071 );
and ( w_18071 , \5494_b1 , \5494_b0 );
or ( \5678_b1 , \5677_b1 , w_18072 );
xor ( \5678_b0 , \5677_b0 , w_18074 );
not ( w_18074 , w_18075 );
and ( w_18075 , w_18072 , w_18073 );
buf ( w_18072 , \5499_b1 );
not ( w_18072 , w_18076 );
not ( w_18073 , w_18077 );
and ( w_18076 , w_18077 , \5499_b0 );
or ( \5679_b1 , \5676_b1 , \5678_b1 );
not ( \5678_b1 , w_18078 );
and ( \5679_b0 , \5676_b0 , w_18079 );
and ( w_18078 , w_18079 , \5678_b0 );
or ( \5680_b1 , \5568_b1 , \5675_b1 );
not ( \5675_b1 , w_18080 );
and ( \5680_b0 , \5568_b0 , w_18081 );
and ( w_18080 , w_18081 , \5675_b0 );
or ( \5681_b1 , \5679_b1 , w_18082 );
or ( \5681_b0 , \5679_b0 , \5680_b0 );
not ( \5680_b0 , w_18083 );
and ( w_18083 , w_18082 , \5680_b1 );
or ( \5682_b1 , \5563_b1 , w_18085 );
not ( w_18085 , w_18086 );
and ( \5682_b0 , \5563_b0 , w_18087 );
and ( w_18086 ,  , w_18087 );
buf ( w_18085 , \5681_b1 );
not ( w_18085 , w_18088 );
not (  , w_18089 );
and ( w_18088 , w_18089 , \5681_b0 );
or ( \5683_b1 , \5568_b1 , \5675_b1 );
xor ( \5683_b0 , \5568_b0 , w_18090 );
not ( w_18090 , w_18091 );
and ( w_18091 , \5675_b1 , \5675_b0 );
or ( \5684_b1 , \5683_b1 , \5678_b1 );
xor ( \5684_b0 , \5683_b0 , w_18092 );
not ( w_18092 , w_18093 );
and ( w_18093 , \5678_b1 , \5678_b0 );
or ( \5685_b1 , \5627_b1 , \5629_b1 );
xor ( \5685_b0 , \5627_b0 , w_18094 );
not ( w_18094 , w_18095 );
and ( w_18095 , \5629_b1 , \5629_b0 );
or ( \5686_b1 , \5685_b1 , \5671_b1 );
xor ( \5686_b0 , \5685_b0 , w_18096 );
not ( w_18096 , w_18097 );
and ( w_18097 , \5671_b1 , \5671_b0 );
buf ( \5687_b1 , \5686_b1 );
buf ( \5687_b0 , \5686_b0 );
buf ( \5688_b1 , \5687_b1 );
not ( \5688_b1 , w_18098 );
not ( \5688_b0 , w_18099 );
and ( w_18098 , w_18099 , \5687_b0 );
or ( \5689_b1 , \5486_b1 , \5492_b1 );
xor ( \5689_b0 , \5486_b0 , w_18100 );
not ( w_18100 , w_18101 );
and ( w_18101 , \5492_b1 , \5492_b0 );
or ( \5690_b1 , \5689_b1 , \5483_b1 );
xor ( \5690_b0 , \5689_b0 , w_18102 );
not ( w_18102 , w_18103 );
and ( w_18103 , \5483_b1 , \5483_b0 );
buf ( \5691_b1 , \5690_b1 );
buf ( \5691_b0 , \5690_b0 );
or ( \5692_b1 , \5688_b1 , w_18105 );
not ( w_18105 , w_18106 );
and ( \5692_b0 , \5688_b0 , w_18107 );
and ( w_18106 ,  , w_18107 );
buf ( w_18105 , \5691_b1 );
not ( w_18105 , w_18108 );
not (  , w_18109 );
and ( w_18108 , w_18109 , \5691_b0 );
or ( \5693_b1 , \5344_b1 , \4492_b1 );
xor ( \5693_b0 , \5344_b0 , w_18110 );
not ( w_18110 , w_18111 );
and ( w_18111 , \4492_b1 , \4492_b0 );
buf ( \5694_b1 , \5693_b1 );
not ( \5694_b1 , w_18112 );
not ( \5694_b0 , w_18113 );
and ( w_18112 , w_18113 , \5693_b0 );
buf ( \5695_b1 , \5694_b1 );
not ( \5695_b1 , w_18114 );
not ( \5695_b0 , w_18115 );
and ( w_18114 , w_18115 , \5694_b0 );
buf ( \5696_b1 , \4231_b1 );
not ( \5696_b1 , w_18116 );
not ( \5696_b0 , w_18117 );
and ( w_18116 , w_18117 , \4231_b0 );
or ( \5697_b1 , \5695_b1 , w_18118 );
or ( \5697_b0 , \5695_b0 , \5696_b0 );
not ( \5696_b0 , w_18119 );
and ( w_18119 , w_18118 , \5696_b1 );
or ( \5698_b1 , \4234_b1 , w_18121 );
not ( w_18121 , w_18122 );
and ( \5698_b0 , \4234_b0 , w_18123 );
and ( w_18122 ,  , w_18123 );
buf ( w_18121 , \5451_b1 );
not ( w_18121 , w_18124 );
not (  , w_18125 );
and ( w_18124 , w_18125 , \5451_b0 );
or ( \5699_b1 , \5697_b1 , w_18127 );
not ( w_18127 , w_18128 );
and ( \5699_b0 , \5697_b0 , w_18129 );
and ( w_18128 ,  , w_18129 );
buf ( w_18127 , \5698_b1 );
not ( w_18127 , w_18130 );
not (  , w_18131 );
and ( w_18130 , w_18131 , \5698_b0 );
or ( \5700_b1 , \5574_b1 , \5585_b1 );
xor ( \5700_b0 , \5574_b0 , w_18132 );
not ( w_18132 , w_18133 );
and ( w_18133 , \5585_b1 , \5585_b0 );
or ( \5701_b1 , \5699_b1 , \5700_b1 );
xor ( \5701_b0 , \5699_b0 , w_18134 );
not ( w_18134 , w_18135 );
and ( w_18135 , \5700_b1 , \5700_b0 );
buf ( \5702_b1 , \4042_b1 );
not ( \5702_b1 , w_18136 );
not ( \5702_b0 , w_18137 );
and ( w_18136 , w_18137 , \4042_b0 );
buf ( \5703_b1 , \5270_b1 );
not ( \5703_b1 , w_18138 );
not ( \5703_b0 , w_18139 );
and ( w_18138 , w_18139 , \5270_b0 );
or ( \5704_b1 , \5702_b1 , w_18140 );
or ( \5704_b0 , \5702_b0 , \5703_b0 );
not ( \5703_b0 , w_18141 );
and ( w_18141 , w_18140 , \5703_b1 );
or ( \5705_b1 , \5273_b1 , w_18143 );
not ( w_18143 , w_18144 );
and ( \5705_b0 , \5273_b0 , w_18145 );
and ( w_18144 ,  , w_18145 );
buf ( w_18143 , \4116_b1 );
not ( w_18143 , w_18146 );
not (  , w_18147 );
and ( w_18146 , w_18147 , \4116_b0 );
or ( \5706_b1 , \5704_b1 , w_18149 );
not ( w_18149 , w_18150 );
and ( \5706_b0 , \5704_b0 , w_18151 );
and ( w_18150 ,  , w_18151 );
buf ( w_18149 , \5705_b1 );
not ( w_18149 , w_18152 );
not (  , w_18153 );
and ( w_18152 , w_18153 , \5705_b0 );
or ( \5707_b1 , \5019_b1 , \5706_b1 );
not ( \5706_b1 , w_18154 );
and ( \5707_b0 , \5019_b0 , w_18155 );
and ( w_18154 , w_18155 , \5706_b0 );
or ( \5708_b1 , \5580_b1 , \5021_b1 );
not ( \5021_b1 , w_18156 );
and ( \5708_b0 , \5580_b0 , w_18157 );
and ( w_18156 , w_18157 , \5021_b0 );
or ( \5709_b1 , \5707_b1 , w_18159 );
not ( w_18159 , w_18160 );
and ( \5709_b0 , \5707_b0 , w_18161 );
and ( w_18160 ,  , w_18161 );
buf ( w_18159 , \5708_b1 );
not ( w_18159 , w_18162 );
not (  , w_18163 );
and ( w_18162 , w_18163 , \5708_b0 );
buf ( \5710_b1 , \5709_b1 );
not ( \5710_b1 , w_18164 );
not ( \5710_b0 , w_18165 );
and ( w_18164 , w_18165 , \5709_b0 );
buf ( \5711_b1 , \5710_b1 );
not ( \5711_b1 , w_18166 );
not ( \5711_b0 , w_18167 );
and ( w_18166 , w_18167 , \5710_b0 );
buf ( \5712_b1 , \4252_b1 );
not ( \5712_b1 , w_18168 );
not ( \5712_b0 , w_18169 );
and ( w_18168 , w_18169 , \4252_b0 );
or ( \5713_b1 , \5712_b1 , w_18171 );
not ( w_18171 , w_18172 );
and ( \5713_b0 , \5712_b0 , w_18173 );
and ( w_18172 ,  , w_18173 );
buf ( w_18171 , \4048_b1 );
not ( w_18171 , w_18174 );
not (  , w_18175 );
and ( w_18174 , w_18175 , \4048_b0 );
buf ( \5714_b1 , \5713_b1 );
not ( \5714_b1 , w_18176 );
not ( \5714_b0 , w_18177 );
and ( w_18176 , w_18177 , \5713_b0 );
buf ( \5715_b1 , \5714_b1 );
not ( \5715_b1 , w_18178 );
not ( \5715_b0 , w_18179 );
and ( w_18178 , w_18179 , \5714_b0 );
or ( \5716_b1 , \5711_b1 , w_18180 );
or ( \5716_b0 , \5711_b0 , \5715_b0 );
not ( \5715_b0 , w_18181 );
and ( w_18181 , w_18180 , \5715_b1 );
buf ( \5717_b1 , \4045_b1 );
not ( \5717_b1 , w_18182 );
not ( \5717_b0 , w_18183 );
and ( w_18182 , w_18183 , \4045_b0 );
buf ( \5718_b1 , \5178_b1 );
not ( \5718_b1 , w_18184 );
not ( \5718_b0 , w_18185 );
and ( w_18184 , w_18185 , \5178_b0 );
or ( \5719_b1 , \5717_b1 , w_18186 );
or ( \5719_b0 , \5717_b0 , \5718_b0 );
not ( \5718_b0 , w_18187 );
and ( w_18187 , w_18186 , \5718_b1 );
or ( \5720_b1 , \4665_b1 , w_18189 );
not ( w_18189 , w_18190 );
and ( \5720_b0 , \4665_b0 , w_18191 );
and ( w_18190 ,  , w_18191 );
buf ( w_18189 , \4286_b1 );
not ( w_18189 , w_18192 );
not (  , w_18193 );
and ( w_18192 , w_18193 , \4286_b0 );
or ( \5721_b1 , \5719_b1 , w_18195 );
not ( w_18195 , w_18196 );
and ( \5721_b0 , \5719_b0 , w_18197 );
and ( w_18196 ,  , w_18197 );
buf ( w_18195 , \5720_b1 );
not ( w_18195 , w_18198 );
not (  , w_18199 );
and ( w_18198 , w_18199 , \5720_b0 );
buf ( \5722_b1 , \5721_b1 );
not ( \5722_b1 , w_18200 );
not ( \5722_b0 , w_18201 );
and ( w_18200 , w_18201 , \5721_b0 );
buf ( \5723_b1 , \4662_b1 );
not ( \5723_b1 , w_18202 );
not ( \5723_b0 , w_18203 );
and ( w_18202 , w_18203 , \4662_b0 );
or ( \5724_b1 , \5722_b1 , w_18204 );
or ( \5724_b0 , \5722_b0 , \5723_b0 );
not ( \5723_b0 , w_18205 );
and ( w_18205 , w_18204 , \5723_b1 );
or ( \5725_b1 , \4672_b1 , w_18207 );
not ( w_18207 , w_18208 );
and ( \5725_b0 , \4672_b0 , w_18209 );
and ( w_18208 ,  , w_18209 );
buf ( w_18207 , \5615_b1 );
not ( w_18207 , w_18210 );
not (  , w_18211 );
and ( w_18210 , w_18211 , \5615_b0 );
or ( \5726_b1 , \5724_b1 , w_18213 );
not ( w_18213 , w_18214 );
and ( \5726_b0 , \5724_b0 , w_18215 );
and ( w_18214 ,  , w_18215 );
buf ( w_18213 , \5725_b1 );
not ( w_18213 , w_18216 );
not (  , w_18217 );
and ( w_18216 , w_18217 , \5725_b0 );
or ( \5727_b1 , \5713_b1 , w_18219 );
not ( w_18219 , w_18220 );
and ( \5727_b0 , \5713_b0 , w_18221 );
and ( w_18220 ,  , w_18221 );
buf ( w_18219 , \5709_b1 );
not ( w_18219 , w_18222 );
not (  , w_18223 );
and ( w_18222 , w_18223 , \5709_b0 );
or ( \5728_b1 , \5726_b1 , w_18225 );
not ( w_18225 , w_18226 );
and ( \5728_b0 , \5726_b0 , w_18227 );
and ( w_18226 ,  , w_18227 );
buf ( w_18225 , \5727_b1 );
not ( w_18225 , w_18228 );
not (  , w_18229 );
and ( w_18228 , w_18229 , \5727_b0 );
or ( \5729_b1 , \5716_b1 , w_18231 );
not ( w_18231 , w_18232 );
and ( \5729_b0 , \5716_b0 , w_18233 );
and ( w_18232 ,  , w_18233 );
buf ( w_18231 , \5728_b1 );
not ( w_18231 , w_18234 );
not (  , w_18235 );
and ( w_18234 , w_18235 , \5728_b0 );
or ( \5730_b1 , \5701_b1 , \5729_b1 );
not ( \5729_b1 , w_18236 );
and ( \5730_b0 , \5701_b0 , w_18237 );
and ( w_18236 , w_18237 , \5729_b0 );
or ( \5731_b1 , \5699_b1 , \5700_b1 );
not ( \5700_b1 , w_18238 );
and ( \5731_b0 , \5699_b0 , w_18239 );
and ( w_18238 , w_18239 , \5700_b0 );
or ( \5732_b1 , \5730_b1 , w_18240 );
or ( \5732_b0 , \5730_b0 , \5731_b0 );
not ( \5731_b0 , w_18241 );
and ( w_18241 , w_18240 , \5731_b1 );
or ( \5733_b1 , \5586_b1 , \5588_b1 );
xor ( \5733_b0 , \5586_b0 , w_18242 );
not ( w_18242 , w_18243 );
and ( w_18243 , \5588_b1 , \5588_b0 );
or ( \5734_b1 , \5733_b1 , \5624_b1 );
xor ( \5734_b0 , \5733_b0 , w_18244 );
not ( w_18244 , w_18245 );
and ( w_18245 , \5624_b1 , \5624_b0 );
or ( \5735_b1 , \5732_b1 , \5734_b1 );
xor ( \5735_b0 , \5732_b0 , w_18246 );
not ( w_18246 , w_18247 );
and ( w_18247 , \5734_b1 , \5734_b0 );
or ( \5736_b1 , \5632_b1 , \5634_b1 );
xor ( \5736_b0 , \5632_b0 , w_18248 );
not ( w_18248 , w_18249 );
and ( w_18249 , \5634_b1 , \5634_b0 );
or ( \5737_b1 , \5736_b1 , \5668_b1 );
xor ( \5737_b0 , \5736_b0 , w_18250 );
not ( w_18250 , w_18251 );
and ( w_18251 , \5668_b1 , \5668_b0 );
or ( \5738_b1 , \5735_b1 , \5737_b1 );
not ( \5737_b1 , w_18252 );
and ( \5738_b0 , \5735_b0 , w_18253 );
and ( w_18252 , w_18253 , \5737_b0 );
or ( \5739_b1 , \5732_b1 , \5734_b1 );
not ( \5734_b1 , w_18254 );
and ( \5739_b0 , \5732_b0 , w_18255 );
and ( w_18254 , w_18255 , \5734_b0 );
or ( \5740_b1 , \5738_b1 , w_18256 );
or ( \5740_b0 , \5738_b0 , \5739_b0 );
not ( \5739_b0 , w_18257 );
and ( w_18257 , w_18256 , \5739_b1 );
or ( \5741_b1 , \5692_b1 , \5740_b1 );
not ( \5740_b1 , w_18258 );
and ( \5741_b0 , \5692_b0 , w_18259 );
and ( w_18258 , w_18259 , \5740_b0 );
or ( \5742_b1 , \5688_b1 , w_18261 );
not ( w_18261 , w_18262 );
and ( \5742_b0 , \5688_b0 , w_18263 );
and ( w_18262 ,  , w_18263 );
buf ( w_18261 , \5691_b1 );
not ( w_18261 , w_18264 );
not (  , w_18265 );
and ( w_18264 , w_18265 , \5691_b0 );
or ( \5743_b1 , \5741_b1 , w_18267 );
not ( w_18267 , w_18268 );
and ( \5743_b0 , \5741_b0 , w_18269 );
and ( w_18268 ,  , w_18269 );
buf ( w_18267 , \5742_b1 );
not ( w_18267 , w_18270 );
not (  , w_18271 );
and ( w_18270 , w_18271 , \5742_b0 );
or ( \5744_b1 , \5684_b1 , w_18273 );
not ( w_18273 , w_18274 );
and ( \5744_b0 , \5684_b0 , w_18275 );
and ( w_18274 ,  , w_18275 );
buf ( w_18273 , \5743_b1 );
not ( w_18273 , w_18276 );
not (  , w_18277 );
and ( w_18276 , w_18277 , \5743_b0 );
or ( \5745_b1 , \5682_b1 , \5744_b1 );
not ( \5744_b1 , w_18278 );
and ( \5745_b0 , \5682_b0 , w_18279 );
and ( w_18278 , w_18279 , \5744_b0 );
buf ( \5746_b1 , \4011_b1 );
not ( \5746_b1 , w_18280 );
not ( \5746_b0 , w_18281 );
and ( w_18280 , w_18281 , \4011_b0 );
buf ( \5747_b1 , \4404_b1 );
not ( \5747_b1 , w_18282 );
not ( \5747_b0 , w_18283 );
and ( w_18282 , w_18283 , \4404_b0 );
or ( \5748_b1 , \5746_b1 , w_18284 );
or ( \5748_b0 , \5746_b0 , \5747_b0 );
not ( \5747_b0 , w_18285 );
and ( w_18285 , w_18284 , \5747_b1 );
buf ( \5749_b1 , \4069_b1 );
not ( \5749_b1 , w_18286 );
not ( \5749_b0 , w_18287 );
and ( w_18286 , w_18287 , \4069_b0 );
or ( \5750_b1 , \5749_b1 , w_18289 );
not ( w_18289 , w_18290 );
and ( \5750_b0 , \5749_b0 , w_18291 );
and ( w_18290 ,  , w_18291 );
buf ( w_18289 , \4270_b1 );
not ( w_18289 , w_18292 );
not (  , w_18293 );
and ( w_18292 , w_18293 , \4270_b0 );
or ( \5751_b1 , \5748_b1 , w_18295 );
not ( w_18295 , w_18296 );
and ( \5751_b0 , \5748_b0 , w_18297 );
and ( w_18296 ,  , w_18297 );
buf ( w_18295 , \5750_b1 );
not ( w_18295 , w_18298 );
not (  , w_18299 );
and ( w_18298 , w_18299 , \5750_b0 );
buf ( \5752_b1 , \5751_b1 );
not ( \5752_b1 , w_18300 );
not ( \5752_b0 , w_18301 );
and ( w_18300 , w_18301 , \5751_b0 );
buf ( \5753_b1 , \4558_b1 );
not ( \5753_b1 , w_18302 );
not ( \5753_b0 , w_18303 );
and ( w_18302 , w_18303 , \4558_b0 );
or ( \5754_b1 , \5752_b1 , w_18304 );
or ( \5754_b0 , \5752_b0 , \5753_b0 );
not ( \5753_b0 , w_18305 );
and ( w_18305 , w_18304 , \5753_b1 );
buf ( \5755_b1 , \4043_b1 );
not ( \5755_b1 , w_18306 );
not ( \5755_b0 , w_18307 );
and ( w_18306 , w_18307 , \4043_b0 );
buf ( \5756_b1 , \4069_b1 );
not ( \5756_b1 , w_18308 );
not ( \5756_b0 , w_18309 );
and ( w_18308 , w_18309 , \4069_b0 );
or ( \5757_b1 , \5755_b1 , w_18310 );
or ( \5757_b0 , \5755_b0 , \5756_b0 );
not ( \5756_b0 , w_18311 );
and ( w_18311 , w_18310 , \5756_b1 );
or ( \5758_b1 , \5749_b1 , w_18313 );
not ( w_18313 , w_18314 );
and ( \5758_b0 , \5749_b0 , w_18315 );
and ( w_18314 ,  , w_18315 );
buf ( w_18313 , \4217_b1 );
not ( w_18313 , w_18316 );
not (  , w_18317 );
and ( w_18316 , w_18317 , \4217_b0 );
or ( \5759_b1 , \5757_b1 , w_18319 );
not ( w_18319 , w_18320 );
and ( \5759_b0 , \5757_b0 , w_18321 );
and ( w_18320 ,  , w_18321 );
buf ( w_18319 , \5758_b1 );
not ( w_18319 , w_18322 );
not (  , w_18323 );
and ( w_18322 , w_18323 , \5758_b0 );
or ( \5760_b1 , \4562_b1 , w_18325 );
not ( w_18325 , w_18326 );
and ( \5760_b0 , \4562_b0 , w_18327 );
and ( w_18326 ,  , w_18327 );
buf ( w_18325 , \5759_b1 );
not ( w_18325 , w_18328 );
not (  , w_18329 );
and ( w_18328 , w_18329 , \5759_b0 );
or ( \5761_b1 , \5754_b1 , w_18331 );
not ( w_18331 , w_18332 );
and ( \5761_b0 , \5754_b0 , w_18333 );
and ( w_18332 ,  , w_18333 );
buf ( w_18331 , \5760_b1 );
not ( w_18331 , w_18334 );
not (  , w_18335 );
and ( w_18334 , w_18335 , \5760_b0 );
buf ( \5762_b1 , \4048_b1 );
not ( \5762_b1 , w_18336 );
not ( \5762_b0 , w_18337 );
and ( w_18336 , w_18337 , \4048_b0 );
buf ( \5763_b1 , \4212_b1 );
not ( \5763_b1 , w_18338 );
not ( \5763_b0 , w_18339 );
and ( w_18338 , w_18339 , \4212_b0 );
or ( \5764_b1 , \5762_b1 , w_18340 );
or ( \5764_b0 , \5762_b0 , \5763_b0 );
not ( \5763_b0 , w_18341 );
and ( w_18341 , w_18340 , \5763_b1 );
or ( \5765_b1 , \4492_b1 , w_18343 );
not ( w_18343 , w_18344 );
and ( \5765_b0 , \4492_b0 , w_18345 );
and ( w_18344 ,  , w_18345 );
buf ( w_18343 , \5388_b1 );
not ( w_18343 , w_18346 );
not (  , w_18347 );
and ( w_18346 , w_18347 , \5388_b0 );
or ( \5766_b1 , \5764_b1 , w_18349 );
not ( w_18349 , w_18350 );
and ( \5766_b0 , \5764_b0 , w_18351 );
and ( w_18350 ,  , w_18351 );
buf ( w_18349 , \5765_b1 );
not ( w_18349 , w_18352 );
not (  , w_18353 );
and ( w_18352 , w_18353 , \5765_b0 );
buf ( \5767_b1 , \5766_b1 );
not ( \5767_b1 , w_18354 );
not ( \5767_b0 , w_18355 );
and ( w_18354 , w_18355 , \5766_b0 );
buf ( \5768_b1 , \4231_b1 );
not ( \5768_b1 , w_18356 );
not ( \5768_b0 , w_18357 );
and ( w_18356 , w_18357 , \4231_b0 );
or ( \5769_b1 , \5767_b1 , w_18358 );
or ( \5769_b0 , \5767_b0 , \5768_b0 );
not ( \5768_b0 , w_18359 );
and ( w_18359 , w_18358 , \5768_b1 );
buf ( \5770_b1 , \4029_b1 );
not ( \5770_b1 , w_18360 );
not ( \5770_b0 , w_18361 );
and ( w_18360 , w_18361 , \4029_b0 );
buf ( \5771_b1 , \4212_b1 );
not ( \5771_b1 , w_18362 );
not ( \5771_b0 , w_18363 );
and ( w_18362 , w_18363 , \4212_b0 );
or ( \5772_b1 , \5770_b1 , w_18364 );
or ( \5772_b0 , \5770_b0 , \5771_b0 );
not ( \5771_b0 , w_18365 );
and ( w_18365 , w_18364 , \5771_b1 );
or ( \5773_b1 , \4492_b1 , w_18367 );
not ( w_18367 , w_18368 );
and ( \5773_b0 , \4492_b0 , w_18369 );
and ( w_18368 ,  , w_18369 );
buf ( w_18367 , \5339_b1 );
not ( w_18367 , w_18370 );
not (  , w_18371 );
and ( w_18370 , w_18371 , \5339_b0 );
or ( \5774_b1 , \5772_b1 , w_18373 );
not ( w_18373 , w_18374 );
and ( \5774_b0 , \5772_b0 , w_18375 );
and ( w_18374 ,  , w_18375 );
buf ( w_18373 , \5773_b1 );
not ( w_18373 , w_18376 );
not (  , w_18377 );
and ( w_18376 , w_18377 , \5773_b0 );
or ( \5775_b1 , \4234_b1 , w_18379 );
not ( w_18379 , w_18380 );
and ( \5775_b0 , \4234_b0 , w_18381 );
and ( w_18380 ,  , w_18381 );
buf ( w_18379 , \5774_b1 );
not ( w_18379 , w_18382 );
not (  , w_18383 );
and ( w_18382 , w_18383 , \5774_b0 );
or ( \5776_b1 , \5769_b1 , w_18385 );
not ( w_18385 , w_18386 );
and ( \5776_b0 , \5769_b0 , w_18387 );
and ( w_18386 ,  , w_18387 );
buf ( w_18385 , \5775_b1 );
not ( w_18385 , w_18388 );
not (  , w_18389 );
and ( w_18388 , w_18389 , \5775_b0 );
or ( \5777_b1 , \5761_b1 , \5776_b1 );
xor ( \5777_b0 , \5761_b0 , w_18390 );
not ( w_18390 , w_18391 );
and ( w_18391 , \5776_b1 , \5776_b0 );
buf ( \5778_b1 , \4026_b1 );
not ( \5778_b1 , w_18392 );
not ( \5778_b0 , w_18393 );
and ( w_18392 , w_18393 , \4026_b0 );
buf ( \5779_b1 , \4173_b1 );
not ( \5779_b1 , w_18394 );
not ( \5779_b0 , w_18395 );
and ( w_18394 , w_18395 , \4173_b0 );
or ( \5780_b1 , \5778_b1 , w_18396 );
or ( \5780_b0 , \5778_b0 , \5779_b0 );
not ( \5779_b0 , w_18397 );
and ( w_18397 , w_18396 , \5779_b1 );
or ( \5781_b1 , \4177_b1 , w_18399 );
not ( w_18399 , w_18400 );
and ( \5781_b0 , \4177_b0 , w_18401 );
and ( w_18400 ,  , w_18401 );
buf ( w_18399 , \5344_b1 );
not ( w_18399 , w_18402 );
not (  , w_18403 );
and ( w_18402 , w_18403 , \5344_b0 );
or ( \5782_b1 , \5780_b1 , w_18405 );
not ( w_18405 , w_18406 );
and ( \5782_b0 , \5780_b0 , w_18407 );
and ( w_18406 ,  , w_18407 );
buf ( w_18405 , \5781_b1 );
not ( w_18405 , w_18408 );
not (  , w_18409 );
and ( w_18408 , w_18409 , \5781_b0 );
buf ( \5783_b1 , \5782_b1 );
not ( \5783_b1 , w_18410 );
not ( \5783_b0 , w_18411 );
and ( w_18410 , w_18411 , \5782_b0 );
buf ( \5784_b1 , \4194_b1 );
not ( \5784_b1 , w_18412 );
not ( \5784_b0 , w_18413 );
and ( w_18412 , w_18413 , \4194_b0 );
or ( \5785_b1 , \5783_b1 , w_18414 );
or ( \5785_b0 , \5783_b0 , \5784_b0 );
not ( \5784_b0 , w_18415 );
and ( w_18415 , w_18414 , \5784_b1 );
buf ( \5786_b1 , \4023_b1 );
not ( \5786_b1 , w_18416 );
not ( \5786_b0 , w_18417 );
and ( w_18416 , w_18417 , \4023_b0 );
buf ( \5787_b1 , \4184_b1 );
not ( \5787_b1 , w_18418 );
not ( \5787_b0 , w_18419 );
and ( w_18418 , w_18419 , \4184_b0 );
or ( \5788_b1 , \5786_b1 , w_18420 );
or ( \5788_b0 , \5786_b0 , \5787_b0 );
not ( \5787_b0 , w_18421 );
and ( w_18421 , w_18420 , \5787_b1 );
or ( \5789_b1 , \4171_b1 , w_18423 );
not ( w_18423 , w_18424 );
and ( \5789_b0 , \4171_b0 , w_18425 );
and ( w_18424 ,  , w_18425 );
buf ( w_18423 , \5131_b1 );
not ( w_18423 , w_18426 );
not (  , w_18427 );
and ( w_18426 , w_18427 , \5131_b0 );
or ( \5790_b1 , \5788_b1 , w_18429 );
not ( w_18429 , w_18430 );
and ( \5790_b0 , \5788_b0 , w_18431 );
and ( w_18430 ,  , w_18431 );
buf ( w_18429 , \5789_b1 );
not ( w_18429 , w_18432 );
not (  , w_18433 );
and ( w_18432 , w_18433 , \5789_b0 );
or ( \5791_b1 , \5111_b1 , w_18435 );
not ( w_18435 , w_18436 );
and ( \5791_b0 , \5111_b0 , w_18437 );
and ( w_18436 ,  , w_18437 );
buf ( w_18435 , \5790_b1 );
not ( w_18435 , w_18438 );
not (  , w_18439 );
and ( w_18438 , w_18439 , \5790_b0 );
or ( \5792_b1 , \5785_b1 , w_18441 );
not ( w_18441 , w_18442 );
and ( \5792_b0 , \5785_b0 , w_18443 );
and ( w_18442 ,  , w_18443 );
buf ( w_18441 , \5791_b1 );
not ( w_18441 , w_18444 );
not (  , w_18445 );
and ( w_18444 , w_18445 , \5791_b0 );
or ( \5793_b1 , \5777_b1 , \5792_b1 );
not ( \5792_b1 , w_18446 );
and ( \5793_b0 , \5777_b0 , w_18447 );
and ( w_18446 , w_18447 , \5792_b0 );
or ( \5794_b1 , \5761_b1 , \5776_b1 );
not ( \5776_b1 , w_18448 );
and ( \5794_b0 , \5761_b0 , w_18449 );
and ( w_18448 , w_18449 , \5776_b0 );
or ( \5795_b1 , \5793_b1 , w_18450 );
or ( \5795_b0 , \5793_b0 , \5794_b0 );
not ( \5794_b0 , w_18451 );
and ( w_18451 , w_18450 , \5794_b1 );
buf ( \5796_b1 , \5795_b1 );
not ( \5796_b1 , w_18452 );
not ( \5796_b0 , w_18453 );
and ( w_18452 , w_18453 , \5795_b0 );
or ( \5797_b1 , \4224_b1 , w_18455 );
not ( w_18455 , w_18456 );
and ( \5797_b0 , \4224_b0 , w_18457 );
and ( w_18456 ,  , w_18457 );
buf ( w_18455 , \5388_b1 );
not ( w_18455 , w_18458 );
not (  , w_18459 );
and ( w_18458 , w_18459 , \5388_b0 );
or ( \5798_b1 , \5797_b1 , \4172_b1 );
not ( \4172_b1 , w_18460 );
and ( \5798_b0 , \5797_b0 , w_18461 );
and ( w_18460 , w_18461 , \4172_b0 );
buf ( \5799_b1 , \4048_b1 );
not ( \5799_b1 , w_18462 );
not ( \5799_b0 , w_18463 );
and ( w_18462 , w_18463 , \4048_b0 );
buf ( \5800_b1 , \4224_b1 );
not ( \5800_b1 , w_18464 );
not ( \5800_b0 , w_18465 );
and ( w_18464 , w_18465 , \4224_b0 );
buf ( \5801_b1 , \5800_b1 );
not ( \5801_b1 , w_18466 );
not ( \5801_b0 , w_18467 );
and ( w_18466 , w_18467 , \5800_b0 );
or ( \5802_b1 , \5799_b1 , w_18468 );
or ( \5802_b0 , \5799_b0 , \5801_b0 );
not ( \5801_b0 , w_18469 );
and ( w_18469 , w_18468 , \5801_b1 );
or ( \5803_b1 , \5802_b1 , w_18471 );
not ( w_18471 , w_18472 );
and ( \5803_b0 , \5802_b0 , w_18473 );
and ( w_18472 ,  , w_18473 );
buf ( w_18471 , \4492_b1 );
not ( w_18471 , w_18474 );
not (  , w_18475 );
and ( w_18474 , w_18475 , \4492_b0 );
or ( \5804_b1 , \5798_b1 , w_18477 );
not ( w_18477 , w_18478 );
and ( \5804_b0 , \5798_b0 , w_18479 );
and ( w_18478 ,  , w_18479 );
buf ( w_18477 , \5803_b1 );
not ( w_18477 , w_18480 );
not (  , w_18481 );
and ( w_18480 , w_18481 , \5803_b0 );
buf ( \5805_b1 , \4047_b1 );
not ( \5805_b1 , w_18482 );
not ( \5805_b0 , w_18483 );
and ( w_18482 , w_18483 , \4047_b0 );
buf ( \5806_b1 , \5270_b1 );
not ( \5806_b1 , w_18484 );
not ( \5806_b0 , w_18485 );
and ( w_18484 , w_18485 , \5270_b0 );
or ( \5807_b1 , \5805_b1 , w_18486 );
or ( \5807_b0 , \5805_b0 , \5806_b0 );
not ( \5806_b0 , w_18487 );
and ( w_18487 , w_18486 , \5806_b1 );
or ( \5808_b1 , \5016_b1 , w_18489 );
not ( w_18489 , w_18490 );
and ( \5808_b0 , \5016_b0 , w_18491 );
and ( w_18490 ,  , w_18491 );
buf ( w_18489 , \4178_b1 );
not ( w_18489 , w_18492 );
not (  , w_18493 );
and ( w_18492 , w_18493 , \4178_b0 );
or ( \5809_b1 , \5807_b1 , w_18495 );
not ( w_18495 , w_18496 );
and ( \5809_b0 , \5807_b0 , w_18497 );
and ( w_18496 ,  , w_18497 );
buf ( w_18495 , \5808_b1 );
not ( w_18495 , w_18498 );
not (  , w_18499 );
and ( w_18498 , w_18499 , \5808_b0 );
buf ( \5810_b1 , \5809_b1 );
not ( \5810_b1 , w_18500 );
not ( \5810_b0 , w_18501 );
and ( w_18500 , w_18501 , \5809_b0 );
buf ( \5811_b1 , \5390_b1 );
not ( \5811_b1 , w_18502 );
not ( \5811_b0 , w_18503 );
and ( w_18502 , w_18503 , \5390_b0 );
or ( \5812_b1 , \5810_b1 , w_18504 );
or ( \5812_b0 , \5810_b0 , \5811_b0 );
not ( \5811_b0 , w_18505 );
and ( w_18505 , w_18504 , \5811_b1 );
or ( \5813_b1 , \5706_b1 , w_18507 );
not ( w_18507 , w_18508 );
and ( \5813_b0 , \5706_b0 , w_18509 );
and ( w_18508 ,  , w_18509 );
buf ( w_18507 , \5021_b1 );
not ( w_18507 , w_18510 );
not (  , w_18511 );
and ( w_18510 , w_18511 , \5021_b0 );
or ( \5814_b1 , \5812_b1 , w_18513 );
not ( w_18513 , w_18514 );
and ( \5814_b0 , \5812_b0 , w_18515 );
and ( w_18514 ,  , w_18515 );
buf ( w_18513 , \5813_b1 );
not ( w_18513 , w_18516 );
not (  , w_18517 );
and ( w_18516 , w_18517 , \5813_b0 );
or ( \5815_b1 , \5804_b1 , w_18519 );
not ( w_18519 , w_18520 );
and ( \5815_b0 , \5804_b0 , w_18521 );
and ( w_18520 ,  , w_18521 );
buf ( w_18519 , \5814_b1 );
not ( w_18519 , w_18522 );
not (  , w_18523 );
and ( w_18522 , w_18523 , \5814_b0 );
buf ( \5816_b1 , \4192_b1 );
not ( \5816_b1 , w_18524 );
not ( \5816_b0 , w_18525 );
and ( w_18524 , w_18525 , \4192_b0 );
or ( \5817_b1 , \5816_b1 , \5650_b1 );
not ( \5650_b1 , w_18526 );
and ( \5817_b0 , \5816_b0 , w_18527 );
and ( w_18526 , w_18527 , \5650_b0 );
buf ( \5818_b1 , \5816_b1 );
not ( \5818_b1 , w_18528 );
not ( \5818_b0 , w_18529 );
and ( w_18528 , w_18529 , \5816_b0 );
or ( \5819_b1 , \5790_b1 , \4186_b1 );
not ( \4186_b1 , w_18530 );
and ( \5819_b0 , \5790_b0 , w_18531 );
and ( w_18530 , w_18531 , \4186_b0 );
or ( \5820_b1 , \5818_b1 , \5819_b1 );
not ( \5819_b1 , w_18532 );
and ( \5820_b0 , \5818_b0 , w_18533 );
and ( w_18532 , w_18533 , \5819_b0 );
or ( \5821_b1 , \5817_b1 , w_18535 );
not ( w_18535 , w_18536 );
and ( \5821_b0 , \5817_b0 , w_18537 );
and ( w_18536 ,  , w_18537 );
buf ( w_18535 , \5820_b1 );
not ( w_18535 , w_18538 );
not (  , w_18539 );
and ( w_18538 , w_18539 , \5820_b0 );
or ( \5822_b1 , \5815_b1 , \5821_b1 );
xor ( \5822_b0 , \5815_b0 , w_18540 );
not ( w_18540 , w_18541 );
and ( w_18541 , \5821_b1 , \5821_b0 );
buf ( \5823_b1 , \4230_b1 );
not ( \5823_b1 , w_18542 );
not ( \5823_b0 , w_18543 );
and ( w_18542 , w_18543 , \4230_b0 );
buf ( \5824_b1 , \5774_b1 );
not ( \5824_b1 , w_18544 );
not ( \5824_b0 , w_18545 );
and ( w_18544 , w_18545 , \5774_b0 );
buf ( \5825_b1 , \5824_b1 );
not ( \5825_b1 , w_18546 );
not ( \5825_b0 , w_18547 );
and ( w_18546 , w_18547 , \5824_b0 );
or ( \5826_b1 , \5823_b1 , \5825_b1 );
not ( \5825_b1 , w_18548 );
and ( \5826_b0 , \5823_b0 , w_18549 );
and ( w_18548 , w_18549 , \5825_b0 );
buf ( \5827_b1 , \4234_b1 );
not ( \5827_b1 , w_18550 );
not ( \5827_b0 , w_18551 );
and ( w_18550 , w_18551 , \4234_b0 );
or ( \5828_b1 , \5827_b1 , w_18553 );
not ( w_18553 , w_18554 );
and ( \5828_b0 , \5827_b0 , w_18555 );
and ( w_18554 ,  , w_18555 );
buf ( w_18553 , \5693_b1 );
not ( w_18553 , w_18556 );
not (  , w_18557 );
and ( w_18556 , w_18557 , \5693_b0 );
or ( \5829_b1 , \5826_b1 , w_18559 );
not ( w_18559 , w_18560 );
and ( \5829_b0 , \5826_b0 , w_18561 );
and ( w_18560 ,  , w_18561 );
buf ( w_18559 , \5828_b1 );
not ( w_18559 , w_18562 );
not (  , w_18563 );
and ( w_18562 , w_18563 , \5828_b0 );
or ( \5830_b1 , \5822_b1 , \5829_b1 );
xor ( \5830_b0 , \5822_b0 , w_18564 );
not ( w_18564 , w_18565 );
and ( w_18565 , \5829_b1 , \5829_b0 );
or ( \5831_b1 , \5796_b1 , w_18567 );
not ( w_18567 , w_18568 );
and ( \5831_b0 , \5796_b0 , w_18569 );
and ( w_18568 ,  , w_18569 );
buf ( w_18567 , \5830_b1 );
not ( w_18567 , w_18570 );
not (  , w_18571 );
and ( w_18570 , w_18571 , \5830_b0 );
buf ( \5832_b1 , \5831_b1 );
not ( \5832_b1 , w_18572 );
not ( \5832_b0 , w_18573 );
and ( w_18572 , w_18573 , \5831_b0 );
or ( \5833_b1 , \5804_b1 , \5814_b1 );
xor ( \5833_b0 , \5804_b0 , w_18574 );
not ( w_18574 , w_18575 );
and ( w_18575 , \5814_b1 , \5814_b0 );
or ( \5834_b1 , \4234_b1 , \4048_b1 );
not ( \4048_b1 , w_18576 );
and ( \5834_b0 , \4234_b0 , w_18577 );
and ( w_18576 , w_18577 , \4048_b0 );
buf ( \5835_b1 , \3963_b1 );
not ( \5835_b1 , w_18578 );
not ( \5835_b0 , w_18579 );
and ( w_18578 , w_18579 , \3963_b0 );
buf ( \5836_b1 , \5234_b1 );
not ( \5836_b1 , w_18580 );
not ( \5836_b0 , w_18581 );
and ( w_18580 , w_18581 , \5234_b0 );
or ( \5837_b1 , \5835_b1 , w_18582 );
or ( \5837_b0 , \5835_b0 , \5836_b0 );
not ( \5836_b0 , w_18583 );
and ( w_18583 , w_18582 , \5836_b1 );
or ( \5838_b1 , \4088_b1 , w_18585 );
not ( w_18585 , w_18586 );
and ( \5838_b0 , \4088_b0 , w_18587 );
and ( w_18586 ,  , w_18587 );
buf ( w_18585 , \4486_b1 );
not ( w_18585 , w_18588 );
not (  , w_18589 );
and ( w_18588 , w_18589 , \4486_b0 );
or ( \5839_b1 , \5837_b1 , w_18591 );
not ( w_18591 , w_18592 );
and ( \5839_b0 , \5837_b0 , w_18593 );
and ( w_18592 ,  , w_18593 );
buf ( w_18591 , \5838_b1 );
not ( w_18591 , w_18594 );
not (  , w_18595 );
and ( w_18594 , w_18595 , \5838_b0 );
buf ( \5840_b1 , \5839_b1 );
not ( \5840_b1 , w_18596 );
not ( \5840_b0 , w_18597 );
and ( w_18596 , w_18597 , \5839_b0 );
buf ( \5841_b1 , \4085_b1 );
not ( \5841_b1 , w_18598 );
not ( \5841_b0 , w_18599 );
and ( w_18598 , w_18599 , \4085_b0 );
or ( \5842_b1 , \5840_b1 , w_18600 );
or ( \5842_b0 , \5840_b0 , \5841_b0 );
not ( \5841_b0 , w_18601 );
and ( w_18601 , w_18600 , \5841_b1 );
buf ( \5843_b1 , \3958_b1 );
not ( \5843_b1 , w_18602 );
not ( \5843_b0 , w_18603 );
and ( w_18602 , w_18603 , \3958_b0 );
buf ( \5844_b1 , \5234_b1 );
not ( \5844_b1 , w_18604 );
not ( \5844_b0 , w_18605 );
and ( w_18604 , w_18605 , \5234_b0 );
or ( \5845_b1 , \5843_b1 , w_18606 );
or ( \5845_b0 , \5843_b0 , \5844_b0 );
not ( \5844_b0 , w_18607 );
and ( w_18607 , w_18606 , \5844_b1 );
or ( \5846_b1 , \4088_b1 , w_18609 );
not ( w_18609 , w_18610 );
and ( \5846_b0 , \4088_b0 , w_18611 );
and ( w_18610 ,  , w_18611 );
buf ( w_18609 , \4473_b1 );
not ( w_18609 , w_18612 );
not (  , w_18613 );
and ( w_18612 , w_18613 , \4473_b0 );
or ( \5847_b1 , \5845_b1 , w_18615 );
not ( w_18615 , w_18616 );
and ( \5847_b0 , \5845_b0 , w_18617 );
and ( w_18616 ,  , w_18617 );
buf ( w_18615 , \5846_b1 );
not ( w_18615 , w_18618 );
not (  , w_18619 );
and ( w_18618 , w_18619 , \5846_b0 );
or ( \5848_b1 , \4596_b1 , w_18621 );
not ( w_18621 , w_18622 );
and ( \5848_b0 , \4596_b0 , w_18623 );
and ( w_18622 ,  , w_18623 );
buf ( w_18621 , \5847_b1 );
not ( w_18621 , w_18624 );
not (  , w_18625 );
and ( w_18624 , w_18625 , \5847_b0 );
or ( \5849_b1 , \5842_b1 , w_18627 );
not ( w_18627 , w_18628 );
and ( \5849_b0 , \5842_b0 , w_18629 );
and ( w_18628 ,  , w_18629 );
buf ( w_18627 , \5848_b1 );
not ( w_18627 , w_18630 );
not (  , w_18631 );
and ( w_18630 , w_18631 , \5848_b0 );
or ( \5850_b1 , \5834_b1 , w_18632 );
or ( \5850_b0 , \5834_b0 , \5849_b0 );
not ( \5849_b0 , w_18633 );
and ( w_18633 , w_18632 , \5849_b1 );
buf ( \5851_b1 , \4043_b1 );
not ( \5851_b1 , w_18634 );
not ( \5851_b0 , w_18635 );
and ( w_18634 , w_18635 , \4043_b0 );
buf ( \5852_b1 , \5178_b1 );
not ( \5852_b1 , w_18636 );
not ( \5852_b0 , w_18637 );
and ( w_18636 , w_18637 , \5178_b0 );
or ( \5853_b1 , \5851_b1 , w_18638 );
or ( \5853_b0 , \5851_b0 , \5852_b0 );
not ( \5852_b0 , w_18639 );
and ( w_18639 , w_18638 , \5852_b1 );
or ( \5854_b1 , \4548_b1 , w_18641 );
not ( w_18641 , w_18642 );
and ( \5854_b0 , \4548_b0 , w_18643 );
and ( w_18642 ,  , w_18643 );
buf ( w_18641 , \4217_b1 );
not ( w_18641 , w_18644 );
not (  , w_18645 );
and ( w_18644 , w_18645 , \4217_b0 );
or ( \5855_b1 , \5853_b1 , w_18647 );
not ( w_18647 , w_18648 );
and ( \5855_b0 , \5853_b0 , w_18649 );
and ( w_18648 ,  , w_18649 );
buf ( w_18647 , \5854_b1 );
not ( w_18647 , w_18650 );
not (  , w_18651 );
and ( w_18650 , w_18651 , \5854_b0 );
buf ( \5856_b1 , \5855_b1 );
not ( \5856_b1 , w_18652 );
not ( \5856_b0 , w_18653 );
and ( w_18652 , w_18653 , \5855_b0 );
buf ( \5857_b1 , \4662_b1 );
not ( \5857_b1 , w_18654 );
not ( \5857_b0 , w_18655 );
and ( w_18654 , w_18655 , \4662_b0 );
or ( \5858_b1 , \5856_b1 , w_18656 );
or ( \5858_b0 , \5856_b0 , \5857_b0 );
not ( \5857_b0 , w_18657 );
and ( w_18657 , w_18656 , \5857_b1 );
buf ( \5859_b1 , \4041_b1 );
not ( \5859_b1 , w_18658 );
not ( \5859_b0 , w_18659 );
and ( w_18658 , w_18659 , \4041_b0 );
buf ( \5860_b1 , \4666_b1 );
not ( \5860_b1 , w_18660 );
not ( \5860_b0 , w_18661 );
and ( w_18660 , w_18661 , \4666_b0 );
or ( \5861_b1 , \5859_b1 , w_18662 );
or ( \5861_b0 , \5859_b0 , \5860_b0 );
not ( \5860_b0 , w_18663 );
and ( w_18663 , w_18662 , \5860_b1 );
or ( \5862_b1 , \4665_b1 , w_18665 );
not ( w_18665 , w_18666 );
and ( \5862_b0 , \4665_b0 , w_18667 );
and ( w_18666 ,  , w_18667 );
buf ( w_18665 , \4238_b1 );
not ( w_18665 , w_18668 );
not (  , w_18669 );
and ( w_18668 , w_18669 , \4238_b0 );
or ( \5863_b1 , \5861_b1 , w_18671 );
not ( w_18671 , w_18672 );
and ( \5863_b0 , \5861_b0 , w_18673 );
and ( w_18672 ,  , w_18673 );
buf ( w_18671 , \5862_b1 );
not ( w_18671 , w_18674 );
not (  , w_18675 );
and ( w_18674 , w_18675 , \5862_b0 );
or ( \5864_b1 , \4672_b1 , w_18677 );
not ( w_18677 , w_18678 );
and ( \5864_b0 , \4672_b0 , w_18679 );
and ( w_18678 ,  , w_18679 );
buf ( w_18677 , \5863_b1 );
not ( w_18677 , w_18680 );
not (  , w_18681 );
and ( w_18680 , w_18681 , \5863_b0 );
or ( \5865_b1 , \5858_b1 , w_18683 );
not ( w_18683 , w_18684 );
and ( \5865_b0 , \5858_b0 , w_18685 );
and ( w_18684 ,  , w_18685 );
buf ( w_18683 , \5864_b1 );
not ( w_18683 , w_18686 );
not (  , w_18687 );
and ( w_18686 , w_18687 , \5864_b0 );
or ( \5866_b1 , \5850_b1 , w_18689 );
not ( w_18689 , w_18690 );
and ( \5866_b0 , \5850_b0 , w_18691 );
and ( w_18690 ,  , w_18691 );
buf ( w_18689 , \5865_b1 );
not ( w_18689 , w_18692 );
not (  , w_18693 );
and ( w_18692 , w_18693 , \5865_b0 );
or ( \5867_b1 , \4234_b1 , w_18695 );
not ( w_18695 , w_18696 );
and ( \5867_b0 , \4234_b0 , w_18697 );
and ( w_18696 ,  , w_18697 );
buf ( w_18695 , \4048_b1 );
not ( w_18695 , w_18698 );
not (  , w_18699 );
and ( w_18698 , w_18699 , \4048_b0 );
buf ( \5868_b1 , \5867_b1 );
not ( \5868_b1 , w_18700 );
not ( \5868_b0 , w_18701 );
and ( w_18700 , w_18701 , \5867_b0 );
or ( \5869_b1 , \5868_b1 , w_18703 );
not ( w_18703 , w_18704 );
and ( \5869_b0 , \5868_b0 , w_18705 );
and ( w_18704 ,  , w_18705 );
buf ( w_18703 , \5849_b1 );
not ( w_18703 , w_18706 );
not (  , w_18707 );
and ( w_18706 , w_18707 , \5849_b0 );
or ( \5870_b1 , \5866_b1 , w_18709 );
not ( w_18709 , w_18710 );
and ( \5870_b0 , \5866_b0 , w_18711 );
and ( w_18710 ,  , w_18711 );
buf ( w_18709 , \5869_b1 );
not ( w_18709 , w_18712 );
not (  , w_18713 );
and ( w_18712 , w_18713 , \5869_b0 );
or ( \5871_b1 , \5833_b1 , \5870_b1 );
xor ( \5871_b0 , \5833_b0 , w_18714 );
not ( w_18714 , w_18715 );
and ( w_18715 , \5870_b1 , \5870_b0 );
buf ( \5872_b1 , \4045_b1 );
not ( \5872_b1 , w_18716 );
not ( \5872_b0 , w_18717 );
and ( w_18716 , w_18717 , \4045_b0 );
buf ( \5873_b1 , \1395_b1 );
buf ( \5873_b0 , \1395_b0 );
buf ( \5874_b1 , \5873_b1 );
not ( \5874_b1 , w_18718 );
not ( \5874_b0 , w_18719 );
and ( w_18718 , w_18719 , \5873_b0 );
buf ( \5875_b1 , \5874_b1 );
not ( \5875_b1 , w_18720 );
not ( \5875_b0 , w_18721 );
and ( w_18720 , w_18721 , \5874_b0 );
or ( \5876_b1 , \5872_b1 , w_18722 );
or ( \5876_b0 , \5872_b0 , \5875_b0 );
not ( \5875_b0 , w_18723 );
and ( w_18723 , w_18722 , \5875_b1 );
or ( \5877_b1 , \5273_b1 , w_18725 );
not ( w_18725 , w_18726 );
and ( \5877_b0 , \5273_b0 , w_18727 );
and ( w_18726 ,  , w_18727 );
buf ( w_18725 , \4286_b1 );
not ( w_18725 , w_18728 );
not (  , w_18729 );
and ( w_18728 , w_18729 , \4286_b0 );
or ( \5878_b1 , \5876_b1 , w_18731 );
not ( w_18731 , w_18732 );
and ( \5878_b0 , \5876_b0 , w_18733 );
and ( w_18732 ,  , w_18733 );
buf ( w_18731 , \5877_b1 );
not ( w_18731 , w_18734 );
not (  , w_18735 );
and ( w_18734 , w_18735 , \5877_b0 );
buf ( \5879_b1 , \5878_b1 );
not ( \5879_b1 , w_18736 );
not ( \5879_b0 , w_18737 );
and ( w_18736 , w_18737 , \5878_b0 );
buf ( \5880_b1 , \5019_b1 );
not ( \5880_b1 , w_18738 );
not ( \5880_b0 , w_18739 );
and ( w_18738 , w_18739 , \5019_b0 );
or ( \5881_b1 , \5879_b1 , w_18740 );
or ( \5881_b0 , \5879_b0 , \5880_b0 );
not ( \5880_b0 , w_18741 );
and ( w_18741 , w_18740 , \5880_b1 );
or ( \5882_b1 , \5809_b1 , w_18743 );
not ( w_18743 , w_18744 );
and ( \5882_b0 , \5809_b0 , w_18745 );
and ( w_18744 ,  , w_18745 );
buf ( w_18743 , \5021_b1 );
not ( w_18743 , w_18746 );
not (  , w_18747 );
and ( w_18746 , w_18747 , \5021_b0 );
or ( \5883_b1 , \5881_b1 , w_18749 );
not ( w_18749 , w_18750 );
and ( \5883_b0 , \5881_b0 , w_18751 );
and ( w_18750 ,  , w_18751 );
buf ( w_18749 , \5882_b1 );
not ( w_18749 , w_18752 );
not (  , w_18753 );
and ( w_18752 , w_18753 , \5882_b0 );
buf ( \5884_b1 , \5883_b1 );
not ( \5884_b1 , w_18754 );
not ( \5884_b0 , w_18755 );
and ( w_18754 , w_18755 , \5883_b0 );
buf ( \5885_b1 , \4023_b1 );
not ( \5885_b1 , w_18756 );
not ( \5885_b0 , w_18757 );
and ( w_18756 , w_18757 , \4023_b0 );
buf ( \5886_b1 , \4110_b1 );
not ( \5886_b1 , w_18758 );
not ( \5886_b0 , w_18759 );
and ( w_18758 , w_18759 , \4110_b0 );
or ( \5887_b1 , \5885_b1 , w_18760 );
or ( \5887_b0 , \5885_b0 , \5886_b0 );
not ( \5886_b0 , w_18761 );
and ( w_18761 , w_18760 , \5886_b1 );
or ( \5888_b1 , \4109_b1 , w_18763 );
not ( w_18763 , w_18764 );
and ( \5888_b0 , \4109_b0 , w_18765 );
and ( w_18764 ,  , w_18765 );
buf ( w_18763 , \5131_b1 );
not ( w_18763 , w_18766 );
not (  , w_18767 );
and ( w_18766 , w_18767 , \5131_b0 );
or ( \5889_b1 , \5887_b1 , w_18769 );
not ( w_18769 , w_18770 );
and ( \5889_b0 , \5887_b0 , w_18771 );
and ( w_18770 ,  , w_18771 );
buf ( w_18769 , \5888_b1 );
not ( w_18769 , w_18772 );
not (  , w_18773 );
and ( w_18772 , w_18773 , \5888_b0 );
buf ( \5890_b1 , \5889_b1 );
not ( \5890_b1 , w_18774 );
not ( \5890_b0 , w_18775 );
and ( w_18774 , w_18775 , \5889_b0 );
buf ( \5891_b1 , \5431_b1 );
not ( \5891_b1 , w_18776 );
not ( \5891_b0 , w_18777 );
and ( w_18776 , w_18777 , \5431_b0 );
or ( \5892_b1 , \5890_b1 , w_18778 );
or ( \5892_b0 , \5890_b0 , \5891_b0 );
not ( \5891_b0 , w_18779 );
and ( w_18779 , w_18778 , \5891_b1 );
buf ( \5893_b1 , \4019_b1 );
not ( \5893_b1 , w_18780 );
not ( \5893_b0 , w_18781 );
and ( w_18780 , w_18781 , \4019_b0 );
buf ( \5894_b1 , \4142_b1 );
not ( \5894_b1 , w_18782 );
not ( \5894_b0 , w_18783 );
and ( w_18782 , w_18783 , \4142_b0 );
or ( \5895_b1 , \5893_b1 , w_18784 );
or ( \5895_b0 , \5893_b0 , \5894_b0 );
not ( \5894_b0 , w_18785 );
and ( w_18785 , w_18784 , \5894_b1 );
or ( \5896_b1 , \4109_b1 , w_18787 );
not ( w_18787 , w_18788 );
and ( \5896_b0 , \4109_b0 , w_18789 );
and ( w_18788 ,  , w_18789 );
buf ( w_18787 , \4585_b1 );
not ( w_18787 , w_18790 );
not (  , w_18791 );
and ( w_18790 , w_18791 , \4585_b0 );
or ( \5897_b1 , \5895_b1 , w_18793 );
not ( w_18793 , w_18794 );
and ( \5897_b0 , \5895_b0 , w_18795 );
and ( w_18794 ,  , w_18795 );
buf ( w_18793 , \5896_b1 );
not ( w_18793 , w_18796 );
not (  , w_18797 );
and ( w_18796 , w_18797 , \5896_b0 );
or ( \5898_b1 , \5897_b1 , w_18799 );
not ( w_18799 , w_18800 );
and ( \5898_b0 , \5897_b0 , w_18801 );
and ( w_18800 ,  , w_18801 );
buf ( w_18799 , \4139_b1 );
not ( w_18799 , w_18802 );
not (  , w_18803 );
and ( w_18802 , w_18803 , \4139_b0 );
or ( \5899_b1 , \5892_b1 , w_18805 );
not ( w_18805 , w_18806 );
and ( \5899_b0 , \5892_b0 , w_18807 );
and ( w_18806 ,  , w_18807 );
buf ( w_18805 , \5898_b1 );
not ( w_18805 , w_18808 );
not (  , w_18809 );
and ( w_18808 , w_18809 , \5898_b0 );
buf ( \5900_b1 , \5899_b1 );
not ( \5900_b1 , w_18810 );
not ( \5900_b0 , w_18811 );
and ( w_18810 , w_18811 , \5899_b0 );
or ( \5901_b1 , \5884_b1 , w_18812 );
or ( \5901_b0 , \5884_b0 , \5900_b0 );
not ( \5900_b0 , w_18813 );
and ( w_18813 , w_18812 , \5900_b1 );
or ( \5902_b1 , \5899_b1 , w_18814 );
or ( \5902_b0 , \5899_b0 , \5883_b0 );
not ( \5883_b0 , w_18815 );
and ( w_18815 , w_18814 , \5883_b1 );
buf ( \5903_b1 , \4046_b1 );
not ( \5903_b1 , w_18816 );
not ( \5903_b0 , w_18817 );
and ( w_18816 , w_18817 , \4046_b0 );
buf ( \5904_b1 , \4069_b1 );
buf ( \5904_b0 , \4069_b0 );
buf ( \5905_b1 , \5904_b1 );
not ( \5905_b1 , w_18818 );
not ( \5905_b0 , w_18819 );
and ( w_18818 , w_18819 , \5904_b0 );
or ( \5906_b1 , \5903_b1 , w_18820 );
or ( \5906_b0 , \5903_b0 , \5905_b0 );
not ( \5905_b0 , w_18821 );
and ( w_18821 , w_18820 , \5905_b1 );
or ( \5907_b1 , \5060_b1 , w_18823 );
not ( w_18823 , w_18824 );
and ( \5907_b0 , \5060_b0 , w_18825 );
and ( w_18824 ,  , w_18825 );
buf ( w_18823 , \4256_b1 );
not ( w_18823 , w_18826 );
not (  , w_18827 );
and ( w_18826 , w_18827 , \4256_b0 );
or ( \5908_b1 , \5906_b1 , w_18829 );
not ( w_18829 , w_18830 );
and ( \5908_b0 , \5906_b0 , w_18831 );
and ( w_18830 ,  , w_18831 );
buf ( w_18829 , \5907_b1 );
not ( w_18829 , w_18832 );
not (  , w_18833 );
and ( w_18832 , w_18833 , \5907_b0 );
buf ( \5909_b1 , \5908_b1 );
not ( \5909_b1 , w_18834 );
not ( \5909_b0 , w_18835 );
and ( w_18834 , w_18835 , \5908_b0 );
buf ( \5910_b1 , \5361_b1 );
not ( \5910_b1 , w_18836 );
not ( \5910_b0 , w_18837 );
and ( w_18836 , w_18837 , \5361_b0 );
or ( \5911_b1 , \5909_b1 , w_18838 );
or ( \5911_b0 , \5909_b0 , \5910_b0 );
not ( \5910_b0 , w_18839 );
and ( w_18839 , w_18838 , \5910_b1 );
or ( \5912_b1 , \4055_b1 , w_18841 );
not ( w_18841 , w_18842 );
and ( \5912_b0 , \4055_b0 , w_18843 );
and ( w_18842 ,  , w_18843 );
buf ( w_18841 , \5751_b1 );
not ( w_18841 , w_18844 );
not (  , w_18845 );
and ( w_18844 , w_18845 , \5751_b0 );
or ( \5913_b1 , \5911_b1 , w_18847 );
not ( w_18847 , w_18848 );
and ( \5913_b0 , \5911_b0 , w_18849 );
and ( w_18848 ,  , w_18849 );
buf ( w_18847 , \5912_b1 );
not ( w_18847 , w_18850 );
not (  , w_18851 );
and ( w_18850 , w_18851 , \5912_b0 );
or ( \5914_b1 , \5902_b1 , w_18853 );
not ( w_18853 , w_18854 );
and ( \5914_b0 , \5902_b0 , w_18855 );
and ( w_18854 ,  , w_18855 );
buf ( w_18853 , \5913_b1 );
not ( w_18853 , w_18856 );
not (  , w_18857 );
and ( w_18856 , w_18857 , \5913_b0 );
or ( \5915_b1 , \5901_b1 , w_18859 );
not ( w_18859 , w_18860 );
and ( \5915_b0 , \5901_b0 , w_18861 );
and ( w_18860 ,  , w_18861 );
buf ( w_18859 , \5914_b1 );
not ( w_18859 , w_18862 );
not (  , w_18863 );
and ( w_18862 , w_18863 , \5914_b0 );
or ( \5916_b1 , \5871_b1 , \5915_b1 );
not ( \5915_b1 , w_18864 );
and ( \5916_b0 , \5871_b0 , w_18865 );
and ( w_18864 , w_18865 , \5915_b0 );
or ( \5917_b1 , \5833_b1 , \5870_b1 );
not ( \5870_b1 , w_18866 );
and ( \5917_b0 , \5833_b0 , w_18867 );
and ( w_18866 , w_18867 , \5870_b0 );
or ( \5918_b1 , \5916_b1 , w_18868 );
or ( \5918_b0 , \5916_b0 , \5917_b0 );
not ( \5917_b0 , w_18869 );
and ( w_18869 , w_18868 , \5917_b1 );
buf ( \5919_b1 , \5918_b1 );
not ( \5919_b1 , w_18870 );
not ( \5919_b0 , w_18871 );
and ( w_18870 , w_18871 , \5918_b0 );
or ( \5920_b1 , \5832_b1 , w_18872 );
or ( \5920_b0 , \5832_b0 , \5919_b0 );
not ( \5919_b0 , w_18873 );
and ( w_18873 , w_18872 , \5919_b1 );
or ( \5921_b1 , \5830_b1 , w_18874 );
or ( \5921_b0 , \5830_b0 , \5796_b0 );
not ( \5796_b0 , w_18875 );
and ( w_18875 , w_18874 , \5796_b1 );
or ( \5922_b1 , \5920_b1 , w_18877 );
not ( w_18877 , w_18878 );
and ( \5922_b0 , \5920_b0 , w_18879 );
and ( w_18878 ,  , w_18879 );
buf ( w_18877 , \5921_b1 );
not ( w_18877 , w_18880 );
not (  , w_18881 );
and ( w_18880 , w_18881 , \5921_b0 );
buf ( \5923_b1 , \5922_b1 );
not ( \5923_b1 , w_18882 );
not ( \5923_b0 , w_18883 );
and ( w_18882 , w_18883 , \5922_b0 );
buf ( \5924_b1 , \5759_b1 );
not ( \5924_b1 , w_18884 );
not ( \5924_b0 , w_18885 );
and ( w_18884 , w_18885 , \5759_b0 );
buf ( \5925_b1 , \4558_b1 );
not ( \5925_b1 , w_18886 );
not ( \5925_b0 , w_18887 );
and ( w_18886 , w_18887 , \4558_b0 );
or ( \5926_b1 , \5924_b1 , w_18888 );
or ( \5926_b0 , \5924_b0 , \5925_b0 );
not ( \5925_b0 , w_18889 );
and ( w_18889 , w_18888 , \5925_b1 );
or ( \5927_b1 , \4055_b1 , w_18891 );
not ( w_18891 , w_18892 );
and ( \5927_b0 , \4055_b0 , w_18893 );
and ( w_18892 ,  , w_18893 );
buf ( w_18891 , \5640_b1 );
not ( w_18891 , w_18894 );
not (  , w_18895 );
and ( w_18894 , w_18895 , \5640_b0 );
or ( \5928_b1 , \5926_b1 , w_18897 );
not ( w_18897 , w_18898 );
and ( \5928_b0 , \5926_b0 , w_18899 );
and ( w_18898 ,  , w_18899 );
buf ( w_18897 , \5927_b1 );
not ( w_18897 , w_18900 );
not (  , w_18901 );
and ( w_18900 , w_18901 , \5927_b0 );
buf ( \5929_b1 , \5928_b1 );
not ( \5929_b1 , w_18902 );
not ( \5929_b0 , w_18903 );
and ( w_18902 , w_18903 , \5928_b0 );
buf ( \5930_b1 , \4046_b1 );
not ( \5930_b1 , w_18904 );
not ( \5930_b0 , w_18905 );
and ( w_18904 , w_18905 , \4046_b0 );
buf ( \5931_b1 , \4089_b1 );
not ( \5931_b1 , w_18906 );
not ( \5931_b0 , w_18907 );
and ( w_18906 , w_18907 , \4089_b0 );
or ( \5932_b1 , \5930_b1 , w_18908 );
or ( \5932_b0 , \5930_b0 , \5931_b0 );
not ( \5931_b0 , w_18909 );
and ( w_18909 , w_18908 , \5931_b1 );
or ( \5933_b1 , \4088_b1 , w_18911 );
not ( w_18911 , w_18912 );
and ( \5933_b0 , \4088_b0 , w_18913 );
and ( w_18912 ,  , w_18913 );
buf ( w_18911 , \4256_b1 );
not ( w_18911 , w_18914 );
not (  , w_18915 );
and ( w_18914 , w_18915 , \4256_b0 );
or ( \5934_b1 , \5932_b1 , w_18917 );
not ( w_18917 , w_18918 );
and ( \5934_b0 , \5932_b0 , w_18919 );
and ( w_18918 ,  , w_18919 );
buf ( w_18917 , \5933_b1 );
not ( w_18917 , w_18920 );
not (  , w_18921 );
and ( w_18920 , w_18921 , \5933_b0 );
buf ( \5935_b1 , \5934_b1 );
not ( \5935_b1 , w_18922 );
not ( \5935_b0 , w_18923 );
and ( w_18922 , w_18923 , \5934_b0 );
buf ( \5936_b1 , \4086_b1 );
not ( \5936_b1 , w_18924 );
not ( \5936_b0 , w_18925 );
and ( w_18924 , w_18925 , \4086_b0 );
or ( \5937_b1 , \5935_b1 , w_18926 );
or ( \5937_b0 , \5935_b0 , \5936_b0 );
not ( \5936_b0 , w_18927 );
and ( w_18927 , w_18926 , \5936_b1 );
or ( \5938_b1 , \4596_b1 , w_18929 );
not ( w_18929 , w_18930 );
and ( \5938_b0 , \4596_b0 , w_18931 );
and ( w_18930 ,  , w_18931 );
buf ( w_18929 , \5594_b1 );
not ( w_18929 , w_18932 );
not (  , w_18933 );
and ( w_18932 , w_18933 , \5594_b0 );
or ( \5939_b1 , \5937_b1 , w_18935 );
not ( w_18935 , w_18936 );
and ( \5939_b0 , \5937_b0 , w_18937 );
and ( w_18936 ,  , w_18937 );
buf ( w_18935 , \5938_b1 );
not ( w_18935 , w_18938 );
not (  , w_18939 );
and ( w_18938 , w_18939 , \5938_b0 );
buf ( \5940_b1 , \5939_b1 );
not ( \5940_b1 , w_18940 );
not ( \5940_b0 , w_18941 );
and ( w_18940 , w_18941 , \5939_b0 );
or ( \5941_b1 , \5929_b1 , w_18942 );
or ( \5941_b0 , \5929_b0 , \5940_b0 );
not ( \5940_b0 , w_18943 );
and ( w_18943 , w_18942 , \5940_b1 );
or ( \5942_b1 , \5939_b1 , w_18944 );
or ( \5942_b0 , \5939_b0 , \5928_b0 );
not ( \5928_b0 , w_18945 );
and ( w_18945 , w_18944 , \5928_b1 );
buf ( \5943_b1 , \3963_b1 );
not ( \5943_b1 , w_18946 );
not ( \5943_b0 , w_18947 );
and ( w_18946 , w_18947 , \3963_b0 );
buf ( \5944_b1 , \4110_b1 );
not ( \5944_b1 , w_18948 );
not ( \5944_b0 , w_18949 );
and ( w_18948 , w_18949 , \4110_b0 );
or ( \5945_b1 , \5943_b1 , w_18950 );
or ( \5945_b0 , \5943_b0 , \5944_b0 );
not ( \5944_b0 , w_18951 );
and ( w_18951 , w_18950 , \5944_b1 );
or ( \5946_b1 , \4115_b1 , w_18953 );
not ( w_18953 , w_18954 );
and ( \5946_b0 , \4115_b0 , w_18955 );
and ( w_18954 ,  , w_18955 );
buf ( w_18953 , \4486_b1 );
not ( w_18953 , w_18956 );
not (  , w_18957 );
and ( w_18956 , w_18957 , \4486_b0 );
or ( \5947_b1 , \5945_b1 , w_18959 );
not ( w_18959 , w_18960 );
and ( \5947_b0 , \5945_b0 , w_18961 );
and ( w_18960 ,  , w_18961 );
buf ( w_18959 , \5946_b1 );
not ( w_18959 , w_18962 );
not (  , w_18963 );
and ( w_18962 , w_18963 , \5946_b0 );
buf ( \5948_b1 , \5947_b1 );
not ( \5948_b1 , w_18964 );
not ( \5948_b0 , w_18965 );
and ( w_18964 , w_18965 , \5947_b0 );
buf ( \5949_b1 , \4425_b1 );
not ( \5949_b1 , w_18966 );
not ( \5949_b0 , w_18967 );
and ( w_18966 , w_18967 , \4425_b0 );
or ( \5950_b1 , \5948_b1 , w_18968 );
or ( \5950_b0 , \5948_b0 , \5949_b0 );
not ( \5949_b0 , w_18969 );
and ( w_18969 , w_18968 , \5949_b1 );
or ( \5951_b1 , \4429_b1 , w_18971 );
not ( w_18971 , w_18972 );
and ( \5951_b0 , \4429_b0 , w_18973 );
and ( w_18972 ,  , w_18973 );
buf ( w_18971 , \5604_b1 );
not ( w_18971 , w_18974 );
not (  , w_18975 );
and ( w_18974 , w_18975 , \5604_b0 );
or ( \5952_b1 , \5950_b1 , w_18977 );
not ( w_18977 , w_18978 );
and ( \5952_b0 , \5950_b0 , w_18979 );
and ( w_18978 ,  , w_18979 );
buf ( w_18977 , \5951_b1 );
not ( w_18977 , w_18980 );
not (  , w_18981 );
and ( w_18980 , w_18981 , \5951_b0 );
or ( \5953_b1 , \5942_b1 , w_18983 );
not ( w_18983 , w_18984 );
and ( \5953_b0 , \5942_b0 , w_18985 );
and ( w_18984 ,  , w_18985 );
buf ( w_18983 , \5952_b1 );
not ( w_18983 , w_18986 );
not (  , w_18987 );
and ( w_18986 , w_18987 , \5952_b0 );
or ( \5954_b1 , \5941_b1 , w_18989 );
not ( w_18989 , w_18990 );
and ( \5954_b0 , \5941_b0 , w_18991 );
and ( w_18990 ,  , w_18991 );
buf ( w_18989 , \5953_b1 );
not ( w_18989 , w_18992 );
not (  , w_18993 );
and ( w_18992 , w_18993 , \5953_b0 );
or ( \5955_b1 , \5609_b1 , \5621_b1 );
xor ( \5955_b0 , \5609_b0 , w_18994 );
not ( w_18994 , w_18995 );
and ( w_18995 , \5621_b1 , \5621_b0 );
or ( \5956_b1 , \5955_b1 , w_18996 );
xor ( \5956_b0 , \5955_b0 , w_18998 );
not ( w_18998 , w_18999 );
and ( w_18999 , w_18996 , w_18997 );
buf ( w_18996 , \5599_b1 );
not ( w_18996 , w_19000 );
not ( w_18997 , w_19001 );
and ( w_19000 , w_19001 , \5599_b0 );
or ( \5957_b1 , \5954_b1 , \5956_b1 );
xor ( \5957_b0 , \5954_b0 , w_19002 );
not ( w_19002 , w_19003 );
and ( w_19003 , \5956_b1 , \5956_b0 );
or ( \5958_b1 , \5645_b1 , \5655_b1 );
xor ( \5958_b0 , \5645_b0 , w_19004 );
not ( w_19004 , w_19005 );
and ( w_19005 , \5655_b1 , \5655_b0 );
or ( \5959_b1 , \5958_b1 , \5665_b1 );
xor ( \5959_b0 , \5958_b0 , w_19006 );
not ( w_19006 , w_19007 );
and ( w_19007 , \5665_b1 , \5665_b0 );
or ( \5960_b1 , \5957_b1 , w_19008 );
xor ( \5960_b0 , \5957_b0 , w_19010 );
not ( w_19010 , w_19011 );
and ( w_19011 , w_19008 , w_19009 );
buf ( w_19008 , \5959_b1 );
not ( w_19008 , w_19012 );
not ( w_19009 , w_19013 );
and ( w_19012 , w_19013 , \5959_b0 );
buf ( \5961_b1 , \5960_b1 );
not ( \5961_b1 , w_19014 );
not ( \5961_b0 , w_19015 );
and ( w_19014 , w_19015 , \5960_b0 );
or ( \5962_b1 , \5923_b1 , w_19016 );
or ( \5962_b0 , \5923_b0 , \5961_b0 );
not ( \5961_b0 , w_19017 );
and ( w_19017 , w_19016 , \5961_b1 );
buf ( \5963_b1 , \5922_b1 );
not ( \5963_b1 , w_19018 );
not ( \5963_b0 , w_19019 );
and ( w_19018 , w_19019 , \5922_b0 );
or ( \5964_b1 , \5954_b1 , \5956_b1 );
xor ( \5964_b0 , \5954_b0 , w_19020 );
not ( w_19020 , w_19021 );
and ( w_19021 , \5956_b1 , \5956_b0 );
or ( \5965_b1 , \5964_b1 , \5959_b1 );
xor ( \5965_b0 , \5964_b0 , w_19022 );
not ( w_19022 , w_19023 );
and ( w_19023 , \5959_b1 , \5959_b0 );
or ( \5966_b1 , \5963_b1 , w_19025 );
not ( w_19025 , w_19026 );
and ( \5966_b0 , \5963_b0 , w_19027 );
and ( w_19026 ,  , w_19027 );
buf ( w_19025 , \5965_b1 );
not ( w_19025 , w_19028 );
not (  , w_19029 );
and ( w_19028 , w_19029 , \5965_b0 );
or ( \5967_b1 , \5962_b1 , w_19031 );
not ( w_19031 , w_19032 );
and ( \5967_b0 , \5962_b0 , w_19033 );
and ( w_19032 ,  , w_19033 );
buf ( w_19031 , \5966_b1 );
not ( w_19031 , w_19034 );
not (  , w_19035 );
and ( w_19034 , w_19035 , \5966_b0 );
or ( \5968_b1 , \5928_b1 , \5952_b1 );
xor ( \5968_b0 , \5928_b0 , w_19036 );
not ( w_19036 , w_19037 );
and ( w_19037 , \5952_b1 , \5952_b0 );
buf ( \5969_b1 , \5939_b1 );
not ( \5969_b1 , w_19038 );
not ( \5969_b0 , w_19039 );
and ( w_19038 , w_19039 , \5939_b0 );
or ( \5970_b1 , \5968_b1 , \5969_b1 );
not ( \5969_b1 , w_19040 );
and ( \5970_b0 , \5968_b0 , w_19041 );
and ( w_19040 , w_19041 , \5969_b0 );
buf ( \5971_b1 , \5968_b1 );
not ( \5971_b1 , w_19042 );
not ( \5971_b0 , w_19043 );
and ( w_19042 , w_19043 , \5968_b0 );
or ( \5972_b1 , \5971_b1 , \5939_b1 );
not ( \5939_b1 , w_19044 );
and ( \5972_b0 , \5971_b0 , w_19045 );
and ( w_19044 , w_19045 , \5939_b0 );
or ( \5973_b1 , \5970_b1 , w_19047 );
not ( w_19047 , w_19048 );
and ( \5973_b0 , \5970_b0 , w_19049 );
and ( w_19048 ,  , w_19049 );
buf ( w_19047 , \5972_b1 );
not ( w_19047 , w_19050 );
not (  , w_19051 );
and ( w_19050 , w_19051 , \5972_b0 );
or ( \5974_b1 , \5709_b1 , \5714_b1 );
xor ( \5974_b0 , \5709_b0 , w_19052 );
not ( w_19052 , w_19053 );
and ( w_19053 , \5714_b1 , \5714_b0 );
or ( \5975_b1 , \5974_b1 , \5726_b1 );
xor ( \5975_b0 , \5974_b0 , w_19054 );
not ( w_19054 , w_19055 );
and ( w_19055 , \5726_b1 , \5726_b0 );
or ( \5976_b1 , \5973_b1 , w_19057 );
not ( w_19057 , w_19058 );
and ( \5976_b0 , \5973_b0 , w_19059 );
and ( w_19058 ,  , w_19059 );
buf ( w_19057 , \5975_b1 );
not ( w_19057 , w_19060 );
not (  , w_19061 );
and ( w_19060 , w_19061 , \5975_b0 );
buf ( \5977_b1 , \5847_b1 );
not ( \5977_b1 , w_19062 );
not ( \5977_b0 , w_19063 );
and ( w_19062 , w_19063 , \5847_b0 );
buf ( \5978_b1 , \4086_b1 );
not ( \5978_b1 , w_19064 );
not ( \5978_b0 , w_19065 );
and ( w_19064 , w_19065 , \4086_b0 );
or ( \5979_b1 , \5977_b1 , w_19066 );
or ( \5979_b0 , \5977_b0 , \5978_b0 );
not ( \5978_b0 , w_19067 );
and ( w_19067 , w_19066 , \5978_b1 );
or ( \5980_b1 , \4596_b1 , w_19069 );
not ( w_19069 , w_19070 );
and ( \5980_b0 , \4596_b0 , w_19071 );
and ( w_19070 ,  , w_19071 );
buf ( w_19069 , \5934_b1 );
not ( w_19069 , w_19072 );
not (  , w_19073 );
and ( w_19072 , w_19073 , \5934_b0 );
or ( \5981_b1 , \5979_b1 , w_19075 );
not ( w_19075 , w_19076 );
and ( \5981_b0 , \5979_b0 , w_19077 );
and ( w_19076 ,  , w_19077 );
buf ( w_19075 , \5980_b1 );
not ( w_19075 , w_19078 );
not (  , w_19079 );
and ( w_19078 , w_19079 , \5980_b0 );
buf ( \5982_b1 , \5981_b1 );
not ( \5982_b1 , w_19080 );
not ( \5982_b0 , w_19081 );
and ( w_19080 , w_19081 , \5981_b0 );
buf ( \5983_b1 , \4425_b1 );
not ( \5983_b1 , w_19082 );
not ( \5983_b0 , w_19083 );
and ( w_19082 , w_19083 , \4425_b0 );
buf ( \5984_b1 , \5897_b1 );
not ( \5984_b1 , w_19084 );
not ( \5984_b0 , w_19085 );
and ( w_19084 , w_19085 , \5897_b0 );
or ( \5985_b1 , \5983_b1 , w_19086 );
or ( \5985_b0 , \5983_b0 , \5984_b0 );
not ( \5984_b0 , w_19087 );
and ( w_19087 , w_19086 , \5984_b1 );
or ( \5986_b1 , \4140_b1 , w_19089 );
not ( w_19089 , w_19090 );
and ( \5986_b0 , \4140_b0 , w_19091 );
and ( w_19090 ,  , w_19091 );
buf ( w_19089 , \5947_b1 );
not ( w_19089 , w_19092 );
not (  , w_19093 );
and ( w_19092 , w_19093 , \5947_b0 );
or ( \5987_b1 , \5985_b1 , w_19095 );
not ( w_19095 , w_19096 );
and ( \5987_b0 , \5985_b0 , w_19097 );
and ( w_19096 ,  , w_19097 );
buf ( w_19095 , \5986_b1 );
not ( w_19095 , w_19098 );
not (  , w_19099 );
and ( w_19098 , w_19099 , \5986_b0 );
buf ( \5988_b1 , \5987_b1 );
not ( \5988_b1 , w_19100 );
not ( \5988_b0 , w_19101 );
and ( w_19100 , w_19101 , \5987_b0 );
or ( \5989_b1 , \5982_b1 , w_19102 );
or ( \5989_b0 , \5982_b0 , \5988_b0 );
not ( \5988_b0 , w_19103 );
and ( w_19103 , w_19102 , \5988_b1 );
or ( \5990_b1 , \5981_b1 , w_19104 );
or ( \5990_b0 , \5981_b0 , \5987_b0 );
not ( \5987_b0 , w_19105 );
and ( w_19105 , w_19104 , \5987_b1 );
buf ( \5991_b1 , \5863_b1 );
not ( \5991_b1 , w_19106 );
not ( \5991_b0 , w_19107 );
and ( w_19106 , w_19107 , \5863_b0 );
buf ( \5992_b1 , \4662_b1 );
not ( \5992_b1 , w_19108 );
not ( \5992_b0 , w_19109 );
and ( w_19108 , w_19109 , \4662_b0 );
or ( \5993_b1 , \5991_b1 , w_19110 );
or ( \5993_b0 , \5991_b0 , \5992_b0 );
not ( \5992_b0 , w_19111 );
and ( w_19111 , w_19110 , \5992_b1 );
or ( \5994_b1 , \4672_b1 , w_19113 );
not ( w_19113 , w_19114 );
and ( \5994_b0 , \4672_b0 , w_19115 );
and ( w_19114 ,  , w_19115 );
buf ( w_19113 , \5721_b1 );
not ( w_19113 , w_19116 );
not (  , w_19117 );
and ( w_19116 , w_19117 , \5721_b0 );
or ( \5995_b1 , \5993_b1 , w_19119 );
not ( w_19119 , w_19120 );
and ( \5995_b0 , \5993_b0 , w_19121 );
and ( w_19120 ,  , w_19121 );
buf ( w_19119 , \5994_b1 );
not ( w_19119 , w_19122 );
not (  , w_19123 );
and ( w_19122 , w_19123 , \5994_b0 );
or ( \5996_b1 , \5990_b1 , w_19125 );
not ( w_19125 , w_19126 );
and ( \5996_b0 , \5990_b0 , w_19127 );
and ( w_19126 ,  , w_19127 );
buf ( w_19125 , \5995_b1 );
not ( w_19125 , w_19128 );
not (  , w_19129 );
and ( w_19128 , w_19129 , \5995_b0 );
or ( \5997_b1 , \5989_b1 , w_19131 );
not ( w_19131 , w_19132 );
and ( \5997_b0 , \5989_b0 , w_19133 );
and ( w_19132 ,  , w_19133 );
buf ( w_19131 , \5996_b1 );
not ( w_19131 , w_19134 );
not (  , w_19135 );
and ( w_19134 , w_19135 , \5996_b0 );
or ( \5998_b1 , \5976_b1 , \5997_b1 );
not ( \5997_b1 , w_19136 );
and ( \5998_b0 , \5976_b0 , w_19137 );
and ( w_19136 , w_19137 , \5997_b0 );
or ( \5999_b1 , \5973_b1 , w_19139 );
not ( w_19139 , w_19140 );
and ( \5999_b0 , \5973_b0 , w_19141 );
and ( w_19140 ,  , w_19141 );
buf ( w_19139 , \5975_b1 );
not ( w_19139 , w_19142 );
not (  , w_19143 );
and ( w_19142 , w_19143 , \5975_b0 );
or ( \6000_b1 , \5998_b1 , w_19145 );
not ( w_19145 , w_19146 );
and ( \6000_b0 , \5998_b0 , w_19147 );
and ( w_19146 ,  , w_19147 );
buf ( w_19145 , \5999_b1 );
not ( w_19145 , w_19148 );
not (  , w_19149 );
and ( w_19148 , w_19149 , \5999_b0 );
buf ( \6001_b1 , \6000_b1 );
not ( \6001_b1 , w_19150 );
not ( \6001_b0 , w_19151 );
and ( w_19150 , w_19151 , \6000_b0 );
buf ( \6002_b1 , \6001_b1 );
not ( \6002_b1 , w_19152 );
not ( \6002_b0 , w_19153 );
and ( w_19152 , w_19153 , \6001_b0 );
or ( \6003_b1 , \5815_b1 , \5821_b1 );
xor ( \6003_b0 , \5815_b0 , w_19154 );
not ( w_19154 , w_19155 );
and ( w_19155 , \5821_b1 , \5821_b0 );
or ( \6004_b1 , \6003_b1 , \5829_b1 );
not ( \5829_b1 , w_19156 );
and ( \6004_b0 , \6003_b0 , w_19157 );
and ( w_19156 , w_19157 , \5829_b0 );
or ( \6005_b1 , \5815_b1 , \5821_b1 );
not ( \5821_b1 , w_19158 );
and ( \6005_b0 , \5815_b0 , w_19159 );
and ( w_19158 , w_19159 , \5821_b0 );
or ( \6006_b1 , \6004_b1 , w_19160 );
or ( \6006_b0 , \6004_b0 , \6005_b0 );
not ( \6005_b0 , w_19161 );
and ( w_19161 , w_19160 , \6005_b1 );
buf ( \6007_b1 , \6006_b1 );
not ( \6007_b1 , w_19162 );
not ( \6007_b0 , w_19163 );
and ( w_19162 , w_19163 , \6006_b0 );
or ( \6008_b1 , \5699_b1 , \5700_b1 );
xor ( \6008_b0 , \5699_b0 , w_19164 );
not ( w_19164 , w_19165 );
and ( w_19165 , \5700_b1 , \5700_b0 );
or ( \6009_b1 , \6008_b1 , \5729_b1 );
xor ( \6009_b0 , \6008_b0 , w_19166 );
not ( w_19166 , w_19167 );
and ( w_19167 , \5729_b1 , \5729_b0 );
buf ( \6010_b1 , \6009_b1 );
not ( \6010_b1 , w_19168 );
not ( \6010_b0 , w_19169 );
and ( w_19168 , w_19169 , \6009_b0 );
or ( \6011_b1 , \6007_b1 , w_19170 );
or ( \6011_b0 , \6007_b0 , \6010_b0 );
not ( \6010_b0 , w_19171 );
and ( w_19171 , w_19170 , \6010_b1 );
or ( \6012_b1 , \6009_b1 , w_19172 );
or ( \6012_b0 , \6009_b0 , \6006_b0 );
not ( \6006_b0 , w_19173 );
and ( w_19173 , w_19172 , \6006_b1 );
or ( \6013_b1 , \6011_b1 , w_19175 );
not ( w_19175 , w_19176 );
and ( \6013_b0 , \6011_b0 , w_19177 );
and ( w_19176 ,  , w_19177 );
buf ( w_19175 , \6012_b1 );
not ( w_19175 , w_19178 );
not (  , w_19179 );
and ( w_19178 , w_19179 , \6012_b0 );
buf ( \6014_b1 , \6013_b1 );
not ( \6014_b1 , w_19180 );
not ( \6014_b0 , w_19181 );
and ( w_19180 , w_19181 , \6013_b0 );
buf ( \6015_b1 , \6014_b1 );
not ( \6015_b1 , w_19182 );
not ( \6015_b0 , w_19183 );
and ( w_19182 , w_19183 , \6014_b0 );
or ( \6016_b1 , \6002_b1 , w_19184 );
or ( \6016_b0 , \6002_b0 , \6015_b0 );
not ( \6015_b0 , w_19185 );
and ( w_19185 , w_19184 , \6015_b1 );
or ( \6017_b1 , \6013_b1 , w_19187 );
not ( w_19187 , w_19188 );
and ( \6017_b0 , \6013_b0 , w_19189 );
and ( w_19188 ,  , w_19189 );
buf ( w_19187 , \6000_b1 );
not ( w_19187 , w_19190 );
not (  , w_19191 );
and ( w_19190 , w_19191 , \6000_b0 );
or ( \6018_b1 , \6016_b1 , w_19193 );
not ( w_19193 , w_19194 );
and ( \6018_b0 , \6016_b0 , w_19195 );
and ( w_19194 ,  , w_19195 );
buf ( w_19193 , \6017_b1 );
not ( w_19193 , w_19196 );
not (  , w_19197 );
and ( w_19196 , w_19197 , \6017_b0 );
buf ( \6019_b1 , \6018_b1 );
not ( \6019_b1 , w_19198 );
not ( \6019_b0 , w_19199 );
and ( w_19198 , w_19199 , \6018_b0 );
or ( \6020_b1 , \5967_b1 , \6019_b1 );
not ( \6019_b1 , w_19200 );
and ( \6020_b0 , \5967_b0 , w_19201 );
and ( w_19200 , w_19201 , \6019_b0 );
buf ( \6021_b1 , \5967_b1 );
not ( \6021_b1 , w_19202 );
not ( \6021_b0 , w_19203 );
and ( w_19202 , w_19203 , \5967_b0 );
or ( \6022_b1 , \6021_b1 , \6018_b1 );
not ( \6018_b1 , w_19204 );
and ( \6022_b0 , \6021_b0 , w_19205 );
and ( w_19204 , w_19205 , \6018_b0 );
or ( \6023_b1 , \6020_b1 , w_19207 );
not ( w_19207 , w_19208 );
and ( \6023_b0 , \6020_b0 , w_19209 );
and ( w_19208 ,  , w_19209 );
buf ( w_19207 , \6022_b1 );
not ( w_19207 , w_19210 );
not (  , w_19211 );
and ( w_19210 , w_19211 , \6022_b0 );
buf ( \6024_b1 , \5795_b1 );
not ( \6024_b1 , w_19212 );
not ( \6024_b0 , w_19213 );
and ( w_19212 , w_19213 , \5795_b0 );
buf ( \6025_b1 , \5830_b1 );
not ( \6025_b1 , w_19214 );
not ( \6025_b0 , w_19215 );
and ( w_19214 , w_19215 , \5830_b0 );
or ( \6026_b1 , \6024_b1 , w_19216 );
or ( \6026_b0 , \6024_b0 , \6025_b0 );
not ( \6025_b0 , w_19217 );
and ( w_19217 , w_19216 , \6025_b1 );
or ( \6027_b1 , \5795_b1 , w_19218 );
or ( \6027_b0 , \5795_b0 , \5830_b0 );
not ( \5830_b0 , w_19219 );
and ( w_19219 , w_19218 , \5830_b1 );
or ( \6028_b1 , \6026_b1 , w_19221 );
not ( w_19221 , w_19222 );
and ( \6028_b0 , \6026_b0 , w_19223 );
and ( w_19222 ,  , w_19223 );
buf ( w_19221 , \6027_b1 );
not ( w_19221 , w_19224 );
not (  , w_19225 );
and ( w_19224 , w_19225 , \6027_b0 );
or ( \6029_b1 , \6028_b1 , \5918_b1 );
xor ( \6029_b0 , \6028_b0 , w_19226 );
not ( w_19226 , w_19227 );
and ( w_19227 , \5918_b1 , \5918_b0 );
buf ( \6030_b1 , \5975_b1 );
not ( \6030_b1 , w_19228 );
not ( \6030_b0 , w_19229 );
and ( w_19228 , w_19229 , \5975_b0 );
buf ( \6031_b1 , \5997_b1 );
not ( \6031_b1 , w_19230 );
not ( \6031_b0 , w_19231 );
and ( w_19230 , w_19231 , \5997_b0 );
or ( \6032_b1 , \6030_b1 , w_19232 );
or ( \6032_b0 , \6030_b0 , \6031_b0 );
not ( \6031_b0 , w_19233 );
and ( w_19233 , w_19232 , \6031_b1 );
or ( \6033_b1 , \5997_b1 , w_19234 );
or ( \6033_b0 , \5997_b0 , \5975_b0 );
not ( \5975_b0 , w_19235 );
and ( w_19235 , w_19234 , \5975_b1 );
or ( \6034_b1 , \6032_b1 , w_19237 );
not ( w_19237 , w_19238 );
and ( \6034_b0 , \6032_b0 , w_19239 );
and ( w_19238 ,  , w_19239 );
buf ( w_19237 , \6033_b1 );
not ( w_19237 , w_19240 );
not (  , w_19241 );
and ( w_19240 , w_19241 , \6033_b0 );
buf ( \6035_b1 , \5973_b1 );
not ( \6035_b1 , w_19242 );
not ( \6035_b0 , w_19243 );
and ( w_19242 , w_19243 , \5973_b0 );
or ( \6036_b1 , \6034_b1 , \6035_b1 );
not ( \6035_b1 , w_19244 );
and ( \6036_b0 , \6034_b0 , w_19245 );
and ( w_19244 , w_19245 , \6035_b0 );
buf ( \6037_b1 , \6034_b1 );
not ( \6037_b1 , w_19246 );
not ( \6037_b0 , w_19247 );
and ( w_19246 , w_19247 , \6034_b0 );
or ( \6038_b1 , \6037_b1 , \5973_b1 );
not ( \5973_b1 , w_19248 );
and ( \6038_b0 , \6037_b0 , w_19249 );
and ( w_19248 , w_19249 , \5973_b0 );
or ( \6039_b1 , \6036_b1 , w_19251 );
not ( w_19251 , w_19252 );
and ( \6039_b0 , \6036_b0 , w_19253 );
and ( w_19252 ,  , w_19253 );
buf ( w_19251 , \6038_b1 );
not ( w_19251 , w_19254 );
not (  , w_19255 );
and ( w_19254 , w_19255 , \6038_b0 );
or ( \6040_b1 , \6029_b1 , w_19256 );
or ( \6040_b0 , \6029_b0 , \6039_b0 );
not ( \6039_b0 , w_19257 );
and ( w_19257 , w_19256 , \6039_b1 );
or ( \6041_b1 , \5761_b1 , \5776_b1 );
xor ( \6041_b0 , \5761_b0 , w_19258 );
not ( w_19258 , w_19259 );
and ( w_19259 , \5776_b1 , \5776_b0 );
or ( \6042_b1 , \6041_b1 , \5792_b1 );
xor ( \6042_b0 , \6041_b0 , w_19260 );
not ( w_19260 , w_19261 );
and ( w_19261 , \5792_b1 , \5792_b0 );
buf ( \6043_b1 , \6042_b1 );
not ( \6043_b1 , w_19262 );
not ( \6043_b0 , w_19263 );
and ( w_19262 , w_19263 , \6042_b0 );
or ( \6044_b1 , \5995_b1 , \5987_b1 );
not ( \5987_b1 , w_19264 );
and ( \6044_b0 , \5995_b0 , w_19265 );
and ( w_19264 , w_19265 , \5987_b0 );
buf ( \6045_b1 , \5995_b1 );
not ( \6045_b1 , w_19266 );
not ( \6045_b0 , w_19267 );
and ( w_19266 , w_19267 , \5995_b0 );
buf ( \6046_b1 , \5987_b1 );
not ( \6046_b1 , w_19268 );
not ( \6046_b0 , w_19269 );
and ( w_19268 , w_19269 , \5987_b0 );
or ( \6047_b1 , \6045_b1 , \6046_b1 );
not ( \6046_b1 , w_19270 );
and ( \6047_b0 , \6045_b0 , w_19271 );
and ( w_19270 , w_19271 , \6046_b0 );
or ( \6048_b1 , \6044_b1 , w_19273 );
not ( w_19273 , w_19274 );
and ( \6048_b0 , \6044_b0 , w_19275 );
and ( w_19274 ,  , w_19275 );
buf ( w_19273 , \6047_b1 );
not ( w_19273 , w_19276 );
not (  , w_19277 );
and ( w_19276 , w_19277 , \6047_b0 );
buf ( \6049_b1 , \5981_b1 );
not ( \6049_b1 , w_19278 );
not ( \6049_b0 , w_19279 );
and ( w_19278 , w_19279 , \5981_b0 );
or ( \6050_b1 , \6048_b1 , \6049_b1 );
not ( \6049_b1 , w_19280 );
and ( \6050_b0 , \6048_b0 , w_19281 );
and ( w_19280 , w_19281 , \6049_b0 );
buf ( \6051_b1 , \6048_b1 );
not ( \6051_b1 , w_19282 );
not ( \6051_b0 , w_19283 );
and ( w_19282 , w_19283 , \6048_b0 );
or ( \6052_b1 , \6051_b1 , \5981_b1 );
not ( \5981_b1 , w_19284 );
and ( \6052_b0 , \6051_b0 , w_19285 );
and ( w_19284 , w_19285 , \5981_b0 );
or ( \6053_b1 , \6050_b1 , w_19287 );
not ( w_19287 , w_19288 );
and ( \6053_b0 , \6050_b0 , w_19289 );
and ( w_19288 ,  , w_19289 );
buf ( w_19287 , \6052_b1 );
not ( w_19287 , w_19290 );
not (  , w_19291 );
and ( w_19290 , w_19291 , \6052_b0 );
buf ( \6054_b1 , \6053_b1 );
buf ( \6054_b0 , \6053_b0 );
or ( \6055_b1 , \6043_b1 , w_19293 );
not ( w_19293 , w_19294 );
and ( \6055_b0 , \6043_b0 , w_19295 );
and ( w_19294 ,  , w_19295 );
buf ( w_19293 , \6054_b1 );
not ( w_19293 , w_19296 );
not (  , w_19297 );
and ( w_19296 , w_19297 , \6054_b0 );
buf ( \6056_b1 , \6055_b1 );
not ( \6056_b1 , w_19298 );
not ( \6056_b0 , w_19299 );
and ( w_19298 , w_19299 , \6055_b0 );
or ( \6057_b1 , \4029_b1 , \4177_b1 );
not ( \4177_b1 , w_19300 );
and ( \6057_b0 , \4029_b0 , w_19301 );
and ( w_19300 , w_19301 , \4177_b0 );
buf ( \6058_b1 , \4029_b1 );
not ( \6058_b1 , w_19302 );
not ( \6058_b0 , w_19303 );
and ( w_19302 , w_19303 , \4029_b0 );
or ( \6059_b1 , \6058_b1 , \4176_b1 );
not ( \4176_b1 , w_19304 );
and ( \6059_b0 , \6058_b0 , w_19305 );
and ( w_19304 , w_19305 , \4176_b0 );
or ( \6060_b1 , \6057_b1 , w_19307 );
not ( w_19307 , w_19308 );
and ( \6060_b0 , \6057_b0 , w_19309 );
and ( w_19308 ,  , w_19309 );
buf ( w_19307 , \6059_b1 );
not ( w_19307 , w_19310 );
not (  , w_19311 );
and ( w_19310 , w_19311 , \6059_b0 );
buf ( \6061_b1 , \6060_b1 );
not ( \6061_b1 , w_19312 );
not ( \6061_b0 , w_19313 );
and ( w_19312 , w_19313 , \6060_b0 );
buf ( \6062_b1 , \4195_b1 );
not ( \6062_b1 , w_19314 );
not ( \6062_b0 , w_19315 );
and ( w_19314 , w_19315 , \4195_b0 );
or ( \6063_b1 , \6061_b1 , w_19316 );
or ( \6063_b0 , \6061_b0 , \6062_b0 );
not ( \6062_b0 , w_19317 );
and ( w_19317 , w_19316 , \6062_b1 );
or ( \6064_b1 , \5111_b1 , w_19319 );
not ( w_19319 , w_19320 );
and ( \6064_b0 , \5111_b0 , w_19321 );
and ( w_19320 ,  , w_19321 );
buf ( w_19319 , \5782_b1 );
not ( w_19319 , w_19322 );
not (  , w_19323 );
and ( w_19322 , w_19323 , \5782_b0 );
or ( \6065_b1 , \6063_b1 , w_19325 );
not ( w_19325 , w_19326 );
and ( \6065_b0 , \6063_b0 , w_19327 );
and ( w_19326 ,  , w_19327 );
buf ( w_19325 , \6064_b1 );
not ( w_19325 , w_19328 );
not (  , w_19329 );
and ( w_19328 , w_19329 , \6064_b0 );
buf ( \6066_b1 , \5388_b1 );
not ( \6066_b1 , w_19330 );
not ( \6066_b0 , w_19331 );
and ( w_19330 , w_19331 , \5388_b0 );
buf ( \6067_b1 , \4190_b1 );
not ( \6067_b1 , w_19332 );
not ( \6067_b0 , w_19333 );
and ( w_19332 , w_19333 , \4190_b0 );
or ( \6068_b1 , \6066_b1 , w_19334 );
or ( \6068_b0 , \6066_b0 , \6067_b0 );
not ( \6067_b0 , w_19335 );
and ( w_19335 , w_19334 , \6067_b1 );
or ( \6069_b1 , \6068_b1 , w_19337 );
not ( w_19337 , w_19338 );
and ( \6069_b0 , \6068_b0 , w_19339 );
and ( w_19338 ,  , w_19339 );
buf ( w_19337 , \4368_b1 );
not ( w_19337 , w_19340 );
not (  , w_19341 );
and ( w_19340 , w_19341 , \4368_b0 );
or ( \6070_b1 , \3487_b1 , w_19343 );
not ( w_19343 , w_19344 );
and ( \6070_b0 , \3487_b0 , w_19345 );
and ( w_19344 ,  , w_19345 );
buf ( w_19343 , \4048_b1 );
not ( w_19343 , w_19346 );
not (  , w_19347 );
and ( w_19346 , w_19347 , \4048_b0 );
buf ( \6072_b1 , \4011_b1 );
not ( \6072_b1 , w_19348 );
not ( \6072_b0 , w_19349 );
and ( w_19348 , w_19349 , \4011_b0 );
buf ( \6073_b1 , \5178_b1 );
not ( \6073_b1 , w_19350 );
not ( \6073_b0 , w_19351 );
and ( w_19350 , w_19351 , \5178_b0 );
or ( \6074_b1 , \6072_b1 , w_19352 );
or ( \6074_b0 , \6072_b0 , \6073_b0 );
not ( \6073_b0 , w_19353 );
and ( w_19353 , w_19352 , \6073_b1 );
or ( \6075_b1 , \4665_b1 , w_19355 );
not ( w_19355 , w_19356 );
and ( \6075_b0 , \4665_b0 , w_19357 );
and ( w_19356 ,  , w_19357 );
buf ( w_19355 , \4270_b1 );
not ( w_19355 , w_19358 );
not (  , w_19359 );
and ( w_19358 , w_19359 , \4270_b0 );
or ( \6076_b1 , \6074_b1 , w_19361 );
not ( w_19361 , w_19362 );
and ( \6076_b0 , \6074_b0 , w_19363 );
and ( w_19362 ,  , w_19363 );
buf ( w_19361 , \6075_b1 );
not ( w_19361 , w_19364 );
not (  , w_19365 );
and ( w_19364 , w_19365 , \6075_b0 );
buf ( \6077_b1 , \6076_b1 );
not ( \6077_b1 , w_19366 );
not ( \6077_b0 , w_19367 );
and ( w_19366 , w_19367 , \6076_b0 );
buf ( \6078_b1 , \4662_b1 );
not ( \6078_b1 , w_19368 );
not ( \6078_b0 , w_19369 );
and ( w_19368 , w_19369 , \4662_b0 );
or ( \6079_b1 , \6077_b1 , w_19370 );
or ( \6079_b0 , \6077_b0 , \6078_b0 );
not ( \6078_b0 , w_19371 );
and ( w_19371 , w_19370 , \6078_b1 );
or ( \6080_b1 , \4672_b1 , w_19373 );
not ( w_19373 , w_19374 );
and ( \6080_b0 , \4672_b0 , w_19375 );
and ( w_19374 ,  , w_19375 );
buf ( w_19373 , \5855_b1 );
not ( w_19373 , w_19376 );
not (  , w_19377 );
and ( w_19376 , w_19377 , \5855_b0 );
or ( \6081_b1 , \6079_b1 , w_19379 );
not ( w_19379 , w_19380 );
and ( \6081_b0 , \6079_b0 , w_19381 );
and ( w_19380 ,  , w_19381 );
buf ( w_19379 , \6080_b1 );
not ( w_19379 , w_19382 );
not (  , w_19383 );
and ( w_19382 , w_19383 , \6080_b0 );
or ( \6082_b1 , \6071_b1 , \6081_b1 );
not ( \6081_b1 , w_19384 );
and ( \6082_b0 , \6071_b0 , w_19385 );
and ( w_19384 , w_19385 , \6081_b0 );
or ( \6083_b1 , \6065_b1 , \6082_b1 );
xor ( \6083_b0 , \6065_b0 , w_19386 );
not ( w_19386 , w_19387 );
and ( w_19387 , \6082_b1 , \6082_b0 );
or ( \6084_b1 , \4238_b1 , \5873_b1 );
not ( \5873_b1 , w_19388 );
and ( \6084_b0 , \4238_b0 , w_19389 );
and ( w_19388 , w_19389 , \5873_b0 );
buf ( \6085_b1 , \4238_b1 );
not ( \6085_b1 , w_19390 );
not ( \6085_b0 , w_19391 );
and ( w_19390 , w_19391 , \4238_b0 );
or ( \6086_b1 , \6085_b1 , \5874_b1 );
not ( \5874_b1 , w_19392 );
and ( \6086_b0 , \6085_b0 , w_19393 );
and ( w_19392 , w_19393 , \5874_b0 );
or ( \6087_b1 , \6084_b1 , w_19395 );
not ( w_19395 , w_19396 );
and ( \6087_b0 , \6084_b0 , w_19397 );
and ( w_19396 ,  , w_19397 );
buf ( w_19395 , \6086_b1 );
not ( w_19395 , w_19398 );
not (  , w_19399 );
and ( w_19398 , w_19399 , \6086_b0 );
buf ( \6088_b1 , \6087_b1 );
not ( \6088_b1 , w_19400 );
not ( \6088_b0 , w_19401 );
and ( w_19400 , w_19401 , \6087_b0 );
buf ( \6089_b1 , \6088_b1 );
not ( \6089_b1 , w_19402 );
not ( \6089_b0 , w_19403 );
and ( w_19402 , w_19403 , \6088_b0 );
buf ( \6090_b1 , \5019_b1 );
not ( \6090_b1 , w_19404 );
not ( \6090_b0 , w_19405 );
and ( w_19404 , w_19405 , \5019_b0 );
or ( \6091_b1 , \6089_b1 , w_19406 );
or ( \6091_b0 , \6089_b0 , \6090_b0 );
not ( \6090_b0 , w_19407 );
and ( w_19407 , w_19406 , \6090_b1 );
or ( \6092_b1 , \5878_b1 , w_19409 );
not ( w_19409 , w_19410 );
and ( \6092_b0 , \5878_b0 , w_19411 );
and ( w_19410 ,  , w_19411 );
buf ( w_19409 , \5021_b1 );
not ( w_19409 , w_19412 );
not (  , w_19413 );
and ( w_19412 , w_19413 , \5021_b0 );
or ( \6093_b1 , \6091_b1 , w_19415 );
not ( w_19415 , w_19416 );
and ( \6093_b0 , \6091_b0 , w_19417 );
and ( w_19416 ,  , w_19417 );
buf ( w_19415 , \6092_b1 );
not ( w_19415 , w_19418 );
not (  , w_19419 );
and ( w_19418 , w_19419 , \6092_b0 );
or ( \6094_b1 , \5344_b1 , \4142_b1 );
not ( \4142_b1 , w_19420 );
and ( \6094_b0 , \5344_b0 , w_19421 );
and ( w_19420 , w_19421 , \4142_b0 );
buf ( \6095_b1 , \5344_b1 );
not ( \6095_b1 , w_19422 );
not ( \6095_b0 , w_19423 );
and ( w_19422 , w_19423 , \5344_b0 );
or ( \6096_b1 , \6095_b1 , \4109_b1 );
not ( \4109_b1 , w_19424 );
and ( \6096_b0 , \6095_b0 , w_19425 );
and ( w_19424 , w_19425 , \4109_b0 );
or ( \6097_b1 , \6094_b1 , w_19427 );
not ( w_19427 , w_19428 );
and ( \6097_b0 , \6094_b0 , w_19429 );
and ( w_19428 ,  , w_19429 );
buf ( w_19427 , \6096_b1 );
not ( w_19427 , w_19430 );
not (  , w_19431 );
and ( w_19430 , w_19431 , \6096_b0 );
buf ( \6098_b1 , \6097_b1 );
not ( \6098_b1 , w_19432 );
not ( \6098_b0 , w_19433 );
and ( w_19432 , w_19433 , \6097_b0 );
buf ( \6099_b1 , \4425_b1 );
not ( \6099_b1 , w_19434 );
not ( \6099_b0 , w_19435 );
and ( w_19434 , w_19435 , \4425_b0 );
or ( \6100_b1 , \6098_b1 , w_19436 );
or ( \6100_b0 , \6098_b0 , \6099_b0 );
not ( \6099_b0 , w_19437 );
and ( w_19437 , w_19436 , \6099_b1 );
or ( \6101_b1 , \4429_b1 , w_19439 );
not ( w_19439 , w_19440 );
and ( \6101_b0 , \4429_b0 , w_19441 );
and ( w_19440 ,  , w_19441 );
buf ( w_19439 , \5889_b1 );
not ( w_19439 , w_19442 );
not (  , w_19443 );
and ( w_19442 , w_19443 , \5889_b0 );
or ( \6102_b1 , \6100_b1 , w_19445 );
not ( w_19445 , w_19446 );
and ( \6102_b0 , \6100_b0 , w_19447 );
and ( w_19446 ,  , w_19447 );
buf ( w_19445 , \6101_b1 );
not ( w_19445 , w_19448 );
not (  , w_19449 );
and ( w_19448 , w_19449 , \6101_b0 );
or ( \6103_b1 , \6093_b1 , \6102_b1 );
xor ( \6103_b0 , \6093_b0 , w_19450 );
not ( w_19450 , w_19451 );
and ( w_19451 , \6102_b1 , \6102_b0 );
or ( \6104_b1 , \4019_b1 , \4088_b1 );
not ( \4088_b1 , w_19452 );
and ( \6104_b0 , \4019_b0 , w_19453 );
and ( w_19452 , w_19453 , \4088_b0 );
buf ( \6105_b1 , \4019_b1 );
not ( \6105_b1 , w_19454 );
not ( \6105_b0 , w_19455 );
and ( w_19454 , w_19455 , \4019_b0 );
or ( \6106_b1 , \6105_b1 , \5234_b1 );
not ( \5234_b1 , w_19456 );
and ( \6106_b0 , \6105_b0 , w_19457 );
and ( w_19456 , w_19457 , \5234_b0 );
or ( \6107_b1 , \6104_b1 , w_19459 );
not ( w_19459 , w_19460 );
and ( \6107_b0 , \6104_b0 , w_19461 );
and ( w_19460 ,  , w_19461 );
buf ( w_19459 , \6106_b1 );
not ( w_19459 , w_19462 );
not (  , w_19463 );
and ( w_19462 , w_19463 , \6106_b0 );
buf ( \6108_b1 , \6107_b1 );
not ( \6108_b1 , w_19464 );
not ( \6108_b0 , w_19465 );
and ( w_19464 , w_19465 , \6107_b0 );
buf ( \6109_b1 , \4437_b1 );
not ( \6109_b1 , w_19466 );
not ( \6109_b0 , w_19467 );
and ( w_19466 , w_19467 , \4437_b0 );
or ( \6110_b1 , \6108_b1 , w_19468 );
or ( \6110_b0 , \6108_b0 , \6109_b0 );
not ( \6109_b0 , w_19469 );
and ( w_19469 , w_19468 , \6109_b1 );
or ( \6111_b1 , \4331_b1 , w_19471 );
not ( w_19471 , w_19472 );
and ( \6111_b0 , \4331_b0 , w_19473 );
and ( w_19472 ,  , w_19473 );
buf ( w_19471 , \5839_b1 );
not ( w_19471 , w_19474 );
not (  , w_19475 );
and ( w_19474 , w_19475 , \5839_b0 );
or ( \6112_b1 , \6110_b1 , w_19477 );
not ( w_19477 , w_19478 );
and ( \6112_b0 , \6110_b0 , w_19479 );
and ( w_19478 ,  , w_19479 );
buf ( w_19477 , \6111_b1 );
not ( w_19477 , w_19480 );
not (  , w_19481 );
and ( w_19480 , w_19481 , \6111_b0 );
or ( \6113_b1 , \6103_b1 , \6112_b1 );
not ( \6112_b1 , w_19482 );
and ( \6113_b0 , \6103_b0 , w_19483 );
and ( w_19482 , w_19483 , \6112_b0 );
or ( \6114_b1 , \6093_b1 , \6102_b1 );
not ( \6102_b1 , w_19484 );
and ( \6114_b0 , \6093_b0 , w_19485 );
and ( w_19484 , w_19485 , \6102_b0 );
or ( \6115_b1 , \6113_b1 , w_19486 );
or ( \6115_b0 , \6113_b0 , \6114_b0 );
not ( \6114_b0 , w_19487 );
and ( w_19487 , w_19486 , \6114_b1 );
or ( \6116_b1 , \6083_b1 , \6115_b1 );
not ( \6115_b1 , w_19488 );
and ( \6116_b0 , \6083_b0 , w_19489 );
and ( w_19488 , w_19489 , \6115_b0 );
or ( \6117_b1 , \6065_b1 , \6082_b1 );
not ( \6082_b1 , w_19490 );
and ( \6117_b0 , \6065_b0 , w_19491 );
and ( w_19490 , w_19491 , \6082_b0 );
or ( \6118_b1 , \6116_b1 , w_19492 );
or ( \6118_b0 , \6116_b0 , \6117_b0 );
not ( \6117_b0 , w_19493 );
and ( w_19493 , w_19492 , \6117_b1 );
buf ( \6119_b1 , \6118_b1 );
not ( \6119_b1 , w_19494 );
not ( \6119_b0 , w_19495 );
and ( w_19494 , w_19495 , \6118_b0 );
or ( \6120_b1 , \6056_b1 , w_19496 );
or ( \6120_b0 , \6056_b0 , \6119_b0 );
not ( \6119_b0 , w_19497 );
and ( w_19497 , w_19496 , \6119_b1 );
buf ( \6121_b1 , \6054_b1 );
not ( \6121_b1 , w_19498 );
not ( \6121_b0 , w_19499 );
and ( w_19498 , w_19499 , \6054_b0 );
or ( \6122_b1 , \6121_b1 , w_19501 );
not ( w_19501 , w_19502 );
and ( \6122_b0 , \6121_b0 , w_19503 );
and ( w_19502 ,  , w_19503 );
buf ( w_19501 , \6042_b1 );
not ( w_19501 , w_19504 );
not (  , w_19505 );
and ( w_19504 , w_19505 , \6042_b0 );
or ( \6123_b1 , \6120_b1 , w_19507 );
not ( w_19507 , w_19508 );
and ( \6123_b0 , \6120_b0 , w_19509 );
and ( w_19508 ,  , w_19509 );
buf ( w_19507 , \6122_b1 );
not ( w_19507 , w_19510 );
not (  , w_19511 );
and ( w_19510 , w_19511 , \6122_b0 );
or ( \6124_b1 , \6040_b1 , \6123_b1 );
not ( \6123_b1 , w_19512 );
and ( \6124_b0 , \6040_b0 , w_19513 );
and ( w_19512 , w_19513 , \6123_b0 );
or ( \6125_b1 , \6039_b1 , \6029_b1 );
not ( \6029_b1 , w_19514 );
and ( \6125_b0 , \6039_b0 , w_19515 );
and ( w_19514 , w_19515 , \6029_b0 );
or ( \6126_b1 , \6124_b1 , w_19517 );
not ( w_19517 , w_19518 );
and ( \6126_b0 , \6124_b0 , w_19519 );
and ( w_19518 ,  , w_19519 );
buf ( w_19517 , \6125_b1 );
not ( w_19517 , w_19520 );
not (  , w_19521 );
and ( w_19520 , w_19521 , \6125_b0 );
or ( \6127_b1 , \6023_b1 , w_19523 );
not ( w_19523 , w_19524 );
and ( \6127_b0 , \6023_b0 , w_19525 );
and ( w_19524 ,  , w_19525 );
buf ( w_19523 , \6126_b1 );
not ( w_19523 , w_19526 );
not (  , w_19527 );
and ( w_19526 , w_19527 , \6126_b0 );
or ( \6128_b1 , \6039_b1 , \6029_b1 );
xor ( \6128_b0 , \6039_b0 , w_19528 );
not ( w_19528 , w_19529 );
and ( w_19529 , \6029_b1 , \6029_b0 );
buf ( \6129_b1 , \6123_b1 );
not ( \6129_b1 , w_19530 );
not ( \6129_b0 , w_19531 );
and ( w_19530 , w_19531 , \6123_b0 );
or ( \6130_b1 , \6128_b1 , \6129_b1 );
not ( \6129_b1 , w_19532 );
and ( \6130_b0 , \6128_b0 , w_19533 );
and ( w_19532 , w_19533 , \6129_b0 );
buf ( \6131_b1 , \6128_b1 );
not ( \6131_b1 , w_19534 );
not ( \6131_b0 , w_19535 );
and ( w_19534 , w_19535 , \6128_b0 );
or ( \6132_b1 , \6131_b1 , \6123_b1 );
not ( \6123_b1 , w_19536 );
and ( \6132_b0 , \6131_b0 , w_19537 );
and ( w_19536 , w_19537 , \6123_b0 );
or ( \6133_b1 , \6130_b1 , w_19539 );
not ( w_19539 , w_19540 );
and ( \6133_b0 , \6130_b0 , w_19541 );
and ( w_19540 ,  , w_19541 );
buf ( w_19539 , \6132_b1 );
not ( w_19539 , w_19542 );
not (  , w_19543 );
and ( w_19542 , w_19543 , \6132_b0 );
or ( \6134_b1 , \5833_b1 , \5870_b1 );
xor ( \6134_b0 , \5833_b0 , w_19544 );
not ( w_19544 , w_19545 );
and ( w_19545 , \5870_b1 , \5870_b0 );
or ( \6135_b1 , \6134_b1 , \5915_b1 );
xor ( \6135_b0 , \6134_b0 , w_19546 );
not ( w_19546 , w_19547 );
and ( w_19547 , \5915_b1 , \5915_b0 );
buf ( \6136_b1 , \6135_b1 );
not ( \6136_b1 , w_19548 );
not ( \6136_b0 , w_19549 );
and ( w_19548 , w_19549 , \6135_b0 );
buf ( \6137_b1 , \6042_b1 );
not ( \6137_b1 , w_19550 );
not ( \6137_b0 , w_19551 );
and ( w_19550 , w_19551 , \6042_b0 );
buf ( \6138_b1 , \6053_b1 );
not ( \6138_b1 , w_19552 );
not ( \6138_b0 , w_19553 );
and ( w_19552 , w_19553 , \6053_b0 );
or ( \6139_b1 , \6137_b1 , w_19554 );
or ( \6139_b0 , \6137_b0 , \6138_b0 );
not ( \6138_b0 , w_19555 );
and ( w_19555 , w_19554 , \6138_b1 );
or ( \6140_b1 , \6053_b1 , w_19556 );
or ( \6140_b0 , \6053_b0 , \6042_b0 );
not ( \6042_b0 , w_19557 );
and ( w_19557 , w_19556 , \6042_b1 );
or ( \6141_b1 , \6139_b1 , w_19559 );
not ( w_19559 , w_19560 );
and ( \6141_b0 , \6139_b0 , w_19561 );
and ( w_19560 ,  , w_19561 );
buf ( w_19559 , \6140_b1 );
not ( w_19559 , w_19562 );
not (  , w_19563 );
and ( w_19562 , w_19563 , \6140_b0 );
buf ( \6142_b1 , \6118_b1 );
not ( \6142_b1 , w_19564 );
not ( \6142_b0 , w_19565 );
and ( w_19564 , w_19565 , \6118_b0 );
or ( \6143_b1 , \6141_b1 , \6142_b1 );
not ( \6142_b1 , w_19566 );
and ( \6143_b0 , \6141_b0 , w_19567 );
and ( w_19566 , w_19567 , \6142_b0 );
buf ( \6144_b1 , \6141_b1 );
not ( \6144_b1 , w_19568 );
not ( \6144_b0 , w_19569 );
and ( w_19568 , w_19569 , \6141_b0 );
or ( \6145_b1 , \6144_b1 , \6118_b1 );
not ( \6118_b1 , w_19570 );
and ( \6145_b0 , \6144_b0 , w_19571 );
and ( w_19570 , w_19571 , \6118_b0 );
or ( \6146_b1 , \6143_b1 , w_19573 );
not ( w_19573 , w_19574 );
and ( \6146_b0 , \6143_b0 , w_19575 );
and ( w_19574 ,  , w_19575 );
buf ( w_19573 , \6145_b1 );
not ( w_19573 , w_19576 );
not (  , w_19577 );
and ( w_19576 , w_19577 , \6145_b0 );
or ( \6147_b1 , \6136_b1 , w_19579 );
not ( w_19579 , w_19580 );
and ( \6147_b0 , \6136_b0 , w_19581 );
and ( w_19580 ,  , w_19581 );
buf ( w_19579 , \6146_b1 );
not ( w_19579 , w_19582 );
not (  , w_19583 );
and ( w_19582 , w_19583 , \6146_b0 );
or ( \6148_b1 , \5867_b1 , \5849_b1 );
xor ( \6148_b0 , \5867_b0 , w_19584 );
not ( w_19584 , w_19585 );
and ( w_19585 , \5849_b1 , \5849_b0 );
or ( \6149_b1 , \6148_b1 , \5865_b1 );
xor ( \6149_b0 , \6148_b0 , w_19586 );
not ( w_19586 , w_19587 );
and ( w_19587 , \5865_b1 , \5865_b0 );
buf ( \6150_b1 , \6149_b1 );
not ( \6150_b1 , w_19588 );
not ( \6150_b0 , w_19589 );
and ( w_19588 , w_19589 , \6149_b0 );
or ( \6151_b1 , \5883_b1 , \5899_b1 );
xor ( \6151_b0 , \5883_b0 , w_19590 );
not ( w_19590 , w_19591 );
and ( w_19591 , \5899_b1 , \5899_b0 );
or ( \6152_b1 , \6151_b1 , w_19592 );
xor ( \6152_b0 , \6151_b0 , w_19594 );
not ( w_19594 , w_19595 );
and ( w_19595 , w_19592 , w_19593 );
buf ( w_19592 , \5913_b1 );
not ( w_19592 , w_19596 );
not ( w_19593 , w_19597 );
and ( w_19596 , w_19597 , \5913_b0 );
buf ( \6153_b1 , \6152_b1 );
not ( \6153_b1 , w_19598 );
not ( \6153_b0 , w_19599 );
and ( w_19598 , w_19599 , \6152_b0 );
or ( \6154_b1 , \6150_b1 , w_19600 );
or ( \6154_b0 , \6150_b0 , \6153_b0 );
not ( \6153_b0 , w_19601 );
and ( w_19601 , w_19600 , \6153_b1 );
buf ( \6155_b1 , \3958_b1 );
not ( \6155_b1 , w_19602 );
not ( \6155_b0 , w_19603 );
and ( w_19602 , w_19603 , \3958_b0 );
buf ( \6156_b1 , \4069_b1 );
not ( \6156_b1 , w_19604 );
not ( \6156_b0 , w_19605 );
and ( w_19604 , w_19605 , \4069_b0 );
or ( \6157_b1 , \6155_b1 , w_19606 );
or ( \6157_b0 , \6155_b0 , \6156_b0 );
not ( \6156_b0 , w_19607 );
and ( w_19607 , w_19606 , \6156_b1 );
buf ( \6158_b1 , \5904_b1 );
not ( \6158_b1 , w_19608 );
not ( \6158_b0 , w_19609 );
and ( w_19608 , w_19609 , \5904_b0 );
or ( \6159_b1 , \6158_b1 , w_19611 );
not ( w_19611 , w_19612 );
and ( \6159_b0 , \6158_b0 , w_19613 );
and ( w_19612 ,  , w_19613 );
buf ( w_19611 , \4473_b1 );
not ( w_19611 , w_19614 );
not (  , w_19615 );
and ( w_19614 , w_19615 , \4473_b0 );
or ( \6160_b1 , \6157_b1 , w_19617 );
not ( w_19617 , w_19618 );
and ( \6160_b0 , \6157_b0 , w_19619 );
and ( w_19618 ,  , w_19619 );
buf ( w_19617 , \6159_b1 );
not ( w_19617 , w_19620 );
not (  , w_19621 );
and ( w_19620 , w_19621 , \6159_b0 );
buf ( \6161_b1 , \6160_b1 );
not ( \6161_b1 , w_19622 );
not ( \6161_b0 , w_19623 );
and ( w_19622 , w_19623 , \6160_b0 );
buf ( \6162_b1 , \4411_b1 );
not ( \6162_b1 , w_19624 );
not ( \6162_b0 , w_19625 );
and ( w_19624 , w_19625 , \4411_b0 );
buf ( \6163_b1 , \6162_b1 );
not ( \6163_b1 , w_19626 );
not ( \6163_b0 , w_19627 );
and ( w_19626 , w_19627 , \6162_b0 );
or ( \6164_b1 , \6161_b1 , w_19628 );
or ( \6164_b0 , \6161_b0 , \6163_b0 );
not ( \6163_b0 , w_19629 );
and ( w_19629 , w_19628 , \6163_b1 );
or ( \6165_b1 , \4562_b1 , w_19631 );
not ( w_19631 , w_19632 );
and ( \6165_b0 , \4562_b0 , w_19633 );
and ( w_19632 ,  , w_19633 );
buf ( w_19631 , \5908_b1 );
not ( w_19631 , w_19634 );
not (  , w_19635 );
and ( w_19634 , w_19635 , \5908_b0 );
or ( \6166_b1 , \6164_b1 , w_19637 );
not ( w_19637 , w_19638 );
and ( \6166_b0 , \6164_b0 , w_19639 );
and ( w_19638 ,  , w_19639 );
buf ( w_19637 , \6165_b1 );
not ( w_19637 , w_19640 );
not (  , w_19641 );
and ( w_19640 , w_19641 , \6165_b0 );
buf ( \6167_b1 , \6166_b1 );
not ( \6167_b1 , w_19642 );
not ( \6167_b0 , w_19643 );
and ( w_19642 , w_19643 , \6166_b0 );
or ( \6168_b1 , \4048_b1 , \4177_b1 );
not ( \4177_b1 , w_19644 );
and ( \6168_b0 , \4048_b0 , w_19645 );
and ( w_19644 , w_19645 , \4177_b0 );
buf ( \6169_b1 , \4048_b1 );
not ( \6169_b1 , w_19646 );
not ( \6169_b0 , w_19647 );
and ( w_19646 , w_19647 , \4048_b0 );
or ( \6170_b1 , \6169_b1 , \4284_b1 );
not ( \4284_b1 , w_19648 );
and ( \6170_b0 , \6169_b0 , w_19649 );
and ( w_19648 , w_19649 , \4284_b0 );
or ( \6171_b1 , \6168_b1 , w_19651 );
not ( w_19651 , w_19652 );
and ( \6171_b0 , \6168_b0 , w_19653 );
and ( w_19652 ,  , w_19653 );
buf ( w_19651 , \6170_b1 );
not ( w_19651 , w_19654 );
not (  , w_19655 );
and ( w_19654 , w_19655 , \6170_b0 );
buf ( \6172_b1 , \6171_b1 );
not ( \6172_b1 , w_19656 );
not ( \6172_b0 , w_19657 );
and ( w_19656 , w_19657 , \6171_b0 );
buf ( \6173_b1 , \4194_b1 );
not ( \6173_b1 , w_19658 );
not ( \6173_b0 , w_19659 );
and ( w_19658 , w_19659 , \4194_b0 );
or ( \6174_b1 , \6172_b1 , w_19660 );
or ( \6174_b0 , \6172_b0 , \6173_b0 );
not ( \6173_b0 , w_19661 );
and ( w_19661 , w_19660 , \6173_b1 );
or ( \6175_b1 , \6060_b1 , w_19663 );
not ( w_19663 , w_19664 );
and ( \6175_b0 , \6060_b0 , w_19665 );
and ( w_19664 ,  , w_19665 );
buf ( w_19663 , \5111_b1 );
not ( w_19663 , w_19666 );
not (  , w_19667 );
and ( w_19666 , w_19667 , \5111_b0 );
or ( \6176_b1 , \6174_b1 , w_19669 );
not ( w_19669 , w_19670 );
and ( \6176_b0 , \6174_b0 , w_19671 );
and ( w_19670 ,  , w_19671 );
buf ( w_19669 , \6175_b1 );
not ( w_19669 , w_19672 );
not (  , w_19673 );
and ( w_19672 , w_19673 , \6175_b0 );
buf ( \6177_b1 , \6176_b1 );
not ( \6177_b1 , w_19674 );
not ( \6177_b0 , w_19675 );
and ( w_19674 , w_19675 , \6176_b0 );
or ( \6178_b1 , \6167_b1 , w_19677 );
not ( w_19677 , w_19678 );
and ( \6178_b0 , \6167_b0 , w_19679 );
and ( w_19678 ,  , w_19679 );
buf ( w_19677 , \6177_b1 );
not ( w_19677 , w_19680 );
not (  , w_19681 );
and ( w_19680 , w_19681 , \6177_b0 );
buf ( \6179_b1 , \6178_b1 );
not ( \6179_b1 , w_19682 );
not ( \6179_b0 , w_19683 );
and ( w_19682 , w_19683 , \6178_b0 );
or ( \6180_b1 , \6071_b1 , \6081_b1 );
xor ( \6180_b0 , \6071_b0 , w_19684 );
not ( w_19684 , w_19685 );
and ( w_19685 , \6081_b1 , \6081_b0 );
buf ( \6181_b1 , \6180_b1 );
not ( \6181_b1 , w_19686 );
not ( \6181_b0 , w_19687 );
and ( w_19686 , w_19687 , \6180_b0 );
or ( \6182_b1 , \6179_b1 , w_19688 );
or ( \6182_b0 , \6179_b0 , \6181_b0 );
not ( \6181_b0 , w_19689 );
and ( w_19689 , w_19688 , \6181_b1 );
or ( \6183_b1 , \6166_b1 , w_19691 );
not ( w_19691 , w_19692 );
and ( \6183_b0 , \6166_b0 , w_19693 );
and ( w_19692 ,  , w_19693 );
buf ( w_19691 , \6176_b1 );
not ( w_19691 , w_19694 );
not (  , w_19695 );
and ( w_19694 , w_19695 , \6176_b0 );
or ( \6184_b1 , \6182_b1 , w_19697 );
not ( w_19697 , w_19698 );
and ( \6184_b0 , \6182_b0 , w_19699 );
and ( w_19698 ,  , w_19699 );
buf ( w_19697 , \6183_b1 );
not ( w_19697 , w_19700 );
not (  , w_19701 );
and ( w_19700 , w_19701 , \6183_b0 );
or ( \6185_b1 , \6154_b1 , w_19703 );
not ( w_19703 , w_19704 );
and ( \6185_b0 , \6154_b0 , w_19705 );
and ( w_19704 ,  , w_19705 );
buf ( w_19703 , \6184_b1 );
not ( w_19703 , w_19706 );
not (  , w_19707 );
and ( w_19706 , w_19707 , \6184_b0 );
buf ( \6186_b1 , \6152_b1 );
not ( \6186_b1 , w_19708 );
not ( \6186_b0 , w_19709 );
and ( w_19708 , w_19709 , \6152_b0 );
buf ( \6187_b1 , \6149_b1 );
not ( \6187_b1 , w_19710 );
not ( \6187_b0 , w_19711 );
and ( w_19710 , w_19711 , \6149_b0 );
or ( \6188_b1 , \6186_b1 , w_19713 );
not ( w_19713 , w_19714 );
and ( \6188_b0 , \6186_b0 , w_19715 );
and ( w_19714 ,  , w_19715 );
buf ( w_19713 , \6187_b1 );
not ( w_19713 , w_19716 );
not (  , w_19717 );
and ( w_19716 , w_19717 , \6187_b0 );
or ( \6189_b1 , \6185_b1 , w_19719 );
not ( w_19719 , w_19720 );
and ( \6189_b0 , \6185_b0 , w_19721 );
and ( w_19720 ,  , w_19721 );
buf ( w_19719 , \6188_b1 );
not ( w_19719 , w_19722 );
not (  , w_19723 );
and ( w_19722 , w_19723 , \6188_b0 );
buf ( \6190_b1 , \6189_b1 );
not ( \6190_b1 , w_19724 );
not ( \6190_b0 , w_19725 );
and ( w_19724 , w_19725 , \6189_b0 );
buf ( \6191_b1 , \6190_b1 );
not ( \6191_b1 , w_19726 );
not ( \6191_b0 , w_19727 );
and ( w_19726 , w_19727 , \6190_b0 );
or ( \6192_b1 , \6147_b1 , \6191_b1 );
not ( \6191_b1 , w_19728 );
and ( \6192_b0 , \6147_b0 , w_19729 );
and ( w_19728 , w_19729 , \6191_b0 );
buf ( \6193_b1 , \6135_b1 );
not ( \6193_b1 , w_19730 );
not ( \6193_b0 , w_19731 );
and ( w_19730 , w_19731 , \6135_b0 );
or ( \6194_b1 , \6193_b1 , w_19733 );
not ( w_19733 , w_19734 );
and ( \6194_b0 , \6193_b0 , w_19735 );
and ( w_19734 ,  , w_19735 );
buf ( w_19733 , \6146_b1 );
not ( w_19733 , w_19736 );
not (  , w_19737 );
and ( w_19736 , w_19737 , \6146_b0 );
or ( \6195_b1 , \6192_b1 , w_19739 );
not ( w_19739 , w_19740 );
and ( \6195_b0 , \6192_b0 , w_19741 );
and ( w_19740 ,  , w_19741 );
buf ( w_19739 , \6194_b1 );
not ( w_19739 , w_19742 );
not (  , w_19743 );
and ( w_19742 , w_19743 , \6194_b0 );
or ( \6196_b1 , \6133_b1 , w_19745 );
not ( w_19745 , w_19746 );
and ( \6196_b0 , \6133_b0 , w_19747 );
and ( w_19746 ,  , w_19747 );
buf ( w_19745 , \6195_b1 );
not ( w_19745 , w_19748 );
not (  , w_19749 );
and ( w_19748 , w_19749 , \6195_b0 );
or ( \6197_b1 , \6127_b1 , w_19751 );
not ( w_19751 , w_19752 );
and ( \6197_b0 , \6127_b0 , w_19753 );
and ( w_19752 ,  , w_19753 );
buf ( w_19751 , \6196_b1 );
not ( w_19751 , w_19754 );
not (  , w_19755 );
and ( w_19754 , w_19755 , \6196_b0 );
buf ( \6198_b1 , \6197_b1 );
not ( \6198_b1 , w_19756 );
not ( \6198_b0 , w_19757 );
and ( w_19756 , w_19757 , \6197_b0 );
or ( \6199_b1 , \6166_b1 , \6176_b1 );
xor ( \6199_b0 , \6166_b0 , w_19758 );
not ( w_19758 , w_19759 );
and ( w_19759 , \6176_b1 , \6176_b0 );
or ( \6200_b1 , \6199_b1 , \6180_b1 );
xor ( \6200_b0 , \6199_b0 , w_19760 );
not ( w_19760 , w_19761 );
and ( w_19761 , \6180_b1 , \6180_b0 );
buf ( \6201_b1 , \4128_b1 );
not ( \6201_b1 , w_19762 );
not ( \6201_b0 , w_19763 );
and ( w_19762 , w_19763 , \4128_b0 );
or ( \6202_b1 , \6201_b1 , w_19765 );
not ( w_19765 , w_19766 );
and ( \6202_b0 , \6201_b0 , w_19767 );
and ( w_19766 ,  , w_19767 );
buf ( w_19765 , \4048_b1 );
not ( w_19765 , w_19768 );
not (  , w_19769 );
and ( w_19768 , w_19769 , \4048_b0 );
buf ( \6203_b1 , \6202_b1 );
not ( \6203_b1 , w_19770 );
not ( \6203_b0 , w_19771 );
and ( w_19770 , w_19771 , \6202_b0 );
buf ( \6204_b1 , \4089_b1 );
not ( \6204_b1 , w_19772 );
not ( \6204_b0 , w_19773 );
and ( w_19772 , w_19773 , \4089_b0 );
or ( \6205_b1 , \6203_b1 , \6204_b1 );
not ( \6204_b1 , w_19774 );
and ( \6205_b0 , \6203_b0 , w_19775 );
and ( w_19774 , w_19775 , \6204_b0 );
buf ( \6206_b1 , \4048_b1 );
not ( \6206_b1 , w_19776 );
not ( \6206_b0 , w_19777 );
and ( w_19776 , w_19777 , \4048_b0 );
buf ( \6207_b1 , \6201_b1 );
not ( \6207_b1 , w_19778 );
not ( \6207_b0 , w_19779 );
and ( w_19778 , w_19779 , \6201_b0 );
or ( \6208_b1 , \6206_b1 , w_19780 );
or ( \6208_b0 , \6206_b0 , \6207_b0 );
not ( \6207_b0 , w_19781 );
and ( w_19781 , w_19780 , \6207_b1 );
or ( \6209_b1 , \6208_b1 , w_19783 );
not ( w_19783 , w_19784 );
and ( \6209_b0 , \6208_b0 , w_19785 );
and ( w_19784 ,  , w_19785 );
buf ( w_19783 , \4109_b1 );
not ( w_19783 , w_19786 );
not (  , w_19787 );
and ( w_19786 , w_19787 , \4109_b0 );
or ( \6210_b1 , \6205_b1 , w_19789 );
not ( w_19789 , w_19790 );
and ( \6210_b0 , \6205_b0 , w_19791 );
and ( w_19790 ,  , w_19791 );
buf ( w_19789 , \6209_b1 );
not ( w_19789 , w_19792 );
not (  , w_19793 );
and ( w_19792 , w_19793 , \6209_b0 );
or ( \6211_b1 , \4473_b1 , \5178_b1 );
not ( \5178_b1 , w_19794 );
and ( \6211_b0 , \4473_b0 , w_19795 );
and ( w_19794 , w_19795 , \5178_b0 );
buf ( \6212_b1 , \4473_b1 );
not ( \6212_b1 , w_19796 );
not ( \6212_b0 , w_19797 );
and ( w_19796 , w_19797 , \4473_b0 );
or ( \6213_b1 , \6212_b1 , \4665_b1 );
not ( \4665_b1 , w_19798 );
and ( \6213_b0 , \6212_b0 , w_19799 );
and ( w_19798 , w_19799 , \4665_b0 );
or ( \6214_b1 , \6211_b1 , w_19801 );
not ( w_19801 , w_19802 );
and ( \6214_b0 , \6211_b0 , w_19803 );
and ( w_19802 ,  , w_19803 );
buf ( w_19801 , \6213_b1 );
not ( w_19801 , w_19804 );
not (  , w_19805 );
and ( w_19804 , w_19805 , \6213_b0 );
or ( \6215_b1 , \4541_b1 , w_19807 );
not ( w_19807 , w_19808 );
and ( \6215_b0 , \4541_b0 , w_19809 );
and ( w_19808 ,  , w_19809 );
buf ( w_19807 , \6214_b1 );
not ( w_19807 , w_19810 );
not (  , w_19811 );
and ( w_19810 , w_19811 , \6214_b0 );
or ( \6216_b1 , \6215_b1 , w_19812 );
or ( \6216_b0 , \6215_b0 , \5187_b0 );
not ( \5187_b0 , w_19813 );
and ( w_19813 , w_19812 , \5187_b1 );
buf ( \6217_b1 , \4046_b1 );
not ( \6217_b1 , w_19814 );
not ( \6217_b0 , w_19815 );
and ( w_19814 , w_19815 , \4046_b0 );
buf ( \6218_b1 , \5178_b1 );
not ( \6218_b1 , w_19816 );
not ( \6218_b0 , w_19817 );
and ( w_19816 , w_19817 , \5178_b0 );
or ( \6219_b1 , \6217_b1 , w_19818 );
or ( \6219_b0 , \6217_b0 , \6218_b0 );
not ( \6218_b0 , w_19819 );
and ( w_19819 , w_19818 , \6218_b1 );
or ( \6220_b1 , \4665_b1 , w_19821 );
not ( w_19821 , w_19822 );
and ( \6220_b0 , \4665_b0 , w_19823 );
and ( w_19822 ,  , w_19823 );
buf ( w_19821 , \4256_b1 );
not ( w_19821 , w_19824 );
not (  , w_19825 );
and ( w_19824 , w_19825 , \4256_b0 );
or ( \6221_b1 , \6219_b1 , w_19827 );
not ( w_19827 , w_19828 );
and ( \6221_b0 , \6219_b0 , w_19829 );
and ( w_19828 ,  , w_19829 );
buf ( w_19827 , \6220_b1 );
not ( w_19827 , w_19830 );
not (  , w_19831 );
and ( w_19830 , w_19831 , \6220_b0 );
or ( \6222_b1 , \5187_b1 , w_19833 );
not ( w_19833 , w_19834 );
and ( \6222_b0 , \5187_b0 , w_19835 );
and ( w_19834 ,  , w_19835 );
buf ( w_19833 , \6221_b1 );
not ( w_19833 , w_19836 );
not (  , w_19837 );
and ( w_19836 , w_19837 , \6221_b0 );
or ( \6223_b1 , \6216_b1 , w_19839 );
not ( w_19839 , w_19840 );
and ( \6223_b0 , \6216_b0 , w_19841 );
and ( w_19840 ,  , w_19841 );
buf ( w_19839 , \6222_b1 );
not ( w_19839 , w_19842 );
not (  , w_19843 );
and ( w_19842 , w_19843 , \6222_b0 );
or ( \6224_b1 , \6210_b1 , \6223_b1 );
not ( \6223_b1 , w_19844 );
and ( \6224_b0 , \6210_b0 , w_19845 );
and ( w_19844 , w_19845 , \6223_b0 );
buf ( \6225_b1 , \5390_b1 );
not ( \6225_b1 , w_19846 );
not ( \6225_b0 , w_19847 );
and ( w_19846 , w_19847 , \5390_b0 );
buf ( \6226_b1 , \4011_b1 );
not ( \6226_b1 , w_19848 );
not ( \6226_b0 , w_19849 );
and ( w_19848 , w_19849 , \4011_b0 );
buf ( \6227_b1 , \5273_b1 );
not ( \6227_b1 , w_19850 );
not ( \6227_b0 , w_19851 );
and ( w_19850 , w_19851 , \5273_b0 );
buf ( \6228_b1 , \6227_b1 );
not ( \6228_b1 , w_19852 );
not ( \6228_b0 , w_19853 );
and ( w_19852 , w_19853 , \6227_b0 );
or ( \6229_b1 , \6226_b1 , w_19854 );
or ( \6229_b0 , \6226_b0 , \6228_b0 );
not ( \6228_b0 , w_19855 );
and ( w_19855 , w_19854 , \6228_b1 );
or ( \6230_b1 , \5873_b1 , w_19857 );
not ( w_19857 , w_19858 );
and ( \6230_b0 , \5873_b0 , w_19859 );
and ( w_19858 ,  , w_19859 );
buf ( w_19857 , \4270_b1 );
not ( w_19857 , w_19860 );
not (  , w_19861 );
and ( w_19860 , w_19861 , \4270_b0 );
or ( \6231_b1 , \6229_b1 , w_19863 );
not ( w_19863 , w_19864 );
and ( \6231_b0 , \6229_b0 , w_19865 );
and ( w_19864 ,  , w_19865 );
buf ( w_19863 , \6230_b1 );
not ( w_19863 , w_19866 );
not (  , w_19867 );
and ( w_19866 , w_19867 , \6230_b0 );
buf ( \6232_b1 , \6231_b1 );
not ( \6232_b1 , w_19868 );
not ( \6232_b0 , w_19869 );
and ( w_19868 , w_19869 , \6231_b0 );
or ( \6233_b1 , \6225_b1 , w_19870 );
or ( \6233_b0 , \6225_b0 , \6232_b0 );
not ( \6232_b0 , w_19871 );
and ( w_19871 , w_19870 , \6232_b1 );
buf ( \6234_b1 , \4043_b1 );
not ( \6234_b1 , w_19872 );
not ( \6234_b0 , w_19873 );
and ( w_19872 , w_19873 , \4043_b0 );
buf ( \6235_b1 , \5576_b1 );
not ( \6235_b1 , w_19874 );
not ( \6235_b0 , w_19875 );
and ( w_19874 , w_19875 , \5576_b0 );
or ( \6236_b1 , \6234_b1 , w_19876 );
or ( \6236_b0 , \6234_b0 , \6235_b0 );
not ( \6235_b0 , w_19877 );
and ( w_19877 , w_19876 , \6235_b1 );
or ( \6237_b1 , \4217_b1 , w_19879 );
not ( w_19879 , w_19880 );
and ( \6237_b0 , \4217_b0 , w_19881 );
and ( w_19880 ,  , w_19881 );
buf ( w_19879 , \5873_b1 );
not ( w_19879 , w_19882 );
not (  , w_19883 );
and ( w_19882 , w_19883 , \5873_b0 );
or ( \6238_b1 , \6236_b1 , w_19885 );
not ( w_19885 , w_19886 );
and ( \6238_b0 , \6236_b0 , w_19887 );
and ( w_19886 ,  , w_19887 );
buf ( w_19885 , \6237_b1 );
not ( w_19885 , w_19888 );
not (  , w_19889 );
and ( w_19888 , w_19889 , \6237_b0 );
or ( \6239_b1 , \6238_b1 , w_19891 );
not ( w_19891 , w_19892 );
and ( \6239_b0 , \6238_b0 , w_19893 );
and ( w_19892 ,  , w_19893 );
buf ( w_19891 , \5021_b1 );
not ( w_19891 , w_19894 );
not (  , w_19895 );
and ( w_19894 , w_19895 , \5021_b0 );
or ( \6240_b1 , \6233_b1 , w_19897 );
not ( w_19897 , w_19898 );
and ( \6240_b0 , \6233_b0 , w_19899 );
and ( w_19898 ,  , w_19899 );
buf ( w_19897 , \6239_b1 );
not ( w_19897 , w_19900 );
not (  , w_19901 );
and ( w_19900 , w_19901 , \6239_b0 );
or ( \6241_b1 , \4114_b1 , \4029_b1 );
not ( \4029_b1 , w_19902 );
and ( \6241_b0 , \4114_b0 , w_19903 );
and ( w_19902 , w_19903 , \4029_b0 );
or ( \6242_b1 , \4109_b1 , \5339_b1 );
not ( \5339_b1 , w_19904 );
and ( \6242_b0 , \4109_b0 , w_19905 );
and ( w_19904 , w_19905 , \5339_b0 );
or ( \6243_b1 , \6241_b1 , w_19907 );
not ( w_19907 , w_19908 );
and ( \6243_b0 , \6241_b0 , w_19909 );
and ( w_19908 ,  , w_19909 );
buf ( w_19907 , \6242_b1 );
not ( w_19907 , w_19910 );
not (  , w_19911 );
and ( w_19910 , w_19911 , \6242_b0 );
buf ( \6244_b1 , \4139_b1 );
not ( \6244_b1 , w_19912 );
not ( \6244_b0 , w_19913 );
and ( w_19912 , w_19913 , \4139_b0 );
or ( \6245_b1 , \6243_b1 , w_19914 );
or ( \6245_b0 , \6243_b0 , \6244_b0 );
not ( \6244_b0 , w_19915 );
and ( w_19915 , w_19914 , \6244_b1 );
buf ( \6246_b1 , \4139_b1 );
not ( \6246_b1 , w_19916 );
not ( \6246_b0 , w_19917 );
and ( w_19916 , w_19917 , \4139_b0 );
or ( \6247_b1 , \4048_b1 , \4146_b1 );
not ( \4146_b1 , w_19918 );
and ( \6247_b0 , \4048_b0 , w_19919 );
and ( w_19918 , w_19919 , \4146_b0 );
buf ( \6248_b1 , \4048_b1 );
not ( \6248_b1 , w_19920 );
not ( \6248_b0 , w_19921 );
and ( w_19920 , w_19921 , \4048_b0 );
or ( \6249_b1 , \6248_b1 , \4145_b1 );
not ( \4145_b1 , w_19922 );
and ( \6249_b0 , \6248_b0 , w_19923 );
and ( w_19922 , w_19923 , \4145_b0 );
or ( \6250_b1 , \6247_b1 , w_19925 );
not ( w_19925 , w_19926 );
and ( \6250_b0 , \6247_b0 , w_19927 );
and ( w_19926 ,  , w_19927 );
buf ( w_19925 , \6249_b1 );
not ( w_19925 , w_19928 );
not (  , w_19929 );
and ( w_19928 , w_19929 , \6249_b0 );
or ( \6252_b1 , \6245_b1 , w_19931 );
not ( w_19931 , w_19932 );
and ( \6252_b0 , \6245_b0 , w_19933 );
and ( w_19932 ,  , w_19933 );
buf ( w_19931 , \6251_b1 );
not ( w_19931 , w_19934 );
not (  , w_19935 );
and ( w_19934 , w_19935 , \6251_b0 );
or ( \6253_b1 , \6240_b1 , \6252_b1 );
xor ( \6253_b0 , \6240_b0 , w_19936 );
not ( w_19936 , w_19937 );
and ( w_19937 , \6252_b1 , \6252_b0 );
buf ( \6254_b1 , \4026_b1 );
not ( \6254_b1 , w_19938 );
not ( \6254_b0 , w_19939 );
and ( w_19938 , w_19939 , \4026_b0 );
buf ( \6255_b1 , \4089_b1 );
not ( \6255_b1 , w_19940 );
not ( \6255_b0 , w_19941 );
and ( w_19940 , w_19941 , \4089_b0 );
or ( \6256_b1 , \6254_b1 , w_19942 );
or ( \6256_b0 , \6254_b0 , \6255_b0 );
not ( \6255_b0 , w_19943 );
and ( w_19943 , w_19942 , \6255_b1 );
or ( \6257_b1 , \4088_b1 , w_19945 );
not ( w_19945 , w_19946 );
and ( \6257_b0 , \4088_b0 , w_19947 );
and ( w_19946 ,  , w_19947 );
buf ( w_19945 , \5344_b1 );
not ( w_19945 , w_19948 );
not (  , w_19949 );
and ( w_19948 , w_19949 , \5344_b0 );
or ( \6258_b1 , \6256_b1 , w_19951 );
not ( w_19951 , w_19952 );
and ( \6258_b0 , \6256_b0 , w_19953 );
and ( w_19952 ,  , w_19953 );
buf ( w_19951 , \6257_b1 );
not ( w_19951 , w_19954 );
not (  , w_19955 );
and ( w_19954 , w_19955 , \6257_b0 );
buf ( \6259_b1 , \6258_b1 );
not ( \6259_b1 , w_19956 );
not ( \6259_b0 , w_19957 );
and ( w_19956 , w_19957 , \6258_b0 );
buf ( \6260_b1 , \4437_b1 );
not ( \6260_b1 , w_19958 );
not ( \6260_b0 , w_19959 );
and ( w_19958 , w_19959 , \4437_b0 );
or ( \6261_b1 , \6259_b1 , w_19960 );
or ( \6261_b0 , \6259_b0 , \6260_b0 );
not ( \6260_b0 , w_19961 );
and ( w_19961 , w_19960 , \6260_b1 );
buf ( \6262_b1 , \4023_b1 );
not ( \6262_b1 , w_19962 );
not ( \6262_b0 , w_19963 );
and ( w_19962 , w_19963 , \4023_b0 );
buf ( \6263_b1 , \5234_b1 );
not ( \6263_b1 , w_19964 );
not ( \6263_b0 , w_19965 );
and ( w_19964 , w_19965 , \5234_b0 );
or ( \6264_b1 , \6262_b1 , w_19966 );
or ( \6264_b0 , \6262_b0 , \6263_b0 );
not ( \6263_b0 , w_19967 );
and ( w_19967 , w_19966 , \6263_b1 );
or ( \6265_b1 , \4088_b1 , w_19969 );
not ( w_19969 , w_19970 );
and ( \6265_b0 , \4088_b0 , w_19971 );
and ( w_19970 ,  , w_19971 );
buf ( w_19969 , \5131_b1 );
not ( w_19969 , w_19972 );
not (  , w_19973 );
and ( w_19972 , w_19973 , \5131_b0 );
or ( \6266_b1 , \6264_b1 , w_19975 );
not ( w_19975 , w_19976 );
and ( \6266_b0 , \6264_b0 , w_19977 );
and ( w_19976 ,  , w_19977 );
buf ( w_19975 , \6265_b1 );
not ( w_19975 , w_19978 );
not (  , w_19979 );
and ( w_19978 , w_19979 , \6265_b0 );
or ( \6267_b1 , \4331_b1 , w_19981 );
not ( w_19981 , w_19982 );
and ( \6267_b0 , \4331_b0 , w_19983 );
and ( w_19982 ,  , w_19983 );
buf ( w_19981 , \6266_b1 );
not ( w_19981 , w_19984 );
not (  , w_19985 );
and ( w_19984 , w_19985 , \6266_b0 );
or ( \6268_b1 , \6261_b1 , w_19987 );
not ( w_19987 , w_19988 );
and ( \6268_b0 , \6261_b0 , w_19989 );
and ( w_19988 ,  , w_19989 );
buf ( w_19987 , \6267_b1 );
not ( w_19987 , w_19990 );
not (  , w_19991 );
and ( w_19990 , w_19991 , \6267_b0 );
or ( \6269_b1 , \6253_b1 , \6268_b1 );
not ( \6268_b1 , w_19992 );
and ( \6269_b0 , \6253_b0 , w_19993 );
and ( w_19992 , w_19993 , \6268_b0 );
or ( \6270_b1 , \6240_b1 , \6252_b1 );
not ( \6252_b1 , w_19994 );
and ( \6270_b0 , \6240_b0 , w_19995 );
and ( w_19994 , w_19995 , \6252_b0 );
or ( \6271_b1 , \6269_b1 , w_19996 );
or ( \6271_b0 , \6269_b0 , \6270_b0 );
not ( \6270_b0 , w_19997 );
and ( w_19997 , w_19996 , \6270_b1 );
or ( \6272_b1 , \6224_b1 , \6271_b1 );
xor ( \6272_b0 , \6224_b0 , w_19998 );
not ( w_19998 , w_19999 );
and ( w_19999 , \6271_b1 , \6271_b0 );
or ( \6273_b1 , \5816_b1 , \4048_b1 );
not ( \4048_b1 , w_20000 );
and ( \6273_b0 , \5816_b0 , w_20001 );
and ( w_20000 , w_20001 , \4048_b0 );
buf ( \6274_b1 , \6266_b1 );
not ( \6274_b1 , w_20002 );
not ( \6274_b0 , w_20003 );
and ( w_20002 , w_20003 , \6266_b0 );
buf ( \6275_b1 , \4437_b1 );
not ( \6275_b1 , w_20004 );
not ( \6275_b0 , w_20005 );
and ( w_20004 , w_20005 , \4437_b0 );
or ( \6276_b1 , \6274_b1 , w_20006 );
or ( \6276_b0 , \6274_b0 , \6275_b0 );
not ( \6275_b0 , w_20007 );
and ( w_20007 , w_20006 , \6275_b1 );
or ( \6277_b1 , \4331_b1 , w_20009 );
not ( w_20009 , w_20010 );
and ( \6277_b0 , \4331_b0 , w_20011 );
and ( w_20010 ,  , w_20011 );
buf ( w_20009 , \6107_b1 );
not ( w_20009 , w_20012 );
not (  , w_20013 );
and ( w_20012 , w_20013 , \6107_b0 );
or ( \6278_b1 , \6276_b1 , w_20015 );
not ( w_20015 , w_20016 );
and ( \6278_b0 , \6276_b0 , w_20017 );
and ( w_20016 ,  , w_20017 );
buf ( w_20015 , \6277_b1 );
not ( w_20015 , w_20018 );
not (  , w_20019 );
and ( w_20018 , w_20019 , \6277_b0 );
or ( \6279_b1 , \6273_b1 , \6278_b1 );
xor ( \6279_b0 , \6273_b0 , w_20020 );
not ( w_20020 , w_20021 );
and ( w_20021 , \6278_b1 , \6278_b0 );
buf ( \6280_b1 , \6221_b1 );
not ( \6280_b1 , w_20022 );
not ( \6280_b0 , w_20023 );
and ( w_20022 , w_20023 , \6221_b0 );
buf ( \6281_b1 , \4662_b1 );
not ( \6281_b1 , w_20024 );
not ( \6281_b0 , w_20025 );
and ( w_20024 , w_20025 , \4662_b0 );
or ( \6282_b1 , \6280_b1 , w_20026 );
or ( \6282_b0 , \6280_b0 , \6281_b0 );
not ( \6281_b0 , w_20027 );
and ( w_20027 , w_20026 , \6281_b1 );
or ( \6283_b1 , \4672_b1 , w_20029 );
not ( w_20029 , w_20030 );
and ( \6283_b0 , \4672_b0 , w_20031 );
and ( w_20030 ,  , w_20031 );
buf ( w_20029 , \6076_b1 );
not ( w_20029 , w_20032 );
not (  , w_20033 );
and ( w_20032 , w_20033 , \6076_b0 );
or ( \6284_b1 , \6282_b1 , w_20035 );
not ( w_20035 , w_20036 );
and ( \6284_b0 , \6282_b0 , w_20037 );
and ( w_20036 ,  , w_20037 );
buf ( w_20035 , \6283_b1 );
not ( w_20035 , w_20038 );
not (  , w_20039 );
and ( w_20038 , w_20039 , \6283_b0 );
or ( \6285_b1 , \6279_b1 , \6284_b1 );
xor ( \6285_b0 , \6279_b0 , w_20040 );
not ( w_20040 , w_20041 );
and ( w_20041 , \6284_b1 , \6284_b0 );
or ( \6286_b1 , \6272_b1 , \6285_b1 );
not ( \6285_b1 , w_20042 );
and ( \6286_b0 , \6272_b0 , w_20043 );
and ( w_20042 , w_20043 , \6285_b0 );
or ( \6287_b1 , \6224_b1 , \6271_b1 );
not ( \6271_b1 , w_20044 );
and ( \6287_b0 , \6224_b0 , w_20045 );
and ( w_20044 , w_20045 , \6271_b0 );
or ( \6288_b1 , \6286_b1 , w_20046 );
or ( \6288_b0 , \6286_b0 , \6287_b0 );
not ( \6287_b0 , w_20047 );
and ( w_20047 , w_20046 , \6287_b1 );
or ( \6289_b1 , \6200_b1 , \6288_b1 );
xor ( \6289_b0 , \6200_b0 , w_20048 );
not ( w_20048 , w_20049 );
and ( w_20049 , \6288_b1 , \6288_b0 );
buf ( \6290_b1 , \6087_b1 );
not ( \6290_b1 , w_20050 );
not ( \6290_b0 , w_20051 );
and ( w_20050 , w_20051 , \6087_b0 );
buf ( \6291_b1 , \5265_b1 );
not ( \6291_b1 , w_20052 );
not ( \6291_b0 , w_20053 );
and ( w_20052 , w_20053 , \5265_b0 );
or ( \6292_b1 , \6290_b1 , \6291_b1 );
not ( \6291_b1 , w_20054 );
and ( \6292_b0 , \6290_b0 , w_20055 );
and ( w_20054 , w_20055 , \6291_b0 );
or ( \6293_b1 , \5019_b1 , \6238_b1 );
not ( \6238_b1 , w_20056 );
and ( \6293_b0 , \5019_b0 , w_20057 );
and ( w_20056 , w_20057 , \6238_b0 );
or ( \6294_b1 , \6292_b1 , w_20059 );
not ( w_20059 , w_20060 );
and ( \6294_b0 , \6292_b0 , w_20061 );
and ( w_20060 ,  , w_20061 );
buf ( w_20059 , \6293_b1 );
not ( w_20059 , w_20062 );
not (  , w_20063 );
and ( w_20062 , w_20063 , \6293_b0 );
buf ( \6295_b1 , \6294_b1 );
not ( \6295_b1 , w_20064 );
not ( \6295_b0 , w_20065 );
and ( w_20064 , w_20065 , \6294_b0 );
buf ( \6296_b1 , \6295_b1 );
not ( \6296_b1 , w_20066 );
not ( \6296_b0 , w_20067 );
and ( w_20066 , w_20067 , \6295_b0 );
buf ( \6297_b1 , \6244_b1 );
not ( \6297_b1 , w_20068 );
not ( \6297_b0 , w_20069 );
and ( w_20068 , w_20069 , \6244_b0 );
buf ( \6298_b1 , \4134_b1 );
not ( \6298_b1 , w_20070 );
not ( \6298_b0 , w_20071 );
and ( w_20070 , w_20071 , \4134_b0 );
or ( \6299_b1 , \6298_b1 , w_20073 );
not ( w_20073 , w_20074 );
and ( \6299_b0 , \6298_b0 , w_20075 );
and ( w_20074 ,  , w_20075 );
buf ( w_20073 , \6243_b1 );
not ( w_20073 , w_20076 );
not (  , w_20077 );
and ( w_20076 , w_20077 , \6243_b0 );
buf ( \6300_b1 , \6299_b1 );
not ( \6300_b1 , w_20078 );
not ( \6300_b0 , w_20079 );
and ( w_20078 , w_20079 , \6299_b0 );
or ( \6301_b1 , \6297_b1 , w_20080 );
or ( \6301_b0 , \6297_b0 , \6300_b0 );
not ( \6300_b0 , w_20081 );
and ( w_20081 , w_20080 , \6300_b1 );
or ( \6302_b1 , \4139_b1 , w_20083 );
not ( w_20083 , w_20084 );
and ( \6302_b0 , \4139_b0 , w_20085 );
and ( w_20084 ,  , w_20085 );
buf ( w_20083 , \6097_b1 );
not ( w_20083 , w_20086 );
not (  , w_20087 );
and ( w_20086 , w_20087 , \6097_b0 );
or ( \6303_b1 , \6301_b1 , w_20089 );
not ( w_20089 , w_20090 );
and ( \6303_b0 , \6301_b0 , w_20091 );
and ( w_20090 ,  , w_20091 );
buf ( w_20089 , \6302_b1 );
not ( w_20089 , w_20092 );
not (  , w_20093 );
and ( w_20092 , w_20093 , \6302_b0 );
buf ( \6304_b1 , \6303_b1 );
not ( \6304_b1 , w_20094 );
not ( \6304_b0 , w_20095 );
and ( w_20094 , w_20095 , \6303_b0 );
or ( \6305_b1 , \6296_b1 , w_20096 );
or ( \6305_b0 , \6296_b0 , \6304_b0 );
not ( \6304_b0 , w_20097 );
and ( w_20097 , w_20096 , \6304_b1 );
or ( \6306_b1 , \6303_b1 , w_20098 );
or ( \6306_b0 , \6303_b0 , \6295_b0 );
not ( \6295_b0 , w_20099 );
and ( w_20099 , w_20098 , \6295_b1 );
buf ( \6307_b1 , \3963_b1 );
not ( \6307_b1 , w_20100 );
not ( \6307_b0 , w_20101 );
and ( w_20100 , w_20101 , \3963_b0 );
buf ( \6308_b1 , \5904_b1 );
not ( \6308_b1 , w_20102 );
not ( \6308_b0 , w_20103 );
and ( w_20102 , w_20103 , \5904_b0 );
or ( \6309_b1 , \6307_b1 , w_20104 );
or ( \6309_b0 , \6307_b0 , \6308_b0 );
not ( \6308_b0 , w_20105 );
and ( w_20105 , w_20104 , \6308_b1 );
or ( \6310_b1 , \4403_b1 , w_20107 );
not ( w_20107 , w_20108 );
and ( \6310_b0 , \4403_b0 , w_20109 );
and ( w_20108 ,  , w_20109 );
buf ( w_20107 , \4486_b1 );
not ( w_20107 , w_20110 );
not (  , w_20111 );
and ( w_20110 , w_20111 , \4486_b0 );
or ( \6311_b1 , \6309_b1 , w_20113 );
not ( w_20113 , w_20114 );
and ( \6311_b0 , \6309_b0 , w_20115 );
and ( w_20114 ,  , w_20115 );
buf ( w_20113 , \6310_b1 );
not ( w_20113 , w_20116 );
not (  , w_20117 );
and ( w_20116 , w_20117 , \6310_b0 );
buf ( \6312_b1 , \6311_b1 );
not ( \6312_b1 , w_20118 );
not ( \6312_b0 , w_20119 );
and ( w_20118 , w_20119 , \6311_b0 );
buf ( \6313_b1 , \6162_b1 );
not ( \6313_b1 , w_20120 );
not ( \6313_b0 , w_20121 );
and ( w_20120 , w_20121 , \6162_b0 );
or ( \6314_b1 , \6312_b1 , w_20122 );
or ( \6314_b0 , \6312_b0 , \6313_b0 );
not ( \6313_b0 , w_20123 );
and ( w_20123 , w_20122 , \6313_b1 );
or ( \6315_b1 , \4055_b1 , w_20125 );
not ( w_20125 , w_20126 );
and ( \6315_b0 , \4055_b0 , w_20127 );
and ( w_20126 ,  , w_20127 );
buf ( w_20125 , \6160_b1 );
not ( w_20125 , w_20128 );
not (  , w_20129 );
and ( w_20128 , w_20129 , \6160_b0 );
or ( \6316_b1 , \6314_b1 , w_20131 );
not ( w_20131 , w_20132 );
and ( \6316_b0 , \6314_b0 , w_20133 );
and ( w_20132 ,  , w_20133 );
buf ( w_20131 , \6315_b1 );
not ( w_20131 , w_20134 );
not (  , w_20135 );
and ( w_20134 , w_20135 , \6315_b0 );
or ( \6317_b1 , \6306_b1 , w_20137 );
not ( w_20137 , w_20138 );
and ( \6317_b0 , \6306_b0 , w_20139 );
and ( w_20138 ,  , w_20139 );
buf ( w_20137 , \6316_b1 );
not ( w_20137 , w_20140 );
not (  , w_20141 );
and ( w_20140 , w_20141 , \6316_b0 );
or ( \6318_b1 , \6305_b1 , w_20143 );
not ( w_20143 , w_20144 );
and ( \6318_b0 , \6305_b0 , w_20145 );
and ( w_20144 ,  , w_20145 );
buf ( w_20143 , \6317_b1 );
not ( w_20143 , w_20146 );
not (  , w_20147 );
and ( w_20146 , w_20147 , \6317_b0 );
or ( \6319_b1 , \6273_b1 , \6278_b1 );
xor ( \6319_b0 , \6273_b0 , w_20148 );
not ( w_20148 , w_20149 );
and ( w_20149 , \6278_b1 , \6278_b0 );
or ( \6320_b1 , \6319_b1 , \6284_b1 );
not ( \6284_b1 , w_20150 );
and ( \6320_b0 , \6319_b0 , w_20151 );
and ( w_20150 , w_20151 , \6284_b0 );
or ( \6321_b1 , \6273_b1 , \6278_b1 );
not ( \6278_b1 , w_20152 );
and ( \6321_b0 , \6273_b0 , w_20153 );
and ( w_20152 , w_20153 , \6278_b0 );
or ( \6322_b1 , \6320_b1 , w_20154 );
or ( \6322_b0 , \6320_b0 , \6321_b0 );
not ( \6321_b0 , w_20155 );
and ( w_20155 , w_20154 , \6321_b1 );
or ( \6323_b1 , \6318_b1 , \6322_b1 );
xor ( \6323_b0 , \6318_b0 , w_20156 );
not ( w_20156 , w_20157 );
and ( w_20157 , \6322_b1 , \6322_b0 );
or ( \6324_b1 , \6093_b1 , \6102_b1 );
xor ( \6324_b0 , \6093_b0 , w_20158 );
not ( w_20158 , w_20159 );
and ( w_20159 , \6102_b1 , \6102_b0 );
or ( \6325_b1 , \6324_b1 , \6112_b1 );
xor ( \6325_b0 , \6324_b0 , w_20160 );
not ( w_20160 , w_20161 );
and ( w_20161 , \6112_b1 , \6112_b0 );
or ( \6326_b1 , \6323_b1 , \6325_b1 );
xor ( \6326_b0 , \6323_b0 , w_20162 );
not ( w_20162 , w_20163 );
and ( w_20163 , \6325_b1 , \6325_b0 );
or ( \6327_b1 , \6289_b1 , w_20164 );
xor ( \6327_b0 , \6289_b0 , w_20166 );
not ( w_20166 , w_20167 );
and ( w_20167 , w_20164 , w_20165 );
buf ( w_20164 , \6326_b1 );
not ( w_20164 , w_20168 );
not ( w_20165 , w_20169 );
and ( w_20168 , w_20169 , \6326_b0 );
or ( \6328_b1 , \6224_b1 , \6271_b1 );
xor ( \6328_b0 , \6224_b0 , w_20170 );
not ( w_20170 , w_20171 );
and ( w_20171 , \6271_b1 , \6271_b0 );
or ( \6329_b1 , \6328_b1 , \6285_b1 );
xor ( \6329_b0 , \6328_b0 , w_20172 );
not ( w_20172 , w_20173 );
and ( w_20173 , \6285_b1 , \6285_b0 );
buf ( \6330_b1 , \6329_b1 );
not ( \6330_b1 , w_20174 );
not ( \6330_b0 , w_20175 );
and ( w_20174 , w_20175 , \6329_b0 );
buf ( \6331_b1 , \6330_b1 );
not ( \6331_b1 , w_20176 );
not ( \6331_b0 , w_20177 );
and ( w_20176 , w_20177 , \6330_b0 );
buf ( \6332_b1 , \4019_b1 );
not ( \6332_b1 , w_20178 );
not ( \6332_b0 , w_20179 );
and ( w_20178 , w_20179 , \4019_b0 );
buf ( \6333_b1 , \4069_b1 );
not ( \6333_b1 , w_20180 );
not ( \6333_b0 , w_20181 );
and ( w_20180 , w_20181 , \4069_b0 );
or ( \6334_b1 , \6332_b1 , w_20182 );
or ( \6334_b0 , \6332_b0 , \6333_b0 );
not ( \6333_b0 , w_20183 );
and ( w_20183 , w_20182 , \6333_b1 );
or ( \6335_b1 , \4403_b1 , w_20185 );
not ( w_20185 , w_20186 );
and ( \6335_b0 , \4403_b0 , w_20187 );
and ( w_20186 ,  , w_20187 );
buf ( w_20185 , \4585_b1 );
not ( w_20185 , w_20188 );
not (  , w_20189 );
and ( w_20188 , w_20189 , \4585_b0 );
or ( \6336_b1 , \6334_b1 , w_20191 );
not ( w_20191 , w_20192 );
and ( \6336_b0 , \6334_b0 , w_20193 );
and ( w_20192 ,  , w_20193 );
buf ( w_20191 , \6335_b1 );
not ( w_20191 , w_20194 );
not (  , w_20195 );
and ( w_20194 , w_20195 , \6335_b0 );
buf ( \6337_b1 , \6336_b1 );
not ( \6337_b1 , w_20196 );
not ( \6337_b0 , w_20197 );
and ( w_20196 , w_20197 , \6336_b0 );
buf ( \6338_b1 , \5361_b1 );
not ( \6338_b1 , w_20198 );
not ( \6338_b0 , w_20199 );
and ( w_20198 , w_20199 , \5361_b0 );
or ( \6339_b1 , \6337_b1 , w_20200 );
or ( \6339_b0 , \6337_b0 , \6338_b0 );
not ( \6338_b0 , w_20201 );
and ( w_20201 , w_20200 , \6338_b1 );
or ( \6340_b1 , \4055_b1 , w_20203 );
not ( w_20203 , w_20204 );
and ( \6340_b0 , \4055_b0 , w_20205 );
and ( w_20204 ,  , w_20205 );
buf ( w_20203 , \6311_b1 );
not ( w_20203 , w_20206 );
not (  , w_20207 );
and ( w_20206 , w_20207 , \6311_b0 );
or ( \6341_b1 , \6339_b1 , w_20209 );
not ( w_20209 , w_20210 );
and ( \6341_b0 , \6339_b0 , w_20211 );
and ( w_20210 ,  , w_20211 );
buf ( w_20209 , \6340_b1 );
not ( w_20209 , w_20212 );
not (  , w_20213 );
and ( w_20212 , w_20213 , \6340_b0 );
or ( \6342_b1 , \6210_b1 , \6223_b1 );
xor ( \6342_b0 , \6210_b0 , w_20214 );
not ( w_20214 , w_20215 );
and ( w_20215 , \6223_b1 , \6223_b0 );
or ( \6343_b1 , \6341_b1 , \6342_b1 );
xor ( \6343_b0 , \6341_b0 , w_20216 );
not ( w_20216 , w_20217 );
and ( w_20217 , \6342_b1 , \6342_b0 );
buf ( \6344_b1 , \6246_b1 );
not ( \6344_b1 , w_20218 );
not ( \6344_b0 , w_20219 );
and ( w_20218 , w_20219 , \6246_b0 );
or ( \6345_b1 , \6344_b1 , w_20221 );
not ( w_20221 , w_20222 );
and ( \6345_b0 , \6344_b0 , w_20223 );
and ( w_20222 ,  , w_20223 );
buf ( w_20221 , \4048_b1 );
not ( w_20221 , w_20224 );
not (  , w_20225 );
and ( w_20224 , w_20225 , \4048_b0 );
buf ( \6346_b1 , \5390_b1 );
not ( \6346_b1 , w_20226 );
not ( \6346_b0 , w_20227 );
and ( w_20226 , w_20227 , \5390_b0 );
buf ( \6347_b1 , \4046_b1 );
not ( \6347_b1 , w_20228 );
not ( \6347_b0 , w_20229 );
and ( w_20228 , w_20229 , \4046_b0 );
buf ( \6348_b1 , \6227_b1 );
not ( \6348_b1 , w_20230 );
not ( \6348_b0 , w_20231 );
and ( w_20230 , w_20231 , \6227_b0 );
or ( \6349_b1 , \6347_b1 , w_20232 );
or ( \6349_b0 , \6347_b0 , \6348_b0 );
not ( \6348_b0 , w_20233 );
and ( w_20233 , w_20232 , \6348_b1 );
buf ( \6350_b1 , \5270_b1 );
not ( \6350_b1 , w_20234 );
not ( \6350_b0 , w_20235 );
and ( w_20234 , w_20235 , \5270_b0 );
or ( \6351_b1 , \6350_b1 , w_20237 );
not ( w_20237 , w_20238 );
and ( \6351_b0 , \6350_b0 , w_20239 );
and ( w_20238 ,  , w_20239 );
buf ( w_20237 , \4256_b1 );
not ( w_20237 , w_20240 );
not (  , w_20241 );
and ( w_20240 , w_20241 , \4256_b0 );
or ( \6352_b1 , \6349_b1 , w_20243 );
not ( w_20243 , w_20244 );
and ( \6352_b0 , \6349_b0 , w_20245 );
and ( w_20244 ,  , w_20245 );
buf ( w_20243 , \6351_b1 );
not ( w_20243 , w_20246 );
not (  , w_20247 );
and ( w_20246 , w_20247 , \6351_b0 );
buf ( \6353_b1 , \6352_b1 );
not ( \6353_b1 , w_20248 );
not ( \6353_b0 , w_20249 );
and ( w_20248 , w_20249 , \6352_b0 );
or ( \6354_b1 , \6346_b1 , w_20250 );
or ( \6354_b0 , \6346_b0 , \6353_b0 );
not ( \6353_b0 , w_20251 );
and ( w_20251 , w_20250 , \6353_b1 );
or ( \6355_b1 , \6231_b1 , w_20253 );
not ( w_20253 , w_20254 );
and ( \6355_b0 , \6231_b0 , w_20255 );
and ( w_20254 ,  , w_20255 );
buf ( w_20253 , \5021_b1 );
not ( w_20253 , w_20256 );
not (  , w_20257 );
and ( w_20256 , w_20257 , \5021_b0 );
or ( \6356_b1 , \6354_b1 , w_20259 );
not ( w_20259 , w_20260 );
and ( \6356_b0 , \6354_b0 , w_20261 );
and ( w_20260 ,  , w_20261 );
buf ( w_20259 , \6355_b1 );
not ( w_20259 , w_20262 );
not (  , w_20263 );
and ( w_20262 , w_20263 , \6355_b0 );
buf ( \6357_b1 , \6356_b1 );
not ( \6357_b1 , w_20264 );
not ( \6357_b0 , w_20265 );
and ( w_20264 , w_20265 , \6356_b0 );
or ( \6358_b1 , \6345_b1 , w_20267 );
not ( w_20267 , w_20268 );
and ( \6358_b0 , \6345_b0 , w_20269 );
and ( w_20268 ,  , w_20269 );
buf ( w_20267 , \6357_b1 );
not ( w_20267 , w_20270 );
not (  , w_20271 );
and ( w_20270 , w_20271 , \6357_b0 );
buf ( \6359_b1 , \6358_b1 );
not ( \6359_b1 , w_20272 );
not ( \6359_b0 , w_20273 );
and ( w_20272 , w_20273 , \6358_b0 );
buf ( \6360_b1 , \4029_b1 );
not ( \6360_b1 , w_20274 );
not ( \6360_b0 , w_20275 );
and ( w_20274 , w_20275 , \4029_b0 );
buf ( \6361_b1 , \5234_b1 );
not ( \6361_b1 , w_20276 );
not ( \6361_b0 , w_20277 );
and ( w_20276 , w_20277 , \5234_b0 );
or ( \6362_b1 , \6360_b1 , w_20278 );
or ( \6362_b0 , \6360_b0 , \6361_b0 );
not ( \6361_b0 , w_20279 );
and ( w_20279 , w_20278 , \6361_b1 );
or ( \6363_b1 , \4088_b1 , w_20281 );
not ( w_20281 , w_20282 );
and ( \6363_b0 , \4088_b0 , w_20283 );
and ( w_20282 ,  , w_20283 );
buf ( w_20281 , \5339_b1 );
not ( w_20281 , w_20284 );
not (  , w_20285 );
and ( w_20284 , w_20285 , \5339_b0 );
or ( \6364_b1 , \6362_b1 , w_20287 );
not ( w_20287 , w_20288 );
and ( \6364_b0 , \6362_b0 , w_20289 );
and ( w_20288 ,  , w_20289 );
buf ( w_20287 , \6363_b1 );
not ( w_20287 , w_20290 );
not (  , w_20291 );
and ( w_20290 , w_20291 , \6363_b0 );
buf ( \6365_b1 , \6364_b1 );
not ( \6365_b1 , w_20292 );
not ( \6365_b0 , w_20293 );
and ( w_20292 , w_20293 , \6364_b0 );
buf ( \6366_b1 , \4085_b1 );
not ( \6366_b1 , w_20294 );
not ( \6366_b0 , w_20295 );
and ( w_20294 , w_20295 , \4085_b0 );
or ( \6367_b1 , \6365_b1 , w_20296 );
or ( \6367_b0 , \6365_b0 , \6366_b0 );
not ( \6366_b0 , w_20297 );
and ( w_20297 , w_20296 , \6366_b1 );
or ( \6368_b1 , \4331_b1 , w_20299 );
not ( w_20299 , w_20300 );
and ( \6368_b0 , \4331_b0 , w_20301 );
and ( w_20300 ,  , w_20301 );
buf ( w_20299 , \6258_b1 );
not ( w_20299 , w_20302 );
not (  , w_20303 );
and ( w_20302 , w_20303 , \6258_b0 );
or ( \6369_b1 , \6367_b1 , w_20305 );
not ( w_20305 , w_20306 );
and ( \6369_b0 , \6367_b0 , w_20307 );
and ( w_20306 ,  , w_20307 );
buf ( w_20305 , \6368_b1 );
not ( w_20305 , w_20308 );
not (  , w_20309 );
and ( w_20308 , w_20309 , \6368_b0 );
buf ( \6370_b1 , \6369_b1 );
not ( \6370_b1 , w_20310 );
not ( \6370_b0 , w_20311 );
and ( w_20310 , w_20311 , \6369_b0 );
or ( \6371_b1 , \6359_b1 , w_20312 );
or ( \6371_b0 , \6359_b0 , \6370_b0 );
not ( \6370_b0 , w_20313 );
and ( w_20313 , w_20312 , \6370_b1 );
buf ( \6372_b1 , \6345_b1 );
not ( \6372_b1 , w_20314 );
not ( \6372_b0 , w_20315 );
and ( w_20314 , w_20315 , \6345_b0 );
or ( \6373_b1 , \6372_b1 , w_20317 );
not ( w_20317 , w_20318 );
and ( \6373_b0 , \6372_b0 , w_20319 );
and ( w_20318 ,  , w_20319 );
buf ( w_20317 , \6356_b1 );
not ( w_20317 , w_20320 );
not (  , w_20321 );
and ( w_20320 , w_20321 , \6356_b0 );
or ( \6374_b1 , \6371_b1 , w_20323 );
not ( w_20323 , w_20324 );
and ( \6374_b0 , \6371_b0 , w_20325 );
and ( w_20324 ,  , w_20325 );
buf ( w_20323 , \6373_b1 );
not ( w_20323 , w_20326 );
not (  , w_20327 );
and ( w_20326 , w_20327 , \6373_b0 );
or ( \6375_b1 , \6343_b1 , \6374_b1 );
not ( \6374_b1 , w_20328 );
and ( \6375_b0 , \6343_b0 , w_20329 );
and ( w_20328 , w_20329 , \6374_b0 );
or ( \6376_b1 , \6341_b1 , \6342_b1 );
not ( \6342_b1 , w_20330 );
and ( \6376_b0 , \6341_b0 , w_20331 );
and ( w_20330 , w_20331 , \6342_b0 );
or ( \6377_b1 , \6375_b1 , w_20332 );
or ( \6377_b0 , \6375_b0 , \6376_b0 );
not ( \6376_b0 , w_20333 );
and ( w_20333 , w_20332 , \6376_b1 );
buf ( \6378_b1 , \6377_b1 );
buf ( \6378_b0 , \6377_b0 );
or ( \6379_b1 , \6294_b1 , w_20334 );
xor ( \6379_b0 , \6294_b0 , w_20336 );
not ( w_20336 , w_20337 );
and ( w_20337 , w_20334 , w_20335 );
buf ( w_20334 , \6303_b1 );
not ( w_20334 , w_20338 );
not ( w_20335 , w_20339 );
and ( w_20338 , w_20339 , \6303_b0 );
or ( \6380_b1 , \6379_b1 , w_20340 );
xor ( \6380_b0 , \6379_b0 , w_20342 );
not ( w_20342 , w_20343 );
and ( w_20343 , w_20340 , w_20341 );
buf ( w_20340 , \6316_b1 );
not ( w_20340 , w_20344 );
not ( w_20341 , w_20345 );
and ( w_20344 , w_20345 , \6316_b0 );
buf ( \6381_b1 , \6380_b1 );
not ( \6381_b1 , w_20346 );
not ( \6381_b0 , w_20347 );
and ( w_20346 , w_20347 , \6380_b0 );
or ( \6382_b1 , \6378_b1 , w_20349 );
not ( w_20349 , w_20350 );
and ( \6382_b0 , \6378_b0 , w_20351 );
and ( w_20350 ,  , w_20351 );
buf ( w_20349 , \6381_b1 );
not ( w_20349 , w_20352 );
not (  , w_20353 );
and ( w_20352 , w_20353 , \6381_b0 );
buf ( \6383_b1 , \6382_b1 );
not ( \6383_b1 , w_20354 );
not ( \6383_b0 , w_20355 );
and ( w_20354 , w_20355 , \6382_b0 );
or ( \6384_b1 , \6331_b1 , \6383_b1 );
not ( \6383_b1 , w_20356 );
and ( \6384_b0 , \6331_b0 , w_20357 );
and ( w_20356 , w_20357 , \6383_b0 );
or ( \6385_b1 , \6378_b1 , \6381_b1 );
not ( \6381_b1 , w_20358 );
and ( \6385_b0 , \6378_b0 , w_20359 );
and ( w_20358 , w_20359 , \6381_b0 );
or ( \6386_b1 , \6384_b1 , w_20361 );
not ( w_20361 , w_20362 );
and ( \6386_b0 , \6384_b0 , w_20363 );
and ( w_20362 ,  , w_20363 );
buf ( w_20361 , \6385_b1 );
not ( w_20361 , w_20364 );
not (  , w_20365 );
and ( w_20364 , w_20365 , \6385_b0 );
or ( \6387_b1 , \6327_b1 , w_20367 );
not ( w_20367 , w_20368 );
and ( \6387_b0 , \6327_b0 , w_20369 );
and ( w_20368 ,  , w_20369 );
buf ( w_20367 , \6386_b1 );
not ( w_20367 , w_20370 );
not (  , w_20371 );
and ( w_20370 , w_20371 , \6386_b0 );
or ( \6388_b1 , \6240_b1 , \6252_b1 );
xor ( \6388_b0 , \6240_b0 , w_20372 );
not ( w_20372 , w_20373 );
and ( w_20373 , \6252_b1 , \6252_b0 );
or ( \6389_b1 , \6388_b1 , \6268_b1 );
xor ( \6389_b0 , \6388_b0 , w_20374 );
not ( w_20374 , w_20375 );
and ( w_20375 , \6268_b1 , \6268_b0 );
buf ( \6390_b1 , \4023_b1 );
not ( \6390_b1 , w_20376 );
not ( \6390_b0 , w_20377 );
and ( w_20376 , w_20377 , \4023_b0 );
buf ( \6391_b1 , \4069_b1 );
not ( \6391_b1 , w_20378 );
not ( \6391_b0 , w_20379 );
and ( w_20378 , w_20379 , \4069_b0 );
or ( \6392_b1 , \6390_b1 , w_20380 );
or ( \6392_b0 , \6390_b0 , \6391_b0 );
not ( \6391_b0 , w_20381 );
and ( w_20381 , w_20380 , \6391_b1 );
or ( \6393_b1 , \4407_b1 , w_20383 );
not ( w_20383 , w_20384 );
and ( \6393_b0 , \4407_b0 , w_20385 );
and ( w_20384 ,  , w_20385 );
buf ( w_20383 , \5131_b1 );
not ( w_20383 , w_20386 );
not (  , w_20387 );
and ( w_20386 , w_20387 , \5131_b0 );
or ( \6394_b1 , \6392_b1 , w_20389 );
not ( w_20389 , w_20390 );
and ( \6394_b0 , \6392_b0 , w_20391 );
and ( w_20390 ,  , w_20391 );
buf ( w_20389 , \6393_b1 );
not ( w_20389 , w_20392 );
not (  , w_20393 );
and ( w_20392 , w_20393 , \6393_b0 );
buf ( \6395_b1 , \6394_b1 );
not ( \6395_b1 , w_20394 );
not ( \6395_b0 , w_20395 );
and ( w_20394 , w_20395 , \6394_b0 );
buf ( \6396_b1 , \4065_b1 );
not ( \6396_b1 , w_20396 );
not ( \6396_b0 , w_20397 );
and ( w_20396 , w_20397 , \4065_b0 );
or ( \6397_b1 , \6395_b1 , w_20398 );
or ( \6397_b0 , \6395_b0 , \6396_b0 );
not ( \6396_b0 , w_20399 );
and ( w_20399 , w_20398 , \6396_b1 );
or ( \6398_b1 , \4055_b1 , w_20401 );
not ( w_20401 , w_20402 );
and ( \6398_b0 , \4055_b0 , w_20403 );
and ( w_20402 ,  , w_20403 );
buf ( w_20401 , \6336_b1 );
not ( w_20401 , w_20404 );
not (  , w_20405 );
and ( w_20404 , w_20405 , \6336_b0 );
or ( \6399_b1 , \6397_b1 , w_20407 );
not ( w_20407 , w_20408 );
and ( \6399_b0 , \6397_b0 , w_20409 );
and ( w_20408 ,  , w_20409 );
buf ( w_20407 , \6398_b1 );
not ( w_20407 , w_20410 );
not (  , w_20411 );
and ( w_20410 , w_20411 , \6398_b0 );
buf ( \6400_b1 , \6399_b1 );
not ( \6400_b1 , w_20412 );
not ( \6400_b0 , w_20413 );
and ( w_20412 , w_20413 , \6399_b0 );
buf ( \6401_b1 , \5019_b1 );
not ( \6401_b1 , w_20414 );
not ( \6401_b0 , w_20415 );
and ( w_20414 , w_20415 , \5019_b0 );
buf ( \6402_b1 , \3958_b1 );
not ( \6402_b1 , w_20416 );
not ( \6402_b0 , w_20417 );
and ( w_20416 , w_20417 , \3958_b0 );
buf ( \6403_b1 , \5874_b1 );
not ( \6403_b1 , w_20418 );
not ( \6403_b0 , w_20419 );
and ( w_20418 , w_20419 , \5874_b0 );
or ( \6404_b1 , \6402_b1 , w_20420 );
or ( \6404_b0 , \6402_b0 , \6403_b0 );
not ( \6403_b0 , w_20421 );
and ( w_20421 , w_20420 , \6403_b1 );
or ( \6405_b1 , \5873_b1 , w_20423 );
not ( w_20423 , w_20424 );
and ( \6405_b0 , \5873_b0 , w_20425 );
and ( w_20424 ,  , w_20425 );
buf ( w_20423 , \4473_b1 );
not ( w_20423 , w_20426 );
not (  , w_20427 );
and ( w_20426 , w_20427 , \4473_b0 );
or ( \6406_b1 , \6404_b1 , w_20429 );
not ( w_20429 , w_20430 );
and ( \6406_b0 , \6404_b0 , w_20431 );
and ( w_20430 ,  , w_20431 );
buf ( w_20429 , \6405_b1 );
not ( w_20429 , w_20432 );
not (  , w_20433 );
and ( w_20432 , w_20433 , \6405_b0 );
buf ( \6407_b1 , \6406_b1 );
not ( \6407_b1 , w_20434 );
not ( \6407_b0 , w_20435 );
and ( w_20434 , w_20435 , \6406_b0 );
or ( \6408_b1 , \6401_b1 , w_20436 );
or ( \6408_b0 , \6401_b0 , \6407_b0 );
not ( \6407_b0 , w_20437 );
and ( w_20437 , w_20436 , \6407_b1 );
or ( \6409_b1 , \6352_b1 , w_20439 );
not ( w_20439 , w_20440 );
and ( \6409_b0 , \6352_b0 , w_20441 );
and ( w_20440 ,  , w_20441 );
buf ( w_20439 , \5021_b1 );
not ( w_20439 , w_20442 );
not (  , w_20443 );
and ( w_20442 , w_20443 , \5021_b0 );
or ( \6410_b1 , \6408_b1 , w_20445 );
not ( w_20445 , w_20446 );
and ( \6410_b0 , \6408_b0 , w_20447 );
and ( w_20446 ,  , w_20447 );
buf ( w_20445 , \6409_b1 );
not ( w_20445 , w_20448 );
not (  , w_20449 );
and ( w_20448 , w_20449 , \6409_b0 );
or ( \6411_b1 , \4076_b1 , w_20451 );
not ( w_20451 , w_20452 );
and ( \6411_b0 , \4076_b0 , w_20453 );
and ( w_20452 ,  , w_20453 );
buf ( w_20451 , \5388_b1 );
not ( w_20451 , w_20454 );
not (  , w_20455 );
and ( w_20454 , w_20455 , \5388_b0 );
or ( \6412_b1 , \5749_b1 , \6411_b1 );
not ( \6411_b1 , w_20456 );
and ( \6412_b0 , \5749_b0 , w_20457 );
and ( w_20456 , w_20457 , \6411_b0 );
buf ( \6413_b1 , \4048_b1 );
not ( \6413_b1 , w_20458 );
not ( \6413_b0 , w_20459 );
and ( w_20458 , w_20459 , \4048_b0 );
buf ( \6414_b1 , \3272_b1 );
not ( \6414_b1 , w_20460 );
not ( \6414_b0 , w_20461 );
and ( w_20460 , w_20461 , \3272_b0 );
or ( \6415_b1 , \6413_b1 , w_20462 );
or ( \6415_b0 , \6413_b0 , \6414_b0 );
not ( \6414_b0 , w_20463 );
and ( w_20463 , w_20462 , \6414_b1 );
or ( \6416_b1 , \6415_b1 , w_20465 );
not ( w_20465 , w_20466 );
and ( \6416_b0 , \6415_b0 , w_20467 );
and ( w_20466 ,  , w_20467 );
buf ( w_20465 , \4088_b1 );
not ( w_20465 , w_20468 );
not (  , w_20469 );
and ( w_20468 , w_20469 , \4088_b0 );
or ( \6417_b1 , \6412_b1 , w_20471 );
not ( w_20471 , w_20472 );
and ( \6417_b0 , \6412_b0 , w_20473 );
and ( w_20472 ,  , w_20473 );
buf ( w_20471 , \6416_b1 );
not ( w_20471 , w_20474 );
not (  , w_20475 );
and ( w_20474 , w_20475 , \6416_b0 );
or ( \6418_b1 , \6410_b1 , w_20477 );
not ( w_20477 , w_20478 );
and ( \6418_b0 , \6410_b0 , w_20479 );
and ( w_20478 ,  , w_20479 );
buf ( w_20477 , \6417_b1 );
not ( w_20477 , w_20480 );
not (  , w_20481 );
and ( w_20480 , w_20481 , \6417_b0 );
or ( \6419_b1 , \6400_b1 , w_20483 );
not ( w_20483 , w_20484 );
and ( \6419_b0 , \6400_b0 , w_20485 );
and ( w_20484 ,  , w_20485 );
buf ( w_20483 , \6418_b1 );
not ( w_20483 , w_20486 );
not (  , w_20487 );
and ( w_20486 , w_20487 , \6418_b0 );
buf ( \6420_b1 , \6419_b1 );
not ( \6420_b1 , w_20488 );
not ( \6420_b0 , w_20489 );
and ( w_20488 , w_20489 , \6419_b0 );
buf ( \6421_b1 , \4662_b1 );
not ( \6421_b1 , w_20490 );
not ( \6421_b0 , w_20491 );
and ( w_20490 , w_20491 , \4662_b0 );
buf ( \6422_b1 , \3963_b1 );
not ( \6422_b1 , w_20492 );
not ( \6422_b0 , w_20493 );
and ( w_20492 , w_20493 , \3963_b0 );
buf ( \6423_b1 , \4666_b1 );
not ( \6423_b1 , w_20494 );
not ( \6423_b0 , w_20495 );
and ( w_20494 , w_20495 , \4666_b0 );
or ( \6424_b1 , \6422_b1 , w_20496 );
or ( \6424_b0 , \6422_b0 , \6423_b0 );
not ( \6423_b0 , w_20497 );
and ( w_20497 , w_20496 , \6423_b1 );
or ( \6425_b1 , \4665_b1 , w_20499 );
not ( w_20499 , w_20500 );
and ( \6425_b0 , \4665_b0 , w_20501 );
and ( w_20500 ,  , w_20501 );
buf ( w_20499 , \4486_b1 );
not ( w_20499 , w_20502 );
not (  , w_20503 );
and ( w_20502 , w_20503 , \4486_b0 );
or ( \6426_b1 , \6424_b1 , w_20505 );
not ( w_20505 , w_20506 );
and ( \6426_b0 , \6424_b0 , w_20507 );
and ( w_20506 ,  , w_20507 );
buf ( w_20505 , \6425_b1 );
not ( w_20505 , w_20508 );
not (  , w_20509 );
and ( w_20508 , w_20509 , \6425_b0 );
buf ( \6427_b1 , \6426_b1 );
not ( \6427_b1 , w_20510 );
not ( \6427_b0 , w_20511 );
and ( w_20510 , w_20511 , \6426_b0 );
or ( \6428_b1 , \6421_b1 , w_20512 );
or ( \6428_b0 , \6421_b0 , \6427_b0 );
not ( \6427_b0 , w_20513 );
and ( w_20513 , w_20512 , \6427_b1 );
or ( \6429_b1 , \5187_b1 , w_20515 );
not ( w_20515 , w_20516 );
and ( \6429_b0 , \5187_b0 , w_20517 );
and ( w_20516 ,  , w_20517 );
buf ( w_20515 , \6214_b1 );
not ( w_20515 , w_20518 );
not (  , w_20519 );
and ( w_20518 , w_20519 , \6214_b0 );
or ( \6430_b1 , \6428_b1 , w_20521 );
not ( w_20521 , w_20522 );
and ( \6430_b0 , \6428_b0 , w_20523 );
and ( w_20522 ,  , w_20523 );
buf ( w_20521 , \6429_b1 );
not ( w_20521 , w_20524 );
not (  , w_20525 );
and ( w_20524 , w_20525 , \6429_b0 );
buf ( \6431_b1 , \6430_b1 );
not ( \6431_b1 , w_20526 );
not ( \6431_b0 , w_20527 );
and ( w_20526 , w_20527 , \6430_b0 );
or ( \6432_b1 , \6420_b1 , w_20528 );
or ( \6432_b0 , \6420_b0 , \6431_b0 );
not ( \6431_b0 , w_20529 );
and ( w_20529 , w_20528 , \6431_b1 );
buf ( \6433_b1 , \6418_b1 );
not ( \6433_b1 , w_20530 );
not ( \6433_b0 , w_20531 );
and ( w_20530 , w_20531 , \6418_b0 );
or ( \6434_b1 , \6433_b1 , w_20533 );
not ( w_20533 , w_20534 );
and ( \6434_b0 , \6433_b0 , w_20535 );
and ( w_20534 ,  , w_20535 );
buf ( w_20533 , \6399_b1 );
not ( w_20533 , w_20536 );
not (  , w_20537 );
and ( w_20536 , w_20537 , \6399_b0 );
or ( \6435_b1 , \6432_b1 , w_20539 );
not ( w_20539 , w_20540 );
and ( \6435_b0 , \6432_b0 , w_20541 );
and ( w_20540 ,  , w_20541 );
buf ( w_20539 , \6434_b1 );
not ( w_20539 , w_20542 );
not (  , w_20543 );
and ( w_20542 , w_20543 , \6434_b0 );
or ( \6436_b1 , \6389_b1 , \6435_b1 );
xor ( \6436_b0 , \6389_b0 , w_20544 );
not ( w_20544 , w_20545 );
and ( w_20545 , \6435_b1 , \6435_b0 );
or ( \6437_b1 , \6341_b1 , \6342_b1 );
xor ( \6437_b0 , \6341_b0 , w_20546 );
not ( w_20546 , w_20547 );
and ( w_20547 , \6342_b1 , \6342_b0 );
or ( \6438_b1 , \6437_b1 , \6374_b1 );
xor ( \6438_b0 , \6437_b0 , w_20548 );
not ( w_20548 , w_20549 );
and ( w_20549 , \6374_b1 , \6374_b0 );
or ( \6439_b1 , \6436_b1 , \6438_b1 );
not ( \6438_b1 , w_20550 );
and ( \6439_b0 , \6436_b0 , w_20551 );
and ( w_20550 , w_20551 , \6438_b0 );
buf ( \6440_b1 , \6436_b1 );
not ( \6440_b1 , w_20552 );
not ( \6440_b0 , w_20553 );
and ( w_20552 , w_20553 , \6436_b0 );
buf ( \6441_b1 , \6438_b1 );
not ( \6441_b1 , w_20554 );
not ( \6441_b0 , w_20555 );
and ( w_20554 , w_20555 , \6438_b0 );
or ( \6442_b1 , \6440_b1 , \6441_b1 );
not ( \6441_b1 , w_20556 );
and ( \6442_b0 , \6440_b0 , w_20557 );
and ( w_20556 , w_20557 , \6441_b0 );
or ( \6443_b1 , \6439_b1 , w_20559 );
not ( w_20559 , w_20560 );
and ( \6443_b0 , \6439_b0 , w_20561 );
and ( w_20560 ,  , w_20561 );
buf ( w_20559 , \6442_b1 );
not ( w_20559 , w_20562 );
not (  , w_20563 );
and ( w_20562 , w_20563 , \6442_b0 );
buf ( \6444_b1 , \6357_b1 );
not ( \6444_b1 , w_20564 );
not ( \6444_b0 , w_20565 );
and ( w_20564 , w_20565 , \6357_b0 );
buf ( \6445_b1 , \6345_b1 );
not ( \6445_b1 , w_20566 );
not ( \6445_b0 , w_20567 );
and ( w_20566 , w_20567 , \6345_b0 );
buf ( \6446_b1 , \6445_b1 );
not ( \6446_b1 , w_20568 );
not ( \6446_b0 , w_20569 );
and ( w_20568 , w_20569 , \6445_b0 );
or ( \6447_b1 , \6444_b1 , w_20570 );
or ( \6447_b0 , \6444_b0 , \6446_b0 );
not ( \6446_b0 , w_20571 );
and ( w_20571 , w_20570 , \6446_b1 );
or ( \6448_b1 , \6372_b1 , w_20572 );
or ( \6448_b0 , \6372_b0 , \6357_b0 );
not ( \6357_b0 , w_20573 );
and ( w_20573 , w_20572 , \6357_b1 );
or ( \6449_b1 , \6447_b1 , w_20575 );
not ( w_20575 , w_20576 );
and ( \6449_b0 , \6447_b0 , w_20577 );
and ( w_20576 ,  , w_20577 );
buf ( w_20575 , \6448_b1 );
not ( w_20575 , w_20578 );
not (  , w_20579 );
and ( w_20578 , w_20579 , \6448_b0 );
or ( \6450_b1 , \6449_b1 , \6369_b1 );
xor ( \6450_b0 , \6449_b0 , w_20580 );
not ( w_20580 , w_20581 );
and ( w_20581 , \6369_b1 , \6369_b0 );
buf ( \6451_b1 , \5388_b1 );
not ( \6451_b1 , w_20582 );
not ( \6451_b0 , w_20583 );
and ( w_20582 , w_20583 , \5388_b0 );
buf ( \6452_b1 , \4088_b1 );
not ( \6452_b1 , w_20584 );
not ( \6452_b0 , w_20585 );
and ( w_20584 , w_20585 , \4088_b0 );
or ( \6453_b1 , \6451_b1 , w_20586 );
or ( \6453_b0 , \6451_b0 , \6452_b0 );
not ( \6452_b0 , w_20587 );
and ( w_20587 , w_20586 , \6452_b1 );
or ( \6454_b1 , \4089_b1 , w_20589 );
not ( w_20589 , w_20590 );
and ( \6454_b0 , \4089_b0 , w_20591 );
and ( w_20590 ,  , w_20591 );
buf ( w_20589 , \4048_b1 );
not ( w_20589 , w_20592 );
not (  , w_20593 );
and ( w_20592 , w_20593 , \4048_b0 );
or ( \6455_b1 , \6453_b1 , w_20595 );
not ( w_20595 , w_20596 );
and ( \6455_b0 , \6453_b0 , w_20597 );
and ( w_20596 ,  , w_20597 );
buf ( w_20595 , \6454_b1 );
not ( w_20595 , w_20598 );
not (  , w_20599 );
and ( w_20598 , w_20599 , \6454_b0 );
or ( \6456_b1 , \4086_b1 , \6455_b1 );
not ( \6455_b1 , w_20600 );
and ( \6456_b0 , \4086_b0 , w_20601 );
and ( w_20600 , w_20601 , \6455_b0 );
buf ( \6457_b1 , \5241_b1 );
not ( \6457_b1 , w_20602 );
not ( \6457_b0 , w_20603 );
and ( w_20602 , w_20603 , \5241_b0 );
or ( \6458_b1 , \6457_b1 , \6364_b1 );
not ( \6364_b1 , w_20604 );
and ( \6458_b0 , \6457_b0 , w_20605 );
and ( w_20604 , w_20605 , \6364_b0 );
or ( \6459_b1 , \6456_b1 , w_20607 );
not ( w_20607 , w_20608 );
and ( \6459_b0 , \6456_b0 , w_20609 );
and ( w_20608 ,  , w_20609 );
buf ( w_20607 , \6458_b1 );
not ( w_20607 , w_20610 );
not (  , w_20611 );
and ( w_20610 , w_20611 , \6458_b0 );
buf ( \6460_b1 , \6459_b1 );
not ( \6460_b1 , w_20612 );
not ( \6460_b0 , w_20613 );
and ( w_20612 , w_20613 , \6459_b0 );
buf ( \6461_b1 , \6460_b1 );
not ( \6461_b1 , w_20614 );
not ( \6461_b0 , w_20615 );
and ( w_20614 , w_20615 , \6460_b0 );
buf ( \6462_b1 , \4026_b1 );
not ( \6462_b1 , w_20616 );
not ( \6462_b0 , w_20617 );
and ( w_20616 , w_20617 , \4026_b0 );
buf ( \6463_b1 , \4069_b1 );
not ( \6463_b1 , w_20618 );
not ( \6463_b0 , w_20619 );
and ( w_20618 , w_20619 , \4069_b0 );
or ( \6464_b1 , \6462_b1 , w_20620 );
or ( \6464_b0 , \6462_b0 , \6463_b0 );
not ( \6463_b0 , w_20621 );
and ( w_20621 , w_20620 , \6463_b1 );
or ( \6465_b1 , \5749_b1 , w_20623 );
not ( w_20623 , w_20624 );
and ( \6465_b0 , \5749_b0 , w_20625 );
and ( w_20624 ,  , w_20625 );
buf ( w_20623 , \5344_b1 );
not ( w_20623 , w_20626 );
not (  , w_20627 );
and ( w_20626 , w_20627 , \5344_b0 );
or ( \6466_b1 , \6464_b1 , w_20629 );
not ( w_20629 , w_20630 );
and ( \6466_b0 , \6464_b0 , w_20631 );
and ( w_20630 ,  , w_20631 );
buf ( w_20629 , \6465_b1 );
not ( w_20629 , w_20632 );
not (  , w_20633 );
and ( w_20632 , w_20633 , \6465_b0 );
or ( \6467_b1 , \6466_b1 , \4065_b1 );
not ( \4065_b1 , w_20634 );
and ( \6467_b0 , \6466_b0 , w_20635 );
and ( w_20634 , w_20635 , \4065_b0 );
or ( \6468_b1 , \4562_b1 , \6394_b1 );
not ( \6394_b1 , w_20636 );
and ( \6468_b0 , \4562_b0 , w_20637 );
and ( w_20636 , w_20637 , \6394_b0 );
or ( \6469_b1 , \6467_b1 , w_20639 );
not ( w_20639 , w_20640 );
and ( \6469_b0 , \6467_b0 , w_20641 );
and ( w_20640 ,  , w_20641 );
buf ( w_20639 , \6468_b1 );
not ( w_20639 , w_20642 );
not (  , w_20643 );
and ( w_20642 , w_20643 , \6468_b0 );
buf ( \6470_b1 , \6469_b1 );
not ( \6470_b1 , w_20644 );
not ( \6470_b0 , w_20645 );
and ( w_20644 , w_20645 , \6469_b0 );
buf ( \6471_b1 , \6470_b1 );
not ( \6471_b1 , w_20646 );
not ( \6471_b0 , w_20647 );
and ( w_20646 , w_20647 , \6470_b0 );
or ( \6472_b1 , \6461_b1 , w_20648 );
or ( \6472_b0 , \6461_b0 , \6471_b0 );
not ( \6471_b0 , w_20649 );
and ( w_20649 , w_20648 , \6471_b1 );
buf ( \6473_b1 , \6459_b1 );
not ( \6473_b1 , w_20650 );
not ( \6473_b0 , w_20651 );
and ( w_20650 , w_20651 , \6459_b0 );
buf ( \6474_b1 , \6469_b1 );
not ( \6474_b1 , w_20652 );
not ( \6474_b0 , w_20653 );
and ( w_20652 , w_20653 , \6469_b0 );
or ( \6475_b1 , \6473_b1 , w_20654 );
or ( \6475_b0 , \6473_b0 , \6474_b0 );
not ( \6474_b0 , w_20655 );
and ( w_20655 , w_20654 , \6474_b1 );
buf ( \6476_b1 , \4019_b1 );
not ( \6476_b1 , w_20656 );
not ( \6476_b0 , w_20657 );
and ( w_20656 , w_20657 , \4019_b0 );
buf ( \6477_b1 , \5178_b1 );
not ( \6477_b1 , w_20658 );
not ( \6477_b0 , w_20659 );
and ( w_20658 , w_20659 , \5178_b0 );
or ( \6478_b1 , \6476_b1 , w_20660 );
or ( \6478_b0 , \6476_b0 , \6477_b0 );
not ( \6477_b0 , w_20661 );
and ( w_20661 , w_20660 , \6477_b1 );
or ( \6479_b1 , \4665_b1 , w_20663 );
not ( w_20663 , w_20664 );
and ( \6479_b0 , \4665_b0 , w_20665 );
and ( w_20664 ,  , w_20665 );
buf ( w_20663 , \4585_b1 );
not ( w_20663 , w_20666 );
not (  , w_20667 );
and ( w_20666 , w_20667 , \4585_b0 );
or ( \6480_b1 , \6478_b1 , w_20669 );
not ( w_20669 , w_20670 );
and ( \6480_b0 , \6478_b0 , w_20671 );
and ( w_20670 ,  , w_20671 );
buf ( w_20669 , \6479_b1 );
not ( w_20669 , w_20672 );
not (  , w_20673 );
and ( w_20672 , w_20673 , \6479_b0 );
buf ( \6481_b1 , \6480_b1 );
not ( \6481_b1 , w_20674 );
not ( \6481_b0 , w_20675 );
and ( w_20674 , w_20675 , \6480_b0 );
buf ( \6482_b1 , \4662_b1 );
not ( \6482_b1 , w_20676 );
not ( \6482_b0 , w_20677 );
and ( w_20676 , w_20677 , \4662_b0 );
or ( \6483_b1 , \6481_b1 , w_20678 );
or ( \6483_b0 , \6481_b0 , \6482_b0 );
not ( \6482_b0 , w_20679 );
and ( w_20679 , w_20678 , \6482_b1 );
or ( \6484_b1 , \5187_b1 , w_20681 );
not ( w_20681 , w_20682 );
and ( \6484_b0 , \5187_b0 , w_20683 );
and ( w_20682 ,  , w_20683 );
buf ( w_20681 , \6426_b1 );
not ( w_20681 , w_20684 );
not (  , w_20685 );
and ( w_20684 , w_20685 , \6426_b0 );
or ( \6485_b1 , \6483_b1 , w_20687 );
not ( w_20687 , w_20688 );
and ( \6485_b0 , \6483_b0 , w_20689 );
and ( w_20688 ,  , w_20689 );
buf ( w_20687 , \6484_b1 );
not ( w_20687 , w_20690 );
not (  , w_20691 );
and ( w_20690 , w_20691 , \6484_b0 );
or ( \6486_b1 , \6475_b1 , w_20693 );
not ( w_20693 , w_20694 );
and ( \6486_b0 , \6475_b0 , w_20695 );
and ( w_20694 ,  , w_20695 );
buf ( w_20693 , \6485_b1 );
not ( w_20693 , w_20696 );
not (  , w_20697 );
and ( w_20696 , w_20697 , \6485_b0 );
or ( \6487_b1 , \6472_b1 , w_20699 );
not ( w_20699 , w_20700 );
and ( \6487_b0 , \6472_b0 , w_20701 );
and ( w_20700 ,  , w_20701 );
buf ( w_20699 , \6486_b1 );
not ( w_20699 , w_20702 );
not (  , w_20703 );
and ( w_20702 , w_20703 , \6486_b0 );
or ( \6488_b1 , \6450_b1 , \6487_b1 );
xor ( \6488_b0 , \6450_b0 , w_20704 );
not ( w_20704 , w_20705 );
and ( w_20705 , \6487_b1 , \6487_b0 );
or ( \6489_b1 , \6418_b1 , \6399_b1 );
xor ( \6489_b0 , \6418_b0 , w_20706 );
not ( w_20706 , w_20707 );
and ( w_20707 , \6399_b1 , \6399_b0 );
or ( \6490_b1 , \6489_b1 , w_20708 );
xor ( \6490_b0 , \6489_b0 , w_20710 );
not ( w_20710 , w_20711 );
and ( w_20711 , w_20708 , w_20709 );
buf ( w_20708 , \6430_b1 );
not ( w_20708 , w_20712 );
not ( w_20709 , w_20713 );
and ( w_20712 , w_20713 , \6430_b0 );
or ( \6491_b1 , \6488_b1 , \6490_b1 );
not ( \6490_b1 , w_20714 );
and ( \6491_b0 , \6488_b0 , w_20715 );
and ( w_20714 , w_20715 , \6490_b0 );
or ( \6492_b1 , \6450_b1 , \6487_b1 );
not ( \6487_b1 , w_20716 );
and ( \6492_b0 , \6450_b0 , w_20717 );
and ( w_20716 , w_20717 , \6487_b0 );
or ( \6493_b1 , \6491_b1 , w_20718 );
or ( \6493_b0 , \6491_b0 , \6492_b0 );
not ( \6492_b0 , w_20719 );
and ( w_20719 , w_20718 , \6492_b1 );
or ( \6494_b1 , \6443_b1 , w_20721 );
not ( w_20721 , w_20722 );
and ( \6494_b0 , \6443_b0 , w_20723 );
and ( w_20722 ,  , w_20723 );
buf ( w_20721 , \6493_b1 );
not ( w_20721 , w_20724 );
not (  , w_20725 );
and ( w_20724 , w_20725 , \6493_b0 );
buf ( \6495_b1 , \6494_b1 );
not ( \6495_b1 , w_20726 );
not ( \6495_b0 , w_20727 );
and ( w_20726 , w_20727 , \6494_b0 );
or ( \6496_b1 , \6450_b1 , \6487_b1 );
xor ( \6496_b0 , \6450_b0 , w_20728 );
not ( w_20728 , w_20729 );
and ( w_20729 , \6487_b1 , \6487_b0 );
or ( \6497_b1 , \6496_b1 , \6490_b1 );
xor ( \6497_b0 , \6496_b0 , w_20730 );
not ( w_20730 , w_20731 );
and ( w_20731 , \6490_b1 , \6490_b0 );
or ( \6498_b1 , \4103_b1 , w_20733 );
not ( w_20733 , w_20734 );
and ( \6498_b0 , \4103_b0 , w_20735 );
and ( w_20734 ,  , w_20735 );
buf ( w_20733 , \5388_b1 );
not ( w_20733 , w_20736 );
not (  , w_20737 );
and ( w_20736 , w_20737 , \5388_b0 );
buf ( \6499_b1 , \3963_b1 );
not ( \6499_b1 , w_20738 );
not ( \6499_b0 , w_20739 );
and ( w_20738 , w_20739 , \3963_b0 );
buf ( \6500_b1 , \5023_b1 );
not ( \6500_b1 , w_20740 );
not ( \6500_b0 , w_20741 );
and ( w_20740 , w_20741 , \5023_b0 );
or ( \6501_b1 , \6499_b1 , w_20742 );
or ( \6501_b0 , \6499_b0 , \6500_b0 );
not ( \6500_b0 , w_20743 );
and ( w_20743 , w_20742 , \6500_b1 );
buf ( \6502_b1 , \5576_b1 );
not ( \6502_b1 , w_20744 );
not ( \6502_b0 , w_20745 );
and ( w_20744 , w_20745 , \5576_b0 );
or ( \6503_b1 , \6502_b1 , w_20747 );
not ( w_20747 , w_20748 );
and ( \6503_b0 , \6502_b0 , w_20749 );
and ( w_20748 ,  , w_20749 );
buf ( w_20747 , \4486_b1 );
not ( w_20747 , w_20750 );
not (  , w_20751 );
and ( w_20750 , w_20751 , \4486_b0 );
or ( \6504_b1 , \6501_b1 , w_20753 );
not ( w_20753 , w_20754 );
and ( \6504_b0 , \6501_b0 , w_20755 );
and ( w_20754 ,  , w_20755 );
buf ( w_20753 , \6503_b1 );
not ( w_20753 , w_20756 );
not (  , w_20757 );
and ( w_20756 , w_20757 , \6503_b0 );
buf ( \6505_b1 , \6504_b1 );
not ( \6505_b1 , w_20758 );
not ( \6505_b0 , w_20759 );
and ( w_20758 , w_20759 , \6504_b0 );
buf ( \6506_b1 , \5020_b1 );
not ( \6506_b1 , w_20760 );
not ( \6506_b0 , w_20761 );
and ( w_20760 , w_20761 , \5020_b0 );
or ( \6507_b1 , \6505_b1 , w_20762 );
or ( \6507_b0 , \6505_b0 , \6506_b0 );
not ( \6506_b0 , w_20763 );
and ( w_20763 , w_20762 , \6506_b1 );
or ( \6508_b1 , \6406_b1 , w_20765 );
not ( w_20765 , w_20766 );
and ( \6508_b0 , \6406_b0 , w_20767 );
and ( w_20766 ,  , w_20767 );
buf ( w_20765 , \5021_b1 );
not ( w_20765 , w_20768 );
not (  , w_20769 );
and ( w_20768 , w_20769 , \5021_b0 );
or ( \6509_b1 , \6507_b1 , w_20771 );
not ( w_20771 , w_20772 );
and ( \6509_b0 , \6507_b0 , w_20773 );
and ( w_20772 ,  , w_20773 );
buf ( w_20771 , \6508_b1 );
not ( w_20771 , w_20774 );
not (  , w_20775 );
and ( w_20774 , w_20775 , \6508_b0 );
or ( \6510_b1 , \6498_b1 , \6509_b1 );
xor ( \6510_b0 , \6498_b0 , w_20776 );
not ( w_20776 , w_20777 );
and ( w_20777 , \6509_b1 , \6509_b0 );
buf ( \6511_b1 , \4662_b1 );
not ( \6511_b1 , w_20778 );
not ( \6511_b0 , w_20779 );
and ( w_20778 , w_20779 , \4662_b0 );
buf ( \6512_b1 , \4023_b1 );
not ( \6512_b1 , w_20780 );
not ( \6512_b0 , w_20781 );
and ( w_20780 , w_20781 , \4023_b0 );
buf ( \6513_b1 , \4666_b1 );
not ( \6513_b1 , w_20782 );
not ( \6513_b0 , w_20783 );
and ( w_20782 , w_20783 , \4666_b0 );
or ( \6514_b1 , \6512_b1 , w_20784 );
or ( \6514_b0 , \6512_b0 , \6513_b0 );
not ( \6513_b0 , w_20785 );
and ( w_20785 , w_20784 , \6513_b1 );
buf ( \6515_b1 , \5178_b1 );
not ( \6515_b1 , w_20786 );
not ( \6515_b0 , w_20787 );
and ( w_20786 , w_20787 , \5178_b0 );
or ( \6516_b1 , \6515_b1 , w_20789 );
not ( w_20789 , w_20790 );
and ( \6516_b0 , \6515_b0 , w_20791 );
and ( w_20790 ,  , w_20791 );
buf ( w_20789 , \5131_b1 );
not ( w_20789 , w_20792 );
not (  , w_20793 );
and ( w_20792 , w_20793 , \5131_b0 );
or ( \6517_b1 , \6514_b1 , w_20795 );
not ( w_20795 , w_20796 );
and ( \6517_b0 , \6514_b0 , w_20797 );
and ( w_20796 ,  , w_20797 );
buf ( w_20795 , \6516_b1 );
not ( w_20795 , w_20798 );
not (  , w_20799 );
and ( w_20798 , w_20799 , \6516_b0 );
buf ( \6518_b1 , \6517_b1 );
not ( \6518_b1 , w_20800 );
not ( \6518_b0 , w_20801 );
and ( w_20800 , w_20801 , \6517_b0 );
or ( \6519_b1 , \6511_b1 , w_20802 );
or ( \6519_b0 , \6511_b0 , \6518_b0 );
not ( \6518_b0 , w_20803 );
and ( w_20803 , w_20802 , \6518_b1 );
or ( \6520_b1 , \4672_b1 , w_20805 );
not ( w_20805 , w_20806 );
and ( \6520_b0 , \4672_b0 , w_20807 );
and ( w_20806 ,  , w_20807 );
buf ( w_20805 , \6480_b1 );
not ( w_20805 , w_20808 );
not (  , w_20809 );
and ( w_20808 , w_20809 , \6480_b0 );
or ( \6521_b1 , \6519_b1 , w_20811 );
not ( w_20811 , w_20812 );
and ( \6521_b0 , \6519_b0 , w_20813 );
and ( w_20812 ,  , w_20813 );
buf ( w_20811 , \6520_b1 );
not ( w_20811 , w_20814 );
not (  , w_20815 );
and ( w_20814 , w_20815 , \6520_b0 );
or ( \6522_b1 , \6510_b1 , \6521_b1 );
not ( \6521_b1 , w_20816 );
and ( \6522_b0 , \6510_b0 , w_20817 );
and ( w_20816 , w_20817 , \6521_b0 );
or ( \6523_b1 , \6498_b1 , \6509_b1 );
not ( \6509_b1 , w_20818 );
and ( \6523_b0 , \6498_b0 , w_20819 );
and ( w_20818 , w_20819 , \6509_b0 );
or ( \6524_b1 , \6522_b1 , w_20820 );
or ( \6524_b0 , \6522_b0 , \6523_b0 );
not ( \6523_b0 , w_20821 );
and ( w_20821 , w_20820 , \6523_b1 );
or ( \6525_b1 , \6410_b1 , \6417_b1 );
xor ( \6525_b0 , \6410_b0 , w_20822 );
not ( w_20822 , w_20823 );
and ( w_20823 , \6417_b1 , \6417_b0 );
or ( \6526_b1 , \6524_b1 , w_20824 );
or ( \6526_b0 , \6524_b0 , \6525_b0 );
not ( \6525_b0 , w_20825 );
and ( w_20825 , w_20824 , \6525_b1 );
buf ( \6527_b1 , \6526_b1 );
not ( \6527_b1 , w_20826 );
not ( \6527_b0 , w_20827 );
and ( w_20826 , w_20827 , \6526_b0 );
buf ( \6528_b1 , \6470_b1 );
not ( \6528_b1 , w_20828 );
not ( \6528_b0 , w_20829 );
and ( w_20828 , w_20829 , \6470_b0 );
buf ( \6529_b1 , \6485_b1 );
not ( \6529_b1 , w_20830 );
not ( \6529_b0 , w_20831 );
and ( w_20830 , w_20831 , \6485_b0 );
buf ( \6530_b1 , \6529_b1 );
not ( \6530_b1 , w_20832 );
not ( \6530_b0 , w_20833 );
and ( w_20832 , w_20833 , \6529_b0 );
or ( \6531_b1 , \6528_b1 , w_20834 );
or ( \6531_b0 , \6528_b0 , \6530_b0 );
not ( \6530_b0 , w_20835 );
and ( w_20835 , w_20834 , \6530_b1 );
or ( \6532_b1 , \6485_b1 , w_20837 );
not ( w_20837 , w_20838 );
and ( \6532_b0 , \6485_b0 , w_20839 );
and ( w_20838 ,  , w_20839 );
buf ( w_20837 , \6469_b1 );
not ( w_20837 , w_20840 );
not (  , w_20841 );
and ( w_20840 , w_20841 , \6469_b0 );
or ( \6533_b1 , \6531_b1 , w_20843 );
not ( w_20843 , w_20844 );
and ( \6533_b0 , \6531_b0 , w_20845 );
and ( w_20844 ,  , w_20845 );
buf ( w_20843 , \6532_b1 );
not ( w_20843 , w_20846 );
not (  , w_20847 );
and ( w_20846 , w_20847 , \6532_b0 );
or ( \6534_b1 , \6533_b1 , \6460_b1 );
not ( \6460_b1 , w_20848 );
and ( \6534_b0 , \6533_b0 , w_20849 );
and ( w_20848 , w_20849 , \6460_b0 );
buf ( \6535_b1 , \6533_b1 );
not ( \6535_b1 , w_20850 );
not ( \6535_b0 , w_20851 );
and ( w_20850 , w_20851 , \6533_b0 );
or ( \6536_b1 , \6535_b1 , \6459_b1 );
not ( \6459_b1 , w_20852 );
and ( \6536_b0 , \6535_b0 , w_20853 );
and ( w_20852 , w_20853 , \6459_b0 );
or ( \6537_b1 , \6534_b1 , w_20855 );
not ( w_20855 , w_20856 );
and ( \6537_b0 , \6534_b0 , w_20857 );
and ( w_20856 ,  , w_20857 );
buf ( w_20855 , \6536_b1 );
not ( w_20855 , w_20858 );
not (  , w_20859 );
and ( w_20858 , w_20859 , \6536_b0 );
buf ( \6538_b1 , \6537_b1 );
not ( \6538_b1 , w_20860 );
not ( \6538_b0 , w_20861 );
and ( w_20860 , w_20861 , \6537_b0 );
or ( \6539_b1 , \6527_b1 , w_20862 );
or ( \6539_b0 , \6527_b0 , \6538_b0 );
not ( \6538_b0 , w_20863 );
and ( w_20863 , w_20862 , \6538_b1 );
or ( \6540_b1 , \6524_b1 , w_20865 );
not ( w_20865 , w_20866 );
and ( \6540_b0 , \6524_b0 , w_20867 );
and ( w_20866 ,  , w_20867 );
buf ( w_20865 , \6525_b1 );
not ( w_20865 , w_20868 );
not (  , w_20869 );
and ( w_20868 , w_20869 , \6525_b0 );
or ( \6541_b1 , \6539_b1 , w_20871 );
not ( w_20871 , w_20872 );
and ( \6541_b0 , \6539_b0 , w_20873 );
and ( w_20872 ,  , w_20873 );
buf ( w_20871 , \6540_b1 );
not ( w_20871 , w_20874 );
not (  , w_20875 );
and ( w_20874 , w_20875 , \6540_b0 );
or ( \6542_b1 , \6497_b1 , w_20877 );
not ( w_20877 , w_20878 );
and ( \6542_b0 , \6497_b0 , w_20879 );
and ( w_20878 ,  , w_20879 );
buf ( w_20877 , \6541_b1 );
not ( w_20877 , w_20880 );
not (  , w_20881 );
and ( w_20880 , w_20881 , \6541_b0 );
buf ( \6543_b1 , \6542_b1 );
not ( \6543_b1 , w_20882 );
not ( \6543_b0 , w_20883 );
and ( w_20882 , w_20883 , \6542_b0 );
or ( \6544_b1 , \6495_b1 , w_20884 );
or ( \6544_b0 , \6495_b0 , \6543_b0 );
not ( \6543_b0 , w_20885 );
and ( w_20885 , w_20884 , \6543_b1 );
or ( \6545_b1 , \6443_b1 , w_20886 );
or ( \6545_b0 , \6443_b0 , \6493_b0 );
not ( \6493_b0 , w_20887 );
and ( w_20887 , w_20886 , \6493_b1 );
or ( \6546_b1 , \6544_b1 , w_20889 );
not ( w_20889 , w_20890 );
and ( \6546_b0 , \6544_b0 , w_20891 );
and ( w_20890 ,  , w_20891 );
buf ( w_20889 , \6545_b1 );
not ( w_20889 , w_20892 );
not (  , w_20893 );
and ( w_20892 , w_20893 , \6545_b0 );
buf ( \6547_b1 , \6377_b1 );
not ( \6547_b1 , w_20894 );
not ( \6547_b0 , w_20895 );
and ( w_20894 , w_20895 , \6377_b0 );
buf ( \6548_b1 , \6380_b1 );
not ( \6548_b1 , w_20896 );
not ( \6548_b0 , w_20897 );
and ( w_20896 , w_20897 , \6380_b0 );
or ( \6549_b1 , \6547_b1 , \6548_b1 );
not ( \6548_b1 , w_20898 );
and ( \6549_b0 , \6547_b0 , w_20899 );
and ( w_20898 , w_20899 , \6548_b0 );
or ( \6550_b1 , \6377_b1 , \6380_b1 );
not ( \6380_b1 , w_20900 );
and ( \6550_b0 , \6377_b0 , w_20901 );
and ( w_20900 , w_20901 , \6380_b0 );
or ( \6551_b1 , \6549_b1 , w_20903 );
not ( w_20903 , w_20904 );
and ( \6551_b0 , \6549_b0 , w_20905 );
and ( w_20904 ,  , w_20905 );
buf ( w_20903 , \6550_b1 );
not ( w_20903 , w_20906 );
not (  , w_20907 );
and ( w_20906 , w_20907 , \6550_b0 );
buf ( \6552_b1 , \6551_b1 );
not ( \6552_b1 , w_20908 );
not ( \6552_b0 , w_20909 );
and ( w_20908 , w_20909 , \6551_b0 );
buf ( \6553_b1 , \6552_b1 );
not ( \6553_b1 , w_20910 );
not ( \6553_b0 , w_20911 );
and ( w_20910 , w_20911 , \6552_b0 );
buf ( \6554_b1 , \6330_b1 );
not ( \6554_b1 , w_20912 );
not ( \6554_b0 , w_20913 );
and ( w_20912 , w_20913 , \6330_b0 );
or ( \6555_b1 , \6553_b1 , w_20914 );
or ( \6555_b0 , \6553_b0 , \6554_b0 );
not ( \6554_b0 , w_20915 );
and ( w_20915 , w_20914 , \6554_b1 );
or ( \6556_b1 , \6329_b1 , w_20917 );
not ( w_20917 , w_20918 );
and ( \6556_b0 , \6329_b0 , w_20919 );
and ( w_20918 ,  , w_20919 );
buf ( w_20917 , \6551_b1 );
not ( w_20917 , w_20920 );
not (  , w_20921 );
and ( w_20920 , w_20921 , \6551_b0 );
or ( \6557_b1 , \6555_b1 , w_20923 );
not ( w_20923 , w_20924 );
and ( \6557_b0 , \6555_b0 , w_20925 );
and ( w_20924 ,  , w_20925 );
buf ( w_20923 , \6556_b1 );
not ( w_20923 , w_20926 );
not (  , w_20927 );
and ( w_20926 , w_20927 , \6556_b0 );
buf ( \6558_b1 , \6389_b1 );
not ( \6558_b1 , w_20928 );
not ( \6558_b0 , w_20929 );
and ( w_20928 , w_20929 , \6389_b0 );
buf ( \6559_b1 , \6438_b1 );
not ( \6559_b1 , w_20930 );
not ( \6559_b0 , w_20931 );
and ( w_20930 , w_20931 , \6438_b0 );
or ( \6560_b1 , \6558_b1 , w_20932 );
or ( \6560_b0 , \6558_b0 , \6559_b0 );
not ( \6559_b0 , w_20933 );
and ( w_20933 , w_20932 , \6559_b1 );
or ( \6561_b1 , \6438_b1 , w_20934 );
or ( \6561_b0 , \6438_b0 , \6389_b0 );
not ( \6389_b0 , w_20935 );
and ( w_20935 , w_20934 , \6389_b1 );
or ( \6562_b1 , \6561_b1 , w_20937 );
not ( w_20937 , w_20938 );
and ( \6562_b0 , \6561_b0 , w_20939 );
and ( w_20938 ,  , w_20939 );
buf ( w_20937 , \6435_b1 );
not ( w_20937 , w_20940 );
not (  , w_20941 );
and ( w_20940 , w_20941 , \6435_b0 );
or ( \6563_b1 , \6560_b1 , w_20943 );
not ( w_20943 , w_20944 );
and ( \6563_b0 , \6560_b0 , w_20945 );
and ( w_20944 ,  , w_20945 );
buf ( w_20943 , \6562_b1 );
not ( w_20943 , w_20946 );
not (  , w_20947 );
and ( w_20946 , w_20947 , \6562_b0 );
or ( \6564_b1 , \6557_b1 , w_20949 );
not ( w_20949 , w_20950 );
and ( \6564_b0 , \6557_b0 , w_20951 );
and ( w_20950 ,  , w_20951 );
buf ( w_20949 , \6563_b1 );
not ( w_20949 , w_20952 );
not (  , w_20953 );
and ( w_20952 , w_20953 , \6563_b0 );
or ( \6565_b1 , \6546_b1 , w_20954 );
or ( \6565_b0 , \6546_b0 , \6564_b0 );
not ( \6564_b0 , w_20955 );
and ( w_20955 , w_20954 , \6564_b1 );
or ( \6566_b1 , \6557_b1 , w_20957 );
not ( w_20957 , w_20958 );
and ( \6566_b0 , \6557_b0 , w_20959 );
and ( w_20958 ,  , w_20959 );
buf ( w_20957 , \6563_b1 );
not ( w_20957 , w_20960 );
not (  , w_20961 );
and ( w_20960 , w_20961 , \6563_b0 );
or ( \6567_b1 , \6565_b1 , w_20963 );
not ( w_20963 , w_20964 );
and ( \6567_b0 , \6565_b0 , w_20965 );
and ( w_20964 ,  , w_20965 );
buf ( w_20963 , \6566_b1 );
not ( w_20963 , w_20966 );
not (  , w_20967 );
and ( w_20966 , w_20967 , \6566_b0 );
or ( \6568_b1 , \6387_b1 , \6567_b1 );
not ( \6567_b1 , w_20968 );
and ( \6568_b0 , \6387_b0 , w_20969 );
and ( w_20968 , w_20969 , \6567_b0 );
or ( \6569_b1 , \6327_b1 , w_20971 );
not ( w_20971 , w_20972 );
and ( \6569_b0 , \6327_b0 , w_20973 );
and ( w_20972 ,  , w_20973 );
buf ( w_20971 , \6386_b1 );
not ( w_20971 , w_20974 );
not (  , w_20975 );
and ( w_20974 , w_20975 , \6386_b0 );
or ( \6570_b1 , \6568_b1 , w_20977 );
not ( w_20977 , w_20978 );
and ( \6570_b0 , \6568_b0 , w_20979 );
and ( w_20978 ,  , w_20979 );
buf ( w_20977 , \6569_b1 );
not ( w_20977 , w_20980 );
not (  , w_20981 );
and ( w_20980 , w_20981 , \6569_b0 );
buf ( \6571_b1 , \6564_b1 );
buf ( \6571_b0 , \6564_b0 );
or ( \6572_b1 , \6497_b1 , w_20982 );
or ( \6572_b0 , \6497_b0 , \6541_b0 );
not ( \6541_b0 , w_20983 );
and ( w_20983 , w_20982 , \6541_b1 );
or ( \6573_b1 , \6545_b1 , w_20985 );
not ( w_20985 , w_20986 );
and ( \6573_b0 , \6545_b0 , w_20987 );
and ( w_20986 ,  , w_20987 );
buf ( w_20985 , \6572_b1 );
not ( w_20985 , w_20988 );
not (  , w_20989 );
and ( w_20988 , w_20989 , \6572_b0 );
or ( \6574_b1 , \6571_b1 , w_20991 );
not ( w_20991 , w_20992 );
and ( \6574_b0 , \6571_b0 , w_20993 );
and ( w_20992 ,  , w_20993 );
buf ( w_20991 , \6573_b1 );
not ( w_20991 , w_20994 );
not (  , w_20995 );
and ( w_20994 , w_20995 , \6573_b0 );
or ( \6575_b1 , \6525_b1 , \6524_b1 );
xor ( \6575_b0 , \6525_b0 , w_20996 );
not ( w_20996 , w_20997 );
and ( w_20997 , \6524_b1 , \6524_b0 );
or ( \6576_b1 , \6575_b1 , w_20998 );
xor ( \6576_b0 , \6575_b0 , w_21000 );
not ( w_21000 , w_21001 );
and ( w_21001 , w_20998 , w_20999 );
buf ( w_20998 , \6537_b1 );
not ( w_20998 , w_21002 );
not ( w_20999 , w_21003 );
and ( w_21002 , w_21003 , \6537_b0 );
or ( \6577_b1 , \6498_b1 , \6509_b1 );
xor ( \6577_b0 , \6498_b0 , w_21004 );
not ( w_21004 , w_21005 );
and ( w_21005 , \6509_b1 , \6509_b0 );
or ( \6578_b1 , \6577_b1 , \6521_b1 );
xor ( \6578_b0 , \6577_b0 , w_21006 );
not ( w_21006 , w_21007 );
and ( w_21007 , \6521_b1 , \6521_b0 );
buf ( \6579_b1 , \4029_b1 );
not ( \6579_b1 , w_21008 );
not ( \6579_b0 , w_21009 );
and ( w_21008 , w_21009 , \4029_b0 );
buf ( \6580_b1 , \4069_b1 );
not ( \6580_b1 , w_21010 );
not ( \6580_b0 , w_21011 );
and ( w_21010 , w_21011 , \4069_b0 );
or ( \6581_b1 , \6579_b1 , w_21012 );
or ( \6581_b0 , \6579_b0 , \6580_b0 );
not ( \6580_b0 , w_21013 );
and ( w_21013 , w_21012 , \6580_b1 );
or ( \6582_b1 , \4407_b1 , w_21015 );
not ( w_21015 , w_21016 );
and ( \6582_b0 , \4407_b0 , w_21017 );
and ( w_21016 ,  , w_21017 );
buf ( w_21015 , \5339_b1 );
not ( w_21015 , w_21018 );
not (  , w_21019 );
and ( w_21018 , w_21019 , \5339_b0 );
or ( \6583_b1 , \6581_b1 , w_21021 );
not ( w_21021 , w_21022 );
and ( \6583_b0 , \6581_b0 , w_21023 );
and ( w_21022 ,  , w_21023 );
buf ( w_21021 , \6582_b1 );
not ( w_21021 , w_21024 );
not (  , w_21025 );
and ( w_21024 , w_21025 , \6582_b0 );
buf ( \6584_b1 , \6583_b1 );
not ( \6584_b1 , w_21026 );
not ( \6584_b0 , w_21027 );
and ( w_21026 , w_21027 , \6583_b0 );
buf ( \6585_b1 , \6162_b1 );
not ( \6585_b1 , w_21028 );
not ( \6585_b0 , w_21029 );
and ( w_21028 , w_21029 , \6162_b0 );
or ( \6586_b1 , \6584_b1 , w_21030 );
or ( \6586_b0 , \6584_b0 , \6585_b0 );
not ( \6585_b0 , w_21031 );
and ( w_21031 , w_21030 , \6585_b1 );
or ( \6587_b1 , \4055_b1 , w_21033 );
not ( w_21033 , w_21034 );
and ( \6587_b0 , \4055_b0 , w_21035 );
and ( w_21034 ,  , w_21035 );
buf ( w_21033 , \6466_b1 );
not ( w_21033 , w_21036 );
not (  , w_21037 );
and ( w_21036 , w_21037 , \6466_b0 );
or ( \6588_b1 , \6586_b1 , w_21039 );
not ( w_21039 , w_21040 );
and ( \6588_b0 , \6586_b0 , w_21041 );
and ( w_21040 ,  , w_21041 );
buf ( w_21039 , \6587_b1 );
not ( w_21039 , w_21042 );
not (  , w_21043 );
and ( w_21042 , w_21043 , \6587_b0 );
buf ( \6589_b1 , \6588_b1 );
not ( \6589_b1 , w_21044 );
not ( \6589_b0 , w_21045 );
and ( w_21044 , w_21045 , \6588_b0 );
buf ( \6590_b1 , \5388_b1 );
not ( \6590_b1 , w_21046 );
not ( \6590_b0 , w_21047 );
and ( w_21046 , w_21047 , \5388_b0 );
buf ( \6591_b1 , \4049_b1 );
not ( \6591_b1 , w_21048 );
not ( \6591_b0 , w_21049 );
and ( w_21048 , w_21049 , \4049_b0 );
or ( \6592_b1 , \6590_b1 , w_21050 );
or ( \6592_b0 , \6590_b0 , \6591_b0 );
not ( \6591_b0 , w_21051 );
and ( w_21051 , w_21050 , \6591_b1 );
or ( \6593_b1 , \6592_b1 , w_21053 );
not ( w_21053 , w_21054 );
and ( \6593_b0 , \6592_b0 , w_21055 );
and ( w_21054 ,  , w_21055 );
buf ( w_21053 , \4665_b1 );
not ( w_21053 , w_21056 );
not (  , w_21057 );
and ( w_21056 , w_21057 , \4665_b0 );
or ( \6594_b1 , \1454_b1 , w_21059 );
not ( w_21059 , w_21060 );
and ( \6594_b0 , \1454_b0 , w_21061 );
and ( w_21060 ,  , w_21061 );
buf ( w_21059 , \4048_b1 );
not ( w_21059 , w_21062 );
not (  , w_21063 );
and ( w_21062 , w_21063 , \4048_b0 );
buf ( \6596_b1 , \6595_b1 );
not ( \6596_b1 , w_21064 );
not ( \6596_b0 , w_21065 );
and ( w_21064 , w_21065 , \6595_b0 );
buf ( \6597_b1 , \5019_b1 );
not ( \6597_b1 , w_21066 );
not ( \6597_b0 , w_21067 );
and ( w_21066 , w_21067 , \5019_b0 );
buf ( \6598_b1 , \4019_b1 );
not ( \6598_b1 , w_21068 );
not ( \6598_b0 , w_21069 );
and ( w_21068 , w_21069 , \4019_b0 );
buf ( \6599_b1 , \5023_b1 );
not ( \6599_b1 , w_21070 );
not ( \6599_b0 , w_21071 );
and ( w_21070 , w_21071 , \5023_b0 );
or ( \6600_b1 , \6598_b1 , w_21072 );
or ( \6600_b0 , \6598_b0 , \6599_b0 );
not ( \6599_b0 , w_21073 );
and ( w_21073 , w_21072 , \6599_b1 );
or ( \6601_b1 , \6502_b1 , w_21075 );
not ( w_21075 , w_21076 );
and ( \6601_b0 , \6502_b0 , w_21077 );
and ( w_21076 ,  , w_21077 );
buf ( w_21075 , \4585_b1 );
not ( w_21075 , w_21078 );
not (  , w_21079 );
and ( w_21078 , w_21079 , \4585_b0 );
or ( \6602_b1 , \6600_b1 , w_21081 );
not ( w_21081 , w_21082 );
and ( \6602_b0 , \6600_b0 , w_21083 );
and ( w_21082 ,  , w_21083 );
buf ( w_21081 , \6601_b1 );
not ( w_21081 , w_21084 );
not (  , w_21085 );
and ( w_21084 , w_21085 , \6601_b0 );
buf ( \6603_b1 , \6602_b1 );
not ( \6603_b1 , w_21086 );
not ( \6603_b0 , w_21087 );
and ( w_21086 , w_21087 , \6602_b0 );
or ( \6604_b1 , \6597_b1 , w_21088 );
or ( \6604_b0 , \6597_b0 , \6603_b0 );
not ( \6603_b0 , w_21089 );
and ( w_21089 , w_21088 , \6603_b1 );
or ( \6605_b1 , \6504_b1 , w_21091 );
not ( w_21091 , w_21092 );
and ( \6605_b0 , \6504_b0 , w_21093 );
and ( w_21092 ,  , w_21093 );
buf ( w_21091 , \5021_b1 );
not ( w_21091 , w_21094 );
not (  , w_21095 );
and ( w_21094 , w_21095 , \5021_b0 );
or ( \6606_b1 , \6604_b1 , w_21097 );
not ( w_21097 , w_21098 );
and ( \6606_b0 , \6604_b0 , w_21099 );
and ( w_21098 ,  , w_21099 );
buf ( w_21097 , \6605_b1 );
not ( w_21097 , w_21100 );
not (  , w_21101 );
and ( w_21100 , w_21101 , \6605_b0 );
or ( \6607_b1 , \6596_b1 , w_21103 );
not ( w_21103 , w_21104 );
and ( \6607_b0 , \6596_b0 , w_21105 );
and ( w_21104 ,  , w_21105 );
buf ( w_21103 , \6606_b1 );
not ( w_21103 , w_21106 );
not (  , w_21107 );
and ( w_21106 , w_21107 , \6606_b0 );
or ( \6608_b1 , \6589_b1 , w_21109 );
not ( w_21109 , w_21110 );
and ( \6608_b0 , \6589_b0 , w_21111 );
and ( w_21110 ,  , w_21111 );
buf ( w_21109 , \6607_b1 );
not ( w_21109 , w_21112 );
not (  , w_21113 );
and ( w_21112 , w_21113 , \6607_b0 );
or ( \6609_b1 , \6578_b1 , \6608_b1 );
not ( \6608_b1 , w_21114 );
and ( \6609_b0 , \6578_b0 , w_21115 );
and ( w_21114 , w_21115 , \6608_b0 );
buf ( \6610_b1 , \6588_b1 );
not ( \6610_b1 , w_21116 );
not ( \6610_b0 , w_21117 );
and ( w_21116 , w_21117 , \6588_b0 );
or ( \6611_b1 , \6610_b1 , w_21119 );
not ( w_21119 , w_21120 );
and ( \6611_b0 , \6610_b0 , w_21121 );
and ( w_21120 ,  , w_21121 );
buf ( w_21119 , \6607_b1 );
not ( w_21119 , w_21122 );
not (  , w_21123 );
and ( w_21122 , w_21123 , \6607_b0 );
or ( \6612_b1 , \6609_b1 , w_21125 );
not ( w_21125 , w_21126 );
and ( \6612_b0 , \6609_b0 , w_21127 );
and ( w_21126 ,  , w_21127 );
buf ( w_21125 , \6611_b1 );
not ( w_21125 , w_21128 );
not (  , w_21129 );
and ( w_21128 , w_21129 , \6611_b0 );
or ( \6613_b1 , \6576_b1 , w_21131 );
not ( w_21131 , w_21132 );
and ( \6613_b0 , \6576_b0 , w_21133 );
and ( w_21132 ,  , w_21133 );
buf ( w_21131 , \6612_b1 );
not ( w_21131 , w_21134 );
not (  , w_21135 );
and ( w_21134 , w_21135 , \6612_b0 );
buf ( \6614_b1 , \6613_b1 );
not ( \6614_b1 , w_21136 );
not ( \6614_b0 , w_21137 );
and ( w_21136 , w_21137 , \6613_b0 );
buf ( \6615_b1 , \6588_b1 );
not ( \6615_b1 , w_21138 );
not ( \6615_b0 , w_21139 );
and ( w_21138 , w_21139 , \6588_b0 );
buf ( \6616_b1 , \6607_b1 );
not ( \6616_b1 , w_21140 );
not ( \6616_b0 , w_21141 );
and ( w_21140 , w_21141 , \6607_b0 );
or ( \6617_b1 , \6615_b1 , \6616_b1 );
not ( \6616_b1 , w_21142 );
and ( \6617_b0 , \6615_b0 , w_21143 );
and ( w_21142 , w_21143 , \6616_b0 );
or ( \6618_b1 , \6588_b1 , \6607_b1 );
not ( \6607_b1 , w_21144 );
and ( \6618_b0 , \6588_b0 , w_21145 );
and ( w_21144 , w_21145 , \6607_b0 );
or ( \6619_b1 , \6617_b1 , w_21147 );
not ( w_21147 , w_21148 );
and ( \6619_b0 , \6617_b0 , w_21149 );
and ( w_21148 ,  , w_21149 );
buf ( w_21147 , \6618_b1 );
not ( w_21147 , w_21150 );
not (  , w_21151 );
and ( w_21150 , w_21151 , \6618_b0 );
or ( \6620_b1 , \6578_b1 , \6619_b1 );
xor ( \6620_b0 , \6578_b0 , w_21152 );
not ( w_21152 , w_21153 );
and ( w_21153 , \6619_b1 , \6619_b0 );
buf ( \6621_b1 , \6606_b1 );
not ( \6621_b1 , w_21154 );
not ( \6621_b0 , w_21155 );
and ( w_21154 , w_21155 , \6606_b0 );
buf ( \6622_b1 , \6595_b1 );
not ( \6622_b1 , w_21156 );
not ( \6622_b0 , w_21157 );
and ( w_21156 , w_21157 , \6595_b0 );
or ( \6623_b1 , \6621_b1 , \6622_b1 );
not ( \6622_b1 , w_21158 );
and ( \6623_b0 , \6621_b0 , w_21159 );
and ( w_21158 , w_21159 , \6622_b0 );
or ( \6624_b1 , \6606_b1 , \6595_b1 );
not ( \6595_b1 , w_21160 );
and ( \6624_b0 , \6606_b0 , w_21161 );
and ( w_21160 , w_21161 , \6595_b0 );
or ( \6625_b1 , \6623_b1 , w_21163 );
not ( w_21163 , w_21164 );
and ( \6625_b0 , \6623_b0 , w_21165 );
and ( w_21164 ,  , w_21165 );
buf ( w_21163 , \6624_b1 );
not ( w_21163 , w_21166 );
not (  , w_21167 );
and ( w_21166 , w_21167 , \6624_b0 );
or ( \6626_b1 , \5178_b1 , \4026_b1 );
not ( \4026_b1 , w_21168 );
and ( \6626_b0 , \5178_b0 , w_21169 );
and ( w_21168 , w_21169 , \4026_b0 );
buf ( \6627_b1 , \5178_b1 );
not ( \6627_b1 , w_21170 );
not ( \6627_b0 , w_21171 );
and ( w_21170 , w_21171 , \5178_b0 );
or ( \6628_b1 , \6627_b1 , \5344_b1 );
not ( \5344_b1 , w_21172 );
and ( \6628_b0 , \6627_b0 , w_21173 );
and ( w_21172 , w_21173 , \5344_b0 );
or ( \6629_b1 , \6626_b1 , w_21174 );
or ( \6629_b0 , \6626_b0 , \6628_b0 );
not ( \6628_b0 , w_21175 );
and ( w_21175 , w_21174 , \6628_b1 );
buf ( \6630_b1 , \6629_b1 );
not ( \6630_b1 , w_21176 );
not ( \6630_b0 , w_21177 );
and ( w_21176 , w_21177 , \6629_b0 );
buf ( \6631_b1 , \4662_b1 );
not ( \6631_b1 , w_21178 );
not ( \6631_b0 , w_21179 );
and ( w_21178 , w_21179 , \4662_b0 );
or ( \6632_b1 , \6630_b1 , w_21180 );
or ( \6632_b0 , \6630_b0 , \6631_b0 );
not ( \6631_b0 , w_21181 );
and ( w_21181 , w_21180 , \6631_b1 );
or ( \6633_b1 , \4672_b1 , w_21183 );
not ( w_21183 , w_21184 );
and ( \6633_b0 , \4672_b0 , w_21185 );
and ( w_21184 ,  , w_21185 );
buf ( w_21183 , \6517_b1 );
not ( w_21183 , w_21186 );
not (  , w_21187 );
and ( w_21186 , w_21187 , \6517_b0 );
or ( \6634_b1 , \6632_b1 , w_21189 );
not ( w_21189 , w_21190 );
and ( \6634_b0 , \6632_b0 , w_21191 );
and ( w_21190 ,  , w_21191 );
buf ( w_21189 , \6633_b1 );
not ( w_21189 , w_21192 );
not (  , w_21193 );
and ( w_21192 , w_21193 , \6633_b0 );
buf ( \6635_b1 , \6634_b1 );
not ( \6635_b1 , w_21194 );
not ( \6635_b0 , w_21195 );
and ( w_21194 , w_21195 , \6634_b0 );
or ( \6636_b1 , \6625_b1 , \6635_b1 );
xor ( \6636_b0 , \6625_b0 , w_21196 );
not ( w_21196 , w_21197 );
and ( w_21197 , \6635_b1 , \6635_b0 );
buf ( \6637_b1 , \4411_b1 );
not ( \6637_b1 , w_21198 );
not ( \6637_b0 , w_21199 );
and ( w_21198 , w_21199 , \4411_b0 );
or ( \6638_b1 , \5388_b1 , \4070_b1 );
not ( \4070_b1 , w_21200 );
and ( \6638_b0 , \5388_b0 , w_21201 );
and ( w_21200 , w_21201 , \4070_b0 );
buf ( \6639_b1 , \5388_b1 );
not ( \6639_b1 , w_21202 );
not ( \6639_b0 , w_21203 );
and ( w_21202 , w_21203 , \5388_b0 );
or ( \6640_b1 , \6639_b1 , \4399_b1 );
not ( \4399_b1 , w_21204 );
and ( \6640_b0 , \6639_b0 , w_21205 );
and ( w_21204 , w_21205 , \4399_b0 );
or ( \6641_b1 , \6638_b1 , w_21207 );
not ( w_21207 , w_21208 );
and ( \6641_b0 , \6638_b0 , w_21209 );
and ( w_21208 ,  , w_21209 );
buf ( w_21207 , \6640_b1 );
not ( w_21207 , w_21210 );
not (  , w_21211 );
and ( w_21210 , w_21211 , \6640_b0 );
buf ( \6642_b1 , \6641_b1 );
not ( \6642_b1 , w_21212 );
not ( \6642_b0 , w_21213 );
and ( w_21212 , w_21213 , \6641_b0 );
or ( \6643_b1 , \6637_b1 , \6642_b1 );
not ( \6642_b1 , w_21214 );
and ( \6643_b0 , \6637_b0 , w_21215 );
and ( w_21214 , w_21215 , \6642_b0 );
buf ( \6644_b1 , \6583_b1 );
not ( \6644_b1 , w_21216 );
not ( \6644_b0 , w_21217 );
and ( w_21216 , w_21217 , \6583_b0 );
or ( \6645_b1 , \6644_b1 , w_21219 );
not ( w_21219 , w_21220 );
and ( \6645_b0 , \6644_b0 , w_21221 );
and ( w_21220 ,  , w_21221 );
buf ( w_21219 , \4056_b1 );
not ( w_21219 , w_21222 );
not (  , w_21223 );
and ( w_21222 , w_21223 , \4056_b0 );
or ( \6646_b1 , \6643_b1 , w_21225 );
not ( w_21225 , w_21226 );
and ( \6646_b0 , \6643_b0 , w_21227 );
and ( w_21226 ,  , w_21227 );
buf ( w_21225 , \6645_b1 );
not ( w_21225 , w_21228 );
not (  , w_21229 );
and ( w_21228 , w_21229 , \6645_b0 );
or ( \6647_b1 , \6636_b1 , \6646_b1 );
not ( \6646_b1 , w_21230 );
and ( \6647_b0 , \6636_b0 , w_21231 );
and ( w_21230 , w_21231 , \6646_b0 );
or ( \6648_b1 , \6625_b1 , \6635_b1 );
not ( \6635_b1 , w_21232 );
and ( \6648_b0 , \6625_b0 , w_21233 );
and ( w_21232 , w_21233 , \6635_b0 );
or ( \6649_b1 , \6647_b1 , w_21234 );
or ( \6649_b0 , \6647_b0 , \6648_b0 );
not ( \6648_b0 , w_21235 );
and ( w_21235 , w_21234 , \6648_b1 );
or ( \6650_b1 , \6620_b1 , w_21237 );
not ( w_21237 , w_21238 );
and ( \6650_b0 , \6620_b0 , w_21239 );
and ( w_21238 ,  , w_21239 );
buf ( w_21237 , \6649_b1 );
not ( w_21237 , w_21240 );
not (  , w_21241 );
and ( w_21240 , w_21241 , \6649_b0 );
buf ( \6651_b1 , \4026_b1 );
not ( \6651_b1 , w_21242 );
not ( \6651_b0 , w_21243 );
and ( w_21242 , w_21243 , \4026_b0 );
buf ( \6652_b1 , \5874_b1 );
not ( \6652_b1 , w_21244 );
not ( \6652_b0 , w_21245 );
and ( w_21244 , w_21245 , \5874_b0 );
or ( \6653_b1 , \6651_b1 , w_21246 );
or ( \6653_b0 , \6651_b0 , \6652_b0 );
not ( \6652_b0 , w_21247 );
and ( w_21247 , w_21246 , \6652_b1 );
or ( \6654_b1 , \5024_b1 , w_21249 );
not ( w_21249 , w_21250 );
and ( \6654_b0 , \5024_b0 , w_21251 );
and ( w_21250 ,  , w_21251 );
buf ( w_21249 , \5344_b1 );
not ( w_21249 , w_21252 );
not (  , w_21253 );
and ( w_21252 , w_21253 , \5344_b0 );
or ( \6655_b1 , \6653_b1 , w_21255 );
not ( w_21255 , w_21256 );
and ( \6655_b0 , \6653_b0 , w_21257 );
and ( w_21256 ,  , w_21257 );
buf ( w_21255 , \6654_b1 );
not ( w_21255 , w_21258 );
not (  , w_21259 );
and ( w_21258 , w_21259 , \6654_b0 );
buf ( \6656_b1 , \6655_b1 );
not ( \6656_b1 , w_21260 );
not ( \6656_b0 , w_21261 );
and ( w_21260 , w_21261 , \6655_b0 );
buf ( \6657_b1 , \5020_b1 );
not ( \6657_b1 , w_21262 );
not ( \6657_b0 , w_21263 );
and ( w_21262 , w_21263 , \5020_b0 );
or ( \6658_b1 , \6656_b1 , w_21264 );
or ( \6658_b0 , \6656_b0 , \6657_b0 );
not ( \6657_b0 , w_21265 );
and ( w_21265 , w_21264 , \6657_b1 );
buf ( \6659_b1 , \4023_b1 );
not ( \6659_b1 , w_21266 );
not ( \6659_b0 , w_21267 );
and ( w_21266 , w_21267 , \4023_b0 );
buf ( \6660_b1 , \5874_b1 );
not ( \6660_b1 , w_21268 );
not ( \6660_b0 , w_21269 );
and ( w_21268 , w_21269 , \5874_b0 );
or ( \6661_b1 , \6659_b1 , w_21270 );
or ( \6661_b0 , \6659_b0 , \6660_b0 );
not ( \6660_b0 , w_21271 );
and ( w_21271 , w_21270 , \6660_b1 );
or ( \6662_b1 , \5873_b1 , w_21273 );
not ( w_21273 , w_21274 );
and ( \6662_b0 , \5873_b0 , w_21275 );
and ( w_21274 ,  , w_21275 );
buf ( w_21273 , \5131_b1 );
not ( w_21273 , w_21276 );
not (  , w_21277 );
and ( w_21276 , w_21277 , \5131_b0 );
or ( \6663_b1 , \6661_b1 , w_21279 );
not ( w_21279 , w_21280 );
and ( \6663_b0 , \6661_b0 , w_21281 );
and ( w_21280 ,  , w_21281 );
buf ( w_21279 , \6662_b1 );
not ( w_21279 , w_21282 );
not (  , w_21283 );
and ( w_21282 , w_21283 , \6662_b0 );
or ( \6664_b1 , \6663_b1 , w_21285 );
not ( w_21285 , w_21286 );
and ( \6664_b0 , \6663_b0 , w_21287 );
and ( w_21286 ,  , w_21287 );
buf ( w_21285 , \5021_b1 );
not ( w_21285 , w_21288 );
not (  , w_21289 );
and ( w_21288 , w_21289 , \5021_b0 );
or ( \6665_b1 , \6658_b1 , w_21291 );
not ( w_21291 , w_21292 );
and ( \6665_b0 , \6658_b0 , w_21293 );
and ( w_21292 ,  , w_21293 );
buf ( w_21291 , \6664_b1 );
not ( w_21291 , w_21294 );
not (  , w_21295 );
and ( w_21294 , w_21295 , \6664_b0 );
buf ( \6666_b1 , \6665_b1 );
not ( \6666_b1 , w_21296 );
not ( \6666_b0 , w_21297 );
and ( w_21296 , w_21297 , \6665_b0 );
buf ( \6667_b1 , \5178_b1 );
not ( \6667_b1 , w_21298 );
not ( \6667_b0 , w_21299 );
and ( w_21298 , w_21299 , \5178_b0 );
buf ( \6668_b1 , \4535_b1 );
not ( \6668_b1 , w_21300 );
not ( \6668_b0 , w_21301 );
and ( w_21300 , w_21301 , \4535_b0 );
or ( \6669_b1 , \6668_b1 , w_21303 );
not ( w_21303 , w_21304 );
and ( \6669_b0 , \6668_b0 , w_21305 );
and ( w_21304 ,  , w_21305 );
buf ( w_21303 , \4048_b1 );
not ( w_21303 , w_21306 );
not (  , w_21307 );
and ( w_21306 , w_21307 , \4048_b0 );
buf ( \6670_b1 , \5388_b1 );
not ( \6670_b1 , w_21308 );
not ( \6670_b0 , w_21309 );
and ( w_21308 , w_21309 , \5388_b0 );
buf ( \6671_b1 , \4535_b1 );
not ( \6671_b1 , w_21310 );
not ( \6671_b0 , w_21311 );
and ( w_21310 , w_21311 , \4535_b0 );
or ( \6672_b1 , \6670_b1 , w_21312 );
or ( \6672_b0 , \6670_b0 , \6671_b0 );
not ( \6671_b0 , w_21313 );
and ( w_21313 , w_21312 , \6671_b1 );
or ( \6673_b1 , \6672_b1 , w_21315 );
not ( w_21315 , w_21316 );
and ( \6673_b0 , \6672_b0 , w_21317 );
and ( w_21316 ,  , w_21317 );
buf ( w_21315 , \5873_b1 );
not ( w_21315 , w_21318 );
not (  , w_21319 );
and ( w_21318 , w_21319 , \5873_b0 );
buf ( \6675_b1 , \6674_b1 );
not ( \6675_b1 , w_21320 );
not ( \6675_b0 , w_21321 );
and ( w_21320 , w_21321 , \6674_b0 );
or ( \6676_b1 , \6666_b1 , \6675_b1 );
not ( \6675_b1 , w_21322 );
and ( \6676_b0 , \6666_b0 , w_21323 );
and ( w_21322 , w_21323 , \6675_b0 );
or ( \6677_b1 , \6665_b1 , \6674_b1 );
not ( \6674_b1 , w_21324 );
and ( \6677_b0 , \6665_b0 , w_21325 );
and ( w_21324 , w_21325 , \6674_b0 );
or ( \6678_b1 , \6676_b1 , w_21327 );
not ( w_21327 , w_21328 );
and ( \6678_b0 , \6676_b0 , w_21329 );
and ( w_21328 ,  , w_21329 );
buf ( w_21327 , \6677_b1 );
not ( w_21327 , w_21330 );
not (  , w_21331 );
and ( w_21330 , w_21331 , \6677_b0 );
buf ( \6679_b1 , \4663_b1 );
not ( \6679_b1 , w_21332 );
not ( \6679_b0 , w_21333 );
and ( w_21332 , w_21333 , \4663_b0 );
or ( \6680_b1 , \5388_b1 , \4665_b1 );
not ( \4665_b1 , w_21334 );
and ( \6680_b0 , \5388_b0 , w_21335 );
and ( w_21334 , w_21335 , \4665_b0 );
buf ( \6681_b1 , \5388_b1 );
not ( \6681_b1 , w_21336 );
not ( \6681_b0 , w_21337 );
and ( w_21336 , w_21337 , \5388_b0 );
or ( \6682_b1 , \6681_b1 , \4666_b1 );
not ( \4666_b1 , w_21338 );
and ( \6682_b0 , \6681_b0 , w_21339 );
and ( w_21338 , w_21339 , \4666_b0 );
or ( \6683_b1 , \6680_b1 , w_21341 );
not ( w_21341 , w_21342 );
and ( \6683_b0 , \6680_b0 , w_21343 );
and ( w_21342 ,  , w_21343 );
buf ( w_21341 , \6682_b1 );
not ( w_21341 , w_21344 );
not (  , w_21345 );
and ( w_21344 , w_21345 , \6682_b0 );
buf ( \6684_b1 , \6683_b1 );
not ( \6684_b1 , w_21346 );
not ( \6684_b0 , w_21347 );
and ( w_21346 , w_21347 , \6683_b0 );
or ( \6685_b1 , \6679_b1 , \6684_b1 );
not ( \6684_b1 , w_21348 );
and ( \6685_b0 , \6679_b0 , w_21349 );
and ( w_21348 , w_21349 , \6684_b0 );
buf ( \6686_b1 , \4029_b1 );
not ( \6686_b1 , w_21350 );
not ( \6686_b0 , w_21351 );
and ( w_21350 , w_21351 , \4029_b0 );
buf ( \6687_b1 , \4666_b1 );
not ( \6687_b1 , w_21352 );
not ( \6687_b0 , w_21353 );
and ( w_21352 , w_21353 , \4666_b0 );
or ( \6688_b1 , \6686_b1 , w_21354 );
or ( \6688_b0 , \6686_b0 , \6687_b0 );
not ( \6687_b0 , w_21355 );
and ( w_21355 , w_21354 , \6687_b1 );
buf ( \6689_b1 , \5178_b1 );
not ( \6689_b1 , w_21356 );
not ( \6689_b0 , w_21357 );
and ( w_21356 , w_21357 , \5178_b0 );
or ( \6690_b1 , \6689_b1 , w_21359 );
not ( w_21359 , w_21360 );
and ( \6690_b0 , \6689_b0 , w_21361 );
and ( w_21360 ,  , w_21361 );
buf ( w_21359 , \5339_b1 );
not ( w_21359 , w_21362 );
not (  , w_21363 );
and ( w_21362 , w_21363 , \5339_b0 );
or ( \6691_b1 , \6688_b1 , w_21365 );
not ( w_21365 , w_21366 );
and ( \6691_b0 , \6688_b0 , w_21367 );
and ( w_21366 ,  , w_21367 );
buf ( w_21365 , \6690_b1 );
not ( w_21365 , w_21368 );
not (  , w_21369 );
and ( w_21368 , w_21369 , \6690_b0 );
or ( \6692_b1 , \5187_b1 , \6691_b1 );
not ( \6691_b1 , w_21370 );
and ( \6692_b0 , \5187_b0 , w_21371 );
and ( w_21370 , w_21371 , \6691_b0 );
or ( \6693_b1 , \6685_b1 , w_21373 );
not ( w_21373 , w_21374 );
and ( \6693_b0 , \6685_b0 , w_21375 );
and ( w_21374 ,  , w_21375 );
buf ( w_21373 , \6692_b1 );
not ( w_21373 , w_21376 );
not (  , w_21377 );
and ( w_21376 , w_21377 , \6692_b0 );
or ( \6694_b1 , \6678_b1 , w_21378 );
or ( \6694_b0 , \6678_b0 , \6693_b0 );
not ( \6693_b0 , w_21379 );
and ( w_21379 , w_21378 , \6693_b1 );
buf ( \6695_b1 , \4048_b1 );
not ( \6695_b1 , w_21380 );
not ( \6695_b0 , w_21381 );
and ( w_21380 , w_21381 , \4048_b0 );
buf ( \6696_b1 , \5874_b1 );
not ( \6696_b1 , w_21382 );
not ( \6696_b0 , w_21383 );
and ( w_21382 , w_21383 , \5874_b0 );
or ( \6697_b1 , \6695_b1 , w_21384 );
or ( \6697_b0 , \6695_b0 , \6696_b0 );
not ( \6696_b0 , w_21385 );
and ( w_21385 , w_21384 , \6696_b1 );
or ( \6698_b1 , \5024_b1 , w_21387 );
not ( w_21387 , w_21388 );
and ( \6698_b0 , \5024_b0 , w_21389 );
and ( w_21388 ,  , w_21389 );
buf ( w_21387 , \5388_b1 );
not ( w_21387 , w_21390 );
not (  , w_21391 );
and ( w_21390 , w_21391 , \5388_b0 );
or ( \6699_b1 , \6697_b1 , w_21393 );
not ( w_21393 , w_21394 );
and ( \6699_b0 , \6697_b0 , w_21395 );
and ( w_21394 ,  , w_21395 );
buf ( w_21393 , \6698_b1 );
not ( w_21393 , w_21396 );
not (  , w_21397 );
and ( w_21396 , w_21397 , \6698_b0 );
or ( \6700_b1 , \5020_b1 , \6699_b1 );
not ( \6699_b1 , w_21398 );
and ( \6700_b0 , \5020_b0 , w_21399 );
and ( w_21398 , w_21399 , \6699_b0 );
buf ( \6701_b1 , \4029_b1 );
not ( \6701_b1 , w_21400 );
not ( \6701_b0 , w_21401 );
and ( w_21400 , w_21401 , \4029_b0 );
buf ( \6702_b1 , \5874_b1 );
not ( \6702_b1 , w_21402 );
not ( \6702_b0 , w_21403 );
and ( w_21402 , w_21403 , \5874_b0 );
or ( \6703_b1 , \6701_b1 , w_21404 );
or ( \6703_b0 , \6701_b0 , \6702_b0 );
not ( \6702_b0 , w_21405 );
and ( w_21405 , w_21404 , \6702_b1 );
or ( \6704_b1 , \5873_b1 , w_21407 );
not ( w_21407 , w_21408 );
and ( \6704_b0 , \5873_b0 , w_21409 );
and ( w_21408 ,  , w_21409 );
buf ( w_21407 , \5339_b1 );
not ( w_21407 , w_21410 );
not (  , w_21411 );
and ( w_21410 , w_21411 , \5339_b0 );
or ( \6705_b1 , \6703_b1 , w_21413 );
not ( w_21413 , w_21414 );
and ( \6705_b0 , \6703_b0 , w_21415 );
and ( w_21414 ,  , w_21415 );
buf ( w_21413 , \6704_b1 );
not ( w_21413 , w_21416 );
not (  , w_21417 );
and ( w_21416 , w_21417 , \6704_b0 );
or ( \6706_b1 , \6705_b1 , \5021_b1 );
not ( \5021_b1 , w_21418 );
and ( \6706_b0 , \6705_b0 , w_21419 );
and ( w_21418 , w_21419 , \5021_b0 );
or ( \6707_b1 , \6700_b1 , w_21421 );
not ( w_21421 , w_21422 );
and ( \6707_b0 , \6700_b0 , w_21423 );
and ( w_21422 ,  , w_21423 );
buf ( w_21421 , \6706_b1 );
not ( w_21421 , w_21424 );
not (  , w_21425 );
and ( w_21424 , w_21425 , \6706_b0 );
or ( \6708_b1 , \5021_b1 , w_21427 );
not ( w_21427 , w_21428 );
and ( \6708_b0 , \5021_b0 , w_21429 );
and ( w_21428 ,  , w_21429 );
buf ( w_21427 , \4048_b1 );
not ( w_21427 , w_21430 );
not (  , w_21431 );
and ( w_21430 , w_21431 , \4048_b0 );
or ( \6709_b1 , \5024_b1 , w_21433 );
not ( w_21433 , w_21434 );
and ( \6709_b0 , \5024_b0 , w_21435 );
and ( w_21434 ,  , w_21435 );
buf ( w_21433 , \6708_b1 );
not ( w_21433 , w_21436 );
not (  , w_21437 );
and ( w_21436 , w_21437 , \6708_b0 );
or ( \6710_b1 , \6707_b1 , w_21439 );
not ( w_21439 , w_21440 );
and ( \6710_b0 , \6707_b0 , w_21441 );
and ( w_21440 ,  , w_21441 );
buf ( w_21439 , \6709_b1 );
not ( w_21439 , w_21442 );
not (  , w_21443 );
and ( w_21442 , w_21443 , \6709_b0 );
buf ( \6711_b1 , \6710_b1 );
not ( \6711_b1 , w_21444 );
not ( \6711_b0 , w_21445 );
and ( w_21444 , w_21445 , \6710_b0 );
buf ( \6712_b1 , \5020_b1 );
not ( \6712_b1 , w_21446 );
not ( \6712_b0 , w_21447 );
and ( w_21446 , w_21447 , \5020_b0 );
buf ( \6713_b1 , \6705_b1 );
not ( \6713_b1 , w_21448 );
not ( \6713_b0 , w_21449 );
and ( w_21448 , w_21449 , \6705_b0 );
or ( \6714_b1 , \6712_b1 , w_21450 );
or ( \6714_b0 , \6712_b0 , \6713_b0 );
not ( \6713_b0 , w_21451 );
and ( w_21451 , w_21450 , \6713_b1 );
or ( \6715_b1 , \6655_b1 , w_21453 );
not ( w_21453 , w_21454 );
and ( \6715_b0 , \6655_b0 , w_21455 );
and ( w_21454 ,  , w_21455 );
buf ( w_21453 , \5021_b1 );
not ( w_21453 , w_21456 );
not (  , w_21457 );
and ( w_21456 , w_21457 , \5021_b0 );
or ( \6716_b1 , \6714_b1 , w_21459 );
not ( w_21459 , w_21460 );
and ( \6716_b0 , \6714_b0 , w_21461 );
and ( w_21460 ,  , w_21461 );
buf ( w_21459 , \6715_b1 );
not ( w_21459 , w_21462 );
not (  , w_21463 );
and ( w_21462 , w_21463 , \6715_b0 );
buf ( \6717_b1 , \6716_b1 );
not ( \6717_b1 , w_21464 );
not ( \6717_b0 , w_21465 );
and ( w_21464 , w_21465 , \6716_b0 );
or ( \6718_b1 , \5187_b1 , w_21467 );
not ( w_21467 , w_21468 );
and ( \6718_b0 , \5187_b0 , w_21469 );
and ( w_21468 ,  , w_21469 );
buf ( w_21467 , \4048_b1 );
not ( w_21467 , w_21470 );
not (  , w_21471 );
and ( w_21470 , w_21471 , \4048_b0 );
or ( \6719_b1 , \6717_b1 , w_21473 );
not ( w_21473 , w_21474 );
and ( \6719_b0 , \6717_b0 , w_21475 );
and ( w_21474 ,  , w_21475 );
buf ( w_21473 , \6718_b1 );
not ( w_21473 , w_21476 );
not (  , w_21477 );
and ( w_21476 , w_21477 , \6718_b0 );
buf ( \6720_b1 , \6719_b1 );
not ( \6720_b1 , w_21478 );
not ( \6720_b0 , w_21479 );
and ( w_21478 , w_21479 , \6719_b0 );
or ( \6721_b1 , \6711_b1 , w_21480 );
or ( \6721_b0 , \6711_b0 , \6720_b0 );
not ( \6720_b0 , w_21481 );
and ( w_21481 , w_21480 , \6720_b1 );
buf ( \6722_b1 , \6718_b1 );
not ( \6722_b1 , w_21482 );
not ( \6722_b0 , w_21483 );
and ( w_21482 , w_21483 , \6718_b0 );
or ( \6723_b1 , \6722_b1 , w_21485 );
not ( w_21485 , w_21486 );
and ( \6723_b0 , \6722_b0 , w_21487 );
and ( w_21486 ,  , w_21487 );
buf ( w_21485 , \6716_b1 );
not ( w_21485 , w_21488 );
not (  , w_21489 );
and ( w_21488 , w_21489 , \6716_b0 );
or ( \6724_b1 , \6721_b1 , w_21491 );
not ( w_21491 , w_21492 );
and ( \6724_b0 , \6721_b0 , w_21493 );
and ( w_21492 ,  , w_21493 );
buf ( w_21491 , \6723_b1 );
not ( w_21491 , w_21494 );
not (  , w_21495 );
and ( w_21494 , w_21495 , \6723_b0 );
or ( \6725_b1 , \6678_b1 , w_21497 );
not ( w_21497 , w_21498 );
and ( \6725_b0 , \6678_b0 , w_21499 );
and ( w_21498 ,  , w_21499 );
buf ( w_21497 , \6693_b1 );
not ( w_21497 , w_21500 );
not (  , w_21501 );
and ( w_21500 , w_21501 , \6693_b0 );
or ( \6726_b1 , \6724_b1 , w_21503 );
not ( w_21503 , w_21504 );
and ( \6726_b0 , \6724_b0 , w_21505 );
and ( w_21504 ,  , w_21505 );
buf ( w_21503 , \6725_b1 );
not ( w_21503 , w_21506 );
not (  , w_21507 );
and ( w_21506 , w_21507 , \6725_b0 );
or ( \6727_b1 , \6694_b1 , w_21509 );
not ( w_21509 , w_21510 );
and ( \6727_b0 , \6694_b0 , w_21511 );
and ( w_21510 ,  , w_21511 );
buf ( w_21509 , \6726_b1 );
not ( w_21509 , w_21512 );
not (  , w_21513 );
and ( w_21512 , w_21513 , \6726_b0 );
buf ( \6728_b1 , \6727_b1 );
not ( \6728_b1 , w_21514 );
not ( \6728_b0 , w_21515 );
and ( w_21514 , w_21515 , \6727_b0 );
or ( \6729_b1 , \4055_b1 , w_21517 );
not ( w_21517 , w_21518 );
and ( \6729_b0 , \4055_b0 , w_21519 );
and ( w_21518 ,  , w_21519 );
buf ( w_21517 , \4048_b1 );
not ( w_21517 , w_21520 );
not (  , w_21521 );
and ( w_21520 , w_21521 , \4048_b0 );
buf ( \6730_b1 , \6602_b1 );
not ( \6730_b1 , w_21522 );
not ( \6730_b0 , w_21523 );
and ( w_21522 , w_21523 , \6602_b0 );
buf ( \6731_b1 , \6730_b1 );
not ( \6731_b1 , w_21524 );
not ( \6731_b0 , w_21525 );
and ( w_21524 , w_21525 , \6730_b0 );
buf ( \6732_b1 , \5265_b1 );
not ( \6732_b1 , w_21526 );
not ( \6732_b0 , w_21527 );
and ( w_21526 , w_21527 , \5265_b0 );
or ( \6733_b1 , \6731_b1 , \6732_b1 );
not ( \6732_b1 , w_21528 );
and ( \6733_b0 , \6731_b0 , w_21529 );
and ( w_21528 , w_21529 , \6732_b0 );
or ( \6734_b1 , \6663_b1 , \5020_b1 );
not ( \5020_b1 , w_21530 );
and ( \6734_b0 , \6663_b0 , w_21531 );
and ( w_21530 , w_21531 , \5020_b0 );
or ( \6735_b1 , \6733_b1 , w_21533 );
not ( w_21533 , w_21534 );
and ( \6735_b0 , \6733_b0 , w_21535 );
and ( w_21534 ,  , w_21535 );
buf ( w_21533 , \6734_b1 );
not ( w_21533 , w_21536 );
not (  , w_21537 );
and ( w_21536 , w_21537 , \6734_b0 );
or ( \6736_b1 , \6729_b1 , \6735_b1 );
xor ( \6736_b0 , \6729_b0 , w_21538 );
not ( w_21538 , w_21539 );
and ( w_21539 , \6735_b1 , \6735_b0 );
buf ( \6737_b1 , \6691_b1 );
not ( \6737_b1 , w_21540 );
not ( \6737_b0 , w_21541 );
and ( w_21540 , w_21541 , \6691_b0 );
buf ( \6738_b1 , \4662_b1 );
not ( \6738_b1 , w_21542 );
not ( \6738_b0 , w_21543 );
and ( w_21542 , w_21543 , \4662_b0 );
or ( \6739_b1 , \6737_b1 , w_21544 );
or ( \6739_b0 , \6737_b0 , \6738_b0 );
not ( \6738_b0 , w_21545 );
and ( w_21545 , w_21544 , \6738_b1 );
or ( \6740_b1 , \5187_b1 , w_21547 );
not ( w_21547 , w_21548 );
and ( \6740_b0 , \5187_b0 , w_21549 );
and ( w_21548 ,  , w_21549 );
buf ( w_21547 , \6629_b1 );
not ( w_21547 , w_21550 );
not (  , w_21551 );
and ( w_21550 , w_21551 , \6629_b0 );
or ( \6741_b1 , \6739_b1 , w_21553 );
not ( w_21553 , w_21554 );
and ( \6741_b0 , \6739_b0 , w_21555 );
and ( w_21554 ,  , w_21555 );
buf ( w_21553 , \6740_b1 );
not ( w_21553 , w_21556 );
not (  , w_21557 );
and ( w_21556 , w_21557 , \6740_b0 );
or ( \6742_b1 , \6736_b1 , w_21558 );
xor ( \6742_b0 , \6736_b0 , w_21560 );
not ( w_21560 , w_21561 );
and ( w_21561 , w_21558 , w_21559 );
buf ( w_21558 , \6741_b1 );
not ( w_21558 , w_21562 );
not ( w_21559 , w_21563 );
and ( w_21562 , w_21563 , \6741_b0 );
buf ( \6743_b1 , \6674_b1 );
not ( \6743_b1 , w_21564 );
not ( \6743_b0 , w_21565 );
and ( w_21564 , w_21565 , \6674_b0 );
or ( \6744_b1 , \6743_b1 , w_21567 );
not ( w_21567 , w_21568 );
and ( \6744_b0 , \6743_b0 , w_21569 );
and ( w_21568 ,  , w_21569 );
buf ( w_21567 , \6665_b1 );
not ( w_21567 , w_21570 );
not (  , w_21571 );
and ( w_21570 , w_21571 , \6665_b0 );
or ( \6745_b1 , \6742_b1 , w_21573 );
not ( w_21573 , w_21574 );
and ( \6745_b0 , \6742_b0 , w_21575 );
and ( w_21574 ,  , w_21575 );
buf ( w_21573 , \6744_b1 );
not ( w_21573 , w_21576 );
not (  , w_21577 );
and ( w_21576 , w_21577 , \6744_b0 );
buf ( \6746_b1 , \6745_b1 );
not ( \6746_b1 , w_21578 );
not ( \6746_b0 , w_21579 );
and ( w_21578 , w_21579 , \6745_b0 );
or ( \6747_b1 , \6728_b1 , w_21580 );
or ( \6747_b0 , \6728_b0 , \6746_b0 );
not ( \6746_b0 , w_21581 );
and ( w_21581 , w_21580 , \6746_b1 );
or ( \6748_b1 , \6742_b1 , w_21582 );
or ( \6748_b0 , \6742_b0 , \6744_b0 );
not ( \6744_b0 , w_21583 );
and ( w_21583 , w_21582 , \6744_b1 );
or ( \6749_b1 , \6747_b1 , w_21585 );
not ( w_21585 , w_21586 );
and ( \6749_b0 , \6747_b0 , w_21587 );
and ( w_21586 ,  , w_21587 );
buf ( w_21585 , \6748_b1 );
not ( w_21585 , w_21588 );
not (  , w_21589 );
and ( w_21588 , w_21589 , \6748_b0 );
or ( \6750_b1 , \6625_b1 , \6635_b1 );
xor ( \6750_b0 , \6625_b0 , w_21590 );
not ( w_21590 , w_21591 );
and ( w_21591 , \6635_b1 , \6635_b0 );
or ( \6751_b1 , \6750_b1 , \6646_b1 );
xor ( \6751_b0 , \6750_b0 , w_21592 );
not ( w_21592 , w_21593 );
and ( w_21593 , \6646_b1 , \6646_b0 );
buf ( \6752_b1 , \6729_b1 );
not ( \6752_b1 , w_21594 );
not ( \6752_b0 , w_21595 );
and ( w_21594 , w_21595 , \6729_b0 );
buf ( \6753_b1 , \6735_b1 );
not ( \6753_b1 , w_21596 );
not ( \6753_b0 , w_21597 );
and ( w_21596 , w_21597 , \6735_b0 );
or ( \6754_b1 , \6752_b1 , w_21598 );
or ( \6754_b0 , \6752_b0 , \6753_b0 );
not ( \6753_b0 , w_21599 );
and ( w_21599 , w_21598 , \6753_b1 );
or ( \6755_b1 , \6754_b1 , w_21601 );
not ( w_21601 , w_21602 );
and ( \6755_b0 , \6754_b0 , w_21603 );
and ( w_21602 ,  , w_21603 );
buf ( w_21601 , \6741_b1 );
not ( w_21601 , w_21604 );
not (  , w_21605 );
and ( w_21604 , w_21605 , \6741_b0 );
or ( \6756_b1 , \6729_b1 , w_21606 );
or ( \6756_b0 , \6729_b0 , \6735_b0 );
not ( \6735_b0 , w_21607 );
and ( w_21607 , w_21606 , \6735_b1 );
or ( \6757_b1 , \6755_b1 , \6756_b1 );
not ( \6756_b1 , w_21608 );
and ( \6757_b0 , \6755_b0 , w_21609 );
and ( w_21608 , w_21609 , \6756_b0 );
or ( \6758_b1 , \6751_b1 , w_21611 );
not ( w_21611 , w_21612 );
and ( \6758_b0 , \6751_b0 , w_21613 );
and ( w_21612 ,  , w_21613 );
buf ( w_21611 , \6757_b1 );
not ( w_21611 , w_21614 );
not (  , w_21615 );
and ( w_21614 , w_21615 , \6757_b0 );
or ( \6760_b1 , \6751_b1 , w_21617 );
not ( w_21617 , w_21618 );
and ( \6760_b0 , \6751_b0 , w_21619 );
and ( w_21618 ,  , w_21619 );
buf ( w_21617 , \6757_b1 );
not ( w_21617 , w_21620 );
not (  , w_21621 );
and ( w_21620 , w_21621 , \6757_b0 );
or ( \6761_b1 , \6650_b1 , w_21623 );
not ( w_21623 , w_21624 );
and ( \6761_b0 , \6650_b0 , w_21625 );
and ( w_21624 ,  , w_21625 );
buf ( w_21623 , \6760_b1 );
not ( w_21623 , w_21626 );
not (  , w_21627 );
and ( w_21626 , w_21627 , \6760_b0 );
or ( \6762_b1 , \6620_b1 , w_21628 );
or ( \6762_b0 , \6620_b0 , \6649_b0 );
not ( \6649_b0 , w_21629 );
and ( w_21629 , w_21628 , \6649_b1 );
buf ( \6764_b1 , \6763_b1 );
not ( \6764_b1 , w_21630 );
not ( \6764_b0 , w_21631 );
and ( w_21630 , w_21631 , \6763_b0 );
or ( \6765_b1 , \6614_b1 , w_21632 );
or ( \6765_b0 , \6614_b0 , \6764_b0 );
not ( \6764_b0 , w_21633 );
and ( w_21633 , w_21632 , \6764_b1 );
or ( \6766_b1 , \6576_b1 , w_21634 );
or ( \6766_b0 , \6576_b0 , \6612_b0 );
not ( \6612_b0 , w_21635 );
and ( w_21635 , w_21634 , \6612_b1 );
or ( \6767_b1 , \6765_b1 , w_21637 );
not ( w_21637 , w_21638 );
and ( \6767_b0 , \6765_b0 , w_21639 );
and ( w_21638 ,  , w_21639 );
buf ( w_21637 , \6766_b1 );
not ( w_21637 , w_21640 );
not (  , w_21641 );
and ( w_21640 , w_21641 , \6766_b0 );
or ( \6769_b1 , \6570_b1 , w_21643 );
not ( w_21643 , w_21644 );
and ( \6769_b0 , \6570_b0 , w_21645 );
and ( w_21644 ,  , w_21645 );
buf ( w_21643 , \6768_b1 );
not ( w_21643 , w_21646 );
not (  , w_21647 );
and ( w_21646 , w_21647 , \6768_b0 );
or ( \6770_b1 , \6135_b1 , \6189_b1 );
not ( \6189_b1 , w_21648 );
and ( \6770_b0 , \6135_b0 , w_21649 );
and ( w_21648 , w_21649 , \6189_b0 );
buf ( \6771_b1 , \6135_b1 );
not ( \6771_b1 , w_21650 );
not ( \6771_b0 , w_21651 );
and ( w_21650 , w_21651 , \6135_b0 );
or ( \6772_b1 , \6771_b1 , \6190_b1 );
not ( \6190_b1 , w_21652 );
and ( \6772_b0 , \6771_b0 , w_21653 );
and ( w_21652 , w_21653 , \6190_b0 );
or ( \6773_b1 , \6770_b1 , w_21655 );
not ( w_21655 , w_21656 );
and ( \6773_b0 , \6770_b0 , w_21657 );
and ( w_21656 ,  , w_21657 );
buf ( w_21655 , \6772_b1 );
not ( w_21655 , w_21658 );
not (  , w_21659 );
and ( w_21658 , w_21659 , \6772_b0 );
buf ( \6774_b1 , \6773_b1 );
not ( \6774_b1 , w_21660 );
not ( \6774_b0 , w_21661 );
and ( w_21660 , w_21661 , \6773_b0 );
buf ( \6775_b1 , \6146_b1 );
not ( \6775_b1 , w_21662 );
not ( \6775_b0 , w_21663 );
and ( w_21662 , w_21663 , \6146_b0 );
or ( \6776_b1 , \6774_b1 , w_21664 );
or ( \6776_b0 , \6774_b0 , \6775_b0 );
not ( \6775_b0 , w_21665 );
and ( w_21665 , w_21664 , \6775_b1 );
or ( \6777_b1 , \6773_b1 , w_21666 );
or ( \6777_b0 , \6773_b0 , \6146_b0 );
not ( \6146_b0 , w_21667 );
and ( w_21667 , w_21666 , \6146_b1 );
or ( \6778_b1 , \6776_b1 , w_21669 );
not ( w_21669 , w_21670 );
and ( \6778_b0 , \6776_b0 , w_21671 );
and ( w_21670 ,  , w_21671 );
buf ( w_21669 , \6777_b1 );
not ( w_21669 , w_21672 );
not (  , w_21673 );
and ( w_21672 , w_21673 , \6777_b0 );
buf ( \6779_b1 , \6778_b1 );
not ( \6779_b1 , w_21674 );
not ( \6779_b0 , w_21675 );
and ( w_21674 , w_21675 , \6778_b0 );
or ( \6780_b1 , \6065_b1 , \6082_b1 );
xor ( \6780_b0 , \6065_b0 , w_21676 );
not ( w_21676 , w_21677 );
and ( w_21677 , \6082_b1 , \6082_b0 );
or ( \6781_b1 , \6780_b1 , \6115_b1 );
xor ( \6781_b0 , \6780_b0 , w_21678 );
not ( w_21678 , w_21679 );
and ( w_21679 , \6115_b1 , \6115_b0 );
or ( \6782_b1 , \6318_b1 , \6322_b1 );
xor ( \6782_b0 , \6318_b0 , w_21680 );
not ( w_21680 , w_21681 );
and ( w_21681 , \6322_b1 , \6322_b0 );
or ( \6783_b1 , \6782_b1 , \6325_b1 );
not ( \6325_b1 , w_21682 );
and ( \6783_b0 , \6782_b0 , w_21683 );
and ( w_21682 , w_21683 , \6325_b0 );
or ( \6784_b1 , \6318_b1 , \6322_b1 );
not ( \6322_b1 , w_21684 );
and ( \6784_b0 , \6318_b0 , w_21685 );
and ( w_21684 , w_21685 , \6322_b0 );
or ( \6785_b1 , \6783_b1 , w_21686 );
or ( \6785_b0 , \6783_b0 , \6784_b0 );
not ( \6784_b0 , w_21687 );
and ( w_21687 , w_21686 , \6784_b1 );
or ( \6786_b1 , \6781_b1 , \6785_b1 );
xor ( \6786_b0 , \6781_b0 , w_21688 );
not ( w_21688 , w_21689 );
and ( w_21689 , \6785_b1 , \6785_b0 );
buf ( \6787_b1 , \6149_b1 );
not ( \6787_b1 , w_21690 );
not ( \6787_b0 , w_21691 );
and ( w_21690 , w_21691 , \6149_b0 );
buf ( \6788_b1 , \6186_b1 );
not ( \6788_b1 , w_21692 );
not ( \6788_b0 , w_21693 );
and ( w_21692 , w_21693 , \6186_b0 );
or ( \6789_b1 , \6787_b1 , w_21694 );
or ( \6789_b0 , \6787_b0 , \6788_b0 );
not ( \6788_b0 , w_21695 );
and ( w_21695 , w_21694 , \6788_b1 );
or ( \6790_b1 , \6152_b1 , w_21697 );
not ( w_21697 , w_21698 );
and ( \6790_b0 , \6152_b0 , w_21699 );
and ( w_21698 ,  , w_21699 );
buf ( w_21697 , \6187_b1 );
not ( w_21697 , w_21700 );
not (  , w_21701 );
and ( w_21700 , w_21701 , \6187_b0 );
or ( \6791_b1 , \6789_b1 , w_21703 );
not ( w_21703 , w_21704 );
and ( \6791_b0 , \6789_b0 , w_21705 );
and ( w_21704 ,  , w_21705 );
buf ( w_21703 , \6790_b1 );
not ( w_21703 , w_21706 );
not (  , w_21707 );
and ( w_21706 , w_21707 , \6790_b0 );
or ( \6792_b1 , \6791_b1 , \6184_b1 );
not ( \6184_b1 , w_21708 );
and ( \6792_b0 , \6791_b0 , w_21709 );
and ( w_21708 , w_21709 , \6184_b0 );
buf ( \6793_b1 , \6791_b1 );
not ( \6793_b1 , w_21710 );
not ( \6793_b0 , w_21711 );
and ( w_21710 , w_21711 , \6791_b0 );
buf ( \6794_b1 , \6184_b1 );
not ( \6794_b1 , w_21712 );
not ( \6794_b0 , w_21713 );
and ( w_21712 , w_21713 , \6184_b0 );
or ( \6795_b1 , \6793_b1 , \6794_b1 );
not ( \6794_b1 , w_21714 );
and ( \6795_b0 , \6793_b0 , w_21715 );
and ( w_21714 , w_21715 , \6794_b0 );
or ( \6796_b1 , \6792_b1 , w_21717 );
not ( w_21717 , w_21718 );
and ( \6796_b0 , \6792_b0 , w_21719 );
and ( w_21718 ,  , w_21719 );
buf ( w_21717 , \6795_b1 );
not ( w_21717 , w_21720 );
not (  , w_21721 );
and ( w_21720 , w_21721 , \6795_b0 );
or ( \6797_b1 , \6786_b1 , \6796_b1 );
not ( \6796_b1 , w_21722 );
and ( \6797_b0 , \6786_b0 , w_21723 );
and ( w_21722 , w_21723 , \6796_b0 );
or ( \6798_b1 , \6781_b1 , \6785_b1 );
not ( \6785_b1 , w_21724 );
and ( \6798_b0 , \6781_b0 , w_21725 );
and ( w_21724 , w_21725 , \6785_b0 );
or ( \6799_b1 , \6797_b1 , w_21726 );
or ( \6799_b0 , \6797_b0 , \6798_b0 );
not ( \6798_b0 , w_21727 );
and ( w_21727 , w_21726 , \6798_b1 );
buf ( \6800_b1 , \6799_b1 );
not ( \6800_b1 , w_21728 );
not ( \6800_b0 , w_21729 );
and ( w_21728 , w_21729 , \6799_b0 );
or ( \6801_b1 , \6779_b1 , w_21731 );
not ( w_21731 , w_21732 );
and ( \6801_b0 , \6779_b0 , w_21733 );
and ( w_21732 ,  , w_21733 );
buf ( w_21731 , \6800_b1 );
not ( w_21731 , w_21734 );
not (  , w_21735 );
and ( w_21734 , w_21735 , \6800_b0 );
or ( \6802_b1 , \6781_b1 , \6785_b1 );
xor ( \6802_b0 , \6781_b0 , w_21736 );
not ( w_21736 , w_21737 );
and ( w_21737 , \6785_b1 , \6785_b0 );
or ( \6803_b1 , \6802_b1 , \6796_b1 );
xor ( \6803_b0 , \6802_b0 , w_21738 );
not ( w_21738 , w_21739 );
and ( w_21739 , \6796_b1 , \6796_b0 );
buf ( \6804_b1 , \6803_b1 );
not ( \6804_b1 , w_21740 );
not ( \6804_b0 , w_21741 );
and ( w_21740 , w_21741 , \6803_b0 );
or ( \6805_b1 , \6326_b1 , w_21742 );
or ( \6805_b0 , \6326_b0 , \6288_b0 );
not ( \6288_b0 , w_21743 );
and ( w_21743 , w_21742 , \6288_b1 );
buf ( \6806_b1 , \6200_b1 );
buf ( \6806_b0 , \6200_b0 );
or ( \6807_b1 , \6805_b1 , w_21745 );
not ( w_21745 , w_21746 );
and ( \6807_b0 , \6805_b0 , w_21747 );
and ( w_21746 ,  , w_21747 );
buf ( w_21745 , \6806_b1 );
not ( w_21745 , w_21748 );
not (  , w_21749 );
and ( w_21748 , w_21749 , \6806_b0 );
or ( \6808_b1 , \6326_b1 , w_21751 );
not ( w_21751 , w_21752 );
and ( \6808_b0 , \6326_b0 , w_21753 );
and ( w_21752 ,  , w_21753 );
buf ( w_21751 , \6288_b1 );
not ( w_21751 , w_21754 );
not (  , w_21755 );
and ( w_21754 , w_21755 , \6288_b0 );
or ( \6809_b1 , \6807_b1 , w_21757 );
not ( w_21757 , w_21758 );
and ( \6809_b0 , \6807_b0 , w_21759 );
and ( w_21758 ,  , w_21759 );
buf ( w_21757 , \6808_b1 );
not ( w_21757 , w_21760 );
not (  , w_21761 );
and ( w_21760 , w_21761 , \6808_b0 );
buf ( \6810_b1 , \6809_b1 );
not ( \6810_b1 , w_21762 );
not ( \6810_b0 , w_21763 );
and ( w_21762 , w_21763 , \6809_b0 );
or ( \6811_b1 , \6804_b1 , w_21765 );
not ( w_21765 , w_21766 );
and ( \6811_b0 , \6804_b0 , w_21767 );
and ( w_21766 ,  , w_21767 );
buf ( w_21765 , \6810_b1 );
not ( w_21765 , w_21768 );
not (  , w_21769 );
and ( w_21768 , w_21769 , \6810_b0 );
or ( \6812_b1 , \6801_b1 , \6811_b1 );
not ( \6811_b1 , w_21770 );
and ( \6812_b0 , \6801_b0 , w_21771 );
and ( w_21770 , w_21771 , \6811_b0 );
buf ( \6814_b1 , \6126_b1 );
not ( \6814_b1 , w_21772 );
not ( \6814_b0 , w_21773 );
and ( w_21772 , w_21773 , \6126_b0 );
buf ( \6815_b1 , \6023_b1 );
not ( \6815_b1 , w_21774 );
not ( \6815_b0 , w_21775 );
and ( w_21774 , w_21775 , \6023_b0 );
or ( \6816_b1 , \6814_b1 , w_21777 );
not ( w_21777 , w_21778 );
and ( \6816_b0 , \6814_b0 , w_21779 );
and ( w_21778 ,  , w_21779 );
buf ( w_21777 , \6815_b1 );
not ( w_21777 , w_21780 );
not (  , w_21781 );
and ( w_21780 , w_21781 , \6815_b0 );
buf ( \6817_b1 , \6816_b1 );
not ( \6817_b1 , w_21782 );
not ( \6817_b0 , w_21783 );
and ( w_21782 , w_21783 , \6816_b0 );
buf ( \6818_b1 , \6197_b1 );
not ( \6818_b1 , w_21784 );
not ( \6818_b0 , w_21785 );
and ( w_21784 , w_21785 , \6197_b0 );
or ( \6819_b1 , \6817_b1 , w_21786 );
or ( \6819_b0 , \6817_b0 , \6818_b0 );
not ( \6818_b0 , w_21787 );
and ( w_21787 , w_21786 , \6818_b1 );
buf ( \6820_b1 , \6133_b1 );
not ( \6820_b1 , w_21788 );
not ( \6820_b0 , w_21789 );
and ( w_21788 , w_21789 , \6133_b0 );
buf ( \6821_b1 , \6195_b1 );
not ( \6821_b1 , w_21790 );
not ( \6821_b0 , w_21791 );
and ( w_21790 , w_21791 , \6195_b0 );
or ( \6822_b1 , \6820_b1 , w_21793 );
not ( w_21793 , w_21794 );
and ( \6822_b0 , \6820_b0 , w_21795 );
and ( w_21794 ,  , w_21795 );
buf ( w_21793 , \6821_b1 );
not ( w_21793 , w_21796 );
not (  , w_21797 );
and ( w_21796 , w_21797 , \6821_b0 );
or ( \6823_b1 , \6778_b1 , w_21799 );
not ( w_21799 , w_21800 );
and ( \6823_b0 , \6778_b0 , w_21801 );
and ( w_21800 ,  , w_21801 );
buf ( w_21799 , \6799_b1 );
not ( w_21799 , w_21802 );
not (  , w_21803 );
and ( w_21802 , w_21803 , \6799_b0 );
buf ( \6824_b1 , \6823_b1 );
not ( \6824_b1 , w_21804 );
not ( \6824_b0 , w_21805 );
and ( w_21804 , w_21805 , \6823_b0 );
or ( \6825_b1 , \6803_b1 , w_21807 );
not ( w_21807 , w_21808 );
and ( \6825_b0 , \6803_b0 , w_21809 );
and ( w_21808 ,  , w_21809 );
buf ( w_21807 , \6809_b1 );
not ( w_21807 , w_21810 );
not (  , w_21811 );
and ( w_21810 , w_21811 , \6809_b0 );
buf ( \6826_b1 , \6825_b1 );
not ( \6826_b1 , w_21812 );
not ( \6826_b0 , w_21813 );
and ( w_21812 , w_21813 , \6825_b0 );
or ( \6827_b1 , \6824_b1 , w_21814 );
or ( \6827_b0 , \6824_b0 , \6826_b0 );
not ( \6826_b0 , w_21815 );
and ( w_21815 , w_21814 , \6826_b1 );
or ( \6828_b1 , \6827_b1 , w_21817 );
not ( w_21817 , w_21818 );
and ( \6828_b0 , \6827_b0 , w_21819 );
and ( w_21818 ,  , w_21819 );
buf ( w_21817 , \6801_b1 );
not ( w_21817 , w_21820 );
not (  , w_21821 );
and ( w_21820 , w_21821 , \6801_b0 );
or ( \6830_b1 , \6819_b1 , w_21823 );
not ( w_21823 , w_21824 );
and ( \6830_b0 , \6819_b0 , w_21825 );
and ( w_21824 ,  , w_21825 );
buf ( w_21823 , \6829_b1 );
not ( w_21823 , w_21826 );
not (  , w_21827 );
and ( w_21826 , w_21827 , \6829_b0 );
or ( \6831_b1 , \6813_b1 , w_21829 );
not ( w_21829 , w_21830 );
and ( \6831_b0 , \6813_b0 , w_21831 );
and ( w_21830 ,  , w_21831 );
buf ( w_21829 , \6830_b1 );
not ( w_21829 , w_21832 );
not (  , w_21833 );
and ( w_21832 , w_21833 , \6830_b0 );
buf ( \6832_b1 , \5740_b1 );
not ( \6832_b1 , w_21834 );
not ( \6832_b0 , w_21835 );
and ( w_21834 , w_21835 , \5740_b0 );
buf ( \6833_b1 , \5686_b1 );
not ( \6833_b1 , w_21836 );
not ( \6833_b0 , w_21837 );
and ( w_21836 , w_21837 , \5686_b0 );
buf ( \6834_b1 , \5690_b1 );
not ( \6834_b1 , w_21838 );
not ( \6834_b0 , w_21839 );
and ( w_21838 , w_21839 , \5690_b0 );
or ( \6835_b1 , \6833_b1 , \6834_b1 );
not ( \6834_b1 , w_21840 );
and ( \6835_b0 , \6833_b0 , w_21841 );
and ( w_21840 , w_21841 , \6834_b0 );
or ( \6836_b1 , \5686_b1 , \5690_b1 );
not ( \5690_b1 , w_21842 );
and ( \6836_b0 , \5686_b0 , w_21843 );
and ( w_21842 , w_21843 , \5690_b0 );
or ( \6837_b1 , \6835_b1 , w_21845 );
not ( w_21845 , w_21846 );
and ( \6837_b0 , \6835_b0 , w_21847 );
and ( w_21846 ,  , w_21847 );
buf ( w_21845 , \6836_b1 );
not ( w_21845 , w_21848 );
not (  , w_21849 );
and ( w_21848 , w_21849 , \6836_b0 );
buf ( \6838_b1 , \6837_b1 );
not ( \6838_b1 , w_21850 );
not ( \6838_b0 , w_21851 );
and ( w_21850 , w_21851 , \6837_b0 );
or ( \6839_b1 , \6832_b1 , w_21852 );
or ( \6839_b0 , \6832_b0 , \6838_b0 );
not ( \6838_b0 , w_21853 );
and ( w_21853 , w_21852 , \6838_b1 );
or ( \6840_b1 , \5740_b1 , w_21854 );
or ( \6840_b0 , \5740_b0 , \6837_b0 );
not ( \6837_b0 , w_21855 );
and ( w_21855 , w_21854 , \6837_b1 );
or ( \6841_b1 , \6839_b1 , w_21857 );
not ( w_21857 , w_21858 );
and ( \6841_b0 , \6839_b0 , w_21859 );
and ( w_21858 ,  , w_21859 );
buf ( w_21857 , \6840_b1 );
not ( w_21857 , w_21860 );
not (  , w_21861 );
and ( w_21860 , w_21861 , \6840_b0 );
buf ( \6842_b1 , \6841_b1 );
not ( \6842_b1 , w_21862 );
not ( \6842_b0 , w_21863 );
and ( w_21862 , w_21863 , \6841_b0 );
or ( \6843_b1 , \5954_b1 , \5956_b1 );
xor ( \6843_b0 , \5954_b0 , w_21864 );
not ( w_21864 , w_21865 );
and ( w_21865 , \5956_b1 , \5956_b0 );
or ( \6844_b1 , \6843_b1 , \5959_b1 );
not ( \5959_b1 , w_21866 );
and ( \6844_b0 , \6843_b0 , w_21867 );
and ( w_21866 , w_21867 , \5959_b0 );
or ( \6845_b1 , \5954_b1 , \5956_b1 );
not ( \5956_b1 , w_21868 );
and ( \6845_b0 , \5954_b0 , w_21869 );
and ( w_21868 , w_21869 , \5956_b0 );
or ( \6846_b1 , \6844_b1 , w_21870 );
or ( \6846_b0 , \6844_b0 , \6845_b0 );
not ( \6845_b0 , w_21871 );
and ( w_21871 , w_21870 , \6845_b1 );
buf ( \6847_b1 , \6009_b1 );
not ( \6847_b1 , w_21872 );
not ( \6847_b0 , w_21873 );
and ( w_21872 , w_21873 , \6009_b0 );
or ( \6848_b1 , \6847_b1 , w_21875 );
not ( w_21875 , w_21876 );
and ( \6848_b0 , \6847_b0 , w_21877 );
and ( w_21876 ,  , w_21877 );
buf ( w_21875 , \6006_b1 );
not ( w_21875 , w_21878 );
not (  , w_21879 );
and ( w_21878 , w_21879 , \6006_b0 );
buf ( \6849_b1 , \6848_b1 );
not ( \6849_b1 , w_21880 );
not ( \6849_b0 , w_21881 );
and ( w_21880 , w_21881 , \6848_b0 );
buf ( \6850_b1 , \6001_b1 );
not ( \6850_b1 , w_21882 );
not ( \6850_b0 , w_21883 );
and ( w_21882 , w_21883 , \6001_b0 );
or ( \6851_b1 , \6849_b1 , w_21884 );
or ( \6851_b0 , \6849_b0 , \6850_b0 );
not ( \6850_b0 , w_21885 );
and ( w_21885 , w_21884 , \6850_b1 );
or ( \6852_b1 , \6847_b1 , w_21886 );
or ( \6852_b0 , \6847_b0 , \6006_b0 );
not ( \6006_b0 , w_21887 );
and ( w_21887 , w_21886 , \6006_b1 );
or ( \6853_b1 , \6851_b1 , w_21889 );
not ( w_21889 , w_21890 );
and ( \6853_b0 , \6851_b0 , w_21891 );
and ( w_21890 ,  , w_21891 );
buf ( w_21889 , \6852_b1 );
not ( w_21889 , w_21892 );
not (  , w_21893 );
and ( w_21892 , w_21893 , \6852_b0 );
or ( \6854_b1 , \6846_b1 , \6853_b1 );
xor ( \6854_b0 , \6846_b0 , w_21894 );
not ( w_21894 , w_21895 );
and ( w_21895 , \6853_b1 , \6853_b0 );
or ( \6855_b1 , \5732_b1 , \5734_b1 );
xor ( \6855_b0 , \5732_b0 , w_21896 );
not ( w_21896 , w_21897 );
and ( w_21897 , \5734_b1 , \5734_b0 );
or ( \6856_b1 , \6855_b1 , \5737_b1 );
xor ( \6856_b0 , \6855_b0 , w_21898 );
not ( w_21898 , w_21899 );
and ( w_21899 , \5737_b1 , \5737_b0 );
or ( \6857_b1 , \6854_b1 , \6856_b1 );
not ( \6856_b1 , w_21900 );
and ( \6857_b0 , \6854_b0 , w_21901 );
and ( w_21900 , w_21901 , \6856_b0 );
or ( \6858_b1 , \6846_b1 , \6853_b1 );
not ( \6853_b1 , w_21902 );
and ( \6858_b0 , \6846_b0 , w_21903 );
and ( w_21902 , w_21903 , \6853_b0 );
or ( \6859_b1 , \6857_b1 , w_21904 );
or ( \6859_b0 , \6857_b0 , \6858_b0 );
not ( \6858_b0 , w_21905 );
and ( w_21905 , w_21904 , \6858_b1 );
buf ( \6860_b1 , \6859_b1 );
not ( \6860_b1 , w_21906 );
not ( \6860_b0 , w_21907 );
and ( w_21906 , w_21907 , \6859_b0 );
or ( \6861_b1 , \6842_b1 , w_21909 );
not ( w_21909 , w_21910 );
and ( \6861_b0 , \6842_b0 , w_21911 );
and ( w_21910 ,  , w_21911 );
buf ( w_21909 , \6860_b1 );
not ( w_21909 , w_21912 );
not (  , w_21913 );
and ( w_21912 , w_21913 , \6860_b0 );
or ( \6862_b1 , \6846_b1 , \6853_b1 );
xor ( \6862_b0 , \6846_b0 , w_21914 );
not ( w_21914 , w_21915 );
and ( w_21915 , \6853_b1 , \6853_b0 );
or ( \6863_b1 , \6862_b1 , \6856_b1 );
xor ( \6863_b0 , \6862_b0 , w_21916 );
not ( w_21916 , w_21917 );
and ( w_21917 , \6856_b1 , \6856_b0 );
buf ( \6864_b1 , \6863_b1 );
not ( \6864_b1 , w_21918 );
not ( \6864_b0 , w_21919 );
and ( w_21918 , w_21919 , \6863_b0 );
buf ( \6865_b1 , \6018_b1 );
not ( \6865_b1 , w_21920 );
not ( \6865_b0 , w_21921 );
and ( w_21920 , w_21921 , \6018_b0 );
buf ( \6866_b1 , \5965_b1 );
not ( \6866_b1 , w_21922 );
not ( \6866_b0 , w_21923 );
and ( w_21922 , w_21923 , \5965_b0 );
or ( \6867_b1 , \6865_b1 , w_21924 );
or ( \6867_b0 , \6865_b0 , \6866_b0 );
not ( \6866_b0 , w_21925 );
and ( w_21925 , w_21924 , \6866_b1 );
buf ( \6868_b1 , \5965_b1 );
not ( \6868_b1 , w_21926 );
not ( \6868_b0 , w_21927 );
and ( w_21926 , w_21927 , \5965_b0 );
buf ( \6869_b1 , \6868_b1 );
not ( \6869_b1 , w_21928 );
not ( \6869_b0 , w_21929 );
and ( w_21928 , w_21929 , \6868_b0 );
buf ( \6870_b1 , \6019_b1 );
not ( \6870_b1 , w_21930 );
not ( \6870_b0 , w_21931 );
and ( w_21930 , w_21931 , \6019_b0 );
or ( \6871_b1 , \6869_b1 , w_21932 );
or ( \6871_b0 , \6869_b0 , \6870_b0 );
not ( \6870_b0 , w_21933 );
and ( w_21933 , w_21932 , \6870_b1 );
or ( \6872_b1 , \6871_b1 , w_21935 );
not ( w_21935 , w_21936 );
and ( \6872_b0 , \6871_b0 , w_21937 );
and ( w_21936 ,  , w_21937 );
buf ( w_21935 , \5922_b1 );
not ( w_21935 , w_21938 );
not (  , w_21939 );
and ( w_21938 , w_21939 , \5922_b0 );
or ( \6873_b1 , \6867_b1 , w_21941 );
not ( w_21941 , w_21942 );
and ( \6873_b0 , \6867_b0 , w_21943 );
and ( w_21942 ,  , w_21943 );
buf ( w_21941 , \6872_b1 );
not ( w_21941 , w_21944 );
not (  , w_21945 );
and ( w_21944 , w_21945 , \6872_b0 );
buf ( \6874_b1 , \6873_b1 );
not ( \6874_b1 , w_21946 );
not ( \6874_b0 , w_21947 );
and ( w_21946 , w_21947 , \6873_b0 );
or ( \6875_b1 , \6864_b1 , w_21949 );
not ( w_21949 , w_21950 );
and ( \6875_b0 , \6864_b0 , w_21951 );
and ( w_21950 ,  , w_21951 );
buf ( w_21949 , \6874_b1 );
not ( w_21949 , w_21952 );
not (  , w_21953 );
and ( w_21952 , w_21953 , \6874_b0 );
or ( \6876_b1 , \6861_b1 , \6875_b1 );
not ( \6875_b1 , w_21954 );
and ( \6876_b0 , \6861_b0 , w_21955 );
and ( w_21954 , w_21955 , \6875_b0 );
or ( \6878_b1 , \6841_b1 , w_21957 );
not ( w_21957 , w_21958 );
and ( \6878_b0 , \6841_b0 , w_21959 );
and ( w_21958 ,  , w_21959 );
buf ( w_21957 , \6859_b1 );
not ( w_21957 , w_21960 );
not (  , w_21961 );
and ( w_21960 , w_21961 , \6859_b0 );
or ( \6879_b1 , \6863_b1 , w_21963 );
not ( w_21963 , w_21964 );
and ( \6879_b0 , \6863_b0 , w_21965 );
and ( w_21964 ,  , w_21965 );
buf ( w_21963 , \6873_b1 );
not ( w_21963 , w_21966 );
not (  , w_21967 );
and ( w_21966 , w_21967 , \6873_b0 );
or ( \6880_b1 , \6878_b1 , w_21969 );
not ( w_21969 , w_21970 );
and ( \6880_b0 , \6878_b0 , w_21971 );
and ( w_21970 ,  , w_21971 );
buf ( w_21969 , \6879_b1 );
not ( w_21969 , w_21972 );
not (  , w_21973 );
and ( w_21972 , w_21973 , \6879_b0 );
or ( \6881_b1 , \6880_b1 , \6861_b1 );
not ( \6861_b1 , w_21974 );
and ( \6881_b0 , \6880_b0 , w_21975 );
and ( w_21974 , w_21975 , \6861_b0 );
or ( \6882_b1 , \6881_b1 , w_21977 );
not ( w_21977 , w_21978 );
and ( \6882_b0 , \6881_b0 , w_21979 );
and ( w_21978 ,  , w_21979 );
buf ( w_21977 , \5745_b1 );
not ( w_21977 , w_21980 );
not (  , w_21981 );
and ( w_21980 , w_21981 , \5745_b0 );
buf ( \6883_b1 , \5682_b1 );
buf ( \6883_b0 , \5682_b0 );
or ( \6884_b1 , \5684_b1 , w_21983 );
not ( w_21983 , w_21984 );
and ( \6884_b0 , \5684_b0 , w_21985 );
and ( w_21984 ,  , w_21985 );
buf ( w_21983 , \5743_b1 );
not ( w_21983 , w_21986 );
not (  , w_21987 );
and ( w_21986 , w_21987 , \5743_b0 );
or ( \6885_b1 , \6883_b1 , \6884_b1 );
not ( \6884_b1 , w_21988 );
and ( \6885_b0 , \6883_b0 , w_21989 );
and ( w_21988 , w_21989 , \6884_b0 );
or ( \6886_b1 , \5681_b1 , w_21991 );
not ( w_21991 , w_21992 );
and ( \6886_b0 , \5681_b0 , w_21993 );
and ( w_21992 ,  , w_21993 );
buf ( w_21991 , \5563_b1 );
not ( w_21991 , w_21994 );
not (  , w_21995 );
and ( w_21994 , w_21995 , \5563_b0 );
or ( \6887_b1 , \6885_b1 , w_21997 );
not ( w_21997 , w_21998 );
and ( \6887_b0 , \6885_b0 , w_21999 );
and ( w_21998 ,  , w_21999 );
buf ( w_21997 , \6886_b1 );
not ( w_21997 , w_22000 );
not (  , w_22001 );
and ( w_22000 , w_22001 , \6886_b0 );
buf ( \6889_b1 , \6888_b1 );
not ( \6889_b1 , w_22002 );
not ( \6889_b0 , w_22003 );
and ( w_22002 , w_22003 , \6888_b0 );
or ( \6890_b1 , \5561_b1 , w_22004 );
or ( \6890_b0 , \5561_b0 , \6889_b0 );
not ( \6889_b0 , w_22005 );
and ( w_22005 , w_22004 , \6889_b1 );
or ( \6891_b1 , \5206_b1 , w_22006 );
or ( \6891_b0 , \5206_b0 , \5382_b0 );
not ( \5382_b0 , w_22007 );
and ( w_22007 , w_22006 , \5382_b1 );
or ( \6892_b1 , \5385_b1 , w_22008 );
or ( \6892_b0 , \5385_b0 , \5509_b0 );
not ( \5509_b0 , w_22009 );
and ( w_22009 , w_22008 , \5509_b1 );
or ( \6893_b1 , \6891_b1 , w_22011 );
not ( w_22011 , w_22012 );
and ( \6893_b0 , \6891_b0 , w_22013 );
and ( w_22012 ,  , w_22013 );
buf ( w_22011 , \6892_b1 );
not ( w_22011 , w_22014 );
not (  , w_22015 );
and ( w_22014 , w_22015 , \6892_b0 );
buf ( \6894_b1 , \5383_b1 );
not ( \6894_b1 , w_22016 );
not ( \6894_b0 , w_22017 );
and ( w_22016 , w_22017 , \5383_b0 );
or ( \6895_b1 , \5558_b1 , w_22019 );
not ( w_22019 , w_22020 );
and ( \6895_b0 , \5558_b0 , w_22021 );
and ( w_22020 ,  , w_22021 );
buf ( w_22019 , \6894_b1 );
not ( w_22019 , w_22022 );
not (  , w_22023 );
and ( w_22022 , w_22023 , \6894_b0 );
or ( \6896_b1 , \6893_b1 , \6895_b1 );
not ( \6895_b1 , w_22024 );
and ( \6896_b0 , \6893_b0 , w_22025 );
and ( w_22024 , w_22025 , \6895_b0 );
or ( \6897_b1 , \5538_b1 , w_22026 );
or ( \6897_b0 , \5538_b0 , \5542_b0 );
not ( \5542_b0 , w_22027 );
and ( w_22027 , w_22026 , \5542_b1 );
buf ( \6898_b1 , \5557_b1 );
not ( \6898_b1 , w_22028 );
not ( \6898_b0 , w_22029 );
and ( w_22028 , w_22029 , \5557_b0 );
or ( \6899_b1 , \6897_b1 , w_22030 );
or ( \6899_b0 , \6897_b0 , \6898_b0 );
not ( \6898_b0 , w_22031 );
and ( w_22031 , w_22030 , \6898_b1 );
buf ( \6900_b1 , \5556_b1 );
not ( \6900_b1 , w_22032 );
not ( \6900_b0 , w_22033 );
and ( w_22032 , w_22033 , \5556_b0 );
or ( \6901_b1 , \6900_b1 , w_22035 );
not ( w_22035 , w_22036 );
and ( \6901_b0 , \6900_b0 , w_22037 );
and ( w_22036 ,  , w_22037 );
buf ( w_22035 , \5553_b1 );
not ( w_22035 , w_22038 );
not (  , w_22039 );
and ( w_22038 , w_22039 , \5553_b0 );
or ( \6902_b1 , \6899_b1 , w_22041 );
not ( w_22041 , w_22042 );
and ( \6902_b0 , \6899_b0 , w_22043 );
and ( w_22042 ,  , w_22043 );
buf ( w_22041 , \6901_b1 );
not ( w_22041 , w_22044 );
not (  , w_22045 );
and ( w_22044 , w_22045 , \6901_b0 );
or ( \6903_b1 , \6896_b1 , w_22047 );
not ( w_22047 , w_22048 );
and ( \6903_b0 , \6896_b0 , w_22049 );
and ( w_22048 ,  , w_22049 );
buf ( w_22047 , \6902_b1 );
not ( w_22047 , w_22050 );
not (  , w_22051 );
and ( w_22050 , w_22051 , \6902_b0 );
or ( \6904_b1 , \6890_b1 , w_22053 );
not ( w_22053 , w_22054 );
and ( \6904_b0 , \6890_b0 , w_22055 );
and ( w_22054 ,  , w_22055 );
buf ( w_22053 , \6903_b1 );
not ( w_22053 , w_22056 );
not (  , w_22057 );
and ( w_22056 , w_22057 , \6903_b0 );
buf ( \6905_b1 , \6904_b1 );
not ( \6905_b1 , w_22058 );
not ( \6905_b0 , w_22059 );
and ( w_22058 , w_22059 , \6904_b0 );
or ( \6906_b1 , \4985_b1 , w_22060 );
or ( \6906_b0 , \4985_b0 , \6905_b0 );
not ( \6905_b0 , w_22061 );
and ( w_22061 , w_22060 , \6905_b1 );
buf ( \6907_b1 , \4960_b1 );
not ( \6907_b1 , w_22062 );
not ( \6907_b0 , w_22063 );
and ( w_22062 , w_22063 , \4960_b0 );
buf ( \6908_b1 , \6907_b1 );
not ( \6908_b1 , w_22064 );
not ( \6908_b0 , w_22065 );
and ( w_22064 , w_22065 , \6907_b0 );
buf ( \6909_b1 , \4927_b1 );
not ( \6909_b1 , w_22066 );
not ( \6909_b0 , w_22067 );
and ( w_22066 , w_22067 , \4927_b0 );
or ( \6910_b1 , \4515_b1 , w_22069 );
not ( w_22069 , w_22070 );
and ( \6910_b0 , \4515_b0 , w_22071 );
and ( w_22070 ,  , w_22071 );
buf ( w_22069 , \4692_b1 );
not ( w_22069 , w_22072 );
not (  , w_22073 );
and ( w_22072 , w_22073 , \4692_b0 );
buf ( \6911_b1 , \6910_b1 );
not ( \6911_b1 , w_22074 );
not ( \6911_b0 , w_22075 );
and ( w_22074 , w_22075 , \6910_b0 );
or ( \6912_b1 , \6911_b1 , w_22077 );
not ( w_22077 , w_22078 );
and ( \6912_b0 , \6911_b0 , w_22079 );
and ( w_22078 ,  , w_22079 );
buf ( w_22077 , \4766_b1 );
not ( w_22077 , w_22080 );
not (  , w_22081 );
and ( w_22080 , w_22081 , \4766_b0 );
or ( \6913_b1 , \4764_b1 , w_22083 );
not ( w_22083 , w_22084 );
and ( \6913_b0 , \4764_b0 , w_22085 );
and ( w_22084 ,  , w_22085 );
buf ( w_22083 , \4698_b1 );
not ( w_22083 , w_22086 );
not (  , w_22087 );
and ( w_22086 , w_22087 , \4698_b0 );
or ( \6914_b1 , \4771_b1 , w_22089 );
not ( w_22089 , w_22090 );
and ( \6914_b0 , \4771_b0 , w_22091 );
and ( w_22090 ,  , w_22091 );
buf ( w_22089 , \4832_b1 );
not ( w_22089 , w_22092 );
not (  , w_22093 );
and ( w_22092 , w_22093 , \4832_b0 );
or ( \6915_b1 , \4840_b1 , w_22095 );
not ( w_22095 , w_22096 );
and ( \6915_b0 , \4840_b0 , w_22097 );
and ( w_22096 ,  , w_22097 );
buf ( w_22095 , \4883_b1 );
not ( w_22095 , w_22098 );
not (  , w_22099 );
and ( w_22098 , w_22099 , \4883_b0 );
or ( \6917_b1 , \6912_b1 , \6916_b1 );
not ( \6916_b1 , w_22100 );
and ( \6917_b0 , \6912_b0 , w_22101 );
and ( w_22100 , w_22101 , \6916_b0 );
or ( \6918_b1 , \4834_b1 , \4885_b1 );
not ( \4885_b1 , w_22102 );
and ( \6918_b0 , \4834_b0 , w_22103 );
and ( w_22102 , w_22103 , \4885_b0 );
buf ( \6919_b1 , \6915_b1 );
not ( \6919_b1 , w_22104 );
not ( \6919_b0 , w_22105 );
and ( w_22104 , w_22105 , \6915_b0 );
or ( \6920_b1 , \6918_b1 , w_22107 );
not ( w_22107 , w_22108 );
and ( \6920_b0 , \6918_b0 , w_22109 );
and ( w_22108 ,  , w_22109 );
buf ( w_22107 , \6919_b1 );
not ( w_22107 , w_22110 );
not (  , w_22111 );
and ( w_22110 , w_22111 , \6919_b0 );
or ( \6921_b1 , \6917_b1 , w_22113 );
not ( w_22113 , w_22114 );
and ( \6921_b0 , \6917_b0 , w_22115 );
and ( w_22114 ,  , w_22115 );
buf ( w_22113 , \6920_b1 );
not ( w_22113 , w_22116 );
not (  , w_22117 );
and ( w_22116 , w_22117 , \6920_b0 );
buf ( \6922_b1 , \6921_b1 );
not ( \6922_b1 , w_22118 );
not ( \6922_b0 , w_22119 );
and ( w_22118 , w_22119 , \6921_b0 );
or ( \6923_b1 , \6909_b1 , w_22120 );
or ( \6923_b0 , \6909_b0 , \6922_b0 );
not ( \6922_b0 , w_22121 );
and ( w_22121 , w_22120 , \6922_b1 );
or ( \6924_b1 , \4920_b1 , w_22122 );
or ( \6924_b0 , \4920_b0 , \4926_b0 );
not ( \4926_b0 , w_22123 );
and ( w_22123 , w_22122 , \4926_b1 );
or ( \6925_b1 , \6923_b1 , w_22125 );
not ( w_22125 , w_22126 );
and ( \6925_b0 , \6923_b0 , w_22127 );
and ( w_22126 ,  , w_22127 );
buf ( w_22125 , \6924_b1 );
not ( w_22125 , w_22128 );
not (  , w_22129 );
and ( w_22128 , w_22129 , \6924_b0 );
buf ( \6926_b1 , \6925_b1 );
not ( \6926_b1 , w_22130 );
not ( \6926_b0 , w_22131 );
and ( w_22130 , w_22131 , \6925_b0 );
or ( \6927_b1 , \6908_b1 , w_22132 );
or ( \6927_b0 , \6908_b0 , \6926_b0 );
not ( \6926_b0 , w_22133 );
and ( w_22133 , w_22132 , \6926_b1 );
or ( \6928_b1 , \4932_b1 , w_22135 );
not ( w_22135 , w_22136 );
and ( \6928_b0 , \4932_b0 , w_22137 );
and ( w_22136 ,  , w_22137 );
buf ( w_22135 , \4959_b1 );
not ( w_22135 , w_22138 );
not (  , w_22139 );
and ( w_22138 , w_22139 , \4959_b0 );
or ( \6929_b1 , \6927_b1 , w_22141 );
not ( w_22141 , w_22142 );
and ( \6929_b0 , \6927_b0 , w_22143 );
and ( w_22142 ,  , w_22143 );
buf ( w_22141 , \6928_b1 );
not ( w_22141 , w_22144 );
not (  , w_22145 );
and ( w_22144 , w_22145 , \6928_b0 );
buf ( \6930_b1 , \4983_b1 );
not ( \6930_b1 , w_22146 );
not ( \6930_b0 , w_22147 );
and ( w_22146 , w_22147 , \4983_b0 );
or ( \6931_b1 , \6929_b1 , \6930_b1 );
not ( \6930_b1 , w_22148 );
and ( \6931_b0 , \6929_b0 , w_22149 );
and ( w_22148 , w_22149 , \6930_b0 );
or ( \6932_b1 , \4964_b1 , \4982_b1 );
not ( \4982_b1 , w_22150 );
and ( \6932_b0 , \4964_b0 , w_22151 );
and ( w_22150 , w_22151 , \4982_b0 );
or ( \6933_b1 , \6931_b1 , w_22153 );
not ( w_22153 , w_22154 );
and ( \6933_b0 , \6931_b0 , w_22155 );
and ( w_22154 ,  , w_22155 );
buf ( w_22153 , \6932_b1 );
not ( w_22153 , w_22156 );
not (  , w_22157 );
and ( w_22156 , w_22157 , \6932_b0 );
or ( \6934_b1 , \6906_b1 , w_22159 );
not ( w_22159 , w_22160 );
and ( \6934_b0 , \6906_b0 , w_22161 );
and ( w_22160 ,  , w_22161 );
buf ( w_22159 , \6933_b1 );
not ( w_22159 , w_22162 );
not (  , w_22163 );
and ( w_22162 , w_22163 , \6933_b0 );
buf ( \6935_b1 , \4978_b1 );
not ( \6935_b1 , w_22164 );
not ( \6935_b0 , w_22165 );
and ( w_22164 , w_22165 , \4978_b0 );
or ( \6936_b1 , \4815_b1 , \6935_b1 );
not ( \6935_b1 , w_22166 );
and ( \6936_b0 , \4815_b0 , w_22167 );
and ( w_22166 , w_22167 , \6935_b0 );
or ( \6937_b1 , \4859_b1 , \4156_b1 );
not ( \4156_b1 , w_22168 );
and ( \6937_b0 , \4859_b0 , w_22169 );
and ( w_22168 , w_22169 , \4156_b0 );
or ( \6938_b1 , \6936_b1 , w_22171 );
not ( w_22171 , w_22172 );
and ( \6938_b0 , \6936_b0 , w_22173 );
and ( w_22172 ,  , w_22173 );
buf ( w_22171 , \6937_b1 );
not ( w_22171 , w_22174 );
not (  , w_22175 );
and ( w_22174 , w_22175 , \6937_b0 );
buf ( \6939_b1 , \6938_b1 );
not ( \6939_b1 , w_22176 );
not ( \6939_b0 , w_22177 );
and ( w_22176 , w_22177 , \6938_b0 );
or ( \6940_b1 , \4156_b1 , w_22179 );
not ( w_22179 , w_22180 );
and ( \6940_b0 , \4156_b0 , w_22181 );
and ( w_22180 ,  , w_22181 );
buf ( w_22179 , \4044_b1 );
not ( w_22179 , w_22182 );
not (  , w_22183 );
and ( w_22182 , w_22183 , \4044_b0 );
buf ( \6941_b1 , \6940_b1 );
not ( \6941_b1 , w_22184 );
not ( \6941_b0 , w_22185 );
and ( w_22184 , w_22185 , \6940_b0 );
or ( \6942_b1 , \6939_b1 , \6941_b1 );
not ( \6941_b1 , w_22186 );
and ( \6942_b0 , \6939_b0 , w_22187 );
and ( w_22186 , w_22187 , \6941_b0 );
or ( \6943_b1 , \6938_b1 , \6940_b1 );
not ( \6940_b1 , w_22188 );
and ( \6943_b0 , \6938_b0 , w_22189 );
and ( w_22188 , w_22189 , \6940_b0 );
or ( \6944_b1 , \6942_b1 , w_22191 );
not ( w_22191 , w_22192 );
and ( \6944_b0 , \6942_b0 , w_22193 );
and ( w_22192 ,  , w_22193 );
buf ( w_22191 , \6943_b1 );
not ( w_22191 , w_22194 );
not (  , w_22195 );
and ( w_22194 , w_22195 , \6943_b0 );
buf ( \6945_b1 , \6944_b1 );
not ( \6945_b1 , w_22196 );
not ( \6945_b0 , w_22197 );
and ( w_22196 , w_22197 , \6944_b0 );
or ( \6946_b1 , \4972_b1 , \4973_b1 );
xor ( \6946_b0 , \4972_b0 , w_22198 );
not ( w_22198 , w_22199 );
and ( w_22199 , \4973_b1 , \4973_b0 );
or ( \6947_b1 , \6946_b1 , \4980_b1 );
not ( \4980_b1 , w_22200 );
and ( \6947_b0 , \6946_b0 , w_22201 );
and ( w_22200 , w_22201 , \4980_b0 );
or ( \6948_b1 , \4972_b1 , \4973_b1 );
not ( \4973_b1 , w_22202 );
and ( \6948_b0 , \4972_b0 , w_22203 );
and ( w_22202 , w_22203 , \4973_b0 );
or ( \6949_b1 , \6947_b1 , w_22204 );
or ( \6949_b0 , \6947_b0 , \6948_b0 );
not ( \6948_b0 , w_22205 );
and ( w_22205 , w_22204 , \6948_b1 );
buf ( \6950_b1 , \6949_b1 );
not ( \6950_b1 , w_22206 );
not ( \6950_b0 , w_22207 );
and ( w_22206 , w_22207 , \6949_b0 );
or ( \6951_b1 , \6945_b1 , w_22208 );
or ( \6951_b0 , \6945_b0 , \6950_b0 );
not ( \6950_b0 , w_22209 );
and ( w_22209 , w_22208 , \6950_b1 );
or ( \6952_b1 , \6949_b1 , w_22210 );
or ( \6952_b0 , \6949_b0 , \6944_b0 );
not ( \6944_b0 , w_22211 );
and ( w_22211 , w_22210 , \6944_b1 );
or ( \6953_b1 , \6951_b1 , w_22213 );
not ( w_22213 , w_22214 );
and ( \6953_b0 , \6951_b0 , w_22215 );
and ( w_22214 ,  , w_22215 );
buf ( w_22213 , \6952_b1 );
not ( w_22213 , w_22216 );
not (  , w_22217 );
and ( w_22216 , w_22217 , \6952_b0 );
buf ( \6954_b1 , \6953_b1 );
not ( \6954_b1 , w_22218 );
not ( \6954_b0 , w_22219 );
and ( w_22218 , w_22219 , \6953_b0 );
or ( \6955_b1 , \4968_b1 , \4969_b1 );
xor ( \6955_b0 , \4968_b0 , w_22220 );
not ( w_22220 , w_22221 );
and ( w_22221 , \4969_b1 , \4969_b0 );
or ( \6956_b1 , \6955_b1 , \4981_b1 );
not ( \4981_b1 , w_22222 );
and ( \6956_b0 , \6955_b0 , w_22223 );
and ( w_22222 , w_22223 , \4981_b0 );
or ( \6957_b1 , \4968_b1 , \4969_b1 );
not ( \4969_b1 , w_22224 );
and ( \6957_b0 , \4968_b0 , w_22225 );
and ( w_22224 , w_22225 , \4969_b0 );
or ( \6958_b1 , \6956_b1 , w_22226 );
or ( \6958_b0 , \6956_b0 , \6957_b0 );
not ( \6957_b0 , w_22227 );
and ( w_22227 , w_22226 , \6957_b1 );
buf ( \6959_b1 , \6958_b1 );
not ( \6959_b1 , w_22228 );
not ( \6959_b0 , w_22229 );
and ( w_22228 , w_22229 , \6958_b0 );
or ( \6960_b1 , \6954_b1 , w_22230 );
or ( \6960_b0 , \6954_b0 , \6959_b0 );
not ( \6959_b0 , w_22231 );
and ( w_22231 , w_22230 , \6959_b1 );
or ( \6961_b1 , \6958_b1 , w_22232 );
or ( \6961_b0 , \6958_b0 , \6953_b0 );
not ( \6953_b0 , w_22233 );
and ( w_22233 , w_22232 , \6953_b1 );
or ( \6962_b1 , \6960_b1 , w_22235 );
not ( w_22235 , w_22236 );
and ( \6962_b0 , \6960_b0 , w_22237 );
and ( w_22236 ,  , w_22237 );
buf ( w_22235 , \6961_b1 );
not ( w_22235 , w_22238 );
not (  , w_22239 );
and ( w_22238 , w_22239 , \6961_b0 );
buf ( \6963_b1 , \6962_b1 );
not ( \6963_b1 , w_22240 );
not ( \6963_b0 , w_22241 );
and ( w_22240 , w_22241 , \6962_b0 );
or ( \6964_b1 , \6934_b1 , \6963_b1 );
not ( \6963_b1 , w_22242 );
and ( \6964_b0 , \6934_b0 , w_22243 );
and ( w_22242 , w_22243 , \6963_b0 );
buf ( \6965_b1 , \6934_b1 );
not ( \6965_b1 , w_22244 );
not ( \6965_b0 , w_22245 );
and ( w_22244 , w_22245 , \6934_b0 );
or ( \6966_b1 , \6965_b1 , \6962_b1 );
not ( \6962_b1 , w_22246 );
and ( \6966_b0 , \6965_b0 , w_22247 );
and ( w_22246 , w_22247 , \6962_b0 );
or ( \6967_b1 , \6964_b1 , w_22249 );
not ( w_22249 , w_22250 );
and ( \6967_b0 , \6964_b0 , w_22251 );
and ( w_22250 ,  , w_22251 );
buf ( w_22249 , \6966_b1 );
not ( w_22249 , w_22252 );
not (  , w_22253 );
and ( w_22252 , w_22253 , \6966_b0 );
buf ( \6968_b1 , \4928_b1 );
not ( \6968_b1 , w_22254 );
not ( \6968_b0 , w_22255 );
and ( w_22254 , w_22255 , \4928_b0 );
buf ( \6969_b1 , \6968_b1 );
not ( \6969_b1 , w_22256 );
not ( \6969_b0 , w_22257 );
and ( w_22256 , w_22257 , \6968_b0 );
buf ( \6970_b1 , \6904_b1 );
not ( \6970_b1 , w_22258 );
not ( \6970_b0 , w_22259 );
and ( w_22258 , w_22259 , \6904_b0 );
or ( \6971_b1 , \6969_b1 , w_22260 );
or ( \6971_b0 , \6969_b0 , \6970_b0 );
not ( \6970_b0 , w_22261 );
and ( w_22261 , w_22260 , \6970_b1 );
buf ( \6972_b1 , \6925_b1 );
not ( \6972_b1 , w_22262 );
not ( \6972_b0 , w_22263 );
and ( w_22262 , w_22263 , \6925_b0 );
or ( \6973_b1 , \6971_b1 , w_22265 );
not ( w_22265 , w_22266 );
and ( \6973_b0 , \6971_b0 , w_22267 );
and ( w_22266 ,  , w_22267 );
buf ( w_22265 , \6972_b1 );
not ( w_22265 , w_22268 );
not (  , w_22269 );
and ( w_22268 , w_22269 , \6972_b0 );
or ( \6974_b1 , \6907_b1 , w_22271 );
not ( w_22271 , w_22272 );
and ( \6974_b0 , \6907_b0 , w_22273 );
and ( w_22272 ,  , w_22273 );
buf ( w_22271 , \6928_b1 );
not ( w_22271 , w_22274 );
not (  , w_22275 );
and ( w_22274 , w_22275 , \6928_b0 );
buf ( \6975_b1 , \6974_b1 );
not ( \6975_b1 , w_22276 );
not ( \6975_b0 , w_22277 );
and ( w_22276 , w_22277 , \6974_b0 );
or ( \6976_b1 , \6973_b1 , \6975_b1 );
not ( \6975_b1 , w_22278 );
and ( \6976_b0 , \6973_b0 , w_22279 );
and ( w_22278 , w_22279 , \6975_b0 );
buf ( \6977_b1 , \6973_b1 );
not ( \6977_b1 , w_22280 );
not ( \6977_b0 , w_22281 );
and ( w_22280 , w_22281 , \6973_b0 );
or ( \6978_b1 , \6977_b1 , \6974_b1 );
not ( \6974_b1 , w_22282 );
and ( \6978_b0 , \6977_b0 , w_22283 );
and ( w_22282 , w_22283 , \6974_b0 );
or ( \6979_b1 , \6976_b1 , w_22285 );
not ( w_22285 , w_22286 );
and ( \6979_b0 , \6976_b0 , w_22287 );
and ( w_22286 ,  , w_22287 );
buf ( w_22285 , \6978_b1 );
not ( w_22285 , w_22288 );
not (  , w_22289 );
and ( w_22288 , w_22289 , \6978_b0 );
or ( \6980_b1 , \4836_b1 , \4885_b1 );
not ( \4885_b1 , w_22290 );
and ( \6980_b0 , \4836_b0 , w_22291 );
and ( w_22290 , w_22291 , \4885_b0 );
buf ( \6981_b1 , \6980_b1 );
not ( \6981_b1 , w_22292 );
not ( \6981_b0 , w_22293 );
and ( w_22292 , w_22293 , \6980_b0 );
buf ( \6982_b1 , \6904_b1 );
not ( \6982_b1 , w_22294 );
not ( \6982_b0 , w_22295 );
and ( w_22294 , w_22295 , \6904_b0 );
or ( \6983_b1 , \6981_b1 , w_22296 );
or ( \6983_b0 , \6981_b0 , \6982_b0 );
not ( \6982_b0 , w_22297 );
and ( w_22297 , w_22296 , \6982_b1 );
buf ( \6984_b1 , \6921_b1 );
not ( \6984_b1 , w_22298 );
not ( \6984_b0 , w_22299 );
and ( w_22298 , w_22299 , \6921_b0 );
or ( \6985_b1 , \6983_b1 , w_22301 );
not ( w_22301 , w_22302 );
and ( \6985_b0 , \6983_b0 , w_22303 );
and ( w_22302 ,  , w_22303 );
buf ( w_22301 , \6984_b1 );
not ( w_22301 , w_22304 );
not (  , w_22305 );
and ( w_22304 , w_22305 , \6984_b0 );
or ( \6986_b1 , \6924_b1 , w_22307 );
not ( w_22307 , w_22308 );
and ( \6986_b0 , \6924_b0 , w_22309 );
and ( w_22308 ,  , w_22309 );
buf ( w_22307 , \4927_b1 );
not ( w_22307 , w_22310 );
not (  , w_22311 );
and ( w_22310 , w_22311 , \4927_b0 );
buf ( \6987_b1 , \6986_b1 );
not ( \6987_b1 , w_22312 );
not ( \6987_b0 , w_22313 );
and ( w_22312 , w_22313 , \6986_b0 );
or ( \6988_b1 , \6985_b1 , \6987_b1 );
not ( \6987_b1 , w_22314 );
and ( \6988_b0 , \6985_b0 , w_22315 );
and ( w_22314 , w_22315 , \6987_b0 );
buf ( \6989_b1 , \6985_b1 );
not ( \6989_b1 , w_22316 );
not ( \6989_b0 , w_22317 );
and ( w_22316 , w_22317 , \6985_b0 );
or ( \6990_b1 , \6989_b1 , \6986_b1 );
not ( \6986_b1 , w_22318 );
and ( \6990_b0 , \6989_b0 , w_22319 );
and ( w_22318 , w_22319 , \6986_b0 );
or ( \6991_b1 , \6988_b1 , w_22321 );
not ( w_22321 , w_22322 );
and ( \6991_b0 , \6988_b0 , w_22323 );
and ( w_22322 ,  , w_22323 );
buf ( w_22321 , \6990_b1 );
not ( w_22321 , w_22324 );
not (  , w_22325 );
and ( w_22324 , w_22325 , \6990_b0 );
buf ( \6992_b1 , \4836_b1 );
not ( \6992_b1 , w_22326 );
not ( \6992_b0 , w_22327 );
and ( w_22326 , w_22327 , \4836_b0 );
buf ( \6993_b1 , \6904_b1 );
not ( \6993_b1 , w_22328 );
not ( \6993_b0 , w_22329 );
and ( w_22328 , w_22329 , \6904_b0 );
or ( \6994_b1 , \6992_b1 , w_22330 );
or ( \6994_b0 , \6992_b0 , \6993_b0 );
not ( \6993_b0 , w_22331 );
and ( w_22331 , w_22330 , \6993_b1 );
or ( \6995_b1 , \6912_b1 , w_22333 );
not ( w_22333 , w_22334 );
and ( \6995_b0 , \6912_b0 , w_22335 );
and ( w_22334 ,  , w_22335 );
buf ( w_22333 , \6913_b1 );
not ( w_22333 , w_22336 );
not (  , w_22337 );
and ( w_22336 , w_22337 , \6913_b0 );
buf ( \6996_b1 , \4835_b1 );
not ( \6996_b1 , w_22338 );
not ( \6996_b0 , w_22339 );
and ( w_22338 , w_22339 , \4835_b0 );
or ( \6997_b1 , \6995_b1 , \6996_b1 );
not ( \6996_b1 , w_22340 );
and ( \6997_b0 , \6995_b0 , w_22341 );
and ( w_22340 , w_22341 , \6996_b0 );
buf ( \6998_b1 , \6914_b1 );
not ( \6998_b1 , w_22342 );
not ( \6998_b0 , w_22343 );
and ( w_22342 , w_22343 , \6914_b0 );
or ( \6999_b1 , \6997_b1 , w_22345 );
not ( w_22345 , w_22346 );
and ( \6999_b0 , \6997_b0 , w_22347 );
and ( w_22346 ,  , w_22347 );
buf ( w_22345 , \6998_b1 );
not ( w_22345 , w_22348 );
not (  , w_22349 );
and ( w_22348 , w_22349 , \6998_b0 );
or ( \7000_b1 , \6994_b1 , w_22351 );
not ( w_22351 , w_22352 );
and ( \7000_b0 , \6994_b0 , w_22353 );
and ( w_22352 ,  , w_22353 );
buf ( w_22351 , \6999_b1 );
not ( w_22351 , w_22354 );
not (  , w_22355 );
and ( w_22354 , w_22355 , \6999_b0 );
buf ( \7001_b1 , \6919_b1 );
not ( \7001_b1 , w_22356 );
not ( \7001_b0 , w_22357 );
and ( w_22356 , w_22357 , \6919_b0 );
or ( \7002_b1 , \7001_b1 , w_22359 );
not ( w_22359 , w_22360 );
and ( \7002_b0 , \7001_b0 , w_22361 );
and ( w_22360 ,  , w_22361 );
buf ( w_22359 , \4885_b1 );
not ( w_22359 , w_22362 );
not (  , w_22363 );
and ( w_22362 , w_22363 , \4885_b0 );
buf ( \7003_b1 , \7002_b1 );
not ( \7003_b1 , w_22364 );
not ( \7003_b0 , w_22365 );
and ( w_22364 , w_22365 , \7002_b0 );
or ( \7004_b1 , \7000_b1 , \7003_b1 );
not ( \7003_b1 , w_22366 );
and ( \7004_b0 , \7000_b0 , w_22367 );
and ( w_22366 , w_22367 , \7003_b0 );
buf ( \7005_b1 , \7000_b1 );
not ( \7005_b1 , w_22368 );
not ( \7005_b0 , w_22369 );
and ( w_22368 , w_22369 , \7000_b0 );
or ( \7006_b1 , \7005_b1 , \7002_b1 );
not ( \7002_b1 , w_22370 );
and ( \7006_b0 , \7005_b0 , w_22371 );
and ( w_22370 , w_22371 , \7002_b0 );
or ( \7007_b1 , \7004_b1 , w_22373 );
not ( w_22373 , w_22374 );
and ( \7007_b0 , \7004_b0 , w_22375 );
and ( w_22374 ,  , w_22375 );
buf ( w_22373 , \7006_b1 );
not ( w_22373 , w_22376 );
not (  , w_22377 );
and ( w_22376 , w_22377 , \7006_b0 );
buf ( \7008_b1 , \4767_b1 );
not ( \7008_b1 , w_22378 );
not ( \7008_b0 , w_22379 );
and ( w_22378 , w_22379 , \4767_b0 );
buf ( \7009_b1 , \7008_b1 );
not ( \7009_b1 , w_22380 );
not ( \7009_b0 , w_22381 );
and ( w_22380 , w_22381 , \7008_b0 );
buf ( \7010_b1 , \6904_b1 );
not ( \7010_b1 , w_22382 );
not ( \7010_b0 , w_22383 );
and ( w_22382 , w_22383 , \6904_b0 );
or ( \7011_b1 , \7009_b1 , w_22384 );
or ( \7011_b0 , \7009_b0 , \7010_b0 );
not ( \7010_b0 , w_22385 );
and ( w_22385 , w_22384 , \7010_b1 );
buf ( \7012_b1 , \6995_b1 );
not ( \7012_b1 , w_22386 );
not ( \7012_b0 , w_22387 );
and ( w_22386 , w_22387 , \6995_b0 );
or ( \7013_b1 , \7011_b1 , w_22389 );
not ( w_22389 , w_22390 );
and ( \7013_b0 , \7011_b0 , w_22391 );
and ( w_22390 ,  , w_22391 );
buf ( w_22389 , \7012_b1 );
not ( w_22389 , w_22392 );
not (  , w_22393 );
and ( w_22392 , w_22393 , \7012_b0 );
buf ( \7014_b1 , \6998_b1 );
not ( \7014_b1 , w_22394 );
not ( \7014_b0 , w_22395 );
and ( w_22394 , w_22395 , \6998_b0 );
or ( \7015_b1 , \7014_b1 , w_22397 );
not ( w_22397 , w_22398 );
and ( \7015_b0 , \7014_b0 , w_22399 );
and ( w_22398 ,  , w_22399 );
buf ( w_22397 , \4834_b1 );
not ( w_22397 , w_22400 );
not (  , w_22401 );
and ( w_22400 , w_22401 , \4834_b0 );
buf ( \7016_b1 , \7015_b1 );
not ( \7016_b1 , w_22402 );
not ( \7016_b0 , w_22403 );
and ( w_22402 , w_22403 , \7015_b0 );
or ( \7017_b1 , \7013_b1 , \7016_b1 );
not ( \7016_b1 , w_22404 );
and ( \7017_b0 , \7013_b0 , w_22405 );
and ( w_22404 , w_22405 , \7016_b0 );
buf ( \7018_b1 , \7013_b1 );
not ( \7018_b1 , w_22406 );
not ( \7018_b0 , w_22407 );
and ( w_22406 , w_22407 , \7013_b0 );
or ( \7019_b1 , \7018_b1 , \7015_b1 );
not ( \7015_b1 , w_22408 );
and ( \7019_b0 , \7018_b0 , w_22409 );
and ( w_22408 , w_22409 , \7015_b0 );
or ( \7020_b1 , \7017_b1 , w_22411 );
not ( w_22411 , w_22412 );
and ( \7020_b0 , \7017_b0 , w_22413 );
and ( w_22412 ,  , w_22413 );
buf ( w_22411 , \7019_b1 );
not ( w_22411 , w_22414 );
not (  , w_22415 );
and ( w_22414 , w_22415 , \7019_b0 );
buf ( \7021_b1 , \4694_b1 );
not ( \7021_b1 , w_22416 );
not ( \7021_b0 , w_22417 );
and ( w_22416 , w_22417 , \4694_b0 );
buf ( \7022_b1 , \6904_b1 );
not ( \7022_b1 , w_22418 );
not ( \7022_b0 , w_22419 );
and ( w_22418 , w_22419 , \6904_b0 );
or ( \7023_b1 , \7021_b1 , w_22420 );
or ( \7023_b0 , \7021_b0 , \7022_b0 );
not ( \7022_b0 , w_22421 );
and ( w_22421 , w_22420 , \7022_b1 );
or ( \7024_b1 , \7023_b1 , w_22423 );
not ( w_22423 , w_22424 );
and ( \7024_b0 , \7023_b0 , w_22425 );
and ( w_22424 ,  , w_22425 );
buf ( w_22423 , \6910_b1 );
not ( w_22423 , w_22426 );
not (  , w_22427 );
and ( w_22426 , w_22427 , \6910_b0 );
or ( \7025_b1 , \6913_b1 , w_22429 );
not ( w_22429 , w_22430 );
and ( \7025_b0 , \6913_b0 , w_22431 );
and ( w_22430 ,  , w_22431 );
buf ( w_22429 , \4766_b1 );
not ( w_22429 , w_22432 );
not (  , w_22433 );
and ( w_22432 , w_22433 , \4766_b0 );
buf ( \7026_b1 , \7025_b1 );
not ( \7026_b1 , w_22434 );
not ( \7026_b0 , w_22435 );
and ( w_22434 , w_22435 , \7025_b0 );
or ( \7027_b1 , \7024_b1 , \7026_b1 );
not ( \7026_b1 , w_22436 );
and ( \7027_b0 , \7024_b0 , w_22437 );
and ( w_22436 , w_22437 , \7026_b0 );
buf ( \7028_b1 , \7024_b1 );
not ( \7028_b1 , w_22438 );
not ( \7028_b0 , w_22439 );
and ( w_22438 , w_22439 , \7024_b0 );
or ( \7029_b1 , \7028_b1 , \7025_b1 );
not ( \7025_b1 , w_22440 );
and ( \7029_b0 , \7028_b0 , w_22441 );
and ( w_22440 , w_22441 , \7025_b0 );
or ( \7030_b1 , \7027_b1 , w_22443 );
not ( w_22443 , w_22444 );
and ( \7030_b0 , \7027_b0 , w_22445 );
and ( w_22444 ,  , w_22445 );
buf ( w_22443 , \7029_b1 );
not ( w_22443 , w_22446 );
not (  , w_22447 );
and ( w_22446 , w_22447 , \7029_b0 );
buf ( \7031_b1 , \5543_b1 );
not ( \7031_b1 , w_22448 );
not ( \7031_b0 , w_22449 );
and ( w_22448 , w_22449 , \5543_b0 );
buf ( \7032_b1 , \5511_b1 );
not ( \7032_b1 , w_22450 );
not ( \7032_b0 , w_22451 );
and ( w_22450 , w_22451 , \5511_b0 );
buf ( \7033_b1 , \6888_b1 );
not ( \7033_b1 , w_22452 );
not ( \7033_b0 , w_22453 );
and ( w_22452 , w_22453 , \6888_b0 );
or ( \7034_b1 , \7032_b1 , w_22454 );
or ( \7034_b0 , \7032_b0 , \7033_b0 );
not ( \7033_b0 , w_22455 );
and ( w_22455 , w_22454 , \7033_b1 );
buf ( \7035_b1 , \6894_b1 );
not ( \7035_b1 , w_22456 );
not ( \7035_b0 , w_22457 );
and ( w_22456 , w_22457 , \6894_b0 );
or ( \7036_b1 , \6893_b1 , w_22459 );
not ( w_22459 , w_22460 );
and ( \7036_b0 , \6893_b0 , w_22461 );
and ( w_22460 ,  , w_22461 );
buf ( w_22459 , \7035_b1 );
not ( w_22459 , w_22462 );
not (  , w_22463 );
and ( w_22462 , w_22463 , \7035_b0 );
or ( \7037_b1 , \7034_b1 , w_22465 );
not ( w_22465 , w_22466 );
and ( \7037_b0 , \7034_b0 , w_22467 );
and ( w_22466 ,  , w_22467 );
buf ( w_22465 , \7036_b1 );
not ( w_22465 , w_22468 );
not (  , w_22469 );
and ( w_22468 , w_22469 , \7036_b0 );
buf ( \7038_b1 , \7037_b1 );
not ( \7038_b1 , w_22470 );
not ( \7038_b0 , w_22471 );
and ( w_22470 , w_22471 , \7037_b0 );
or ( \7039_b1 , \7031_b1 , w_22472 );
or ( \7039_b0 , \7031_b0 , \7038_b0 );
not ( \7038_b0 , w_22473 );
and ( w_22473 , w_22472 , \7038_b1 );
or ( \7040_b1 , \7039_b1 , w_22475 );
not ( w_22475 , w_22476 );
and ( \7040_b0 , \7039_b0 , w_22477 );
and ( w_22476 ,  , w_22477 );
buf ( w_22475 , \6897_b1 );
not ( w_22475 , w_22478 );
not (  , w_22479 );
and ( w_22478 , w_22479 , \6897_b0 );
or ( \7041_b1 , \6901_b1 , w_22481 );
not ( w_22481 , w_22482 );
and ( \7041_b0 , \6901_b0 , w_22483 );
and ( w_22482 ,  , w_22483 );
buf ( w_22481 , \5557_b1 );
not ( w_22481 , w_22484 );
not (  , w_22485 );
and ( w_22484 , w_22485 , \5557_b0 );
buf ( \7042_b1 , \7041_b1 );
not ( \7042_b1 , w_22486 );
not ( \7042_b0 , w_22487 );
and ( w_22486 , w_22487 , \7041_b0 );
or ( \7043_b1 , \7040_b1 , \7042_b1 );
not ( \7042_b1 , w_22488 );
and ( \7043_b0 , \7040_b0 , w_22489 );
and ( w_22488 , w_22489 , \7042_b0 );
buf ( \7044_b1 , \7040_b1 );
not ( \7044_b1 , w_22490 );
not ( \7044_b0 , w_22491 );
and ( w_22490 , w_22491 , \7040_b0 );
or ( \7045_b1 , \7044_b1 , \7041_b1 );
not ( \7041_b1 , w_22492 );
and ( \7045_b0 , \7044_b0 , w_22493 );
and ( w_22492 , w_22493 , \7041_b0 );
or ( \7046_b1 , \7043_b1 , w_22495 );
not ( w_22495 , w_22496 );
and ( \7046_b0 , \7043_b0 , w_22497 );
and ( w_22496 ,  , w_22497 );
buf ( w_22495 , \7045_b1 );
not ( w_22495 , w_22498 );
not (  , w_22499 );
and ( w_22498 , w_22499 , \7045_b0 );
buf ( \7047_b1 , \4927_b1 );
not ( \7047_b1 , w_22500 );
not ( \7047_b0 , w_22501 );
and ( w_22500 , w_22501 , \4927_b0 );
or ( \7048_b1 , \7047_b1 , w_22503 );
not ( w_22503 , w_22504 );
and ( \7048_b0 , \7047_b0 , w_22505 );
and ( w_22504 ,  , w_22505 );
buf ( w_22503 , \4960_b1 );
not ( w_22503 , w_22506 );
not (  , w_22507 );
and ( w_22506 , w_22507 , \4960_b0 );
or ( \7049_b1 , \6980_b1 , \7048_b1 );
not ( \7048_b1 , w_22508 );
and ( \7049_b0 , \6980_b0 , w_22509 );
and ( w_22508 , w_22509 , \7048_b0 );
buf ( \7050_b1 , \6888_b1 );
buf ( \7050_b0 , \6888_b0 );
buf ( \7052_b1 , \6903_b1 );
not ( \7052_b1 , w_22510 );
not ( \7052_b0 , w_22511 );
and ( w_22510 , w_22511 , \6903_b0 );
or ( \7053_b1 , \7052_b1 , w_22513 );
not ( w_22513 , w_22514 );
and ( \7053_b0 , \7052_b0 , w_22515 );
and ( w_22514 ,  , w_22515 );
buf ( w_22513 , \7049_b1 );
not ( w_22513 , w_22516 );
not (  , w_22517 );
and ( w_22516 , w_22517 , \7049_b0 );
buf ( \7054_b1 , \6929_b1 );
not ( \7054_b1 , w_22518 );
not ( \7054_b0 , w_22519 );
and ( w_22518 , w_22519 , \6929_b0 );
or ( \7056_b1 , \6932_b1 , w_22521 );
not ( w_22521 , w_22522 );
and ( \7056_b0 , \6932_b0 , w_22523 );
and ( w_22522 ,  , w_22523 );
buf ( w_22521 , \4983_b1 );
not ( w_22521 , w_22524 );
not (  , w_22525 );
and ( w_22524 , w_22525 , \4983_b0 );
or ( \7057_b1 , \7055_b1 , \7056_b1 );
not ( \7056_b1 , w_22526 );
and ( \7057_b0 , \7055_b0 , w_22527 );
and ( w_22526 , w_22527 , \7056_b0 );
buf ( \7058_b1 , \7055_b1 );
not ( \7058_b1 , w_22528 );
not ( \7058_b0 , w_22529 );
and ( w_22528 , w_22529 , \7055_b0 );
buf ( \7059_b1 , \7056_b1 );
not ( \7059_b1 , w_22530 );
not ( \7059_b0 , w_22531 );
and ( w_22530 , w_22531 , \7056_b0 );
or ( \7060_b1 , \7058_b1 , \7059_b1 );
not ( \7059_b1 , w_22532 );
and ( \7060_b0 , \7058_b0 , w_22533 );
and ( w_22532 , w_22533 , \7059_b0 );
or ( \7061_b1 , \7057_b1 , w_22535 );
not ( w_22535 , w_22536 );
and ( \7061_b0 , \7057_b0 , w_22537 );
and ( w_22536 ,  , w_22537 );
buf ( w_22535 , \7060_b1 );
not ( w_22535 , w_22538 );
not (  , w_22539 );
and ( w_22538 , w_22539 , \7060_b0 );
buf ( \7062_b1 , \5510_b1 );
buf ( \7062_b0 , \5510_b0 );
buf ( \7063_b1 , \7062_b1 );
not ( \7063_b1 , w_22540 );
not ( \7063_b0 , w_22541 );
and ( w_22540 , w_22541 , \7062_b0 );
buf ( \7064_b1 , \7050_b1 );
not ( \7064_b1 , w_22542 );
not ( \7064_b0 , w_22543 );
and ( w_22542 , w_22543 , \7050_b0 );
or ( \7065_b1 , \7063_b1 , w_22544 );
or ( \7065_b0 , \7063_b0 , \7064_b0 );
not ( \7064_b0 , w_22545 );
and ( w_22545 , w_22544 , \7064_b1 );
or ( \7066_b1 , \7065_b1 , w_22547 );
not ( w_22547 , w_22548 );
and ( \7066_b0 , \7065_b0 , w_22549 );
and ( w_22548 ,  , w_22549 );
buf ( w_22547 , \6892_b1 );
not ( w_22547 , w_22550 );
not (  , w_22551 );
and ( w_22550 , w_22551 , \6892_b0 );
or ( \7067_b1 , \7035_b1 , w_22553 );
not ( w_22553 , w_22554 );
and ( \7067_b0 , \7035_b0 , w_22555 );
and ( w_22554 ,  , w_22555 );
buf ( w_22553 , \6891_b1 );
not ( w_22553 , w_22556 );
not (  , w_22557 );
and ( w_22556 , w_22557 , \6891_b0 );
buf ( \7068_b1 , \7067_b1 );
not ( \7068_b1 , w_22558 );
not ( \7068_b0 , w_22559 );
and ( w_22558 , w_22559 , \7067_b0 );
or ( \7069_b1 , \7066_b1 , \7068_b1 );
not ( \7068_b1 , w_22560 );
and ( \7069_b0 , \7066_b0 , w_22561 );
and ( w_22560 , w_22561 , \7068_b0 );
buf ( \7070_b1 , \7066_b1 );
not ( \7070_b1 , w_22562 );
not ( \7070_b0 , w_22563 );
and ( w_22562 , w_22563 , \7066_b0 );
or ( \7071_b1 , \7070_b1 , \7067_b1 );
not ( \7067_b1 , w_22564 );
and ( \7071_b0 , \7070_b0 , w_22565 );
and ( w_22564 , w_22565 , \7067_b0 );
or ( \7072_b1 , \7069_b1 , w_22567 );
not ( w_22567 , w_22568 );
and ( \7072_b0 , \7069_b0 , w_22569 );
and ( w_22568 ,  , w_22569 );
buf ( w_22567 , \7071_b1 );
not ( w_22567 , w_22570 );
not (  , w_22571 );
and ( w_22570 , w_22571 , \7071_b0 );
or ( \7073_b1 , \6892_b1 , w_22573 );
not ( w_22573 , w_22574 );
and ( \7073_b0 , \6892_b0 , w_22575 );
and ( w_22574 ,  , w_22575 );
buf ( w_22573 , \7062_b1 );
not ( w_22573 , w_22576 );
not (  , w_22577 );
and ( w_22576 , w_22577 , \7062_b0 );
buf ( \7074_b1 , \7073_b1 );
not ( \7074_b1 , w_22578 );
not ( \7074_b0 , w_22579 );
and ( w_22578 , w_22579 , \7073_b0 );
or ( \7075_b1 , \7050_b1 , \7074_b1 );
not ( \7074_b1 , w_22580 );
and ( \7075_b0 , \7050_b0 , w_22581 );
and ( w_22580 , w_22581 , \7074_b0 );
buf ( \7076_b1 , \7050_b1 );
not ( \7076_b1 , w_22582 );
not ( \7076_b0 , w_22583 );
and ( w_22582 , w_22583 , \7050_b0 );
or ( \7077_b1 , \7076_b1 , \7073_b1 );
not ( \7073_b1 , w_22584 );
and ( \7077_b0 , \7076_b0 , w_22585 );
and ( w_22584 , w_22585 , \7073_b0 );
or ( \7078_b1 , \7075_b1 , w_22587 );
not ( w_22587 , w_22588 );
and ( \7078_b0 , \7075_b0 , w_22589 );
and ( w_22588 ,  , w_22589 );
buf ( w_22587 , \7077_b1 );
not ( w_22587 , w_22590 );
not (  , w_22591 );
and ( w_22590 , w_22591 , \7077_b0 );
buf ( \7079_b1 , \6886_b1 );
not ( \7079_b1 , w_22592 );
not ( \7079_b0 , w_22593 );
and ( w_22592 , w_22593 , \6886_b0 );
or ( \7080_b1 , \7079_b1 , w_22595 );
not ( w_22595 , w_22596 );
and ( \7080_b0 , \7079_b0 , w_22597 );
and ( w_22596 ,  , w_22597 );
buf ( w_22595 , \6883_b1 );
not ( w_22595 , w_22598 );
not (  , w_22599 );
and ( w_22598 , w_22599 , \6883_b0 );
buf ( \7081_b1 , \6831_b1 );
buf ( \7081_b0 , \6831_b0 );
buf ( \7082_b1 , \7081_b1 );
not ( \7082_b1 , w_22600 );
not ( \7082_b0 , w_22601 );
and ( w_22600 , w_22601 , \7081_b0 );
buf ( \7083_b1 , \6876_b1 );
not ( \7083_b1 , w_22602 );
not ( \7083_b0 , w_22603 );
and ( w_22602 , w_22603 , \6876_b0 );
or ( \7084_b1 , \7082_b1 , w_22604 );
or ( \7084_b0 , \7082_b0 , \7083_b0 );
not ( \7083_b0 , w_22605 );
and ( w_22605 , w_22604 , \7083_b1 );
buf ( \7085_b1 , \6881_b1 );
not ( \7085_b1 , w_22606 );
not ( \7085_b0 , w_22607 );
and ( w_22606 , w_22607 , \6881_b0 );
or ( \7086_b1 , \7084_b1 , w_22609 );
not ( w_22609 , w_22610 );
and ( \7086_b0 , \7084_b0 , w_22611 );
and ( w_22610 ,  , w_22611 );
buf ( w_22609 , \7085_b1 );
not ( w_22609 , w_22612 );
not (  , w_22613 );
and ( w_22612 , w_22613 , \7085_b0 );
buf ( \7087_b1 , \5744_b1 );
buf ( \7087_b0 , \5744_b0 );
or ( \7088_b1 , \7086_b1 , \7087_b1 );
not ( \7087_b1 , w_22614 );
and ( \7088_b0 , \7086_b0 , w_22615 );
and ( w_22614 , w_22615 , \7087_b0 );
buf ( \7089_b1 , \6884_b1 );
buf ( \7089_b0 , \6884_b0 );
or ( \7090_b1 , \7088_b1 , w_22617 );
not ( w_22617 , w_22618 );
and ( \7090_b0 , \7088_b0 , w_22619 );
and ( w_22618 ,  , w_22619 );
buf ( w_22617 , \7089_b1 );
not ( w_22617 , w_22620 );
not (  , w_22621 );
and ( w_22620 , w_22621 , \7089_b0 );
or ( \7091_b1 , \7080_b1 , \7090_b1 );
not ( \7090_b1 , w_22622 );
and ( \7091_b0 , \7080_b0 , w_22623 );
and ( w_22622 , w_22623 , \7090_b0 );
buf ( \7092_b1 , \7080_b1 );
not ( \7092_b1 , w_22624 );
not ( \7092_b0 , w_22625 );
and ( w_22624 , w_22625 , \7080_b0 );
buf ( \7093_b1 , \7090_b1 );
not ( \7093_b1 , w_22626 );
not ( \7093_b0 , w_22627 );
and ( w_22626 , w_22627 , \7090_b0 );
or ( \7094_b1 , \7092_b1 , \7093_b1 );
not ( \7093_b1 , w_22628 );
and ( \7094_b0 , \7092_b0 , w_22629 );
and ( w_22628 , w_22629 , \7093_b0 );
or ( \7095_b1 , \7091_b1 , w_22631 );
not ( w_22631 , w_22632 );
and ( \7095_b0 , \7091_b0 , w_22633 );
and ( w_22632 ,  , w_22633 );
buf ( w_22631 , \7094_b1 );
not ( w_22631 , w_22634 );
not (  , w_22635 );
and ( w_22634 , w_22635 , \7094_b0 );
buf ( \7096_b1 , \7087_b1 );
not ( \7096_b1 , w_22636 );
not ( \7096_b0 , w_22637 );
and ( w_22636 , w_22637 , \7087_b0 );
or ( \7097_b1 , \7096_b1 , w_22639 );
not ( w_22639 , w_22640 );
and ( \7097_b0 , \7096_b0 , w_22641 );
and ( w_22640 ,  , w_22641 );
buf ( w_22639 , \7089_b1 );
not ( w_22639 , w_22642 );
not (  , w_22643 );
and ( w_22642 , w_22643 , \7089_b0 );
or ( \7098_b1 , \7097_b1 , \7086_b1 );
not ( \7086_b1 , w_22644 );
and ( \7098_b0 , \7097_b0 , w_22645 );
and ( w_22644 , w_22645 , \7086_b0 );
buf ( \7099_b1 , \7097_b1 );
not ( \7099_b1 , w_22646 );
not ( \7099_b0 , w_22647 );
and ( w_22646 , w_22647 , \7097_b0 );
buf ( \7100_b1 , \7086_b1 );
not ( \7100_b1 , w_22648 );
not ( \7100_b0 , w_22649 );
and ( w_22648 , w_22649 , \7086_b0 );
or ( \7101_b1 , \7099_b1 , \7100_b1 );
not ( \7100_b1 , w_22650 );
and ( \7101_b0 , \7099_b0 , w_22651 );
and ( w_22650 , w_22651 , \7100_b0 );
or ( \7102_b1 , \7098_b1 , w_22653 );
not ( w_22653 , w_22654 );
and ( \7102_b0 , \7098_b0 , w_22655 );
and ( w_22654 ,  , w_22655 );
buf ( w_22653 , \7101_b1 );
not ( w_22653 , w_22656 );
not (  , w_22657 );
and ( w_22656 , w_22657 , \7101_b0 );
buf ( \7103_b1 , \6875_b1 );
not ( \7103_b1 , w_22658 );
not ( \7103_b0 , w_22659 );
and ( w_22658 , w_22659 , \6875_b0 );
buf ( \7104_b1 , \7081_b1 );
not ( \7104_b1 , w_22660 );
not ( \7104_b0 , w_22661 );
and ( w_22660 , w_22661 , \7081_b0 );
or ( \7105_b1 , \7103_b1 , w_22662 );
or ( \7105_b0 , \7103_b0 , \7104_b0 );
not ( \7104_b0 , w_22663 );
and ( w_22663 , w_22662 , \7104_b1 );
or ( \7106_b1 , \7105_b1 , w_22665 );
not ( w_22665 , w_22666 );
and ( \7106_b0 , \7105_b0 , w_22667 );
and ( w_22666 ,  , w_22667 );
buf ( w_22665 , \6879_b1 );
not ( w_22665 , w_22668 );
not (  , w_22669 );
and ( w_22668 , w_22669 , \6879_b0 );
or ( \7107_b1 , \6878_b1 , w_22671 );
not ( w_22671 , w_22672 );
and ( \7107_b0 , \6878_b0 , w_22673 );
and ( w_22672 ,  , w_22673 );
buf ( w_22671 , \6861_b1 );
not ( w_22671 , w_22674 );
not (  , w_22675 );
and ( w_22674 , w_22675 , \6861_b0 );
buf ( \7108_b1 , \7107_b1 );
not ( \7108_b1 , w_22676 );
not ( \7108_b0 , w_22677 );
and ( w_22676 , w_22677 , \7107_b0 );
or ( \7109_b1 , \7106_b1 , \7108_b1 );
not ( \7108_b1 , w_22678 );
and ( \7109_b0 , \7106_b0 , w_22679 );
and ( w_22678 , w_22679 , \7108_b0 );
buf ( \7110_b1 , \7106_b1 );
not ( \7110_b1 , w_22680 );
not ( \7110_b0 , w_22681 );
and ( w_22680 , w_22681 , \7106_b0 );
or ( \7111_b1 , \7110_b1 , \7107_b1 );
not ( \7107_b1 , w_22682 );
and ( \7111_b0 , \7110_b0 , w_22683 );
and ( w_22682 , w_22683 , \7107_b0 );
or ( \7112_b1 , \7109_b1 , w_22685 );
not ( w_22685 , w_22686 );
and ( \7112_b0 , \7109_b0 , w_22687 );
and ( w_22686 ,  , w_22687 );
buf ( w_22685 , \7111_b1 );
not ( w_22685 , w_22688 );
not (  , w_22689 );
and ( w_22688 , w_22689 , \7111_b0 );
or ( \7113_b1 , \6875_b1 , w_22691 );
not ( w_22691 , w_22692 );
and ( \7113_b0 , \6875_b0 , w_22693 );
and ( w_22692 ,  , w_22693 );
buf ( w_22691 , \6879_b1 );
not ( w_22691 , w_22694 );
not (  , w_22695 );
and ( w_22694 , w_22695 , \6879_b0 );
buf ( \7114_b1 , \7113_b1 );
not ( \7114_b1 , w_22696 );
not ( \7114_b0 , w_22697 );
and ( w_22696 , w_22697 , \7113_b0 );
or ( \7115_b1 , \7081_b1 , \7114_b1 );
not ( \7114_b1 , w_22698 );
and ( \7115_b0 , \7081_b0 , w_22699 );
and ( w_22698 , w_22699 , \7114_b0 );
buf ( \7116_b1 , \7081_b1 );
not ( \7116_b1 , w_22700 );
not ( \7116_b0 , w_22701 );
and ( w_22700 , w_22701 , \7081_b0 );
or ( \7117_b1 , \7116_b1 , \7113_b1 );
not ( \7113_b1 , w_22702 );
and ( \7117_b0 , \7116_b0 , w_22703 );
and ( w_22702 , w_22703 , \7113_b0 );
or ( \7118_b1 , \7115_b1 , w_22705 );
not ( w_22705 , w_22706 );
and ( \7118_b0 , \7115_b0 , w_22707 );
and ( w_22706 ,  , w_22707 );
buf ( w_22705 , \7117_b1 );
not ( w_22705 , w_22708 );
not (  , w_22709 );
and ( w_22708 , w_22709 , \7117_b0 );
buf ( \7119_b1 , \6812_b1 );
not ( \7119_b1 , w_22710 );
not ( \7119_b0 , w_22711 );
and ( w_22710 , w_22711 , \6812_b0 );
buf ( \7120_b1 , \6769_b1 );
not ( \7120_b1 , w_22712 );
not ( \7120_b0 , w_22713 );
and ( w_22712 , w_22713 , \6769_b0 );
or ( \7121_b1 , \7119_b1 , w_22714 );
or ( \7121_b0 , \7119_b0 , \7120_b0 );
not ( \7120_b0 , w_22715 );
and ( w_22715 , w_22714 , \7120_b1 );
or ( \7122_b1 , \7121_b1 , w_22717 );
not ( w_22717 , w_22718 );
and ( \7122_b0 , \7121_b0 , w_22719 );
and ( w_22718 ,  , w_22719 );
buf ( w_22717 , \6828_b1 );
not ( w_22717 , w_22720 );
not (  , w_22721 );
and ( w_22720 , w_22721 , \6828_b0 );
buf ( \7123_b1 , \6196_b1 );
buf ( \7123_b0 , \6196_b0 );
or ( \7124_b1 , \7122_b1 , \7123_b1 );
not ( \7123_b1 , w_22722 );
and ( \7124_b0 , \7122_b0 , w_22723 );
and ( w_22722 , w_22723 , \7123_b0 );
buf ( \7125_b1 , \6822_b1 );
not ( \7125_b1 , w_22724 );
not ( \7125_b0 , w_22725 );
and ( w_22724 , w_22725 , \6822_b0 );
or ( \7126_b1 , \7124_b1 , w_22727 );
not ( w_22727 , w_22728 );
and ( \7126_b0 , \7124_b0 , w_22729 );
and ( w_22728 ,  , w_22729 );
buf ( w_22727 , \7125_b1 );
not ( w_22727 , w_22730 );
not (  , w_22731 );
and ( w_22730 , w_22731 , \7125_b0 );
or ( \7127_b1 , \6127_b1 , w_22733 );
not ( w_22733 , w_22734 );
and ( \7127_b0 , \6127_b0 , w_22735 );
and ( w_22734 ,  , w_22735 );
buf ( w_22733 , \6816_b1 );
not ( w_22733 , w_22736 );
not (  , w_22737 );
and ( w_22736 , w_22737 , \6816_b0 );
or ( \7128_b1 , \7126_b1 , \7127_b1 );
not ( \7127_b1 , w_22738 );
and ( \7128_b0 , \7126_b0 , w_22739 );
and ( w_22738 , w_22739 , \7127_b0 );
buf ( \7129_b1 , \7126_b1 );
not ( \7129_b1 , w_22740 );
not ( \7129_b0 , w_22741 );
and ( w_22740 , w_22741 , \7126_b0 );
buf ( \7130_b1 , \7127_b1 );
not ( \7130_b1 , w_22742 );
not ( \7130_b0 , w_22743 );
and ( w_22742 , w_22743 , \7127_b0 );
or ( \7131_b1 , \7129_b1 , \7130_b1 );
not ( \7130_b1 , w_22744 );
and ( \7131_b0 , \7129_b0 , w_22745 );
and ( w_22744 , w_22745 , \7130_b0 );
or ( \7132_b1 , \7128_b1 , w_22747 );
not ( w_22747 , w_22748 );
and ( \7132_b0 , \7128_b0 , w_22749 );
and ( w_22748 ,  , w_22749 );
buf ( w_22747 , \7131_b1 );
not ( w_22747 , w_22750 );
not (  , w_22751 );
and ( w_22750 , w_22751 , \7131_b0 );
or ( \7133_b1 , \6822_b1 , w_22753 );
not ( w_22753 , w_22754 );
and ( \7133_b0 , \6822_b0 , w_22755 );
and ( w_22754 ,  , w_22755 );
buf ( w_22753 , \7123_b1 );
not ( w_22753 , w_22756 );
not (  , w_22757 );
and ( w_22756 , w_22757 , \7123_b0 );
buf ( \7134_b1 , \7133_b1 );
not ( \7134_b1 , w_22758 );
not ( \7134_b0 , w_22759 );
and ( w_22758 , w_22759 , \7133_b0 );
or ( \7135_b1 , \7122_b1 , \7134_b1 );
not ( \7134_b1 , w_22760 );
and ( \7135_b0 , \7122_b0 , w_22761 );
and ( w_22760 , w_22761 , \7134_b0 );
buf ( \7136_b1 , \7122_b1 );
not ( \7136_b1 , w_22762 );
not ( \7136_b0 , w_22763 );
and ( w_22762 , w_22763 , \7122_b0 );
or ( \7137_b1 , \7136_b1 , \7133_b1 );
not ( \7133_b1 , w_22764 );
and ( \7137_b0 , \7136_b0 , w_22765 );
and ( w_22764 , w_22765 , \7133_b0 );
or ( \7138_b1 , \7135_b1 , w_22767 );
not ( w_22767 , w_22768 );
and ( \7138_b0 , \7135_b0 , w_22769 );
and ( w_22768 ,  , w_22769 );
buf ( w_22767 , \7137_b1 );
not ( w_22767 , w_22770 );
not (  , w_22771 );
and ( w_22770 , w_22771 , \7137_b0 );
or ( \7139_b1 , \6769_b1 , \6811_b1 );
not ( \6811_b1 , w_22772 );
and ( \7139_b0 , \6769_b0 , w_22773 );
and ( w_22772 , w_22773 , \6811_b0 );
buf ( \7140_b1 , \6825_b1 );
not ( \7140_b1 , w_22774 );
not ( \7140_b0 , w_22775 );
and ( w_22774 , w_22775 , \6825_b0 );
or ( \7141_b1 , \7139_b1 , w_22777 );
not ( w_22777 , w_22778 );
and ( \7141_b0 , \7139_b0 , w_22779 );
and ( w_22778 ,  , w_22779 );
buf ( w_22777 , \7140_b1 );
not ( w_22777 , w_22780 );
not (  , w_22781 );
and ( w_22780 , w_22781 , \7140_b0 );
or ( \7142_b1 , \6823_b1 , w_22783 );
not ( w_22783 , w_22784 );
and ( \7142_b0 , \6823_b0 , w_22785 );
and ( w_22784 ,  , w_22785 );
buf ( w_22783 , \6801_b1 );
not ( w_22783 , w_22786 );
not (  , w_22787 );
and ( w_22786 , w_22787 , \6801_b0 );
or ( \7143_b1 , \7141_b1 , \7142_b1 );
not ( \7142_b1 , w_22788 );
and ( \7143_b0 , \7141_b0 , w_22789 );
and ( w_22788 , w_22789 , \7142_b0 );
buf ( \7144_b1 , \7141_b1 );
not ( \7144_b1 , w_22790 );
not ( \7144_b0 , w_22791 );
and ( w_22790 , w_22791 , \7141_b0 );
buf ( \7145_b1 , \7142_b1 );
not ( \7145_b1 , w_22792 );
not ( \7145_b0 , w_22793 );
and ( w_22792 , w_22793 , \7142_b0 );
or ( \7146_b1 , \7144_b1 , \7145_b1 );
not ( \7145_b1 , w_22794 );
and ( \7146_b0 , \7144_b0 , w_22795 );
and ( w_22794 , w_22795 , \7145_b0 );
or ( \7147_b1 , \7143_b1 , w_22797 );
not ( w_22797 , w_22798 );
and ( \7147_b0 , \7143_b0 , w_22799 );
and ( w_22798 ,  , w_22799 );
buf ( w_22797 , \7146_b1 );
not ( w_22797 , w_22800 );
not (  , w_22801 );
and ( w_22800 , w_22801 , \7146_b0 );
or ( \7148_b1 , \6910_b1 , \4694_b1 );
not ( \4694_b1 , w_22802 );
and ( \7148_b0 , \6910_b0 , w_22803 );
and ( w_22802 , w_22803 , \4694_b0 );
or ( \7149_b1 , \6811_b1 , w_22805 );
not ( w_22805 , w_22806 );
and ( \7149_b0 , \6811_b0 , w_22807 );
and ( w_22806 ,  , w_22807 );
buf ( w_22805 , \6825_b1 );
not ( w_22805 , w_22808 );
not (  , w_22809 );
and ( w_22808 , w_22809 , \6825_b0 );
buf ( \7150_b1 , \7149_b1 );
not ( \7150_b1 , w_22810 );
not ( \7150_b0 , w_22811 );
and ( w_22810 , w_22811 , \7149_b0 );
or ( \7151_b1 , \6769_b1 , \7150_b1 );
not ( \7150_b1 , w_22812 );
and ( \7151_b0 , \6769_b0 , w_22813 );
and ( w_22812 , w_22813 , \7150_b0 );
buf ( \7152_b1 , \6769_b1 );
not ( \7152_b1 , w_22814 );
not ( \7152_b0 , w_22815 );
and ( w_22814 , w_22815 , \6769_b0 );
or ( \7153_b1 , \7152_b1 , \7149_b1 );
not ( \7149_b1 , w_22816 );
and ( \7153_b0 , \7152_b0 , w_22817 );
and ( w_22816 , w_22817 , \7149_b0 );
or ( \7154_b1 , \7151_b1 , w_22819 );
not ( w_22819 , w_22820 );
and ( \7154_b0 , \7151_b0 , w_22821 );
and ( w_22820 ,  , w_22821 );
buf ( w_22819 , \7153_b1 );
not ( w_22819 , w_22822 );
not (  , w_22823 );
and ( w_22822 , w_22823 , \7153_b0 );
buf ( \7155_b1 , \6571_b1 );
not ( \7155_b1 , w_22824 );
not ( \7155_b0 , w_22825 );
and ( w_22824 , w_22825 , \6571_b0 );
buf ( \7156_b1 , \7155_b1 );
not ( \7156_b1 , w_22826 );
not ( \7156_b0 , w_22827 );
and ( w_22826 , w_22827 , \7155_b0 );
buf ( \7157_b1 , \6767_b1 );
not ( \7157_b1 , w_22828 );
not ( \7157_b0 , w_22829 );
and ( w_22828 , w_22829 , \6767_b0 );
buf ( \7158_b1 , \6573_b1 );
not ( \7158_b1 , w_22830 );
not ( \7158_b0 , w_22831 );
and ( w_22830 , w_22831 , \6573_b0 );
buf ( \7159_b1 , \7158_b1 );
not ( \7159_b1 , w_22832 );
not ( \7159_b0 , w_22833 );
and ( w_22832 , w_22833 , \7158_b0 );
or ( \7160_b1 , \7157_b1 , w_22834 );
or ( \7160_b0 , \7157_b0 , \7159_b0 );
not ( \7159_b0 , w_22835 );
and ( w_22835 , w_22834 , \7159_b1 );
or ( \7161_b1 , \7160_b1 , w_22837 );
not ( w_22837 , w_22838 );
and ( \7161_b0 , \7160_b0 , w_22839 );
and ( w_22838 ,  , w_22839 );
buf ( w_22837 , \6546_b1 );
not ( w_22837 , w_22840 );
not (  , w_22841 );
and ( w_22840 , w_22841 , \6546_b0 );
buf ( \7162_b1 , \7161_b1 );
not ( \7162_b1 , w_22842 );
not ( \7162_b0 , w_22843 );
and ( w_22842 , w_22843 , \7161_b0 );
or ( \7163_b1 , \7156_b1 , w_22844 );
or ( \7163_b0 , \7156_b0 , \7162_b0 );
not ( \7162_b0 , w_22845 );
and ( w_22845 , w_22844 , \7162_b1 );
or ( \7164_b1 , \7163_b1 , w_22847 );
not ( w_22847 , w_22848 );
and ( \7164_b0 , \7163_b0 , w_22849 );
and ( w_22848 ,  , w_22849 );
buf ( w_22847 , \6566_b1 );
not ( w_22847 , w_22850 );
not (  , w_22851 );
and ( w_22850 , w_22851 , \6566_b0 );
buf ( \7165_b1 , \6569_b1 );
not ( \7165_b1 , w_22852 );
not ( \7165_b0 , w_22853 );
and ( w_22852 , w_22853 , \6569_b0 );
or ( \7166_b1 , \7165_b1 , w_22855 );
not ( w_22855 , w_22856 );
and ( \7166_b0 , \7165_b0 , w_22857 );
and ( w_22856 ,  , w_22857 );
buf ( w_22855 , \6387_b1 );
not ( w_22855 , w_22858 );
not (  , w_22859 );
and ( w_22858 , w_22859 , \6387_b0 );
buf ( \7167_b1 , \7166_b1 );
not ( \7167_b1 , w_22860 );
not ( \7167_b0 , w_22861 );
and ( w_22860 , w_22861 , \7166_b0 );
or ( \7168_b1 , \7164_b1 , \7167_b1 );
not ( \7167_b1 , w_22862 );
and ( \7168_b0 , \7164_b0 , w_22863 );
and ( w_22862 , w_22863 , \7167_b0 );
buf ( \7169_b1 , \7164_b1 );
not ( \7169_b1 , w_22864 );
not ( \7169_b0 , w_22865 );
and ( w_22864 , w_22865 , \7164_b0 );
or ( \7170_b1 , \7169_b1 , \7166_b1 );
not ( \7166_b1 , w_22866 );
and ( \7170_b0 , \7169_b0 , w_22867 );
and ( w_22866 , w_22867 , \7166_b0 );
or ( \7171_b1 , \7168_b1 , w_22869 );
not ( w_22869 , w_22870 );
and ( \7171_b0 , \7168_b0 , w_22871 );
and ( w_22870 ,  , w_22871 );
buf ( w_22869 , \7170_b1 );
not ( w_22869 , w_22872 );
not (  , w_22873 );
and ( w_22872 , w_22873 , \7170_b0 );
buf ( \7172_b1 , \6571_b1 );
not ( \7172_b1 , w_22874 );
not ( \7172_b0 , w_22875 );
and ( w_22874 , w_22875 , \6571_b0 );
or ( \7173_b1 , \7172_b1 , w_22877 );
not ( w_22877 , w_22878 );
and ( \7173_b0 , \7172_b0 , w_22879 );
and ( w_22878 ,  , w_22879 );
buf ( w_22877 , \6566_b1 );
not ( w_22877 , w_22880 );
not (  , w_22881 );
and ( w_22880 , w_22881 , \6566_b0 );
buf ( \7174_b1 , \7173_b1 );
not ( \7174_b1 , w_22882 );
not ( \7174_b0 , w_22883 );
and ( w_22882 , w_22883 , \7173_b0 );
buf ( \7175_b1 , \7161_b1 );
not ( \7175_b1 , w_22884 );
not ( \7175_b0 , w_22885 );
and ( w_22884 , w_22885 , \7161_b0 );
or ( \7176_b1 , \7174_b1 , w_22886 );
or ( \7176_b0 , \7174_b0 , \7175_b0 );
not ( \7175_b0 , w_22887 );
and ( w_22887 , w_22886 , \7175_b1 );
or ( \7177_b1 , \7173_b1 , w_22888 );
or ( \7177_b0 , \7173_b0 , \7161_b0 );
not ( \7161_b0 , w_22889 );
and ( w_22889 , w_22888 , \7161_b1 );
or ( \7178_b1 , \7176_b1 , w_22891 );
not ( w_22891 , w_22892 );
and ( \7178_b0 , \7176_b0 , w_22893 );
and ( w_22892 ,  , w_22893 );
buf ( w_22891 , \7177_b1 );
not ( w_22891 , w_22894 );
not (  , w_22895 );
and ( w_22894 , w_22895 , \7177_b0 );
buf ( \7179_b1 , \6572_b1 );
not ( \7179_b1 , w_22896 );
not ( \7179_b0 , w_22897 );
and ( w_22896 , w_22897 , \6572_b0 );
buf ( \7180_b1 , \6767_b1 );
not ( \7180_b1 , w_22898 );
not ( \7180_b0 , w_22899 );
and ( w_22898 , w_22899 , \6767_b0 );
or ( \7181_b1 , \7179_b1 , w_22900 );
or ( \7181_b0 , \7179_b0 , \7180_b0 );
not ( \7180_b0 , w_22901 );
and ( w_22901 , w_22900 , \7180_b1 );
or ( \7182_b1 , \7181_b1 , w_22903 );
not ( w_22903 , w_22904 );
and ( \7182_b0 , \7181_b0 , w_22905 );
and ( w_22904 ,  , w_22905 );
buf ( w_22903 , \6542_b1 );
not ( w_22903 , w_22906 );
not (  , w_22907 );
and ( w_22906 , w_22907 , \6542_b0 );
or ( \7183_b1 , \6545_b1 , w_22909 );
not ( w_22909 , w_22910 );
and ( \7183_b0 , \6545_b0 , w_22911 );
and ( w_22910 ,  , w_22911 );
buf ( w_22909 , \6494_b1 );
not ( w_22909 , w_22912 );
not (  , w_22913 );
and ( w_22912 , w_22913 , \6494_b0 );
buf ( \7184_b1 , \7183_b1 );
not ( \7184_b1 , w_22914 );
not ( \7184_b0 , w_22915 );
and ( w_22914 , w_22915 , \7183_b0 );
or ( \7185_b1 , \7182_b1 , \7184_b1 );
not ( \7184_b1 , w_22916 );
and ( \7185_b0 , \7182_b0 , w_22917 );
and ( w_22916 , w_22917 , \7184_b0 );
buf ( \7186_b1 , \7182_b1 );
not ( \7186_b1 , w_22918 );
not ( \7186_b0 , w_22919 );
and ( w_22918 , w_22919 , \7182_b0 );
or ( \7187_b1 , \7186_b1 , \7183_b1 );
not ( \7183_b1 , w_22920 );
and ( \7187_b0 , \7186_b0 , w_22921 );
and ( w_22920 , w_22921 , \7183_b0 );
or ( \7188_b1 , \7185_b1 , w_22923 );
not ( w_22923 , w_22924 );
and ( \7188_b0 , \7185_b0 , w_22925 );
and ( w_22924 ,  , w_22925 );
buf ( w_22923 , \7187_b1 );
not ( w_22923 , w_22926 );
not (  , w_22927 );
and ( w_22926 , w_22927 , \7187_b0 );
or ( \7189_b1 , \6542_b1 , w_22929 );
not ( w_22929 , w_22930 );
and ( \7189_b0 , \6542_b0 , w_22931 );
and ( w_22930 ,  , w_22931 );
buf ( w_22929 , \6572_b1 );
not ( w_22929 , w_22932 );
not (  , w_22933 );
and ( w_22932 , w_22933 , \6572_b0 );
buf ( \7190_b1 , \7189_b1 );
not ( \7190_b1 , w_22934 );
not ( \7190_b0 , w_22935 );
and ( w_22934 , w_22935 , \7189_b0 );
buf ( \7191_b1 , \6767_b1 );
not ( \7191_b1 , w_22936 );
not ( \7191_b0 , w_22937 );
and ( w_22936 , w_22937 , \6767_b0 );
or ( \7192_b1 , \7190_b1 , w_22938 );
or ( \7192_b0 , \7190_b0 , \7191_b0 );
not ( \7191_b0 , w_22939 );
and ( w_22939 , w_22938 , \7191_b1 );
or ( \7193_b1 , \7189_b1 , w_22940 );
or ( \7193_b0 , \7189_b0 , \6767_b0 );
not ( \6767_b0 , w_22941 );
and ( w_22941 , w_22940 , \6767_b1 );
or ( \7194_b1 , \7192_b1 , w_22943 );
not ( w_22943 , w_22944 );
and ( \7194_b0 , \7192_b0 , w_22945 );
and ( w_22944 ,  , w_22945 );
buf ( w_22943 , \7193_b1 );
not ( w_22943 , w_22946 );
not (  , w_22947 );
and ( w_22946 , w_22947 , \7193_b0 );
or ( \7195_b1 , \6766_b1 , w_22949 );
not ( w_22949 , w_22950 );
and ( \7195_b0 , \6766_b0 , w_22951 );
and ( w_22950 ,  , w_22951 );
buf ( w_22949 , \6613_b1 );
not ( w_22949 , w_22952 );
not (  , w_22953 );
and ( w_22952 , w_22953 , \6613_b0 );
or ( \7196_b1 , \6749_b1 , \6758_b1 );
not ( \6758_b1 , w_22954 );
and ( \7196_b0 , \6749_b0 , w_22955 );
and ( w_22954 , w_22955 , \6758_b0 );
or ( \7197_b1 , \7196_b1 , w_22957 );
not ( w_22957 , w_22958 );
and ( \7197_b0 , \7196_b0 , w_22959 );
and ( w_22958 ,  , w_22959 );
buf ( w_22957 , \6760_b1 );
not ( w_22957 , w_22960 );
not (  , w_22961 );
and ( w_22960 , w_22961 , \6760_b0 );
or ( \7198_b1 , \6762_b1 , w_22963 );
not ( w_22963 , w_22964 );
and ( \7198_b0 , \6762_b0 , w_22965 );
and ( w_22964 ,  , w_22965 );
buf ( w_22963 , \6650_b1 );
not ( w_22963 , w_22966 );
not (  , w_22967 );
and ( w_22966 , w_22967 , \6650_b0 );
or ( \7199_b1 , \6748_b1 , w_22969 );
not ( w_22969 , w_22970 );
and ( \7199_b0 , \6748_b0 , w_22971 );
and ( w_22970 ,  , w_22971 );
buf ( w_22969 , \6745_b1 );
not ( w_22969 , w_22972 );
not (  , w_22973 );
and ( w_22972 , w_22973 , \6745_b0 );
or ( \7200_b1 , \6694_b1 , w_22975 );
not ( w_22975 , w_22976 );
and ( \7200_b0 , \6694_b0 , w_22977 );
and ( w_22976 ,  , w_22977 );
buf ( w_22975 , \6725_b1 );
not ( w_22975 , w_22978 );
not (  , w_22979 );
and ( w_22978 , w_22979 , \6725_b0 );
or ( \7201_b1 , \6723_b1 , w_22981 );
not ( w_22981 , w_22982 );
and ( \7201_b0 , \6723_b0 , w_22983 );
and ( w_22982 ,  , w_22983 );
buf ( w_22981 , \6719_b1 );
not ( w_22981 , w_22984 );
not (  , w_22985 );
and ( w_22984 , w_22985 , \6719_b0 );
or ( \7202_b1 , \6707_b1 , \6709_b1 );
not ( \6709_b1 , w_22986 );
and ( \7202_b0 , \6707_b0 , w_22987 );
and ( w_22986 , w_22987 , \6709_b0 );
or ( \7203_b1 , \7202_b1 , w_22989 );
not ( w_22989 , w_22990 );
and ( \7203_b0 , \7202_b0 , w_22991 );
and ( w_22990 ,  , w_22991 );
buf ( w_22989 , \6710_b1 );
not ( w_22989 , w_22992 );
not (  , w_22993 );
and ( w_22992 , w_22993 , \6710_b0 );
buf ( \7204_b1 , \6708_b1 );
not ( \7204_b1 , w_22994 );
not ( \7204_b0 , w_22995 );
and ( w_22994 , w_22995 , \6708_b0 );
or ( \7205_b1 , \6897_b1 , \5543_b1 );
not ( \5543_b1 , w_22996 );
and ( \7205_b0 , \6897_b0 , w_22997 );
and ( w_22996 , w_22997 , \5543_b0 );
or ( \7206_b1 , \7037_b1 , \7205_b1 );
xor ( \7206_b0 , \7037_b0 , w_22998 );
not ( w_22998 , w_22999 );
and ( w_22999 , \7205_b1 , \7205_b0 );
or ( \7207_b1 , \7198_b1 , \7197_b1 );
xor ( \7207_b0 , \7198_b0 , w_23000 );
not ( w_23000 , w_23001 );
and ( w_23001 , \7197_b1 , \7197_b0 );
buf ( \7208_b1 , \6760_b1 );
not ( \7208_b1 , w_23002 );
not ( \7208_b0 , w_23003 );
and ( w_23002 , w_23003 , \6760_b0 );
or ( \7209_b1 , \7208_b1 , w_23005 );
not ( w_23005 , w_23006 );
and ( \7209_b0 , \7208_b0 , w_23007 );
and ( w_23006 ,  , w_23007 );
buf ( w_23005 , \6758_b1 );
not ( w_23005 , w_23008 );
not (  , w_23009 );
and ( w_23008 , w_23009 , \6758_b0 );
or ( \7210_b1 , \6749_b1 , w_23010 );
xor ( \7210_b0 , \6749_b0 , w_23012 );
not ( w_23012 , w_23013 );
and ( w_23013 , w_23010 , w_23011 );
buf ( w_23010 , \7209_b1 );
not ( w_23010 , w_23014 );
not ( w_23011 , w_23015 );
and ( w_23014 , w_23015 , \7209_b0 );
or ( \7211_b1 , \6727_b1 , w_23016 );
xor ( \7211_b0 , \6727_b0 , w_23018 );
not ( w_23018 , w_23019 );
and ( w_23019 , w_23016 , w_23017 );
buf ( w_23016 , \7199_b1 );
not ( w_23016 , w_23020 );
not ( w_23017 , w_23021 );
and ( w_23020 , w_23021 , \7199_b0 );
or ( \7212_b1 , \7200_b1 , w_23022 );
xor ( \7212_b0 , \7200_b0 , w_23024 );
not ( w_23024 , w_23025 );
and ( w_23025 , w_23022 , w_23023 );
buf ( w_23022 , \6724_b1 );
not ( w_23022 , w_23026 );
not ( w_23023 , w_23027 );
and ( w_23026 , w_23027 , \6724_b0 );
or ( \7213_b1 , \6710_b1 , w_23028 );
xor ( \7213_b0 , \6710_b0 , w_23030 );
not ( w_23030 , w_23031 );
and ( w_23031 , w_23028 , w_23029 );
buf ( w_23028 , \7201_b1 );
not ( w_23028 , w_23032 );
not ( w_23029 , w_23033 );
and ( w_23032 , w_23033 , \7201_b0 );
buf ( \7214_b1 , \7195_b1 );
not ( \7214_b1 , w_23034 );
not ( \7214_b0 , w_23035 );
and ( w_23034 , w_23035 , \7195_b0 );
or ( \7215_b1 , \6763_b1 , \7214_b1 );
xor ( \7215_b0 , \6763_b0 , w_23036 );
not ( w_23036 , w_23037 );
and ( w_23037 , \7214_b1 , \7214_b0 );
or ( \7216_b1 , \7148_b1 , \6904_b1 );
xor ( \7216_b0 , \7148_b0 , w_23038 );
not ( w_23038 , w_23039 );
and ( w_23039 , \6904_b1 , \6904_b0 );
or ( \115_b1 , \113_b1 , w_23040 );
not ( w_23040 , w_23042 );
and ( \115_b0 , \113_b0 , w_23043 );
and ( w_23042 , w_23043 , w_23041 );
or ( w_23040 , \114_b1 , \b[9]_b1 );
not ( \b[9]_b1 , w_23044 );
and ( w_23041 , \114_b0 , w_23045 );
and ( w_23044 , w_23045 , \b[9]_b0 );
or ( \207_b1 , \205_b1 , w_23046 );
not ( w_23046 , w_23048 );
and ( \207_b0 , \205_b0 , w_23049 );
and ( w_23048 , w_23049 , w_23047 );
or ( w_23046 , \206_b1 , \b[7]_b1 );
not ( \b[7]_b1 , w_23050 );
and ( w_23047 , \206_b0 , w_23051 );
and ( w_23050 , w_23051 , \b[7]_b0 );
or ( \340_b1 , \338_b1 , w_23052 );
not ( w_23052 , w_23056 );
and ( \340_b0 , \338_b0 , w_23057 );
and ( w_23056 , w_23057 , w_23053 );
or ( w_23052 , \339_b1 , w_23054 );
not ( w_23054 , w_23058 );
and ( w_23053 , \339_b0 , w_23059 );
and ( w_23058 , w_23059 , w_23055 );
buf ( w_23054 , \b[5]_b1 );
not ( w_23054 , w_23060 );
not ( w_23055 , w_23061 );
and ( w_23060 , w_23061 , \b[5]_b0 );
or ( \532_b1 , \530_b1 , w_23062 );
not ( w_23062 , w_23066 );
and ( \532_b0 , \530_b0 , w_23067 );
and ( w_23066 , w_23067 , w_23063 );
or ( w_23062 , \423_b1 , w_23064 );
not ( w_23064 , w_23068 );
and ( w_23063 , \423_b0 , w_23069 );
and ( w_23068 , w_23069 , w_23065 );
buf ( w_23064 , \531_b1 );
not ( w_23064 , w_23070 );
not ( w_23065 , w_23071 );
and ( w_23070 , w_23071 , \531_b0 );
or ( \541_b1 , \328_b1 , w_23072 );
not ( w_23072 , w_23076 );
and ( \541_b0 , \328_b0 , w_23077 );
and ( w_23076 , w_23077 , w_23073 );
or ( w_23072 , \426_b1 , w_23074 );
not ( w_23074 , w_23078 );
and ( w_23073 , \426_b0 , w_23079 );
and ( w_23078 , w_23079 , w_23075 );
or ( w_23074 , \532_b1 , \540_b1 );
not ( \540_b1 , w_23080 );
and ( w_23075 , \532_b0 , w_23081 );
and ( w_23080 , w_23081 , \540_b0 );
or ( \553_b1 , \545_b1 , w_23082 );
not ( w_23082 , w_23084 );
and ( \553_b0 , \545_b0 , w_23085 );
and ( w_23084 , w_23085 , w_23083 );
or ( w_23082 , \551_b1 , \552_b1 );
not ( \552_b1 , w_23086 );
and ( w_23083 , \551_b0 , w_23087 );
and ( w_23086 , w_23087 , \552_b0 );
or ( \587_b1 , \585_b1 , w_23088 );
not ( w_23088 , w_23092 );
and ( \587_b0 , \585_b0 , w_23093 );
and ( w_23092 , w_23093 , w_23089 );
or ( w_23088 , \586_b1 , w_23090 );
not ( w_23090 , w_23094 );
and ( w_23089 , \586_b0 , w_23095 );
and ( w_23094 , w_23095 , w_23091 );
buf ( w_23090 , \b[11]_b1 );
not ( w_23090 , w_23096 );
not ( w_23091 , w_23097 );
and ( w_23096 , w_23097 , \b[11]_b0 );
or ( \657_b1 , \652_b1 , w_23098 );
not ( w_23098 , w_23102 );
and ( \657_b0 , \652_b0 , w_23103 );
and ( w_23102 , w_23103 , w_23099 );
or ( w_23098 , \529_b1 , w_23100 );
not ( w_23100 , w_23104 );
and ( w_23099 , \529_b0 , w_23105 );
and ( w_23104 , w_23105 , w_23101 );
buf ( w_23100 , \403_b1 );
not ( w_23100 , w_23106 );
not ( w_23101 , w_23107 );
and ( w_23106 , w_23107 , \403_b0 );
or ( \689_b1 , \687_b1 , w_23108 );
not ( w_23108 , w_23112 );
and ( \689_b0 , \687_b0 , w_23113 );
and ( w_23112 , w_23113 , w_23109 );
or ( w_23108 , \688_b1 , w_23110 );
not ( w_23110 , w_23114 );
and ( w_23109 , \688_b0 , w_23115 );
and ( w_23114 , w_23115 , w_23111 );
buf ( w_23110 , \c[7]_b1 );
not ( w_23110 , w_23116 );
not ( w_23111 , w_23117 );
and ( w_23116 , w_23117 , \c[7]_b0 );
or ( \764_b1 , \762_b1 , w_23118 );
not ( w_23118 , w_23122 );
and ( \764_b0 , \762_b0 , w_23123 );
and ( w_23122 , w_23123 , w_23119 );
or ( w_23118 , \763_b1 , w_23120 );
not ( w_23120 , w_23124 );
and ( w_23119 , \763_b0 , w_23125 );
and ( w_23124 , w_23125 , w_23121 );
buf ( w_23120 , \c[5]_b1 );
not ( w_23120 , w_23126 );
not ( w_23121 , w_23127 );
and ( w_23126 , w_23127 , \c[5]_b0 );
or ( \837_b1 , \834_b1 , w_23128 );
not ( w_23128 , w_23132 );
and ( \837_b0 , \834_b0 , w_23133 );
and ( w_23132 , w_23133 , w_23129 );
or ( w_23128 , \c[3]_b1 , w_23130 );
not ( w_23130 , w_23134 );
and ( w_23129 , \c[3]_b0 , w_23135 );
and ( w_23134 , w_23135 , w_23131 );
buf ( w_23130 , \836_b1 );
not ( w_23130 , w_23136 );
not ( w_23131 , w_23137 );
and ( w_23136 , w_23137 , \836_b0 );
or ( \942_b1 , \940_b1 , w_23138 );
not ( w_23138 , w_23142 );
and ( \942_b0 , \940_b0 , w_23143 );
and ( w_23142 , w_23143 , w_23139 );
or ( w_23138 , \941_b1 , w_23140 );
not ( w_23140 , w_23144 );
and ( w_23139 , \941_b0 , w_23145 );
and ( w_23144 , w_23145 , w_23141 );
buf ( w_23140 , \d[5]_b1 );
not ( w_23140 , w_23146 );
not ( w_23141 , w_23147 );
and ( w_23146 , w_23147 , \d[5]_b0 );
or ( \1071_b1 , \1066_b1 , w_23148 );
not ( w_23148 , w_23152 );
and ( \1071_b0 , \1066_b0 , w_23153 );
and ( w_23152 , w_23153 , w_23149 );
or ( w_23148 , \1069_b1 , w_23150 );
not ( w_23150 , w_23154 );
and ( w_23149 , \1069_b0 , w_23155 );
and ( w_23154 , w_23155 , w_23151 );
buf ( w_23150 , \1070_b1 );
not ( w_23150 , w_23156 );
not ( w_23151 , w_23157 );
and ( w_23156 , w_23157 , \1070_b0 );
or ( \1112_b1 , \1110_b1 , w_23158 );
not ( w_23158 , w_23162 );
and ( \1112_b0 , \1110_b0 , w_23163 );
and ( w_23162 , w_23163 , w_23159 );
or ( w_23158 , \1111_b1 , w_23160 );
not ( w_23160 , w_23164 );
and ( w_23159 , \1111_b0 , w_23165 );
and ( w_23164 , w_23165 , w_23161 );
buf ( w_23160 , \d[7]_b1 );
not ( w_23160 , w_23166 );
not ( w_23161 , w_23167 );
and ( w_23166 , w_23167 , \d[7]_b0 );
or ( \1334_b1 , \1303_b1 , w_23168 );
not ( w_23168 , w_23172 );
and ( \1334_b0 , \1303_b0 , w_23173 );
and ( w_23172 , w_23173 , w_23169 );
or ( w_23168 , \1318_b1 , w_23170 );
not ( w_23170 , w_23174 );
and ( w_23169 , \1318_b0 , w_23175 );
and ( w_23174 , w_23175 , w_23171 );
buf ( w_23170 , \1333_b1 );
not ( w_23170 , w_23176 );
not ( w_23171 , w_23177 );
and ( w_23176 , w_23177 , \1333_b0 );
or ( \1391_b1 , \1382_b1 , w_23178 );
not ( w_23178 , w_23182 );
and ( \1391_b0 , \1382_b0 , w_23183 );
and ( w_23182 , w_23183 , w_23179 );
or ( w_23178 , \1385_b1 , w_23180 );
not ( w_23180 , w_23184 );
and ( w_23179 , \1385_b0 , w_23185 );
and ( w_23184 , w_23185 , w_23181 );
buf ( w_23180 , \1390_b1 );
not ( w_23180 , w_23186 );
not ( w_23181 , w_23187 );
and ( w_23186 , w_23187 , \1390_b0 );
or ( \1443_b1 , \1407_b1 , w_23188 );
not ( w_23188 , w_23190 );
and ( \1443_b0 , \1407_b0 , w_23191 );
and ( w_23190 , w_23191 , w_23189 );
or ( w_23188 , \1410_b1 , \1442_b1 );
not ( \1442_b1 , w_23192 );
and ( w_23189 , \1410_b0 , w_23193 );
and ( w_23192 , w_23193 , \1442_b0 );
or ( \1487_b1 , \1485_b1 , w_23194 );
not ( w_23194 , w_23198 );
and ( \1487_b0 , \1485_b0 , w_23199 );
and ( w_23198 , w_23199 , w_23195 );
or ( w_23194 , \1177_b1 , w_23196 );
not ( w_23196 , w_23200 );
and ( w_23195 , \1177_b0 , w_23201 );
and ( w_23200 , w_23201 , w_23197 );
buf ( w_23196 , \1486_b1 );
not ( w_23196 , w_23202 );
not ( w_23197 , w_23203 );
and ( w_23202 , w_23203 , \1486_b0 );
or ( \1501_b1 , \1499_b1 , w_23204 );
not ( w_23204 , w_23208 );
and ( \1501_b0 , \1499_b0 , w_23209 );
and ( w_23208 , w_23209 , w_23205 );
or ( w_23204 , \1240_b1 , w_23206 );
not ( w_23206 , w_23210 );
and ( w_23205 , \1240_b0 , w_23211 );
and ( w_23210 , w_23211 , w_23207 );
buf ( w_23206 , \1500_b1 );
not ( w_23206 , w_23212 );
not ( w_23207 , w_23213 );
and ( w_23212 , w_23213 , \1500_b0 );
or ( \1649_b1 , \1647_b1 , w_23214 );
not ( w_23214 , w_23216 );
and ( \1649_b0 , \1647_b0 , w_23217 );
and ( w_23216 , w_23217 , w_23215 );
or ( w_23214 , \1648_b1 , \d[13]_b1 );
not ( \d[13]_b1 , w_23218 );
and ( w_23215 , \1648_b0 , w_23219 );
and ( w_23218 , w_23219 , \d[13]_b0 );
or ( \1669_b1 , \1667_b1 , w_23220 );
not ( w_23220 , w_23224 );
and ( \1669_b0 , \1667_b0 , w_23225 );
and ( w_23224 , w_23225 , w_23221 );
or ( w_23220 , \1668_b1 , w_23222 );
not ( w_23222 , w_23226 );
and ( w_23221 , \1668_b0 , w_23227 );
and ( w_23226 , w_23227 , w_23223 );
buf ( w_23222 , \d[15]_b1 );
not ( w_23222 , w_23228 );
not ( w_23223 , w_23229 );
and ( w_23228 , w_23229 , \d[15]_b0 );
or ( \1859_b1 , \1857_b1 , w_23230 );
not ( w_23230 , w_23234 );
and ( \1859_b0 , \1857_b0 , w_23235 );
and ( w_23234 , w_23235 , w_23231 );
or ( w_23230 , \1858_b1 , w_23232 );
not ( w_23232 , w_23236 );
and ( w_23231 , \1858_b0 , w_23237 );
and ( w_23236 , w_23237 , w_23233 );
buf ( w_23232 , \d[11]_b1 );
not ( w_23232 , w_23238 );
not ( w_23233 , w_23239 );
and ( w_23238 , w_23239 , \d[11]_b0 );
or ( \2035_b1 , \2033_b1 , w_23240 );
not ( w_23240 , w_23242 );
and ( \2035_b0 , \2033_b0 , w_23243 );
and ( w_23242 , w_23243 , w_23241 );
or ( w_23240 , \2034_b1 , \d[9]_b1 );
not ( \d[9]_b1 , w_23244 );
and ( w_23241 , \2034_b0 , w_23245 );
and ( w_23244 , w_23245 , \d[9]_b0 );
or ( \2224_b1 , \1954_b1 , w_23246 );
not ( w_23246 , w_23248 );
and ( \2224_b0 , \1954_b0 , w_23249 );
and ( w_23248 , w_23249 , w_23247 );
or ( w_23246 , \2223_b1 , \2031_b1 );
not ( \2031_b1 , w_23250 );
and ( w_23247 , \2223_b0 , w_23251 );
and ( w_23250 , w_23251 , \2031_b0 );
or ( \2324_b1 , \2322_b1 , w_23252 );
not ( w_23252 , w_23256 );
and ( \2324_b0 , \2322_b0 , w_23257 );
and ( w_23256 , w_23257 , w_23253 );
or ( w_23252 , \2323_b1 , w_23254 );
not ( w_23254 , w_23258 );
and ( w_23253 , \2323_b0 , w_23259 );
and ( w_23258 , w_23259 , w_23255 );
buf ( w_23254 , \c[11]_b1 );
not ( w_23254 , w_23260 );
not ( w_23255 , w_23261 );
and ( w_23260 , w_23261 , \c[11]_b0 );
or ( \2432_b1 , \2430_b1 , w_23262 );
not ( w_23262 , w_23264 );
and ( \2432_b0 , \2430_b0 , w_23265 );
and ( w_23264 , w_23265 , w_23263 );
or ( w_23262 , \2431_b1 , \c[13]_b1 );
not ( \c[13]_b1 , w_23266 );
and ( w_23263 , \2431_b0 , w_23267 );
and ( w_23266 , w_23267 , \c[13]_b0 );
or ( \2574_b1 , \2572_b1 , w_23268 );
not ( w_23268 , w_23272 );
and ( \2574_b0 , \2572_b0 , w_23273 );
and ( w_23272 , w_23273 , w_23269 );
or ( w_23268 , \2573_b1 , w_23270 );
not ( w_23270 , w_23274 );
and ( w_23269 , \2573_b0 , w_23275 );
and ( w_23274 , w_23275 , w_23271 );
buf ( w_23270 , \c[15]_b1 );
not ( w_23270 , w_23276 );
not ( w_23271 , w_23277 );
and ( w_23276 , w_23277 , \c[15]_b0 );
or ( \2739_b1 , \2737_b1 , w_23278 );
not ( w_23278 , w_23280 );
and ( \2739_b0 , \2737_b0 , w_23281 );
and ( w_23280 , w_23281 , w_23279 );
or ( w_23278 , \2738_b1 , \c[9]_b1 );
not ( \c[9]_b1 , w_23282 );
and ( w_23279 , \2738_b0 , w_23283 );
and ( w_23282 , w_23283 , \c[9]_b0 );
or ( \2901_b1 , \2869_b1 , w_23284 );
not ( w_23284 , w_23290 );
and ( \2901_b0 , \2869_b0 , w_23291 );
and ( w_23290 , w_23291 , w_23285 );
or ( w_23284 , \2892_b1 , w_23286 );
not ( w_23286 , w_23292 );
and ( w_23285 , \2892_b0 , w_23293 );
and ( w_23292 , w_23293 , w_23287 );
or ( w_23286 , \2900_b1 , w_23288 );
not ( w_23288 , w_23294 );
and ( w_23287 , \2900_b0 , w_23295 );
and ( w_23294 , w_23295 , w_23289 );
buf ( w_23288 , \782_b1 );
not ( w_23288 , w_23296 );
not ( w_23289 , w_23297 );
and ( w_23296 , w_23297 , \782_b0 );
or ( \2928_b1 , \2921_b1 , w_23298 );
not ( w_23298 , w_23300 );
and ( \2928_b0 , \2921_b0 , w_23301 );
and ( w_23300 , w_23301 , w_23299 );
or ( w_23298 , \2927_b1 , \2728_b1 );
not ( \2728_b1 , w_23302 );
and ( w_23299 , \2927_b0 , w_23303 );
and ( w_23302 , w_23303 , \2728_b0 );
or ( \2966_b1 , \1487_b1 , w_23304 );
not ( w_23304 , w_23308 );
and ( \2966_b0 , \1487_b0 , w_23309 );
and ( w_23308 , w_23309 , w_23305 );
or ( w_23304 , \1186_b1 , w_23306 );
not ( w_23306 , w_23310 );
and ( w_23305 , \1186_b0 , w_23311 );
and ( w_23310 , w_23311 , w_23307 );
buf ( w_23306 , \1184_b1 );
not ( w_23306 , w_23312 );
not ( w_23307 , w_23313 );
and ( w_23312 , w_23313 , \1184_b0 );
or ( \2968_b1 , \1209_b1 , w_23314 );
not ( w_23314 , w_23318 );
and ( \2968_b0 , \1209_b0 , w_23319 );
and ( w_23318 , w_23319 , w_23315 );
or ( w_23314 , \1482_b1 , w_23316 );
not ( w_23316 , w_23320 );
and ( w_23315 , \1482_b0 , w_23321 );
and ( w_23320 , w_23321 , w_23317 );
buf ( w_23316 , \1202_b1 );
not ( w_23316 , w_23322 );
not ( w_23317 , w_23323 );
and ( w_23322 , w_23323 , \1202_b0 );
or ( \2972_b1 , \1204_b1 , w_23324 );
not ( w_23324 , w_23326 );
and ( \2972_b0 , \1204_b0 , w_23327 );
and ( w_23326 , w_23327 , w_23325 );
or ( w_23324 , \1210_b1 , \1200_b1 );
not ( \1200_b1 , w_23328 );
and ( w_23325 , \1210_b0 , w_23329 );
and ( w_23328 , w_23329 , \1200_b0 );
or ( \2993_b1 , \2979_b1 , w_23330 );
not ( w_23330 , w_23332 );
and ( \2993_b0 , \2979_b0 , w_23333 );
and ( w_23332 , w_23333 , w_23331 );
or ( w_23330 , \2985_b1 , \2992_b1 );
not ( \2992_b1 , w_23334 );
and ( w_23331 , \2985_b0 , w_23335 );
and ( w_23334 , w_23335 , \2992_b0 );
or ( \3028_b1 , \1501_b1 , w_23336 );
not ( w_23336 , w_23340 );
and ( \3028_b0 , \1501_b0 , w_23341 );
and ( w_23340 , w_23341 , w_23337 );
or ( w_23336 , \1249_b1 , w_23338 );
not ( w_23338 , w_23342 );
and ( w_23337 , \1249_b0 , w_23343 );
and ( w_23342 , w_23343 , w_23339 );
buf ( w_23338 , \1247_b1 );
not ( w_23338 , w_23344 );
not ( w_23339 , w_23345 );
and ( w_23344 , w_23345 , \1247_b0 );
or ( \3030_b1 , \1272_b1 , w_23346 );
not ( w_23346 , w_23350 );
and ( \3030_b0 , \1272_b0 , w_23351 );
and ( w_23350 , w_23351 , w_23347 );
or ( w_23346 , \1496_b1 , w_23348 );
not ( w_23348 , w_23352 );
and ( w_23347 , \1496_b0 , w_23353 );
and ( w_23352 , w_23353 , w_23349 );
buf ( w_23348 , \1265_b1 );
not ( w_23348 , w_23354 );
not ( w_23349 , w_23355 );
and ( w_23354 , w_23355 , \1265_b0 );
or ( \3034_b1 , \1267_b1 , w_23356 );
not ( w_23356 , w_23358 );
and ( \3034_b0 , \1267_b0 , w_23359 );
and ( w_23358 , w_23359 , w_23357 );
or ( w_23356 , \1273_b1 , \1263_b1 );
not ( \1263_b1 , w_23360 );
and ( w_23357 , \1273_b0 , w_23361 );
and ( w_23360 , w_23361 , \1263_b0 );
or ( \3055_b1 , \3041_b1 , w_23362 );
not ( w_23362 , w_23364 );
and ( \3055_b0 , \3041_b0 , w_23365 );
and ( w_23364 , w_23365 , w_23363 );
or ( w_23362 , \3047_b1 , \3054_b1 );
not ( \3054_b1 , w_23366 );
and ( w_23363 , \3047_b0 , w_23367 );
and ( w_23366 , w_23367 , \3054_b0 );
or ( \3103_b1 , \3102_b1 , w_23368 );
not ( w_23368 , w_23372 );
and ( \3103_b0 , \3102_b0 , w_23373 );
and ( w_23372 , w_23373 , w_23369 );
or ( w_23368 , \b[15]_b1 , w_23370 );
not ( w_23370 , w_23374 );
and ( w_23369 , \b[15]_b0 , w_23375 );
and ( w_23374 , w_23375 , w_23371 );
buf ( w_23370 , \c[15]_b1 );
not ( w_23370 , w_23376 );
not ( w_23371 , w_23377 );
and ( w_23376 , w_23377 , \c[15]_b0 );
or ( \3120_b1 , \1316_b1 , w_23378 );
not ( w_23378 , w_23382 );
and ( \3120_b0 , \1316_b0 , w_23383 );
and ( w_23382 , w_23383 , w_23379 );
or ( w_23378 , \b[11]_b1 , w_23380 );
not ( w_23380 , w_23384 );
and ( w_23379 , \b[11]_b0 , w_23385 );
and ( w_23384 , w_23385 , w_23381 );
buf ( w_23380 , \c[11]_b1 );
not ( w_23380 , w_23386 );
not ( w_23381 , w_23387 );
and ( w_23386 , w_23387 , \c[11]_b0 );
or ( \3135_b1 , \2979_b1 , w_23388 );
not ( w_23388 , w_23390 );
and ( \3135_b0 , \2979_b0 , w_23391 );
and ( w_23390 , w_23391 , w_23389 );
or ( w_23388 , \2991_b1 , \3134_b1 );
not ( \3134_b1 , w_23392 );
and ( w_23389 , \2991_b0 , w_23393 );
and ( w_23392 , w_23393 , \3134_b0 );
or ( \3151_b1 , \3041_b1 , w_23394 );
not ( w_23394 , w_23396 );
and ( \3151_b0 , \3041_b0 , w_23397 );
and ( w_23396 , w_23397 , w_23395 );
or ( w_23394 , \3053_b1 , \3150_b1 );
not ( \3150_b1 , w_23398 );
and ( w_23395 , \3053_b0 , w_23399 );
and ( w_23398 , w_23399 , \3150_b0 );
or ( \3213_b1 , \1316_b1 , w_23400 );
not ( w_23400 , w_23404 );
and ( \3213_b0 , \1316_b0 , w_23405 );
and ( w_23404 , w_23405 , w_23401 );
or ( w_23400 , \b[6]_b1 , w_23402 );
not ( w_23402 , w_23406 );
and ( w_23401 , \b[6]_b0 , w_23407 );
and ( w_23406 , w_23407 , w_23403 );
buf ( w_23402 , \c[6]_b1 );
not ( w_23402 , w_23408 );
not ( w_23403 , w_23409 );
and ( w_23408 , w_23409 , \c[6]_b0 );
or ( \3270_b1 , \3213_b1 , w_23410 );
not ( w_23410 , w_23414 );
and ( \3270_b0 , \3213_b0 , w_23415 );
and ( w_23414 , w_23415 , w_23411 );
or ( w_23410 , \3215_b1 , w_23412 );
not ( w_23412 , w_23416 );
and ( w_23411 , \3215_b0 , w_23417 );
and ( w_23416 , w_23417 , w_23413 );
buf ( w_23412 , \3269_b1 );
not ( w_23412 , w_23418 );
not ( w_23413 , w_23419 );
and ( w_23418 , w_23419 , \3269_b0 );
or ( \3293_b1 , \3102_b1 , w_23420 );
not ( w_23420 , w_23424 );
and ( \3293_b0 , \3102_b0 , w_23425 );
and ( w_23424 , w_23425 , w_23421 );
or ( w_23420 , \b[14]_b1 , w_23422 );
not ( w_23422 , w_23426 );
and ( w_23421 , \b[14]_b0 , w_23427 );
and ( w_23426 , w_23427 , w_23423 );
buf ( w_23422 , \c[14]_b1 );
not ( w_23422 , w_23428 );
not ( w_23423 , w_23429 );
and ( w_23428 , w_23429 , \c[14]_b0 );
or ( \3311_b1 , \2979_b1 , w_23430 );
not ( w_23430 , w_23432 );
and ( \3311_b0 , \2979_b0 , w_23433 );
and ( w_23432 , w_23433 , w_23431 );
or ( w_23430 , \2992_b1 , \2982_b1 );
not ( \2982_b1 , w_23434 );
and ( w_23431 , \2992_b0 , w_23435 );
and ( w_23434 , w_23435 , \2982_b0 );
or ( \3324_b1 , \3041_b1 , w_23436 );
not ( w_23436 , w_23438 );
and ( \3324_b0 , \3041_b0 , w_23439 );
and ( w_23438 , w_23439 , w_23437 );
or ( w_23436 , \3054_b1 , \3044_b1 );
not ( \3044_b1 , w_23440 );
and ( w_23437 , \3054_b0 , w_23441 );
and ( w_23440 , w_23441 , \3044_b0 );
or ( \3366_b1 , \3287_b1 , w_23442 );
not ( w_23442 , w_23448 );
and ( \3366_b0 , \3287_b0 , w_23449 );
and ( w_23448 , w_23449 , w_23443 );
or ( w_23442 , \3288_b1 , w_23444 );
not ( w_23444 , w_23450 );
and ( w_23443 , \3288_b0 , w_23451 );
and ( w_23450 , w_23451 , w_23445 );
or ( w_23444 , \3346_b1 , w_23446 );
not ( w_23446 , w_23452 );
and ( w_23445 , \3346_b0 , w_23453 );
and ( w_23452 , w_23453 , w_23447 );
buf ( w_23446 , \3365_b1 );
not ( w_23446 , w_23454 );
not ( w_23447 , w_23455 );
and ( w_23454 , w_23455 , \3365_b0 );
or ( \3479_b1 , \3102_b1 , w_23456 );
not ( w_23456 , w_23460 );
and ( \3479_b0 , \3102_b0 , w_23461 );
and ( w_23460 , w_23461 , w_23457 );
or ( w_23456 , \b[10]_b1 , w_23458 );
not ( w_23458 , w_23462 );
and ( w_23457 , \b[10]_b0 , w_23463 );
and ( w_23462 , w_23463 , w_23459 );
buf ( w_23458 , \c[10]_b1 );
not ( w_23458 , w_23464 );
not ( w_23459 , w_23465 );
and ( w_23464 , w_23465 , \c[10]_b0 );
or ( \3480_b1 , \3470_b1 , w_23466 );
not ( w_23466 , w_23470 );
and ( \3480_b0 , \3470_b0 , w_23471 );
and ( w_23470 , w_23471 , w_23467 );
or ( w_23466 , \3478_b1 , w_23468 );
not ( w_23468 , w_23472 );
and ( w_23467 , \3478_b0 , w_23473 );
and ( w_23472 , w_23473 , w_23469 );
buf ( w_23468 , \3479_b1 );
not ( w_23468 , w_23474 );
not ( w_23469 , w_23475 );
and ( w_23474 , w_23475 , \3479_b0 );
or ( \3493_b1 , \2205_b1 , w_23476 );
not ( w_23476 , w_23478 );
and ( \3493_b0 , \2205_b0 , w_23479 );
and ( w_23478 , w_23479 , w_23477 );
or ( w_23476 , \2112_b1 , \2206_b1 );
not ( \2206_b1 , w_23480 );
and ( w_23477 , \2112_b0 , w_23481 );
and ( w_23480 , w_23481 , \2206_b0 );
or ( \3514_b1 , \3513_b1 , w_23482 );
not ( w_23482 , w_23486 );
and ( \3514_b0 , \3513_b0 , w_23487 );
and ( w_23486 , w_23487 , w_23483 );
or ( w_23482 , \2910_b1 , w_23484 );
not ( w_23484 , w_23488 );
and ( w_23483 , \2910_b0 , w_23489 );
and ( w_23488 , w_23489 , w_23485 );
buf ( w_23484 , \2814_b1 );
not ( w_23484 , w_23490 );
not ( w_23485 , w_23491 );
and ( w_23490 , w_23491 , \2814_b0 );
or ( \3515_b1 , \3508_b1 , w_23492 );
not ( w_23492 , w_23496 );
and ( \3515_b0 , \3508_b0 , w_23497 );
and ( w_23496 , w_23497 , w_23493 );
or ( w_23492 , \3514_b1 , w_23494 );
not ( w_23494 , w_23498 );
and ( w_23493 , \3514_b0 , w_23499 );
and ( w_23498 , w_23499 , w_23495 );
buf ( w_23494 , \2926_b1 );
not ( w_23494 , w_23500 );
not ( w_23495 , w_23501 );
and ( w_23500 , w_23501 , \2926_b0 );
or ( \3534_b1 , \2979_b1 , w_23502 );
not ( w_23502 , w_23504 );
and ( \3534_b0 , \2979_b0 , w_23505 );
and ( w_23504 , w_23505 , w_23503 );
or ( w_23502 , \2992_b1 , \3533_b1 );
not ( \3533_b1 , w_23506 );
and ( w_23503 , \2992_b0 , w_23507 );
and ( w_23506 , w_23507 , \3533_b0 );
or ( \3547_b1 , \3041_b1 , w_23508 );
not ( w_23508 , w_23510 );
and ( \3547_b0 , \3041_b0 , w_23511 );
and ( w_23510 , w_23511 , w_23509 );
or ( w_23508 , \3054_b1 , \3546_b1 );
not ( \3546_b1 , w_23512 );
and ( w_23509 , \3054_b0 , w_23513 );
and ( w_23512 , w_23513 , \3546_b0 );
or ( \3575_b1 , \3566_b1 , w_23514 );
not ( w_23514 , w_23518 );
and ( \3575_b0 , \3566_b0 , w_23519 );
and ( w_23518 , w_23519 , w_23515 );
or ( w_23514 , \3567_b1 , w_23516 );
not ( w_23516 , w_23520 );
and ( w_23515 , \3567_b0 , w_23521 );
and ( w_23520 , w_23521 , w_23517 );
buf ( w_23516 , \3574_b1 );
not ( w_23516 , w_23522 );
not ( w_23517 , w_23523 );
and ( w_23522 , w_23523 , \3574_b0 );
or ( \3667_b1 , \3664_b1 , w_23528 );
or ( \3667_b0 , \3664_b0 , w_23525 );
not ( w_23525 , w_23529 );
and ( w_23529 , w_23528 , w_23524 );
or ( w_23524 , \3665_b1 , w_23530 );
or ( w_23525 , \3665_b0 , w_23527 );
not ( w_23527 , w_23531 );
and ( w_23531 , w_23530 , w_23526 );
buf ( w_23526 , \3666_b1 );
not ( w_23526 , w_23532 );
not ( w_23527 , w_23533 );
and ( w_23532 , w_23533 , \3666_b0 );
or ( \3676_b1 , \3671_b1 , w_23534 );
not ( w_23534 , w_23538 );
and ( \3676_b0 , \3671_b0 , w_23539 );
and ( w_23538 , w_23539 , w_23535 );
or ( w_23534 , \3673_b1 , w_23536 );
not ( w_23536 , w_23540 );
and ( w_23535 , \3673_b0 , w_23541 );
and ( w_23540 , w_23541 , w_23537 );
buf ( w_23536 , \3675_b1 );
not ( w_23536 , w_23542 );
not ( w_23537 , w_23543 );
and ( w_23542 , w_23543 , \3675_b0 );
or ( \3738_b1 , \3735_b1 , w_23548 );
or ( \3738_b0 , \3735_b0 , w_23545 );
not ( w_23545 , w_23549 );
and ( w_23549 , w_23548 , w_23544 );
or ( w_23544 , \3736_b1 , w_23550 );
or ( w_23545 , \3736_b0 , w_23547 );
not ( w_23547 , w_23551 );
and ( w_23551 , w_23550 , w_23546 );
buf ( w_23546 , \3737_b1 );
not ( w_23546 , w_23552 );
not ( w_23547 , w_23553 );
and ( w_23552 , w_23553 , \3737_b0 );
or ( \3743_b1 , \3708_b1 , w_23554 );
not ( w_23554 , w_23558 );
and ( \3743_b0 , \3708_b0 , w_23559 );
and ( w_23558 , w_23559 , w_23555 );
or ( w_23554 , \3710_b1 , w_23556 );
not ( w_23556 , w_23560 );
and ( w_23555 , \3710_b0 , w_23561 );
and ( w_23560 , w_23561 , w_23557 );
buf ( w_23556 , \3742_b1 );
not ( w_23556 , w_23562 );
not ( w_23557 , w_23563 );
and ( w_23562 , w_23563 , \3742_b0 );
or ( \3818_b1 , \3769_b1 , w_23564 );
not ( w_23564 , w_23568 );
and ( \3818_b0 , \3769_b0 , w_23569 );
and ( w_23568 , w_23569 , w_23565 );
or ( w_23564 , \3770_b1 , w_23566 );
not ( w_23566 , w_23570 );
and ( w_23565 , \3770_b0 , w_23571 );
and ( w_23570 , w_23571 , w_23567 );
buf ( w_23566 , \3817_b1 );
not ( w_23566 , w_23572 );
not ( w_23567 , w_23573 );
and ( w_23572 , w_23573 , \3817_b0 );
or ( \3873_b1 , \3870_b1 , w_23578 );
or ( \3873_b0 , \3870_b0 , w_23575 );
not ( w_23575 , w_23579 );
and ( w_23579 , w_23578 , w_23574 );
or ( w_23574 , \3871_b1 , w_23580 );
or ( w_23575 , \3871_b0 , w_23577 );
not ( w_23577 , w_23581 );
and ( w_23581 , w_23580 , w_23576 );
buf ( w_23576 , \3872_b1 );
not ( w_23576 , w_23582 );
not ( w_23577 , w_23583 );
and ( w_23582 , w_23583 , \3872_b0 );
or ( \3890_b1 , \3887_b1 , w_23588 );
or ( \3890_b0 , \3887_b0 , w_23585 );
not ( w_23585 , w_23589 );
and ( w_23589 , w_23588 , w_23584 );
or ( w_23584 , \3888_b1 , w_23590 );
or ( w_23585 , \3888_b0 , w_23587 );
not ( w_23587 , w_23591 );
and ( w_23591 , w_23590 , w_23586 );
buf ( w_23586 , \3889_b1 );
not ( w_23586 , w_23592 );
not ( w_23587 , w_23593 );
and ( w_23592 , w_23593 , \3889_b0 );
or ( \3894_b1 , \3891_b1 , w_23594 );
not ( w_23594 , w_23598 );
and ( \3894_b0 , \3891_b0 , w_23599 );
and ( w_23598 , w_23599 , w_23595 );
or ( w_23594 , \3892_b1 , w_23596 );
not ( w_23596 , w_23600 );
and ( w_23595 , \3892_b0 , w_23601 );
and ( w_23600 , w_23601 , w_23597 );
buf ( w_23596 , \3893_b1 );
not ( w_23596 , w_23602 );
not ( w_23597 , w_23603 );
and ( w_23602 , w_23603 , \3893_b0 );
or ( \3903_b1 , \3894_b1 , w_23604 );
not ( w_23604 , w_23610 );
and ( \3903_b0 , \3894_b0 , w_23611 );
and ( w_23610 , w_23611 , w_23605 );
or ( w_23604 , \3897_b1 , w_23606 );
not ( w_23606 , w_23612 );
and ( w_23605 , \3897_b0 , w_23613 );
and ( w_23612 , w_23613 , w_23607 );
or ( w_23606 , \3900_b1 , w_23608 );
not ( w_23608 , w_23614 );
and ( w_23607 , \3900_b0 , w_23615 );
and ( w_23614 , w_23615 , w_23609 );
buf ( w_23608 , \3902_b1 );
not ( w_23608 , w_23616 );
not ( w_23609 , w_23617 );
and ( w_23616 , w_23617 , \3902_b0 );
or ( \3909_b1 , \3906_b1 , w_23618 );
not ( w_23618 , w_23622 );
and ( \3909_b0 , \3906_b0 , w_23623 );
and ( w_23622 , w_23623 , w_23619 );
or ( w_23618 , \3907_b1 , w_23620 );
not ( w_23620 , w_23624 );
and ( w_23619 , \3907_b0 , w_23625 );
and ( w_23624 , w_23625 , w_23621 );
buf ( w_23620 , \3908_b1 );
not ( w_23620 , w_23626 );
not ( w_23621 , w_23627 );
and ( w_23626 , w_23627 , \3908_b0 );
or ( \3925_b1 , \3914_b1 , w_23628 );
not ( w_23628 , w_23630 );
and ( \3925_b0 , \3914_b0 , w_23631 );
and ( w_23630 , w_23631 , w_23629 );
or ( w_23628 , \3921_b1 , \3924_b1 );
not ( \3924_b1 , w_23632 );
and ( w_23629 , \3921_b0 , w_23633 );
and ( w_23632 , w_23633 , \3924_b0 );
or ( \3939_b1 , \3932_b1 , w_23634 );
not ( w_23634 , w_23638 );
and ( \3939_b0 , \3932_b0 , w_23639 );
and ( w_23638 , w_23639 , w_23635 );
or ( w_23634 , \3937_b1 , w_23636 );
not ( w_23636 , w_23640 );
and ( w_23635 , \3937_b0 , w_23641 );
and ( w_23640 , w_23641 , w_23637 );
buf ( w_23636 , \3938_b1 );
not ( w_23636 , w_23642 );
not ( w_23637 , w_23643 );
and ( w_23642 , w_23643 , \3938_b0 );
or ( \3967_b1 , \3914_b1 , w_23644 );
not ( w_23644 , w_23646 );
and ( \3967_b0 , \3914_b0 , w_23647 );
and ( w_23646 , w_23647 , w_23645 );
or ( w_23644 , \3921_b1 , \3966_b1 );
not ( \3966_b1 , w_23648 );
and ( w_23645 , \3921_b0 , w_23649 );
and ( w_23648 , w_23649 , \3966_b0 );
or ( \3977_b1 , \3914_b1 , w_23650 );
not ( w_23650 , w_23652 );
and ( \3977_b0 , \3914_b0 , w_23653 );
and ( w_23652 , w_23653 , w_23651 );
or ( w_23650 , \3921_b1 , \3976_b1 );
not ( \3976_b1 , w_23654 );
and ( w_23651 , \3921_b0 , w_23655 );
and ( w_23654 , w_23655 , \3976_b0 );
or ( \3981_b1 , \3978_b1 , w_23656 );
not ( w_23656 , w_23660 );
and ( \3981_b0 , \3978_b0 , w_23661 );
and ( w_23660 , w_23661 , w_23657 );
or ( w_23656 , \3980_b1 , w_23658 );
not ( w_23658 , w_23662 );
and ( w_23657 , \3980_b0 , w_23663 );
and ( w_23662 , w_23663 , w_23659 );
buf ( w_23658 , \3883_b1 );
not ( w_23658 , w_23664 );
not ( w_23659 , w_23665 );
and ( w_23664 , w_23665 , \3883_b0 );
or ( \3987_b1 , \3972_b1 , w_23668 );
or ( \3987_b0 , \3972_b0 , w_23667 );
not ( w_23667 , w_23669 );
and ( w_23669 , w_23668 , w_23666 );
or ( w_23666 , \3983_b1 , w_23670 );
or ( w_23667 , \3983_b0 , \3986_b0 );
not ( \3986_b0 , w_23671 );
and ( w_23671 , w_23670 , \3986_b1 );
or ( \3993_b1 , \3988_b1 , w_23676 );
or ( \3993_b0 , \3988_b0 , w_23673 );
not ( w_23673 , w_23677 );
and ( w_23677 , w_23676 , w_23672 );
or ( w_23672 , \3989_b1 , w_23678 );
or ( w_23673 , \3989_b0 , w_23675 );
not ( w_23675 , w_23679 );
and ( w_23679 , w_23678 , w_23674 );
buf ( w_23674 , \3992_b1 );
not ( w_23674 , w_23680 );
not ( w_23675 , w_23681 );
and ( w_23680 , w_23681 , \3992_b0 );
or ( \3996_b1 , \3914_b1 , w_23682 );
not ( w_23682 , w_23684 );
and ( \3996_b0 , \3914_b0 , w_23685 );
and ( w_23684 , w_23685 , w_23683 );
or ( w_23682 , \3920_b1 , \3995_b1 );
not ( \3995_b1 , w_23686 );
and ( w_23683 , \3920_b0 , w_23687 );
and ( w_23686 , w_23687 , \3995_b0 );
or ( \4016_b1 , \4014_b1 , w_23688 );
not ( w_23688 , w_23692 );
and ( \4016_b0 , \4014_b0 , w_23693 );
and ( w_23692 , w_23693 , w_23689 );
or ( w_23688 , \4015_b1 , w_23690 );
not ( w_23690 , w_23694 );
and ( w_23689 , \4015_b0 , w_23695 );
and ( w_23694 , w_23695 , w_23691 );
buf ( w_23690 , \3906_b1 );
not ( w_23690 , w_23696 );
not ( w_23691 , w_23697 );
and ( w_23696 , w_23697 , \3906_b0 );
or ( \4928_b1 , \4836_b1 , w_23698 );
not ( w_23698 , w_23702 );
and ( \4928_b0 , \4836_b0 , w_23703 );
and ( w_23702 , w_23703 , w_23699 );
or ( w_23698 , \4885_b1 , w_23700 );
not ( w_23700 , w_23704 );
and ( w_23699 , \4885_b0 , w_23705 );
and ( w_23704 , w_23705 , w_23701 );
buf ( w_23700 , \4927_b1 );
not ( w_23700 , w_23706 );
not ( w_23701 , w_23707 );
and ( w_23706 , w_23707 , \4927_b0 );
or ( \4984_b1 , \4928_b1 , w_23712 );
or ( \4984_b0 , \4928_b0 , w_23709 );
not ( w_23709 , w_23713 );
and ( w_23713 , w_23712 , w_23708 );
or ( w_23708 , \4960_b1 , w_23714 );
or ( w_23709 , \4960_b0 , w_23711 );
not ( w_23711 , w_23715 );
and ( w_23715 , w_23714 , w_23710 );
buf ( w_23710 , \4983_b1 );
not ( w_23710 , w_23716 );
not ( w_23711 , w_23717 );
and ( w_23716 , w_23717 , \4983_b0 );
or ( \5423_b1 , \4063_b1 , w_23718 );
not ( w_23718 , w_23722 );
and ( \5423_b0 , \4063_b0 , w_23723 );
and ( w_23722 , w_23723 , w_23719 );
or ( w_23718 , \4053_b1 , w_23720 );
not ( w_23720 , w_23724 );
and ( w_23719 , \4053_b0 , w_23725 );
and ( w_23724 , w_23725 , w_23721 );
buf ( w_23720 , \5422_b1 );
not ( w_23720 , w_23726 );
not ( w_23721 , w_23727 );
and ( w_23726 , w_23727 , \5422_b0 );
or ( \5461_b1 , \5460_b1 , w_23728 );
not ( w_23728 , w_23732 );
and ( \5461_b0 , \5460_b0 , w_23733 );
and ( w_23732 , w_23733 , w_23729 );
or ( w_23728 , \4252_b1 , w_23730 );
not ( w_23730 , w_23734 );
and ( w_23729 , \4252_b0 , w_23735 );
and ( w_23734 , w_23735 , w_23731 );
buf ( w_23730 , \4251_b1 );
not ( w_23730 , w_23736 );
not ( w_23731 , w_23737 );
and ( w_23736 , w_23737 , \4251_b0 );
or ( \5574_b1 , \5572_b1 , w_23738 );
not ( w_23738 , w_23740 );
and ( \5574_b0 , \5572_b0 , w_23741 );
and ( w_23740 , w_23741 , w_23739 );
or ( w_23738 , \4156_b1 , \5573_b1 );
not ( \5573_b1 , w_23742 );
and ( w_23739 , \4156_b0 , w_23743 );
and ( w_23742 , w_23743 , \5573_b0 );
or ( \6071_b1 , \6069_b1 , w_23744 );
not ( w_23744 , w_23746 );
and ( \6071_b0 , \6069_b0 , w_23747 );
and ( w_23746 , w_23747 , w_23745 );
or ( w_23744 , \4172_b1 , \6070_b1 );
not ( \6070_b1 , w_23748 );
and ( w_23745 , \4172_b0 , w_23749 );
and ( w_23748 , w_23749 , \6070_b0 );
or ( \6251_b1 , \6246_b1 , w_23750 );
not ( w_23750 , w_23754 );
and ( \6251_b0 , \6246_b0 , w_23755 );
and ( w_23754 , w_23755 , w_23751 );
or ( w_23750 , \6250_b1 , w_23752 );
not ( w_23752 , w_23756 );
and ( w_23751 , \6250_b0 , w_23757 );
and ( w_23756 , w_23757 , w_23753 );
buf ( w_23752 , \4134_b1 );
not ( w_23752 , w_23758 );
not ( w_23753 , w_23759 );
and ( w_23758 , w_23759 , \4134_b0 );
or ( \6595_b1 , \6593_b1 , w_23760 );
not ( w_23760 , w_23764 );
and ( \6595_b0 , \6593_b0 , w_23765 );
and ( w_23764 , w_23765 , w_23761 );
or ( w_23760 , \4070_b1 , w_23762 );
not ( w_23762 , w_23766 );
and ( w_23761 , \4070_b0 , w_23767 );
and ( w_23766 , w_23767 , w_23763 );
buf ( w_23762 , \6594_b1 );
not ( w_23762 , w_23768 );
not ( w_23763 , w_23769 );
and ( w_23768 , w_23769 , \6594_b0 );
or ( \6674_b1 , \6667_b1 , w_23770 );
not ( w_23770 , w_23774 );
and ( \6674_b0 , \6667_b0 , w_23775 );
and ( w_23774 , w_23775 , w_23771 );
or ( w_23770 , \6669_b1 , w_23772 );
not ( w_23772 , w_23776 );
and ( w_23771 , \6669_b0 , w_23777 );
and ( w_23776 , w_23777 , w_23773 );
buf ( w_23772 , \6673_b1 );
not ( w_23772 , w_23778 );
not ( w_23773 , w_23779 );
and ( w_23778 , w_23779 , \6673_b0 );
or ( \6759_b1 , \6650_b1 , w_23780 );
not ( w_23780 , w_23784 );
and ( \6759_b0 , \6650_b0 , w_23785 );
and ( w_23784 , w_23785 , w_23781 );
or ( w_23780 , \6749_b1 , w_23782 );
not ( w_23782 , w_23786 );
and ( w_23781 , \6749_b0 , w_23787 );
and ( w_23786 , w_23787 , w_23783 );
buf ( w_23782 , \6758_b1 );
not ( w_23782 , w_23788 );
not ( w_23783 , w_23789 );
and ( w_23788 , w_23789 , \6758_b0 );
or ( \6763_b1 , \6759_b1 , w_23790 );
not ( w_23790 , w_23794 );
and ( \6763_b0 , \6759_b0 , w_23795 );
and ( w_23794 , w_23795 , w_23791 );
or ( w_23790 , \6761_b1 , w_23792 );
not ( w_23792 , w_23796 );
and ( w_23791 , \6761_b0 , w_23797 );
and ( w_23796 , w_23797 , w_23793 );
buf ( w_23792 , \6762_b1 );
not ( w_23792 , w_23798 );
not ( w_23793 , w_23799 );
and ( w_23798 , w_23799 , \6762_b0 );
or ( \6768_b1 , \6574_b1 , w_23800 );
not ( w_23800 , w_23804 );
and ( \6768_b0 , \6574_b0 , w_23805 );
and ( w_23804 , w_23805 , w_23801 );
or ( w_23800 , \6767_b1 , w_23802 );
not ( w_23802 , w_23806 );
and ( w_23801 , \6767_b0 , w_23807 );
and ( w_23806 , w_23807 , w_23803 );
buf ( w_23802 , \6387_b1 );
not ( w_23802 , w_23808 );
not ( w_23803 , w_23809 );
and ( w_23808 , w_23809 , \6387_b0 );
or ( \6813_b1 , \6198_b1 , w_23810 );
not ( w_23810 , w_23814 );
and ( \6813_b0 , \6198_b0 , w_23815 );
and ( w_23814 , w_23815 , w_23811 );
or ( w_23810 , \6769_b1 , w_23812 );
not ( w_23812 , w_23816 );
and ( w_23811 , \6769_b0 , w_23817 );
and ( w_23816 , w_23817 , w_23813 );
buf ( w_23812 , \6812_b1 );
not ( w_23812 , w_23818 );
not ( w_23813 , w_23819 );
and ( w_23818 , w_23819 , \6812_b0 );
or ( \6829_b1 , \6822_b1 , w_23820 );
not ( w_23820 , w_23824 );
and ( \6829_b0 , \6822_b0 , w_23825 );
and ( w_23824 , w_23825 , w_23821 );
or ( w_23820 , \6828_b1 , w_23822 );
not ( w_23822 , w_23826 );
and ( w_23821 , \6828_b0 , w_23827 );
and ( w_23826 , w_23827 , w_23823 );
buf ( w_23822 , \6816_b1 );
not ( w_23822 , w_23828 );
not ( w_23823 , w_23829 );
and ( w_23828 , w_23829 , \6816_b0 );
or ( \6877_b1 , \5745_b1 , w_23830 );
not ( w_23830 , w_23834 );
and ( \6877_b0 , \5745_b0 , w_23835 );
and ( w_23834 , w_23835 , w_23831 );
or ( w_23830 , \6831_b1 , w_23832 );
not ( w_23832 , w_23836 );
and ( w_23831 , \6831_b0 , w_23837 );
and ( w_23836 , w_23837 , w_23833 );
buf ( w_23832 , \6876_b1 );
not ( w_23832 , w_23838 );
not ( w_23833 , w_23839 );
and ( w_23838 , w_23839 , \6876_b0 );
or ( \6888_b1 , \6877_b1 , w_23840 );
not ( w_23840 , w_23844 );
and ( \6888_b0 , \6877_b0 , w_23845 );
and ( w_23844 , w_23845 , w_23841 );
or ( w_23840 , \6882_b1 , w_23842 );
not ( w_23842 , w_23846 );
and ( w_23841 , \6882_b0 , w_23847 );
and ( w_23846 , w_23847 , w_23843 );
buf ( w_23842 , \6887_b1 );
not ( w_23842 , w_23848 );
not ( w_23843 , w_23849 );
and ( w_23848 , w_23849 , \6887_b0 );
or ( \6916_b1 , \6913_b1 , w_23850 );
not ( w_23850 , w_23852 );
and ( \6916_b0 , \6913_b0 , w_23853 );
and ( w_23852 , w_23853 , w_23851 );
or ( w_23850 , \6914_b1 , \6915_b1 );
not ( \6915_b1 , w_23854 );
and ( w_23851 , \6914_b0 , w_23855 );
and ( w_23854 , w_23855 , \6915_b0 );
or ( \7051_b1 , \7049_b1 , w_23856 );
not ( w_23856 , w_23860 );
and ( \7051_b0 , \7049_b0 , w_23861 );
and ( w_23860 , w_23861 , w_23857 );
or ( w_23856 , \7050_b1 , w_23858 );
not ( w_23858 , w_23862 );
and ( w_23857 , \7050_b0 , w_23863 );
and ( w_23862 , w_23863 , w_23859 );
buf ( w_23858 , \5560_b1 );
not ( w_23858 , w_23864 );
not ( w_23859 , w_23865 );
and ( w_23864 , w_23865 , \5560_b0 );
or ( \7055_b1 , \7051_b1 , w_23866 );
not ( w_23866 , w_23870 );
and ( \7055_b0 , \7051_b0 , w_23871 );
and ( w_23870 , w_23871 , w_23867 );
or ( w_23866 , \7053_b1 , w_23868 );
not ( w_23868 , w_23872 );
and ( w_23867 , \7053_b0 , w_23873 );
and ( w_23872 , w_23873 , w_23869 );
buf ( w_23868 , \7054_b1 );
not ( w_23868 , w_23874 );
not ( w_23869 , w_23875 );
and ( w_23874 , w_23875 , \7054_b0 );
endmodule

