// ...
module top(\A[0][9]_b1 ,\A[0][9]_b0 ,\A[0][8]_b1 ,\A[0][8]_b0 ,\A[0][7]_b1 ,\A[0][7]_b0 ,\A[0][6]_b1 ,\A[0][6]_b0 ,\A[0][5]_b1 ,
		\A[0][5]_b0 ,\A[0][4]_b1 ,\A[0][4]_b0 ,\A[0][3]_b1 ,\A[0][3]_b0 ,\A[0][2]_b1 ,\A[0][2]_b0 ,\A[0][1]_b1 ,\A[0][1]_b0 ,
		\A[0][0]_b1 ,\A[0][0]_b0 ,\A[1][9]_b1 ,\A[1][9]_b0 ,\A[1][8]_b1 ,\A[1][8]_b0 ,\A[1][7]_b1 ,\A[1][7]_b0 ,\A[1][6]_b1 ,
		\A[1][6]_b0 ,\A[1][5]_b1 ,\A[1][5]_b0 ,\A[1][4]_b1 ,\A[1][4]_b0 ,\A[1][3]_b1 ,\A[1][3]_b0 ,\A[1][2]_b1 ,\A[1][2]_b0 ,
		\A[1][1]_b1 ,\A[1][1]_b0 ,\A[1][0]_b1 ,\A[1][0]_b0 ,\A[2][9]_b1 ,\A[2][9]_b0 ,\A[2][8]_b1 ,\A[2][8]_b0 ,\A[2][7]_b1 ,
		\A[2][7]_b0 ,\A[2][6]_b1 ,\A[2][6]_b0 ,\A[2][5]_b1 ,\A[2][5]_b0 ,\A[2][4]_b1 ,\A[2][4]_b0 ,\A[2][3]_b1 ,\A[2][3]_b0 ,
		\A[2][2]_b1 ,\A[2][2]_b0 ,\A[2][1]_b1 ,\A[2][1]_b0 ,\A[2][0]_b1 ,\A[2][0]_b0 ,\B[9]_b1 ,\B[9]_b0 ,\B[8]_b1 ,
		\B[8]_b0 ,\B[7]_b1 ,\B[7]_b0 ,\B[6]_b1 ,\B[6]_b0 ,\B[5]_b1 ,\B[5]_b0 ,\B[4]_b1 ,\B[4]_b0 ,
		\B[3]_b1 ,\B[3]_b0 ,\B[2]_b1 ,\B[2]_b0 ,\B[1]_b1 ,\B[1]_b0 ,\B[0]_b1 ,\B[0]_b0 ,\I[7]_b1 ,
		\I[7]_b0 ,\I[6]_b1 ,\I[6]_b0 ,\I[5]_b1 ,\I[5]_b0 ,\I[4]_b1 ,\I[4]_b0 ,\I[3]_b1 ,\I[3]_b0 ,
		\I[2]_b1 ,\I[2]_b0 ,\I[1]_b1 ,\I[1]_b0 ,\I[0]_b1 ,\I[0]_b0 ,\O[19]_b1 ,\O[19]_b0 ,\O[18]_b1 ,
		\O[18]_b0 ,\O[17]_b1 ,\O[17]_b0 ,\O[16]_b1 ,\O[16]_b0 ,\O[15]_b1 ,\O[15]_b0 ,\O[14]_b1 ,\O[14]_b0 ,
		\O[13]_b1 ,\O[13]_b0 ,\O[12]_b1 ,\O[12]_b0 ,\O[11]_b1 ,\O[11]_b0 ,\O[10]_b1 ,\O[10]_b0 ,\O[9]_b1 ,
		\O[9]_b0 ,\O[8]_b1 ,\O[8]_b0 ,\O[7]_b1 ,\O[7]_b0 ,\O[6]_b1 ,\O[6]_b0 ,\O[5]_b1 ,\O[5]_b0 ,
		\O[4]_b1 ,\O[4]_b0 ,\O[3]_b1 ,\O[3]_b0 ,\O[2]_b1 ,\O[2]_b0 ,\O[1]_b1 ,\O[1]_b0 ,\O[0]_b1 ,
		\O[0]_b0 );
input \A[0][9]_b1 ,\A[0][9]_b0 ,\A[0][8]_b1 ,\A[0][8]_b0 ,\A[0][7]_b1 ,\A[0][7]_b0 ,\A[0][6]_b1 ,\A[0][6]_b0 ,\A[0][5]_b1 ,
		\A[0][5]_b0 ,\A[0][4]_b1 ,\A[0][4]_b0 ,\A[0][3]_b1 ,\A[0][3]_b0 ,\A[0][2]_b1 ,\A[0][2]_b0 ,\A[0][1]_b1 ,\A[0][1]_b0 ,
		\A[0][0]_b1 ,\A[0][0]_b0 ,\A[1][9]_b1 ,\A[1][9]_b0 ,\A[1][8]_b1 ,\A[1][8]_b0 ,\A[1][7]_b1 ,\A[1][7]_b0 ,\A[1][6]_b1 ,
		\A[1][6]_b0 ,\A[1][5]_b1 ,\A[1][5]_b0 ,\A[1][4]_b1 ,\A[1][4]_b0 ,\A[1][3]_b1 ,\A[1][3]_b0 ,\A[1][2]_b1 ,\A[1][2]_b0 ,
		\A[1][1]_b1 ,\A[1][1]_b0 ,\A[1][0]_b1 ,\A[1][0]_b0 ,\A[2][9]_b1 ,\A[2][9]_b0 ,\A[2][8]_b1 ,\A[2][8]_b0 ,\A[2][7]_b1 ,
		\A[2][7]_b0 ,\A[2][6]_b1 ,\A[2][6]_b0 ,\A[2][5]_b1 ,\A[2][5]_b0 ,\A[2][4]_b1 ,\A[2][4]_b0 ,\A[2][3]_b1 ,\A[2][3]_b0 ,
		\A[2][2]_b1 ,\A[2][2]_b0 ,\A[2][1]_b1 ,\A[2][1]_b0 ,\A[2][0]_b1 ,\A[2][0]_b0 ,\B[9]_b1 ,\B[9]_b0 ,\B[8]_b1 ,
		\B[8]_b0 ,\B[7]_b1 ,\B[7]_b0 ,\B[6]_b1 ,\B[6]_b0 ,\B[5]_b1 ,\B[5]_b0 ,\B[4]_b1 ,\B[4]_b0 ,
		\B[3]_b1 ,\B[3]_b0 ,\B[2]_b1 ,\B[2]_b0 ,\B[1]_b1 ,\B[1]_b0 ,\B[0]_b1 ,\B[0]_b0 ,\I[7]_b1 ,
		\I[7]_b0 ,\I[6]_b1 ,\I[6]_b0 ,\I[5]_b1 ,\I[5]_b0 ,\I[4]_b1 ,\I[4]_b0 ,\I[3]_b1 ,\I[3]_b0 ,
		\I[2]_b1 ,\I[2]_b0 ,\I[1]_b1 ,\I[1]_b0 ,\I[0]_b1 ,\I[0]_b0 ;
output \O[19]_b1 ,\O[19]_b0 ,\O[18]_b1 ,\O[18]_b0 ,\O[17]_b1 ,\O[17]_b0 ,\O[16]_b1 ,\O[16]_b0 ,\O[15]_b1 ,
		\O[15]_b0 ,\O[14]_b1 ,\O[14]_b0 ,\O[13]_b1 ,\O[13]_b0 ,\O[12]_b1 ,\O[12]_b0 ,\O[11]_b1 ,\O[11]_b0 ,
		\O[10]_b1 ,\O[10]_b0 ,\O[9]_b1 ,\O[9]_b0 ,\O[8]_b1 ,\O[8]_b0 ,\O[7]_b1 ,\O[7]_b0 ,\O[6]_b1 ,
		\O[6]_b0 ,\O[5]_b1 ,\O[5]_b0 ,\O[4]_b1 ,\O[4]_b0 ,\O[3]_b1 ,\O[3]_b0 ,\O[2]_b1 ,\O[2]_b0 ,
		\O[1]_b1 ,\O[1]_b0 ,\O[0]_b1 ,\O[0]_b0 ;

wire \69_ZERO_b1 , \69_ZERO_b0 , \70_ONE_b1 , \70_ONE_b0 , \71_b1 , \71_b0 , \72_b1 , \72_b0 , \73_b1 , \73_b0 , 
		\74_b1 , \74_b0 , \75_b1 , \75_b0 , \76_b1 , \76_b0 , \77_b1 , \77_b0 , \78_b1 , \78_b0 , 
		\79_b1 , \79_b0 , \80_b1 , \80_b0 , \81_b1 , \81_b0 , \82_b1 , \82_b0 , \83_b1 , \83_b0 , 
		\84_b1 , \84_b0 , \85_b1 , \85_b0 , \86_b1 , \86_b0 , \87_b1 , \87_b0 , \88_b1 , \88_b0 , 
		\89_b1 , \89_b0 , \90_b1 , \90_b0 , \91_b1 , \91_b0 , \92_b1 , \92_b0 , \93_b1 , \93_b0 , 
		\94_b1 , \94_b0 , \95_b1 , \95_b0 , \96_b1 , \96_b0 , \97_b1 , \97_b0 , \98_b1 , \98_b0 , 
		\99_b1 , \99_b0 , \100_b1 , \100_b0 , \101_b1 , \101_b0 , \102_b1 , \102_b0 , \103_b1 , \103_b0 , 
		\104_b1 , \104_b0 , \105_b1 , \105_b0 , \106_b1 , \106_b0 , \107_b1 , \107_b0 , \108_b1 , \108_b0 , 
		\109_b1 , \109_b0 , \110_b1 , \110_b0 , \111_b1 , \111_b0 , \112_b1 , \112_b0 , \113_b1 , \113_b0 , 
		\114_b1 , \114_b0 , \115_b1 , \115_b0 , \116_b1 , \116_b0 , \117_b1 , \117_b0 , \118_b1 , \118_b0 , 
		\119_b1 , \119_b0 , \120_b1 , \120_b0 , \121_b1 , \121_b0 , \122_b1 , \122_b0 , \123_b1 , \123_b0 , 
		\124_b1 , \124_b0 , \125_b1 , \125_b0 , \126_b1 , \126_b0 , \127_b1 , \127_b0 , \128_b1 , \128_b0 , 
		\129_b1 , \129_b0 , \130_b1 , \130_b0 , \131_b1 , \131_b0 , \132_b1 , \132_b0 , \133_b1 , \133_b0 , 
		\134_b1 , \134_b0 , \135_b1 , \135_b0 , \136_b1 , \136_b0 , \137_b1 , \137_b0 , \138_b1 , \138_b0 , 
		\139_b1 , \139_b0 , \140_b1 , \140_b0 , \141_b1 , \141_b0 , \142_b1 , \142_b0 , \143_b1 , \143_b0 , 
		\144_b1 , \144_b0 , \145_b1 , \145_b0 , \146_b1 , \146_b0 , \147_b1 , \147_b0 , \148_b1 , \148_b0 , 
		\149_b1 , \149_b0 , \150_b1 , \150_b0 , \151_b1 , \151_b0 , \152_b1 , \152_b0 , \153_b1 , \153_b0 , 
		\154_b1 , \154_b0 , \155_b1 , \155_b0 , \156_b1 , \156_b0 , \157_b1 , \157_b0 , \158_b1 , \158_b0 , 
		\159_b1 , \159_b0 , \160_b1 , \160_b0 , \161_b1 , \161_b0 , \162_b1 , \162_b0 , \163_b1 , \163_b0 , 
		\164_b1 , \164_b0 , \165_b1 , \165_b0 , \166_b1 , \166_b0 , \167_b1 , \167_b0 , \168_b1 , \168_b0 , 
		\169_b1 , \169_b0 , \170_b1 , \170_b0 , \171_b1 , \171_b0 , \172_b1 , \172_b0 , \173_b1 , \173_b0 , 
		\174_b1 , \174_b0 , \175_b1 , \175_b0 , \176_b1 , \176_b0 , \177_b1 , \177_b0 , \178_b1 , \178_b0 , 
		\179_b1 , \179_b0 , \180_b1 , \180_b0 , \181_b1 , \181_b0 , \182_b1 , \182_b0 , \183_b1 , \183_b0 , 
		\184_b1 , \184_b0 , \185_b1 , \185_b0 , \186_b1 , \186_b0 , \187_b1 , \187_b0 , \188_b1 , \188_b0 , 
		\189_b1 , \189_b0 , \190_b1 , \190_b0 , \191_b1 , \191_b0 , \192_b1 , \192_b0 , \193_b1 , \193_b0 , 
		\194_b1 , \194_b0 , \195_b1 , \195_b0 , \196_b1 , \196_b0 , \197_b1 , \197_b0 , \198_b1 , \198_b0 , 
		\199_b1 , \199_b0 , \200_b1 , \200_b0 , \201_b1 , \201_b0 , \202_b1 , \202_b0 , \203_b1 , \203_b0 , 
		\204_b1 , \204_b0 , \205_b1 , \205_b0 , \206_b1 , \206_b0 , \207_b1 , \207_b0 , \208_b1 , \208_b0 , 
		\209_b1 , \209_b0 , \210_b1 , \210_b0 , \211_b1 , \211_b0 , \212_b1 , \212_b0 , \213_b1 , \213_b0 , 
		\214_b1 , \214_b0 , \215_b1 , \215_b0 , \216_b1 , \216_b0 , \217_b1 , \217_b0 , \218_b1 , \218_b0 , 
		\219_b1 , \219_b0 , \220_b1 , \220_b0 , \221_b1 , \221_b0 , \222_b1 , \222_b0 , \223_b1 , \223_b0 , 
		\224_b1 , \224_b0 , \225_b1 , \225_b0 , \226_b1 , \226_b0 , \227_b1 , \227_b0 , \228_b1 , \228_b0 , 
		\229_b1 , \229_b0 , \230_b1 , \230_b0 , \231_b1 , \231_b0 , \232_b1 , \232_b0 , \233_b1 , \233_b0 , 
		\234_b1 , \234_b0 , \235_b1 , \235_b0 , \236_b1 , \236_b0 , \237_b1 , \237_b0 , \238_b1 , \238_b0 , 
		\239_b1 , \239_b0 , \240_b1 , \240_b0 , \241_b1 , \241_b0 , \242_b1 , \242_b0 , \243_b1 , \243_b0 , 
		\244_b1 , \244_b0 , \245_b1 , \245_b0 , \246_b1 , \246_b0 , \247_b1 , \247_b0 , \248_b1 , \248_b0 , 
		\249_b1 , \249_b0 , \250_b1 , \250_b0 , \251_b1 , \251_b0 , \252_b1 , \252_b0 , \253_b1 , \253_b0 , 
		\254_b1 , \254_b0 , \255_b1 , \255_b0 , \256_b1 , \256_b0 , \257_b1 , \257_b0 , \258_b1 , \258_b0 , 
		\259_b1 , \259_b0 , \260_b1 , \260_b0 , \261_b1 , \261_b0 , \262_b1 , \262_b0 , \263_b1 , \263_b0 , 
		\264_b1 , \264_b0 , \265_b1 , \265_b0 , \266_b1 , \266_b0 , \267_b1 , \267_b0 , \268_b1 , \268_b0 , 
		\269_b1 , \269_b0 , \270_b1 , \270_b0 , \271_b1 , \271_b0 , \272_b1 , \272_b0 , \273_b1 , \273_b0 , 
		\274_b1 , \274_b0 , \275_b1 , \275_b0 , \276_b1 , \276_b0 , \277_b1 , \277_b0 , \278_b1 , \278_b0 , 
		\279_b1 , \279_b0 , \280_b1 , \280_b0 , \281_b1 , \281_b0 , \282_b1 , \282_b0 , \283_b1 , \283_b0 , 
		\284_b1 , \284_b0 , \285_b1 , \285_b0 , \286_b1 , \286_b0 , \287_b1 , \287_b0 , \288_b1 , \288_b0 , 
		\289_b1 , \289_b0 , \290_b1 , \290_b0 , \291_b1 , \291_b0 , \292_b1 , \292_b0 , \293_b1 , \293_b0 , 
		\294_b1 , \294_b0 , \295_b1 , \295_b0 , \296_b1 , \296_b0 , \297_b1 , \297_b0 , \298_b1 , \298_b0 , 
		\299_b1 , \299_b0 , \300_b1 , \300_b0 , \301_b1 , \301_b0 , \302_b1 , \302_b0 , \303_b1 , \303_b0 , 
		\304_b1 , \304_b0 , \305_b1 , \305_b0 , \306_b1 , \306_b0 , \307_b1 , \307_b0 , \308_b1 , \308_b0 , 
		\309_b1 , \309_b0 , \310_b1 , \310_b0 , \311_b1 , \311_b0 , \312_b1 , \312_b0 , \313_b1 , \313_b0 , 
		\314_b1 , \314_b0 , \315_b1 , \315_b0 , \316_b1 , \316_b0 , \317_b1 , \317_b0 , \318_b1 , \318_b0 , 
		\319_b1 , \319_b0 , \320_b1 , \320_b0 , \321_b1 , \321_b0 , \322_b1 , \322_b0 , \323_b1 , \323_b0 , 
		\324_b1 , \324_b0 , \325_b1 , \325_b0 , \326_b1 , \326_b0 , \327_b1 , \327_b0 , \328_b1 , \328_b0 , 
		\329_b1 , \329_b0 , \330_b1 , \330_b0 , \331_b1 , \331_b0 , \332_b1 , \332_b0 , \333_b1 , \333_b0 , 
		\334_b1 , \334_b0 , \335_b1 , \335_b0 , \336_b1 , \336_b0 , \337_b1 , \337_b0 , \338_b1 , \338_b0 , 
		\339_b1 , \339_b0 , \340_b1 , \340_b0 , \341_b1 , \341_b0 , \342_b1 , \342_b0 , \343_b1 , \343_b0 , 
		\344_b1 , \344_b0 , \345_b1 , \345_b0 , \346_b1 , \346_b0 , \347_b1 , \347_b0 , \348_b1 , \348_b0 , 
		\349_b1 , \349_b0 , \350_b1 , \350_b0 , \351_b1 , \351_b0 , \352_b1 , \352_b0 , \353_b1 , \353_b0 , 
		\354_b1 , \354_b0 , \355_b1 , \355_b0 , \356_b1 , \356_b0 , \357_b1 , \357_b0 , \358_b1 , \358_b0 , 
		\359_b1 , \359_b0 , \360_b1 , \360_b0 , \361_b1 , \361_b0 , \362_b1 , \362_b0 , \363_b1 , \363_b0 , 
		\364_b1 , \364_b0 , \365_b1 , \365_b0 , \366_b1 , \366_b0 , \367_b1 , \367_b0 , \368_b1 , \368_b0 , 
		\369_b1 , \369_b0 , \370_b1 , \370_b0 , \371_b1 , \371_b0 , \372_b1 , \372_b0 , \373_b1 , \373_b0 , 
		\374_b1 , \374_b0 , \375_b1 , \375_b0 , \376_b1 , \376_b0 , \377_b1 , \377_b0 , \378_b1 , \378_b0 , 
		\379_b1 , \379_b0 , \380_b1 , \380_b0 , \381_b1 , \381_b0 , \382_b1 , \382_b0 , \383_b1 , \383_b0 , 
		\384_b1 , \384_b0 , \385_b1 , \385_b0 , \386_b1 , \386_b0 , \387_b1 , \387_b0 , \388_b1 , \388_b0 , 
		\389_b1 , \389_b0 , \390_b1 , \390_b0 , \391_b1 , \391_b0 , \392_b1 , \392_b0 , \393_b1 , \393_b0 , 
		\394_b1 , \394_b0 , \395_b1 , \395_b0 , \396_b1 , \396_b0 , \397_b1 , \397_b0 , \398_b1 , \398_b0 , 
		\399_b1 , \399_b0 , \400_b1 , \400_b0 , \401_b1 , \401_b0 , \402_b1 , \402_b0 , \403_b1 , \403_b0 , 
		\404_b1 , \404_b0 , \405_b1 , \405_b0 , \406_b1 , \406_b0 , \407_b1 , \407_b0 , \408_b1 , \408_b0 , 
		\409_b1 , \409_b0 , \410_b1 , \410_b0 , \411_b1 , \411_b0 , \412_b1 , \412_b0 , \413_b1 , \413_b0 , 
		\414_b1 , \414_b0 , \415_b1 , \415_b0 , \416_b1 , \416_b0 , \417_b1 , \417_b0 , \418_b1 , \418_b0 , 
		\419_b1 , \419_b0 , \420_b1 , \420_b0 , \421_b1 , \421_b0 , \422_b1 , \422_b0 , \423_b1 , \423_b0 , 
		\424_b1 , \424_b0 , \425_b1 , \425_b0 , \426_b1 , \426_b0 , \427_b1 , \427_b0 , \428_b1 , \428_b0 , 
		\429_b1 , \429_b0 , \430_b1 , \430_b0 , \431_b1 , \431_b0 , \432_b1 , \432_b0 , \433_b1 , \433_b0 , 
		\434_b1 , \434_b0 , \435_b1 , \435_b0 , \436_b1 , \436_b0 , \437_b1 , \437_b0 , \438_b1 , \438_b0 , 
		\439_b1 , \439_b0 , \440_b1 , \440_b0 , \441_b1 , \441_b0 , \442_b1 , \442_b0 , \443_b1 , \443_b0 , 
		\444_b1 , \444_b0 , \445_b1 , \445_b0 , \446_b1 , \446_b0 , \447_b1 , \447_b0 , \448_b1 , \448_b0 , 
		\449_b1 , \449_b0 , \450_b1 , \450_b0 , \451_b1 , \451_b0 , \452_b1 , \452_b0 , \453_b1 , \453_b0 , 
		\454_b1 , \454_b0 , \455_b1 , \455_b0 , \456_b1 , \456_b0 , \457_b1 , \457_b0 , \458_b1 , \458_b0 , 
		\459_b1 , \459_b0 , \460_b1 , \460_b0 , \461_b1 , \461_b0 , \462_b1 , \462_b0 , \463_b1 , \463_b0 , 
		\464_b1 , \464_b0 , \465_b1 , \465_b0 , \466_b1 , \466_b0 , \467_b1 , \467_b0 , \468_b1 , \468_b0 , 
		\469_b1 , \469_b0 , \470_b1 , \470_b0 , \471_b1 , \471_b0 , \472_b1 , \472_b0 , \473_b1 , \473_b0 , 
		\474_b1 , \474_b0 , \475_b1 , \475_b0 , \476_b1 , \476_b0 , \477_b1 , \477_b0 , \478_b1 , \478_b0 , 
		\479_b1 , \479_b0 , \480_b1 , \480_b0 , \481_b1 , \481_b0 , \482_b1 , \482_b0 , \483_b1 , \483_b0 , 
		\484_b1 , \484_b0 , \485_b1 , \485_b0 , \486_b1 , \486_b0 , \487_b1 , \487_b0 , \488_b1 , \488_b0 , 
		\489_b1 , \489_b0 , \490_b1 , \490_b0 , \491_b1 , \491_b0 , \492_b1 , \492_b0 , \493_b1 , \493_b0 , 
		\494_b1 , \494_b0 , \495_b1 , \495_b0 , \496_b1 , \496_b0 , \497_b1 , \497_b0 , \498_b1 , \498_b0 , 
		\499_b1 , \499_b0 , \500_b1 , \500_b0 , \501_b1 , \501_b0 , \502_b1 , \502_b0 , \503_b1 , \503_b0 , 
		\504_b1 , \504_b0 , \505_b1 , \505_b0 , \506_b1 , \506_b0 , \507_b1 , \507_b0 , \508_b1 , \508_b0 , 
		\509_b1 , \509_b0 , \510_b1 , \510_b0 , \511_b1 , \511_b0 , \512_b1 , \512_b0 , \513_b1 , \513_b0 , 
		\514_b1 , \514_b0 , \515_b1 , \515_b0 , \516_b1 , \516_b0 , \517_b1 , \517_b0 , \518_b1 , \518_b0 , 
		\519_b1 , \519_b0 , \520_b1 , \520_b0 , \521_b1 , \521_b0 , \522_b1 , \522_b0 , \523_b1 , \523_b0 , 
		\524_b1 , \524_b0 , \525_b1 , \525_b0 , \526_b1 , \526_b0 , \527_b1 , \527_b0 , \528_b1 , \528_b0 , 
		\529_b1 , \529_b0 , \530_b1 , \530_b0 , \531_b1 , \531_b0 , \532_b1 , \532_b0 , \533_b1 , \533_b0 , 
		\534_b1 , \534_b0 , \535_b1 , \535_b0 , \536_b1 , \536_b0 , \537_b1 , \537_b0 , \538_b1 , \538_b0 , 
		\539_b1 , \539_b0 , \540_b1 , \540_b0 , \541_b1 , \541_b0 , \542_b1 , \542_b0 , \543_b1 , \543_b0 , 
		\544_b1 , \544_b0 , \545_b1 , \545_b0 , \546_b1 , \546_b0 , \547_b1 , \547_b0 , \548_b1 , \548_b0 , 
		\549_b1 , \549_b0 , \550_b1 , \550_b0 , \551_b1 , \551_b0 , \552_b1 , \552_b0 , \553_b1 , \553_b0 , 
		\554_b1 , \554_b0 , \555_b1 , \555_b0 , \556_b1 , \556_b0 , \557_b1 , \557_b0 , \558_b1 , \558_b0 , 
		\559_b1 , \559_b0 , \560_b1 , \560_b0 , \561_b1 , \561_b0 , \562_b1 , \562_b0 , \563_b1 , \563_b0 , 
		\564_b1 , \564_b0 , \565_b1 , \565_b0 , \566_b1 , \566_b0 , \567_b1 , \567_b0 , \568_b1 , \568_b0 , 
		\569_b1 , \569_b0 , \570_b1 , \570_b0 , \571_b1 , \571_b0 , \572_b1 , \572_b0 , \573_b1 , \573_b0 , 
		\574_b1 , \574_b0 , \575_b1 , \575_b0 , \576_b1 , \576_b0 , \577_b1 , \577_b0 , \578_b1 , \578_b0 , 
		\579_b1 , \579_b0 , \580_b1 , \580_b0 , \581_b1 , \581_b0 , \582_b1 , \582_b0 , \583_b1 , \583_b0 , 
		\584_b1 , \584_b0 , \585_b1 , \585_b0 , \586_b1 , \586_b0 , \587_b1 , \587_b0 , \588_b1 , \588_b0 , 
		\589_b1 , \589_b0 , \590_b1 , \590_b0 , \591_b1 , \591_b0 , \592_b1 , \592_b0 , \593_b1 , \593_b0 , 
		\594_b1 , \594_b0 , \595_b1 , \595_b0 , \596_b1 , \596_b0 , \597_b1 , \597_b0 , \598_b1 , \598_b0 , 
		\599_b1 , \599_b0 , \600_b1 , \600_b0 , \601_b1 , \601_b0 , \602_b1 , \602_b0 , \603_b1 , \603_b0 , 
		\604_b1 , \604_b0 , \605_b1 , \605_b0 , \606_b1 , \606_b0 , \607_b1 , \607_b0 , \608_b1 , \608_b0 , 
		\609_b1 , \609_b0 , \610_b1 , \610_b0 , \611_b1 , \611_b0 , \612_b1 , \612_b0 , \613_b1 , \613_b0 , 
		\614_b1 , \614_b0 , \615_b1 , \615_b0 , \616_b1 , \616_b0 , \617_b1 , \617_b0 , \618_b1 , \618_b0 , 
		\619_b1 , \619_b0 , \620_b1 , \620_b0 , \621_b1 , \621_b0 , \622_b1 , \622_b0 , \623_b1 , \623_b0 , 
		\624_b1 , \624_b0 , \625_b1 , \625_b0 , \626_b1 , \626_b0 , \627_b1 , \627_b0 , \628_b1 , \628_b0 , 
		\629_b1 , \629_b0 , \630_b1 , \630_b0 , \631_b1 , \631_b0 , \632_b1 , \632_b0 , \633_b1 , \633_b0 , 
		\634_b1 , \634_b0 , \635_b1 , \635_b0 , \636_b1 , \636_b0 , \637_b1 , \637_b0 , \638_b1 , \638_b0 , 
		\639_b1 , \639_b0 , \640_b1 , \640_b0 , \641_b1 , \641_b0 , \642_b1 , \642_b0 , \643_b1 , \643_b0 , 
		\644_b1 , \644_b0 , \645_b1 , \645_b0 , \646_b1 , \646_b0 , \647_b1 , \647_b0 , \648_b1 , \648_b0 , 
		\649_b1 , \649_b0 , \650_b1 , \650_b0 , \651_b1 , \651_b0 , \652_b1 , \652_b0 , \653_b1 , \653_b0 , 
		\654_b1 , \654_b0 , \655_b1 , \655_b0 , \656_b1 , \656_b0 , \657_b1 , \657_b0 , \658_b1 , \658_b0 , 
		\659_b1 , \659_b0 , \660_b1 , \660_b0 , \661_b1 , \661_b0 , \662_b1 , \662_b0 , \663_b1 , \663_b0 , 
		\664_b1 , \664_b0 , \665_b1 , \665_b0 , \666_b1 , \666_b0 , \667_b1 , \667_b0 , \668_b1 , \668_b0 , 
		\669_b1 , \669_b0 , \670_b1 , \670_b0 , \671_b1 , \671_b0 , \672_b1 , \672_b0 , \673_b1 , \673_b0 , 
		\674_b1 , \674_b0 , \675_b1 , \675_b0 , \676_b1 , \676_b0 , \677_b1 , \677_b0 , \678_b1 , \678_b0 , 
		\679_b1 , \679_b0 , \680_b1 , \680_b0 , \681_b1 , \681_b0 , \682_b1 , \682_b0 , \683_b1 , \683_b0 , 
		\684_b1 , \684_b0 , \685_b1 , \685_b0 , \686_b1 , \686_b0 , \687_b1 , \687_b0 , \688_b1 , \688_b0 , 
		\689_b1 , \689_b0 , \690_b1 , \690_b0 , \691_b1 , \691_b0 , \692_b1 , \692_b0 , \693_b1 , \693_b0 , 
		\694_b1 , \694_b0 , \695_b1 , \695_b0 , \696_b1 , \696_b0 , \697_b1 , \697_b0 , \698_b1 , \698_b0 , 
		\699_b1 , \699_b0 , \700_b1 , \700_b0 , \701_b1 , \701_b0 , \702_b1 , \702_b0 , \703_b1 , \703_b0 , 
		\704_b1 , \704_b0 , \705_b1 , \705_b0 , \706_b1 , \706_b0 , \707_b1 , \707_b0 , \708_b1 , \708_b0 , 
		\709_b1 , \709_b0 , \710_b1 , \710_b0 , \711_b1 , \711_b0 , \712_b1 , \712_b0 , \713_b1 , \713_b0 , 
		\714_b1 , \714_b0 , \715_b1 , \715_b0 , \716_b1 , \716_b0 , \717_b1 , \717_b0 , \718_b1 , \718_b0 , 
		\719_b1 , \719_b0 , \720_b1 , \720_b0 , \721_b1 , \721_b0 , \722_b1 , \722_b0 , \723_b1 , \723_b0 , 
		\724_b1 , \724_b0 , \725_b1 , \725_b0 , \726_b1 , \726_b0 , \727_b1 , \727_b0 , \728_b1 , \728_b0 , 
		\729_b1 , \729_b0 , \730_b1 , \730_b0 , \731_b1 , \731_b0 , \732_b1 , \732_b0 , \733_b1 , \733_b0 , 
		\734_b1 , \734_b0 , \735_b1 , \735_b0 , \736_b1 , \736_b0 , \737_b1 , \737_b0 , \738_b1 , \738_b0 , 
		\739_b1 , \739_b0 , \740_b1 , \740_b0 , \741_b1 , \741_b0 , \742_b1 , \742_b0 , \743_b1 , \743_b0 , 
		\744_b1 , \744_b0 , \745_b1 , \745_b0 , \746_b1 , \746_b0 , \747_b1 , \747_b0 , \748_b1 , \748_b0 , 
		\749_b1 , \749_b0 , \750_b1 , \750_b0 , \751_b1 , \751_b0 , \752_b1 , \752_b0 , \753_b1 , \753_b0 , 
		\754_b1 , \754_b0 , \755_b1 , \755_b0 , \756_b1 , \756_b0 , \757_b1 , \757_b0 , \758_b1 , \758_b0 , 
		\759_b1 , \759_b0 , \760_b1 , \760_b0 , \761_b1 , \761_b0 , \762_b1 , \762_b0 , \763_b1 , \763_b0 , 
		\764_b1 , \764_b0 , \765_b1 , \765_b0 , \766_b1 , \766_b0 , \767_b1 , \767_b0 , \768_b1 , \768_b0 , 
		\769_b1 , \769_b0 , \770_b1 , \770_b0 , \771_b1 , \771_b0 , \772_b1 , \772_b0 , \773_b1 , \773_b0 , 
		\774_b1 , \774_b0 , \775_b1 , \775_b0 , \776_b1 , \776_b0 , \777_b1 , \777_b0 , \778_b1 , \778_b0 , 
		\779_b1 , \779_b0 , \780_b1 , \780_b0 , \781_b1 , \781_b0 , \782_b1 , \782_b0 , \783_b1 , \783_b0 , 
		\784_b1 , \784_b0 , \785_b1 , \785_b0 , \786_b1 , \786_b0 , \787_b1 , \787_b0 , \788_b1 , \788_b0 , 
		\789_b1 , \789_b0 , \790_b1 , \790_b0 , \791_b1 , \791_b0 , \792_b1 , \792_b0 , \793_b1 , \793_b0 , 
		\794_b1 , \794_b0 , \795_b1 , \795_b0 , \796_b1 , \796_b0 , \797_b1 , \797_b0 , \798_b1 , \798_b0 , 
		\799_b1 , \799_b0 , \800_b1 , \800_b0 , \801_b1 , \801_b0 , \802_b1 , \802_b0 , \803_b1 , \803_b0 , 
		\804_b1 , \804_b0 , \805_b1 , \805_b0 , \806_b1 , \806_b0 , \807_b1 , \807_b0 , \808_b1 , \808_b0 , 
		\809_b1 , \809_b0 , \810_b1 , \810_b0 , \811_b1 , \811_b0 , \812_b1 , \812_b0 , \813_b1 , \813_b0 , 
		\814_b1 , \814_b0 , \815_b1 , \815_b0 , \816_b1 , \816_b0 , \817_b1 , \817_b0 , \818_b1 , \818_b0 , 
		\819_b1 , \819_b0 , \820_b1 , \820_b0 , \821_b1 , \821_b0 , \822_b1 , \822_b0 , \823_b1 , \823_b0 , 
		\824_b1 , \824_b0 , \825_b1 , \825_b0 , \826_b1 , \826_b0 , \827_b1 , \827_b0 , \828_b1 , \828_b0 , 
		\829_b1 , \829_b0 , \830_b1 , \830_b0 , \831_b1 , \831_b0 , \832_b1 , \832_b0 , \833_b1 , \833_b0 , 
		\834_b1 , \834_b0 , \835_b1 , \835_b0 , \836_b1 , \836_b0 , \837_b1 , \837_b0 , \838_b1 , \838_b0 , 
		\839_b1 , \839_b0 , \840_b1 , \840_b0 , \841_b1 , \841_b0 , \842_b1 , \842_b0 , \843_b1 , \843_b0 , 
		\844_b1 , \844_b0 , \845_b1 , \845_b0 , \846_b1 , \846_b0 , \847_b1 , \847_b0 , \848_b1 , \848_b0 , 
		\849_b1 , \849_b0 , \850_b1 , \850_b0 , \851_b1 , \851_b0 , \852_b1 , \852_b0 , \853_b1 , \853_b0 , 
		\854_b1 , \854_b0 , \855_b1 , \855_b0 , \856_b1 , \856_b0 , \857_b1 , \857_b0 , \858_b1 , \858_b0 , 
		\859_b1 , \859_b0 , \860_b1 , \860_b0 , \861_b1 , \861_b0 , \862_b1 , \862_b0 , \863_b1 , \863_b0 , 
		\864_b1 , \864_b0 , \865_b1 , \865_b0 , \866_b1 , \866_b0 , \867_b1 , \867_b0 , \868_b1 , \868_b0 , 
		\869_b1 , \869_b0 , \870_b1 , \870_b0 , \871_b1 , \871_b0 , \872_b1 , \872_b0 , \873_b1 , \873_b0 , 
		\874_b1 , \874_b0 , \875_b1 , \875_b0 , \876_b1 , \876_b0 , \877_b1 , \877_b0 , \878_b1 , \878_b0 , 
		\879_b1 , \879_b0 , \880_b1 , \880_b0 , \881_b1 , \881_b0 , \882_b1 , \882_b0 , \883_b1 , \883_b0 , 
		\884_b1 , \884_b0 , \885_b1 , \885_b0 , \886_b1 , \886_b0 , \887_b1 , \887_b0 , \888_b1 , \888_b0 , 
		\889_b1 , \889_b0 , \890_b1 , \890_b0 , \891_b1 , \891_b0 , \892_b1 , \892_b0 , \893_b1 , \893_b0 , 
		\894_b1 , \894_b0 , \895_b1 , \895_b0 , \896_b1 , \896_b0 , \897_b1 , \897_b0 , \898_b1 , \898_b0 , 
		\899_b1 , \899_b0 , \900_b1 , \900_b0 , \901_b1 , \901_b0 , \902_b1 , \902_b0 , \903_b1 , \903_b0 , 
		\904_b1 , \904_b0 , \905_b1 , \905_b0 , \906_b1 , \906_b0 , \907_b1 , \907_b0 , \908_b1 , \908_b0 , 
		\909_b1 , \909_b0 , \910_b1 , \910_b0 , \911_b1 , \911_b0 , \912_b1 , \912_b0 , \913_b1 , \913_b0 , 
		\914_b1 , \914_b0 , \915_b1 , \915_b0 , \916_b1 , \916_b0 , \917_b1 , \917_b0 , \918_b1 , \918_b0 , 
		\919_b1 , \919_b0 , \920_b1 , \920_b0 , \921_b1 , \921_b0 , \922_b1 , \922_b0 , \923_b1 , \923_b0 , 
		\924_b1 , \924_b0 , \925_b1 , \925_b0 , \926_b1 , \926_b0 , \927_b1 , \927_b0 , \928_b1 , \928_b0 , 
		\929_b1 , \929_b0 , \930_b1 , \930_b0 , \931_b1 , \931_b0 , \932_b1 , \932_b0 , \933_b1 , \933_b0 , 
		\934_b1 , \934_b0 , \935_b1 , \935_b0 , \936_b1 , \936_b0 , \937_b1 , \937_b0 , \938_b1 , \938_b0 , 
		\939_b1 , \939_b0 , \940_b1 , \940_b0 , \941_b1 , \941_b0 , \942_b1 , \942_b0 , \943_b1 , \943_b0 , 
		\944_b1 , \944_b0 , \945_b1 , \945_b0 , \946_b1 , \946_b0 , \947_b1 , \947_b0 , \948_b1 , \948_b0 , 
		\949_b1 , \949_b0 , \950_b1 , \950_b0 , \951_b1 , \951_b0 , \952_b1 , \952_b0 , \953_b1 , \953_b0 , 
		\954_b1 , \954_b0 , \955_b1 , \955_b0 , \956_b1 , \956_b0 , \957_b1 , \957_b0 , \958_b1 , \958_b0 , 
		\959_b1 , \959_b0 , \960_b1 , \960_b0 , \961_b1 , \961_b0 , \962_b1 , \962_b0 , \963_b1 , \963_b0 , 
		\964_b1 , \964_b0 , \965_b1 , \965_b0 , \966_b1 , \966_b0 , \967_b1 , \967_b0 , \968_b1 , \968_b0 , 
		\969_b1 , \969_b0 , \970_b1 , \970_b0 , \971_b1 , \971_b0 , \972_b1 , \972_b0 , \973_b1 , \973_b0 , 
		\974_b1 , \974_b0 , \975_b1 , \975_b0 , \976_b1 , \976_b0 , \977_b1 , \977_b0 , \978_b1 , \978_b0 , 
		\979_b1 , \979_b0 , \980_b1 , \980_b0 , \981_b1 , \981_b0 , \982_b1 , \982_b0 , \983_b1 , \983_b0 , 
		\984_b1 , \984_b0 , \985_b1 , \985_b0 , \986_b1 , \986_b0 , \987_b1 , \987_b0 , \988_b1 , \988_b0 , 
		\989_b1 , \989_b0 , \990_b1 , \990_b0 , \991_b1 , \991_b0 , \992_b1 , \992_b0 , \993_b1 , \993_b0 , 
		\994_b1 , \994_b0 , \995_b1 , \995_b0 , \996_b1 , \996_b0 , \997_b1 , \997_b0 , \998_b1 , \998_b0 , 
		\999_b1 , \999_b0 , \1000_b1 , \1000_b0 , \1001_b1 , \1001_b0 , \1002_b1 , \1002_b0 , \1003_b1 , \1003_b0 , 
		\1004_b1 , \1004_b0 , \1005_b1 , \1005_b0 , \1006_b1 , \1006_b0 , \1007_b1 , \1007_b0 , \1008_b1 , \1008_b0 , 
		\1009_b1 , \1009_b0 , \1010_b1 , \1010_b0 , \1011_b1 , \1011_b0 , \1012_b1 , \1012_b0 , \1013_b1 , \1013_b0 , 
		\1014_b1 , \1014_b0 , \1015_b1 , \1015_b0 , \1016_b1 , \1016_b0 , \1017_b1 , \1017_b0 , \1018_b1 , \1018_b0 , 
		\1019_b1 , \1019_b0 , \1020_b1 , \1020_b0 , \1021_b1 , \1021_b0 , \1022_b1 , \1022_b0 , \1023_b1 , \1023_b0 , 
		\1024_b1 , \1024_b0 , \1025_b1 , \1025_b0 , \1026_b1 , \1026_b0 , \1027_b1 , \1027_b0 , \1028_b1 , \1028_b0 , 
		\1029_b1 , \1029_b0 , \1030_b1 , \1030_b0 , \1031_b1 , \1031_b0 , \1032_b1 , \1032_b0 , \1033_b1 , \1033_b0 , 
		\1034_b1 , \1034_b0 , \1035_b1 , \1035_b0 , \1036_b1 , \1036_b0 , \1037_b1 , \1037_b0 , \1038_b1 , \1038_b0 , 
		\1039_b1 , \1039_b0 , \1040_b1 , \1040_b0 , \1041_b1 , \1041_b0 , \1042_b1 , \1042_b0 , \1043_b1 , \1043_b0 , 
		\1044_b1 , \1044_b0 , \1045_b1 , \1045_b0 , \1046_b1 , \1046_b0 , \1047_b1 , \1047_b0 , \1048_b1 , \1048_b0 , 
		\1049_b1 , \1049_b0 , \1050_b1 , \1050_b0 , \1051_b1 , \1051_b0 , \1052_b1 , \1052_b0 , \1053_b1 , \1053_b0 , 
		\1054_b1 , \1054_b0 , \1055_b1 , \1055_b0 , \1056_b1 , \1056_b0 , \1057_b1 , \1057_b0 , \1058_b1 , \1058_b0 , 
		\1059_b1 , \1059_b0 , \1060_b1 , \1060_b0 , \1061_b1 , \1061_b0 , \1062_b1 , \1062_b0 , \1063_b1 , \1063_b0 , 
		\1064_b1 , \1064_b0 , \1065_b1 , \1065_b0 , \1066_b1 , \1066_b0 , \1067_b1 , \1067_b0 , \1068_b1 , \1068_b0 , 
		\1069_b1 , \1069_b0 , w_0 , w_1 , w_2 , w_3 , w_4 , w_5 , w_6 , w_7 , 
		w_8 , w_9 , w_10 , w_11 , w_12 , w_13 , w_14 , w_15 , w_16 , w_17 , 
		w_18 , w_19 , w_20 , w_21 , w_22 , w_23 , w_24 , w_25 , w_26 , w_27 , 
		w_28 , w_29 , w_30 , w_31 , w_32 , w_33 , w_34 , w_35 , w_36 , w_37 , 
		w_38 , w_39 , w_40 , w_41 , w_42 , w_43 , w_44 , w_45 , w_46 , w_47 , 
		w_48 , w_49 , w_50 , w_51 , w_52 , w_53 , w_54 , w_55 , w_56 , w_57 , 
		w_58 , w_59 , w_60 , w_61 , w_62 , w_63 , w_64 , w_65 , w_66 , w_67 , 
		w_68 , w_69 , w_70 , w_71 , w_72 , w_73 , w_74 , w_75 , w_76 , w_77 , 
		w_78 , w_79 , w_80 , w_81 , w_82 , w_83 , w_84 , w_85 , w_86 , w_87 , 
		w_88 , w_89 , w_90 , w_91 , w_92 , w_93 , w_94 , w_95 , w_96 , w_97 , 
		w_98 , w_99 , w_100 , w_101 , w_102 , w_103 , w_104 , w_105 , w_106 , w_107 , 
		w_108 , w_109 , w_110 , w_111 , w_112 , w_113 , w_114 , w_115 , w_116 , w_117 , 
		w_118 , w_119 , w_120 , w_121 , w_122 , w_123 , w_124 , w_125 , w_126 , w_127 , 
		w_128 , w_129 , w_130 , w_131 , w_132 , w_133 , w_134 , w_135 , w_136 , w_137 , 
		w_138 , w_139 , w_140 , w_141 , w_142 , w_143 , w_144 , w_145 , w_146 , w_147 , 
		w_148 , w_149 , w_150 , w_151 , w_152 , w_153 , w_154 , w_155 , w_156 , w_157 , 
		w_158 , w_159 , w_160 , w_161 , w_162 , w_163 , w_164 , w_165 , w_166 , w_167 , 
		w_168 , w_169 , w_170 , w_171 , w_172 , w_173 , w_174 , w_175 , w_176 , w_177 , 
		w_178 , w_179 , w_180 , w_181 , w_182 , w_183 , w_184 , w_185 , w_186 , w_187 , 
		w_188 , w_189 , w_190 , w_191 , w_192 , w_193 , w_194 , w_195 , w_196 , w_197 , 
		w_198 , w_199 , w_200 , w_201 , w_202 , w_203 , w_204 , w_205 , w_206 , w_207 , 
		w_208 , w_209 , w_210 , w_211 , w_212 , w_213 , w_214 , w_215 , w_216 , w_217 , 
		w_218 , w_219 , w_220 , w_221 , w_222 , w_223 , w_224 , w_225 , w_226 , w_227 , 
		w_228 , w_229 , w_230 , w_231 , w_232 , w_233 , w_234 , w_235 , w_236 , w_237 , 
		w_238 , w_239 , w_240 , w_241 , w_242 , w_243 , w_244 , w_245 , w_246 , w_247 , 
		w_248 , w_249 , w_250 , w_251 , w_252 , w_253 , w_254 , w_255 , w_256 , w_257 , 
		w_258 , w_259 , w_260 , w_261 , w_262 , w_263 , w_264 , w_265 , w_266 , w_267 , 
		w_268 , w_269 , w_270 , w_271 , w_272 , w_273 , w_274 , w_275 , w_276 , w_277 , 
		w_278 , w_279 , w_280 , w_281 , w_282 , w_283 , w_284 , w_285 , w_286 , w_287 , 
		w_288 , w_289 , w_290 , w_291 , w_292 , w_293 , w_294 , w_295 , w_296 , w_297 , 
		w_298 , w_299 , w_300 , w_301 , w_302 , w_303 , w_304 , w_305 , w_306 , w_307 , 
		w_308 , w_309 , w_310 , w_311 , w_312 , w_313 , w_314 , w_315 , w_316 , w_317 , 
		w_318 , w_319 , w_320 , w_321 , w_322 , w_323 , w_324 , w_325 , w_326 , w_327 , 
		w_328 , w_329 , w_330 , w_331 , w_332 , w_333 , w_334 , w_335 , w_336 , w_337 , 
		w_338 , w_339 , w_340 , w_341 , w_342 , w_343 , w_344 , w_345 , w_346 , w_347 , 
		w_348 , w_349 , w_350 , w_351 , w_352 , w_353 , w_354 , w_355 , w_356 , w_357 , 
		w_358 , w_359 , w_360 , w_361 , w_362 , w_363 , w_364 , w_365 , w_366 , w_367 , 
		w_368 , w_369 , w_370 , w_371 , w_372 , w_373 , w_374 , w_375 , w_376 , w_377 , 
		w_378 , w_379 , w_380 , w_381 , w_382 , w_383 , w_384 , w_385 , w_386 , w_387 , 
		w_388 , w_389 , w_390 , w_391 , w_392 , w_393 , w_394 , w_395 , w_396 , w_397 , 
		w_398 , w_399 , w_400 , w_401 , w_402 , w_403 , w_404 , w_405 , w_406 , w_407 , 
		w_408 , w_409 , w_410 , w_411 , w_412 , w_413 , w_414 , w_415 , w_416 , w_417 , 
		w_418 , w_419 , w_420 , w_421 , w_422 , w_423 , w_424 , w_425 , w_426 , w_427 , 
		w_428 , w_429 , w_430 , w_431 , w_432 , w_433 , w_434 , w_435 , w_436 , w_437 , 
		w_438 , w_439 , w_440 , w_441 , w_442 , w_443 , w_444 , w_445 , w_446 , w_447 , 
		w_448 , w_449 , w_450 , w_451 , w_452 , w_453 , w_454 , w_455 , w_456 , w_457 , 
		w_458 , w_459 , w_460 , w_461 , w_462 , w_463 , w_464 , w_465 , w_466 , w_467 , 
		w_468 , w_469 , w_470 , w_471 , w_472 , w_473 , w_474 , w_475 , w_476 , w_477 , 
		w_478 , w_479 , w_480 , w_481 , w_482 , w_483 , w_484 , w_485 , w_486 , w_487 , 
		w_488 , w_489 , w_490 , w_491 , w_492 , w_493 , w_494 , w_495 , w_496 , w_497 , 
		w_498 , w_499 , w_500 , w_501 , w_502 , w_503 , w_504 , w_505 , w_506 , w_507 , 
		w_508 , w_509 , w_510 , w_511 , w_512 , w_513 , w_514 , w_515 , w_516 , w_517 , 
		w_518 , w_519 , w_520 , w_521 , w_522 , w_523 , w_524 , w_525 , w_526 , w_527 , 
		w_528 , w_529 , w_530 , w_531 , w_532 , w_533 , w_534 , w_535 , w_536 , w_537 , 
		w_538 , w_539 , w_540 , w_541 , w_542 , w_543 , w_544 , w_545 , w_546 , w_547 , 
		w_548 , w_549 , w_550 , w_551 , w_552 , w_553 , w_554 , w_555 , w_556 , w_557 , 
		w_558 , w_559 , w_560 , w_561 , w_562 , w_563 , w_564 , w_565 , w_566 , w_567 , 
		w_568 , w_569 , w_570 , w_571 , w_572 , w_573 , w_574 , w_575 , w_576 , w_577 , 
		w_578 , w_579 , w_580 , w_581 , w_582 , w_583 , w_584 , w_585 , w_586 , w_587 , 
		w_588 , w_589 , w_590 , w_591 , w_592 , w_593 , w_594 , w_595 , w_596 , w_597 , 
		w_598 , w_599 , w_600 , w_601 , w_602 , w_603 , w_604 , w_605 , w_606 , w_607 , 
		w_608 , w_609 , w_610 , w_611 , w_612 , w_613 , w_614 , w_615 , w_616 , w_617 , 
		w_618 , w_619 , w_620 , w_621 , w_622 , w_623 , w_624 , w_625 , w_626 , w_627 , 
		w_628 , w_629 , w_630 , w_631 , w_632 , w_633 , w_634 , w_635 , w_636 , w_637 , 
		w_638 , w_639 , w_640 , w_641 , w_642 , w_643 , w_644 , w_645 , w_646 , w_647 , 
		w_648 , w_649 , w_650 , w_651 , w_652 , w_653 , w_654 , w_655 , w_656 , w_657 , 
		w_658 , w_659 , w_660 , w_661 , w_662 , w_663 , w_664 , w_665 , w_666 , w_667 , 
		w_668 , w_669 , w_670 , w_671 , w_672 , w_673 , w_674 , w_675 , w_676 , w_677 , 
		w_678 , w_679 , w_680 , w_681 , w_682 , w_683 , w_684 , w_685 , w_686 , w_687 , 
		w_688 , w_689 , w_690 , w_691 , w_692 , w_693 , w_694 , w_695 , w_696 , w_697 , 
		w_698 , w_699 , w_700 , w_701 , w_702 , w_703 , w_704 , w_705 , w_706 , w_707 , 
		w_708 , w_709 , w_710 , w_711 , w_712 , w_713 , w_714 , w_715 , w_716 , w_717 , 
		w_718 , w_719 , w_720 , w_721 , w_722 , w_723 , w_724 , w_725 , w_726 , w_727 , 
		w_728 , w_729 , w_730 , w_731 , w_732 , w_733 , w_734 , w_735 , w_736 , w_737 , 
		w_738 , w_739 , w_740 , w_741 , w_742 , w_743 , w_744 , w_745 , w_746 , w_747 , 
		w_748 , w_749 , w_750 , w_751 , w_752 , w_753 , w_754 , w_755 , w_756 , w_757 , 
		w_758 , w_759 , w_760 , w_761 , w_762 , w_763 , w_764 , w_765 , w_766 , w_767 , 
		w_768 , w_769 , w_770 , w_771 , w_772 , w_773 , w_774 , w_775 , w_776 , w_777 , 
		w_778 , w_779 , w_780 , w_781 , w_782 , w_783 , w_784 , w_785 , w_786 , w_787 , 
		w_788 , w_789 , w_790 , w_791 , w_792 , w_793 , w_794 , w_795 , w_796 , w_797 , 
		w_798 , w_799 , w_800 , w_801 , w_802 , w_803 , w_804 , w_805 , w_806 , w_807 , 
		w_808 , w_809 , w_810 , w_811 , w_812 , w_813 , w_814 , w_815 , w_816 , w_817 , 
		w_818 , w_819 , w_820 , w_821 , w_822 , w_823 , w_824 , w_825 , w_826 , w_827 , 
		w_828 , w_829 , w_830 , w_831 , w_832 , w_833 , w_834 , w_835 , w_836 , w_837 , 
		w_838 , w_839 , w_840 , w_841 , w_842 , w_843 , w_844 , w_845 , w_846 , w_847 , 
		w_848 , w_849 , w_850 , w_851 , w_852 , w_853 , w_854 , w_855 , w_856 , w_857 , 
		w_858 , w_859 , w_860 , w_861 , w_862 , w_863 , w_864 , w_865 , w_866 , w_867 , 
		w_868 , w_869 , w_870 , w_871 , w_872 , w_873 , w_874 , w_875 , w_876 , w_877 , 
		w_878 , w_879 , w_880 , w_881 , w_882 , w_883 , w_884 , w_885 , w_886 , w_887 , 
		w_888 , w_889 , w_890 , w_891 , w_892 , w_893 , w_894 , w_895 , w_896 , w_897 , 
		w_898 , w_899 , w_900 , w_901 , w_902 , w_903 , w_904 , w_905 , w_906 , w_907 , 
		w_908 , w_909 , w_910 , w_911 , w_912 , w_913 , w_914 , w_915 , w_916 , w_917 , 
		w_918 , w_919 , w_920 , w_921 , w_922 , w_923 , w_924 , w_925 , w_926 , w_927 , 
		w_928 , w_929 , w_930 , w_931 , w_932 , w_933 , w_934 , w_935 , w_936 , w_937 , 
		w_938 , w_939 , w_940 , w_941 , w_942 , w_943 , w_944 , w_945 , w_946 , w_947 , 
		w_948 , w_949 , w_950 , w_951 , w_952 , w_953 , w_954 , w_955 , w_956 , w_957 , 
		w_958 , w_959 , w_960 , w_961 , w_962 , w_963 , w_964 , w_965 , w_966 , w_967 , 
		w_968 , w_969 , w_970 , w_971 , w_972 , w_973 , w_974 , w_975 , w_976 , w_977 , 
		w_978 , w_979 , w_980 , w_981 , w_982 , w_983 , w_984 , w_985 , w_986 , w_987 , 
		w_988 , w_989 , w_990 , w_991 , w_992 , w_993 , w_994 , w_995 , w_996 , w_997 , 
		w_998 , w_999 , w_1000 , w_1001 , w_1002 , w_1003 , w_1004 , w_1005 , w_1006 , w_1007 , 
		w_1008 , w_1009 , w_1010 , w_1011 , w_1012 , w_1013 , w_1014 , w_1015 , w_1016 , w_1017 , 
		w_1018 , w_1019 , w_1020 , w_1021 , w_1022 , w_1023 , w_1024 , w_1025 , w_1026 , w_1027 , 
		w_1028 , w_1029 , w_1030 , w_1031 , w_1032 , w_1033 , w_1034 , w_1035 , w_1036 , w_1037 , 
		w_1038 , w_1039 , w_1040 , w_1041 , w_1042 , w_1043 , w_1044 , w_1045 , w_1046 , w_1047 , 
		w_1048 , w_1049 , w_1050 , w_1051 , w_1052 , w_1053 , w_1054 , w_1055 , w_1056 , w_1057 , 
		w_1058 , w_1059 , w_1060 , w_1061 , w_1062 , w_1063 , w_1064 , w_1065 , w_1066 , w_1067 , 
		w_1068 , w_1069 , w_1070 , w_1071 , w_1072 , w_1073 , w_1074 , w_1075 , w_1076 , w_1077 , 
		w_1078 , w_1079 , w_1080 , w_1081 , w_1082 , w_1083 , w_1084 , w_1085 , w_1086 , w_1087 , 
		w_1088 , w_1089 , w_1090 , w_1091 , w_1092 , w_1093 , w_1094 , w_1095 , w_1096 , w_1097 , 
		w_1098 , w_1099 , w_1100 , w_1101 , w_1102 , w_1103 , w_1104 , w_1105 , w_1106 , w_1107 , 
		w_1108 , w_1109 , w_1110 , w_1111 , w_1112 , w_1113 , w_1114 , w_1115 , w_1116 , w_1117 , 
		w_1118 , w_1119 , w_1120 , w_1121 , w_1122 , w_1123 , w_1124 , w_1125 , w_1126 , w_1127 , 
		w_1128 , w_1129 , w_1130 , w_1131 , w_1132 , w_1133 , w_1134 , w_1135 , w_1136 , w_1137 , 
		w_1138 , w_1139 , w_1140 , w_1141 , w_1142 , w_1143 , w_1144 , w_1145 , w_1146 , w_1147 , 
		w_1148 , w_1149 , w_1150 , w_1151 , w_1152 , w_1153 , w_1154 , w_1155 , w_1156 , w_1157 , 
		w_1158 , w_1159 , w_1160 , w_1161 , w_1162 , w_1163 , w_1164 , w_1165 , w_1166 , w_1167 , 
		w_1168 , w_1169 , w_1170 , w_1171 , w_1172 , w_1173 , w_1174 , w_1175 , w_1176 , w_1177 , 
		w_1178 , w_1179 , w_1180 , w_1181 , w_1182 , w_1183 , w_1184 , w_1185 , w_1186 , w_1187 , 
		w_1188 , w_1189 , w_1190 , w_1191 , w_1192 , w_1193 , w_1194 , w_1195 , w_1196 , w_1197 , 
		w_1198 , w_1199 , w_1200 , w_1201 , w_1202 , w_1203 , w_1204 , w_1205 , w_1206 , w_1207 , 
		w_1208 , w_1209 , w_1210 , w_1211 , w_1212 , w_1213 , w_1214 , w_1215 , w_1216 , w_1217 , 
		w_1218 , w_1219 , w_1220 , w_1221 , w_1222 , w_1223 , w_1224 , w_1225 , w_1226 , w_1227 , 
		w_1228 , w_1229 , w_1230 , w_1231 , w_1232 , w_1233 , w_1234 , w_1235 , w_1236 , w_1237 , 
		w_1238 , w_1239 , w_1240 , w_1241 , w_1242 , w_1243 , w_1244 , w_1245 , w_1246 , w_1247 , 
		w_1248 , w_1249 , w_1250 , w_1251 , w_1252 , w_1253 , w_1254 , w_1255 , w_1256 , w_1257 , 
		w_1258 , w_1259 , w_1260 , w_1261 , w_1262 , w_1263 , w_1264 , w_1265 , w_1266 , w_1267 , 
		w_1268 , w_1269 , w_1270 , w_1271 , w_1272 , w_1273 , w_1274 , w_1275 , w_1276 , w_1277 , 
		w_1278 , w_1279 , w_1280 , w_1281 , w_1282 , w_1283 , w_1284 , w_1285 , w_1286 , w_1287 , 
		w_1288 , w_1289 , w_1290 , w_1291 , w_1292 , w_1293 , w_1294 , w_1295 , w_1296 , w_1297 , 
		w_1298 , w_1299 , w_1300 , w_1301 , w_1302 , w_1303 , w_1304 , w_1305 , w_1306 , w_1307 , 
		w_1308 , w_1309 , w_1310 , w_1311 , w_1312 , w_1313 , w_1314 , w_1315 , w_1316 , w_1317 , 
		w_1318 , w_1319 , w_1320 , w_1321 , w_1322 , w_1323 , w_1324 , w_1325 , w_1326 , w_1327 , 
		w_1328 , w_1329 , w_1330 , w_1331 , w_1332 , w_1333 , w_1334 , w_1335 , w_1336 , w_1337 , 
		w_1338 , w_1339 , w_1340 , w_1341 , w_1342 , w_1343 , w_1344 , w_1345 , w_1346 , w_1347 , 
		w_1348 , w_1349 , w_1350 , w_1351 , w_1352 , w_1353 , w_1354 , w_1355 , w_1356 , w_1357 , 
		w_1358 , w_1359 , w_1360 , w_1361 , w_1362 , w_1363 , w_1364 , w_1365 , w_1366 , w_1367 , 
		w_1368 , w_1369 , w_1370 , w_1371 , w_1372 , w_1373 , w_1374 , w_1375 , w_1376 , w_1377 , 
		w_1378 , w_1379 , w_1380 , w_1381 , w_1382 , w_1383 , w_1384 , w_1385 , w_1386 , w_1387 , 
		w_1388 , w_1389 , w_1390 , w_1391 , w_1392 , w_1393 , w_1394 , w_1395 , w_1396 , w_1397 , 
		w_1398 , w_1399 , w_1400 , w_1401 , w_1402 , w_1403 , w_1404 , w_1405 , w_1406 , w_1407 , 
		w_1408 , w_1409 , w_1410 , w_1411 , w_1412 , w_1413 , w_1414 , w_1415 , w_1416 , w_1417 , 
		w_1418 , w_1419 , w_1420 , w_1421 , w_1422 , w_1423 , w_1424 , w_1425 , w_1426 , w_1427 , 
		w_1428 , w_1429 , w_1430 , w_1431 , w_1432 , w_1433 , w_1434 , w_1435 , w_1436 , w_1437 , 
		w_1438 , w_1439 , w_1440 , w_1441 , w_1442 , w_1443 , w_1444 , w_1445 , w_1446 , w_1447 , 
		w_1448 , w_1449 , w_1450 , w_1451 , w_1452 , w_1453 , w_1454 , w_1455 , w_1456 , w_1457 , 
		w_1458 , w_1459 , w_1460 , w_1461 , w_1462 , w_1463 , w_1464 , w_1465 , w_1466 , w_1467 , 
		w_1468 , w_1469 , w_1470 , w_1471 , w_1472 , w_1473 , w_1474 , w_1475 , w_1476 , w_1477 , 
		w_1478 , w_1479 , w_1480 , w_1481 , w_1482 , w_1483 , w_1484 , w_1485 , w_1486 , w_1487 , 
		w_1488 , w_1489 , w_1490 , w_1491 , w_1492 , w_1493 , w_1494 , w_1495 , w_1496 , w_1497 , 
		w_1498 , w_1499 , w_1500 , w_1501 , w_1502 , w_1503 , w_1504 , w_1505 , w_1506 , w_1507 , 
		w_1508 , w_1509 , w_1510 , w_1511 , w_1512 , w_1513 , w_1514 , w_1515 , w_1516 , w_1517 , 
		w_1518 , w_1519 , w_1520 , w_1521 , w_1522 , w_1523 , w_1524 , w_1525 , w_1526 , w_1527 , 
		w_1528 , w_1529 , w_1530 , w_1531 , w_1532 , w_1533 , w_1534 , w_1535 , w_1536 , w_1537 , 
		w_1538 , w_1539 , w_1540 , w_1541 , w_1542 , w_1543 , w_1544 , w_1545 , w_1546 , w_1547 , 
		w_1548 , w_1549 , w_1550 , w_1551 , w_1552 , w_1553 , w_1554 , w_1555 , w_1556 , w_1557 , 
		w_1558 , w_1559 , w_1560 , w_1561 , w_1562 , w_1563 , w_1564 , w_1565 , w_1566 , w_1567 , 
		w_1568 , w_1569 , w_1570 , w_1571 , w_1572 , w_1573 , w_1574 , w_1575 , w_1576 , w_1577 , 
		w_1578 , w_1579 , w_1580 , w_1581 , w_1582 , w_1583 , w_1584 , w_1585 , w_1586 , w_1587 , 
		w_1588 , w_1589 , w_1590 , w_1591 , w_1592 , w_1593 , w_1594 , w_1595 , w_1596 , w_1597 , 
		w_1598 , w_1599 , w_1600 , w_1601 , w_1602 , w_1603 , w_1604 , w_1605 , w_1606 , w_1607 , 
		w_1608 , w_1609 , w_1610 , w_1611 , w_1612 , w_1613 , w_1614 , w_1615 , w_1616 , w_1617 , 
		w_1618 , w_1619 , w_1620 , w_1621 , w_1622 , w_1623 , w_1624 , w_1625 , w_1626 , w_1627 , 
		w_1628 , w_1629 , w_1630 , w_1631 , w_1632 , w_1633 , w_1634 , w_1635 , w_1636 , w_1637 , 
		w_1638 , w_1639 , w_1640 , w_1641 , w_1642 , w_1643 , w_1644 , w_1645 , w_1646 , w_1647 , 
		w_1648 , w_1649 , w_1650 , w_1651 , w_1652 , w_1653 , w_1654 , w_1655 , w_1656 , w_1657 , 
		w_1658 , w_1659 , w_1660 , w_1661 , w_1662 , w_1663 , w_1664 , w_1665 , w_1666 , w_1667 , 
		w_1668 , w_1669 , w_1670 , w_1671 , w_1672 , w_1673 , w_1674 , w_1675 , w_1676 , w_1677 , 
		w_1678 , w_1679 , w_1680 , w_1681 , w_1682 , w_1683 , w_1684 , w_1685 , w_1686 , w_1687 , 
		w_1688 , w_1689 , w_1690 , w_1691 , w_1692 , w_1693 , w_1694 , w_1695 , w_1696 , w_1697 , 
		w_1698 , w_1699 , w_1700 , w_1701 , w_1702 , w_1703 , w_1704 , w_1705 , w_1706 , w_1707 , 
		w_1708 , w_1709 , w_1710 , w_1711 , w_1712 , w_1713 , w_1714 , w_1715 , w_1716 , w_1717 , 
		w_1718 , w_1719 , w_1720 , w_1721 , w_1722 , w_1723 , w_1724 , w_1725 , w_1726 , w_1727 , 
		w_1728 , w_1729 , w_1730 , w_1731 , w_1732 , w_1733 , w_1734 , w_1735 , w_1736 , w_1737 , 
		w_1738 , w_1739 , w_1740 , w_1741 , w_1742 , w_1743 , w_1744 , w_1745 , w_1746 , w_1747 , 
		w_1748 , w_1749 , w_1750 , w_1751 , w_1752 , w_1753 , w_1754 , w_1755 , w_1756 , w_1757 , 
		w_1758 , w_1759 , w_1760 , w_1761 , w_1762 , w_1763 , w_1764 , w_1765 , w_1766 , w_1767 , 
		w_1768 , w_1769 , w_1770 , w_1771 , w_1772 , w_1773 , w_1774 , w_1775 , w_1776 , w_1777 , 
		w_1778 , w_1779 , w_1780 , w_1781 , w_1782 , w_1783 , w_1784 , w_1785 , w_1786 , w_1787 , 
		w_1788 , w_1789 , w_1790 , w_1791 , w_1792 , w_1793 , w_1794 , w_1795 , w_1796 , w_1797 , 
		w_1798 , w_1799 , w_1800 , w_1801 , w_1802 , w_1803 , w_1804 , w_1805 , w_1806 , w_1807 , 
		w_1808 , w_1809 , w_1810 , w_1811 , w_1812 , w_1813 , w_1814 , w_1815 , w_1816 , w_1817 , 
		w_1818 , w_1819 , w_1820 , w_1821 , w_1822 , w_1823 , w_1824 , w_1825 , w_1826 , w_1827 , 
		w_1828 , w_1829 , w_1830 , w_1831 , w_1832 , w_1833 , w_1834 , w_1835 , w_1836 , w_1837 , 
		w_1838 , w_1839 , w_1840 , w_1841 , w_1842 , w_1843 , w_1844 , w_1845 , w_1846 , w_1847 , 
		w_1848 , w_1849 , w_1850 , w_1851 , w_1852 , w_1853 , w_1854 , w_1855 , w_1856 , w_1857 , 
		w_1858 , w_1859 , w_1860 , w_1861 , w_1862 , w_1863 , w_1864 , w_1865 , w_1866 , w_1867 , 
		w_1868 , w_1869 , w_1870 , w_1871 , w_1872 , w_1873 , w_1874 , w_1875 , w_1876 , w_1877 , 
		w_1878 , w_1879 , w_1880 , w_1881 , w_1882 , w_1883 , w_1884 , w_1885 , w_1886 , w_1887 , 
		w_1888 , w_1889 , w_1890 , w_1891 , w_1892 , w_1893 , w_1894 , w_1895 , w_1896 , w_1897 , 
		w_1898 , w_1899 , w_1900 , w_1901 , w_1902 , w_1903 , w_1904 , w_1905 , w_1906 , w_1907 , 
		w_1908 , w_1909 , w_1910 , w_1911 , w_1912 , w_1913 , w_1914 , w_1915 , w_1916 , w_1917 , 
		w_1918 , w_1919 , w_1920 , w_1921 , w_1922 , w_1923 , w_1924 , w_1925 , w_1926 , w_1927 , 
		w_1928 , w_1929 , w_1930 , w_1931 , w_1932 , w_1933 , w_1934 , w_1935 , w_1936 , w_1937 , 
		w_1938 , w_1939 , w_1940 , w_1941 , w_1942 , w_1943 , w_1944 , w_1945 , w_1946 , w_1947 , 
		w_1948 , w_1949 , w_1950 , w_1951 , w_1952 , w_1953 , w_1954 , w_1955 , w_1956 , w_1957 , 
		w_1958 , w_1959 , w_1960 , w_1961 , w_1962 , w_1963 , w_1964 , w_1965 , w_1966 , w_1967 , 
		w_1968 , w_1969 , w_1970 , w_1971 , w_1972 , w_1973 , w_1974 , w_1975 , w_1976 , w_1977 , 
		w_1978 , w_1979 , w_1980 , w_1981 , w_1982 , w_1983 , w_1984 , w_1985 , w_1986 , w_1987 , 
		w_1988 , w_1989 , w_1990 , w_1991 , w_1992 , w_1993 , w_1994 , w_1995 , w_1996 , w_1997 , 
		w_1998 , w_1999 , w_2000 , w_2001 , w_2002 , w_2003 , w_2004 , w_2005 , w_2006 , w_2007 , 
		w_2008 , w_2009 , w_2010 , w_2011 , w_2012 , w_2013 , w_2014 , w_2015 , w_2016 , w_2017 , 
		w_2018 , w_2019 , w_2020 , w_2021 , w_2022 , w_2023 , w_2024 , w_2025 , w_2026 , w_2027 , 
		w_2028 , w_2029 , w_2030 , w_2031 , w_2032 , w_2033 , w_2034 , w_2035 , w_2036 , w_2037 , 
		w_2038 , w_2039 , w_2040 , w_2041 , w_2042 , w_2043 , w_2044 , w_2045 , w_2046 , w_2047 , 
		w_2048 , w_2049 , w_2050 , w_2051 , w_2052 , w_2053 , w_2054 , w_2055 , w_2056 , w_2057 , 
		w_2058 , w_2059 , w_2060 , w_2061 , w_2062 , w_2063 , w_2064 , w_2065 , w_2066 , w_2067 , 
		w_2068 , w_2069 , w_2070 , w_2071 , w_2072 , w_2073 , w_2074 , w_2075 , w_2076 , w_2077 , 
		w_2078 , w_2079 , w_2080 , w_2081 , w_2082 , w_2083 , w_2084 , w_2085 , w_2086 , w_2087 , 
		w_2088 , w_2089 , w_2090 , w_2091 , w_2092 , w_2093 , w_2094 , w_2095 , w_2096 , w_2097 , 
		w_2098 , w_2099 , w_2100 , w_2101 , w_2102 , w_2103 , w_2104 , w_2105 , w_2106 , w_2107 , 
		w_2108 , w_2109 , w_2110 , w_2111 , w_2112 , w_2113 , w_2114 , w_2115 , w_2116 , w_2117 , 
		w_2118 , w_2119 , w_2120 , w_2121 , w_2122 , w_2123 , w_2124 , w_2125 , w_2126 , w_2127 , 
		w_2128 , w_2129 , w_2130 , w_2131 , w_2132 , w_2133 , w_2134 , w_2135 , w_2136 , w_2137 , 
		w_2138 , w_2139 , w_2140 , w_2141 , w_2142 , w_2143 , w_2144 , w_2145 , w_2146 , w_2147 , 
		w_2148 , w_2149 , w_2150 , w_2151 , w_2152 , w_2153 , w_2154 , w_2155 , w_2156 , w_2157 , 
		w_2158 , w_2159 , w_2160 , w_2161 , w_2162 , w_2163 , w_2164 , w_2165 , w_2166 , w_2167 , 
		w_2168 , w_2169 , w_2170 , w_2171 , w_2172 , w_2173 , w_2174 , w_2175 , w_2176 , w_2177 , 
		w_2178 , w_2179 , w_2180 , w_2181 , w_2182 , w_2183 , w_2184 , w_2185 , w_2186 , w_2187 , 
		w_2188 , w_2189 , w_2190 , w_2191 , w_2192 , w_2193 , w_2194 , w_2195 , w_2196 , w_2197 , 
		w_2198 , w_2199 , w_2200 , w_2201 , w_2202 , w_2203 , w_2204 , w_2205 , w_2206 , w_2207 , 
		w_2208 , w_2209 , w_2210 , w_2211 , w_2212 , w_2213 , w_2214 , w_2215 , w_2216 , w_2217 , 
		w_2218 , w_2219 , w_2220 , w_2221 , w_2222 , w_2223 , w_2224 , w_2225 , w_2226 , w_2227 , 
		w_2228 , w_2229 , w_2230 , w_2231 , w_2232 , w_2233 , w_2234 , w_2235 , w_2236 , w_2237 , 
		w_2238 , w_2239 , w_2240 , w_2241 , w_2242 , w_2243 , w_2244 , w_2245 , w_2246 , w_2247 , 
		w_2248 , w_2249 , w_2250 , w_2251 , w_2252 , w_2253 , w_2254 , w_2255 , w_2256 , w_2257 , 
		w_2258 , w_2259 , w_2260 , w_2261 , w_2262 , w_2263 , w_2264 , w_2265 , w_2266 , w_2267 , 
		w_2268 , w_2269 , w_2270 , w_2271 , w_2272 , w_2273 , w_2274 , w_2275 , w_2276 , w_2277 , 
		w_2278 , w_2279 , w_2280 , w_2281 , w_2282 , w_2283 , w_2284 , w_2285 , w_2286 , w_2287 , 
		w_2288 , w_2289 , w_2290 , w_2291 , w_2292 , w_2293 , w_2294 , w_2295 , w_2296 , w_2297 , 
		w_2298 , w_2299 , w_2300 , w_2301 , w_2302 , w_2303 , w_2304 , w_2305 , w_2306 , w_2307 , 
		w_2308 , w_2309 , w_2310 , w_2311 , w_2312 , w_2313 , w_2314 , w_2315 , w_2316 , w_2317 , 
		w_2318 , w_2319 , w_2320 , w_2321 , w_2322 , w_2323 , w_2324 , w_2325 , w_2326 , w_2327 , 
		w_2328 , w_2329 , w_2330 , w_2331 , w_2332 , w_2333 , w_2334 , w_2335 , w_2336 , w_2337 , 
		w_2338 , w_2339 , w_2340 , w_2341 , w_2342 , w_2343 , w_2344 , w_2345 , w_2346 , w_2347 , 
		w_2348 , w_2349 , w_2350 , w_2351 , w_2352 , w_2353 , w_2354 , w_2355 , w_2356 , w_2357 , 
		w_2358 , w_2359 , w_2360 , w_2361 , w_2362 , w_2363 , w_2364 , w_2365 , w_2366 , w_2367 , 
		w_2368 , w_2369 , w_2370 , w_2371 , w_2372 , w_2373 , w_2374 , w_2375 , w_2376 , w_2377 , 
		w_2378 , w_2379 , w_2380 , w_2381 , w_2382 , w_2383 , w_2384 , w_2385 , w_2386 , w_2387 , 
		w_2388 , w_2389 , w_2390 , w_2391 , w_2392 , w_2393 , w_2394 , w_2395 , w_2396 , w_2397 , 
		w_2398 , w_2399 , w_2400 , w_2401 , w_2402 , w_2403 , w_2404 , w_2405 , w_2406 , w_2407 , 
		w_2408 , w_2409 , w_2410 , w_2411 , w_2412 , w_2413 , w_2414 , w_2415 , w_2416 , w_2417 , 
		w_2418 , w_2419 , w_2420 , w_2421 , w_2422 , w_2423 , w_2424 , w_2425 , w_2426 , w_2427 , 
		w_2428 , w_2429 , w_2430 , w_2431 , w_2432 , w_2433 , w_2434 , w_2435 , w_2436 , w_2437 , 
		w_2438 , w_2439 , w_2440 , w_2441 , w_2442 , w_2443 , w_2444 , w_2445 , w_2446 , w_2447 , 
		w_2448 , w_2449 , w_2450 , w_2451 , w_2452 , w_2453 , w_2454 , w_2455 , w_2456 , w_2457 , 
		w_2458 , w_2459 , w_2460 , w_2461 , w_2462 , w_2463 , w_2464 , w_2465 , w_2466 , w_2467 , 
		w_2468 , w_2469 , w_2470 , w_2471 , w_2472 , w_2473 , w_2474 , w_2475 , w_2476 , w_2477 , 
		w_2478 , w_2479 , w_2480 , w_2481 , w_2482 , w_2483 , w_2484 , w_2485 , w_2486 , w_2487 , 
		w_2488 , w_2489 , w_2490 , w_2491 , w_2492 , w_2493 , w_2494 , w_2495 , w_2496 , w_2497 , 
		w_2498 , w_2499 , w_2500 , w_2501 , w_2502 , w_2503 , w_2504 , w_2505 , w_2506 , w_2507 , 
		w_2508 , w_2509 , w_2510 , w_2511 , w_2512 , w_2513 , w_2514 , w_2515 , w_2516 , w_2517 , 
		w_2518 , w_2519 , w_2520 , w_2521 , w_2522 , w_2523 , w_2524 , w_2525 , w_2526 , w_2527 , 
		w_2528 , w_2529 , w_2530 , w_2531 , w_2532 , w_2533 , w_2534 , w_2535 , w_2536 , w_2537 , 
		w_2538 , w_2539 , w_2540 , w_2541 , w_2542 , w_2543 , w_2544 , w_2545 , w_2546 , w_2547 , 
		w_2548 , w_2549 , w_2550 , w_2551 , w_2552 , w_2553 , w_2554 , w_2555 , w_2556 , w_2557 , 
		w_2558 , w_2559 , w_2560 , w_2561 , w_2562 , w_2563 , w_2564 , w_2565 , w_2566 , w_2567 , 
		w_2568 , w_2569 , w_2570 , w_2571 , w_2572 , w_2573 , w_2574 , w_2575 , w_2576 , w_2577 , 
		w_2578 , w_2579 , w_2580 , w_2581 , w_2582 , w_2583 , w_2584 , w_2585 , w_2586 , w_2587 , 
		w_2588 , w_2589 , w_2590 , w_2591 , w_2592 , w_2593 , w_2594 , w_2595 , w_2596 , w_2597 , 
		w_2598 , w_2599 , w_2600 , w_2601 , w_2602 , w_2603 , w_2604 , w_2605 , w_2606 , w_2607 , 
		w_2608 , w_2609 , w_2610 , w_2611 , w_2612 , w_2613 , w_2614 , w_2615 , w_2616 , w_2617 , 
		w_2618 , w_2619 , w_2620 , w_2621 , w_2622 , w_2623 , w_2624 , w_2625 , w_2626 , w_2627 , 
		w_2628 , w_2629 , w_2630 , w_2631 , w_2632 , w_2633 , w_2634 , w_2635 , w_2636 , w_2637 , 
		w_2638 , w_2639 , w_2640 , w_2641 , w_2642 , w_2643 , w_2644 , w_2645 , w_2646 , w_2647 , 
		w_2648 , w_2649 , w_2650 , w_2651 , w_2652 , w_2653 , w_2654 , w_2655 , w_2656 , w_2657 , 
		w_2658 , w_2659 , w_2660 , w_2661 , w_2662 , w_2663 , w_2664 , w_2665 , w_2666 , w_2667 , 
		w_2668 , w_2669 , w_2670 , w_2671 , w_2672 , w_2673 , w_2674 , w_2675 , w_2676 , w_2677 , 
		w_2678 , w_2679 , w_2680 , w_2681 , w_2682 , w_2683 , w_2684 , w_2685 , w_2686 , w_2687 , 
		w_2688 , w_2689 , w_2690 , w_2691 , w_2692 , w_2693 , w_2694 , w_2695 , w_2696 , w_2697 , 
		w_2698 , w_2699 , w_2700 , w_2701 , w_2702 , w_2703 , w_2704 , w_2705 , w_2706 , w_2707 , 
		w_2708 , w_2709 , w_2710 , w_2711 , w_2712 , w_2713 , w_2714 , w_2715 , w_2716 , w_2717 , 
		w_2718 , w_2719 , w_2720 , w_2721 , w_2722 , w_2723 , w_2724 , w_2725 , w_2726 , w_2727 , 
		w_2728 , w_2729 , w_2730 , w_2731 , w_2732 , w_2733 , w_2734 , w_2735 , w_2736 , w_2737 , 
		w_2738 , w_2739 , w_2740 , w_2741 , w_2742 , w_2743 , w_2744 , w_2745 , w_2746 , w_2747 , 
		w_2748 , w_2749 , w_2750 , w_2751 , w_2752 , w_2753 , w_2754 , w_2755 , w_2756 , w_2757 , 
		w_2758 , w_2759 , w_2760 , w_2761 , w_2762 , w_2763 , w_2764 , w_2765 , w_2766 , w_2767 , 
		w_2768 , w_2769 , w_2770 , w_2771 , w_2772 , w_2773 , w_2774 , w_2775 , w_2776 , w_2777 , 
		w_2778 , w_2779 , w_2780 , w_2781 , w_2782 , w_2783 , w_2784 , w_2785 , w_2786 , w_2787 , 
		w_2788 , w_2789 , w_2790 , w_2791 , w_2792 , w_2793 , w_2794 , w_2795 , w_2796 , w_2797 , 
		w_2798 , w_2799 , w_2800 , w_2801 , w_2802 , w_2803 , w_2804 , w_2805 , w_2806 , w_2807 , 
		w_2808 , w_2809 , w_2810 , w_2811 , w_2812 , w_2813 , w_2814 , w_2815 , w_2816 , w_2817 , 
		w_2818 , w_2819 , w_2820 , w_2821 , w_2822 , w_2823 , w_2824 , w_2825 , w_2826 , w_2827 , 
		w_2828 , w_2829 , w_2830 , w_2831 , w_2832 , w_2833 , w_2834 , w_2835 , w_2836 , w_2837 , 
		w_2838 , w_2839 , w_2840 , w_2841 , w_2842 , w_2843 , w_2844 , w_2845 , w_2846 , w_2847 , 
		w_2848 , w_2849 , w_2850 , w_2851 , w_2852 , w_2853 , w_2854 , w_2855 , w_2856 , w_2857 , 
		w_2858 , w_2859 , w_2860 , w_2861 , w_2862 , w_2863 , w_2864 , w_2865 , w_2866 , w_2867 , 
		w_2868 , w_2869 , w_2870 , w_2871 , w_2872 , w_2873 , w_2874 , w_2875 , w_2876 , w_2877 , 
		w_2878 , w_2879 , w_2880 , w_2881 , w_2882 , w_2883 , w_2884 , w_2885 , w_2886 , w_2887 , 
		w_2888 , w_2889 , w_2890 , w_2891 , w_2892 , w_2893 , w_2894 , w_2895 , w_2896 , w_2897 , 
		w_2898 , w_2899 , w_2900 , w_2901 , w_2902 , w_2903 , w_2904 , w_2905 , w_2906 , w_2907 , 
		w_2908 , w_2909 , w_2910 , w_2911 , w_2912 , w_2913 , w_2914 , w_2915 , w_2916 , w_2917 , 
		w_2918 , w_2919 , w_2920 , w_2921 , w_2922 , w_2923 , w_2924 , w_2925 , w_2926 , w_2927 , 
		w_2928 , w_2929 , w_2930 , w_2931 , w_2932 , w_2933 , w_2934 , w_2935 , w_2936 , w_2937 , 
		w_2938 , w_2939 , w_2940 , w_2941 , w_2942 , w_2943 , w_2944 , w_2945 , w_2946 , w_2947 , 
		w_2948 , w_2949 , w_2950 , w_2951 , w_2952 , w_2953 , w_2954 , w_2955 , w_2956 , w_2957 , 
		w_2958 , w_2959 , w_2960 , w_2961 , w_2962 , w_2963 , w_2964 , w_2965 , w_2966 , w_2967 , 
		w_2968 , w_2969 , w_2970 , w_2971 , w_2972 , w_2973 , w_2974 , w_2975 , w_2976 , w_2977 , 
		w_2978 , w_2979 , w_2980 , w_2981 , w_2982 , w_2983 , w_2984 , w_2985 , w_2986 , w_2987 , 
		w_2988 , w_2989 , w_2990 , w_2991 , w_2992 , w_2993 , w_2994 , w_2995 , w_2996 , w_2997 , 
		w_2998 , w_2999 , w_3000 , w_3001 , w_3002 , w_3003 , w_3004 , w_3005 , w_3006 , w_3007 , 
		w_3008 , w_3009 , w_3010 , w_3011 , w_3012 , w_3013 , w_3014 , w_3015 , w_3016 , w_3017 , 
		w_3018 , w_3019 , w_3020 , w_3021 , w_3022 , w_3023 , w_3024 , w_3025 , w_3026 , w_3027 , 
		w_3028 , w_3029 , w_3030 , w_3031 , w_3032 , w_3033 , w_3034 , w_3035 , w_3036 , w_3037 , 
		w_3038 , w_3039 , w_3040 , w_3041 , w_3042 , w_3043 , w_3044 , w_3045 , w_3046 , w_3047 , 
		w_3048 , w_3049 , w_3050 , w_3051 , w_3052 , w_3053 , w_3054 , w_3055 , w_3056 , w_3057 , 
		w_3058 , w_3059 , w_3060 , w_3061 , w_3062 , w_3063 , w_3064 , w_3065 , w_3066 , w_3067 , 
		w_3068 , w_3069 , w_3070 , w_3071 , w_3072 , w_3073 , w_3074 , w_3075 , w_3076 , w_3077 , 
		w_3078 , w_3079 , w_3080 , w_3081 , w_3082 , w_3083 , w_3084 , w_3085 , w_3086 , w_3087 , 
		w_3088 , w_3089 , w_3090 , w_3091 , w_3092 , w_3093 , w_3094 , w_3095 , w_3096 , w_3097 , 
		w_3098 , w_3099 , w_3100 , w_3101 , w_3102 , w_3103 , w_3104 , w_3105 , w_3106 , w_3107 , 
		w_3108 , w_3109 , w_3110 , w_3111 , w_3112 , w_3113 , w_3114 , w_3115 , w_3116 , w_3117 , 
		w_3118 , w_3119 , w_3120 , w_3121 , w_3122 , w_3123 , w_3124 , w_3125 , w_3126 , w_3127 , 
		w_3128 , w_3129 , w_3130 , w_3131 , w_3132 , w_3133 , w_3134 , w_3135 , w_3136 , w_3137 , 
		w_3138 , w_3139 , w_3140 , w_3141 , w_3142 , w_3143 , w_3144 , w_3145 , w_3146 , w_3147 , 
		w_3148 , w_3149 , w_3150 , w_3151 , w_3152 , w_3153 , w_3154 , w_3155 , w_3156 , w_3157 , 
		w_3158 , w_3159 , w_3160 , w_3161 , w_3162 , w_3163 , w_3164 , w_3165 , w_3166 , w_3167 , 
		w_3168 , w_3169 , w_3170 , w_3171 , w_3172 , w_3173 , w_3174 , w_3175 , w_3176 , w_3177 , 
		w_3178 , w_3179 , w_3180 , w_3181 , w_3182 , w_3183 , w_3184 , w_3185 , w_3186 , w_3187 , 
		w_3188 , w_3189 , w_3190 , w_3191 , w_3192 , w_3193 , w_3194 , w_3195 , w_3196 , w_3197 , 
		w_3198 , w_3199 , w_3200 , w_3201 , w_3202 , w_3203 , w_3204 , w_3205 , w_3206 , w_3207 ;
buf ( \O[19]_b1 , \934_b1 );
buf ( \O[19]_b0 , \934_b0 );
buf ( \O[18]_b1 , \940_b1 );
buf ( \O[18]_b0 , \940_b0 );
buf ( \O[17]_b1 , \960_b1 );
buf ( \O[17]_b0 , \960_b0 );
buf ( \O[16]_b1 , \1067_b1 );
buf ( \O[16]_b0 , \1067_b0 );
buf ( \O[15]_b1 , \979_b1 );
buf ( \O[15]_b0 , \979_b0 );
buf ( \O[14]_b1 , \1068_b1 );
buf ( \O[14]_b0 , \1068_b0 );
buf ( \O[13]_b1 , \991_b1 );
buf ( \O[13]_b0 , \991_b0 );
buf ( \O[12]_b1 , \1069_b1 );
buf ( \O[12]_b0 , \1069_b0 );
buf ( \O[11]_b1 , \1004_b1 );
buf ( \O[11]_b0 , \1004_b0 );
buf ( \O[10]_b1 , \1011_b1 );
buf ( \O[10]_b0 , \1011_b0 );
buf ( \O[9]_b1 , \1018_b1 );
buf ( \O[9]_b0 , \1018_b0 );
buf ( \O[8]_b1 , \1024_b1 );
buf ( \O[8]_b0 , \1024_b0 );
buf ( \O[7]_b1 , \1033_b1 );
buf ( \O[7]_b0 , \1033_b0 );
buf ( \O[6]_b1 , \1041_b1 );
buf ( \O[6]_b0 , \1041_b0 );
buf ( \O[5]_b1 , \1047_b1 );
buf ( \O[5]_b0 , \1047_b0 );
buf ( \O[4]_b1 , \1053_b1 );
buf ( \O[4]_b0 , \1053_b0 );
buf ( \O[3]_b1 , \1059_b1 );
buf ( \O[3]_b0 , \1059_b0 );
buf ( \O[2]_b1 , \1061_b1 );
buf ( \O[2]_b0 , \1061_b0 );
buf ( \O[1]_b1 , \1065_b1 );
buf ( \O[1]_b0 , \1065_b0 );
buf ( \O[0]_b1 , \1066_b1 );
buf ( \O[0]_b0 , \1066_b0 );
or ( \71_b1 , \I[1]_b1 , w_1 );
not ( w_1 , w_2 );
and ( \71_b0 , \I[1]_b0 , w_3 );
and ( w_2 ,  , w_3 );
buf ( w_1 , \I[0]_b1 );
not ( w_1 , w_4 );
not (  , w_5 );
and ( w_4 , w_5 , \I[0]_b0 );
buf ( \72_b1 , \71_b1 );
not ( \72_b1 , w_6 );
not ( \72_b0 , w_7 );
and ( w_6 , w_7 , \71_b0 );
buf ( \73_b1 , \A[0][9]_b1 );
not ( \73_b1 , w_8 );
not ( \73_b0 , w_9 );
and ( w_8 , w_9 , \A[0][9]_b0 );
or ( \74_b1 , \72_b1 , w_10 );
or ( \74_b0 , \72_b0 , \73_b0 );
not ( \73_b0 , w_11 );
and ( w_11 , w_10 , \73_b1 );
or ( \75_b1 , \A[1][9]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_12 );
and ( \75_b0 , \A[1][9]_b0 , w_13 );
and ( w_12 , w_13 , \I[0]_b0 );
or ( \76_b1 , \A[2][9]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_14 );
and ( \76_b0 , \A[2][9]_b0 , w_15 );
and ( w_14 , w_15 , \I[1]_b0 );
or ( \77_b1 , \75_b1 , w_17 );
not ( w_17 , w_18 );
and ( \77_b0 , \75_b0 , w_19 );
and ( w_18 ,  , w_19 );
buf ( w_17 , \76_b1 );
not ( w_17 , w_20 );
not (  , w_21 );
and ( w_20 , w_21 , \76_b0 );
or ( \78_b1 , \74_b1 , w_23 );
not ( w_23 , w_24 );
and ( \78_b0 , \74_b0 , w_25 );
and ( w_24 ,  , w_25 );
buf ( w_23 , \77_b1 );
not ( w_23 , w_26 );
not (  , w_27 );
and ( w_26 , w_27 , \77_b0 );
buf ( \79_b1 , \78_b1 );
buf ( \79_b0 , \78_b0 );
buf ( \80_b1 , \A[0][7]_b1 );
not ( \80_b1 , w_28 );
not ( \80_b0 , w_29 );
and ( w_28 , w_29 , \A[0][7]_b0 );
or ( \82_b1 , \A[2][7]_b1 , w_31 );
not ( w_31 , w_32 );
and ( \82_b0 , \A[2][7]_b0 , w_33 );
and ( w_32 ,  , w_33 );
buf ( w_31 , \I[1]_b1 );
not ( w_31 , w_34 );
not (  , w_35 );
and ( w_34 , w_35 , \I[1]_b0 );
or ( \83_b1 , \A[1][7]_b1 , w_37 );
not ( w_37 , w_38 );
and ( \83_b0 , \A[1][7]_b0 , w_39 );
and ( w_38 ,  , w_39 );
buf ( w_37 , \I[0]_b1 );
not ( w_37 , w_40 );
not (  , w_41 );
and ( w_40 , w_41 , \I[0]_b0 );
or ( \84_b1 , \82_b1 , w_43 );
not ( w_43 , w_44 );
and ( \84_b0 , \82_b0 , w_45 );
and ( w_44 ,  , w_45 );
buf ( w_43 , \83_b1 );
not ( w_43 , w_46 );
not (  , w_47 );
and ( w_46 , w_47 , \83_b0 );
or ( \85_b1 , \81_b1 , w_49 );
not ( w_49 , w_50 );
and ( \85_b0 , \81_b0 , w_51 );
and ( w_50 ,  , w_51 );
buf ( w_49 , \84_b1 );
not ( w_49 , w_52 );
not (  , w_53 );
and ( w_52 , w_53 , \84_b0 );
buf ( \86_b1 , \85_b1 );
not ( \86_b1 , w_54 );
not ( \86_b0 , w_55 );
and ( w_54 , w_55 , \85_b0 );
buf ( \87_b1 , \A[0][5]_b1 );
not ( \87_b1 , w_56 );
not ( \87_b0 , w_57 );
and ( w_56 , w_57 , \A[0][5]_b0 );
or ( \88_b1 , \I[1]_b1 , w_59 );
not ( w_59 , w_60 );
and ( \88_b0 , \I[1]_b0 , w_61 );
and ( w_60 ,  , w_61 );
buf ( w_59 , \I[0]_b1 );
not ( w_59 , w_62 );
not (  , w_63 );
and ( w_62 , w_63 , \I[0]_b0 );
buf ( \89_b1 , \88_b1 );
not ( \89_b1 , w_64 );
not ( \89_b0 , w_65 );
and ( w_64 , w_65 , \88_b0 );
or ( \90_b1 , \87_b1 , w_66 );
or ( \90_b0 , \87_b0 , \89_b0 );
not ( \89_b0 , w_67 );
and ( w_67 , w_66 , \89_b1 );
or ( \91_b1 , \A[1][5]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_68 );
and ( \91_b0 , \A[1][5]_b0 , w_69 );
and ( w_68 , w_69 , \I[0]_b0 );
or ( \92_b1 , \A[2][5]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_70 );
and ( \92_b0 , \A[2][5]_b0 , w_71 );
and ( w_70 , w_71 , \I[1]_b0 );
or ( \93_b1 , \91_b1 , w_73 );
not ( w_73 , w_74 );
and ( \93_b0 , \91_b0 , w_75 );
and ( w_74 ,  , w_75 );
buf ( w_73 , \92_b1 );
not ( w_73 , w_76 );
not (  , w_77 );
and ( w_76 , w_77 , \92_b0 );
or ( \94_b1 , \90_b1 , w_79 );
not ( w_79 , w_80 );
and ( \94_b0 , \90_b0 , w_81 );
and ( w_80 ,  , w_81 );
buf ( w_79 , \93_b1 );
not ( w_79 , w_82 );
not (  , w_83 );
and ( w_82 , w_83 , \93_b0 );
buf ( \95_b1 , \94_b1 );
buf ( \95_b0 , \94_b0 );
or ( \96_b1 , \I[1]_b1 , w_85 );
not ( w_85 , w_86 );
and ( \96_b0 , \I[1]_b0 , w_87 );
and ( w_86 ,  , w_87 );
buf ( w_85 , \I[0]_b1 );
not ( w_85 , w_88 );
not (  , w_89 );
and ( w_88 , w_89 , \I[0]_b0 );
buf ( \97_b1 , \96_b1 );
not ( \97_b1 , w_90 );
not ( \97_b0 , w_91 );
and ( w_90 , w_91 , \96_b0 );
buf ( \98_b1 , \A[0][2]_b1 );
not ( \98_b1 , w_92 );
not ( \98_b0 , w_93 );
and ( w_92 , w_93 , \A[0][2]_b0 );
or ( \99_b1 , \97_b1 , w_94 );
or ( \99_b0 , \97_b0 , \98_b0 );
not ( \98_b0 , w_95 );
and ( w_95 , w_94 , \98_b1 );
or ( \100_b1 , \A[1][2]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_96 );
and ( \100_b0 , \A[1][2]_b0 , w_97 );
and ( w_96 , w_97 , \I[0]_b0 );
or ( \101_b1 , \A[2][2]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_98 );
and ( \101_b0 , \A[2][2]_b0 , w_99 );
and ( w_98 , w_99 , \I[1]_b0 );
or ( \102_b1 , \100_b1 , w_101 );
not ( w_101 , w_102 );
and ( \102_b0 , \100_b0 , w_103 );
and ( w_102 ,  , w_103 );
buf ( w_101 , \101_b1 );
not ( w_101 , w_104 );
not (  , w_105 );
and ( w_104 , w_105 , \101_b0 );
or ( \103_b1 , \99_b1 , w_107 );
not ( w_107 , w_108 );
and ( \103_b0 , \99_b0 , w_109 );
and ( w_108 ,  , w_109 );
buf ( w_107 , \102_b1 );
not ( w_107 , w_110 );
not (  , w_111 );
and ( w_110 , w_111 , \102_b0 );
buf ( \104_b1 , \103_b1 );
buf ( \104_b0 , \103_b0 );
buf ( \105_b1 , \A[0][1]_b1 );
not ( \105_b1 , w_112 );
not ( \105_b0 , w_113 );
and ( w_112 , w_113 , \A[0][1]_b0 );
or ( \107_b1 , \A[2][1]_b1 , w_115 );
not ( w_115 , w_116 );
and ( \107_b0 , \A[2][1]_b0 , w_117 );
and ( w_116 ,  , w_117 );
buf ( w_115 , \I[1]_b1 );
not ( w_115 , w_118 );
not (  , w_119 );
and ( w_118 , w_119 , \I[1]_b0 );
or ( \108_b1 , \A[1][1]_b1 , w_121 );
not ( w_121 , w_122 );
and ( \108_b0 , \A[1][1]_b0 , w_123 );
and ( w_122 ,  , w_123 );
buf ( w_121 , \I[0]_b1 );
not ( w_121 , w_124 );
not (  , w_125 );
and ( w_124 , w_125 , \I[0]_b0 );
or ( \109_b1 , \107_b1 , w_127 );
not ( w_127 , w_128 );
and ( \109_b0 , \107_b0 , w_129 );
and ( w_128 ,  , w_129 );
buf ( w_127 , \108_b1 );
not ( w_127 , w_130 );
not (  , w_131 );
and ( w_130 , w_131 , \108_b0 );
or ( \110_b1 , \106_b1 , w_133 );
not ( w_133 , w_134 );
and ( \110_b0 , \106_b0 , w_135 );
and ( w_134 ,  , w_135 );
buf ( w_133 , \109_b1 );
not ( w_133 , w_136 );
not (  , w_137 );
and ( w_136 , w_137 , \109_b0 );
buf ( \111_b1 , \110_b1 );
not ( \111_b1 , w_138 );
not ( \111_b0 , w_139 );
and ( w_138 , w_139 , \110_b0 );
or ( \112_b1 , \I[1]_b1 , w_141 );
not ( w_141 , w_142 );
and ( \112_b0 , \I[1]_b0 , w_143 );
and ( w_142 ,  , w_143 );
buf ( w_141 , \I[0]_b1 );
not ( w_141 , w_144 );
not (  , w_145 );
and ( w_144 , w_145 , \I[0]_b0 );
or ( \113_b1 , \112_b1 , w_147 );
not ( w_147 , w_148 );
and ( \113_b0 , \112_b0 , w_149 );
and ( w_148 ,  , w_149 );
buf ( w_147 , \A[0][0]_b1 );
not ( w_147 , w_150 );
not (  , w_151 );
and ( w_150 , w_151 , \A[0][0]_b0 );
or ( \114_b1 , \A[1][0]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_152 );
and ( \114_b0 , \A[1][0]_b0 , w_153 );
and ( w_152 , w_153 , \I[0]_b0 );
or ( \115_b1 , \A[2][0]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_154 );
and ( \115_b0 , \A[2][0]_b0 , w_155 );
and ( w_154 , w_155 , \I[1]_b0 );
or ( \116_b1 , \114_b1 , w_157 );
not ( w_157 , w_158 );
and ( \116_b0 , \114_b0 , w_159 );
and ( w_158 ,  , w_159 );
buf ( w_157 , \115_b1 );
not ( w_157 , w_160 );
not (  , w_161 );
and ( w_160 , w_161 , \115_b0 );
or ( \117_b1 , \113_b1 , w_163 );
not ( w_163 , w_164 );
and ( \117_b0 , \113_b0 , w_165 );
and ( w_164 ,  , w_165 );
buf ( w_163 , \116_b1 );
not ( w_163 , w_166 );
not (  , w_167 );
and ( w_166 , w_167 , \116_b0 );
buf ( \118_b1 , \117_b1 );
buf ( \118_b0 , \117_b0 );
or ( \119_b1 , \I[1]_b1 , w_169 );
not ( w_169 , w_170 );
and ( \119_b0 , \I[1]_b0 , w_171 );
and ( w_170 ,  , w_171 );
buf ( w_169 , \I[0]_b1 );
not ( w_169 , w_172 );
not (  , w_173 );
and ( w_172 , w_173 , \I[0]_b0 );
buf ( \120_b1 , \119_b1 );
not ( \120_b1 , w_174 );
not ( \120_b0 , w_175 );
and ( w_174 , w_175 , \119_b0 );
buf ( \121_b1 , \A[0][4]_b1 );
not ( \121_b1 , w_176 );
not ( \121_b0 , w_177 );
and ( w_176 , w_177 , \A[0][4]_b0 );
or ( \122_b1 , \120_b1 , w_178 );
or ( \122_b0 , \120_b0 , \121_b0 );
not ( \121_b0 , w_179 );
and ( w_179 , w_178 , \121_b1 );
or ( \123_b1 , \A[1][4]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_180 );
and ( \123_b0 , \A[1][4]_b0 , w_181 );
and ( w_180 , w_181 , \I[0]_b0 );
or ( \124_b1 , \A[2][4]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_182 );
and ( \124_b0 , \A[2][4]_b0 , w_183 );
and ( w_182 , w_183 , \I[1]_b0 );
or ( \125_b1 , \123_b1 , w_185 );
not ( w_185 , w_186 );
and ( \125_b0 , \123_b0 , w_187 );
and ( w_186 ,  , w_187 );
buf ( w_185 , \124_b1 );
not ( w_185 , w_188 );
not (  , w_189 );
and ( w_188 , w_189 , \124_b0 );
or ( \126_b1 , \122_b1 , w_191 );
not ( w_191 , w_192 );
and ( \126_b0 , \122_b0 , w_193 );
and ( w_192 ,  , w_193 );
buf ( w_191 , \125_b1 );
not ( w_191 , w_194 );
not (  , w_195 );
and ( w_194 , w_195 , \125_b0 );
buf ( \127_b1 , \126_b1 );
buf ( \127_b0 , \126_b0 );
or ( \128_b1 , \I[1]_b1 , w_197 );
not ( w_197 , w_198 );
and ( \128_b0 , \I[1]_b0 , w_199 );
and ( w_198 ,  , w_199 );
buf ( w_197 , \I[0]_b1 );
not ( w_197 , w_200 );
not (  , w_201 );
and ( w_200 , w_201 , \I[0]_b0 );
buf ( \129_b1 , \128_b1 );
not ( \129_b1 , w_202 );
not ( \129_b0 , w_203 );
and ( w_202 , w_203 , \128_b0 );
buf ( \130_b1 , \A[0][6]_b1 );
not ( \130_b1 , w_204 );
not ( \130_b0 , w_205 );
and ( w_204 , w_205 , \A[0][6]_b0 );
or ( \131_b1 , \129_b1 , w_206 );
or ( \131_b0 , \129_b0 , \130_b0 );
not ( \130_b0 , w_207 );
and ( w_207 , w_206 , \130_b1 );
or ( \132_b1 , \A[1][6]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_208 );
and ( \132_b0 , \A[1][6]_b0 , w_209 );
and ( w_208 , w_209 , \I[0]_b0 );
or ( \133_b1 , \A[2][6]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_210 );
and ( \133_b0 , \A[2][6]_b0 , w_211 );
and ( w_210 , w_211 , \I[1]_b0 );
or ( \134_b1 , \132_b1 , w_213 );
not ( w_213 , w_214 );
and ( \134_b0 , \132_b0 , w_215 );
and ( w_214 ,  , w_215 );
buf ( w_213 , \133_b1 );
not ( w_213 , w_216 );
not (  , w_217 );
and ( w_216 , w_217 , \133_b0 );
or ( \135_b1 , \131_b1 , w_219 );
not ( w_219 , w_220 );
and ( \135_b0 , \131_b0 , w_221 );
and ( w_220 ,  , w_221 );
buf ( w_219 , \134_b1 );
not ( w_219 , w_222 );
not (  , w_223 );
and ( w_222 , w_223 , \134_b0 );
buf ( \136_b1 , \135_b1 );
buf ( \136_b0 , \135_b0 );
buf ( \137_b1 , \A[0][3]_b1 );
not ( \137_b1 , w_224 );
not ( \137_b0 , w_225 );
and ( w_224 , w_225 , \A[0][3]_b0 );
or ( \139_b1 , \A[2][3]_b1 , w_227 );
not ( w_227 , w_228 );
and ( \139_b0 , \A[2][3]_b0 , w_229 );
and ( w_228 ,  , w_229 );
buf ( w_227 , \I[1]_b1 );
not ( w_227 , w_230 );
not (  , w_231 );
and ( w_230 , w_231 , \I[1]_b0 );
or ( \140_b1 , \A[1][3]_b1 , w_233 );
not ( w_233 , w_234 );
and ( \140_b0 , \A[1][3]_b0 , w_235 );
and ( w_234 ,  , w_235 );
buf ( w_233 , \I[0]_b1 );
not ( w_233 , w_236 );
not (  , w_237 );
and ( w_236 , w_237 , \I[0]_b0 );
or ( \141_b1 , \139_b1 , w_239 );
not ( w_239 , w_240 );
and ( \141_b0 , \139_b0 , w_241 );
and ( w_240 ,  , w_241 );
buf ( w_239 , \140_b1 );
not ( w_239 , w_242 );
not (  , w_243 );
and ( w_242 , w_243 , \140_b0 );
or ( \142_b1 , \138_b1 , w_245 );
not ( w_245 , w_246 );
and ( \142_b0 , \138_b0 , w_247 );
and ( w_246 ,  , w_247 );
buf ( w_245 , \141_b1 );
not ( w_245 , w_248 );
not (  , w_249 );
and ( w_248 , w_249 , \141_b0 );
buf ( \143_b1 , \142_b1 );
not ( \143_b1 , w_250 );
not ( \143_b0 , w_251 );
and ( w_250 , w_251 , \142_b0 );
or ( \144_b1 , \A[1][8]_b1 , \I[0]_b1 );
not ( \I[0]_b1 , w_252 );
and ( \144_b0 , \A[1][8]_b0 , w_253 );
and ( w_252 , w_253 , \I[0]_b0 );
or ( \145_b1 , \A[2][8]_b1 , \I[1]_b1 );
not ( \I[1]_b1 , w_254 );
and ( \145_b0 , \A[2][8]_b0 , w_255 );
and ( w_254 , w_255 , \I[1]_b0 );
or ( \146_b1 , \144_b1 , w_257 );
not ( w_257 , w_258 );
and ( \146_b0 , \144_b0 , w_259 );
and ( w_258 ,  , w_259 );
buf ( w_257 , \145_b1 );
not ( w_257 , w_260 );
not (  , w_261 );
and ( w_260 , w_261 , \145_b0 );
or ( \147_b1 , \79_b1 , w_263 );
not ( w_263 , w_264 );
and ( \147_b0 , \79_b0 , w_265 );
and ( w_264 ,  , w_265 );
buf ( w_263 , \B[8]_b1 );
not ( w_263 , w_266 );
not (  , w_267 );
and ( w_266 , w_267 , \B[8]_b0 );
or ( \148_b1 , \I[1]_b1 , w_269 );
not ( w_269 , w_270 );
and ( \148_b0 , \I[1]_b0 , w_271 );
and ( w_270 ,  , w_271 );
buf ( w_269 , \I[0]_b1 );
not ( w_269 , w_272 );
not (  , w_273 );
and ( w_272 , w_273 , \I[0]_b0 );
buf ( \149_b1 , \148_b1 );
not ( \149_b1 , w_274 );
not ( \149_b0 , w_275 );
and ( w_274 , w_275 , \148_b0 );
buf ( \150_b1 , \A[0][8]_b1 );
not ( \150_b1 , w_276 );
not ( \150_b0 , w_277 );
and ( w_276 , w_277 , \A[0][8]_b0 );
or ( \151_b1 , \149_b1 , w_278 );
or ( \151_b0 , \149_b0 , \150_b0 );
not ( \150_b0 , w_279 );
and ( w_279 , w_278 , \150_b1 );
or ( \152_b1 , \151_b1 , w_281 );
not ( w_281 , w_282 );
and ( \152_b0 , \151_b0 , w_283 );
and ( w_282 ,  , w_283 );
buf ( w_281 , \146_b1 );
not ( w_281 , w_284 );
not (  , w_285 );
and ( w_284 , w_285 , \146_b0 );
buf ( \153_b1 , \152_b1 );
buf ( \153_b0 , \152_b0 );
or ( \154_b1 , \153_b1 , w_287 );
not ( w_287 , w_288 );
and ( \154_b0 , \153_b0 , w_289 );
and ( w_288 ,  , w_289 );
buf ( w_287 , \B[9]_b1 );
not ( w_287 , w_290 );
not (  , w_291 );
and ( w_290 , w_291 , \B[9]_b0 );
or ( \155_b1 , \147_b1 , \154_b1 );
xor ( \155_b0 , \147_b0 , w_292 );
not ( w_292 , w_293 );
and ( w_293 , \154_b1 , \154_b0 );
or ( \156_b1 , \79_b1 , w_295 );
not ( w_295 , w_296 );
and ( \156_b0 , \79_b0 , w_297 );
and ( w_296 ,  , w_297 );
buf ( w_295 , \B[7]_b1 );
not ( w_295 , w_298 );
not (  , w_299 );
and ( w_298 , w_299 , \B[7]_b0 );
or ( \157_b1 , \86_b1 , w_301 );
not ( w_301 , w_302 );
and ( \157_b0 , \86_b0 , w_303 );
and ( w_302 ,  , w_303 );
buf ( w_301 , \B[9]_b1 );
not ( w_301 , w_304 );
not (  , w_305 );
and ( w_304 , w_305 , \B[9]_b0 );
or ( \158_b1 , \156_b1 , \157_b1 );
xor ( \158_b0 , \156_b0 , w_306 );
not ( w_306 , w_307 );
and ( w_307 , \157_b1 , \157_b0 );
or ( \159_b1 , \153_b1 , w_309 );
not ( w_309 , w_310 );
and ( \159_b0 , \153_b0 , w_311 );
and ( w_310 ,  , w_311 );
buf ( w_309 , \B[8]_b1 );
not ( w_309 , w_312 );
not (  , w_313 );
and ( w_312 , w_313 , \B[8]_b0 );
or ( \160_b1 , \158_b1 , \159_b1 );
not ( \159_b1 , w_314 );
and ( \160_b0 , \158_b0 , w_315 );
and ( w_314 , w_315 , \159_b0 );
or ( \161_b1 , \156_b1 , \157_b1 );
not ( \157_b1 , w_316 );
and ( \161_b0 , \156_b0 , w_317 );
and ( w_316 , w_317 , \157_b0 );
or ( \162_b1 , \160_b1 , w_318 );
or ( \162_b0 , \160_b0 , \161_b0 );
not ( \161_b0 , w_319 );
and ( w_319 , w_318 , \161_b1 );
or ( \163_b1 , \155_b1 , \162_b1 );
not ( \162_b1 , w_320 );
and ( \163_b0 , \155_b0 , w_321 );
and ( w_320 , w_321 , \162_b0 );
or ( \164_b1 , \147_b1 , \154_b1 );
not ( \154_b1 , w_322 );
and ( \164_b0 , \147_b0 , w_323 );
and ( w_322 , w_323 , \154_b0 );
or ( \165_b1 , \163_b1 , w_324 );
or ( \165_b0 , \163_b0 , \164_b0 );
not ( \164_b0 , w_325 );
and ( w_325 , w_324 , \164_b1 );
or ( \166_b1 , \79_b1 , w_327 );
not ( w_327 , w_328 );
and ( \166_b0 , \79_b0 , w_329 );
and ( w_328 ,  , w_329 );
buf ( w_327 , \B[9]_b1 );
not ( w_327 , w_330 );
not (  , w_331 );
and ( w_330 , w_331 , \B[9]_b0 );
or ( \167_b1 , \165_b1 , w_333 );
not ( w_333 , w_334 );
and ( \167_b0 , \165_b0 , w_335 );
and ( w_334 ,  , w_335 );
buf ( w_333 , \166_b1 );
not ( w_333 , w_336 );
not (  , w_337 );
and ( w_336 , w_337 , \166_b0 );
buf ( \168_b1 , \167_b1 );
not ( \168_b1 , w_338 );
not ( \168_b0 , w_339 );
and ( w_338 , w_339 , \167_b0 );
or ( \169_b1 , \95_b1 , w_341 );
not ( w_341 , w_342 );
and ( \169_b0 , \95_b0 , w_343 );
and ( w_342 ,  , w_343 );
buf ( w_341 , \B[7]_b1 );
not ( w_341 , w_344 );
not (  , w_345 );
and ( w_344 , w_345 , \B[7]_b0 );
or ( \170_b1 , \127_b1 , w_347 );
not ( w_347 , w_348 );
and ( \170_b0 , \127_b0 , w_349 );
and ( w_348 ,  , w_349 );
buf ( w_347 , \B[8]_b1 );
not ( w_347 , w_350 );
not (  , w_351 );
and ( w_350 , w_351 , \B[8]_b0 );
or ( \171_b1 , \169_b1 , \170_b1 );
xor ( \171_b0 , \169_b0 , w_352 );
not ( w_352 , w_353 );
and ( w_353 , \170_b1 , \170_b0 );
or ( \172_b1 , \86_b1 , w_355 );
not ( w_355 , w_356 );
and ( \172_b0 , \86_b0 , w_357 );
and ( w_356 ,  , w_357 );
buf ( w_355 , \B[5]_b1 );
not ( w_355 , w_358 );
not (  , w_359 );
and ( w_358 , w_359 , \B[5]_b0 );
or ( \173_b1 , \171_b1 , \172_b1 );
xor ( \173_b0 , \171_b0 , w_360 );
not ( w_360 , w_361 );
and ( w_361 , \172_b1 , \172_b0 );
or ( \174_b1 , \79_b1 , w_363 );
not ( w_363 , w_364 );
and ( \174_b0 , \79_b0 , w_365 );
and ( w_364 ,  , w_365 );
buf ( w_363 , \B[3]_b1 );
not ( w_363 , w_366 );
not (  , w_367 );
and ( w_366 , w_367 , \B[3]_b0 );
or ( \175_b1 , \152_b1 , w_369 );
not ( w_369 , w_370 );
and ( \175_b0 , \152_b0 , w_371 );
and ( w_370 ,  , w_371 );
buf ( w_369 , \B[4]_b1 );
not ( w_369 , w_372 );
not (  , w_373 );
and ( w_372 , w_373 , \B[4]_b0 );
or ( \176_b1 , \174_b1 , \175_b1 );
xor ( \176_b0 , \174_b0 , w_374 );
not ( w_374 , w_375 );
and ( w_375 , \175_b1 , \175_b0 );
or ( \177_b1 , \136_b1 , \B[6]_b1 );
not ( \B[6]_b1 , w_376 );
and ( \177_b0 , \136_b0 , w_377 );
and ( w_376 , w_377 , \B[6]_b0 );
or ( \178_b1 , \176_b1 , w_378 );
xor ( \178_b0 , \176_b0 , w_380 );
not ( w_380 , w_381 );
and ( w_381 , w_378 , w_379 );
buf ( w_378 , \177_b1 );
not ( w_378 , w_382 );
not ( w_379 , w_383 );
and ( w_382 , w_383 , \177_b0 );
or ( \179_b1 , \173_b1 , \178_b1 );
not ( \178_b1 , w_384 );
and ( \179_b0 , \173_b0 , w_385 );
and ( w_384 , w_385 , \178_b0 );
or ( \180_b1 , \143_b1 , w_387 );
not ( w_387 , w_388 );
and ( \180_b0 , \143_b0 , w_389 );
and ( w_388 ,  , w_389 );
buf ( w_387 , \B[8]_b1 );
not ( w_387 , w_390 );
not (  , w_391 );
and ( w_390 , w_391 , \B[8]_b0 );
or ( \181_b1 , \127_b1 , w_393 );
not ( w_393 , w_394 );
and ( \181_b0 , \127_b0 , w_395 );
and ( w_394 ,  , w_395 );
buf ( w_393 , \B[7]_b1 );
not ( w_393 , w_396 );
not (  , w_397 );
and ( w_396 , w_397 , \B[7]_b0 );
or ( \182_b1 , \180_b1 , \181_b1 );
xor ( \182_b0 , \180_b0 , w_398 );
not ( w_398 , w_399 );
and ( w_399 , \181_b1 , \181_b0 );
or ( \183_b1 , \79_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_400 );
and ( \183_b0 , \79_b0 , w_401 );
and ( w_400 , w_401 , \B[1]_b0 );
or ( \184_b1 , \152_b1 , \B[2]_b1 );
not ( \B[2]_b1 , w_402 );
and ( \184_b0 , \152_b0 , w_403 );
and ( w_402 , w_403 , \B[2]_b0 );
or ( \185_b1 , \183_b1 , w_405 );
not ( w_405 , w_406 );
and ( \185_b0 , \183_b0 , w_407 );
and ( w_406 ,  , w_407 );
buf ( w_405 , \184_b1 );
not ( w_405 , w_408 );
not (  , w_409 );
and ( w_408 , w_409 , \184_b0 );
or ( \186_b1 , \182_b1 , \185_b1 );
not ( \185_b1 , w_410 );
and ( \186_b0 , \182_b0 , w_411 );
and ( w_410 , w_411 , \185_b0 );
or ( \187_b1 , \180_b1 , \181_b1 );
not ( \181_b1 , w_412 );
and ( \187_b0 , \180_b0 , w_413 );
and ( w_412 , w_413 , \181_b0 );
or ( \188_b1 , \186_b1 , w_414 );
or ( \188_b0 , \186_b0 , \187_b0 );
not ( \187_b0 , w_415 );
and ( w_415 , w_414 , \187_b1 );
or ( \189_b1 , \179_b1 , w_417 );
not ( w_417 , w_418 );
and ( \189_b0 , \179_b0 , w_419 );
and ( w_418 ,  , w_419 );
buf ( w_417 , \188_b1 );
not ( w_417 , w_420 );
not (  , w_421 );
and ( w_420 , w_421 , \188_b0 );
buf ( \190_b1 , \178_b1 );
not ( \190_b1 , w_422 );
not ( \190_b0 , w_423 );
and ( w_422 , w_423 , \178_b0 );
buf ( \191_b1 , \173_b1 );
not ( \191_b1 , w_424 );
not ( \191_b0 , w_425 );
and ( w_424 , w_425 , \173_b0 );
or ( \192_b1 , \190_b1 , \191_b1 );
not ( \191_b1 , w_426 );
and ( \192_b0 , \190_b0 , w_427 );
and ( w_426 , w_427 , \191_b0 );
or ( \193_b1 , \189_b1 , w_429 );
not ( w_429 , w_430 );
and ( \193_b0 , \189_b0 , w_431 );
and ( w_430 ,  , w_431 );
buf ( w_429 , \192_b1 );
not ( w_429 , w_432 );
not (  , w_433 );
and ( w_432 , w_433 , \192_b0 );
buf ( \194_b1 , \193_b1 );
not ( \194_b1 , w_434 );
not ( \194_b0 , w_435 );
and ( w_434 , w_435 , \193_b0 );
or ( \195_b1 , \95_b1 , w_437 );
not ( w_437 , w_438 );
and ( \195_b0 , \95_b0 , w_439 );
and ( w_438 ,  , w_439 );
buf ( w_437 , \B[8]_b1 );
not ( w_437 , w_440 );
not (  , w_441 );
and ( w_440 , w_441 , \B[8]_b0 );
or ( \196_b1 , \127_b1 , w_443 );
not ( w_443 , w_444 );
and ( \196_b0 , \127_b0 , w_445 );
and ( w_444 ,  , w_445 );
buf ( w_443 , \B[9]_b1 );
not ( w_443 , w_446 );
not (  , w_447 );
and ( w_446 , w_447 , \B[9]_b0 );
or ( \197_b1 , \195_b1 , \196_b1 );
xor ( \197_b0 , \195_b0 , w_448 );
not ( w_448 , w_449 );
and ( w_449 , \196_b1 , \196_b0 );
or ( \198_b1 , \86_b1 , w_451 );
not ( w_451 , w_452 );
and ( \198_b0 , \86_b0 , w_453 );
and ( w_452 ,  , w_453 );
buf ( w_451 , \B[6]_b1 );
not ( w_451 , w_454 );
not (  , w_455 );
and ( w_454 , w_455 , \B[6]_b0 );
or ( \199_b1 , \197_b1 , \198_b1 );
xor ( \199_b0 , \197_b0 , w_456 );
not ( w_456 , w_457 );
and ( w_457 , \198_b1 , \198_b0 );
buf ( \200_b1 , \143_b1 );
buf ( \200_b0 , \143_b0 );
or ( \201_b1 , \200_b1 , w_459 );
not ( w_459 , w_460 );
and ( \201_b0 , \200_b0 , w_461 );
and ( w_460 ,  , w_461 );
buf ( w_459 , \B[9]_b1 );
not ( w_459 , w_462 );
not (  , w_463 );
and ( w_462 , w_463 , \B[9]_b0 );
or ( \202_b1 , \152_b1 , w_465 );
not ( w_465 , w_466 );
and ( \202_b0 , \152_b0 , w_467 );
and ( w_466 ,  , w_467 );
buf ( w_465 , \B[3]_b1 );
not ( w_465 , w_468 );
not (  , w_469 );
and ( w_468 , w_469 , \B[3]_b0 );
or ( \203_b1 , \136_b1 , w_471 );
not ( w_471 , w_472 );
and ( \203_b0 , \136_b0 , w_473 );
and ( w_472 ,  , w_473 );
buf ( w_471 , \B[5]_b1 );
not ( w_471 , w_474 );
not (  , w_475 );
and ( w_474 , w_475 , \B[5]_b0 );
or ( \204_b1 , \202_b1 , \203_b1 );
xor ( \204_b0 , \202_b0 , w_476 );
not ( w_476 , w_477 );
and ( w_477 , \203_b1 , \203_b0 );
or ( \205_b1 , \79_b1 , w_479 );
not ( w_479 , w_480 );
and ( \205_b0 , \79_b0 , w_481 );
and ( w_480 ,  , w_481 );
buf ( w_479 , \B[2]_b1 );
not ( w_479 , w_482 );
not (  , w_483 );
and ( w_482 , w_483 , \B[2]_b0 );
or ( \206_b1 , \204_b1 , \205_b1 );
not ( \205_b1 , w_484 );
and ( \206_b0 , \204_b0 , w_485 );
and ( w_484 , w_485 , \205_b0 );
or ( \207_b1 , \202_b1 , \203_b1 );
not ( \203_b1 , w_486 );
and ( \207_b0 , \202_b0 , w_487 );
and ( w_486 , w_487 , \203_b0 );
or ( \208_b1 , \206_b1 , w_488 );
or ( \208_b0 , \206_b0 , \207_b0 );
not ( \207_b0 , w_489 );
and ( w_489 , w_488 , \207_b1 );
or ( \209_b1 , \201_b1 , \208_b1 );
xor ( \209_b0 , \201_b0 , w_490 );
not ( w_490 , w_491 );
and ( w_491 , \208_b1 , \208_b0 );
or ( \210_b1 , \95_b1 , w_493 );
not ( w_493 , w_494 );
and ( \210_b0 , \95_b0 , w_495 );
and ( w_494 ,  , w_495 );
buf ( w_493 , \B[6]_b1 );
not ( w_493 , w_496 );
not (  , w_497 );
and ( w_496 , w_497 , \B[6]_b0 );
or ( \211_b1 , \104_b1 , w_499 );
not ( w_499 , w_500 );
and ( \211_b0 , \104_b0 , w_501 );
and ( w_500 ,  , w_501 );
buf ( w_499 , \B[9]_b1 );
not ( w_499 , w_502 );
not (  , w_503 );
and ( w_502 , w_503 , \B[9]_b0 );
or ( \212_b1 , \210_b1 , \211_b1 );
xor ( \212_b0 , \210_b0 , w_504 );
not ( w_504 , w_505 );
and ( w_505 , \211_b1 , \211_b0 );
or ( \213_b1 , \86_b1 , w_507 );
not ( w_507 , w_508 );
and ( \213_b0 , \86_b0 , w_509 );
and ( w_508 ,  , w_509 );
buf ( w_507 , \B[4]_b1 );
not ( w_507 , w_510 );
not (  , w_511 );
and ( w_510 , w_511 , \B[4]_b0 );
or ( \214_b1 , \212_b1 , \213_b1 );
not ( \213_b1 , w_512 );
and ( \214_b0 , \212_b0 , w_513 );
and ( w_512 , w_513 , \213_b0 );
or ( \215_b1 , \210_b1 , \211_b1 );
not ( \211_b1 , w_514 );
and ( \215_b0 , \210_b0 , w_515 );
and ( w_514 , w_515 , \211_b0 );
or ( \216_b1 , \214_b1 , w_516 );
or ( \216_b0 , \214_b0 , \215_b0 );
not ( \215_b0 , w_517 );
and ( w_517 , w_516 , \215_b1 );
or ( \217_b1 , \209_b1 , \216_b1 );
not ( \216_b1 , w_518 );
and ( \217_b0 , \209_b0 , w_519 );
and ( w_518 , w_519 , \216_b0 );
or ( \218_b1 , \201_b1 , \208_b1 );
not ( \208_b1 , w_520 );
and ( \218_b0 , \201_b0 , w_521 );
and ( w_520 , w_521 , \208_b0 );
or ( \219_b1 , \217_b1 , w_522 );
or ( \219_b0 , \217_b0 , \218_b0 );
not ( \218_b0 , w_523 );
and ( w_523 , w_522 , \218_b1 );
or ( \220_b1 , \199_b1 , \219_b1 );
xor ( \220_b0 , \199_b0 , w_524 );
not ( w_524 , w_525 );
and ( w_525 , \219_b1 , \219_b0 );
buf ( \221_b1 , \175_b1 );
not ( \221_b1 , w_526 );
not ( \221_b0 , w_527 );
and ( w_526 , w_527 , \175_b0 );
buf ( \222_b1 , \174_b1 );
not ( \222_b1 , w_528 );
not ( \222_b0 , w_529 );
and ( w_528 , w_529 , \174_b0 );
or ( \223_b1 , \221_b1 , w_530 );
or ( \223_b0 , \221_b0 , \222_b0 );
not ( \222_b0 , w_531 );
and ( w_531 , w_530 , \222_b1 );
or ( \224_b1 , \223_b1 , w_533 );
not ( w_533 , w_534 );
and ( \224_b0 , \223_b0 , w_535 );
and ( w_534 ,  , w_535 );
buf ( w_533 , \177_b1 );
not ( w_533 , w_536 );
not (  , w_537 );
and ( w_536 , w_537 , \177_b0 );
buf ( \225_b1 , \174_b1 );
not ( \225_b1 , w_538 );
not ( \225_b0 , w_539 );
and ( w_538 , w_539 , \174_b0 );
buf ( \226_b1 , \175_b1 );
not ( \226_b1 , w_540 );
not ( \226_b0 , w_541 );
and ( w_540 , w_541 , \175_b0 );
or ( \227_b1 , \225_b1 , w_543 );
not ( w_543 , w_544 );
and ( \227_b0 , \225_b0 , w_545 );
and ( w_544 ,  , w_545 );
buf ( w_543 , \226_b1 );
not ( w_543 , w_546 );
not (  , w_547 );
and ( w_546 , w_547 , \226_b0 );
or ( \228_b1 , \224_b1 , w_549 );
not ( w_549 , w_550 );
and ( \228_b0 , \224_b0 , w_551 );
and ( w_550 ,  , w_551 );
buf ( w_549 , \227_b1 );
not ( w_549 , w_552 );
not (  , w_553 );
and ( w_552 , w_553 , \227_b0 );
buf ( \229_b1 , \228_b1 );
not ( \229_b1 , w_554 );
not ( \229_b0 , w_555 );
and ( w_554 , w_555 , \228_b0 );
buf ( \230_b1 , \229_b1 );
not ( \230_b1 , w_556 );
not ( \230_b0 , w_557 );
and ( w_556 , w_557 , \229_b0 );
or ( \231_b1 , \169_b1 , \172_b1 );
not ( \172_b1 , w_558 );
and ( \231_b0 , \169_b0 , w_559 );
and ( w_558 , w_559 , \172_b0 );
or ( \232_b1 , \231_b1 , w_560 );
or ( \232_b0 , \231_b0 , \170_b0 );
not ( \170_b0 , w_561 );
and ( w_561 , w_560 , \170_b1 );
or ( \233_b1 , \172_b1 , w_562 );
or ( \233_b0 , \172_b0 , \169_b0 );
not ( \169_b0 , w_563 );
and ( w_563 , w_562 , \169_b1 );
or ( \234_b1 , \232_b1 , w_565 );
not ( w_565 , w_566 );
and ( \234_b0 , \232_b0 , w_567 );
and ( w_566 ,  , w_567 );
buf ( w_565 , \233_b1 );
not ( w_565 , w_568 );
not (  , w_569 );
and ( w_568 , w_569 , \233_b0 );
buf ( \235_b1 , \234_b1 );
not ( \235_b1 , w_570 );
not ( \235_b0 , w_571 );
and ( w_570 , w_571 , \234_b0 );
or ( \236_b1 , \230_b1 , \235_b1 );
not ( \235_b1 , w_572 );
and ( \236_b0 , \230_b0 , w_573 );
and ( w_572 , w_573 , \235_b0 );
buf ( \237_b1 , \228_b1 );
not ( \237_b1 , w_574 );
not ( \237_b0 , w_575 );
and ( w_574 , w_575 , \228_b0 );
or ( \238_b1 , \234_b1 , \237_b1 );
not ( \237_b1 , w_576 );
and ( \238_b0 , \234_b0 , w_577 );
and ( w_576 , w_577 , \237_b0 );
or ( \239_b1 , \236_b1 , w_579 );
not ( w_579 , w_580 );
and ( \239_b0 , \236_b0 , w_581 );
and ( w_580 ,  , w_581 );
buf ( w_579 , \238_b1 );
not ( w_579 , w_582 );
not (  , w_583 );
and ( w_582 , w_583 , \238_b0 );
buf ( \240_b1 , \239_b1 );
not ( \240_b1 , w_584 );
not ( \240_b0 , w_585 );
and ( w_584 , w_585 , \239_b0 );
or ( \241_b1 , \153_b1 , w_587 );
not ( w_587 , w_588 );
and ( \241_b0 , \153_b0 , w_589 );
and ( w_588 ,  , w_589 );
buf ( w_587 , \B[5]_b1 );
not ( w_587 , w_590 );
not (  , w_591 );
and ( w_590 , w_591 , \B[5]_b0 );
or ( \242_b1 , \79_b1 , w_593 );
not ( w_593 , w_594 );
and ( \242_b0 , \79_b0 , w_595 );
and ( w_594 ,  , w_595 );
buf ( w_593 , \B[4]_b1 );
not ( w_593 , w_596 );
not (  , w_597 );
and ( w_596 , w_597 , \B[4]_b0 );
or ( \243_b1 , \241_b1 , \242_b1 );
xor ( \243_b0 , \241_b0 , w_598 );
not ( w_598 , w_599 );
and ( w_599 , \242_b1 , \242_b0 );
or ( \244_b1 , \136_b1 , w_601 );
not ( w_601 , w_602 );
and ( \244_b0 , \136_b0 , w_603 );
and ( w_602 ,  , w_603 );
buf ( w_601 , \B[7]_b1 );
not ( w_601 , w_604 );
not (  , w_605 );
and ( w_604 , w_605 , \B[7]_b0 );
or ( \245_b1 , \243_b1 , \244_b1 );
xor ( \245_b0 , \243_b0 , w_606 );
not ( w_606 , w_607 );
and ( w_607 , \244_b1 , \244_b0 );
buf ( \246_b1 , \245_b1 );
not ( \246_b1 , w_608 );
not ( \246_b0 , w_609 );
and ( w_608 , w_609 , \245_b0 );
buf ( \247_b1 , \246_b1 );
not ( \247_b1 , w_610 );
not ( \247_b0 , w_611 );
and ( w_610 , w_611 , \246_b0 );
or ( \248_b1 , \240_b1 , w_612 );
or ( \248_b0 , \240_b0 , \247_b0 );
not ( \247_b0 , w_613 );
and ( w_613 , w_612 , \247_b1 );
buf ( \249_b1 , \239_b1 );
not ( \249_b1 , w_614 );
not ( \249_b0 , w_615 );
and ( w_614 , w_615 , \239_b0 );
or ( \250_b1 , \249_b1 , w_617 );
not ( w_617 , w_618 );
and ( \250_b0 , \249_b0 , w_619 );
and ( w_618 ,  , w_619 );
buf ( w_617 , \245_b1 );
not ( w_617 , w_620 );
not (  , w_621 );
and ( w_620 , w_621 , \245_b0 );
or ( \251_b1 , \248_b1 , w_623 );
not ( w_623 , w_624 );
and ( \251_b0 , \248_b0 , w_625 );
and ( w_624 ,  , w_625 );
buf ( w_623 , \250_b1 );
not ( w_623 , w_626 );
not (  , w_627 );
and ( w_626 , w_627 , \250_b0 );
or ( \252_b1 , \220_b1 , w_628 );
xor ( \252_b0 , \220_b0 , w_630 );
not ( w_630 , w_631 );
and ( w_631 , w_628 , w_629 );
buf ( w_628 , \251_b1 );
not ( w_628 , w_632 );
not ( w_629 , w_633 );
and ( w_632 , w_633 , \251_b0 );
buf ( \253_b1 , \252_b1 );
not ( \253_b1 , w_634 );
not ( \253_b0 , w_635 );
and ( w_634 , w_635 , \252_b0 );
or ( \254_b1 , \194_b1 , w_636 );
or ( \254_b0 , \194_b0 , \253_b0 );
not ( \253_b0 , w_637 );
and ( w_637 , w_636 , \253_b1 );
or ( \255_b1 , \201_b1 , \208_b1 );
xor ( \255_b0 , \201_b0 , w_638 );
not ( w_638 , w_639 );
and ( w_639 , \208_b1 , \208_b0 );
or ( \256_b1 , \255_b1 , \216_b1 );
xor ( \256_b0 , \255_b0 , w_640 );
not ( w_640 , w_641 );
and ( w_641 , \216_b1 , \216_b0 );
or ( \257_b1 , \202_b1 , \203_b1 );
xor ( \257_b0 , \202_b0 , w_642 );
not ( w_642 , w_643 );
and ( w_643 , \203_b1 , \203_b0 );
or ( \258_b1 , \257_b1 , \205_b1 );
xor ( \258_b0 , \257_b0 , w_644 );
not ( w_644 , w_645 );
and ( w_645 , \205_b1 , \205_b0 );
buf ( \259_b1 , \258_b1 );
not ( \259_b1 , w_646 );
not ( \259_b0 , w_647 );
and ( w_646 , w_647 , \258_b0 );
or ( \260_b1 , \136_b1 , w_649 );
not ( w_649 , w_650 );
and ( \260_b0 , \136_b0 , w_651 );
and ( w_650 ,  , w_651 );
buf ( w_649 , \B[4]_b1 );
not ( w_649 , w_652 );
not (  , w_653 );
and ( w_652 , w_653 , \B[4]_b0 );
buf ( \261_b1 , \260_b1 );
not ( \261_b1 , w_654 );
not ( \261_b0 , w_655 );
and ( w_654 , w_655 , \260_b0 );
or ( \262_b1 , \104_b1 , w_657 );
not ( w_657 , w_658 );
and ( \262_b0 , \104_b0 , w_659 );
and ( w_658 ,  , w_659 );
buf ( w_657 , \B[8]_b1 );
not ( w_657 , w_660 );
not (  , w_661 );
and ( w_660 , w_661 , \B[8]_b0 );
buf ( \263_b1 , \262_b1 );
not ( \263_b1 , w_662 );
not ( \263_b0 , w_663 );
and ( w_662 , w_663 , \262_b0 );
or ( \264_b1 , \261_b1 , w_664 );
or ( \264_b0 , \261_b0 , \263_b0 );
not ( \263_b0 , w_665 );
and ( w_665 , w_664 , \263_b1 );
or ( \265_b1 , \111_b1 , \B[9]_b1 );
not ( \B[9]_b1 , w_666 );
and ( \265_b0 , \111_b0 , w_667 );
and ( w_666 , w_667 , \B[9]_b0 );
or ( \266_b1 , \264_b1 , w_669 );
not ( w_669 , w_670 );
and ( \266_b0 , \264_b0 , w_671 );
and ( w_670 ,  , w_671 );
buf ( w_669 , \265_b1 );
not ( w_669 , w_672 );
not (  , w_673 );
and ( w_672 , w_673 , \265_b0 );
buf ( \267_b1 , \260_b1 );
not ( \267_b1 , w_674 );
not ( \267_b0 , w_675 );
and ( w_674 , w_675 , \260_b0 );
buf ( \268_b1 , \262_b1 );
not ( \268_b1 , w_676 );
not ( \268_b0 , w_677 );
and ( w_676 , w_677 , \262_b0 );
or ( \269_b1 , \267_b1 , w_679 );
not ( w_679 , w_680 );
and ( \269_b0 , \267_b0 , w_681 );
and ( w_680 ,  , w_681 );
buf ( w_679 , \268_b1 );
not ( w_679 , w_682 );
not (  , w_683 );
and ( w_682 , w_683 , \268_b0 );
or ( \270_b1 , \266_b1 , w_685 );
not ( w_685 , w_686 );
and ( \270_b0 , \266_b0 , w_687 );
and ( w_686 ,  , w_687 );
buf ( w_685 , \269_b1 );
not ( w_685 , w_688 );
not (  , w_689 );
and ( w_688 , w_689 , \269_b0 );
or ( \271_b1 , \259_b1 , w_691 );
not ( w_691 , w_692 );
and ( \271_b0 , \259_b0 , w_693 );
and ( w_692 ,  , w_693 );
buf ( w_691 , \270_b1 );
not ( w_691 , w_694 );
not (  , w_695 );
and ( w_694 , w_695 , \270_b0 );
buf ( \272_b1 , \270_b1 );
not ( \272_b1 , w_696 );
not ( \272_b0 , w_697 );
and ( w_696 , w_697 , \270_b0 );
buf ( \273_b1 , \272_b1 );
not ( \273_b1 , w_698 );
not ( \273_b0 , w_699 );
and ( w_698 , w_699 , \272_b0 );
buf ( \274_b1 , \258_b1 );
not ( \274_b1 , w_700 );
not ( \274_b0 , w_701 );
and ( w_700 , w_701 , \258_b0 );
or ( \275_b1 , \273_b1 , w_702 );
or ( \275_b0 , \273_b0 , \274_b0 );
not ( \274_b0 , w_703 );
and ( w_703 , w_702 , \274_b1 );
or ( \276_b1 , \95_b1 , w_705 );
not ( w_705 , w_706 );
and ( \276_b0 , \95_b0 , w_707 );
and ( w_706 ,  , w_707 );
buf ( w_705 , \B[5]_b1 );
not ( w_705 , w_708 );
not (  , w_709 );
and ( w_708 , w_709 , \B[5]_b0 );
buf ( \277_b1 , \276_b1 );
not ( \277_b1 , w_710 );
not ( \277_b0 , w_711 );
and ( w_710 , w_711 , \276_b0 );
or ( \278_b1 , \86_b1 , w_713 );
not ( w_713 , w_714 );
and ( \278_b0 , \86_b0 , w_715 );
and ( w_714 ,  , w_715 );
buf ( w_713 , \B[3]_b1 );
not ( w_713 , w_716 );
not (  , w_717 );
and ( w_716 , w_717 , \B[3]_b0 );
buf ( \279_b1 , \278_b1 );
not ( \279_b1 , w_718 );
not ( \279_b0 , w_719 );
and ( w_718 , w_719 , \278_b0 );
or ( \280_b1 , \277_b1 , w_720 );
or ( \280_b0 , \277_b0 , \279_b0 );
not ( \279_b0 , w_721 );
and ( w_721 , w_720 , \279_b1 );
or ( \281_b1 , \127_b1 , w_723 );
not ( w_723 , w_724 );
and ( \281_b0 , \127_b0 , w_725 );
and ( w_724 ,  , w_725 );
buf ( w_723 , \B[6]_b1 );
not ( w_723 , w_726 );
not (  , w_727 );
and ( w_726 , w_727 , \B[6]_b0 );
buf ( \282_b1 , \281_b1 );
not ( \282_b1 , w_728 );
not ( \282_b0 , w_729 );
and ( w_728 , w_729 , \281_b0 );
or ( \283_b1 , \280_b1 , w_731 );
not ( w_731 , w_732 );
and ( \283_b0 , \280_b0 , w_733 );
and ( w_732 ,  , w_733 );
buf ( w_731 , \282_b1 );
not ( w_731 , w_734 );
not (  , w_735 );
and ( w_734 , w_735 , \282_b0 );
or ( \284_b1 , \278_b1 , w_736 );
or ( \284_b0 , \278_b0 , \276_b0 );
not ( \276_b0 , w_737 );
and ( w_737 , w_736 , \276_b1 );
or ( \285_b1 , \283_b1 , w_739 );
not ( w_739 , w_740 );
and ( \285_b0 , \283_b0 , w_741 );
and ( w_740 ,  , w_741 );
buf ( w_739 , \284_b1 );
not ( w_739 , w_742 );
not (  , w_743 );
and ( w_742 , w_743 , \284_b0 );
or ( \286_b1 , \275_b1 , w_745 );
not ( w_745 , w_746 );
and ( \286_b0 , \275_b0 , w_747 );
and ( w_746 ,  , w_747 );
buf ( w_745 , \285_b1 );
not ( w_745 , w_748 );
not (  , w_749 );
and ( w_748 , w_749 , \285_b0 );
or ( \287_b1 , \271_b1 , \286_b1 );
not ( \286_b1 , w_750 );
and ( \287_b0 , \271_b0 , w_751 );
and ( w_750 , w_751 , \286_b0 );
or ( \288_b1 , \256_b1 , \287_b1 );
xor ( \288_b0 , \256_b0 , w_752 );
not ( w_752 , w_753 );
and ( w_753 , \287_b1 , \287_b0 );
or ( \289_b1 , \210_b1 , \211_b1 );
xor ( \289_b0 , \210_b0 , w_754 );
not ( w_754 , w_755 );
and ( w_755 , \211_b1 , \211_b0 );
or ( \290_b1 , \289_b1 , \213_b1 );
xor ( \290_b0 , \289_b0 , w_756 );
not ( w_756 , w_757 );
and ( w_757 , \213_b1 , \213_b0 );
or ( \291_b1 , \180_b1 , \181_b1 );
xor ( \291_b0 , \180_b0 , w_758 );
not ( w_758 , w_759 );
and ( w_759 , \181_b1 , \181_b0 );
or ( \292_b1 , \291_b1 , \185_b1 );
xor ( \292_b0 , \291_b0 , w_760 );
not ( w_760 , w_761 );
and ( w_761 , \185_b1 , \185_b0 );
or ( \293_b1 , \290_b1 , \292_b1 );
xor ( \293_b0 , \290_b0 , w_762 );
not ( w_762 , w_763 );
and ( w_763 , \292_b1 , \292_b0 );
or ( \294_b1 , \200_b1 , w_765 );
not ( w_765 , w_766 );
and ( \294_b0 , \200_b0 , w_767 );
and ( w_766 ,  , w_767 );
buf ( w_765 , \B[7]_b1 );
not ( w_765 , w_768 );
not (  , w_769 );
and ( w_768 , w_769 , \B[7]_b0 );
or ( \295_b1 , \79_b1 , w_771 );
not ( w_771 , w_772 );
and ( \295_b0 , \79_b0 , w_773 );
and ( w_772 ,  , w_773 );
buf ( w_771 , \B[0]_b1 );
not ( w_771 , w_774 );
not (  , w_775 );
and ( w_774 , w_775 , \B[0]_b0 );
buf ( \296_b1 , \295_b1 );
not ( \296_b1 , w_776 );
not ( \296_b0 , w_777 );
and ( w_776 , w_777 , \295_b0 );
or ( \297_b1 , \152_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_778 );
and ( \297_b0 , \152_b0 , w_779 );
and ( w_778 , w_779 , \B[1]_b0 );
or ( \298_b1 , \296_b1 , w_781 );
not ( w_781 , w_782 );
and ( \298_b0 , \296_b0 , w_783 );
and ( w_782 ,  , w_783 );
buf ( w_781 , \297_b1 );
not ( w_781 , w_784 );
not (  , w_785 );
and ( w_784 , w_785 , \297_b0 );
or ( \299_b1 , \294_b1 , \298_b1 );
xor ( \299_b0 , \294_b0 , w_786 );
not ( w_786 , w_787 );
and ( w_787 , \298_b1 , \298_b0 );
or ( \300_b1 , \184_b1 , w_788 );
xor ( \300_b0 , \184_b0 , w_790 );
not ( w_790 , w_791 );
and ( w_791 , w_788 , w_789 );
buf ( w_788 , \183_b1 );
not ( w_788 , w_792 );
not ( w_789 , w_793 );
and ( w_792 , w_793 , \183_b0 );
or ( \301_b1 , \299_b1 , \300_b1 );
not ( \300_b1 , w_794 );
and ( \301_b0 , \299_b0 , w_795 );
and ( w_794 , w_795 , \300_b0 );
or ( \302_b1 , \294_b1 , \298_b1 );
not ( \298_b1 , w_796 );
and ( \302_b0 , \294_b0 , w_797 );
and ( w_796 , w_797 , \298_b0 );
or ( \303_b1 , \301_b1 , w_798 );
or ( \303_b0 , \301_b0 , \302_b0 );
not ( \302_b0 , w_799 );
and ( w_799 , w_798 , \302_b1 );
or ( \304_b1 , \293_b1 , \303_b1 );
not ( \303_b1 , w_800 );
and ( \304_b0 , \293_b0 , w_801 );
and ( w_800 , w_801 , \303_b0 );
or ( \305_b1 , \290_b1 , \292_b1 );
not ( \292_b1 , w_802 );
and ( \305_b0 , \290_b0 , w_803 );
and ( w_802 , w_803 , \292_b0 );
or ( \306_b1 , \304_b1 , w_804 );
or ( \306_b0 , \304_b0 , \305_b0 );
not ( \305_b0 , w_805 );
and ( w_805 , w_804 , \305_b1 );
or ( \307_b1 , \288_b1 , \306_b1 );
not ( \306_b1 , w_806 );
and ( \307_b0 , \288_b0 , w_807 );
and ( w_806 , w_807 , \306_b0 );
or ( \308_b1 , \256_b1 , \287_b1 );
not ( \287_b1 , w_808 );
and ( \308_b0 , \256_b0 , w_809 );
and ( w_808 , w_809 , \287_b0 );
or ( \309_b1 , \307_b1 , w_810 );
or ( \309_b0 , \307_b0 , \308_b0 );
not ( \308_b0 , w_811 );
and ( w_811 , w_810 , \308_b1 );
buf ( \310_b1 , \309_b1 );
not ( \310_b1 , w_812 );
not ( \310_b0 , w_813 );
and ( w_812 , w_813 , \309_b0 );
or ( \311_b1 , \254_b1 , w_815 );
not ( w_815 , w_816 );
and ( \311_b0 , \254_b0 , w_817 );
and ( w_816 ,  , w_817 );
buf ( w_815 , \310_b1 );
not ( w_815 , w_818 );
not (  , w_819 );
and ( w_818 , w_819 , \310_b0 );
or ( \312_b1 , \252_b1 , w_820 );
or ( \312_b0 , \252_b0 , \193_b0 );
not ( \193_b0 , w_821 );
and ( w_821 , w_820 , \193_b1 );
or ( \313_b1 , \311_b1 , w_823 );
not ( w_823 , w_824 );
and ( \313_b0 , \311_b0 , w_825 );
and ( w_824 ,  , w_825 );
buf ( w_823 , \312_b1 );
not ( w_823 , w_826 );
not (  , w_827 );
and ( w_826 , w_827 , \312_b0 );
or ( \314_b1 , \245_b1 , w_829 );
not ( w_829 , w_830 );
and ( \314_b0 , \245_b0 , w_831 );
and ( w_830 ,  , w_831 );
buf ( w_829 , \237_b1 );
not ( w_829 , w_832 );
not (  , w_833 );
and ( w_832 , w_833 , \237_b0 );
buf ( \315_b1 , \314_b1 );
not ( \315_b1 , w_834 );
not ( \315_b0 , w_835 );
and ( w_834 , w_835 , \314_b0 );
buf ( \316_b1 , \234_b1 );
not ( \316_b1 , w_836 );
not ( \316_b0 , w_837 );
and ( w_836 , w_837 , \234_b0 );
or ( \317_b1 , \315_b1 , w_838 );
or ( \317_b0 , \315_b0 , \316_b0 );
not ( \316_b0 , w_839 );
and ( w_839 , w_838 , \316_b1 );
or ( \318_b1 , \245_b1 , w_840 );
or ( \318_b0 , \245_b0 , \237_b0 );
not ( \237_b0 , w_841 );
and ( w_841 , w_840 , \237_b1 );
or ( \319_b1 , \317_b1 , w_843 );
not ( w_843 , w_844 );
and ( \319_b0 , \317_b0 , w_845 );
and ( w_844 ,  , w_845 );
buf ( w_843 , \318_b1 );
not ( w_843 , w_846 );
not (  , w_847 );
and ( w_846 , w_847 , \318_b0 );
or ( \320_b1 , \136_b1 , w_849 );
not ( w_849 , w_850 );
and ( \320_b0 , \136_b0 , w_851 );
and ( w_850 ,  , w_851 );
buf ( w_849 , \B[8]_b1 );
not ( w_849 , w_852 );
not (  , w_853 );
and ( w_852 , w_853 , \B[8]_b0 );
or ( \321_b1 , \79_b1 , w_855 );
not ( w_855 , w_856 );
and ( \321_b0 , \79_b0 , w_857 );
and ( w_856 ,  , w_857 );
buf ( w_855 , \B[5]_b1 );
not ( w_855 , w_858 );
not (  , w_859 );
and ( w_858 , w_859 , \B[5]_b0 );
or ( \322_b1 , \320_b1 , \321_b1 );
xor ( \322_b0 , \320_b0 , w_860 );
not ( w_860 , w_861 );
and ( w_861 , \321_b1 , \321_b0 );
or ( \323_b1 , \153_b1 , w_863 );
not ( w_863 , w_864 );
and ( \323_b0 , \153_b0 , w_865 );
and ( w_864 ,  , w_865 );
buf ( w_863 , \B[6]_b1 );
not ( w_863 , w_866 );
not (  , w_867 );
and ( w_866 , w_867 , \B[6]_b0 );
or ( \324_b1 , \322_b1 , \323_b1 );
xor ( \324_b0 , \322_b0 , w_868 );
not ( w_868 , w_869 );
and ( w_869 , \323_b1 , \323_b0 );
or ( \325_b1 , \241_b1 , \242_b1 );
xor ( \325_b0 , \241_b0 , w_870 );
not ( w_870 , w_871 );
and ( w_871 , \242_b1 , \242_b0 );
or ( \326_b1 , \325_b1 , \244_b1 );
not ( \244_b1 , w_872 );
and ( \326_b0 , \325_b0 , w_873 );
and ( w_872 , w_873 , \244_b0 );
or ( \327_b1 , \241_b1 , \242_b1 );
not ( \242_b1 , w_874 );
and ( \327_b0 , \241_b0 , w_875 );
and ( w_874 , w_875 , \242_b0 );
or ( \328_b1 , \326_b1 , w_876 );
or ( \328_b0 , \326_b0 , \327_b0 );
not ( \327_b0 , w_877 );
and ( w_877 , w_876 , \327_b1 );
or ( \329_b1 , \324_b1 , \328_b1 );
not ( \328_b1 , w_878 );
and ( \329_b0 , \324_b0 , w_879 );
and ( w_878 , w_879 , \328_b0 );
buf ( \330_b1 , \324_b1 );
not ( \330_b1 , w_880 );
not ( \330_b0 , w_881 );
and ( w_880 , w_881 , \324_b0 );
buf ( \331_b1 , \328_b1 );
not ( \331_b1 , w_882 );
not ( \331_b0 , w_883 );
and ( w_882 , w_883 , \328_b0 );
or ( \332_b1 , \330_b1 , \331_b1 );
not ( \331_b1 , w_884 );
and ( \332_b0 , \330_b0 , w_885 );
and ( w_884 , w_885 , \331_b0 );
or ( \333_b1 , \329_b1 , w_887 );
not ( w_887 , w_888 );
and ( \333_b0 , \329_b0 , w_889 );
and ( w_888 ,  , w_889 );
buf ( w_887 , \332_b1 );
not ( w_887 , w_890 );
not (  , w_891 );
and ( w_890 , w_891 , \332_b0 );
or ( \334_b1 , \95_b1 , w_893 );
not ( w_893 , w_894 );
and ( \334_b0 , \95_b0 , w_895 );
and ( w_894 ,  , w_895 );
buf ( w_893 , \B[9]_b1 );
not ( w_893 , w_896 );
not (  , w_897 );
and ( w_896 , w_897 , \B[9]_b0 );
or ( \335_b1 , \86_b1 , w_899 );
not ( w_899 , w_900 );
and ( \335_b0 , \86_b0 , w_901 );
and ( w_900 ,  , w_901 );
buf ( w_899 , \B[7]_b1 );
not ( w_899 , w_902 );
not (  , w_903 );
and ( w_902 , w_903 , \B[7]_b0 );
or ( \336_b1 , \334_b1 , \335_b1 );
xor ( \336_b0 , \334_b0 , w_904 );
not ( w_904 , w_905 );
and ( w_905 , \335_b1 , \335_b0 );
or ( \337_b1 , \195_b1 , \196_b1 );
xor ( \337_b0 , \195_b0 , w_906 );
not ( w_906 , w_907 );
and ( w_907 , \196_b1 , \196_b0 );
or ( \338_b1 , \337_b1 , \198_b1 );
not ( \198_b1 , w_908 );
and ( \338_b0 , \337_b0 , w_909 );
and ( w_908 , w_909 , \198_b0 );
or ( \339_b1 , \195_b1 , \196_b1 );
not ( \196_b1 , w_910 );
and ( \339_b0 , \195_b0 , w_911 );
and ( w_910 , w_911 , \196_b0 );
or ( \340_b1 , \338_b1 , w_912 );
or ( \340_b0 , \338_b0 , \339_b0 );
not ( \339_b0 , w_913 );
and ( w_913 , w_912 , \339_b1 );
or ( \341_b1 , \336_b1 , \340_b1 );
xor ( \341_b0 , \336_b0 , w_914 );
not ( w_914 , w_915 );
and ( w_915 , \340_b1 , \340_b0 );
or ( \342_b1 , \333_b1 , \341_b1 );
not ( \341_b1 , w_916 );
and ( \342_b0 , \333_b0 , w_917 );
and ( w_916 , w_917 , \341_b0 );
buf ( \343_b1 , \333_b1 );
not ( \343_b1 , w_918 );
not ( \343_b0 , w_919 );
and ( w_918 , w_919 , \333_b0 );
buf ( \344_b1 , \341_b1 );
not ( \344_b1 , w_920 );
not ( \344_b0 , w_921 );
and ( w_920 , w_921 , \341_b0 );
or ( \345_b1 , \343_b1 , \344_b1 );
not ( \344_b1 , w_922 );
and ( \345_b0 , \343_b0 , w_923 );
and ( w_922 , w_923 , \344_b0 );
or ( \346_b1 , \342_b1 , w_924 );
or ( \346_b0 , \342_b0 , \345_b0 );
not ( \345_b0 , w_925 );
and ( w_925 , w_924 , \345_b1 );
or ( \347_b1 , \319_b1 , \346_b1 );
xor ( \347_b0 , \319_b0 , w_926 );
not ( w_926 , w_927 );
and ( w_927 , \346_b1 , \346_b0 );
buf ( \348_b1 , \199_b1 );
not ( \348_b1 , w_928 );
not ( \348_b0 , w_929 );
and ( w_928 , w_929 , \199_b0 );
buf ( \349_b1 , \251_b1 );
not ( \349_b1 , w_930 );
not ( \349_b0 , w_931 );
and ( w_930 , w_931 , \251_b0 );
buf ( \350_b1 , \349_b1 );
not ( \350_b1 , w_932 );
not ( \350_b0 , w_933 );
and ( w_932 , w_933 , \349_b0 );
or ( \351_b1 , \348_b1 , w_934 );
or ( \351_b0 , \348_b0 , \350_b0 );
not ( \350_b0 , w_935 );
and ( w_935 , w_934 , \350_b1 );
buf ( \352_b1 , \219_b1 );
not ( \352_b1 , w_936 );
not ( \352_b0 , w_937 );
and ( w_936 , w_937 , \219_b0 );
or ( \353_b1 , \351_b1 , w_939 );
not ( w_939 , w_940 );
and ( \353_b0 , \351_b0 , w_941 );
and ( w_940 ,  , w_941 );
buf ( w_939 , \352_b1 );
not ( w_939 , w_942 );
not (  , w_943 );
and ( w_942 , w_943 , \352_b0 );
buf ( \354_b1 , \199_b1 );
not ( \354_b1 , w_944 );
not ( \354_b0 , w_945 );
and ( w_944 , w_945 , \199_b0 );
or ( \355_b1 , \354_b1 , w_947 );
not ( w_947 , w_948 );
and ( \355_b0 , \354_b0 , w_949 );
and ( w_948 ,  , w_949 );
buf ( w_947 , \251_b1 );
not ( w_947 , w_950 );
not (  , w_951 );
and ( w_950 , w_951 , \251_b0 );
or ( \356_b1 , \353_b1 , w_953 );
not ( w_953 , w_954 );
and ( \356_b0 , \353_b0 , w_955 );
and ( w_954 ,  , w_955 );
buf ( w_953 , \355_b1 );
not ( w_953 , w_956 );
not (  , w_957 );
and ( w_956 , w_957 , \355_b0 );
or ( \357_b1 , \347_b1 , \356_b1 );
xor ( \357_b0 , \347_b0 , w_958 );
not ( w_958 , w_959 );
and ( w_959 , \356_b1 , \356_b0 );
or ( \358_b1 , \313_b1 , w_960 );
or ( \358_b0 , \313_b0 , \357_b0 );
not ( \357_b0 , w_961 );
and ( w_961 , w_960 , \357_b1 );
or ( \359_b1 , \334_b1 , \335_b1 );
xor ( \359_b0 , \334_b0 , w_962 );
not ( w_962 , w_963 );
and ( w_963 , \335_b1 , \335_b0 );
or ( \360_b1 , \359_b1 , \340_b1 );
not ( \340_b1 , w_964 );
and ( \360_b0 , \359_b0 , w_965 );
and ( w_964 , w_965 , \340_b0 );
or ( \361_b1 , \334_b1 , \335_b1 );
not ( \335_b1 , w_966 );
and ( \361_b0 , \334_b0 , w_967 );
and ( w_966 , w_967 , \335_b0 );
or ( \362_b1 , \360_b1 , w_968 );
or ( \362_b0 , \360_b0 , \361_b0 );
not ( \361_b0 , w_969 );
and ( w_969 , w_968 , \361_b1 );
or ( \363_b1 , \86_b1 , w_971 );
not ( w_971 , w_972 );
and ( \363_b0 , \86_b0 , w_973 );
and ( w_972 ,  , w_973 );
buf ( w_971 , \B[8]_b1 );
not ( w_971 , w_974 );
not (  , w_975 );
and ( w_974 , w_975 , \B[8]_b0 );
or ( \364_b1 , \320_b1 , \321_b1 );
xor ( \364_b0 , \320_b0 , w_976 );
not ( w_976 , w_977 );
and ( w_977 , \321_b1 , \321_b0 );
or ( \365_b1 , \364_b1 , \323_b1 );
not ( \323_b1 , w_978 );
and ( \365_b0 , \364_b0 , w_979 );
and ( w_978 , w_979 , \323_b0 );
or ( \366_b1 , \320_b1 , \321_b1 );
not ( \321_b1 , w_980 );
and ( \366_b0 , \320_b0 , w_981 );
and ( w_980 , w_981 , \321_b0 );
or ( \367_b1 , \365_b1 , w_982 );
or ( \367_b0 , \365_b0 , \366_b0 );
not ( \366_b0 , w_983 );
and ( w_983 , w_982 , \366_b1 );
or ( \368_b1 , \363_b1 , \367_b1 );
xor ( \368_b0 , \363_b0 , w_984 );
not ( w_984 , w_985 );
and ( w_985 , \367_b1 , \367_b0 );
or ( \369_b1 , \153_b1 , w_987 );
not ( w_987 , w_988 );
and ( \369_b0 , \153_b0 , w_989 );
and ( w_988 ,  , w_989 );
buf ( w_987 , \B[7]_b1 );
not ( w_987 , w_990 );
not (  , w_991 );
and ( w_990 , w_991 , \B[7]_b0 );
or ( \370_b1 , \79_b1 , w_993 );
not ( w_993 , w_994 );
and ( \370_b0 , \79_b0 , w_995 );
and ( w_994 ,  , w_995 );
buf ( w_993 , \B[6]_b1 );
not ( w_993 , w_996 );
not (  , w_997 );
and ( w_996 , w_997 , \B[6]_b0 );
or ( \371_b1 , \369_b1 , \370_b1 );
xor ( \371_b0 , \369_b0 , w_998 );
not ( w_998 , w_999 );
and ( w_999 , \370_b1 , \370_b0 );
or ( \372_b1 , \136_b1 , w_1001 );
not ( w_1001 , w_1002 );
and ( \372_b0 , \136_b0 , w_1003 );
and ( w_1002 ,  , w_1003 );
buf ( w_1001 , \B[9]_b1 );
not ( w_1001 , w_1004 );
not (  , w_1005 );
and ( w_1004 , w_1005 , \B[9]_b0 );
or ( \373_b1 , \371_b1 , \372_b1 );
xor ( \373_b0 , \371_b0 , w_1006 );
not ( w_1006 , w_1007 );
and ( w_1007 , \372_b1 , \372_b0 );
or ( \374_b1 , \368_b1 , \373_b1 );
xor ( \374_b0 , \368_b0 , w_1008 );
not ( w_1008 , w_1009 );
and ( w_1009 , \373_b1 , \373_b0 );
or ( \375_b1 , \362_b1 , \374_b1 );
xor ( \375_b0 , \362_b0 , w_1010 );
not ( w_1010 , w_1011 );
and ( w_1011 , \374_b1 , \374_b0 );
or ( \376_b1 , \341_b1 , w_1013 );
not ( w_1013 , w_1014 );
and ( \376_b0 , \341_b0 , w_1015 );
and ( w_1014 ,  , w_1015 );
buf ( w_1013 , \324_b1 );
not ( w_1013 , w_1016 );
not (  , w_1017 );
and ( w_1016 , w_1017 , \324_b0 );
or ( \377_b1 , \376_b1 , \331_b1 );
not ( \331_b1 , w_1018 );
and ( \377_b0 , \376_b0 , w_1019 );
and ( w_1018 , w_1019 , \331_b0 );
or ( \378_b1 , \341_b1 , w_1021 );
not ( w_1021 , w_1022 );
and ( \378_b0 , \341_b0 , w_1023 );
and ( w_1022 ,  , w_1023 );
buf ( w_1021 , \324_b1 );
not ( w_1021 , w_1024 );
not (  , w_1025 );
and ( w_1024 , w_1025 , \324_b0 );
or ( \379_b1 , \377_b1 , w_1027 );
not ( w_1027 , w_1028 );
and ( \379_b0 , \377_b0 , w_1029 );
and ( w_1028 ,  , w_1029 );
buf ( w_1027 , \378_b1 );
not ( w_1027 , w_1030 );
not (  , w_1031 );
and ( w_1030 , w_1031 , \378_b0 );
or ( \380_b1 , \375_b1 , \379_b1 );
xor ( \380_b0 , \375_b0 , w_1032 );
not ( w_1032 , w_1033 );
and ( w_1033 , \379_b1 , \379_b0 );
buf ( \381_b1 , \380_b1 );
not ( \381_b1 , w_1034 );
not ( \381_b0 , w_1035 );
and ( w_1034 , w_1035 , \380_b0 );
or ( \382_b1 , \319_b1 , \346_b1 );
xor ( \382_b0 , \319_b0 , w_1036 );
not ( w_1036 , w_1037 );
and ( w_1037 , \346_b1 , \346_b0 );
or ( \383_b1 , \382_b1 , \356_b1 );
not ( \356_b1 , w_1038 );
and ( \383_b0 , \382_b0 , w_1039 );
and ( w_1038 , w_1039 , \356_b0 );
or ( \384_b1 , \319_b1 , \346_b1 );
not ( \346_b1 , w_1040 );
and ( \384_b0 , \319_b0 , w_1041 );
and ( w_1040 , w_1041 , \346_b0 );
or ( \385_b1 , \383_b1 , w_1042 );
or ( \385_b0 , \383_b0 , \384_b0 );
not ( \384_b0 , w_1043 );
and ( w_1043 , w_1042 , \384_b1 );
or ( \386_b1 , \381_b1 , w_1045 );
not ( w_1045 , w_1046 );
and ( \386_b0 , \381_b0 , w_1047 );
and ( w_1046 ,  , w_1047 );
buf ( w_1045 , \385_b1 );
not ( w_1045 , w_1048 );
not (  , w_1049 );
and ( w_1048 , w_1049 , \385_b0 );
buf ( \387_b1 , \386_b1 );
not ( \387_b1 , w_1050 );
not ( \387_b0 , w_1051 );
and ( w_1050 , w_1051 , \386_b0 );
or ( \388_b1 , \358_b1 , w_1053 );
not ( w_1053 , w_1054 );
and ( \388_b0 , \358_b0 , w_1055 );
and ( w_1054 ,  , w_1055 );
buf ( w_1053 , \387_b1 );
not ( w_1053 , w_1056 );
not (  , w_1057 );
and ( w_1056 , w_1057 , \387_b0 );
or ( \389_b1 , \369_b1 , \370_b1 );
xor ( \389_b0 , \369_b0 , w_1058 );
not ( w_1058 , w_1059 );
and ( w_1059 , \370_b1 , \370_b0 );
or ( \390_b1 , \389_b1 , \372_b1 );
not ( \372_b1 , w_1060 );
and ( \390_b0 , \389_b0 , w_1061 );
and ( w_1060 , w_1061 , \372_b0 );
or ( \391_b1 , \369_b1 , \370_b1 );
not ( \370_b1 , w_1062 );
and ( \391_b0 , \369_b0 , w_1063 );
and ( w_1062 , w_1063 , \370_b0 );
or ( \392_b1 , \390_b1 , w_1064 );
or ( \392_b0 , \390_b0 , \391_b0 );
not ( \391_b0 , w_1065 );
and ( w_1065 , w_1064 , \391_b1 );
or ( \393_b1 , \156_b1 , \157_b1 );
xor ( \393_b0 , \156_b0 , w_1066 );
not ( w_1066 , w_1067 );
and ( w_1067 , \157_b1 , \157_b0 );
or ( \394_b1 , \393_b1 , \159_b1 );
xor ( \394_b0 , \393_b0 , w_1068 );
not ( w_1068 , w_1069 );
and ( w_1069 , \159_b1 , \159_b0 );
or ( \395_b1 , \392_b1 , \394_b1 );
xor ( \395_b0 , \392_b0 , w_1070 );
not ( w_1070 , w_1071 );
and ( w_1071 , \394_b1 , \394_b0 );
or ( \396_b1 , \363_b1 , \367_b1 );
xor ( \396_b0 , \363_b0 , w_1072 );
not ( w_1072 , w_1073 );
and ( w_1073 , \367_b1 , \367_b0 );
or ( \397_b1 , \396_b1 , \373_b1 );
not ( \373_b1 , w_1074 );
and ( \397_b0 , \396_b0 , w_1075 );
and ( w_1074 , w_1075 , \373_b0 );
or ( \398_b1 , \363_b1 , \367_b1 );
not ( \367_b1 , w_1076 );
and ( \398_b0 , \363_b0 , w_1077 );
and ( w_1076 , w_1077 , \367_b0 );
or ( \399_b1 , \397_b1 , w_1078 );
or ( \399_b0 , \397_b0 , \398_b0 );
not ( \398_b0 , w_1079 );
and ( w_1079 , w_1078 , \398_b1 );
or ( \400_b1 , \395_b1 , \399_b1 );
not ( \399_b1 , w_1080 );
and ( \400_b0 , \395_b0 , w_1081 );
and ( w_1080 , w_1081 , \399_b0 );
or ( \401_b1 , \392_b1 , \394_b1 );
not ( \394_b1 , w_1082 );
and ( \401_b0 , \392_b0 , w_1083 );
and ( w_1082 , w_1083 , \394_b0 );
or ( \402_b1 , \400_b1 , w_1084 );
or ( \402_b0 , \400_b0 , \401_b0 );
not ( \401_b0 , w_1085 );
and ( w_1085 , w_1084 , \401_b1 );
or ( \403_b1 , \147_b1 , \154_b1 );
xor ( \403_b0 , \147_b0 , w_1086 );
not ( w_1086 , w_1087 );
and ( w_1087 , \154_b1 , \154_b0 );
or ( \404_b1 , \403_b1 , \162_b1 );
xor ( \404_b0 , \403_b0 , w_1088 );
not ( w_1088 , w_1089 );
and ( w_1089 , \162_b1 , \162_b0 );
or ( \405_b1 , \402_b1 , w_1091 );
not ( w_1091 , w_1092 );
and ( \405_b0 , \402_b0 , w_1093 );
and ( w_1092 ,  , w_1093 );
buf ( w_1091 , \404_b1 );
not ( w_1091 , w_1094 );
not (  , w_1095 );
and ( w_1094 , w_1095 , \404_b0 );
or ( \406_b1 , \362_b1 , \374_b1 );
xor ( \406_b0 , \362_b0 , w_1096 );
not ( w_1096 , w_1097 );
and ( w_1097 , \374_b1 , \374_b0 );
or ( \407_b1 , \406_b1 , \379_b1 );
not ( \379_b1 , w_1098 );
and ( \407_b0 , \406_b0 , w_1099 );
and ( w_1098 , w_1099 , \379_b0 );
or ( \408_b1 , \362_b1 , \374_b1 );
not ( \374_b1 , w_1100 );
and ( \408_b0 , \362_b0 , w_1101 );
and ( w_1100 , w_1101 , \374_b0 );
or ( \409_b1 , \407_b1 , w_1102 );
or ( \409_b0 , \407_b0 , \408_b0 );
not ( \408_b0 , w_1103 );
and ( w_1103 , w_1102 , \408_b1 );
or ( \410_b1 , \392_b1 , \394_b1 );
xor ( \410_b0 , \392_b0 , w_1104 );
not ( w_1104 , w_1105 );
and ( w_1105 , \394_b1 , \394_b0 );
or ( \411_b1 , \410_b1 , \399_b1 );
xor ( \411_b0 , \410_b0 , w_1106 );
not ( w_1106 , w_1107 );
and ( w_1107 , \399_b1 , \399_b0 );
or ( \412_b1 , \409_b1 , w_1109 );
not ( w_1109 , w_1110 );
and ( \412_b0 , \409_b0 , w_1111 );
and ( w_1110 ,  , w_1111 );
buf ( w_1109 , \411_b1 );
not ( w_1109 , w_1112 );
not (  , w_1113 );
and ( w_1112 , w_1113 , \411_b0 );
or ( \413_b1 , \405_b1 , w_1115 );
not ( w_1115 , w_1116 );
and ( \413_b0 , \405_b0 , w_1117 );
and ( w_1116 ,  , w_1117 );
buf ( w_1115 , \412_b1 );
not ( w_1115 , w_1118 );
not (  , w_1119 );
and ( w_1118 , w_1119 , \412_b0 );
or ( \414_b1 , \388_b1 , w_1121 );
not ( w_1121 , w_1122 );
and ( \414_b0 , \388_b0 , w_1123 );
and ( w_1122 ,  , w_1123 );
buf ( w_1121 , \413_b1 );
not ( w_1121 , w_1124 );
not (  , w_1125 );
and ( w_1124 , w_1125 , \413_b0 );
buf ( \415_b1 , \414_b1 );
not ( \415_b1 , w_1126 );
not ( \415_b0 , w_1127 );
and ( w_1126 , w_1127 , \414_b0 );
or ( \416_b1 , \256_b1 , \287_b1 );
xor ( \416_b0 , \256_b0 , w_1128 );
not ( w_1128 , w_1129 );
and ( w_1129 , \287_b1 , \287_b0 );
or ( \417_b1 , \416_b1 , \306_b1 );
xor ( \417_b0 , \416_b0 , w_1130 );
not ( w_1130 , w_1131 );
and ( w_1131 , \306_b1 , \306_b0 );
or ( \418_b1 , \190_b1 , \191_b1 );
xor ( \418_b0 , \190_b0 , w_1132 );
not ( w_1132 , w_1133 );
and ( w_1133 , \191_b1 , \191_b0 );
or ( \419_b1 , \418_b1 , \188_b1 );
not ( \188_b1 , w_1134 );
and ( \419_b0 , \418_b0 , w_1135 );
and ( w_1134 , w_1135 , \188_b0 );
buf ( \420_b1 , \418_b1 );
not ( \420_b1 , w_1136 );
not ( \420_b0 , w_1137 );
and ( w_1136 , w_1137 , \418_b0 );
buf ( \421_b1 , \188_b1 );
not ( \421_b1 , w_1138 );
not ( \421_b0 , w_1139 );
and ( w_1138 , w_1139 , \188_b0 );
or ( \422_b1 , \420_b1 , \421_b1 );
not ( \421_b1 , w_1140 );
and ( \422_b0 , \420_b0 , w_1141 );
and ( w_1140 , w_1141 , \421_b0 );
or ( \423_b1 , \419_b1 , w_1142 );
or ( \423_b0 , \419_b0 , \422_b0 );
not ( \422_b0 , w_1143 );
and ( w_1143 , w_1142 , \422_b1 );
or ( \424_b1 , \417_b1 , \423_b1 );
xor ( \424_b0 , \417_b0 , w_1144 );
not ( w_1144 , w_1145 );
and ( w_1145 , \423_b1 , \423_b0 );
buf ( \425_b1 , \285_b1 );
not ( \425_b1 , w_1146 );
not ( \425_b0 , w_1147 );
and ( w_1146 , w_1147 , \285_b0 );
buf ( \426_b1 , \272_b1 );
not ( \426_b1 , w_1148 );
not ( \426_b0 , w_1149 );
and ( w_1148 , w_1149 , \272_b0 );
or ( \427_b1 , \425_b1 , w_1150 );
or ( \427_b0 , \425_b0 , \426_b0 );
not ( \426_b0 , w_1151 );
and ( w_1151 , w_1150 , \426_b1 );
buf ( \428_b1 , \285_b1 );
not ( \428_b1 , w_1152 );
not ( \428_b0 , w_1153 );
and ( w_1152 , w_1153 , \285_b0 );
or ( \429_b1 , \428_b1 , w_1155 );
not ( w_1155 , w_1156 );
and ( \429_b0 , \428_b0 , w_1157 );
and ( w_1156 ,  , w_1157 );
buf ( w_1155 , \270_b1 );
not ( w_1155 , w_1158 );
not (  , w_1159 );
and ( w_1158 , w_1159 , \270_b0 );
or ( \430_b1 , \427_b1 , w_1161 );
not ( w_1161 , w_1162 );
and ( \430_b0 , \427_b0 , w_1163 );
and ( w_1162 ,  , w_1163 );
buf ( w_1161 , \429_b1 );
not ( w_1161 , w_1164 );
not (  , w_1165 );
and ( w_1164 , w_1165 , \429_b0 );
or ( \431_b1 , \430_b1 , \258_b1 );
not ( \258_b1 , w_1166 );
and ( \431_b0 , \430_b0 , w_1167 );
and ( w_1166 , w_1167 , \258_b0 );
buf ( \432_b1 , \430_b1 );
not ( \432_b1 , w_1168 );
not ( \432_b0 , w_1169 );
and ( w_1168 , w_1169 , \430_b0 );
buf ( \433_b1 , \258_b1 );
not ( \433_b1 , w_1170 );
not ( \433_b0 , w_1171 );
and ( w_1170 , w_1171 , \258_b0 );
or ( \434_b1 , \432_b1 , \433_b1 );
not ( \433_b1 , w_1172 );
and ( \434_b0 , \432_b0 , w_1173 );
and ( w_1172 , w_1173 , \433_b0 );
or ( \435_b1 , \431_b1 , w_1175 );
not ( w_1175 , w_1176 );
and ( \435_b0 , \431_b0 , w_1177 );
and ( w_1176 ,  , w_1177 );
buf ( w_1175 , \434_b1 );
not ( w_1175 , w_1178 );
not (  , w_1179 );
and ( w_1178 , w_1179 , \434_b0 );
or ( \436_b1 , \95_b1 , w_1181 );
not ( w_1181 , w_1182 );
and ( \436_b0 , \95_b0 , w_1183 );
and ( w_1182 ,  , w_1183 );
buf ( w_1181 , \B[4]_b1 );
not ( w_1181 , w_1184 );
not (  , w_1185 );
and ( w_1184 , w_1185 , \B[4]_b0 );
or ( \437_b1 , \86_b1 , w_1187 );
not ( w_1187 , w_1188 );
and ( \437_b0 , \86_b0 , w_1189 );
and ( w_1188 ,  , w_1189 );
buf ( w_1187 , \B[2]_b1 );
not ( w_1187 , w_1190 );
not (  , w_1191 );
and ( w_1190 , w_1191 , \B[2]_b0 );
or ( \438_b1 , \436_b1 , \437_b1 );
xor ( \438_b0 , \436_b0 , w_1192 );
not ( w_1192 , w_1193 );
and ( w_1193 , \437_b1 , \437_b0 );
or ( \439_b1 , \B[9]_b1 , w_1195 );
not ( w_1195 , w_1196 );
and ( \439_b0 , \B[9]_b0 , w_1197 );
and ( w_1196 ,  , w_1197 );
buf ( w_1195 , \118_b1 );
not ( w_1195 , w_1198 );
not (  , w_1199 );
and ( w_1198 , w_1199 , \118_b0 );
or ( \440_b1 , \438_b1 , \439_b1 );
not ( \439_b1 , w_1200 );
and ( \440_b0 , \438_b0 , w_1201 );
and ( w_1200 , w_1201 , \439_b0 );
or ( \441_b1 , \436_b1 , \437_b1 );
not ( \437_b1 , w_1202 );
and ( \441_b0 , \436_b0 , w_1203 );
and ( w_1202 , w_1203 , \437_b0 );
or ( \442_b1 , \440_b1 , w_1204 );
or ( \442_b0 , \440_b0 , \441_b0 );
not ( \441_b0 , w_1205 );
and ( w_1205 , w_1204 , \441_b1 );
or ( \443_b1 , \276_b1 , \281_b1 );
xor ( \443_b0 , \276_b0 , w_1206 );
not ( w_1206 , w_1207 );
and ( w_1207 , \281_b1 , \281_b0 );
or ( \444_b1 , \443_b1 , \278_b1 );
xor ( \444_b0 , \443_b0 , w_1208 );
not ( w_1208 , w_1209 );
and ( w_1209 , \278_b1 , \278_b0 );
or ( \445_b1 , \442_b1 , \444_b1 );
xor ( \445_b0 , \442_b0 , w_1210 );
not ( w_1210 , w_1211 );
and ( w_1211 , \444_b1 , \444_b0 );
or ( \446_b1 , \136_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_1212 );
and ( \446_b0 , \136_b0 , w_1213 );
and ( w_1212 , w_1213 , \B[3]_b0 );
or ( \447_b1 , \104_b1 , \B[7]_b1 );
not ( \B[7]_b1 , w_1214 );
and ( \447_b0 , \104_b0 , w_1215 );
and ( w_1214 , w_1215 , \B[7]_b0 );
or ( \448_b1 , \446_b1 , w_1216 );
or ( \448_b0 , \446_b0 , \447_b0 );
not ( \447_b0 , w_1217 );
and ( w_1217 , w_1216 , \447_b1 );
or ( \449_b1 , \111_b1 , w_1219 );
not ( w_1219 , w_1220 );
and ( \449_b0 , \111_b0 , w_1221 );
and ( w_1220 ,  , w_1221 );
buf ( w_1219 , \B[8]_b1 );
not ( w_1219 , w_1222 );
not (  , w_1223 );
and ( w_1222 , w_1223 , \B[8]_b0 );
buf ( \450_b1 , \449_b1 );
not ( \450_b1 , w_1224 );
not ( \450_b0 , w_1225 );
and ( w_1224 , w_1225 , \449_b0 );
or ( \451_b1 , \448_b1 , \450_b1 );
not ( \450_b1 , w_1226 );
and ( \451_b0 , \448_b0 , w_1227 );
and ( w_1226 , w_1227 , \450_b0 );
or ( \452_b1 , \446_b1 , \447_b1 );
not ( \447_b1 , w_1228 );
and ( \452_b0 , \446_b0 , w_1229 );
and ( w_1228 , w_1229 , \447_b0 );
or ( \453_b1 , \451_b1 , w_1231 );
not ( w_1231 , w_1232 );
and ( \453_b0 , \451_b0 , w_1233 );
and ( w_1232 ,  , w_1233 );
buf ( w_1231 , \452_b1 );
not ( w_1231 , w_1234 );
not (  , w_1235 );
and ( w_1234 , w_1235 , \452_b0 );
or ( \454_b1 , \445_b1 , \453_b1 );
not ( \453_b1 , w_1236 );
and ( \454_b0 , \445_b0 , w_1237 );
and ( w_1236 , w_1237 , \453_b0 );
or ( \455_b1 , \442_b1 , \444_b1 );
not ( \444_b1 , w_1238 );
and ( \455_b0 , \442_b0 , w_1239 );
and ( w_1238 , w_1239 , \444_b0 );
or ( \456_b1 , \454_b1 , w_1240 );
or ( \456_b0 , \454_b0 , \455_b0 );
not ( \455_b0 , w_1241 );
and ( w_1241 , w_1240 , \455_b1 );
or ( \457_b1 , \435_b1 , \456_b1 );
xor ( \457_b0 , \435_b0 , w_1242 );
not ( w_1242 , w_1243 );
and ( w_1243 , \456_b1 , \456_b0 );
or ( \458_b1 , \260_b1 , \268_b1 );
xor ( \458_b0 , \260_b0 , w_1244 );
not ( w_1244 , w_1245 );
and ( w_1245 , \268_b1 , \268_b0 );
or ( \459_b1 , \458_b1 , \265_b1 );
xor ( \459_b0 , \458_b0 , w_1246 );
not ( w_1246 , w_1247 );
and ( w_1247 , \265_b1 , \265_b0 );
or ( \460_b1 , \200_b1 , w_1249 );
not ( w_1249 , w_1250 );
and ( \460_b0 , \200_b0 , w_1251 );
and ( w_1250 ,  , w_1251 );
buf ( w_1249 , \B[6]_b1 );
not ( w_1249 , w_1252 );
not (  , w_1253 );
and ( w_1252 , w_1253 , \B[6]_b0 );
or ( \461_b1 , \127_b1 , w_1255 );
not ( w_1255 , w_1256 );
and ( \461_b0 , \127_b0 , w_1257 );
and ( w_1256 ,  , w_1257 );
buf ( w_1255 , \B[5]_b1 );
not ( w_1255 , w_1258 );
not (  , w_1259 );
and ( w_1258 , w_1259 , \B[5]_b0 );
or ( \462_b1 , \460_b1 , \461_b1 );
xor ( \462_b0 , \460_b0 , w_1260 );
not ( w_1260 , w_1261 );
and ( w_1261 , \461_b1 , \461_b0 );
buf ( \463_b1 , \297_b1 );
not ( \463_b1 , w_1262 );
not ( \463_b0 , w_1263 );
and ( w_1262 , w_1263 , \297_b0 );
buf ( \464_b1 , \295_b1 );
not ( \464_b1 , w_1264 );
not ( \464_b0 , w_1265 );
and ( w_1264 , w_1265 , \295_b0 );
or ( \465_b1 , \463_b1 , \464_b1 );
not ( \464_b1 , w_1266 );
and ( \465_b0 , \463_b0 , w_1267 );
and ( w_1266 , w_1267 , \464_b0 );
or ( \466_b1 , \297_b1 , \295_b1 );
not ( \295_b1 , w_1268 );
and ( \466_b0 , \297_b0 , w_1269 );
and ( w_1268 , w_1269 , \295_b0 );
or ( \467_b1 , \465_b1 , w_1271 );
not ( w_1271 , w_1272 );
and ( \467_b0 , \465_b0 , w_1273 );
and ( w_1272 ,  , w_1273 );
buf ( w_1271 , \466_b1 );
not ( w_1271 , w_1274 );
not (  , w_1275 );
and ( w_1274 , w_1275 , \466_b0 );
or ( \468_b1 , \462_b1 , \467_b1 );
not ( \467_b1 , w_1276 );
and ( \468_b0 , \462_b0 , w_1277 );
and ( w_1276 , w_1277 , \467_b0 );
or ( \469_b1 , \460_b1 , \461_b1 );
not ( \461_b1 , w_1278 );
and ( \469_b0 , \460_b0 , w_1279 );
and ( w_1278 , w_1279 , \461_b0 );
or ( \470_b1 , \468_b1 , w_1280 );
or ( \470_b0 , \468_b0 , \469_b0 );
not ( \469_b0 , w_1281 );
and ( w_1281 , w_1280 , \469_b1 );
or ( \471_b1 , \459_b1 , \470_b1 );
xor ( \471_b0 , \459_b0 , w_1282 );
not ( w_1282 , w_1283 );
and ( w_1283 , \470_b1 , \470_b0 );
or ( \472_b1 , \86_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_1284 );
and ( \472_b0 , \86_b0 , w_1285 );
and ( w_1284 , w_1285 , \B[0]_b0 );
or ( \473_b1 , \297_b1 , w_1287 );
not ( w_1287 , w_1288 );
and ( \473_b0 , \297_b0 , w_1289 );
and ( w_1288 ,  , w_1289 );
buf ( w_1287 , \472_b1 );
not ( w_1287 , w_1290 );
not (  , w_1291 );
and ( w_1290 , w_1291 , \472_b0 );
or ( \474_b1 , \143_b1 , w_1293 );
not ( w_1293 , w_1294 );
and ( \474_b0 , \143_b0 , w_1295 );
and ( w_1294 ,  , w_1295 );
buf ( w_1293 , \B[5]_b1 );
not ( w_1293 , w_1296 );
not (  , w_1297 );
and ( w_1296 , w_1297 , \B[5]_b0 );
buf ( \475_b1 , \474_b1 );
not ( \475_b1 , w_1298 );
not ( \475_b0 , w_1299 );
and ( w_1298 , w_1299 , \474_b0 );
or ( \476_b1 , \127_b1 , w_1301 );
not ( w_1301 , w_1302 );
and ( \476_b0 , \127_b0 , w_1303 );
and ( w_1302 ,  , w_1303 );
buf ( w_1301 , \B[4]_b1 );
not ( w_1301 , w_1304 );
not (  , w_1305 );
and ( w_1304 , w_1305 , \B[4]_b0 );
buf ( \477_b1 , \476_b1 );
not ( \477_b1 , w_1306 );
not ( \477_b0 , w_1307 );
and ( w_1306 , w_1307 , \476_b0 );
or ( \478_b1 , \475_b1 , w_1308 );
or ( \478_b0 , \475_b0 , \477_b0 );
not ( \477_b0 , w_1309 );
and ( w_1309 , w_1308 , \477_b1 );
or ( \479_b1 , \136_b1 , \B[2]_b1 );
not ( \B[2]_b1 , w_1310 );
and ( \479_b0 , \136_b0 , w_1311 );
and ( w_1310 , w_1311 , \B[2]_b0 );
or ( \480_b1 , \478_b1 , w_1313 );
not ( w_1313 , w_1314 );
and ( \480_b0 , \478_b0 , w_1315 );
and ( w_1314 ,  , w_1315 );
buf ( w_1313 , \479_b1 );
not ( w_1313 , w_1316 );
not (  , w_1317 );
and ( w_1316 , w_1317 , \479_b0 );
buf ( \481_b1 , \476_b1 );
not ( \481_b1 , w_1318 );
not ( \481_b0 , w_1319 );
and ( w_1318 , w_1319 , \476_b0 );
buf ( \482_b1 , \474_b1 );
not ( \482_b1 , w_1320 );
not ( \482_b0 , w_1321 );
and ( w_1320 , w_1321 , \474_b0 );
or ( \483_b1 , \481_b1 , w_1323 );
not ( w_1323 , w_1324 );
and ( \483_b0 , \481_b0 , w_1325 );
and ( w_1324 ,  , w_1325 );
buf ( w_1323 , \482_b1 );
not ( w_1323 , w_1326 );
not (  , w_1327 );
and ( w_1326 , w_1327 , \482_b0 );
or ( \484_b1 , \480_b1 , w_1329 );
not ( w_1329 , w_1330 );
and ( \484_b0 , \480_b0 , w_1331 );
and ( w_1330 ,  , w_1331 );
buf ( w_1329 , \483_b1 );
not ( w_1329 , w_1332 );
not (  , w_1333 );
and ( w_1332 , w_1333 , \483_b0 );
buf ( \485_b1 , \484_b1 );
not ( \485_b1 , w_1334 );
not ( \485_b0 , w_1335 );
and ( w_1334 , w_1335 , \484_b0 );
or ( \486_b1 , \473_b1 , \485_b1 );
xor ( \486_b0 , \473_b0 , w_1336 );
not ( w_1336 , w_1337 );
and ( w_1337 , \485_b1 , \485_b0 );
or ( \487_b1 , \111_b1 , w_1339 );
not ( w_1339 , w_1340 );
and ( \487_b0 , \111_b0 , w_1341 );
and ( w_1340 ,  , w_1341 );
buf ( w_1339 , \B[7]_b1 );
not ( w_1339 , w_1342 );
not (  , w_1343 );
and ( w_1342 , w_1343 , \B[7]_b0 );
or ( \488_b1 , \95_b1 , w_1345 );
not ( w_1345 , w_1346 );
and ( \488_b0 , \95_b0 , w_1347 );
and ( w_1346 ,  , w_1347 );
buf ( w_1345 , \B[3]_b1 );
not ( w_1345 , w_1348 );
not (  , w_1349 );
and ( w_1348 , w_1349 , \B[3]_b0 );
or ( \489_b1 , \487_b1 , w_1351 );
not ( w_1351 , w_1352 );
and ( \489_b0 , \487_b0 , w_1353 );
and ( w_1352 ,  , w_1353 );
buf ( w_1351 , \488_b1 );
not ( w_1351 , w_1354 );
not (  , w_1355 );
and ( w_1354 , w_1355 , \488_b0 );
or ( \490_b1 , \118_b1 , \B[8]_b1 );
not ( \B[8]_b1 , w_1356 );
and ( \490_b0 , \118_b0 , w_1357 );
and ( w_1356 , w_1357 , \B[8]_b0 );
or ( \491_b1 , \489_b1 , \490_b1 );
not ( \490_b1 , w_1358 );
and ( \491_b0 , \489_b0 , w_1359 );
and ( w_1358 , w_1359 , \490_b0 );
or ( \492_b1 , \487_b1 , w_1361 );
not ( w_1361 , w_1362 );
and ( \492_b0 , \487_b0 , w_1363 );
and ( w_1362 ,  , w_1363 );
buf ( w_1361 , \488_b1 );
not ( w_1361 , w_1364 );
not (  , w_1365 );
and ( w_1364 , w_1365 , \488_b0 );
or ( \493_b1 , \491_b1 , w_1367 );
not ( w_1367 , w_1368 );
and ( \493_b0 , \491_b0 , w_1369 );
and ( w_1368 ,  , w_1369 );
buf ( w_1367 , \492_b1 );
not ( w_1367 , w_1370 );
not (  , w_1371 );
and ( w_1370 , w_1371 , \492_b0 );
or ( \494_b1 , \486_b1 , \493_b1 );
not ( \493_b1 , w_1372 );
and ( \494_b0 , \486_b0 , w_1373 );
and ( w_1372 , w_1373 , \493_b0 );
or ( \495_b1 , \473_b1 , \485_b1 );
not ( \485_b1 , w_1374 );
and ( \495_b0 , \473_b0 , w_1375 );
and ( w_1374 , w_1375 , \485_b0 );
or ( \496_b1 , \494_b1 , w_1376 );
or ( \496_b0 , \494_b0 , \495_b0 );
not ( \495_b0 , w_1377 );
and ( w_1377 , w_1376 , \495_b1 );
or ( \497_b1 , \471_b1 , \496_b1 );
not ( \496_b1 , w_1378 );
and ( \497_b0 , \471_b0 , w_1379 );
and ( w_1378 , w_1379 , \496_b0 );
or ( \498_b1 , \459_b1 , \470_b1 );
not ( \470_b1 , w_1380 );
and ( \498_b0 , \459_b0 , w_1381 );
and ( w_1380 , w_1381 , \470_b0 );
or ( \499_b1 , \497_b1 , w_1382 );
or ( \499_b0 , \497_b0 , \498_b0 );
not ( \498_b0 , w_1383 );
and ( w_1383 , w_1382 , \498_b1 );
or ( \500_b1 , \457_b1 , \499_b1 );
not ( \499_b1 , w_1384 );
and ( \500_b0 , \457_b0 , w_1385 );
and ( w_1384 , w_1385 , \499_b0 );
or ( \501_b1 , \435_b1 , \456_b1 );
not ( \456_b1 , w_1386 );
and ( \501_b0 , \435_b0 , w_1387 );
and ( w_1386 , w_1387 , \456_b0 );
or ( \502_b1 , \500_b1 , w_1388 );
or ( \502_b0 , \500_b0 , \501_b0 );
not ( \501_b0 , w_1389 );
and ( w_1389 , w_1388 , \501_b1 );
or ( \503_b1 , \424_b1 , w_1390 );
xor ( \503_b0 , \424_b0 , w_1392 );
not ( w_1392 , w_1393 );
and ( w_1393 , w_1390 , w_1391 );
buf ( w_1390 , \502_b1 );
not ( w_1390 , w_1394 );
not ( w_1391 , w_1395 );
and ( w_1394 , w_1395 , \502_b0 );
or ( \504_b1 , \290_b1 , \292_b1 );
xor ( \504_b0 , \290_b0 , w_1396 );
not ( w_1396 , w_1397 );
and ( w_1397 , \292_b1 , \292_b0 );
or ( \505_b1 , \504_b1 , \303_b1 );
xor ( \505_b0 , \504_b0 , w_1398 );
not ( w_1398 , w_1399 );
and ( w_1399 , \303_b1 , \303_b0 );
or ( \506_b1 , \294_b1 , \298_b1 );
xor ( \506_b0 , \294_b0 , w_1400 );
not ( w_1400 , w_1401 );
and ( w_1401 , \298_b1 , \298_b0 );
or ( \507_b1 , \506_b1 , \300_b1 );
xor ( \507_b0 , \506_b0 , w_1402 );
not ( w_1402 , w_1403 );
and ( w_1403 , \300_b1 , \300_b0 );
or ( \508_b1 , \442_b1 , \444_b1 );
xor ( \508_b0 , \442_b0 , w_1404 );
not ( w_1404 , w_1405 );
and ( w_1405 , \444_b1 , \444_b0 );
or ( \509_b1 , \508_b1 , \453_b1 );
xor ( \509_b0 , \508_b0 , w_1406 );
not ( w_1406 , w_1407 );
and ( w_1407 , \453_b1 , \453_b0 );
or ( \510_b1 , \507_b1 , \509_b1 );
xor ( \510_b0 , \507_b0 , w_1408 );
not ( w_1408 , w_1409 );
and ( w_1409 , \509_b1 , \509_b0 );
or ( \511_b1 , \446_b1 , \447_b1 );
xor ( \511_b0 , \446_b0 , w_1410 );
not ( w_1410 , w_1411 );
and ( w_1411 , \447_b1 , \447_b0 );
or ( \512_b1 , \511_b1 , \450_b1 );
not ( \450_b1 , w_1412 );
and ( \512_b0 , \511_b0 , w_1413 );
and ( w_1412 , w_1413 , \450_b0 );
buf ( \513_b1 , \511_b1 );
not ( \513_b1 , w_1414 );
not ( \513_b0 , w_1415 );
and ( w_1414 , w_1415 , \511_b0 );
or ( \514_b1 , \513_b1 , \449_b1 );
not ( \449_b1 , w_1416 );
and ( \514_b0 , \513_b0 , w_1417 );
and ( w_1416 , w_1417 , \449_b0 );
or ( \515_b1 , \512_b1 , w_1419 );
not ( w_1419 , w_1420 );
and ( \515_b0 , \512_b0 , w_1421 );
and ( w_1420 ,  , w_1421 );
buf ( w_1419 , \514_b1 );
not ( w_1419 , w_1422 );
not (  , w_1423 );
and ( w_1422 , w_1423 , \514_b0 );
buf ( \516_b1 , \515_b1 );
not ( \516_b1 , w_1424 );
not ( \516_b0 , w_1425 );
and ( w_1424 , w_1425 , \515_b0 );
or ( \517_b1 , \436_b1 , \437_b1 );
xor ( \517_b0 , \436_b0 , w_1426 );
not ( w_1426 , w_1427 );
and ( w_1427 , \437_b1 , \437_b0 );
or ( \518_b1 , \517_b1 , \439_b1 );
xor ( \518_b0 , \517_b0 , w_1428 );
not ( w_1428 , w_1429 );
and ( w_1429 , \439_b1 , \439_b0 );
or ( \519_b1 , \516_b1 , w_1431 );
not ( w_1431 , w_1432 );
and ( \519_b0 , \516_b0 , w_1433 );
and ( w_1432 ,  , w_1433 );
buf ( w_1431 , \518_b1 );
not ( w_1431 , w_1434 );
not (  , w_1435 );
and ( w_1434 , w_1435 , \518_b0 );
or ( \520_b1 , \104_b1 , \B[6]_b1 );
not ( \B[6]_b1 , w_1436 );
and ( \520_b0 , \104_b0 , w_1437 );
and ( w_1436 , w_1437 , \B[6]_b0 );
or ( \521_b1 , \86_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1438 );
and ( \521_b0 , \86_b0 , w_1439 );
and ( w_1438 , w_1439 , \B[1]_b0 );
buf ( \522_b1 , \521_b1 );
not ( \522_b1 , w_1440 );
not ( \522_b0 , w_1441 );
and ( w_1440 , w_1441 , \521_b0 );
or ( \523_b1 , \153_b1 , w_1443 );
not ( w_1443 , w_1444 );
and ( \523_b0 , \153_b0 , w_1445 );
and ( w_1444 ,  , w_1445 );
buf ( w_1443 , \B[0]_b1 );
not ( w_1443 , w_1446 );
not (  , w_1447 );
and ( w_1446 , w_1447 , \B[0]_b0 );
buf ( \524_b1 , \523_b1 );
not ( \524_b1 , w_1448 );
not ( \524_b0 , w_1449 );
and ( w_1448 , w_1449 , \523_b0 );
or ( \525_b1 , \522_b1 , w_1450 );
or ( \525_b0 , \522_b0 , \524_b0 );
not ( \524_b0 , w_1451 );
and ( w_1451 , w_1450 , \524_b1 );
or ( \526_b1 , \521_b1 , w_1452 );
or ( \526_b0 , \521_b0 , \523_b0 );
not ( \523_b0 , w_1453 );
and ( w_1453 , w_1452 , \523_b1 );
or ( \527_b1 , \525_b1 , w_1455 );
not ( w_1455 , w_1456 );
and ( \527_b0 , \525_b0 , w_1457 );
and ( w_1456 ,  , w_1457 );
buf ( w_1455 , \526_b1 );
not ( w_1455 , w_1458 );
not (  , w_1459 );
and ( w_1458 , w_1459 , \526_b0 );
or ( \528_b1 , \520_b1 , \527_b1 );
xor ( \528_b0 , \520_b0 , w_1460 );
not ( w_1460 , w_1461 );
and ( w_1461 , \527_b1 , \527_b0 );
or ( \529_b1 , \136_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1462 );
and ( \529_b0 , \136_b0 , w_1463 );
and ( w_1462 , w_1463 , \B[1]_b0 );
or ( \530_b1 , \472_b1 , \529_b1 );
not ( \529_b1 , w_1464 );
and ( \530_b0 , \472_b0 , w_1465 );
and ( w_1464 , w_1465 , \529_b0 );
or ( \531_b1 , \528_b1 , \530_b1 );
not ( \530_b1 , w_1466 );
and ( \531_b0 , \528_b0 , w_1467 );
and ( w_1466 , w_1467 , \530_b0 );
or ( \532_b1 , \520_b1 , \527_b1 );
not ( \527_b1 , w_1468 );
and ( \532_b0 , \520_b0 , w_1469 );
and ( w_1468 , w_1469 , \527_b0 );
or ( \533_b1 , \531_b1 , w_1470 );
or ( \533_b0 , \531_b0 , \532_b0 );
not ( \532_b0 , w_1471 );
and ( w_1471 , w_1470 , \532_b1 );
or ( \534_b1 , \519_b1 , \533_b1 );
not ( \533_b1 , w_1472 );
and ( \534_b0 , \519_b0 , w_1473 );
and ( w_1472 , w_1473 , \533_b0 );
or ( \535_b1 , \516_b1 , w_1475 );
not ( w_1475 , w_1476 );
and ( \535_b0 , \516_b0 , w_1477 );
and ( w_1476 ,  , w_1477 );
buf ( w_1475 , \518_b1 );
not ( w_1475 , w_1478 );
not (  , w_1479 );
and ( w_1478 , w_1479 , \518_b0 );
or ( \536_b1 , \534_b1 , w_1481 );
not ( w_1481 , w_1482 );
and ( \536_b0 , \534_b0 , w_1483 );
and ( w_1482 ,  , w_1483 );
buf ( w_1481 , \535_b1 );
not ( w_1481 , w_1484 );
not (  , w_1485 );
and ( w_1484 , w_1485 , \535_b0 );
or ( \537_b1 , \510_b1 , \536_b1 );
not ( \536_b1 , w_1486 );
and ( \537_b0 , \510_b0 , w_1487 );
and ( w_1486 , w_1487 , \536_b0 );
or ( \538_b1 , \507_b1 , \509_b1 );
not ( \509_b1 , w_1488 );
and ( \538_b0 , \507_b0 , w_1489 );
and ( w_1488 , w_1489 , \509_b0 );
or ( \539_b1 , \537_b1 , w_1490 );
or ( \539_b0 , \537_b0 , \538_b0 );
not ( \538_b0 , w_1491 );
and ( w_1491 , w_1490 , \538_b1 );
or ( \540_b1 , \505_b1 , \539_b1 );
xor ( \540_b0 , \505_b0 , w_1492 );
not ( w_1492 , w_1493 );
and ( w_1493 , \539_b1 , \539_b0 );
or ( \541_b1 , \435_b1 , \456_b1 );
xor ( \541_b0 , \435_b0 , w_1494 );
not ( w_1494 , w_1495 );
and ( w_1495 , \456_b1 , \456_b0 );
or ( \542_b1 , \541_b1 , \499_b1 );
xor ( \542_b0 , \541_b0 , w_1496 );
not ( w_1496 , w_1497 );
and ( w_1497 , \499_b1 , \499_b0 );
or ( \543_b1 , \540_b1 , \542_b1 );
not ( \542_b1 , w_1498 );
and ( \543_b0 , \540_b0 , w_1499 );
and ( w_1498 , w_1499 , \542_b0 );
or ( \544_b1 , \505_b1 , \539_b1 );
not ( \539_b1 , w_1500 );
and ( \544_b0 , \505_b0 , w_1501 );
and ( w_1500 , w_1501 , \539_b0 );
or ( \545_b1 , \543_b1 , w_1502 );
or ( \545_b0 , \543_b0 , \544_b0 );
not ( \544_b0 , w_1503 );
and ( w_1503 , w_1502 , \544_b1 );
or ( \546_b1 , \503_b1 , w_1505 );
not ( w_1505 , w_1506 );
and ( \546_b0 , \503_b0 , w_1507 );
and ( w_1506 ,  , w_1507 );
buf ( w_1505 , \545_b1 );
not ( w_1505 , w_1508 );
not (  , w_1509 );
and ( w_1508 , w_1509 , \545_b0 );
buf ( \547_b1 , \417_b1 );
not ( \547_b1 , w_1510 );
not ( \547_b0 , w_1511 );
and ( w_1510 , w_1511 , \417_b0 );
buf ( \548_b1 , \423_b1 );
not ( \548_b1 , w_1512 );
not ( \548_b0 , w_1513 );
and ( w_1512 , w_1513 , \423_b0 );
buf ( \549_b1 , \548_b1 );
not ( \549_b1 , w_1514 );
not ( \549_b0 , w_1515 );
and ( w_1514 , w_1515 , \548_b0 );
or ( \550_b1 , \547_b1 , w_1516 );
or ( \550_b0 , \547_b0 , \549_b0 );
not ( \549_b0 , w_1517 );
and ( w_1517 , w_1516 , \549_b1 );
buf ( \551_b1 , \502_b1 );
not ( \551_b1 , w_1518 );
not ( \551_b0 , w_1519 );
and ( w_1518 , w_1519 , \502_b0 );
or ( \552_b1 , \550_b1 , w_1521 );
not ( w_1521 , w_1522 );
and ( \552_b0 , \550_b0 , w_1523 );
and ( w_1522 ,  , w_1523 );
buf ( w_1521 , \551_b1 );
not ( w_1521 , w_1524 );
not (  , w_1525 );
and ( w_1524 , w_1525 , \551_b0 );
buf ( \553_b1 , \417_b1 );
not ( \553_b1 , w_1526 );
not ( \553_b0 , w_1527 );
and ( w_1526 , w_1527 , \417_b0 );
or ( \554_b1 , \553_b1 , w_1529 );
not ( w_1529 , w_1530 );
and ( \554_b0 , \553_b0 , w_1531 );
and ( w_1530 ,  , w_1531 );
buf ( w_1529 , \423_b1 );
not ( w_1529 , w_1532 );
not (  , w_1533 );
and ( w_1532 , w_1533 , \423_b0 );
or ( \555_b1 , \552_b1 , w_1535 );
not ( w_1535 , w_1536 );
and ( \555_b0 , \552_b0 , w_1537 );
and ( w_1536 ,  , w_1537 );
buf ( w_1535 , \554_b1 );
not ( w_1535 , w_1538 );
not (  , w_1539 );
and ( w_1538 , w_1539 , \554_b0 );
buf ( \556_b1 , \555_b1 );
not ( \556_b1 , w_1540 );
not ( \556_b0 , w_1541 );
and ( w_1540 , w_1541 , \555_b0 );
or ( \557_b1 , \193_b1 , \309_b1 );
xor ( \557_b0 , \193_b0 , w_1542 );
not ( w_1542 , w_1543 );
and ( w_1543 , \309_b1 , \309_b0 );
or ( \558_b1 , \557_b1 , \252_b1 );
xor ( \558_b0 , \557_b0 , w_1544 );
not ( w_1544 , w_1545 );
and ( w_1545 , \252_b1 , \252_b0 );
or ( \559_b1 , \556_b1 , w_1547 );
not ( w_1547 , w_1548 );
and ( \559_b0 , \556_b0 , w_1549 );
and ( w_1548 ,  , w_1549 );
buf ( w_1547 , \558_b1 );
not ( w_1547 , w_1550 );
not (  , w_1551 );
and ( w_1550 , w_1551 , \558_b0 );
or ( \560_b1 , \546_b1 , w_1553 );
not ( w_1553 , w_1554 );
and ( \560_b0 , \546_b0 , w_1555 );
and ( w_1554 ,  , w_1555 );
buf ( w_1553 , \559_b1 );
not ( w_1553 , w_1556 );
not (  , w_1557 );
and ( w_1556 , w_1557 , \559_b0 );
or ( \561_b1 , \415_b1 , w_1559 );
not ( w_1559 , w_1560 );
and ( \561_b0 , \415_b0 , w_1561 );
and ( w_1560 ,  , w_1561 );
buf ( w_1559 , \560_b1 );
not ( w_1559 , w_1562 );
not (  , w_1563 );
and ( w_1562 , w_1563 , \560_b0 );
buf ( \562_b1 , \561_b1 );
not ( \562_b1 , w_1564 );
not ( \562_b0 , w_1565 );
and ( w_1564 , w_1565 , \561_b0 );
or ( \563_b1 , \136_b1 , w_1567 );
not ( w_1567 , w_1568 );
and ( \563_b0 , \136_b0 , w_1569 );
and ( w_1568 ,  , w_1569 );
buf ( w_1567 , \B[0]_b1 );
not ( w_1567 , w_1570 );
not (  , w_1571 );
and ( w_1570 , w_1571 , \B[0]_b0 );
buf ( \564_b1 , \563_b1 );
not ( \564_b1 , w_1572 );
not ( \564_b0 , w_1573 );
and ( w_1572 , w_1573 , \563_b0 );
or ( \565_b1 , \95_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1574 );
and ( \565_b0 , \95_b0 , w_1575 );
and ( w_1574 , w_1575 , \B[1]_b0 );
buf ( \566_b1 , \565_b1 );
not ( \566_b1 , w_1576 );
not ( \566_b0 , w_1577 );
and ( w_1576 , w_1577 , \565_b0 );
or ( \567_b1 , \564_b1 , \566_b1 );
not ( \566_b1 , w_1578 );
and ( \567_b0 , \564_b0 , w_1579 );
and ( w_1578 , w_1579 , \566_b0 );
or ( \568_b1 , \563_b1 , \565_b1 );
not ( \565_b1 , w_1580 );
and ( \568_b0 , \563_b0 , w_1581 );
and ( w_1580 , w_1581 , \565_b0 );
or ( \569_b1 , \567_b1 , w_1583 );
not ( w_1583 , w_1584 );
and ( \569_b0 , \567_b0 , w_1585 );
and ( w_1584 ,  , w_1585 );
buf ( w_1583 , \568_b1 );
not ( w_1583 , w_1586 );
not (  , w_1587 );
and ( w_1586 , w_1587 , \568_b0 );
or ( \570_b1 , \111_b1 , w_1589 );
not ( w_1589 , w_1590 );
and ( \570_b0 , \111_b0 , w_1591 );
and ( w_1590 ,  , w_1591 );
buf ( w_1589 , \B[4]_b1 );
not ( w_1589 , w_1592 );
not (  , w_1593 );
and ( w_1592 , w_1593 , \B[4]_b0 );
or ( \571_b1 , \200_b1 , w_1595 );
not ( w_1595 , w_1596 );
and ( \571_b0 , \200_b0 , w_1597 );
and ( w_1596 ,  , w_1597 );
buf ( w_1595 , \B[2]_b1 );
not ( w_1595 , w_1598 );
not (  , w_1599 );
and ( w_1598 , w_1599 , \B[2]_b0 );
or ( \572_b1 , \570_b1 , \571_b1 );
xor ( \572_b0 , \570_b0 , w_1600 );
not ( w_1600 , w_1601 );
and ( w_1601 , \571_b1 , \571_b0 );
or ( \573_b1 , \104_b1 , w_1603 );
not ( w_1603 , w_1604 );
and ( \573_b0 , \104_b0 , w_1605 );
and ( w_1604 ,  , w_1605 );
buf ( w_1603 , \B[3]_b1 );
not ( w_1603 , w_1606 );
not (  , w_1607 );
and ( w_1606 , w_1607 , \B[3]_b0 );
or ( \574_b1 , \572_b1 , \573_b1 );
not ( \573_b1 , w_1608 );
and ( \574_b0 , \572_b0 , w_1609 );
and ( w_1608 , w_1609 , \573_b0 );
or ( \575_b1 , \570_b1 , \571_b1 );
not ( \571_b1 , w_1610 );
and ( \575_b0 , \570_b0 , w_1611 );
and ( w_1610 , w_1611 , \571_b0 );
or ( \576_b1 , \574_b1 , w_1612 );
or ( \576_b0 , \574_b0 , \575_b0 );
not ( \575_b0 , w_1613 );
and ( w_1613 , w_1612 , \575_b1 );
or ( \577_b1 , \569_b1 , \576_b1 );
xor ( \577_b0 , \569_b0 , w_1614 );
not ( w_1614 , w_1615 );
and ( w_1615 , \576_b1 , \576_b0 );
or ( \578_b1 , \104_b1 , w_1617 );
not ( w_1617 , w_1618 );
and ( \578_b0 , \104_b0 , w_1619 );
and ( w_1618 ,  , w_1619 );
buf ( w_1617 , \B[4]_b1 );
not ( w_1617 , w_1620 );
not (  , w_1621 );
and ( w_1620 , w_1621 , \B[4]_b0 );
or ( \579_b1 , \143_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_1622 );
and ( \579_b0 , \143_b0 , w_1623 );
and ( w_1622 , w_1623 , \B[3]_b0 );
or ( \580_b1 , \578_b1 , \579_b1 );
xor ( \580_b0 , \578_b0 , w_1624 );
not ( w_1624 , w_1625 );
and ( w_1625 , \579_b1 , \579_b0 );
or ( \581_b1 , \127_b1 , w_1627 );
not ( w_1627 , w_1628 );
and ( \581_b0 , \127_b0 , w_1629 );
and ( w_1628 ,  , w_1629 );
buf ( w_1627 , \B[2]_b1 );
not ( w_1627 , w_1630 );
not (  , w_1631 );
and ( w_1630 , w_1631 , \B[2]_b0 );
or ( \582_b1 , \580_b1 , w_1632 );
xor ( \582_b0 , \580_b0 , w_1634 );
not ( w_1634 , w_1635 );
and ( w_1635 , w_1632 , w_1633 );
buf ( w_1632 , \581_b1 );
not ( w_1632 , w_1636 );
not ( w_1633 , w_1637 );
and ( w_1636 , w_1637 , \581_b0 );
or ( \583_b1 , \577_b1 , \582_b1 );
not ( \582_b1 , w_1638 );
and ( \583_b0 , \577_b0 , w_1639 );
and ( w_1638 , w_1639 , \582_b0 );
or ( \584_b1 , \569_b1 , \576_b1 );
not ( \576_b1 , w_1640 );
and ( \584_b0 , \569_b0 , w_1641 );
and ( w_1640 , w_1641 , \576_b0 );
or ( \585_b1 , \583_b1 , w_1642 );
or ( \585_b0 , \583_b0 , \584_b0 );
not ( \584_b0 , w_1643 );
and ( w_1643 , w_1642 , \584_b1 );
buf ( \586_b1 , \585_b1 );
not ( \586_b1 , w_1644 );
not ( \586_b0 , w_1645 );
and ( w_1644 , w_1645 , \585_b0 );
buf ( \587_b1 , \565_b1 );
not ( \587_b1 , w_1646 );
not ( \587_b0 , w_1647 );
and ( w_1646 , w_1647 , \565_b0 );
or ( \588_b1 , \587_b1 , w_1649 );
not ( w_1649 , w_1650 );
and ( \588_b0 , \587_b0 , w_1651 );
and ( w_1650 ,  , w_1651 );
buf ( w_1649 , \563_b1 );
not ( w_1649 , w_1652 );
not (  , w_1653 );
and ( w_1652 , w_1653 , \563_b0 );
or ( \589_b1 , \472_b1 , \529_b1 );
xor ( \589_b0 , \472_b0 , w_1654 );
not ( w_1654 , w_1655 );
and ( w_1655 , \529_b1 , \529_b0 );
or ( \590_b1 , \588_b1 , \589_b1 );
xor ( \590_b0 , \588_b0 , w_1656 );
not ( w_1656 , w_1657 );
and ( w_1657 , \589_b1 , \589_b0 );
buf ( \591_b1 , \581_b1 );
not ( \591_b1 , w_1658 );
not ( \591_b0 , w_1659 );
and ( w_1658 , w_1659 , \581_b0 );
buf ( \592_b1 , \578_b1 );
not ( \592_b1 , w_1660 );
not ( \592_b0 , w_1661 );
and ( w_1660 , w_1661 , \578_b0 );
or ( \593_b1 , \591_b1 , w_1662 );
or ( \593_b0 , \591_b0 , \592_b0 );
not ( \592_b0 , w_1663 );
and ( w_1663 , w_1662 , \592_b1 );
or ( \594_b1 , \593_b1 , w_1665 );
not ( w_1665 , w_1666 );
and ( \594_b0 , \593_b0 , w_1667 );
and ( w_1666 ,  , w_1667 );
buf ( w_1665 , \579_b1 );
not ( w_1665 , w_1668 );
not (  , w_1669 );
and ( w_1668 , w_1669 , \579_b0 );
or ( \595_b1 , \578_b1 , w_1670 );
or ( \595_b0 , \578_b0 , \581_b0 );
not ( \581_b0 , w_1671 );
and ( w_1671 , w_1670 , \581_b1 );
or ( \596_b1 , \594_b1 , w_1673 );
not ( w_1673 , w_1674 );
and ( \596_b0 , \594_b0 , w_1675 );
and ( w_1674 ,  , w_1675 );
buf ( w_1673 , \595_b1 );
not ( w_1673 , w_1676 );
not (  , w_1677 );
and ( w_1676 , w_1677 , \595_b0 );
or ( \597_b1 , \590_b1 , \596_b1 );
xor ( \597_b0 , \590_b0 , w_1678 );
not ( w_1678 , w_1679 );
and ( w_1679 , \596_b1 , \596_b0 );
buf ( \598_b1 , \597_b1 );
not ( \598_b1 , w_1680 );
not ( \598_b0 , w_1681 );
and ( w_1680 , w_1681 , \597_b0 );
or ( \599_b1 , \586_b1 , \598_b1 );
not ( \598_b1 , w_1682 );
and ( \599_b0 , \586_b0 , w_1683 );
and ( w_1682 , w_1683 , \598_b0 );
or ( \600_b1 , \585_b1 , \597_b1 );
not ( \597_b1 , w_1684 );
and ( \600_b0 , \585_b0 , w_1685 );
and ( w_1684 , w_1685 , \597_b0 );
or ( \601_b1 , \599_b1 , w_1687 );
not ( w_1687 , w_1688 );
and ( \601_b0 , \599_b0 , w_1689 );
and ( w_1688 ,  , w_1689 );
buf ( w_1687 , \600_b1 );
not ( w_1687 , w_1690 );
not (  , w_1691 );
and ( w_1690 , w_1691 , \600_b0 );
or ( \602_b1 , \95_b1 , w_1693 );
not ( w_1693 , w_1694 );
and ( \602_b0 , \95_b0 , w_1695 );
and ( w_1694 ,  , w_1695 );
buf ( w_1693 , \B[2]_b1 );
not ( w_1693 , w_1696 );
not (  , w_1697 );
and ( w_1696 , w_1697 , \B[2]_b0 );
or ( \603_b1 , \104_b1 , w_1699 );
not ( w_1699 , w_1700 );
and ( \603_b0 , \104_b0 , w_1701 );
and ( w_1700 ,  , w_1701 );
buf ( w_1699 , \B[5]_b1 );
not ( w_1699 , w_1702 );
not (  , w_1703 );
and ( w_1702 , w_1703 , \B[5]_b0 );
or ( \604_b1 , \602_b1 , \603_b1 );
xor ( \604_b0 , \602_b0 , w_1704 );
not ( w_1704 , w_1705 );
and ( w_1705 , \603_b1 , \603_b0 );
or ( \605_b1 , \111_b1 , w_1707 );
not ( w_1707 , w_1708 );
and ( \605_b0 , \111_b0 , w_1709 );
and ( w_1708 ,  , w_1709 );
buf ( w_1707 , \B[6]_b1 );
not ( w_1707 , w_1710 );
not (  , w_1711 );
and ( w_1710 , w_1711 , \B[6]_b0 );
or ( \606_b1 , \604_b1 , \605_b1 );
xor ( \606_b0 , \604_b0 , w_1712 );
not ( w_1712 , w_1713 );
and ( w_1713 , \605_b1 , \605_b0 );
buf ( \607_b1 , \606_b1 );
not ( \607_b1 , w_1714 );
not ( \607_b0 , w_1715 );
and ( w_1714 , w_1715 , \606_b0 );
buf ( \608_b1 , \607_b1 );
not ( \608_b1 , w_1716 );
not ( \608_b0 , w_1717 );
and ( w_1716 , w_1717 , \607_b0 );
or ( \609_b1 , \118_b1 , w_1719 );
not ( w_1719 , w_1720 );
and ( \609_b0 , \118_b0 , w_1721 );
and ( w_1720 ,  , w_1721 );
buf ( w_1719 , \B[7]_b1 );
not ( w_1719 , w_1722 );
not (  , w_1723 );
and ( w_1722 , w_1723 , \B[7]_b0 );
or ( \610_b1 , \127_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_1724 );
and ( \610_b0 , \127_b0 , w_1725 );
and ( w_1724 , w_1725 , \B[3]_b0 );
or ( \611_b1 , \609_b1 , \610_b1 );
xor ( \611_b0 , \609_b0 , w_1726 );
not ( w_1726 , w_1727 );
and ( w_1727 , \610_b1 , \610_b0 );
or ( \612_b1 , \200_b1 , w_1729 );
not ( w_1729 , w_1730 );
and ( \612_b0 , \200_b0 , w_1731 );
and ( w_1730 ,  , w_1731 );
buf ( w_1729 , \B[4]_b1 );
not ( w_1729 , w_1732 );
not (  , w_1733 );
and ( w_1732 , w_1733 , \B[4]_b0 );
or ( \613_b1 , \611_b1 , w_1734 );
xor ( \613_b0 , \611_b0 , w_1736 );
not ( w_1736 , w_1737 );
and ( w_1737 , w_1734 , w_1735 );
buf ( w_1734 , \612_b1 );
not ( w_1734 , w_1738 );
not ( w_1735 , w_1739 );
and ( w_1738 , w_1739 , \612_b0 );
buf ( \614_b1 , \613_b1 );
not ( \614_b1 , w_1740 );
not ( \614_b0 , w_1741 );
and ( w_1740 , w_1741 , \613_b0 );
or ( \615_b1 , \608_b1 , w_1742 );
or ( \615_b0 , \608_b0 , \614_b0 );
not ( \614_b0 , w_1743 );
and ( w_1743 , w_1742 , \614_b1 );
buf ( \616_b1 , \613_b1 );
not ( \616_b1 , w_1744 );
not ( \616_b0 , w_1745 );
and ( w_1744 , w_1745 , \613_b0 );
or ( \617_b1 , \616_b1 , w_1747 );
not ( w_1747 , w_1748 );
and ( \617_b0 , \616_b0 , w_1749 );
and ( w_1748 ,  , w_1749 );
buf ( w_1747 , \606_b1 );
not ( w_1747 , w_1750 );
not (  , w_1751 );
and ( w_1750 , w_1751 , \606_b0 );
or ( \618_b1 , \615_b1 , w_1753 );
not ( w_1753 , w_1754 );
and ( \618_b0 , \615_b0 , w_1755 );
and ( w_1754 ,  , w_1755 );
buf ( w_1753 , \617_b1 );
not ( w_1753 , w_1756 );
not (  , w_1757 );
and ( w_1756 , w_1757 , \617_b0 );
or ( \619_b1 , \118_b1 , \B[6]_b1 );
not ( \B[6]_b1 , w_1758 );
and ( \619_b0 , \118_b0 , w_1759 );
and ( w_1758 , w_1759 , \B[6]_b0 );
buf ( \620_b1 , \619_b1 );
not ( \620_b1 , w_1760 );
not ( \620_b0 , w_1761 );
and ( w_1760 , w_1761 , \619_b0 );
or ( \621_b1 , \111_b1 , w_1763 );
not ( w_1763 , w_1764 );
and ( \621_b0 , \111_b0 , w_1765 );
and ( w_1764 ,  , w_1765 );
buf ( w_1763 , \B[5]_b1 );
not ( w_1763 , w_1766 );
not (  , w_1767 );
and ( w_1766 , w_1767 , \B[5]_b0 );
or ( \622_b1 , \620_b1 , w_1768 );
or ( \622_b0 , \620_b0 , \621_b0 );
not ( \621_b0 , w_1769 );
and ( w_1769 , w_1768 , \621_b1 );
buf ( \623_b1 , \621_b1 );
not ( \623_b1 , w_1770 );
not ( \623_b0 , w_1771 );
and ( w_1770 , w_1771 , \621_b0 );
buf ( \624_b1 , \620_b1 );
not ( \624_b1 , w_1772 );
not ( \624_b0 , w_1773 );
and ( w_1772 , w_1773 , \620_b0 );
or ( \625_b1 , \623_b1 , w_1774 );
or ( \625_b0 , \623_b0 , \624_b0 );
not ( \624_b0 , w_1775 );
and ( w_1775 , w_1774 , \624_b1 );
or ( \626_b1 , \127_b1 , w_1777 );
not ( w_1777 , w_1778 );
and ( \626_b0 , \127_b0 , w_1779 );
and ( w_1778 ,  , w_1779 );
buf ( w_1777 , \B[1]_b1 );
not ( w_1777 , w_1780 );
not (  , w_1781 );
and ( w_1780 , w_1781 , \B[1]_b0 );
buf ( \627_b1 , \626_b1 );
not ( \627_b1 , w_1782 );
not ( \627_b0 , w_1783 );
and ( w_1782 , w_1783 , \626_b0 );
or ( \628_b1 , \95_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_1784 );
and ( \628_b0 , \95_b0 , w_1785 );
and ( w_1784 , w_1785 , \B[0]_b0 );
or ( \629_b1 , \627_b1 , w_1787 );
not ( w_1787 , w_1788 );
and ( \629_b0 , \627_b0 , w_1789 );
and ( w_1788 ,  , w_1789 );
buf ( w_1787 , \628_b1 );
not ( w_1787 , w_1790 );
not (  , w_1791 );
and ( w_1790 , w_1791 , \628_b0 );
buf ( \630_b1 , \629_b1 );
not ( \630_b1 , w_1792 );
not ( \630_b0 , w_1793 );
and ( w_1792 , w_1793 , \629_b0 );
or ( \631_b1 , \625_b1 , w_1795 );
not ( w_1795 , w_1796 );
and ( \631_b0 , \625_b0 , w_1797 );
and ( w_1796 ,  , w_1797 );
buf ( w_1795 , \630_b1 );
not ( w_1795 , w_1798 );
not (  , w_1799 );
and ( w_1798 , w_1799 , \630_b0 );
or ( \632_b1 , \622_b1 , w_1801 );
not ( w_1801 , w_1802 );
and ( \632_b0 , \622_b0 , w_1803 );
and ( w_1802 ,  , w_1803 );
buf ( w_1801 , \631_b1 );
not ( w_1801 , w_1804 );
not (  , w_1805 );
and ( w_1804 , w_1805 , \631_b0 );
buf ( \633_b1 , \632_b1 );
not ( \633_b1 , w_1806 );
not ( \633_b0 , w_1807 );
and ( w_1806 , w_1807 , \632_b0 );
or ( \634_b1 , \618_b1 , \633_b1 );
not ( \633_b1 , w_1808 );
and ( \634_b0 , \618_b0 , w_1809 );
and ( w_1808 , w_1809 , \633_b0 );
buf ( \635_b1 , \618_b1 );
not ( \635_b1 , w_1810 );
not ( \635_b0 , w_1811 );
and ( w_1810 , w_1811 , \618_b0 );
or ( \636_b1 , \635_b1 , \632_b1 );
not ( \632_b1 , w_1812 );
and ( \636_b0 , \635_b0 , w_1813 );
and ( w_1812 , w_1813 , \632_b0 );
or ( \637_b1 , \634_b1 , w_1815 );
not ( w_1815 , w_1816 );
and ( \637_b0 , \634_b0 , w_1817 );
and ( w_1816 ,  , w_1817 );
buf ( w_1815 , \636_b1 );
not ( w_1815 , w_1818 );
not (  , w_1819 );
and ( w_1818 , w_1819 , \636_b0 );
buf ( \638_b1 , \637_b1 );
not ( \638_b1 , w_1820 );
not ( \638_b0 , w_1821 );
and ( w_1820 , w_1821 , \637_b0 );
or ( \639_b1 , \601_b1 , \638_b1 );
not ( \638_b1 , w_1822 );
and ( \639_b0 , \601_b0 , w_1823 );
and ( w_1822 , w_1823 , \638_b0 );
buf ( \640_b1 , \601_b1 );
not ( \640_b1 , w_1824 );
not ( \640_b0 , w_1825 );
and ( w_1824 , w_1825 , \601_b0 );
or ( \641_b1 , \640_b1 , \637_b1 );
not ( \637_b1 , w_1826 );
and ( \641_b0 , \640_b0 , w_1827 );
and ( w_1826 , w_1827 , \637_b0 );
or ( \642_b1 , \639_b1 , w_1829 );
not ( w_1829 , w_1830 );
and ( \642_b0 , \639_b0 , w_1831 );
and ( w_1830 ,  , w_1831 );
buf ( w_1829 , \641_b1 );
not ( w_1829 , w_1832 );
not (  , w_1833 );
and ( w_1832 , w_1833 , \641_b0 );
or ( \643_b1 , \619_b1 , \621_b1 );
xor ( \643_b0 , \619_b0 , w_1834 );
not ( w_1834 , w_1835 );
and ( w_1835 , \621_b1 , \621_b0 );
or ( \644_b1 , \643_b1 , w_1836 );
xor ( \644_b0 , \643_b0 , w_1838 );
not ( w_1838 , w_1839 );
and ( w_1839 , w_1836 , w_1837 );
buf ( w_1836 , \629_b1 );
not ( w_1836 , w_1840 );
not ( w_1837 , w_1841 );
and ( w_1840 , w_1841 , \629_b0 );
or ( \645_b1 , \118_b1 , w_1843 );
not ( w_1843 , w_1844 );
and ( \645_b0 , \118_b0 , w_1845 );
and ( w_1844 ,  , w_1845 );
buf ( w_1843 , \B[5]_b1 );
not ( w_1843 , w_1846 );
not (  , w_1847 );
and ( w_1846 , w_1847 , \B[5]_b0 );
or ( \646_b1 , \127_b1 , w_1849 );
not ( w_1849 , w_1850 );
and ( \646_b0 , \127_b0 , w_1851 );
and ( w_1850 ,  , w_1851 );
buf ( w_1849 , \B[0]_b1 );
not ( w_1849 , w_1852 );
not (  , w_1853 );
and ( w_1852 , w_1853 , \B[0]_b0 );
buf ( \647_b1 , \646_b1 );
not ( \647_b1 , w_1854 );
not ( \647_b0 , w_1855 );
and ( w_1854 , w_1855 , \646_b0 );
or ( \648_b1 , \143_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1856 );
and ( \648_b0 , \143_b0 , w_1857 );
and ( w_1856 , w_1857 , \B[1]_b0 );
or ( \649_b1 , \647_b1 , w_1859 );
not ( w_1859 , w_1860 );
and ( \649_b0 , \647_b0 , w_1861 );
and ( w_1860 ,  , w_1861 );
buf ( w_1859 , \648_b1 );
not ( w_1859 , w_1862 );
not (  , w_1863 );
and ( w_1862 , w_1863 , \648_b0 );
or ( \650_b1 , \645_b1 , \649_b1 );
xor ( \650_b0 , \645_b0 , w_1864 );
not ( w_1864 , w_1865 );
and ( w_1865 , \649_b1 , \649_b0 );
buf ( \651_b1 , \628_b1 );
not ( \651_b1 , w_1866 );
not ( \651_b0 , w_1867 );
and ( w_1866 , w_1867 , \628_b0 );
buf ( \652_b1 , \626_b1 );
not ( \652_b1 , w_1868 );
not ( \652_b0 , w_1869 );
and ( w_1868 , w_1869 , \626_b0 );
or ( \653_b1 , \651_b1 , \652_b1 );
not ( \652_b1 , w_1870 );
and ( \653_b0 , \651_b0 , w_1871 );
and ( w_1870 , w_1871 , \652_b0 );
or ( \654_b1 , \626_b1 , \628_b1 );
not ( \628_b1 , w_1872 );
and ( \654_b0 , \626_b0 , w_1873 );
and ( w_1872 , w_1873 , \628_b0 );
or ( \655_b1 , \653_b1 , w_1875 );
not ( w_1875 , w_1876 );
and ( \655_b0 , \653_b0 , w_1877 );
and ( w_1876 ,  , w_1877 );
buf ( w_1875 , \654_b1 );
not ( w_1875 , w_1878 );
not (  , w_1879 );
and ( w_1878 , w_1879 , \654_b0 );
or ( \656_b1 , \650_b1 , \655_b1 );
not ( \655_b1 , w_1880 );
and ( \656_b0 , \650_b0 , w_1881 );
and ( w_1880 , w_1881 , \655_b0 );
or ( \657_b1 , \645_b1 , \649_b1 );
not ( \649_b1 , w_1882 );
and ( \657_b0 , \645_b0 , w_1883 );
and ( w_1882 , w_1883 , \649_b0 );
or ( \658_b1 , \656_b1 , w_1884 );
or ( \658_b0 , \656_b0 , \657_b0 );
not ( \657_b0 , w_1885 );
and ( w_1885 , w_1884 , \657_b1 );
or ( \659_b1 , \644_b1 , \658_b1 );
xor ( \659_b0 , \644_b0 , w_1886 );
not ( w_1886 , w_1887 );
and ( w_1887 , \658_b1 , \658_b0 );
or ( \660_b1 , \569_b1 , \576_b1 );
xor ( \660_b0 , \569_b0 , w_1888 );
not ( w_1888 , w_1889 );
and ( w_1889 , \576_b1 , \576_b0 );
or ( \661_b1 , \660_b1 , \582_b1 );
xor ( \661_b0 , \660_b0 , w_1890 );
not ( w_1890 , w_1891 );
and ( w_1891 , \582_b1 , \582_b0 );
or ( \662_b1 , \659_b1 , \661_b1 );
not ( \661_b1 , w_1892 );
and ( \662_b0 , \659_b0 , w_1893 );
and ( w_1892 , w_1893 , \661_b0 );
or ( \663_b1 , \644_b1 , \658_b1 );
not ( \658_b1 , w_1894 );
and ( \663_b0 , \644_b0 , w_1895 );
and ( w_1894 , w_1895 , \658_b0 );
or ( \664_b1 , \662_b1 , w_1896 );
or ( \664_b0 , \662_b0 , \663_b0 );
not ( \663_b0 , w_1897 );
and ( w_1897 , w_1896 , \663_b1 );
or ( \665_b1 , \642_b1 , w_1899 );
not ( w_1899 , w_1900 );
and ( \665_b0 , \642_b0 , w_1901 );
and ( w_1900 ,  , w_1901 );
buf ( w_1899 , \664_b1 );
not ( w_1899 , w_1902 );
not (  , w_1903 );
and ( w_1902 , w_1903 , \664_b0 );
buf ( \666_b1 , \665_b1 );
not ( \666_b1 , w_1904 );
not ( \666_b0 , w_1905 );
and ( w_1904 , w_1905 , \665_b0 );
or ( \667_b1 , \644_b1 , \658_b1 );
xor ( \667_b0 , \644_b0 , w_1906 );
not ( w_1906 , w_1907 );
and ( w_1907 , \658_b1 , \658_b0 );
or ( \668_b1 , \667_b1 , \661_b1 );
xor ( \668_b0 , \667_b0 , w_1908 );
not ( w_1908 , w_1909 );
and ( w_1909 , \661_b1 , \661_b0 );
or ( \669_b1 , \118_b1 , w_1911 );
not ( w_1911 , w_1912 );
and ( \669_b0 , \118_b0 , w_1913 );
and ( w_1912 ,  , w_1913 );
buf ( w_1911 , \B[4]_b1 );
not ( w_1911 , w_1914 );
not (  , w_1915 );
and ( w_1914 , w_1915 , \B[4]_b0 );
or ( \670_b1 , \104_b1 , w_1917 );
not ( w_1917 , w_1918 );
and ( \670_b0 , \104_b0 , w_1919 );
and ( w_1918 ,  , w_1919 );
buf ( w_1917 , \B[2]_b1 );
not ( w_1917 , w_1920 );
not (  , w_1921 );
and ( w_1920 , w_1921 , \B[2]_b0 );
or ( \671_b1 , \669_b1 , \670_b1 );
xor ( \671_b0 , \669_b0 , w_1922 );
not ( w_1922 , w_1923 );
and ( w_1923 , \670_b1 , \670_b0 );
or ( \672_b1 , \111_b1 , w_1925 );
not ( w_1925 , w_1926 );
and ( \672_b0 , \111_b0 , w_1927 );
and ( w_1926 ,  , w_1927 );
buf ( w_1925 , \B[3]_b1 );
not ( w_1925 , w_1928 );
not (  , w_1929 );
and ( w_1928 , w_1929 , \B[3]_b0 );
or ( \673_b1 , \671_b1 , \672_b1 );
not ( \672_b1 , w_1930 );
and ( \673_b0 , \671_b0 , w_1931 );
and ( w_1930 , w_1931 , \672_b0 );
or ( \674_b1 , \669_b1 , \670_b1 );
not ( \670_b1 , w_1932 );
and ( \674_b0 , \669_b0 , w_1933 );
and ( w_1932 , w_1933 , \670_b0 );
or ( \675_b1 , \673_b1 , w_1934 );
or ( \675_b0 , \673_b0 , \674_b0 );
not ( \674_b0 , w_1935 );
and ( w_1935 , w_1934 , \674_b1 );
or ( \676_b1 , \570_b1 , \571_b1 );
xor ( \676_b0 , \570_b0 , w_1936 );
not ( w_1936 , w_1937 );
and ( w_1937 , \571_b1 , \571_b0 );
or ( \677_b1 , \676_b1 , \573_b1 );
xor ( \677_b0 , \676_b0 , w_1938 );
not ( w_1938 , w_1939 );
and ( w_1939 , \573_b1 , \573_b0 );
or ( \678_b1 , \675_b1 , \677_b1 );
xor ( \678_b0 , \675_b0 , w_1940 );
not ( w_1940 , w_1941 );
and ( w_1941 , \677_b1 , \677_b0 );
or ( \679_b1 , \645_b1 , \649_b1 );
xor ( \679_b0 , \645_b0 , w_1942 );
not ( w_1942 , w_1943 );
and ( w_1943 , \649_b1 , \649_b0 );
or ( \680_b1 , \679_b1 , \655_b1 );
xor ( \680_b0 , \679_b0 , w_1944 );
not ( w_1944 , w_1945 );
and ( w_1945 , \655_b1 , \655_b0 );
or ( \681_b1 , \678_b1 , \680_b1 );
not ( \680_b1 , w_1946 );
and ( \681_b0 , \678_b0 , w_1947 );
and ( w_1946 , w_1947 , \680_b0 );
or ( \682_b1 , \675_b1 , \677_b1 );
not ( \677_b1 , w_1948 );
and ( \682_b0 , \675_b0 , w_1949 );
and ( w_1948 , w_1949 , \677_b0 );
or ( \683_b1 , \681_b1 , w_1950 );
or ( \683_b0 , \681_b0 , \682_b0 );
not ( \682_b0 , w_1951 );
and ( w_1951 , w_1950 , \682_b1 );
or ( \684_b1 , \668_b1 , w_1953 );
not ( w_1953 , w_1954 );
and ( \684_b0 , \668_b0 , w_1955 );
and ( w_1954 ,  , w_1955 );
buf ( w_1953 , \683_b1 );
not ( w_1953 , w_1956 );
not (  , w_1957 );
and ( w_1956 , w_1957 , \683_b0 );
buf ( \685_b1 , \684_b1 );
not ( \685_b1 , w_1958 );
not ( \685_b0 , w_1959 );
and ( w_1958 , w_1959 , \684_b0 );
or ( \686_b1 , \675_b1 , \677_b1 );
xor ( \686_b0 , \675_b0 , w_1960 );
not ( w_1960 , w_1961 );
and ( w_1961 , \677_b1 , \677_b0 );
or ( \687_b1 , \686_b1 , \680_b1 );
xor ( \687_b0 , \686_b0 , w_1962 );
not ( w_1962 , w_1963 );
and ( w_1963 , \680_b1 , \680_b0 );
or ( \688_b1 , \200_b1 , w_1965 );
not ( w_1965 , w_1966 );
and ( \688_b0 , \200_b0 , w_1967 );
and ( w_1966 ,  , w_1967 );
buf ( w_1965 , \B[0]_b1 );
not ( w_1965 , w_1968 );
not (  , w_1969 );
and ( w_1968 , w_1969 , \B[0]_b0 );
buf ( \689_b1 , \688_b1 );
not ( \689_b1 , w_1970 );
not ( \689_b0 , w_1971 );
and ( w_1970 , w_1971 , \688_b0 );
or ( \690_b1 , \104_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_1972 );
and ( \690_b0 , \104_b0 , w_1973 );
and ( w_1972 , w_1973 , \B[1]_b0 );
or ( \691_b1 , \689_b1 , w_1975 );
not ( w_1975 , w_1976 );
and ( \691_b0 , \689_b0 , w_1977 );
and ( w_1976 ,  , w_1977 );
buf ( w_1975 , \690_b1 );
not ( w_1975 , w_1978 );
not (  , w_1979 );
and ( w_1978 , w_1979 , \690_b0 );
buf ( \692_b1 , \648_b1 );
not ( \692_b1 , w_1980 );
not ( \692_b0 , w_1981 );
and ( w_1980 , w_1981 , \648_b0 );
buf ( \693_b1 , \646_b1 );
not ( \693_b1 , w_1982 );
not ( \693_b0 , w_1983 );
and ( w_1982 , w_1983 , \646_b0 );
or ( \694_b1 , \692_b1 , \693_b1 );
not ( \693_b1 , w_1984 );
and ( \694_b0 , \692_b0 , w_1985 );
and ( w_1984 , w_1985 , \693_b0 );
or ( \695_b1 , \648_b1 , \646_b1 );
not ( \646_b1 , w_1986 );
and ( \695_b0 , \648_b0 , w_1987 );
and ( w_1986 , w_1987 , \646_b0 );
or ( \696_b1 , \694_b1 , w_1989 );
not ( w_1989 , w_1990 );
and ( \696_b0 , \694_b0 , w_1991 );
and ( w_1990 ,  , w_1991 );
buf ( w_1989 , \695_b1 );
not ( w_1989 , w_1992 );
not (  , w_1993 );
and ( w_1992 , w_1993 , \695_b0 );
or ( \697_b1 , \691_b1 , \696_b1 );
xor ( \697_b0 , \691_b0 , w_1994 );
not ( w_1994 , w_1995 );
and ( w_1995 , \696_b1 , \696_b0 );
or ( \698_b1 , \669_b1 , \670_b1 );
xor ( \698_b0 , \669_b0 , w_1996 );
not ( w_1996 , w_1997 );
and ( w_1997 , \670_b1 , \670_b0 );
or ( \699_b1 , \698_b1 , \672_b1 );
xor ( \699_b0 , \698_b0 , w_1998 );
not ( w_1998 , w_1999 );
and ( w_1999 , \672_b1 , \672_b0 );
or ( \700_b1 , \697_b1 , \699_b1 );
not ( \699_b1 , w_2000 );
and ( \700_b0 , \697_b0 , w_2001 );
and ( w_2000 , w_2001 , \699_b0 );
or ( \701_b1 , \691_b1 , \696_b1 );
not ( \696_b1 , w_2002 );
and ( \701_b0 , \691_b0 , w_2003 );
and ( w_2002 , w_2003 , \696_b0 );
or ( \702_b1 , \700_b1 , w_2004 );
or ( \702_b0 , \700_b0 , \701_b0 );
not ( \701_b0 , w_2005 );
and ( w_2005 , w_2004 , \701_b1 );
or ( \703_b1 , \687_b1 , w_2007 );
not ( w_2007 , w_2008 );
and ( \703_b0 , \687_b0 , w_2009 );
and ( w_2008 ,  , w_2009 );
buf ( w_2007 , \702_b1 );
not ( w_2007 , w_2010 );
not (  , w_2011 );
and ( w_2010 , w_2011 , \702_b0 );
buf ( \704_b1 , \703_b1 );
not ( \704_b1 , w_2012 );
not ( \704_b0 , w_2013 );
and ( w_2012 , w_2013 , \703_b0 );
or ( \705_b1 , \691_b1 , \696_b1 );
xor ( \705_b0 , \691_b0 , w_2014 );
not ( w_2014 , w_2015 );
and ( w_2015 , \696_b1 , \696_b0 );
or ( \706_b1 , \705_b1 , \699_b1 );
xor ( \706_b0 , \705_b0 , w_2016 );
not ( w_2016 , w_2017 );
and ( w_2017 , \699_b1 , \699_b0 );
buf ( \707_b1 , \690_b1 );
not ( \707_b1 , w_2018 );
not ( \707_b0 , w_2019 );
and ( w_2018 , w_2019 , \690_b0 );
buf ( \708_b1 , \688_b1 );
not ( \708_b1 , w_2020 );
not ( \708_b0 , w_2021 );
and ( w_2020 , w_2021 , \688_b0 );
or ( \709_b1 , \707_b1 , \708_b1 );
not ( \708_b1 , w_2022 );
and ( \709_b0 , \707_b0 , w_2023 );
and ( w_2022 , w_2023 , \708_b0 );
or ( \710_b1 , \688_b1 , \690_b1 );
not ( \690_b1 , w_2024 );
and ( \710_b0 , \688_b0 , w_2025 );
and ( w_2024 , w_2025 , \690_b0 );
or ( \711_b1 , \709_b1 , w_2027 );
not ( w_2027 , w_2028 );
and ( \711_b0 , \709_b0 , w_2029 );
and ( w_2028 ,  , w_2029 );
buf ( w_2027 , \710_b1 );
not ( w_2027 , w_2030 );
not (  , w_2031 );
and ( w_2030 , w_2031 , \710_b0 );
buf ( \712_b1 , \711_b1 );
not ( \712_b1 , w_2032 );
not ( \712_b0 , w_2033 );
and ( w_2032 , w_2033 , \711_b0 );
or ( \713_b1 , \118_b1 , \B[3]_b1 );
not ( \B[3]_b1 , w_2034 );
and ( \713_b0 , \118_b0 , w_2035 );
and ( w_2034 , w_2035 , \B[3]_b0 );
buf ( \714_b1 , \713_b1 );
not ( \714_b1 , w_2036 );
not ( \714_b0 , w_2037 );
and ( w_2036 , w_2037 , \713_b0 );
or ( \715_b1 , \111_b1 , w_2039 );
not ( w_2039 , w_2040 );
and ( \715_b0 , \111_b0 , w_2041 );
and ( w_2040 ,  , w_2041 );
buf ( w_2039 , \B[2]_b1 );
not ( w_2039 , w_2042 );
not (  , w_2043 );
and ( w_2042 , w_2043 , \B[2]_b0 );
or ( \716_b1 , \714_b1 , w_2045 );
not ( w_2045 , w_2046 );
and ( \716_b0 , \714_b0 , w_2047 );
and ( w_2046 ,  , w_2047 );
buf ( w_2045 , \715_b1 );
not ( w_2045 , w_2048 );
not (  , w_2049 );
and ( w_2048 , w_2049 , \715_b0 );
or ( \717_b1 , \712_b1 , w_2051 );
not ( w_2051 , w_2052 );
and ( \717_b0 , \712_b0 , w_2053 );
and ( w_2052 ,  , w_2053 );
buf ( w_2051 , \716_b1 );
not ( w_2051 , w_2054 );
not (  , w_2055 );
and ( w_2054 , w_2055 , \716_b0 );
buf ( \718_b1 , \715_b1 );
not ( \718_b1 , w_2056 );
not ( \718_b0 , w_2057 );
and ( w_2056 , w_2057 , \715_b0 );
or ( \719_b1 , \718_b1 , w_2059 );
not ( w_2059 , w_2060 );
and ( \719_b0 , \718_b0 , w_2061 );
and ( w_2060 ,  , w_2061 );
buf ( w_2059 , \713_b1 );
not ( w_2059 , w_2062 );
not (  , w_2063 );
and ( w_2062 , w_2063 , \713_b0 );
or ( \720_b1 , \717_b1 , \719_b1 );
not ( \719_b1 , w_2064 );
and ( \720_b0 , \717_b0 , w_2065 );
and ( w_2064 , w_2065 , \719_b0 );
or ( \721_b1 , \706_b1 , w_2066 );
or ( \721_b0 , \706_b0 , \720_b0 );
not ( \720_b0 , w_2067 );
and ( w_2067 , w_2066 , \720_b1 );
or ( \722_b1 , \104_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_2068 );
and ( \722_b0 , \104_b0 , w_2069 );
and ( w_2068 , w_2069 , \B[0]_b0 );
or ( \723_b1 , \118_b1 , \B[2]_b1 );
not ( \B[2]_b1 , w_2070 );
and ( \723_b0 , \118_b0 , w_2071 );
and ( w_2070 , w_2071 , \B[2]_b0 );
or ( \724_b1 , \722_b1 , \723_b1 );
not ( \723_b1 , w_2072 );
and ( \724_b0 , \722_b0 , w_2073 );
and ( w_2072 , w_2073 , \723_b0 );
buf ( \725_b1 , \724_b1 );
not ( \725_b1 , w_2074 );
not ( \725_b0 , w_2075 );
and ( w_2074 , w_2075 , \724_b0 );
buf ( \726_b1 , \711_b1 );
not ( \726_b1 , w_2076 );
not ( \726_b0 , w_2077 );
and ( w_2076 , w_2077 , \711_b0 );
buf ( \727_b1 , \715_b1 );
not ( \727_b1 , w_2078 );
not ( \727_b0 , w_2079 );
and ( w_2078 , w_2079 , \715_b0 );
buf ( \728_b1 , \713_b1 );
not ( \728_b1 , w_2080 );
not ( \728_b0 , w_2081 );
and ( w_2080 , w_2081 , \713_b0 );
or ( \729_b1 , \727_b1 , w_2082 );
or ( \729_b0 , \727_b0 , \728_b0 );
not ( \728_b0 , w_2083 );
and ( w_2083 , w_2082 , \728_b1 );
or ( \730_b1 , \713_b1 , w_2084 );
or ( \730_b0 , \713_b0 , \715_b0 );
not ( \715_b0 , w_2085 );
and ( w_2085 , w_2084 , \715_b1 );
or ( \731_b1 , \729_b1 , w_2087 );
not ( w_2087 , w_2088 );
and ( \731_b0 , \729_b0 , w_2089 );
and ( w_2088 ,  , w_2089 );
buf ( w_2087 , \730_b1 );
not ( w_2087 , w_2090 );
not (  , w_2091 );
and ( w_2090 , w_2091 , \730_b0 );
buf ( \732_b1 , \731_b1 );
not ( \732_b1 , w_2092 );
not ( \732_b0 , w_2093 );
and ( w_2092 , w_2093 , \731_b0 );
or ( \733_b1 , \726_b1 , \732_b1 );
not ( \732_b1 , w_2094 );
and ( \733_b0 , \726_b0 , w_2095 );
and ( w_2094 , w_2095 , \732_b0 );
or ( \734_b1 , \731_b1 , \711_b1 );
not ( \711_b1 , w_2096 );
and ( \734_b0 , \731_b0 , w_2097 );
and ( w_2096 , w_2097 , \711_b0 );
or ( \735_b1 , \733_b1 , w_2099 );
not ( w_2099 , w_2100 );
and ( \735_b0 , \733_b0 , w_2101 );
and ( w_2100 ,  , w_2101 );
buf ( w_2099 , \734_b1 );
not ( w_2099 , w_2102 );
not (  , w_2103 );
and ( w_2102 , w_2103 , \734_b0 );
or ( \736_b1 , \725_b1 , w_2105 );
not ( w_2105 , w_2106 );
and ( \736_b0 , \725_b0 , w_2107 );
and ( w_2106 ,  , w_2107 );
buf ( w_2105 , \735_b1 );
not ( w_2105 , w_2108 );
not (  , w_2109 );
and ( w_2108 , w_2109 , \735_b0 );
buf ( \737_b1 , \736_b1 );
not ( \737_b1 , w_2110 );
not ( \737_b0 , w_2111 );
and ( w_2110 , w_2111 , \736_b0 );
or ( \738_b1 , \111_b1 , w_2113 );
not ( w_2113 , w_2114 );
and ( \738_b0 , \111_b0 , w_2115 );
and ( w_2114 ,  , w_2115 );
buf ( w_2113 , \B[1]_b1 );
not ( w_2113 , w_2116 );
not (  , w_2117 );
and ( w_2116 , w_2117 , \B[1]_b0 );
buf ( \739_b1 , \738_b1 );
not ( \739_b1 , w_2118 );
not ( \739_b0 , w_2119 );
and ( w_2118 , w_2119 , \738_b0 );
or ( \740_b1 , \118_b1 , w_2121 );
not ( w_2121 , w_2122 );
and ( \740_b0 , \118_b0 , w_2123 );
and ( w_2122 ,  , w_2123 );
buf ( w_2121 , \B[0]_b1 );
not ( w_2121 , w_2124 );
not (  , w_2125 );
and ( w_2124 , w_2125 , \B[0]_b0 );
or ( \741_b1 , \738_b1 , w_2127 );
not ( w_2127 , w_2128 );
and ( \741_b0 , \738_b0 , w_2129 );
and ( w_2128 ,  , w_2129 );
buf ( w_2127 , \740_b1 );
not ( w_2127 , w_2130 );
not (  , w_2131 );
and ( w_2130 , w_2131 , \740_b0 );
or ( \742_b1 , \739_b1 , \741_b1 );
xor ( \742_b0 , \739_b0 , w_2132 );
not ( w_2132 , w_2133 );
and ( w_2133 , \741_b1 , \741_b0 );
or ( \743_b1 , \722_b1 , \723_b1 );
xor ( \743_b0 , \722_b0 , w_2134 );
not ( w_2134 , w_2135 );
and ( w_2135 , \723_b1 , \723_b0 );
or ( \744_b1 , \742_b1 , \743_b1 );
not ( \743_b1 , w_2136 );
and ( \744_b0 , \742_b0 , w_2137 );
and ( w_2136 , w_2137 , \743_b0 );
or ( \745_b1 , \739_b1 , \741_b1 );
not ( \741_b1 , w_2138 );
and ( \745_b0 , \739_b0 , w_2139 );
and ( w_2138 , w_2139 , \741_b0 );
or ( \746_b1 , \744_b1 , w_2140 );
or ( \746_b0 , \744_b0 , \745_b0 );
not ( \745_b0 , w_2141 );
and ( w_2141 , w_2140 , \745_b1 );
buf ( \747_b1 , \746_b1 );
not ( \747_b1 , w_2142 );
not ( \747_b0 , w_2143 );
and ( w_2142 , w_2143 , \746_b0 );
or ( \748_b1 , \737_b1 , w_2144 );
or ( \748_b0 , \737_b0 , \747_b0 );
not ( \747_b0 , w_2145 );
and ( w_2145 , w_2144 , \747_b1 );
buf ( \749_b1 , \735_b1 );
not ( \749_b1 , w_2146 );
not ( \749_b0 , w_2147 );
and ( w_2146 , w_2147 , \735_b0 );
or ( \750_b1 , \749_b1 , w_2149 );
not ( w_2149 , w_2150 );
and ( \750_b0 , \749_b0 , w_2151 );
and ( w_2150 ,  , w_2151 );
buf ( w_2149 , \724_b1 );
not ( w_2149 , w_2152 );
not (  , w_2153 );
and ( w_2152 , w_2153 , \724_b0 );
or ( \751_b1 , \748_b1 , w_2155 );
not ( w_2155 , w_2156 );
and ( \751_b0 , \748_b0 , w_2157 );
and ( w_2156 ,  , w_2157 );
buf ( w_2155 , \750_b1 );
not ( w_2155 , w_2158 );
not (  , w_2159 );
and ( w_2158 , w_2159 , \750_b0 );
or ( \752_b1 , \706_b1 , w_2161 );
not ( w_2161 , w_2162 );
and ( \752_b0 , \706_b0 , w_2163 );
and ( w_2162 ,  , w_2163 );
buf ( w_2161 , \720_b1 );
not ( w_2161 , w_2164 );
not (  , w_2165 );
and ( w_2164 , w_2165 , \720_b0 );
or ( \753_b1 , \751_b1 , w_2167 );
not ( w_2167 , w_2168 );
and ( \753_b0 , \751_b0 , w_2169 );
and ( w_2168 ,  , w_2169 );
buf ( w_2167 , \752_b1 );
not ( w_2167 , w_2170 );
not (  , w_2171 );
and ( w_2170 , w_2171 , \752_b0 );
or ( \754_b1 , \721_b1 , w_2173 );
not ( w_2173 , w_2174 );
and ( \754_b0 , \721_b0 , w_2175 );
and ( w_2174 ,  , w_2175 );
buf ( w_2173 , \753_b1 );
not ( w_2173 , w_2176 );
not (  , w_2177 );
and ( w_2176 , w_2177 , \753_b0 );
buf ( \755_b1 , \754_b1 );
not ( \755_b1 , w_2178 );
not ( \755_b0 , w_2179 );
and ( w_2178 , w_2179 , \754_b0 );
or ( \756_b1 , \704_b1 , w_2180 );
or ( \756_b0 , \704_b0 , \755_b0 );
not ( \755_b0 , w_2181 );
and ( w_2181 , w_2180 , \755_b1 );
or ( \757_b1 , \687_b1 , w_2182 );
or ( \757_b0 , \687_b0 , \702_b0 );
not ( \702_b0 , w_2183 );
and ( w_2183 , w_2182 , \702_b1 );
or ( \758_b1 , \756_b1 , w_2185 );
not ( w_2185 , w_2186 );
and ( \758_b0 , \756_b0 , w_2187 );
and ( w_2186 ,  , w_2187 );
buf ( w_2185 , \757_b1 );
not ( w_2185 , w_2188 );
not (  , w_2189 );
and ( w_2188 , w_2189 , \757_b0 );
buf ( \759_b1 , \758_b1 );
not ( \759_b1 , w_2190 );
not ( \759_b0 , w_2191 );
and ( w_2190 , w_2191 , \758_b0 );
or ( \760_b1 , \685_b1 , w_2192 );
or ( \760_b0 , \685_b0 , \759_b0 );
not ( \759_b0 , w_2193 );
and ( w_2193 , w_2192 , \759_b1 );
buf ( \761_b1 , \668_b1 );
not ( \761_b1 , w_2194 );
not ( \761_b0 , w_2195 );
and ( w_2194 , w_2195 , \668_b0 );
buf ( \762_b1 , \683_b1 );
not ( \762_b1 , w_2196 );
not ( \762_b0 , w_2197 );
and ( w_2196 , w_2197 , \683_b0 );
or ( \763_b1 , \761_b1 , w_2199 );
not ( w_2199 , w_2200 );
and ( \763_b0 , \761_b0 , w_2201 );
and ( w_2200 ,  , w_2201 );
buf ( w_2199 , \762_b1 );
not ( w_2199 , w_2202 );
not (  , w_2203 );
and ( w_2202 , w_2203 , \762_b0 );
or ( \764_b1 , \760_b1 , w_2205 );
not ( w_2205 , w_2206 );
and ( \764_b0 , \760_b0 , w_2207 );
and ( w_2206 ,  , w_2207 );
buf ( w_2205 , \763_b1 );
not ( w_2205 , w_2208 );
not (  , w_2209 );
and ( w_2208 , w_2209 , \763_b0 );
buf ( \765_b1 , \764_b1 );
not ( \765_b1 , w_2210 );
not ( \765_b0 , w_2211 );
and ( w_2210 , w_2211 , \764_b0 );
or ( \766_b1 , \666_b1 , w_2212 );
or ( \766_b0 , \666_b0 , \765_b0 );
not ( \765_b0 , w_2213 );
and ( w_2213 , w_2212 , \765_b1 );
buf ( \767_b1 , \642_b1 );
not ( \767_b1 , w_2214 );
not ( \767_b0 , w_2215 );
and ( w_2214 , w_2215 , \642_b0 );
buf ( \768_b1 , \664_b1 );
not ( \768_b1 , w_2216 );
not ( \768_b0 , w_2217 );
and ( w_2216 , w_2217 , \664_b0 );
or ( \769_b1 , \767_b1 , w_2219 );
not ( w_2219 , w_2220 );
and ( \769_b0 , \767_b0 , w_2221 );
and ( w_2220 ,  , w_2221 );
buf ( w_2219 , \768_b1 );
not ( w_2219 , w_2222 );
not (  , w_2223 );
and ( w_2222 , w_2223 , \768_b0 );
or ( \770_b1 , \766_b1 , w_2225 );
not ( w_2225 , w_2226 );
and ( \770_b0 , \766_b0 , w_2227 );
and ( w_2226 ,  , w_2227 );
buf ( w_2225 , \769_b1 );
not ( w_2225 , w_2228 );
not (  , w_2229 );
and ( w_2228 , w_2229 , \769_b0 );
buf ( \771_b1 , \606_b1 );
not ( \771_b1 , w_2230 );
not ( \771_b0 , w_2231 );
and ( w_2230 , w_2231 , \606_b0 );
buf ( \772_b1 , \613_b1 );
not ( \772_b1 , w_2232 );
not ( \772_b0 , w_2233 );
and ( w_2232 , w_2233 , \613_b0 );
or ( \773_b1 , \771_b1 , w_2234 );
or ( \773_b0 , \771_b0 , \772_b0 );
not ( \772_b0 , w_2235 );
and ( w_2235 , w_2234 , \772_b1 );
or ( \774_b1 , \773_b1 , w_2237 );
not ( w_2237 , w_2238 );
and ( \774_b0 , \773_b0 , w_2239 );
and ( w_2238 ,  , w_2239 );
buf ( w_2237 , \632_b1 );
not ( w_2237 , w_2240 );
not (  , w_2241 );
and ( w_2240 , w_2241 , \632_b0 );
or ( \775_b1 , \616_b1 , w_2243 );
not ( w_2243 , w_2244 );
and ( \775_b0 , \616_b0 , w_2245 );
and ( w_2244 ,  , w_2245 );
buf ( w_2243 , \607_b1 );
not ( w_2243 , w_2246 );
not (  , w_2247 );
and ( w_2246 , w_2247 , \607_b0 );
or ( \776_b1 , \774_b1 , w_2249 );
not ( w_2249 , w_2250 );
and ( \776_b0 , \774_b0 , w_2251 );
and ( w_2250 ,  , w_2251 );
buf ( w_2249 , \775_b1 );
not ( w_2249 , w_2252 );
not (  , w_2253 );
and ( w_2252 , w_2253 , \775_b0 );
buf ( \777_b1 , \612_b1 );
not ( \777_b1 , w_2254 );
not ( \777_b0 , w_2255 );
and ( w_2254 , w_2255 , \612_b0 );
buf ( \778_b1 , \609_b1 );
not ( \778_b1 , w_2256 );
not ( \778_b0 , w_2257 );
and ( w_2256 , w_2257 , \609_b0 );
or ( \779_b1 , \777_b1 , w_2258 );
or ( \779_b0 , \777_b0 , \778_b0 );
not ( \778_b0 , w_2259 );
and ( w_2259 , w_2258 , \778_b1 );
or ( \780_b1 , \779_b1 , w_2261 );
not ( w_2261 , w_2262 );
and ( \780_b0 , \779_b0 , w_2263 );
and ( w_2262 ,  , w_2263 );
buf ( w_2261 , \610_b1 );
not ( w_2261 , w_2264 );
not (  , w_2265 );
and ( w_2264 , w_2265 , \610_b0 );
or ( \781_b1 , \612_b1 , w_2266 );
or ( \781_b0 , \612_b0 , \609_b0 );
not ( \609_b0 , w_2267 );
and ( w_2267 , w_2266 , \609_b1 );
or ( \782_b1 , \780_b1 , w_2269 );
not ( w_2269 , w_2270 );
and ( \782_b0 , \780_b0 , w_2271 );
and ( w_2270 ,  , w_2271 );
buf ( w_2269 , \781_b1 );
not ( w_2269 , w_2272 );
not (  , w_2273 );
and ( w_2272 , w_2273 , \781_b0 );
buf ( \783_b1 , \603_b1 );
not ( \783_b1 , w_2274 );
not ( \783_b0 , w_2275 );
and ( w_2274 , w_2275 , \603_b0 );
buf ( \784_b1 , \605_b1 );
not ( \784_b1 , w_2276 );
not ( \784_b0 , w_2277 );
and ( w_2276 , w_2277 , \605_b0 );
or ( \785_b1 , \783_b1 , w_2278 );
or ( \785_b0 , \783_b0 , \784_b0 );
not ( \784_b0 , w_2279 );
and ( w_2279 , w_2278 , \784_b1 );
buf ( \786_b1 , \602_b1 );
not ( \786_b1 , w_2280 );
not ( \786_b0 , w_2281 );
and ( w_2280 , w_2281 , \602_b0 );
or ( \787_b1 , \785_b1 , w_2283 );
not ( w_2283 , w_2284 );
and ( \787_b0 , \785_b0 , w_2285 );
and ( w_2284 ,  , w_2285 );
buf ( w_2283 , \786_b1 );
not ( w_2283 , w_2286 );
not (  , w_2287 );
and ( w_2286 , w_2287 , \786_b0 );
or ( \788_b1 , \603_b1 , w_2288 );
or ( \788_b0 , \603_b0 , \605_b0 );
not ( \605_b0 , w_2289 );
and ( w_2289 , w_2288 , \605_b1 );
or ( \789_b1 , \787_b1 , w_2291 );
not ( w_2291 , w_2292 );
and ( \789_b0 , \787_b0 , w_2293 );
and ( w_2292 ,  , w_2293 );
buf ( w_2291 , \788_b1 );
not ( w_2291 , w_2294 );
not (  , w_2295 );
and ( w_2294 , w_2295 , \788_b0 );
or ( \790_b1 , \782_b1 , \789_b1 );
xor ( \790_b0 , \782_b0 , w_2296 );
not ( w_2296 , w_2297 );
and ( w_2297 , \789_b1 , \789_b0 );
or ( \791_b1 , \479_b1 , \476_b1 );
xor ( \791_b0 , \479_b0 , w_2298 );
not ( w_2298 , w_2299 );
and ( w_2299 , \476_b1 , \476_b0 );
buf ( \792_b1 , \474_b1 );
not ( \792_b1 , w_2300 );
not ( \792_b0 , w_2301 );
and ( w_2300 , w_2301 , \474_b0 );
or ( \793_b1 , \791_b1 , \792_b1 );
xor ( \793_b0 , \791_b0 , w_2302 );
not ( w_2302 , w_2303 );
and ( w_2303 , \792_b1 , \792_b0 );
buf ( \794_b1 , \793_b1 );
not ( \794_b1 , w_2304 );
not ( \794_b0 , w_2305 );
and ( w_2304 , w_2305 , \793_b0 );
or ( \795_b1 , \790_b1 , \794_b1 );
not ( \794_b1 , w_2306 );
and ( \795_b0 , \790_b0 , w_2307 );
and ( w_2306 , w_2307 , \794_b0 );
buf ( \796_b1 , \790_b1 );
not ( \796_b1 , w_2308 );
not ( \796_b0 , w_2309 );
and ( w_2308 , w_2309 , \790_b0 );
or ( \797_b1 , \796_b1 , \793_b1 );
not ( \793_b1 , w_2310 );
and ( \797_b0 , \796_b0 , w_2311 );
and ( w_2310 , w_2311 , \793_b0 );
or ( \798_b1 , \795_b1 , w_2313 );
not ( w_2313 , w_2314 );
and ( \798_b0 , \795_b0 , w_2315 );
and ( w_2314 ,  , w_2315 );
buf ( w_2313 , \797_b1 );
not ( w_2313 , w_2316 );
not (  , w_2317 );
and ( w_2316 , w_2317 , \797_b0 );
or ( \799_b1 , \776_b1 , \798_b1 );
xor ( \799_b0 , \776_b0 , w_2318 );
not ( w_2318 , w_2319 );
and ( w_2319 , \798_b1 , \798_b0 );
or ( \800_b1 , \488_b1 , \487_b1 );
xor ( \800_b0 , \488_b0 , w_2320 );
not ( w_2320 , w_2321 );
and ( w_2321 , \487_b1 , \487_b0 );
or ( \801_b1 , \800_b1 , \490_b1 );
xor ( \801_b0 , \800_b0 , w_2322 );
not ( w_2322 , w_2323 );
and ( w_2323 , \490_b1 , \490_b0 );
or ( \802_b1 , \520_b1 , \527_b1 );
xor ( \802_b0 , \520_b0 , w_2324 );
not ( w_2324 , w_2325 );
and ( w_2325 , \527_b1 , \527_b0 );
or ( \803_b1 , \802_b1 , \530_b1 );
xor ( \803_b0 , \802_b0 , w_2326 );
not ( w_2326 , w_2327 );
and ( w_2327 , \530_b1 , \530_b0 );
or ( \804_b1 , \801_b1 , \803_b1 );
xor ( \804_b0 , \801_b0 , w_2328 );
not ( w_2328 , w_2329 );
and ( w_2329 , \803_b1 , \803_b0 );
or ( \805_b1 , \588_b1 , \589_b1 );
xor ( \805_b0 , \588_b0 , w_2330 );
not ( w_2330 , w_2331 );
and ( w_2331 , \589_b1 , \589_b0 );
or ( \806_b1 , \805_b1 , \596_b1 );
not ( \596_b1 , w_2332 );
and ( \806_b0 , \805_b0 , w_2333 );
and ( w_2332 , w_2333 , \596_b0 );
or ( \807_b1 , \588_b1 , \589_b1 );
not ( \589_b1 , w_2334 );
and ( \807_b0 , \588_b0 , w_2335 );
and ( w_2334 , w_2335 , \589_b0 );
or ( \808_b1 , \806_b1 , w_2336 );
or ( \808_b0 , \806_b0 , \807_b0 );
not ( \807_b0 , w_2337 );
and ( w_2337 , w_2336 , \807_b1 );
or ( \809_b1 , \804_b1 , \808_b1 );
xor ( \809_b0 , \804_b0 , w_2338 );
not ( w_2338 , w_2339 );
and ( w_2339 , \808_b1 , \808_b0 );
or ( \810_b1 , \799_b1 , \809_b1 );
xor ( \810_b0 , \799_b0 , w_2340 );
not ( w_2340 , w_2341 );
and ( w_2341 , \809_b1 , \809_b0 );
buf ( \811_b1 , \810_b1 );
not ( \811_b1 , w_2342 );
not ( \811_b0 , w_2343 );
and ( w_2342 , w_2343 , \810_b0 );
buf ( \812_b1 , \597_b1 );
not ( \812_b1 , w_2344 );
not ( \812_b0 , w_2345 );
and ( w_2344 , w_2345 , \597_b0 );
buf ( \813_b1 , \638_b1 );
not ( \813_b1 , w_2346 );
not ( \813_b0 , w_2347 );
and ( w_2346 , w_2347 , \638_b0 );
or ( \814_b1 , \812_b1 , w_2348 );
or ( \814_b0 , \812_b0 , \813_b0 );
not ( \813_b0 , w_2349 );
and ( w_2349 , w_2348 , \813_b1 );
buf ( \815_b1 , \597_b1 );
not ( \815_b1 , w_2350 );
not ( \815_b0 , w_2351 );
and ( w_2350 , w_2351 , \597_b0 );
buf ( \816_b1 , \815_b1 );
not ( \816_b1 , w_2352 );
not ( \816_b0 , w_2353 );
and ( w_2352 , w_2353 , \815_b0 );
buf ( \817_b1 , \637_b1 );
not ( \817_b1 , w_2354 );
not ( \817_b0 , w_2355 );
and ( w_2354 , w_2355 , \637_b0 );
or ( \818_b1 , \816_b1 , w_2356 );
or ( \818_b0 , \816_b0 , \817_b0 );
not ( \817_b0 , w_2357 );
and ( w_2357 , w_2356 , \817_b1 );
buf ( \819_b1 , \585_b1 );
not ( \819_b1 , w_2358 );
not ( \819_b0 , w_2359 );
and ( w_2358 , w_2359 , \585_b0 );
or ( \820_b1 , \818_b1 , w_2361 );
not ( w_2361 , w_2362 );
and ( \820_b0 , \818_b0 , w_2363 );
and ( w_2362 ,  , w_2363 );
buf ( w_2361 , \819_b1 );
not ( w_2361 , w_2364 );
not (  , w_2365 );
and ( w_2364 , w_2365 , \819_b0 );
or ( \821_b1 , \814_b1 , w_2367 );
not ( w_2367 , w_2368 );
and ( \821_b0 , \814_b0 , w_2369 );
and ( w_2368 ,  , w_2369 );
buf ( w_2367 , \820_b1 );
not ( w_2367 , w_2370 );
not (  , w_2371 );
and ( w_2370 , w_2371 , \820_b0 );
buf ( \822_b1 , \821_b1 );
not ( \822_b1 , w_2372 );
not ( \822_b0 , w_2373 );
and ( w_2372 , w_2373 , \821_b0 );
or ( \823_b1 , \811_b1 , w_2375 );
not ( w_2375 , w_2376 );
and ( \823_b0 , \811_b0 , w_2377 );
and ( w_2376 ,  , w_2377 );
buf ( w_2375 , \822_b1 );
not ( w_2375 , w_2378 );
not (  , w_2379 );
and ( w_2378 , w_2379 , \822_b0 );
or ( \824_b1 , \770_b1 , w_2381 );
not ( w_2381 , w_2382 );
and ( \824_b0 , \770_b0 , w_2383 );
and ( w_2382 ,  , w_2383 );
buf ( w_2381 , \823_b1 );
not ( w_2381 , w_2384 );
not (  , w_2385 );
and ( w_2384 , w_2385 , \823_b0 );
or ( \825_b1 , \518_b1 , \515_b1 );
not ( \515_b1 , w_2386 );
and ( \825_b0 , \518_b0 , w_2387 );
and ( w_2386 , w_2387 , \515_b0 );
buf ( \826_b1 , \518_b1 );
not ( \826_b1 , w_2388 );
not ( \826_b0 , w_2389 );
and ( w_2388 , w_2389 , \518_b0 );
or ( \827_b1 , \826_b1 , \516_b1 );
not ( \516_b1 , w_2390 );
and ( \827_b0 , \826_b0 , w_2391 );
and ( w_2390 , w_2391 , \516_b0 );
or ( \828_b1 , \825_b1 , w_2392 );
or ( \828_b0 , \825_b0 , \827_b0 );
not ( \827_b0 , w_2393 );
and ( w_2393 , w_2392 , \827_b1 );
or ( \829_b1 , \828_b1 , \533_b1 );
xor ( \829_b0 , \828_b0 , w_2394 );
not ( w_2394 , w_2395 );
and ( w_2395 , \533_b1 , \533_b0 );
or ( \830_b1 , \801_b1 , \803_b1 );
xor ( \830_b0 , \801_b0 , w_2396 );
not ( w_2396 , w_2397 );
and ( w_2397 , \803_b1 , \803_b0 );
or ( \831_b1 , \830_b1 , \808_b1 );
not ( \808_b1 , w_2398 );
and ( \831_b0 , \830_b0 , w_2399 );
and ( w_2398 , w_2399 , \808_b0 );
or ( \832_b1 , \801_b1 , \803_b1 );
not ( \803_b1 , w_2400 );
and ( \832_b0 , \801_b0 , w_2401 );
and ( w_2400 , w_2401 , \803_b0 );
or ( \833_b1 , \831_b1 , w_2402 );
or ( \833_b0 , \831_b0 , \832_b0 );
not ( \832_b0 , w_2403 );
and ( w_2403 , w_2402 , \832_b1 );
or ( \834_b1 , \829_b1 , \833_b1 );
xor ( \834_b0 , \829_b0 , w_2404 );
not ( w_2404 , w_2405 );
and ( w_2405 , \833_b1 , \833_b0 );
or ( \835_b1 , \460_b1 , \461_b1 );
xor ( \835_b0 , \460_b0 , w_2406 );
not ( w_2406 , w_2407 );
and ( w_2407 , \461_b1 , \461_b0 );
or ( \836_b1 , \835_b1 , \467_b1 );
xor ( \836_b0 , \835_b0 , w_2408 );
not ( w_2408 , w_2409 );
and ( w_2409 , \467_b1 , \467_b0 );
or ( \837_b1 , \473_b1 , \485_b1 );
xor ( \837_b0 , \473_b0 , w_2410 );
not ( w_2410 , w_2411 );
and ( w_2411 , \485_b1 , \485_b0 );
or ( \838_b1 , \837_b1 , \493_b1 );
xor ( \838_b0 , \837_b0 , w_2412 );
not ( w_2412 , w_2413 );
and ( w_2413 , \493_b1 , \493_b0 );
or ( \839_b1 , \836_b1 , \838_b1 );
xor ( \839_b0 , \836_b0 , w_2414 );
not ( w_2414 , w_2415 );
and ( w_2415 , \838_b1 , \838_b0 );
or ( \840_b1 , \782_b1 , w_2416 );
or ( \840_b0 , \782_b0 , \789_b0 );
not ( \789_b0 , w_2417 );
and ( w_2417 , w_2416 , \789_b1 );
or ( \841_b1 , \840_b1 , \794_b1 );
not ( \794_b1 , w_2418 );
and ( \841_b0 , \840_b0 , w_2419 );
and ( w_2418 , w_2419 , \794_b0 );
or ( \842_b1 , \782_b1 , \789_b1 );
not ( \789_b1 , w_2420 );
and ( \842_b0 , \782_b0 , w_2421 );
and ( w_2420 , w_2421 , \789_b0 );
or ( \843_b1 , \841_b1 , w_2423 );
not ( w_2423 , w_2424 );
and ( \843_b0 , \841_b0 , w_2425 );
and ( w_2424 ,  , w_2425 );
buf ( w_2423 , \842_b1 );
not ( w_2423 , w_2426 );
not (  , w_2427 );
and ( w_2426 , w_2427 , \842_b0 );
or ( \844_b1 , \839_b1 , \843_b1 );
xor ( \844_b0 , \839_b0 , w_2428 );
not ( w_2428 , w_2429 );
and ( w_2429 , \843_b1 , \843_b0 );
buf ( \845_b1 , \844_b1 );
not ( \845_b1 , w_2430 );
not ( \845_b0 , w_2431 );
and ( w_2430 , w_2431 , \844_b0 );
or ( \846_b1 , \834_b1 , \845_b1 );
not ( \845_b1 , w_2432 );
and ( \846_b0 , \834_b0 , w_2433 );
and ( w_2432 , w_2433 , \845_b0 );
buf ( \847_b1 , \834_b1 );
not ( \847_b1 , w_2434 );
not ( \847_b0 , w_2435 );
and ( w_2434 , w_2435 , \834_b0 );
or ( \848_b1 , \847_b1 , \844_b1 );
not ( \844_b1 , w_2436 );
and ( \848_b0 , \847_b0 , w_2437 );
and ( w_2436 , w_2437 , \844_b0 );
or ( \849_b1 , \846_b1 , w_2439 );
not ( w_2439 , w_2440 );
and ( \849_b0 , \846_b0 , w_2441 );
and ( w_2440 ,  , w_2441 );
buf ( w_2439 , \848_b1 );
not ( w_2439 , w_2442 );
not (  , w_2443 );
and ( w_2442 , w_2443 , \848_b0 );
or ( \850_b1 , \776_b1 , \798_b1 );
xor ( \850_b0 , \776_b0 , w_2444 );
not ( w_2444 , w_2445 );
and ( w_2445 , \798_b1 , \798_b0 );
or ( \851_b1 , \850_b1 , \809_b1 );
not ( \809_b1 , w_2446 );
and ( \851_b0 , \850_b0 , w_2447 );
and ( w_2446 , w_2447 , \809_b0 );
or ( \852_b1 , \776_b1 , \798_b1 );
not ( \798_b1 , w_2448 );
and ( \852_b0 , \776_b0 , w_2449 );
and ( w_2448 , w_2449 , \798_b0 );
or ( \853_b1 , \851_b1 , w_2450 );
or ( \853_b0 , \851_b0 , \852_b0 );
not ( \852_b0 , w_2451 );
and ( w_2451 , w_2450 , \852_b1 );
or ( \854_b1 , \849_b1 , w_2453 );
not ( w_2453 , w_2454 );
and ( \854_b0 , \849_b0 , w_2455 );
and ( w_2454 ,  , w_2455 );
buf ( w_2453 , \853_b1 );
not ( w_2453 , w_2456 );
not (  , w_2457 );
and ( w_2456 , w_2457 , \853_b0 );
or ( \855_b1 , \810_b1 , w_2459 );
not ( w_2459 , w_2460 );
and ( \855_b0 , \810_b0 , w_2461 );
and ( w_2460 ,  , w_2461 );
buf ( w_2459 , \821_b1 );
not ( w_2459 , w_2462 );
not (  , w_2463 );
and ( w_2462 , w_2463 , \821_b0 );
or ( \856_b1 , \854_b1 , \855_b1 );
not ( \855_b1 , w_2464 );
and ( \856_b0 , \854_b0 , w_2465 );
and ( w_2464 , w_2465 , \855_b0 );
or ( \857_b1 , \824_b1 , w_2467 );
not ( w_2467 , w_2468 );
and ( \857_b0 , \824_b0 , w_2469 );
and ( w_2468 ,  , w_2469 );
buf ( w_2467 , \856_b1 );
not ( w_2467 , w_2470 );
not (  , w_2471 );
and ( w_2470 , w_2471 , \856_b0 );
buf ( \858_b1 , \857_b1 );
not ( \858_b1 , w_2472 );
not ( \858_b0 , w_2473 );
and ( w_2472 , w_2473 , \857_b0 );
or ( \859_b1 , \459_b1 , \470_b1 );
xor ( \859_b0 , \459_b0 , w_2474 );
not ( w_2474 , w_2475 );
and ( w_2475 , \470_b1 , \470_b0 );
or ( \860_b1 , \859_b1 , \496_b1 );
xor ( \860_b0 , \859_b0 , w_2476 );
not ( w_2476 , w_2477 );
and ( w_2477 , \496_b1 , \496_b0 );
buf ( \861_b1 , \860_b1 );
not ( \861_b1 , w_2478 );
not ( \861_b0 , w_2479 );
and ( w_2478 , w_2479 , \860_b0 );
or ( \862_b1 , \836_b1 , \838_b1 );
xor ( \862_b0 , \836_b0 , w_2480 );
not ( w_2480 , w_2481 );
and ( w_2481 , \838_b1 , \838_b0 );
or ( \863_b1 , \862_b1 , \843_b1 );
not ( \843_b1 , w_2482 );
and ( \863_b0 , \862_b0 , w_2483 );
and ( w_2482 , w_2483 , \843_b0 );
or ( \864_b1 , \836_b1 , \838_b1 );
not ( \838_b1 , w_2484 );
and ( \864_b0 , \836_b0 , w_2485 );
and ( w_2484 , w_2485 , \838_b0 );
or ( \865_b1 , \863_b1 , w_2486 );
or ( \865_b0 , \863_b0 , \864_b0 );
not ( \864_b0 , w_2487 );
and ( w_2487 , w_2486 , \864_b1 );
buf ( \866_b1 , \865_b1 );
not ( \866_b1 , w_2488 );
not ( \866_b0 , w_2489 );
and ( w_2488 , w_2489 , \865_b0 );
buf ( \867_b1 , \866_b1 );
not ( \867_b1 , w_2490 );
not ( \867_b0 , w_2491 );
and ( w_2490 , w_2491 , \866_b0 );
or ( \868_b1 , \861_b1 , w_2492 );
or ( \868_b0 , \861_b0 , \867_b0 );
not ( \867_b0 , w_2493 );
and ( w_2493 , w_2492 , \867_b1 );
buf ( \869_b1 , \860_b1 );
not ( \869_b1 , w_2494 );
not ( \869_b0 , w_2495 );
and ( w_2494 , w_2495 , \860_b0 );
or ( \870_b1 , \869_b1 , w_2497 );
not ( w_2497 , w_2498 );
and ( \870_b0 , \869_b0 , w_2499 );
and ( w_2498 ,  , w_2499 );
buf ( w_2497 , \865_b1 );
not ( w_2497 , w_2500 );
not (  , w_2501 );
and ( w_2500 , w_2501 , \865_b0 );
or ( \871_b1 , \868_b1 , w_2503 );
not ( w_2503 , w_2504 );
and ( \871_b0 , \868_b0 , w_2505 );
and ( w_2504 ,  , w_2505 );
buf ( w_2503 , \870_b1 );
not ( w_2503 , w_2506 );
not (  , w_2507 );
and ( w_2506 , w_2507 , \870_b0 );
or ( \872_b1 , \507_b1 , \509_b1 );
xor ( \872_b0 , \507_b0 , w_2508 );
not ( w_2508 , w_2509 );
and ( w_2509 , \509_b1 , \509_b0 );
or ( \873_b1 , \872_b1 , \536_b1 );
xor ( \873_b0 , \872_b0 , w_2510 );
not ( w_2510 , w_2511 );
and ( w_2511 , \536_b1 , \536_b0 );
or ( \874_b1 , \871_b1 , \873_b1 );
xor ( \874_b0 , \871_b0 , w_2512 );
not ( w_2512 , w_2513 );
and ( w_2513 , \873_b1 , \873_b0 );
or ( \875_b1 , \833_b1 , w_2514 );
or ( \875_b0 , \833_b0 , \829_b0 );
not ( \829_b0 , w_2515 );
and ( w_2515 , w_2514 , \829_b1 );
or ( \876_b1 , \845_b1 , \875_b1 );
not ( \875_b1 , w_2516 );
and ( \876_b0 , \845_b0 , w_2517 );
and ( w_2516 , w_2517 , \875_b0 );
or ( \877_b1 , \829_b1 , \833_b1 );
not ( \833_b1 , w_2518 );
and ( \877_b0 , \829_b0 , w_2519 );
and ( w_2518 , w_2519 , \833_b0 );
or ( \878_b1 , \876_b1 , w_2521 );
not ( w_2521 , w_2522 );
and ( \878_b0 , \876_b0 , w_2523 );
and ( w_2522 ,  , w_2523 );
buf ( w_2521 , \877_b1 );
not ( w_2521 , w_2524 );
not (  , w_2525 );
and ( w_2524 , w_2525 , \877_b0 );
or ( \879_b1 , \874_b1 , w_2527 );
not ( w_2527 , w_2528 );
and ( \879_b0 , \874_b0 , w_2529 );
and ( w_2528 ,  , w_2529 );
buf ( w_2527 , \878_b1 );
not ( w_2527 , w_2530 );
not (  , w_2531 );
and ( w_2530 , w_2531 , \878_b0 );
buf ( \880_b1 , \849_b1 );
not ( \880_b1 , w_2532 );
not ( \880_b0 , w_2533 );
and ( w_2532 , w_2533 , \849_b0 );
buf ( \881_b1 , \853_b1 );
not ( \881_b1 , w_2534 );
not ( \881_b0 , w_2535 );
and ( w_2534 , w_2535 , \853_b0 );
or ( \882_b1 , \880_b1 , w_2537 );
not ( w_2537 , w_2538 );
and ( \882_b0 , \880_b0 , w_2539 );
and ( w_2538 ,  , w_2539 );
buf ( w_2537 , \881_b1 );
not ( w_2537 , w_2540 );
not (  , w_2541 );
and ( w_2540 , w_2541 , \881_b0 );
or ( \883_b1 , \879_b1 , w_2543 );
not ( w_2543 , w_2544 );
and ( \883_b0 , \879_b0 , w_2545 );
and ( w_2544 ,  , w_2545 );
buf ( w_2543 , \882_b1 );
not ( w_2543 , w_2546 );
not (  , w_2547 );
and ( w_2546 , w_2547 , \882_b0 );
or ( \884_b1 , \505_b1 , \539_b1 );
xor ( \884_b0 , \505_b0 , w_2548 );
not ( w_2548 , w_2549 );
and ( w_2549 , \539_b1 , \539_b0 );
or ( \885_b1 , \884_b1 , w_2550 );
xor ( \885_b0 , \884_b0 , w_2552 );
not ( w_2552 , w_2553 );
and ( w_2553 , w_2550 , w_2551 );
buf ( w_2550 , \542_b1 );
not ( w_2550 , w_2554 );
not ( w_2551 , w_2555 );
and ( w_2554 , w_2555 , \542_b0 );
buf ( \886_b1 , \860_b1 );
not ( \886_b1 , w_2556 );
not ( \886_b0 , w_2557 );
and ( w_2556 , w_2557 , \860_b0 );
buf ( \887_b1 , \873_b1 );
not ( \887_b1 , w_2558 );
not ( \887_b0 , w_2559 );
and ( w_2558 , w_2559 , \873_b0 );
or ( \888_b1 , \886_b1 , w_2560 );
or ( \888_b0 , \886_b0 , \887_b0 );
not ( \887_b0 , w_2561 );
and ( w_2561 , w_2560 , \887_b1 );
buf ( \889_b1 , \865_b1 );
not ( \889_b1 , w_2562 );
not ( \889_b0 , w_2563 );
and ( w_2562 , w_2563 , \865_b0 );
or ( \890_b1 , \888_b1 , w_2565 );
not ( w_2565 , w_2566 );
and ( \890_b0 , \888_b0 , w_2567 );
and ( w_2566 ,  , w_2567 );
buf ( w_2565 , \889_b1 );
not ( w_2565 , w_2568 );
not (  , w_2569 );
and ( w_2568 , w_2569 , \889_b0 );
buf ( \891_b1 , \860_b1 );
not ( \891_b1 , w_2570 );
not ( \891_b0 , w_2571 );
and ( w_2570 , w_2571 , \860_b0 );
buf ( \892_b1 , \873_b1 );
not ( \892_b1 , w_2572 );
not ( \892_b0 , w_2573 );
and ( w_2572 , w_2573 , \873_b0 );
or ( \893_b1 , \891_b1 , w_2575 );
not ( w_2575 , w_2576 );
and ( \893_b0 , \891_b0 , w_2577 );
and ( w_2576 ,  , w_2577 );
buf ( w_2575 , \892_b1 );
not ( w_2575 , w_2578 );
not (  , w_2579 );
and ( w_2578 , w_2579 , \892_b0 );
or ( \894_b1 , \890_b1 , w_2581 );
not ( w_2581 , w_2582 );
and ( \894_b0 , \890_b0 , w_2583 );
and ( w_2582 ,  , w_2583 );
buf ( w_2581 , \893_b1 );
not ( w_2581 , w_2584 );
not (  , w_2585 );
and ( w_2584 , w_2585 , \893_b0 );
or ( \895_b1 , \885_b1 , w_2587 );
not ( w_2587 , w_2588 );
and ( \895_b0 , \885_b0 , w_2589 );
and ( w_2588 ,  , w_2589 );
buf ( w_2587 , \894_b1 );
not ( w_2587 , w_2590 );
not (  , w_2591 );
and ( w_2590 , w_2591 , \894_b0 );
or ( \896_b1 , \883_b1 , w_2593 );
not ( w_2593 , w_2594 );
and ( \896_b0 , \883_b0 , w_2595 );
and ( w_2594 ,  , w_2595 );
buf ( w_2593 , \895_b1 );
not ( w_2593 , w_2596 );
not (  , w_2597 );
and ( w_2596 , w_2597 , \895_b0 );
buf ( \897_b1 , \896_b1 );
not ( \897_b1 , w_2598 );
not ( \897_b0 , w_2599 );
and ( w_2598 , w_2599 , \896_b0 );
or ( \898_b1 , \858_b1 , w_2600 );
or ( \898_b0 , \858_b0 , \897_b0 );
not ( \897_b0 , w_2601 );
and ( w_2601 , w_2600 , \897_b1 );
or ( \899_b1 , \505_b1 , \539_b1 );
xor ( \899_b0 , \505_b0 , w_2602 );
not ( w_2602 , w_2603 );
and ( w_2603 , \539_b1 , \539_b0 );
or ( \900_b1 , \899_b1 , \542_b1 );
xor ( \900_b0 , \899_b0 , w_2604 );
not ( w_2604 , w_2605 );
and ( w_2605 , \542_b1 , \542_b0 );
buf ( \901_b1 , \894_b1 );
not ( \901_b1 , w_2606 );
not ( \901_b0 , w_2607 );
and ( w_2606 , w_2607 , \894_b0 );
or ( \902_b1 , \900_b1 , w_2609 );
not ( w_2609 , w_2610 );
and ( \902_b0 , \900_b0 , w_2611 );
and ( w_2610 ,  , w_2611 );
buf ( w_2609 , \901_b1 );
not ( w_2609 , w_2612 );
not (  , w_2613 );
and ( w_2612 , w_2613 , \901_b0 );
or ( \903_b1 , \874_b1 , w_2615 );
not ( w_2615 , w_2616 );
and ( \903_b0 , \874_b0 , w_2617 );
and ( w_2616 ,  , w_2617 );
buf ( w_2615 , \878_b1 );
not ( w_2615 , w_2618 );
not (  , w_2619 );
and ( w_2618 , w_2619 , \878_b0 );
or ( \904_b1 , \902_b1 , \903_b1 );
not ( \903_b1 , w_2620 );
and ( \904_b0 , \902_b0 , w_2621 );
and ( w_2620 , w_2621 , \903_b0 );
or ( \905_b1 , \900_b1 , w_2623 );
not ( w_2623 , w_2624 );
and ( \905_b0 , \900_b0 , w_2625 );
and ( w_2624 ,  , w_2625 );
buf ( w_2623 , \901_b1 );
not ( w_2623 , w_2626 );
not (  , w_2627 );
and ( w_2626 , w_2627 , \901_b0 );
or ( \906_b1 , \904_b1 , w_2629 );
not ( w_2629 , w_2630 );
and ( \906_b0 , \904_b0 , w_2631 );
and ( w_2630 ,  , w_2631 );
buf ( w_2629 , \905_b1 );
not ( w_2629 , w_2632 );
not (  , w_2633 );
and ( w_2632 , w_2633 , \905_b0 );
or ( \907_b1 , \898_b1 , w_2635 );
not ( w_2635 , w_2636 );
and ( \907_b0 , \898_b0 , w_2637 );
and ( w_2636 ,  , w_2637 );
buf ( w_2635 , \906_b1 );
not ( w_2635 , w_2638 );
not (  , w_2639 );
and ( w_2638 , w_2639 , \906_b0 );
buf ( \908_b1 , \907_b1 );
not ( \908_b1 , w_2640 );
not ( \908_b0 , w_2641 );
and ( w_2640 , w_2641 , \907_b0 );
or ( \909_b1 , \562_b1 , w_2642 );
or ( \909_b0 , \562_b0 , \908_b0 );
not ( \908_b0 , w_2643 );
and ( w_2643 , w_2642 , \908_b1 );
buf ( \910_b1 , \559_b1 );
not ( \910_b1 , w_2644 );
not ( \910_b0 , w_2645 );
and ( w_2644 , w_2645 , \559_b0 );
or ( \911_b1 , \503_b1 , w_2647 );
not ( w_2647 , w_2648 );
and ( \911_b0 , \503_b0 , w_2649 );
and ( w_2648 ,  , w_2649 );
buf ( w_2647 , \545_b1 );
not ( w_2647 , w_2650 );
not (  , w_2651 );
and ( w_2650 , w_2651 , \545_b0 );
buf ( \912_b1 , \911_b1 );
not ( \912_b1 , w_2652 );
not ( \912_b0 , w_2653 );
and ( w_2652 , w_2653 , \911_b0 );
or ( \913_b1 , \910_b1 , w_2654 );
or ( \913_b0 , \910_b0 , \912_b0 );
not ( \912_b0 , w_2655 );
and ( w_2655 , w_2654 , \912_b1 );
buf ( \914_b1 , \558_b1 );
not ( \914_b1 , w_2656 );
not ( \914_b0 , w_2657 );
and ( w_2656 , w_2657 , \558_b0 );
or ( \915_b1 , \914_b1 , w_2659 );
not ( w_2659 , w_2660 );
and ( \915_b0 , \914_b0 , w_2661 );
and ( w_2660 ,  , w_2661 );
buf ( w_2659 , \555_b1 );
not ( w_2659 , w_2662 );
not (  , w_2663 );
and ( w_2662 , w_2663 , \555_b0 );
or ( \916_b1 , \913_b1 , w_2665 );
not ( w_2665 , w_2666 );
and ( \916_b0 , \913_b0 , w_2667 );
and ( w_2666 ,  , w_2667 );
buf ( w_2665 , \915_b1 );
not ( w_2665 , w_2668 );
not (  , w_2669 );
and ( w_2668 , w_2669 , \915_b0 );
or ( \917_b1 , \916_b1 , w_2671 );
not ( w_2671 , w_2672 );
and ( \917_b0 , \916_b0 , w_2673 );
and ( w_2672 ,  , w_2673 );
buf ( w_2671 , \414_b1 );
not ( w_2671 , w_2674 );
not (  , w_2675 );
and ( w_2674 , w_2675 , \414_b0 );
buf ( \918_b1 , \412_b1 );
not ( \918_b1 , w_2676 );
not ( \918_b0 , w_2677 );
and ( w_2676 , w_2677 , \412_b0 );
or ( \919_b1 , \313_b1 , w_2679 );
not ( w_2679 , w_2680 );
and ( \919_b0 , \313_b0 , w_2681 );
and ( w_2680 ,  , w_2681 );
buf ( w_2679 , \357_b1 );
not ( w_2679 , w_2682 );
not (  , w_2683 );
and ( w_2682 , w_2683 , \357_b0 );
or ( \920_b1 , \919_b1 , w_2685 );
not ( w_2685 , w_2686 );
and ( \920_b0 , \919_b0 , w_2687 );
and ( w_2686 ,  , w_2687 );
buf ( w_2685 , \386_b1 );
not ( w_2685 , w_2688 );
not (  , w_2689 );
and ( w_2688 , w_2689 , \386_b0 );
buf ( \921_b1 , \385_b1 );
not ( \921_b1 , w_2690 );
not ( \921_b0 , w_2691 );
and ( w_2690 , w_2691 , \385_b0 );
or ( \922_b1 , \921_b1 , w_2693 );
not ( w_2693 , w_2694 );
and ( \922_b0 , \921_b0 , w_2695 );
and ( w_2694 ,  , w_2695 );
buf ( w_2693 , \380_b1 );
not ( w_2693 , w_2696 );
not (  , w_2697 );
and ( w_2696 , w_2697 , \380_b0 );
or ( \923_b1 , \920_b1 , w_2699 );
not ( w_2699 , w_2700 );
and ( \923_b0 , \920_b0 , w_2701 );
and ( w_2700 ,  , w_2701 );
buf ( w_2699 , \922_b1 );
not ( w_2699 , w_2702 );
not (  , w_2703 );
and ( w_2702 , w_2703 , \922_b0 );
or ( \924_b1 , \918_b1 , w_2705 );
not ( w_2705 , w_2706 );
and ( \924_b0 , \918_b0 , w_2707 );
and ( w_2706 ,  , w_2707 );
buf ( w_2705 , \923_b1 );
not ( w_2705 , w_2708 );
not (  , w_2709 );
and ( w_2708 , w_2709 , \923_b0 );
or ( \925_b1 , \409_b1 , w_2711 );
not ( w_2711 , w_2712 );
and ( \925_b0 , \409_b0 , w_2713 );
and ( w_2712 ,  , w_2713 );
buf ( w_2711 , \411_b1 );
not ( w_2711 , w_2714 );
not (  , w_2715 );
and ( w_2714 , w_2715 , \411_b0 );
or ( \926_b1 , \924_b1 , w_2716 );
or ( \926_b0 , \924_b0 , \925_b0 );
not ( \925_b0 , w_2717 );
and ( w_2717 , w_2716 , \925_b1 );
or ( \927_b1 , \926_b1 , w_2719 );
not ( w_2719 , w_2720 );
and ( \927_b0 , \926_b0 , w_2721 );
and ( w_2720 ,  , w_2721 );
buf ( w_2719 , \405_b1 );
not ( w_2719 , w_2722 );
not (  , w_2723 );
and ( w_2722 , w_2723 , \405_b0 );
or ( \928_b1 , \402_b1 , w_2724 );
or ( \928_b0 , \402_b0 , \404_b0 );
not ( \404_b0 , w_2725 );
and ( w_2725 , w_2724 , \404_b1 );
or ( \930_b1 , \909_b1 , w_2727 );
not ( w_2727 , w_2728 );
and ( \930_b0 , \909_b0 , w_2729 );
and ( w_2728 ,  , w_2729 );
buf ( w_2727 , \929_b1 );
not ( w_2727 , w_2730 );
not (  , w_2731 );
and ( w_2730 , w_2731 , \929_b0 );
buf ( \931_b1 , \930_b1 );
not ( \931_b1 , w_2732 );
not ( \931_b0 , w_2733 );
and ( w_2732 , w_2733 , \930_b0 );
or ( \932_b1 , \168_b1 , w_2734 );
or ( \932_b0 , \168_b0 , \931_b0 );
not ( \931_b0 , w_2735 );
and ( w_2735 , w_2734 , \931_b1 );
or ( \933_b1 , \165_b1 , w_2736 );
or ( \933_b0 , \165_b0 , \166_b0 );
not ( \166_b0 , w_2737 );
and ( w_2737 , w_2736 , \166_b1 );
or ( \934_b1 , \932_b1 , w_2739 );
not ( w_2739 , w_2740 );
and ( \934_b0 , \932_b0 , w_2741 );
and ( w_2740 ,  , w_2741 );
buf ( w_2739 , \933_b1 );
not ( w_2739 , w_2742 );
not (  , w_2743 );
and ( w_2742 , w_2743 , \933_b0 );
or ( \935_b1 , \167_b1 , w_2745 );
not ( w_2745 , w_2746 );
and ( \935_b0 , \167_b0 , w_2747 );
and ( w_2746 ,  , w_2747 );
buf ( w_2745 , \933_b1 );
not ( w_2745 , w_2748 );
not (  , w_2749 );
and ( w_2748 , w_2749 , \933_b0 );
buf ( \936_b1 , \935_b1 );
not ( \936_b1 , w_2750 );
not ( \936_b0 , w_2751 );
and ( w_2750 , w_2751 , \935_b0 );
buf ( \937_b1 , \930_b1 );
not ( \937_b1 , w_2752 );
not ( \937_b0 , w_2753 );
and ( w_2752 , w_2753 , \930_b0 );
or ( \938_b1 , \936_b1 , w_2754 );
or ( \938_b0 , \936_b0 , \937_b0 );
not ( \937_b0 , w_2755 );
and ( w_2755 , w_2754 , \937_b1 );
or ( \939_b1 , \935_b1 , w_2756 );
or ( \939_b0 , \935_b0 , \930_b0 );
not ( \930_b0 , w_2757 );
and ( w_2757 , w_2756 , \930_b1 );
or ( \940_b1 , \938_b1 , w_2759 );
not ( w_2759 , w_2760 );
and ( \940_b0 , \938_b0 , w_2761 );
and ( w_2760 ,  , w_2761 );
buf ( w_2759 , \939_b1 );
not ( w_2759 , w_2762 );
not (  , w_2763 );
and ( w_2762 , w_2763 , \939_b0 );
buf ( \941_b1 , \412_b1 );
not ( \941_b1 , w_2764 );
not ( \941_b0 , w_2765 );
and ( w_2764 , w_2765 , \412_b0 );
or ( \942_b1 , \560_b1 , w_2767 );
not ( w_2767 , w_2768 );
and ( \942_b0 , \560_b0 , w_2769 );
and ( w_2768 ,  , w_2769 );
buf ( w_2767 , \388_b1 );
not ( w_2767 , w_2770 );
not (  , w_2771 );
and ( w_2770 , w_2771 , \388_b0 );
buf ( \943_b1 , \942_b1 );
not ( \943_b1 , w_2772 );
not ( \943_b0 , w_2773 );
and ( w_2772 , w_2773 , \942_b0 );
buf ( \944_b1 , \907_b1 );
not ( \944_b1 , w_2774 );
not ( \944_b0 , w_2775 );
and ( w_2774 , w_2775 , \907_b0 );
or ( \945_b1 , \943_b1 , w_2776 );
or ( \945_b0 , \943_b0 , \944_b0 );
not ( \944_b0 , w_2777 );
and ( w_2777 , w_2776 , \944_b1 );
or ( \946_b1 , \358_b1 , \387_b1 );
not ( \387_b1 , w_2778 );
and ( \946_b0 , \358_b0 , w_2779 );
and ( w_2778 , w_2779 , \387_b0 );
or ( \947_b1 , \916_b1 , \946_b1 );
not ( \946_b1 , w_2780 );
and ( \947_b0 , \916_b0 , w_2781 );
and ( w_2780 , w_2781 , \946_b0 );
buf ( \948_b1 , \923_b1 );
not ( \948_b1 , w_2782 );
not ( \948_b0 , w_2783 );
and ( w_2782 , w_2783 , \923_b0 );
or ( \949_b1 , \947_b1 , w_2785 );
not ( w_2785 , w_2786 );
and ( \949_b0 , \947_b0 , w_2787 );
and ( w_2786 ,  , w_2787 );
buf ( w_2785 , \948_b1 );
not ( w_2785 , w_2788 );
not (  , w_2789 );
and ( w_2788 , w_2789 , \948_b0 );
or ( \950_b1 , \945_b1 , w_2791 );
not ( w_2791 , w_2792 );
and ( \950_b0 , \945_b0 , w_2793 );
and ( w_2792 ,  , w_2793 );
buf ( w_2791 , \949_b1 );
not ( w_2791 , w_2794 );
not (  , w_2795 );
and ( w_2794 , w_2795 , \949_b0 );
buf ( \951_b1 , \950_b1 );
not ( \951_b1 , w_2796 );
not ( \951_b0 , w_2797 );
and ( w_2796 , w_2797 , \950_b0 );
or ( \952_b1 , \941_b1 , w_2798 );
or ( \952_b0 , \941_b0 , \951_b0 );
not ( \951_b0 , w_2799 );
and ( w_2799 , w_2798 , \951_b1 );
buf ( \953_b1 , \925_b1 );
not ( \953_b1 , w_2800 );
not ( \953_b0 , w_2801 );
and ( w_2800 , w_2801 , \925_b0 );
or ( \954_b1 , \952_b1 , w_2803 );
not ( w_2803 , w_2804 );
and ( \954_b0 , \952_b0 , w_2805 );
and ( w_2804 ,  , w_2805 );
buf ( w_2803 , \953_b1 );
not ( w_2803 , w_2806 );
not (  , w_2807 );
and ( w_2806 , w_2807 , \953_b0 );
or ( \955_b1 , \405_b1 , w_2809 );
not ( w_2809 , w_2810 );
and ( \955_b0 , \405_b0 , w_2811 );
and ( w_2810 ,  , w_2811 );
buf ( w_2809 , \928_b1 );
not ( w_2809 , w_2812 );
not (  , w_2813 );
and ( w_2812 , w_2813 , \928_b0 );
buf ( \956_b1 , \955_b1 );
not ( \956_b1 , w_2814 );
not ( \956_b0 , w_2815 );
and ( w_2814 , w_2815 , \955_b0 );
or ( \957_b1 , \954_b1 , \956_b1 );
not ( \956_b1 , w_2816 );
and ( \957_b0 , \954_b0 , w_2817 );
and ( w_2816 , w_2817 , \956_b0 );
buf ( \958_b1 , \954_b1 );
not ( \958_b1 , w_2818 );
not ( \958_b0 , w_2819 );
and ( w_2818 , w_2819 , \954_b0 );
or ( \959_b1 , \958_b1 , \955_b1 );
not ( \955_b1 , w_2820 );
and ( \959_b0 , \958_b0 , w_2821 );
and ( w_2820 , w_2821 , \955_b0 );
or ( \960_b1 , \957_b1 , w_2823 );
not ( w_2823 , w_2824 );
and ( \960_b0 , \957_b0 , w_2825 );
and ( w_2824 ,  , w_2825 );
buf ( w_2823 , \959_b1 );
not ( w_2823 , w_2826 );
not (  , w_2827 );
and ( w_2826 , w_2827 , \959_b0 );
buf ( \961_b1 , \358_b1 );
buf ( \961_b0 , \358_b0 );
buf ( \962_b1 , \961_b1 );
not ( \962_b1 , w_2828 );
not ( \962_b0 , w_2829 );
and ( w_2828 , w_2829 , \961_b0 );
buf ( \963_b1 , \560_b1 );
not ( \963_b1 , w_2830 );
not ( \963_b0 , w_2831 );
and ( w_2830 , w_2831 , \560_b0 );
buf ( \964_b1 , \963_b1 );
not ( \964_b1 , w_2832 );
not ( \964_b0 , w_2833 );
and ( w_2832 , w_2833 , \963_b0 );
buf ( \965_b1 , \907_b1 );
not ( \965_b1 , w_2834 );
not ( \965_b0 , w_2835 );
and ( w_2834 , w_2835 , \907_b0 );
or ( \966_b1 , \964_b1 , w_2836 );
or ( \966_b0 , \964_b0 , \965_b0 );
not ( \965_b0 , w_2837 );
and ( w_2837 , w_2836 , \965_b1 );
buf ( \967_b1 , \916_b1 );
not ( \967_b1 , w_2838 );
not ( \967_b0 , w_2839 );
and ( w_2838 , w_2839 , \916_b0 );
or ( \968_b1 , \966_b1 , w_2841 );
not ( w_2841 , w_2842 );
and ( \968_b0 , \966_b0 , w_2843 );
and ( w_2842 ,  , w_2843 );
buf ( w_2841 , \967_b1 );
not ( w_2841 , w_2844 );
not (  , w_2845 );
and ( w_2844 , w_2845 , \967_b0 );
buf ( \969_b1 , \968_b1 );
not ( \969_b1 , w_2846 );
not ( \969_b0 , w_2847 );
and ( w_2846 , w_2847 , \968_b0 );
or ( \970_b1 , \962_b1 , w_2848 );
or ( \970_b0 , \962_b0 , \969_b0 );
not ( \969_b0 , w_2849 );
and ( w_2849 , w_2848 , \969_b1 );
buf ( \971_b1 , \919_b1 );
buf ( \971_b0 , \919_b0 );
or ( \972_b1 , \970_b1 , w_2851 );
not ( w_2851 , w_2852 );
and ( \972_b0 , \970_b0 , w_2853 );
and ( w_2852 ,  , w_2853 );
buf ( w_2851 , \971_b1 );
not ( w_2851 , w_2854 );
not (  , w_2855 );
and ( w_2854 , w_2855 , \971_b0 );
buf ( \973_b1 , \387_b1 );
not ( \973_b1 , w_2856 );
not ( \973_b0 , w_2857 );
and ( w_2856 , w_2857 , \387_b0 );
or ( \974_b1 , \973_b1 , w_2859 );
not ( w_2859 , w_2860 );
and ( \974_b0 , \973_b0 , w_2861 );
and ( w_2860 ,  , w_2861 );
buf ( w_2859 , \922_b1 );
not ( w_2859 , w_2862 );
not (  , w_2863 );
and ( w_2862 , w_2863 , \922_b0 );
or ( \975_b1 , \972_b1 , \974_b1 );
not ( \974_b1 , w_2864 );
and ( \975_b0 , \972_b0 , w_2865 );
and ( w_2864 , w_2865 , \974_b0 );
buf ( \976_b1 , \972_b1 );
not ( \976_b1 , w_2866 );
not ( \976_b0 , w_2867 );
and ( w_2866 , w_2867 , \972_b0 );
buf ( \977_b1 , \974_b1 );
not ( \977_b1 , w_2868 );
not ( \977_b0 , w_2869 );
and ( w_2868 , w_2869 , \974_b0 );
or ( \978_b1 , \976_b1 , \977_b1 );
not ( \977_b1 , w_2870 );
and ( \978_b0 , \976_b0 , w_2871 );
and ( w_2870 , w_2871 , \977_b0 );
or ( \979_b1 , \975_b1 , w_2873 );
not ( w_2873 , w_2874 );
and ( \979_b0 , \975_b0 , w_2875 );
and ( w_2874 ,  , w_2875 );
buf ( w_2873 , \978_b1 );
not ( w_2873 , w_2876 );
not (  , w_2877 );
and ( w_2876 , w_2877 , \978_b0 );
buf ( \980_b1 , \546_b1 );
buf ( \980_b0 , \546_b0 );
buf ( \981_b1 , \980_b1 );
not ( \981_b1 , w_2878 );
not ( \981_b0 , w_2879 );
and ( w_2878 , w_2879 , \980_b0 );
buf ( \982_b1 , \907_b1 );
not ( \982_b1 , w_2880 );
not ( \982_b0 , w_2881 );
and ( w_2880 , w_2881 , \907_b0 );
or ( \983_b1 , \981_b1 , w_2882 );
or ( \983_b0 , \981_b0 , \982_b0 );
not ( \982_b0 , w_2883 );
and ( w_2883 , w_2882 , \982_b1 );
buf ( \984_b1 , \911_b1 );
not ( \984_b1 , w_2884 );
not ( \984_b0 , w_2885 );
and ( w_2884 , w_2885 , \911_b0 );
or ( \985_b1 , \983_b1 , w_2887 );
not ( w_2887 , w_2888 );
and ( \985_b0 , \983_b0 , w_2889 );
and ( w_2888 ,  , w_2889 );
buf ( w_2887 , \984_b1 );
not ( w_2887 , w_2890 );
not (  , w_2891 );
and ( w_2890 , w_2891 , \984_b0 );
or ( \986_b1 , \559_b1 , w_2893 );
not ( w_2893 , w_2894 );
and ( \986_b0 , \559_b0 , w_2895 );
and ( w_2894 ,  , w_2895 );
buf ( w_2893 , \915_b1 );
not ( w_2893 , w_2896 );
not (  , w_2897 );
and ( w_2896 , w_2897 , \915_b0 );
buf ( \987_b1 , \986_b1 );
not ( \987_b1 , w_2898 );
not ( \987_b0 , w_2899 );
and ( w_2898 , w_2899 , \986_b0 );
or ( \988_b1 , \985_b1 , \987_b1 );
not ( \987_b1 , w_2900 );
and ( \988_b0 , \985_b0 , w_2901 );
and ( w_2900 , w_2901 , \987_b0 );
buf ( \989_b1 , \985_b1 );
not ( \989_b1 , w_2902 );
not ( \989_b0 , w_2903 );
and ( w_2902 , w_2903 , \985_b0 );
or ( \990_b1 , \989_b1 , \986_b1 );
not ( \986_b1 , w_2904 );
and ( \990_b0 , \989_b0 , w_2905 );
and ( w_2904 , w_2905 , \986_b0 );
or ( \991_b1 , \988_b1 , w_2907 );
not ( w_2907 , w_2908 );
and ( \991_b0 , \988_b0 , w_2909 );
and ( w_2908 ,  , w_2909 );
buf ( w_2907 , \990_b1 );
not ( w_2907 , w_2910 );
not (  , w_2911 );
and ( w_2910 , w_2911 , \990_b0 );
or ( \992_b1 , \857_b1 , w_2913 );
not ( w_2913 , w_2914 );
and ( \992_b0 , \857_b0 , w_2915 );
and ( w_2914 ,  , w_2915 );
buf ( w_2913 , \882_b1 );
not ( w_2913 , w_2916 );
not (  , w_2917 );
and ( w_2916 , w_2917 , \882_b0 );
buf ( \993_b1 , \992_b1 );
not ( \993_b1 , w_2918 );
not ( \993_b0 , w_2919 );
and ( w_2918 , w_2919 , \992_b0 );
buf ( \994_b1 , \879_b1 );
buf ( \994_b0 , \879_b0 );
or ( \995_b1 , \993_b1 , \994_b1 );
not ( \994_b1 , w_2920 );
and ( \995_b0 , \993_b0 , w_2921 );
and ( w_2920 , w_2921 , \994_b0 );
buf ( \996_b1 , \903_b1 );
buf ( \996_b0 , \903_b0 );
or ( \997_b1 , \995_b1 , w_2923 );
not ( w_2923 , w_2924 );
and ( \997_b0 , \995_b0 , w_2925 );
and ( w_2924 ,  , w_2925 );
buf ( w_2923 , \996_b1 );
not ( w_2923 , w_2926 );
not (  , w_2927 );
and ( w_2926 , w_2927 , \996_b0 );
buf ( \998_b1 , \905_b1 );
not ( \998_b1 , w_2928 );
not ( \998_b0 , w_2929 );
and ( w_2928 , w_2929 , \905_b0 );
or ( \999_b1 , \998_b1 , w_2931 );
not ( w_2931 , w_2932 );
and ( \999_b0 , \998_b0 , w_2933 );
and ( w_2932 ,  , w_2933 );
buf ( w_2931 , \902_b1 );
not ( w_2931 , w_2934 );
not (  , w_2935 );
and ( w_2934 , w_2935 , \902_b0 );
or ( \1000_b1 , \997_b1 , \999_b1 );
not ( \999_b1 , w_2936 );
and ( \1000_b0 , \997_b0 , w_2937 );
and ( w_2936 , w_2937 , \999_b0 );
buf ( \1001_b1 , \997_b1 );
not ( \1001_b1 , w_2938 );
not ( \1001_b0 , w_2939 );
and ( w_2938 , w_2939 , \997_b0 );
buf ( \1002_b1 , \999_b1 );
not ( \1002_b1 , w_2940 );
not ( \1002_b0 , w_2941 );
and ( w_2940 , w_2941 , \999_b0 );
or ( \1003_b1 , \1001_b1 , \1002_b1 );
not ( \1002_b1 , w_2942 );
and ( \1003_b0 , \1001_b0 , w_2943 );
and ( w_2942 , w_2943 , \1002_b0 );
or ( \1004_b1 , \1000_b1 , w_2945 );
not ( w_2945 , w_2946 );
and ( \1004_b0 , \1000_b0 , w_2947 );
and ( w_2946 ,  , w_2947 );
buf ( w_2945 , \1003_b1 );
not ( w_2945 , w_2948 );
not (  , w_2949 );
and ( w_2948 , w_2949 , \1003_b0 );
buf ( \1005_b1 , \996_b1 );
not ( \1005_b1 , w_2950 );
not ( \1005_b0 , w_2951 );
and ( w_2950 , w_2951 , \996_b0 );
or ( \1006_b1 , \1005_b1 , w_2953 );
not ( w_2953 , w_2954 );
and ( \1006_b0 , \1005_b0 , w_2955 );
and ( w_2954 ,  , w_2955 );
buf ( w_2953 , \994_b1 );
not ( w_2953 , w_2956 );
not (  , w_2957 );
and ( w_2956 , w_2957 , \994_b0 );
or ( \1007_b1 , \992_b1 , \1006_b1 );
not ( \1006_b1 , w_2958 );
and ( \1007_b0 , \992_b0 , w_2959 );
and ( w_2958 , w_2959 , \1006_b0 );
buf ( \1008_b1 , \992_b1 );
not ( \1008_b1 , w_2960 );
not ( \1008_b0 , w_2961 );
and ( w_2960 , w_2961 , \992_b0 );
buf ( \1009_b1 , \1006_b1 );
not ( \1009_b1 , w_2962 );
not ( \1009_b0 , w_2963 );
and ( w_2962 , w_2963 , \1006_b0 );
or ( \1010_b1 , \1008_b1 , \1009_b1 );
not ( \1009_b1 , w_2964 );
and ( \1010_b0 , \1008_b0 , w_2965 );
and ( w_2964 , w_2965 , \1009_b0 );
or ( \1011_b1 , \1007_b1 , w_2967 );
not ( w_2967 , w_2968 );
and ( \1011_b0 , \1007_b0 , w_2969 );
and ( w_2968 ,  , w_2969 );
buf ( w_2967 , \1010_b1 );
not ( w_2967 , w_2970 );
not (  , w_2971 );
and ( w_2970 , w_2971 , \1010_b0 );
or ( \1012_b1 , \824_b1 , w_2973 );
not ( w_2973 , w_2974 );
and ( \1012_b0 , \824_b0 , w_2975 );
and ( w_2974 ,  , w_2975 );
buf ( w_2973 , \855_b1 );
not ( w_2973 , w_2976 );
not (  , w_2977 );
and ( w_2976 , w_2977 , \855_b0 );
or ( \1013_b1 , \882_b1 , w_2979 );
not ( w_2979 , w_2980 );
and ( \1013_b0 , \882_b0 , w_2981 );
and ( w_2980 ,  , w_2981 );
buf ( w_2979 , \854_b1 );
not ( w_2979 , w_2982 );
not (  , w_2983 );
and ( w_2982 , w_2983 , \854_b0 );
buf ( \1014_b1 , \1013_b1 );
not ( \1014_b1 , w_2984 );
not ( \1014_b0 , w_2985 );
and ( w_2984 , w_2985 , \1013_b0 );
or ( \1015_b1 , \1012_b1 , \1014_b1 );
not ( \1014_b1 , w_2986 );
and ( \1015_b0 , \1012_b0 , w_2987 );
and ( w_2986 , w_2987 , \1014_b0 );
buf ( \1016_b1 , \1012_b1 );
not ( \1016_b1 , w_2988 );
not ( \1016_b0 , w_2989 );
and ( w_2988 , w_2989 , \1012_b0 );
or ( \1017_b1 , \1016_b1 , \1013_b1 );
not ( \1013_b1 , w_2990 );
and ( \1017_b0 , \1016_b0 , w_2991 );
and ( w_2990 , w_2991 , \1013_b0 );
or ( \1018_b1 , \1015_b1 , w_2993 );
not ( w_2993 , w_2994 );
and ( \1018_b0 , \1015_b0 , w_2995 );
and ( w_2994 ,  , w_2995 );
buf ( w_2993 , \1017_b1 );
not ( w_2993 , w_2996 );
not (  , w_2997 );
and ( w_2996 , w_2997 , \1017_b0 );
or ( \1019_b1 , \823_b1 , w_2999 );
not ( w_2999 , w_3000 );
and ( \1019_b0 , \823_b0 , w_3001 );
and ( w_3000 ,  , w_3001 );
buf ( w_2999 , \855_b1 );
not ( w_2999 , w_3002 );
not (  , w_3003 );
and ( w_3002 , w_3003 , \855_b0 );
buf ( \1020_b1 , \1019_b1 );
not ( \1020_b1 , w_3004 );
not ( \1020_b0 , w_3005 );
and ( w_3004 , w_3005 , \1019_b0 );
or ( \1021_b1 , \770_b1 , \1020_b1 );
not ( \1020_b1 , w_3006 );
and ( \1021_b0 , \770_b0 , w_3007 );
and ( w_3006 , w_3007 , \1020_b0 );
buf ( \1022_b1 , \770_b1 );
not ( \1022_b1 , w_3008 );
not ( \1022_b0 , w_3009 );
and ( w_3008 , w_3009 , \770_b0 );
or ( \1023_b1 , \1022_b1 , \1019_b1 );
not ( \1019_b1 , w_3010 );
and ( \1023_b0 , \1022_b0 , w_3011 );
and ( w_3010 , w_3011 , \1019_b0 );
or ( \1024_b1 , \1021_b1 , w_3013 );
not ( w_3013 , w_3014 );
and ( \1024_b0 , \1021_b0 , w_3015 );
and ( w_3014 ,  , w_3015 );
buf ( w_3013 , \1023_b1 );
not ( w_3013 , w_3016 );
not (  , w_3017 );
and ( w_3016 , w_3017 , \1023_b0 );
or ( \1025_b1 , \961_b1 , w_3019 );
not ( w_3019 , w_3020 );
and ( \1025_b0 , \961_b0 , w_3021 );
and ( w_3020 ,  , w_3021 );
buf ( w_3019 , \971_b1 );
not ( w_3019 , w_3022 );
not (  , w_3023 );
and ( w_3022 , w_3023 , \971_b0 );
or ( \1026_b1 , \984_b1 , w_3025 );
not ( w_3025 , w_3026 );
and ( \1026_b0 , \984_b0 , w_3027 );
and ( w_3026 ,  , w_3027 );
buf ( w_3025 , \980_b1 );
not ( w_3025 , w_3028 );
not (  , w_3029 );
and ( w_3028 , w_3029 , \980_b0 );
or ( \1027_b1 , \769_b1 , w_3031 );
not ( w_3031 , w_3032 );
and ( \1027_b0 , \769_b0 , w_3033 );
and ( w_3032 ,  , w_3033 );
buf ( w_3031 , \665_b1 );
not ( w_3031 , w_3034 );
not (  , w_3035 );
and ( w_3034 , w_3035 , \665_b0 );
buf ( \1028_b1 , \1027_b1 );
not ( \1028_b1 , w_3036 );
not ( \1028_b0 , w_3037 );
and ( w_3036 , w_3037 , \1027_b0 );
buf ( \1029_b1 , \764_b1 );
buf ( \1029_b0 , \764_b0 );
buf ( \1030_b1 , \1029_b1 );
not ( \1030_b1 , w_3038 );
not ( \1030_b0 , w_3039 );
and ( w_3038 , w_3039 , \1029_b0 );
or ( \1031_b1 , \1028_b1 , w_3040 );
or ( \1031_b0 , \1028_b0 , \1030_b0 );
not ( \1030_b0 , w_3041 );
and ( w_3041 , w_3040 , \1030_b1 );
or ( \1032_b1 , \1029_b1 , w_3042 );
or ( \1032_b0 , \1029_b0 , \1027_b0 );
not ( \1027_b0 , w_3043 );
and ( w_3043 , w_3042 , \1027_b1 );
or ( \1033_b1 , \1031_b1 , w_3045 );
not ( w_3045 , w_3046 );
and ( \1033_b0 , \1031_b0 , w_3047 );
and ( w_3046 ,  , w_3047 );
buf ( w_3045 , \1032_b1 );
not ( w_3045 , w_3048 );
not (  , w_3049 );
and ( w_3048 , w_3049 , \1032_b0 );
or ( \1034_b1 , \412_b1 , w_3051 );
not ( w_3051 , w_3052 );
and ( \1034_b0 , \412_b0 , w_3053 );
and ( w_3052 ,  , w_3053 );
buf ( w_3051 , \953_b1 );
not ( w_3051 , w_3054 );
not (  , w_3055 );
and ( w_3054 , w_3055 , \953_b0 );
buf ( \1035_b1 , \758_b1 );
buf ( \1035_b0 , \758_b0 );
buf ( \1036_b1 , \1035_b1 );
not ( \1036_b1 , w_3056 );
not ( \1036_b0 , w_3057 );
and ( w_3056 , w_3057 , \1035_b0 );
or ( \1037_b1 , \763_b1 , w_3059 );
not ( w_3059 , w_3060 );
and ( \1037_b0 , \763_b0 , w_3061 );
and ( w_3060 ,  , w_3061 );
buf ( w_3059 , \684_b1 );
not ( w_3059 , w_3062 );
not (  , w_3063 );
and ( w_3062 , w_3063 , \684_b0 );
buf ( \1038_b1 , \1037_b1 );
not ( \1038_b1 , w_3064 );
not ( \1038_b0 , w_3065 );
and ( w_3064 , w_3065 , \1037_b0 );
or ( \1039_b1 , \1036_b1 , w_3066 );
or ( \1039_b0 , \1036_b0 , \1038_b0 );
not ( \1038_b0 , w_3067 );
and ( w_3067 , w_3066 , \1038_b1 );
or ( \1040_b1 , \1035_b1 , w_3068 );
or ( \1040_b0 , \1035_b0 , \1037_b0 );
not ( \1037_b0 , w_3069 );
and ( w_3069 , w_3068 , \1037_b1 );
or ( \1041_b1 , \1039_b1 , w_3071 );
not ( w_3071 , w_3072 );
and ( \1041_b0 , \1039_b0 , w_3073 );
and ( w_3072 ,  , w_3073 );
buf ( w_3071 , \1040_b1 );
not ( w_3071 , w_3074 );
not (  , w_3075 );
and ( w_3074 , w_3075 , \1040_b0 );
or ( \1042_b1 , \757_b1 , \703_b1 );
not ( \703_b1 , w_3076 );
and ( \1042_b0 , \757_b0 , w_3077 );
and ( w_3076 , w_3077 , \703_b0 );
or ( \1043_b1 , \1042_b1 , \754_b1 );
not ( \754_b1 , w_3078 );
and ( \1043_b0 , \1042_b0 , w_3079 );
and ( w_3078 , w_3079 , \754_b0 );
buf ( \1044_b1 , \1042_b1 );
not ( \1044_b1 , w_3080 );
not ( \1044_b0 , w_3081 );
and ( w_3080 , w_3081 , \1042_b0 );
buf ( \1045_b1 , \754_b1 );
not ( \1045_b1 , w_3082 );
not ( \1045_b0 , w_3083 );
and ( w_3082 , w_3083 , \754_b0 );
or ( \1046_b1 , \1044_b1 , \1045_b1 );
not ( \1045_b1 , w_3084 );
and ( \1046_b0 , \1044_b0 , w_3085 );
and ( w_3084 , w_3085 , \1045_b0 );
or ( \1047_b1 , \1043_b1 , w_3087 );
not ( w_3087 , w_3088 );
and ( \1047_b0 , \1043_b0 , w_3089 );
and ( w_3088 ,  , w_3089 );
buf ( w_3087 , \1046_b1 );
not ( w_3087 , w_3090 );
not (  , w_3091 );
and ( w_3090 , w_3091 , \1046_b0 );
or ( \1048_b1 , \721_b1 , w_3093 );
not ( w_3093 , w_3094 );
and ( \1048_b0 , \721_b0 , w_3095 );
and ( w_3094 ,  , w_3095 );
buf ( w_3093 , \752_b1 );
not ( w_3093 , w_3096 );
not (  , w_3097 );
and ( w_3096 , w_3097 , \752_b0 );
buf ( \1049_b1 , \751_b1 );
not ( \1049_b1 , w_3098 );
not ( \1049_b0 , w_3099 );
and ( w_3098 , w_3099 , \751_b0 );
or ( \1050_b1 , \1048_b1 , \1049_b1 );
not ( \1049_b1 , w_3100 );
and ( \1050_b0 , \1048_b0 , w_3101 );
and ( w_3100 , w_3101 , \1049_b0 );
buf ( \1051_b1 , \1048_b1 );
not ( \1051_b1 , w_3102 );
not ( \1051_b0 , w_3103 );
and ( w_3102 , w_3103 , \1048_b0 );
or ( \1052_b1 , \1051_b1 , \751_b1 );
not ( \751_b1 , w_3104 );
and ( \1052_b0 , \1051_b0 , w_3105 );
and ( w_3104 , w_3105 , \751_b0 );
or ( \1053_b1 , \1050_b1 , w_3107 );
not ( w_3107 , w_3108 );
and ( \1053_b0 , \1050_b0 , w_3109 );
and ( w_3108 ,  , w_3109 );
buf ( w_3107 , \1052_b1 );
not ( w_3107 , w_3110 );
not (  , w_3111 );
and ( w_3110 , w_3111 , \1052_b0 );
or ( \1054_b1 , \750_b1 , w_3113 );
not ( w_3113 , w_3114 );
and ( \1054_b0 , \750_b0 , w_3115 );
and ( w_3114 ,  , w_3115 );
buf ( w_3113 , \736_b1 );
not ( w_3113 , w_3116 );
not (  , w_3117 );
and ( w_3116 , w_3117 , \736_b0 );
buf ( \1055_b1 , \1054_b1 );
not ( \1055_b1 , w_3118 );
not ( \1055_b0 , w_3119 );
and ( w_3118 , w_3119 , \1054_b0 );
buf ( \1056_b1 , \746_b1 );
not ( \1056_b1 , w_3120 );
not ( \1056_b0 , w_3121 );
and ( w_3120 , w_3121 , \746_b0 );
or ( \1057_b1 , \1055_b1 , w_3122 );
or ( \1057_b0 , \1055_b0 , \1056_b0 );
not ( \1056_b0 , w_3123 );
and ( w_3123 , w_3122 , \1056_b1 );
or ( \1058_b1 , \746_b1 , w_3124 );
or ( \1058_b0 , \746_b0 , \1054_b0 );
not ( \1054_b0 , w_3125 );
and ( w_3125 , w_3124 , \1054_b1 );
or ( \1059_b1 , \1057_b1 , w_3127 );
not ( w_3127 , w_3128 );
and ( \1059_b0 , \1057_b0 , w_3129 );
and ( w_3128 ,  , w_3129 );
buf ( w_3127 , \1058_b1 );
not ( w_3127 , w_3130 );
not (  , w_3131 );
and ( w_3130 , w_3131 , \1058_b0 );
or ( \1060_b1 , \739_b1 , \741_b1 );
xor ( \1060_b0 , \739_b0 , w_3132 );
not ( w_3132 , w_3133 );
and ( w_3133 , \741_b1 , \741_b0 );
or ( \1061_b1 , \1060_b1 , \743_b1 );
xor ( \1061_b0 , \1060_b0 , w_3134 );
not ( w_3134 , w_3135 );
and ( w_3135 , \743_b1 , \743_b0 );
or ( \1062_b1 , \111_b1 , \B[0]_b1 );
not ( \B[0]_b1 , w_3136 );
and ( \1062_b0 , \111_b0 , w_3137 );
and ( w_3136 , w_3137 , \B[0]_b0 );
or ( \1063_b1 , \118_b1 , \B[1]_b1 );
not ( \B[1]_b1 , w_3138 );
and ( \1063_b0 , \118_b0 , w_3139 );
and ( w_3138 , w_3139 , \B[1]_b0 );
or ( \1064_b1 , \1062_b1 , w_3141 );
not ( w_3141 , w_3142 );
and ( \1064_b0 , \1062_b0 , w_3143 );
and ( w_3142 ,  , w_3143 );
buf ( w_3141 , \1063_b1 );
not ( w_3141 , w_3144 );
not (  , w_3145 );
and ( w_3144 , w_3145 , \1063_b0 );
or ( \1065_b1 , \741_b1 , w_3147 );
not ( w_3147 , w_3148 );
and ( \1065_b0 , \741_b0 , w_3149 );
and ( w_3148 ,  , w_3149 );
buf ( w_3147 , \1064_b1 );
not ( w_3147 , w_3150 );
not (  , w_3151 );
and ( w_3150 , w_3151 , \1064_b0 );
buf ( \1066_b1 , \740_b1 );
not ( \1066_b1 , w_3152 );
not ( \1066_b0 , w_3153 );
and ( w_3152 , w_3153 , \740_b0 );
or ( \1067_b1 , \950_b1 , w_3154 );
xor ( \1067_b0 , \950_b0 , w_3156 );
not ( w_3156 , w_3157 );
and ( w_3157 , w_3154 , w_3155 );
buf ( w_3154 , \1034_b1 );
not ( w_3154 , w_3158 );
not ( w_3155 , w_3159 );
and ( w_3158 , w_3159 , \1034_b0 );
or ( \1068_b1 , \968_b1 , w_3160 );
xor ( \1068_b0 , \968_b0 , w_3162 );
not ( w_3162 , w_3163 );
and ( w_3163 , w_3160 , w_3161 );
buf ( w_3160 , \1025_b1 );
not ( w_3160 , w_3164 );
not ( w_3161 , w_3165 );
and ( w_3164 , w_3165 , \1025_b0 );
or ( \1069_b1 , \1026_b1 , w_3166 );
xor ( \1069_b0 , \1026_b0 , w_3168 );
not ( w_3168 , w_3169 );
and ( w_3169 , w_3166 , w_3167 );
buf ( w_3166 , \907_b1 );
not ( w_3166 , w_3170 );
not ( w_3167 , w_3171 );
and ( w_3170 , w_3171 , \907_b0 );
or ( \81_b1 , \80_b1 , w_3176 );
or ( \81_b0 , \80_b0 , w_3173 );
not ( w_3173 , w_3177 );
and ( w_3177 , w_3176 , w_3172 );
or ( w_3172 , \I[0]_b1 , w_3178 );
or ( w_3173 , \I[0]_b0 , w_3175 );
not ( w_3175 , w_3179 );
and ( w_3179 , w_3178 , w_3174 );
buf ( w_3174 , \I[1]_b1 );
not ( w_3174 , w_3180 );
not ( w_3175 , w_3181 );
and ( w_3180 , w_3181 , \I[1]_b0 );
or ( \106_b1 , \105_b1 , w_3186 );
or ( \106_b0 , \105_b0 , w_3183 );
not ( w_3183 , w_3187 );
and ( w_3187 , w_3186 , w_3182 );
or ( w_3182 , \I[0]_b1 , w_3188 );
or ( w_3183 , \I[0]_b0 , w_3185 );
not ( w_3185 , w_3189 );
and ( w_3189 , w_3188 , w_3184 );
buf ( w_3184 , \I[1]_b1 );
not ( w_3184 , w_3190 );
not ( w_3185 , w_3191 );
and ( w_3190 , w_3191 , \I[1]_b0 );
or ( \138_b1 , \137_b1 , w_3196 );
or ( \138_b0 , \137_b0 , w_3193 );
not ( w_3193 , w_3197 );
and ( w_3197 , w_3196 , w_3192 );
or ( w_3192 , \I[0]_b1 , w_3198 );
or ( w_3193 , \I[0]_b0 , w_3195 );
not ( w_3195 , w_3199 );
and ( w_3199 , w_3198 , w_3194 );
buf ( w_3194 , \I[1]_b1 );
not ( w_3194 , w_3200 );
not ( w_3195 , w_3201 );
and ( w_3200 , w_3201 , \I[1]_b0 );
or ( \929_b1 , \917_b1 , w_3202 );
not ( w_3202 , w_3204 );
and ( \929_b0 , \917_b0 , w_3205 );
and ( w_3204 , w_3205 , w_3203 );
or ( w_3202 , \927_b1 , \928_b1 );
not ( \928_b1 , w_3206 );
and ( w_3203 , \927_b0 , w_3207 );
and ( w_3206 , w_3207 , \928_b0 );
endmodule

